/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
l4gSYexUXlM7ifAaBP6t2MLRFhQaRe7Sma+zo2L28DiA8DDFN158h0/DaBr1OsRaQKqTpiBWurc1
Kc+8TD5uaOBbdGAOqQnBtAA+GhRIwIir9IbLuxBMnT/JmOaK4MUYPqvoRzrgYyXFE5yrJmMkU220
b8Arh6+dyt3Bh0bC5r9kA89v3D+ja9uQnY/8oodAq0Q20j5GmOBNL7A1mEvLof/A0UYhDRCv3pRO
FKF8KrYOR3RN8PBeGCM1EFnr+wW3J99nOfKe+v5+if1arByO/0BxWK1JYTBdcxntFYOrk/8juzWe
cyuQA25yLLNZSsEfw7pTdA4YqggvIwnYX+4CfA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="nooMg7GjkDsMTPG3DLODBuXednbZgjpzUjgowzton6E="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52400)
`pragma protect data_block
OIw4y6hn7TeoR9JbrM9EZGVOSQ8RnwJcq3UTN0ZQEspziLZmwWO83l9mud2+eh6A3W5BDM+VE/sq
5XVTEeQXt3wqLYeYfWktw5CWxajAk3scDhRmpzDrc69/YUansoEmGA7OKydBKp7ojGgYCMpBqwQh
ohTEnLUYDBO9sMHkW0vFUkvnnqtye/AUotH+GvUhgmbTtskc0fumOZq1CpebvvjdBXXKeJVSYHuP
VLgEJ91XDl252Gl+tsQQ9NBhcRtfabzKS+yadazwXTW4jowBYtywKR16p1PU9xnGcFaU/yNXokH1
ilgVaOPxR0jcW1O8YZJ8P7eEfSUtXQ+WCzkJNGi6i5tqbb9VdzFm1FckcRfDuWglQDZfVGeHsBa9
Kw/RwZFdK4djZBVRmPiYqtjD6qsdoE1OB8SP+SzqS9apXMrQ1S5Zh8Pfg4bYewWvT4nfT/e7o7Im
iq+yoavfjn2CLfzAGk8nuD0ujsO5BjjyMSalxuLpiJ0ZLdMPKIk1VjI7bWEc01GPxvk4tdhBX89z
DWf1qkB6mixpuMinljxaiR81jR3gDILrSLchgLXc5VUGtgiNU3BXT8KI6LslMvgADW67ZtGvNfeq
3LMeFQ5CP7xMGH5BiD2NAvBOlnmnkkcY48+EPBKpNRWqVh86dM7S1nP/1Zmj98cbcSFOzIWE4DHB
KHNTX+4/xdtvcUPEBYhAPZP0wiNp1rwAnXccnDUJdRQutox4Sz/rPi4LjpFZY+Bw1h+djt+RX9js
DJX6EerAxnKY7sU66r3AXoCEB7JlbtI/X3wQU+1nezKxcxUJzyHHL2+sYU+/IaNodKoylt1yTc7f
xO64cAgz7EC3YM9MyXK3dJk4Zmjh9nXvSIV+KtMCFw27HODI0u71J5RtmesXL4wssZ1JPylD1tOl
qmyQ438dF2mkuwOpZHYVD6zJhz9r4b5BIOKg7UG68uGKiL5UCOIbMa+/NzGX5CIbqOjqCdnB1dno
+hqqpONN8UgpmDBv5y28c5BLH9/DNzrGi+yPdVn2QNz1ds28WTJWpkaEcls3nU7zW1bWzoqr3yHH
HlK+H6BFDaARkHi/0UhgmUwTI4QurZS3TQ/Bi7qao1Sabn04w2isKO3K5N0inQCwLdU/3mtJN5pz
4+y6EPAlEwqSBsABOmA12Jhvk8jSkJYmAIIoBltfgp8mH/bxeGX1HA4HnDKpJwpNN/pIYuo8MVkU
RFr4KPImv+skcB016YTPB3ck8cqszIHdhCfbLi/Wmo4L7iyl8DcbeBLPCKLVQfVpn5W8LpmlfPFJ
sXDRek0+AsMz4TUPQgSkJx86TGdC9iRal/X/YioCAFuA711z1ptxxbrrnOWG/l+bRnebrm0aB3a9
VjqnWSVl/DXM0mdqjy+d2S2XZPeeDNjDTfOf/dSqsgcvlkjgotBCVQF7PGQGe0+dLfBuTp9yFyOZ
tM7VmqJ0GvkXtAlLf6eYgqGdJxCPZ0fX+TLHyv0wJxuhf19qoRJCXihhCNwVREg02Pn8d012xfLd
RG1C+y98gSDFAR4kdeeVpwYdowYIt1AYpMAlwpxE04rSzrA9x1j2D/cWZ9ig6Ic0FWyaBVYv2SY+
mh/rt1xL1YBPfC6i+VfB+Nj1Bk3yVkJk6K48nM2UkouTxNMj7vfEXgIY6+ygIpNkVpIkOK6K/75u
vUQG44O/mSU3zgtz6U3uR8bZ1q9MV7CIY9jLl+QrJz1PaZ68Jh67qBVprgWOG0cYIxDmt1/WjAMS
Ls/vFdc7RplUHA2fB0UUYmZqj1ZJpqj5uRwps893E/1sZQ772unLYAMuHYBeJMbkJu0nIqt32zhQ
Ht0S0d51GpqRJ3UzM6QIWekAg8lx/wzRCgUpUslAH10txoua6GOxYSgzlQvpxJH+zzyCojKbc4rm
RVPoB5JlUp4P8Iz9jHQfBROUCzPjqwrB/gxMLuPcRMqo2e+/pTOyISted94NsKC4rWfGjnuthhO2
5LkUm7UnbXSUeh0845PyBqIV8JkHx2SxbrcK8F70HPY242BiZVu88MuvIkBviGc5Q7+YnsKlMDoZ
y8DQFkejLb5ZVx5KBfWbyRw5QP8S2YU4s3xAfCLK2ATadrpkdvUdG9ocePWGa+flYHxFphrx5FE4
lcGjD4JXEkCHGgg0AfnS1w4hdFY4mAV9JnlX4rKdUbPslYKD8XdWFmE31jl31Axm2RaPvGZ7vp6c
W67OoqmXgulHRjcLRdpN9D/zUljgVXuLMfiM2q64KSVt4eqtkMT9zPeLEkT8nPGtLMFUBkJ2M5lm
iXSUrPg5fmG+OD7bmD+7Thn+Bx4dVNlGwNGaOdmxLH9qGNmxGccDSJJOgikMbCpTAJHYroW0FmFU
serbuKpreQM3Z6EccJ8KOLi3YNvErUtEdOaHt58rsLfqfjinbvjkQcwRGjmZlaZylSlkuiT2yn42
x4S8YO2k/dh41RwITcQZ+7tj3dQdWd4BxQ7LvAvpyOmKiWEJ9/5oYgZ/PDxaI15GEVYDLKwa3+KR
VFFfYWho3nvjVNCDSbdrqblkYUsNLjeQLcF45wU7H7diTxAZOta2AfUY7Mf9n8zwK39yfk6j2jSH
hFtSDRLXCpTtsfuP51t1NrrX7UNq9efCEUvJLj7h62jSEMY9LkAe69yt4vTFqZyKI0sDe88H3PzH
wVWifUmbwvRmFx1dEzBFvMYVsT/MhsMWa7dWfqJRKDohGhR+e/6lPNY6aWgipOLIikj14Kcf2HPP
/NRhYGWRgcMa9UvjFr7bp2mc3d2vSueQhmE5L/u+poAqal7l98vUA+VPsVse8wHfj6CX4tcOi0oV
KW5majNDQZFRvKP724R+m/Myx8+hpS+lS5hRgvDk0M9FQIf7M44W7H85BlJQGtbrY3OHPdqcI0D6
Wi7wWSPzStrKuJifXRl7zCCbh9y+MjyN1/ROhFO/SLgKLP6vb5CEEW/7s1x4+444P4Fk/9GhRDEJ
Q/LY94MwLo7KS1W98gYTHSwaT7SUu8v9Tu0z3b4V43dpKgbzlo0h0poNVLliY3GYdcyjrEAmPDSo
kypE428l5lR6zVd1hrjhoX7vHUjAyOckciZHJd2SrZUvoAFswX9yDmot70wvlInc72edR/ADVDbT
wxWdYvE3/p1HXl0S9pDPkGhl8SjJWfOtfhqEcm/9RLfmVHvuIzJmrZmJBG5YqUc9frkkO435mXx2
6RRhRD+CTnZlz3u84f5JVcVCe7zeju7nZwEEHdvY0ObuwmEVW/UNROKrbZXQPTAmOFDvdPZCLJHh
N3CaWs1Mj6rhZsPkPmaubhDMUsXyvX06crrNn30o9jjKUpgaDXe6GiRzQ9cTjak/Px0YeAN5Zq+u
ZXFMWJvuj21Yza0KaHQ9yTqMgUvHJMdVPUCt2ixpcS+GFFCVvoyAKRyEOuLkR/TjX0D3pke+/FO7
jTjs7DIoJFeG4sqsZznio+2AjhOrm/KKW10f+sDMHEoTO2UP0gA4Ch2Sdx7kTqoIDDlscPsGy/ZX
bszjxaNBqZIfDw+19bfJM95jfeVaULEbjTW3XBLb5zBGEQcWcPOM9uskrR+glgipBXBtyY7L3C6R
mxHErDTw9ljxPAcFV51dcoCG9nv1ur5goXyuOe8XyeocdlpsitqQeZjAZ2snL2woYMBINE9ezoWw
uHwT45KnaDn4cLeuJ/d0aZuhzC7nk0TMRraV+nTjbSAyjVUvwjPS6yDi+N7tM83ps0AFrR74oHW5
dTGADbf3hMgYnXPYoHWymbS1Tvf72TKQrEYspgEh6q6XjPyqF+f+5wj5KrkXVHmq1L2JZc86+CIa
YanGlfZpwjqqQxSFWEzrPYHhF0J7R5yyjOMmi0/Q0a/zQp5NqViDNjiHKsBUPhVsGFBfc8xUSBJa
nO1yr0t3fXAM2fhFH6sawDi21yYzcRnFX6Zil5FZ8tQysA1lIkV//H2nJISrfLOPC+R7tzEAOHPo
cpKQNP4ZTSUBQyyZ6G+RxkOXxGPiBrPaC2PWslcW+WKELuXVBUKO65mT2k4Hy8ySAOo4IU7Nx1Vg
lyaYQ2UL5ofil//FiRn9Y7IsKXOPYYXDKFFiBUZ56PPiWu/WHHPspxZGHxCwrKMZaDlzMH8h3CPZ
/7bJpURIQIQkuBq/JnhxaXalkI04aCEM4dir824A6Y4H9eYGlX0G5HUy71+3osklClrzXaNLUtW+
QYKzIivE1kFsI2fpAxHBN3ur9O1QrEM6H5nFaTvB/VBEuPXPRSniREbY3wQ9nh1NRnc5Ym3qL00U
Cogy6VBSXAvpY+N7G/jnwiNmouKHzQa7Ldx4V63MPv2LDJnFZjc1tUJDCKzhMrsdKovNPxsNycf6
1ZblINhiAdyrscWlbn+hXdJjRmrptbiqr0Vtc1uOzFkW7k8v/Q/hCWNLSsECXZwYtDuZ1FZbH+ig
LHM/8SdEoB/r/3uXV34xtrUVkrcuMo5tT6VTdRwF/zkZGZFsn5GOj9rBqEB4y3AgbR3NtXIcIGw2
SD2Ub3Rc+HyFgCbYSfM6Pch1netyJ8xA5L10nJ8NHvmD875bu/YvhDnwFs8z36deJfe+guCuhMFI
Ug4tCZejW38JuA98tjOA/ZrgPZ0U1XtpUI9TxKlhs1lRL33m70jvKZQGYY0LypjfqqfVeNjbbAWn
9xFDksgWy3fWxoDpYuQ66u1WbnT9ouHkDWggUIUbx3Vv7ibutXpRB/16PSe+eKKQjd0vwXVPg+En
xdW5m/gYQqE2Wi9qNvl/YbeCWGbla/QYxeQOOnvsDgr0ZCsLlWue/v0e6nyDWcmRon9rbRDR6R72
8QVCQld9ZY18dXyZFfVDqHYkNj0XGBsBS3YofQEic5JI0Ry1bH793+pnjxNexT4RaFJcLhHiV/OG
CqxDDoYqwlHToOFwPpnxuYppO5pziT3vsqgnfhD6URB/KzgMWDnnGtue8UfWVLNJcTx5Om3zivV6
/VL4f2GF3k/PzPh4jV4ySF4VnGoe0UPby6NlXhtyb4hbe+54FSKNoIMGI3URj016oRFgW5RUXOWG
e1yLh5VO/l1P1SmHhjTPvOJ8P5/7r8RvzljMw2cK61mrYR0rPRNJJ3xUbbpsINBDtryGOoCkWvnt
bRWjJ6ZIPrUX/I9YRTfpO9j1jUslkUxCMig2iBXJCsBwIYUL56/k6e3QFmC4OVCiyFMB8tpUzChk
VEXkgto32li6XMy2i+EI7dFQmjAQLGqUpPAPAslpXq0nfszLdPlNIAY+L0BehADCpkS/7M43CQZK
yK7lViIe9lVI38YaQO4KKzC1X+CPsOnke9HhGekLFgsvXUC2TVFqMCXFiZfKtjI4+bTadUQnD6Zs
EDRpU7GM7LHUC+s1LjjGsT5yX4GdYxj5wK6Jp+ctxgyY0GjKAa6+b5UyNLgDLXvWvt+fSMmfU0Bg
odyktV8mbRhcrL4p0iz09YZN3bxB++dLYPh60uMX4Rl5XpK/rMHSu6nCyGJxxa4+eJW65SlFtkNj
WOCTJonIqFd+2pnwT7Qp4qshOLd44ZyeKt25q3wJCgjWwJm8fkZ+yEOsqmhXt5NcXCAMDEfySp+p
L69NheSoqk08g2gTDLRHFifOsL68oySXLK5Z5LpVSFDhWHem5XMkJGuKj31D1AWLJvgnBkzHnxWl
obDW70gIOh1ol0VpSN7vvBEHpeMcDqmKffTcleLfbNxTh4fdbqe4Vj3je8RevwvoNKzO2nFfqYcF
mkrXVRzcj7xluKuYFa61pSYynTqoiokNk12MdTlo6YGCV2Gq5BWhw4YBHO2TFQ0LJuJQn9jqCfui
jDnx0U9vqGgvjozJSRlGCC2NU6J71r84xkB4QRU8EcmOt/qhGCyEYEmUdCnMwKLBpNtr/tcSZuQz
KiT8Xl6hxDG6WdwryZtxzIo8f9i4Z6RZPUeJzl3Q5xmTvm1GuoWs7F+Uy8iGJcdwpr+2rRRHboS+
h5zYgGCMJXhBzBLiQ2rQmNFB8AVnVDXxstGMgM+Javs+hccm7i+JrpCaPGUVFAM3t56yP/o2K2EC
SGXAD/3vPZd4BWnYhLpfw6NtPnTiF0QyIrSALMmD13XLy80GAggvZaptxsDiWopXfFL/6yg5foVl
XeO2c+3H1S1i+pom5tOj3C9AspYLwibHx55Q90WKqlM8Fs9FF70U/8CTLDaQCPxaCKbw+OgQBhAT
Z7bZoDXTBR+DHpozpwsdwEOyNW284Chgp+DiAR/eW2VUVICD/N5U6WwXgNzKBFEveBMipQfWq8+P
87Q8WQplZVzEzIIEJYUu3hPJe94dseTYZiPnSUSEiWet0qC6Ep9DyBh7IDEquZdCBhfEW5i9eKag
BXFlxfz/+ezwqhiqeesjp/UV01jaSzNq82BVF/OrAMgTmi8CK0Pw47y7raOw+CSeMuaV9LLJLk6Z
S1Rmucsq0VmgIzAnDo7h78U1au7eBs704OCRksUSzMobjaNh7wM/XZxdARRe8wsiM1qRo7+l0Uv/
1x9F2R75RtRFDxXNxhPJEfop1oBOf1hhy2ALvSQGjhQIfvs2YN/3OoXYjrZ5Qeuutk9CBIkgXxF3
kv4crn8efUGKRYTZRFn5h9lRTesWQtH1ehAsK9U1Dl2zMvp8OcFerbH/xEb68RxAIWQ/j9j1d6TW
J+ZV3VFayIvnzHg/DkbCgCRTq9S6pgRCyubzz2pQh526RCyhnPSXDuTkWO4xhnyenu+O8wNm1Bov
KcX6PrIIFSt0rk8IYaw5bShFHoH0LgahzAcqerSzQ8AGqIqFcw+GXY0QdLrdhdmxIUm4BDZ6wBAD
Hjq8XqvQGWZYgEUNG9/lTDTfqq0GJpfq8Ao6w7LzBQudH0SN82PTqv6BGMDVsdVuaucXoCS/c22i
YmsKT+NjJRfZu4kVx+ORfoh+a07qemSMwnwFYqtw+sCbkCaPsTeLc1ERiHotBpdBEXi0KgqP6DiF
qgb2JN7ibNJ1XFuJMXVjOdC64chN/Rpbo31VYrQaJ/8QSKj7Ddk9DfM/D5P11yNtMlMsL01xy+ua
zKhautRFYsFW3KBisL37RTzd4az3d6nACVol1GYZPWafQgjSRD8sY1V/9p2wbV3PTq+UkUZv3O3I
VJQ9CfxXqH94xFtl160CNsTkZ54Blynow8KMfVMl2hsJcR3AWhssK1QpssU76R10cRCcZfmySFWI
v9b/Sw2Q910huhyWGBk/0S7eWzeVKte4qSNcbimMnqZXWKepGdBfiTNPItAqij/Pb/l4FuPShAaG
4Ac4qZ+uDpdBG49idWJz2VV9gFnZ2Wm7uOMbBGdfYYypYdu2tTUOtBFl5VrzIXzrhdY3CCB3N57Y
nBYpCIo0OlxOU7Lguu+O/zjYachvkD6aiSYeP/v27Hzp0Bb7XmsH4KwKZITyFimpZI55zCnMr3LX
/1dGJxh7io/NwzPIIf8OhZGPHH6MpvZ9SJrvHyAV9eeK5vL/FJn+Ww1zJORFCWPo1CKEA6ZD7Kxd
YsNGecy9Ns4g7DSQmjFSlxbnB2LpEeOpQshHKiikOllCVP6dASzNzyzRKTxkh1ZaC0N1ZESh1W5y
POFXQbt+gKjJ7LIrhdLv2eShfp96k2CH4mmD4yDdkBa0izCcvdRcFhruZj2En5PZ4mwnuIoe7c35
AZKfjaw6dVPaYiQqTkdKyA0+XR2biJh4ICCBYxc4UFYximWOxGMKGLHvHtak0l8ZzguV9hkndc48
R0/l2Dn2QgGew6cUm6USN1GzjrDyUkUrHlOY0SAuBpcCFSSBA1VNu+7+d9Fc/1aTYGMqSIwvavp3
HniEKMyoz1tt2XiT+C7nEN2uCymWf/jDBMz+zQ3diArdabHvBVCWLzlPr+FOK8YTl0TT399TWWOt
hXp+tBasHyAWibEMai7bvkw+2Yb50d+ImeARMjLrCmdSbUOeraOrM+LVzjaRsYaG8D6MsfEDCuGA
5gQdWKCjT+m3xj5nsSOPXyolEEDRJcWTsM/asPiXO06fxj9hDa7zmlnk0WBwK+U7p8XgxfA01bRt
E6bE6qXRFPsLcBPzyauuEHZvXZk7GlNQHEPr12Wxdq3fmLXPeV+rs8qznDioPsH1bRmlWdy5Uhw3
GYUtFEz0o7Bfuv+VF+mjK6CVhm19+S0WlsaYvDpVDeGRT567dsGrqpWqkEwHfV3YFoVddyGtC/Do
nevm85AdBRFOx3HzoExz0pqP0Fz9kGq24vWh86DjfuBUdnawGNd5759QBNmX9dwkg1hAySHCnT/O
/jmi6+vjGiX8kbr5fRr8u/k/VmwcE4JXXv+ppokUaf3ZTUt8UmTMu/dp1Pmis4kXvNIw7EDFEBzZ
YrZKGQ2Jo/8ye0jd5ipyx7Bm3IWMd+LwkBuOVfJqhc3Wb0Fuh+uiXkovQuh7i73CzfFwOTg208BD
f8hObrw+Wd03sqpjFtlVkqBGAc+ngFN5BN4RqhYd+JQj/KuEVNwo/r2yzF9hSWZSKMspxJw+mJMi
Tt+SHz89s9YCud/lKwBuokq575FFtlE3Kzv7EpaE1EuvC2lBveYVnmhVyGbtfgkxRUr41wW4JinH
+ul4/HpsuVJyYYSR/lF4myh6YNu0cl7QuNVaKriUPxcCNUT9+vG73vMYwi3MKew91Dx/O+xyDbS0
kRciWVcCHmTJB4roouAEIbeDLOzl/ik1W3FCRD+7M9QwKWwP8Dhge5HxzJinb2w133Xr5JYukF7B
EMwVrlyzSH/CB6oGh+fR8qu8RnzK69x67QfSfV6xlq/N1EHO9foDjlTBFW8ukloopjrqr+6E3Sv1
cVZh2wAHAWe85KEV6bP9kthm2Ea+bGNqr3o/xsychsJ0MU9htdSwswucKXx4pw42JXu7OaCI1/pw
W0VSmulqPmhpi/YzzZa0jTUHlI77jA5S6lN+2g90tKaj47GzR/7fW/4DBY7CHcPlOTAs3GhfeeHU
y4Ax+2timiUY/UspsPU70ORoyBgi/fBFd3oJp6rCdzpOP+aTJPp4Ybqkd9NAYQl4laFP8u/BpGik
zLawVWVXIgyNuv736tQe+TjMGukC3v9T6zr26HBVJ6i5C+0e70fufcHyXdVGOFCnk+oF6AdHPx9K
HYR6a3B19zCxUjyTwS1fQCA9QUgE2hizmtsNygwPXJx15DKWPMi4gZg2KNqmC+eysbX71eiNzBMz
P/dQrJvl1kY85mpmOqLH6gF+DUzXxZkUxmKzInLknJDAlV0upp3iFTGNp5C0T0eH4P9hGOG719dG
KYT57j1pttrOFa/cgOWXt6jDQDVaUSKuANDZn7Eb1IkCvfOp+/I2mIVRCz0jpBsbVwiD+VIOLruw
IgETixyHoKPlDzpOkeV2KeXoKqegQCSoCuE+Qtj518Kmgv45BSiJDhqGm3zAIIxjw2E1sIjtDr0h
X8+M9oYT818KPofXGKDn5rOVeGZUb64krxVCVAAyO5SmJyaZZ5PEgdWhh0E0F5IYk5y23JN7Tt9T
R3cq9JwXFa6mOHFzvfRgs37c1MdL9EIwC42z8jS29fdRqRzSIXNUgpEo5WDq2W5HTq5sn2cL0/Fu
TAyy4R94PYZTeAdrXKOThDRKVTUTbk+eSp9bBRcop8xYVNT+tLRtjjhHB+5dNneJ8t4M6/41/gPa
xpmNXWeaeIClFmOsaUKIOs/VzLRiJwQyX1OLBp8gd+rNcHxA5C+mktISiPq2xDKYDOkc5iFOTCgq
AZgfRDS088qzYpT79pxfDH/IKzHELXwE6KFluhqnv4m5hEdNhSavkc5ngSVD6L8rkGD4dAAefAAh
sgfOW4Jo0GBseqMyZBkaTjFygtrU4RMv3c88szzmwsqhuD8k45e7Lg9dzkt2Be2ZRVPe30M8z+1N
36mAdm27ldN5nBQmu655GSKo7qy1ofkEnY86hFqVIBfX+snSS+ci9r0XW/46a5lra1ZOcD6mzr2k
QMtsEdUWepfyr4smWyHkn1kiDOjitYY3fCsyKvr/C7uUe+7mP9fPN53q1FhV7FeASfIajAZq3ZbF
8uOkWN7ntWNuZWGOScZK1yxU/XQerh6ggll96okLapR9u5nASar/29GuE3QKZqE9FCghxaNzd2aw
1Em2RJGf0duT6kzazI6BQfsdumoZM4muETXQK/T0VTYnVeZMaML4jnQnRlNrfTQ8dY4ZJJVVCiIk
427agBRcfcqMG7TNtAfmmOIj1P4wifr5Y9yX4UetiDDunhl03H/Ku3SFB847lH9U5d3/bMybXLLd
y8AEzXSNbHeuMCm25Z4KvxBnaDUrcWL9sJWZIhVPP6lU5AC+tI3366GiIzGEJl2RotUTtkX204EN
L34W/u0BeRvT7n61yGI4E0/jDvkpagsta/EJMjcnrO/4kWVOlaEfKe+BVtEUtC5gtDWVdEuZ7rZd
3MMwoZx5iaQZ7vXJBwdfc8zydS211ZSe2XSxPLXevxiYCg6eYcEvI45hDPf9rBjJ2BPTYTeElPg6
IFl2OjBztR1anEzBEDjtKSqFHriezm6no7cGM75UH2d4MtlHkIwzAwILeg96rPpOI6HwBuMYgr94
QatsvBpehUeCigxYP7lTKTDl4nuA3m14Leu1NDthAJlTOY5/HaJ9GBMdAflDVkMzWmfon9csucXA
ooGS9EB8wzO5UbT265mV6dPX0H9mC24i4UMdF29YUYLRYzlqXSzMH/Tabp4HvvqIZAcV7Rm8hLt+
bEHQeQWfo/LUnYJWV1UbiuGqEHPfqlfYfVEML2dvK9VPq5Yi1CuyzrGHJsx18d1GNQf1snmvTMj1
vgNrmNyjDtmjtPSNvU78tbxQ7G1qcYKu9dNZ06zX1omqNMdqCmydMcVZEPyz39d4Vpcl6OolJa5D
8mld2sMW7Orx4VoXWKRpb2+aC27zmloH615qWCVdnYE1nFJij57HMq5yPgpN8st5OcPYwCmdsee5
tookJ+N/l2mh9z04QQN75NgWJGPlioT2m0Dues/tyHkLM9aJgLuTc7wX+1mKYHYwLGrUBQp9Na9e
4pjVpPsjjz4j86GPbPA+DdKA8kA9x9vxFaCYv0Ppx/9R0RUerWolupkhIc+zaqxQ1yGu6f4Z1N6U
j0lRdVQ8ygpeCKgZVUJFB39uWZ9lVVsOMgd+iu0YghGd9KSVhrB+WpoInJYNfcaaspiQov2uk09/
ikTBiHO+Vw0k6vfPzWnJM4nhWtVcq1ojM2ua8dTCcdg5fUGWcaiULsANTJFSw5WyodJezzvZ77vm
ZumUh6jDAanmo7hSw22k7YKdLv2b4jMb2ofS72txxrw9nA+m30yR/KX5rAtHFzlhALWOq05/8GRS
kt04IX+XClzSDrm03WwISsmKuYJn/idVymnpCyHvLwvZkAbUoTyGbjja8PUS3Ooa/DKkfwsElUI8
YpsefJS3dCvmlr/2FOGSun334YtCbLH21joW6vrFLK8rfcstorzJ+13Sn94jcCFSlqogk4VJwEJc
NpbmRbahanxg218XEe/v0qHtBbB+IyBeR8jbGUpofboWpMgFz+Hn66JJBLw3SCQblvF8QlUONcYX
1M23LAwVhj2pCHsaRca68ZYMdfvhuAZ055PMd0uPGyWqQGtmNiniqjSkLrjuTGND+EWZ3IcjeQFk
91bNR9lMVVd4Q0ml/9ZztP25iweF6ES1uQQvctHnTJ1I7cClO9VO/xKlwAqEpRHUyyHLCUr1e1ar
I4nkJk+MJ6gqTNA9lKHqAWma/Vgp43/GMwdXHAPXM//sHuY3JB2INgzoUapjB6bXqm+MzmIgoRUK
1vZgm8s8KOm82jSPf9HAsI/dQ33GxiKNPGPZ/J3dEK86Ai2MlXZyVaUpvs0eoqT1DUN75eN9Bb3Y
r9IIqvS0u3hkDBd7+4XEcYh3qUAuvg3eCJ68pTAGg2Rz4AD+nt2xGrUHSVRkRQpKaMgWYJtZtNrp
hy1QjrjqGx2u6PDk1pAaIiMKyh1QASIEdvZbCZHilD0o9XfYHgvJp4YWxAud1n/9wY2FSsBgnxX9
md1ZESbs5fMhqztBODtXB0mtipJsaoA6xGoJT861UWuMLRN33TDSUP1D9FpSrjj7jJ9b2YeSIsYQ
Tvde1ChLx3DJfcQxT1hrBO2WgCpS9uXjzWCtddaYV4JAjhAh7fZtZGD7J8rF0Esom5m5tmZfm/zJ
mcFMGnhy1QLMm0gc3GdKANzRUngTPoLHoOApJR/j4M9het4Zm0xzA9mwgf081iofTLZHRXCtsqRL
DjOA/REAM778nx8n75UnkSjwAg5QvV8rT+4EByJJoaOwzWpUyJtv9i6scnUJMGiY7qjK6oxjbKbY
k+oZ4Cm2QCx0oOXUOIW2sWfFTbw7oxPky3j6YUXQZXEe0uoamNh4HjZO4QyUQEqnel49yFIBFjaw
Ee1oOAhcySnYOmfH/Heds3XZ8Z00jQf+VJo1ED0Z6ep5uf6nBw8t7Z4dDEhpugL93/q3+7mOIbSv
ZZa0f/ulBmjgYdyXit4nBfJIMPOGZ0M98+InMJk3tilhHwuNVSF1hJKPM8r9whmzH3hUlEWr1uqq
6l9kwYcMOBjoWHP9KRyWwSgAL6o+mSmgjMSqcg/b/u9bsr+yTpWjCIYZd/g+dskJxLTavbxKRqQF
i2mtamYGySSjen4SfOAV0NdUrRzA+4Hn5sFto48ZS5r7a0TzDEKhlsCz+Y3/MlTwxu0cPhz031zI
amG3SJLYYe1HO2+DVWroYjsTBet487sb5tB7roDVVR8jycNTWK7Qoc2C9/k7pd0xiGFv8uFga3eo
tiG11jyt8HggwSbegCjhDEmwKqGfiH01Z7d4x0NE9XISYSIDTui7tQt+sM1ihbrRpgv9vJIlL6Ue
eSKbHRpAQVFpxFwCsTe8ZNmdSIjqK9cVmlkJR6ns+4pJ/wy+YPvCCp+3NVLRRLaDBodBlBfhNPas
cftnKf3lE1wxWPgJrKRNCsP32QLR1Rto/HB2piJ37Yd8m2i1h5kjJO+IHHxngxxQmA5OJF46MzbF
QACIFzi6UJjJnHwm3SWSmH9dSsrnMEDfPXjs6HSACCZUbNz6vsdZj6QJ5Oa1Ihj1pF8m58U6GRcl
Nbl8azi98ll/pBw9nCVUhJGfngg2mGeBWaQrHf8ozofCgYIqh89JEp9FxX9TkCfVqlFGFYZ8l6lD
dVfgi4Yz+zFLu5LtZaTghgsGgfz+jVUSrZ7Vl3EEL9V1DS3BA70EDDRkamuNh3fMPP3P9L7NZCZn
YzvPAu5iW0Vs6gRUVmHog4ENe2YHGqZkHYJARxrT2YBzsNk+odt534dU4JoRefyIO3KD8lK/6YDJ
zTcXaiHk8PDZQIDQubEbPfZFC1+AOLB9MSqkwd6yWlQviBS8H7xColhBYdIV41zgz3p3ru0pF4f2
SQC618y+U/HWI1pSVvo6Uqv5E0eCUq054PeIliopRsZV/jXdLh7ijmQOIDZSD1mEBPqG4aFBkMJF
5ql6rtjl30F0x12O0dbKZHapiQCJrI92x6lkUKR0VuMxf261orexduYaTz75gvS9yKaXpMgDlk6E
/bPEJFilLsrc2mJa/PLWAzeXxxWhmD3HiaeBFp5izGb0G92nGbJXJh4d01xi2pl/ja/a5XPBNeSL
38asRZ3dY/wBjTxI3ecFqh6q39b1BSTedIcsfnyxkbathdBUDb5ff1CXEPo7TkzTOgTq6fe8xRLc
srsiAIejuuWpXUs39uP8p88Uk3BqCWeRUqylIuebB+iSlFRjHWn5h9f8qT30JYjwwGPIPxRmTjj7
LqZ3Gqqno2GnhpCV4NzKM+pMpl/232aSoh+H9g1jPC6X0VJpdPliDLZezlHs7OzAC1V+L3C2eAj2
/2cBclLIPF8h8pc1u/LvKOz8C6UCHVOkEwSIFvRIXzxYIENy9CgglTZ7di/f+gbD778fiyqi2kbI
aco07YFqBr0gyfNkN0EgDRi8rtYRMhPCaS+JprhY6Xx37Wvj1joy0LovDQRiYkiJl3UEnH3oMW+P
HNzt/FbFyBadBSZy1RQbPzFUXrgaE85d3PSmYXRIT753NrabD6bkhJDxhnBwPjW+aQyd8ub34y8q
HM0yA5xBu32o5NHPpSfAg81jtjAEPx/v0PdX/UHxVhI9UL5ccwpHzttCbcwYDFUdCbM9eV+SqL3e
0o4UIDDKkLOKWcge/fJKxP75dL8j9mDdnW4OWnIa3RacZMOw3D/KJWM7CGIm8HSLDYTQ2kmvaAXt
nbsWHp4Q/z+eeGRtHWpmETkerYKxPvCqDwTlMv3EK/JhwaJjmCTj5A4j9di5+BtIGJF8PbI3ondW
NkxDtPbTlmr9ZWmDts/ZkrxLPolgdG49l1dRG2uzpliyKw2QdD8dA/jNzesWvKJGgq8u9fVEST1s
WXBdeZNdDMuHg4Cl4Ai00uT+5vM44Jm5rQ528B3hzSZ0AE4v+sRR4qRVp55J7sOmYEQ6G281b4EL
rmb0QnYTBDooKTucIRnKMAH3FQHuORpnujyb8yJxmtPHTfRwWcKS27yVXvpD90YtfRbBzLGrwhX3
DOrCR1ylcIEKoU9uKebOVP2eG2ue0P41ps85Hie+Fuynuhjh3aPrCL8qDcv9O8XxI9zSaysslACm
cfEbnmHpYPZMV2OX/jpqG1VDosngLOg4flTNFbVARkBB4S2Sqrz5XaueMIRAVhVLUJ/S2bg20FS8
elcL8fAe/hnCZYdXhLpsyKzi6o8XkVCLZFf0C1dUCOXoO9kEPq9LwaLOoHAB1k/C6wkObmtR1gwh
IzH4Vf07iAsfnW/hRRekg9AP3af6+7Q1lDid1nmMz8sAk0qH4lGJdtfcaInM+b/thuxdPQmjxFvd
2FxYMbiKsSfhfZjtiSikJWNNk7BnrcJu9PIiMUCMfaI+UZ4ZbTapN7X0tJyZWjeNR43uSauYBSGH
rBqr5eMx5qIRc5I81iY4VXF8+jRAg9arPr6CIJ6pe7PALm2f8dLd9ImBkYqge7FosU6NJzbDsJOD
hPyE1V1edasx2vsHJwqOJtoXWe9O/Ije38e6zZBr3NNIil2fZ2RMKjvFsyZWuF3tfpXO7wbVyma0
9XQfBBmM0yuuf6mtAAJbXEtiq1wUf12EIw+9gQDxmTjQfVjXN3vQsU1GldNREqlAcuMbkFoif51o
d4hYYL7gt8iG0GPUCTv0cCs1rkGyvqJJEplrVS6OfKtB5MPucrj8ubMikuvyJSVtqxkC3GhBmIot
NDNZnCcga4R+Id9V+x5b/JUstcveGqwN3TW/vpt9UAjVpY7F6IjTD6DrbpABHEqi9/BW+6jzjage
bfKtiOXm5QJfjmYPlTO+LO7uEFkhA6qS/zh8s/n/3hgWrH0BVqn2RMdkmJJrRpHZ7sGyddPjrHc1
nx5QZ6JYsyPw8CeNqHnT+0TFJNI3OC7/HpHvkGbt4ynINhCBXAl2/5soqPIqC4ePt6iHD1UUWUva
S+u7/TX8tefB0+/qVvpR4I7w3HdjWzurS4riLY4t+TmJ9DvjiQK2xQExn6xe8ZXiZECYZUkperuP
CIpkvtBXaIvTi1djp0xvoKnOIC8xNCLHvkrDwghsbS8PTCVqJ3PiIhnANVZv9yuAgpsPUdDkTA1b
ByjBg+aeTPVHqL9Pn8rfMkjJed/obqebsTrkEe0+GSiVd2FJGaxgkVNbL31kWjfCMWRYOZFBQ5sG
ZN4jTHN/F3TLh63vweoCDOwR8lCr+rzS+hEqSsn140NFfzzSGwzh7/ajdbHUMOXtwgjitULieiL3
McnJ7Ay2Hpu/s0OLMkTVk+SecQfg/fRryujCtGGrFg2a/2eMcU6rRi0gevpWSwcWNZnKyHq22Wei
5hIbB+cFUWTqIeSK+twsdlTX9ZQGoibElErCPMUpsUNt6/x5S60/XyJax//BmUus95g4s1DkFy6N
/P6q+Zme8r02HajpVjcNCrWIglYzlMLQbdVTDzgVcfEDYXGLV+kSgBMqYATPN1OP3IhzPioLx8mO
qMJ2rVbz6MqUQ/XB9Mdzr+cpRtc6Ym1U4xtrEDRCWHoc5QOMN8CkKuZ0Rfqpkpj5p9kUJkRkH78L
ca0pu1f3NqgSCvb0IK8scvpMh+Fn0YEm0KRvQy5s0eDIuKt1XU/crOKDM0Ma6rXzHCffPNIkIJEh
XLSgLQ2SGEhUEDZHEKY0wfvvg5HPEaH9USCrlFldFpuJ/iCAA4gK9MUm8Ym814oGIkxxctxUc3Jl
1cx4te0f4wMom2la/25f0lQaaxqXj36+HfzFaVmITTJkm4LNaljq/akyr+ct5cWEo4syo62MCHeB
7wWIrV1J9Y2R5RWH7CQby/+fXu1b9E/y7Q3yFnEd3UTqQOOICOMej1ye7jkpMwmT8T712+eiYegl
T2TyaShZ90bMZIIqfzDkL9gOZTSkNKJl+kSopEL608U0wIQQl/TuW+hl4mfN4lCNzm/HJdB4qQc3
mTuh1zk5pwxnLQ1Y9emHsTLe3nV3VYPOK8zPptV3FQebycoQJITG/eT5PLthBzaxzkWexSK2ij+p
nk1yJOS0weyXUZnxe4nzQvtgCMzK1PHn63EBOjA2fai2IrtA/YrCQ6KEGGY1+Nj9XTrz3cNQNMc7
rBHXLAFexu3v38m3fqK/TriENTok7Mzs3ByETApSD/OGSYzGMX0tgCq8x/mJGrivU6VeVg+DveCa
PkC1vN8Idduv7oGmrZhHE1dpI5C/zz3zfQEYXVTaUfsLWOLH/+1K/Qe4ebh/FP6BILWBgU59jdZU
J8Tg3M65EEBc+SX+c1c45gX3Qcx7ChCS2Iohly0lSNvdZtbh9CUoQZuhZqdi03CKc89d8UBpzMRh
lxRUXhfH3m+WxrNSKlf2Sw/NAk8zBk3AMr9+BCJ0BHXj3f6c2iGGwca1qbL7bW4rzEYUkmFtTtnQ
aDAF9zexIoikQdfh6LRmwQQnvNYfWub+D3gdb4mrHvrfUzPnFSzZkg4tZvxcBaxIa7nSGtPAo/kX
AIO4D1EYhqzMoeMEija9IU9Vtwo81SSiMGESuhPLWKDsAVN/j7qn4Ul+ESYUFGApEjfEIw0FMFEG
ZZpzXdlX1FeRZBfuv2VNgxE1dD7CIkhnqRL5+DYAIxrhsGEsjLmu8Ckingzfp2FIT9tLYNgaRgtb
okOcfw2wpFj6GWStJeZEbrBCHY/pq31lTnidjo2ZwKIm/r/SOov954BoVzPlfsvXHCEpAfZM6azF
HModnPFcGBe6vy9cAU7HqZtHMc4Gd8xJD2j2FE5q+2uNRymwYf+/8S3ZtWkGuWzyysxD3z8E+Mnr
JqUmipXP4QsxZ6lAcZQI4QdFgWKuedbt91ovO2msjLYhx6Qf4qn1vezG8ZbwON0Jf0bpZ2Owy9tz
pgDaH0hRsbMqd0h3HBbO4uG4PLeKuUX6B7S42CesTQN9BPlKWEPB6a3clBIw56gch7rri6gxARbk
UiLCBpDBpxRuA2NAxP8CWsrI/0Q6DPe9U5t+aEwODVmF3cMbu+8wXG5vE5vV0Y/chM0LO2HoOO2A
+88XZJSRN+pjZf231QcDCySGOjV/ieWC2mggJHIa7xlZIq1RMFbn6KjFC6rOAB+Y4NIhooRe/7sV
R88MHU/8BLsEREK+0q5Dr82uV5l7IH6OkPrb4JNIEnGCWNPaBCR0uU1Y7ZMav+h+ITviHJloLzDd
yNyxE907cYCMJqa8Rr+3wmdgB7FcKL7QVCbVs3ka5nmEgf7lqW+YJ/LlQuspsUILSVk1ubyMrRMJ
1KiOm8SmLUQhlOwlQbd9JkPav3NB5u3VGlCwqChntBsKHXfzofqObesGmlYOfTabXr5zHtSrdMQ5
Xg0HL1FA9JAqokULHdJoXkk2fLdxzVE03gqoagKx8qOkwCpTh7KddN7acMWnwU0Xvy1KI9A5MXCE
7CK3hrd5XnX6Uns2mzjGL6utIQFbYU+/kASxZsZwpaXH2k358xZbKsM+X2XSG0e4irrPWt7NZqP2
HTjypX4l3ymJ/XBREe8zYHRiCUw195DFAcgjiYjj6dS1BX8v6LM0MhUjM/6/SSnrAwP7qUVA/bcU
myBrZmzyv8ZLUCC9ebUOkRdktVYZnNz4d/QcpiT8h0x5Jgf91PZDZ1CRQx/oVraEMs7kAskggLTJ
XGhAYjlr6p0Hyk/+igMlN1p1Wh88jWfSc6cwLWOHR7nFNTK0GfegUy5QLnmrdIwEWrgSOYaBMYr5
658i4EKTy7mqLy2phMJ/dW9cE/TYIlxtI9vYByZJ3tWJCryvSocoYbG7P/o3TLSX/wc4MZJSK1EW
KC/7yYy58RDXI3PzVjHDIE4/2F55OP1K+1Ng+KqnPDmTVe4yl0AOOpaGvI/tdJTaVcME1vJAVIzM
cdo+GXi8vrkjg19FCrUA/qOf4qNEL6irQQ3Pf1VCPC0UMoC9ecDuaBV97SBwuBkqTopfGtjp4MeU
Fp5M2yXCIgLybf6TiKZj3fiPyMYh0AcpoQIvEZg9KUFfVWc4AG7R9H3rS2bxMFTX9lGbw8SLON2A
g7lxOEZheEXda1o2/K9qvHVF5hMqT2n85WkLgX+hmTchOe4JoUcD6YOx7ZoTgmXnoKV8QEPYFCMy
KW6/lmH5tNVTynLgWkMWo3/xnC3HbzoK+X2qjSNnuPXL80SKBE1vfpG0/vGnei1m9QN+nVxUPYHY
DrlDMPJbDRQaioFUAbuURmNHW4aaSOFPQAJjyJ7CiAY3flGkuSutL0c5ej2Xyz3d9o0fyS9vp0OT
sEkJgQnlrhhfEfZdIrcdsxm0c8vP5xmHCP2wlhCfHOM422eTisCM/gk9k49DsKYTO90lnkDL2uON
Ohi7QF5PwgUxL1arVFvPp8Ymsmi6T+fhC4NyMFEE+SJ7cDaHlzJnCAJi1B+9jRxvoKK78BH3iUIU
I0JuhUBpFy4ym0d5IEthpeGOAONXga/n5QpfFi44svgpo9rCmiLn0k/lDn2hcVkFPfZkx/kKIr2O
WIHKmmhjNvf8Ow/r/iXGnpG//z/zKW7copHq+Uxn3dCnMnpZmhkWsOmIEDVf+f9LRzvQtaYzDz9S
U4cU3DIleYy5o5VX1TrReE9g8bF8kJxL6JHdkW3QdZDGQAy8koKcAsGxKpueunpF+MrjuPhcf6Sc
tjLia8pXDYfeMrs8SRvPtMcEx53Lw0yCsTfgvNLA8GPns043COwS/wyPv1pNd7+9LAnLloZt2g1y
TmHvxfKYHfcRCw6uRnGNbTkSIZKbAtyHYXmFAJxUhYxk+drIp/iMKdo6J39qi2TMlvNoDOvffr5n
bAZ8WKTYEmzlawB/vYGajm63jRSZ3Mu6DIcgvYv3DEKH/lFy7LO1PLMVUHcx1yj34nBx6RkmTyt3
EmANYy4Qm6s+sw7Lt1vb4tlvnjEqf9zWJY5LMsbsSBiYi9VpcyNSj/xuveFQVUpFIm7GjmRi8AAz
MiPchfwcVd2gNgv9e3lv+WmXe5JMWMhhiobW6AvF5NEn/N3ldML1kG/DJZZYocX/3pjgUMyNT6ip
QSW0hVFN8q2ATdArfI4Zu+7QKBmlO/oqH0uAcizhoiUaSLpV/mS62A2DRYiMdMn5jnK0lwU9FhxG
5dkeZEc6fGumLVOxk3PeybTGbhj3Hff9SXbauT7fMpFZaj4HOfXQIElhn6UUOQxjH+N2F/MfUPFn
Azy8dsUY04WFtd5S9CA4T43tkxfMJYCGbrQ0zolQvL0MSOvCsX7c9jPDEDAjvyosjyAsboRRRDmO
oYcuWvd8IgqixNOycSWwVnefZ2YStCDjQHjr2lcG7zNzjuTr7GJGoSW9BsEU3l+puK/6Jow6/wU1
t8qovXqcAkifxARrJ6Qb7L3Yt/iOnJUEQteU6wcObDNqZFeP8kJhFk4UO3aG1wXaqUelwurx1avw
VACd8gNMWp9N4O9vNOjtzZtZeS5FG5KWshXsyhXkK83U413keqNGMS1zU5VgPerZViaMg+eHyCOb
joKMVJy5LTwjXNzJPm6W0nuMzGQXWOaHcujE3pVy7E5tAheiDL9Ewq/9go94miv+m1GxYT1r8Q+4
DPDjDqZLqcNeuwm0MQnhniWnyXcnRx1b9pWFAvrBWajSGNQF1GXf6dAWh1AbTeQlU//8C1oWyLBV
TSKNJtzMSKfokaLCi3xHsWOzjxDzWOQGpPxfYtAb1f+xdzm4xq102CJm3vZiPCGFpJ5oH2P6ArZ8
d7HZw1pQUHYW0sHTK55u9r7pxhbzZB7330SruGu8tU80ZofM5tW+zhKXLTkAKeF0unr2P4mtpVPY
uLBOu1KQkoKdUhpIf9fUx4rXeB7aydqobgV+bbAoEMq+5y3KWR6PsnJ+GcspQ8q/TMlopJjhozb1
hx9GXIRwBxZaq+456nmKoPbZjBTF7Cu4ZPGjXCFYjz3XO8F+mSvc+fGCzV3CtXW/tIesea4sKryI
qrLhOpFDA2uDWen2YafhrAxUJ9zNG04wDswcImLXfs4WS2RxUCvJthWqA8fN+O/54sddfyEBLfpD
iu339PqiU4795uTK7tNo1xMbYMTSTIOQksPrVip/2fG/MVt6W9mD5n5usvP0nOWpVWbb/aqMy2Yr
wbNW6B3hJuQZUSfKnlLlRZM8j2ph5gWPk5YieqGac4ws0ryWknqRUrMFktxekd2Tvvwevzg7sfSv
p9SHLphZABuus0R1p5qNagjNmZGWBe29e6bpEJynPrm8L3xPfyqUxy8Oo8+AIGTOe3kyqJl29Ms2
ylxDUMo70K7FTMkL2rrKHMGvgDqWJpl3uoF3/nIKp2hkDmxQA47ov0ct4kM4uDjMtBCiZqOJcE9m
aMKqQmu7iYthkXTWm1wMw76XDHnJ4eI8/jZVmmV94hlEYDtg9e58KkiO/1aNmYBhMQWR9ezQyMYW
DxS+6nwoRdyLE55/aqX981xsK3AFnSu3T+3TwX/s92M8/kjiAUqdFdpak6o5tUyzrGVU9M0v7VDW
ewS5M+zTCvqhyuy+DYLWTA1xK8hiT24mg6jwPJVsNr+rJMxschd0ujWtzovVApD8VuWhsv/tkD7z
smoBzcmciVLMF+W923x8HStOlbiMzuJ72kLsQFx4Omg37jHvE43IFtjivVkmHOcm4uPJmR0WZXy+
b+6zXfnP+yx7O4xu0/gx1pQvfuQBc7i28Ai6Mw40fz4005t8IvvG4KrrK3pAdsR0owOT7QYLjDKP
p3qMKzgNUfkLTIzTHy/JUYla3OS3uwrz4tndiAQ65QvzR9gcAVMpKWGx5fKp2JPQ5UCaB4Inw0Fa
0r4pFvfZ1T/BVkQQEGd0uh721v/N1KvasjkaH8uNZFn589KJst+95PSVz9WTQGpgmIzzwFz7jbK9
Qgd9C1cxUIMiUoshbTx45TPw9QUnAwmJ13mXGw2pyZK688PTKwJDDLddyoME4N/zOeUj8xgKCpy0
nLsseKoJqMhVdyTK1lG2QRKX+1f2AM3tEWqfHHHf5nBH/y77Wcl1idtVSPMw9aN5Dem9Ku8CDXHu
84S2WgF4lFg6y0uo5uBFxrY3ljmfpLNoIF9Xj2VbIegwpe5M3WlSG3gIDpGK10gBTo492EZG6COU
3QGH2+1c5sZIFZuLSxNNsw/AzpJIHwWGkd6MYr+PH4CKCqWT8lUMPbcdq8V+fOyd0p7uuRKEV0yl
sTBzAgaseWCHrLfratdygBLhXUXSEQ1bWYBTCZB3UtSBQQ53+PXi6ikK3/9cKmeDHg5fbj9IpqOD
+Eg+9YaHvWdx9q9UB0BHL/t3tBvCcKrc+1jzYf4+2SUjrm/3hE9cjgYETuYCI4FpnWjwHkLhOfKg
aZtSDh1JYtQZO/F0gUvtp5FRek0vALvx8ASsHBHO2lv3MR7RFA1IBIkIctX9t5/bprQ7CulWEd7J
70Xf9Lv8HY8B7eAf0ln8lG8IFfiAzVXjuh0DGBxMOBEZN/tvvohHWwDW7/Mq0NWNuQZvO8d00us1
3BsDHB7t+zAu8tEkMpM/5s7zCZZ4lZIw4nDNN1zVqFfZSrSRJQ1bFXZAYcqO6BtEVryycaamXFvq
+6nD3AallzvtIG074SOk82f0loES6EMyODxR5mzZsk4CNK8fIMvL0F981Cg5i58gDihKmnNSGjXl
WMwTRoN+C+Jq7y3Pa1I57Wde1Ddh15nx7K/abuud8pLbjUyv3GRrJZkIqbeW5j+Xta8BygyDcEKN
dIRUikCEKr0VNfnMyyBJQPnN/1q5U0tuKOCNxYP3VhK6qeDifEti/c6o3WTnfClq3k0RyEP8nGVt
OvNE6jYKlg+sx4H5U9hnu76CLsWyY1fZZXB+RqKS+emUBa7ZCk2u2IY5V5EFtgcjwUhOnQdNbhw/
RdnRIrz8FJ63PhTrM9NJBNkMa800ekU/x4PhSc71EqJvvObon1p1tB401T77Ofb2ytNdcc36e/XI
JnSdpCT1sQx5KWDQzqSDrQwDu8LAhjqZV7DWVf+pUdRMRPB2VKmDarzUhy2M1rQxTaiHaYZSl7Rv
38kUkSVBal7XYiWtjSGVbDzB007abTy+rXhUuOzUPqPrB1OqMNwh+jJq6s/KYMemhBHp/bC7FncA
7tDRVL4wOhH0k29AowTYef9Hs1Ufy1+jmDpS/E0sGb58YTdGqfcXnU17DLWHJK+KSb5GsghTnJIv
oRTJUNKMnwLMnl2ziSQu5ZaPjOqAtc6FO9l24/1QYeRGqVlp+Z4Z/Yn8fVVLZyKnjdfSooR+ZFx8
DETeyxBSAs7regc3ByRx1aSdefpC4uUOrLdmrjSP+XX3/37Ll3L1+zA9tf1Mpc4Ovzegah2+fXft
jYkHk9ab5gB5EBGQJs+f6Oc2YNgPpns6Onz1Q5V+EhVWmwv7RRTqk0xv7N6PInfbI1iYJ8iPWhNs
r5piojsyd8AT5yPiyfzd9sZLQlVUi0ONSjEijOFEG2ZZnn4f+QATiYydPVIh3x4MCGg5b8JGJw+p
7bKEwQx3q1VuiVe25v7mcoZam62RrbnPhnOhnGBIjbZSdvbubWP6nenuZe6EkdR89C4vkTkkT6C4
O+uibtE9kyQh5EdSbIS/onzjwN99fkVwMJUyfKHAFh9+PFWalb2efdm/MC0sbZ0tozw49LAQt+Jl
m/HWtm8hbd9ZWPBG/o30V9EPIjv3HRudh/fXlbPTXqzOHmyoFbKH4hY4ZLnYuek5lxDlYECoCXrP
klDBeaQ0hNz/36yX4uuutQSAR8wc5SRfx+Vu04RBpnPAJF+Fan88z1RcnOSEmqiOfhsylbiJcz46
Stl+CYdcsT5BCyoJHT7d9bST4KBLG+uOnEklWfFNz90zQI4p603TEKezQAQoetg3nEeQ5sm4wXFQ
uzKujnpDvwZyuxdMTa6tRWb8tiLhxlBjxxzN9PELZ2sLw+0hLzfNsz0fubO+9SXwqMFefj2ZAR5d
GHavQoBXG4eWwfjOsezcmXjdd3YjXeE9tMr+/nA4s+Z/ADhvXqqarFdlQVgeF5Aqf6D1dmvL+nPb
U49oNK4TJkk/3hqfUmNsNxXEoGm83zTCDWPFrS9YIRTCD/OKXOzaZlMIYjpdG30Ul1hFsa3iyaUk
PcUP7PgfQcIzMMJBIuLT4bU4pgRQuwOQ6S10oosqEPPO/0YXZSkPwPnQwIC6/EKVNTjCecAUO4MN
1Rwg5NXNdfs3IpCqUwZLD1U/raoGTI0ACPg6TP7X0Acd8gJEFiWQrSOYnttfdDoO8iPYdkrD82Yx
XQ7vrlqsMrMSy703gy3hpkCP8bGhqJ+q/fndGY9IUwg1rob3NRTVLNHPyWgOGBfvx1yAYWgpxOZf
HgqJD0RjlNA2i0gMc3+BfC3IFVd+K6Sfqz+/Im9QByMmfUhUItOmTlafrt5MH6DGuAZGnPrzJtEg
Eok5ZBMdudaHo+Ez4k/6av1plNHUcUQnaB1BN4mmQpC2rRy6nrBrEGKR9QRv6WBLJvQe9NIBy/zf
qSmbgdXiC99CmA53dUr7/ww1b4akaKSQOuheAMOgJj+JX9lVr0ZRdrcyuqWLdE1/9m3IkW2ABz5v
HAWXXaqtnVBaRZXvieiylcYUEcCY4+YsRK4m/H+qAy0AQNG6uaA3npt5NdlvyrfQQXtUfc8s34y9
tXJkWr9wSF+idCewS7CWaM4iuDg95jy0R6Af8WzCyv22GJiad8XhFWbIGxliTw/T+ZmrL1LIkkJc
myGQxGr3N5lgk7ysjQZzA6Onsf4FDVGNgw6DvUjXh32dVZi4f8VEojvBAXGhdTuwTD+Y8AUiqIsc
K/xTp9HxlXLr49RL+wN/9adqYHcKbECUFKP0wMrOUnMqJ9k2KrwZtsyfzd5VyJ5UQZHByQV6NNGB
YOWrBhsyHG2tR1hoLhyKuvFWuoGL/yhrh0zrvFvxDqcUD8nSMnD7FgnhtNQ5N+Kd9HE132uKcXob
P3FagjrkRUo7OXuw0OmA+GDoiYzuin4RwyeFWU61uqxwjIdVdh7CdKgpLBf3f5j5utwPByqGgvar
g9sCn8TsUscURmcG3YLgO8uOQVDEymwqopQrHkLEFHKvXlt7YIdcpB6ZCuaGDsNgQttEN3qxoyuc
1wwnfm28WzInmuWftY+naknU0Mx8sZ40W4L0AkXLOrCfIpy+VntqdwDhoemjjRIiMbqvwqFTm5Xi
7NQiZP0u2Iq4wnUZ2n0q9N6QrX5OS/y/+0+fdwZtrPeZOZXQU9bKrz+QAd4DR2kkf4C9G7xjGYXC
zJRzWuZwnTsMCJkt8rWRMG1zNElNHLxHZBxevgJi5teaGjnRctPV+/KlKPh46N1U0doZg9HUQF1b
5OvajuWpZxDmGlZQSg9e6a3LBO/qBjJoggXmhL9/ioH/c5NtFagIP9oBLkh/3zXW9+AvV4g53JPr
+XDdVGlPwqFweLxs0ZMgOqtX4y4grKEs7KlaCcJt1AozN4HYDRcWxtfyyzaxr1bjhDK04Jp4V+Pm
+ghzYuIc5lto4Qvqevsoxbdwh8UriJWerbPQ3bls7kQUSqTumyodRiN6lzUQXqHTWWdUV7wjyoB7
diE/jmSKpSZCW+ps9gdvBANRg2cm/LptLO7n0KIRh1WCasDmLwr6YD2vDtfUblduge002IDEoJ+w
55zCXuYIJRdAbvI4VGNzi+BY1IYPjupMqGyGk2wJ2fTJVVnZ9CVhITwoo9YhY0qzm/zLJ8GF9kwX
9uwXszw4DT6siCo5cQvl0pPUMl9+tlgTrVXW9rcBDQTLoh+R1hT5NBMzxD42WPENFLD5PtgUhQ0K
eVW9ZRktbKFwKgTe8nQlMR3oF4tyzWL3Hoolc78LZv1wScGDcsIomfsDgfhreYOWImyUl57+GkiQ
5Sq7sJDoaV8lqBgH2k6dfkiyDHd7nL0Kg8m4fbRZbdGeJporWsu3oDnG6OLmrTIuEfn75nomEO3T
KSeHvlKGLvOC1ewZRXIWLU8dpJUzMHv7FMzwxwT5+UusggR3bCYO/GyYrc7zhBOEWfX5Edr8JxKV
K/XuNShbjU49iWmnBgh8J3yu7AFzo2FyZYpupTXXp+6WPFOC4RKmmCs5VuzWClY/Sapz/yH5j7Wf
5xvjSRf/jNdCREodkMOi0RlvabcU5eVDSCdwz/l+AKGDD0ONajYnHPJEtavcrr0lGvGwsWBOwE7J
OKIMwTMPU/6WIc2PwoiLvTCsFetfedZrA/mheipvmI+1nN+NYgLWzBV1YLSXzrNBHcsSYDk1SUXB
/nwta3363LDkR4oT5DtT91/27e8wfOknXnvDmI4H93LIkFTAjBuhXvgI+hvieXH9MUa5eB1UojSE
QZUS7kG86JTiHxLJWJ5pSS5ZB77FLY2dxPu1wtYvBZU4BeHImgOS9ZyRbcInlBt9zu9u+1vgIUu1
UCxH8LmLH34TZ4nncmzDUUdlms38PvjKj+0k/pnzVBeprUyfqT1a7pGZRJu2P4893c65RccPyJA6
zsT9hPHwm+WpSmI75nhYP7KnmCnYmnDPlo+Ls26P+Vdkc0YQGWzQ0LAfPPLx7IAaGAZyhvgzRh4g
vMKu/H+k0HKafT6Sx81OJCzNgvnBNBIwOyotTlGwRQJWRk9symQYj+JFm4zl6rdw70Dv1eO0PKi0
e9ui7BeVROvZOll2g7YeoFDBiwzn6I6E/24BWAQbeCQUac2zq1sHmn5mQm5HQoTB3v82uFm/4Ev+
ytucre3p4LpAtY9q/Ie02jLtWvBtgQe+kddCgH8/fN+9kYwmG1D546KenfMAA5Wzk6PXjzzWPAnX
zHxb7nPCZAno6/wu2IjbmD5EFrt4mGqsixrvrp3LuCzRJL0phajPWsJVd+T1e4z2xVXnOG46K2bK
vj0hPNDGHHMKQXcLZi4xFc8hPyTT3UXI/cyuU34A3IV1D4caFWX93TRl62WQYwDyfqFC79JPpKHb
K1qEj3gJaoi4sMdElpr4KALpU2bET9L499cyWtZFnbW9fcJvqXw1f6rbLU6LNm7z2A/4zfRW81f7
n5AbzGYWBcVxn/iszRyzHVRiESOOkeCuITVtmQJkzn4XjSnAU3VsvEOWDpo98FdmL01/uU4vLzfg
ph4tmzu8pMgekFGUt9LlPH/tmv9lumiFAgPpQfnpheqAgm0+K+vHGuQRXr1F0E9fS0feHklY3cXm
yjT5dwKiD+8xiC9YGQKjxUWksng9VKa92XPYBrPTykg0/kCLFypqfMFNFAu3CdM/m829BbWvDCdH
dumvBSL+nIXaohBll12KD36VTjA1DI+jtAFKq4pFhEkaI7dBjm8cTdgoKax/17LxackEtHPNvBbb
mx/x8DJuUUymJkUR6/Z5C5tTWXVU8tZ7V/H3fKTNKH2Wcpx5F2K86ItJmhsB2gLOJ2ry5R2mLXAw
z3Hk4Rhe/V1zeeedYjdJ12kcBmtNuigux7x0v7B+jcIOVx55c112aCeeAcDn+Z6pbw5kb030QvXe
Di3lryOaZ0uo0QIiAyL9tyQprlgJLBwMfl+X0AUfZZe8pzBxvc+SzvEdmXmoze1nFybW4YLvBnMf
Im9wicyTwnfZy3t3XXCJb7yFaecGoPNS5PMaI9i6jSJSwIbVWgl+Mbljz82PRn9MPecV3eKg+MJ1
wq9+xru3VIY9WJg1l4HgKZfoe0NnCAQPJ4xO1Br0/2IO/wAW6Ee4yFLQeQtXTYbpvnOwnED1D/MF
D7zjlARI0pvnQ3umGlORp9ng1YklvtxrUDzxoe4MePn6JYojTNCLxJCxC91J4jGL54tBFPDce79k
r9P4+MuFCMjZqQPQ66lTzLnU1m0rV/78QhIISwCL97lvBirkDgSmZOSpwT+v9cdSWqXn4vdWRJsC
87Fh187ykPuX1IUDuz6RDjigOqTkjlDQmcbuISpb7FQMsrZ1hxfmdEq2IsvtuL0xNOnu8b6Bw+Sr
4CyEYxRVi4x3NmAi2A6JHRrfDbBob63vEblRSpQYT5Y4v6RN7UrIg5M4S0zG+G6UeAl4XC5rFgNu
SkpGKje4Ftas4P1Hih0ngmEeiFWMIG1LMGfCguNYPqNCb89Ak2G04z9My2L330v2w/3aVaNJXifs
wFDUCmebGqY985NsQzTV6WnUzDU7bR5hS1lOBwUmQ1oAbTJucLYP1aLoLgU3V2WnbnqL7OzUeVrI
X1mMr0X8qnsWtQPfMasSDHypLG32HF98wCfemnDEl4uOvkziXU94E/L3sisTewXH//S61K2NaXn9
05cUkPUm7aru5XVGSVRX8n9P+rgsyvaaM1E8XyZmgg7dh5mOF2YVGkG/hHkPhXpcAOQ3jHF6elKT
1iDT0oG0hZj1T25aqfgcvVzVzVjYnjsrPj77kLYYWm1QqqRfTOZnmy8qAUhSXSFIXu1Q00mMqZK/
fc6k2AIHoYbKLp1f2CJbNtE05ppnhBccaUWCzK5938o6w5+wMps7iPl22yUFcl/y1KKwFN3xH6aX
0AewDmJ1IwRSnIbtqgZpiNtowJS8ML8qxjdSkj8NMw+yjPigyZEMd8RpG9NHpUxhZ/p2unjAqunz
LTrCTpzcMPZBKsA5DtKjmNWs4kPtxrGz3MX39xISjUWeSsUqRTYsT1WGkN9V4YrrDmGiOzP+9WLQ
Dq6s2Bow+C1NtS6yrGhjXyXF4C5djB9gNb/XUAc0Ay61caoXmVHz50n7hK8rkzmsKnZxwoSO4ggK
7byhJ3Du7X6POeyKKarhw5ZZUt/vbjU5de2hFlWXaaweBKhsmx/5+3MFAjrayHGSzmgKe3J3cL1c
PAh7vHtOMZY9m5CgqpJXK3S6Uesw5S02GqZ7Q1WH2WS2jz2g2Q9ldPp25WCEl5B8skd/y75EWnND
3+or7TEVflSZbsqDlCnoe1rj+vf97DP2CnMBMTdV+A1+wawCnDwAezVPjQ7lB/uoxmx2WvoAopAB
5I/Rpyp46bH4oUzPEXRxXFQwzFxmkCuQ/ddCHj/AZrof1BCm3G4XtXFQO97YiYjNfjP10RSQzjje
VmN/mt4TrV+SVpO+SjGRmetpH6+T9WYOCdUfgA7RaJ5yrSYFepV56jOTwFg2TcNY2QZd7Mma6Qj4
UCwuLGLz7c9rYzT7eNXMBNOCH33JEy3BsTHan9BEZfE3R5MztNREUbYon8l2HKFIKtUj0x2yghYw
8/dVzWOu+G7bPvpDZ5hGHNH0r7C2uEHCC5b/g7niParbZrylsREPQ3F7LbqacpKlrrY5L1jgLbFy
jKAh9j5mar05Wk338/HcLy1fcuQNg1FN6rwId2r80c4GehWx/05GpdE0Ov4oGPj090TaxfmG2oKl
G00ZsKBcQ0aQpdjcwq6+YLrvETam7WIBApW0hqOlYcHqm+iuHPGuWsaFaH1metsylEquuN7txGe5
bNqPsQcc4AuZupoB5lgrckW0D5Qmqb/asrv6Y/GRFMqxm7Ch0+Y/qNwOBOePqTzV4O2CipiIozXy
0l+b9JlrDgpvCSGuSei+WAjkpt0NWU2DN8emzAb8i+qQhicnmmKpz8F5Ro18FDeasFBwrPlwzm6t
p5byYvEhG3uYNFO361oYhIDelzEHjUcqq+yXBvRIOsyXfeTYXZPh6a4Rh9ZP62rHn7epJarwCS0O
JXPFEOFv5wzrUo6P/A6pUQJwvlDwHfjGMe0ud8CvyfJlLve8hdW0/0zTp0eVv1oVc66cEUtn95y4
yA9wKKuVqLOHKj4XDx5DMPSxfJ8g4kr0wDkAA7yIcHg5ld4VO5m+gnpKNA4TPOC9zk9LTVKGaYJY
+xqEWhrMw9GQv7ObqoHpwIimJcrStN5EZG2V/8ZzRuJLeL5zc0PYSU6bA+JQHmCkquMLTZ48Wh3e
rFYO+297c4x+STJS212cTRK+kJq+WdQANn/lHeSvD4CUraPKXIfc0fN+r3torPOfZ5GM1YhyIfX/
ymKKMPvt4QK/9ly9zlTPo2UMpAOzcvLHjrbibyuT0pSm1+P+WUpzqsuefJnVScXdsgragkUaC3Cd
1gd0DoMKB8hO+I0RvwgbpSp6Oip7LZCYHobC+vQwVYf/wyQsK8h2bhsj6iauCZNsP2NqnxYw6MfC
o3jx0dlw7g67U9SSJol9zylpvdDadEZzcf+v9fK3nuPxaKsOh7QCay3eHLU/bXN1bWXKw8LhlX5o
ToIUgyqrrUeaPgcj+hehBLOvrev/NqHgF11RdZQd9OayBPULYJkiD1A0nf+9fnTB5Jn7itGi3rHs
59MVMy/65hw9kAXhyd3LhRPGIV4xMye4i6J89B0XXdxg4w/7iq4hvnglKsqweObn3DaooEXnsS6X
JIhDGNEZkVIBDUa8687cB200dkHwFshWeBnEkpzFgiU3ks8g4UMwKeSbEvdev8Xq6aD10vHFO2JZ
9lINbkNjIGtFO95h1Mh30GRKTwUDpsw5ec5Yk6JGIM30fMf137buqVfOjIHntqw4vRs403QOfslw
f4vhBm06pjx+ae4SVfib3sfKRVPCf7kL60Fh7FqYzDWZQUnqmS15m9NVqs09NgmBDWBNLNtHBs6x
HHhnsbNuE9vQAjoF5FEmOZnUZMbZFi2rrCGXXDMAQteWpMHcu9SahgZTr9HCZQMMTpuSw+L6CPog
kTLwRiRrg+LyuENI+gVNCMexje2CUs6G5D1Xghhuyd79di1a+HLDjD/VgSPytu2qrTmBkGAGon8Z
3CzXkT0/9CY0okRMu17LfLmeSOoplzGcgIp7fm5ZHUnmF1t+SCF2GoCnmz9+XvoVZTAvuOMfTmOm
e93PRcNoD3zHKba+1ySVXYDJkiXmeAj1UgOfhhnS0gyOD0jFhcqv9g6mZxeaeq3xqpQY+G6KL1WO
1PYLSfFYHo3x/rvKwUljdIQIhhfbk7h2bzFmEEo5+b9gNDnt+txD7a4LOmkKj31onYhiMb5kNXJU
5qzjwsMyRAIILhx4JxspsrbYfTRDh/ovUJCxGd83iNWsnTrWAe/yWUKOhiaQa3yLuEdOenHOB4rx
DvT62WW2dXE3IPV9Q6xS93puqz+zXFCWOyZKhv4EDbndsP0K5DO3ywmJNpD5K4FeIrUdFhDL80rT
4/RBeUKCs0F7IuHiJCvntOoXv1GscMKa/FPVhQK+NgS7E7R2lKRJrzcv7VuH0eKcajSUNeVxAIXD
B30E2SegaZdJDGslHEFWwHCjRYBrUnqpdw/KrH0/WIQIzfoSG254ygbYalF7BEEkmCERn3yz2rM3
R+KkMsW93KxYaCbeE0xIDTS5Bq8cD6t1bnl/JG6ujha3XnR96ZUn8jnhwKhColtZ/edLr4q3jfqT
iCJjbp9fdz104vJzEx0MohveCsz6wA8n7gSg+pIClF9PqaCf3DLKsXfhG7O6fR+hpyskoTCWS1Lu
YebU5NKRQR7lAQti6GyZZmenlTA9RoaOFOXTY8e9XKIjXoI7CJUV578F7YmoGBX+fWxuPVD2x5DG
neHvTPoql3M9iIGevPVoyhjT1eXOQE4tBzc8YhcKEuowJuZXwGTIVziv/OtESuGR5u7lmd++ymn7
4p8lsIZwA4OomU5aI+Xh+AEbKKr/UI+p/Dprkxgr1Vzi1LJFs27FwlU74qIF/QJBF2BRSoSONcKX
8dwL54+Nc6uuCD8qMLzoIs3OIoeXIffw6YIvNoquMrwVc0aQpvAy2B8Rz4wr+Yj/jaBcUu6FzYWw
uRRS/8myEBBWxVKhUwDDcxt0BKmuPDhO1h7czijHkFKaB5W8PNksaZCI7Vgm0CpB/pTD/CB21s/h
7BL+TIzr4H867GRXow/LkOu+aYxxXdKt59BPYWERWWbOqmEGHBA9e5PTkxfs2p9WSyg+EGTxqH+6
XJsMCiUv2UDL+64Bywqb+UdVD/ozG4V8+Janq/TnbxZYtoTlrLyCGD3wtNKKbvS6C42liUEJv82F
FWXEJv1J5tOd4CE9EUg75P7vCC+muf4P+8mZLpO6xDh7BI1NfFiUTFtqZtXCzdQA4mOBkRvaoaNb
DIk0vw3Tar5OdIV15j0lmws/i47vv89024dNo0edBSzquTduqj08lTqAc6PNo6YFocwguo06G2RN
4ioCB614UCW/P1zE1PF4neKOz9Qgb5vVHVjVurG8pE/cmnRXXcMaq9b9AR2QdJldnM7APLuSxPwP
XJfly3vPIRbBoF6ryk4BkFJ1P5qZfABP7RTJMG6d/FZvYjrQu3GqNxlgWz+qXsUkqt/tEUJnWuAB
TXTQYw58MCn3W5f3WSn0zkGdqygsJNCP45YNaelfXoAoKoss4oM2fS2yKtAz0eaTwasjku7rK3eM
hLPw1FqHzvqmQaeYchJSglsTlCi5iopuafyemvVVxyuFTuedeQFt6hZw0VTAMuYSGfuh7LO6O7Ll
sJLeMbcFl7HX1ULLbikuZ8L0MTsm8iV7jBXpoGfxzMJe2r6QP86OZWJekztnC/Gd/65lu6XK9Mih
iUfkThp5jrEdFeyr0/5/OrwCtrrC+6gxPOBqh48Tzasyretr8gI22IiIYXTJcmkr7Jth6Rqu4gxa
XchDXRn0PxJXhCEjqDgMBEuNkGc4Pn8R6VZfhrcMJEQlD4DQv/0VC7qRVOoS3+KtVLpOpjGsco7x
+XSgnj6bE3OqaLFopUpc0d7OngB1z7tpuqxDG/wz4er2JKSbTSZvhZLym5vMsuuVgp0c1Bl6hgpb
2/xpttxtBT5SJ5PwK3TY/WKYvAH+Vx/eTDOe4PdYgC+fBWUFT08GgixjgLgaUkz7ixAtl86fbckh
g8l0ptmQ+zxfJXMXv1Ozz+SSwNxSThfBlAm2KlvLxOVVUp5cfuTZrDtDlXpUTITfYX0Sd669+bSL
7PF4nVBwKX6pV9KeZmXeJ+iStip9ZaF+g9jpL1bKhArRmSZ/9TzKBrJtZw25LavMsgWrjPOXU9Gn
HmLv9C+jHNmkxN5uePZc8fLH6u3nTragZd+iJLLcFoxOOBYqfS7Ket9OjQUXsHP1b2eKogwAzqPD
WFLfboL69Z65bfyLaGmcgW8e4oX+dOI6bJCxi8xWhh/kbUQUz8zEauEmqcUxxrZ0sK16G87gH1EE
xI7TkgsS7uEhzXxh0xUYpfVcrBtMKhkBhonJBmoHfcfi1ukkKFyBy7is0DkW649sIFuDjwosjdzG
hwaGPaqm2k08sys64s61sjvJM3xNkR2xMSY4/68rVGGCNZqO36vdztLP9mSh2diB1cVdKxvtFuSK
1TcLopA/uorQw7y9WndKmxZ+lu8qYKUfT2tN1I3yt05z/T7DSipz9/CpyJ3Ss5e0KZeRYZRKhKqm
8pyCZRAVgJ0HQJX0by7X5P4G+0H6nL1O0MpLUDzjDapJenuC2F5wdp3NMOLoQYFd3Gyr+M7fjv5q
nIP+oX5hLk1emUpbPbRZHe4AFwN2GKRRPsRjTsMGPsVuxUkTuRH+djHWnP5LLL4xChKpMFZpjYWb
9gXMiRHoPu1RxOuWyEP1IWchU+4jcUU2Xm7aliUT5igDDT6f8FF2i27hSopAhKDXwU4QpCqiiSPL
T6WEFmNwa7JxhGrAhvaClLSr/v3f21ZSNm24Et5vndVMP+yUZbQSV2aCqrwUw5mICKG9TxMNb55v
d/MMOPKFd9OQNkUzXCBS6t75hhCyB4+QMF1TvNxnO+NhsmBHJOdc/DBaUm2QKy8aGlrpXvm4B4Lj
66qiwZTQ6YJIonRcdEbqtVVHAw9m3LuuFSTtGvZ6i/7ci1EliNq+dTVMMSFEQAb6jiirsOBYWVSy
aQCoAv6NR8vhdM3RSIyeNrtO9gfYf6SOkPh+WcCQuFMZ6M5x2AawCnZiWagjQ+s8x0hXhEXULRHN
iInLcBHlnaZqQ1bxTvNUiPghJb3as6mZhlWuoPNzq0XZSlFKIbCmxr4Zlfb5aboUIpBRIcpRzTvZ
03tp8mhxayHCBT3nyoI+PuzUtpsq9rt8UAdb3g+EH9BNFCw7v7VwmMraEuo7l5jKD0z5YPFiu2+g
zvCEQzDvbCgeTABf1WOj8+c2HrDmsqgUUuRniDoj9tHYvwI+z2gr77lgt8eDawGlO21T1RzjQi6X
TX2wzFw93PuL7/ghNfxOndvvLjal2pqDwFi5LpIlCh6ECZ9seG/gZ5B4efhAHU/fSLj6iSM+BU4e
zOJmVzRPZYCn/lSQkplZ/xfspfYosATgDh168cxXZ04yuAozOlOUTUBznvqhCHri+K09GZ1El3Yt
jU+urygI1LbFDxdHLZyPi2xlhQgt7GDsUyMg+mysz9C5sZucgrb+xBSsrLazYUgVhaelkVPgbI4c
5ocJBswpx+15QhDEp7LIpKtqUmUV3cqdYAAL9RrAfcbgm7b3mkshjpPLl3IqmmIN4ugKzxoLjPrE
hDS1TkSzt5NYfESQzn/VJ5DiMkN3Sq70NmWk5Id383/vxP2QcTnleTj9XqbabaUIkudGpJLwZnPH
mCs+ADlFYxBtoW1lBwgsx4c/hn88P6dfCCPxRUxF2qXNC7N0EXPTL8G2+SMJBuoaDLq7BDIBrbF+
A1XfOJgKVzpGJHD1F24SC9r/tOwV7bOiOWMx3aB+HWGZMPweSkE5pTChcsU61IkJ9YKTXp4BFrxH
4ao965i4qoxIELBRVeZiBvwlA6QurBLHJFQZ5Ty2+D3XVioQdvFBuOgjL0dl9vQYrnWsq/YlFD7p
dIUtZjIs1PPHBfE8fYuEJHiHcIzQ1Nooa7gXiHtPzmZFY+bffQNIhX1iOvNe4E/G3h4PjBLNdXas
u9caxkQHYUGvC9nU7Rr3QPdsyZqZW4+cA54l4+vEEoqzxmavSewmM1WjErNzPJV3XduATqf69djB
ByMSQbPCklCDn3bC3DaKerbIG4T33UN/zSdScuWfr6ruZe3jt5MBUNfqCsmwr2BuXzN6wu5GsubO
JQMYhTagt8pC15Enst0V0nIgduH4BUkYNB/r4RZcfBHzxYiSR28FfhlYewwIwzkUqRHtebUAfG0C
WBT6edqNTTvzohm1Cn0AoBsBCQqVFFtFAuLzUokFE+PCvnsckyMi/tmTnjSoPmlyNrupe+Cofe5j
HdprpVHUTmOsxkM3Y2UcL39X8PUrcmCEpwLR8wJrraglt3cXNmNHbGwXPEwM8yPHP02wHUnNhrAe
4EqwqwITFqSfSFvNN5CkdWiEHHGN6l1qwV69J34oizE+FcMuLZ+AA5G3KTp4Vt0TV776C7v/Jc8v
05YPMAeiJwjRpDdQLDDHjurNVg1CeRXZ0n5IQaU9PCyhZNDkeFkmIDtwtA2cNZ0dnu/3f9eCZ8ZB
WvdcOWEAOYkpLqFd6MMhBhlUYzLROXhi9pJ1RK7VBUadhui0QBIRXkVcYHW5RlUexGTCHunvFFP7
qPUX164xFO7rMkQhS9AzW+hlv6a3wXEgagIXRLtC6w9iodIIjMyYF3p3CSFOaq2LVNot/ELVUM7W
+ov8lAnaJhou9fwtpJQQeM6AahQR6ZaaMPjLU4NgQKUjUP8ukYjRTyUPe/ou3NHBqez6GfoNJ8K8
6cGcKSOzV5Wd9FadagFi8Mz2RIqWz4XRKHP6GgGIaiEnSMVs/h8DQ/uM5t17rE+atgf37AlO8Tha
dZ0aIPYlTlSWGGyb4RnOoKTNIpC8Ocj07qdhECb+IzCeMLPpmHTtgdvYDy58BY2+HSbpYwfzrC1o
09SDX9PeDF9sLYpzCx27ybygCqpUpxlAt7jIEPWzCnO1gHDLCm1vLHAZ2fAXVtcmqVvUyjtiGLci
5ixH4YV6XfbUwqxRPK/Tm3byWvyxSJR+RiqvMIdC2poKUMf/EvalYOjf7bOnYvMGg6SBPj3ulqVA
WDQ8gHxlR8EBECnH89R/IGtno/fTlaJvkENYLaf5LtClXZayi74GMt4GLrSU7I0sdVBBkvth81b/
9/daHXr3FW1JEkTYUK09SzZaabENOGDrFaMEAFWNyag//MQZDpDCqUk7y3z+W9nYFc8fN8b9bq32
vGITpcKcyJt3riCJeG6aH8DhcJQV2fdc/Sdc/c7O1jey+XZoE9FNLWb4TtZLUgl+y28WSX19hIvt
Hj5bCZTGAqdTGl7dFDZg1pBA98DvQsj3ZivuaD+0Y5iKQunWQsAYlYuU8lqZUuiPXSZl+V5pllVo
2bVQQJiCcJPvIcil7Fey1dkxgvDzYAMfwVfKb/Tjw2lX9jW5K6xOpV12nBRVRul+89ZitQ2l/90l
NkBr8jCV+b2RecNaJnbcgauoj3C+SiyRjkYcIEY5ApdspjQvnyiFYWThjwv9r30W2eahF3GO24Wh
evWWILqvQqO3MPw0NMpT7caqHPO/dMg14ohcQLFY0Zc8LK6ZQPsW1w/qvu1Q3+s9iHiSagUQPGRc
QfaRLPLqhfPr04p7dFDoQSNZEcabB38KX6HZXkhYRAaTAGtTUg8wPA64lNd/0iIVwKvvTrfmjcel
oYoPzZeWI4JBqVaEA7zpEZQCg1mY0emASkzQQJ13+w83AVaE7dxOMj9KJJRt2LbQpRsXaEm9ADw1
YD9XNqjE08JOtYVV6S/8vdisADjfzKORrcDFPjx3VY8q6zHkjdVgNjPhO2knL1K7jWFuD/LUHylf
EWXBs5AbxxD4EMjUjge1St+qhKEIbwBQ9Ov1tac9ksHGuqGOP6frys/Klt6u5WdcUFu+USUo57O2
DCBd0FQAKnvYpJM4zY7Yao9VpKYJ8KV0g+BII7w4RLA/AHH4KhUxh2eEUn6dO8/zF7P2Zb8dINPg
ArrYF9n/8mF4+DMmLWXFlPpd40LAlFjnxTKJiTAU9EknHpuo1hma3JyPC7IjNz3hTcn/gC8s2KtL
XAop2FgsXR7/NZ5WqyOvnq/wcKJxbsjywwBqo7x+MTOX/dX/jEIgYK1eEMzeMCLY/3dyEhAWTlKg
US7rA/jSKBW2S+C/Cr+WdgjCIwdtrQQqZlmKhjCc1CC44E1sqEBvOlTudG1GVVaXJjvvMLkOK9hH
nhLzmzPnMpC8LRmEiEBt68oM08dkBe+MqYFkloXQZYKBJDOHPdjx5hjU79D0wrAcoaMbdHgxXlmG
Ne/AJMmpn4cFdxf4Y2+h1NbttXAEBIf2p5ApjBhE6+d7VDBq4IFRoNNFTIA0sp4znY5gk4M61RTC
wHyAt9gHuJX3RyEAi3HQjbKHbW7TZ5qu2agZCck/FeXwo7Sd0i0TLbUxOmNHhlFSBfV1CT/gBurD
mq3eZqfjtDw83h73amX9V7P8heuhs8jS25WKNYU3BSqrJjJf4MxesQl4KPpsz1m+KPe6tZ1V5sdc
d+bcp8ytUdeWxOSdjRAsE85LWKlercMjOtiu1vFkn0q1cLIikHa6dhCCw75IZh4YFsI9TuBuHoho
ftVlHYsBJsBApChCat80afv0I5H4REXZ8384cQffcXWutRoxcU3r98i6+FtCboDVf8euQQHKrC9+
yei0q4VufZVcJxvC4chNLCpR2xeKaqCo6Qag+BVzoXgY1ec6kEcc3P/VN/c4nhooIVQMckI5BwhP
aYz1rhdQDFy3cNT1YaAzubcwb7MtXBXR2p4IOofgxrAvSBvaKeowvLCQLBF+x7fEf1ci9hsM9iw0
QuQtQPg5o9jcoKBIMk1l3bmrSWvsVDLACQCPZvbfFTU/jMFoyzqCoTBUta8Qamr7Y5urDj481kZr
DQRZ8v0qu+8ldZAWr5Hy1Q9WeObtbpRCUR/+jxy0waQzOWxgyqMiKS/c02f4KWyM2Jx7qFFbORdq
RiErP6Ass2uSfDx0GZ5baKgoGoQEZA9ZCrgXH+kwP+Bel2rbOEeQjfpZRJkcn/SUIMcUylz1Dvf7
0IrGJ4lXYUqcR21rCV+tCWg+xsIhyDlEFWlbRrXT5TUKWG+YXTJX2uHhuYG12BQ1dp3TazQ8UlRK
P078CUwWyonn509fax1FxUeuQanZ2oGDzPUhHDBlmf982Tp9poB9Q/J4dcsHNda/4bN0yrluz9vB
fKoOMmw+07Z8xIPqQPsVMTccjdylS7zF/hKRctyGHXjutXecXbBH6mQEDH89PVllEUTaCBWfniOa
0wRBX0p74wyWgd1I7srjbnLb/0xw+YXLIq515rSZtxg+me/vsfiz1wAJHZCOq0BxAnhpevnRhXju
nvve6DEP3LEopxzxVXvEjHPN7i/ejkythZr633+H4y2BhWEnfHak4XvyReh3jJVq1/98si3LQeQz
u5Iat/sRcEXAvAHlDOf1gpeB5Xcm/GhDNB0V9LGElBwKWytnmpOCrirT6ka0BSOmWz5Rne0DTxgB
jmTB4s/8UkTTzpSInnQ4eyozrprEtJJQHRDWZFGrJTxwthqn00+1DsN4JRHBzd4k/KLcG/bafoke
GmGlxO/+fKONWwUG6+vpcBxkEiX+qfBhlzvRvrzfjaCTHUH3R7ME/AvJvqsQEaejwgImP4q2xD3r
qE18+nEL5jKHUVm9jD2kkedMVfIKwIvhQc2d1QX9h4DEPSHDY46NIvN0lp5fWakKS19ddFUdEHVc
J8guDL4GD6orHoAvDFxrUTqnPea+uKHrFm+ojmQHQWD6uGzwehdsZ7bcfAgKECb+yRAL4YyAuqGx
x9eXOjrD9A3/KfosncJq0XrbX1Pd1aebfZwOnROJQesPx7xzOhc0Y/IAMtw6nAstswVGmvjRW9Ad
jtKwFX3+GIbnnKwW7Rihqj8DKDtXZzanLxYvf6fRPB1072bAchh2sl6PIMx3YeCzElcc5jvqwSBX
opoc0dJ25O/nb4owqX+faF9ZAEkWkE1fKYihcfEfHb+gA4bpf6Fgw8YBVyCxAkSa4yud5r8ba7wF
23shNolpNIVJ/4A0TyExiJ/QlIJTiSid/Iq9OpQPD+94Y026md3OpcnxN8Fd+gtDt/NCFAJKPpIj
DWNegt2gHN+xKBpEgwa0kCGWa0H50ZpV4ZZcGoV7c1u62NOP0fhPp9Yie2x4TG2C2h2zo4D1uNIF
4XkCrI5mQzDE/g1mAr6nhdzoaMHQKW0UCPOs3hYe3p48mjJsLYWxUi1R1BQUfTFpdSjTMtUrFzec
8iuuzbNw5M/pcih5B4mhgRTdcDyE+AUzYezBJ1RW74Dmu4IbG7cMuBKVmm+h+do7gPM3Z2L4rATr
HYsnCZOWEZ/cXLYsqvH2TkxjeHonx3yJU7wYBiZhCeGuUeIuArVZ+aNq5yR43i0QApDCO2uzxVhd
zJhigU2ezh0IIXeRkmW0J/VcyK4QPw3ptdIwgK463aTUz0vghrk7OU5xr+M2Q13ZmvGZ4d952XHb
T7DQyB6jgtdRUvB5NHZpfpJjnmoxDfH1AVknYNlm0eOUWJDR4LhN925X0us6LUD7SM+LzOJS66FP
S870ABkmU+tlRE06APuDcTEvqBeO0y6y8+1ZBvzggCuWHFUPHz7KukEEb2HqjTPFyAiVAOJRSjAW
55WsE59nWDOkaewGcNnrUXK6EEEoWQm8xnMfkAuhOtOFBGL+T9PQxxnj+rrrcrFkLfkYhRMJlu6b
SmUv3WrQDxC+sgCyjfcAIqlZIEt+/iexKGGilkhGG32jiyQ7En12tDbqHGKPJO8PcClHTPX6+/bU
+arGlm6aZvKCuScVfZTWIUrASSvn3i43IYgobYHDnSTPTHeCgWtY7/1gDJkrNkV895reC4RQBIWi
inpJNmEVQdvxDwYQgrsBlOdjYCa7hLuzV3IKXBbjzJcY7vsElaAe+ry4ClizunkDnb9HQ6lXoUXc
XoDrsPW+knvW6jW1vwU1yqvjClx1GxjslbxZ+WAmZWnGElCtbvEsXzztyzZgwDPc6V6TISXca6oA
Bq+ZVPFbID54CcwGiCvrQjR708iFUCzdhHDTCIXbyx0p4l9kPNaZGPGSjDYCWxoW7bxma33urhjs
S31Ds04PSU77mfbXw1CmkHmCmaUR/71SMl/oOM8ODIIO3cDtcr0LJfGzVEkpSaInbQKwZOEAgqEw
ct05/4zK8oITGqv/1yhm97btASE7vbrTJ+hyE0Q6gmOOVJ+n7QS9oE6nPphYefUmh3f6gMPdbylU
Uilq1UY5iuHC717SF88/kreZ4rfSSnLqf73z/S1vjqB15Afn4MjxH0F32VhU+r4KtyASAKaucca7
SYT9hrcHW49QmU9PFJiBeUm7pgvjae2qs/281BR7P4Ib85NqbKDNHMRP08djS8t1nBJSY8aQ4U76
q6A1w4SHyzCH2/tIrTIy3q9nHzP6603jseLA6ta+SqVfzoUdg1OhsHWUnDP72vj3x7q9k35aKU/V
hf3/BRVio1VZCtvD0tapJnnBxK+LLqSiG67vblAj0Wh/YquuceGZj0jNzoN/mITMZyI5GYys+4tX
FvlCkCLkVMshrMwwTWdloQtdTRy/QUqFIG5rdzTloXcO2MugtG/wLkI5J1I4Haa3I80aORxmiaUN
pBe2h7yXoozIaROYAbxySS1Paae9u7oEIMHPd/4CJwlP1iPfpu4FevONjfqz9Fn8UDvTdzjHF8Y0
YQZeyT2dtQhfgr8wjbkzmqe/mVot8ZuKLVrT3QbavBxB46F4+LwOCD94JpM5fw55LRVm6YAtGnSR
rkxDEwD4QSEiseCv40pQwSAShXKnuybhb8HazaEu6TTPN8tBj63csNUVPisyag4Zm4nACribH8o5
LBzJH5quRWzu3j23Ak4P1ymjuMgsX7KLjbTc3xLoVqoZZfJrU9yPtN4T5nBPLGWla53XA+P5QhuU
paQJi+Qve9oDhoPY1QjylPJpzJO293XX4UPY2GCpsRk9RhQ634BN0UsenDrlHK6e0MMfBBb4LR6v
NBFC+iLWnqhHE8/eyHoXmqKrKzzbCPZ3/3VQ/Kv9o8k8tsdK4NXAdRIA9E0iVYQdojkpeRXnj108
yJs9yJ2LIq+9Lj/QSr1VSmVh3i+8KLis25nrhAE0bfQ0hvkBP0O+6VPGdsk2JlTksnX5ZrxEfppT
pyKnN2KsvU7+kmuoJd1/jy2VADPAg/wCYrjUDBtqa1gDfckATxU/ftHkXmNC/23wvqvtIEZhohKj
pMvKegORBaZLGcx+qc11oNxs7TMaN9xiSSyqL6ZpDlw6vTys1H0cMJC6b4trKjsUumiwNsFR80nS
p3Naf7OXCzJvdOSgvfwTcnuyxvF4T0xUm31im3KqXftoOeOfShFiIfRUuMq4uW4aP8MAEKz2ThFu
yynXFq2HbR3WJ+fjWu/zf6K2LO7fs5t7T066Xee+OWwW8G68kBSbfMBSgXkd0NTUhiXXon+HF0G8
rWJAr6pvi0Il2QoKo4zYfC3q6I2iMiMWbh6snfYQgn7jhKOYDrlPq2ndFCIIrq5VM7g1GYfnBqy3
KUlVub/i1KO5y8D1a+nlnKeB+DsrQkacqmRs0TLZrH9BeSidCF+XUG8jBBNF9SuM1vz5Y3CLjALB
PZ+cH456gep7tu4Un7RtvzyKH1IlRXhG7BB9v2b1Yr4Jb0lXXcQfiiwPRdNKhJg945WVyFFDCXY0
37h8s90YtamVZ5WyL9dhuodB9UgOuJVD2fz30dZgqI2gga2in5d7x4iQQWA8emsHJuER/piw93nb
Ae544eGnEk27SR+2UtcaqEeDmfHIlHPsEtNo4V19TIfJ1aqKqvr9BiWNm4jCX9AQzyFb7jRUb9g1
KpTsC2a1Wf92knoBkA8q2OWDdIvqhgYXqjNlx+Zkr9VrAKybI6XWE8IUgjPkDcBjcVKUsbYlY54c
XkNK3wll3Pxr5toAfhzieHS81S8gs5U8C0sBJCylSKX8YkBw8IFQwvRcHC4ceiqs5uPMQcTESswP
1oqZ12BOZ/sswDoU1ticC+2K1Dyxbqvg08rPmTvieW5R5/jDp54KsUBHNENGE85LoWuTKgSpqEOn
xZ0hx94lpvZgoGcqhBckYDaGkDgtaYVWzPUXSdVxAQQq8YnVT72tJnLOakFar3dwVWEP0J8eoYTU
QNuEZpOhKV/kzjhO5tZz9Pn9ps30MPjpagHPur3yVrldPDPokljFOKLgHbml49RHWCGwDlm/BjK5
/WqhgU25eSuhscA4/sRD3FYmNBQ/xj+oVJIQo7K/pAPYuj7+8yhzdYy6sSm/PqrOeo0LkzQuEHPx
97yFD6EBrD84MupdxLCAe44UxbMVyJ1arlR+7d5M45sYkcZ5d00dsMPYl4w1qCJgMUGbuQubk+UC
u0xOyncEYvaeD5dqKVAATIwBTNAqkvnAfHMsfOJxRcKSFqT02Mhqc4Qs4r/t3U9LQW/ORAu0xfLN
hW/28eGlfK50PbuvNCmx/7mPgdpCDDdmLfLAa7q9a7HOqwGuFWDADBOufr6TrlYlPXijDWgPME67
FudW0cuQXR8eDoCbTUKpodvEoY65CWclEyZQ6ErOr3Kx4eGOkE2gOaZ7psCt9rZ/zGiEs6PhLSF2
ojzYE4aziJ7k8H5x3h8NJY2iw0+SgN+KgOLoLcMhOcIKnGqE0Bb2QO6XQE+S+ENLxBBjaeIOXA9/
H7Zmo6aylnCQehSh22STWThikZ8JouDVPUJ4zLXCGsnNdTdeScutZ718s35lIdGe02FMYpZeER62
+7S8x7QlcMj7/fXfJlwTSlY/j8lluInN7t6rJcBJkPYtnjMl16rSOearJQ/RJ1KAy1O+/A/xFBW1
XY4zTDSUdx70ncn2NUMYRW1zNxxChBcLeddz8GGCz+b9JqbIy1Nrt+55HHLCK8dtsamEMLySyqV/
NtFtbZPRXwrXTtrKJNHToDuxm2xjxKbkC//oJE5u1O/nPT1qZIcpDplhYHZZl8DVZd8TW1OshUl5
aetxeB1fG5UQfKkuj52+xOOUwFz9cDcebJ7+yvyE0u+7p7LFtGWgO0B44VP15p5S5flSEGWvn5Sf
SYTA8VhOcpBoRkyrb5h0HU1lgkGn9K4bbNMs+WZjnAV/t4o5n7eBhE7U95SRmbAPiT4NyYfevjWu
aJxtqQWjEcH0jE1Zp7cKZgcLhkuoTQpCe+X2+AjTRxToCBgs5jU9mNbRX+7/aCKxNoxAlgLxs2LM
BWM3bPTlhOiZ6hLzX6EzknHnMFYy9+tOXQYt9zmc4lHRcgH32Qb8LRNqSbBcZWAVjzs0kN21kOmw
HSS9o8qI4zwC4pnxNqAd+8jCHyBA6mqeCk57dlGUf0b0mrgXWeOiwl6MXNIbOlBsofBcDXa/Rjvg
dIGJBr1EGb7XlX5Gb5G/aR1I14vehyfe+ufhJa9Be+tSBxw3nFSVOFFu6xkldPoUzw8/6Afv/Y4a
RD30zhkjnX3yPvfqxxICKPCt7AP9pFZ09acZ68nRDBtxKDypT8c8TXJaqEMl48EeSU8ESMXB+QQN
uyFXsF2sSHuLZrrEo9vvPPAgJmBMWaZ+gPYEpmSN9eQQIy2bJ7wlkIMcUcf7cl/2OhSqAp/AgLcp
b+ajcZbzlwv6+izPOcMEYwagPqn2ulRfp/xMqxwEKtFqazlbbuUKc1PoDN/uqDQfVB2Fx/HXaJOo
FPi4qC8o/8tsQKeqIU7ZLvdz5RkrCeToyAcAQceydMxG5CwvobDuAncQfuI7uK+NgfS5xwXZxlS9
JEVrGo3E6AR1lYqNN1tPNqyvlLn49ubOH0hmwKv0vClE1azoJkWRdEJSFdypvXGOW95zcnmUNnQx
a/XSwQvRdANVM3y0MJ2xYmP1y4p9nShxQkXQPLoxlZNK6iQHVjGsGRmV5Wh7x298YpSIN4Gtiq33
B+J62j5vw7OrQ8axAviNL5EJ1leTW9l0NV00wb9/EojyRZrm+EkuLI8BA4Rpr7Y66i4dZljUhQ70
Y03B237WcAyCdlnJ89obnN9lwuvlh4zqsbj1O6kJXZERozQqM5eYwIMkF6AE4kV435rX0IlG2GF3
sUneY6e2UvNYn4d7fY9WnydRcmPzlJKGr4Nxd4911wq9q2h3FqhkGFflHVKXdJEonPaKJAyZV+cH
+nbMtPAIqTpt1HG8VIqY1J7PDWh9UVOJh4iby20qf8skySugoK+Zw0BvHuQSOh6Z1pORJjnrB3IX
nHFMQCxOG4frWeMP6jsbJocpcgXSPZV/pQR6p4g+UcyHHC9/sJ8MbA4MRFju5rrW4vGR51DALz6A
aPPk4wrTFIHiLf4yxvT3k3Gz2XEsG+yuqylwrdRByiqG8LU5b4zdbzIbFSL8bq1qQW23buXHuQP1
cl7gp0nJ5BKBBkgp9KTK06+pIx5ZwogaV+89FMLfHcTEOe86oscZ4owh8wIJWUeaEgvbKn3DrqF2
eWSzoFuNuUj8Dl/Inrz7/asCIYXVqy5Mi/6VMkYbTC1HODCFfRXFhdW9S5sqTq6X0te+n7ycOAyc
t5wCWK//L822LEf5Ov46sOKk5zvxELBmimWFyZjlI4fdFbLT4ovGq1UGUtL70hP69ZRNcxRGEdno
mtqfKebg99LiJ7bE8cYHHdIVebIZrWQgbzBDSXh3nzfaKwOJy/rhlsuHg6+ZS+2KGmcxr3tQk7au
DIugUsCrFeHMq2yUxC4JSwRWo5sWuM7HVH8mKUtUglOc5zr1jqzUrPwY24RQtBzlXA3BM6Dgplje
AizuCHEqVIfLfco67H/YtNNLb7yvJhZD3TovXxKpr1IKUHKmyn2ClaBVSnce4yAWWhOV2/s7kToB
o4a4Oh2CseEh19+mhy1aQ3+wASkd02YLCANOhxpfmNe6pttJ/ZxDftxybZZeTDKgQijOmC5Zf3sy
dj6ScVJRKm8UedEBcaFkwqFLo3h4KdlB78XjCqSrc7dDQv/SHmn1HLSponWuTFU4jHe3IodyDMk9
YmbYrNNwzpqEE4TsEpnDTERX8Uw+WIptOUpGu/n4Hf1MFnow9kormRW8id5BaPMPFsKWcC8x0OqK
Ky7loZYDGIfCBeC/2bkQdJZlUv2WMs2/hf82qTAKsiBpd00+mYw6lYa8dzcTt0YyWa1BBc3MX37X
t2ca+uwgmfQZaJ8NS5P5No9tCUe6Bt72zLwUkB9XCxtwFJUg4sGUL8v3DytJXL0BN2mh2LIi2+49
9/0qjhahU9gah4nJmLlIM6o8USForXMxPxcb3J/Ik3SaFXakPLbs81X7Bi0pPVcX1AXhk4detmHF
Gru7UFROFdhOdE06ygt38xGM35g1QaVupF0I2lf7EHEq+DTYDOSa+OSwoXIyC80L0D3grgSCvnEm
gDC/3ytdTBdaYz1kDjggnvekTZlUxaVrRVd25zfPkTJID+f8/H7j7YZn51tSNw07trUdb0i8FhEd
xBLebFmkmyt9pT+k0+oG9xTSb1rr3HZQEEr+d3aILoOEPgI6MIjVac7CtKveaJvZENs7btgczuvZ
JcLyAFCnl5iEPIBxPMpeyfT80+ptkR+DpD1M8geEieKaExybTDWKxDJdxU3PKbYREmHCuyUQeH6L
2aopUvmdh5LrGsL1DSkYHEjDTBTUVy0R2kKp8H+zVtFzawFp41TkllZ+h+NxB/pTMT6OVZxXYniw
R6KmLZ1Dy+hQ7Qwnh8z5ph3NbwDxkcOtrdwSnqy+tKoJWdR2PVsRiFyY4IRrSX7vlLDdMP2zo0en
HSj93VOmmwAizUZoRftOSte22IYnwOPHEXnd8lOFsS3xLYnBKTWspnr1/iTB0kfWPN3TznB0ntsX
Je/B0JPE8qNEb19cp2NCIul7Tc5HL1AHB6yQQ1wBfXATiFTGyhcGTcLdI+AZneW8QtPqQPkIhyxg
TzGxUw7GAL/KlMPAt5dnu71vkl8jiyTjePEr4Ub+Ilr659LQKUv6hq4vjE4Tse2LoJXho/b/S5/u
GnSa8YmyyppZIZ8SdofijzoRf3UpVcJDzBd8WwldyHv8QQPwM/twcUm7+WuA5Y179qq0kbc0MQgv
W8bOjbtFfaGqvcEZwDma0/oqxzFvryV0iuiB61il79TtW5XECnkzPYyhhEf04SlbEuKXRwAxi/7t
3bhaVJoNqODYItX8PFCqmCcoV9UKYtEQ88J5y93LQOYhgVv85mqCkzIIFiDxf0BeVe4vSvi8tugu
YUvA7oJQXfSH1E0BmwVBVsLCUl9A4KlzJFzbO8u7Pj1PyNexzHm9qF4sXDFsHs6qz7mwHsp9IL5S
rQ5H3rdpZezVGtuF+pGaHGu4l7tq5An/bjDI9j5YSVCoaEWTC74E1+FEYFyECED4PThX1qVBcBg0
+Y4+7jGsu1rzgQ5UypGX3OIjdtSteopzgN2Fu75tcLcjaQRp5XBR8FPPXmumU0Ar+Q4f8Q8wwN4E
LriYrV2c0tQS7Y8V8DWuCznSIxOFJnvnxlkAXhT1NGmxeF9uQ1Buf/ie4DlIVy7c7K3YOWtStHl1
yBYdd1JNCu3zF1v9vcDxGHT/rqVIdJK+dNZrB04egro+QNbJkWLa4MewStUSZU0/viZi/1v7Axkt
3mD/oEpjVSZzf9GRBZVvYrUAd4515ZeFW4FcjOBbsIXjwVdddPDh+5XBrcDIDbty1WRrM/BPuJeW
L6jd/GE9FZLhyil+OZUqS8Z/KDAnxBqWSKuAu83LxnTMvVt/CQWxz32tu8gpCv5XRoj1vtsNri/F
RmR7f8Oop8l68ZrYguTnEaObnEch9nQf1h4/AWYdv/QMzZ3hvcXNaAc9ss2f0Tpw5OfAxBSDU1Ia
yOTZykARDmVxUw0Uz/l0spRIuI7DTPjDtYIoEpK9f2yjwB1cbZkyw1y2+eEpRy0y+geu2TMaMtYV
Q5H53Qmo8DTXdC5XYydx3dvgvkZ4zhp4DeaCPgjaQ8q7Iz+wUlTWUNi+7ZPKTCO3VijX6Dwozrbl
51h/QmES7RZm5JpUfVyxuwP4/zFs1NDZGlpFNfODzs/tF51ThmkYUNhPMtKqxlJ8+SAiUH9yqUl3
wQVh15XNwcQ7Wn8HG9e6M1TmDyWxkFvJrfenUSszbvvL3U+p/hdaa7f/WTHElrgVL1ddKKKJyUhd
/wI7rJzCDEsbGg37lmJ/SzXCupwZRL1qXtOaCQloNrTy3GxY31ofISwGchy5X9Sy3+zaDd8+yZFf
H992xkqxWQ+Z/2dscC/Y9pC7e66ZPbxNR3B2kxf8IZ2xR/zRMJcA/KGG5OqMaPBiix5rX8yQo8gJ
twIk2bElG+nA8nXcpr2a+nDC8Tfu89ciDKQ9365vhcdcgXPJHo9lQaIOT7y2TEuKymb38T3sY3li
98ZnoxmA8+8NBDk9SlQGGG03jqPLavTa4CUOxGGZHEAXZBKL86C/LDLsJObBPYg8XmlYyshyeHpc
pdcwFZbD9pj+sTlfol5TQXWUbarIP6QwASJxc6Eyv5YWZgGkjjC1RIBQHNqpGNW7ezeP//RR2/RN
h/rBUPPcxqY7XyP+uy+OjnTfXzuBiFKsTr8hEAlnAowUR2eHLRq+hH/VJQ0lapLQy0g/47jXC512
Bjeoi7kIcAJMmqPKhRToTPUfERYgRpWBUuMvKKe9TXVbS9RXv7Sg/xohEnmUbdgdrVP9yjjetG5E
p2RceEd4aQJESvq5e3dZiOnMJA2fXM64KKOkdzLhP88xhkFfEGI0WHP7BmMEq4ZFL8psUt9ZUesC
SbpXqTnezSnI+Lsdfr+L5Ip7Fq4FHUCJbYn088HX8Mjf/Yc46/n43q8R76IMCuD1C1D3A3PBiZ9F
9M39vLHcSihzdCeKvAR5Z8SHjSKychdqRpk0faKsbzCx66tEiEwuZ70yY1tNahCx1udg4sCwvjBq
DTK1+0Y9NIu0FDPYkzpsh1518m9/RZluvxV4kN2a4KjQ3uLn7oujnbWb3rYpil0iNoW1+E3p2PqU
ekQQRbNlVkPdLcSlkh44/7vS3yGH7HuT7kukM+oKTiSNgVoQ5L9a1KpDBiGPIekoLOB+bHSTh5dm
wtbOEL0Y+BxrCgrL3oxzQei6IfZ/EON5/2Sa+Gww/D47kw9V19gQu3fgFlRW+P0w8tZFiq51jj39
PWQOPwx1JQGtL+wjUY93pbJnhtcgzfvYvZwNpvJNBAHi9SRKfr+91QObYMbH19QDLpLAerHuaYzD
+CFvVo5iI7Ttnh525wm49Ygl5dfTVia7p0hjeTXXTOqZvtONEhq3cUSGcGotaPWaO2k7lC7CoalV
hq3ZlynSaJiwnPRprXZoG57EKkVUhYR8o9WiXRb7zpq4NA0IRhtoa03drbBnvbfLZvMhQU6THfVJ
5QpnTkuKRtQbMSr4ks8luvcxFnbLQIXJmC97FQj/VlQ9e0e4FIc1OqoUFzj3JrWh7OxqAoYTchMS
vveUGynnRhQKel0o4rY1l0OyP6e43xZlT+9nBrqNDo1ICGQXXadzLrdVHUuLqJjfZxeiiywIiuSz
GAPf5xBqUT+5lJMQ8TNFNgLTWc+LoRaZgJAQ3zqLxfZTll8Kg35rmIeIbDMidQvitXos4boJrwxh
GgfFakO7ut19YlF6fjd2jN9v1MAEOwaTwADZ1q1IsB1aYUNJmOjEM9XyIfxD7pUIuuBzOmn9Gqh0
SENYobJJuoHNS9dn0z0a4ETUgdP65QtcPaXWZ+DrjlyBvQ0sW4t6eSvSlrcAGPtWsjXzjxP1c+PH
8jrexhAKvl8b6Uz4bWCD8zO77JGRNGXKCHo124fhiOi/c+LZtLSJ+G4+IBjHJUK5SQJsHKPh2Awm
zQ/BPW5o8Htn5gL4MFoqmQIQZ2GnEQac7JXWguKQCBHfDDZen3X/05RHHZvP8ndeTmDADFl+qm9c
VhdaXsKAtXEFKNZqoGBLyMXXsVYHyycrdJDnmVklIlteSEF6rnYbLzZ9V26oxPtuc7HKK66OkdM8
kXwQeXsJbTz56R1snCaz6v+LMMH67AX/t1Vi0rezAUn/WtCC03cl+l0nRz6eiLIc8rsQzpxyeYhO
nSEaJ8FrtzA8CJLk0wcvsGBeZxdzcv6K1Ubjc+vmLxWoOVbBDaS+il7ZSDV/HzsJRRJi6WK+XJbh
G/hG8it7aqJAYbCx4CVBodbmsgFZW6g/N9qMb26U+thZA+/pJNPiWtHc9407JLSYBYodjWopNBZg
H26tLN8a1r3rzdwnhmhP5SdlS2m7lNwkVv0u+tkd5zjAmcLTYzXgpVMHCLuPZy6LIsqwi0J7+NPo
HTOWqwWdLBK9DKwru6EYGOMKxUKm+zI0tNLvDGw/VWUSDR1sn6Vj1Lm5cH7yhBi2M+8OlJXgAjyB
wQzzCRgdbXN7ZuiXba1H25TA19Mq04vsVt5VQktSAd3pGVgeyJ/2FwcaepOBLYILDJEEHmHexNup
SD05cD6/eyip/Ek3TUEkaBujZSo+2+J2/SCUc8DKyw4chQ7GsPjm0zZ2NzFkRRjj8lWGL/fQ3hkJ
Hpa1Z9GEQtjb4csTKICHiasaPXgrUIbf2DoIe2mHp+WhgX7eRA0VEoU8ZacHZjyxm/J8JhKBNtAR
7waUGTHnDbngJ7kF4J8r89WtviItX8IdeDw4EXfd43FYrkas/jFScHGRKZE++yFJWsXiCkmhjD99
Cy2eAWO9mKV71y55RIL6dLWUxHUpLzKvg1dSPGJbLwJOBEudf4/gTYhxQwiTXhvXgWabqCqWmDhU
b1IPURu9Armv+VNb7Ovf7xQx+xMxR5KW9H2CVS3kn2lqtC8CntEBPLYxE8RLaJjIavwPxeFBUtId
hbHeVMxI/acb23naz37IbBGpuEfTHcNBc5LbpgWA5cOXJUJa3AvH8g/U9hGKuYoPmhxUx7fekfRW
6LVe7slmSldCCTAaOacXSo7RrfkXKRSTHmNPO8wvWAmQh07jViVqN0mWh1XrenOMj5XYN4BgVoyk
lxcSUkPktDCXHMabtQvPI00HA5sdVUyL/WSgi+0bB+3Omc0UVYPu2Wy6KRMYB9c14GcCLqLu/cum
S0M0vbmwO70nj1NhJ/XQQE5huUZnFpuvnmMnrLsAsRyWoPlF2RLA2Z0YUH9rHPL8AQje9Pi2fnUJ
8g38T7PXeHWY/Lklsi4r9OMJqxGBFCIqdi4iXYDmSKRdhIcb/kqtbgY+tSKDn9x86V+Q+sjPvD/Q
ahobxukOBlGO1i0y2Z6R7rdHOhbeMb/XWn769hBOHbWebQB+Yd+r99O2kD8T37NMjG/+kd3ye46s
XKw8SJwspQLFcsj0R5yt5/iO8b/xsjGfxW0LFxmQt0ZzXake3IWFhTFlQARtS/NN+37tw+eV2Vx+
tsPVqj4sil7PCNfxdXvoOKnandO0vHBXcSS/gwKA+wrgoVDc19gqrhUdaY9xmzhxEp1zUWz6Jaij
AH3+4WJs9fYGXFwLz6c3Fu7D72zuXVgNzYo6H1w30s+w3JJRP746cjVbDG9s+cuhNOFL/IE37/WN
13ND7TYg3V4dQLT153DcgYAe/3IW8Aeaw4UpCARofaLERLDCG6mdxUHXpMajl6dclob/7PC0+Vjj
T/t8JQVGvGGnlGTt1/j/B9Ch/ulWTZ3MRlPQrBLix9r946hB4UtshqhuwGmsdTGp+xHA3cGRn8KN
+EtuzgZOxEkBuUdXI3dPkGSGpWtmr3uMZYxvFi7RSfFrQ5b0kHD3+ArlG/maBh2RqFkTXjCrRwcU
/Pjn+K/9DR38IDVF05+lHwperxh8xtL8Fd2hHGZsaaB1SR+Sb535pYLvsmhNiJmT+R7qI01itIJA
cYqy3nvaG/RtarUKHTQVzeFZnHBVwdoM6zXdiNYH2ak8EW87Xikj/GYrMhTPurqdGooav+Uck0Aa
1j7yGDjxHB+y9r7qxtJCc6cugX9LZs3e60BVwhzd86cEq6I/14GCGJ4mvU9GABkcRr+rYH90tozt
lZYlcmLUXorOnLCZwrcHfvsTc/e+131zow5D3mq4/ioDpylv4LDF7Y6WJNLckYIMuNtiqFOLrDoG
9a9uaBITupMETa6kOJTGtHeCKGlikxsDBOL0y/EiXpNKpXiviawg5X00nXLaj/JBqy7qwwb2Sq1b
w8iaDRTAUDY75gQKyj1R9FWPRqh/EWqPirrtkpRavQgZs0etDvdirtuZaoYeyjorQECCLab/FKNm
ft/OHgIP1dWH8iQOks6fcWZJy+R77JsyHoQCaa53gwp7/45hCZlb9uM+J8sjQRbSb6vQ//h3ZAvD
apgGaLvljmU1fqPUUPDYqPQnT04sFeA7+ZbYSJ1CZBK4y/wAFUuBQ+AhD/cTzpSlgUpYp0rQSRWS
1fb8z9bS8JUqXxUomDvSRP3lgkaKCTYKb9eLN3KpMux0J2lCsv5QE7h2yJ4HFeSAL6yEgjnq2rKv
UfGCnRTguoh224sYyGw6pkKnICV+Hl7f+b2REmi85dCaWM0/vGiKxcNGYKiDCN9Um+dyP9Q3BsOT
2PUEJLzccohbmEaGLn/PShOX0WyMctMxnl9Y9IjYuX+UZMDoRWNFkuRGaY0t27O9ee7f3XYGMQZu
9Rau6IoMZUpYmCYwr9HzzKFNeE8kSUOfafeUre68coXFwAE/HNlfJ8THbcMU3a70CwOghBHlWLGS
rQppnfoxgKbLxOdz+bpGMwQkt8nvNX3xmagC2g5H8nBMZgaSrHQ31RBqPM4Wb9M6Liz400ow1LHt
Mkx1c1n5j3XRI5hIMrhTevSY9hCSP5cpUULIkE9mFD0joraA4Q1PLR1NKqmfBdcSn243TBr+KS8M
7dvGNjd0xkLBLdUAMP/dptcF1JLtj+H+XmdkNu4h/7XTp3eVLfMpDHwr9V2CSi/CJC9Tkdszn1X9
H82FVQg8JSd+VFGWMW3L0oyZ3hHFaBPMu15ylxNV5CZGQ8AdCR3fgc+rwbnUaz6XI16zGnB5T2eP
+mHPLckk9f0dYrtovt/j8zE4PMCvi2nbkIP4oGX3YwxGJHhm+wyNkxI1LPZ24JzlhF9DuhJ/Bo+u
5doNqBjtbxCaxukt5yj9NFATzk87P6OtFxdmnwWWFnwNr9xhLFgSGw+MExPlUSAM5gVPmdKNIAzk
XgYfhNYEbZDi0gtn3TDjKkVO2yK3CaOat8d0/LEtUjKdv7/yB16s1JcKNZgfHr+oIXyz42swclcy
poofybnpkGLXXAc2dgIQZoGWqmpTSyDz84oEoPX2aQu68ihk4VkJ+RQvQ2VKWTECXWKWAyst/oRa
S646mbTPbZSucZ5wzZrnNJ0QTkPYHL6fw1qwRrpEC8mJE3J12kYp6bWSG45w3CotWHTeAihQx50m
8ssUvgRB3Yd9NEcjhMmNZUoHPmswluRNBI3OkackvwZSzkUKjJGoNEyzxt2sDSjF29aFOWmGtUwM
M4g3+lsIlEugYJzYxgY9Bd2iCOvUynbv0QVZgIdf07LZfx4x0SuvYYC6l39RKzVsRWH5YDDglt9p
5BJCttBKZ0ifP/AAvDaipFvRXcDDpRDemmk5e3+++E9Q2ms8HDnCk2bLBBNJoMwnv49KpA0wsyfY
GdVfjaqs0iPk+gkP2/4/d0Jza8gZ+XZcmX3Pq23wO3rQPxhjjm1lFrxYCciu+VbM3wuBfHI6SxiA
YTvXhtblRqZVeBScuRRrAebDCAt9wSJou4EFbyA92r3+SHmJWpm1CDpftLZTREYWIHtwUQFL3t8h
nzU+yLFEAx2PNSb5T9Bwq2xuJjumAGjelQSmiSSj9yLxcmc6x0advmOCO92wiIMCzo1MSA2aiLxX
1Nct4WF3FoHsHX54x7dZhEva/eBVIyRILgJY+DLQMBYQnrtiPPLYUfRcj8tSJIUonFeF1GXCmKNE
tc3P4xGWp/AYL+XEayFiNgHIlwfT3Gdi2V1EYdPiporNM7znCB0tRbEIHIu3bc4fDh0ls2oHETru
w1R5lctPrvcjC4pG6/Vw2du8x1qMXOg3t239RKkeC2uIjGYCVmHJn1kkjj4s1qP4X7OTM3uW7Nqb
TNy/k8RrWcLCh+3iMGE6U5Kihbgb1835rG7XXgV6y0mKx5v5Yu9Kxf775qN4KF9NFUYw8yUq/whv
BPjT+npL/aMjxDhQK6UE2dqiy5chmBc2n9FYB3aBDs1yxFssNlneEgjoYn0VoDlSZk8fOIDQwWnF
Y9oM224n7BxI2f5hJ7Oz9sVL6lTCSl2XU+qThXOuDCZemaO2BWfHRpBz/gw91PAgnC/uUtc2oRRg
/M9AZDBubOqzgw5/ARDiVje2GP/YDLJNFklDo+KhsI7e3VGiOSHQRGSYbb/XO/5x2gb6SZG7UgZ/
yDshCoD9LVOGc41Y3pOCJ/0TXHBgLDMBFcJM7yKMXc3PXTZzPoZiDZPmwysQPn/zozZJR4UKBG43
c24y+oByv69vC+SBsDTcsyyE6YvL7/qNOqGIju+1B3mCKs7LwBtNfoCB1eQQkQjoOUkFGBsSPM4p
tqRb1IVPV7QpJI5R6NxNTaUfwL/kcMZptR1W7ksNX1xmQDvToPt9jMi6lXq0h6dMCR9HLxDahTK0
q5gqwOWHVWJaO74pR6w/OIAjQWY9phGb2Z1/iqBkOMa32C6+g29eWejXSAUmoQy4KCO/aouWn2NB
p/GC/uCGRUfL75YTFvDbuy1Xboozwkanuv1pzoTVEV/MNc7ljF2IHItoYyFAJ2dfwBpLUovm6NGG
ZVSr8Z/rABxBlp49yr58kVsBpoNIbgV4rcc8/C5tYguloM9bOyhHMXQrEfAc4JzrR4YdkFXIkMNG
bYxiNHgBezy8cj2TOC/gb8oHdeo+dYbEQKlui0uv0IIxCsv8y2ArrlW5J9/MajXho/mciNWTEY1d
h+yHHaeGNKAtWQz/iGkHPRIuAembnZPT56sbQMbWOWl//+GyNpCeU3TTyr0ejvt/A5qCr43GZzhf
hW9AAdGnSQsM01N0wrcprTOOt1zWjeDt5KtCXk+V0tpds86UJ9WRrOd3ozimUw1Z3lzo2ImheWFb
aJgk/aHXEv0IrxPYGAyLvdDnCB5wiFH8wh/4qfNmbZR9FeRMrW/T0ld8KNPVCSs4NTCq+2pODNs3
7v9QxS9ZnSD8+FbUFmfIzNrTLtNOBENkRLDyPrgGdIusgiVSEX9Mxv8eLZFTVZlgqqtHmHJV22zM
/cXHF1DyMv33Oovkvnb8Z4H9Y8IzjbYaIK3gq78XBvtsqa/PkoNng0mrLQ4VoLacJe1aebqhvZzJ
egA6UvQbeuwNj5VYFFAwszeVY5wkYAoYS2TWi4B5rcu3VyY1kKNJg6ubc61bns0lAyJuRfPOiK9o
wTHCMSylxke5p+liJ91dM2UURKS5xDdA/jLNCQXy8f25NoWpYCk/3C/wQ2e2W5bF5ZpuLy9sfA0z
ao1FOqZwbRqNuDIYuU64ncEuKwyzMuO5xsYe3rVlwWqzanHCloh9A2XdF6/ZwxWUlJhMyUTpH0pL
OEcwRmDzYcCeacLI5veE5YgGdEXhplhdLCkknW+2Ykwl0axyVkEToNAXofaq2/MbL99xEi4AzUX9
4rZustWALfYeZuLLFOaFwcIntU7MknA3JLmKtaPsv5xioJowKWN0E2OohAd5W/cEHnM0MYWoHze+
KGycje/3G1H90B7ay88C914nIKnZ6hr5Jg4fEsQeuaIUOwqpi+NGDunEIFKacX4FccO3in9aTvM5
SQ2HM5KLr61owEoPvZmKcHBRpiQyYGBWMNc7kv+QePhxqi02pE/fcM9Z9lzANURgKVRealnr3yp0
P+gZ9e+gQO18PVOqFexIsdphg+ZGVqAdYXJICV5oCrB5YzWI5OFsBp2GxWiIr4SkGl7hNIdlO9ov
DS6Auzemg93BNzGbHGaQLHzxDhOYVxUkEvgeu2VVmajIABinuaf7L5TBRZIAWkQygUxMZOhOxKIl
Yt8EW7hS8uPwUGj5WH3Ow+B/Bb9WCYJ/j8EbOlEVR2qSXM65S/8m8qZTUoz4eGIFxADdwSbrDEpm
q/JwlQ5t+GljU/EbzlnPGhbbsgqtAP1WY1FTE1Ot88x6UrBray3WsrWeEK+sKQXVeyfpvqi25ce7
3oOo5s1ZTTMvbeFZxi6Bupp6caAN/kMqVE0IxNNuqsqUhBxwDWShaM5vFug0d/ozjwjvT4Kr8cii
jcrAgaXUXkRyahaJEhG8jQRVWQdTfS1rnUEk9GGNbPIhkNtalRsyTLbUN0aTzgcTrt+GntQCIIwD
cWAkYVH095UU4Luh28QKRt5/4d64ruzx5rj11d0HYTbOZXLYILUtqnhg37p4DCqj0JhZorpzZAmw
pxAXFuMeCmCKIJTCpYD7HISLBIZR9+FhXmOiSPhVMV35smT8jt1EBD4ppZihC6YQUeWI52t/FT8I
9cc9eVAETWTHRzq3+hpNGciJc0KMcmukTkUWWSDn5foGvBDQHS1IqXVcazq0mzdOMLBw4Fuq4sqz
8MsX+q8HyKYe42AT2XXeRZWdJG3/90h076vaZPlOe07U2jyAg/D+UIfFCcxSVWBrscwE3BTCyyqS
0YBqjHd0rkSaAxvl0d5giHadvA6hDyW+maIkhFsPoa4XVky93YQeVI/tCPyAd4bw1pQXabdQua/g
zpXv8Dy5ibDNiM4BNxid07dc04YDEF7nJcMW5yjCUv8dEowRlMRbt1qO451JN/fWIs6v1d4GhSSf
1O1ACxMXsGEOaQvx0MVjAMRVlBlp1eoj+33okkgcTDOTU1KEkGVVFUC1ge+RlHlakofVIHE35iNS
BbBiCy2WrOOMMiut11fkwxXRFPTJFR+qkN42SfRa2r+guJo97R8NGWzGkSDncy7E3y/TpB7xljNj
inTxpFfchjQM2FOV5zpvNOYpXRxaLwWUH0LjlIGsFky7wxWUID/KGE1U4Tpfs50nTzAQNBqnvjNX
MoenioNZDENNPqn1QBXbidj4eNuP/V0SaycWwhCQYvpP9w7MkBfqeuEZFY4gMrK1FIdTOLTkwL4Q
qRLdbA50y6GMp6H1zoBD4wID537ZNzD4BYOSpVnBnBN0j5pymoI/Cbs6jFHpm2BL5ssPuQ4PswgM
rR49kj+8xfRvoY3bQK8Inu9XImN5739NpcS7bCz/Phsk6j0Y2d2D+aDbBCKGqBlSju/zcbdFn9kn
EvK8Y96Hw7jwRHbH5vpgAoT/Jh6C4jPi7bvAyYkO0QMesVT0X7nHGcHTTMKFpCJY14vPsgLhspP0
XlXt7/DJvzBxDnPB9bbLQeiw6HgFDOhhy4uzg/hqMYvjyF7bE0Nk6FI+XYrbxlc+bY8prFbnjnzL
7FZNQc2WNJ65CNagnpl/Sz++v/u98Km18oQN7gmR/+SDsN0nIn0WsXKttAjXpK+NG6HiLTn7mkl6
7uFGCl23KgUP8wLu5wu7ck2VYjWpUM9oww74YX8vyiHM3zwX2Keo/fcaExAAQhSPIbct9mJ6R0uh
7FtgYGmcGpA3iFcVRjAqyAAvTuwhhetxU/VTbQJfoTPhsAPlPpXc6e+I6rE7CDaGW6XIRKzFTx+f
y4wFL9LO9GpYNvO8CEbxAXXUlxFtC+fi4D6+sOevIBht2o4yaRF/2H/0B69zylamQyyPOZaTa3M0
4z5lT3WpRlDUFY3GKSC4TGTszQRI6Q8BLNDeNcBOuSI5azaxos8FafjB+skvdPGQKzU9QlWAXln0
rlDphd+c0COEBovm/9nKEMYoEAEtsb4nNRQVbYJprdgi6Br4w6yJu25+29yXYfsPlAERU5rudSpM
U06zr7husYUj13j1ahPirgj/dWmneKHi3bGtyGpdTfGiByo88jjb1XH7zjeHzYgdvbQvyf9+PsLm
qtc14mbcuTGoCLiqtS8slolKWgTZfoblcb4zxJ7pq144q6ZhxOINID1mvyw3/vgwUz+ix1OPoZy0
P6JeO0o0/O2ZU9R6/N8e+kzm9DK3yZIOrKiiMJzVeO4+WdAGXfE4vX5lmb7gP7vsVMADJRv4guT+
/5a0TZ/SIM5aKCN4Q+pVH4XJgNoyv9MBnC/vdSBeCERvNhF05yo5ebtlpz78twCZZXUM/Zb+R/Xc
N1EeSI2LM4DhVp/26PkSAz8U7aOQovn3YhqS694w47PHAsz8R6l8H1EtGp3YTz8SnY5FlwxCB98S
ixe3agjQF3UQo52VJ5YtoNjRU390HtrbOCBq3QP1glCH+46cgw8eyPh0rQ2zRXUG9NxZ4RujmJNx
bS8C2NFYKD5FTdA2BM1REyVhJj3H0ZHuQa9xq2ZLOXj903VPyevx+oTCd20YzZKAFPsVENKh8NNy
ep8BeiiHEOsFL1GjnTCg/TBesBpIVJthf9xX4BQNsOXGvTeQarKKLmGvzVDR0LI2U9Z0u3e6TqP/
egCHqD1d48MGB1tDeruC6VPx/2JeDyOOKRI5z+HcXlq4B32SUnThsMeOf9L9a1/8cPcwhWGIdSu5
Cq9MyA3pOBv0Lb0MP/VNJyrSoaH2VE4i2RxDuPIiI8VMkEKgQpg9ogXGL/sbIFPxkOGrroc1OPtY
52Ei79PB3DlThhD8z/SWgq8NsodjmDhMao1fHRajnhdwtoAJQZu1I/ArplE1Vq82te7+fZdmjsJt
nKom1DDNJtLb/QwTBqk9x8H4DiLOYbTmBnp9R1DELiKTGDxXOzvYSRHFGVPuxA8/5fxRkEBQrFpT
EcVhOGo+mYWUApY7OxI1r8fooHV5tHlHGbQMAUK4eNQWqeqJ0Kjicd5wvuNS38B8jMpvlh1NCgVq
0N3LasAp2hEB6hbiySRx86QsnYpjG8tjxWQbLfe9BAZ7/9mA5nuIti4olFdJvWpDquTr4X9RGM99
oEbssYLG9wUqct1HkXYS0k30R3Xeovf5qe7+IYyHzqv3QxjwTuoyZCfgdK03UJ2MMAZSHWuVbWpa
96aYWwFIho2eBGGw3hC4qeGm6eHcUA77gMBBfyL5YcpjAWZLYd+J4/1odPFWIfqpZ+TgIzjiNHEN
Q2hUNPhnCmTSxBznwbgrCoi0Htf3zEKqfNjPze1G8Etuy5KI9eypbwI5i3K738BiyF39QTQOaUis
ASs6Mq8qE/9AzpM+OkMROA2/HFK6WJ2n/GR8uoLb/UsPlhS3l22OLRec4loWCrp2IdLk+xdMTonG
FfFv9mG5+hR98Zwgz2GTa19n7QQNPjD+N7hKGKuTBQcBDABXAUNV7fcuZBQGkmn7F6nRKjhuwmx3
y2clAiu70OJJRDFDt79l972m5ZQdDBx8OaYgjCD81VktUd/gPsPDUzKGQRlC/5k5wvQN+wg137Xb
LxCozXLYjhajO4noJFrtYt046PVBaclcd0wHBqNwOTxlQEvderrZEuWahOwFLqSFtDIGleIQmiSz
kbhHCwkwxAjqn3+Z3vhFzCJDHZxF+Su9jsWXCNl0lMgv3mk36SpPa9XOJMSMeMP/M2Pacb6Qu82u
zzg7CFDxUdXrQ7PD+m/IbVMrvHATakTLJkE2z22PSPEBeKdAOse+aswQ5LwAGujywT2IQbpT3AVC
xG8J3p63S7R8BB0WRj6BuuE9wZWkUdjQqQKyvWN37RRQT0R/Q/cOnGmJgJIg5EHdzoEilF0ULrEL
DKOGFMWGdRDJ68Lro4gtgYU4UiIbuursauVFgYexvWUe6SuFZBSd/REdzekYTLZWOPXIUHpjHaPW
oV69f0OWjBmHmgpyYY3TOmtDPXUDTHqePBW0l95oWMr8fww1qI0jOkMbi02OTEjHHGEFeAHCP9fT
B+X2jRXNhakPvsJ88C4MYNXPb5cxbsXu0Jy7kGP2S5G57IUUnPhGOUkWpLELN+fYz4P4Fe4FZnSZ
5fMTIo2/JbcW9tHAbUOtN0Wn0oUK66vfRBeYn0Qy2vxk/GrdfpHG8z2RxKiqkIS1sigyfoapqDL/
M4YPMXp04q5O+Fi/kl0urhI4CxtVQXURiYwXA0dysqe+q7YolMJdkRZ2NrRdT7S9kDbgALXeqkbt
ZeZ/1u2xayS7BhUfSKq+JTUuYfOF4jG7L4UoTnVixpzBPz+G3Etz+pWblR1sAVL5trUyG7luLv4s
VecG+ajqzPDbpYz+RTM9Qg26PxNxdbLL/gPwdAZt6pT3FZsrqhd9hQ0HiX595S2H6L7hc/O4hN8m
D/W4DYJiGUnXhbLg+atn5KobzRpSwzpDo/XOWuBT1T4G8TlLi+xYRjQ57rKXQ8EO2TRfpRqLVfbR
Z7s33+hZhjJsKxUypDEsH9HnKZ5gbMfWdlGYEj4mkC6B8NKirm+cvvuCvb7DQrVqj9/CUBbr5hsp
eZhiV/Y4FC/LlZkTAEiLBt1RCXEzVU8XzMhifQZzhCanbnYRBMONPgVbzt8i3MglrpyXCQARlPVP
2o1XN9L1gp+dSmTkm2ifRj+Ytqi7fsBlsh7qyjOSBzvNkmDXf0d7NUPVZjRGRHt9pig/Wk2ifOCh
ufs444fW6RbkNbNCbHvY4R/lg0G0+EdF0jd49cTZtx7LKuRjmfEgQfz9SlMfNQpU6w3Pmv5jASoM
4bLIsbnhsr8RenDkbEn3urqS4EwkosL5zO2/93+BjLm0dE+HGDV8qyZGGeH3mjtlsKiUcFKMB3KB
Lc3uFp1xbV1UT/U8oVwCQQHhpO/RPU9paMbw/ad1jtKDiokcScL74fIXeqHKrdTl7urlLDYiJroA
CigO7ReScWGQquDUgBvcbC3vujUrvRg8ixeBoAGhekf0eq0KUfkPKty6Ie4bjVtcXD9esXy33Jvu
8eLgDxMJlvyARWgdk85itlF8G8kWQKi5IbaV0fLje7v7kdh3Xfz39QzrUl95oJPyxv+Dg/w7i/BA
yRr3RI8SF5wSL4lF3/77YyOqIrYm0w2Z0LEV1MgIjplEH5vcwAqDWs4uC3kn8vr69J5A/N64shyj
zyZz5zyPbYp09cLTid8DfKWz4GQvTgxUNoQ92EIwTuquxzSeAA+iKHfR0hvs/liVbytcIQQYz4cS
fnOqgdgF5Yxp2LSzWjPzPcq1haA9HxJ0p4oQEMewjaBEAYqvMsO4FFBuLZaI+ygFvCh/gZ6dTHhg
bj6gmF09IpJYh1616oOFpNrxim669LldxxN3ezPQhk9C8/iV5pUlmJMluECqC6U+SrMnq3cDphna
CXwHMXud6ZMcCzAImZSg+9P2QlKZsqTKDWWoaI30T+4DeACfbvh0GoBrhWoLKhWWLmj6v5XRCSEH
oK3kL5ob64Tn0tOFMH45frIX3nDldR/iCbTcy1Um/KXUWMkK06FpFW2D4bBgkA6XyQ7abZGu6PfI
qe4xuphhbrAMlFld8AkJP7JPEN9TAVsJuUNcazVgFLZHWpphoMUmMnAcPJw3z08GRUOwMei9Mmpl
JNoRSBsjNmIThTcky7dFIQ0ZbQMSZZ55jKgxFUewGsPS0Q/8Fycg5JNUjWYDK3uVy3voQz5tqt6Q
DjmAvtcsOS2uNzLQHaBaG6C9niwc+onOAGA4P5aqg19rV2xPFHUIzBQWmMWtQN+e4tYuJiZzZTyn
io3RTci3bg9r/a4j4Vj4If9vjoRKuq1rmV3RcoSnPIwypqVeIh/syGZN3+muDYem5N6Vqb6JSm+F
3RaqWVTX4LrCy0s6RxMPO1C8/LUXmIbX72y7ANfWyXMReEWvAUDyNqyhrweCneoxWv/7uYK6Y1Op
JMMAJjQkoDL3LW2oJppwYLbiEiyrWnzl7rP6ltGKoA249nxipbHVRntVkmc5lxeOZ5J/MJdhc/VL
FDegOR31R33cYaEPmGU5G5IwcXCGXp/FBcJnv0IbiF4xQhw+UThS9nDklZo2R254YOG+IQXkAJnO
cHquJrPUx314Rz7RugYmE7iWwGHyTZ1DW12oMx6vYqn0RumubpcgCC0dlizRT5XluGlKHWMEymja
6bMx325VvqddRrB1HJD6qCeiirzbFzw/z9Q/sF12m5a6wN+clO46tBBtca3PjOPKBodaJZd819k+
Is4dKB7jBPDY8VuAmhlw9emxVgPJFvlKzMEcNvcBz0F+rSfdV4SIvduCo7jLlIzhkR/IsVWo4QBY
IwXKM9Y1bKz4q9apgBIC6Kt3zLT0aw6QSAQnzRhhN8e0iuM3scoNt2Q0209aQkKjnDkDwqK4pqty
M2IqC6uHsFZRToMlYabrwcsO5bfU9B/qWokwWZfxL88ywbGWPMUhkJvsd7mzt1sw6fAOpuJI2UP8
HQEkfUzzvmMo1A1aOxvWg5GXSkDmLbpERDXpZNkC7fCjmXkTsZxHKm1qucAxWzRJY/8akF9yLSSM
aum85qx1kgY/CQuE9imR/1JId+pX50Kj+tCBmR4/S0lfm0K/gyJ7t3yLG/Oa++vBBqwKYlZH9FZQ
CC9vKLdCDQ8NJ5vH96oBGCr1bLviE/DIx8qquZ46JcMkotwrWZY99b82vQOLc5/YT2lNi+M8sxT4
713oxdb8+sDcNiWxS9wZSIIeqcNK7VvN1DZSL5MJnR9+ayZ6SyTLYn6HU+ljn5DrVAjAxuowpNVm
Was0Hl0+6gU+Py7ZduQ02EHk1NwPmWqb8kRFCTc9MSacs2Dm/mRmzy/s7TkmYK0icU29XwK+X4+F
+efOP8nenDc8vaJU8RcCqd9e0R0NCRb/LAvXSu0cxUMNtxXNaJtJp6+yfQ3KPSsaU/uJBgZlRVsJ
IDBNg4Ip0NYq/T9L5/vvMPsbrOhg2NBnpGHOnxaFFJ14Mbgd6iOjn438/t6qHipis303vg2IslpQ
GQZE9KNLjUOHCLpI9Bbqo9AqeW5m3WjoUGYUbLJ6qtsKNH8TjoRzGzsyhY22WQOvBF2BRFv6rNif
mWiyyXUElNiCTARq7OjoUukkyjbXaPyyACRRGD3BTZDV4Z2/lWbUYgDN1pDQAf1ZKMsNDdTsA9op
dr+0YmtYuO+neGFCSTE2vjEU2muOaFoOc7qIsHvL8+QjBGtftf7I4GcE6mhdyfY4stDpvP4yJ6Jx
TIWH/r+L1/DJtukCVT3f9vpIj607PEK1iLLia7xFtIdl9c+fmfdsTONPwyt2ArcmxDjOtiBECRxn
Ot3qbVDxSsdXpMjGbLkepITAta1nMdzlipR2evoVSo9FeuKAe/c/s1W8ugdR92z6oBWF9TfoJJ31
D5BR9VLFW0+Swfa0WzZatjCBz9ocq+mKhFB9mgdfwza3+0gBO3eMZMptHuJQD7zpeaNsyguFM8xR
YhaGaxe2xIVsXY4B8o0kOka3RFnSjHsINVHBORNCcJ+cvsDS47OBs9utl94VtL0JzvgKMhT/aAuj
wm5h71tKYA1+LomdnY8TOScESpqM23oGUffjWtXsiDtJWoMdlZjNba7HHEaUWmc2Ikw/N9l6GXY3
8I7VwycTuy7ng5A1viD5GhiILcxKaCut8TXxmxPCmrscJY/nkZMWtmSgvs3nMUEnwgF7EQ+6ALqY
/3isWnKz5m0AJypEJher2sEEYNyLtvbXdPFiFkegnOMcgX0lM9cBPQMpt44+MQIALfgqdr7WaLNI
sidka8lahMeQkFwxdIP9LfKu2Bo8iJu9c3quIQ0fscYdfbj79FwpqFLjGDtC4y+2sEWusBRO5VGY
lqlWcQPzzeOKYayweB1kXV38IjvYFgEbdjA8shfTO2mvtvbR/auelxdJ/UnNzzJ9TbwyfACjL8ra
0XLxUNKKpBI6MC8IfJvGr/kbOpWcnBLh8NZH2pGzFcavLgebDV51i/qFRToA48EtYyoLjyogLacW
eT7pniWPv+qVhvYug37klBakOR0JeI5m2YGPM+aEfHn0vRYXm7dxtSa8iCF7Cw5umlTIc//UOGoH
8Ei3pdJFMuj86s55e0ybhupw8Tmrf0Ps+JmRv5Gn/rGUqdoPg03Tver+goC8r6RLMo/YJYYq/ouB
kiWV0hg4gxTBuuKr+Ps/jjyueqgT/0dPHwfEPlEq5d938M1bRHYHZaYdFVBVDds6TNv4tF//Cifr
AF+aClmsfadZ9iHxg6DgJZrt6Kz8mbRj1Amb9HYkUYwdSJC5+NMHUjQELwhkjvLkBG+5TQa3GjO2
l7X8uNVxeQJ5z5PiJgJF5nygxPvOnyyERJzSonqS6UoGW5OjSMvz3kVDVDphr3CPCdBnSjYCbYpt
KUexmiFKzWenObw/HiFm9bc3OlHV7GZMd1F/wH6JlbjkyTMbaEjgeRIIAcsEK1HViy5ncL3eolLD
/dfKn2B6UnW/PZLkXuYZSF2iuFChtexUod5zYO5DGzVrkklZSHeahWw9Sp3RxSvUeSpncldQQwmx
NL8lH3qQwn2xi4N/lWQommg5ZS1mQqDKmXy5W3UIjwmEY1p7luY8p6vHaVTmKlbawNnChQO/v6Yc
BI8E61w2p0LrlTVcwTScPcnqnb5E4VTmMYqha7qubseJmZ/0JXD4FA9qLCcBp319is3uWRbLsJgO
C7VcwA3aFLbx7sxAi9aRLYCYguzvr5whDQ5+fx15Yj5vKkmKk3mTl9VJMMk3WCulqlmZCx9v21iS
saA2jt54NUJiZfftIYLFH4nrAWpFUJB+kduvjBj8OHjEIZtK72vh1Me3DpRlUhrnQMCpCBen6yq/
wsscDEwXX2B4CxXmA7kfOx9/XxrlGZ9lRqAz3bcE7T4/TWwxrXWGYckLavasjLc7M26wL9ZDLqic
djYOiFQNq9Z9oUiHwWX6B/3m8Gjg8fJ7C3v3t59I1uRWaPTJKxczsEKZn8M05JghRntfDXXT+Hmr
kmWzPtznIxzDC/i/FGHca6zSxek6204DLVMHU+MBD8SyivRFBqj/FYArzamFnUkHtUxEhsAJ8Rma
zqBDwTvKnvWZGoQKr6jLfIpmzeTeKfNSmP6syhJ4vi0V/4dlvidzZy6BYgVZD4P3nO0EowMQiXS5
ZueAbcf/6Im12MY7K1/7SAOmx1lDHUBBTEFVPXo+E1ood0yUrxhvc49cSimYWy2uoCwQNoW+8uF2
2s0vGCt8a15Mxt4ofsvfzmVfUfy4R2DULWkxGsiFYmKB+hIWXipRYxEqajVQ4pjPUk2ufsPsFvNp
9dq9jZNpiRPhUYOMMZ5vvhkSdqWK2l1Nj+w2NIJoZuu90xdrLXRWp/b9boX6DXgRLCCFTK5BMXwj
RLvE5sQrBKMn2mSXqs82ZOkQbkZF15trzTs0pQrkY1TwJNUZXiJ5TfRxdwxI+LEZPftoSzmAGNVe
z9UxbSE21nHuUvZN9c9sUrvI1CandmRi5IUyuobeT63X5exRuQhcP+SfSGKbQRgKlAWW501MYBzk
pnUWbVbBzcoezQsfggXBPwlQWD+NUpCP187gyLEtub0IX4hpFr7gx1R5BzTxcKOAzm6rvtf+dk2w
ErfJIi9Hj/cNwTUWKNcoTKRzuHRA8glWs2AEPKIfqAGviEQmp/zVKcLmbC6hvETIeLFH65O6P0mS
phH8R7a1y+k0mJYnUaZamCX3LlDge/gwzZ9EX1ry57XV7Pbis/V6aFVK53g6mLVAJKSyR2ewSjA6
997GVqFGGzi2NRw1IGHiUhWh2tEEnSMj1j+8mGBEOmBVMQr6G2f/90NGb3/l1YTX14Dqlv7WMA4q
w+zmMU5+UmcfpREq/UJIMA/7Svy/my8WvPx5peLTGvSh4KfKhShtDxhZyd9x8SoYwaEijrsr+SRl
rszBWewvMu5sNUZ6vdyMiEqNlRIt6KrIRf4bFql8Egj491BPe12bn9bzSDSPTaHzG2N0qTfaJqas
Ud799ObM/QhkbDeyzAxf1xQC70MO8xIKIwGivqjehQe3tB8zplYn9djTA6y65ZSezlOhDtbOfxtR
cp9XzYFgQt5a29+lYtT6M3ZbmKGQBTxcPCFy+z3PTzzRYhklVQ9kyezMCB2UrVqkSLnpclFfT6tK
w6yXSPhl79QzqrpkSXrnOf+ElBLED1fKDsIUQDMJ+Lm1iDSkj/xAfBIfr3A0vFc/Y+06oNHY6agB
6cmMiZO+8/p11dzv2y60DR/cJvUDkSXE4at4V1n4arGUQ4o5+CTF8p5HPkaB8uEMGEzFTqP4R9xJ
GOOxiM5O2ROkG6DQh3UjCmsVgdq46jBqvDYuHC0b0I+2e56ZxyE0XuiaRoZ9/m0ubtGxiyhh1CGN
BYEAfPJ9YBoisD1F0XMJvANRM0WK8GNEzZaooPIuXPWilkju9CyIwBIlxGCR3OuKJiMcgHvM2Eo9
1WgUJpzBfCwzuN8feJjWzlJfZbz8+29yAtVdRnSMw7FRpXDrm1IBWkRySu3V6roXNpB89S2ANbk2
9ZBZFt5BYsPnSXqPN8EjIfonhc8G/1P762Jw+yZaOlYBp55GH5y3Dar0MsNS3XiTnNNXH9BXJNk3
cRDnAj2rkTLGY13QyOdTuKUuYZUy05o9PAaJ0/b0W/+fNjaj27ZPszCgW8A9t/xo6adBrD7oBisf
ETYr0g2zfVrkMZS//vI65hgCfd2I+UFdx4rPehF5Z/OVh915rf9yOZj4W7pq8Yiod2SAOTDVsRei
5BzElR/wBhyy/Vt4BiRymJrTCPh/iv/fkdnUDR/Kun6FO/OA7KW4SzQ0C9Ahgk+eLF8mIC0YTC+a
E8jn5SrESJq7EG7TzcJb5YyYbblvs+ehK9vwxuTG+E/haGhWr8m38XSFUmSjeWSWtresgKGVPKrS
vfbXodvXnzajK+vmi0iEN8JHCDFz/1uCwcxvrA2+xAp6obAJDntjaJD1xQ+9bwyJSA0kYru0Yifv
Jvx+h9sNIbGRxjqzjlJeHwAiOHHZlwWCJUcK/2bR0blyhNo/Vo9I7LfC/ktU34NVtpKutIm5C3cJ
tbE87kIdx7VGbmbEUhltYCEO6L0y0ZIFEhAW6oNuozw2fzVVZTa42yvCVfKp82oIYB3V2ExPTOZF
paN5jql1dk9KfwlsXS+aCxF7U0G8s33ci4jDn3jCVizQ0xDdJ0zD2qXGWp6fyhQW/IbAOUQDLwRA
zIamIrx2zGKyrP20MUFGgtT94gfRUVHfezgoxqGZwk0dFXEYINRBRo9tCWFWHpREZbTEKRDrk/+Y
Nk+rZmhBoyJEdJLtytrdO1f9D5BoQNoScthGhY5YNQBWmG7pOX2isgW0+SpQmWPi5DJFHNcz3sPL
YqNNSxAOyVx17sJ49upHertJWYT0DtstC1gKuyG/vvLmCoA3PZRTMPdCvUzQv4hT1DdmlYUNAEgy
06TPCZjuKlqTJmENwecfQVdV9UF8e6eRNswLkpCBQeXUXEWYimr7/e0xfONX+lOfTn+DMipH+gUG
+Z5rVrKEYgS9k0nv2Gi8UE2RuKGuqDQG5AItC7QjfCpniw/49nK27RatwdGggM9891IhnpfeZLgu
cLZ3YZw79vocqKeK96szhPGCl/EqHNfkfBMQY6CcVBiBvtOljIjEpzuL+ojoW84RVbAanr5cR2QF
VoJoW9L0WVpDgWnBjgwDn0HEcsFjIx9YqXfdzg2BEbY7n6zl81yoQI5LHVGzQUQ1F79vjz+omDZs
DEtl30gE9zACYvhl2AlxLXsKbHIOAIn9VKd5bIMiXFjfQkAO8uDZTU2QZwqmkaPNedK3gNCNn6Tu
Ei3asLKN1LBvokQnq/jJu0Tx3sFTZFweB9RAswzUWGb3EtaXSF1a3vWnFPXsjeyce7GFseRlY7Rp
+8udg3e/D49DEYGvOI3OGkj315KNZZpuurTcyx1lfKjZVqguUINxX+wsHEDi/tE3BLtVmAdqjSIu
snA/9yNWwlNV+/R1NFHyJeQ25dKnQo/VxhRnT1j7z4Yb399SEjdcewdMwF4cdpmw1hTYzLHLpslM
f/oAsdtrBqFvfCB5lF5zLTvKGVZrbmIi+Gzs83rvLKjFMEijx8GkmoasT+ezh7CigoxS4+vKOXKK
4Ig543Jzx9yzKejisi59yWGL9hz1jIvH0YazIuSvpONYZDzuEfJZmxueEwdHu17rzZFT7rz9hKiN
JigE8Og6MyxYU+ZusCyFPFnfaHM51sP4O9qXFd/fOIFD/GlLS5WRPX17QzjOl/cHlJTR63CDXp3r
3cio1QfKYYyl03vKe6OKgTlnwPpcAyNtup2REInpfOrSk0viVXGQb0tGsL4xG4H9qbNJIC4u3BJO
g43KVNL82lyZowwuEN8qw8Zt2yDw+DJyxJMYKMcJXCPXXO5WKZlUEc8/Wc3gU1rqjlPu066KmAv3
mI42mQ8POjIY0mXqEfj/zHNkZ7J5k+JcUFQvsfWZJjUmAtfhtw921R/s+JMGLMXkGpV3Kpm4Bo51
xk4XnK+ZZN4XE8YnCxqqaZn4/wjoJ57g+gWNcECuj7QxRPnGSgUH7S3iSs19NYtsm6kMUI8k5TE3
sLlfR419D/vSHfIYhjjacIxRCtmXpaAXKSY6+f9V/djenLnfUNABaltOO6CoZuINmvEsxkQKqyc7
N+70MfmC8S7OQeV7WOjLE9oQL/LoL7gw9vnJePiIU6MAAfJu29YgzuDNiocYhGf+abj2NDZ7Rdo5
PmEtHOkoCbqFqX1BnhFhLg7zdhSujWKnSCep7TrcW7fADeE+H1cbBKMDvM+m90Hf8k31FAWrAFKw
dIEgHNgJ1bNyKCq2AS0ojnt4HL+Fg5xUHEIAEkRfO2ap3sgvocrYSiXf4CzLdh0bQl75ZYsynpiu
q99uBo1RWSRZzx/N8Bsq+GXu3MQzNhe8EAB6VTOZTfYx6L6SQlLvxYlIyHrB5OqGr9DZDN+/aQgn
PRO+Nu8dZVpIlvmjBEMgQVb/PPCtywKiQ9NbipIryVCORcneMdccjID+bf939xDJiWevzTcE5JGE
vK5TVNTqwTCkQrWtXAiRnSwwOOUkOr+XXXRnP7YsaeAFS+PhrwFWMPohlyqQc+vvwL2K2cLrsULW
S49aYrHf1O1SpOWFCJfzcqiZAkxnTY7P9bSB6f3CZg2MP6GrOt+vCGGIFvYopJFegRSUVtahUlTE
nudh5zKIf9YzEbVnO5CtE0x0fCsRAIy/FYmUtCG3T1oIBGJvkBGnwKBuplKfOJZDNcbn69HTlL6O
99KDkj1HcNVHhLoUN7UPuSJx6tTYSIoLhRau4wqYTzWjV4kAzsAA30asZW3YUOY2h7DFBuD9nwIQ
BcI2qMREOCfWFKzYwlsSyen6F6LYGnnKI7I0r4o3AlnzrStMS/6v+zTF5reoTDscuXu2hLrpGBL/
Goo0ahCEmbYEoER6NIktdEZw6r6ytDvlxDkueievBrzZFlC9bHKHQDoItYrfENo7f5YWVpC/nJrU
vZFJz1y2OhSUVrVpJGUSylBAsEcAJf8lNAv42QUF1aw8U27VruG87NldmTOOWbecgqtmAE2xun9V
ey9GlhNGRWnLo1ry+VrHKCyFY5gu7e0kUwkdV8yXZcQWP/8Mvn7X82ZDNmsp2NxzAimKOWgNkKCI
60nX8qFvuMw5g6T35wUYvwsTyF2DcuAojUw5tg6qgXhUTmnb4UjZklleRnyrvBFdAKlrgq86DN0d
aQkTtTfD+Uwb3/Am6AAYNLrs22+LrBkeyge7IzRSUHNx+oNDQChWQan6B1EdyyAKIyXnGhqyw+uY
r6DQp9lAUROpTV+3ewBJ2Qkou3bJ3ztiaavBTcVjH4HltAMnw0kGdNWmL5vAWEY4xiWIhllr7P7I
lJB2gE65OJmruIQjPxv8qkOFRfuYBf3KZLPVHOleRW/zjUU3fmgs33XYJ6gRm1gExvBh4PyesQ3Z
JgKYTv5trRrz3apgzvaGVSzV7kNrGcce2l9qKoS7wAzNMsk4Mfrfsk8TcT0ER0CINsODIocr03ch
DcKQupQ2ZxpuzXnHzpb2fuqFp7HyhYjDmNMmVkjXeirEwUNDE/wuTifDRJXgP8wHBPSxcbEDwzJG
ClKCT3NgoqRHS3DnxoqNJttDdGc6JkyjTfM+iSXIDLrr6J96PDMJUvGmRepl3erATfjhITXVaCD3
QGppt47U3kx2+fEMwZjwYlGfmp+3nOgywf7ew14mRLCTlu+4CYc0ChIcxptA32ygDTSwoFiWbz1X
VLlQt7WxoQpqYcrqJGqRQI0r1vo9d/Ugbua4OJPGd+m6CRuTCDYrW7ydowhFYVG7BU8vM6Jk8xUk
9GHk6n0N60O/yNqG2Z10D1BlyisRG8l4aWTIy8Ocva/2oA3d3b08IEL+Ld3tdfhi/HWTqY+sAptC
mABw3y/l9gK8PBB/42V2kXyPA5QPaytRalHH9PpBq21L69X9r18nn5vliYUY5QtwcT93NhCzJwRx
r8Q/SZpEAbb+4u+I5jAcxVpFayHa+ZtmS9VCYVbANPUwpg4RK2RHImYO5Yhz7sbKz3ykJ1ND7kuh
ej158M1av+SjFJmKhs/UjU4voa7Nb1jW4QY6qeFa4VPpytJvCsHTqpxnJGZu5bw+gat9uNHNOMHJ
OWMU5VDXBuHmuK2gsvVEaarxkLeC7CaXdeG2PAIXeS7IMAVKmOyuR6ch7I4lxLTJNozXO7QdB13A
XirL+lVKUgA5+/Bxxa4wIqB1cZxgxDI1MuhrL+7YKdZfu1LJ22s694A7mdDGpbnT0v6Am7G5XQws
y7NNfupvOBBSJHkSslcuac0gK9s4P1ufvNfx4kx9UAfu8BkzDVqm+dmRUi6HI/eSUeFEDFDyodeo
XbFQq9oZabDbuCgGVfQxQ4F9Tyn+K37BsN5CIDmMrWyWZlncsvq6pETlGq8sQ0VTR2JN4Kz2eKF5
vvtFaroDn5tH/n7cEsBeshFGp6QwhYAZpSQsdBjTaqcfhGL2049FWLe7TRhbG36dnnxDyYOf935F
SNrwZqsAT1eRvB1sdhIV/vYc+6cKuh0grGuMrKOUrRRbUv9DF3bsK2E6GnnpwtKAB8wrPXDgF/AH
/QMhbqDrnfeUjUcgnlVuyW0yjwVAu4RZHRI/DGSem0R83SYB4I8y7YCQYnsw2heEvi6HNmRW4H/Y
WBO8oJ3z1AZoqmpsNzGtzqzQt8XCN72gmeSg+WoOUD0pWU9DbVoun9ZNIQb6iyVGjfvfufxhQy4U
2hnuyp2S+aZOa3uS9SZqgvrSTLbOzY3r1PyOvnbFHg1yIA1szdFQwDqvmC1S5x6FvHF4QrbuqG+o
uD9Q3Wg7kb085IwaEcjon2OaK4bumIbzwtF/kMxsJGZPw1l8t0ViLh2aHQXy6kBp4/PtZ6Gw2Dj9
B7myFwfQaA2NPI+XtdhiGUxW3rRuar/IEVA1fHJ0w1VhO6xAoWbGxILzm1hE2Uuz1ZWHHSLtB/8N
HCDpyF/5h/8L44bkiBPNx6oIhL3xsPI3KuoRjC+hr/T05EPEa9XGPYh1Bp+xFQQ2RP8dHAMtn2sn
dHFLZgVla/z0uHFCCC0Zs6Qx53AhZAhYQDHqwNdaxWz7BbJlIcKdqLFK5l4YPybpEwz7DBDYYQPf
Nl36Is0p34I6jaqwIn+uoKVO4TqmIUIPGjpVIZgS1F3Hd81yGSLp63sKKLCRd+v8B5nCh1ouayXm
ItaAbenQ3uoG8WS28s6p6yGeHqDsLN3Gg4jaGscJszvVxbu8T7JpPWgwLEa1pQxMlfOfD0JnbyFu
qpuiwCt6z2+4JF/QfP7Fdte4yJzEgKWv9HTnu/FtB0bQcumYF4BZ1JgLySTkr6rsfhwsxZCKBn8e
78Z8OmaJsT+oxoOADKOpMTDPaTpsccyNOCnaGtHN35Rk+OupYbkFAn/RDRzgaB7Zo2nqLsJmbVfD
+JALejzGX+kquuV6ULmyt5rJgoQCbr1Fgckb4deEu8ElrLsxKiqoNBr2IaadfNpWCV44dKof4ZEJ
wwxWE74UV686buhvf1PLnUQkDBcPe2DKO2ThLb55nhycSxGE30O+YgibIVGzxjM8hsSmdQQz5GNr
2aHLGwuBa+pqy0sB/BHsj2Zzvs0I4tZ58xng0Ng1JwtP/mpeDhCCBtQUrlO+qfdBVzAGzLipvhtF
0C5iTuL+Kj+uMX3GVpnVyp5lWnXBp9N2UiEMafVg8CQX1xQ2AvWNiUEBOje4/j5suatwOHn5apKC
svv6AEAQKTlIYWS0aRKpDuCQ6Ogf9Wg7zaR/uA8TWUP4kGD25NWnItrd1vYjqSbnC2u06zHqhtYJ
MrcRQtoljLhdNXREV9lnTmI=
`pragma protect end_protected

// 
