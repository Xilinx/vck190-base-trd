/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa", key_block
WnUYD0g6/qDSYmWHmuZSsLHluSdi9+myTeKuKMxZY1YiclF8fPuiqftouQOib18cBMrk+rhxXYqY
YxxEMkXifSggXUrW22+E+kt/etsSl4zJseXz6n9xUwZYg3xlqNjifu0w0ji98CtnXurauen1JNyx
O3YJAh7IDwn6xZR3LTGYOPxMj1rA3ndIEld9FoiPlSfzRSRuhh7ozr80Ea1y9ZyRdn6UvlSGNFWa
K+qWQ9v0fQI5P76f/h7qmdvfXu9BKunBkypsT5BoGjV+yipSZpdDPJFuKi8ZALQ4AfQwwQQ4W9Ow
ic2MhxBJty6sWw08okzuCC7DdaVW8+sh3E0SQA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="GeeiI2S+0qmTuse/FWjb6tqEZItAqGIcIYeurwykgk8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1168)
`pragma protect data_block
1KvCHb5eogwPJFXkT9BICzMxzNH+vrV26b5lOwPoY9M0sYVnE2KsmsRg210SBURV0M30hwtf7pfj
XyWOmX35FQ9DwsUPUplUUfy5Cluw8mrrx8eZ6mmYz/XAP9UJVt9w3LO2fy3etx8tFEJq8wqqnzt+
nO/bBjvdzZDFyqVJvEulnR/1VWZmGkXijJmgekS488ZWlLAZLfcwoNZDprBViIASOO0UmdLCZVY+
mJq5QtvSKAa8lBszx/3827n3LVeWw05RpzQPKJQKC29FZB6jkij0I3g4Hkmd5SAapVbVbt3P9aTK
4x71BlL8QXWZQqR5vnHUx1Pa3RE971hcin2m+d1PcOQwxrUA75Sz/8Jy5V75olxQb/VZ941umwMG
PS/QqjynhuUfnvmTBh83pPwYMt2i2e+G7jfYgQcJFN4N8JyAb7+LQPwK+frpK5ST3jgTIGplB+d0
owN7Q6I9mU3rRY4D30OUwFkAYZOFD4bCpIOjsXxYHtr0SUYn+a6KhtWb/5RchxYO45Xw8k+M+eZw
faI+UB++sE63obGA8yoAagIP3cJAUV7WN/SGHJaAYXNzpGx/LB1K7ef/9WRD5MoQZZM43HOFwsV4
VeC40idOJ+CwnUQ8LhEyeCPy7xCpjljLsb/zKy7BWaU7v1ewi3c53QJQMgxT/Cwd4MCUXFIG47nm
7f4lTws4lvCel9k/fyhVGCZ0WQOMiTzuqVTVwbRr9t9gK5qL/haHgpywn/QBss/OV2L9kYh58rcZ
6Ea+jCtXRDabeJ4T5TKqNeiOSyRYcDsKBMHpW0L//WfkPGoHRNq/UyC/2TTP56LDRlc+IizKFnrw
s/uNncGl2Szun2tjfYLCKEZj4KOTmHdYEu+FG0rgO2Ybn1k5oe14cnKYvx/X5+r0jUPdWH55c2ja
I7jB1BIYCyoyCy1yE1KL9NmmKi7bFCplQV7gvxuVn8Hp6yq6v0Ig0665ujTPPG6xxz86OnjJ3rNu
ZxhbtFEaPjTLCjDUSgRWiyHeWRYZL8GN4lfdyKWgR3FD/E4nIIGWj+AxmfNwf3kSKMcsqBzpBf6h
A/jJIeYARRfv9xb6LyAlybS34LAfWpt8gb3RYoQFmdN4+hpjTGyVn1CCP03DZxCZexnikUXzvXhk
425A590SFW9/XCXFrT0cwipPR20UKVBoURfsG/V6UkGxzUpH9OW/nuJ/4ItL30sNZbH2bBQDx8r3
U64Ju/4q1IQeL+RRdXuUsUbKE49HzPuw8qNncSC+iDYd2iqg99olhKAtg0/ynW0lSZu2QvULuDwf
ILr7lYSSQ9AfmMWa9fs1NaQWCXpndSGnFxMGb61Qnxj5FNqur00DdJKGP4wdLTQL0+2XYsEAvlVL
mR14/xUSQNjJ+m8PDuZM0FQzpm+KYA3MshdpN8GdhHpr/U3GwSYERWNxVOvt7eNVsmt0wlK3NGuv
kvBDcLSP5fhTyAcM7EMP12KkvwNuNKx2C015n4eW/YMs2R6cMrmiLpUChdXSsnnpPW/qAWGBGOyc
P+1mmRZuiGuWiue+Hh/l23+3GsX+ahAxfPGgDw==
`pragma protect end_protected

// 
