/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Fgcvq9yodAEyu7zsWWZ7LwHLqer2uRdIROgj+b6me/wmyj6mu+r4+a1EPBMoGlf2Rxb0wqrGm/yl
7FT0a+0gf6RIUa901Ug60cEq5l3MsNjnNX0EuQ9QHnbWnPHO5sk3W38XYr3s1DoIymcMyzWSb3j7
DAgt+R0iGXGbLJHe2UuAgwrybNhjpWacbybFOYZoLu5Z50wmOHt3p6J+gVbTwfuHK/f+KnS4VtSD
EJxx9+hQNEvkukNe5IcvkATvsJ495o97/SdF6+o/UvTHUZ0m3la3MPtrbbqjxbRc5d/SBaUYwJ/0
DSKgI3IBXs0nO4MGwCQX4Cy0xa1KtNy17Uqy4A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="YyF30NSJW4xBU1bz6CmJ7uDDg1utz4oEiyNQAWYk7H4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1168)
`pragma protect data_block
3JkMrY1IEAXvStruy6C+3uh/9WhMi9+PGUwiTLF/rFT8/uU5PEQzLn2D0tCvB008AeSkVify/pjC
2VhGBc+u0ll/erzEDw3YAzB5kcOOClFu1/zuXOS68KBd3Jh0xm3ZtAp9WVR7/4CVtWC7oXfs810X
rBPYAy0/qC2BxTHs52AcmyAJWnc+VWhZh59YZR5DwCQZc0mt7G4JD5EyStzAchxWEOoi4PY8xuJC
/d6UGS1lM3urB3uBjA36XbhRsbfzTAZdC1aPYDT9WSa4h5ihQRC0fOt4iuZ23vRafKstHHprcKeN
oW5OCZ93TSgo1BYsAR0o+cgoj0aVHoyhf7IXmXCk6/4Wjanhh3lH375oWZPCfDhqzqELsxku/NYD
E4d3z76yPPrMh/HhjN5GtehwMRuAtbQsv3UWAj7Bju/UuWW9VabtzzqjKVe/wEw5BS/9Bd0LAL9n
CAYjrwKKRxAOfBmZYfwkoxpeZ66sgt/cPu9H2FeFgtO9g02K7pFQs8DGoGQEuQ1X+N2bz3jmYl/1
ISgYO5rtU4vkzeNcIBU+IhJP5fGIE3L7zdsBpmmzGxt8H9uNddU6Fz7pD7D8pycuSx/aLgr2/Vbv
qmHPVV203ydw3wO5O4wPW1EQKgROIY/xgwqE0ZagsmNqbivhgB7s2eAHHGFgcEklX3E099gMSyvH
UHknSU85mQ3GIZ7Emhl+60cfDJZEB4BKHMTPjT6UwCKEj5q6by3vk3gWCpB/KiS1Z+J4Li1NZd2X
LrkMdGHwzEolxAdCELRfV+q2Qg1MlIrgmYxxnksgn9vRsxK1ATt8ryExcOaAJFTZyOo+e7iTo+U4
GSATeeo7QmUusUPEjDYdrj3iiuroz3lBEYd/X0ksLELm9r6xiIQ88F0PgYhP/3po7OdVlWrrPS/P
oMd2D65tO2UDgV2/cbvtsJ4cJORVy7JFHJzG0qZkubHFb3DtnPq0nKtCRnh+xci/DbUSnYnxKg8D
V4cd3ZU8+2jYIJ5HggcGQce/sPdQc7k/IsR2/nangKbxC8ZNIV0O2KfESiC+NjRrK5+QgiPyXP1X
PEkvixUNA6/rqL61PXYKHQZgmjSoj2t912kWsRdOr7uAbUt+RKKiOQh5IwPgj6HElBgQeoohjmiB
XnqnScR+r8W+W6RcoK7DTeGSnlWFIP1gKbUmWc1BvkptY3Q8byTzFahztQW8OxVLh0qZgFUVJM6u
c7O5eAi+6WRtUncIAPvjkhfXs2ccvQJsnWzdJzECT24I1i1bOTlkYuON3odYBOK5I2uGk8ySaQKa
iQP+aXYb5GXHCukRzcYQ/vma32Zh6LnZHbtJPpUZDFnuPWwu5AUJ1xrCbv9CKLJQrv4Va6eQuX2F
pwhEEqASuiDErfjk0KJa8772t6m/7Gu+5bh/91VUhvVqejXwkfUCZdmrUHMgda6Z1yHJu+8Mb/K7
g/tfRulgZqTLcVeMt8DI8QD85yq56SQN1t6jp0xtDURF+uEDPQNhmH2eZJijqCyTI8OwNcv5Pf7p
GQBawKSoLvSx3/B+fO7Xn9GET7WWgLDfaTMgKQ==
`pragma protect end_protected

// 
