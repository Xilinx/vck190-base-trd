/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
l4gSYexUXlM7ifAaBP6t2MLRFhQaRe7Sma+zo2L28DiA8DDFN158h0/DaBr1OsRaQKqTpiBWurc1
Kc+8TD5uaOBbdGAOqQnBtAA+GhRIwIir9IbLuxBMnT/JmOaK4MUYPqvoRzrgYyXFE5yrJmMkU220
b8Arh6+dyt3Bh0bC5r9kA89v3D+ja9uQnY/8oodAq0Q20j5GmOBNL7A1mEvLof/A0UYhDRCv3pRO
FKF8KrYOR3RN8PBeGCM1EFnr+wW3J99nOfKe+v5+if1arByO/0BxWK1JYTBdcxntFYOrk/8juzWe
cyuQA25yLLNZSsEfw7pTdA4YqggvIwnYX+4CfA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="nooMg7GjkDsMTPG3DLODBuXednbZgjpzUjgowzton6E="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1136)
`pragma protect data_block
OIw4y6hn7TeoR9JbrM9EZHSSqwf8hSPKkPsRR+/FodPRcDxFSc4dIItfhXP6BWnOLi6NTlihVecl
3N3qAMpEAFR+7a5h1FYFtbm+mYfrwcT5ILzALwlwtcppKEKPpqG511GWoS9euy0YYjUm0SXDMyIz
1/stQwRex0D6dR//n2OES+8Qa+RRw5RFC8TyANgLDjDMu+9c8pme/1g5ll2lFqai7Jr5UhvtSKOq
wGn2GkFudPnORxAAkboL1Ozpdf8M92J62JnFbVVjqOmTF5hfHIRDEj8QF15F9ah1/qHyJLlifBfn
npB9MhesTwTARartC3sf8Jwv45OFn3b2NbR7qn86QWT8FRpd0UfSJks+aHsWcAiifMcTcatQHBMi
fl68q/KVmvZVNq6sSxhJsW3A2UE/OhUc2J14aGlSm5vKFD7l0d3bV+a7bmUhccar00LpdeHiE8ca
5s6c+SpMWzmot0ayWME24l9/zOEDfyWdEZQArcxm3RlwVxHoVl1oPEMQYE74pRCxuBbxn+/BLMTf
E1B47RAmiSRQkgGVaPMxKTQXeRFUDyDsyp00cwmXwBcJ5C5bb8KxQijejj7XV2nBq2eOOEsW+pO1
cWWYdGgXajjm/YHMW4blUl+WDKOlTolo+midWzT9HRnaikP/BdYU4ni4H+OLzHZJxxynebOl1wms
bqOScQDM9oOiKS7ZeCPWAF9eruUo7oRJY4BEpj8rbG6fsJB03ZxBeQWePCWu1Em3IVDyXKe3FXix
ewRAF/Pt2dlVtxb6wqvA80IcQFBckiKAxe/noowB56hSnzOiIvkhjD/r7uSt7x8xre/bKbe40EBC
MPHJxPJBTdpG9M5a6iqv9D+yWWX4HvNFWW0ubTL9vNhLtD08ak4WPbwwLkNBjc8D6+OS8Pm24GE5
62HeRphvMMXqI/B2Hw11pBcaM3FdPalfVQtjkUyYfWJdIRI8x7Flsx4CY95g3DktRnj3ngvL3TIE
cHdXLfCYU2m1nMr5tXjPN7XTAQI8ymKNbWqHOBfp4CL5DWeSjxiKPYmcOO4lV9zkfH3N9TDwxGlz
ldMItefDoDHYxffV6RVOTIVUF+C5Hl6+rpImGaHqDt37jZjSKY5aGMhj/oLwtaoZjILtLiLbX+s0
V9kJ+sgJoP9NSiWGsVuLKk+bnJhzv8qhV5jie23G6/DGMJhaw7p7/RMiGhNwIHfed92Obzj6vTZ/
UqZYiy3I49+g9MSM+3h2xxpJQzCgzLN7MySnM/n99L2L85/3Pz78Uoyo/pjGwsg98rxwXtfI2wUo
ILWbDXqH20qkotVNz2xThkEejUf2AsovAZKB9U1lSwVLT8+CfOhG07H1h/GqY/dCZeWw6jHoA0a5
/PA8nj5aCIrtzlNXn2GJspo1+j0PUg3YX2BPYIE3UbCxYyx9r3BfGO17K9D4N9Cc1GvLu3/73EIJ
M0IYkx2w95RqJl9sBDr9e8AMTFE6Gb224XgYo+PQKpnfrs82v1S/pJ8YtB2at2q6zQ/IKfo=
`pragma protect end_protected

// 
