/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa", key_block
WnUYD0g6/qDSYmWHmuZSsLHluSdi9+myTeKuKMxZY1YiclF8fPuiqftouQOib18cBMrk+rhxXYqY
YxxEMkXifSggXUrW22+E+kt/etsSl4zJseXz6n9xUwZYg3xlqNjifu0w0ji98CtnXurauen1JNyx
O3YJAh7IDwn6xZR3LTGYOPxMj1rA3ndIEld9FoiPlSfzRSRuhh7ozr80Ea1y9ZyRdn6UvlSGNFWa
K+qWQ9v0fQI5P76f/h7qmdvfXu9BKunBkypsT5BoGjV+yipSZpdDPJFuKi8ZALQ4AfQwwQQ4W9Ow
ic2MhxBJty6sWw08okzuCC7DdaVW8+sh3E0SQA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="GeeiI2S+0qmTuse/FWjb6tqEZItAqGIcIYeurwykgk8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
1KvCHb5eogwPJFXkT9BIC66Z5d/vD8Y0LoXeLRDd9RkF0v9jeeyleY7h3UQcs0WLQCH4KDyTl/gj
afHwBubGWTMlAHO2YdYkjhXKvWErPpwasTAXkodJImT2mSqrn/N6qvL2hS3EtsqLMpZkC3zH436a
W0lqRAyQatRbKxUUeCnuEkZGbGO4g4X+heuIH9J6kko5+HMI2AX80rukZ2iLtSpuAi/4VcOghT2p
CdkY3/vTU8Wq/W8a44wkFa7tsyjuMAdaGnP8sjAgXmu1rvoElNEd2HGb9pbYZNtwxpq24TagiY9O
zR4T/jxlGFXZ5ug+Bwu5pLL6N3RHyy3ua5JgWofftQbIXYhZhuv43XAIE1upfmOFk6qoMNTKLcLC
CHwpG7UDGmze2Ne5ZzU9f9pS3nLXVslsh/UABAADzL7O+4qhXjnNEKNQ7YYki2Ms0mjIHdCyhW1d
VHDSj8XXP5R+7eyUL392G9gcgZF6yoTnUhy9ZIs8ae9KJDe3iLL1hN9aWHc5jyouvx8cCLcrw4er
Mh6tBTmEytOSe9WzFWc1efQkQYA0bj5VG6oHDK4gC8XbD0KwOik1nr9z6pq57yQ4U70sNBMn7fza
erTlzVRMjdkkjEWF1R3j4Lmkl8sZOlB0QJlLLWfhZXsPp0xuFeSaMwbWqk48oo5WHLivSAeD7dNU
G5Z/PU4S637Pn+7fTQvG6hdoQ06sMGRmYkbc2MlDCkcnFMKQwUu8zey7GjDYPFP/r3esr1zUzZac
1P8q9svN8I0Uoc5BsfYpJiIFHHJpirJScHDtejLUnNhR7WZN2ade8ESyEftondv3rKdPG/MxXReG
q3GwaMp4OPYETejNxXHW/dcTZv/6b7tDCciYZw4Sic0C8YYmgVrNCjts45vjpAIW4t6pHSvY8/wb
GenseRU7tkyYU+B4bjhJs4+M50E+pnfQ9Y4RmX0IqfB+yeElt98IYvRL7qXicZti2AaDVECmEPkw
jA/UtzQki31mGVrqUWBBKzFLvN51BTEM5jTiihXQwaTpcVqEZrf4G+fpLFUowCb5WCubzsFmCIxP
0tZImm4dpMTUCZqsfFBebBgC5YFzTbSjEhJDHK0R+7pFYkg1fwcEvnOId7sNK4IskyJFRNHYRFk1
Fsr9x8hx86LkWh3eC6D0+5JjBbEw8TBC5UR2NVDDZ1kTkKd3C7DDBQE4uVwivXkwhbcRhvkK+SRa
o/X5GzcQiP63tNC1y5j9QiLnI7kK3xwMwJYCdmtXnUZyAmPGdiPb5zq29ltJzP8ItBC1vdVr5N6d
CRu1oLvWOwNdFA7+I+WxFlRRAJLRzLBv5x0cUYtIeJ0cOAZss/SPwz/fGMjsJzynHgbOd+7ZHltF
Azy+lfk0dd5zB3wIqpa25bFcgkUEBpMLYrGItM9l238VeS+INKoYlQwNMuCvxwgmomVckQ15iWiS
5CFl70Y=
`pragma protect end_protected

// 
