/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa", key_block
WnUYD0g6/qDSYmWHmuZSsLHluSdi9+myTeKuKMxZY1YiclF8fPuiqftouQOib18cBMrk+rhxXYqY
YxxEMkXifSggXUrW22+E+kt/etsSl4zJseXz6n9xUwZYg3xlqNjifu0w0ji98CtnXurauen1JNyx
O3YJAh7IDwn6xZR3LTGYOPxMj1rA3ndIEld9FoiPlSfzRSRuhh7ozr80Ea1y9ZyRdn6UvlSGNFWa
K+qWQ9v0fQI5P76f/h7qmdvfXu9BKunBkypsT5BoGjV+yipSZpdDPJFuKi8ZALQ4AfQwwQQ4W9Ow
ic2MhxBJty6sWw08okzuCC7DdaVW8+sh3E0SQA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="GeeiI2S+0qmTuse/FWjb6tqEZItAqGIcIYeurwykgk8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5952)
`pragma protect data_block
1KvCHb5eogwPJFXkT9BIC4y5w7VLpxCd0K4dh/GMkc67+ESWWoQ3xHPJaaYdsIOM7r7oOGfRnj5i
N1slRX80fF1mQ4dWW0iiSvVuFou6uQ8XOPNI0YDlSX2AisKnF3Ls0BmIjMNIwGnPQguitkEfISJN
KkXa497XGpF4/wjvTYr75dCsuHeaeHtmTPNAP3IsYrqkYDnujDHEtZ3wMZxepjA/1jM0wZaR5PjK
EJrl2aRbar1D+uYw3HeCqe+dAtXZs4/U+LHTsh4GvFDKSP+DrXMNR21IwjDVmDQd8FX+UBT/bgh7
G+j+iOq6gO7f0RBWH23dbSJ/AktHoXxK+T1tNpeYk0uxeeM6HPfjcRAPjq4XpJ7RDPCChoJjDI0T
323SUX1XObn3SAOObX47ZQ0RFsz1G360R1jRE4AHGnRyEIdBrWJKkE0n8FWvgw+FTyLhriVg8huB
UqVYznxHR5qiVG2z9/rzGCAoEJBqKT6n18SHHYjtZQMHxxpuYtBHxJTsFOvTv3hsD/kaU953DvD+
o6GIQQp03dIzn51BC2kpaajW07ExDhT0sa0NsVuQ00jW+Z98PDlhTGvoOSXhkDR1FmxthASB18DG
dE1+eaLKNmSy8z5lKFPFBRQ2cJHvgs3FJD4TfOhnz+3r6Ez8iFVegfQnV/744VXh3FZwiR4SoXZS
8RykxuJwz4yJQlUvdV8P9H8JCwu2b/fxisZkJufaqjjJ0Oh/L9rLoCRPyQsEnBOuRaqUjO7LTCWP
kVN9ydmN1Jj013BWoGb3FGFONnYVej555LqNg7nyKSv79MCxobp2rJh57foiHpu7oBrDm3okYVfA
TmErrgXu04T5p8PR4PCxilhsYXfs6gQBkVnL1iy9764XSbIui9ftf498rh8TSG95BEFowSwCrlCK
Suy7F1nMZ/ZQbvAsvzZMnVhp0i9dRGrqFEhhMLzq27BxIjPFNkiQD/PHZJ/biDfKh8hCG8fNXIJB
9sWhbL7PHjl7jZfAfu/imA7VD7UEGgcZaFJmAfJjHVQ6/HB693QOFUP/4GDu/QL4dZS2ervP2nVL
G2eI0NmHhaYX8MkQzBJ/hsQrC2sUrgcMgavruRV8fgrMkvZ18WS9RJ35HHW3KCqDrLMv3IAmjNV8
XnTyyVvQyXLI7Pal9KKGsABKTsx6ZlSG+AVlZuxfzAxQgz3Q+BeczFYwXr9BWfG9WM5g+jKfWvFi
9SJ3NwaR6Q0w18RgNiRD10BzD47d/H/h6n+pluN0viX1m0zp/Pbv7qbdYyBbF9ETRZszswlVnuoS
lqKNkfGEBpfkefV5mn/8REqMnEofs0llsd3cpn3McI8B5yheP0X4XgvTF7dlOokMj8XsPDh0QhOE
oBnxyB9zIFrvfnMwovyF844wkxFjd8AyiAD3WQKzrxHfD8QKHp5FU9uTqmrJExWfTcQgbpMiy3Y5
Jt7rgmS0bunR5LCxTmrtbyWv77HOkdU1tIhlcqsbfmUchLOqh4sc0QvFXQDoL5S0EmE6bJSzbvFI
SaAhOMvv42Yfw8BhRL5lC7uAXv9Gm+MAq2zwxPmMsFqmB5+Nb3+EV1BfAKlh9RYptCGW2gNSmJPH
yslvp6qjpwhVVzpBl4xuh41fMo8iRwVDTqNhA5dtCv90TMgUwsvoUjg+d/KyUmMzofJIdvertrvp
6nsOVO5Kvmi7tQuFed/N/5pgzczbSrP+QwK8XMKEmCD6IEKaoB59lfm5oJlmo9ph7K4hG1a9U+u/
dbcUuD2XrsGaOW5KVyB3zBiwXyDeECz4iGbaN93z4KzD4inoZlH1POdsUlZczTqdJue41yvVJJ0e
yXsNsS4MSHRqOoX2mckiH3FtY4inSM04yewJ3cHBxtSIAsirjxXIlb0WT8zXIgjpK3el3na46Utu
nprGcT52wLHCsHsx2bzYjf49i5Rhb2VUAv/9nYPb+RQKldjsAeKtfJOXoHEIkrGJOsgrlw1le7v4
QqStPXhTYrbZee/phwTmpmZF7EBdOum7a5oa4yZWnH8i5HekgN5a15XMZrA3NYlaSLoOK2VVZ4FJ
mlOHbU9rs5fKUmaKDX5EcSI5nYXQg8JwgpXqtVnv632JjTJU5Rv96G72DFun9WbZ3qrk+/PsKpiJ
mhxMHMZElz1QbYW365bCQub0OC4cz/6kCwFXM7Qowlwhl4pETveoA3OTWwYcLMaVw1WbytaXQb2v
V1VIC6RmA81sATp0WR7nXBNh25TjdcmlvVydkMUbji8trCik10/YR5PXjW/JMuz4TQPQAnRzJdsK
NVeLYuZijzc964oQ4/m8R22MDU71GpP9SUM5sV6MYuBeF+Rss7R9X35cpqODwPawMXd5YYfIOjDN
s4EyCb9F3DOqt8ELeie1j7OQSdVA7TJdbxA/DSoC7/HPOkrJvpAq3p+P2853hNJgkMZDssdc9SVZ
sGPIvyB/OgeHMcggfugGcf5tDoYM0gEejEnEeNTYeSwIqzMdy6JhG7uB/EcNLKyguRH4YIEgFqgE
wyH992cw9jjYbzjj+rb5pJ/bW1q2URcbSappwrg745r+mSApyYioysGKeQma0Pnd4G+5Rz4MSEpK
ULd6CNI4fJgq1oxEcYBo23o8IOBKE+eiyLWUz3wcBme6EUiB2wIwZWLYDAw07lds9Bk5mKbJgVZ1
iS8C3FqVK8+nvZe+uUimfCquIHnFg5F3L/h+yzeAtka8W725njaVhHKiBmJ/+N59y4ipRUfa1og0
R7yJFXx/U01dLBGqtXpTCPyH51lkegEOx89Vh42FYCiIzj94Iwdu71rEhGiTKrIeQlKOOe0RQkd0
+udj7y+OkyhGoV5pY0u0KfGM6FFPkA31bO3TBwFkk5LKc/6eUSP5W9KUw06QZsS/Dmu0ht9JrNMh
MFqAvSX5nJXCBLnvpqvkopoF+Pmqt5LOwP7yVsdBrUmJfunEXsCyhxF4n5Ka6IUuammqoPf10Vv1
KWoTn3IwKpNlH2KQLCEx3M/6/YMC3+j34pJSmtel3p6xPbLNYfjEsHXGmcxI4yr6ipi+hXCAYttv
zzDon4/45h7Qx295Ip15XWSmptbSXaLHFnR9uOMU03AatQvlKpAMgyKLKHvb8xqTzXsmWfVbvj1I
bqRbO27FjUBX00FB/m2QQvTFYSjKGMp2flnI7MlNRyx8j+vQMEw+tXad5LsD478mHYzB482aR1Dx
rTesxpz0cy8BIgbhsq+wWxXcE3o3mvGPRLk8VogKzowo8xAI0SjU/42/uOzEcoZG7qe0d/p8Vk3s
3tWfkwdYM9p3Ch0FF+x8VSmeBSlpdiBn4wGMbCW0oyV5ufDsyE9xawO+14XuC0gk8fxm5NlwYNYG
eCutAps20wZsRdmVtblPMP4rFWfgrH8NQAlCZjuu+F775COJc2TmZ5HjCSfY3mkAbYXfUhSfCXkD
biim7WsQ5B6MV0DqfG+MHU3Pn95je99Zm3NTEOcxfyLp4WnjcmzjBx+ioXxi0ARNAVhc1ZE9u7dK
LGnasXmnQkpRNTNnbwFVDZ2V/o50svGJK24DcKrSZ58iVWQtGyaX2+aa07gU6pl3sVYRBlQEDQkV
T0Dtsar6wOhf0MwnhcaZJjobcqfDeVyMUctlshe3mCgbfV1P+lrUaz+Js0iYXb2+qJO3Hjc7xR5o
IWhVitVOZM3GKDMZpUIs/3Ozj07FkzQuDj9onRoZ5NaUnUpul7Ab/oWPXFnUkZNCqYMPb0B7NL9d
gjPpywxxzoOULNuChJNQ7ytc5Mcdv4OoTPMmAu0P2SS75YG6h+yZ/7Zryi9hnCGv48sdAV4rGKwE
OlcBay3vXTVu4+kF2sdFhtAkpCTwmXGCPxnn90B15Hqz0QoHXyZKl6u305t4GtZe4dRWoWhjv32I
gKuHsIh8iloAsU0HZJVLGzZttMK9GW0L0k5/yDPTOIetyZe9UEsKd4AtGRGr+pZSZ3vpzP63/e76
R+HiiaiRv70hDw37NABHBG8Z4PB2BOtpEJvpZJvT57PoU+QmCl1QZPzXoWQyyv9/krHOQTyFGvNz
Do37w77+T6MypdLpZWO/YLiC9nqO8tHWpzmQECOa7tyzZ1ONoBRBxzPGBJUVfMX5D/R03D2IlsAz
HpCDOIIQ3+vhNFzGSRWVL8gj5TfT+wGywgcTFUxaNLxMUEghn8zcybUP9datAKv22BNKUFaO+pdi
kbNIiw1BDpTgj6HfLIFP6L2K88iAwR/1NChmIaw77kLG0kjZQ6BgK/eYc+9fsN3YPQci6fB7BGHi
/MYPwcZWsu6i0N2DzNQMHaBP+a6qqCV0GSP0VPFtOm13ACEFP0oIuEa1IvsRIuMeb2QRzQBOkYcE
5oBdQyf+w9hQAFxVAx9+iCmdrSj2Mp25yai9GMlaOqqopDKmynAHNsEscz2DXQ889GVuNYUsDy+X
ejvnnrhzwQkAVsGMPT8zFDnAANL0sRA0eaHcJUyEWFURNQHEdNVlFvlLrVhQWw9IWv2/qy0ok++W
9mP/ylfaILxPHO7bBObahDU7VWbdrrrmKpx0LY6S85ygdurpkt3MwNqkg8/+AF7/JxAQuOpglSwz
hY3yHwtgqvbs12zrxc1XuN3I58blwOPMH1YnVGBBY/09EwqC1+wbr76Hq9Lehog6tjNf82U5sxe7
hXDDaATrljiWUf9MDBmiq4l71DshRngtDy91YiSISPZC14zeWzvLxC/ZKgB6MneGEIiL5lVRsGRy
asF2CHSVkVtwD9SCsBiQr+jXtMED9wl7O5eYMXd3Kj1QAK+H518Xc5N3khmQ+8ttT6KUCncLpXc3
BauFEbLMHm2TMUSbN+fm1TYjowbfOX9yw6AesvBk3ECGdZiBzq0jFmJhkdL6DCrwkhlPFYlERqbW
DQF0u01EIi1oK5V3CSkKl2d3/6TrCcerD7MmsE4SHnFCRXV/L6/DsUtVt7XmbFY6BJZpTMHsrvTh
3WRS+5tbnuVfVuGNr8Z62BpOO2fyYFLIPYZ2Pl2Yj6mbwM1RB8U+0cIFD9M2hU015ZqKwqx3TvU+
CSguc9uTFbaA2qhk3BvXiphcPzgS6b5nKYN4dSPQ+cmxsVSFUh/Ys6f0O82UFP3Uh8+J6p9TELTb
QQSmTUAW6nqCPjp2AaNIFq0Hq6ibiL+7dv2s5/SxJfC919mjx1t8kboaFpWyzqyZlIWdWcjQ3mkR
94EfwofG9l4udblrCJ8dPT4IViN2JAwNAY7n8uNdRFxyshhggzs/C+hI4S/8noM+YdBcJcBox/l8
YbfuLvgcur/7GqkhKMyLYmKA97CEzJSLm6NerIbgV3pBCIKogILVP9ku18zLKJUls2EYNSgs9hI2
uFVlqNWH2abIyi3mhbsjIwEGlK2lH8ro3U6/5KZB4lOx/BbRfOrxMAN7G8j2wGjTf6XaxNiJoqhE
2X7zQvnVDfDB2JjsFIsDqUe3UC6FKe+zm/NmEdgMJVNXZH2ACeHoEqeFTD7d2GNU6czBEayAQ0Tg
DCMdA01rvxVmEdwTIgY3bWlvQUvBPWH81nBz1dprTS37ShGekCkpIduroCw6D7a2+i9COyB2n9dy
dVvGU7Dr4PVKV7Ishzhewt/OxHcWQTsHAvtXp7ppo69M7RRCRJVXqdq6m8JmBKeobtjHWmzFTCWb
CDqOgYhTlIRslXr151Qoei5LcgcYQF3yynCmnfOK4DEp+8+UNaf/p/aCMzUNxGE1q9/PSoclY8S2
ySw+93f3jxFQeH4+9Z64EpHFpkwR8q7KxudASL1RVoADA8Ks6yGgZxX0ExKn+UM13DOhwpKk2TXl
XFnHUF4CkzhcphRnRX7YwzUHq8fp1jJwEknDeUDzmfNtSp9D95q4135jV6JKASRzjN6LmQXZD+FM
JkjHIRctJYK1pduXW0LnKZ0ZA5fP+fuiq1xXalpHKPGyj6NFQL1x4Jigmx8kqyOdx8nolhXs0pfc
bPwTpjBElLap0VVYlcRSKxtCr/FXygfFsmQ15vjPVGBfa6WbCJm5nQ6UXGECZ3Hhvg5bgf37Dmyf
F601WTNqoMqIy6X7Sxi+H2LbYGBp96G/uMwqhVJRSzTlPETMXOaE7A9l1XA2gJdb/O5sREOLsLGC
IqSlg+0l8BZ8723jMa9rU0I5WcrE5exs83dFv4ykLA4upUk/OqsOdSn5iJqIUxMNMxR2PbhT/DC4
NsjfzqAWDWYQ/SIBzMbQsiNbyq56rnbTosfKKsG4KCxBoqlODPJh1H7Gc21U1jvgRNSW4STqftyA
6T9xQUxXB17+rWTZwzFlg2wW4LMhcPIZNmnGwDO4XgE3Ze2sVmMGaJetXgC22GOQpDqJkxqTpFxJ
hB9N7sqv6RDdU33mLSyQOjieN00liRaykBzYanjti1vVsRQQ/2gxvrH5U2jnnkSvXHVvfkWLWBUO
W6/4YdHvutN5+fIB04eR164A5ke31bya1O/E0d625tb6PitPSgBUtNfHsyNs3a/yR1LeZIt+FRQE
ig61H5iyc0a+OdFHPE2GmuERv2TD21/ZASNvfcLFTGB5V3CX+NYi2451SPIsWN9HLMCThEeYtBMe
bQr6q02k26uvWKMsb4DAaGEmHOFX1guC+fOKqzCSrjrSQDMhRXQrBZfINQN7UoyAjavxmNXS+zfc
SicNVNsIt8Ak0tb0LissisrdKqQjFeHxIn90zyrpDNKpM3sd+t/c8KGw3ztXCvNOxv76GGnNg0mB
dA1qi/92biU4AwubOaWcgXudENnNHiV2LWX7GUCsd6p2eF59O40xcQ7ksWp0iHlAzUYxHRIZL4L5
s6t3x+zLmJYD9B9zFqJ1uIyDfdDpCSPNfIedIruyKukoAbgVkcCqtjWpdgPc+jauxFTrA7GTu6kD
yxkXIpyznCIlQ+OXUesXqYzdtsWzB/NeeNBGDH3lKNyuQMHe835EY4uhn82ZR2VAVuMtQrMtjY4g
S9g0CKmAnbi5MiAkJ6KOKYmHBSxI6s6vLulPqegsp9ymcPZyX0ACa+rZqoZzRjNiG/NvICM+X5Wx
MnIb3e1d6T2UlEKD4D2zTj57bQJJe8RIA9qToc3RU4Oz3npbil+2/LxOVE5e9Go07MK6bVjC2eZ6
plNbwzyzNiEeFOTVdV/8F86OerYB+k2FVKBE6TXuh0DkKp4eTu9cH/XwRDNbEO0SFFv0HWLH73sQ
9RzDK2L846BkgwD2mBc4QxWq3sncf140O01XDW6P1LyYSCYwTg7mRT3F3HF7BeT3m4RzWHWNumVh
INvtBmKeK1cFc4IPw+K9niAMrAbac55XDRFEedBh0gBEHto6d/UQnACEKXmmNE8GawTEGF4z8Bje
HPh0AxysZyAhIV+mxRozgutY+vE4PDSGxc83hEcnJSVX4omEuBdHnAYxFLI6PUJJjNYH1S3Tsech
jyMQ5SHy+ub6eMEsG+yt2ID6f/pZJuBM1rtdCPTs3CdRiDn6e5kWrm5OnDWMm1BEo42oLUgpWemE
Tc33SUwgVPCJPdJE+sWCFmIsGdwrJG3i7H61TZplYak3cJ+DeDJPaKBIcCIF5N+BVbBiRE1L33Ci
Q5v+JuhsYQeS24nlLcYnnMZnIjJa/7CLz71/jadegT1b3JbH8CYqneeyERD372pwuCL7Cn5DoWor
ihuFMj8fG+/YD1AI5SxlEoOU5Me5sQTarj8e75QEFYKQrpJHyYsUhkzn+YhBfsJwMiDUdstfrsSC
irdoFAH8iuIqXeBLr3CJ1XwuTD24k7E8JupPLB8XPh3pE9mtxU1KaLkp1tlzDOjVmXEshVTe/PDR
o/T0ThXYAKH9od/KjbOFT2O0To/Se574ehyIobJMX/KCjvJ7ZC+bCLMceZoL+ig437M6dRLUS1dx
dyt7uxSbRCq6UpjzWrB/s8SrRBlUDOzNKEvHhF6fXwbV4ftOBhhshNWSxY8lJ3/uxiyAgfwZBbW4
ljk6s28RlNYpDSVTGKDaR6o+bdOH9rPl
`pragma protect end_protected

// 
