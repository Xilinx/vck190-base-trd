/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa", key_block
WnUYD0g6/qDSYmWHmuZSsLHluSdi9+myTeKuKMxZY1YiclF8fPuiqftouQOib18cBMrk+rhxXYqY
YxxEMkXifSggXUrW22+E+kt/etsSl4zJseXz6n9xUwZYg3xlqNjifu0w0ji98CtnXurauen1JNyx
O3YJAh7IDwn6xZR3LTGYOPxMj1rA3ndIEld9FoiPlSfzRSRuhh7ozr80Ea1y9ZyRdn6UvlSGNFWa
K+qWQ9v0fQI5P76f/h7qmdvfXu9BKunBkypsT5BoGjV+yipSZpdDPJFuKi8ZALQ4AfQwwQQ4W9Ow
ic2MhxBJty6sWw08okzuCC7DdaVW8+sh3E0SQA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="GeeiI2S+0qmTuse/FWjb6tqEZItAqGIcIYeurwykgk8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1486576)
`pragma protect data_block
1KvCHb5eogwPJFXkT9BIC2M3N7PuMQaTXKJRnoq6xPfXm+VJ64XSDTljyNSnzwmuy7B2qORrSMcP
BrSqzCnZtZ7tbngy1CsOKvatG5/2QfUz8E7nF9H0pd92IdwEEXUA/smxHi9eiB2xlQOHV+ZGW4p9
3c2NhaKjPrq401WOF2X5sdP2zuL+dcdHIOm22GrNt1s/jw6/jW7mfAnEkIEPM9Hl4t/ZSGxD4pqq
NqpKQ0Kdj2LD0/CfMAaup/ua9Ypb5dx4EUGLSOOrLM2UBzLwRsCWDUJ9/VVewV1REXFjgzAYtUbG
ZL+FlsX4RAqKtLW6v3GXXpA+qpWY8aLDbWueKRNp2RmJLB4WFw3kAT/EJUZk01Ne/wch0awSo9Oy
3gZwQrLFPCY5DAPqGLJgZdBz23qRLcEaJEjt7VIkGGYA8szEVAZHQW2w6Hl3bNvRXqx1xsMOCV64
/VWe18KqTRy2u+cXRRdEEjVWRVv3qm0X1yP8PsHC3hV3uk0dC+Ntb7Q52CD1eXDMnE3mrufe1FYU
SQ2PGr071FZkMc0NYnHjlohSYx3tMYoHGAYvJHY1gbwzZhi/k+1MnIdIjmf3cZ300cfDND3GWMZd
UCo8YOXKnHjsIk477Reh7cIV/9iARj3ZE7yFwXN8E6Z5ktxJq0ZuCB9YQ8/QB3O77rjn+UxoKXaO
LJIdsPCL02HJhCzvo9ZyhDII0DqA8F3UD5TIa5d4hDJev/Qpwy3ux4vUVympnD/Y6UBrPi1RF9I1
VrlZMh2tpQ/ZIj5aEGEMA37ue0Ge0qPaxadZmuqMeZIJjjJApT39vErvzpFTfImk1u9N5zzclIlb
tXlDEElE/9BIGhVjiDVwqc73CoPG4vcj3IRfr1jzgOhP1SG6qs4MMzgBfmMiKTkm6B983pUQHbIo
uPkRsAYY/JpcWkaheMF3v2C4eDAx55m6Y3cCNCwWv9LRNG5Slo6XpTcEspr/Y9kMznmryi/coAPc
/eonG+WMeaxe8Dq7xBgeKk3/ugWpbQw5FJBnk66R4zt2yCvkRc8nz21To6/pU3lgCRfBiLc2HVoc
HDXOP76nxyM4mjcESbaWblH7En4j18C8yaHT0qFF/0ECthnGg36VYW/RjAUPOQDQZowbzlmRT4O0
eae45hkHf6HIF2AR6X+PHj5fsqdOBmNA5noo59UKXZ1QiG4cPo/KVHbjn5slcvkCGEo3wCQCFrqN
a5sNCcAFbRQRA+2eZlk2NncDJdNvGLlqf/JaCXJYvc3NQ4uUmCnp024FQFNcBPFKMoZUHSkKGsHP
WkIDvysglAkz0+hoMH2ilXsJ6i1Bg+vvlbEjdQ9iz/vevhPRDRnkXRbjnkQZ0Bb4hLXR/PrDbPRN
HGgSPFc2jUiOMqyyaju8Ynk/DhBmiVrUvSoEklh6nqKVmTRUC32vxkOB0v/MpuH2YpLHdugXrXC1
bOTplp1QdKxwttMD8et5engV5RTvsYcJVMgQjTVSSsoxylzMQ1IP4lfQJYYCR/YGHSUixejYUerA
DDZkk5c/CXhgU72a3+/AUuFoqZHlP5kmv45V0uB+FchmNou1LGTAHQ/rvwCaZtUpdF08HnQNM6OE
ouPSnZJspWwcEyGlxu3M9uBpS56iumAsvv1/KNDtMwqFL7WyKBPSDtXDb7K0A4azkfHjttdeBNhr
T8RlQPqpn53L53fJlzXn2bw0+fnjMfMk4wbiEZJEBt0RVr7ioW8wlUFOvyqYVL3YIa3/a9oM+UgQ
vQuRSIMLcnqfkgMrSCLQicJoUYAT8zCdw97tSwpCBf/jv4hL2wtyMTVJK3ZSIbKQ3NW8OIoMW342
pvqBAlutcS9LYpovBiS79+PxtCXJSWX8v1JaVNYWSTMJPQhNXd3bTYnZfH+q+4mF6o0yXQ718QK/
BSc86/feejazqFqRL79HUuydawSeJswyj0nC0mla/lmFXmb90+PGT8hpD/O6Qqsb6Cj6k78vuB2g
ySGBd8zmS0ccScnjRXnLundDXf8qysmqvLJ/uY+mOVNsitE+X2MYPS8Hnoc2ITD6mFPsfw88efJs
6tnUOpuVoDB7zwEI7lMxlIIhd6qp7KwKi7+F2TbDJB4taszyEPZ17r8Fdef6bmqySePd2PWEENHC
yWeNx4NzQeCn+XurRpEqJoh4l5U4jq2SUHfcTNDYwdGDx5IUp2Vc1WyllSU2+T/zkIBwi4vhjM/m
nmna7rvFYocYyHzuKK4nUIHy0TdvBx4eoW6/zw39cwLyp2/ADGGz740FJDYyWAMMJx51FQn+XxVX
kzTfy7/3g/bb0KJnlhES2rkyu9dTy3zx+QshIkddaLW9WWOF8Qg32yVmgIxoD24y+jm+C9blpume
8FGHTk/dChD5dIMyLbllQGiN5LS86UpGNliLaQI+MWZm3jw72Fttqq1yF64N87O91v1FsF040SOs
Z2kL/9OhnNz6AAOLNcYE6QLB7wWWtLwK9tbvADIU7mUEcFWW+0SOY/yUYgv6QFRcJf3E8v/rdvvg
JeHUkFDpBiRy2buhnCbDWtob97t/e1DgiXhAJ5JAyLcyRa3KNEB5kk4GOJWxTlJZvTs9qMA9x8Cm
QX6nthaOZFHLei/Mgfx2DqFAxn4vJfLNIt3SBO8ft9i2gl/o8n3CewKKIvEBuqQxiuEM6yt0Y/n7
rB4LJGDvf86egm7yDT3tWD4GsqA7ESPMM1xUSOqfalLySM48WP2yFU0mlN50/czv9W/R3/QGbXqV
Doxf8RxwcTZaKKyodOMS3Uho8G+FOvK7mizVNOtAVAX6t5Isp6qVs/RrJLRUq7tY5A5ThdOJ8Blo
1gxGBMO0iBfSwx5vpGaI3mEBI5eVyVubB8mqCWP/SQRSWXCY1nmiRsZrA8zx2q6FJCCzYVjRpO9b
u+182yHnvpPF8xM3duP3D1wik9Pf/zx5/on/E/A3DfTS3TLsStlsSy6pYBMtuj3H33h2v/jT99oY
nXu0y5Cfuapg9Zhc+OhBld42wE/JgS3NBP9++MIiRaq9wdyMSjdUIJ4kpaXxK+rWMIpHftOqrRBu
rdf5EGp3x/qhcHQipZSM7Xu3Vw4im8vH5XHIUdls9sgtv0YGfINnFVNa7M1vfixZHQTW2r5AjfXH
+zKyI35cp7Uthx51MkB8TEMZGg9TCeSNShV4If4vMr7v5KnY2QZiCwx3nmM5xzT7e057buY/uEjQ
6AUla3w9/67lLPp0UiRC4yJZwGw0ysOKWnMVPY+pP0AFUoKUmqE3IWQE+D7hiFmOUZWNAwqlxhHR
UVSoQ4qXZR7vPKuZ2xv2O8LB7LegNTHT78WpDUSKVa9ScKmhiwZZEFMcdhRJAH8z2G2yuEuXwd5D
GE7yHT4ex/Bb5ZRtUXJwWHcwMs7jUMc2/4BCdsSnfXDYXdIRAQ/jQ9ie0OySI74KQ8YZdzAcqXav
QHeIWDUxn86+hjqv+jZlgVne+gXfGcCQthw1MgBNuCntwZZKqmYmFz2fCWT6R1Wecyf0en8c+t0D
BFGTniKOMbXZb9t6XDAfb0xk9JPcur/Qpyumg35ZBg7u9yvuINklDNeGmlIylAn3GGK3pplhZrJz
38AHQaAAtr1cau9Sp+tu3geuiB+IeC1ys0FOg+PotUpInw+c2NBcupLd6xiGf/nRauAzVJ56ai2w
cf7ZS23s6V+dSWrHmBwoFr/XnLKKYPG16lyrbMkN3i/5sdPwj0EZj/xDTlp53Yv65Xyidyoym1Ab
cBIUE83vQO1q0gqEuEvPVD0PtVZYGOI37lYcT35F6hkdgvPDt3fTIntvdmDeVE3V9Jzoapp793m2
8EzdMa2RZ0OXf6TA765IWtZE2uf20FEiaBzXTIh5ihQ4LGxwYeMmwuHRZ/6RfnYWsOzdIGBCAskb
+cLN4AQI0s+1KcRtwUqCmbtqVOKoLrjKr8Bb4IcHxpLIH24W0L1GbzzgCukGc/AJOpMRQikkn3bZ
W3dPT+AIQHsqdsWQzXydn6VTdGqhmtWKL6412bYjrZG7uodttKGSPgl7H1jWanRqNRKbJmkwLtR0
MrS3B7vNwtPrNMx25ag6PjG2MFB6FcTaDdWFNwE2mwnLihkOrzJi2LpJXqyvVO2wt2y0w6kJkW7P
2dbPYduuvL7H6ssIggUx1CRfBRp5RWQwza2aG8H4WTQ6yv85E6mwIVuXUg3NQanSl03wU/XebJto
B9YoHCUR2cv9DeFCzI3CtWMra+HlvoP0WpRV8f43Pm+1I5wFyHem3WmE0E9X+7qGyhB9gvvuXg60
5sB59ISBh8P4M9Bg2gjy76fkh1c+gaOC9wUziFqhf//POd2txh/+fTNxLw9ljWrMmkSLcARkFiOu
nScnBY++qDdgz3jmun6W9knFxyrFvIfyPZDmrMao6pgLt9vno2AZ1/EBpwqcKig8sdZp+TNbZvJE
zDf/i2gOOHgIq+70mMXzanTXWZiUjS2VtUqnN86oE8Shi27UATtH2wZP8TOO9CmPyAHSsmAizUTf
cX9c61gH1lLjSPc0YOlxEaT5bD5Lmo8ruXSwVmSd9vIM+Pq/6nfGrp19HcFXty8JXkKtY2u8z3dq
QIy8twaJmHy+tZOBzoGgXXbarPCw4xN0hm11Vo68MrECgKivQiaZD1ifF+xxhhSqR/uDkhmqNGKF
dYo+OC5SDLSzky4pIibSoIBzPnHc6MWNTaGFXst3tdqZ2a3kriEDiZaqBMAtlVFC8ZUqMt2Kea37
ldKVleXB8bRP+L7K4mhkJ4YohshDeX4ern9sbk38bVdfltVYrVP6HMCsR1z4MNOas61i9gpwOIuX
TNvbrS2i4LBzKga8TnRgl2+32RIb0UuT+VwxykwnlhlcBnh4J2Wha1MLZPmO/0lD40yiMV8PQKSm
z/xeSi0JARAg4QmaHdr1LPbPccIe1nKwc+J30sNHTso4MjWNlHgqlSGXRBriYIZHx5Gfvwbr8pXL
ESNE2pZQcwc//7FXjHlA1FQhOQUOlgqu1EVSDwZ7KYEXouIGaxUhz7D4ew7axBFZLwQAwbJSJAEg
CAC/0WODox2T8D+A0CyYnOWrUNnnKcBk85u35bTHgmtuEvzd3OWBbpppNB/HuSr1FJYK+uyACMiX
HbXa2lKYHNLjhhm3koWqoLvPHODCR7syHTqOmZrFftLwxd3tt1sCCFY17GJvKezlq/2bOWGDbLvv
dTC2kZnihuDtAhpJZsB8t7OrM1kAGMOeVVij7eIhEsT/jPMjXzK62j6aAU0oK7rs7KPoG+Umit7b
moifATqjqus9teA2fUcBTHkgc5E5mF0a2ks4RZ8drDUSGmpVYE8fugv9UK2Huf4bNkg518X58k/Z
EX6x1h7UMHFA2QYhU8P5UnuMtog3oVR+C0wYUcwK/+4m9Ms+AKM4U+x/I/fwdkW2W6tN5ZNiM6US
PftiUAFCfyGkKoPgipDj8Tl/Jh/J4wxeBDcJsUv5FJKoutU2Ua+cQqDMWnK6ypfztwXgcA9NUlDq
8erw2xu7OECnPANLFfG1VhfTVAZud3mjZ7DAe/Tuw7kHTFF3NXHVT+FVMw5U382BEqDFr0GS6IRX
DD2FOlky9nu0OThkTVaNTz0b6PZ5SXbGu9o4YnG1CUw4fzR2nCdGyFYxcGSr/z3dO+ZBJT1qZuT9
cEonPKLKx3dhnUzXC9P5oOFlzLjs9xmEPwGh8RLNTUtJpGt3b7kT3YbEVK0zhb0NMl65f2ex3JKm
+fwHZN5Rnw2W5TXKQH1uAyRGWgGk4ZQbucRnX/o3DULPt54THW3AUyWjPWqAzASdO9FMfIcFX8Sh
uxviDULej4gD37DEfSsSqZQ5glNNWQ494t3+H96sB9jEzL0ei16dRZGZ1Zr4OWOV7HdXlO9MJk/6
pE/xBYMjRGhs38yffMFDTJ57qW2PUxg9OPiZf+oqc5R4lHimS93+TSugzy5rQD+LRdXD1Xh6t0W7
LL7UnBByGzDTpoIJPVtTErIdHVAuP//3SVdpD6fCcYy5rWjP6CakoAJVKKgs0cYrA80+EcM12Efy
tw9SzYW2M0vwDdaDDAoT+PXWPcBpDDg0RD5BI1IYk2dqFGSJsdGxZe8GRxDB6ksSFY5KX2PsCfbq
74itCqF2ByjKjFIlmp+16mp6m0338hk7WrY02K/VCtjN1jJMkAv4uF91FSCX6TuL6cFEsPqKBOEn
qFu8LzkcHn3Xi4PX6E/izSPihxuc9ykdKflbu9UrOEh1WXXuv4Mo4o8hqNUF9eXqfwnuYMpbEHyQ
gp6YucelHxAjuBaGxlMqe7tAqjTWBoIU7AePzOZgASAjZqm5Ea7x+qauFo2AHJqsAHEMkXsx7HhK
RBoLS1kKDeSyqhMs/9dyEaNKsydX/5nm1VBdPEA4C07Z/lKGk1gK1NpdSZFn2E28qbbcMFBWaMHe
C9Iasfhg9A1yk1D0sOUe7jlKd1igQCgdFpIX7kwjVSajMj9OWgdC88eVqhiJiYuSFxfSwK/WdBQJ
r5JuFvnMtuKAt9a5f+nWsOihjg2nGjGo13/YTCo7zBweEu4HMBbGxAiW6riY3S3+uJuCGTtyISBT
ziA5R3HlhuIUypvLCN4CxBuRMD8mkjmdw4PXm8aqp2OEwL9PE1oIqSTRUAIrAInEzUWBt3MNg0ji
TXGdaj+i6ini+aHkGJgahDG7E4KTkHVcspczOO8H+fIRVhryPhoFt5xgDsltAPnkVNIT6fy4szGX
OCqGDRoGWWbVa/jIaNPagsnKwR9WDfPVrwj2+2qBX/swe8jEpamo2J6qdZ4SLomTCT2nzxAKDp9l
eecWDGcNarRiLtK/i1DTsgylOUF6UvPlmL2tzsvBrW5kFzeW1VcC9maGfj7BeGXLnHwgylouZddd
Zf035J4wCxnJbxhmg62ih4hwU7qCZaGughxXm8ipflJLcgyEteq5ZE/o86l1o3qef+oeotiji3Vl
eDhmOXWp0E2k8Hu5mY/27DgxU0V9fp/cOlniUZW8f+hEAe7ZKo3Uep9DLDDpgVTAMEiUpU6MYKIc
8oaHZOJr4rZl0gQ0PZS7+PtYsq3y4EQUVxPHN3O0GHbnk7V7YW+AYYJedaz2gpyctKKcs06ARxQs
0HzHxZl/boTsocdSqJqBuFCn/x5YJXNnF4qSai+Gm0OW0D9t9PypQXhBDr8Yqp+RRk7G/65Zr5Mp
+9qcmAP3nBtlgvA5qCvY0wv6nLZsekOmbQYT82nWDAFyELFDZOFbIF+Wm6CDO8FFq7exOk+BnPlu
QIf/8yLMbFsYqd4S9+WRq73UwJ+z+xjGU5pC/y+JMzdsgNBERoROhAY6iP7FTlVEyLzS1HZ1Giut
NUCqHMoHL7Oy0KWnW4j7IpA6hwUfI/Pm44P6z6MFcYGHgRbza8OnAv6eVEue4fTbrNLzU8ArN0OJ
1/fLRtMDDL0qdm/CcZcn79VpStK+Tn9fCZKoVly+26Yy2WE+kcdaJ8opuEI6Fne8/IGi+7K2PsQc
0eVOvtAWqsdVeyXETXxMGPyZ8JphwfbMetzFUPWdBjxvWvPWRD7UEXC5H+MYMx97RzqnUYGDC7pn
uLn8AaSlLoMhQWatUMzOWhncjrmbxI5Rlgyw+7JxVJbTXuRgYCJyh5uCf2rquvd30/e6cDP+YzbX
PsDHn059vFUA4NT/79iHAPxQclkqrpDZBXZfHMauYxJlEVVv5M4CQ6y9l6jOJ8YC/R3G8JgBOeXs
Jq8oIU0Gcklg/4EtDKT8kDLJtcigE6K1NmjFAZWuV0i46W0jVoK286PEf6/ykyzVjf+kCoMc5Jm/
M2Jwj5Z68foHPjV9gA0h3Np4XkK6JM5skhyEjEVxP46gYNShbw5JF5UG6hACT5835zGhkllRDWMs
qX0zIu604deIhhCpm1fAxXoWhKmLoTXBeB4brKGfQ80+RocnHTGTyZyhNCAEmuKgS0xCaWCQILOa
cSe2XU6S5RgPEkCSUbmq3cm5ZLeyIStYepTRp/i+4j4p/aA5DIVj72msq+ckdaUc8Cs8ohstZdhp
1OB/NFc2+iq/vieHkCqf9Juj160AKsExJAX3v4fIx3f0qi6HM2pO7xooAad1VCwUexBBLduf0cQK
k9getgugqY5mBl79er5XlFLIc3FsiNUa6Q6wC6OX5VcjumLwVoWHScYAVYH/uQoLlBszzIhHZTYY
nbbPU639n7ELmh5zygdIyIN9RCfXhp2Ziov+GloeVMMveEadiruOOigmXGpgrQT8ZnA4NSDMbvky
gOJeOV4FggoNw8aBWQg+LAixrLzzqDn+MKu3JNE1yBbixkBqvcXhwIodB7hlFlh58PDZW5L1HiNI
V+W1eeXEjAt0KQKR6GfuygPc4KPH5e0aUaZDenBAC9vVokeE9VMTN1z5IOQLsk7Xc4NYmQ/wTWSw
TT2hl5Zvb19VvHzLEIu73PqQbT3fARGAZqnGQiwaJfJl74jlBO0xE3OxYwmpOBuTnxggcXm3ZnDp
b3/6u42fET/axKDJuDRtHE/YAJXwT0GGzBKqLy/niQ5aooVqmr/hzkOcygB2ZGio1rc/sEIG0Cdu
aN3kwAq6y/i/aeatlVobcCupzmeev1eAhs2e+NJf8bTB9PzWheZXTpze7bsndOTEePl/rt7cXQKF
g8BCPr8MXnK2ddGTfPF4Df1qkrq9F/wgK9HbVk9CgJfh680AA3L2DfnPTP3CVAb3WNBkmWhBY3iF
9AtbhE4kZzoPn7gkzBgqBET+jhylFBpsmx7pE9IhzNyz0Va09clOBdtaLjbuYtjfvnnrcEi03yFq
VLjQnzXG6aIg1K3eNWX18Xbcn+T6aBPv2V43luRIMvVkBM/cDWMKZqrT6H1ybPW/Qy3mfCMQ9Lbm
tg/25OQ/bMStoJEOcC4mSHUK/4bnK8H8D1x8cn1Q7hQHaXnRZqP9tusSnMpBHdrP6DFY0oi3/DEY
cwaNCWJGg5mSP1fFThgGQ5/EyjLY2cM1II8Tl3Yl7buD0trT0qL25QMNG0vtcXhBveSily8BKDD+
QKs3+X2LC+KtsB0AxidUym2kvuViWLPg5+namw8N0qUdoi0pUS7lDACrItd7U6xAsrIP84QzdNU1
tsR7lkDFmFkb4Clk92Up1+WhKxnZym3lpHrqDZHjKw5/9wPKob4mAf0ePSVfzVC0bjG0PkDN14Hz
3HHi4all1S6whrPAk8rxkiRatcLcryhiQyuNZlXMhmnaoIp93h5E3SwgUMYNLbe7mOvNkb6Z3zJg
2zKg7Sffyh2SvaaHznzSFDJTRvDxZCC+DAUqBjgZYo8NxbrbC1Y9B76O3KlmdxL61ZkUWthLEdPd
x8c1s1daNQUdmPLKdtdLRKuQM4/FffZIo+4jGo1JB1LrFJR4yet4mvKW1g+6gDBBQ0rD2g77KHzA
aFqUbZbliq+Dkj1ERjhfrJ7g+UUdalxHTUxAYWpWxMGHO/bHByqftCLnC8Lu7WnPo9o3fuPxoY3j
EOUbVV98dCLh7YPvrYUIzMsfz0G7BuBdlL/wxrUrOPV8ZwIamxHdYmfi5eJzQ6ntXVM1gqELwpep
WppeHro2HmgoIqenwcBbMHVJN+3qu3ZyFxWUlvRP3x8WYY9N4Yf4Um26xyoROlWzHCwMdOV0ryvW
K48qd8pi9lFIJQEhXlswk8fEWdox7BYwmtJeNAMeHCgkq0wf+mG8DtedNNxIywX8/XWCf4WPIe4x
HRZzTI6n1MIYbzyrj2V+5w5eMsXgKJGziB8PagWyi8twfD6qe8dZWgbAVwN/gaFL5IzcdeTH3vPI
vGL9j8h6bAvT0hK7cEfwjoQvcT3DtKW6ooN4i5UmvFntTfMNUzt+nFFI4I5WohChuPnRDw+NFutc
6H/Ut0fKFhXMdRHYQUkf9HWgaSam7Gx01F8kaBQv+6+YqeDnmEv17T5IIpL1IPnmBdhnhYkFktbB
pWsv2lQdD80j6SpuNl+9Qf/W2NOkCaP5RhIGQqOoTlbgmDM2wEV8OykDFvwqybzf1UdNTUxQAJJ4
AegVAC/cNA9Lo+eZcA8lfmnO7iBaKHH/nyoXb1XFODnGezAKl98GbAjbKAv5RhfBFZVijl4cBI3/
am/b9LueFZF0GePC5vVGy++P6KRwodap4+YUh9V/Q30yUU6Y563cyITVwB9JJm/MeY3EpTaDnZsT
zS7Kqxkn76QwRpwYhF8h/OtUSoJwlUr73CzO9vK9x5vcW97z2l9lOpvrceXpDh9jfiSUTa9mDFHl
htJNm4sT4fk7eDAWk99boKolk30kUI5gSKpXE6LkCkRJKeXwTGDbr9pl1XXwMwdHjEonmprM4Vpf
a53RgmcaUx69wswcMczSUD1QsfHR7gGOuH6u2C1FyHFK+5bp6nneva/9T7Duu785HmsLO/P4s9Tn
HkCOQNPUUigMQ6aahMePapqhMnN9P2P9NAvtohrFY/Ro9Rf3U2YkepB9CASFWobO8Iao0bczRua6
XhNJbEps1967WM9LeKhrFthwpldvPHfY4w6WiQD35/PcdehjI6tQUZYcIP/mlfVz+ifaqtMddAa3
6ZjPLSjgjTASmzCej9pYigNkUnB9nwPlll9k81rpdWg9LC0mmoo+WymTyJDceyPFaJSd0sk8IJWE
aT/ARs3dYkzVeu09ZPMOsLDSQTMDvyCGAgoe092Wd9qHupsIxdhJF5Kbx+F1FW85eEtDGMKK4NoL
Me5ajcRG6dRxAtJlSgE/v+pByFfLcdiRMOIQdbxRJ0ZJjmZ63DeSMBNzOK2+ffZ1FCf1AYMm3F86
QDzl0QyQ5i6Hud7PXSVi4oX2GKGA7DWVVuFSwYYLlPz4118KjSVUG6ihNjKrJzLEWVu4irLCHJ3C
t0RSqUUc1L8Ygc/UR2XvE0bR8poTHA+aiHpeaC/mmSb9v/wRhRoUD5YlKxOF7DUjlbA275FDLuTU
PebjOhfRW/tw4o3AvAH2At5VFlbtueNZrMY//g+e1V6270f9fP+1yFLSYdVFfUp+AupY1mjilpMx
MJ2twsNQyqtAljqa7FArcG+pbLRp/AZI+eML3odFZCeALc3yMdg0SKCsy8/lfD5T7TxrbJQg+4vB
/soAt9duK4MS2ybUSHmojm4uz6vlLkI+P/9OS4ZSFF4qFODGPJhQoZSx4sdoW/IPF45lY4GjTxVG
GaRPzOiNZ2ctgdZtE8d9ksRCHu5PgJRIFC3wbizI+kCvps5JBCPHiqn3LRwgqSYbZLDxvrznwyoD
IGS0kohFP780I+SuCpfweENuux9Nn5Sikp4xEHKm8UZGBuxMgy5d0Nr9IJ/rKfJkQC6NmWLIz7Kb
5t8QQhmbG0AxuDX/ADkPMxgXkVwlTeS4Rj6gmZanzX1bn3Yrc460cgVFMte6qeaCbLJO/rTOrkVU
L3rFKitxV6Q+julD6r92mkwJBrPudAtStt4TV6HZuiH7oOlRMwAG9wuHyooeIOco1G73Lt30Giy4
JWZ3H4Z/sSHEbla7D/9VxTrCtqMgdEHLlS0DuVsj9nEFEyk2Mj3bei2u7mywhoUeMn3a8Ju3cayy
yClbhWZqRpRiNM0tB+Nash67JFHYAAHf58P0NNm9oOuNNJyKiEAcC+AJX4jhLPabgeqXqbwaPo4a
Q0dt3thsKgW98GbHhNrBydSMHZwwApssoyvw6BVbdYHSQ5HRBwTN1MH7gdlnLZEDw8CmRM4i5hC6
NWxBFWuHtU5fNEuKAtSHsNctwvArj1zFUo5gih5gdw+JShXhlvJ9H1rSj+7c+Mq/vu+AahYPXlib
QKsO+ypVmPxkU1Z2D1GZ8MHBiKSuq5gSixOa4iZVP1TrY8L9/Zc76wgRCEcTSfvvj+KXgZiSoCoN
ACjwT/I3lM0VWE89ERybYiCsIyV5BBeEOncehu85CStAS9c9KlIX7yy9ANbdtO6xqaaeM8PLNC5w
pharboGpORY37Fnj+tsdM1nnN7c5PcHS1QZQ7MxKT4fyZsF0WvuzeUTMMQPFFv0+8DdJF/3A2uv4
eK7sAfc1yWOH0QeqzWNvLrVY+OGRMfZBzT5MwL/R2r9g/8931RbsbuPNPflRUxheaRa3PhXHHDf7
nDefFCPFtGfRE8Q4LyAh3mj+2X0n2xmPVK4neI2wMJagNQquL/dRFSgK4QrMWbjlZMYWffQRbJOS
UB54qVdUdudxSy2MguV88Yz/yQ0g1X6QJslX4RufTHjXkRKyPOof+EFywpLorfbQ0IJnmQsCDV5M
WGlbExaLb3PtAf2w5eTiAWmmdvHezNZ1fXxH8yelegftyVJLs1JhA1pj/Tm2YZwNiW/4EzjneZFL
LMEeo5k07vK8CxB9c9cxFePkz310hdMV//ZmlAqVrQHLweB4CX7vPkwb17oNZz9l4aS+AcIPLSKT
0XfscHstbcrtL8eOTyTkcu1HhZlPpCQTAN6fAMfc3vN3Td3uLPMxmvcfAHv0xLOQdN/LEjeJYi05
qAHEXPti63UsylWvz2wIhZCFA4H0HTHWbVvJttBlMPQ7g5/orjee6kCjSumnEzMnb2lNePKFGjah
dKKwWMYBkYU3Xbp/vxiHGs8L96zqgGY15hvWqkkRvplmoNVE9xgppPYVqD6r6Oro8AKw54H91OeU
o6j5UbyTocF6+OtedpzxAPLTZ5MsPfHedeGGqqH3iANLdgYXLMtz6fHMPRKLUvhYgmboZVjl78aS
EavkBaYnslV94nUCJkUzArzxaKEfU2z33FBCgCgVFZylduyU0tEkIZ+en2sQG/afQSaLEc43rXd1
G+rRk5af33USoFhSnyAGVn9oW9kyrI1U9M6s90njBKdAYS/CevJDB8o2gYeAQ0HLP4QRoaGKWBPW
MdozvUAtCDw8PXVEfdGfVjErXrOy8Ie7zMODRy1RqJPSwyYrkbE2c3vVguRYJ9PHt8YBzaAvEywB
EPtpNbrJTHSYnDsADpmb1BveL1tHrEWyDW8oPdcbZC1BlEPYU6M2PC4x0edCCuy08EOXTOk1u7ft
3Tiqd0kcf37SL7ZKGHUjBYlKUf58Iw43TfVVmVpigPuk0gJLyPvg+TcxT707GCNKQfOnNkgJq2BT
yfWUbkby12GxOKe+OVcir3KJL0yzgd3NwnLVoq/vadRVXv9DRhXBjMrUc/vAJpItv6oC764CDF+y
jFfV5FjNsyb5XgfnqlM2wTT8UItbihdE+3BBpdGPQ6gQ5Jhvgf/iisPRF6vyZ6e3eTCqttRCStOe
amnc+8Pudt5aDM3pQhkH58spT8psampVwp49GvqyHlPr37XNbHIIVtliXnCwnhuVpQuliCzurkgA
GoNSGBcX6y0Mok6LhkIAQcxfULVeFl8aU0habRO18TNN92a3XUqo1kCvfrEiMhsFjl/qcs4Q1eoQ
lWE1k5x1ph9yOImWoJcCweoRIYhLbkqZ7u9hQ4Zcy/5rDxfW6ZqssSp+kqKeQX7GN6ghUDdbdZ71
0ch0MB1reH/EyaE05es62riV4dx6M7E1IOAKbJhR1TAWM2jCFYUP8dkLfBi5PFCONejUdoZt3uza
kwvgOeJ6WilnhV3lv90hFbi9os0mOSJCn0FNbD2y5K/RRYn8z8RNfrfQqbNi2cDS1ZcdO0HCoztu
AcFUiKtnBBFrVylalrsfFQnMMhM31M8MdnUtORuDVt9QJPv5cF1PoI5mZU3YMoBvkjg2YKc+qZ8j
5sIIwx8SongIDvnJWzXwZrLR1WDHE2M52VKJl6T5qGFAWzoO9iXpW9LHdVBdxmsMf9cSSpWcVfoS
6Xe1wobR5+ufLjxHGL2K8OKgVEpyhfh7X/dh0ctr0V9nWuFD9bZ4lxAcl8fK+2pFTET4KH+On6de
amEj6+or0PZcZKqj1/YExW9vnD6zxyh3hijIyCVekl5UJC44YLJcVZ/nEfCVy6+59SVfecKjHEtA
xR5QHZYTXvEDQbVg7luvAfs1EnvJ/chVKLFH4Iq6f/NB/HKxkEbOpMjVik7OXet/7ZO7rb8nW5EL
4IkauiYouJmCs7pOsv/OWkwjGB47Wi3xmTiUQ3gPUKBqCEy6L6ymvKP4BSryPLC+yUToDHOWxfnA
PeXNPA4CRwG9Qe/wwvvveIZ4LwjotBLqJQbucb0F33eINtryLQQwtiXR/Kgdv3isf1kZHrT1+5ej
RCsgTyIR603JtKA2nSN0C/pgKtck9j8gCqdeY0Mw7fWXLzoEZBt7CREzTXoqJxZeOuh3ztkNastI
dwy5ba7b7umjdr9yPOEbkpzYmiy/9UXizlOr+64Gs0Dtnn6yC8LhcuD1jWBDK86PlQ/cMHrGM89X
Sn4ofmUzcBYsmSL5oNix0C24o2IYxZDuElQ8aEYZNopU3TQq+k/z3VGPcfr40EIWot2otkQf66eD
pGtxTZvHvsgRwMVBrLV8ErNdhNpRaYrnRnn4Aj4aGXYwmm3tWUg/4odgV1fJCDBW9UGTF+tdxqEL
8l+9mzocQvlG8RVSPMODD1ZxY5KRqgv4FBqt91ooTrqXohD9kxBTowxaXbLVddcR0cPOx1hEvmmT
1O0vJ1OwVx8ATDVICWhC198BUQQq27PlTLT9rXDzLWoOQSTM4g4zVO9QUNfKJrqjmeZbqg6+gvx/
ccHqUPpCUGpl9pxOztLo68DnmcJOfe+8W0AGGX++jGEw6CNxWQeUBqIB8x5xQY2gIW5/pbSQZv0U
fTZw+Jv/V1D/mRHR7/ewdt7i9LHqXgPSPDh+WJ33Y+Ov1CAYxe5RlNmY1BSLloo7CjDexIQyYBam
q19gPeAwToFlf0ytw3HkilNqu6WF6QdCleMk68vaQs0IKG71IZI1IUTxX2YQ5c4ECWf3zUFhHfXI
OE1WODAUNJNJaOkJUb3Rau+eq6Wl7msRL+0+KcQula5wp07+6yQX5spFqqafdAPfw2+ggDAEKEN4
vC5SS5jW2EmaalzbN/rQtTQASsMRzOdWe8ofNwed/wKCNsLCqV5sbimgQEIFpSBWD6odS6l7EupL
ZmK/SrR5vp8NymC+zflYVc/BI1HU8PHC7Dl/KrhLVpjqF7GK1AJJdPkwggl3LoNroysWiqCaiqhF
ThwQbS2VTxZAmNZ6cpj495f86xJ9l8yLtQeE1qjMqPDtnxJLYDQLXwL2CpwdDlNDsfBYl/bI9Tmy
lEbQv5UmcunVuSJW0kLqcYVwRqWfEoKUTiRdkDv6ZYoekwTc72tqiMKoJswsXycyYP55LG5QkAxh
/4DSiBGdNGpi5Ej80LrNHaeybWcSXQoroUnRZzKfHJFsoA+UzZwj/ki5nSeBL1xPWy0hKetF9Z0S
X51+8RsEEt1gDv/zF7EMRKiRCRrHvc9BHnsLJ2CcNk3dze7/cYuWGReybtcIbaYHAsxV3uiJ98Lj
sDEn2I7vY4t1HW/glcFcAkorVzHkkGL5iJv3ijo3gWQD64fo6UeDQT0YdxVfyYbtl4soy6PG96oK
TUxrfOwr1xi1IdVgz6BS//jDhln3wRVqIauwRqgrS4/nL5p8Y/5OUj093zxrES2ZBQ8VRoFzeMzG
dmaHeKvTgdKmUuUP3+dzscCsIPmUJHpRgmza2l41QM/8VScQ8t0qR1gzXZRvXKHejWq/dlhfxaE/
j1zOGFGMPvR+UgQBnukH/Co/6dNlsSq19uk41qWNTntc+zz/05TBaUNARqlZ5tTyJCzffvBOStyH
GUACQjZdy52oDGT9HsDHvF6mv9ob6Ituzl4A5sVehXkKycJdnu75vv17hW6RgOghpMMafR6sBWc7
hQSATkVvb5pfKqwvtTXSaYhWCXk3Yt6imLRpVE+Mx7xnX0/M7tcWY/4n19XG8FkcLrEWPtkxoBwT
m9zUYjlxMUGTYBHcFB/OpfPojo7sziabmC8uOSZSp+GuYpo7+HIyNaaXH2xVnZXxFP+u3m/XoH9m
0Nc3c3GdmUT9B9sYyiuc1rbQ2pRQBSHbDCICnGbjJjm2ZAQ5sLlb8UIznnkWRKJYyU8GGZBZJvhn
GhmKlUCg4Av5y2SmKqQ7pBMpEZY7p9RlaM2ngV0EY1T5RFkgu9MWEpgF8YgG0+d1e7QZwlVJysGQ
AS5n8MvCZc1Ru0PC6uRHgZiBf3Fc0C9WrRMZTwmdn4FuwIBmF1wDLZ2cdnrGbIh7+ZLR9i34GUKc
wbOUQyk2xegl344DE7sVi8D2Pb+rbAVkLkneuYyigaHvbCubSbmKUO8vTLIVnuX7K7iP4G65NE8m
2ys5t+2bc8seh+W4+ulJVZWnswPvapTeMrGaKUMB5lrIOcu2VJxjXFzQ4fccQ3LzfZQPgMzjzNzn
F44y1GxZBLqN8cywdswIm4W0YNs2Tj7DYJJDHDd2BnqRqb/7rCGtSmhBwcVM+kFG34NY58X2XnIs
Kf2kQwtOT7DU5h3SgGwJ9hkbQhK/bYGULthdGOxBRKpLyE+ZpXytwcZJMa6nToo9rhXpIZ6M71Lv
DvMCyeLPDypxIvali42Hte76SlKPHyjtxO5LXyNF6b9GF0db2WBX4P0MsXpTyze/qgWg3j6K8I3h
T03iWF4ZHQtlS4UA4NtRhmvZHDMkJbDzbwWJpSkX/1tk7HVqqDI/+52yPa0mcfnj0z9PdIQy7DRS
pB8FyfFdqwFO1gFPAaGMEogPQ7XvsL2a8SbgPO6yrjSz1MzkWgKFDBAT9L/pyr6IFOTOtTHblydY
xhMOjJBWni+5bjZ7ZaGyWCYgVCYcwtEgoC9YX0EavdEjPMWDYdIR9iDcv3vGWkeIzX1/TFPoz7gk
6+V1fAnmq9qEhsIGKG5/5bD+xl7nBCRhVe9AM+ntWydlxt/Mlq7IZYL7jJ5eyKWpcFHIeNw62O3/
m1Q371WAHbnPSElhg0eXuBl5WD26cp1Y85dJsqfPLPTL14f5KqjP8qiylv9fRCZ6dIgpDpfxf6uX
wQhgsp1YiajPT+8s5lnlQTrtAScKdiHn6C3cvc1hdZWxGSsD1+BkKnGezNYe/AcvQakun3+84e0O
VioJ0iyuAYOVYm47JKitaZW7R5NrIIF2FVG9sedj59APRfhXVjYBVhYQK/l4Aiuceu/Obej8QQEN
psTdnLP93x6KUvd+N7QTl+E6NvWm4zJr3GvCvHx1CkgzBk2+CpaMWLA23xL2MAj8fHjKFZZNOWcV
xq4bRkGFhnKdaNU41YeSy1mgnzsy/hMLh2XgcsmDc9kSzowajBDZh3971Lyu+ezDAKI6juC4Lsjb
HS7W7M51Z5c+XWTS++CROnAu4RxcIFzkPdFvMx81KOSPJWcpEANnNBWXnQGgB976EiskipjK3KdM
VTAdpZqZqlc4tHV2GzDANPTfBYoC7sCb43iYh+YpVONfig375qVwoMOp8ICEf+QhtwxLMIexc8Ek
ghbbJTtY0em5iCQtm4ya5IzDsN0E4Y9XnuW+AnsQUYzsUz4/GfrlCRjOIgLNvqBQ8MeCOHkgOUNW
zpchV7DyawjkFUz5XzxGPi/pcNtNGJpOR07OMqcAVjpOlE65LNA/LnVrZ/aWO3MHPxYoKEDdQVzE
qSq4412iRmOH9KclLJn/kc6gh+8PA/iAWAjtBQc7QZLNAcFPhbOphh4+US+xUplsJRsa5HMQP9a6
UAFZhV9Wx7aYENVaQiNp6wBU2G5Mj7xGwSDrE2hEMUFSG4Yvb7+jM92MqtHXyUy3fB5VEoM8YDba
EiWrl4JTp7u0t8iXQaP7lUyxFwkuxMqawiTKKQP48XOfrCt449MSdy9ju/oisONy62xpB6fPUHrE
SN8q8XT714svt2oqMkb2AePgq2QLr88c62RGkcmsH7MCpDJDLREHSwHHIi1BHGcTYsKo0DOgzbB9
rbZ1dUqIpRghekeOcXJJq0x29DTyVeLUwLdDkEVipeq8cPzttsDM2Hx/SVx3dewARn++gfZKmrvI
W2zy1fYnEkBbFEGqiycoXnDV06+dH7Kp8zK+gIgUz2bdMQHWBZxbDmq1Ht9ktYFeoyJ3zen5FnI+
9bmVeQyX88nUCDpYiMtnXBePLo9yEf3qDX4j3VvIa9plyiCjX29K9cfvwMP072IPzd16BTemRNB0
bxCZxQVTG22dZseiwVlIBe9uMOyl6nI069Y5pXShfly+RiAHjByHRW2MnoM68PXdz5mnOTm1UdIL
UTK9P/86wTTGbatxYuR1PFowt7USDb+mMa3eEK2UQG0rcZwyvkr5HD8DDLTolAWyDoiI0Nu7kJvR
RiFU7K8pYb1WBUlRdg+9jQMx3W/DyMpmqCQIH84tdqDZ2GGuNj3QFKP7L6d0M8mykNLGBAAku99T
gbGvz17Ml4Y/hSwWfWQlIwY3M8gt3DMSNNhPkeKNUQf+f/jqBtwT7IuWXMuluZPUtidJ5Fymxp0M
VqUX9MjJ0m5MTXHIQ15s8oCBL5z3T+VdKd4wggDJPVZIgqZUBSoFN3IZltOECOHOqmMG7CNEJFUr
cqMiApZKl3O4MoYnTrzAxoGyxl4pIDCMDexmXS4ZqkOtT+yVCzWQ3YDtYm02Ai6fFrbHgZToESvU
a8iYZ7eXYuVqWVYUzYh3WKF9a235Cv0VwiOmvcleF/0A3J0fcXZSsOJqAL+l/cgmtwDjbp9G+qO6
zFnimRm9l/phniTDzBMpOMqMXDfOf5HDQh2yJ7QF1veQ/VJ7/rALxLiPUxBI9t/Z0OUUt38v5U4e
fQWkxEbDIty+MOMMNcjdzf6iyPnoIHMVAkuxwtw2awfaJL7qyaKi4hg8lNBXqWrZugZjcCOYyWbT
CS34HJz0vVmj85ZxfGgeghrW4RVWWvWDfTliAOnJMwmHE2yD3dya/avMQGHVT/ljvydCC6eMVY4l
zykifKYFwYZ/5x/WpJadW7UV2QjpAsbz/94IVs1yjREtHaATg6ocTE3X+vw5saW2OTnQ1TgRkfmS
I4yAJ6+3rhkXp/FrDDLTNsQNugnWgvBMi6JrblEVmvKXvyGhzG0gluQIBl4gN0AZEk5+bJmT2TuN
fKwk++3KPY17MpnuqS+Pj0Eobxw77x1qDw065KEMjWo19FrAUtfwAMc4HfgPip9A8HCbHwvOKQNl
P2Gr4LGCTWZID65Jhm8H13Jy9RcUnaZkxlIzr/T5pla4rIYw8sIx/3ZG15sJ1Zlr6FftG+2nRDkv
0k9Jw0oTGPENtbzzV7Wyrxh4Vx+ufVvvi55WD17wHeWKOVSIgqFmr1XC5ExqDvRjRTkC3/0XI0yZ
eK4oRUH0v02Dls24VuJL+78+U6zo7sL1nrhFBFnpZc/XS5RFFK1paOOn1gLRSnHKt8ogu8SIJzyo
hIA27pV5Tl9JxxbUCWRB7TDezxdnWN1YSz2+Bt0LV7D/kP7iZQJduPNzDHqoDbnHEuN5ddo0qzGG
yk1aRsTA+AfxCjl0xjmKpCkpGUEX13h/QeV/YW/OGpmxXARSXTE1wkpxcvjGYnfCBeFDhhFdM93O
iTLP5yxDUU+7xGLshA+GVE0+oYRJm/UodzxERkcJf1wl8W9EeeSyww5W+II1OVGm2zfN0uge04v8
+/A9U2GtPmrBi4WQayHWvq4IHR+UrYKjxwd1iMigzGJDES2iiWnJrVwRdPWmE51EvQ7Oi3ApHlHI
+Gms6Xv0Lc+G94GmVNVjy4CZM9x++w1JRhynIinLlczJIxuOCdTI0AorCw5ntZofHr1FcansV60h
O+EDDD0kwV5mHm6DujNdsZ43szhQz/WFGrzWfETOKGvYzbvzpqVdEqA+A0bjLIk6eaCsr0/wzrS/
srD/uvORaIw4vVcE/KRPUyAeXmMVIr8suVE9J3yk6TMhY68/sr8JI4v5cbQ46W8a8K3OOMzWThnK
wJ29xHx5gXNF8ZANSCiZJEL2E/0uabow8bQCf4F/DEP2MLRcKPWzNd60Pj6VuIR7vSdqntUtG06G
oUxsbPrhU0hBGb3ssTFxJDeNYOkpXVEuf+VRqPDkdbWBYdWZYhjmWpSIJgNdjuITuGmLDx74BnuP
kRbvLyrL7PNKa33lOFEbmeKhneEJZdcQWDex27Scw3wzFvYpMzTUu3XqWiWfj3E5/vswtEGi4rKb
d0qFVTTwyLzYQP7Vu9yA0laGWem73S5uOlyutb4wvAetY+7+1bG2xJHC+5BaJMDu+1f9lNEn9S8Y
wxjTWCxANv0r6M3s85/CcauCqfKaKAb2k3+wP6aPo2/bF+/722Z9qzYehQuxv9tpWJ01PMR89beo
7h8xIEg6/NY46iATL5X4sXRH5ot3ece2WCdMrH1iNcNzca04T3iAaEeltT/hapydUIhE+zK4J8NI
jHQMLtG7tKcLWaToZ+w6cyESjFDQWk1QRVoPxnqG+nQs5BoMznrldhjeQKBbYUpQJaDz1yp2r5G5
SjCAOMqIgJki8Z9g0NOO+OyhY+HlY0ZnJf3jDBdxO3JlMqViKu6n//kLSu/+4ykO1iUyWPmecSnA
WixgL+6dfqbmOnkek6R24eI8+WHmSNffAl5wuWRociosTsFxtG9bX4G83XVfClrcg2sIoFeBi/TU
+KhIPyWuFaBIqDcGa01GcBK0kzFBNZncQRsTQO0SfRvcK/OH2wDFUUQJSCJOrV6uU0FiOA+COcyi
ME5Q64/d6TMyZgUjY3ufdoc4CD6H/4uxVcot6IFIpMKi9h5VnUgi6Ek/otUFpMDKrZLqi1r1qElg
+T4n9MEN6K3U0AAEjeS7zqObfhDhepyK1wV09estep4JY0Dw0zPtPgElvmNu3EWaCjaq1G42dOam
p9YRFiK52mPop/h50fwufndnjkyGzbHgQ8jW8euQQAHmJkCq7RkZm4tSS86duQnMNE13d1fkXwAw
V99SZC2siN+8QO61pTstNoLIzh9dJrQ0tWkfPmcnzre0mZRsf1XsCQ1VZZUeRwAbFyoAAWS6j3s9
h4a3fx7HUT2hh0ThSyS9b/8lr11zSLHn1NfkFFajJl2ScUS18SnrUYvRqZQXe4luDx0vNC+QXpkb
H3AKQyEWRcD6T/kPoOA0+Xm9Ko5S514Wb2XxFqeGFa8G4adzF5kyBJf4qMCRz5OZCjwVsUIkPN+/
+PUe/DQmAuWkyNp6gaJI7h0jGLuzidGMa0A3jtAoobhtMU9d1x6gHQkP7pvdD3QLB/3C19bF+eGu
1K2LjKMZq6xRkNvfMXMpWCGOsC1xFeY4lyz4+0ZzVvakWVbpEZ1SI+Gbg0GYUrF30k5LO+AT8yl0
MqJ1zVB6QlXVljyhJlNBUI3WVn/JLbPToa4Ny82+ev9CzhUW8qdPkXcjBsxuDEshLdVIoadwoyXg
fPYiqXhzkcpmrlBtPtHqh+mOX1yefoFZovbi2vUTxLK6j6DNP9AQ51CjKPKawo60uobi8XSX34vu
6TG5x4hYQZOns3hegQrO1O963+qY+OER2uRgM6Ha91jbBf1NJm781g0UuMYo9dakbfkGS6C7Rorh
BPDXW5SCEi+tAKl5zPLwmrz2adLtEOznjqSQwhrBidjbCZ5hDmHP8dvk3eVJpbjCOVbGCp4QLRRP
P7q1rfkdakhZ5AIY+VgW7rgjqVmLjS8Z33Yg789+vLbsS7ccs6HHMGPUTaa21DiPmudZN1qe1yKL
Gxe3NJOqQ4sWRohKHBzHrYiKbQgjBLUftK7sy1/MojNX5iN0PXIOX0CgXI+Oxv+r8LBfMMZRB7ou
FDgBCXfizxIYCQ/2vEIRSMD+DiCrAGvKHTg0Tfv2q9G/YUNO1pLWYqh1k5SF2fiJK/o4w0j6sUZD
EZUkgv29fiYS8j94tai2ndqHP56tWnxuuw6z5255koWf4Yda66J76qkYsVn+kjgvYeB9ewkAC2ml
ZYbtuTUHK+/CJjCXFWRlS7/pWSw3xUWC0ImEg0UwISLb+bYhgbPkhbIg4pZ6erPWSLqM7fEQ2Miv
P6p7nLjlsb7Rnncri1DCxBOpd4Y9MpyTK5ZgMRaD3/i3hoPsoiRcG3KTwrWN6SbzQe7gYddllxgq
0irn/xGhLep0tKG3XhPfdesJ7rv04ze4bu8BiJP0tnJhOT09Ea6vH6yAiKarIpittiCOF2dFuRj4
WpegxZckSrUD3EWXs6l2lLERHgMo+tXojD9eDcQISnXcS2W1G5J+H/vC4q6ERl/wZzKuxGJBuEEZ
pXTVf05tM27oeS23g2hda/p7bcONPQzKq4Het5AOy9D57C+ULcxmVDML31onjIzOtt1oXyjyUYhb
n53Gt2OXDG5HfvlPD3oBTMBBvloFjh4YEglY6cJxky+dcCqAuIakKkwBFPaagJ3n9SMct9pZvrrB
2MStWUGD/DKvK8uTUgYIOezcA3ljyDtWl8Vc80ll2l4gfUtDnc2OEnihOgEJfd/AZAr8nlB+Enww
L86KJ2iKJQrAF/lwuc+TmWX4HMj+I2iuZo2/7ipfne0rD0ImqHEETxHvIPX2F2RoGuaREy9qWBwh
Kua8gQDqQjP13OxqoGHX530TphYZCWfEiVc4BRkzh17Dc3WBREscUt0pNashewex/GAj5tJPHi9H
BjH25B/qxONp3q1LzaAmIbNhcSZIINSqR83/74e0xY+BmiCu7yLsht9uyPQQKP/Uvl6EavOtpgJV
6tXWKuHM+U5NzNHoxjQbUemKnGfT73V4vqn3vDJvXMgG9ozOxC1ssnHIbZ/Ij/Ti8DRlL33vjAgL
sPbgpAm45RVs1qCHOU6bBOW5vBrRLb2C37EGp9moikVQLt0ZqsmKbY+bB1VTveQk87CjuJwdABLO
r18xw6FrFmP9Egnvtj7PY4ub7K5BrGyxFh1B0ihOPp6D9HQtF9PhlxRtk5fRNpcOkQoj3+6FEQcq
oVb8vbFoSlkJpqtqUT9PKnr8V1FYWNHJhPw0ur6Q39v03Qu1rVPPrOUnr8s1A5i16VvrQluVpuvI
oivoM9BoMOXtdsDzYMhEDqDSE1dtBDyZTOSIcZvnuOsMFx5OhlxO0fjL69BfaO/x3/EcQjSNdi8m
3b8043Y3ZD55mRsysLZMxDwg4+q6yZuN1+vpTpjXVcy2noLVaVkI3i96Tjy6B09ubhA589tp3Ti/
Fva1keqxokUBS2EW+fFqng1Aahtt99m+M1ZlHCeG/GkP4u5+IC6KjCwAjJqjOoDCbpC91GTqvQLe
AZ386mgls3+Oeezm3nA6CaM0dHseeF1bH6JrE6DegI4acNREfKLo+EwUwcJe4f5ovYDaOHzJmNH2
w1VtVPVgFqpvHB9d8y0WvH6j3CNVZR8jQsJPFimVLJ4vxtsJswaBH7CPIrWd99FeX6vir1ut/nOn
GpxU248K7lgDFpSjdV5+X4VjHCaJWWhhhDcyNFxFVb9f4vIJA79hZt7p1qxljqK9HO3GTiLW+FE1
QK2fFXiYnCafnHwQbWfTlniFNR4sHQ/ZbZTThR3ESMuguyAjaiemOqW5dC1jvPKuO4kWTKvipSCO
iyLPC0kNZgMrty/WjXzkJZbfBV1iQ5QPJPE9rAcaSpUAdsdiDBP1qqIzMV+ZBjDRMMq+yl04tdrU
tNHacxHmDykNf4TphA9r1gIWJVpp4BcZevNI9jvtvIr6ilzESeeVi5SIPSohRuhBMWCR/E6kF9Zu
p6iv8T6Sti7icOF5uW09Q61LOv3qlnR9ngIe6pW+MAjQzNc1dKKEFXYTi6fcuqf4jNUdoSWEzTwT
Tdmi9UQJsAH4oGD5e8FKq5GEgEgel+6T6ZllAvF5/E6A30WxMrEtuZ0KU5eiI31KN7504232aNoi
a76VYe7YvNQD9MxljEXYmrVT84LtnPgtty2JFwmHAG8fITYP4D1A8oGsYQ8EgP40GotTrUOyvuep
3bUCGJuirUqnhVWQc6O5RE3NT/kjXErrJMGOQmbL2kdHpRV2aCcH7ufmE1gHrA61ptiBw6iwX6ha
a83CfutdbcBnHLul3TBhd9bp/A6/JcBt2XQTq2+GR9po2mYizBt0aVmv8budoykAAvRvYAJwa45G
AvmRuvxZUjYNBJXy5+KWfd3HorsdHpOLFcDyb5X8iInGW2qQqhRh8uMN8sqKZbANKpcmVfHJnqgh
Z3BIWW+l3v9ts8LPtJGnKzlYsljB896vMUdlPG4zN+dhlNvjAv/px0VlwctkbNAI36s9oWiVvO1r
5TskB31G0p5TpSPGhjhB06Etqtj7t2PhiCBBcPk/1gy4npE+M7eyryQLAf+AGFMudbgPmjCTR5iI
akEr2QMUzhORsq5QuhEjr5Hvdi8EeP/c3MWXd08zZDCEu8PcV76IGLkoM93VkMspplFkTbUnejzr
5sOhbUBgj/gAEHiYSuvIUGjhoaEYiOejAU6Schu5f4moNt4mEVj/PfHhYT7+giXyS9O4SlntrZMF
6K8JCAyxgxmntbHcAYx5L1CgCJcKfckLKHpqEGOk4GoxI89NbkuJcruTSv0SKvwfjQQ4ySESaxC8
Br2m97IRQPgZtHLhRy06D5jnltiGVpRvHEg2MhbG0QA1/hj/yPgtrrl4M4JSEtSQ7VMe9iED7mYn
wGS4Q0ne5dmP3eBgDKm2/mQmNKoSEaXesabudBxtJhHw5oN9p9CSAKZbrHJWV/6NwEzLCQNOPtcG
aAW6R64KmyZVWPjIe5yd3DiZZN6yJGv5mQ3+wwaMy9GaVVbZxhdK+17AQzzPTaOvss/jOu7+W2ju
pFlruFZOHjoAExNH6v6HH/VW0abmQYLSyVfN3LmWyXxslWmXoZFfhDty1CT+UOX8m2QgHpw6WUIu
ZIiiXnP2Gs5rkFfb55GrbO/vjaaV98YFWkHC9WwHYAKRQN1N6NbPjQoIW9cHrIkvD2bgecBk9m4E
ueZXRvRk8BdzLB/67HdYVAvYdVuf8Kv4P4hHooqxfDvkbyE3V+LmbvoDIZ18579Jf6X2REHAylp0
2TlM/QWmeqx9NrXHxabV2CL9YaAfFn1Ub+MuG9aA+9h90acBrW/jUJfRYoMyFWza/8BF9YFY1jIv
To8o4ZA4cr+2ogjKtcFZ4YYqznTo5/KnK8zFVGM7ymA78Cx1b6KkhMC67wCQE70Qfsx8p9lEIHga
j6U/Xjapxp+C82MZSmtXkhtB6c6v0uWkX1zA+jpCMKukmFYccx7XfN8YruWRsy9E4Sb8pqsufeqp
9Sk2PBrc6uj2YaemTwvxnnNfVXWI+nR+AYLR5jlbI/1p1yg3GRG+2344sW9/rc6MM+AyimPcVsly
a1gnAqfY7D6OtNViOe+hTEzARF3ZipCpFhO1AgmGPGnWCXG+x2ITAe4XnxIQhhaAfbatBkFxSpoo
pqtCFO6XcrL/hVRXnXZvpZJEYGA0yUwP3e4n2eYV3T/13cA0dNYNPlQgQcTDmVKaqkh2dNPkILXk
YUwEl6jhwke4pUGVaV3pNh1IG1Qua5rFor0I4UbbdoowI11DXlxwVZoDWhH9I2erO2+MfXAzvN20
WF5PM7sXo89/ix1AXr+yvgP1jzzrVnNjs3AQ3KQYK7ZoIywAP1X5zHmROb3fv5wA3xp8E7JKDaHy
iTCf4oSuP7AzXQrbbCsLGQdhL3r7WEhowpBWoXLD3aImKh3tMNBy8HtuvxFjNmqoc82s0dtSnLac
Og35S0t5/UWBx92QfQvPXWmO77rWFtBhjFtozS3r1xtk6yP6Hn7RbIMTbQK6E8rJrlaXlIpH2WIc
uGj1NFkF2ZOWfPqOrfQfcgXkGlgR1/KGWg9bvHGURvpE7+VaKCfO77tMM/2ulZeDSyI+l0uQJxJJ
DGwpMHODYs68BKKzk3ljanCg2L/BfLd65TztXXt3JTd9xaVG+8ajbQdLWrvIXHb81c03ceK8QN1A
y458lOVmwnpf5catNYOe721Vl+tbZojxNiBfHLoC8TQ0VTJEwAzkarEJJubrCL8HyMcmJvSWyJRd
KiiqebgxLE8PuyKuNQY9/i6H5ILO9rSaJw5zEr7XCObYnPTIzTjZOxSoMzvOk6qx6/RcblEoTKfm
ybnkmyEbUCMP7hO/jBatej4Ng1tff0zR2BjgjNLMo80pDKyuutrr2gMmQjeQTcIiHh+tPJ7dUwSG
xoLhYYQpp90H2PxkZbUJ6EHBdmcmQ6hSTGCdzLxah22CKkn+T+TsLXMRJ52PpHuQ9T8YLXJk4KbD
K0FbEfeTyIKH2J5GEtJS/K9xOeJ1BtO8GIEjJeqZG7AxY+YFK4OIX6l0ohYC9GRfAyMFLg7gd5aV
2WqNwfa8YpXaF9Dnqht4WbvqpHUfvEffFAzIrw1H4XJjtStPIZ3l8vTNYVwLh/x83W1OWgeVkmC2
fVCumXImf7eITw2TtMsD79Qj1mzw6C0MJ2YB5L1z1K33Q+77t7h5wxTfV7awY84UaAV5GQqvm0+H
52Gqc08gTf03xQ8Ebx3SDJAQJSOCS9ot2Z9vjxbHVdrs+a3Wu5A6wi+9kUK9luVKbH9EetIP3Cbf
QUlGOrk3PtKqcvUqzWxMBCLoHtIyiorMEKJFevZ8+EKe9Wu7cLcYk8/AtNYhkOjep5vp7lQ22XfK
ZxRGyCSNao+9u3/DwLDEtG+ob2EOY23Luhs68E/6lTOjLB5vSyZ682tQT4/I2FZfEAykRM/zf8JB
tCXxGY8QiMJFhMKIIOa3N9CnkPLVC3ai8E+Sf7y8l/O5MXzLPsDXabf/ohEqrDSPUmHZ6cMHCMW3
Z9cR06+42Jj7lwLk3EIlS1o3UrMbOaOIjScc4IFGE50CJSVkiqAHvCm9rOeRpOycKU22lj7twPPW
0YuHopaQWFjfg9+t9wHSXphsTspkl3q6R4gD9SAlCucZN07JlBPUBRKfHxLwsWqpPfYju7w8byvq
lSsxHoSg/ogR7/qZ0D6KpXUNnL9ncbRzlE9uU15tJfIIXk27nHN9yQf+pt7tCxwi2gEHT1LhZlIY
l/lMSEqfgdiWS3rPTEEYNwB8G6z89HXMzGhgHxDcfkv6JdPUn/uX54KsrxnEN/XWl3PBqTc1yw/8
PwtZJaBeXs9z5Z6UumYLpLlA0OIdWEv/aEN1GXdMVEQEpmvu1DRsNL23AkhJzUQZ+FO0SSkOrvvj
yHHQM3WJYZkWR9v6rOqyFcY956CVFDVMlZ4hRy9TkGwKouLdtKCURSCLyf830r/rvp7GJGPVs0+A
JrBuAynvwfL265UK9tDRlq2+cBn99fvZekoSx9oIrUYEWRYeo8VKZ2zuRfJGH2Co1Smls8B4UxEu
JlmMma1FsH06sxlE7gxTzmouA8v3na5iefdLY4qpaaOM3uXE8dJkdxeUV7nusnUqaogv3OWOSp+1
vUzGKUQ3llswTbmxN/o/PjJrjVvJoZcGTW74ipADG7prYHspJvj9oWyRBehGs5kmxQIQxEe5+KUc
U8EfClShlt53aYhnVWPz3tfWh2uI7yhq3vaiNq8PyxfKgAHWHyl81HFryQ50nYAOLUZ2vFPkbQ8u
7d4FDjcgY9EDYjynC1PiO14RxV/ep5TOtfMfrByey1PzmPEkunsJjAncWAcPTT/qm+54puwIVBN4
mjbX2up8VA4WmpkS7vsYil1tmc9rSMYgCio4TMAp/r8XgKzUUWQSf9Q++a0THZkLyL61+VsFEvbd
TEEEkpcijwLecVu3GmNR50ZTuPQKt9nZArQjErrxH1wvG0uq5qD4MXIbvZp6Jc5N0j+Pf6+cbBZ2
GCVoqFeEfCZ5ykiRZDY8fiy3zxf+qzwhn/6YaiRv6bm+bgVwtV0KZjG9XPtuESKeTYNyL29+bUuG
5sCNItfeAqyY4oCbZLpM7l8vIEvk8qyrGGRNNTK10shcay1+3AjkbdzWXh/XxiPd1aIJFT0PnJOA
daiOzfsizGYsK29ak6SLqmpgGzYhNFPkHOyjEkxzvXG5waUT1hHTx4phXE1F5WON7+v53CvH9Ajw
YXUzYbt2pcGadWc1W4aRiiyGcja7jr6buciOvjNIPL9iXCbsdkmBQq4YN0vR7G2BkjetEo/aMwpp
XsWXfglWcKOOHdGY6xMMEbfJ4ak1mbTjTwf4DK5hOY6bdnV6y3g4Ii6laH+DGEI7p2gOtLqlYSLs
gLEtCLJ6VsXHzZnFdhSokukzrkMGNPD5and+ty6n7y6Eu2mYlhVePDl03Ym0nr5FR0w4H8Ri9Hwz
jT3WCttEaUPjaD4aNijPw/EdynqnnFEzkJobX/Fmz2FdykwVhUZmH+J1dz2APJU7XUR1CZz8M1H9
Mn8umgexfG0BoSefRbeTCmEaGUuKxoIOncxwGtx4fh5CtIuA1kO51fOUK7UQYNNm0FKTsI0FZywD
HBTB/2es404fauW6tdNrRwAo/7Mcr8Uoa4fCXN5NU96i4rrtwlAf1LCZuOIrxnKYjKTZakMIdluz
IwS/Sdb3BuWGNu8XYV+e7WZyuZz1sQ/Wlp1+ceSHf4cbXsIos504lRe7yZHgcmEgaPSICyI6dMyc
puN2BsS8kjtyohUOvLfLH0VcqeQ4YtwSiFfS9/ekWlH0TWtzBHxayos/FrTKaRJxMGbZCvBCZuzd
G2qSJMH/oy72CVnwkJ9K8//9Td66MGlv2l3lwbEExhFR5LwpR49IOhcVZx/PVG5j8qScBYfTkxHD
j0W5YkGwPJpNAbicjWNTQSH2J/XbUNdsryCjV7Aggqh/Gd9Un9ZDk4Fn448jlj0Ut2ll5NfKnC7P
sehWWn0HTKgbLPQZhVgpHvBtpikensnmXQMXj3yDgw1VjFMJQUjKMRRHqFDMf3vQwh7+wOMFAvlg
XqBxCunw2VNnhFEDZdo0qsInEbC3yJY6aBiu95Ybzx2/jXLFycIWdYdb3Xf5GMMCY20mFclrYX2v
pBxSjM2B7sXzN9+ozAOxHcjJOENIe3e24OMOEYC/46DO//ayswZNpE5bRv5N8D78H9Z++Vg7tpOJ
x4uv2ksyiQUiV2rYux41sTzmnioxckJOomlRlYUS7t8xe5V6mVkd36h6eWBx0oi4ZLW0tG4T/jFq
EunthOqf918qHuD7M0pJB7tTnfpXo37HH+TwMzyt4q0++eFmevP2zdmMnLd8g5UkP/wKmdhAa5dU
QsQeAZo/SJaelcHuWm5bhEDFnyuWg81nWvPpzSyNjS6JX8lLOoWpr1omnag+koVelB0emEaN7Em2
OjhGKUgCi4sy+9KNlWy+AtlPPe67JeVxsqRbU8cODRdQNBuYmbyQ2jy0Z2cZtMrieIEkKCOu+kcD
CkNO7XKq8+UIFrv1N6SCSohGWjoBzS1icMp1FJ1/ACr6AWy3ye/F3Wr4+0vUYgPDsHEN+f3vgF1f
LUzjgjENqswpd+dFmnW83p3oj/xdaFbpEL5q5eJ+EX3H3uI4Gkpt5IycUxqP8lMHfUyKrijg4iKz
LP/jIJqwg8kuo3GSkHVKqqcHr1iKg4wZRt23NSJWzcZ1IFVxu4uqKFdFwOLpeJMW4DeUBGon+RI+
IP7nMksQ78dsTGk3A6LvP7tINlHWhxNBG89t5TuEb8HKOUap7CeRyj5Wf2gJ7hPuuhUplKWtTqBG
7faJUtMphLVumYB49zIwy5vFcYEdZkaKtqVu1CgMKZXR9azbITL3uswxfOJIxzKYNbPF0bdAY4IM
5g2skI7Lu4UIt+KWBoRJlC8UPzMeT6+K6JQwClBmqi+qZDM87oD9O10uFuL/eOVoNoMe8DirTLt+
vDEdM/G3aqzoJ537LaA6I5WjRIMMsKfTr1IuXIVufeqDxT5SS9GvX7ybvvre4ZoVnwF6AKba9ZNE
5GhiqQ0lyLgLF3GzZXTQtPMgbPdh+rWq2H+U4PefGOuaNF2staGCwF2ylMvV45IP4oUg6Y1cq6t/
BcHZLLMRQ24PVDE0+h/IoJ8Qu47vA0cHWgl5LMFgOhZGNzcpel9dy6DXfWxrR88tBGhxj3cAwtQT
Tp5Sm4PPJC36FRuM2sV7NI+dJepUFbfvykmqzWrDnUhz6THAz4OZAnWrT1CjUEYjkTy7s5mSfajn
qCjhAEA8sbKC/a5rlN+pFPr2UTOxBRP1B2n//PQb4wqB3EEfr2/ZlwpUyqLaBfcsHSbP3XRiyjOn
/on89GnbaL6u49uyDNHJBI6J80uU+k8Jr1lLeS6M21a6uP9vQHWKlAk5/hUAKNOtk9/jnEDLpMLn
c539v9wKNWPfXJxCRLZHREmGmXVniSg3ZGP39lTai7qgIKunI9nHYqUhGo65jLGVaEI7a2S+RvdM
JXs0DMDr1150ySKGX/F71JwUbZ61cLWkYlygOR91XWl4r86Q+gVJH52k9CxAgW7jV2658f5qCnl9
NNEBKfZQtnwGZbfU+St1T+li3sAGGJu5CaDrgF6KdFP7RT9nDnpOn1eu+Nqdg5QhjKEbIes4Acgc
M/XpWbg672pF/tdb5gxk3XtKXe+aiIuOG8E8kXEt0BpN5iMDcbhTWKA9xK2DtofW/ImBc8ZiVP5Y
UX+MAVnoueKGe+GspuTHJw9peoOYIlB1Xs8358NAj9XDV33SB8Qkw0g2OP6CJpsrL44XTq1eXg47
Zp6fLxITIM2YAuDgcZeiDRUT7CaLZxqkW7388rHbVjYIigjdlSbqfGyoB86angdm0PAj7ZBf7Fre
xpTuIxUOp6vDfkWPKGcVWUC4Y7OHDJzow/2Zd7xh3p5+9WaAvUXRx1x1Aeap1CwIMAM31ER8jM/x
3Y48tfwpBtYdU1bFUHOE4+JtldtZR+sb+VvacKc9PvQBxovxckamQG4s3K4dSKUY9PJ/19WABSyU
75vazZQu1Qs9Ldfm76FyGBFuAqot21eniNmTQ0uZjGnTfWiYS1KDDcdhVntQSFPOqD08jSwNAHzd
LRMjpJiCgVo4yvuozcoazFr2Sm4wsFBcE5JHQ3m3jRnT6/SVZcx6mbE9EnYmacQ0J69aT1+oi5r2
9oYVc46Zz9DLk05Jp5OEMVuNh06/kqa4WuY6gg3kiq3mbnM52UPJMfpelUnDYg5b7W2sIH1DxSQ1
OG1iVPsK8+UqzjJAS3E0lfsEikaVhnRD3UOOYXmiPl3111PNLmJ7mmiwoVxFI8ZZvu7f71h/BkD4
E8pYuffT8oU8O/kcC1JW4XOiYpzQkrwm5f5tqSSnDzx6Lj40fnHPruMs5HvJI/QW0ZRV/fhAI+TJ
/GlDtsur5pr4cr7OZ2zyPa0jwQFbsdpR7cDwE4DEZDCR9c/00X41YjhcGoFgvPGtN5I02hgel1wH
HId/6aF8cKHX4abRYLw2n4ogorshmNgokXmD2zScWPQdTXy1PM1tvNc4CPwTHMgZ2v2bSiM/D4GV
TsOKovo8PfbqOuLqjcZ9tzw8zS6DkKzuD69tuyyeA9M7M0UNALN1oSU2t9BSIq5rzkZbnSwTG3ge
qVmDCuAYTCoLSZHr738ertnOw2iy6x3SPuvQ58/I5VEpro3R5MJcKbEU6T17f+z2fVe8Oh+9v6mc
xKsC2NgEnhGHAq64xO3WE9YUBssfNl3OsdbQZ809VBfFKU9DERhw8H3ZH9pJznj5VVLiMgIRTJia
zYaSzvpHtuRuy21xr0YEba2yOGHE2YvOP7d/7bMAmjjK6PxnxzT3nzLzsv8QjqNoHWB/lWzw0bbS
VrPppt2m5PoQcQHmeQonVuagijZYkGAeh9PWk1IEs3nvwrp+7w7+omYUyhxwtQRP9CJS93aCKN94
OSWG+F20A7JTuZMJjpDn0KhPr5iPZHhV8cWkMvnvbT7kvuAp0Nc1zkrlfDJ3gV1gQfx6ryldcT/8
pv+rYWYyJ+AhKrCZichU4mD34bu5Evy0RWNNZtD3vhgnuFmhd6nnHAZwXzUD1XeTpuf7FCv123sQ
Wni6wcfJrzZokTf2SfEr0vrwIDNdH4Jg47LPo9i4wCgVRRnZfpflmaLbWkfTCfFcSNDszgVyZBce
yb1323XX5kOjhYV4o1qme3+95OXAaWPgcwP2f2/rYtGevTR7Kbj5EjBGWXqHcSW7ukkk5bVKd8dZ
AMkCxWUP/1j8gdyvIFxeV+hvLgtnyOlaQJ44PAl889w9vOlwEXK50IPgpcJI81uOSv6S6TJ6N2AN
2V9dz4+HQq7Wlt8H2VPNhecMNUobhWaXh6SfTbvAzlESKUxCBIJhGsb2LxB4rGTJDGFvASl6t/Xu
vFNtY97ujfFeaL+NN55GAxd+NfJpmn52s+o86yUD8BAeGTuUkM4Q3+COYa21ykoWnZY/Cf4fQsrH
iTHMa9PMw4d+IByh+p0LP+6niBnRnBayVaU0yDW9Q/+L7D9q/jZ/jYulpLpQopDx7XGRIdGLvxV/
3jbqnOesi3l4pUtRkE1l5amPI8UfgXwCAtqYpcIF9NIMvkkSNOU4XLaACjZJdd7k8qJQtAa04pgA
/BlwdqGwtqVlzgCugrF7PJq/MIzFDxCxpRtEv5ZFJIqSndp5/LirASRhw1hgxNf3IXHRDIMSokhE
LGOQ29YgEa+Qmcb1WmS3MvzfnaS42LSyyUTq+jtknRCNH/xFeOOTZRwtfFAaYsM01wtJb/X5DmFc
V+M1vUGeQN23YBTzbGLqwY1dbGLawY2SAt2I6G0s/ZP+C5KmpwPse4goSwy1Dysg8D/kowV4dGuG
h9xC4XVHxuZ0IqiY8htOKy2rCjY78RYEnvyhF7S6sNZcgGG5DtOOk0KfwRhJqUMvaHiDTIKXJz69
grRRWZYvyripsthh3mJvb3VoJEu5gJXoWcqS06baqP2HsWMhmOxWMh0XrHMrxdSqulcL7TqCEvCT
yZDWLOqtXCINO6LKS2YkZ01RDxr0CEIPPT8R2UR6r/jLKpI6COXJjRvOOJXz1HqxfjDh+Eryn6AS
2xoCKMFzr627B5olMINwmUcdS6xPMGYxjILkB1jaxYIzEPaCCzmGiAeLkr34IgiFQY4vDQie9xde
idrzOsomqYexhb3jltAbHQy9yjgLJwQODK5gBAJ99chDvVUzpLsv6E5w3zkGBEaUNYw3rj9b+Cpl
nZzT/rWUqjDyYXdXAm8QKXSah0T+4Ikmvq11GvMMSvdXNkYv3FX9eSChgBUquOX/TaPFtRXG7dmi
6eckrpB9F0b8i/+mFmUdbiWMrxZesK1awGygXGPvuv4IMKE5bQUgNG7yEA3hhPQd2vCebGVDjQ/B
Wcfzu69+uD2ZNwS9d0L2eYXsdUvHPOrawlINaKdt3aX93dIgGeI/e4WkVw0f7BBZybQNfmaE44pE
Dfvrg46BcNfPIC6jxx0Re4xMWaSPw5RZ0VTCNwncK5LpW6pLXzE2+mh9naU96QAlN1VpA2spFHwA
ZZ+Q7kZkTufyRHWf3BEATkwmOCAEltH2ewEwFgHIcA7v60sT+9T+6dHqZtVit84vUzcxeoDb2GKd
uyeu0MWmtWdmAESQUm5/zoR7VfeVy8Bi7dAI09JrysrlPhfFQPA9d30ccyXoolSkzzWQ+YgZxHB5
7ekgNbjKQ5gpgpfhWJbcXp/oi9qe3JykiCR2KFuGKcWneWYQM3YhWQEJFnVNtXn2xmkAZyGAs7qI
FHfxrFl1b8UiQTNG0mFdyd8LAquY+I91hZwuYGNhVEil/092psaLeOUSAyLlKEEg3M1MMuch71H5
/gTYIrZQcjS18zZLEA2L6NmvesxmOvCySskLC9I5YjhkqMg2RNzpV6Q3M14KFE+vWLWbc2PAyYTy
Lw4Hk9/idPTQiE6lIZl7Wr/LJjRAM/DbhqUnj60XpRaLw+FEYbqa4FB2zDKBS9HzLguZ7H43SO8Q
/QBD0BQXy+cWoY14h6FT6PJ0U/tHtf5K4Skk2pFv3qUJ07ssGRKoGpyCgWbWHgjR+/FMIvAs4QIH
i6zesZkKVguidzaD+GfM59djElXfaNi+9baeH0WldQZmZgeT5PXrq1VuDoIbuMG4ga1oSqe+pjQP
ep5sjlQZ5VvkWxhi26gam+HD8f2dENFZhWg26HLopm9WiuVuQRcJhMA9NnMO40DwJ4EKFBwhiUwE
kOymz3nFtIrTuEg1+3Jnp0dkfX7YOPdfeRAhFOXm91dnyh7Y6IJUsTbEJ4nNtl7szsQZ+7TolJP1
ujUKUeL0kVa7ilJV9I8LBZNXjJfcO2VJMTJ5V7gt1eSwPLG95yzdRu7F5FQk0plRL9O3Cc7N+R3o
EMitaZTaEwYWhhvKtqOgW7sSxpl+CZJCZA6eI2AFHxsxruM8sFVZiX82O93t8OALvu2ZwaeL1Y6g
plDYXBNUe2wgEPoyORzDmtY1PFfi78z7+PmTTQutYK7zpbxicOEfxe9S2O8MYnOY/d1lu711rtXo
W0NozY8uWJhXkqCA0iGUpi3fJ10rkwJhqQj+SSG4GeqUyxZ3Q3HAQzcc7Nk+WSDKw+RgIq5UuHJU
tWuJzEySnQhyU0b12cZqvObSX4scSvkFSyUzBt7AqPkvjQ8TS5xFTUk5KOSZ039909sq3drowfaz
bFBCskcQqVssHy8rDCeoPYAnvM7eXr39WyvPmyPhg+1ns3KOa1/HPJoaI/qft77qrpagqcY35FNT
UNmwpKfZbOoOIuorvW/veJq4M3q0WUbHkxJ3/s5SQiJBa+Ax482fqxv2qK1Tuf1so1v0q8aGhVF0
McF/DAAdxB+xAZGZysytFnnlhQvFW+YJ2jL7BfD3y79odW3pJ38INTXVz6A5N0RobNxXvbHexwhm
8vEIieDHT5a29bf3ax8bgqP8iFBUaSTUtO/PFCQcBdhHJoT+Ox8rMqrblWKd8DXtdxW+cELHx880
eGf4Kr08Kjy6bOSTvC2lVueXFIJP34dwA/ddx6xV3Hhkc8VoOk5M8cwdvkL7GyF4CPWbB80TaFFj
4ZSCH0nCAMTQQ7dOzb1nvZbV5eGWP5+vETZHoiiEcBqRb69/MRylpEFYZPyWlZc1CqhxhKRwkFC0
GbDTTv8OTz11xAv5PBImQAbFYfuMDXTpKtOsCkyNuHz2xyNz0nEbbvZt1ONgR5FgXbWqPwAPCda+
6EUe10JWdXhql9eFDCBBJBUngcjh44dFnExRvhsE2/sUMpkZ0Qx30988D+T5H8DinOZcM6svpecJ
mOWzNTFTDA2upJ3ZZbPCBxy0wLwadW556PNHdhrYwXcyw3Xs6IM7o5uogt5xlh/oANFFak1+TjTt
ZSHUdveCt1bM9FaQPmaDGiVIIr6eHYUaEYdi2lhksURMAkWeTZPC+4Al+2njXBjyrLqdTVC1IHVJ
ZB7s8ihFpj+KKxaHxgZymlJJDSBO14CHa+rE/nN4OyLKQosWmxfkJb3Exva7mToWSHpe8rQgjlFN
B0lswJ4LX8/tz6lkTHDxZp7M9YAt+7dhV3cAa/8tmlh+PxlIzVe4X9xvcusektdHaNJU9uuHYotm
y1jSH7tOWo0walgwSJG91xdjhylCnawTgGDQ3b5ISvPBxigcjwcmhExdR540Jssc4QdQPHqJHmEb
AVReqUJ/qPR4IFqcOhZRtq8NwNG9LO8Ves8kRn5/QfAFi06oUUY6/FvTBDlvirM5XlFeLgSQqlK4
RiV9ywuCNzhz6+b+YB6yW1Ox8xpNQMi9zj0XjhvYFdV86npYpgPmY+dBP/WpUsnwAzmtwaYq77sb
osBjOWxFbup0y+M2jgVmo1Srv+ODx8kScg5DFd+ia4CZESS/BC5lofCLoDaF4m4U7B4y6Pul4+vo
QWklnDi4sD+FLjtVhvbpZsr6RusturhQziYsLylL44u+yOIPl3ZLSZhbQkHO20AuSf4eaDitutJS
ZFFoZdmVv+b7yTha0W7TBsQXt+RASjaxic29X1j0GS71/yDZaf73ohxmPAJdzrRXz0d71D5ubeAx
tyOKwBqoLXXIB0d8g7dJn+is+ztUZiSEaIhFv7q72o5GRWT0S7i6kRNincc2vA5BTsKoovmGO2hH
40N7KtvRvHdmzrVy4T2IwP3e/z0yHpkbgt4rbdhiRLPz8S2CKS8ZfcU9UF+0FuLsge8Uf845AUBt
nx5aVGB4yNTLjdqOWF5KCDmwncI4kiflHWxPCZPzr4oc0/lZTP6cEXwrlaTMY/Xi6Qs6D1eakds0
4KRXj3HqKAx5gHIAL4ukvnrlzMQiOUT1iczM7LD0OpvkfV+ZOeniCiL0xQ7SvD5pYW/YyK/kejON
TMues+QtEI/mcUXPA9AdT14JEZAoDdjKmraULwZFZGByTMdWKqLHtMXV4aPGkETUyPFG2F9mICnj
AXvo1yho0D8HfcGYXT1y/qAUyT7HJkl7HU3QaKzfQh+oLetIg6oTt+BXrozPxYHSBpPBGuGHrUcG
FCeOzrZzni/F7A8mL9Yl7JlNPo9ZRI+yUOJponUVmbLcDGLVQdWVOIjOu2yoFURXzJpR1hf/n5aZ
eO1S44Acz7hP5UK7FSLFtI2Vo1E4OrLBIKXEt466UjWnyBX+i6n1uL0zwPH6kYHyZuA1cDyaBRTk
DvjfI7aCu0u5CnlePiY2wodtdqB/QZVNWAFaxXWv6e2L0frxMqi/qhWAFEsSNOiZGXT7qTaJCfbY
ljtUOoPDFB3DSkXk5QdQ7wHbmVG2sBZqmmeO5pYkyDnutNm94g+fR0T7FpYjEYumJZeqgZcZ8pJ2
UtW1NNlGeGl1qX/5aSXYIqZ02ec339uNUPkHvR2fQn/W/e67pNPjuNIotAlnNQVzLHCojHsoC8De
ETEUeU0QZ6VlBGdy0fyeB4Armb0cJz2MMCRtu6SiSydMRmfgmkVbMxSduNNkHegkSwH3Nh3GoFfQ
BR+Hk5nKpg/7SwVqh1kJCllzHbDjY2BqA/Ti8/Yc5fBmnfkoA3ZEwDp6ohw+elP4p5LXHfbzt7bN
XU2gBU04mbeUGpJZKGzFWCwnIfN9zBdIhjv7ugYYLkv+fXfmxgNBViauWtjfCy8txhAzRstzsEAB
js/KMr0vJzOgO7Rmkh+4If3tb54sOOk0rAf8TAyJ6BwE2KaVFwiLN6MQviP6WGjgUoux1PHMfBDN
9c+brStsySbmZOghuifFh81rE9XBMpo/BDJ8xSJuH8DG5VZ2mVdyMOSIfZUqNIY2zB10F33aLt2G
MKPT7k4M2/STkAetDdrC4kEGMTJiRTX7PW/Z46dHozefTIBolgjgMnudxw40+Hmf/m9vLbqBBQM0
5VaxtZIcU/xpMbD+MB/u1BTugLYU532L4mrSaZL4hopEV/sk6m8ZCajvQZQpYNvLt20Men/5WQq0
CqPvgIhoTc5cgtmzmjTT3TdVMpBRt4ADzVo2jCnk7118EtZkejKuhmgIF1oCFtBJ9LXwIyesbvqw
qThzB79cudgXObpJfG/Ckb7qn/dVdkw4JSEfvKh+jInaMkaLy/ZS+S8S6+Ai6kSTP3FWU4P0yAP4
WWfqarvKQJQA6XcJv9yAoZBQNkwFo5lezBI9+9WTt04pv+se1NwHYSSUjqfnXWWwV7YxciTlLCWt
278Dckno0FBC/HQurVthrBmBz20G5Q5etdGMszZDRL3AqGHFu9des0TsQ6Y0uLLjUkRQn+eDZPfm
KGNuVie1TFacB0Px25WlAcTIlNIKJp4jLBhlOhZCdpABGoJhNOIVRdjNFU5e4TWXhVW+SNjgp4MU
6A0QFXVmygwJYziaO6rxsS7RcrWmEdftOnVrbsHI+CVck5HjvhAgb42FU5nDdros3j1+mOCBQd43
rDKOtbili8QFWO8CBZlMyp0dFyBcHrEv5FeN/+oICm5j02MWEURAMGGnF3aG4wi2e7e2tBlioirF
ju7wrF2Wyz94jnX9gB6rVGkogeNlKIeYMiWGGlvjr9V9av1dKJxEFZWV0rtBDXMlkrvZjU4ngtoD
BQuhyu5rwVLPVW6HgCYS1QKN3OVouhOEepmUIjzXU1npvvdaUU0R/ujB7lB2FKla3898y6CUew8k
d/bevDQ/B1duVQmYPvpHGFJw145/Tlp5CB0cWfiWxrD+J2ivBEIjX1LxKbSBMIxhXkRlygLW9BUs
k6g7EPINoqZTZ75QB/1Ve6vsoV97s43WMVAEG/CpBssbyIpB2x+FsrtJ4eoEi1qTPbCUZ28x2lW6
LgdyUe00K3EXtaE4pTO5QxZIyc9hVyeWWcVAgXrRhxXocduPCC3o0TDUlUaj8Zu5nJt8xpEvM7cm
VOl2Lpdh9K7PAHglRiblWIJhUtEo/zeGvZ0qDfzGTOuc4KbuSVxTGwVECmCyXV1EGD9tTeTuHoqI
W0IVoDdkIDmuywja9zzvNQu2ELAZfr5c6sViO6Q484SSVDgepm1e8ePpGE/bKbhVBLAoM9espl2K
7BzglX3R/q3v9SErQ29JqYhpATaLN3xENoSxW0oZLdOKA4g6VIef/09+v3JE2nJSHBaF+cLL2FXs
bd+ZsRe6DASfRo9YDmdGFEupd1goWDaitMJAMJBUcbC8HHAchtquteOuUBobTo5G1NCX+fEUaZi5
DIpWD/BV/sD01n47GduJeUeU0ymHBVxu5HBI0FTp+jU/73SASxPxCJHW014OXJ2xhZY1eV7KN7p1
TDKgMiHEXrkmqNoSASiNqyKh6BIMUGsw7DdUxiRl8QhHxTm3gy0u32pihDMwa59FW3CsQuU+cK0w
cGQUHgwUMUGsGn7kAnB/riq6UNNLguNoZz6BzFrLp4ob2knD0MymmukWQ3XUOHDqW2tcWml7Z9vt
OsyfKW+LcyyuwnQPPHestNpD3e+U0lY5jYh+PoaoIVfUeMk6DQresi7ilpoawBGUv8JjG7lpB9/0
a7e4EGfFJy0yhY0isB0Rxaax3ZF0MmxCLGtow8eeJ75hwciuP1+1HFiVuI+VqmDe/NQBmIP7+foy
RmBGPZ2FqVZDTcYurb94xiZ4mXrWDr9HZQnKrnY1Z0IS23wdPwUQjnuPsOqusg/Ywq7iTLY+clYW
xCjejQrVz/mUJi+FqyW5F4QY3oUgV0aGEiqMzJcj3rjZq8DG/no5N9epZOM8hZiRLC/axJYfpXHs
39HjX8K2Yr+8TDxLo57c3QeDLfCSZBsLCR/WprC/7XSlcxLnh6sAMvedjBjIRi8LTVmmG/JmuNyY
nA+dhr//kijn16zLrKITSGRkOWtdEEAzVDtFgNBLbDZHbiTDkf5DQu7ma/o7UjhtkNOHME0qcZIr
K1xY8wYcU60908pfXN3qI6yhxtPLFEgakNNa5jaGKGDg16sRupcOdRgUxKmnUNIoLcNj7VXDE9Ph
sDUKyUwRhrRNso2EldXHLbqbnAtWCnH/lYVAXgrbK244BdQjVMfs6qGZ13gtba7mJstZye1PrE9O
NhKn2GhKFhmtebsxq7J0B27BPnyQA3mp6mCV42bRiNUX4pnTYBHsujPyr5ovtdr4RnipY4n5c7pO
E4osov7zDC4wqf5b2PqaXOxqpCaj4JQtJUq3H4wHnk8A/K68mSsEqq7OPxPKWIte+5SIEoxBdfSr
R/ebbw9tDpEKQqeg0jb95CwUCCBur3ZkKaX4d8bG7njenZByx69tyBdoBm1EfYjFTk07YnOkMj8k
jFe9uCvXVfuu1YbAPRC44Bvtac/KoFJS3vPa4H57Bm1dlpqKds/g3s457sjUEyWqhCwdQRLMu8Iu
1OiXaSJNA1F6wbcFjruvmTH3auUrcM17u5l8paqymAPtWWYhsXce5oC/2x8SvHUHzMea/NiuCH5k
k+szV5MuvzGKhYHvAGys911pX8voBGoyy6TUmgazKEUyvVzCKbTFtuAtwrqGMV9uHXyBzpjgi3e3
iljSux8EUcQveI6npkkj2o9OR4uV9ix2FMlQZmvRRgeu1Melrxy0mwZE7IZ7kP0Foqp0K8hVj/Yn
2bek/NBSfyWEy8AOVOxtNF3yJDGjVS4oBinvKc3qXIQROmcVKOT3BIxxEXOYaDP9eafWcHPUqd3D
+iaavZtJbRs98yHe9NiaxxnFN5nnEWo/zTXaWaRgSKwceH9QHuSQpQC0c+nNDM3DR2wj0Kb+9x34
KSNEkCR1r0+CJ783czWMkgs4Rsr5tAPVhgkjwKyfbsTCgZp5bJl9FVGko/Xv0KHvL7rBJUU/o3eL
kei1pWFPVcDO1ElzKlFufHA4kyv9Ewl3yQHcBUWhKVaFcWhwLkFqpBeNXtDK90D2C7uiWqqzNjYO
EiBsURF4GzltTA/MjToBU3H3a0eRkfMV8ITkl36Qq2dcIj6H+GEaKbFIT7aM4o8Y8X2hVk3XEdwH
iePqKpgLvourXIbc6+qODKy+z77o4iCmwYGL+S3R23AiqBMvu0FgGcWo4dBlOVY0VD4bTQfN4F+M
imBppQY/+Yba1/2+ZgPKxN4gbyNrnBYnRr1bIWyEsncxrBSET0GK7yzQ3lh1AzyQ2UdObmLC4/er
RuMO62BfTzpDlLqNlVKaGRykfpQJCI2IfRqBamoeae1Ndc9athb0dieHgUthRhGCu7gIZhSvSWpM
pNUk5pPhWEHFaoAuxEwql5xlWSMxeoxmutOqUVDqBZtAuwAUabWKi5Z+FKjCWtjOjmTzjJ2WFDX/
AL1wMm2hOFQmPw61VBYNHttZDQ131K9f00FdP7mXqxJtXIIVIZftZHQtylzLEoSf8Kdb4xoyGar6
dMo5Oul6PqHBPK50XdEDK40TH/zvo299C1JsYnIiTPEOVYH+/GC5k7C/si4IJe7PcHoYgmT1VOWW
5zs2p1aeWqJnl1ITm2/glIA9gkjvZFP5HvLDXiOjaq+/b+RnUeglS4Z6Bi0/fLaoKmmySkX1wkUP
+4V7sIPepJoscZBAGOr93qbe5VtOpUrrz9mwN+xhiRqzOgDJkyMCFCX4OUmNBHArBOFF2+4ffBsq
8l0eClseJeytuWpzzsH+ySPHQHqbIvD43rBlIYirJx2teSGIfqJM1NNuH/zE2zYtC0byNFoqk7yM
XOrhZ8ByvP/WQKUG5wbMQvQzG366wkwmM3waQpDjkKsPPuxFmzGBn9qyX1yF+26a3poBFUxOMHzH
/PWFnNxNPl3EoDvPLohmpzW9Eq7AowCj7UVi/145LIaWkB6LlVF7RY5qFg4YqtsVGsHZKe36RJM1
AwvDiW1GM7MInvAyR7ZPK0v2auMFHR7xQjOUMGbPtJeb2P4vOXeqoT0K550PqFX7dAjH1bpii7My
P98/Fw6aQ9Qk6k5Rulwbviw0//SApb9cLru7Tu0/7cIA1IECLiS9k1xdYiETwA7K4SH4jNTWydXR
yygIrhCFOdnGt5o1GpPIe7auRAAMMuaLAnGC9ka74ERopj2IGP/ld0h/MKbqigvyNYlst8fkAAia
hW2mHPK+Twkpe5beU48ERvXguHyG0j64e9ZrPRN++HAahVTa8h9R/UO8JK4fGsZ2zwlnBN2K2XWx
Mg9l4uT/cxvxlFLKQntwkPgO9ER8eyFwfEIlXNPIXF10Z0I0EcbAT0GGc2Y4yc9RXn6+bw+fE0CN
up3t03iFXlSUn0vxW8ZQqxTSu1/HvYIJUO7CVu1E/2zsYL2OYEG7tuBfCWdTu5hKbIclm2pGfFee
A5J0RR2SOZgoqE6DnwhAg6kORcMn1aRDiGR+NZLZvz5aHIlImlkFsa0Ptw9+EThyhVJdkcrtG3Up
XqlrFEvBKrwCkBGXRfjGlEaf12otxMK+hg5Eh0P3H1/xcfkCgupO6Kv383Ki7OEFMS+rK3qJ2eQU
hqjuMUHcRvIADW11M9c2gVhqfkaDEVJf1VtYoetrvTYmoqsWfg1rrtK/P8VOBYHBzPvdncr1g7s/
mx8X+4oc3I7vEY97UnQoV4NwvH5uZeXWyLAFQxsWnoS9uXLeVmFJVDq2qiYCx2F2ZJ41aMaITOQl
FAAuxsqAPXCsMe8czqs/kcLfoxlZHsvRCIENDK1SA0JboLpsEy5F7vHkw2ZjbTJIQIGuYJQFSK5b
+eMcN5Yywo02XmwwA3U4HjtT4ANqviYv3a8z5c7PG6/rTUyG0x9rVJfG9kvmj78a9+Vba1iFqOM8
ALeD0HVwmFS+Ur1h9KA8bO2wdtgovV+YQ7Mg4fYN3yDiFIsrO1rfDSSCMPP42SzP8KwZ+17E4QBq
icEwQe5x/YSpKI/WOIRBvLfuqv+KD3mqTChXoTSmvnR7XfDomDtmiByS1i/PXxTDUuMFyX5WtQDe
Jo+hE55PoQvumNY6+vyGNcsePGWJ7nb98UpZ7vRU8gri/2bxPBIFV58T2CpGRsxRsmiN//THKYYn
7aK0QqwuBb/1xPQvltzpBH0ZpJMfbrJahB49cTKIFzCUDZyWfuig4n1aGsGJdqfECYVvcllBWJo7
0b1dTBRjCN35JGU9+WH1z0sIfYH8FJlpEqDcQTFYmbhPLL6rsF21sorhTN/SepeVHLgCTQFSKkof
DxkekchZzgxByWKUhpwQ2AMEdU/4481Ypr9CqsmQKJ8OHcel+1zN9gK/yHANhzgAqbDeKVw9GwRo
duKUyEX9ve3OlssNLwOTAQYUQvgpb+zZnocaq5Fk9TkfHPlQJBUOkCuqD1PxDVFMjSeT8cgAW3Ja
pjFlqKlTg9NMQH1yfttETjPhn6373bfy/3rjQpUc8KiE95GGQpp8fxw8p2YJ5jeJkJp8a+h9fihi
5dcUq2ZnH84HJ/Zt0yauSxUX/4nmGmThiWDLXNskWRbOuwoYAsEwuL58TSQeWk+wRpVveSjAdmOz
CWnD7A4zP/qUTwctsjmmXaGZpw/1zMKRMjEaoMQtk2JCh3WAAFjy2FDgKVFxXlDfDyCkhSq8mEqr
tLQt0SpsU/zGSdF2sAzVeje0BcnP/ic3i1J8jBweYaLXVML1UChX7PSmZWpWwdhZQSbWqvRuuuiz
vnTvqNQVxj1Aswza+TzP1wSESGnwO19l6YciljFSlZIeIhRGZMMohhJtx8T2soGT7Z2/VB+EPqza
U9TPdOdvKXwBC9ASui8PjjIA7B0ZVIaloIPDu3b9+1CytPxctznfZ1J6aurTHlf7bV1Wls2x+C4+
l/AnJOLSGi4umOD3Xbs1s7OgZAo/li1MZO6PXwYQRjajoUI0kli3niIAHcdzi10I/pzv/JfpCFwL
pob+AcQ5D3hTZqIwwuc9335IQmekgSNXefWuaS3AhI1d5FV3zhxHMJqBAlEnfyebsj/1O4ibkESe
OTVKnNvVQ7PEOBo9OfHHCMPIzSrq23JoimUNR5k7QpYyQu1L6nw1jaZ91/5zVeyjvClNOB3k4OUr
7RpktlvO7R/gQiS+W8o+biK3h37zm29lLTiQ3siEqfgAjFDvzRyDH3b3i8hyvzd1uQJef2v5+GQZ
2sOi4I/q0lidikrK4i/hkeu/vl5664XcE+ov92stiDdwS+SsvT+7XXRxclftTeqIId9HwPiTf+yk
2NEUrzhAbj+Wpioylu9/dmI18+Wz5FqDXcgwwPFiWR3jog9Cu0h4rV57Gv2951bzRZSer0sqU8uS
KvAigXdcgkMk8SHBlEJu1qyh50+8jyXYPz+Br9mLG+1L920HIa4PrhAN7XgPcM0cW+Y+GLLD8byh
rMlt1v61/G/OsLUKJMHocYjilHrpjrQRP20mE5OEYZSRfazH0jUJMrxJ7mLF3qkEUmp9n3w6CvCO
rsL1DsEr9UkBPY5p6hDtClgFePtLwpZWKzPWOd8JSr/DgG8UwwRvr7PgYADhwblTptTbtZZJFwOV
S0LP36jS2YrF6KftOHgdUDHsVvKgueNLi+Q3WbPnGEgfWKYZjA+gTwkVAOlX0RkPoH0XobkYtD53
pzOLl4mpApLTZnSImKk37yIoQo0ddcmlr38e3uMMgXEnLcXcODHRUf3Onxtf9gjF3/HxReq62J5T
sd3+0O4gLWjs2MEqpkb9A7zCcQhK2hSlJW+PRIkAe9DjXcQj8/tqJyfWRJYEa+h1D7yzMEs9nn/R
pL8GxF6CGhnTjVMiPOgVwOFNvmQUw6wUYZdLXFnebFAf3EjftRa4xfMY+cj95tOiKPLAk+gIBBRB
VwW8cyOuEqFTX9bGpfKdEK4UUSGmoSZPNyUzsmrqWfGOm6CfEbnqi8vA4Fe6il2tDFw3Iq9taOMc
LkvUy5i9ka/uAzV2uKLgcoijADrkf7/3akAaOtDMdhoMzmRqDBqnVJlCAHmybcKnNQemLnS2OkA6
0tGYdcfMYO8WvbJf56ZpnaT++6lIVOR85150kUBt/UGtNZd28DPCBMEXedZwNvekPy6UdVhTuJNU
EEK8fypCzntX/AjOz8aCEGu8w/a5qYlowV0JH9Q3zjkPvYbmij/kt83JnrIIi7EJSKwhqv8JtGWO
tAyiOcFzLaMOz/MnK+Wxr8KvcU4cK/zYjD+I/9bq6oWJHlMOhEi6Dq7CdjcIKtV2ZHdvzJI2+PFn
9AVkc0kT6zbdJxF5jkUgCqTBmWnNIyM8w7oz7p649f/mKStFTo83wWjQmoJ0pYA/qqGf0xs+357Q
OaFi0smLHTk59vW9/T5Mj//Qw2g5NkxFLj+IqT0pxji7c93GgDFBBkkPH/55dKqhCMOWw/0Fhcbg
yO/l32gELLwCfH6+jdvhyeQ7d0g6UpeXSHcQ8CkzYTNWYqNcJB3SZEg1NfQr5bYrFFavNq+w5dPB
/Ifn/7iQNQ2aAmEhO/t1zX/7TYhiFY/NoPFg6UWiRKmnPYZ1nIHrNaQtVqoYs9JOjPpSf0vIGXZw
Aqi+RwFidOeqw4UixfmfzbdDRTmMDgZ951QnamyaEZgJo5tLeXfJfB4hWYJTkKrYzzWt9V0OIdbh
KG6GrT960kJb2rlJiT9Swj77wl9FSpdQPPbMn77OY5Y8KmcNIhdo8bYnTdRVsa1JWFKoP6D/ec/J
U/AC4UyX7f86v7JudqZRrxjHhLLpWMh9AiC6GoEB5GupGr04CF9yKx90B2EEwLCCUQDG81dgr3Sq
3C0OGLfsQheIcquR49jS5EMK8MDJiS+JekXPnhwY1t9NQ3iyrR3PWef371xIEJlMwyI8hS1C/h3z
0Hfdu4JkhPnvEW8LMsb8+vx2Zr8lqrywmpzWjRRbTzxcMKCN17J35zPOqmp2hNoFYZlTr079kgmQ
3pkWbrOfCEYqEN7n9gR1U8G8sVu5sxQn+SZZKWHhVDWaW4gSkbE8bPxcp+bTqcPlCYKNpPu7a6a6
WMdtvJJ8+zql7BU4DL5hUJdWK47HLkFRsM/F4i42ZxF6X5lm/p6ybekgvhNp8B17lmkWiK7AApyV
8MOM7iMo3mK/VvVm5TqyGBgExWYNaiQOxCg3OtoxdAc88s2LS7y0NVpHsklOUitQMspxDFLfNP0X
p7RdyKaz8sLUoQxOxdsr/6t1uZdM18/GMsvALU5zjfAq59UfR7Cc5RS9vme1/R5Ey2nJE9wgSzUt
jOvsgOWcHwi1ByezC2rRoKpnzG+GGxB7SrL6bPsjn2lolvvI5w327+FvVK641toj7PFquQ9CyjtG
+e/twCojxVZ/vuZVEkoNwr0BACYqMRAD5miBleztPeLnVK5WQ727Sr0HU+BKeLmfuYmX+scTcECp
75QfUKIp/cXViNPDDznkNOi6NBKSM3MXahcVIFwSRYmC8m3PhZbjuV+l8sJbQP5hfkgIvkMWbJyn
NNc09ziXro1N6gPPqeVNfpH+Rnso9z0/wGhgQf+RhH0o1WDE50smMC2kRBjVw1g0DUsW6I/HA3Z4
Bp1ELoOa0y5wE+KHI0BvNIGmq/zCZtzM1nFYvf6uLrp71FZPfNiTqZyD8WLqqFV0uVhB5s/L3SXy
PYahgFiGaLS2nluV6FLEhk48wlJZpM+0fdTVBpLlp4pbUUjnv3GuZI9eUlip3br988jw7aiQbwi9
n7p4eQ627hbA4yWn6Vi6/lNJ/ZxPEKVrHw5HL3u9QiQzIZWLIPS/YZvwukPXyDK9BeXm6DiB8qPt
BjXckBi8IvxmFQyVOhoj9wU098OF3lpHBvj82UPWYR/aiuKCfUt9ZKCviJfuE188yBQpffdm4CXt
MNEWkkUbvAZgfkGUi0JoEg32IKPYTTmFxplkFNe6jRRHmMKauqr/SsOAVGEl8weeX9pwBq5xxsrV
9qtQ85+D1fWx+9/a508b/SA1QZzAadzgvWzBg3sHBztGQCdtsGk8WCYicT5+HamybtfsjDxk6lWn
rxD+woC558T9pg1cJTGpDfPcaY5EfHUCCfmEKHewb+ScVoKnQav/zfaMagZM9PhnEvNQzJQZGN4r
OHp6CI521Qw42dIjBRIH3yjsaW0rPIYwtOOdkRd03dqcKNbq135b6shlsApLBlHYvVtdUOleV/g0
bK8NOXA6fcbdhwOREOeHF6lW38WpAb4iOqrsT1vzh7oj6ZHV/Xwv94Fj4cEnopZ02etlIfB/GoZY
jVCxs+gBV32J2jvneU7qo+6SQ+p20fOH1VszgcY/1qHsCWgqT4rdYfzQ36gGXaZQ51LZm6poZJt7
j+Xgge+geWJ1H8LlYoNxixRgrYkUn/99un3wVyJ3+X47FsnpuChVa4Dsgh8Kv3NjcaPAOemzWus+
lJ6xRpwMj83doeRQRSxk9bBIOSed0QOP3hAznO0HuhqcMPOeleRxM+tmH13YWxMLFUVQZtm27Ukm
Eq0PY62yrRHcXzd/5NPLORketyXFdzT5dfD6JIZTJ48Zzi4fCtxRLZtA0hpwuIHPzZfqPmtfcwIM
w6510QPerqoDW4BYU0yT1FvsmNWYj+0mVS42EK4R44M0yGMAT3ojubSn2+t9R4HeKImSXTc+wwFi
ckHzt93tqU6bqIOmrr/bGm64TtHN/ZwiWhUb8arthabSmqjQtUzi0CqTcNQkww5HYm7lx13q78Fk
guD/pwu8yAuBZ4iELXNWbNGrMabkv3AqSFSHZAbdOETUe7PKtNbup86hT3DLg97QljDsRnf2QHtX
YENnrB4zWMwabrr9RBjWcTjlsVoPTB5cZZZ55GtQUACs0n8mNmV1xv4yfO/dR7CKfVW8r/z6BtPt
Xx4kAjyR+sa5Hav1an90vbX3OyKHCnQF1ZF7zoRgfeBo0hpRBwlHS26WnvFq/vEVFg8wc7t40O9S
DhI8dBafwO4bMd72Nijf6GTXwCU1cnIQvf2f+w8B66qlzgaKzR2G1mHEj9+gKZEAUBH1DURsDPnH
AR6zIEPhtFhoGUJXCnCjKIrQloJMhOnbj6KgYpUfrAoWKr9Xl3MEd+hDG8U5f8J5oPk8mQNBuz5B
XZgE3p+y6AHJ58NssPZEHIjWMNfqXf5V5NRA1j2RUh5nEWrnzU6yDFHtcRkRyxU2rzi8kuYKEeqg
GWDfMQ0fQU25FyoZ3vc4Fob35AJrj+dwTf9Y3J5U6Htl8hT81fn14Gu5udn/PqDWT5M/H975DoDM
QN7C7ZuQ6dDg0ynshcARjcE/Nlwk3tgrBxP3m6e7T74XZgWF6xxiuwC2ten0Z3RYK5bMbBdCN8Ur
iv/lIG4BmOFHPG9woJX8DjR5yL/J5XkEsH0qDMz+/NIBYNa9PnBHkbGUmwxeiFQ/vjUwHUgcZTGx
Z8QxaYaABlOzKCDZ/ZUSQyAwkVy1tZMWJcrawLqYrLHAYgL8b78pMCENMQFaLWkwiR87pc68jprr
g4sSUhqfqdL2rSdthewnAtrwGHFVeNa//8wwn90aRQlSjbM+Az8FlXCINkuNMgCuDjgtRVtIe2SG
bFViH7/sIMv+W0Qugw5lbOhPmehLuUjGPlwY388nprrD1R/Ps26Nev9phdro2yljaJqP8Z3nt7K2
Mq3wg54m2xaEWI8sZshZiNxHIqFqc0K/NJcF8BbQ/x4I26ce11apEHblmeFC5aCD9y2wLbMEUjNV
6SdUctA9YejMmb+HdyKCOSHTKmyyFCMHKD8oKtmVmJJzWZ6OnANiF7wPbHkLPQOJeCVjW98mqjmI
BUHQgCNuPh/pb8pWrCzhQa7jf8BKKPbkj2JTSaZSiE0JdymoX9QqVVXkzpOB0Yw2qZmuNbitylbN
pzCG3HPb11qFyLFVisMUoztyH6/GXMin+/BRUQwu2lmszSaikf0uUiaWDzwgQE4+fZx1W/SWnst2
pM98Uilj1v/px9FZw8uZclEnJ4V0lexJ2SGQI2Z8zb40naO5ZbsQMymHTdQNstRMjAzFWsSHImPF
OPx+LiSypotj6sAD3fbH8ixx8EU9fi/oy00sMzqsyMScXDVy3tSAlDlpURRjnkRKbsl8+lLPyHlI
xKmkHMAxGrAemHeYAteFMSmlbh2lnZaae5LOIsqE6n/51M/ymPqyKjCnhDkJTtIZnu8cbw4M++dA
rIqpc0WlP4HTgRnxWYuVuv9/fs73rye5zq7A3ncVMKcSOliUHVbYGZdHtzT+Y3/w2QD9tgkW5ulQ
1kMXkGGdieIJh9ATzqOePWEKAj4TLrVVLO/PDEr1zo2v9LTu+nmwIsnY+N5SefSnqGqpikTuglC7
u/jK1CoQ6hVIRjKOwonhHMysFmroivFU7Hw1xQTmaCnqwFcsJXAVhOpGwvg2tcb0eq8oi5e4QlbH
Uu/Ff7XaR5dAgPjUJNkjjayKhvK0i+h0/susnA9DVaWfaaBLb2J/eTqFAMh53Rf7cRYkm43P2/Tr
YTN0qJMA8RKmY90g7knDG3YwiGYYkTwh4b1HAI0pCcsFxLbmiZI9HExhWBg1Q1NApvpdM85hyLH0
BBXdL0GQUuJvjRAZjKxI/uFDajpkhZH9aWDHaFQb/izfWTwVha3JWuLmnRZSoXSDHlPn+qdkWbQn
Ue1wuQSu4GiA8iuUr/Z5Gkyhzn8Ftz+tnTlwnuzJTiA9531Zu+f/5D14DgWN6RC2oB/TZV2ZTsRL
2sg7k6EMHEyAm0yt7+QQntxBXHD+QCjYH/CkD46dlxmZSeIkRpDIr3lX2tSz0h9MS8zaMBDW6NuR
r1dK83odcV9nG8QcOpbI04SenJcpwHdxpaDWHCEl1OkKPAyaPGRNK1miwBNCmbr1YPqKSM0D3Bww
ZYKs9gbcqY35ZIE0a70XJHz3NiPogrQ7cVfdqO0YvWHYS7O8E09a1kpBQuRUEVTwoZKsrj/Y8OgL
9OhFVmvGfyCUJJe5wnKh0FVGzy7ys5Vr6aiF1utSsp4HIDm9AZ7h+pQevKbWnKfJhm6lhDokGLbF
FxfWqTq+Z8fuE8EcIXXXZckJNJfMWcblkpH4dpAjfnN8sX1WPViDENOT/30D+THUoV6QtlC3hZpd
sN0l9FdzABVux4hSbcTPWpnZ9YEHxi35g4b2+EXJcejrtDIFpjAS8EnoJL45jjs7C+AWiMYTh/f3
pp05XjqxEzCzDkncgq8dc9YKKr5GhuqEDiZedFa8KQ/ieb5ctG5vbYwegGc2p/GHwpSGl/Qc2J6U
viBPAsNI5557up/94/KL0ghlNEr+vhUWMLbTKDv9kNwGc1XXMF4BsN4FJvtldNllDcyUyqEiD0tx
ZqdTY5B97G1MUEeLIl6oGjyEjaicBmF+z2243D1LNbb77EdiIsTQL8ZySeBF8rUT+oD5wvbmOGJU
q9juwRwiRBy/2jd29RebzcYs4BhDkU0EZdOMqQCDWmkZ/ZqBH/8cg/OBtDFo9g7Y2t87EkuhTwb5
rynBnKbhVMYYy1O2s5lMd5fdqdLzgvKdwGgM9+LvYpobFQtHGDMvJtu0YewjtB1L09xxUH+rcLPM
gddukquGTPbUtYxRuFjizYSPo26Uycvjyg23PCGhtAb1hkwRX8Wc67F2sOgkTnsWNqEzo/RORKux
Jb4XRtsW/LY9mHsRCvsel8uqI0uCcw209ndNKROhnqDAr9HQnbbllaXEZH+VuMY5TgP7EcIC2pHa
oGQ4qt2la18G17ad0e77Nts+EJ0PY8kD9aYpiTzcpHfDZmOaB+v+DUbE/VvbzOutpGJzzPlThNC9
2JTrYxDvkWX5ftPykx/dzFkxHWnkjWmkWsPd4FQnmCz+kP8yZmgmayPKatAPmJMkVSZIaIQR8V9k
peys8dOIg+ecYusUAsLZlTNk7uS9iXMVBlX9UkbOaHn5ARKOZ0m1oQNd0EfZPAqqwvcNc3NIexlU
BP/kR8vfVZFAq28cK3ost9e4s9hG7vcw3TY8vlqpJjWu/ujmNmZK0Uhno3QtEyy8qEPEX5w8VCtd
UUZfmxxXIktxWJuvwFoen3SKI3zp45SZ1zUJjy4dJ3DNzzzfuAc72+BzFyd9vgEQAnzffHrMtQCT
VfnC5ShRbd73P2z8COIn4Z1JLQfJYcGPCLXTNltXWL0j7BmOjNql42BVVEL8hNAXVJXQDhLmHhGy
Q2qPJ27CzFWWAe3DKKIGFSFk+k431I1osWTsE4FSsOmYiKop2nQKQTHhPgu6ZWMOz4mXZzDQBpqX
o6AGaOeWPwTKSojzrccNTXD0FnTWn4m2ieU1PPv5O5LqeoF7271G1UvK1aLQX45vQF89GZAv6wug
I5wFg7GeaxYBa4Ht5AwNn9434C9+3RcxOD4IfrDTdzj012Gxdj/JXSkbOvgtYeYulRk1gRfaFzRA
rEaLK2ahg5+eY65V7ahPWC4bWkUcJ9tp8pArbnzNjka1APQy5It0Uk/V6/SwTtXoAAYxUOB1NUCB
V0TJrbpLpFpJ2KZbimvk7cfwjgX8YtG5y1nunAoqlFtrL+xQSYyrqRArdCnPlo/rGZS8ulUTF+vH
xWs9tFCq1H0fFI8l1gyUHWbYXOBfFCwd705XSKCzOy1T/QBtq/RgKCyWXXV0MUKAnlHpOB+1gPLN
YG8hiYyCOArqysplWR81r7fshmeJUqGa/i9Rvqceb9EQ2CCH7S+4G/J755KSNJIr86IwV+GV8Bp3
UYcDhp1ZQG+srOSv/8FwJ5ihr/ijB/u5lvPZk3c3k2ZgC5tWg7tivHa83SyjfrePga4yLZNT+gZC
qy0M7Uv+sB8/ZA20ru8MQlM5TNbXDguRsEL3ovXf6F4+iH6hFrbX5o1wfyzrMKi5oKMj5P0i+rwr
RHcNevcbZQp/XQCI1iEAT9m7dWut0CesyYlnmlIdRE+XZZbU79m4I9dI/06XUii1nrY+hVEoWGMZ
UOdwwJm4WkmiNikt14ChtugPwBgsdPzYcGiJf1WHAjIelOoDtOwqcJC24K3pRxWOBSUFk8J7i2NF
I5shgkU3wBTZCzuX+ZRzErg3HnnCvPI5keJhg+v3VMj/I4VpplIl0hWDiWPGu04m9UJ4VhXkGPM5
Pwio+PFblf/VE1Yx7O5TjdtdcBh9MHEVxDOeyGct06TCUbVzuPCaTwerg690WNHlDqjrOrq0T8hF
YJ0P1WCD4jys3fYOL93qG8bMelKmfQ+jvm4/AYbuVL//6ukGmF6/YUuzdFpKR9oyACy0JztCV+c3
8BNFpvtvWwnJf4+scjouNo4Dqx7KwSsliK03br9psnichu0imp6wxR4Wwbpd78/0pUaGLCCSNe82
2WD5d+Dwykv8h6ezEZ/rU0yy8EkQwgk2R6cTvEZ7Q/f1UKtBXDzohrZVUlsFLHwpIbUceqZ6YJtY
eAcCQhnTgQqB4njhJmv5EP9ASKyb9Z2gnKkOc4Rd3TE3rb+/RaESWHTFVbIXBkaar3c9KuMwSFG6
ULAmKjIy+pGozjA73FZd0H6MBulPbSAV2OxEO8oTd+RaW719gWRUhGkgQH19bOI0RsjQXAaSECEr
kkBtDINBnQhrFzSjtv/rgBtBBByOEl5mhwUsT9vqSoo/i0/PfEZprLdK7Yiq+ffqMAswIwN1Pehz
//wZeqYrW5SAtWP8dHlKFtEEDeI88iTlhy5TEtLfbpj40ha39xfy6eP33jaPtp93oakmfjYXEhuw
6POcGIOsENHO1AHL/t+zCrrLyJdTwoM7ouHQ2BAHEKUXtLaH+fplOf0S+0pgEtHQavDOM6sz6r/o
YxeVio8GgWVJeXHT/Sh0FZsV5E6Yw/TLHCfpgeL70buT6eNvlMdiawSr4xI41E5Ys8pnoq+V9Ri/
Q7DaFloMQZZ/qhEsbSMhwLjoXG1xE9NOLDZ20r7mI6J2Cqofm6C87o6jVGcY5BOSnuknGpbvTyhX
UqQKYVekwf/qrGXImcvTODBEsMczB3TFR9adKR1oNvS67FhVdeJ67vs5FRqkh3h/ko/r1gE4BVIc
Le4jppLhpg/htSvOQUkIavOn0R3R7Jdsi3O6chIqIjO+HJV/u0twnTvqxLNrjbTxEZ1G0xPzE5S6
V3e6ld82Pu9XbvGOMzdokJOuc39GONNvN4BYNnBXooW65oGSB23OSM/lZtXjBddBcjEy8lbl3Rmj
coFrza1vmzsnJdQ1xAo/DvCXEcB0IiL5yIZ3s9Ewsj7neO9a/xpO5WSNC15fvGtzKwFplzIDteqm
vItDlMRxl07B7oyaoSVkUzaAMaez1o104Gr9pYizqmea90yXbFVuDmJToRgIHER5NipAWKzRiXqk
trFhyn+cuJ1EAOZVnVDHokZ7yIFQq+ZeQHs34mUwC4qwQpbwgmDp9ACNG9HQ+Fb/QaJTf1LkVZp3
NsQIgVyIYeedv+cInJrxMgWup7NFViURr6fofNGfsADA/07K1k5wyS6Vfp0Eb32hQpkCr2nhFl4h
3jaqp+JFOYhScxaHSWEoIkQ45pADVx3e9jmUHMYW3SRRMyn+hFJaFAiULCcG+edJqYOulhuyeroY
QoXXVZCzADay4GUif3KNrt2Zs0uuMstWCzNbF20LGXdLbLKmsc7KBlyszivQQDCQFl5YbIuDAx2k
q0IZ4t/1ozwk4k0+DKuQS1gftZ8kAYhMqA4ql6/GnlZkrfVDyVcLnq+o81G/oBB3s2T2Eja47y0T
vTpe6GmqdeX/OrwULTEt6eTiJgYpe+zx+8FPp8hmUOiwESdCN9SGWolMDbrYCVblot+x70mTgE6K
Gmiv/iNPmRt3HP8ZNKVsRwrIsRHLObwcmwz4z+vIOhu7guQXau9fNQgZLRM+IfkjPgLD5HKB0em+
YdT5vf+hmlvVA0e8HBdpRG+R/HcddWw5eofk6dvblyoLrDEFRQPCCxR9bgRk6Ms5Gc3SQxgCRXzn
r5NF9H5KlhRjf4fYlfDDuao77uSZy7yU4gEfX0dkUyrFL1ncgWQ6XFOkFDYPFkU+lk/h/G5S9tzN
KyjrVLJjkwBU6uVaGVDjvOCIJie3GBIZpriV8KMJoPiFCK0TmKBx3Nm1PN1JA64cC1b7tSrSFRss
kZksc0N4KDZkg0r1quEU6b0YixqQOakelHpn00zozrfB9DBI2ShlGFLj57wFv3JP0R4wiZ5J+lLL
N3UX1Wcc7fFtVm18iY7qkjvdfG7nAiqoKsYUTodUl+BQP4r4v78ahW9bqfyqdJeCAGDNV3Vl3DKh
3onxrwrEmtbcte+PIZHeYhX9FIMUigQ/zcxiVTgNkP2OEA+xy0MqZlWRfS4GddqSAfM/2hDdk3D2
gmT6ofsr9jEFLxyVBpR9sDJWeqEWq5RBYY78vkQ1vKsyLvwcVhWxjQO6fO7VOqNO1IjrNJ2wrwsd
ugJKv8I46FFMwHZDHIN7d1yOhRHneJ7rwbvvida+cnK1pfmN63ADOGCTfgLyKlilTPAcT6KM0WMB
5v/YeeP40f2avx1TNYonK+oh+5AzJ5uFNdIXJjEP0+N78bCV12SdFL2NkoDHg+jU8ZM6pNceFhJJ
AakvThfN53VEJbItp6STxR5tUD3QDIKKHwq0u6d+VQ0yrBihWGXcyYfZOEH8P8EeZssYsa9xvuic
DNdqH2E3gfy+uZ46ykGkChKDMvv8RuoR5SvBdwarlOjzQezJj8a3RUUOlmKMI6T+finmZaRyiMwg
YHspviBXpR4p1tf63UJoyN8XFOTxh25hz5T8KISvwHFhlWIETyexuXcgVG+JfM+EnNLqg7Fv9U6b
ThGz01dQFr6H8II6wefD3fxWTA7UM1tCVOret7GVN2yTLgST4fAR+1XpUWsYKVc634oOHOb1Gkrj
fMm6ioHMZJLDGaAqUcCT6bKG0kRLhPN5l3L6lCa/HDM54X1a5a2JbUgs9NyeQwL4IQuQbWMG3Y6w
DKIbe2yI5MqwqSadR1CKuuQLQoBhfXrNozRHqnmmy2MynFCKDbmU4PlNJA+uv3LQC8A5uA/8snyT
UMJVwMZ3vFSH3hQMaH/owhFYJjGOdgnCg27MTqRyfdFVEuCcc/Le+hx2D5L8geyFr4+UQE/5nAgh
8y93ltHApfQStFlorJQvFIMhuKCaY71QtdLkR61T445rKsIpZEzWtt1B92xnk7QvwfFUgsALb4YP
1KorfaFDA+51U1ycWSwCdG2ly4wJ3C5hzVv2xZGAHv+M8ItqmQuYevRE+SIrKHzPMV+4qQt/NRJR
PrfnNbystbB/TmI376kz+AfbJuL93POYK4NLirJFx2Z/0YP0Ajti+ABaZeuot/pQ23XpkcSwNym0
psUotkEz7StJeqYV72eYEDMKb96wPp0bmF5dNoCMKUpuk0LMeNMnfooUV1eNnX3gdOslWx9YkI8O
nrP8id57SmLnaO6LRMFH4wAPqZ0+oAmfEZZJZMGetOvnYIS0lnMbP/CQOrXueLNtwTy/nx7QdgNT
gpkHE5UrBgY3MsoW/E+N4MYbUh7FMWs+Ks9RDQYHnH9qVHIoA7LbSOtIr5q26PpD98eIp9aeb7m/
FKsPmRogG1tYOpiAhjNRHZZ0kYdT38oqwFz9i+Y4jY7zdi7pefdLrTWNozczJJ8Hoy9fdwURug8V
5CtAheWXE7YbZt/1K//dV9xo37iybYx6FLOfQkKOeYbx/6o/2pIRVmKhRVNffryOEgT6GxYGBFd5
Ir2tdCn61v1axszT2/Ai12ZGsnUOfyMjpWoGcbaiigg7ARIqcp0eGpmQpom3HmxaQelwQSonIJpC
F3V/sOTaO/fMrezL3C0pLbMEvS4Q6OIWpwYRV4fmLq3kq6Ve+IxEKuFHAmmcNm8qZHwIx37V2gx/
NcxDJjZbpKZ4kxTDVdFnBYKgNGPngX/UkyrSmbAmA6pVEcg8rtjS6g1EVVrx46Ra8sMg9VbUV4J5
r2OHABGO1K5V2H+Chl+jwyGq7fWcgwHzqr5Owvd4l4WLZIxd4LXkh5Itkn1VFNmoR+y7Ul0cthfH
XumqQZ/jUnPycTas60nfMe3wno/wff7NEmZLAnmUFw/JJt4PJiBF1ScfskzY+lT1MfLP2p1CBKNx
r5i8vhA9jCjd7oh1yGSdppjLDy052u+2LUSSEcp1wxWgEW08SGu9eCOVgFLWq2EWSehp4aZIE+aY
qhmSy01l2IfQIKGVOAwlccbVxyb+u+oXzCdkiXc4BOMk7hl5ZMx/5qPEsbg+hCX0GSHaUgp7ZmrY
HBPf88hmMIn6kxrj1j5rQIWzknE621kxN4Fy8OPS0zhPOlLsyR+LkBda+LcE9FG5PvTCTA8gzbwk
XH/1CUgfoMdBM8q6RqSQPRtNOdXrGYm/gTknxYT310INfKUUH1A0VIZIai6lmUzv8E0U1pOvjyXn
A/ndscHVBcWUXNMiTMoZNGo6kUpb+8vlu1jd25yFgymhpbntce59LaRagDFaaWotvaOTGQrj2m8e
zYE1ha8BXrOgx+k2fnXBNvPpXRTmwWdpbt/XmkPwOuoce0fEmsDnaInCIGEtqB2hM9TU+ay+Qr89
uhVL/X0nLvFREhjWeR+D7vi+Q282QyBfbnUjnZkeI5aojE25xlFyLTUSrEy8yMdBluwHRMZ7vkBh
jpLieLEeNuBE1zqvecz9zVGfMeIms7J1/O84X3KQHXHFUB1yx2YraevGpkL9CYyB5sPMwy/gWJ4i
MC+irhZMTiAEYejV5DFea8mRpVu4qYHCsHNYi/4vpZfs8iCY+Ke7DPHFUaKH2mRLRMlWDpNXkIPZ
GbrjKY5hcPOPQkwqcP8ViEWkz5g12koo2W6O8K1L3yLFVRq9fRwuelOx3kiMqTMCfSGwXbIP7i8G
COtmMpK4zEw4mk5qOrDX5G7W13LGA5BBX0qzEFIJpafP8Big2cosFOLm6xkFpYzOqyd5QZjn4aSb
LtpQ/t6TpN48hIew7tduHVwVSHilXDdCqgcAxkIap+aX6wL3Y8iNNARUm7PhAhOOwCofwKgDUE8M
JcENJCEE/ThRTweUf66S8Z06gPYEaQYO0TWxrtgcMoZ11B5lZ9L2b52HVWc8X/kg4iLvjDctHrT9
Hm4+FfVf0KqcnZ+tFA8/zfsAIEFUMPA2vjRiDMxVexPBEIPtMCX3VyeU1zvOA56TVu6Y/q65ew5n
ny+j8LckQoBEypC7Ke0GlJaJLU8ViHdMdWx7x1r3So51pwMA3N/x9Yb8UUhUx1qv8RXQcz0bAH03
xd2u0OjRBHI9ufNshgfeMd/OrjBFlyk3A+JaS9ZkWOX8oY7f3kcVhsZ6FiVNP4c+YA3tIPquJxlW
C5Up7f97jFuXDF0E8Z92fWIgBpj62294DBat5h/IQj+MVQvADI9NRkNqaSVAqoxDs1hK4XisZGRz
89wD7EVqmqUMtXgnJp+dOIjCGjj85RUZq2VNA0w2T7s1umRim92rSE3k/D2IWJvb3u8MgNLUqVhm
djkVL1ttUx2VemS3o7j9awsULrHo8ux+pu/PBJuRPs19XabDjm5MI0F2gbXcX3Oyp3V1z3gEFzbc
AusfQoQVMCHBwCpTXFTVcqbIoxZS4DhM+yEbH7qJlI2vkFUu9sMHSTqPvhBi6pefzJQentszDYXn
XC7xi1RW9d/3QdWHZe1nCnBuu+qnEsUDkEgqwlMUSJSZpNv4ry9lbyFYRpnmX9FeGOhLKD2nKfh0
mr9qGkn1z3A/OLCQn4m0aM1haw95STHFw9bYVscpY0D5zkL6n/DjW/CEVQR9w9/TjFH24AMoy9+p
em788bEUfjXr1AowjyixXxZyhwxYp8Cw6e5NkuoeJScv2RM25G1BvfHiYR7sKCjwqpATvBKceW7w
HqSLk0ACcH6mYmYTvvUhdgzz10gK8ui3wiTDhDMfchy1CfILMrPguAphLYyFMP2utfU63tntrrMD
fcsxmwNdGZqDshwkO6HPZbZwI4xXVNixtVPwR7VJ02PM1trJTRpgl+8Yb/SbMUbeJu96LlaCmyoE
baRu6eqyHW636G5ybCaxdBobnQKlJLQ5BrcwKw80aDPPCTNWhkIfy5BqEamebyBt9qcypMs96P37
sF+OmL359YpetLOP/mkPohrka/HxHpOWMAsJQ7+uPGTwgEZeIIEGpeWgbFjwQX8U7qa8ROuNKIzi
jSNUcVrtI6zEk4wZpC58I7Uv2UeAOkCzb6sNPNKOQfM6Qo77ug2waz1+BrsLt74vgWfb4dROnkbM
IPzmo425Sz0d7z9ycgdiUYEnSK309/6w9Y5HHyBewA+qMtz1N38EChSWco0ssm1BmIb+Mt/TrA6p
VpFv6vnlvFu4WF0yaqCpxGRL4fZTBGc7ZobRoNq7tk4k0NUzt1/4Uwi3a3p/tGddKvWZzKZpDEBy
+tt8o3dA/a4CaeBe7nUME/hPzPk0wRepC4CJ8HkKre9RUpjx9T3ZHq25sg3HW5lNnhqE8lXTOZOU
oJJS1qiEy4OhJzMhXHyVY9COUC9yKaV+3JzQA6YyQDsm3Nze9q9D68RYLT7Wa8GJEBpASUFfOZ/k
rHh7HTlTWBnfynrL8ZMZvoLTWLPsKhLRPOrxzungIx5xhJI7WvAn9cGVmr1PKzSqrIqvSNyC5ffx
ZnBt6paCBwdWRUJRVLa1ZtSaDOFnW2xpEZrCwgrk8BN365LUhYe73qaKkyJZEtwW2lkam7omNt8m
sS2b5eRqaV3YP7pjB/dMRXL0YLJNKB28hv8bA1fM3hOlR7QSdL2XzgDbCDeaSARuOB2uH+U8fb5m
BRUvZy5IR98bx0CShC0MdC1HT9EXpqmUuuV7hKVjbLVbMlf38vs3M/wspeDh1KvR0NZonIZpd3mK
TAHUl1Ckt/9u2hIyB0fTQ9l/t4aQurkPFlZrZa17RA5tg6lSY5Tae7faLEEQ1epb952VRgTJMgC1
OL3ttFunwMmhOLCd3Y1sWyPChmPUc0HFoobmBs/eUXPD0bot8eOULlSD2wekEgXVrTTppZwwm58P
ETq0Q/sfE+V5XcOyPs57P8jpwJQpV3JvpZY5XjFrqEacxGx5h+bQ3onzXQCe6g9hjuA7b5f/0hQT
gt+vjyzVwmq4FjGWUkvjMEQwaA1m5ThocjLjnV0ze4rmG/qpqfAH+6TTQDv01u+6EeFfxwwAR5KC
7bgmk5YSaI8eAIUmvsvVjM9vrNtyabRXoCEX+efRsWVV6gRxaXZtlSxFz3Kj5tm9EtpWbMmjspVJ
3AHU0+V4Ko5EcNDZ4l4w9n6Kw2jnr+WZMKJSBNkNRpHIM7gm92/xUCkmyb4HEHuvmGDqycY227Uo
iAmzaM+cj8aoq3sqCuQ1sHsTzIVUrggfYCofPPXiKsq148GUiDcHKl4jCi04CJG4g1fda339C/s/
MKgiZFemCE+mV6xUNt32q+H1oEtZh36K4ENF6cx/SDMWjLsQ6lzDs13bh4pINkkTVtq4G8mrAj4m
cib8639XhixFO/obfqvmFGJ/WtjRRWQSeIqi3wnVOXCqpb7ZDkd3sy3LjlQx7uEDT5eAwlAdvAcv
lE68iKfh5yO2PObzm6j4RrqoAP0QnnZiOqn/0haAn8N5aydCt6V6Cvb9mCn2cipPPSc1Bd8qee1j
oXQEct+V6l8pKX7NORoIw88FYSJyfT8qikeEf3qZcW/e0swutza3yyOggqaa663LlcJn7B50KjeH
/TSkdbVmUnYaewyoDytiW82OZUbn2qx32fgP4bwb8Wn5moTEsATMnlcuUGv8tmVVAYF0rR/1AqvJ
aH0nEAwCH9AMUCTzBOAsoW/JDRcwHgSB403mnQzstc/fCMfHuFR+6NHz07N3NJT51ISwQfo/5Qak
fUt6/s22IQx0FPBKImWvYVkpEVe8h6FHnSVNvuc1YQpttTr3E0YEMRoNrxiWMDrAEa+IPu07MgiD
IRu1PDh4QFXstHJ25Ss9m0DiEDAfhl/D8xgFfvdNB+cm8o/95iXILcVBv8PEMgkkBCTz/fbVdD9R
aCwEjeVzq5zXDZ2HrTgVHPnvG4yl8s8XdLuMz2ujNS/WiyBxZb2pdEtCBaF4X5Q7WCCzdSFC0TD6
c57UJBFPtvKxOs1nAKJvJ9x+y6LUWasiuirqh/1NXjz6E620HsLv96XpbdGwTt380WJYUfBqGxQN
4XB2rsDh0AL8VDpPx9qy7p+CMp3bDxNVNzVIrJnrQ4xvaEC5UpQQ/MIOfw3C57RstXlTEmKR+2Ni
R5nIHFH7WlTfFCaQJ3GMoe+M1dyPH4dLpfJmw0DGmBdvmqV9OdyiDzMzYI+631l2uE7hPAx9YYIH
KvnKmBRzuw8BDYQIq1f7z0WVsa2hSVZ1UaBx9ILElh6hlN4UIzITtvXBxUgRgE5iVojjlQ3RWY68
8K30WQtWFXoQMd97afmnECQPtoOASJpAAXWeMwDSWsIlbhE06j3QbIhxBBamhJDVuK5O41lMiCuv
JPQWzemtEqRXdqxjWcp2rSALcsnP6swKIVbHIOhuegNJm2Wz14hHxSCaXi9ok9LjO1327id4N/t1
ToODe7doETerSSPXJS3vt0j1avTjPw49Ho0pt3rN4yRDa90drng2+HKRUm/RHbqJI9EUDqCrxfJy
ozNSD6YPJ7LuKbz+v+z82QN7XmEHyGt095czBxotJD0SM7KY4TGF4y50dIMWiRkqWSX8qStEcKf3
tIV7+nScpotWr75jGFTujN26Xrcmke9uiekv+V3U+dgf5FQXpg3fWyHfGsgqMf+yAQ5MyFf5bCBj
HjFdm2o5b00vS/8uzGPjW7tgRbdDZI1bWsRn23ZZebcMnyrVvoxvE5HAuLdsG/HpBFXX7ro0/cQL
bw9CiG6kcrV9wZoLszKZGkhwGgn7GOs0ra/KBRInfRiuVHSL+IDj9XCRuB8IJRyWZeCX4TbSVI6f
5Kgl3y8uJ4WNGP8SANVkj4aeTUOaclNXNDiE//myu4ujMx+Ha9SV/WjwHwsf6O9y/oTfQtYPZBsP
ZYB0O2r3Z1O6Gf1U3p1bLIpkg1sPGfu8dEi53oOFcEMXVE9Q+D4deUsqq4FqfAa2vwaphJ3fFGoQ
3pmorbiyuE+61snS1VTDo5mNu1FnFOZHtxsRqNmq1ESMIYf/ueGgKznh6NwYlnS1MApLjt8z0PWI
3zd3Qr9KZAB9RTQaaBMsPRdCUeBRDX+1WuDWq2QcVvKVqKPv2C3MQ1LW2J+jDT6/yCiToEoXaGRp
knRnT2IlF7DWCzWAr5MHMoHyeiZcp5QJNr5Ld3y9CokAtkb0NDFTGIJKZsoq2ymJxhr6NUlyGftu
4dT0tjANc3EAV8sHr9m+c+JnUdQ4bsmDmjjV4QTDbS7pn/PJnUzArVOIuNVzDS1hF+mnxKIQJ2Bl
SpmauiWiqTaB/sv9hpO/cLdAOa7CYKNCDLNaCBTyxfjB33aGX8/F5swyXHYgdm9vP5183EC69oOc
NRjtuBFutRWDYTg+tr188/UYtLRyyBw2maEkhVT/7qtnCyNpD3BnLi19F9g0VlqXcCgy3SHd6yVg
toFrJrqX668+e4Nrsm72kDCZ5QX1HbNpc0U78FG4cFIITBNsCUtehysLHwyi2UnXughs3nuh4LRg
zM65tbhmmfL3CNbzOu8yISI/DwO1TZr/2AXumUhMSH3lkkLnxPzJDzhtMsoy1acIW7+Sveb1E5+S
AKjQHpIMahRHrPL4dOI7+hf8o/4tcoeFAuw3aOO9bOOkC1mbyCPqWuiCsEBxagbZRpCBDmleCP4a
v4hr9ZoBAnfrtmXK7Zbeqe9hH2Z7r66pLbDw8XZgE4Go3j2q7AS3rPyttDwNiCzmJNb6qfkiiLZB
fqAkNhkn5HXfOiFRnPO9t/52EJMM54HbJXi29PhfBhEoHtAf21cu5YDdo5AcZ6mX/bgyn8/TXSgw
DYKti5zbEygE778x5KqyKPn8duksydZnz7XkzSObh5P0Bh3uSikV3x7DsBpQgXJisw0eJwFMbVHJ
5D3DAV9KDxVMi90xqpl1eOfN1/HY25fPDUtR07hmKQECQeeXsVJnWkwUL2oyWHYQyn6WnQ8kLSMi
K+bIfl6uJ5jgeABZ/Jm/q5xO/0iWxuq2qFvy8afV0NoETTomq9mFxiPTmisT6qzjgmD5tEy0lRZV
dTIR9SQ8dTOjjzyuMB8JXV2a8N0qs9/1E0khXzfkpbiDZQ/kPLGq7ydLtbWjmwbB4U+8xuDk0El5
U31S8xcLq5cwICxiKxFB4ssarvQBYQIi8tgJ1icX0r3xwjsn66d3WE9uFNkKp97k63pNePojE1Wc
3bk2QQqxtKc2VXxdy5OeHFbpuKVU4aiUgrwnmHP2Mp/zWGh4LHNdqViFxal6tGc0sK1SkvsAxhtB
43v6Aty8IQp8Ah8BPzLKogKz4FYLDsjlJIidQR+N5K26NqJDt+w9oQFaGtwMiHFxiXUsvcD70PP5
0UdOvoBwx/0dXLoT5bYqk9i2xF8hKXWlN1jhmoqArK/HYk/V5x5dOssAQ39k/t0YoIeFZwVQutRt
CGech1vE1XAk8yPELwTdXAMIm/GEt3b6YRAOYTKDcQMEUipedkHc/IlX8ujoyzsNTEcBIOoeUv4c
CHVybzix0EyE/e+/X8D0PXxhAbO72XU1cwM5LlJfcdRv5bkazHMbeRbK0U/NrM3nmQqqoUuiHOdr
WRJgqglBMtYDlg8ghsV6SX6lC8sLOr7Uw7Nv5K8WA7wg5fa08GQLRREOpodiYCIWJ5LtJH2CpjEo
4ImGXRrAIKshbi18GiXasqrzaaqb9pwX+Pdeb8m0L/Gpj5cGOv9Lny2s+ccRvjJdbkgCaTj1kBoB
gSOk/EK/nwsRJapXokZxv87YqbyCnjEg/ndt1Y+/V2beGytYMWpGVPBTACfxH0sGEtxDDEyxO45a
5l1QO+bNuMlYGM202yR8pWrUKGFHOvtI4YsB1h3Rpn5bh1FIgrdu+6QjxIFL/6A0uBdlDncEgR5w
BAg0yZsb91ISDSsDtLCJGZpBQA0Cs6RsZofDHae+wSTikSqwYmjRydKcEP3l+jeMgVCAkNWppRZS
40Df0zS9t5Mhxlp6obH65IUZPUSLdR+yY6ZmmlJ4PZrc+N8Y/hMUbfYarOSgP3sj8d9wvmlg/9OU
T7uUqy7DsU27H4JvFEUTJYwp4fDup4Ep7bNoaewqKRrdVeoTIq7X20y1WAOjeP62HeIq2ms7dzU0
72WE3ncvzJzVbzrvBOpeTULmTEoPgS96zDAjw+0VyxIG/Ii4L64snNdkbkZp65FqwzCkXNflTwdi
g9wjlP1Q0Zpfu05ppaq/nyGhmWbA1/kyrkOt5/pghRfZuQdohVW1S5pUCu3M5bwWrahs6Fg8ClvM
FL4Kd5S/f82t+RapTOIfRy4pErxK9jfr0yd/p9yghNB6terrsQwmnjveDBmvopv4PpiZG+i1cfVl
1/HrCzrG6sAtD0NKr9wuegpAWXvFl9Vds2JdHvoi3u4TkIL04Rn0Cs3FD7mTFNlhhyf2zLSUldSn
leI3pAMF3yDZYe2INzws8bSU68WBITlAM5Oqy6gmdsAV/xrEeaMmcdpz6hFAquAbz8B6NUBf8jtz
MYe1A/xjOuD68BXdnUZu8/snx+XtegXjpW5FvZfEUCTkLg2rJhKAhjnfXzsFSaZZfhMp5obcCEbr
T2piEbgwjyaJY9WomsakoJL1Nd0c4weNKzAWO+FsKC1gRSQL0iQR3LzW8g942dBo+ly0mqwbi83L
oSIil26ESamU0joe9Wag4uoYMiV4hUGiNhAn1sWRu8qHW1sQ7VGWwjZlZgzrgRnTrFk7PqaV/dHi
V3t2phvkYaAlRiRMAk6SPzmKdQr6CAGSyM0LFZC4tByt0LP0s6HiBfaTEAJwTEMj26waYdfKgeEn
IVdjiruwfIzznzf6knLAvyTscw/LwKU1og9UykYS6lixDgWiOQO5Pz8rThiJOdJViTfQyEoECnuL
EHw7/2GhH9Lp6iyNffAJbrZn0jzcMpd5P4DDmNiSonjwE7W+vdhHnpSh9r10QT9sEknOxUtOXXyz
u+9V8O8v/HVd5wEOVGqDR8aq1aqZyAdEl7fZDaiI89o7G7XjrWQMfjgcOJe1LlTUtfBTIj2SKpI7
jhyBOU/Vo6lrfwrA0BS3YE2cA99jkLhz/ttZBM1S9e4p0Iciu91AXf14gBP95RaPny63rmUAh+bH
PyXa4kO1vkuiEnkFbo/y+wm/qIGah6wE7EkatFKdqwWxB9Zi11soKCsACmTiBzydr2QPOoKjd5et
8LFSsT+BUcgzP9OSTgvEkVNtnVfyZ3Pnuj2Gd0lBHUX/vP67VOcPgJ8B7G54WYL62+jtGvqKjS9h
nKeo58Kj0Wax6ILcd0pzT08m+c9BLYEs77338pZNrSL+W/iKwG038aGLmv/GWV5lLPuHj+InfmBK
YSY/YxnDpAObl8Sdz1IuzUs5Cfp5laVqLchGmjLPvylY4vuQZin65Au1vPLRiM3m8ECX9c+COnco
dNayi/W82LJmlQEnx6l/vJE7z5fEvjhaAfvGpMtYCfVCzRqq0i5p8pukCECeV49nhrKjIbwU2DEU
u47Sl07gU2k43VRjU7tLO2Q6Hx8AnJ2r5Iggnl3gghvv1XncB0Vb1MEpa60Fq7Yv1C3RsJliZbGB
u3fHEmDTNzkjnd+ZJwFPvz3bcFhmbHv1yIXGZxQy7DS5+qL74G+nsZSuFMa7tgdKFOig6YfaLomN
F8G9uISghErKpJ8FPYreEW27v4AedleOObGS/YiINnPFKJNI1/EhO1zpSRQzZQIJLp1uDEn230oh
abI/HTfmY8zf4VGi0OJ1Sn21ff/l6F7cU6uZqvSkvRMGQex1JiTslbKOwYhuOhCDyjHWs7mYr5gm
UKscCGeq65uUMDbL3Jgy9q2IEGqWwER609mrnFD56Z9mvF4TEyEvNOfm79S5e4ofoFklWFmPyHk0
m/XFqew/6EX/TgPcFY2pkviLBr55mWC2wryrWSX2w0WXtKpavNOj3q4Gj0v9bFro0r8OfPZw5CXm
TDYnk6QPAI4YSMFZGOA17iARvB2+xRynRp8pGIuHg6nOzsOnWgLswAMVOdr/eBiYcfaD+2+7qB8k
FRmiWLb4TxvyODE7Jo7THAOe2t6Pg7W4svB8eG8S2+p09/XvR0aQ9CdnLXCX/cTXdOjKCr/2YdPq
6N2IH4pUEeSbHfC0uWbuhWnia9OU4/lgCOEk7yxZlGG3jaOq84q+lQUxXO6Em1JzJJbX77nVZdR+
qI+9rUZobu2CHiZ+QV913uoUsl79OExhpIM6lUd1MZljU6o1Zd6fnFfIrmq62/YoTQjd7fa5NKRz
ChbXwnklVUQGdum4NJFieXY+Pa9qLdqN1nUyJasIi+O4D4A3oAT0eJ4+kNNmkX10nrmZmcBLS+kB
Am3Mk04uWPkKVj3oK18kKSzTjCGFhIgWdnPNR6H0uRuRf3qoNy1PC27MVlQK3ZopaWN6PnyciTgt
MPXJOwafR1OPyMVp5zeN30/u1M8WoX4iZxMmagH7F++P2U9AtNq9ik3uoTTT5XY5jT0pvwHYC2GZ
VoBLOvklMomSr7sgSuAwqNoYVX0OX7caUKY3qkg1cJE+9J7EoOjZELz1/FvxeHXXCBcpSfiEqu+Z
1j70wBn+USPIY8AwTpxziAf/XZyPdeBI7L+vdxB9HYsV+C3nhKje6C7Kl7eDXAIG/tu9g3bvVG2C
6usrIlAhU+1mnFmQBhLeraTh8pMLWjRAuzjSGHnbFKz4i3Tsn2aUr08GcJJ//RpUZdIXMJtyMXsn
IuhV4BAo3RbdLR7HNRgXujjea3coiOL2j3BoOWJJVmXpdNESUVRrUv4nxhofnrghWbEvKneSEJwJ
QByElIx5pQ7q/AmPILESnlK/BiYrflCFSPjrWbSKM1btIIz91Kc5geMvBL0m+JwezQ7/ssgHcYUm
et/c4GOspsI6SmAfXbpU/4bBbquuaAtP/T7k7yUKtaKNG0s3zibiyr4KtXQRYkneTd7c78KH/1Vo
93ZuNWt+fJCe7dgwwdJG4j5WMUXh7tw1TSkFdTge83retq+VQZurbM1pADvaHrTAdaWKVDAIi1KI
YxCHaMk0RNt5uPEZHOlLarY8EtxTWE6mDRQmhaCK8rYhmuuraEaJgGMVH2B9KdQ5xG1YxIcedotZ
ejHQynyx6Ww1j758lsw+Y+Y62gBkMRtinx2hzaH/v86VfKwr5VIE85EA/stOFwhIsBrLyMCKBcnb
xC41fhRo0s5a4k82m7XZDfX+hHEEwXU8L76Olu8Lb92uthS+wxox0/YDyvM5FXRoqY5pUZt2vMmx
+b59uF0WqYyrkD/ghiUQUg4uZ5xxoprKfOGn/ddHu2v7xqTkSSxmbXQas72EM3eXLfVVkdpPl3Go
zt8aunC93g0IbRtTysnVkukn2bXXRaDeUGPsvsopscG17m//7yaxBplIqFnYNKyiZJDUpnyS5aPu
56Ytt55NP64ut0So3GltBuudhczh0GaxUIPkkVQUZLUKXlounhNR6QHJROqR0Q9jDHektGYQp6cI
4wFmotFWlQraS4DeFwsyJRYIU2y4jVTUxyH6HZ5lrFzc5aul5A66y2J22rTGqfumhOOaYKZURf4H
ovxzGWbZ35i9Q9n3J5tJ5sox36NhsxCPhVvP+ToUAQ6vn1BXwWexe18JdoEP4Q8BL2drzMuuUBTM
FCuxu+Rpq4Sf8LJGj+vZR1sc0/Arm0Onx+mLIEM2fiaMVJquDDzdY3tdD95k6Zp1u4TW1nerFMt4
080MD2ArzmeQVjB8TVDepOjTBS/QnlZMvt1bXn9y3PmRe1Szb/pg9pKaAFXtbvJ9D2eMlxNpw85i
73H34kjNjtrNd+DPFYST9j9b7ksEHDLZTmJn0JYLbr4yASzbNP9JPFHWg0kP7mEkRs3kzFvRMV6a
a8j++JURRWHwk+Gum442pNxRNeIjZd9CQ09LeY9A9vF7gd9eJrR/DqUnfyvyQ7e4itufwg0W6ro+
JxilSQKpz9vcYaAbHjwvIhUqSi2EFMKUKpudL8j7hbHD2aiwxVaCrBb/sNXGEo6XyMFEW9d90KmJ
ciTNKdHddMnDqt4UXIymCXxHA5O74DXYRxenuuysQADcRjsm62JGIRzIppxz0Y2/hqHS9glOrwdX
weHpif2rufFzDCvWXv22oCrvidYOGI1tkGGj01VfiLl8WglCqm7ieqUIvGWRi4yq16LTr6nwhIm5
9KoUOLFWNrdaKeCkA2zxGrpEfgCuus3PANc1OSaHxuUg+syIiXF5JVz7otetSL8Shqr6wkDUP2WR
MoNhQwlVwHuhz+2ddksQYrXCBJxft9bkJ+smYLm7oRyWlIk654VObrX6SDb51VioUVYO6B84gifW
qNHKHxud7OOpVPvGo/1+4xp+wwq6Hvc2HHmDYCYg/ia2Ja9wC4B7c+kueSDC7PWvHoLHRZK1D93N
HDTv/9s1RUNVV+IV3u6hTuYY9z7rbhMca1Aipuu4bSAe+gMKxXFyKo7RuaXYolFS4ePBxVQv/Z0v
usqoxLrbTn1ylCuhb31Rsx0xqtVGDEH93g8BSqSQeKfaIFNwSsWr5H9LagXrBZ5dY3BIHPz6XxYH
9urdxsw4njQhxyHXBEHjwvLrGM5B6x58CPVdcz9g78e6B37HQ4FiiBWteEbWsVNcIULx6Az7UzzK
MvQwJ/0I5Y3AYIVZCgH3SgyJxsrQ3tXhzk0kgZsYFz6UPRZEDSMUkqTSC49ULwfhyvpnWyH+8z5Z
sU1zCxsseT4s6MIXByen6Y+iW/S3sEv0cZ4ZAuVVoi2QlywmYgIUo+MkpWhV5XXtpjqXLWWzCnUM
jyt7+JxdF2TBPDbX42wzr6/CiOGhCk0S0Rhy9+wJeQxLfWZxoOwO+1V5/J9X/s/4PY+WucJ+HzZL
dT3LMeRbZ3HTqaN1fL6jfsSX/UJA8lfM8kBH8mr2P0yLIiLQIq0bKcKgP9mX//QXvnQd7Q9GsyyR
Q88v4bCSQvQ0Gqd9ZX+s9gke3+lRRFU4PbQr3BlT6fFqenIJjE+/50J3mg8wKGGhIRx8HQmd0U6H
DFLu56TZE+NWd49/wHb4o4909TIgMBr22t9w9EaTwimUZM/Uvjfu4tQoYzq0Mm9OEtq20k8VEyMY
MWKgHchQ0qZZQ+XgF3/TOeBmjfJ8x4zVmj74tnSXgqj5uwtbec5FU5Ryo5b2EgiAvhX0Ymm22b4F
K6RVSP4H/QK5NKoUGdKE2iRa5Q8twtS7FEVTufraCaJIPh+gG2YrnNZkPFu7XAYOnQgD8Ws5hw9p
VRcffgt0ZY7T4VMZtalCuE+ULIn41upCU/f6EhK0btQy1n081QvxUbWy4gBs6hUa81EOcTyOhfeL
RqWaXUZcK5smPS38+f7YZzOtlx5b6GyfIySmSDKe+Z+J9k1N7MPUYRHgCJl8hK4RwSfa5gL/ccmw
WI0n8ijs85AOQ1BkZd+d8h5czRK9wvCMY2Y9xHcqubRBzek89ECDrlUtKikZ1h53mLfb9HGWC5Lp
K2Nzh70qNmQ+/lJL/E6l2sbd17ZEaK84Fv3Eoru4ALxBRGbvd6aA2ZR+Xf7gyv/cnQF4HGOdCFhn
qDxK0i12RCU9LD5lIIa6aGxV+yQQdifXcnAGrXhdvqLisRpnXZFF9lwnh6YAWqhmF5d17a/UbGID
rJU1zO1y/7EFZSzETcOyZBYC1cpZwEG805v+iLo29H/DYgJzHff2T9QDwVnAzhZmJJpSUpVcd/om
6uXDyaWTWTDQ1MA6h5t6rO5c2DVIdJA7AGu1OhNw6rd7RiByKUKcsNfWeDDroSiT9dL4YH9brbWC
2IeoBL3A6/awc9wXYE+toHnyw/QWelDIs/qQ4iLyNgCAyk89P1GBZwP0CdByl36XfDvyCJlnQCHS
yznGJgT5t1xz4zguKhtjLxmFqo1xW2tZwdjafJGNuuXmoyy/vA1F7+XGjGT6nr71YEdCMHbZgUWB
Iw3t+Zi/RVCdfTYPJ2iqJdB6bt/kE0lgOuFNRI90AWRoas7ApaC/ZVzLBf0LIQmNKaj+hThiCijE
6A1krsQsTdQQdn03BRHkJVDPCpjKMWfgf7gwf3xJM6NgaOdVZtf7h2DRya6tYsljuhfh6Glm58i0
1KK/ibYxXEC70YkaGy2C77Wjrhh4/tsP0jZKnFpw5q3f6t0Er8Nl5jKTAMC807nee35/uTr3qD7c
hIh3u62TsQrWKaSMJrNNiRUmCg3GyMHyYjSPkpx5S96nYSivlK6HchWDNPuvPDRUVuVf8Ioc+oCe
rogmYVqvJvMNaY6ee++xMcMly4teWz2T/ghtntKWpYcYojM6OdIFrb5H1y98arMTLWspV36oEvUO
1Em1hNPyOfYbOsJvcg7yc8StLp36PBNWm9XvrVzVpfs7RLMVjb8jHyCUksIXuW7chJEASRRlWlvD
UfRlVAJJzieFG1pCSPTW9sXEJgDvKgRt5r2pZBS5uRZaz+dGFv/KT/3DclPVLZk9dWdJzrH0Vovy
Eo5pstPcR7ML6WApaODc16os98w5CQO1ibpLCvM6fu159eDTQFIwB3g4hpJvsvQcCxrP2Hl5f2wY
b/WIMKz4mm5+qDH0uUexFFOvLhgVH/aFWUdrTfgNOsAI5LsYIvYubSCyB71TdvruuaNqY9CobVVS
d0ASj4RYoo25Qvk/vygPsIEa3+jZltcoA5tGyx1VRStxKTmVfZeZNvLdwTf+fqI7aiiNmcaj6zi4
3BoUL5G6/k9W9dz/j/HqEJ/9UHCkjGSDIB5LlAuFKmTJtZl/hGJgD7YJu4QXrP/FRHpSW7b4KkrG
+4fXHU8Cv/tZGJW8jW6DiBzaog0PpHRiAmbQDZfFdfj03qi9h/gsFdpqgaBIf79rgv2bfEgnKU9D
L/8pwYX8WvWBxXsqJ3ALvge9DRtuZvg4SctinUOn8cclAoj9/QCfb/9peXW2ulY4RIrb/iZkzECz
1yTD/8VuBk2aZzkrz7sCEeLMEdVLO8KjhfHhb7WNQ6kibroL81Y2z+tzcZZ4yy0fYnwRMSuRGlJc
/5gV+XtkjFsDM75AKFIkGKejzajDh+2PuCRqFCBXnc8CDlOI2ktKdV8+44ovZ2QMvK/8AGW8mQxv
AgTurus3rVOucKg5oonKV406q9ggvVwYoBiEkJaT7NvEW2MRdh4rcAz0Vqp9b48zu4in3zf+gTLd
N65TneAcLC4OBqAeD2AUpVP7byPDQRevW5HKRJC80y1xP0DZUhnUROHDXzaXjddCfKJWq1n6fE5A
6S/6ymz4CZ1JEbYrclrZGmohyB6SwTLAVPaerkQOYZOg5XFp726WrU+Q2LTBQFCNjUz9bmvvFSFE
zEzDETvS/eK9OGb1tp7AImc3yBZeurPTs1Hu6uvFoxpeERDLvF5gXkk2SBo3Wu04oeAGuelLiJjg
ie8fLTetvP6zwRnQe3uS/K3cj8HE96C5fFWZHTZKd2kq7D7TrAA9wTYWGcNwyO5HFdvNGyHeMu5j
4wfufJBJochLrRnvNNtGkhbFQb+irNuAn9YxtgCddLb5a1tBTM6AIGLlsW7ARXWVRbNJlLK0T2+u
MEMfeOciC+XOua+Oro/ngFgdEmMKRRaArhMKmFOe+CbKvpC0kTVXLWZVI9an5gYeDZYGnsjBlbMf
JctAi+I8Ryt6CXuJG4rtR6GFL/DAI1qG+HUaQzy5YSMWL1UAbxeGHVrZ3E/pDMIamBBgqid0cJS7
G75efQ57suzYKxBQgW0aN513WyWQPIfTq7y5msDJig/L4xD49M54CSe2TRfpZd8uSioAAwQ7K3Fh
zCbDgXlbcn0ViNQjbihB7B53oRC4tdMMO13li+6rymO0J9yhaTHGaqS/Wo4tvb8L88C3+USf3d/l
tm0crp2WQThW0wYFUvKoUI8KrBYDHHcWmjKhUHnEVApTQPM4KupZL7nPY/smmJTM4juqF0MXQJg+
unHsRJgLLw6HVnqTy2zjjdR509yM6ZTfJc7VQvmk5eH6NOcW50W9hv1q8FgTA/927uuTjBmVCvDN
P22PJzNidFaP8JSSXR+2rVqnEKGHAqDnxjRgMRBlzNVOYfSii4a92bzgBYjWs3gp6wwlVyNlPHjD
AWATJ9hAUyz+P3LHyPgUiIfpSiEtBDU7qTYgY/0fOURmfXx9/kxy472JhcIfz2tQCofm8p6hL8/K
42XAlfbNr3Dhwb4+fMnWmDw78SdlAIh1qq6jbmSLL5uQWTBdiNPeg4AOzCVzfZdAsXNR6OJYKAtC
9JjvB05ybKJC1qugmv/sI+f5G9zxUg5J0l3KY74yRKMeFy45XBouMcneNld7Bz6DemnInMOOsq7l
QJcoCrudTPXUzDbHH6DfgxVcM7T27CCXEdsrog9nvyINRoknvUMPOz9ysWYO/2eR8sJ9wOfxEjiu
QQk0CHtlLrwEet8DsAuNOk3/FAPEcdGLYPKulMMuYZkv8EXJE9M7hdvJo0s8dkm5t09RrQp9Yunw
axkAH0L1ajT15gLMJ/dv5YFQVnxllz3bKP69FFL5Ap8wpOAJDh0azTrUIOEgybyCGP9MXwgNxJx5
IzTbcVoM8qqDmy6ZcZeYbB/S4OWhChMy3IU/T1cTH/i15t6/DA1nAlzLcrD1sK+WZhOuxyQgA7Rl
3RHGNyongPaFXNieA8pui0cINEf7+YJlOGsVj5fGJqteIK5tAoTb8C4Am5r7H/MbK9QWrpZ2vy/g
MJvtsRfJLb0MFMOk58NJ4fEV6uJ/54KNDBJiveAFGjqWMSxmpmhMCTRrljdR72PGNEHcXxtXI246
Veh3gLeFWlwLlaZ5vOv1oCoZ0cG8W+zL0m5vAO4PVFF6USbfHuolm02GQb5W5ROP2rXag8VEaI5C
XnktLZYYGr5Ra8KLooGBCA8ds0T3cN9/n8iO/x1ChkwS5GulOF/QxLzauBZm+CTQdOY/7G7Laj5f
IhltDIqk7Iy+L1QqD4173YabK/kDot/Pui2R1SU3oOkVhkGIawFoR6I6hL0GZAANHoT60k/8osdi
SegjG38Wi7WXcOFfWXeFgyp319lz9/BfCXXh2ZnHP3Yux+G4QRc90nGqHB62S5tVWqZ9rEFAQeOc
dzoFRHpzVlCZCLOJ2vc/sv55Gmk+NheOTM1AWEilDgw4PglnSWkZ/VMrNsw/wmHMbhB1uvUYAzvs
rPpNA2BdK8dZKuS7fpwhtiIvJz5SInQT5OeTgEax7Q+lwVRSQd0gQld2zRbLA6Ti8bphMEgdvh9i
N/fjYRj89+snQZod810VxrvH77uEBnDIqmBYiHQnnNFrpnDMZ6wpjxqDh3gDi6fkc4sMImZV1Eyt
+bzfavUBbKcp8xKnebMHUSBGYXBaVeUx5np4I+5ZZMAuk+snYGVoME+sbzmMfMcVfCK0rbchosuD
EKKHfUvzzpEzEWx3Q9d3FvDKqcfhvhRIOEwjc8VnFgQS5x2ILQHzc5F9598RetFNrOVR7mzYI5LW
uuA7mF9iqK4uNVehprgGZSgWUmv3WoFRlt/udqw4tpwbkR10Fvezow5OjZSmfzfVmWxZ/GfBV7aN
SSkwlNC1p3Qe8Fi13vdVMvubFM+2if8RrlbKQWl5jMoYbxMUT9oihKKha7PupUaqmCDhqjvJ0zdn
bopV9pv+1qSsCJjXML27whhHvhrA+F+mIQMglAlV0qYWLYBTMptMjdExNNSxTKAvNSEezI2RSTyr
URBEJASsRYTpRzLgDTZmlqGhrPYVSvz5I6NoUhDMqSAVC/BEDDLDcaIJEDNS4vu6BwP3tD9k4Fd9
jAm9zmF2o9oMnmk1UmQ0Zzs6P9WtJl4CmwBhdl6XgC0FWo62KAepaBengrqXua9LShFWebHpOzbj
LyPkULNjqTLXzP9iFkZeH5+LcR9LuexuR9oVlQ+h1tt0VCbkV/YKt36YRqrAmBby02QLb4fMN5Fs
Ryy3dy/AhYe9FbtImcVdjJritV33MFnZwAQcLiAMgFM3a/z0koKtx+AYaymIPSg5Xk0BIdXt4vB2
ZcoT6ne3ACUyrUj2GOeCrzoPVDCEfvUAMusGSnt9LBiwqRCB0OHtBy8J7d8yFN6vkX6AkNkJFr8n
qU7npL1aFNQTKlHeKPdMlBkvV4OKMd8+/KesnQP8lzvTXz3M2GsmTGwAJMOb35B1/bgb/M/YaSx9
8hHIh82PY4tb58AFjUdt/q8Or/wbRR8XL8yLqEYLECm3Nf0eyJ2HrBEoCRqsNYcteF3lH1AkC1GR
SpB3VZGxvltaDSzviYNP7VagBqhYmP94kyIBMtLBhK5GrrnGM27dhywmx2NuPxNB2l7oZj5GTQfC
C5Cx96MlyIbTMpV9wJvZ9R7Owjv14rNgnUk/K+b+rRAmcoLaPfik9jhprqw8wUdW41ES6DpoAVAm
kvULf3bsdkRJHpfBx4jJy8hJeIYYSg8KKx+OFgNVLvAJ/0JmW4qQTKPW056+swAJcPSEv8wxIpZH
7b4aUnJDWbFltrwChdihP0Z+1oQiBSkQ78cmnRP16Mi7vcrT6Wtkn9hIhLtfOthDMMDk6Fma1RrL
grAwnecydkIx9pPJTG41PBJQfk3YVb68QKrtPxgxkY3H3qP4FJdAlX6IssmrGErGG4l9JHlUDeGk
c9SEi0MlEVfz8kSSK+dRjiIl1zGEd8zKKccAEFTnwHF/g9cOmhYq0gz1FXaEf9kBkRQ9HzkG9SEm
9wm+Ppws6D22t0qZUU6De4mkg/RSOjMlzb0/N70IPT1NQYkVWqjRL5cSNQ6dAdjxPJtZek+BoYqY
KC9Jb5Gm0Pn9+NfypPYLRxliEp8E4OKIDd/qiSBYwat8zWBoq73qUoPecKUBx1S4UJQRWHAtZVce
Gl5hKJnT9KEzN3qIlT/Bmebh4P5inXoWzBy6FlWccGwCwhCT6h3/FYpmjubmZj7IuHilaEyfPtjx
zt8CSJQAHSymX97Bs+MyjZuFfg71IRG/4CNjltPnH3EbbgMKr+la1w9pmygtURMVHw5H/vpHC1F7
08vzFqiVkBFhJ7d/Rb7JtbC0KbUFFOiRh2yXTNejl0u15FDo4lBf0hKbmZT0yhJh+9aik0p6HF+d
Fg7865A8IR6+Yy5eKgQCu/ylU+up/8jc0Ix/Txh9jMZtk+Xj1NwZc/5xlmkFQIu7iV3xz5GIq47U
61apfw7NeVzT065dX6sw/jbfd+RYpru08WlHeqtji8zINMHU4gzObO7I98qNUVhnUkxKjfMSJff2
pJzRRcU24nrTlElrLYWmrqwebCWrJr1lj59jq3EJYP0qm82oZfvpMjee37CI1bKd3qyqy2+CxS61
bczM9sa+vsAzGr3x9EvOR0GKMzVZcpKvkjkK9UIk8kp/2C+2snCVv8rgNrAcaJ0hEiFJPdlHBN5E
AHwd/+li6TVlR/E38/oTiHIX0kIFT5JRLHVdZzIUABcgsquI6KYz0K7AjmB7JucnNqs60p4L1NMy
OkyY7qQ0pypUcVe/N6OjUhqhCNgNlvEh5KWYDcfqkzT0RMfr9SPpMM9eu72sz8bONK0hLOc4gZ96
6b6W6HBWpIYCWujIf0x/16mNZImqS4ZN+trn3oJD102KHskskPWA7cx2+oX9A4q7KSqmRKU8ARgT
BGXTzflawy4aqhHKfzSvSwcc4KgJRBp5w6nZUPJvttgkwCMqAlLthlqVUliguvTc44CvJS2+Q7/c
VqiyE8bWtovrcvCr72zrYCS6o/jubxN8ZEG5qP7t11WBewk8DlZwWcIe0p/pQsr3MBp/ek8ifq4v
AmDLlKq5EKV69MtPfxB0oBzPTXisBrB/Y5joSSNQX6YA/cIH6qwoVSeWxx+PoADLDT0sz9/VmocX
EK3SbHa0s2MGq23nnUHlOBBWEDCt5+yucmDlMdSyjzJqt9MlFjJOBO480JqBPMWKsE7V5QzF0gQi
RT7sTuymur8UE3wWA9E95rN/yvNHlTp2kXoCJp7vbsbah0Xf2gt5RFlxWNNF92EHKzbrHyu9Zpg9
HC/r7a+hfnbSuCdjFM9tTt6cPz/Bpo4Dp0lmAkzkNnwz5yRw1C9nC8FspVE/q0I34lG1EvQtx+vQ
a0QT5SMN+dSbds13UVX77s++8CU89xAK2As/Xr19MF+fRzp1qMQ3Fo8i6QDL5S2c3o8mQ2BiYZCo
2groUldBm9xpVZKIqnJdA1maCy4D7fkxdPCY1R95dXB1DhU3kyaDgurs1vpXbAwqh+eD+l337Xuz
EHRFKHXndL8eZjX69D3kRHTLhQReaREZh3H2LkZttfabzmFcClkAcuvcFTD7oH8eQ0NmHyl2CDkH
Ah7cy2KMRdy00yqzCM35SRvkHjCEZb5oIlkQSve1fqgvHEPAEBURIcJEiCt2Aa08jeyw4vfIUKc2
TTE2JA2ZeNGC+MM5bV2BpNuoY04aaOh6pDRC4CkwnUXYOzoTy2gT89kXBzoqCJFfowP3B808GHSW
AdQlCfTYpt1ng5F8SGXw6cxMnYGiSEVAnBCiSRVWMwemvd2xVUUXPpKQEO/XhvaEgjyQLmvL9FLK
Xpv6uLG3XSKjvOpAAIkEl780EIkeOA0y66F6a5qtX8UQKKs2DMgLQBKwA8Y0NDPINezb67QroNW1
6beWD8up5ubMwy2XZO+tT8+xmmleBqn4qpXq1uE8KTSFtdQ1qJkspN2V8tpmRknZGsSEwrF0KSVZ
Egci/1SYQoZ0bpBDL3Jpb8emHKoa1aWNyxGx6mUjj3MAsvB2+UNmeamstDwsbqPShqIax7beAge4
rUC+FSrIZ1sOKetsOAal7u6J5Vh4zC0Qr34qzl4SxROEPNUmpPeyOCJwn2oSqyTXOmaM3MZuGGp/
ut8ihwTMWz4QzPr0XGicTZPK2ncCBGmY8HPVSiVzyYhzsAE1p50QevXkq9BXP0cKsN6PYt7cxUX9
sRRZ4uJyQnR+7VfqNIazr95h0O7uMVkoTfvIaw4t8pqx72Z1uXNHaWzEBFR3WRH3Az2XTP0nX3VF
jYosoVF0opV/KDG+OtolZSsGjxCNEF8fWIt1OLSRdzYjX2MKNxB+lZGCr+HLw0H35bMVeG2a0N/x
9V97nwb47fmQ0UOAxMwKdO0cGDQYEkrlix6W3HDO3l4xNUJlYH+MFGMYMMGo0UDoNO4C6WjP/NgA
ClP/pNwG3aJP75ckq5rZosrEiHYjdpVhC5jOobKEcHcU2ayOWtpC7B0z1zG0cXT1mPd0CGY3budI
4/ZVpvH/844cLd0iigM0dh4bgq1dHTccKqXRW8jmbEbszWKjKUwk+Dx2XNTgBq0KFkRx5CKRxbgr
TMabBHZK3tadzEepoAFknpxjagAermv8EGtrlQf6J56S0196WWYouwqPu7lYd2bx3zWMR2gtQvdt
e2OCw86Bxz6vOUOh3re63GF73+1NYAufFt99A5NSzaLVVFcOsfOG7Ldo3OyuQoj0x2guyXJPdZVH
EmHFtdKDC8tHzvIloWqLTnONr773myWjVZyt1Y0d4FZFbtuKwhWLZ5utyVw8KijfYFl9P9IuG0wc
bexVM/vUizdFC9m1qm6Yu24xNyZ4hHwepPYIT90nb6jc4IelnmHXKMPzz8Lk+ljki0jJNYnDSUK9
F44UdMFWBwvKc/GMWOAAo581aUKCW5CwzbVZmfoQce+vicBwJCnA+0c7g1SZFDONaYCuGYG0/jLF
IC35uxeHfgol8yR6tTVZUW7yJrUrO5+V4B+m2gstqGlC1zCtjIUtwmg8gDtKHM1Z7oThOMk80vAp
VgazfvmORP9jz4mbIqqJOBJc0m2v3dp1d8wMPme0StjQVH15k+ndatYwJjsGJ7Wrj/h0ce2ETsRR
E/cj5kaMFShxQqIyvzuele07B8YLbhPRijyK/GvQ80u3Sx9HrJGIQxEGmN1qmz5EXRs9QAFTiTPF
j2edOCR6ZY3hV5C/9nEAZF1+fn1rxVSYJCWT8ot1VH4THSxq+FyaoXExHa1LIBNnVJE4LK+SP6J3
Bd03weU7UfsaOhU39fiCfbg0QDM3iE6k3H/9yBD9yF2BkI1Ez1vZFc1XqvjpiMJr6DaWoOqdh2Ig
l0FnnyjxM3bPbtseg1q1vLdC08Dz9xUa+WNpCJmyQP8OKgr2gljSr4GvnVy7UCalhl3NqdHOuFdx
Ctq1sWWVWNb6iM0gnJCFdFc4zKsSetvEGkbyZvDsx5wA+DEp2tQM0PxozmfTuBSNKYUVbuKRyXJB
35bESSBKjIr9baSsCkj36OShjNikYkS84nU1lUWjjDV/gCt7UkiAdr0aw1wC1s4pwbjUeHz//lkx
w5ZMvh4d9osHgDnVDriIWWf5n9/IyFnWWW10wlKNa+X/9jq0gnKGzIFzAyCt7vxCEIUwnGZWFZJu
rKsFqVjHJllAEyF2cbYL/28rL4U4CGqdUHKfV7gmvmh7IfTkkEWRRgI/DwExYIPozOioREhbQBl6
lQT2shY+qpmKbefa+zCve5ge56JX2oa9DKdatdhmR2WhA99bL3ADXDaYX9ymnkJDEAO6JwkgbZCe
8zhvlc6lSTHgeFQta6M86SLddgjWSFbcnu4SuP61wRhpZrjtVsV3oCRQZHk0Z/J7STA26CXTMS2H
CEyDjoLKwlJCUyYZPFZvUGp8chIOZk63NFTe7hAxJPBVAdUTS6lhmPeemE2q+VW0KF1YYXSod4g9
6mYDwpoVaIF5Z24d1CRmC5z8Z3VmpCdg75EElGpl7Oz2gRZ/RLG46wkWcOWWmjUNoU5bm+FsUE6/
oIgvAHyDejkyk4VnsU0X1bZIuZChbeeHt/ZUtuPD7PHCn9yBZRh6tBVkfwNCg7PL7q0i+UqZK6f3
MF2t4AEROPrNHtbSgTzMYaZJy8BA7fSKK/yFEr2KKIccjtKe+y+Z4JlD+vo/gf8pYTC9+bkgNOgN
I/doscMpZlbZ16z3SvuNFuTS90ldf8QANi8Cuz2OGKvfwGZg2624u3GpVLZWl6Sd8tJIP8XkDZ6L
Pys7v+XEqq1DgeAHFaaPLKKP5fwLFgSdhkEgN+oth5Uwiho7oZeHDOcz6tCytbo+PiHkp9t3hnrx
aJBMMUjsaU0BaqQIoxuaCbV2goazag0++UwPiVnm8JfEiRFTnqd8cXSaV1qWEfJqmcrswLmQUNzA
ixb0Y+inAjI0/eI0IbwYs20GYVDBcX1MEc8Ed1106XI7dFGfqQGLfRRIfZ3+zR7wLPR3BYs//yk2
MaFJMcxX49ZzxnIKY8vk7LOc32Tp3nK8cy/fYSmiQPl9c+45U8bM9QaPtGszYHq8FFTc0K7F1NxR
MLAOeLuyj9PJnxiQjNhIuEtBgV7MDEYqB+xNjO/psMOuzzYjFucFVzu847peOhqKjQsP0Ej1/yqN
67/j/xsSIs6f6i7iifaLKJc0/hQrmOyQDH25nUVXNwPeJMi96WVbGBWc0bUhWLG0ioq64CieTf+T
uTFEoRH9JgqDFzxsRUjhWiAamYHIgdaJw9R8aiGWia3cJZHLFo32fL8j6Y7zccdTsYOXkD3XxbmT
CNn5KKqi3o1OdNfcpanIn1iPKYoWS8RS7lcj4uicL1D7oekGx7D0ym44ymCTPhtNrymnpy3RKDnL
MSZN0jSad/Tk010UuAVAXDzXcvFROpaPZyxnotTg2tsEeXbXHcpdw9IT5pZ33C17b/iT/GDgWjIR
qW9fDTVq+TIB3LVWn0SrVRLU3Y2dQahbe+OAZBS5zRPgfgppZLSRQdzMkbKihjXgYaYUe2JBA9SA
qcZTPdU0IjtGFxEhbPeFuWNA7wvDnPYCcz7y6TyPWvJTJbmMM+JOPWenXKmLceM1TXexcP0bGxkp
Id9crs2EF0PZeoWRfQrPSsLrq6ssOCaHx1P8oyLP0TpjZ7mQMGB69qIjrDBLYxzY2U+cWyzM3Ump
Gr0Yc4jYbQfRFELzfCye6AcTaVlKTMxhbYAbldkHym1LrW0Z8FXiM+tASFey8fDHT8PUnEu7+v0k
YZy/3j0pt//G657FXimK5Yi85dNO7tBYi1ENZSYHy75rHFsxG20EkNpMRfvKOJasahp+Y/SQ4tFV
a6pGMf0sHm9BnkoE5CGfJqPR8Ois+LhaeIJAp97XRy8f49JqRdOIcqMYggyTtHgQ3JQ3Hzb/u0+2
YkF5DZ5MWJO/lNnrc3jHlJIrJ2A9bDHy/Ki96CMbMxFSPol7UcNxJQ0d/0hPCCLINDcJSFgjUyr9
sh26wa0uhYR2pepmKW7nFQw2exKsN67OA2GbY7bKeK4b8TvCJyaBAB7Nmha4i9zRKxRRcYnauGca
UtQq8gnP8dH5Co1qVTvQX9HNJtSAskM5TTn8hzatHBcu6UScfDU4py6HM5g2Ij242qIOE9wrb05X
xIcwTAvCcu4oEgPJHgHXzHStUMQc6XJi7N3NCxqRUp5/C6Uqu12kMXMsGvh+EcXkBcv3hxlPvu2o
fIoqXXGsxn6I38WENbCF/JyDcR3u50lbhEBrb8vNXSY+GGRXaECx44rOHPKsyk4ve/jy181zFRQH
44PSCPlNDIajE5PnkdlAhVcHSf8p68C/PBsiEXTQ9n6OalYp7aVSQpYh/5HwS3YTYqUgjgNPKP2M
fxJI2j/VGM/vN/xPviVNtaVggR42PgIJ6I9BwGL9K+P5yowmfaVW6mw7lt5U5aC8vrBiWBP5m4LJ
HUF8mu5WXaGHR3DCplO0N5LdBFUjfoPoNGQ9w2jux58uZbmrNMj4QN9aOV8RpVmSLIJlN8NosrK1
u/l3M2dRFCH/tm5rl89ltJZboRRO0mi/qF2Msd/y8hJY+5Pe+RmHGV8yMCEnLKDDgKz21IvEzjS8
BbC/+enhssOtR5hR4dRZltdj40asRa952yH2JlmaNDaaPFkjKr5ZJzwvsGWo2po9jKcyLBA3futy
tZXKxZhq9yhM/gbSZM0B25uUos3H+ZFx8JwiuEPuXwkqEgmP0k+JFseNwKoQ7H9ziLOtmPndbrKv
PrMVziYZitaY/g/4yLquJV4Rh6DslBgKeBUuVSSl8G31m0ZQC5TQBItGgr6cXRfH+37NoygmU0hw
SlDCj01GvPtn3zHdtury1EWNUuPoKX3qGOBa3r1/ZLMGBT8kLpNQFHF/gmdQTU0eLgYK0r3iVxQA
3wCyGMcnUTD0KqbSUdjHwHh/o0yNhd2papl9jAlTbk5k7Bp5+10jSBcAS3rpUNQczcsuoWtN+ghq
qihREMsl7ETZAAByx4Z3Hb6zQL4kN9KMIlxAzBTSwgWXjrnawC14YILdRB8uKx0YlnVYgNaUxt3W
y8vk9ouDlwbAA9nXzgsAOulpC/KxH92h0UAfExs0LLUhb/RV1sSshPU9sEcFo8U5AVF9+yDg1+3L
HdoAr8rdBv5qSIoBhe0U4EaS3FZyga9CPOo3AZfKlUhiN6Ec1d07NxZyc5xN0ZFS1DwHUE7rZy/+
bopNSycKaUwlPiO8KPSOt6ffNTVYDNlXz0ND50jdqGTv2f9SMWAtBn77KIZOO+M+MZOnBtQtPIIt
K0R9GM3NGkivO2lS3Li2PG9rjDQBFHoMiPZbjga/twhQ3cdC4dCPu33is24Ihv3Fa9Sk2deAclaA
Zwekt3nG5/+rklT61ByreQEtTvptds3N50XKqjMtxbtwCdKu7BPgO1VLXDggvnyF1gFZ09WVzpJT
zwc3FEJe6shTxCRhsnTQGkiT++uVZoUBquJCKj9ny7wVyupQdF2+4XAeoIRQtyDaNs1T+XC6CCKN
gVPwg4vnxRJvY7w1IrZ90TD+m6ly9Y1fnHy96xONvqJDdeWyZAq1CxNnkogWaEORH9Y58K0Zm0Dg
VnyHszXHU8o8OwF+SVfCDv+Bwl4YRZakm1vGcmZuTfsY380lce+jV4ENGVubtKnT3eVb7LgTYaPj
l4rgxJ9JLQ9l1RvotT4fAN/ECIq7/wFEWJxmfWCkpkI9TIhvJ/gx9UP1MWv47MgMONZiLYVtoY8N
shnPUsxm0C+ua5uBNdaTClfiYsVIofF/GJBQVtu0q4oGA/em+eQiwHr1ZvpRVh0TYR0bAeITRYeb
39x5bfUDflcpIEL3Map3jwCnY9j6N7ARurJ/wm5msTgt+gHVOtfFdM30Yo9o8Macpa/6H+arCsrE
g9YFR5BeEjEZDMS5PVBnBZ3eWflO5z7iEhm8fFjsHhdW15tZ63mbAcOwY61aweW5rvB2/0czkOLR
N/l0QyIjJ2JDPyxvN8NH/a6VxmhQPDbJoReyYBnv/Pfr8Sa2vSvxDU+7MTo6tEjWufAYWcYbcAfE
Hxw1ycWMbQLKrT1lZUUs2zEVq6PcWlApwik9jSTnhfv359rv0nbWaMiGN6fzT3R06tEiNIlU0iUv
ZOPgC4K+o/ufuPuub3RcByv/k8PP+r3HCW5yT9O5KKJtJcA5HxhTbWh/jIANusb5QEGg1F0YR4z9
zs/4+Gfdq0qp0iR7lLJN1S2xIsc4qWmisqfcgr+RQi2YZ5S/XNgaI5cTXUtzC1xCxp0MQnRiXf1Y
wyLIjXRffmqmudHP6qSTq8cVerpQQMIo9RVJbjeSyRK9/vjWQyzMA+VZpiAXwrTDax66cofJYzvf
0jlc9H8jEj8Ch4It3dwL475Cr6t+1vhvib3YBO4BS9+gNHQylVokdf88L+VyqWolJud49w+7HjcL
TXq1qegKYUSe5+fxxFH5qEOfDV8d4xSo5P/fX6cYgV7Wjdx3KC83N4eo8nk5Zx7W9c4V5M/tY10v
hMbCvhLuNewM028nkghflTt349eiM5UMtO4j5bX9RysewPjTKvf7MfKHqyXSEPqJYeecPgd5FKdB
0q+geRI+9iYEo/ESnQN8AqCwVnXvOjvT5RPCQXRXffn8O1h4K+fOggc36D5Om4OJHzHGUlluOWhJ
7/4SuUsaKTGmn9csb3hkx92k2+Lcwi3aMKN2xW5xfCZpms3M7kfUDeimgmABcJdf1VPfiD30UUlf
XonS3ZYIFABNZ9Bbc3UC0Q4A40cy2vKcQa2/X8nvXGIxw8C2JawQEJWTAK0dHDxIijwbfU/QjEBb
M+XEkpvfH3y9gIbkdr4kk8Fq2CDG7npl2Mvtuvp41mDgmuDc9P6Vvep65eNcAwfYCgKdHdp6Ky0p
72GtSmbr6YIjK0TqOReRyF9xw3P8LXKCAs6iEl89zHxoprKQ8GRMEsuMjKPA6/MwVb3YrIOMboDh
ft56paSLhq7ajVouNRc9AeZ8B7yrA8qeMAbKrkxgDmSSfi4P6+dPfo8AFlGJ6G5OEV6sCAqSgBJ3
4oN03txr/XHHCNRR9IZO+tPfcZrymLiXtcs+hq+0sDDeOw6avnYlUppX4vrU+R7P9RzVuqJVIfcC
ERi76BFrCd5Clx6wQ0gOpD4LstnRN+Z/Ha6ym1sqjdhOvSLJTeRclLKYi6wD3s1/RbVvVjmIKbHi
sXzdR0oHg1L5SDAXl9i8l1plE2dzI8LT2/cx+k8ZTFt5Hm+omQgAmR0QVBBxM5XKnQgaypzY5f0U
VFH6fIHvtTHiK8IPzNzdxJ1vLnusfPS8JzsoZS1XbeSlVE9rMePDZr48/1NOkF9MGy3bw46/4Wn0
2twp/23/UaZlbB2ap710Xza3tH9Kb3ppeBQjeeEpGxLuKhmv5P/z0Y4Cay3r10lt1RH8i81/b5uV
sWNVNQ7qc4CsoHc/V0I+SwGLndEtOqQJX7QPn9WM5fOezIRFj+mp/3qvcSJi1XOTCJY1MFJMnB94
jsuNOQ8dypXl2BE3Iuhrn3DeyT96972xpL4J7JHsqgAzDlkZlfapJFun3jAm8iFSv5aqk0bjkZ50
3e84lLzguMgLVk/Irxa4OFaABxA02udZwFkdT8oakWpmRSis1y4pSIJ+5U8ZAsX27bJMMHaQ2nqM
g+pIAy9VnEVHsZL2Oe+w1a3JGGj6vgN9s09JrG3CeVSr36Z60IV+FmvAUOXzpnIeVEvJhEA7LnyX
UrJOjhqzgwuZJID6vb/rrklhhhWGSQ8PIUgFsLzFLS6VVm9dlPuVDpOZMkJ7Oh1FBuetijD1Vy2w
8mxwdeuijSqvUoxBvvbSFV+6mpfGS9qHvOLdvpM+boDe9Y0rRt7OB/K0DuL0PXdz652prTe2+aRh
JE+iPsErWn+RDj14E8VjQglTz+0tbhl2t2YCQHK7m7q43xJiSE39n/SybqNwW/xQfawi6iEzHA3U
6xQvx1T5FubIS6Zf45qvW4URssiRerULS1L7DM2TtTXThpJyq0aXZ5wBCo2y0Q0VCct3sEOfpZuC
A+/QB/19w2haG3bczP+woHD3rP7Hyo8KM1q1iQcpsXWxcpMhSeKMyWW9M3bFKY3ezBfqoX2oMIZy
2JaRm36Bmlpf3rXj9ctQ59BU61gU9/t2TOIeZKoHCV0w94O6dUP/1yGFKDAobxmSGo8uIAByySlU
cun99IxvQZrS8ffWWMON72+SAO2fDh873p234mso+LTTK/7C5qqVv74PLR95txhbWgG9lnMogxAb
BlODlNBnJQmjgKOcp/GqQQYs5ZYupLoNA3K4cbbsvWYD3qlW0wk2S8RCRd64CaBF/DBqeItyiHZs
C8DOga3aZSe4na+hiNzqRnY/HGNHZzGt6HNkazdY7zlT7QCCpKJrWaVb5Qg/BHbEh4HN2/w5dFIh
axbMPuAnQU1b1XkiN9/r1MGJS/3orkoWkudIWGqz9RYGMfVc6L900d5VQxc9zH8y/E6VfowNNAQh
epB7j4SNVcgQaxmYF2WrWivAOxdcWsTDbQwAFzYvvNuc8TVf+VAASgNfrTlCqrg7H4eHs9Rl0eqG
gEmp2jhZxBAOwUJayUdrNgTQ06nM4FTBJDxWJ9egkB+EoHc5uZcHMlna2ja6+dLZ0rCc+H76PkAH
QNmQRstFQ+Kgt7jsZEewnaRegbkm+V+IqYWEdUKkGX48143d5tRb6SgKyHFckx/6USoNJOQce3wh
hddWRVhrJm6e4Ms78Zke0ljaO6Sf7C7ujs72gxWf7Qu1jMgiSgUb/OWkA2WKV2ZnPb6JsuNMIH+8
FILSC+XcVp68hAH0fJ03IwLofCblDtCfqf5ypmra27nFoCiFFB84StOkP8kHNeYUP67vt+il4N+v
wBgi194Tty134/rmmM9G6Lc+eg40WfSRbyBRlY0yS5C/P0clRDLGVzVkYQA5T6H41mBp+gQ6xqkn
DJcG743qdrXESE/8u3g7APNmA/dvQDXzrInmVI5dOF5RBJeUDVGWrd62Kwxa76n4iVFG65Dytpr7
737T0z/kO3C9aaoo71bYiW0YGDHKAuweo/KLURIIzypj5oYWZTeRfLOKZanhYdeWAZPOi2rw4Uad
AIgwlcON7KwSeVeXP24u0NtkiLJBL+MneRQBxkZipLRLhO8cpDZhy3JzjkeuFBb/1iIzUaYiyy8c
/tmgqNeZTBlT1ZitIpaDmJsQZv2afqFHEVnikectofKZNb6r7+D6K2oBJVLx0uBozas/6LsTK0xH
4gcP9UeM/HzoaHabdqyEeGZUU1hq6J+TP14fmtnL5cyNDCzoJOfk3n2uclkODYs8Wvz3hsqTA/QD
gxpSRr4OGQGsZKTCFnyiK1AAhhswp8fj4RIngjkZprHHZUTn3fXXlwDBXg7xwv9Q+W2by7pAXmp+
ymBbwiww/SiePH0qRag9OwyqeUeQ5U4lgVcMfn4Q9OIwvJwW9NYz3opG8eJH2/qCIpNj7x6ohd/t
6q0rpllLzxopULUV3pJcvSaNfC17SvD6IYOeeUTU2mCs06vvXKqsufXOxE9t7HEv4UumHw/fLaLd
lwsVecJbKuBYoBau1LUXs/mL04GyW12AQ9y2d750sWjBEbAt1hOJMWoHGNB16wfzl8iRsTkFH15q
cyydrO3W8SUQDsPsUhYl6odw7OpydskH5pdmeLHcnTPMn+aHwTXkR2upOSW+Ih4BcV/ZuqnBrOS8
IPMDjOg78aJSdN5Fi+U7rxvYRlflcPhoWLrnWfdn+5liriB3++HVCOd19738UxQ/6L7PgzfZJKgK
a35ajWjvAZbR1/o58lsUlyTwNBCZWat96n0GxZiXaYIP/92RYB+RQE0nRJXIzOuYeTk3UnpbE8tn
CFfKWARP6gZdWEFftSph7LxK7EQ8hHRc2lG9of4DzRg4HDhwuAy6bZhIvirOlP33PEOby6TdSNjn
/rEwIKPhlzoxhWRK7De9xWk4UKjGeK5RIXGGZhyrFkY6MF7WQ1OED7xqcMAFbGNvfr0E7fZZ2syI
EkF6invWeoAQEra4M5kLnzYJOF+Eaw3R1f73WgPyf48DlmEd+IU1LwKLhksHqupwhxFXzuXoydux
oV7JS34Exoqx+XiLsKOfVwSe2EU/VeGp75udKmDWMNXI+mIdkSXmooTcjflzXDfR3kIgIOhEqZbk
PDDJBPjy0H4DymtdVsgcZyPvCUtf4Z+jFEhfmtGMtK1niyRM6FoiwLkW7W1ETk9fpqOuu1ME16yu
cfXvrxpkCTVYdkbkZCUDSoXhaq8MSf/QbS5O19IGQuAAfdVOaTuGzrE8qq9FGiJW+SulTcMJvrZC
PYL2uF0CL7QVu88DJo9ryf002QQlaOO8OK/Nuq2+CRQF97yXPIoREIpdrN9uCYX3BlhH+IdOnNg+
cJC6Oeq+pcWJo2eFGrZzraoRGg2EkZ3A5ZLpNE44HW54Y3157IdmDsaFC6mw6NIcORSYF1N7BSrI
MwYhbB6IIYzrvExQpgb2SdBT3EBOC+rgt/AahcOyrVEorHGYR12UTy11j1thzwkQnZa7G2IHuCGI
7DLb5G2ISjcNJTg6/TfJOfCx3DYagMp4UXeNAKGOqwTM13aEg4e4eIS1NznLswWPLFSAwvc+Up8+
Yf21A5Nr+5ZnWiYVS1O0Ymeeo+0zO3CUdPRtv/qtdnMjmT2YvO0ca+FuwyyzgmIh5G7kXVYr/ayF
azXomED5Xri2maQSWMJOFpeEZAt76jktbUEtGLkHz8d/OBqgiIc5MfJi1am0MOj5A1LkuX4HIy32
Vk5Vls+Ynk5YyhFvetClspNh3DBijBQyYlcytDr5svR1PoihBsZbVIu8WUhV2rJHNWi6ER6f2LJ+
gH/pXb8lWnstDLJ/sfnDOLQc46+fDUeOsm5ssH56F+lvu4wcx7+3J13egQW+C4cT+/zdgnw2UIM5
RaSxHw36OKk8eVuCweIxDxwCpcRaloE7c71WLn5PzfPyQ00aEiu5dZaRln0/atHB1ae5MGeTTLWC
u6YMsyKIRxabcGatjEbDd250ke0d1phMvIh40OnJnqR7Py/suP0VGbcqRHP76o9LDy/zp75FzhlC
boy2sA60BZQDXzZrXT1GeP1bNvBtj8fl/KvXs95v4NqPID8lUIxksjWX9K9MyeTasJOi564vmz7R
IK22ExVybOQJkOCJ/KySE8JLVKeyxowOSMTFAxNRTSuLzCjusvFVbLh2yo0jVsuevILQzZlmO2Eu
9HXClrDE9I8oHsVu61y9/VZhbx6ixo8Q9vA9B/kK304HJpAWk/jdmP8RPZWxxg/VsI0xKK+sypgR
mi3GFxdWuRUhpSu4WSLtTrm0iMixI1vmOlgUPaXMmVT+B+G3cAwMS7xqdzQZYA5+CtOhvLm0rEMO
bkx4LmKa+MKWprBcNk7KPZD2bNFs0pedH0N9WnBvuuTYtR2KYhpUYaFgNx4CCudfpTZcCK6rEeX+
GTG81IomBBbtVz9N31PdcNv/4+8dLUqPjutLhjPrhRN9WZJ3wkN5tRNCRbhhwr+8m0h+N4vKXQ6C
xrK+qvbYq8TLh3IpLw+iCScl4uUcxM/Dt3NYhnZTYMz+PNotNHnzMRe0mm0p/BIvGJbO62FTJ9hO
6Ze+/sDWzjaUBBIckOjzWgM5RWKG02Y4wuurPn+teTmfNJMlnNJqspln0WQxYMBUhui43QOmeUSn
qiGzcpeguMrRzaaA3s0u7cNYsVRLgO6mwFcE8RiDTk8hWoP3b88ve5NTJe+zlonPcYW0b1CLMMCT
RfAv3jDulSgUG7eX4ky/plgzd7rAj1jlz9MmdMUXvw5Hl6v6Bxaa7ypQXWGvJ2AQEHRZcDNW7FVb
hZKrF8K+Bln+H/nP7JtWK7dOwbG3FogVOtY85wgBh+14ke7lsqda4Ewp8i6bynSrK/PmC5j7cHRz
QfGleLLVej4LkLK7T1tsyf7FEEuTAo2kkh6uG/X2VaNBuQ2WDMJdhDAeHcICoGXklBUJ3OPkDIzE
tB6oMMVVXUyQRoUXbYhw5re6Igvs/p+mIvbEcTfJBTAhVrJgAExL4BxF0Y/1TELF36q4r99fHjdf
xpG0rgcytJS1HkRGUBKnh2M9+8miVlgtN+ST6uDsduxrpaipNcq4DXltufs6xpj0QCnwUzp2S2wl
DhC0EFgjehh7fdnUXQdKeFD9gPPagqBGX+eErx4MaPAcuMJmR61swYz3h+Ezv2XmmwAQBnwyWz01
zgGM7YSaIELo4P0EL7cHtYEWz1BiL8HUovlyebWWQq6udmkfUBx2xslagpD7PgH/kuyXzcPnAAj/
11vLVA6WJhF46eT5kmJX6Df3YdF0fTv24kZDGWHn85VnEKCyvX69cRcCoSuZY6o3HbBZATgcE+Wn
DsATRrH+k+nTihMiYT1CZPWvT5KZ5HUMlwCe2vWNg15hIUxVUYYfDnIgwfCh/URqlC7j30Sm5YfV
dMyxOfoTxRnoCsRwF78Y4vuRzqRHTuqKmD/ldz7w0C3M9BxULITnuu2oxd9zmR0bF9+7nQXMuPPF
NWJ/YvAW7MKPrEJ8wlsr9buOytm2QtkMCGiCW30Qi6R+wf2nkk4OhQxrknLQsXpqoeBQNm5HniVf
mGEOv9IwasedqPo91q2X1++W+krNuSHOC8wYr/cVgpiYcrbE96XuKcEEpIhynpm2qoX3hL5+g3NE
8SsPshy8jbHeww8BZHl8sF7l9btpTH8Jlx6lsQttMX3zk2CJbp0iefzrkWx34JWAtvF+Z++EtjkP
gsqXKmL0gK/hU3naUUCHxMvgj2viJMSBFRGQVEUqsM1lmJLtkWPwrZK8E/07KngyTgYGAWCX3Ak8
3lckEThpL0SCCcsPyiq2Us2prT2XHbzrtD6Tx1o/XppOm+4y7VW9S1ViQjDDEOzsjwjZBIq4ycj8
nSQpvVYJM80ozLjHWMN8U73D1UfoBrHI3URPIXC0KBDBtRYf7r7cEKrj7PIsja7kjIcFmn3+8XJJ
wDPKVvKMSlJ1t+nJbxgWQZqWEHG7IMkYSxZF6Ww6NO+SB6VUj/JsGqvaCYEFtFw0HEAFqjexA4VZ
ffP+cnbi1O6AmJUaar11xQvd3UU1VtL0GvQ2Q3yg0CZf31kQzS1NhhJKQ4G2pVIXRP+z+dYCgC/h
leejxjR8Tde9KRoKp4awBfAGSc20cX3pgvE+EUE5rRrWvCKQr1ZJ4JlVNTseIdpmRkYjBEGltfEq
D/gLDEvAmjDc/oQ2+Z8xUM0T9a03V2zu7vBbz1N64wilZeZGsx999KU+Hu+z26BnhkFTv5Osy52W
CwRRIEOgwd1yf3hUNaeWd817dsg2MIzsgky+l5lH04LGdRc1R+ZDyj8ZcCDEpyImkKp24wsdw2w5
CKrpZ3vRKKvaPfs16+nNg94aABObokIAxaXbupl7ZQUOgpPoTmPm64LgMkDlwOLLiYVsD8/oFlwG
+5mAjneUoWOS2q7c8VwT/wWmegsyjetfDjwSlNX5ZxTQoNmdpNOgY0rfiBh0gX+Md5+kgYjcw8uy
UbOjZ24agxvXv+1u4Un4AM8JbmXTlRdQhd0cq/54aL+XKSrDsFvBz1bzki/c2tCOP2nRSFxac1b5
J5e+RWVbrTKH87ClngVJYG74Bcyv4lPxOZEm03KOf6G4w6mZvYT+2zm0lS7Cvdyby7aQLcOKfz/+
o98KxvPf5SbZJYKYyGyiJMxRVYH835SuoO4KyO2XEkPSAm8U+KLkohJYuBKWCPxQrGvDI1bqKauI
xSO3X9tbcppvybeGPa56Y5EVF/0VV/zWjL+uDR/OQmoy2wEW3wR+/8K1C0mvjYNTCzYBBSUljsJh
GTD74Nf/AXg1NrbU+dg5CTU+cmMnfpu3JHo7e3QZOk5USUH7nOV7C1LUbwkM1mn55LHeu9U7qEL+
Ujrc89xDm2dJzIfFWJ0ApJ1PhdUxEi3rzJG8B6qTTKPjUPfiRl+dfl1jtI3lBiu7B/FdLPmmW1Cs
64IfXYBht6BLGiftvHkElAkY70bx63NCqp8wrMM0It4CPT+dpJWuv6tHpkn63dSIxIhhMNkyxJ+k
iUU2CopWzOfFMZXpmW6Pbg6mKkfTBTwqOkLspDrWG9GfYWOXpJjaZaT/z9qlZAwg6lu8i2sJTGQl
YUuX08sBd3WhBqdS8nFA7F5gFhEAMsMU2s1OFzWhdOFAcR6Q63tRS4J2b8fLQS82v6MG9WGwWtFU
V4XASZk9JaHD62Odbwv7iDx5QtJ6kU1DVJy/uhcVOuAt02LdMwxmqHw6tbBBxuJesLURa+9BWro0
smz26XkOb9ppLWYB8uoSHoFFWoezr8w79/v0T5oqXS3cM+eukimTncFQfZC030KovOQL3u8jRlR+
14VUBLMuhG9bOFNIFTqrUk0PyzONHxBLdislCohEiPTISdLeQTBfZ2/i6J1AB5Qoz5PE9Nl4l0vI
CclkRmoVD6jWTPtTE+j6uj0g5LukEv88G9Y1YPrayz4NkdsL8es5kxx0QX/HfxOC9HggNm0YQDx6
S6J4KX85qdw1bzK2QEruf0J3pacAyz0cTd1YuugJebEvIU53+X0sFG/XgZBiQ0JZgNLZ8h9U1RYh
5wAZIuFXm5rB8qHb7dyWuf27f7jhQCsNHAfFYxwKfH6KrJ9Ao+73VHwN7vOPkFdO03a1bnidD+Xg
Y2H7uY4GPnqaThSyH0+x0QMi+tbHkq9dAvywWtx73tz4NaSnQo93zAKbqS72JmHBpo+SNlVvWMD4
nECrfjzCXHUE3878G7vAlb+jnRS0Lwg8TxePnUxAJSb8a584tqmQIcQG0whnB47netopEXTGH7z6
KO6qyULgH+vwIVv+1TkVMaz3RCo1T0WdcVo8Z/ZldTUIKCxS76RFW6MWE6QgtwSum+9DyjrN0as8
T7o7+JC6UkE9La69ERjyv60UXtVbWGZPhzTIEX2sYPJbePBN9PNSpdJ+XgKBHZP8s9RRvYQGlLmU
sV0Y05Kl2AY2QNFYMifgaxoVdhpxQyIYJa3ABT3rFzoxB8Vq0fzLnB46nz9xD4VVVua66x6GWy49
ZVBsjP11DgOPrW8F9Q6+Emq+Ov1hT4hSJEGlvpj8ZoCcnFWjlvcypGCyQ0L+jiOWj8L+SPjy1xA5
vzXnCWMaDipMscpS2NmARQIVizICkYxEdeuvG1nX+y3zu/vsc1GeBQSZ1+jAFwxl7IyI7aHxlIjZ
RkTvOPS8hRsE/T6oMOCXyCBDMQz8RodDM2TltaeGMGTl3Nws8sKwJEgWkDnna36w/L7suvhfFZQ4
G/nsOnFWsKMm/OztzexI9S0GpudVak7Qeyn2FCNcaRDVpwkiuRQ9MuL4Gvc7AGrS4v2Eg4IALSt/
il3iD+4KiuYTiwTHCVDpnGq0wQ5++ecXSRINrPEGkT86Sw03poeF+5d2qgQI1MxdqRtthT0TozII
HCVvsAYCqGJAnPe5KQr/3Ir3TMTm9gpVTPkJeNIZnKTVwLBfo0bhGeV86sf9A2D0MqyrSPeezuUq
pTaXEE8JE8Irdz6Q7XO8KRf6t6g/v0Ur77iwpZHsjSJYK4RkQP8JYVyuOza6v8tiK4sT0z8ZgP81
QTPtQkCGhe1YlVDTdSnzWfJWqF1LTVO67vhwMIhQQLxAeMN41huInnIaozlIYjUAPtuEeibrzAh6
8GAHVRsQ4L2NsLxvEEu7PDvsFjTcukvZbgPXv+7hAD+2UwmRKDuivxTV710QFYkKUOmOfsjjTMUu
F9oBheAfljDVdllnMU8YRU5k8THzZUfq124NIGGqXeIRVloBcfbu6LNGvXYymddnGwUU4Fk3c8QH
IGhU8h/FsjPB2HYR1pyh7XyMv6ZBu/xYK0gEawQMNev6sVwvgWLmEcmhr3IaRKLapSIIhuZr6cH5
v81CtxcYeLgms5UHB3tELmEnPmVERJ6BUJ8JLnDkPzAke+io2qKspWZGEFUNh7BNUY7+LzxJVXmQ
2i79U1S3Ce2L7+4B+F7jGhHziKk70ZX0A4Ds6BC2/7Zjm3kFDzxZefVQ9TZtOy8UBHH2GfGDWWoU
N2z89J+DO+8+4lCe+MhFN+6b4qJDYCUn8DQQfMnENHkkIyeG4AhnzSvflanWAHl0uCBnJK3RoTbD
OwsH/Eq9c0TN9oB3gVABF1OxJyVlmLgNUV6rucxpOOxp5w5b3GNfJt1x7ACHtMzsjDV8UnMJ+Qxb
6rN+x+N6U0TNKvW13p4VQj2fsbpfSThfeXxQEIB0EiHK+9yH1epjI+QFmwfjVSiOnrtO5eUQYM8U
q6oIFPKWEAdqIMTFNMVtkA98gD2qxnZWvRB0hXO/0taz1pZ4eU9soICk2hkOW2CpnBrNtrp//jK/
KwKt06cE76EPiL1XmSjIYpPvbje0onXxmJj6E6A0t3hePYH1ZxWFhfPStaDz+xKpvK6rCu+c/jgy
GR4b8NQ+rTJ9seHICXT+Z6DJy0tpSJmrybR4tkYQw9HFrI60o8bENBdmM0iNY0oh9BBiy6sQIf7T
Ttgg5VjnzNpqLeuj5BAyLdJzaelCEQMpuYd5Ix0STxKFsFJIRU1fVNN2VJ/rG/XjlhkazZqdEfvP
ysdnwVKb0defLklmilM+RczztdASx4++Vuco7Fhzqrm28wH02m0PWvehkm+j/1E1qILNvs0PidwF
1B6TodtS/+KLXXE6EdfYAaSe5svzUgr10CwCz9B5LWbmrawbnWmcBAVPaReFznTN7K57YB4xAB1P
GMByoDPgNy4xgVGqMSWPECl30AZbDNCsBk8V1b8NthnyQU/j7wT4ucGE0cicK4C7jZk9iQvDcd6o
UC/kjAmDI0V/Md5AqdH9m0PivEqGUdL8TdbIQddZSbIcmpUnh4oqM2NKi+/4oSiapaKR00DFLua8
hEQgoqU2eIQu0J/tvJrk0fI0VEqQVPbx2xgi8BiyL2QhKinv/gR0YW8ypI2OEP9KXX11KaChHf9E
9YlIfWHSUFxh8Wf/PMrsZzL7/MP4/o4+q/Fg/Yyo+PfKdo28jX4OLCsZ8VRa9KaxHxwMyf/lTQbA
BfO1/PtWUD77WcMDFH77N2Y6HhbeL65yENUJFh516WXUpzaOnFCBWItxf+3X1rMLYSoiV85Yz7tT
Oq5bP9RgB846nqDAg2Uugs0yDJgp2LXWhNhJ0ohB+zdyh5fC9Naoh7e7NkvjbZuS8Du9fLXJPm3G
AwbtB1JB7nFr9TwaDQqXDDAwKbI63jITR14xtGdN2h//fi6jCgR1vrJ/8rMVz+GkL22Thtt/eLo5
3mk/xbFvIxMqB9J9YZfc5wdfH+pmbbwLYGOD0AjT1t9F8JUaoqtgp8QxWuhA5+yWRRvMASd9Sm/h
k1W8p+gq1A/VQv5Q8Ky7Pwtg2pyXnk62GQJD2GTryeR8w0Ne2Q1xom1T0kKaNc3ks9sFKyCTbLL8
WP/tjAhBLNihCNtNvoN0a4XF5Hs/87ss4fGyb02CXpOnAM6c/BvDOrw91MQG7U1bK9XyX50SE02Q
RPoB0A4fvTeDvNtwFjklzqpRDCMHsbMHqy6iYvIO8nKk3VQ7zDq2UHeBpwycUz5cqM8hp6TaDjuj
ymVncDpo032raEQ+Pe0/1Qko7Cpbq3BS6YeeTLJKjsH8C8Z+nNfUWJuGaphjxHKWaZuiaqC3X13t
NA/8cxE5auFqzxyBVbo/oJlTGEhfWMXre84i/70ornBtVbhCsevWN/+7p033SEekXC/BlSddYSWm
QfGAiKru0YA9iDiJbwGhlAJVWlwA/Ail3iltt/cnEwAfm+cm2bcZe/bjRNMB21tdbTShpXbNh0k/
xHVqSiora61yQXNoVOWI1cxR+rA53hP7MPP3YPPyDNP9CGbTHY7zhQirSicj9bTuHYtzArvMCkQi
qnS2Y/YhGHs7UFwPr5sF2POINxyaZarv3bnCP0KFRPyrS50ybdeOXFyeqJBAte5cI8JwpbgElAXO
J+Y/jT4d47XhMTG8fRLITsoVnsgpVgf0hLuhrMLcE1eK2+ZYM4ZtKJaZiT15oHAmNda0odL9pXwG
tem0c2z4mZ3StdSruj0zraKOZ4B7i/PMTrqaFVe27aqNf+dMUXNF7tPWn09VUH88Ykdj1VxFtvk0
p7Q1zfs39I7pLFkb7aOoY2B+dKgbGJS4+bpA6hQCTWOh5qa9SyEoLXwSJb6Eu4uwxXxQwxqOyz1b
mkX1+r2x0BRhRo30pyL47IZK0gxBErZ9aGkO506tZ4p6I4cvkcyVntlinuvwqQSjlcaQxJAaSm9x
PF3szBCG07z3jUzekMBmh+ycYZzMV0zolVr+Et0ExkYn3sV7KBBjkaxiqtJd/hp2sWO3sqqC6t9y
n9N+OlWPaxMWtoANKSn54v2uqV+8+AgplseF2AF8wuRqfewCLYrmw9h22nYylLnJFwKfaRYQmzUw
yJO4jvDoHvh55TYMgBbJNVOEcIgGJ2dp2ZaUMhDhDL/LVstw2N+lmZAe5+XOCwy6Qkqx+tK8Q1Y+
PL9XbnYvXjFYnIKss5gVKGk8WEpeiMCbWPBmIsBxRlRlXivSVlLjqlP8iLVWFSJDfwAEJ3ZEK3Ug
pK7imfLRfDkhBQry8vDGQO1tPlNbEgUjj4m63x9yNewbDcOOwlPKmf10IIwgom8lCNWNWlPM7CaA
lRI335YLUVyt+d/EHYVJ244nyMbQeDJld6TBIJZ7oUCHTBM7r0jvFqtNIb6VST7+omMZHkVrarba
1y2thTnJM1GqXAu8u+F4C+TkZbaNxvz6IRTaWSWTv+MGepSAK4JqbPLj4Pv87I+QzBp9+4cFjNoN
nR6x1QgZSDLiCcT6+ItdxehaZG+zeud1owaP/+gnO9k1MtQGMOXfipg5ZSNH7DAGSr46shBoLBUS
p2rm12VAqCXSPWp/sB27Bofy506ie9jckkJK0COrcOyuapiXTEJIwpNV6tGNnHzkbqxZz5hgvJTk
qZgV0cZ71Gj8Gfs+eYK0zji+KUdsiSyuJWMnil5pe5fIKrttlk4o44kYeIZRqcNpXzKwqKc638ar
w+3S585DfLdxS2RFjezpusIJp4tFz+gotqba/KxqXHKoTP77aWq8yO54tVhck7o+1TsoeWFKepn0
fJzqxmFFx91kQvb7N/IcgcjwjtBzG5rDng6/G7BO4a7CBzk5u4n6YFSZfB+7QqffBNuO8cgDedc3
l+PwCwTW2bXFQLDO15EETrVvKYSY61hzB1flLGqKpFt7pCqEl48JM/AsgskISCNt4v6/gITwzhe/
p5uDRBWe6eChkSSI0XtKGiJXiWh5tTty4rHjW0T9mmZBIuV1/h9l52lv06zPtI9b8HfVnXSHs/os
qYJPwg6u73ZMIxz+b2pOmogBM+of87RsbdLBmh8XYjoc4/tVHNQVIvgKb3QDlENhdtRNzhlex9y7
rSM9LVwu79vUNuEuTtm6XEYFB+6pYDyyXAhZ7if9zzTqSYiTWTxr+kQeoG4lhCbfjwWyk+NXyslh
Jc/QU3f8bYwdzooW9ldApZgHXSpTTboAC0VYWUYuINXMjIIwmYasbNRiHcGKlt4QZlYCYApABEDE
YQZPXxUIZV7xFJpKRApHj1cgvQSAmRnrL8StfbkoEnCkmG7f674qD/8bbFwKwgiRCihlbz/fAK+B
DGzntjhncHSyq0LcWXbWkJpL+uBFMo3vTzlZsbEU+6faHCK3FvWwflsyeRtIL5JQKez+GYb7MsBH
80o863PsWlq3oAs8zrD4n6I7yBe3mqzW4P+oYlG5mqBfp9679/C144a6ZqRzeBjwZEYfY+tNeoJ6
+Kk9LN5uAehxt7X5BYCPfScaXVT9/5Ng0x6EQnUj4LWeZ6tBqJ0rhoBbmeFOZVAUB5Y/ERzP3mkA
w74UN4axFfAv89sLa09vb+FxrO9ydm0+orxl633ooJQ1bI5C6zTNNm7m9eWmYcbFLIyQ6IEQO2rI
BzM5qC+NBeG5r4wSbe5sceq7wPb6P4GofB5F1XT3LLlJRnGjdWjmn/x/TTigXi382tbai+pgHS95
vffBwizJWWBiIefayuhTrxJny2HuMva9gx8ArvaCdxpyJNhft1b5eixaX9jjFeuJTzjheq/FPyIb
1iTB/bQwFsrN/7zVJFjlBFUc7OUFLq9jqeewhmIbvABJZAG8b7I2P63LiJnAUyA47S9I++HCR2kR
q4Wga0+JTxrE+/iqwOHrHpB0Jtu8zbmwf6j0oe6xd2Gkp8nSsG4qNWHlFwcq0n65gj3tZwDk+jtN
PI/XOGnJgiHss6QdAVpvPC12a46ZsNIROeCodxP7u1XOpY+2JE1WS+pqFUnvM6j4kIMVbRGRMNaV
aSnyo5ewlC6Dr9JK+aIF8aNtsm88muVFxX3QeeXd9SWUP76qzFg+mr7Ht7dBydnfHxNDVqm5kmcy
ugzk1ZvkjpseU18msGOkT4TyXRv264KMmv0yhKsmEjt7nNYYgekvJac9DJjPyNjYYNG00OoLpR5e
UdDbE0IOqN73MJwe+b+FFnYB+VLDT++WpntbKXhbYFPUAo5BV3/VwFYgKHGYCFR/b0s3QoHlzbpR
XgDu+d60iytL1utDZn7CGuzFgodRng3R7hFsvdBq44xjB4WeUcbYGucxFDeDb9CPSCCMd2EtZMcv
uaOFYyiiCUMUknjKS/woEa4R9LebH/Ypwkk2GTkK40f9VJ0b/iIqCG/b4nQaTHcNWSeSlSj4YbsE
4vu2DsJ9RqhHCnHQJc/JCAQvkCPRk8QmzFUDEXuEESd9Uj1b0m2MwA7pF22k2aGy1UWZ9jthnMR6
W/P30E7rND09dFJ0xiXxFj6eEELMV9OhsHtijueZ9bxogm/GOCUnpkoIdIFVY/ZhA6MX6e+Ynq/j
94oawuOHvA/KICmUlehHcvMIt0hTPrs4OfbIgYrAj0lXweW513EeqDcTaM12aRxzDye37BsEjJL7
Q0fxiuOx/SDd/DHeSbim+6hM3QMUSUOoyMO/vfUbRE9B7HQKfbEkgWxpbwwDdMX266lRaTDGS7qr
BsGPxezYzadxGM7Grh0Y0dswLAXWIMiwnsP9c40jgdYGgzUmsmvL2DYFeX2/XGCooVA5s6SHvkP5
Gl6a7lxdIElUxfczRMi2OuHIkFmlbUvr5g+I0APGlL1sKssnn1ZDh4HEP1VX7qc++w/zDxLx4yhM
z0pxfwidlNAxlZVtTadcz4MgfVVl0t/5nPeZ/cjiEWA5ge/HNZBpRdMgUTFxlpHkV4yOmdWng7Sl
wozIz6kr5WEo5AaO/daqd358EpcPbEx779oCEsE/MQEOkkB8O+uZLlNcxJ/YnU/ElvBRIy+fGMUM
VBxUvaXL8hDjHuLe8H+EA/GC9HpReqnSdQpPR57zclhtJG92NKtduAcebEWQLIHxPWf62GEYJSn3
FC6B+aREv/QW+AeZ9OjAxF1cRiODSriLd4B+x+4qTJgy/gTe5smRaPRQ+iOOL2Osk1jak9gjfTwC
vXXGfB6qYzs/f7TdTquYeIL1I70y5UQTuf7dCPf+CNnuKyFmfZqoxoZP1zRPH18FacAVyReTkjkL
xhJCkxE9GUWUjS4zpXeEqK7lEiqF0EGsAYeeRErKvUneqX4Ev+6Ns2rjj9wmhuzAx0vUXjbetjye
jDXI3CwFy3SZj3atLJVrcnl8mHOXUeVJsKCiWS6spsLgWW5a2InnVdXDjJpDu1fyoMuFxolGL+4t
R2AM/BDwRMh33qdccYM21bbyLayRd+U7MQ03D4qLGnzK0ImLHCvXfAGQWkPepOT4dHTYcNJgBLpk
5ptGa9wnJhU8kXiIAiRJq1y6WA8S0cR3dBHtzFA7ps3oDCngpX+cq/ePy4lZ57Vs6/T6ddUl5ojA
oKlGqudIsWAGqzblZEcAZHgriUbT9TP4RKbzASieQKaAODriS8FGmaxxLLxbZQwMEDSxTkQS2jrz
xlOh54lQQEsSjiQaFfSTaQjSDW2Jj/C/l8SJdUqbttHCO6r9PU/QDK7atq0MR+g7XhhJGYRZnW3C
bkHFM7YZ2bRLCk4gduQwpdrQVJSe7o4P91EJ8nYKY7RHiQ/u4KPIXRdi3L+oov1MOuKlonE6v58S
Xud82pmzcFqZCZ/YaZJZjczYViF4Eh+nPNU2ycmgryJeGgXAqbNCWuZDLfKDGeGuhIsEje6sb2Rw
6nbu0Veu98I0bktXOIgvfEeThJt7P2PfhsP9hm7hdaLYyCqM2sqL5PBgJAUGiBhPRRwrGbCvhgC1
hGZ9mWEQ4QFQt6QpSL9WhWeYeH8DZhvbYVJuqv1VOXr+fyTsc0ZXoBOOm2tpSIDAD+fc5eUaY4AT
ZMlk6vsOKeTfQ/3aN2MYC3G6HdxFxc1s5PVuR5xMnlmxB0vJ/dyY2RasAgpTJyoor2mTnyAlEoA6
uRDOitS13yIbSC38OGZbK4gWdvlizSg7l4AKKfGPOKf0e2rbjmRPYgVBs1y2i0j5Qvh4w6fL8bj3
VM9/3Rj7D56rAcUPqti6SQI57D4CPLrN2wDYtSDjjQwMpmQgr+HrZ+wMKji3eg6QMAsftxVW/8vE
IAcwc5zv+AEs3y9/B3zlyWSh1XlsqwyMdhWTyuBMR3Khesd5ImGHYIOhYiIa4emt4Vs8+fjiZThm
vFqdSVhY7TNhdnXaohrzBHhJm6+k4dYiGy7HKMEWVDMAFao9f2E2wqySN5kMQXgkbBjiGoUCEXhs
/+WvX5trVdtutIwg4qN/cE+1YneAyL4ECwrB60AQg7YqDTeDEHxrZLzR0nthQpa+vCh3+S31r9i0
d41T/i/QPEUAx8ZHydqKliLv50BiCRnC+jUJWo13Iv2rqALfOnUDSILpJ9G/WVvkCQ7blcN5bEGW
jjOKDnRmf+Vb0bb4b0NrWBvdTcO1978ZQH95WaU1H7YQQ3rmOknijlq4EEBLbZEr6zxE0MfkXNSI
bs2ZkLXuQ1qaFY7UPCJ5BJKpa4LaPfJaYvzWUAXYosrbUVb/ner955bN3DQD9SrtXmECGZOMwbEb
Azcg4KshgeoySriSSzvOQ8cfwVuM0Xoerri0o5PKGqUlk9ysBCdsBLg04X66nFZlQkePpAAFSoUz
73cKr9rHHB/rVq5qFa0F8Ttpg0lS4kB3CSfnohr/QPLWq6nb5x+ECWynNVbahef3r8g/bCAQIEFi
71ryrcTKwadwHfYnLDTzhm0gwhy7oeQyD+1f52dpEjwqNeinyGW4HXuAGBsWydbrHsLiRO2xEEgg
cf1C4UMjVt7G4ylc6beOjvbHdnfApEYh0cXNVBL5VOkLVcLzRTxzqPHYqAfQzE6nqeLrX5gN54mV
BRYUyV17v2qLRJHBFvuuTx+TYzCYdn81UVvsrN17YgAivxerD0ep5J1yPVLsGRcl57x9RJdWAgHY
sAzCrCB0DXOOE0yoBf0BJssKYkw9hYUVZw0TtLUNK7pmKH6mumSsLOsWTpbzNcrt8Y6HL0SkFO6d
y6KN5wG7yC4tAw4hBFu2Kx6TaRGMuVtj2aTK93ypqwPw8/cIfuVmU2UFIX7G8AgUajH79TvLXxHm
o4p4lnpvKJu6lIskgwkneVUSmAAClJg0I74X9BsixNdz0m6/6Fy2uLaBQOpzOjG1MdUq1+r3YJ5m
kvPkMUvVNr882HejtXzey0Ngt/KDHifINmEZUbi08FyncT7neDh6TdCCSVUxQdfDTvLdpWq3N4Tq
z9UqZhrmBISkYvnrmS9esnzJkcuqkpnMQoOIa1YXDr9TjNrQ3bkCozvc3RiloWe/VePl60qwtzT4
uPnw1NKpAcZp+3ZlkN57Ec//5Kb/P0Ph2qL2i9J6rKn76VCGpdH6+uuNq4d9OBKcH8FHl+vrqOAy
1Z0OlgQ2NVmdbT33iBB8pwkCMxfOy/wWiteNg51P7BHCnOo/UVO947ncdKZNkmjx086BpL2Fm9UB
weA8KQlV1UKQQcbMXWKbxLU63oCxNUTzq0u+hQUCz98qly5S4a1XGZ0ty6pGjclpdLlDW4CftbSb
zQJ/9mm6I9SIqK26CmuX42KxaZwYqnh0lK8kIp0Tbr9SgN6OthQDSUzj5D4y3UXUBxKL9YNvDVvu
Np164WybmJwJjzR6WmaLAAL/LR7sD4aOjiqP0PRapRqknrtvtgsYhQbuHQe47Is7qf7OhPyoLRRN
4drAroldw82Wb1OBEJtIP+qF90MCVD2o21qV4gSYMpzRbPku0p2xAFYI7sI0eu97Kdey6owunK0U
nmzj8HS8fI41izW/sYpDRYnNz0snVkW5pLnV6s7b8NMIk0LH4lXY4CdF4Rk0NWXBEs8+3BY0rKZh
XZawwF6uMb96IWBwWZGJgvApbYFJG2LyJEXveQ6ptCPbf82SBta+21IK1YUcWdtYWwJEvsgt/UqD
wykoyhzRNuiJY28y+ccMVNKVLtshMx1aQPPsYaSToQWSITZVO6XFSaJArDbV/VnFnumXFpLjQCGy
rBz6Zk9wpz++k+QuDtA/MNqQEzYzfMi4JBiLBAg4Zh2M73nm9pQFIcqVHXZGyDBlJ0jtIKF4SyEC
dz2ArgE7VvH6XGo1RYtOalrnjm+9Uoaok1d9rPuH37QXHsH3zwoYVClrmo1SYRIttZyTZCXJiQKh
7+FN9VvaPr5lfYF8EHtcW65UsKsO3o1Yx9fJvS7a5pKww+uhSuIiyGlw24jTvKlfjKRrfPnh5bxq
9s8W31xRMfE+jEdmem+iEPd2U7Xmie3iEsRVsP+56AwNTojNoMf3I8LFEt1pKAlaBI5ZJQtr1I29
mnHbDgKaJR3nC8jTfXOrgV6q1yT0PyiL9MHVzRGcWaXqQPFhBy63MTuw7Jf2OrYkIVmO5jJPWcag
+a4MX0AFfnwnGXvh1T3LIsA0xI6PtXxzIuqWYtXw7bnHrTiTb31Kw0HyAVNWulrXSs5ZfZx4m13T
s2YH9dVWoj+RIYvFafXtuhbav6gVDtl3cKFTLQvXzOanxAYAxxugsMhuprhQy7HYlOmwBmDojffv
PA6nfsi84L9OtUfSK3X/RI+FKx5ahYY0HwUbs4TK6bKQhls0YZFzna3zVG0qNhQT2EcHJn1n26g7
dSFu1/3kBaI9yq34Oed1yOLzu7wkDEgf4bYiFzlXj5Y5EzCoL5AzqYdwtH1Eb7zxt7m5RzzUSisL
Yq9KpZUkXOPTbKtaS+27i0jxmK2FER0ZVs8jIz5/t/6SaKC3DoDww71XtHCOBGVXJBEix+F6dEsK
wW6YQPwJsiMJ/R+3+RQ1/Fv4HCeTe42DyQQN/RvuPaA803ZmOQPOLlBXIOEiuZt6FYwQBWs0iQl2
yShHwYs2/q/aTQSzHV256hnEKctk9sIgQ7ZmMpa+Q5HRaE8TSPJ9f+CUPfPOYS9n3rn+yEfEG+Ll
YHQ+3212QJE2m4sX0xsz0T5thUGtuvdI9nT47mUfhPhvFW/EFp6qMsyzL4tMGylbZFvcCgfiSF6w
lqVebObZ2C+bMSmJGiOn8pE50UkRIv192Ur4/vo8gZo35um5wZ6iI1eYPkyH48fBe1dCvG4HhxVy
4i3gRtH6mZApwIcItkzdm7egzm6vpfZNunA4dpPWQnp/dRBIzmkNI/dykgUQHNe/FIFdsb9804nt
z4MLj/uR9DsqrcQN3u9JGHI4VAJxCqI4xTWEkwLZzcdofh8AhmJ8UGPGoOXc/jq1j1G98kkFbzMn
Lf3u9DqIJ87qBI0r0lo/zrk49frZCDjBakN4PbvrXInMsy36pt8/5a/nqoGIAxXaJoBWuxFJCcjV
iZP97gYj1n0Mf+ZLHB+6IVNp4IyLxL4XdyDeZ1tPGm3vPLcsglC2Tq9cldiIRvxK6PaThk2+yrZs
aOjck2oAVZEssyKWMj3Zrc+4kDIiw67t14NBw8eOZ3+75vBXGNCnzLyB8BN4TcDWk0enTk2HbMxo
nr2kgUVN7uTyI0Od9z9KrdsYSQtNbfkVWsEhZkH0YmeZ9zXn+IhwY7gl2WzdoOE68ngm70q9KR5v
rGR2GeglbYZcIp+41+JRxRoceS/cykJkxvfrCzEskqMNZsNUlAKm0LB37+gMpjSbP9zgAsV+1Rgs
IxOl2UxDfIhh+zL8w0AHpgUvtUljoRx1Iea5bGI1gjKT8jR/KMdIwXUC2MoorGqjbn9sS3rq2BBN
E4gKwGj9NTZpzu5B0dJJms46Q63cXItf4ny969Hgp66mAhnrBmHwlms0D3ls5F/KwCFZnwUCrc5V
T52KPGp2kNbJn6Kg3BJ/r21QN7DZY03nyEJUfeJ3KNS1OoSSvl6FNiOdlYvN1fGyW3AZq9NqKz/S
bvgKa061LbTFycgS3VgUp1c69GpNM9TM0YX9NcvkrcERpA5uwXYKV6a8+YePDT+HREcCmDp3WflX
BS2FYd5Dj303KerMpWcEBBBaHlLO0+uh/n8bSVfE4fCDs7vu60pv3xtGtWd9HBepiWHtzNnc4Pyl
eHDejqzhf8RALOVVUhZ46CS23dqe4eEeXgm5grwuG4dKrPKZRCHlpeVae1yR6YMIvxsjFyUTur57
SrKr3xyf4w1A+5EwV652OZHRByC5X0VHK3zyeS3TDQ2UsqEUeP82YmaawMgGiw/4WKpt5dWqFGzC
imM77sG1iOqneETHT/rqOICCExTJnXZ3KcJJtMhcx7FP7DNM4rHtgZJcBC0czAgCfKeEKWczkXv8
fxYdhHV1S8F/CEqjY98GLtUxan7EtSsvAWj6FE3XLYNsnuZvgqy9SfL5bFOBOxkKzieq+nkMmWSy
dwfm1JY57lVCVIgLou7fIkmkPcDSl7gsEP4NzTMLYfOjXkZEvxRzShK4PeKskjwZ4Hbb4ZdemATf
5zyH9GNsAsPYQFU0oA6fm6gopQCr748GkZqXj3SK/zc1YKBKsxmqyV9qo7Sq3REvGOPbCZUpQA5+
UPeh4KPP5OSt2Io3VCMX1GnDRBnvkOw1DYmkOsWQv2ByqsP/X8bJw2m0/FM55boLQ7lV8maOHCVN
T7gNiok0SJn1B07iK5Nv1BowqCg8PVms1qUKalpkvCOP6P2whD5iwb2AX0aD42IHocVsqjXzqznT
0tpNxjDvcYKdAnw5MVONrCsH71g03EuDJT7YJCVSjZ0U+ytuYty3PurZ7/68XHUVOKiRbW5IGOEl
ls5zBAFnvvJHfJP9fvrs/zs61yEZeHSLyQ1PaBdVUOm3gVPBgKrRw+9YCTZlb/Xe09QfXcBTkRRZ
Ef9AOzgJsu/68fyAqdBfk63AQ06y4OFEL8wLmEw5FHjxpHS6Kid7oC2hirGTqSO28/AC/reweZRS
Ro4TdpXOupY57PQnqvyNmXzmbHAZWAiJ7bE2h7ftOe5OGMuZKer4x/fCQBJLCKCbvQJLIdFs9xX9
YFDZYj5SuzbsO31cWJcn8BFblg9OcwQ3+G3VQA1mfhfcyV6gkOR0LU9ZQKemLMQoMIHWWp6/n+Eh
N2RbNMgzcpoxnzZS0CDzKflY7K/HaRQ3tjgv6w6kjdDX/eIf1OUY6OuDqCa+ZLcwDQI5r98DFDWV
nX8jQJiGfqTod4AmErz8b4nsoAfDYeqquUQ3FEbu4AtUcQARkBriuq1qv+AO/ZvZwtrs4r+2g8Qv
HN5Fpdu/qacWiC7it/wRD1JDv5dy+BxZZvIxMbnuPiFISu+U/TnvbNIOfX5LN+s/Bj189U2gLWf0
p4OUZXa/nbwE1WWDdMUwTDboKcjv6acyuPPwusS8kjYHBXn7B7RNboSgJdQP3gFvtHIQboawGCj5
q2hcry/ibsl+hiR2vRgyDhiW1cm3YuKf5Knfiu2xDDO0y8MTXsruBeAVI+jgQCtGc+lpkAmwE6mi
qU7U/h/sKESIONeOb4XbAOPpGT8TRjBTvRWRl3KlSmAbCgU23ORRSvSUy5g9fVqElToJ6bYelP4R
xYEtYlGRTvoFPei8Aa7XH+XMl0aV2zWck3IOxJ/4Wh+ik4LIn4vnIKsPXp+o7Qb7Jihtc22gjAC5
4uHLI24B8n9yjktS2UWoq0JevaNc20kc87ozw58KsSHnHl/8F/jC+8ZZLnuSg9TX/eTQweb4YxPe
O7Hlh/FMqrhDS84L6Lfq1z6kh5M6upucjloGXqwhInEHzBbve+JRLH+iY5HIUrjULsh/1VwBz5zz
zAenPaniexyceXncNM3PohoUkgZ0FpH4t3jAci8KKb8LbyMSA06LZuVOMOkXq9ANpuMBL2tdMTdu
nFRZkicKaN1CrnEXPBHRgop770qR4E+mIumwVQFu5A6LzAkZRSQmF4nJ9Le0jVG3xNdXoiTB5SwQ
mofBM3AKMBXX6UxV7rUqxpfxZo6+zJ07n3bqAjrI0pcYtpoY+USzg2Sv/Niy1MImue65HR5oHU3V
t5NfpC91yHloaDkqZcHlxNGGJpBV7vJdsMKgMhhB9ZW3UCer2Co8m30sb2jAbIJUw7/j4PNybpfh
4lN1bYXeBdSGuDej8w0Ts7x1CJRSA5/9tUoBG0bEWUdUJQmkscC8TlybhO6uXo8znOYgR+sllVrA
NaGQ1wPfrlBmeINQekWrBtLkUONi8EGHYh/S8DY91WoDgGahjkHIUvPJsH+aPTqEjPpt/gJKLsR/
kJD+0aBNy6eTrpWGdF/YHhfPgJjfwl7X64YunizobRw1K+T8kLIKt8wwGLh2GjFMaofT2DApA8Ph
hEKXmnuZMmMYLZW5e/q2ldYlj3oqLgn/nfkCaP7uFA02JqhYAwkrkA7axSNhivPgdnRq9tw2WFOT
voVLx6ONoWxOB/xSHvakvil3lHdKctPL9SfIFQdVD5yK2uLkV0QpQz1i/KXPkV/qLYjaErHE3Z++
1mGYIqKCZ7tYLzXggo5+Jqtcl7rwmLdOT2dDDAss3+B65zuS/7VZDQTiJCkvqmmSqjypYt4cT+8b
b78slMZnHRnoi9EU7J9lSfKnUPteTPDs7FTKQm0gNyqJ0rFkDZ9QxcSp6U8fAnqg/kqEH8AzYOwB
2f2hAOVqrtsAoiLeLJD1v0nL9KI1VsXBF2NNAtKTHDDHnRoqi+tmAqzgXxsHL29dGXd61dqChGwQ
S0djl0+mAQNp52L3x82W5XpdUWOjdunWTEsPOAYY7jVuaGGuxIssk3EMRG+saWMnn5ZuwzDrOnRg
twIKbABFxxLJUGJGg6R2i+/WVWjlcu2q5kkFyTRKm5XC6cOC9EM64DvwisBIfCdjG3wvFJJZIn7X
iDzkqRe/BzMhJCtsKo+pR6LCDkrW9MmZpw39gTyAb8wk5uny5WHKXbROk1OFkz+pWaaLUyOSgzzV
z5b+cUVpTNzwN5mOYj4YPFMtCsBUMezT0HDt4N4rhmt6eqWXPFmsComADInIQeUiPlg3DguqMbcs
N9V/GdaV9s3xw/HxnV5ac/LnJmxqIMdk0JlYGVgetbpGgYBKRDV/KUv8gR9iP0t1+2OiOCpFJIyi
x5oRzWUHsgoKSVT9ovp3ISjvgLxZq2fv/j6IwZ06zpy5RkzHmOPEdsq6OFt7zheBmmYczpIX2pBy
mzMleK5a9RSNUG3wn3GmVAfWvfcVLIStBemngSbMSPvwNNrp1XeHEki8YPKWDBeugLx9Nl0dPOQH
1MZm1GPGG2H5R5z6WAfq7exUccZE9ORGn97NHq6oL8icTMJsHdgiI49m1Idt4sQhNLa/JjCBBTn+
jNWKtZdpbEl3mB1qHiaM41/U3qulUNOQH8oUp2pL99alVGPP+XiLBsrQJ3zoh8rRvqIb08BzQHg2
seVA82SqIeZNIZblBwa2jA3jzWBhGa6b6oVbZ1Cx+aBmM88Cnm4iCJUeQxoQeTnMueFRQrRWtR6d
jm9P0EqQ4SzjctN+U6LoAicpfvZ2CvjDENNl7msI48NR2072ynlX6NXV/unZyd0dF/sIGQPYVqMn
vc8oLlDU1Va1C467BSMwagNO2OfeivNiHq8nC11dCIXvtl7Z7AmGUadNCvacV+7gSE6gW4LxmobX
JsmCa/eEYA0iSZQ3x7RNkIrzqedW7uD1isg/hWm4RQ34mvG/nxp3yDckXfyYdLRDLtPOi2auOt48
ZmZJ8I9gMaPYbtRqA0TCXEu1eEbWLhTSL8/zkeJBxIgUWrgTpFE5gDTcVLjke5ghjUE9gAEtSjN2
Flz0vBps4P5/ckUC0SgWgsx4zQaIi+a2D9Ml/ZWsBwKSYmub9WQRo+XRjB/WCVgVvLWcmT7vwhq5
ZDJPrJfJ6qOHoGoC83gpmmwK3DQArTbK4WcHjFbzOiRqZ87rBFq9X13UkOdrVtEVE7+v1goqrrDJ
7ybc381POz6E+p/aq5cOjPep3Vv/im7WN2Q5oCgPO6BxQNaa1v7Lbz5fHzVPDpCY8uQvWR9kDMpq
h6kAtCUsgIqf88ROUPkiSBZZr0zpd9jY5mlLna5cBcTt6WNzDczC96El2lennmNA5AvpZSM4LsFh
zIZa9N8xKXJRXPesj0QE7n3a0QZgc1EKJIInYyEj3gA4ckJyKh+baOVT9qqm5ruG3pboE2Ef3zuf
M+vfqM6UNrOiwd0SdhH5C5UoZcC4ctSXhrYd3oi928QaC8Doc4wTdZofyrxrXXyor9B1AI0a1PmY
VRvnMS6ubacIFH3NLGVW4CNpy5A+Jgol/xuz0InNNbusfwXLAIe22cwXwW4HZLf/JeWhdplH/auv
kqEbOJ/YfB5RckTPk5Cv+EGjmdcTG77tVrx5zTPxWGGGV4/42KMD1k/sPNEP68azq+9H4neO1/EX
SLonWs3GEcf1pU4tGdOqW/Xl9TOxuiAmxr9WCpvDvOq44n2h8qDlu9wvhiSivQ12gbwVbsihtNBb
I/z5JU8KAqULaCR/IE4741UnUCwXh9WtDzeWarj0g/bnXtZcjsPxgYhH9Aw7SS+a6U5T7H3XKGR4
wVOFS952k3oScp1pRUsTX4bYR8/PDpKdknuXbcZuQPF80OnE3rqO7o38O/oWyvCF2Xb3u1WxsnPn
3E0M/3xUNz5QwVV41xnC/wJhtgyS2CDuSgFfivyTXLWPUosDANz+tnRuORwmULP6lLbuyhsyJ/7A
vxBvIY2EOGNzyLsOatH56f4BYs+G8kO98kk6QWjstE4w53J1xFIuY1AnTXgTiowPCccf5HhevRr4
XwteBtlmvYFFvQnjskFgq8uwEpGLy2VtkvAz5nNUn1sUhnpQJirpEup5EZsT+Vy1RJ5wnjPy+JBq
7/z/JfIRP8hL3/32mqwT2JjsiexVgc/h0JDY1GG1nGqX4uxHoaJormhyYJbPG0kovGlcxzm0Vp94
46GvxXz/Sc2UMkq8C0QSAB8OJgCzTyvaNffhroE0MUb2wuK71oN2PSY52f2z4oX18+6DUwacZgp9
wLEQNOlusBY1FXh8whrDhjYEZy8DOp93KWVfWnCeIQdzSg95EBG4mxRM6HXxuKgLTT/nLQZymlkM
naHyT4PXrmWkDRYo94uMpkWQgQwRSa9l+BG2u5ZAOmjY1pz2uAdLWKY4v/p8BmP2Z59scw6ZqG8L
RidQQxs6fMxn7/jisi2y5i31oZeitlLpUmhgiMsen9KjzftklXSmLvmT07J+x7IYSfJoppaFfli/
pm9AeciA/DJpuZacLpi0YhDeDVYRM8MBLzEUPfN1M1cZiOgra0PzhUkrWkV24EzYedNnGkzlFJJg
zSMYRUfEkNrNEF3Q7QcEXEmlhyOfNsbYpwFhq2VJ7AqsSHum+NGSMLMxNE5Jpe+MkeNn7ZggYRmi
QPvDuQkflbO0ZXkT9b5AyrP9HXnOGZwfUAsgnBUJGeckZOwvfyJK2KLkGKFYC+D5Sg091y+HNFOV
f4vriw5hpCcIT2uHgsSN7iBSLHbZTkaAMZz5GMACr2618nShWZZHuJxV3DxmFjBULBBUk/akTcMq
RWl++GhoCsMwZHIX2LNJ96mRmUTzqQrPxVYYXhbLNG4d7jzI/vA1feQv4+YWFc94mO8D5ai8j3lJ
G2bUWZeyQtwXaaxt5MYrE33xKLi9gU477klBLPfsSp+j0dpb46rM+o7xq/m09dyGxYmAforry3JL
0kC9NiqALlYKxtsyPIb9Mcwvm32lHMRw0FmNkJgcuEhGwiGaIkzqDnysm5mgpZDzkqF4CSp74wP0
vZJ7ckx0VBTsTxVraiA5EGQbsLWvRSXS1oQvlF/ZQ0YqXk234hBqvJrr2YKr3rNPaKGN7OUY0gN1
3qTaAmaxnSgxMfpTcMSmuWjeio2vWuPBvXae1TO3sqJw4Tw9cOw+VbYJqVKLpODno5Bl1DmIIKu/
+DnMkvnY6gBaCc5F4mRRXpk32uL+jtUAW9LbcCMVndqWgyGrC37oy00lwqg4E+BmSExnUct8ix7/
y7DX/9HAzG23DqsR7Q/Pv44Wpq9zKTEFSyHUZ2kCpf0vqavccM+WNc7Novgm/j5NAlkdoHi9b/ya
8EZa1sC7S/8NDqR4AZxM9aZjzXJYT1PM+BtzV7zkuUCKJBjZnFSiwm5bF6nXvkXD7xsCS8ib0R5n
PQ1fUWMUyc5b6/xMmBMN9puaWYjHyVP3ctWGGvAHCJHTgcdRFFSuIp5wd8rd94SmAAgbVB8jqL3R
ExbccJHdTebIMfB61j249O1dLlxhX3SPjOBAu+ezh+sbK+5R5DCeb1Wqyrm3mHYY+CbVGrTK+Fi6
LgrPLLmm4sLDF6WLWwGOz3fDJScQNY/mP/BwnKBAIR9t1Cickq7LdgZDDEcggY0C+Clee07/j7MQ
As0ySuri5pc6tNz/XqqiYwha8K8UqUaymvoiD4amKhRyKaePrEmzoZlk36w1uLIYqOCWfGuzYT+g
4Gl/kfzf8KRVZ3uMeSq75QvF3k3C8orFC2DVSBzaZz4F702PhDB9h5d/Jl+9hfEKjOm0VlBUZnSi
Hr7d2/x9yTcrP0y8rPUI+kjpVkGJaAmVscsZnt7N8dWgtO4soCLvIyP0+wqAtOQ+gO0govF1fg+N
r2Nf58Nqi/TQwMYOx89sedQz/jihS8Zq1hQKCAqwBUiPfBWSpH/I3XpauEgkcPOJBYd3gApSvh+y
usBZnqFgVJYnqEieB9wANsM+z2f8Ksz83DDrC1ysaWI2tOOvfblnpu53GWjNkt+62Ye0mC3rDwwe
g+/PcP4C0GRBypzLNd0ywjAKspGk2Pgn9mRj5Eni73nwR1QTcP33nllfMgLSlIoW2yZB+VZnkrZf
9cYwtjpmZjAI/8soWLW7WAb3mMgIWcvLO/j9x6k35RxY7Iz3A+82GJFMkBNReOpPRlhsJMCvkOhl
a+LtnodQDw8SI40fZwR3N1fnvWjfoPUqG7E3zjsyXro5e0jVA7i/nWAtRBBLkC/K14wUZaewiKk2
poIFbVGYSMl+yl5oq+sZzEqERUCuqhW6+GccsHEFVQpJ3B7dr5cVCVQqdrHYBujHPPdwLyFogDSQ
P2VDSd/7n4xYy4dF6DzGPLYR2nqESNh1WmRE7A+6JPZMcP36ns4kjFspot/8rlQhXn+3cvXGlVJb
4Ej9uJnMCh5EB79LI94u0LRfMXoNn/s1i/eiGmh19O8l+peut2lxiNNyrg8r1drMzq+WlcjwxWTr
PXvUpyNZpKc0wMjBn1/VOWzf5szceL8NOkii4iilFCSSO9vDuytLHoMn+jmy8W8oO/+hFAuPeQLC
kyxC+rAHypoxMfyRwihaADfW0dAarwj1A+MY9DFxp4yFyWwKKiz+ggwWbKShkThEYD1na3CAXMmK
3FOQbUrs2TXpXVw3fZ7yTrzI4e9ayzgZFmQtQIjGheLRnZ6gDoGP97EXJ0/MFYog9f5jGppxF1X3
eoWgaMvmpJpA3C+yhXvFjOQPqxh7SverUunJ+AHwDff5B7CR7qQAl9f3XvGATkvp/EwOWvtn8IRi
QsjLqMmVDtydC9NbEJO4pP8wN8cU1WJyizRTp1au46KTZLp2mgcZEHwQadDAwV1a036hSzWhMJjf
RbQHadoKsAGj+x5B9qzKsIp4zlPg1VkM8pXvQaWf5zkPuqvAVqHNfMtyE5lSSFS+80jkS/Gn3iHy
yBaZgy+OVLbXKJAkeCnKUrpdEWgb5qtPz+pLywlW8/5pHH/jxZMmDsvESbkAQv5q30MzGf1frrSV
VMD0RHWitm7+/kxA+xU2+RPR0W5VxG9l/OS65LpiTPie0aVMlQK/tHI7xuQ6ot9egNOAHNx8ClDw
J4l1emjJHP9EZ5vAe0Ae74DQoL8euwAsR7rNRGUS20pZEmP8nfOyQwqTXAsYV0V/H8cQdOpIOj9Q
c9IXFRYmxJokBgmVE3pS+OvD0kCQ4Qp5fAp7JCmWP/V42oc/ZayEc+av0/x7A0RY2eJDcOWB+Xyt
8+RKz+qWAgJjhaz6VsdoA3EvtCj3vuqDkyny7FLToh3IhqeUMiNL5lcklfatgbOnGmCUxEy5bks2
h3IPxExmkYS1TU4e5Yshw8RtXuZ56tmKLOcSWntMarAxOCtWhkE7HztywbVYFOBwkWcOeC7Rfxsh
Lx18G3eG+O3h+n8MkAgOXqprD6cFqzLO4ZxEDadNKYUP9fRpGuPUxTBUhA0ljKv74rHPfLs+afQw
E9/we2lER58G2eDKW9XKdZB3dYqTsMqOPAZdByWuJAieyfkFuMfccgM36AJjfnmkY3vxmGVY5utx
d94nHNmXzi9AWPvMdx8JxoB8Bky3sDuqEVIsr+LAGdxblBsqMlKN6j3TPguOpajsC4leQUYNMGeJ
vx4lehx+aIjxuRKwmhWR0DFuIjwgy98crCYnq0C6kKMRnhavrh2tw0RaotsbTp9hoQ6qNXUep1Jo
6OvB91robgGinPFYI+GcmUShjLt9L+dbEQqY9y4S2KgKZsz7YBqF2yyNNnfPdEeRjK3rniuDYShA
M1qEYFeBlM0O6YX+MGNPi+ouWYbz/qjXPKK/JRR52ODxDYn9U/CQDvuTr7uKtobbTFqDMOiI9rjm
2uafrahdh9MbU3Oku/cR1j3P64FpT2gYVWvQsSNRe7WkZHaq2c3eFR2ob7/TBsyzFcfXkvuOcQ2J
mu5SeuQZCqzXMJ7AiGsDc+GHAKcp808a/6UR2vFlAQ4GSkyFH9FZGmtcQ1Z09sGeeFQWLxRhzxei
UqSu+xiT/wuciVrL+gQHyMbWUXzoCQlbr+gQs5eVJdCVcK1SWcvIcMevlViYf2OEPJQCuUrFyeM5
bW1VJAKFRX59EP47z4DRdD7c5lr1vAg2J5dQfJj2fSvJ/XIfpukBjltQBq9K/aieFlYg9AJ/8JZ5
XgjiI4VRRh46wyg6tLefiGlsZx7C11NBlkMX/d2diMXAcAXR9+Y2ILo63S7wbJuyI7fdSGLIvH/y
m9RR9nPv8QyMOVKrayEI+XhiistlbyD1werTXKqnEBAdWGRF3pajui80YVv+H44BQXRIgBOZYCqC
D/+rNhQgvLiqiuEqzuHt5+up3qoHbiCfyB9Kv7evMP1WMHKUozVS/FH34/AY5w21SOZZUVcifXIA
2ZsgC8M2FJ9CM6eQSODNH4jYa8UT9AFddvH+lnj9fCZhLKqe0OUPfYzcMo8AbURwOvBa5Io+P7wg
4o+g6AsEd0V4mhu2YnqKFK0ab1ITP8o3Eun8UkkFK6xda9krWXyVDvlJmw38OUSlHHqI/q5A19lt
E85YAe39v1ztuKpjpgbrKrC3R39G9g1ILSuziBP+RLchhvJEBLv3o3x28MynAOveaKNa5br2Mrx/
1HoyVXCsATiK0HMGuohowweF6KRmTYAkKfrdqzK1KTIsjrcXK4WER5uhVRAyhy7rynBRJXuHiTEe
XIYqWhVisyljblL3EU8wvx1vtZAgQFA9Xj7zBfF6k3FYACHuW+gUyNUtzZgUs6qOj6mYPrcecyzL
PL/3tzosFA9vxRTLn4HrfT6CjQH21ulQdKH1wtUJa9f/s5Xgyg2E+mV49uzlDKu1hhseThuz+t3D
owRtu/vIjQTmwPs5MfvXesE6nO4nxgpShszyNYSLESbxQcoKfnrKjEDoUu1UrvbGLCoQ+tAu1+oW
W7K8eoe2A3Vo7B4WfvghI3MfKFTA+BT5+88THEr3AqJXIZejHfHGW6gfKlaXu/LZVjh/G3FIdAjh
6ZCVGLbOo1oyphalSpgp/kThFHVDogeMLjySEZHR3GvuyjE0k8908emuFoi82RvWzqUvM4XgtnOm
DzieYMiVzrIRtLVDp2r9eWT8YHcWOtiMYH3SGTOisSKDNJ7fccq2MHTVo1dn5eR8yOqrfgAxHu1B
YfxIW+OqTwu+hep3p/nzlRQYvXL3szpS/vRPeJiITNXrGTW67LaFJhHMW917zxVNrug3U1ZkX2+M
P4xd0JhVsqk4KaryIRLrnKCZKsgRahR1AlYrg1irUAvfl8v82MQmV+KjP3T684k9ERQo6dRnVT+r
f75WOJ3Xv7/eqpi+9uGT4WF7wvYlKYaJMZ5Wa4HIO1WkyYOqyp10DxX7t/gBbx/BLCxbjeWH0M6W
VixicoChxw3xmPC/ZuvFYZXOPZAmZ9xLms+Z1Zi5WXpdw31LWcQDr22T0tV+VgW9iYI7x+ZDCtMT
043RSKy6TT+ewo+vsQkuFLYTZ+4OFovVfSitzrMxBf938c6/4p0juwq/pKFb5NEzv6332jtbI71h
4ad1BmzPrpDBB4DiF7J+kRYPXMB7m5sq5Ot0E+dX3HO8gxbpXEYZeXJzdkdnuivJ4bQ5z7t8CD2P
tCvnt7HNn2UeZBriLvtRj7icPQprsUi4AoDfMJOsiKBDn7yIxfXMA0Zb3sXM58axrQNU5THGyZn/
BWp6hwe6zOggpkZqo4oCV5AwY5S+jaNxJt9cShO1r6pnALUD1x6kxqr4YfBs2W2LbCxdMiRRHesA
jlsk5ikidebp9EQkdEyjvpP9pgM4YnqqqTWHy0BrgZzK6hCfq4GQ3uOXBfFLldKCCms1BVCqGX83
5toR8PDBQQe4R9t2SQAckeTpDWe+RChYu55RWkC5G4G7HpWuzFCGXCSik2NGlgRA7t72LFOTdn22
1AeMbS5RUFtctMBT4SozfgRo9fFZVujKLfeVxXVjXnLtW26CX6NfxLsEOumKlOaesWPd4QmLbTTq
j5ij2XmWnlp4IipQqUloqbe3KOS3tOk2865PGmEYFu8c8925jPUiNkMOrOSuHXsECgLdXQL930Av
83nqgqhQ1OUIaI8tXS//rTB6Dq4lCjBQjZNUj4xK+tTa59dCW4bQtzR9Uovqh05GkAV/RKqNUfu4
I3e1tl2Cx20PvJnGwZQwxdUeVjYmsCTGjaEv8s7zqW2+Dhd0QQw+ohb8aaWrGPwdQatbZvmKDDzn
jKdZhhSFT7ReNbCsdYrUixtr7oNWdMOy0Zn8jB6xlFH+BIO1cFnr1Am5R/eKRtJhiMXHxZRePurt
LW4f8rF4A/0fvCj8/gYMfK7+fEUM27pLnvX+khKgykY2IX4YRw5IZy/vdRB573NpZOcT+/5grZFd
y2Vv/z88L7AH/QZnF2vPFet8P9wxLHE/IOJWPXwCpf6JtzDPIf8cOUErnSm9zOOIC7rTOZdI6woF
LSR2WE4Z3NGmzMZTop0eGTAE5x0barnIbW3Uwcm7okGmH763llEgoElYvNckOYd5vmdjijFt8DVt
TFOkrvb4NLLb/Gcu5ticxG2mug5dYmcHVkjM1lKAyCPu7hmivrEeFhbCrqjZN7c6AIV0IMCbWl3w
Tqe5LubdgPN+gr4hOwke69A7mdD0OfQePxD7dk2oVMY4v1jXOKqf6lBDX66gnE/3Qb8WaqZXyw5h
4EdBjlXNRayHQkN9CxmscNBNJW0J84YXUVcp/zEmQNSGaT8eA5nuLuIRo3HOTa4mrbe/fyzdekEy
ywMRVr8HMzsaFW+q5BHGM5M0J3Y2Oen/yrJPWto4ekYb8J8friaObirCcGnUQkdC4pUcyTAUnIeH
N9gew1azD38spvvt6K9SCnmm3zDOR1tISLjfS7JmHdCVkRsgPsVAp/UBq9HvMtj/I9vpHUGkTDhF
B6xxK5XUcOq/wItS+3UQ9v3CLjUzuqFUFcdvmK+U46gUXzNCFriTjn4ks5j9Tnd7jI9C/cyJ0q08
AF41mWDeiA/xcgA4jIGSRgJ5/8iXuvkgugC+qI/YuPVH3uACZQ4wanA7lUeHi5HAoQ92nEAfTOvC
WO7MixIs4w9rVbPNJxw6VSSV3gvmjXwNxqKfWHy7KXC4qzX6y8MqzB6HRgqM4Mzh0MC/b1v4Pm3l
G8EjDHMB7pHSnKPEV/T0CoD1fEKy6A8VAwJM91mt7cSdAEo1VWh/reOB2egAfRlClXBsX3UqOIs5
KS0MPmkFQBL9pPI3fKmAbHxXraHNyOWkefNXjJFrxcBCywj4E8YbrJJu9E6UAH/inn5TNNG44yW1
yrrQHt69YWxcyBAtEYhbZmymY1idvD6he6U8wL7qWSASmfg+ZDqNzMEAnHRyH8n5IPjLglipvyDE
iX07msl2F7leh3Y0bhRTpDAE0rsvY2BpTadMh8/24iRNBJzhXV6twENqt4pnp+WosB28Mmnmlw+z
kgHSYjNhKmCzjSKQeOpl1CllcFC0D8sYXeZvqv20EUlVEX+SnsRybsUSrNLt2zjupY7z32aYC84u
lDROEAdFzmrGh+77Blq+OED8iYfvf7FpRPq47PGkYhpL93hda55lDOULxMwGTaeQNBF7HaOP75HL
tsVvJD0TZbN1252tuhutC/j0C4m/5ReD5o+e6rHE4SznIlPKu0zGc+KMME2rCMtXfYyL3vnsw/Tl
f1RW/rcL7qb34dXL9NU3oD9g4b8lU2DphybYy9+xevbdddKTCMDt/Z7aelZiN+8+WsrxnG3ebSAe
TF0V5lyGOuqMeOQbwvBPlTOW6KiiHtiQ6v5UanvnjPGIGyq8QdQ+2WOLtJCVjrwjTw8tcZyNrsnB
O8zTrWOg7Yp38/Nj1heREfxdqp8uaXC+71xEpZSxu5Ki2EcgXlug5fIUZbjynLzjGL+pRAOmt3Dk
/nKCaIppYRRB8SiSktax6xmEF8REBz1pfe4GzFaejFv+PGMqeQW8g137XpzJnJW++GwNKTbRpP+b
6mIIy4rbFGjVGPwFEH6VNNifk0Dhc76gzVvCRPdgmFGKNFeQzi603OFTA9CCRJlSdzVNlsgZGK+V
s3J6YZHGWwqoFq6IEuUPzQv/xH5Sel0Px2R9RS7kii8LUOT8wURFpw4BgD6Y0kxY74tPW7Amh2bI
bvZNomkZ/IOYLm7YgxPnZ4OGk9mz76XBkuGJiD1raJmfBfKBb3GI3Tp6q4sHv2KWPnbicWodsPYf
mS9EzSxibcxxkoj2rPDGXzYhnUUAgv8Koe7lWOFUj2u5yk0JSMCAfqLL2+GO6PxVm88e21yH3KHq
K4fbaiTQiut5V9uOzn8GykTYEntVP/C8/fb5MQD280iaGfcW88eyjwFapFmQYa3f5y/stM51wnI3
e6HXYIclsqYEhOI1NVreCmG9RpDs2EsC4qfT3mkoDVGdc5UHXu74I74iuYK77ePRJmsoKCtEgTs6
cmp2L3q0PGZm7mX7fjdJr2sJ1idFeOhwXeE7lJJeXqWaFq5d5CdVBCjyoXd2Kiu71pMYYiaaMhxe
saKIxsXY5CyUK7ayHywQSNr5RrsZVghttEcS2aM032RCyCzcwP/jvD7RzVdZDWq/RnpDjBVxmPfx
fJat/XkW27bxES7tasQlXLYjpbNwPNzZC0nNsL1zgdcFLWz90XWe7Is4JDfkAXiUe2F63kickBvq
8M5bDx7yzCJk6VSB0vDqnv3C27Q2OGFsX3rF9teOzoBwERLqCo36IWj988PtEbSCeXgTseWHA378
yOJbxy9bb9VdojS/x6UPm4ezem4nhUdHdIPEDJ47AbcQMARbsdUbCAicDPB1Bvn/y/URTkCcpneQ
FnD4PEUqC3O5eBlkbN9yq63xzY4cHiVc3gIjBQd4WPBoqoL2XxgtSxE1MEYsAOWiPJp+e3nhY6Ys
6Jww1/ERvsSgaxgNpol5ZrVRI7gksIOvstFFny1bMdRRMNOH2sqduj26y+EI7/GYkzQWltA1dfL4
sRRgN/xtrgaoA8EBmKm+ePrUvP57MH7esVjpLibbGiOSF7Ipv3R+8dpSuSi4yOe0wv1uGFs5whNb
WrZ8O1Omou9nYKWCGhibZO0nEDeHBIswEwvPZGSmFln+D8kvXQ9tZjiI9Qfr2AtPXDED5xIHTFGr
735FA90Jw77zeXnIdAUHwgwoN1eBP4pC6w9OJM+Z4v+yK1lNlrIJjP3ehyxL0UNZKfaLTTWkIyPW
T1Pi/KN/X7LNy/N74GT2/TnwSWfJhcRIxc9z/JfHRPy5XYWvCywuNMI0ZF3EB994BmdblwxLlMUo
8C8vY8Sv+ZkBPpQjIRM4ZcGuBP2xbBZgynAAAxH13rEdRUxe+ygbS8DAW/Os8m9gdT5XiOXAj57v
FwgQi9tUx9zbtrIHvgNnoYOz7VVsV1RS/Yy/wFcoohp59RftaNiKcMxb9W5GYDOF/nxFDfJrwv6+
4fCOqmCYKlXT5aYLNMXbVy6ueCHl1nn6m2KAj5LhUYP3tniWSTQizSBqBazSN8RgxAWRtEXlfRxT
OH0BKdFSUjS/FyADlLhRQw1GDtfy8FkuAUsFhGW19ogvOb1EoTe8E3HVa5aUPZF7fVZobryKM219
KY0XMUzVfiAhvFZ3R8bSvh3vmG4GIrjBi720SXN1CXPUUeGzMQhuEss1q+X0YdwVwevIlSGZsMwf
k7y/FD4Hv+sTektbcwPyjnXUYZ+Z7T8rH0FiCUm3/YVI5Y5GT/n6ZdAPuqCgiJ+TT1qba72J46AN
qBjGaYo39clwSCqJmuGhqgh2SkEyiqhUX/QYjxYz8rnQS/JxVU+Cd8UdBNKjzo3vISimEYzf4Cs1
0co/tYH/CHDrwVEnGdTrUDc2O/1yJKsCb4mbc68f37fRfABm8Ue7z7LdEnKVbwSCfDwVEHQ9WPwQ
KJqxT13OFjz4QyCopPuda/BN1n+JqNuOABm/swOm0jTA/uXTpF7ogWKX2hJWkz/aVBeILfjah0NC
k6eCSZMAVLmmsU7FScomrWxX7aG/It9noEJS4tIFt3D+ShOrE55fjQ6OXFzZEDRsqkAfesxHyO11
DL2iN2CdUI72HCzaS+Se4nsR59V3UxYSSDKsB6K6RCwLkt3sHhzZCJgklmIQJTBn5mBW26Me/ypT
I/LzktXfsAhA23Qm1OyRGXKTfPB+uBAUMCv9UxX36AoRC+SUdXak2CHSwRNEdLaeKtxo0RG4Hv2d
xJTPFf9S+jmRCEbFp9dMgtPkXz1MpWD6FNr5gGJjmmHMd2b7Ek5BasE/hdwKyXAeeRlEREo2MgxT
Hte/f8xwKScD5qPQlITAiUqAxA9ShAMwyF0WGBaYIoaRP4+F0Zj7lapwebBgDy5HybgbRzKIJaTh
df9GZKRgXlCiwatUWCXvzD+rF9N4G230rUNfUxIqmNlRe9AzLo3Q0HxJYxuD1Jj5rd24ay+vBafF
xn+XDHcUgMVBz6zXBqmohivIxPVmJhFf6WEy82nOFPbMsxHnCRELGiNgmbsHoZXksm6rJT9nbN4G
ql31X9oGaWY89Wm/a6/8AWjjngIj75/tfIYs3PNgZvLoGkS325LI0ULlrUiQVBCy8XBuRhF8AMtv
zCqlJziHJ/1mIdP1c8/UydlXfM4PVD0L3jbNvxPuqTFpdm6ISxEvPsTp4EEJycNmq7baMa4Da0Xd
AMfM34HKN7O4R604ycDB2LhW/qVhoU6t3AU+lHTBvJ/TUHfGqb7mqlKh/WaHu/TpxadUnsPre2Ar
QrzGPpm5hb/PfWKINYODrofPZ145FJDEZHlFpTM6DyE06FY0qYBOgbs6KL+lhJeKtcPdYG+7/WKM
BeJqjQ08i9/iA8Td1aYqJ5LYUCtLY1m1OW9EuVTTZvz4ggtaMI5Brnb8qPV2imhafhJSu60Ag3ep
wjLK9KKAkZb2mkDGEMFBI8id+ec3VtuJ5zpBdNyVLt5ouOQcg5dtYwWxTIcaQe68k+nkGU68mY2g
zEdd+QTMSMwgc8CXfR8J06EIBcVjRP5G0O42tKkwyGTdoZ1RZPkeZL2Xhk+ip/zFOhVR1dhyInsc
Z8feEGQNy+SZIcmZYh71LGE8N40aSgigfqLZ7fDJlmCrUnqviXrato5xjzffJ5XmyOV/NEH+iDT9
UvO3Jexznapcb2lnleRcV5vY4bbnKWUCnrBlkxKwOrs4/j2/yfLd5vP4qVCWIV5cU6Mbt7F3eND0
ifEeOvROora9djVQpF/A3tc9zYSROtzWStgftfY0TbEeCMRFV/FUDudOSsGao6kTaunaSWASHyhw
O4BwzpGmnn2N2L/8tD+WUC2+o+HZtDLXx+nI+t4eNPjRyiTDlVt6UpsJR2oSXhXGy052P/SMM3o2
kzFZF1JF8J72Jne0RQ/3+J+CnZN52GykVJGRhYNEAO9JhNjxN1R9oUg5A6eHQsQaNTtnvK8RDmwf
ejB77sJvaYdq7r9T9whNjiAxQYu5xKJyQsVIL5OLbcV0PCx0mz6W+OvGclRFU6jByqMODtsRv7AR
wL1xxY/vmwRGnXadP4X2BjhnwwR4sG4inaHvqsikCO5e/GGXPia+hvNX+jHzflJYTaO6PnxL1blr
Y4VQEqQPDmYXu7UrFBiLQK3GeyltJSF35kvQTeFMpSt42+Wy3wYdox0dDlBD2n749CCikvkJAQAz
93pJ6FKFJLbG3ltqGMvgW8QH2tpq4Yu2LoyIIc+jEi2xHA7a9kZGm4VqSEA31mT5zjekWVQbeMBv
acUt2qOez2Wz0E7Yt2IrJDhakelcoYpqdXKJ+FNz2vQusy1Xa2PMeS6x1S+R37hyy5QhIm9j3MnQ
tlhsukvtMgOQtgTPD0ULbNIXCAjIDPp85O66/FVhnoogTenNs4gZTLbMu/yeSWHokX0lou6lgyns
AQ/zYonYzYJ4JS5caSirrtqdSQPLiHNA2DlcbveCuQ9CXBmitF1Ruv1EitkvJi+NxM232u8irceO
ugxfX1w0JGXPW/lhHUi68Wdg/wwCOiJ5BpujSTuorY947i2LTJx2ey4Hn7DQi39dzjOdiacdA4bN
zfoEMqFvl10rpbfB5YcVf6G87JUWxhVDBEQLutohK/95h3rf9jei+Xr29Te3bNHGaVEk70rWpRud
HsRVg5h7f14E/f1fthGDky6vsIpeXpMe+k48QAnXnYiVSQTKXmzWYVXfNm2cKUwfJt/iaM70wjYN
PgDLrS9Xis4XZIfpN4lJADeYXSn2Lom1Nt/YzEB2LoBiFTbzeGNmaAyUd9JDJh4zIeQc7ewKtOtX
nomoENf/EzAG0mfJu4LlPFKR0CG9DZbB0B1U5i2JpHWJ2jW2mOjoYhP/qcWhcybfdG9vleldiayK
WmmJ8q2SsTL7XathwK9Dj8ZqyL0AGPOsw+GFp78dRk3asKJKlQ1xhTtKLf/f+ga8DsDVgMwXWnCu
Ltkhau2EUg7QJyllu+ZE20PASRkdq3ubI7idPXoGC0TrTrDkkMaZkJQyBdLRFqjqSTUxYebenTUv
aA8XQozQs8noc23b01nXzaZJwfSUfEtnEvSm59RyAOuDPy0QYej5SNhRTT50U0c3uyJkno8ekoTx
uJwqrL5Q7UCFw8Lp2R5+dBYH2SbJb2p4lb/mnL2X9M/zzfesVQtaQJ+/Zdb2Ttdou5BQKyGP5bWo
cAgNXVhzt19stWW9AtnWOjY7muOocKQVn2XvReOj0ZAfDQ0MGBQ1KMVJ+kQPl+gX4GfyGeKyjqj+
9XFUVpK9tOc1pfshpnKlScXAIPPUCd+TCLUTlnoXaMRC5RQ0BBjDd/biX8gh0WpvYMn1zjHb8Sjm
AGtwezuyMuH/scnKxpnTdzGVkR4e8AX0YCwVFaRnAEFSdgIbhRJT3DoE+lH+DZAmWbQGeOQuy0Ab
Wa50qq655+IbW/jgbU4PewHzzEMXGskgcFFHExO3n9YHv0V7a/kZa4c7hVAnKikwV23hoySGuvre
/nfeEj6eRMOGHU7e5bSwBAN0aU06QT3mrruF+Ws6oPDwifSiecTXMB9SNt4AaXv/33H4v1saTiHX
eutLU6WbsIz7k/HqlVQbKTZgRRJGM6L1s6NYwK0zJv9oZWPpbMQcB6A3xR1/eoMt9CRIDywCc/B4
70NKi17irq4vtbuH+t1YrzuQeRT4BVKa3+1ZxMT/+nm5NP+5yxgbdPwTpSTfTndlyekcpzF99wmN
i5clJ9LisJIDflTTxdwAU/yY1Q/MM8zksyF9DtxZnfyUdciqUHkTdxwovw9VnoK07sWhkw5LppUE
vzOVSYoEHbfkbYitx2SAoM7KQgSSrRYiQIyTX1BbSLZWPifuO70iMklLqLeS6z9LQQxDg9s60PIA
Y61Z5uPIIsaUDSuOW+SuOQ6faEK7g6pY/jfTGTFmE01VIXe6xpajKZQcRPiLAb1cs/9nvowsA6ae
eBAKJYjRFy5udm8J5ed8t4USDtHWBdTJfZ4ZpFCuaa1r/dCJ0SYiy4TwAzsfFIt3DVyZfVij0pUe
2hIMkGIpNcYaCTQKkifHPNOT/UVwLvM5DjTMQXOO+XeQ7XlRLUsX0hV2cXbEAHY4D0O42ehfVmPz
k1Vbi8v83LEcUwg8VJqwD/SOGcI63lZSJ90pAjIj0Vm8CbuBUg94ZAfQFXdn67v7kwl0EgJ2tuPX
OmsYQ/cuL6ebl1T1qWCCP8RScASPZ8MrQJ8yxm/aCbd9UWenKw/XEWX0eMNiDxYHAG3MiQkLqIgf
DUH3AKnWFsV3D4fz4z6KpuVLPcT10ZtcfguMI4EOt0F9GZf1jqLmYJKZGwwsAzVLGrCaSjAMZpwE
4EeErP63RmA4/Hzn683JkSh3chAIJkyPTO8oL/zPp3QzqluJ00q04lsVl+wXVeLTg1xcUeWYt89g
i+S2bjpaAvXCVgZLsbIPhSFvfhaokgZ5kn2ixVsHU/IK0UC4dTT6WYPnBSUcQJYGSMO1cP/mjLMM
n8x73rnynM6oMcg0lXkCUwLHr3FTbOlgcLrzG1uFQUGr3eiUEnpVaitQP7rhcMWwOtWuZXRdcCgs
boI2J9sLEkCUEidiApGf80rl/7onITbUAFAMU4cQbSTdCFtdm6SekUgJkC5xxhSMkIZB7S1UZaMV
V3PL2k1k1LjDetBft8qB7zmSBAjFayZXPhp7xOpsy4sUO+vnqbWU8GVPpel/oXWEYnjLMz2JVn6/
ywJ2WIF88xpMjraBsGas9Shd6kMCaWK5Dy5ptyAuKWt5RBzRqMdE7t0TruKRMtMwvd3USEgr0+VK
I+it/Uu8d9lpAN6InjdO0ezxM40cgBAz6zQzbJc4xXMjFRgGqACv3CnOLIb0TI1OqOOei2XnYsmL
gDfi96qHLlhm4Pn3wBWhRFei65GQ/4IBHzrVFMzlDv5pFiNym4pWw//PEaxaFcSK4vE9FTIEPf5Q
0kuEul/8WQ89OoZM4iaT1wMd+2qdaJQZU3TX6QMbMFwHxj599cVofkI3LhBmJC3O08wB6iIUNC6J
tFQCXbU19Y9YcEwlNsYpdQuSNDSkDikTx5hFa1MBTSwAeVa3QX6yycxHiGwbq/RzDLbfaFGybZrw
BK9sDmvwCAR2IkwiIVMyOOap12RpFu9c1/lN/q/jHQRPxioR9uC63vgfQJviMeHkFTkIq3MlwoTM
meyf0dz1Bd+AUgkPfkd3rtxAvJbrU0K14GJgKalz5gz8leo6x3v9/dnJlmMx5rLToSlvfJaUz9cp
9TTmZDN8JFyVVaYHvK6wkHUFejW08QoICELWCkw0unZvH+r8vSeUH12259U7qCSTJk7Fico6y80H
EqFFb2oED6fu7CGRK1/m5aBJRox4qPBN77ewtmIWDPFSRJJJGUIHY0ukCjFXivQHy7VbbMk3q05G
R0Hf/XHg0B1wlzggiO8Bf4f9IDMi+GIQlsrOjZVImXgzbQS1GATwkY2Fh/ZorMMTfo673Aby+cyO
0uD7frIVRH8dQ7EZUAvnY8Xu0qQKOoKe/0wPR8RQ+tvq56Ol0Zo5YYwe+43Lan6yRP6iCO7r9B9o
Dq+E3LlSzzxudH6eap9bNkNyZz/9/s3Pw9rOyD6XKEO1tq/vbwywPryoeGbv/204qPIuAjSo1vZI
0YeTwPlkVnbR8j6gjJy/V8EC54kRVzSK+AT7h8yWrCVo3bTaVp4GYpItUW0tQYFNnSugBoUnFYQi
2rzTKExvjQ7/lvotwjm16JZT7kQRtUsUUmM2Qg6ykjDlPjnbj95VIE4qU2JISY/RE3gwsBlaD4b/
QXK49DNzLN1FAxRb2KSSRG93zo8/RTdfZOEJjeIfdLZQTbcThYEqr64lD+/jWo1FVjI8JssYJek8
gGbu2lBWutssWcqnXDRWz9kOGLsuyqsPJMcSaja4xT0uNSgeKa6DSKkTcxKPIDmdptCpIJMnAE/7
3BfqryaSNScYjLlwqPqHmaPsXN5AAOSQ0/B6nPLlD+F3rqKvCfn5DQjqSuj61jRotRnwtcv7539+
mf7fvA0j39/bEtu3LC7fcoITYL49XAFM9TdE3DS1ukMeljbpLThMG/yHqhx6ptmEW3Yt9brcY7lv
rxEJW0xe+tlJsyhT2kUgOk1csJ7GzDmH2VfLplm4oK6mJh9SmNS6nIT/ekyF2rqoOG3hODnoDOjF
zlblKPzDIbP36wYgU4/OAJvS//HMeJhf5pjgISEDDBJmovhtMwXeq3yXXuyD1ixn2vnIA9BM+Tog
OXK0Pdg8/54KiHn9AbPdoDzx0SxpGZJYia/Zb7ZCPTm7H0Gno4VSyMBXH9cufegEY5i/gDMqTUwp
8dbqD643r2+HYCCPUZVVDLvUbZDdkFtBUXGEgbg4akgFyIMfsUGcUPrLiApPguMrdH1AYaUU29TP
mdnIzoin9GbnhwaANAmnIrJj7unum+2McqNkK9dWg/QsHlahL/pKuVdfcFEAvJyyjRHaCG1s2QTG
WVksoMf5KL/pa/OkN78GJz1LgTfl2dF7I/9sHRh5S5x93rr2kcR+q71XaoUrFQJw7E4jeD45HWyu
DsgplOG/bqOqkEVFO94X4goPLpTFBYAgj+yQxWK2yQykZElWGkwVfxGGXSh0PQYCW8U3ym+qy/0M
llGN9o/9Ad7a6pxlFdKGk0blZxwxK4WS52HSnJRaU9XR7wdjHBY4A7BhOOkHIsncwXEZHMtMmrUN
IvT2GUlENxchnOXEAFaCZybUmaY/fSjBivRbT5EN3WuvGUDTBGo5mkfAmCmruTNAMNcZ0ja8d7Vz
ThgbRLhVcU3o8Nm39BceQuovd13UBl8Upg1mUoXKvNjGRO+qaKbqVFPcWMvRBo6E8MowYL1SIdIb
+64mv8YGOAVuIirmib2jZvZW+oF7FRPgHnP2B7DC41Q7/p4PUaxs4CdlpX4S3zHGoyPE1MWQpVJ6
H7TtZeo+AN70rKG7txJjv0pDYiJ44arjKz//SMp7uD71UnDJRQQRaaebw9FSUQ3aOOgIxiMrE5gF
tdnIIcJjHFWMbGxhb8cT3BGPO17FgAFTbZE8CAEB5sLoACxtDaqq0b5vxDsYj48zszap3hszDVpK
QbnOBECaLBZlwMbeHF4r2h7Y1YEkrsupj4vA6NvprzXv7iIy6jrGiNBxw1U89xp6NePt6+1NQDiI
FsukUZVtDF2LmC2LdeO8XWIr9VyTgldKS028J65nRMOa4exiSNxGTpMg51kBUZVLpk4Dxorm8Ni4
Ur+yk+1pb3ybdcGPCyeVQrrOCcJjbJ/CXomLLyOuKKSR7IyBzggjpETfdeg8pLpr1b7spV0S1nRA
d1xLS1wMaxduwzhDmHPTlA8uG4y8EqjeQdgUvYjDdw0B+WQ2Vz3Vo0oUKWtTJZityPppzLIFZ1OS
EAxrP9SA+OUNMZPIdE4MzM/g4/miyq7tHFo5LDNIWRFG8quZWBPHkpKAvBW5FU/06kVkPyY7SNDE
i69pYXTnQcnVbFE3GZZeqZ62uKgTUThhJUSrYfMZAD33ozJJW4/GRbpJSjjVVlMnRzx/qfemOQSs
89Jjw2h7yZUDwzXm2zU9kXV63ZgZNL3eBGdwK7k4I9v+7IquAvOZodUFi9rXSOVR6zRJh8O/ealu
VAIzYA/k8D6HGZIckonAY00b1EXsu6HnOJ1URiPyhXfvuOZHiEa5S7SsKjm/uO1fw87jf7htEAKJ
T/Gorff0W6GfukAfuFiHbMZ4E+NfabzPDtaaJBSjDsQZ2KtkwjzLOEZltUErxPglnS6GFunkmYhH
LuSjQLoGmII+g209AuI4JHhGlxi9xQXTjOoIcT4oK0zikyNkd+2qEN54382X25wBY5Ti0vaiKH8R
cLY6cNO+qXXBghlpaYTdb8DxdPYmSYUm9YQGS6tsvMGv47pYnJrqXjjOwW5PQRypk+TtvVRWMeSG
KDUcz43oti4wfJVtiZqNbL8W8X1c5r1taoB/khSHuUQCF5gdD5dsschNmdOLaYzbEYGa6MI4bz4z
nbRycQBYxY6bpEn+uQuHrNXeyvrVXj1xT+i0RmY2I64y4fn7gL+cIzIPnzZLw2RdUHdhF9IPyJkS
/HcQxryxhLCxK88yM69VPBNwwx+iLSWzPOvxj+L/zKgnzNd7rZV08G/HOBv3C7s8YGtnPXqJS3W9
qbKy55nOa3dYosOA86erJCXnJZZvqz5Kj4tb66cKcXyu3Yz+OK95JHakBhD7N9mHgV7b+L8q908S
UI0eAf5gL+ZkQTTLIdyBRwXRONnUFWVHAxU19JC13yXlkB4aSx3B3fhNCU49UzxDK29Vg05pjnd3
nD6i+lpTWsTd56mnLbm+3Ni8tzG/qMLX+j0+J4TeXDKr9jtM60KSvzQGYITrzzBKcivvR3ifWYuP
JuBeTJWghCeodWYIPcjuiqvrN1wWbKHKvoxckUFRKdNA+WbvdynosB//EEG6moen64yOLYN2MPre
8CV9gbry4kVjJiJxVgTCTkwLBeLFGmxLcifnlz5Qxme7G0W8yCdnkQROQ5pgX7xoHbz4lULKEsgn
Hj4iA7UTjfrpK2pzS/BzF85LM31ndWmmbYxeSsoks4GBKrFc9UhXDuquCXJExhscGKtuy3kNPqgY
SVCoO35riLp65HetuoLTBRqACe7l2GpOkZbxsgUbjKUa5tKueO6pZhIdkasiBmbHxviMqyYZZAvS
4nd0Z5g5O5A19U/4aeqET0164mpOqKwX/dCngYNkbhOzqIrHAg4YqyoBmvUOkrkHv3843RAN4Wsl
rFGC7ZYfflaNM/L03DEHIBwnp9364PPiNOMB62E59JL+8R8LxemWGqVxzJ3rRQdIt8n8nojOlPYu
HKfGtYptZQzxKZPkupQQikPYgArt+eP6Xl2Bhi1V1ZaifZt50q8yLjVE4r11AD/uITTy4Kl7LMsR
GXYajb/BgNDWolXIRqFeh5BFZjKIUzcIEBjSKaQyE2EFBtYRonnqONiG39nKy9b5/zLyWLr17a/C
Xr8HFfzbeoav2UHZCYPhJwXvgAFp1DnPffOTh2U9vnRFLbPn/f22tLYesn4rFTUyYkTb3MyY4joh
bN4pkPGp3KeRpMEohaRPNKCJs5hibBtN8a5pN1F9Tu2wIbmr12NRfUj6iyzwsZVNtrotCKwYViIV
OHwqXOzPOuo2KnF2H5H6pocdRk5xFen6jq4aoWXKuqasaiRP6wzT3hgU44NAj9P331YKiTrcQWBC
6jpGIZO8cO6cCwR9Z2sMJwnXK4VP8muP3g7DwZAEhE+LBN3ExrSMWEi8DjwthYbWVTLVT0lCATYH
E3n2U4cmj/TmFOCHGDwQSYP0cIdm2SExK5MgpuBHZsULrK0RHPOeagJ3YC0iqmYGQH0rNPEEUL9I
8oOrU4ySmmBJtJfO+9v+L/KOxKFqigDHzbTAi2MR+hwJhxnWRXSUyxEJgjV0fszgH3HDsV1aNbC3
UVFpFePWDkyJDBHBYh493mSo30KhfTP2nkeFjQS8J6v12qoBenXVPaQnF9RMnk9Y/pNLk1eI9/Wv
08RbJTZ1CsSKtyC2SaH7b0JWJZk2n5XX/fQWcL03zXhbZOzQxTTVc4nP/LDV7kA/4Y5317lTo564
B19VKHURsvwFvLCjwxelqq0fKJYSY0wZ+uVT3O0R4aH7B/gfVfMpn9xh3jr5JpR7p+jZJuyPyrWZ
Sr1FRujE1vISN0B3xMkh/BGiN465rAd+5loyF6uWIB+59DpzX4++peAOTXRT1OTYZcynTMzBzgm4
hRbmoa1Z+/u5nTAtZ2jACo9ojppJ2lT4l1zNeRtDMM7j9FU/ZfWWFlBUOnzrlXM/Nuy4JDKAN24i
SZt8x+NK4VnxICb8vISz9EyHI3xZH4QlipAo1rU3bw/JDsxbcFYI/o4DIyEd2GIehqqP29FAaoD/
ijvPYg0exEzwnUk/kCBeUoxqziRFMIiSTzDcniSgVBEXkOsuxuyxQ4TUbCvn6JynmwI4/J/vWJnI
+ErizvnFcmDXZSUPA+Emzgo1kL1BgwozdoPklRrPUuMiY7oq3T7AA3mF+HDth9vM4uVfGBKMyCHr
GYIY2BIKNbM40V8uQW4WudZ1H3xoJuxG8Ioxvh+lXZ2056iBp/Ai7+NBKFfLCsTa+8rT+A+PIDOF
3JLtBGRDTj7lSEGULjFJo9BmLSehXGckCZtdsZjh74T3mBs03Lk5N8OR8MQZhYQe1hsM3w0aAKUe
8+fc6RhgvXCu10hNX51wjWaYsmhjAUBH7dl+8JDWjVaGUPanXDJx016F5H2sLvl+HR5weQfZCHQd
F0t2ASepLUksdqIVcV8DuU8//bHT4GL8sOlXsPiAao2OkePbQ1lVSRCMnpNl2uksH1OOWMj/G3DD
kM5UQYOy0vNah1Uhia/NHy3+TnqeZmvsNYZwxu94YspzXA7eLyiQ3Ns0dJIKIOYhPwyaw6N2q/yO
M+frmYbR0iE3m5yqOVQ0hlDjbBfe6CuEKbfxIwJB94pDS/rdhaAua/iJz+8MSNIuKjihvcK2IeJy
TXyC+WIRkGmDb7EYIiFnnoOOy1u4tdvzIWmyKR431/BQxdtR5fdhk2oqOsHTpMTnoO6Nj4UMF1e7
yDMDPra1vWqqn+XdxlSXFciTsJ7beCcg8WCdkPO9PEJunrE/Z7KkvvRSlAYO3aXAUnhkNjE3aGR/
2uqAJBYZMaCyvR60qhP8GkXWFUazmHU8Rv66NcNlAgWcrlfFHNfL83H67xVzmuxZFKdjDyHM6gAZ
o6DW3Zx2T6Db5xKd0aSmbOM5GT663mI01ljThYDwVF1TCG6JYB/1F1UmX5HgJB2NcGnRCgQ5peLa
m+oUBqA8pvjFAFQTWg1K55lhHR6eZD431od0bAp4Dh2FJNPLyrnHzWhxjogVRPWQ6RJnNiZrG8JO
992O3Jd1Dq2rmTaZpU2XdZAh03HH3Kw7aBpqSRWd8a2f8euOB/rz4P8lZXHF68ct4DKktdf5a9mq
gouVyfzBNa3bVoaVEyNcSHfefJc01cFCRd3DEOp7BsYJ9v5WtCSUeoG7tW2rzma35huTsFwHZg3l
3425kUIR8W/H11GD6EVSFF2JDhoPjWvFZSgwBhx/60OUjE6nY+suMDBI+UB+1fvkDPB0P5qrZxtY
SpyGeFHe2/QA4DR0U1zK6zT/4zQ6oUzTbIpSTowZSPvUOmkR3ZUO39RYPAjNehKp+4G/OEIlTQ56
gXkqRSaEhhBa7JmmfEjUouhULa7IpJVh4l02jNFSNvXQmbVTM++rql8z5VLiRizkL6v6uV9ikC+D
eVU7XQjxg7/rQzGVZBzQMM/3iWeAmTiZHK3+4ZUK6ij4BVhCWXUX9ZrkbFtzsauDvf+jzv4jxW+m
yj1OaChxazCDn4CrSoapdFaqPuHlmq/nM7QO6CjUrEcFqt9qmW6jQzxQvGljA0fKeNKuUelHfFs5
VHHzro3TYorfJtMVTZHsk1ipLYqF7HxBCfUDaFgdiK2nf2C3oJCIWDm7tRXzfiU4FmN5ZZklVSOZ
28bFIMRxlFigQqnHnjU0hasHcxeGyf+bpFkF0ETL+ExWaabj7cHJZb/3hd16r6gDfns9ZnB9JCQ6
/I2tyz+I4De6Df4zZsFKhnn85kWfuM6+jf6t+0eYMpwKENqfATw3gejqRXUgjENcL9eDsZots4vE
fQRPFxX1H1WJy83lk+AZLh3hNalgsjqMtCEr64TpzxPi5C4bC3DX5Uk/gpEo9anJNRsXp9aHaB6C
2R4JgilI/FvEBNr09u/5ok2fjj9Z+C0YSXEKSQTOFkP/0hrDUoA8vs2BrKxpkz68ZEBd9NGIyJt1
KehP5gHdBU4kwREQpF5Q5gUiXE0Tp4WUBRxdgbpvQkd2ThHeqE+lLB/dB4W4nkhKPYwNY+pZXFDU
WAp4ODxiF/Ck+rSoUVjSqp6Lx4YndgPWafWUhyOi+6byjVGR0v3eZV98uckXD1JhvQslC4paya4S
rrXBLD9gKTGYJsKTrgmVaqOSBXVj3CigjHCON29Y0pz5N6rxF7PeI5KUVeoPJKLRXX4A4gLzgA51
zGXn1RyI9PJdhlqmsTSqtb5mZqDaYCrVEURj0jd5+U0/CA5cp8Ll4aHETYyfHNF6KxvAgy9pieQ/
F3muKlf10MEYq8gmwCYe3eQuOAVjSOps4jKBfU4qXsvDLtG0/qjqNSFsECTmA9z6PMLk4O93Ok1q
NvRzHnvwptyWelu6zZc4KYpz4ifP7m7vSEJM7y/EbmCq0gVORSqoTO2Tvf6qBYOk0xP2c+uMmmij
m5KDJVciAoU+3D5sS20XgdD9FhNsbOU3xs08Ktd2hiUF9wuu0Q4AaHeUVhh79YBmBR5naW0cllBK
rYzIXpPIYG67cCal3b9VHSp12rpPAzlpz2Eg7PCDulbvO/iWTGUbt7pT+vuyn7FUbfml1HUXKUl3
5Zqzb+jgHeNjpizD4PTtqDU+1nZ/73/AWBmUkNHdGcijT5fqRwlu1O/hz/sit7yORq0oqkUth2le
GMbHFAfYM8jDdIZXHw1qI+Z+zM9gB0e+j7HdH4W6TJFf4vLGQQgnYLAVfmiRuJTpAiXknU6yrZsk
h5Y7557EsaM6TPR+B6QwzPSzXkEPJGBIjGPR5i9iZYNL5SdORSPY/JrxXZYi38BMbi0eDM7o40lV
7593wv5d9cgLMI7VU/1X2ap0+FF2v3uiYRjcJJ20Dt6QCedCxWOL/IX5752kCTm81vG398FKCQwR
vUb0pG5TYyvio9YfsmMvWlZBZzaTP2M9HLAaZl8+qkIi93RBnhZyZ90nMbuvqp7K+E/DIJYd++pE
lo7HIqqFSOaRrcoKdrFbgdT9DoMssAFESxiJUX8sAeIWC7PovqzQd80X7qe3ah8bqpVJi7t72O7D
0P9jCCNH9m6lvk2gnkncHuGgS0POmpBhwWaE3cy2k4D4FVki4jx09YDTlh6sRisxxXpGAoXRWlfO
JmOAO3BeBRs8vIpfZLjPexjIbsyfDI8RAOTFxin/TfIQE0DH3uCpZM8SHMtbB9SlvBTq++7ykuQJ
QK+WCX0ayRhgRw2JUDphnUXFoVutP5NRK61Pd9l3gCvMxT8VYnVvxj9mnzgkC7NmaW9kJq0BhUAj
riSBstTkOQGLiSstCbYlH3px8EgKCCZPrIhc1r60l68Eq6M1xhG96l46KQDSn7KuXw6VWQPWiIhl
OiIZrKKsxZ13imySEnh5HJLXAqeb7aairHZZVJoEOH++dsE1sH/FQM/a2TybcbEoTzQyL616ByTr
o3salJqo/5v+dSROhGZFHbAWwSlHf2iyYpoxuBqKlXKPlxi0pmwhFjkr3etlKvcbfO1wwm3LETXW
cS8kyh6DWkR3Ra6LsX/Vc1F2vdd99tJFsxUTdjtG/V+qAJ1Sc/lcr16jasxa0UwL5ZhsTa4G4n9H
avpy25n5IiQNkjOQR4n1+k/heGhQUv6pisMZP9UU6VKEGUGSRLE7OZLWn421hU6yx8of9SdtJ6sy
0xC4GY3a5CcTBibPQpivIDML3iSmmATQwYWbfLCzmO/a/XsVTkIszSqnb/Zp6ryaZLw8kkeULhF6
eGgAxHR3Psxtxk75kMVAYBfcur610w5FaLgaZu3gLIeg4wt3QMV9vH2io1yXbqA/YktXCyVpzVsb
Y/Aod5ikNRW6TnIidwS29Ch0rfibN3WOCb6ScEtkoS+HTHkNVwLJeXVpeIXS7670UJ3Xagpu/EQO
4OfwLgUQlmT8WZS0KdFEy2kuWtVM4SRB7FVd4KVSOSKAixFhyE6Lnp3lW+z/Or6PCz/tri5iTAo5
gsaH7khFerU6KOn/Oi/YA8BoQ+xJ8Ufpcr8mNeqwYIeHc/suU70S3fbgBe7j9EMlSW6teqTwaQVJ
J3FT8j0I2+asK9z6e7R28uew9zTcH/FNxSN9MklxZJe4ePNXqxKYLtBlnqZ3x8+kWrJxrsgB0gn3
jxNpCntl/wDJQmLo9AIx24IxH3oNGApp7JNa5hbJgFNk+XV76okk3cphUqaOLjIpLQQT6OQ1Gp/5
/bNgHvCN8AIq6c5zHpBUgGwxYLLMpL+6qdXXDdwQ3BOMdOo6n4vKEz6LplkI/7sNcH/INk6xF2VJ
HMBPei4zGesbKPhUes4NjAc1Vo492pdPMeMwIQnZMhoPMbA8Sb7/rSOj3Qw9Qzf2lwWGOwYdi8Cu
BY/vbxDO+syGihHoq95GxAI1IeKsziuUXqE5NEBCsmJCh7c+WJ/wCOTjccS2csI6Lu7GqfHlU/Mu
7nno4HkTRgpMtdt3fg+9eeSCgM9wzZ+MdAn53IqL7A6janJzQN848o3A4fuVcAkJvqi7MlsaTNEd
xZ2755tROBx2lotyVrYPErhQw0LdNwRak5kwoTmKP/FGSgfffl2/QhB0XSUW7tcJj8VmOH7NpA1+
s0OHAbwuMWk2oZ++e2gxdKjQAo2wVB15F4PjEHeaxC5r+M/WydXR0api8MLOQZzy0+hB1lKie0BJ
u9YI0HaGGrMAwtIP5XA9LaGbbUjK1rihBbe85oRNN4NInhB6HWdpPBZRgi5IHjWsu7lqTf23o5T/
flMg9Ty7LxVkvchfQjZFmemLOwP0c7YORHLnOWcejmj2fqt4bYNXNQAUaZb9vdk56jJlKEPj6Zq+
GiU86+wx+W+TUs7En6ujnjF0hlIR68iY3GLvYa70mCiGVPJs1CTnRpYg36p40pEtCeVTAHUH41eC
5y4Jyw4ofZFeEhIf83DsfZACrIhuVpI1GK/A73skT1Q3oTCGtNscxUpvJXFyUoafrz9l8wnfdjV2
I4jJDYg3NSlKESPD29VNps1HKmYVXA1KE/ewa29vreyWJ/r0RC60JwRPInyq7cfX65hDYyNbCv4R
QC+icPgG7Q8CsXRTjvEy/72TlEGvoubZU0641O7+YnPAeM5BsK/JfGef8JZgNxaZ8uHflCgHEMww
05pPkgM4FPZRNUnqg/vfE2JNWhowXBxyS8OHvXdldXc25Oq8k2UGalmzut67SbOxEQ1UB/v0nzu5
n0jWgvHFzDbigP0ZRmfuZTXl7MEou/5cY8EAPjsTpkM9gwdVkBp1hXM/p3oza3WpohygIcX461zH
Oq1bVEvLB7aNYN2EbI4pgRFhzvz/oyhmS7Hl3JMPeyzEq27SFdkhIae5XNB5j4Vi7+DRNfc7Kk6m
jOKwQglEtYT1Y/O3ZrhMj6FfG9gbeV15l+Mr7/Gu932sdOQOsCaw9JrHyf2r/9kRfLHj56QBiEkB
Wd81hWrVv1aJ0oA0HT0LUGifIVZVcnHF3RjNmA14h5d+yacFSNca1602rf3p0KIca9Vn87naWqSo
DXHKGJ2cuhVX7emDQWem1gSXTENnwuE3U8cesI9zLmR1AAfpQ5oudodlGp1QkE82jPsXq89AWloz
QihDtXqvDeBLvOrUjicp09bHq3BIgpzfXtQEd3ncxM1WJEhopXoYjcpSLK6bKU5qZhwItFMF6S5v
JrGD6lW7ooxNeKRpLosT/u2svycbpB9Q/MOhGOt4MVQNgvJKlwCAucfg/BrKQrFZHKHIOa4ZTCBw
UeqJj8cFvzAd+Te467qnuJha7Do2db6rKUhYiBboaWNPgyM0N65jzwAVMt5geqwRSv2XaaVn+1kF
bXgAqlkfJp51CQ5EjiNE9dQv/MsmsyZIwGzFiphte5y3XBxzJ11eIS8eV/lAkPa7o0vYvNEPZEKP
5A9lu1ZdwnyFTQR932efhvngqlORMGExnK5UbGpGactwk0lYXziW+CErWv3LFSlBoFB16psgxKeA
l3fgpbxKD+y18afJmoA3NFj1sB45BGpkCIq+R+HkhOt1JuU8ZWtxyU9CnBMvElr2Eg46dWOPZqTY
6xNZAp3zr2X3dLtxi6ij+AceyqcQsGeku5T4IowrKmsX7NysNA8wo4pNYRAApyfmrSRxUBk6/vkB
h2M2jbMwJHqyNBcZ3YzgMmYYkW3xzD0mnTX9KyeV4OpHS8iA4lIZdBhMkrGTjNV4DN1ZH+VD91UZ
56AgXYLSfK1XdMujIm7T0JzXFNumZDkr9QJQwWKhacvnbgbJYTo8CEHwnld4/EcxfRwBzOJxnpjV
Stn1i3OruL6kol9Mz9ClmUSfP0/tZZNsgkEXW+hyaePu3+FGIbPdcIAlupDl071YaICpT8fO8Ag4
KmWS4QC0tRLk1/fwr6wG1dKK0sTuHj31yEx8ki2caouIEDQIWCVj2+feHp7LhzEdpEMxk+sfPSLZ
DJxIGHR/YK27MAwNSCC0plBgdu3XpTf8pMYs/9NH6FTTtvDR14alD0ZTdcG2jr5HZZhqJrDkVfX0
CF8X5GpHt0B59MRBM7KysSSUsdNJmaxe4jahjS3Yi3XiGbnOv3kI1lmB3wX9YOYTrrilyI+2XkIn
35+aDhHGHI3+5NCGXQCzFAc31Grau8b0XP2Y4ilkdJLFz6zuGaEtIv07NnBNedTVZw19q0sLpa6D
TMC4gnCbsbdJnB6ZsNmBVRee9Y2RmSSzlovRg19K1cnP4Z4utJoQO/9ZQsZECWZ10fFYUPhR85ui
2GEQBC7AioRGYjKnFKMb4/LuYmBOKYOSal5rhnnDX6CFHJXVAy9qruJnLQXoiw3u/LhDmXRvbsGp
nv5mOqYd2uqf5mVQ4K/BqLPmtJEJIirevsXt1u+OoAw3434COTml43FybBpz3cQIeZCKFObi4g+v
/ta/UA9XwT/xCXvGYf0fbpUynDHEPwEHwyVFNFZGZKeIZKpIwmtQ2MbjwrV4Y5xn9sSQ/S1GRojw
khtZdaT/323+aDDa1lhvMfHbs2YGEr8z9BQgTJ2pdKx+5RnBnOrHESg5mix1LCGChloEhgZ0IkCI
3RAwd4r+cDAlnfNYKNo5Blj1xnLi64lVWd+nu7gtK+JuVAf52V3qyaixekNEezovE0uBk8a1eOkU
GQasx0KFcEmGOewQcDZKYo4cSbLVVWvhErAiniicGfNiO0Yzwx3pGdYfKGFeMqM+cbiv2/0p6/0/
4kfJ5mYO42EHhjnqBMYko4SlPM/RchKCrTMdixDuxYOFXieMPxrRtpQvsw5fOKoMvJHakzjM8k5Y
hiQPlZQQqQ0ru9qoOH6c7Lqp69S3K5fwd2A6Q5Aiq5qVqF3CQgZVv1Iba4Cb+wn7CAPny6plac16
+kixpqX3E1d/t1MyRiod77QCsALzvNarcgrtIKqXKcQz/x9X3wiebTt2GqLTiQBlFLf2G6PI/KoH
4cFwjuV1fkT02BkO8EfyvzX90AgS4sC9LJkJcDYqmtM1UaJNreKN71jNZMO7u8glUmQSNlhN/Thx
+VrhXT1WEemWgRlE+Ph5NQ+azzU5bKnU70yp+V/WkJG/DyRWjum6/KGZBO6+tagjIOAukr/e8I8p
rZS+uQRhyso7CKA2F+UXSVk+xOhE93yZ4ae6yq434IFHEWcJDAUOwEVxFhaDIOn75kyTUuJD5R1W
sxBp1mfY4fSqx/dzEQ8nNcmBR54aSPWocbSDJsmJNNvlN//rUYsTeL2P/Gxl4gHKl+OfxDqaZvA4
Uwv89IUOdJxeAy/FGB2vrakOT8p2RPzaay2/OvVjorWLADQWouZFPwtGFTSPgWTxoQQDQNg9/f9i
FfThHrl/qkkLq1uVBFMQCkMV/Q5fi/SoXmqGsQ+H6JUBRm686/71P54uGfIY9vjfh3Y6gcCx6J/t
gjW9Tjns0VEd/+Il+iQUK2xdltolwHGqCOoARc295YW42cI/X/KI3Z+ZGwstgYPoSjy+ENfbcyjH
t9IFF8keExN1j8lqVBYt2lbTGNDKly8BmV4sIJwkg8rUd8PpLbBtu1hO1QX0NwaYlPVN20m+9BZB
K46xbiWznLRa5NRzfhK3KM+VQRyvWrA5fnisSa6Kjj0T8jXGAMUeXKBUoIHojm87SlmB4GB6yt8P
Ja8gOnbfihQ9Sy7nyXakHG8Vx1WqC8Gbws+K3AOS8p+/skP0q80RCCly3xsKbZFlCTri3XTBIZ49
uHGJMyb8MtVtf7K2laC0p15Kz9OLaLmfZCGdxOVmBezlzYbfK35X/Iqc+OCer0l4ZssSXEQhfxCS
lJ9h0fpOQPGLrl5TwU7TQIZJh8N7B/i53IBT+1IeXgQU+tQyfhAU7qfayFR5De59JRZBhbsyqTGZ
fUBEeAIri/3BSA/1ltbIjWRYgtKZElV80bdxGipaCDTAy5QT6mq4gVL96aBRWUYJPGgdG8+5eD2q
JOX+E6IxhY2ya6M+Vcne8IkrxhA2EE87izqZWzYLF/acNGgt9xvifizQEgM8AKrkV9X1gA1itKlp
n6Y0MY72L9+K8eX5vYK43zXqB2HJYwME3ikS20BBEU0JGyiIiu5x4PCHOnXWSkyIjd0ddAyVdeZw
eyqt/BKhaSLCZNowGNGBSjAaOH3qlpIT4fVODqFg0n/131i7JP7mW8njjKgda0vv97k4otj95SeG
D1zxc3Bi0CRzCFc6TnaGHU71ZoKV0cxbdIQRbgw2lM5LkNdKeM2ekIzH7ijXJ0mvkTRrTwAyLf7H
bYmeUL+22CeWeY89LVl3iIitUtSpL77ejJNf7MQNVfNi4aUlreluPp/QIbvLiXHRaBsAqBY/kppZ
/9Y34VYCx49PeGS5Bim5q5c29nGg/CY7S/9UHfrDarrWIcYLjLNl/MMVvhes8D4BsEc6TxH24q9O
qgyQm/r0XkE3l/73C/75rwrKRAYvcMXSzQ788rVJmDwTebUrvvLIrRJDus3yKdBCHPkQzZnHIqBn
wtUWTTnaAsJA/wIc2B07e8Z2VqVjTKf2xEZbenYJvSDFRDB+TgcFLvbil5wIlfDTb/jNOKSfR0uj
rwjBmDzclzKgZHhXADW4Z2IEjUlEc+DjUSOkB4EoKbmJGfnfkesV/TqVUd6LeYy2D5fqdTEThYHn
vmWXMsce+t7/JFUIrMEd4ypIv9uflggb4u08hax+RZOeTgySqiooRpve9k/qMXgWHwNKjTSANceZ
6ePedeNgKmWkQ5nf6EG9jCNSKVYEWfSIqoS+UGD/3Z7pABMWK5v5H9LBYFZOSJuwhvNCXH2m3eQ8
OKrJVF6dulix9ITkqcGk5Nse2aV6diDKstKLy7fK63Iv0Ph6T/HbH1tyA+/LOlHAbEMKp9QDDtWy
jJMrhfJ6fe++WCD8WoZLuvN4GcxQGmYPgVMM4afcnlcJya0LIKhYm0SNXFYwg08NuWONd9Y4IkZZ
pqPqASlexLoPCRloB18QJSXO1to9OoEnslagqsZrGNW3+7bAQCG6Czy0tWJC4fMuZSQEcZOLOKxA
j/2OoM4Vzg7xY/MgfePT2zZVsqWJWJgHAq4n71PN9U8aOrEofi1yr3uAcdTzDaKEa3goc9vpWe2f
1qzU2VXBs57QEv1ecru1hrI8yHJ+GerGsM9/jdOydO38ujBymuZil+tk7+W/UnEFXtfmJZ74Xyg0
enFWr8aFZTKa5BoXO7eSxQAR75ALYnZUXs7uvMpqz+UqEYe1SvT3+iaaaJPco7ob5slflQQ+HKKu
r///13Lm71xGdbv3cABXVrlpdxwL3OSlauMgptoiZxr8zarHeRWFhalwL8TI8k5NsMpRnLCSsCeO
nC42w1yauxRJ3+zSQHPS2TXZeI2kbnku5qT/x9lOpPEG9CoAgM2zcMlFcW7Vq5kjKKjbNu9ixizV
fAeSREB3yUkRI3GUD7qDFSoRL4mgGLUhztSM5SKF9HbWqdiAtKBrrTFZMpv+NWJbCeJVsSSeD+bz
Zlt2HwGNfBsK936DDvK399rfDvwtfLT3PCVk1fyIxQtNSdGZqPfuG9WL430ST1B2dp+jk2lrMiaD
BbuCMj+jhXWIiJZTuL9QMnZX4mK0HzUyD+N06ySgxdGXRYizl/R9LKOlmlklWX3V2SHmC36grj9q
x0kL117qKV6WK7YfQqnD+rkSxC66msODVcOei1TFQmn9viF2FntfxA33RSU1WoBvFdHSberVjwxo
8a4+jR4mc5NXwKMLKDhY/6eoOOWfdm4Y2o0QZF3OsFWbHFUWWJXWQRcNXR8hhevTW3JLBl818p6d
SCNtNRuyO5FbUP4imdcyJ+/wlMylMzJvSq0am0jARezeD7z7F7vhcNHydlHr1XNP/Owq6+Fg2Vdu
I53886Hxxm586+hy3d7nzcOvycx+JZq55UeM4h56gsqWgCRtQ1lLrK64Diq67pybS+dsodpWgJLF
a7BPa/vdgLgsIBsUgK/E4TrlGH/XCPDkdjvhGDlXyFOjf6C0n54fFMyf+3awSae2BFhy6Z6YoTUU
+zCUoXdivt7DRu5y258pv8E7CoYUt0oJk7IxB03SUgxAfV0WM3Y2u4wbWYovvAIKClOlwsmIQIiz
B6z02DR5hTGHMCVhLXRmaHY+osVKVQuag6rogyv4miAHymMpKs22srz5+j2743/G4XV3UQaoGgt6
htsEHN5FVBdWYmAKz7tb2JkM3T7cJIYG7Ljlwk/WzLeDDaTR8tSNCoKgj6ElLD6PH2e6RB8rWp60
5n0JjjtlfgK4sNK1t/v/hjG+RlQsaAVkJvNR/BJ/L9avyH+x/3Yq2i667XALhys9kAfCBY2+ARl9
KOaurLA5PmBUs3/ZItLimE5zS0lW+qwTCspCYCLasUxyRDD6N8OATZiPvo0zWVPteDc/DV4Qprpp
iOSzblXwzqZ0DONi4yI1tKihRUdk5Ndm3ECIftv5KC8a2j3srDigIYtqufas3ClB9kHxL8/KCMJM
9YVFONWINpio+fAQp/8srngMNT9FO9yavw6nuwKCfspAd+YnaW3RgXPg6YKvbXgieUP+P73v3Rkf
3ymqllHR7Bl6WBh0NZNdOoei/nH+S4vxc+3O57dz+Z3Kod8p1oeydZcVqc6zZOPD7LbpmBXRVNtG
u4oW+lQQ6qnAwUE9JkxRtsxn7YGg6Gyc95m05rvysqjR0E+SOWYRA87tquITxmTydqH4GAsZFNhD
nFgtbYNGSTH9X+PqLoFqn1Df0z5Wx8P6mlWqpwk07YsskmeK5Q6Vljv1/W1lbiHPN0RehGqDXTcj
l8NkpgqKsWmvc+cnJ/og7wqys7tJZhcBdWbpfbgxp3UEO2h8Rkpk0jXeIEKPocAjl0EK7JhNuilf
tLHfudifkOUa9p8tid0G9RbYwiUz5KkpniK1cZDsuDlYIqT8SB2NTQ8Zuu8KH3sAyPt5OeMSc27W
ft5LBEEgV4KnW6Fp+KlfYgF+Vxrwmbo6YRvIzfMILfU79mWWZ9QhhODTP30FHp5VtTVIO+mNrEGZ
r+3X54h9y885ahqJU8qS3R+jwz4LdOy1dF5a2si/UW1u+N/CEtDRJEn1aTbZzz0KJ6bG0nx2MJKy
9PB9aG0RRrsatzAiUYCic4uOg7xEPK/FYXyarhubBiUo2NGWBgQmRwo834XMWwinUxBjR8mxiR8S
RjT/JQTiLWsNWsdhMQUzFfjwLAGPtvRUh42bZ3mXzB7sftBfbrn2Je3T2Wfbbuk/Ppc7W5W0U/uf
KPW0o1wpDft8CrEAFV+R6LoB1cq63I7Yi51EmmIfT/7rVegDiBBm1JmRVrlLSjd+XNjtGUchWTm5
OGIia287nbV21y7qJrHN3VDm9yEGXIpxqpVeowpy6zkjLQ3yH5guYpUcvybZeje2NnW1pmo+97/D
sG19p44IUjtqTfBOg/Y9omVxrc4KbBoczvIbBy1qa8Z2h4gtONxduaNOYa0i9BavZD+qkh39Edho
qfF+1kIEzRwAOW7AsGuR0lm3fmSceBjH8syU4sVXR8LeaWuk5d8dCQlFPd3b71d91GNQbvijxkGq
vpOHPgISU27U2l3odYywniwLbXisAXZOU5leCEWTcKOow+C7dkiVOuZsJ9EO3JVd++lWH3UoLAmX
yBJ95Y2mR+dgpDm6jCH7rVnM2cxSe423PjXQizSEQPjG9eRlrn8+n+s9ARmGOlZlsHiVyezhl6+E
UXHTNfTRiJIXFIqdmrwxb0zTPGdVONdHm3QMq2HXWRK0ZX2yAUJYPJm/JCyfcTGvjXCRFlaAtTZw
+OFMAq+cgpRA8RkU3TtJpgFSNpf1Up/QDOUegFpLXBf6+n+RNJcXAHlKHW05j+mC4UeWP170AJMU
oRF8FDyAzzJOmVvKqOyhH009galGuxNPUwBBJZrtYyCXMpGEC4kd/IkGDUJOKoyP27CGhN3aNVz0
TVj+ys2JM8a/HyCSiLc84jbrtYDDBpKbVE+cLwCtutmqzt0iNqUqzbS5gUTzYcsTJLWheTnafY+t
UQsttwxMLdPTuGeee2UtOnRt1G9DSIWIQlj9H2GipId2XLoA21j6fzqQ4V+VztzOcctUhfWcYVjx
c0B/C9qjPxu9lgVAOiSOg+3wU3sV3TEQVf2g9BohiPie/kulJ/xsOLVBuE52eWVkvZe3iwBg/ESc
xjrCwSz/+a3vlBbZQP3NknLdqL67b0qbwJTF8LW6efIypID6LQv0Ol2o3dvdCx8wOb5ZPtJV/U/l
EuP+fiTEz8WOuKURgT8cMqjF1nheHbLb7eHhVOvCNy9wAhlN+IL3ldBl2xdsKi23P6xP5Qp8hkNo
vxOsKJ162qiKwpyemCG0JMHWeDbBa8RQainUv3nf5E5eVpO3ah0MWirtunnY8kB7IKOeOe5GYoWS
DWsg7G7z4vlhh9+nKKhp9VPlUtFamvDRGkWpP5vVsZ6AF4KCfzUwz3fcT/OOPVf20sbyBLVMFmlP
txBIVqVrYkpHo7BcxoV9s2x6kMw5x/0ziMwu6GXMS8bjvCcvTK88EONx1muDM3k/V9192chaxxyP
TPtxO3KBt5DfScExW0BMdtuTrQu38TWZUuEk2hP0AfXkZ9xaKRJrahFGrJIlwGMWvnEKTCOjhq4V
RoQL8vQ3iCuFO6iPQ7RF3pC5I4htywrWTrWXjVVQUNWGHdjA5dbKzqe7r8+3GbGivvEoxmG8tHiX
bJJ7rfOHLYaC6fDoMfuTAu7g1B7lTDwVdQDcyj8KSsWp0+Rtzgyl6b4POlcEJ16QQmYamHt03xrk
qU9m9isqxgUHqoLeLpgwE4PIx6d+A08f8NSpWWC4CuLUk9xZS1GcLoSoOcHSzXPQ0/G/Ayneyjyx
Opft/yyL581PbrnP57o9lsL0mO/CEDsbyG1orZD8lWTrZt0dMSoDDGUi79lHj4QM6bfCCskTW7pZ
4p0dLydkJYRGtNHiY18bxObtkaivt+0w+So23qVt3Bb94panFUXEGiQVX9GErFCOoWEqEtcZ2bG5
LLo9tRWf9XLnlHeViu8YSEq1ysSdE0vUBTJsopOkbsAUDmAhc/lDLqVyOWdA8DK7BihNf2gePnWY
kOVceTQkJ8wCfLRN6Ds7L1EL9RraXrUpTtt6cmU6SmUHPFRLgcwOWawpIXLZpCrJhtLcOTk/om8b
DMf1Ls7XFnYFqXi+JmMRiJzIRLvxOeqgVqn1lkme22nYftBk9V7WAJ672L90cj8KkoNbQ/LMwQzw
dKs8Jw7DewSoYsx4jC/ayPYU3NbpI1P2WQT0aZ7FK0/ElaFZXDwCVS9hghG4ezjOEcOmyGGK9l4d
qvTcgYNc31KpVbyfkDV2Qp0gmlSWCle3w/iTXO/m7vbqs3kNfL9OkGL96Z5mysjtuev1PihREzgg
R3ArE9tB+XshhS2r8vIoGOfyKcVNQahXsLSV2HI4PMl+Cn4TGQDPbyoCvvG67xs1FuGQ4GDKpIQR
oddYVxp4BoSV0hQQehIsSplNAI8BOYfRN8BQ5xNdypMUhgV7UJvSUxzhSb1HkdOdsOrW0A78kCmO
Ra0mCvpo8aOpcoG0vvCHWOcESRAyE8K34CeBXXFQ7d6EGM9Qi/0HTrnxW55zXij/trUBmPezDeC9
4nB5w9LjMrW+trJNWRLeY+DHR6dbHhgESVNyO1admDJFmEZ+F58jVslCSavt0JZpz5xDqn29yiRL
Et0UHOLSt1wA4XjBp6ba0/rOc8F1BU3v9YF+46JLLpsYdxYo5dJymfVOzIqOhxLlpEr9y6ZCq5Gc
DmUNmQi34yN3SKceIszDiyM2Utlel2Pg30j7fi+nMs5F3VsIQom9hmJYuCOHUHIHeH1uNJYx8QXT
xV5Xb8kAb/7ewE37Xn9+9m9+gm3ACRGLY4TUrys0eXhfE2E7wLOOk8OEQmMx/fnMRXfJBMGFmP9C
tnfM+wJ9pOt1uUe27GItagkv2gSHNSedq1MtzEKAJye1d5O6H7mxTteTPEQRxpf+qeu8iUSz7u7S
JCaIwQhUrwtFhqBi4ZFZ362s+CQgEaTZ8V0j5nOypI+JfM3Tz6qUgH0IxBcaw9haqbwo0rfYvOie
1DlniHLumYGec6uy3D+2vQM6lKq1QjGnQkLUjjPjEjpXttBpcm31NBdIuNk07bj1wNcli5P16Q/3
RTufLv4A3G9tgApQTEDzF7LkDvHxBk3oISFVhYQTIDMRV7lX+m1pkw1Vkul9qyRz91w65z23KOxa
8iET57ozveK0OPgK/sYEaczgDF8IYJFPXWkRTUm9kn/vGqFQe8pU216JUMtGhrSts8JxGWALQRyO
w3JlGImXS1Rrj5hdUOLcC/6N7o/UKitZpejStikMbEfdWrA10p5AqkvbLvk0B+NItpIDrfbwran7
bJ9kSu4y3iHmO4pjkNclj5oFbTFnu3D5On6/Wi0Ag5reR8rsrYmXQdailefE1gRYcUiOWeiFg9fa
mlFCEa+33nlNMPftLtNDdACAhZQlU66ar5mgzMK+ivyooqkQR4XoaRVaq9E5exY7387cBlBn0mBW
Ew+zBKi9lwztbauUZuC7GNXuQu7vsNtVkiZxoRTLTMvmOpw3Lq7Akl4Ah17gsIy2sfcAG0FAadeN
o/SF2+axLS1JMsYk798G5JNiBSSvoGHZJIdu+iudxBJRLFBBt5LXBE3HMlYQmh/q+ciR/0uTnJOB
0mz3+1fzeut7AAGMyWCqHErRhKOQXj7u+skOUiPTk0BJXn1NsDK7WzMUmJrqXyAGiE1S25oZl458
aJRa7qF3MohV6/ViiP1WgH9VDZAN7H83YQfmwwV8MujRBWbj6xUpI5zjMRMD8OH7TnDB7AaZuHNK
aJ9Ld/nli/v2BzXbMqnNxS46MMCnJObjFyL/sAU5ds8Ql5bKpd3tEpHDMEKG1UmM8WDI7yJDFNc9
V5VP/d5IHPYNDfFQ2+e9sRJofbLRfTfmF/wH5p3OP9LvBdiK9vufXbP7D8/n7nf/k1L5Z3YORzvO
9NkT1xBnjXF1uoo1WW+02ZMsy2Inxq3DG3sIXhBW5BrQaNyyh2QEXW9Pm3iVLE7YvYiWudfAmGMV
mOrcYoEfzVEHnikeuEYGH89iKtgv2HMkm9i3Pn41HGkcuU9CtZkHFJPkmPrA+3xhUnaDx/qGVesj
ZmoEbY7nSCSaJQRADAf9HJTyCFknGnf4HAu0/B7Nv7n8X4BO91mMOX34PWK+98iYJ1S8ea9pY2sk
Zx3t/zOwamF170cLlITSktSQHerwVe9ic9TMAoQejtXTygS3c22VKMivoH+g4NhA4rz7X8ZMqo2/
60IiBPWENthhuaM8WZ7ZIRlUYp/Fmo9eTaRgdsHPraPnvR8vqr91OWG5tPFSxpckZs3eOZdTwSrk
Did8Sfe2yt9mNrFrlaZ/+LyoeIrg1MMxKdsJRKdJxHM9woOnXkdOyDB/tR16mKf39vp5kGwNZLUu
Y5N8GMCdY2ROPJHnABK+EPtCN+AE2+mtotZWpiG7zMYws3aEaNbjofYGFTtB34Yvk5uyZilEZVNg
HrTAdA695Ai34cvyCOQwRFkAmYa+FRWi+b2xHtD6Su1IZg22yyb2jkkESDklqRf0N71eHetXBgGt
bOzlorWPyxicXYUNbrWDm7RUdhA2cKWcQ40z7bSJTSUIDTiZYvDlJ9dwxx8p3MY/mQYvVt/2Bd9H
6qytv8a7Q+LbMwQi5mphjzCkCRcUeCg9mkS8YQ3YZdOB42SO5Gxkw9dP0ofXK0BqYbYiSBxl1XLI
EPB5gqnv3EFxeuKKAz7yayXzyL7mOHA/g94Us7FWpSVSMLwXkfC1IjJmlm29x++NoquYaTld/8sc
SKaajEzQe+iuOUjonS+in6fZ008/5J7vrTQwBTFvZczl/plK+JEBi7m/KG4CSUd8Gba1pEq8gmT1
VQBhrRu480PQM9yi6Z2WPKNsCTo82hoqdwjVMXPlQqPbIhsFVj6/I0PYW3ZlcLXyV73dhu5/ciFJ
xMgcxGRpLG3FosyaealAdH9UYed6Qe8nvDg2K5bfUYHzXJtuGeHDj6FbcjEb8c2JTMu36hqjIxyq
IZ/7elA64AU1jPVAP1i/K1ZosUwjt7dFh/pdHTOefglTynQaqCeq29QB/BupQYYsOL6uFg+oAFVu
c8EvlyjGIIR17efqDS/caXLfKTxvSQd9C7GsaVWRySzHdBUZ6AckR+4YYeb7IgynO/XKcWywLOXL
ITht996N4dAX8WF9s0Tl3YzDKj0oDAOtgC6hDC8RhlTSvoEOn2+fdSDnewSwWbyL4ZhrPkCmvh0u
Z//EFe773T1+iGMMrlGOEc23qYhYP7Rx8Yet5M7+Q0e/WXHxemgvlhX8UwksxgV23BgDrKpO0Krp
3pKfMd3nsirP5C/IW008Ez4KoxMwfgb+NAVtfdqMpNQXzA72/iUuqNJb8Y68gU6Ky17/lKQJK8+t
sJ8t/tZQ6wtYHyg58fYql1CEBg3W8yyr40NJ+RSdbkTC6vsxyMbvBKsFEXDWbB4Kt8U5shy9rZjr
JpipquKdyleDCTRpRhY89ofAVz2e7FnZnnEz2ZEMv44TNkXZMR0tvLHxafLoZ0WkqEaq9bfQ14fL
q3rLqWAhGzQuprNK2RG8+8aZyOn0AnxYOs2GJWgYL9JBd+VJbhw2B49CGJJUuXF4IaJ6S5cdfK6P
ZNvTHft0lKxqvoR9YSejgzua+Fpj9P2FpEAY2B1lT5/QZWipc3uFfsglGfgbKO/GfDbP+T2ZH9pP
O+q0FdjJHtDZbn2s1YFNHQDvOS2RhPVYnDGChZYLeYm7S926YL2wloTOc28rV2FDLQhkmAjYCL3x
DjGiqWFC/F87D1ZqTMr/QDpdIVkH4UzIh6X76I00+pKhPNVDYY0nOKuM0Gb2DsvKSGgx6s9Hyqum
JMPBGMGWWs6p6XGIbvJ/lTlZcar0s5lJP9DJLkwZQwSsVjwkXsaN8v7MSiHeNlU6KN3+hyRThiFf
0I/DkNeotlRIpb35SWLb4b+iNsJmcgo/sETIazoZ/NLBntsgq1XsxVvDTtYxgz5BEEV8m2OXxzTk
hQZn3Sx4R8l13jBZXLEFLLerv/pQhEl4OCAcztoOlcjzCsSql1JvA8pUPFfatHIsnagJTM5v3Vpq
laJfTcqP1pYY7nk9/Eq5ETXS9sTDzsIGvZxEKW5WKZc4FpKXeukNrywqP1192hVbaa8Os7b7l5MY
PWu5IcVnLJ8vepD1neV2EBlIh/CwC6vkffyUuZz9ae6taChikc9nT52isqvRUhMvDD8litTrYzOl
mIIQ/ZTEDM8KdB1EKFdie5zO/AowcUuVuUb9j9wO/Q+KQjTBdl8ORlJ1FftN+t3Ec8fvgii7aJwX
Thk9eqTiIFnQSCFWmpuO4yaqRdyeK+Ubwhw8MpQbOVFnlHmg8pCxPHcvX2uawm271Xm//lCyMkL2
SIv5e+ghUQUoWWSrLoHHHPHi8nEmqHTry/Q7dJKSXWhb2k/KqlXGBA4pG+IZ4dKDrBKb+Bkbx1+q
wP0ly07A0u9xQARPiKw3R0AaqVWvZ6OfNQ0SOyPqFURxJCUgvURGyy6HJ4JC92ApHmhV40toCOkj
GWdQD+3lA170uCc0q6HbYbIA2OL3Sxlr4oW0IFhM5xFNC+Kkhn2mYXF0sYAkjszJQiegk+oZ/QSH
ntFyfHcN6KYqvmF/1kGaewK12ab2/0/+Kn88eOoAxsxMLznYG3gGGKRDe6bktb3Mpuc5YOwq4JwT
qs45jvAE5V4h+RHZ5Ke7lkn2JUX6hsVY21+Ie9lO6TJklS0iZSDL6f/sj1aLeDS2G/J190bf3U/g
k40mxm8/tAvZU8bKFeGkbcRtc6sL8HsxbX31SfBe5iRYyE9M3TFuRN2oEzG9oEchWqtxFUeh0EFB
JR8zeknAQqOTbl/AzBSxP8q2Xamm7zbD3XR8Xa7gHiQvS9vAuDoBInHi4URBndl8PPDwtQ4+ezFv
kKI2gm+NeMxt2DmNdxk10MeUZxiqLNZjXz1E1JwjpRIsSXZbn2QiMVEMknSkuKXtBkfr0+rL28Lb
jGf0+Ph8X7siHOngLDD3kV0uuFzrH/OTTQsFeVu2Usai5fQXDgSOeww9/YVHuqQCz1EFx/UyNTT3
cPiejNk7HzsJMFyV+yEf/v21PVsqrQoICVUxcyfo1+80675Y4oKvEaCz1OtiOojA4x83EQnoy0ut
ez6/Sdi7jqiPnz98ceBfS3EBGjXjhDassj7eZqAmP+bX57nP8xJ35G+FVOFqjeO0BfmuqnOCEpP5
JTawdkPN9f1vg2QJiI97U3Ia8v7XS8hbtwjKfnWH08uMq5wFJuUFfJv7XMLVkarFdd/K7m55c7UR
pPArr4/HVay5CIIysRnWuAWnk7kM/3QlELgJ2mImH64UOUy3rspDLS3CpqPlu1pFlHHT8mdwKIin
WhYAkKFU7HbB61TmdG5rL3JWEMmZyux0k8IGj8PVwlVRYAs9QZhufKd10gyquYktSWW/ZsOlNJll
j5bq6gljXRN7dOAxjFFknsISRNBxYgtiaOmsI4gVJC3bvvIyrKMM6nsSAVWFeuFzATfwIar70Jiy
o0kMizPZ9At5jkm/Zs68Jiw7/K6omwx43qcHaqEW/ifqThcQW5nc3Ts2ag+cOQrP/Nqtns5YDWM/
t13JrkNLgAL6sKoOcJ24sXJyVMxXftyGVgyd53S7FW4sMsuBL3Hqv5xG0brpQodCCc2cmXE9yued
qiFHFVReATB02YzFUgbY/zrH72y0NaYIhA54OHbPLjeKXQ+pKNte690SQrARnoM880PfHmv3HhrX
cDu6m757mrv+aw0X2fghtC1ehanQk5wUzISwxeWziPp2Wihb5ppI7CMKY/hdBs7mckDXK3kc3+eT
wmLj6Z2MT0jcuGGD7b658EE+1ZY6gvd59He7KPC5vGut+AYsTZf72I6Y50SHKcv5Ev7xZqBpUXMC
Z5bEXYjKcWLAJtbVIBy6Doq6G8yqmwi2I4tu9vYcnbsdzL+KJYs4XUFSNvbMS024p+znhAImKNk3
oag/p7UIpN8RlDCLrthSREDDo5EalqXTzfASc3vsLWh3sFpYxDGulJef2vedPkeqapH1Mp5iLH15
dlD45iORKL8WXIx7zcH0FforfbfmscUQrj24C12oGNkU+74BLqsBwCbv3uCRZSzsSWAs1j6OpvRb
wP+9+dvywAi9mwXmHrnvqM9s+EkXyVahn12xc61bPvo716I796iXZhOOpZXKBGc/tKbxgMDR2jar
Ukyk0ZkqI0uQ86NaLIBpy4ULcn72ChTcuXoZsUljXkY3JX97X86Ns5F9CvwofA4MmXL4BwkdQltx
HuQxiXdKjFnrEt+xXS9ZrdF7T596ON/sqs7AWiMGNgE5cYn/3WKY4/YrPhIeB6o0TizIIKT3uZlV
MzUs3f9Pp7gfIgeMJ9FF9tnoY9+FpHA4w95CLXzP8K7LMDZtTLs3Ie64lSfeMR24l3KsmjrkeRyX
V2yARhHzBaBmk7/c8V0vgVUsb8KWl8RicYxKhd5+WSQH/esa/0QbknqYiiPCqk305egWBYt47mIn
aO+QhafXUPZ9JmkCbNRVBeg9d28NuRmZRPkMk2u7Pu2RFh89tBrPQaGQkN9pbJq7hbmhsDPOH+1C
0uBFf5jgYnSEuenjQBChHgp7LzfP4sqn5Mn23C/WFatwfNEi+YUOTMDheTjB7WATuaDWB3YAqTSa
gKJaRmgmSASKkOBT+LOxf5BRYcUH8vKZxEtK7fZxAjC8R53in3Wn9IhaopufyNGlNyqXqKFR7OXL
sCKpDW/YPrNc7caiIMgzns2tuXN57wi1r4fvH31Rgcq3NZ2DMriD4B5x3T0lAPezYvAK8gAeZZ2q
FXxlfaXpKRQjVcBg2ZG+WLGnOa4zyUaM5Psnzk2ljpomFVEyneac8PF5eZ3Qi7mRKqlPXnmazXEL
zcD6NzhZi943DkqqXrgMWPKc08uDlxA5Sba5opjUGaIoyA4jq0iChp7JQ9aJIfycF3KW3SSepFc1
0S8RxOaKqd4NMW86ELcS/g0v4uMCJUDcKoNcIQl0L5+AzZy1vGqqgVF5HPdR+qNxVZHRLKNIhXT4
aysF1s9tw3HPfqJL91VxSUo2aPCDjHIbcKUfn9YC/4846MD0s1QZyquu6KWdcT3OQK53tyAPERGd
c8GilQm6HLCnB+2+i1DGw7KtGsnLytpC653RjNqSNFd+6xYQAmyQFV5Q17DBaQmR84zpEGjbt3HX
vdjmjFrlXNsidulAWXhO2xJbS4Y/vOWqOH1Xpzx8M/MAv0VxEZ36Xnk6JmTzVv5qsEchf1D9ftV0
KdDjmnJZ4p/LeEMo2+pj0irAa4uCUeTJ2M9FCrdGBEyb+bgeesaQoYFiA8738YZRs1GCC5y8aPvD
NJKYuiG5iSz7UCwtPUbNu3xFLvQFprUsjUBgI6gXJt6PdZ132nQfYf4JcNfQNgmVkCCv0FrPp85F
veeTPP3HwbElU6QxQVHrFyRPFvir0BOJe7XgxLQvEuRPlsOMgv7DfMEPBfoyKVLT8BjEEtEs8sM8
TCoKgRQtuPiC4/RMlnb6IA21FOnan/zaTeOHN9T9hlshbRikkhr1p6lzQcNDKPxnneCzpADGJBqb
8X8U7h608gCZAv6KobScpa71Nd57r1ZSfo/hAHHUOIxj9vhjl4Qk44iy0zBHKo6hz//dB+euo8o+
u2oZ7HAxS5LERUn5m5UnoUdKpxaANiA4KwFLDeNfMv0PvwZkbHXRy1I4QmNp3ooeGaahecKqFBUD
pRbRQxA7TbLl/NlWKt84AsU+pDRvKBT9vOEw6ZdP+2MUoixgU8EylLiSabRxkX8mqYIaxsnkYWHL
v316ykz+QqGzHfhPOuWuwBK9Lr6HRGxnnIcMj51DPzOucoWlgM2nfwaIpaVl1niwl7i9+akWbaU4
SRMry9bbV+xMV3Z04/Tp4G5XL3KDSO1F0DMwhvjjC5PQH/OnhZmIN4VssUUi5f8DMIBRDsy898fg
rgxmS6lzUVEH4w7QiuQEHNuPz+sNxW6++s84FQDhQyIbXlf/RfmaMZEDnZHstc0qMbhbpExgtSqT
aPq+GbyRuilN8vbc1UJ+QqkzlHpa8H+ui9Yz9spMxz74kWTZKRs8ZBGdR4kP7pv8Ud8E9dP6MSH0
VC6GYtpKlxT1V2CnR9DJJuiZOgGlxe03sDjrEtmya6yg8PIhuQcIOKgCTgwjHw1H0UeI6cWFt5/i
sEMvHV85I6FV6vUa5/FKW3JBECLxjy/kh0wbgfRdmENk1pxoMp0XWM97k/E1xfwwf0Xd5zizNLkH
8JTnBTGcYzAnA8Y7HMla9+xGb1os/Nr1cgyLVkg4UuihTuEC+Zkh+YTPNSPrP4E5FgPpL77TNE02
mHfY9vj6GVRq6P93lPY38ZMOGlw1XNW6X/V0EPdVomW7sLHCnTOTXg0agA4n79wnITTcbv8wxEoY
g730oq3FIddC/4vI27cgQDVgv/SwifpfXdsjUh4QIG3aHk7v+4aJM+P+A5ayXfK/zQB0cS+GqEIk
YmLslTMc3/+QmSX5lnnW9IcWUVF+6i3wzzyHbE268/O3Pz0zC9bYEQThpC3jjwF2+D9g+QjpHADq
rZcXyAAlMu7FGgxUyf7V6agtnNFgi6giPTi5dWrdySH+AapH8GPz/Uh7WdGMmFjs1bmL16ClIzB4
cOOGm9RaCtX4dV7rHbEoVAuBIImOsX8PT2FqDEPYZOLIDZNjwGYfVwrsZsjhnst6e8VI2b3zMYG5
HwLrU8yd2xl2xHkTC6rB0Wtz27yHBJelg2wBrhx8QPBsQsbwA0i/z/aF8mwLuTXDTLgAF63kINbL
rR1ZiK+C4Oc+4WYwioCKDdJyqNQ59DmlKyo5Ojlaq5EoTxRw+7ow8YbKE3eTgxwF6pO9QrWYO4zy
tuffQ2UoB9vstZJQj7+6vjuwxql1RdCfWJL0FHBLtMZ0U8hHGYFGCVH1N2m11WC1hQSh9qIhTNGi
cTcYPzH20xUC1KOXkgEr4slaEVbsG+rl2KMp4kEvDUetMJsprDriZ07U4kKvp/f+Yz+LRgOgRk+F
QRHYaYjjc1pHNwkGzWoBi4lnVkH0WNkWEh8xWrglua6/7aIiFYqezM6tLnE6/Jpp/xFUIuHbCelm
AaXPyAkYlRTthNGKFW0pLK4+GVJ/fqMI80dN/Kf5VduZyZ/rohQBv0lQcqPFCm9Q1psNv2gNBxE9
S1bO+UUoqDaNVQ/vDv3gn2EQ5EP/cPQ9iFt8V+lhsFyyiJj7oGWBO7YTrG1SAYuhh4/chnpIyWbU
GvvaCqdK71jP7Jg1jMy5QlanPm3/lb243dD2yvEUp5TW6nYUaevehZPY/fVYXhvI6xVpKkCpaBKr
gYOkYDsVCbNsN+RFEzWJZgH4PKguV8fFj9NuBqm/maAvNyceCiM3bzx+VQvQkhCikcqQHoA1/8Z0
LMZhv5TKHs/R4ViuafiNne5iWbfYvZsLv0+4JINW4dlnCgpP+QD1wbf57q8hex2QUMDoMTNb9wVH
y9OrhznwMKhso93YNrC7SaAWUJ6155e/iG4chuSNM6WR7dW3a0hgUU7sHQhAIrTG1yc6/rynsAuz
MP+9gzFzyjig5dP9nkXZ6DDMIg2pKbWufnNkSJp65NEWqgZ112IIOGbvpXjx9V86BcmpD5gW6gBs
z9BugnSjTo4+w1YFeq5aGwczUqx8YDQYNjUbElAO+2xas67Ba97TqPYC+WTcXVToMBpJemFTD6z7
I29S+lzd6RipPlYu419aJUMFXrfHmZZiNFL55g2L/MxKyZ59DXOifqheMqZvLA1KSDoA5PQQSAvX
Ahu69WT3NPH9J1J5YSNRk5jk6wPiJiKmyQBpOkHg/CK3kS5gpUOHWcXZZsCyrWouHnFluD3+e20n
TX1/omXyutQNqrRxoCuaFi7AZ2Zb6Y1GMJ656P0rk+ybNIzUQUI2gmj0aj8GfZ2/U2vov7HKDKpc
LeyyIPyKpB5cEYicI+BEkHIPNqnlOeFvH9drg6W7ykEUVXxwp0KwdPkYZf4ym0gVbtfgl6wmTTiz
QdPq7/EuRmJATotFL86Ah/Frbf+NRuEvwh58R3vlpAlrVnqooeAcJ85xrU19u/j49Row/UuZOMj6
1HEBy3bAXQleiQL0RX2A1P2IxYVeVAGRb/3rVsSYIw4NdvCOdhLycPqdTMzTDSW+iZcBwIBFu5v5
7ZvXTJ9kxHmSIFZOH+/jlcFdG38+VEr3zM6cqPO2VYxluIpphxRB80PCrJL6gqnatMoAiFzRRfBE
QPX1GNuvmuH8zDCJc7GIV9fikePD9z/qkzARwbDsqcD/9nOI3JNrqJKH0Va7gyiSearPVDOQlUHX
n8OG2mrCRAhkisSIKALogJiygXYApGZqGw4UHJBA0H9Ei1xzY2Bckz3ntrDZDWP3VIp90Ge4leSS
Y4Ddm8YoU24se0XcYjUjXqpQER/nyMi8lAIxqGqRqV7S3x/hxZqMlxgaELabIZbO2gyMnlyrZ04t
UNLdqR3w7MsF0B9FDW1Mj6apVFDH7B6MEtFxTRHF2vzhO6AD+ZO2O2HItoF0AuFGRLOV24inYlnc
C5azyFSLe1iys31ErEjksn6cJQP5NcEqy6ZYkVfdciAFCCSzw4Kw7fMEHGFk24oXHSZ1/Qfcju6l
HGCoXVUxCFRknHKEr+cVfgA3y2ttAzxyFKwVYoyZRHuYo3cE3D9m9RST/YSH7b7jugBD6DSYtOFd
R2R7rBD9BHqaPV7/QqfpbGhk9/qSlc/33/xFshehQ9VYI3eOPqik9MrmXkam+HuZupRBsavH7xkD
ke+UZ8P+SMJDDDZPhdpZCitvDtMDavfocn+2brVvFTf4Yy5EgJPeDFRavM4aKSyg3CmvfnHJL4H6
lspp9n62HOGGM4LaOlECt+iDAoco90QmWYVAoLobeb4O60qXhppr8rnZiGoeNchB8DHaIlZ1gk2Q
4nySOWVoUCCMaoJ62kt80BTrxeRMT74qOFPM+bNLkn4B9/APWP78F657rX1s3K8d3G6PlZRLXdIz
m4y4p+u728CpgpKYY1ddQ+UPcy4mIcNGZQETgabpJt6jJkait2ASwjlysH/gxlw92T8otXot72Nt
qtWsPLs6skZNFMFQ6bIjIf8t8iJfx8o+xtH2T71av9qDBJKS4l8Y3CI+CzTOt+ljS0HARGhZkhlQ
k4IBKIX2Smzrlicz18juxaPTaBRbMj0Cjvkg7VaRa/RDweifLhCamBRAttiBkONbZm4Ef9APtm1a
Y702zJ5H2viFbocix8v6WOxdXllg9qRGsgLFlAN9qyujWmhQFF/FBE039VIuH7BtcJ98fLrpqnsP
E7AGc5zM1Z2YNM/9l9zMzDtsyTqwXCEdZwn5u809kV3p/PCbs+qmve8hOIOBg7shyXyTGXgirith
C3YgCLgX+eLWev9rgatUvES4Tlk5Bim3cJTteDZ+T2kSK2oxcU64VJ50S01kyLpHhL1dCHGEpLRr
lzem1f/xYh3orbUA0wbIfeywxt6ezIHXenciw//MZ0tOsevQYncG7n1lFut7BEhrKhJNrSTyR3mW
UcOWT+osWBwJQWSPUB+wp2B6rRugJOSDLHMvP1cf83AdCtVAFceaXgK+hgOAkIo5ZWja3jiMwHol
mAj7sobqoz+/SLN66fL4FyZnYdqNY8tpUZrGT0BK3L55W8urCZbLh3yfU6n5LeC/+635xPIY5cvn
P5HvBlh/N6buaAUqnMJrPRKcPN0+jQWq55o8KYq2TU5D1ODQkERMEMQYVbQexTmYQtoS9pdFxcnN
P63+fzucJfPQvlPoO5KocAwFVgyTH/pMXL9Bbz+VKFRYqChoB+76y5LTlzRv70aiZOyckH0tdG++
zD4in3IUzE+JKaqDCH9NytydMIzQ+gkvZOFMkAQsRl/JT6oIfrfkGcAx9dqZPIxGC8U3q4Rp+Cd2
3X+COka1X/QYPcgANgefzeciMGFK3PKTxeokYptVWLUB3p3l0oIjMp8gB6CorXZcAYwXgYI2FgWO
gu2yPdi5aJMee1AZ5sGvwbHOlYbr2kxJ63zT/3jS1FaXhVu4ZE4eck/S2Q+D6r5fIKt7kA6iZ4wX
dYSPa2AJwtRa+aonq8u7lxOVpN2LjcMw27PmbGFKWpig6ZBvgF0jekBhQMPGK5hb6HFIiDCULU9F
ITf1xWbSCmhh4Qu0XVJHhVwhLw45G7+LPsoEMpUdpTsD0SFkev31CbUv6nykVhcs1F/sPbBglcRH
t31yPQ9cP6poz18ZF2PkZS9Mn8UnSkjEnXVp0QPmhKvJH/DV05eERTfZsjFXyycof9jW2bKZ6BbW
dke6rtcz/+bw4mB7LQyJ/+53qtUBGVZ3qm9Z4qjUmtlirA9P5br5drakIG8lHQ3QA63eBwO2W2C8
er8FbA2sEcquozBXA2Svgux2AHZxHPsCODVkMUe+kd7CAtXq/0/wd5B+5YM5XiQWgsPSKU74BzRe
AKi9O8b17YAXus3xdspW7QCZrxMli7nlwzYvbT/cZwutLOZqOt7+dB12IwTtlOstIAUwjDxDiiIA
vnQ0YJVV4uWsZaul8lW8gUqZRdNKKJyhtKdSyba70XT/EGwz8TcqQ3Aa4iknzMLumTKmusLEKXpg
hEXLKTQdwowKMiZxYAGsKVELVMD2j1v/EK669O02R9GO0tNgXRkqo/OvyhmrPxEoBnrINEViGguE
wnoRlaKXL6WOP0Se2d0vUCd8BeDcM02Cj9wLE4zYpVplWQwlXxe1ajqD0+5ikqiurx7o3i/ZZkko
diuKvKtiDDRSiw9pKyMW5Qv6GZ7ojNtlU2al0OF7rkXB5qRohn82xN5UiGAmRPcP3rjZxEkh/PFc
HrnsihQhALgRdEyAiKrCQd/4kQgxKBnJM/2DvwypGS/zLO3VxvadueymYuaZrWqrK8SUTSJbo4Tg
d6hWopAsiVsOTp+zUG0xZSA6PUS/QCT6uN7Yb96i0epUIk1+gFF2+ae+DPw0YpsRBostzNcDVCR5
4cfhUfQ8OKlBW3bJwVOGgbewm6SJ4i1hwAIMLGd5d8Dz5XbkkNja/v14Moa8CLAkDWJgzn+RLNhh
0ssO1Ip9HFJ8E0R2Flo3gTHN3mJXwyXgnfbZpYPteMRsGVvNqS3+7HJ2L+XmXGk7igZ4ADvswjgn
kwghv9mqOHRDNqEFjDz9Jlzj6ufk9NPQNQdcHONczjFMEoVQ3FMVtAttgKlFRGbINZUFhMgYQ6sA
2sr0jVsrz+P98kJfWO+eazkz7iq1VYqDLsX105yoQjsEUFm6lLRaJRNmSDU+ShErMblstwgBQkd5
z4zZsElYuIoDzNZskbrb49uGwERY2cnbsq3TBUvVyzRi0ma0ueZUkUTJjvhLp/y4rYK9HS0hAA8Y
ftW3pXvmFdzIE5iCkYB87GVfo2lVPtpUZb+CYPQ5hTa6b3HfgTHsKi3D+6cgBFk+meeS0AqKKh30
2S4rlk+tGe/97pwpOkcwFHKOUYTHHR6lOlbptKgN99IWyC8vJEyGi6iQVUWHKo4Gi310vRen/isQ
X5BNd7afs38gFeQ+7iLg72uv998TfK4ktUZItWz/TqKgTDdTjwNNXJeaXXBFRpmuJ/wdzL9ihJvP
wFAGpBed9SRq30VkbJdpVRPtFpJFZnJnYI/YXUoCbfYc5ZmlSO4IbFn07JRai2oiedYcff0RVUGn
U5QhchKSRbP5Y93ervjvm7rRA8dPuHKo7uKl+xXTtds0eww3I8ydBMN/Vi6+oRv0jbLHT6Cj57p7
P4thUUihRJBR1JgOKmHtie0Jon1vVOoqQDfMKcqa5DFC5OEJd+ECGN54R/uYz5dApTw76tSQEI3E
yTSjMYqiXtZ7i+bc4XXwYoAEK4QKgS+uRnVeGhYwEhSsB0DoPa5uTxdI5JRrSpIHGmgnnmFC21xa
a2on9aNW94vEp0ej3p0zjFS65S7yoeOJEpWPx6KZGe+dxIszVr/7SECNB+m3UvUIrt52E8LpBZz3
bzRsgBsKm6g0lHWGWcrwjufbHhotR9FnKNFsU2CWQpyUP4S1Yz6zMiRbBdTsF2FoAgVx4MtCWELx
kg6ZN12sPvSygPJ16yvjbYYpmSR0dhQYyk3DBIcjK8FoLqh8w/JDVWG9o2PQqknHmaAxhFzbOXG2
QrNgjZ3vtmrMNyEymfD8AX+2icNfHv5S083k6a7uthP1DiHtt1yC8Om8pt0wDKU3eavHYSspfH6u
SGlvN6Ns6ybZuzLVGevc90Wo0gBhQesD08vKN7J2rDspFH17qin47dMrk9NC3Jngj/vgLuNuPQyp
ygEcC5v+vcso7o+5kjeQuswSkeVyGK8U1jY6MNaZkR2yh94/pOLEuOin0YP0S5rnScLBo4zPIoAG
zEvrefWiT2FvhaJjIo0T/KMA0PH++f2a3R5xEJV4usPB7NfzC8/mlIQkd27tCEoEdjc2m4vrkB+F
lFoqA/vs6m42YZ7TO4AACwNZINUtE94Ndqr0nncSrua9osm8u2J4MzKUIhmoAFQSfmECIid9aEu9
jxtNuao03+Fo3looiu8KSNekoDS3xuqpcszESDF8A/jWaE5qL8/lXsPMLeY/OOkU3Ppx9SVEH7tm
W8/lMfTdkYn7+QWQ717m/rCF9JLaXhwsM4Ti4EiuDTwXGn+ALhoI76CIi9lG/kidfD3k4BS1nqGW
WMGLegG3YquOv2YOpC25EAjXvcNhe5+ic+ETBfmdGAKoGVp43xucCLVvnHC//QnjoQObW4BuQkdj
Hyg44zCRE9qWwqIbgfsIK3v3C04B01WQ4c6rJ6QNPqSJ5WALzjp7ZI+AoaRuN1zSBMvUxKTKjE9f
6dccw0ZUnEL4PL/zWgzZJjQrAeN9n2wNb9p0ROzP5uGxxqoORzhOzAsKnc/b0TFPOWSevzl/Gp1y
/02BHZ0LIWCG9IGsyWc+y0DDXmHPtnsCZwv7LeD5tGAWiy17NGNAwOOUfWFdyJL3hSnKmaQTSpYp
e5lueqh8K18CpkFo3PQP1yBb2S6vj03DBE0xunAzlI1oZktHmQDK2nLEspd6mx8O+IQXc8sTV0ys
Bvz9s83v8RxK0Slgh9lh9hJf9gZF+rRNpbBotenmPAxK5XQVOJ+AKRlDdTJTMAG1GFcsXzpbcwH+
DqBni06cVAcizwJxE/a8EfOuqhIE2aMQftIxfyBs4LOMQQ0bx8a2gV/eyFxOeLk7xIs06xtq3nHa
bfGWBQziIB0vKBycpeuFjg7xJna1mYO1JGGV01l60tYfu92IDlhFhnWGzVRv39t3N5KtPB/aXD1d
cYOGGw+KqQjTUHAfM8S/gGs/6jIcbI0eq0pnA2csbBSrxRM6uQlYHDIUepzBV5u4HT11EhPZn+JA
fsDWCW4/5frMZBefEoHDpVIlXIqIXN22ksyTLI6iqDruwvtTvpYUe5prMHgP65forC6BiqibZEHn
IQnna7oTmj8nomEf7JwglR7gFJ3cJOd3fF7mhKQonUcrsLuDwprN9WtUHGOY1y8uQTfNSuymhlvp
mcPymDqedishcU0fuVRhXJW9PRQCQzsaH9SAT/ApIeSCFa2kD9SqMwfbocf2oStfwAMjyHvqq1fH
vP3nVwUDQDj4DA+9u9YHEPd3XVKm5dH/hqolljbm9VsmSQzkCJWDL6WJ7IyyjCgiKD18v3bsFgsV
2duL5ySRaM4ioQKBsJ0uC8fx89crPKCCX+iSTrqS0fEPQZuqNu7gSBwZJo3DAfZOs8dwUVoVmL4X
PE2LOKegYtsAIt/xhhjkkna4Mc6/x0otMw3Rfn+LHdI3ecZYVlC1JtSp7zFPkx5W9BKGBUKeBeEZ
w9QVzAI/fvY1z1Z92GtlcpszPS4lwd36aZu7OM1R3REI3Tc1Ceih3SmLh/9+Cm2XO37+riEXLMc5
22tdvX6Y43UY1yTWovV6B5fmdDJcJpWPelZDTBfnvlr6BXVfuStHsN4ibkhcpnSoaxHoJy4Dv34N
mV3snyPpqgmPLWQhdmdS5JTCDyhaJP1EYKX+lEP+qGJRDNP+ij/o6aev4dx9eIgilzyeT8aJtvvd
wAUaDoeDd23LtQcNf16i/lcR4Vdnlm/TbEWFOlvEjhiEJhIDOvRgu19CoNuNi2tqZNDJrEK+HpoY
PGoYpiED6q0nyzc37dR0jKTqGgtOnIGRVVjH/8hnMDyy1TCBHdGatxvl1X/m66i24lqPSCuk7P2u
cc5gaccdZ+oFSY2u+JBpG2+jqUv8yDOHjKL+DvwMJJEp2bOJ/xjFplsSaA0UMn0r7DszCyWTaQTQ
DZDUr0kFCFZfFpfqJz3TXT+ZyHC0ppF7msYNdADbyeRbu0j5VhjldPtNQE/c8Ec51gXuaHwTKuRD
tcOi2inSXYfqCOb+sw8JL011UT+TdfhGJeiULeMKidaPrm/n3w+0JzzG/CCiQXVKrv90kvbV10wu
5/6cfwuiKriRSktvrA+5l9DmMvZ0CB2P+4IKE1pQ0Kji4uqRovK/f95G3HOXZ4MGTNAseFiYTteV
0+actObX/ubBBmUbpGTEA7oVr/zwObHUYH7MSkpFNALidCpCCGK2QBkwIV9HrVpwNVV3VPr6oEM+
KabovYgpL+u4JlKXenbFt/HgZ6JapuZ2PM4PkMomWHWVS3TnEzt9TWOhu/xZpth6oiyV0BM/Oc/6
By9UjypCpnUwzURUO5z7xc+0FtIik8t33O/h8woDz9m5SkH7xHU837A4KBP64c0yGM+2MHgLry8u
uG8qO/1dLieVJd0lN4CdAxIZNvWU/DskFFyJvMSqKDtvHX8nVjq6E7jQ+rk7HoedZQh8sJ816erH
ntcNhbc5rU5y8i87HrDjjQ168uh8oD1OO5gQU8heDk4txbsBpzHSSjVD8W2IO6s+7YraDoGzPzmR
oDqV2pZalHuJNBjksczFFHiS71HkxTvP6pmLJ2KvVoVAzSQ9Rm8C3b3WTtz6webHkPbShOQMdSl6
2MB6ns2rJS15xoqL1JAv46jMAWs9aU7kVMWMwQSfyy30NNbtOwX6sgOaNQzJhJFOJ0pFv49l+mJB
eDjK4w54rd50cvsUpMbywPLIf4q6ZmnD9EoFNeMjW2ill/49g05zzmR5UFtZSil5+L4qKhkmohMy
BR7pUAgpY+bLPDKZCvSTQ5Ix8VMH45z8TuOK5vCK2kYwkjg8ctnejIwScJGNusuuiU+gnRq4TILF
jdgO0nyqB1c4HFgjZoaBlYKNN7XY/fVCemsgadI1g008JWFsLcpK8IgPil3FHlp+ciS/PJop2wdn
xGUqv8BWV9+PsrmUGnhivj04+7FbQ439Xt6rTZHOPSY+OrJcQhkQ4t+8sbK5iaiHfvaGs1FV/Sym
/yRA2HhGRYQETvlWMbzBN1JH4oyfOOXpGpYR/cL6pxvxSAC+W7PqYzbqzzTE5zSBHL2Ia7sKRWvV
0qOADpmQbW8hyMH+lTqINcbgBg48rqJeNV3V4AibYxGZlyjcUgSl/6E2WGnlQQIGax629o33hXrK
ndnjhw3S4DiwF8IQOa9Ky+ZA7Nt0idY4/m5nzwlYB4sFUcwFf4fVruQ9DGpvZFpL4PQKLXmM9kBl
UHwo3nwWw06RTfW8h20kFxSxLybL+uQZih/1v2J9wk0eL+f5ikMKICG+OpaptEqeBf8EKNJHroUf
z86t3oM7LXtkI3Veq5cgvENz+QaE8v5TOMX36L2TdHU2grR341JG6K+jTmjysLLhHjICKJ+eldrf
7rfiz2dkIio4TVsxH4a71VUs2yOQ7/GfODW+fymRUReZZIolSXXhKspSbFG9AFASJpXQjOkLA+dI
/fjyZ3Y+NEHjnhHeABDOEHNfCk7Ujk5rseUGYwLyBZ8E5F+f8hn4Y4LuthqJXrD3XmnoAM9eqMss
5BRD1cloHVIdSQXhie6fMcKA1d9Q3mTznyw6P6IPeMzvkuJdFg9kzVBadKfWAzAdZF+cyNOCll6D
u4qc1HH27GPpkMAwOjD/CwtluiQG8cLYpwRV8ZB/xJ5BioHZZUngrYbFg8B7Ce0HSuxajWsS1MZM
Omp2VeKH+5Ed1aMxxQtVU/SzWv3anOO0k6sw/bm87pHS5glMMI9Pwjo/K7rQDLdrSM+1R6pgMfUD
RYdxcBjMfyXiHeWgGfW0jdUzJ31Q/ECqf+6Q1DX+w2xyer2/XrjXe6SHGTAb2XVoubxxiljJWKJr
+wtK75qx7MtBC5uUHxIDMTB5DO/IzzCB6D1Oynmiumw7356aHI/oMMh+05cZ9vLcsvOjKyr9HFe5
aT3iCYExio5Prw5Pt+zMXLjnTrkK4K55b7YugCyOtGK/l3AKyY5AhrwtK8TTCa1/E/L3zyrfHLGJ
AI25DGY7/k79TH3dOPI+tE0t3ngIJjtpUf510CZsPxZhPvIqrWsBjA5c7aYD252gOvXy1PuD1DFE
LwAIF+HVLLIXxPKWvtnBUhgkZPzfL2VAuPFQBxXzPvIetH/0OnfVte/u8JJklfN+/vC2Wg1tpWIJ
PhBabpYkJbcw63mkCaZs/HdfxzFoD12VFFZK6gOxaPzckwmZ+6nS1BdIJcCejTtNJapIP0auGQY3
nnwpR/FZokWPf/KnVwtExxSRUeDFqTZdqrvL6NbfTQXP1ScSks/WCmTLv4I4B8/fA6Vx4FM+dSvJ
Ux5JcTyRVOszDa2kUcl7Isx4V7/gqXWCsSfC4sCZr89iBETOAjUlMm0ovDSxKMtSdX2oSW5fA5tg
aEfItJiSYmnLneXzjFpcKx36vcoh6euosC9w4ncmjg7P0GHB8w5CelsyNkp34A/gVFpvhIJ9Tnfh
fJRm9wPh7IJ2m8NxqYlD07aRIjaEa9jB0sGxFaVZFMp6X6cc0lDNk+pxXi3ateoHKB0IupaE/gsN
3nJhTkRx5p3jEKXOWkKWco8gGkIo/5DntzFgzxyvXDvXUf3tKVXA2OlUZtt582hGHbGhhfnI7UHs
PwEPkp6B4V+fvYO1Gfa/U0d1a6dt0TX7AiONnCZx/tfibAVWV80Rf7eSxZrMYywlf2tXLXKz2bTD
6G8LbadsCfg4pPDvgGHu7gkpEnaNczk8BOwPu2FkZYi0UTIg/b5NQnj0RZbgP7wFMlijyUwGPGSC
wyHfY6598wAH3DCzqJ2fiNhNNa5gjYQVt0szYPXjJ85YCgZvQLWk8WyZBbHKGHwdVhjEYEaXxgOE
resQ3F8dGnFjJ0oLVG9s8ENVVOZzm95P1lUusozJsHx9R5sF49iO4B37rXqA0vw1pFoIhyC8qxH/
G8ovHyVR6hrOKVWztCM2j/Qp/QXV1kLbugVn2nn9mab1DfnY5thTeq0u7T9mvhkrwAtTk0cXlTcq
bRtUVif3bhfkhXsIsCQEGRpVp4rODPcsx7/+l5FG1L2hMrhy0YcA4lXmlfp0W8xCeiHKDvQcYnYz
MxvCMjfwOlMLyE5p8msJmSv953KyvoJjgCZfB90cZBkGOoxBiyaYAETsOS1IXir9zTHr/f0sBFmT
kiqmBIxIlKoh+n6EQw+J0SS9Lfek+c7gACgiwpmXWJpyLGg06LpDQG60aDfGpTpT3F2EfDiijrHE
h0uVntQfHx9Rp/vZ/ZJY8pIHIb2JvQaDboXPYqb9lcbD1TiBz4qDAu53j0MWedHRvVKm78El6Biq
eT3njc25z391Scr5fEXH6IXqo1xelnqU27x0jvyo+D1g1PBskb/kySxFsa+Lq/as5DBXsv0Jj5/g
M/6CsUOCnVy8INS0eimvjXjIACC/dgaw/NrX+pzFXxc5HHYh9Xw9b/Mur7NDP6QgU/E6il6js7DE
rs/r6qdFOUlQ79tglx/vLrGA/9mzEPMIkNeaffMc4BSR9vBEUKTDXUNqrjaJZS3b3bNNGpdXU3sp
3diDh1zr0R90xJkeSMrbzSrvwdb7nORa+pYNQUiwa13Y2grsoGXtKt0xPRVXl1Opq/Lbqszldi5S
/xaAK9VBrE2PPRU4m/F0CxABvUZrus/uwLd68BifMRITV3RJhGB5ZEGUqRIBoe0BSZdnjNornldD
wc9ZjHY/YEJCDxIvNrUTJ0bswi9t67UNKwdi1hRmlZPq6+RYToX/3DXsKSCH5Pjy9/jlEGSNE+Nx
zn4OFEObjwr8T6T7+fBXze4TxrpvS46fywWFkdXB+x5QZW78RHFk3j0uQiXt2E6uFYDxyodyG8N1
lSUgQIxqpLx2QiTlAAtfylN3q1VNRPXpMtZU6fjwSDb2M5qv26WfCfs4+e3fmBuf7BHOfyiNj+2H
eslDjachP40X2lla+5pYbgpbTlxGkV0wdcsPB04OCa8jcyzmpdHy6wgy0jPtcYPstNp2xmslbfql
zE8rGSFcEOtlxqAK6qsZSSC4TJ33sOBBAVbQQJndVYvx+zNmH7+02L6CT42bskbmLlFFexETYdML
LYxKQ7aUZF0vHzX4Qa04DKytY44t1PJc6w80BhDMx0nzZ7fcD9Or3uPK4EpPHnlpFRj56x8HjQqK
kIMvoFVA2I0tMcL/XRM+tnbesKqV4uOCoKw4KKEsyxSzHFMa2ZaunS4gaZgaG6jku7PJJ6klR9QH
FpHiDspS2XxCM06V7URdH3QxZGrnIz60MuXFfAlgqml8mUU1an2RLCXWR6th7yBajjnjGZPFkQaM
e3cUyhBrPJbtQuGMm/jFIhKhg7tqhpVqjiajA87y081g5KHDKrxvmtR/gcMzfxXaSaAkfrBrMCv1
UAiVdCNqSCUXvYrh2cXjyzx/b1SZi0UJ1FdKRVugQXpWQ6/90ynUULvj4CAiSOaKuvrqZw+65fZt
SqfWrVY6+JIn7SoaEJvVgbktVFZ2wMdJd+doyvBU9iIsxQDNNo+TRt3E77W0tO3a23bsWXuVMiTd
BfNL7HxH/GpqDU6/AHLbTllzFmZzONM9N+rOnA/nBPANpeipu85Z5U6jU3iUVY2i5oxrQtoZyKtx
0b+TOkzPykdt1gNvLlAcPAma3Hb+wuWt0U8sRXZKQP7klop6KX3gPZ7RrzCGlZBIZKfh/qu8bDA4
FzGmUwSYGhHXUlj6rD7fzMWI5SuuCx0mRClHR3YLfLwyoAY9gXZz+Gu5kEEW3224BG5WLF93IJFH
k4HSZ7KaKflFebB1YfpuwI7smb89STZQRt5z4ebHPby04QFU06HdCrJsjw2gBinkGqs9GdSEqK/f
cu+ozGxLioDoN87WmngtfHOH09NYXgORRvQaOnYqwghpKruXl1l+moK4W9I4J0UzkDUGjfc31meb
5l+CVAkSNcpseuDYb5QyTB+XMqfXfHStnWbJwLwjJcx2ihJmR3jQeVu85hX2W9WEZA0BW/q5jlTG
3VbmRIoLCcVC3UDAKFtqzTQ15vuZY1bZ4cNoE/NZbLYO6AtL6+rk9UAufwjuKtnCDHs0jaRFdJSr
Tmfh+rry5QO8gthVhYyluivSNPnxFcBZ9WArrIOjX1td/E8suhWfc9zCEXEWIO8UDmI4OWOqe8Ya
iQpnLL7N+VR+li3h6jrmEMfoNgH53UngqRC62yB2iA2zJusK3fAZo2tM5iWgA3UGUpq4Hd8C6Sy7
I9eHnijgTIfPfdWwBFgufcjKDKQP8zQ4Csw9xMdxUP/EVKN1BhA+U3EIfHjq5DVjDN4He7GZdm9V
bG7Dd4Vyqv4OGAKQdYic5qL1HCRTGmrpNolaIoHVEdb1KtBLLJQagkE7Tsb/hE1gBztZO6hY68rm
21huGMFhzFcbmm65v5ppO82/JeHfQEBKSntTUlwJeWf24XcKzN5OMsIkaK4UDpIx6g1eMNVwht08
mXlK7ieEgiDkU4u0BaZGi6XRB1qvsgIbiiqh4YGXiFxh9/PfxvPF5ZtnA7DyHCJzhAg2AhDmC3Xe
5q/SJAEw/U0gLTWwlkzIFYaVA6TOSJuyPGqEzv4rBbrY1K+/ZzAln6c5aA51S+oF1jwWZZhvsFMG
6FjV3s6v3h61oqo5bww3zWLyoEVe293c4CPhQ8dY9s34nyyuoFOmWtgIWbTbJzc3jSZyd8kdZ+HP
b2NPdOYKCaOluGXYM7eDHO+IS4GOy7BqM6bh2c/LWsP5FDY+7lmPNhGiZ37ifftorQM7wAcvtI7S
G9N5x5HuwOmZNgSTr4YtzvzGMxK+I08vD/Rn0Br/TUOWyXgg+VuslS/XyVRjy2HjVmgsCNjr2XXO
pPziStsOCbXaPyclK2qszZQgCFwpnmia2yAozS1Fswto+lB6o2paehMIkDOTHsQkFakeTQb3Jntx
3WyralbQ3ZNd8iGL8tivlojiaPATpP4q29He18WX29pys/K6ITKMbDsiCMITNhLv6OjMb92UYvQD
O75agmh7Rc0Hc2zhXYqNOYUffPFwxgCPtJR2KQAuooLL+WZhzTm1ox231UayU30rReJPM3xe1awr
lX2/LTcgY07iu+zOAuNxIYzKqvxZkfG8iEoSY2yMu6ALAGMcq49io3gqWcgWJC9tqB0TXL+ediez
zTiopjbGwvzV11McWGX+kKSAWFjEQ2Lb30k3wrOv7c1lrFda+/0fc4tvYC1+OiEWbxieQWGRjKqh
NPa0VbhlRxq/YnY9scCtpyYBuGZzri7wqdh2SeU0kskOYNzL6JCO/QGe8H2RrgpzJS7tUAk6trKw
KDz78uYMUmfkWEGn7l90ekGUZOBowZ7nwr4cOPVjoiE8dN+zJ3Pp4aV7NYc/YILFZxPY5MB+/qCA
RhqZAB5lbV/wmqm5ps7WozSr3XVR9BDcJVd4d6CAaDgzoRIYR9n/bAR/U/LHiqZ6vdfKPBWBVYoy
HOT5cIpHprFe5COAHyi8rQ2D6mQxJz2C8jBZg9ov71eWx4Mybm5nbVbQRSpFtAIdD5d4RsLW01rc
u0zSB01RKxxCENItzbFTcfJZ6NgFS9vSD1iB1zeiyiuOzOBITUNtDWL2heMZ1FGjxul3ScKDPBJ3
B6sE0oU7I8IenxHF45wFAdLiACkYz52zNV1vC7bA+u0naiXjhuq0Ax88efwr6QWbsRJUrFzrE86U
BSDMgLg96rrZePbqLQLgwbbHXfjy9oPskMxKMGN2vQvpqq0eE+OFGUyFApHJgJddLL+48GkQ24A/
abj66tWiYpJhHwap4e32OqCqkcK9ssAMe9jorXL97R6ytdKSvFq3RfNch+kr1SaJoQ7kRBde/J8l
BST35yW17BuBsyYt3PFhzaFXVJF5K3q06KymJwMvc66a2Z5QM4+hTTYzkJ/rZYNHxZ7WOIvMefYM
0iRhhb7vSH52/T/gRwBtTiOs4q9U6iNA6r5DH7ddUWVZsosRyFgE0poBl5/660EH3AtAutVCQFDc
mePWeoAZQZsXFOO7ZSLvl80SGUBXb+377RbogqtHlVB94zj/dEJGeFw5RhSnXDhlAXBiaZUwNBRx
1YvMYhqki1u2fmVl0j/Ptk5UtHox9n1RJ/CA7GMZtAe+uln2WY/kwxuJ9Btetcx/GKBubjpeX+Fi
mHLD87H+l5j9jOoc1vsb7Vq87LdEnxFTzffj8/FFJ/Bpav4mPDbzrglOlm3uwb9i7nFt3rVHrHUe
ztxeOZYRa9wLQCxPxMOTVFX+mT6kwIfLWiAg2RkUkFkRAouJtywNCU0Fo2wHm3LU671aGPuvX9a8
05T3h1VJOmwoi0o9qaZZjA0HBAHz83vmHM32q07Iwn57iODNRfuKGUnoJE/qx3nOKAf9urMnqZqy
iADVWdDBUnsf1IlpNs2xqCwcUQBgydaUfz8Lgi40AkHsWS8U4d4+94PAVAd8y4SLHfNFGpStbzx3
0NUi2yRyNyDq8l9IPoMjt3V/ota5B7x+5/uIz8US/PEYim8/67LFAkCglmjfNI2hQRAbQ69AwC+d
5VnbTQvAk7yHfCNV0PpUCUH21vZPT9cBMWB1KTsfMf5aKIvhci0D6Mxh4uqoBttJg+VpJ9cJ15D/
wud9iO0B+tfv+8/BxjaPWH8axDkWhDW8WiBFb8fQ51usaP4UxitBXCNO7iQyVanRr2f7nK8dSNAS
VmeSl2XK/L9u6BDCe6TeMVr59N17LeJ5bydPMQNjMg0JJjjF6t9aJf4NtIITN79POfbjxUcK5d+9
dIrGftubY5rDlKBs82tLzF0REpgta/MMjGNt7nM3ZEoUIXiya03wb8b65PpiEgVixa8WmUxx6GUi
WvRIFdATRaj3bZneRdK1UGA+4MAymXsMhlK8HOXATIgZLDpo1sGxtHlwhnvE3U4OfitrEhZnJcw0
JzptI2aG6nlWmq+/QnTYeXaBK5d0qYOhT1duqNn9ukiFAzk9HD+oXyDyAM8Hw96Sb/B9+sF7E08M
Vxw6q/nj2l3SvQ4QsuPhsT1Th0DUV0yHXoym2lqYDdG4f1y4JUURigJqKGrea9GBzltQ/AR/06RS
tw+oB2ExuarimN4ibZwidCPBESTF8F0KqQiHPICr1d4Jtvx8Coz7UdxQKbB3YZOGDzsRiT7yqZDb
G7Lv0UOHl7IYA4vxcHXOD3yp3Gq1WnkMLzpKsyO4vykUWEj0BDdWtessYPiLATnKPS8WvymyRj6h
oLvwIgXgLRBWv1LLOePdVFyi5hYf9CNKPSCqBT16WFMPBLLSjAcQzbnNw9rtSV8EckJjCi5KBTM7
a4oEvEXQQg2eiZjUkkL2bTH1EIyzAY9+BzG7CxLvh+XlINzDV9bUVnJ91JgbmlaWSojfZuYek+NP
zbubymPUo47YI4EouXmYQVsJYmUt1SmsC13Vh2/I9u50Eud6jEMvkrQrZftMlwlLHmRx5YPg9rYp
lPo9H+Bj0Z2pWoDD0hfaowIou9t7PN4qj6HSdtsjPYFws8D7LmvHPIp1+gnTqOUtQl6R58LFPYCK
Pktx2Y0kmHgjmURHIJUje6DxThO2dDv4sACg7x80NvkKCw/z2Ovz3fy+/3qfhbtBKchAFns+oVQD
W7e9ckVj2U+viohsOWtEILB4IEZSrIMECemtjUi64gNCV1RlxXmwWTCP8pRCLB328Ejesf1IdzJU
Q+q7IdJl0xWbD0mTXFT40rlfPOc5GW5h5FvD4Ar+pQyrw3NMD+BQbc8u2BdMC7mJM6epquHPf5bH
VPEOOQHBeBqV7HN6/5uPHg3gVZRshinMSM65oYPwhCoDLq8nnitDGDond/oHn8XFao9Oy2K3oJQ2
zFHEaD+/T5C/UI8Sq249NQApgp16Maf/0Ot4pRr9BJW/3I7qP1DnvRQfWAH9NDugwDyHk+ErHfnC
TMU0ZpsqbD7s2hLSbVh3oB+nyXUniK1LbBqSDdGXBIpRy8/Xv0XD8apjhcVFCF8r9AsWJzoB4J8r
3q2hX6zcA5GC/ozFh8ggcwhg4znmJqxHDPy54y9YDLpZKBkNg4X+rwRFcCVGEYP2K/i6cI8yT5fx
RRCun99WgIyasyIiY9CTjJmncV6O3ySsnWe92lHj261kpPvo9NvZKNWvL9Gt4HgH+XCuiCA6C1E5
/kmCYB1t/5xxl78/gLbNzi79seFUi8w9QuwGEI7I4zP0bDsZQnOaCCQDcokICshX9taFY+qRI/Al
LpegqU8+pRMo4/EouWxs5AbxjBj0sRGit4W8s33xjMDHZ2VQ7HlHbcpMLVUaRRVusKcogi5i0rvM
nqKbdS0Gic+fB0JIZ/CB86Ye7b5aq7JbB5T4vrgoPZFI6Dse/U94fpgDAL+xtxkYl57Z6lcy3+E3
owTJ29JJ2nsRxuC2DmFUmzsv4ff9qiw9NLP2Pwla5ml6SHCglkFX52oeuI/6/GKlYaIFW0mnLHOF
nepI6wO+IYewuSkFe9ncUe38UcdsfQwkqxOm+c8afvVoL0VF1ljSCRRXPGQ+zDazMh12u0kX0yIK
pZ48NtaYakumf+M34o0wfhiUnY0i7iMAmJZZg0ZIs0lYVfoj2/1xiohPtuRCm9/UJBHevgpX7uoS
I7tICtZTTVe84w90EjZv8AjVjLJEq4HMLjy4HuNnKLSgB3Mp5nnL2lQBhZPAqKuWxgW7qJjfKpLG
fo+IHWNLS7YQt+E3YdO/bi9BPLIMTOMeIUj2TIGoxny88fjSqYcxDhluzrdyWl3QDtAtgdrXRHl/
xXd7ymjCYS0eXudcHW1PWOCs9RClx8A4YhSHjooaqNvXFaqJ0VRdHAD/C73TZPWQoTQ/IDI2GznE
S4ysvxF5G2yxwNEhSOg+1FzBUh26oZkfiX7xtviugV/WuRhMKSGLNR8Ci5EP6AfEu1wxtcxRTHAu
5LONdQ4+8yfigP00YuGqRg+4XsNpNtaN3/0Rp3GXpJTNtdIqZlbZfuay8HpumiOwXNJWdITJhS36
aHJnxC6CAigdRn7xzlsMAyOe7pKYgg1MPvklNm3xZesdR4V9uGgIBd2P6MM719RqwjJB4wl9Mdkp
Gfl4jU0Bh93uWhSTtqGFuFsWYeKZW8Bazc9RSr1jWYqX4W+7hQKxIM3Ee6YPR2HnInkTdqBDBist
KRaUQyhubP6/Mc83IdGvSpC8f7pAunvyK0XQr2QgYDtMpNwOMA1KqaiGsIHXdGLk0FryD8ukFl8d
yK3GHZJXt44eEd/PfaNuSfA6t9TnrxId9YImZK3TfMS8Lf+A9WpnYepV5Vbkyg6fLgcYj4Kt4BHJ
SjITe+PeDLvVBextA+aEOBNJ5OpJV8yEHtpG5NCAizPvG9iKZV2MnGkiTlplAApNZREKGo2kX8ET
PknZOk+NQG5TjCB+Kb3jFTjGdK9rEsscfC/0Ky5BRmRpliktXClT/at+xkTQ1eF/RX/hM6CFE1Fe
mNYhKuid2I0ov+0gXbUCjyl7Uq1Faa6lkkUn785iS1SeWmLLXEYSQ2GeeKA0JmtHPgGgyt/jaVHb
zeVa7OBF2kNHvv1fbKS0FyN6q9NV8SNmCozlnF9Yk6tI1bOJuzeXl3mgGP93k88iBB0iDFcKP+G1
VVfpXD01VrXrBzxo0spyz6D5BEcx7hTGM5n6oPUBxZvb6t2tnT6PQtD/uLwMAnZsP+Byuvf/YSd2
SZZO93DxgsaZTWzSKKmZseIwhmUI6eZu2bESG28rBN0u76lnSCLa/UGY9Hhymzq7jIlWAEYicIAa
Z26Hc39jDS4wo2cTUZsncKq8P425xsNa0yHCIgi+KM8EXQRGeAGnk2Fuf1GCRRHHgkjN7g2meSp3
qUrMXbPrVIgfFXdUwj1k5K30MP9VBFn8mJPOdWFdV6u/Qb048V+0lfOzj5mAG3Cbon/6FbEjnll9
bw5bWw33gu1DZ/KtPCdgShIrvprNp3t+ZyWjN74VcyhX+5bUyZDkXwVFsw+gRcLcpQXRqbyZons6
EPy/ZDlogj4VmGZnypuiYH2+EV68gmHHnj5EqPdVPN/kVlhPdqXVz8Me4xD5eIuH5DV7/qFBDdoc
XyLw7gVnZga7TyHHbgvLcY8fi2OckPv811h4OahpF25BU9rsUbhyK56OEvuvn2qAPRlsWdov76BF
G7t7IRliIopjXBwU0l7wlgcund2bqHsmdLP/nsrydLz6jLsMTk3H1Kf1O+oe52b7C9pZnk8vfOKq
6poCWbgkjlverYqkdF6VESCYKMtmk+J51BkASG5H0XKosCO+F4N7rQYLhC8CXTvQfg77kovjRIzT
/REc0K571hSc5r5GnXMvfEyJLp+k4BANAv/OLAPRdAbDWSNRI3fhp/h5FzozZW6qDXrv/ZvSn+FN
SuFppTvdGqv7yUltyg682+8xVvJ/yZttjL/CUG44h0FWICuzRRfgSjy6Gv3vj4jZ8ljlmohCakLl
YKkVHTtwLM848JH9KEkW9fdP10Dt9ni+6uVkR7TkhnrL+vtFn0GtS6J6RqB1IxGCiuSnMbinvqld
KD+mwjYUBIvKx03zuoP+UAUYVPE7k64ajD1nREtMDXfhtlKj0cN6ugVUT0ZtbFfFRUYT5hL/T+j2
GCE1UXqkGw7lRzbsXjZi6NFfzrjZAyy1fPxTlLi0TXlEecYCkLV5exgTsmtAX7+/spQZ3d0ZnjJD
9OpEPf91NW/Ze/0yYMGrEAhCG1xpuWbYqkC5QN7xRSMalZWV1ZjQPjx/1n1spJRxfmelUJaK5RJQ
H7REtTyvIQiPnoBVQPeGP2lk65DWlLl3adyh9svXgxsGU54lbtOX1qXeupr6f3S96K1Od/0lfi6e
nkagIqiVuO+w03V20ISVOKDdPSEhoDR081iTfc8k8lmuYuDTGAE7UoDFP6ZsbybXMly9BfwAC0yw
zxibMr3Hn3SYWIqn8VCICp068JZmpMtGe8+4cQhcoe8cUVV3/dFkWu5ceMJH4L9Dp0Lf48IA5PT8
kwFbJzOeuHgdVwL8+5EWgK4tdiLL0JCxn6cmhNyWE35fWOwQfjwmo3Fxh4IZRCVM2ogKnBi7ybvC
cHoj4i+W9CHaAtMFeiuQdbiL4TT/QIyFbMmxC3qRDGuX2xVz4OmxooJ9Y7GHoEa+KMUUthM2PaiE
msD5LXS4K9vZuK2VhCbVXhyqAKQh8lPKgtFaqMW3WV3WLVKYOhfMqySnelAZ5nTlKWjOAr1ugqKe
1WdWDCCnhsGSxQubq41Dcs2sHPegWewvSqziAb3geKACNAL3NPgIlUIqSW/Cb9uz2WP9KfRnpdTN
afHjGMDnmGRxzYKVyrl4XDYPQg5wU3TYei7dtgheZ8iUDRy0yOqV3vf5ln2evNRvtXZXCkkvVRIF
5cxQJ6NXjS3GK5duHiv+IP7yY900blEdNFH+rMQEN7ein/PSkiyh0RqiFNBjaXjM4aZulBXD+2ow
HvW/1Ukddwiwz+kXiEX7wdZs6FUCdpOhovb51F8JqCOt2Bh+fqhwIEtVoDyK3HpQAVDpAEQO+DA9
eZHh1yKVMsc2S6RpP7bbQDaD2ooz0LDf6zf5LbJwB3g9JErilfjLvhWgv2VfPr9+QF8jP1bbc7z9
vsNK3DMIuBLSpZRztFmiYzLo+GBG2a9o9vVTfi5/QaxirO/PWZqkNdVI7oD5a8A+Cg0Q1tiGp/VP
l/G+4pI0DrD5mw+AmnufOS5DpX0d7FA7kHO/2NzJtKwU8NwBQk+VEaJZePVLoOpuZvqxBKgfAgl6
2sWZNd/KO98/p0ZIpourPysIzi7TqqF+C6ICi04oOCtVY7de/beWjm4Z+FxZIOsCAbor+4BdLSPO
sZvkoWe/2w+poy5uK5q0KLR2i3NVPB8EgVL0iCLcLKUcrxRYPD70hmZtY+qlOhhfCFf/okeqWIxC
VnCbKGANsa2tWRlmkfQRkrm0ACEn7dIu26rboN18qE/cCQ759dg4Qp3wgM6GVGjCV1FMmE0J3VBo
xUyBB3G6aQYdBNipO/n2PQjoojdbWRyhPyEwDaEkfoYOO2ibfq7YqLTvAeEmk3XHfG3lHkljGI0N
Us9ucx+qQdranE3xVE49C30alYCu64xhS5F+qMYby+aeL4ldiRuEIK4VPmOfoueUhQWiuw4s1jAr
ISktvDrYXOyS3eOMylG3KmF4zkVc/AmYdKXsQY1NSBdshQKLJ6yO2LbE7cM+k2NJfvAThTTUoGR4
wDIaYyGTmiYxYI+oa/aAeMWJZqvgBDD4Y4cHFa8y53O00PiTLfhlfCtcCI3VQ7yfydqivUNGHcj1
3WOW+vNNRMCU2EVVTSQT0qQAAkdXm4wy/MKwDXcmIhwwU7xv41BlSuoogBDvtMjmtssHZ2p3puPP
Fsd8jtZ9ShVaWAHDWDykQqTkoshZcf11rJAhnZzw8i2ytTfcrC+Lb2DrArBfhCerltqGvpM5vk7C
LwCJcMvletFPJjhtD8KrJ1iAB8oFkUaU55A1HccSdGhrcRPxqpGVN7j8o2gr+/eRRIflEu89/to0
gaqyad8zzK3aT78DiAUrzuZ8fe4/eyzNx5wIO3zlOs2AyYcqIbHaFXvdo0KZGyjDWZkkU6m4yrMl
pTHj1klV3LVAV2J/2Kqx3UNvUmNFfa20rJ8JzjwMTIqq79KQsFAAysDYzkGLdLOjgOnHMH6C9A1B
hh3gfCAhNgT3bwXVs6K1hH4JZJslIZat6y7Cm2qLQmc3249GEHH9U600lfrSUT6uEurOA3ggYxKI
SGnDSv001Z2AW57fANhx7Xe4xCDBMKHwR7DSl5yMStX2XrflZjI0QVvty7dxrsgelQ+A0e2VeISx
EMPNleV0HwogFHBtNx3+Gek5+5Nltisoe3weka/+PICIFhrZ9n9vVWSKrptM8RbCE5XOAL6kl5lW
GYqT0RAqMFg2xpf+a2J6us+cRfmUlSbp+aA+JIrxQhraXc77wV8mlkrPNxAV+iHNZERCxwL0fMeX
SXXf+MwUlqxcBn5EY9zak1mxZz6VOnospoEQIBWXWfryjBLLi3xLv0v6STb1LktjeXxOnS+WvpkX
42TmU9v+A9Vww/DVHsczTLYSPxLlfUw5IG6cNgVAoACr8VrwGJkGZ6yBvSUbSR/ZYAM9ro+9ZxDn
JTis600HaVFFqhyIBQE85F5sfqBnPMTWlnIIC1CdJ8OGSWrd0Mt9ZzLeSTyLiNvu5mDnnk1G+d0j
G8H13gsr5PbjefdjM/+HUZhy7wPXK9G0Cs60IdEnQ0V/eK4ZSzHemc6ng0pr2kY0lxjSEgF1uqiD
6n7+E9ACQH/h5aS/H3jx8UsjytU0msz9BH8ROXH1ygxWR5S92Zl6DOpcZZnzcbmnrwja/PN5PsD8
ScXRl4QHBi8KAa2EpQ+PqOtmR/p+sNHJ83HBXerA1UOufJzqI57R5SbLfX7ZmdJSK/cy59QwaZza
xFokSLyqtDUoDuJe8eEOXwjeUxP/itrTt+SUyp2tohqu3UEAwVqI2KUye4H54CvX305Sv1pg7Kit
+HVEZTg4QTCr+n7PVmwRv1ZgoaaPGrgDx7Gc4ALNKjzdtsdtLM5xWWtofMVXtT3VV1mLKpqEKTJp
WDxlIE6NaWRJsGQ8DSE3hKnQ/yOhY/S5O5dtsu15/f4HTqV+7iOddYa7UYA3SUB6XvwHikjh8Cst
K8wqlCMe8chYYHLs4uep7Qyatl6uY9DV1zZHUKvfQ1LbVehY6ED0dQQdogKt3aCaCs3sFBY8EyLi
RCKCwAjrp9f41UtlabHFx/pe/1qcmT9PZdVT5buvgMaBYOlZVHrSeimfpB8899OQh5JEfGTf1AgC
BidmHBF/SkVDV5dzdK1JCh47kN4TU2Mt2d6Nqpcm1X+Pxwag2WzkDBcY5sbNvMk1cyExTlQ0O8X4
a3RmGnl2J3E4MM37LbKWe13UuVeJxkw9n3fHPTB9iUECgVE+FkXUtJX6Y5YNIxYh0CGNuwAOgxl2
bIUwTlIX1VshzWp/H8N2yn9Xh1PgoVY5OS2/ZG/wChTCUGv5nGcR0ykkjbcsGQZQdMnZydWjBjW+
EYCHq10OvZ6UUhwzpKA76Pu3iGLnMCuILXRyTfcVLoSNTIvJjgXWcP4Umuc0gFPMcQuKPM/b3RPe
+xUmyBh7GZUOPcpFRdmuP5b5oUYmaPlm0HiF1p9Kyyo2DpC5BZpTZvedJVMAGFHlQl9b246x47HC
tbqssB8AdKfHalvMOXfZNPYo8nuvGlgvLrxigY5AEQ3AoO7qg4tbroNbruQZXL7HHuNgVQ1eB2dY
uA05FnpgR2CjV8WgiPQ++55oFSH0yidyjY3PCgEyLHqpWwkoKOww8RlymEhHZB1emSo54m0+sPjW
5LWz4ErcvjQMeXn4l7MMl11/lkGmkz6vnceS4+Z/M/wl4ob4s4mTxvYIhGfTm5/EvZMzPM01/DFc
qA5KX+emqMRpIGZ1B090j36nOC/Sup6YAoTcYl1V/FezNV3BxWHD07uWRGbow1cMJuuED1K4tPM4
tZzN2QT1KT5ZdS4lofbn+C2tGWJWBl7LZ4gK4/ieQLooo/Pgtm36UfGREBNapaB3Gk2LyyW7Zo6W
rJ0vfCMUimP++TnU/TM+TCv2YCTtwRUQRRXbCZTUnW51/lQZOdv1rklwJ0QbdgBh/d17daQC32cS
O3yaN6gR7aBMHXrjr967hfCAGiDSPI3DD3gSJPdixz20/S+xlUc6v9NkVwSUG3IW1YW/yT5oUO8W
pSP6vssZ6u60s5MgviKyEFFzrMKZAYzVNbLiby1uwuWinUaneWhT0Mp2jwcisYGC6ALb1pkKzEpf
XmetVjamytDTpobFjPQnJ2VwYsfIbYPb6rPralgfQpv0DHN1+Obt13YJKWuzTAfEHC16PGIBAjm7
wNu8WUSM3OfPuEwUkIisDhcVQlKLmbMxL98v/n0IjUurk6eaRuh53gWJeE7jfPG96kaFxWrEjHhi
U2Zo3cKAFOmNweB5j9tOobdlE0BHP4wFWbgjlYobcNmzKmMuiVXX2wf4AfDfz/cGj1dQgfvOcMOd
5osqWCYn3cjGCit0q4shaeY5QuWn0RnkbtF79XWUOIuY4YKuIBis//d9A6FrL0qFrov2kY7b5PWL
X9Z+NDC4eWd8Gfv0EGhE3eKhXMAEeLgBWjhcf2rX9sXZKsfA1AA/5ql9b0Uwvk458rqtb9qV11VR
I2dCc+kDD3JE4AjmABywG9zkdFlFc8KDOsAWEoK8LdAv/qBR/vU5mQv4UCislruwcwMPe/WQlZhN
YYj1NUC3aqa2NcmVFbHFbkiL8OOuMf5HX7cHTy3oZeoyFD/G1Pn1JAIdaMPjOgcmqxioSPzifDjw
HVewhACW1GYFAOZ1Rb/b4BjXr24LneQz8koNIvExiVpPbCDWMjDUo7Vljxwbcvgvjgnj1S2ZENuz
oQ+irJoT+P6qaSOmDaF0jzG09LWowgAwkE7TFCxY96Vy0UOsuKFTR3/58lJFs1WMyt3jKQY3ze31
s7SHvjon24sVKsfQOvpJWhD9QtzEwoobNhe071FH+ObEuI4t3a3ujORHOIDFtBpdIqfRIOZl9UOn
Mq5vQpxrnql6j7OCP2SHTl/nCkYWkEWeagAsh7/SdfHgkDgkB4HAEIhJ9jM/EJQOwjf7uOWqGHG9
ZHjKBUPErmR1BfGA3dQw/hPw6gvUI46kK9SvyoZZIog6BFEKtfGVgpFFhb+Rb9ka6LFOeru5XBLg
LZsYcAkp41ouYoSNEqMLcPSg8FsQBbq1kEPDM5o/X8Fb4LoozIRKQHWHnaF4+bZA53FmFtXYI61/
Df6XLTIYGylfdw192qvIHewWxD4Yyt2LOVWitr2VpTf+smaP1qjQAvOyuIzWyZw4M+yQShqr2oAx
EjRdFF6xSZcoNwDrB6/BjHtL8JyNvXRMhnJK3yy4e0pXvntoxGOu7VMJ4ME1e+Xd2hJDcbPuGlcQ
fFcUPLIvw/3eSvclOCL642hPESwR4N/UJQ/oH4jwnMskfHwnjb31XK2Bbg9zPmQBvbvSDieZZsyf
zIrKs4NBGjdMuRyjTOiZZN1S2xjAemtOD260kL/sjo+f/ykqM2bIkDc/NIEN0wQj6rhftboilhFz
IcniKnpdat5JFKdwnvpIIY1dSgnDKeQruEAoTWNAj0aFzfQJWcrBN+jCmW7dcdpfRC/K1/+AwUDh
q5yfEj4r8pj5QK9t//4nIZuzs6iEtlGJIW0OTY8tWR+/lRLr0DBC+ZW/rnYgRbXiad436KvY+g15
j/GXZJGriRyVQL2XMcKTWtfeXkBtBiC8jydYnNveT1Xd5QJ8YAwMztbw0kBqqdwYDM7L7aIB5u9r
0UB1jpWGVUbZ8R6yBoAmVpBD5PSVI9g26ErCeM46RVDesISUNbYnBe3sabMvByydwdwuiNB2LMRY
xNAHT03bMjmrmA0aI4Rpo/g8pzhz8wFJyBpObNHurAPrb4PnSTsKvn7fBQBxC1/c+mSWVIGwmx7M
TxTu1X0Mo+7crn7nMzV0B2VjhsoNf0mhpwsXBlkLencO9iHjki9pyr0U/BmBUKQyj8JrsulwPS5+
5xFcbUeJijeign7PZYAyPs2FdQ+BP/zf/oOERuPzQEdtbnJG+Ot4HK7jEX1a2ebU+8vFfCWAuMJ+
Yu09zNit9KN1sxO8D1KJFViuS7xJLKCaJuvqAIcidhmMKz8JDNgOOLwadO2MGxgaMuY56rM29kCu
F5M1BGsnKIFM1jG2Lm+yYdA/hdBqwcJHM0cJlaonTQrwJEeNL9aNS8Jz3O13FKDvfDk2eDjgk3yI
xb4avPdKzasjbT1amVcIQeqpCpLITE/CaLv6oDEmfHhZS/KtSfYIBRbFnosQJMYi+2zZTM5J1KFY
1saMOzfzMTE0vLPk2OMQ4ZCf1UOB6Wqahh9vMBDtqNxfdHDfkM65S1B52BKdz16mg0t6DUWZSJdW
Va6a+pwQgji3WJn9WgNckjCA/vAJLZxRX9MQOTXZW6RXhDPP9dkS09W9sR8DodnAsZG5msCBSH3h
nvjkQKCxaS494ooiXr8plaQzuzUvqQvc22JXEcc3Or76HJIHTCkNz3C9V7ApHKqg3J00kA9xoWEe
0biykw6JR6JS4HkBbr6fWZU/LokwVlzH33EX9e47xgrbekde2oByf8Nf/QnAqIcmIbiQEWUXEZrh
/TFDOzKtWh+0GWf3/2SUx98PEIVRrBiYHsZJmmXklOgszrrHkad0L43sA6SD9m0qmJc6zBinbC9u
Wh10/d5eXWoOhjiQuwuib2ZeTcTmw9zN6eDIEntO9HhIyMO415hRa/FtYu/xtzXU8UbCd/JwbYp2
3Je5OpKwS7+rih5o8rxugOx/2735N1ovQXB1ALcCx2UpLxciVBPrgzzDZ70aSUlsFIoEkViVXM3t
PaeGQE76bRGK/xxoY5tHEFnZunWcD7E+98TnSz7qAlFml7J/YlKfgpXekwduRgV2esyPJCB/Z5X4
T9I2y3QfKrWYIcJ09qq+Ja/nzsd2W3wgwykUf53fwkh6Hn412nG9Zu6eDkvqbT6rslpeEs+AH9JQ
zucOtx+SRovznOrP+p0gxMYUX6VfnNCufttZKizDFvKrWXuSWy7yk+lDvIIppOWnXYXTMrdeOBuX
5MLiUkLEfGVHJScWReH3DXiWhA9muTjMWkVPnrI7TUc2sGxiwBuq+GMOLOQI5ioL/iJ+iJajiYFG
H2NKG2G4f1BY5M6VdjxoUbC0jqaZxOzt6DL++nWfKlRNIrPv0n/1JM77QywbYCwEbIrWUmq0R0nR
b+ckcxxJRlZxZDmrQAr3yURPFAr/s/+qKm0XjIowYTMIi12dLQOFtlM0PT/9101HbZfZ8INdVHQX
nubDNojU+LPdusj9cxRcgLEx4AnNmgIm3o/vXEqOQk0sC0TA7Mer6dlsmV7CqePlpyajvDldSHWV
3NUyomRu/j5XCgtJ+aJFcRoKyntajYqpM5rt1aIgX19w6ofiftf+bY7aksCqp0heOfExlYWrSBM9
SloXfyAogymErTlMa/Dqepx5oYYhrGq1eIY4TPOqOh0Cj9dqMWCVSdU8I2DD4ShGDqzlZUYT7AsZ
HfXemtntzPS/vvQHBlOmx6YKdgOZ4PWhUUPGKwaEhulhN+g29IgMyFDsmeYwZ2/sHa0Rw5pwUzx7
Uw8M0m9t+UNI9Sgh5lI99lAC61i8NnVta1qoYKNeTnl6nF/7HTVPPiKDSKk4CPHs58HHy1RmW9RZ
b7MxqDIXhfp1M6tLnMjL1pXLnxrbXYbJZ61WLb8aZ0hVOLuF9J9238PG3Fqn5jeIpKWrSskYAnkj
y0yPGNvTCxb6KxKCv/rcOt4lg08OartYDGTKpkdTPc82Q2N2iOpVce3zQHFL27uHS+mLXZyjTe7k
sYpkSEZQxfeKEglGOQc3Jl5+cE9H0tARLDhdDEHMGt584sKi8gBsMx5pG4WOSzqSMf2BetVVm0vK
vKXkOrzUR3nRDTIwv47C1/rAZFdggYwBCGVlZDUT1J9HnoNLrCx3tnL3tCk+I0G5Wv0abTnnZig3
WHvdn3NSEw0uFPbkH6KfTcOJVomsV0U4P8HbfDHAnouD5jLoWIyM7rziAQLnY6uw4J8nOCKsN2S/
H0L1EbPB+oJD9RmsPBlYNj6JV21JIR38WN9vuOQH3akUgOUjOua9UQjTDPGBxDGE6j+a3kXl+IGV
1GkgK8GXudL8v+OiQUFBXFhnO2SZqGWcqDJZeUIVRdMnVmrLJnwMy56LjaEQ50MpJ56zyD0zIUr2
VvFwZa8/JBiAsVQEkWzaZi2zWSicLwOrSW/mW6QGRj8HVMRMjnm0bWYBGCG2WtgftPcyy2Ru0qKA
G6+2mzgKkibnZ0FHjrkEgRNadOTAsBStjWhm60AVAxG2XI6c7G9Gf4H9LqSuHtkySg9Afv7CmGbh
DHsf0q+TQqHbCcMBJcL57ueBuLa32IFVu9iNiV2VgwOHnHrJIjD5VVgJMfy3VflUnFBjTfp3zfgh
gPbuZLVxIct0pvsNB/W3p82s0ZPF4rk9xPl0xfgqtpllr2QFb4hWpjLGSASnT7qaGXXLKLGCxVBu
2uzZQMhk5P2YrLBdwrlo/PZoTqml2CUc61mXGE4JHDAZW28PyvDFM7nixxirPWsdlTCuKrigdW68
sq2zmeH3UDq/4wfjgvqkF9gaI0vO32G2O5/gjIikenUG5UFgjl1UiSzw9PGYCHtnGd/WWAJAR6tW
sgsB4PsGzp/LtFHvnG/Iv4xktS4IcCEI/xHwqdq9w/2xM9ienPqJcet37Uj0ydpa7Xaq4FHSlhAk
gF3eNYo5cLhGILZJ9QmEPGGrWGkCHHV6E4TlFmZ+X6aHytjqTY0LnFxcwj33elQZs8xP3/hxC0B5
/1pag85e8+3LyesCBDENN/IBWcYgkGiJAo/T2BS2Cw1psUgUXVo4AXP0KsB1fNc/1DZvKC4j1Ba+
pY+rYduLP9yr8r6d7Zvi+HNhjBD4ILJ7nwe3PgawvafJwN97t4+QsafWjKJ5RFg5elbYTBMaMbEm
dL8EPTkb1kaR0qkZZyFl46Qf/i++hEP5H8U2LK+mc2QMFzIzt1pclkxT5rWRXiPjO65PJxj2rj28
JWjsCI5QlwSfl2vabOxByjnTluuOdqD1X45fFTlsVHLgMVVq/lNG3Jv3XBNMS20bJS5zi3gOaEpu
kAATkGF8H7nVnOkoeLCdJv845Sa4hziDqqDvXLaanr+RyBB8/HozGwa9MKiwHkCOGiG821Frkeg2
LvD4IoM3bgV5RUeiq+slNY1ykfdRlRgXTvqXmmkrrpT4NNk77vlaJAjGT3JYGAQpPBo1lq9579Nn
Bh5nG2lxIkl+/8MCly9IxfCScq/BfwmK4xP4NcnhuvHrC8ya/IGYsn2zRG1YS5kOlWNbsciwLQ0Y
wGQKp9+9yKd/uPvSN9+SL7Nzw6JwBRqUD11Yw7U6TXiWQlycFciTzDYUZOE1uMtUUbK2nCzpYFpk
ClKLypHUwrdd/JHvHGbKSRp3DOeUjZX+5kOrm62DGqQ1s3+tXJsZYJ5MTOfJYIUF0X9AZzKGFTEs
w0cykVdF2dZCgKqP3sFsBEQlInD0CP6FKCSx554wtETnqQMGYfLr3ZhhGLKlC0t0nUlfudI89Nny
53MTsz+2Zvo1fXIaSFfLB4wH5tabLw+1gxTSRrfvT0q31iRwWqZKZ+5I+FHsegsjO3aWnz4wP/Gc
mTQPJu4lk0UQGx7/GR/Fk6m2f4fFH4jxHMJwCwMH6AW3UCrkDybr6HtPOAdOuk1bd6ORUr7sCfaH
yE8GiSiaNsVNGegzeVyMA76bHIpq4ubXoGCXtlFkYwgNvTxzYR2+y15/D7ET4zk/sqCu4CtBT/Bs
vjDYbUD5h+AS3VyVcdJFjb5AOSMrDRi8b2WokGonghwh6V5R4lMAzVC9Bm0UzoBW5TrlUZv6JBJZ
ZD9I9+t8q5IUmOk49u96dhI9FXYq5LBCZDCdCLFqC9l8xLLNA3H1YNNHUyMpAz8vIIAGiBcNDeYI
WcBDIk1m+OBl5wJM/QIdWVKG5n8gFJG1IZJFNUkAR91qldVc+dvr+pPBCcBtrH2EmeD80t3/m/Rc
5Eq0GoBZ006RBwt9/NuLoJe99bE2eJtkHniseyYRQmAuTp8XKvNfjf7PJCmu5jAZiC08tj4h/qZk
CjqCTb0H/vamXaQ7byIUrbUMQxPsrsDm9Bd9ffSWzBb9GEjD3EKxdwOyvXV7/z1qOZzIgqr71Eys
RQAfkXuweHTlxO6Tmy5hGcVpGCiYT2HhPQGSx6Fea8gGKgwWfjRW22Mg7lW0k049EQInEdM+hair
3lTawcqIwzXKlkU3eleHl3dyyuMI6/oNy8SRCvR5JS27S0s2i83YqmwLUVcA4sFd82MfdNyBaFKa
IlvsnFo2S51rBwOCliix9HNwvxxH4IMw+bEWkgpy+jW5K3IlNcAL/jFNz9V+5/7+sEFcphcrEdXR
sjBFs1Me4BGRiWWR/IFtxxio6SD46dUXWRySNY1MQK0s53VcUnapowGNkDPSp9JT4+TcTCIibE7p
ENANN+QPO+ABcRs9MEazeEyyCyahfFZ9nemLBTPfL8Dbv3A0hWfnYhzywHG1/g6rr4ue1HcIu0OC
2t9/dePUWBCZRvDg3JKO8msZJ93VXq/aWFRvYxeHn3TWIeTorgu1RfxKzFOmVv55kB7Yseo9aXpa
8bCZaC+PfMC73DxvBgbevdM9pUS9I+XSRQ72ruLzGxW9NLEiVAsNlzNh39qdnCumcnTtVnYPBZGh
4JMLnwS2uwRhkgG6C6YNTmWVlwIuK7k3nd4wZRvuFqnXXPI+KoUyoyu8moX84fCMdBXMrOPkRvTG
Q05qS3EU/ldY7kK7JgwQN/layLzzgBVk61YSeNSmQL5hKZqb2fND+pPh1kWuJmclFWlw6i4/Bgoy
l+18z03TeVQkqJftxgvq7TSKlaR44Tjc0NApOQkw/TkvbsWdrW9I4cckg3tDVKa96p2eN9y9WiNq
VWPtx2zJgvmQ/4azzc/wBBFwVsHWkKEKMB8I8C5MUgCkKJR1Txk/q1S140GjuMIbbWHWqzId2exq
EOYxZDPfojz+XMez4Mx5fZeN5vMDyPTbrknddGp2vzxImB9asDRrZVQ+kLJVhNksvpls2oc41ajZ
KrOQT8nFKUR/68X1t5AnQr63tocpdWM5SW7xg0zI1gPk4Xd8sYajVWKp+k5dHCX01BeDff1C9NW6
e2oRWFV6v/PVvOK0ikobzoCjKk+DNSqsYvYAZYCj5+HrNRsO/g60VwQ/h15R2c25KTGVCiNpD09a
ICnzZtBBmVQgjgMMLtgXA4wmhv4I0NsgK2BJlWbJaqTXJLUdX5Pi6XlnVF0ZbsRcikI8hqk5+/Nr
7iypaRk+DcxWj4WwVtIXkz+VVIObAwQEiP14YRiy1/x7T6YFKWZ8T8i4u8Fnsb3gzuAQ2eHVOO3W
aNEVCsWZICOypiMCzcaJPUB29t7/7ajuE4fc9oI/p7BV2xltD4CQFwlJ98z0hFfWxPmg5kxIrEVl
jeuMKd73PdDt2Ue91NzTSPdlnbVZM7+/RDLPAkCMxGFtTDUqo364HlU4xK6qG/bOWQXbLq68X6Dj
AaaYOGU68ZQm13YPmcMhAO1q7+fOzEX7F/sAb5LlloqjePQIjzblBWvipIi7V9RWoSfqbcQUpUmO
ZZjg/+istA+AzfiqzEXlvK20EfEk1W2ZZTzfxeuG73NNqH3uW5zLX5ExjlAG6tbRAhicMm+cPr9p
TUVJwbHwNkNezQH7bPmkNkS/9TtnCZiELCAqINHWaRRvCVvsh9YuTGwJxmrKpEwTOdc9pokDS0Ha
GD1dZO1RoDKO1n/S1xORh/C08g3Uev4IXfVzl+KS99KitNN2YZ5xdr5ELH2DVTsruo0zg1t4nakO
BRMjMAispbfxY6H6s3FKkN7jBP9AqNP+6KZqv6ELNnRDUwVRrODEUBH0zgu75MmDgCmjI4EzoXW7
2vFikkkU14KKDyT09zHwG8CL2RQd0cwJa+pdysv1xQWGcw9ZCP/iqvAhlkZhee3MLSeULuPeUyu6
9KggcVPuWiM1Qqr594EZQxocP4uWCbhCNnSu31LeSR/eTKDDQm0aqKGBewVTF05bxOIeY0EPXxOi
zaY5gE7Ew7ejuodqfNXjcTYTzC7l1v42Z3e6NyeQw54VJjM2bRLysuvA859bhWo2bAmDce2gSzbp
pkv26uY0cgZhiJ67Hk6FUz7YWS6dDw60CJ2dYdlxtGi8UmhFsn143CxY5huqt3T+76CrfqVMcB5y
0c8o81vvFarfE/wwqzabd8NG3nmjgCl8Dv+PF+NFLi9mR4regBjox1ari1BCs7E2faIEscmHvkif
p+o2lxJSdyfubP54my9erwWnBCrtUz+yQRRo/danYknYd9hTj5lW0r19h2UkC2CgyfZmxItS0AQ6
OlbZhP7/fvb55p9KsSjdt2JTWyI+LwrziZe6oqZINqmvYmnThlR78/dCn8XFxS/2VyCGXR3WFw80
qAG5h4xriuMtWoxtlsBcHAhHvQoU59LzkVfZzLn63JK+7ptZSKo+Eyp/4f0GX0KoIHmLY3dk0epR
yR3Oc4QDN+piojo6Ds3AiFIlro0PFbj0A83ah6R2QlUzGle/sH4qZjmJ4XknyGcH/Rqt0SXLxs9g
x69AjKzA+P3Um2Vz21VTTVq9QPephK192MCkVWt1W7GwF42/TQM/adQt3rbqS1GIn8ts5/4+49pU
LRnzPtuQCTW9Du7RcgOmGQBD+5pzqJm+cKl9qS7e+74OptGL39s67DBoOx4qVjaQLMLLcJI2s1sw
w4ZZAOQtd14OLFbiSUYXdUtPAfcxnTjaRZqHscpuwy8qxw266wpTc7kYELA7UE7Pii08l6wmfIns
BTMTY4ghDbnByJGlDODzH9oPIR+4UHyQcL5+SirWweashBKUWFXZvAiKNbPFp/zNuY9FffxA3R1Y
Svby1+eXgeCPu35uF40gg6LxtIw5tc426b4qm9bXGYGI20HaKhfDs99V0QnNMtboDGEfj8+BRyHT
csix9jlt7s2i5SMqOzj55ewakQn47kf5kAVZdmvGFIPPlMYWyrRtpWqIQGmALAc3/nc1M2dSt0/L
TGXBOqL7ZTyzc4LxvfO7Ls82ikv5h/mzohyIBs6PR8aE6ZJacIaxTI2Z2QfIOeOzucfXjqe4Moir
yJ95fTSc04RafVMNoCjHQP+HmCfoCxg2+OycelNndC90NHsCBxL3B3unr9rlrwDQnB/YOFxwjlPa
lPIWFh97iXTH2x90bLkv9CI4gFcCBuDSrpTexd0tB4I301NTkpB16qroLl6/2fOEJ+jTKVwQqWdj
6VEpv5ED1aqs+rHN30EhnL62qCPGC8FB8aE/WpHS4p4tVpTt1zOgwUhKqy59oBX02ot7VPJrA6lx
VAxRioDysnZQdTsOP9Oj9EWJh1epLnAXmUZE2Dm3PAWariEUlY8MbStm7JNeG7IzBJeGys3AzgyD
KeQoKJl+78jIn7vbR0BXyd63BAv4vuOKTgivy6x32rvMyR3WCIAjcb9t10sUWijsHNMwBksRjaY0
spF0Sd9m0YflZhXxpkx7hpvkEDYXKH+QNcM2BTXotzrQJUTv/aJ58GcTCkG9r0AnT1fCCbbTy3Lg
vCOYSvt3lJAcd4tdOdd3vgORTdOwK8DXlW+PR+AFmBqgatCqQ7hRu0zob0vSIBvIS9H4lbFxi82G
qQcUWdr2h0NFzHQZTUTQfRoj3QE/5hp883/5VPIh2VmtH4ZixL4vpJ/NyOSqsvJsefGlI0B1bLrZ
EQPFLeRYGEH9JQ5oDbIGByLITI014ARpDvruB3GifgUleKnXeS66ZmKrRJC1led0ZFfPajFn7eY/
F4r6sGOSqH2ErIYM8opJDRAOBN7iafoY3KuITZhIQ/GRnwKpBUQoeiBCr66Q7c/kw0N8zSSf9VVr
H3MDB3mlNKXWegB6EpOYttqGbbnw1I3CbILQzSB8QIz+A0SvpAFQ3hCIuYsKqGi48shYf3REkeba
Y+kwNfoiU1dEiqtAQY84A+UXhQsofv/LS5QQJAQ3MXpkQPrKNu0qO0JfVZdsCXayK/ImbaAWto1B
fSMgCjCLWXpKTB7vCipjos5JE+1bdcIS5VpEjbjLG01koYeL01LIJAe2yRAcL5mMy6/RZmdF/81h
MOCIUPgWHag70+Yl4doLFw/N/7X6bw3nwvlshSrhTRj0XvF2y1JOwd5HwTqAqrNpWCkfheqlkuxA
0DTcWEr72zIIko/TnZqw86l5BJTWaH163FohrhdFGwpk0Zl0ZKcGymEq0W9F50Xy/KHDUg4qbFP2
miJAMgLGW4hFEEDhixDiCcCshTZIZpSCYP9vTCwiQGRJu4urRVsdRIdVFIio37OXD3MLHr2/wAOx
69l3NNH1BVxwtI2FZyWaJXFbdxWlD2XgHvJ2endgRKR294hEG67E1ZO0hRG1+zAPKrn9YrVSUpm8
LxQpdI8RPicXvdeo9LWaeHxHAeY0p0v8QCrgi6F0siqdzLfLrFHgf8ArHbCp4+pmbTNL8YeX90VL
E+btKb5+1kAqpMntFySgFhavPlU4+aSpnVHZT1bkXzc/gi7oiQEDmBI5IiHGEVAoLbiDE2454N02
5kdrOH0eYJargvkGuyrDk0EWlgwdAi9+F9yb4Uis1CEclfSjChsSB2uhL4b85KHY4cG6Jr5yzBQc
4I/K1zLm4eEjIWcuyB2tfLfqUQfd7g9Ihr//C1AoJmwongY1teMnqTAhaIljoyQvEWkFEC52S6wD
0UnOlupXxVlTcBI0RXITJxg/OefSDwiU1bOm3kwVgopu/2lFwT8+JshqPPXGr2lZn294fdpiSSH8
V62GRLLBCcEHPe4oS9RkL3mwIjL986AtU3GzTuVtC6JrVilA6uG5+Ep6Jj6XTAyZajlGm+UHGzh0
76kcvbAu+KKzuXtzVq8M37Jg2ry9U52mTJy/USBlNCxKpcw5qHZjAnw4bkIiReVUgUI3nsyJNuJS
iRIsujH+g7BELEAj2sdjrWqVhchNIJ5uE1G/bnF2BVqHOaUi/2TO1OoXiVn85SltLBKzoViBpQO7
yskZ1RDf89dbd+uXoiB+oHkotBSz6B7XCnwtYWBsCkzz15j0Y2thIRYf+acwyFsy3CBZLPpjqrbP
Nd76IjfhI5n6yJLcPYPzzI2Amqq6NQo/P/Ldllf119QpetmYrV2NL9I3jnuK8e7WVyFq/EBqp8Fe
Bxsir+EdSYivizRv3hqGL5D5TUSvfK2EwOcD5kEU4pKgrmOMbZDjrM7PGzcSyIpMbng5ApzWOrGZ
qk8R3hDkCp+5cFAalCH0DU6LkMPN+cPfJ+UB6UtP8rco4czaNT8AZmMSSVMCVPAJX1xo3V3f/tsk
hZANgIHOLJ9734tes8WzZZrITdqvGRvG4mYe1UNl6jFKMWJ29HOWmbkXQeKYdXDrXiAT12iHrTVX
LUztQ5OElwL87LACdwchCKxHhV8roeVLJTuRbbEufQdSwMvhmvOFe9YYLSJ8MCLSZ/EB4O7iI99/
xJboXx3tmv0jQRizYJHH34kWzff9DqEO2ZAWJ5dLTnvAPGiZoIsM22lFWmE2siR2oCE8vr1YlK0/
bbVUslXruc6LyV0BXHodY6rHod32mL8OXUHEEVtv+zqEzsaVdg2S7SSwkCWfeWcrpXNj72h2t/nu
dC0o9scAF3XQoZ5De9vy9FwQthOOlu/8mxM3NS3d27wsRhRPUAFDBBhCvzhUYq7IDO4we9W2whtc
05xqQ1vTOqEe53fpJy3/F3GSfJdWqBQImUa7hbkr95OJeN08Fpt0SG4+g75KL+C/rri1KhoTOqkc
QmfE3+xB3y8/PUl7Xspz4+YEnuiMXS3Jm5qAg2bR/dtshOYKghx1ln+YDLTpwtVbWS2v5i2qo1KV
durMXyRTHfF2mIfdFPAIJ5bYIfb7IEDkasnAK37GNNFBFR2dWXQkBqdC+1PUxGq7aMWY0o2ZGpJm
vzH0llRh45erKiDjrt640DnQ1t21BSdI6ZsMPZbA/KmJtLVrFT4OHzRUDMQNwKfekyEDmYDJmBdt
hzBdd9FvgaY80qxWq+hTJZI6k+baJenz8eoqTkdfKpBV0zBHwVeJkVwAR2C8rev2JL9bUGbeUkWO
7u/NAj+t5HIn77n2ZOCipF9RazXYvPP1KDydgwyMUTdFxrjl2aIuTsIQWLTJaxvBgIW2sPc5LXp7
mTVq/x451R5Gfj6xikp2wx+yMN5CtrokApC2vUrhOaIesFn7CjCxC6N+E0G8ulnU37yeAuOWAytz
jBCH3AMy0p+GvEAf7dr6sQ2/HUJiCoJ3yqCuIzNbeYQlrtDe5G9QDyXv2HVqieWxA9/hEPX/4EFQ
FwyPxUvfwZbEh0APvq/p0kBTjb7swR/OipuQ4SG3Hv/CA5Xcw1I/BW1UYT5wSsiuBpGUprx1MRjC
K/3Hz+QzH8fvtczzO4lIr0tsHFSxM4LHShSrcULPjbyxQVnjfuGE6Mui71lSL03Y38EiLmwV+7mV
QpydwYDdOzq9bn8P7VR38KgkF2bUHpeH9a5Ww5YwUYsUInSSARLcY3dlyqlKOMeE8oy9iMHgzMDj
pI9EmwwYnPmDg0u5bSTbJVAdgGqz6mSN8/e66Toe6Tu54Y79MJ3FI2l/elNg8RSY3yGsXxhQOjKX
zQ5JBMyr4GWDYaXPj1Tu8V09tIFnQLtL7QIfhVrTkWLz3mOgSsD4w2JTwp0/XM2IED7QV/y03q3C
kIqnL8C2oPWvf/cLTWPQQefrwq+LdUHst6j7fbytDKFDOkkVIxwpu5oh8V8AY84zArJimIJqpacW
8CKXoGsBmhUMHIF3uuxvM1k3Wzcqp3XI3E2EkVNuN0ybLhu9uBxwFeRznzNSpSE7+C4L525+GSde
Yr7aJIwUgU0ehuZTawJYOYAGVWLZakocCCMvOVdGHvTjhJgs8a3nPA9pHmvU0lNdDJUb/FbF0J0N
BgXoMLJnPZ79WKzdWPTSfMKvtAm6QerCUX5hcCgh6XVR9VYosMKf32lf7ptWsKBrhqren+5HZFC3
sxypwxAxu1CmQfVNj62BbruNJ/GvLdlwUZlrbJOL7vCWYLS2rB2CSPPE4BW3cShC7VE9gzQJu3Uq
YGqIm8aK0LDAkfMRmAEn9x52DUsUSZr9m58Iob85wCSNQhvRrl4zi7XSzKTFq6foK8Y2dQUsMsZw
dgEumLSkiAukF7ad1bT48NgWvDALcmU0H3Nmdg5rsnTj12atizfUJm3EApO/y9CkAAi3hEOhz7Cr
7aomnYbkl6HnxX+BsvW7/AUL4ZNQgo/PjUDlbgaxnNQuzO2i4MCI19JAeQguPkTaES02rPN1G5K7
+Z/RKl3Lth28HFPrHXr4jNrxWbjEoKfSxJKGDJi0iX+WhWObMQypevi5V+vfHfUpFuzmA15XSWEN
4QhTTLCVUVEaYxPQioBtkVi9I5VUjnguV19vidP8BS4jvMbWGnrvoZTr97FnuXTegG0Cyj1kfyaQ
2obsvSUMtHh8y5QOvFwkhF/LlXB87afZQYV0c6qFP8IncbfsTOEdym8RuhFItURZETcDgUz6MPui
PtSbHFQ3MtT/Z45LKKm9C11QnWIrzt9H6QWg7ltDQvpdShfBpRPVXXCEV0oz8uTM9UNIGf2pDwn3
ZftG9CWDCl3u13MW1Y3ZR9NJAV2K4MYhGoCakuvSfnXYbZkwvmVknNQLg9ptIgsULYpWs6XFz7Lj
GIl0cZuO05BYl4m2918cD7kepcFTqj4WH1wqWOU7b/BAcOMSxNJvmufzqt+xVYSbbhFyp/0HhWDo
o2tYkU3lnaw0MTaEvFqHe9IEQZkjYY2Xt0OUpSZFoV29iVOVps6uvkCWWHss4lGxPICvTlGdsAGR
4mZhoKEKCMh29xNIqHQyCWKE9H22Z2Y1wcn9snlRgkYjefQxptXt31X9w1ryvSQKqb34KRs6ddxX
NbHXpkgjq1XwfUISeP7jFcCZuRdFx74E3DQX0HoXbMXcj2VDENgYrCd5G96LRFevBzKnbEZmhCM6
bDJ1SET55K+6o9p8XXVZdj9OnEiCMCu6aLXeUvmq98MyPMWE5yLb94ye2xECPGOFfDZuU3ojqDKW
q3IpFzM6sM15NF9RkblwJ6edr6I9lV4+Cymzp+d9ZhfcGJ33LxHdoCfPcrLxtQ7yOf00FYefKlHt
iw/5LKy1Y0fwDK9xwiUvsdS94DguK7eotL03C+nX3SS2MoE6kZ8LkvZmtrgZiyYTZCQov9N3TGUF
abay+ngnWq17EUoKyCwOLGHyL9cnGHV56DELYW9+05zDq5HyTwtFHvClpf0kqkPU1N3zntDllZHd
IEPT4YJQQIb7xhDdX32M5gbKi1My4G7vo+mXx+o3nRaPFztppET0FxzRwwxA2e3fnnUZ8EG6Xh70
1pKacdYlUwTsAT3vMbWb7OyfUes1FYBGYB21OkJ5OYPzqgm28wKw/RHlTAUXlN/G5edGnH/sCeCx
EzwzgIxNEGfjSg90Pvl5QC24bWcYFRpNE/1ui8Jcsamz2x6TvODpgZVrsBb1m2ePlDfTa387h7EC
HV7w/aDspDJXAi6+qQSf664q081OU7iYjy6wAqpFgmPAg6qcf9aCw4XbUYjlTDkOK2EOGuDMEiTC
50S2SjDSpHJ0wnUC4F4L/PdExmz7ZN7KKxFsXBE3PJH9IbTwkofoTZe9KN2S02u+ooeKM8OViFvJ
gUxCIZ3/uwIIAwJxoLfgGj6vCeRC79gcrRrsMj64ZTvDsrsrRpmD9OvQvfTMaHg/ZJVFhEY/jSzB
sFJnlTpMGO0M5xRaEVMpDCfBSF8OhMF/cS/pg/JhqxefcHz4uNkWnS6ION3FSl3w6JHdxB1DTsw6
Moin9d9xV8jf8QVkTOWrjOyNkTV+TVJOxrZ5WfYjycVcGUMDwoyqtQqfLAmZe0tV3Ftyw946o7dY
/wfvb4Dx+bu2SxEPP30+YNBRrcVMEjHLU79sIAGYTUIsSd/4CTKdJ20aKyykC9FdGMaKUkEcFfLG
CjiUrWbf2MH+Mn6g6QNtfmFbTMUa5t/b0ThzvE19SULi23EDZv+k2mnEuR9hnEtApNde3Ykn7e20
oC4zuHUgmPZLgsWhh6VwQgh5rc0A4tQZu7C3MtMbuUBjvnuTH5dZK2mLih9PBaQuH5F0yh8P5PKd
nYV5ZUE4yokUOJdJCE04TVU7aSCx9mAHJXKvaGOZa3nSkNR2pZl0oi3gMzGLRJNXSWAPYqX51B1l
tS1nB4V6UgBFkm40uxFqeDzR8/umrYOT1NknN+i8YNY5GIN6ROVXrwCAD6uBevLmGRERzmpevOoD
Lk+JqQ/4d9haBRTtK4TUwGsHxFqoOhyac6THMWlH4ujNlBpxQULzDGEHNNd/6szR5kcxB0DJpk2Q
pCabR0Wgfi5+DOOgtWPZQZzVymJDaRYVtLCnfZB8Ix4SjNMQrkKLcKlAzmCERI8PMecUVD01y9bb
XUspGvW9vAOIXn9xSxxzI3wN5cLGcLF4lNBoKj9L3NBK3C+5p+QNQ3KIU7oiRegr+aAguHjIkjAh
t8L/0YJO+r5TBSj5hiJ8BIFI8VGMmew0KzuQgj0BhUYpl06rRjjM3X755u1QQP5brDv3ATaL11oZ
oIvxVbqiwDxkgVHvq+qyObfBub9yHL0XW0g3b8J9LfmwnCfxcD1KJWdPYLm4iEhsWIDyeWUAevMf
eGojTpTYWqSuYFZdEO1I+wV2gaIsicQsvdyrh89FyNhrH7FitPaX9Dl1qVQGcj4ThY03DWqL5s28
e3vnPRwSs4rQX+DFpjyh5MDT6pYq3bfR/KdOIVf9I8EZr0JnR48K2h6FIeZSxBcr3s9pLValjsZ7
8xKZloyHrVISFpdtVeAd2Y+gc1rcFpKyyzuAco5GOCGA4HHH6oUsTgr8tvHGGeFpi5UFNGs84y/P
Rj+wIrCcPmB9gJ6xixqggMFzFWVutXwQjL52dnQ9ZRVjerOdHWpSwUlIclvt/J7dafU62z4TQNPq
bHI0Cb8GRZhabN4qDGHUEUz5yZ7chaBNSJO6ftNFmt5q3gQe8saZVgusS5C3Ny871/XkvxziSnJZ
pbOg+hj72AOGKwx+pNSpOvGYtKxktjAJbOm47kO54gJkk4qYXo+MJEl4UJ/49EvR+ZN3o2l2WxuL
6oCKPndzbtfhMfyqz+Ij+nZueAzkWen/+EyoP432lD/ii2jWQI6M7sx9rQ03WDqC3xH9me8O9TUy
SE28aqxtxcA8B4TnZOpj1XRFcuhqiElnzFu/6WGWWXh9ten+aw6gXMhZ5+9EYWp2NMkMmeUuIfyM
IxGVKypeYYgOFcmqG9M5sTmg1BUlILy2KwgkfD/zN+TUwI2e9WHlT6Yv8qEK3sJ6+6mf4cOb0q+s
KnZ/ESsq/i89w7/bxxsleH28/MI032VinF4NJ+7roagP95mK9o2jyUyZhJFQBmACVBiwQ5e4hNff
HgbNjuYZv0qxLNoonljDyAUYme1Xj+KbSZ4yiAXyrN3ISAC36ccWPvQLETyYE92QneG5F09ruOL+
uztqJMyuLxH37OH2z/AfL+hayhbb8mq6c/kP5Xd0PlA2yME5xd3rYEE6LmF3Horw7qAQ0RNgpmuv
wy9/ommyaU6hK4yUXPrlqVPEW28kyFM9f8us+o33Hn4PnSfwakEXmeQboKPfCOXyEvhEo16yTiGB
k6c8v8RhIGLC7yiVQ5W6zqEHhdo5NZQVZAX4L2/qxs8YQLReedT0tJTAYbHNfZXY5nUivGIFdXiv
O7R8hRI/5DqY3e0rvnWc+FPTC15260r5afC65tXMxQT9TjkLKCTcQ9x6ldWJcnkLLWMS07w5j+pu
T/JXZmgmeJ+ERmfSNnHxUHuUd8AI4h9CsfSIfx08lzOd+oGlNxS3a5WN/dTw7q3EXowwlz/PQwSJ
wbnbmzX77wLR2vaHv2SV6rJk/ToJ0ifkzjvjpoNvZogGP5Xtd62Xf/OborZ6jtmId6iZwoWEOGtt
5LoUntHOZRYmuVhLfD560c2/i97OeLVAtmOFLC49qyvJQSUrLA4hsIW+3zUfZlzMMIPNTZAytAzl
CkxSpPQJghWYj510dbFCWqOY9UngvAuB4PNRc68aEjlJ9SRFsxnCVt66ZXtDLdC+pBhdpDEGwTLn
Xjln9OIbJ9defYpMdeOaoWcYrDZCJb3jCbODdPXZ4gBf2pKMZz2+dmRh+LLX490iwuSA4N7K5PZv
0QHoYEIjXFl+H8ff8LCd45kA3og6jbH4k5e4gjcdy1IL+IFDw2470WsVbgkK+o8Z03Eu4TmHQz/2
Tb+Magaif0aU/z9EhcOMCnqzRRActdft8BD1glc5/4QbriXLM3hhAXsRlpcybXTXvjSsSIbox0PQ
2IVIPNJI35Pw40CqnlFlruycl7YJvVnQnXGCMJB9ofrFcJzdWr1gXtMeEs2AXZrT/0oF4FpUg7Bp
uIkTl1VoceEUXiaXAvzrEH1EmcqSosoZOVE+sTH+CXFw7pns/qwCPHeGj7ztoxWOJPxFnC1YdfOS
iknjvfvk+/brFnzifvTMdJCPt97bLY9jOnij3ax1bbl9rSKjsx/MjFI3X4O3S4cj66JPSVK3izBI
21qEn14N2tZSGp1JfkNdAEPlT1FOPP8F+dwHG5CtPE2Zdw80+ov8fdFmttB40jU4sklvSwFyNLDT
S/IoYNWA0Ivr9MDqN9vCMcyV/HmJeU+BqIbYq+1gHApBfgaudYyVTBLWOtM3nQuUXRV36MYYY+Bx
sMd6xfHKUaWlnVZzSC2EqfRcsVnelmyoiLvKQb+RwnQc7/d8PLERcxPDvHcCXFfDdxKNdPSZT7MD
fnD0bFdSgyiE4LwoTqDlfO6xtFl7wjLcTOcoAnb6o5q5LedELkubTs4ZK4a6V0+8Iqv3ggHk+Khn
jzywiCcFriq9AXXdxUQF/0NaNFVDu/LHojqNvs/GCGvKpmvBwQPOwUD079h72w/TuUZnYlnIqR/V
ZF3VLPZy7BUgTd+EPP4T92p8NdooVhCJelgLxdfp9XuUywmqjbAFvjZ/crKwgdjknkGUtz/pmO40
b60bmRpyhlHJzwHfao3f1MV5F/oHaz6mrrpDosPMIVaFIQBnf5zx+OpVqDRY4Vei1nZ0h/FvTnFM
sqfC84W7iOrKlOvrmdsKZGE4rdwVy0a/sZJEucfA/ZR7nW85WloRNbdBVVgGE3lz4EzeOoGEkXeE
C3g241sMfidEUgMFZcHaseeGXA3QHvVAauPjLF875AWRTNQy2f4rdif1rPkwS+mrnYtg69NusfNk
HIdqKUg1vtEtJiEugoYIZ13mDx+frgDnGt5BmWo28rwnQWZQW33aZ8urjIRozjoA62w9UgM/r72N
nkAi10Wk/4iiNq7PDV3PeXCY8tzfa6elmEWixwnWO4eivbpnZh8ggXn8vKdBw5uS7zxFrx5uYo1G
30xwhJcdaNrUBsjdIix7kAawnivF8DLKAUm+CseYyd1wQL+VWNah6yiPtJSHCqDEK0ki/XMbRGEy
UgKBELtaMfZXoOfcQxc4hMUgguWsmxh2F5A4moXfUOFMbBgK7fLJsbatvN3qQ6zUTFfaQzN4anHw
rBf+CpYa+o2g7YLkO+rucDWTEnGpCckSFBynt0bJK4k4PKIi96paFbnp+FnT+GEiioBhPGm6TbUr
6Py5Fx6UZd0d2YOFikoBeJKk6r3acx8vvt7WrotSowXAW7STI7jPoOosI9FaYBWlo4lHlUr4chyL
qJuaWxQE72B26aric+8We0WXoNRSxYIQ0juwwKsM6lQd+c2uRb1TOEFS6uBQJyM55fPU4B6+q4wi
M4sZ0ifNv2q8lzsIJ43WZ6zNcTaRIesREximhPBntZFpH1RW8RMHq9kBko5PwUgRITYN4vqEXjlf
JRPaVNJsRRmLciGJU7t60+K+awaucNiGTa4CifaPWfzPspMHmKsOwOkiyEfif7589AB41lekDd1N
f1Z3X3U4A3V5qKQNcavk7rmHHrCIFAxyo3/+N/h5l6Ycg3Fytlc1mk61FMH4K0GCdn0D0fiDsQAt
dkMB0nK/z4pKGhjouuECRJfTo1JrkeQ/LobT3VQgnALMOIkGqWLaChvHL4vOY/Z4StI9lOxHIyrZ
hsrwqhqXQPbyodvn0KjP8tdkLyi1aEWD9SHvS8O4YbvoqmDWLhYfPMgPuAFotxt+vLYWpf3Stkki
GcDNVRxKSb5Sr8yW6GH2UsmEGihK+YByiAncX6bxv7750unOoWKWXnp05RaFxB1b2gw1Q2KWdLz4
dYjusM2QmwP7CLbFZzp4oz3VpQIFzjOWxlE4RU6GuyD3ulwnQVC5vDNbItPDeshLeMQf9wrUvRI1
4re3cOy94NNNy4ZoI69sSI9vhvMZnjqcJVlHNRFF95wXKe7wK6f88Vlk8qsrEqkp4vNlwmuNujBM
MzRQ4lP0TKqcoVGP+koX57nVKAqMjpD7GYYC0yAwyMRX1jXSqeNsXdTCRbFOiXpFAP3YeNLWxyv4
2hYc+esYbXqZuNuIaPApEQlhujGKI6VIDOuM9LJ+Kfmwfkft5xBL8yyrWO6jsF5uLrS7ueljYzWO
ElQ8NI7YXtb3z5PwwejCBQmYJ3aFQhQnyrlEbsV/HnpuA+Ax6ay4v4B+pVSv8mKHGwVut/MyW0TN
K+y9QrbryVh1bk1UyHRPW9dNK6S499/UKi3qjcUL1UD7RgK6aTrhKcdMhvTLshWVkJvgcJTlHX6j
c9IjvIJ5Nu01cNnlShn9XrW2GbtHmcTKhMbfiRQWEf7HgEc06bUolYD0FwgUn49JZRZ6JapYKXHL
0y4ag/Eweyi1H93Z23W6kdeYFD6U/0506CXCC1gSS5raVHASBqkmx+zJuyQff5Vd/3sWG+g2NS0C
eb6leOjJtFP3jG4wqaKCj/jQTqUm+wuujP58paMNP4o5kF2xSxuj4SZg/xMLDlBxJ6N7pe7e4X6c
dNZaAevtu1Gco9umLxv7H5BQB9iww2sN9Y3M7ePLWrcMLlmCP3WXptsZbLY9HlSHRtmu7L7DSm0p
C+nrzl3qRUFXeXdOpS/JwM6xEvDu9c8rRP3720TzmrruzTWoqoEBYC7OoeBEUd1eM1rUVqEdcPey
FxOpta9yEexyElhQw0NNTdorrCj3s8ALIVPHJyZpR0sYYy3iMXcwB7dnxBTRT5PCy7Z9ZF1O/ywq
6nKG4e+3fbLIen9h8s5QOUF+pNUK33LmJNiXJ/kHxppW3PcriIiVVw7xB/NlMbVMPLH8MPK1XKda
wpBwQtr53FrisJogqyQGGTXv8d6rwfQJ74M3kLnxTRxaRi/KQzcXwVSth3hc1SOn82LlEKE/zGtC
8y7I8HAUFau2zsDh2QKJe05tdiVEQtuBOoIFF3FSa8RMnn/NOmIDjwx6HBP/2w+PuxAppQqFKfPq
hXO6HtQqN7lRe8GJfSyHKUU/lkaP7Lbw0M5sjArIrORwsUSUUXHVYfXkHG84bfapdcXyBI57j5RJ
vqvTZqZ4cFy2irOd6ywbrRpXi9VgA3VQgu2Aq5tejWPGraePMLCCzWS6zq6HgfHMGRGVQgfS0Lt6
PLpnalVe7S8TRsF/e6kcWGWwxwAi0Z5SGZ01sUhE720eGzJ6qRpYXXvOePWe9NOP6jqhHU5u76Ka
o0KtMdUAdJnXSdfineKJQjTsjrE6ZVoDXL/kG4S3puACrQhwRU8j8tIuv+vhPBRNd94G5Je3e9JE
kDNg6oKDqDBYgRMHgjDInQoo7GQHg+pevKKZwSeNpGKy0o9prXIP6kx/Df9fsD0IHk9+CL3236aH
iFgtGRrzQaZGUXX0N1s+d0BsqE997MRbz0m9+7i7HQttEcwPh0dnaTZmJiNKqpPf0r77Xat6crVw
5xQTwPmhvR4YNFXQ2XgAKwxGAfYdtGYdDeVF4/biGJG1o6VT6i7KyhHC+gOz5OHNDCpzRRtJcR+f
VkpM4LRh1lpL7YWWq1yu/JgdP4Cnh6OTrEaeY7z3KLdqJLO6pmNmSH2qNz48DSB8smTmCY6i81i9
tKKrVp50ccfuEoY7axtP9aZgow8j/LUQubgWPn7an2LsmyLjRNQQ7URZdfRMI1S2+8+Icn/UcIrJ
u0ThTNRmgkoFcMZR1ZhP4kokopownnsiEi3XGOoBI7uFm6ZrNvk7itecmIDdDSN+aIah5KkC6XMe
10wVi3OYWUJJxVH0K/4jyJMqenfDewtot00Hjr9LH622JEVvp6JaPg4adFHE8r/5XXYFOEEgxj6M
gZhgxsXnAb/XxlhPMP4GCtgWtxubhcEOSW/H+TAPyMCYXmxIz6qNGWsffNb3PNFvTgHI+qbfGdlS
6kICKnJrVPv999tr0p2xrj9s0t90j073xl82FZAi/VZcVKSgSAlGzfJ5WMgdUkXDDn2lvaVdsIKZ
aTJh5CMVolkipWlkw8TgGhud7UHvFB5u1iU6Kyu3ur51NL6ALXhnwWzmr6hpuYVS7w7D0Zo37WD9
a+QsJ2Q041znNnPLfTZlTzIGWjJp6uTSBqknRsjMMgBRqxaOgwfKXgrzgUhg657mb90uxQ+XmgDZ
Mz0z1zTxOYEj+7JUr7jlFxv/5HWSSu6AuIWaObGRJi8SlWQAst3+PRcl+eJcb8xzSFDDTMT955aH
Lbv1u89m8UOThAe4CitxBIVBc+sH+TtZ0Uz3JvHdZ0KvDP9mE7KC7DHt7NO92Ln/bBHDwvmupbkX
6YhIfCoDK/DPkyhOgX2fOLuoWBmZTPkWTd9N0RbZC+5JWTD8/bsIJ0ssZ7aMEIh3PS3EWQhibVe0
bOBBtSOHb0tv9x8rWVz5rygmT1AA6CwgfQWc0tQq4bER1UOZ0XlDiUN5M+0oOPBOUG95X97rXBzD
Hn5t3xXVVr3da/3z6T23uysJDL3Md9/4bNYM3Pmkn9dFbcRV5/HEy3ATRzJ318I3quThj1WhnNDf
6TfLvwJgC2Hzgt7cCwiuYu2LXYgiZrbmQ0q++UxjnrpxfkSLjJc+67Ov1v33g72D0ROI+uLxBVQr
+bZMJQ40Zi+9wM5V+bvwran9BQ6Jk/CJh+cIIWNnqckKcBcSNM35shB5V3yWOpG0GCHVyNQmQO0w
tg2xIolUZuQlXjczB8i27I8USkIUyO6rCEmoYfUkV37gPoTiebTzD5eywt8nIpw89UXwxMTLYiLn
MGQ56HcQIJrmwPpt9kr7RiPFQ4H9qJ1ZdfLms1q/shb7I7UT+eoGvx7AOEWz8Cm4d8L8f6UVYSNz
lZD4QNK8aeTxANBaZIjcH6Cr3mza66HV6hzvSLqSE4YSlsEls33Z7dOd/qIJmaYc9ihefS+4WGH8
vZBDmSbpVYpxmvDrNxwLeY9QT4+ZZMReLHMEuuMyHHlT08uFqBH09i3b4lMNi3AM9pZNipmUKtYs
ySDIhxctmYMSsmLNDMyfDt6+5uUzcMv+1Pl+qadwBZMybxnq/9G9HNDNDYHJO+dVgOH1gp79Rf4d
j9UkGjzScKsxYXxCyKK7JSbmtTGkL0Dmh/LGHpBREt5NScggBBEnyJPRrqrZKKpIyNe2AT9VyqmJ
bQscKFiJJUsG8SFDZ4OD92MjTmjVYQ6kVrbt0bhFwtJsurmAhZBBetMKD6uNkilu265hSoLcSUD5
zIT0VGeefCkobSRVsXuzAV+RESsH68v9Mm+OReyhqsoYu4E8JDJOIM36bf9f8HteWNmqEn6l7jtZ
c3kGZbWjSFKX0j7G4wQkHfz13FcSSu1vafUs6RNUMRtvfSBAskbw0n9N2iJalY4kPUGjovMywCK9
Kop08llCIIFPv4KVitfgzwPCTMQCQw3vGwRU6ehxYLDnV7pF/ZRB8806sp0BIDa51pkLYCy/kqEm
d1r//NkKOBfc229EPTg7pq7FhGWVU4Urd68d/MWKkVvKtGBw5MrRGqx4itTpQ6d0ASHOeEekjh4K
+RvYDB2A/SkOVJbMKmcLfLcFrHNZtaVMnFmTbXP0r8QsMdDC8K2nMPrpKfled9b9LxX/JCTisfT6
PfWWsOdN3dmVJkpK34HhA9dwJug+k3RgLb4oGunY/hI9VA8RXXavKHSHhq0/UD+iQNEwF3p9I6gf
V8RcreGM43Jinp35B6ewMJvjUDMECoM7/yp+unSg/Ee37ey1CHUsQKnMtipw1WXUNGvUYUZq3c91
Bzq1Om3YCunE28KMUWGnqyc0MGpW23EwxX1em6qCZ90POcVYiodSuWOZRDcn5FCXe5cT8f0fXp+u
Co8PNbmYk+f3SxWRJq1gk6aPU1ABMkNbbjpoRmfIlWT+LKU+tsCPGj9wunv7aJdKMNrsW1T9mcff
NliIqc5DUvfCBAgpxfzVIldKEDK6l4DlbjVnWblRazBWiXEzdyq+agXf2oSjnAptJrdGg7Bsg4k7
hMf1cNV6v8U2AZTb2FgO/kwYNCKCoq/bsPJMx85KQawjo223rjTUoXxqa9xQtqLbPg6DMVNQ8fAQ
ZisD7Bbi+ALhDeQW4jImgP621vwHKExgaETHHNtwYTy0JZ3KEODdZxGBeFzKpFYjG5rR96j83NmN
t3UPkRio7GQaj2i2TuETQRzHpXxXkzPy/WcmoP1CHO2CRS4yGa9bJ5ZgPATxiCrxQns8pZQ8/IzL
TEtV6wn9gza8V55ZkJiu26/UY1jLdP3KAQr8qdYAtS5pwCST91ZOC6Qheruq4x9tr7M3CceoR3Mm
A7S04K0bKMmxIUEWyIF93fneyzjwsO58Hqu9fNlhsxMinFbVr8YxBOyEMimC2OjhjWxdt6CucZ3c
WmoQEMMmHsTQz0uWV/9v/Uv758kqygp6r5o9y1Z0akuPSl1bt4g3joHnxd2an+VKYcUg/sB3oGSZ
Ou0XF+rU2GFP42cdhmJX9jL1GQQeHAipDmqHH/ulWdD0k2eqLBlH4KQ+ocQFgIx6JngmzEi7ZUYO
BFs+J1z0wBowva0SiB98cnMwaUABKUp3/Pn5YgPZPTt/5wM2tluD+hQMayPvQPM09kYHdMaglIb4
YqXfTrej5I0wQWa3gQPb+2ZUXbb4dndOJStvA3blkUWDALrOvyJjzQmm5K674wzbT2HlEZaZ/ZUi
mbvzmdLdH0O2vwLZMKb/pugwJUogOT8xbqlKLfKSLX6YzyRqfLU72P2X4beXYg5HxO0bzzubDcAK
oT3/Gwq870+R1BZ4xq35EsTh6Mj9ioyDb+RFHYG2pIK9rqQL7jBzw6nRV2zAu9+21UAlgxrkm7Ak
AMX9caK9qMzD5Jw/WY8wnTF5DHGvHBVk26RU/uuVpR55n9b2JlxushTF8UHW4SBhiB5K6iez/YYl
DTtaSjfYZyKQFKXfz0AFkJBn/5I1HH1E4JFsXg8PKhFdGArTfiF2z6uKUzKj9AwAiaqwu+8hPeVp
jIuOiM46JQBAr34qM4GLSzMHuog5u2TmARrBP4d2z/RJ24ok7C0HUs0KoQ0+lmWhoGRCXPXJIAQB
hHUkPaKsfm3tpoYw28Wryy8YWy7Ylk+iL+RvMi4bNsaDngA67qJSy0E3PwNN1laCK8THKmVRr6Yd
gEPyCEe68hpQC1nyyVbHczzYUOQwMEVs8RmY9P3mSCV4WFFDqKIM2RVzMPbX2CAonVm2rPzkr3eO
0XHwMs09kxznlZcc86Z4dtuKeatn9aJ06h3AxoX80rBz5ka4s0MNbV1kUQgeUKB/1uq8LRHwahbn
VVqutOXC5vuHeIyj1oImjc7kUW1xHZXILRRW9wMBsqJgjATArUYj21jMS4S7JX7WqBJw9Sk3fJQ3
fNdy9nZVzgH5ZXAKVN/4oIOqDxQC2fpiKgRIfj7gDcfoUPExFPmJt/MHpCQVQCesNRrxKw384R8Z
BTafpxRS9+zkWRpmqRtfq4yHbdsPq2ja5WTrh1siyG5tTI0rgVuiGzpDlz7smf3HsCc5t8YH3aqA
/0hY2ewZIllPX0Y+OVBnDR0sj/LmWcfRhj29hNDUicOByH6WqqGELIicS07Qi+Sz2mlStFLAUoWu
KOEorPFzvvYNl77GYo9zVqsqLtRsaIVoMyAtswqZKcGsV3lfCcky6BKHRBFhw7lByNHyY5dIhu/x
9i1Zm4fIGULuIHac3ol5r+DE1J5k0M7JXQTCL+Pzaw8rY9u7fySYksrxO/nR8WL494DP5/psQL74
N7xP4zYgNHoFkDVaj58YLhUNoMHatVNJEMnBSDT5fNYXzIpLYszovkpUIoujVNFL2OG4WHa6qAnF
19UBem5mSxu+N+Rl9fJWeKOJkCcbFBnhy70gnrbStLhQYfiuUA4RKMB05+FUdKugqEu2xTJdBtF0
6rh6OsQ2ruKdXyScXA3qdef6NzurlDU7C8u2ExbCK/pFdpZAa1CHYlCx9jL7+kjSQFVFJjCNccyi
CqJeix97yL5OWajghPG46kAEI8Eb81nd42WfQBKKnKZr0DVZ0vtsMbhQYdfGBvjm3ikbthH/jBH/
AjLv5acMdVjsDrwR1huEYFYUnvHzk22Zbak0gqbx9qgdqvYg0EAgS5g9mbcZmNrJKOBhYvmjQGca
1nIoM67sQdlmVB5Jw4PdM7Dlhq6egKoqu+VJcsgdPJJtgFq0l9Jb7k0FfXniJ3IN4mP8Qpm0cOwv
HPVwGH7Gkfr/wGi34021MYuQv5RZQqe72DWhgYIz0OtOprPwTg1hbpHYa7RjEdyUs3bvpTi97U0L
JZC/p1WzO5kTkH+u00lIF7gS6D7lVhu8ezQTQ8PDdqrehrUquVFNfwZWxTEeUcm0D1k+BU8Pbn+q
eesutZ1jBbs4frDt6xa27SmEcZbgAn9OR0L/0VQXZNMVgzUwzL25gAgccjEf0u31k6Wj8AHJ/3g7
zG2DfdhVeIHM4TtvAWhtB9H2Ggu7LKVmgYzGVvxMNFrR/6e94gw3XfLDc+7OblljO8m01zDXR/wG
B2fm1K1xp91f7pmEsHnKCF0Ayd2yBd9IwETh8DIy22q+2GEsEFkCvy9T1H+H+pte9fPiu0bXnjPn
4vGlEuy7TJUsuUPCzEPAawb5gvDG9wVH45s15yUQHKERA4WeiHwrdJT824ddvhkpwUJA1hegOlI7
+D2OrL7jpmq8ZxvHuisiUsHHM7I7jgU7iGyyuyuPdazgYvJ63hW6Z21u8AAFOPT605UQDlND67Oo
dANJMO4pDEqP+77VbVx1mwYNG7RfJVgaFvtKAvdRD1uI6fgtRzAIPupZvxCWe/SCQ3byHJ0YCtY2
am2enqHyH+kKdsJ5VOd8QVovQEKcu0WNkN8o2qjqGwQDXJcyMCHdAbhcpnFLWD3jnEeoefs26bDt
fN+sxB+mmDM1S85JO01RHZi1jdeoUX64sOU3nzUPWKRNKFWkn3R7SKf0swWjPKzjaQfrdf3mLPBD
V2aatRCIo+xzqAgF74wV9wnTKg36lZjapzS0/JdjFmnvFxvdxbTjTAvnVfLiy9FLohRn+kRsTpha
tuyVzvJQYUakgHxRVYqh0vI14WM0dk6tDiNa5wRXqKaPhqcFC7xXe7avZpHFrbniqV+oZBatuEJb
8SbK0EPpXupqqPUOIvYA2lIMaeNT44j2HaWcr3TaV25xImqEui7uC7v4ZCA2VHeFL08dVwmhNIti
nIIOMTqZ3qXN2hPejys8mns5zJaEpj/zqzp02LARIZ3Od7IkxZjtjdSFfbDUS5F52504M5GsgrCR
TYJs4pfRdjvUr3CSA54jSALsGQb1f2iZ9frVs7FDiGIFObWfYMLza+51Evl2S+LvGvL9CAsyng3H
uWRtJwHKn3ImDKk6481drLvqiNuSxcCHomazGQw20AUT9pzt4v2uICym4Vhw4GWNXe/vmuWeC1fs
HcR6guxTeCU1OoAkYZeECgS3WMJ03VqP/LnWDvwn1g7IiF8duMD3pLVqgFiHT5AMv8ydtpfeQy5Y
FnGFrBQCKn82cU/wBudaAlbV0EP9GnCyi/u//AmRFjNfEKHwLhW/qC8oLStbiRwZcfDbjsTsCB2J
X6zec3a1h8//7YWlP2HYKxisLvHPODgMGjTyYUR/WvcB3o2yHq3QJ2OekAHSZo4Nz/1p/U3CYAlU
8FbSt/LPNvaHr8lYBSDDOeZAz1PX6xZa9rhfQe/DijPGQq2rQqQIJZUJm/xEEecJiEt2hAgqoUgI
ltoC/sh6eTjaO6Loz1VOcHsR8zBU9a+TK8MwJKM6EEmWh9eqkMN5e6/SY06J+r1ghobpcRrN9753
R7LNNMCFBSqb9uAF/97+0R11RFpPFWJ8G57Rp8LLFJOlG0dsKWNUwvywy8lUOJfEGCd20YVrv8jz
LnvZX9bGp8UIHIYhA4zGHi/auWHb5wiyiyLIQTL6gtUa3DRe6wrpgzDLI3rtuN5fTwkol/IYfpJc
+dJCPrl4gWHf/8Y/YqsmVom23rgSpvYH4Hzj3GaDigsaXo5q4RVyn8o34e/Dh4Oeq+QKmDvUoycb
AbgonZYJoxo8JUdcRsonLB3Dd5zjB3tP06p54gWIo0ajAJJ6RdMNdymP5tT/0mcwU3E1FhvLuqPY
Wvwg9cBfwSS7SM8e1faK5Ye9w8M0ddB9sATKF8GRPg8L04Y773Clh4WDfuMBc2NZSD89RCT3/HnT
VhdXa4P1eeFiYA0/DTgcp0KXqJZOl9M61VU9HKKnGVi+VvUu+ueCVzYzvzhfOqOBzFhSDe1IL3P3
47GLdsXbdmSYC/w+PJGnQSiWeGbJLfRuh3FyQj+u1/jOgRZUVFxhOco9stK/wIGRW3ngmlZ7WJd2
LmsjiSn3KAEtKQ7+oOW43wFyANg3DS7fHS/9NZvZnas8+4D0CkNgPL9jWmorkMk5nnOnS3CIQuV9
DP+xDQINTIhfj1F6nKAXSIg8BqNQXn9hRld+Vi+tmlHKTuQTrLT7/v4d5GehSu+EFFYOjuwnuJqQ
9ileTHrizx6weffemPAyT5Y1Glvutk+Yn8hx55LggQaGkJSgw8xWdndUTcoXK+BBWo4+tjqITWX5
2xkNc9dFTWncNxuNIZ7Kv28+A+zK/J5CkpeaMvYjY0tr+2BOxF/5T2IAyKELsNTpFQqrGn2KQt//
bIjLKmihalE0QifMq3+vwNsafG72rBl85ZaKykGP7WaH0UukBPIfhn84qpKQ2g0EPIGCSJgCSzpN
ib1pL9j2SVLOpndmsCEwyj4lP9Y86H/Flm9Arxpe0iIw8Fdc0592oKsfsNpwDKDTC9WqUC1+tGOY
0MdxpMDEnpX2/U2fA0CEMXe8bYTeANA+/XNX8JfahaJLuVWHrOmX56yhbPINAkxpA2wBpuRsdAt1
xbEhXjjWjM8CTirzPgzOss+XDCy1VicE7gmpfIuFyG8Ih2tO5SRZortEOmZMEtGUznRBokBJqtxU
+vEgV1l97N+vAneDq9Ph8EdljK0PKkrxhcuEk59+jHnfVse5vTTxl0zX5GPHWde9ywHPYj+VIW23
mJzluWVuODMUgn57+l6m/Cb0I1UpI3wQ+nujGjcC7QbMPmuC/EPHfhe1YyihRwYO+wxYXHwK5XT4
XsPTmQxlF2pdeS0eFzR08OCPTYTYflyjILUtXjeH+QqyUKpwJdqoTgrz+PNcp8qGIhJpcVnuP6vA
0KmQquNCc7FBpRdJl5ItWbymGCF634B0N/Yfk0MPeoOxYxrIh+1AA9khUE1wC23pXv2nfUBXI9cn
FuQFruxoAyQ1zo4XsgF1InPaz1Nh0p4mniHFEW338HJ1c+u1kDn5kC5E2MDO5jUCJHD6qIieMW3M
BOQaP+nInrTe5YFsqE8Y4s8IZZQhfCFnjdV3JFvO5ti9J1ZA4+b9iZDFTJHclNJtr7hI1B2va36m
zVfnD0UCfhxhIvZWfP1lR6JNO1u/ZuHHyx4LPUG7CFKmYjAM+N7SeHwJe7TkNp1TWrKlTdVn2PDq
wY8VweGmPUGFjYjrvimp2swZP0achsCXG2iv0+hPv9L0Q/JUzhLv+aA4rOonqjL9/dM7BoISkxwy
TXrwzG7boGesByFsaxY8xIBwGiH3ym9q5FgOej8qaIxh2XgeYVdp4g97Y0/5uqZ5TN0HSvBib5Ku
fpy1/R0as5VJDGz7NLUbK/lW1e0CH0wUd67dIhQ+rv8Cg8wkLCzWt2rASlFKYOr7pl7Fcbz+1qM5
8wG7wdVB0t8DLtL785el7x2ZD63iDMO7USWpYpGdjtAsDpc61vRofsCVKYMOWWsCGhY9VfBxH7Vy
KRroussTeel+pNF7n86RCO8JBtJHyXoFLON2IobIXKffQGlJ5MjBVENCRuJyaS76baqwbrg126UW
KVWW4cSFXpiOLjUoQpJsiDwUy02xNiIK9DD+0XMLEjNDFFVaTBv91a+b5gPlZoU52sqWYdo4OCm6
q5WBjhj8go93lq5lG5Bfyug2u9BG++A+PFZM/FBNEJB1VyOrZfUkPKGv0yfH8erSeeS/CB3BAa8B
yliiWv3k8Svt5GmeYFXNZkFFxaAaiPlPU17GMQj7g3PO2vwJiDW642/Yh8dvtxouSsi/s8PJ4Rlz
81yyYtZU7x01kl6kzLVScCtvZmF8ZDuR55KUMhs1xcgQcxOSn6qrtbiIEMXkuDVYYOETLAu6/gKO
Kav9F2UaHLAUImzDUMOK26vdfCeoLO9m9iZ/DvOcxdtCjJHG4u0PQOdG717MhmvA5fveipxqAOuD
XUkMXeIdwmf0aff1uKpywx0Bz1VwZ2UM9c1hmIRJEfgm4aGAhVj5PLlp65U4vfOGCQIBStL//ZeO
2A9o7xyCkMXlyG82G87aeCYT4o7udtKStKi6LYYoe1w8aCd0g2/3C8n+wK4TzDgKeqzpaYCo/noT
Xs4p46TfkfmyIIEDzR64v0c/58yn8mmY9TozMqs7zF5yhx4+mC4ZL4QuHaXAAd7MmWd38oHBWKNo
6XlsSHCEACUF8mPmt8aYGo4/9mmXyvDw2idm5oUS7t8TShFKdI4A7Lhc7YbHzJvJGVbMiJVHaMc4
llG1Ksxll9HPzh7CBmL1MVvEu+m/KS5vXpSM1hzJsFZKknzbZBjbxWTGz/8oBrJ4OkfMBdUXLVin
MCGyPL1rv7vXsE0pGXmkaAHkNgCjFBI7Ri6vHMYk5fP7k3lzVjkym373QYxQGbkr9dkE26/tuw/S
gex8LWh7eeBtgqYit9XhmlhVzaELcmgv5D7SnVuEo1jZDv+yBs6D1bRA6xBa4pA0rXyAu5wycnNa
Eot3CmLErX4gxXulAt/1A5trBCecsXSkXlhdKpSwMGBcCGO1CYndwXQdENDcRbS4a1OV95wXPk5E
dq8qJXOPPCQ4nMM5MgL1jHvI4mo7kooDMIruPJDDt1a86u0C3+ykl1AK0DFUqcbpeLjzJN9Yvw6C
QDoniuu4bo6GPaebXlpGV3YNyfvrs+OOvYQATkDecK+KP4Qxz2Dnvx6KZHwV2zZwm98nzsE3t3LB
RQo/CfXVs6ftr2LWTdCFQB3sO69ovs6G8MYLO7OlQWXvGbVQ0s8t69DRXGfJf6Jk/9RbrmUvGFUV
z2n7BSAzzE8zIVxKt2dvyKVKuDrKzYG1ViSP7mUvOlNZ9+8HUX/dZbHo12wY5dJfiLhven2OJTMo
OKnEuDSSPN203WjJ1pPYzuCZLOns6+uTHLRZjz4148/HLpvPw+0pWQZjAjertpodCqi2YU8ki+5A
25DMz/aXTPm0qtCCZAv69dgDdmHBYRZ9iTZfQheXTOPRFSPYL9LN03ha2pfEstWOMxubAw/a8c/H
k9acAIP85vw5u+S3NZlimVYnmNYLqMusIyu0+jC02y0xn6DzKT8urYcYn++7QFa5qQ9dw4ZxZ7jz
bZYcR/6MC6ev/SSEKya96a7bVF046Ao1ty/4y3CRN2X3Io0n0arM2jL5/MKB2nywk1Ng1gGzvdiZ
TMyl2s0WXJdFK8WSnWR0+T68HLlOOBDT43QgS9R5zt4sEyyeGS+lcEUtcw65VIDfWUAfyyv7AP5y
+u1JebqaB6xcz5Bxq1YT4AsdvpLK103mE8PdDwpVdsslC5hdK1H+tFF0tQIzCiph118I99cLrhfU
LySyemIlM3Cu+tG5TOXwaqeegif7dBrr74AFzAH6xisfNuUo//6eXtvYs34fG58Y2VYFHnVv178g
ooOJ00FkvFH68ZwSHPXvy0AyD5IqVTAJNh49B+wZrgzDQY05JFryQ9BZP6i3DBf6ye2hkdxLuVM9
3pwKnmD6rZJMpIhLuSwz3TiZNcv8/bh7/f2SWAP/IsjNyBX4kLusV0MB9/0j6vq+YelqCTbiTwDn
dinO9Ei7kXyO1/VPSngaiT1548i87LvgKOjO7gmGmzgBGyu+nAA1YSovsOOgetBdPH7ajFzzPJTE
JDuD5phSkq26b+hmlvEl0JcC1rAnGXAnUM+5E3ljD3dc2bkCN7Vbt+BSISp+Y6G6YchvBal5kEn7
elWsmj+KFaUSwnU0QQszM6jCljS9m08YeoZQqvCAd4ibZWi/SU/U4118/XSuYrkleudkOvdFzvGU
r+DDX4mRhkzqeVbmV5Chl4dr9RUo1gapvF/t71KjFWK/qd0XnF53bicDQeU1cJBNO69ELileoQpn
z4Ugwic+OhsFCcLwIlf7LE0KWyrzmt+MDvlWd6IapdRDhYeubIySbI/r6gA3gevu86ngBSFTwoXp
qZZbm1pYQRuDSOyP4p7QbV8Bc/2dQPqbaCzk8ife58ZZx/taGiqS2frC0XlgabcffYUU4TqLEOF2
B2QypXbi0XPCQOqZ8F09ZthbXrIpsBXPMcVJugfh1MsrGd3bXpjUhepH+XuIeybIvd56pfaXfaz6
DUHPLNmEDshjN5Eukl/R65rvKob4GxagnXAaMmqovVUz454iWsXLbhCMEkkNR7QmMrviPUFeMdOP
YnBqtc8IzWjYNbuB0TWPBT8T3vdtplF88dN55cL52UweTKR1WEliP1Cn0zk8F5UErZdKcgKbxpXO
bOLi6YPOodU+KbutyoIpZxh1rmu3UmSE2FN7d5U+atP9XofWytQm9JowthjO0bnqmfLSjSjShY4e
3/U/hnryWuUAgP28oceGBwviij2RbbzB7UxWNKz1fdFmiGuQVKTdWuEfNJpV5+A0xP25bgM/htRf
VNC7vgbg/DTZPpuD+QfSToZs6o3toDWXcXQo566rhZIFU1jLNZaF+WwKzEF9PylPHWyTuCutZo1+
YdOGB9ldpqfjF0US3bb5KnLqMM08eawO0rm3obIEWwTN9v4u3GldtdHzENu8RnAjm4+g7BGoPQr4
2qj1MxIqAO2DRQ+aJZCQhnNNTi5INJL9Xy2XF2RVkczA1RSKeSMYMBDQKhwCSv44iB+ov3FLITn4
N4XOmpi7AME6V82xj4gutrhoYAM3GqkRRll22J6BBhECSDzrW+ANz2AOZMDO2B1n/DzTLH0jKkLy
OMS5W84QBBjked1Na+Z9sBwR5u/9kqLgh89ISauZX+lgIopxF++jLMHrmD1NRewQIENdyGnLUMmL
b2cEmRpcyk3iFeMXqsho8IfIGDVNIKdHa5x6bNLS0xVfWYrovM89zuFhYk6lRa0RjuPq6F6+d/rP
VjEMfQctI4rvY1A53ZDolfypFexVgQfomFcvnHn/N+HnsSrxWwtNkoF4pAbKPq4H4e0yMeOldKo9
DpJkII07a25vb6fjUQwzfS8+gFfNzTzepJ4sEd/V8Ep7GVONocGJgQijjiaBggh3L284dp2vGvJS
I1Snr8B5zWag+EsQeFmbQHyfkMcWYwMhFEN/qW7WxgG2bytitGYQB3d/vzxYpJ/MrVc5UDQU7xHA
7wQOEI+FWfzNRGiNo/2/Rfn/n6LO/4dEU9Oy47l6rbXiAMb8Bpc7+fDUV04jxCsrfpv3fd++SojU
cSL2GV0wSmM9fwhds1+IYogR229fgzZ9pisnsxbf58FXQdRhkckMKaWJVRaLfsdqDIGeu6HneyqD
jHpLMOMJSdH5i9m/lglxAUE6BkMnzUJP9yllww3AEOyfEt89n45f4gUlWEGKqBKY7LjNIB5QabqW
xOyngc+vM2WHQBN+tHocaHXliUUFhW79XGTSIJHK2vrpZMdJgDX9/7zQEAp39WrvOwCGB3tF4JKj
HVhGxSZIVVLZQKr+EiXfXeUWbDLFhPu99TePtVh/Fwvh+YXAGUWZZHO0v0BZXPFIhiemD0xaDDGT
+3Z3ulP/dblST9eBomXd/rqlVkTLnC5e99AeNUfD6hEFYSvu7IkVtNfzbzB6A0THHjFxrsmn7/mE
/JbUEthNbyIsV6POsVmh78NC8mdRUAOxV3yXaYHh4Zh39xEkioX5hlbiT55rmV9TDywydlzjRvJM
NGs6p4pSAfT0uJ02aRKOSPE4qcBbAYBKlBoX4nZuPFB2HYQ3q1H00byA4vz/BAz1OsBU4qZ6idDP
/UMfFlC0+nAdrTEguQJoeyvdpGiVAZpdQwBIHdwMw5dYq3wjbCVEajLsp8jqYI9Rkvkihp27Yviy
mMrMzMIfDxQ06a4eyRPXN0KMoThOhVRmAhtlAsMTfzhotkFoljV24zyeaNGa0sDTq50yXSYy+2oM
52oWVqKK67HrJjOY5staxRXnRz/tOEeIw7A2EeFJY6fxKPglTYCJzV32c8UZmAINA5H33szCGisq
PDvsURerN3nc3se1Th/O9vYfVJRBX0HqaLuHL9VHTabTsJhlHihHHay5zEybnHkgp4H9hW1La9Zz
ZwVg96ktVDfAxkk++UhS83PBN5vj5L6xzhPDOaknP5KklF6Ytegm1d6cxBnS4VHz75x+zS6zw5+U
0JYVJzHI84AEXQBkeK9IpWbZ98dnPVQhRwBMrolUvw6JWsAjy6VoN77cQXQxUo3+M1E+ojb1rVHX
DB+p469lIo9MNKTlo4/3TsiV0hsa57AfuIZBh5D0tF24v7GOX5L4horMyNMB4odkqktsdlMR659x
LKaM//g9oQ+MoZ+/1G6hShiHEQQZjm80GyIQhTQok2DNtuXN9zfCqtrMbJ2uUb51H7SCMKpb5sLV
jlL1D+VyuXLQjMnyQi7RjTy5GLU6YP8Kofh4yQhsqeRaA8aPTWLOlqeFpV3/LZD41yKYDnaHZjTF
CAxgeuq3bdTByJp/lddV0Iu0u8XoVA/vkZwXU27iUjvqDLdgWh4g1kq9F7vInKUv+Yizy+cnFNgT
eDExfkAerGIO24OnGwMxRhgRjyB8dTGLZaPdIZDZbScBi06CSZsuYFF8bphRelbHs2YAngOF85VG
LeuFaaSLsxpL23oDIrfq/xL/lIGS9yMHS5a2oNUjEC1cd8oKYKS4212SHgNJ9dlv/p8O33TbzJ8Z
cvA2ix+6MRq3bkx6JO6oq6UNoP3gDcAMEwyHibnIcCTh1bRkubug7gYdRW9upHAqQG8qUMC1Qc2y
iJTG6VfC+xSMqD0ln4cj6l4H48Gv56VQPNEtOEXnTQ7UUqzD+DW4PcZs+rx7O7+iBj4PW45WL282
i6RE+K/o1GZjBzpiupggQaqA3QxkIYY5fRJfTzCSONG0TRCBzuXvVuloCchNHxPAS9Zbj6gGtnBO
tGwTy3wmMTKw+1/qLaQ8f1tibRn7Qqt+9O4LDGPx8RIN9E5l5UdVjlpT/oXgZ0Hs4Pa2+Mot/CCL
GmemrMQ+1/jqIfaBAq+SPzB2diJGou4mC/5vvMY5Pq7/Kz5CuhrzYQqTdcyxj0oIUXMgl+kG8uTS
BxWLEtBybI4fZqD5XcF6JAYOia/oqgxWE02BGfbJ/8j44fr1xrAhwlGrg84wmH/8vZhX+Z/gimwA
4o6npeG2DCA66cftasDf3zHV/fp/7wgA/3DKBLsvKYp8Z/pU17/cx0Dn5jkDrmdpPlH/x1hdrnBZ
7XVE9p9BQNj4l+s6ukZ1CBt1rgrgA3pNmc+DZeVXb44TJqagxiNVh4HJadc9wHWi9hQbLKrHXkEx
CnLIj1We3Fyk5fSZYw1BhMrIxU5VLZph+mOHDH3qy+YW3hKpzhGKcVWjAOX9/ZHoImW3q+KlDC82
o9CoGBp36AY1+ego45yHED6wnZxh00GG9yinqy/AEwGxWXEVekxo1xMvdHHBMI/hTSza1xkM65R7
2dNGFNaHOqE8SUA16qURgCxURGskAmssIjnUZdD5yV1sZFse2E3BlgNsMGn/73NHvvSvs/SYXXlm
GSCIBW9MkyIO/vovPAdy0hdAWJ/+qgmxq5ot+ZUdemJDuO4e1Usnn2H2slO+YSNgXzWRwOJRukwz
3FB9EvWyEl9od9oEo8SGl0JiEkpsq2OP6oRGPEOKSfdopGIfB2NGW3IlmIhk0Eoho6MAi6yunOgt
gkz+CB9EjQcCzjELMCzhjt5PjYVCiwHWI+ECS6b9p/DUglu7H+Vs/AuRnS2weVYGwpbVl/C2IgJ2
tOFzTgGVsRiOYzCwIlzUAOFUpUM+Azp9JfHTQcgK0VT6wKWrOpIKpcbc7jhWXdCc5UnPPyOWOZvi
KiSWtyIxNDwiGdzP0/u477paAiaWrksAwcDt+f7AJJe/STuy7aE+qgxmtFMtTGZnzasUy6MTFpJe
/jDWBAOjjxlAfAGJWTMHyXHinPxo0lrU88P8u7nF6XYj+0lcU1erOzME/JhvTHr5wxLEwLqdyN8P
M6bRbou6uY1ud/4dvlVGQFM666010/pXYgMS653CP9OmxgrHD2yLNaBzmhAhoFuHsY5p3mfX4ZqL
AxZJ0pZD5Ew66utoKg0jXFWXYy6QuLgl77XSusX1HpKCb3DlnSqpEEqalm0dUpNqiOaaPz8sWE9q
30XmWLoN3I4TfUG7tevRz6LsKfZEIPtKYuWYz3QezZDNYA6UIQucxYi5Gf55UJK9iZfCnn6tgm+x
i3r7RPqCavmUszl5R5flcO6ZriOas3QgIBM/Dnipzy4rsxnw8ka0sIq/cyJfMaoRN87KBiSGdJKP
YdbKMRBaagrktgWMaiciwxc9AJn+pl9oKom621QDoUcfd2rsEYAExgYcRxmrGm3nDQhytbvnmeIv
W5w0U+hvS9pHzHVToJcvtr5TF2+A2/V0Hd5JaLRk/IeV7wkaYKJkuk2Ssq9aP+IFN55Lr0dqlGab
uRX/goAcJk5jUchD5BpPyNTH7cdpjgyyE0JLqYint2BJcv+rIl8+b2rvhpR7b5RBQKbK2+8quP5e
F6IvTc/e+0bd6Ll/LCFDFg4PhbQKkCs0Xp/iosYlXE3JRNcCARI/1K506jh1JVOoAc4A9sZuaqNJ
CcpioBUI6xAFnjgVk5mtTILcCbn3nh4owvBpTa3m2za/9LQ5g5AmZkY2pl0d6ylyYRmQSpwN8zj8
kWtp+7LBFlo7GOuvR+I1k5xoNWjSOAOI/iCt3I91sV27F6RNBOyq7FPGChsJ9ll2m6yboLT3vHL2
GXeltbsOW47ar9r5e/44+qDB8N9CqIjp8lKF7TOH0/dqhJve0IKKo+YO6KYL/JjWkd4wPvrv23qV
SiaedUIbyC5IBisvp0JKYxA52ZRIrn9uAiAnpACT0TNGV7lGkMnpeHcv2SndmxdPHllncecjuiG9
AcXRG/NrOqy4sgIoYSpD1eaXMb2FPvVSiWfjX98IXWEdRCGtOgo4dL7JqYaxSucC45Pa1YezO1qh
3H7sn8gANdBJ5HOlJOVhW+/UOtFDO7zKYXNNvlxFXPctGWe4Y16KSocgMl4wdlrcTSskJegyu+Hh
FSgv2Lfopfut7W72cddYXhcOAktTcpNpw56ii7LVeXqc+W7bsj219K/Jo29Jre6RsMj5fjyYeOpx
7Dg43dXFqBa+pqE9sOMMYVo35f/xELVVVRXOp9vaFSme+Oewns9UEerCQUXr4JtkF8RcsXzS3fT9
is2QCfwSDqrkNnbQUez+m+JLZv2jiqxcQAUBjB/neQh/6Oib5+BCWZ1fEb2+UHuvYlkW0Qox7x9p
GEVIhGLEj3yngKl58YrbPtJBfhQgSMQjprUZb7DqdfjuVbVs+4CSLDg/cGiF7Y43WX9d12Q2M4IK
OhP4g947mYmSdgIXkCQB7wguOYj7wle87zBO8U5tZGdTMpr8isfzBwx5n0SUF+jQExzo5L2yYdTu
RAqmFFTOe+tyJMNtvyoAv0qVgfw4A17myOqwC16r/PQXQXGh5ZjlYaWWS+2rGv1QIl+r/3KXCXds
enteep9fZ+XBIBgim4XzJb5X5Lb4ssCyRYwt/dyldf+nhKQLyKJSrKs0QkNLDxibVb4SC8hBMe7r
mTsZh35rAqzqnrPiyaT/Y0bNCEBkt+ojPWyJHhKLalS6mxn33d4BuxlL9fHYTF9KkWUeba+Metil
gVO1mzyvWFybtt7HDy5hJgV3Y/AESn9/ejAyvVOlZqV/n+IAJT9Cw6igDeCzGbG1fSwNv4IhY9v3
buY/IN0IKqXy3ySwizb1ninsXPWV1ERbTX0PmGthwfcn9r5qSHYrMsJfWHliPf1GpvpvaSt3yfaW
HRsvujCo14sq6lLrz+iG2cscD3M6VqCgHeBiQL72pVrl90Um13/SVFVHwU/hJTEtCXWgWixoyS7m
/J7Xh4tlGwaMFZ+a1UHO8t5NieqeYRrH1s384PfupUTS0Irp8Us3w+j3OS3sc8a1CJPzRicvzW3m
qZv94w5SjrcG+Dt35Te8F5OgkVnbU1wzR92Emuv0qeNLhb5FoEI5vBjuMcJ2mnvrdVBC7LgVtfBY
zLuHlzqrNIfqN6ZcCVXI+wmoCs/4bzW3wE2Bxpe+Y+RhFnyczsaWLecGb+E5dGz3frqF99hB+nXu
vy9Q1SuH6AQ0G72fm1hJuLChNVRxM3Q96Sb/BjLWDeglatCef73IKyZyslgq9sJMis+QsabNGBeZ
zRIYeyAVNLXPDpzIJFYTOHo4OPqWPHWcxzt159FB1b7e+a9Ije/l8NUdhKdF+aLi6DxVC/Elj49+
mJb4Rfe7DIYdDlKWquQm+vJMwFqdCiGyxlDeLgfY6S/j6DUyThTJKMor5iJoJ7KWOOkXUUgyE8DC
fMjRfgIiTdWO5+HmFPsDbRK2RPwDUzFnPwfBHjcEqyCpSBTOuFX7h48mm7ThBcEVrJ4vWqFXlSKg
NkczaVt+N6535d3CCVyWNb3v9fS6/nxn8fcf6SH8aQ/XvAVibq0lVUS5XPtRkUwyqAy4tg8/gq7L
yvrmR4g1IiltVW+YmCZmYj+rlXPC/z6KCz8zUHhQgO3PefFZmww9UcICSPbbEiU3gb0/E1RdFoGX
/IojQVo4xs6WBv1zbKfUEw5PryGx4+VJ5VnjQ5u4cdO4U1ziumdy7SSg4hMYdAvYCZrUAZ3Y2BQK
A7XTGD5OO00spMzCDCZpNo998/fFSRx3jqMS58oQgIaDoWYQk1y5BkA/V8esnAf8rrBB0shHvFQL
QLpR5ysBHPQUO5zlbseGraL+WY6BMBfWh1GZUkMWz1BZWmMAR5bh2Muv5BQFM4k3Kthxx055gDCS
ORQeJRROHu678bS/PdwHP+uIM37zUhhtLYCIXt3zbSsOUosN69kYxoepSKKGiSDzrZ34LG/xEnRr
Rl93DWPadGp/5Fj5JY9DEUIC70loRipdHtGZzCxeADaPsFfJcjPOtEAF562LpAhgQiiNNxnwCnxG
NeSasvTJHgL9OY2M8Xinh8bJqjqd2aWhODRXCEac2jtHAl2+fCO0cYRjejgYIaL82CILXVllk1f2
dOahowHNo0kUI7TwM5bVhpGWrvofM+FfEuQfERjBVI+cMFLnjBX6DMatiKfrYwNQ7goK35opaKxu
zZ66HctF4j5dM908qJX/Lac50crBGUMMhcxeqrVT6Eaxy3PmzfnJE2ORd3VraY9Br9wBAxx75t43
pMLBOPPbli2cb+NI9/OoBS5tQ7CW9sXnG6dGT8rVuzyLo+Ca6g2EmX3i1FE6wSCGKEYT/Bugw+v+
AmaPi4Y9VglOpofJh9nNz2jhjIaQaZciCWaIf7b6cZIbdMj9BSErADszobYu3gT8NYYDWtOZueOr
pxeJgMDb9NVsrpgrSqbswHGKQwjNd9SYRcfeYr0EtVJmQvW4xhfKVeFPddksqqyj0AvKOmVDhpHU
hHGIqybuUGUot2Bc136AoRH9DA2pVGXA8yuvH/a375b117CdvrXcJ09mHqOGRFFpiBJ2vF5cla20
Sx2jAfwnz1MQYfzExYScVBaDKnvvir9ViN3IIOX28BJtFhdztIi1dG82NWPwr2UunxFnkKDRTiOU
1X8eUrCgqGrIQHQKfLSSCdrUlB+FrW5cyHqb0Ah6Il2gQWTqDMNY8njPd1aSiZLwmEmKB6yCgwXl
42BajnArkAFoY2wUGEqUHD2fpkwr+qTOkvQ51dhtNWui5kbDN9quWowPWAgJC/O8kC55puL35Hqb
1h1m4wFEriv5JhH1AQWQkim045nBr76XU2V8rWLxwRUOQ5mEuskOMd39hLsjfXTYyShenysqnDOV
qV3meK3FGs6LRiFppd6l7RFZQkBoKDJ3JSKIrDF/agzpP3pzQSOyJjN+sxR7P7OQOmpWcmFR3qrb
O4uZ4HaEie5uesET5d3BBeHb73d8H13OLx9HgPkLdF5OeTQ3zb1xav8bZfMVi20m2/lWJbugw1pu
bmvDwKLNgYn1IeqKhMg22Oz5Jl70Fk7PJClpSprddgPt15GNBKmGikTD0wqPCGI4eLMHgxCtqQii
4qG36yQuU5Bc4icxO0ixtJJOD2csRgSwy9p4mdjoMioWEYE8kFM1upaII+xVIxWhwE9smVhl5Vs6
7fWH727pTNp3vI524HCNE9ySaxumvnMuIHttoYtPo/puZhvqDCW5q/tolwL/q2lOYBLDclLRMgeV
zLd3t3XexrjtrcluET3t6rP2FGsI7uNDfvieu6GmYeQpz/qxxRW4+FOYopebRxEqj9VG9oqr5JaJ
OHmyXDmsBiNAwcSp2AmHgOkKVlwjRdHTFh7Be8MyP8nTBPSEdDwaPAb8lYmTq3QVbdinR8YVpd3D
7kY+DobcgIk015OzRy/MgjuMD7gvTBh+A+3pyyqckQJYIva57lkc8nY/zViX0ERhfTKj/guQGuS0
KAfE8/c0rWRdxY939IgxnU05zW0jshSFkACt4t/CwiwMxgWxu+NFr5qREC31zsFTzVHT7EFv1yQu
dtoAkrb6S/2mirf9BrocvSOrpd1AnmuFViD5CFSIr3uKxAtcD0QCh8CadcEwvfPzZw9WA2wYfy6B
DVEyLv7p80DWymyaUK2/4XE5nOrKtaa1vl+nwEyuj9M0HeEkAY3WNHi5YFLqX1v5IobO973unlSr
EecnIrPPwo4mcfrcjZxwWLXxWRgRTIc4YTkUGNBMTkfBf6Y1nlk8IAqdAHsm/fYEnj9Ljj7BYvY/
AlB7PO2qfFs0FzYFHBIa10L7bg1CilRPWbCNQaBv5uaIVa1lDeaA6qADo6guMKq9WZWxHoX6sMG/
O11LXBway/fSyGIOoszOIVNqVkO4zzhrO1++sjMcrSqROT1iCUw4ehijfXjn+jo4rZQf3jaIg4Qr
ezFF2v0GaS+AzRK429CU8QzR4XKKDig0e8NFHxFY+dxjAcc0vOM/0uuI7NHUGv+l37IOY+WiSEEh
qxZmF747S+kvHA2WygMwwOrTWniDKeZ/0NXsZeNwaSILcOPPHmZiw8IFxWBwhenLKmQIJ77A4esd
KHnsT1EqkcOs7yRE6Q+7h0xiROK+Q1dgfi4cPE7rAYyf50yR61ZJN99+IwWWHK7w63a4dxpuPK0m
iO1XNbSMltXbdYseoLSkEiKwDQEGFyZ+97P0DeuP1v+rab86SXiyHl3iTNb9se/9iqfjiMOHiB4f
OdIyXwNbyIi0aHVkwwd8j35yJ/p6hdblDzDebGpmrIjkw1kQhF/t7Y+f6fQ0Kh6dDcY21iVH1Ze6
DGPAhmZRBXJ72dER3H9H+V1h6iX7NZ2VgiKFkdgWJpqO4tR1Wy6vt84hvbNP/PRWalTfI935QXki
rKM0g9lRQqxacD/tBVHCfc2yN5K6TGUzmzCtGncvnh/8zC203ZmAhotnrJYxn2AFF3EHfNw2QOEe
sii0/OrcZ65gi7IF+KwDJGb9sG213SS6HuxNi+9NrqrQ9jY7m3mia9THeszXGRgBwZDBT/RQcLGi
8jHnrzKMsnw22pM6csRiPTpdG6/2Y3Xb+At3LehoMiCGy4PA8rfG+e/uH86Juo0J3wDJz3nmYsSo
N/5Ldxq81s5yxjJ75d/HWk0+7s1gWJRVITt937ERQpe/XC3w62HOQ7rom0TJz9BEhFZGL8UxGJM/
5qk1+9GvRM0WFBvTTXHSey79A8w3sa1Ly+PQZAjD8/bzZKqdy3iWBb9DNMV1XJmSqdM34kRZ6A73
B4pAJ8A0GVk2vTLjsv23LvPaCpd8sXiC5GPJk1GbZxnFIeU5ukmPbEmgHWcrg3D5J07hz3tv1lkb
9okWHecQy0x4BWFJaqpvfDy3A7jnDCqjJFBjK5lNkOTDrCkpS2n5SYZ4xCuyxHJEJqtdYof/AhCB
DbV5JtbsaIKaftnqZZmHc1tBXMKotXW8zUIuLnAkrOW4eAf8/i3R+bVGmUn7zXrlScpxSncI43Qq
CCn+NFofQp0KBbwzF+fUTy86pH6oYzfP3Qh1+gH+59yca52inMMX840PnAxSaFtp7n5TseYg8rBz
70ILHGHScsKdPjlrV6vhkyUV6VZ3BUOUhPGhkSZt48xU4e4zMaIT3BWk2uUY9/JE6+hoom8Fl8tE
ZpvdssmVxLGCiI7rEUmNkGF5QLlOl5WN4x8b7woPafikeFdgo5VQEwuuSiK7w1AlAJmMzhAdiu2E
l4diyw5F4cxdOoCS+31ifLbpQ0vP9MEZW0nRrSj4G8G5Z0F6roeI7Vhoc8fiII5MRqkPYRqL9i0F
iUbbJ8ygH6QKEt4NyxT4rHf3fS9DjOg63L9cwIcWm4MJmyF0Em+GK1ooIocagDZYF+U9DIpoPo4p
MmLfmOokAZNNZKzjxNNc+TwC7Ea3pqYwY67xzpVV/ucnkgK/vxhBccihKDfomkfBRowNzohIBAxQ
BDUMRnw2gkTX68SzQfNhskYAke1XnWUHLWNYiPT3JuPzajg366FpW/UBwioMhyBl4eppqM8kkc/C
RF64hP3bH7r5fomi2IutnBam5PU3KSoTodZww1O5sK0XOmZwL5bvZf1iPuijDGkAkAUXwTxxKx8s
4Sybvh3j3x2on8RXA8Nr+jEKbhfAKgMnwjrxNPWbljlDf8pm/FV/cPQ9dUXQYV2PHMSZN3yxuj5G
LG02m42w+iMGp9A3kirrKX8CwhZkaYl0FD3GxkHb5++FEFmSQg2vL1DGbjjmScLIvQCtTnY3q2hG
R4SVbr98O58AhnWRY2sP69Tmz8ACYko3nd6OzM+jCEFi42m2CAh7CdnXNsDGwRRwYyExRw6GNC21
FHE25EWsL9i3Ejk26JWPMv0e2RuU2IC0/1ukH58kcqqBcIhB7CEgyaKE7qrFj7SpGaW8feU9BlhH
AGJD5A4WPlhM+AYaV+U3HTzwmKLeX8XQwbbIwP09s+ILCZsezZEIsSX+WpyrNp/XSqa73S0gOe+U
d3LAwFf/7BvszF9ZsM+fr0yrJmTVuZesgjXpkFZ5tuz92P7Q4KJpWHibwoxGaiTrWma081n9rSb2
HwAI9orajG4VVh7l4VjcuUtQd4sMXp7djWwSr538NYQ8ngIbjsaD50HhOqKHvUaPJ0vwNu+qSXu3
mMoJhzDK4jEDRjkXdCfV9zOeX867XESw+vZy4r7uLxMP75Wp6ELuy8L41dq71AGbTeYhsiFrAXxw
39LjYV/TzPFG8VNVXPwbo32pzWUOhmyrwtxc7Ny2jeLoqERsHEVSFKPgAEI4SDNXII3ZIXVBlHnQ
JRb/7K7NiiBTk3AauuFd4fNp8EwAmc2P8CsqSPwPdvdPO0g21hihyacgeUu04zeMXxcG5wuO/Djs
i/Y9SRZrA3eEn3e739gYjl17yhXgwEDl/xV0ZuWEOIzJ87+3c5Xt5JYwHEQWKa4213xVffN3ye4H
Q33S2GO+b0VC8EL4rZy389arLgELjq86bqImR/sOyJTQc13RGB/SkUDGXSMCWDPcGTEHx7KIMXyI
+OdBRb1Sn5kKNoEoB1RuIzdwzdLFpoMR8hsn0tvBG9sqoKEyjiN7SLdil3h1kCJIMkjc5qpRZiSC
JXzbOgQexVCb87NtfWTnGvkyqltzHdPWsYsQLBaAbNzNsKKEJtfteDpw0uODaDzDF86NW2IC1JeT
dT1sqAT3U6YeSPF1qx63JWXDnOJD80+9roALKiSIwnUQU+RlfAR05HSJSET273xusVOFa5sKiCN3
u+5DljdIovGelpbk9oQto2qF/ANBNM77KdpjC47l+r475n5xAiVsGYoGYx9ZFbfgOPPcsQE7RiyT
83nLdMcvMweOiaXfPW7SqFhLxHU4uIXyohP9M7XVAxilbctm3yzYyOeZKM0wnl25yMwpNBAoeZb3
oOFM3WsXO7Yvv2PILaKj04hCp7fg7Qc3aHbsERLpjD0raKHJrRA0QDMN5medKkic9B5uDDdOEh0q
JSCGFaKXddZqRhyLBzMeHvc657nJN6wNKhA+aoIQDbJ6sP3KCoeczm+ackxA2YMUYD3CXqgTc7QD
6PkwnM/c1QDKOsDy+wW4ZmJWF3pgJt5ByPsnqfbWGSJGxz+cvV+dh1hL43s6FNEs9GWTqNmJ8mVR
P1inD2yuz7Wenp89E75hdzr9vKtxgHFQrbqDwVUPd5wj47eBwgZi9WDtIfYCIvJ1vROCeQpMvvli
oWcZBVorgs3pQ0gmFsfzm3KzBfZWaWpdPevQ04I4lkO+/pRxV21zMtgGtTwo9dgPWwU6oLmR7vZ5
qhQqrwrg35pXF7/6dzyGp6SUIDnhoOteEJR1FM35kuZwQrOcIyrAVPgWabMw+35B6qQPZ/swGeZE
8nOhojK3RNoOv+idHDH8HVmwrAB87kjQbf+zrfmFrhZCqetfQ+ii4t/R+N+u5p4vvY5ZokYD3Kgg
9G/HHKJK3UZt/ptl7j2hFZWW6eY5hQFQXsPdAJivMvU0FMLLcqHMWrSwdUoKdfn30LB9OqFjP1Ob
PQrj6wDk1KevssfUYEn3QVVcJVanvaSCX97kLKhHczqfg3DBn0IErQzYMZ2OhF9oQ5XPw05OZN0t
Quq/y7MkLiBZqWssWO/Q/WNSDt/8pmsoDjcu5NV54laR8iHQm6dlQNwqkbsoVe7Haguw4fyhmpsH
M/yBiaLROSPJI5sDTajGaXRD6yXOZQaOVnNZmgyIu58JfP2YotyoRKlPSNtmkC08OrQq1fCIF0PT
ghON1VbQHonUxY7bBg4f0j0FwDjjxPGCFQ6a8QV3Kpxe/zseXuP36KsRUMznbnHWAkzysRca0bTe
LgCrK/hIjoi8v7SjUY/eINVQh8ickwP61+N0OX9OL08hY2GbLGJUhpQIGaSFKpbyat1nOyuOgE/3
dppa0f+AjbZrKnGzwZSfUZlT1d6DGPhzd19Po9iXEyuWajnavdvr8mYwUT/ufpG2w90+ebmq4Akl
jb+x3gD0n9//+ZkIb9xtnxnoUbEV1EwUuNzXASktKr6hyJ9U4lmfIQ8tkrZ0HxyMHTBaG4QkNF+l
xINEXgJz10GsEMYXsP6wvbyInU8iReK7oo082zaUI4t2Pu+Nbn9cHG78FOPDDr4fyXiKlA10655A
vRMWNAMCYI7x0foh9yUY59JfP74AT9O8Fb1CT1VJUq9r5H9BQM7pjy17HIkkLgSVQG469PrkJydC
wdoXV7Bw2idxZ+8sPDni5HU4Uw0iwM5Vv1gE/hzcj0RNKU9sxnAQB+Tw7zBV0f3baO2HG+fujJ3s
BUB6S69b7B7yyGS5XGl+tG7GLWa09oUpvLvqbbqsjCchJftS8RtK9BW6wOidzFo+Pk9HFO3wRa+h
c/92VoGrdAKnUj5yv++1StamVDdVaQibbCgGGGK039JXgMLOwMx6SRvnuiApxRGjb61MDLiX8Rfq
hnMLKyxWKtG9YMFgrjrnESLHlyOQLLEvOCo1dSq8IkuR0z2RvJfun7UlxjBx78NBnU43bUalXAk3
v3Xn8d1y70gqNO17w9GUHQ2ncJeJeP1CeGXKv8k4rVJtQBGBAL6tjYDTZL4fDUR03TRfy0UIvsAt
GJeYtQRQ3kWDM/Wv0TS9IaMj7uDIleaMNKMBntJajjbncbOn7o2mxHLJVnkgPxzlW29HH5vfcxwg
8fxi1h3hZNt6oLegO3yNGPz9XMpJGXmljh+eDQSeNzDSJl3WhWgNmJNL0Msp3qLIHnJtZuJANDnL
tAdEFHXJuaYLYjINlFD8mM4WEaT1hCOf8AY90r91I9wLs3LsGBxEXYCy3tcWJqhJqmV/MZSJZMvZ
WzZyJYsptG7C4LRmcUDxA3TPu29IMSOc+RRiL1iyCCmRC63zjm4Jrpdz0nSGhzJPKfFXRKAYBj7d
lyPCkDf80MZxr3LCp1GNVM+CZxyu2qFVXxOSiRz3+YPyfcgMLjW1lxQjL+V7W4k/OdviUHyaBAuD
Kypz9F12GtyD6+nqHBj1w+tnmpz34e5CuYT0qbZ85d0EaETFaKl/u7msQCJgbl/6//QKw80iWq6o
bGAP4d7WAevRNCQLMUcyd1RXmlNCF7Z56wnw9CEq8xv4wIwOJ2u09qrl3fQsrOSz/1c+1MiBsF6O
1aYOKeDMxafL7zCcLrmxt29NHS4OaPJ+V1ursQV5THkA7qNCqCN1tGBV98TqsGUl/pwgXQ8HAKxQ
jowf3Jv1vOrvA8dMjGBU9RQ1flWhwWyFOU3ektsaI2J15Hc5z0uxzNrumaj9lGG+BnnLeDvHSKMV
AV+S/NHIRAp8AxsXNURG2rb/JpCmyc6SoffwHN9ID8roqZeT4bhLIuUjQd8XRbuVDE3zf84QhTX/
30Qg37pwPCZ7qvuNFytBK8o83/v/jor0m6j5s+imHoDKpLrU+Ht186g3tMGKxwz7lTGQK+tiQYit
DyUi1BuPeop3dnBkhqnDYd4QsYL+O9iUFn/P3bArxERtS8Pp6GS6/UVNYy3GnnBpET9DWPH93dpn
T9ZeeuleB4vlzmlLHb3P3P+jOkvu7vXQNshW2e12BVi8yCVvHPzYdK76YMJ+3k77OgFn1cs4Ihmg
qC0KUsxFAxZq/C02yNERXKVrkHF/lCqB2UTjb4YOPpXVwVWdiCoVGJqdPqTe7joDMG8OXgq4/k72
HSL0nicEFq5buk4CTwaK4sKzv1cpruN4kwSDD0wXsy9I3jdMKfafglnSNhSC742v1NuffOgX8icT
ciPHjRuJdUcjfG+rsJtW1+gnGkL0pQUMbQree6KuRkuJ/odHdqd6MkXNkCE1smSHgqZEEgD1Ms7T
dgnowr7H9/vFeIh0zS7lXtKZ32eo/BmcSkZNxBxrAnPOF9htfO+HTOFtGFECfvSJGa9l/TlLk+q0
Noo31zWSoGQnCcHimKi86WrCfJs8EOxdOUHOn2g2XE7322cWhkkZcwTLe+ROcEeikB+1AEL61GzP
2sXqvAaQuDy1FrOrCGdoAnc4FmghMD7wRdGbJrV91u2nmWFkbDHjcb3V0vOUi4BJIjLBA73sqd1r
/gw7+M++ynAS5G94okGe6DWuYNgY5DKpEXBl8JfLMg9lCLn44cplldydwDOCCkUWDx2aMOxj1E/E
PCvRI2BPS4QJ7pQboGEyoH9bTY70DBlM9NQa9SwWAOhud9x+A9jqT7hXTNj87+TF7bwXsW5bDx9L
WZ8zUGNiEwyfRf/E1JszMgOUCNSMvDymN5UGh6t4O+qKuwRFGH9xNoCAjZXCC+DPOGq6VSMxcQ6L
Pah8OjPXG+Bi9RftBLaB64+pgCNmK+MZGVNDkUpySXs5ktmLi/Fwjk9SYNVM2N94JsCenGTOU25x
4l6sz0Wweu7beGtJLKbbjRd/47BVmZNDsmVbH5Rvz224KPHKmyFVOqCeMLhTFDSheUaaOgjkeGmH
1QMLb1dmyo1qwquNApz5AbqXjLuy5U3Tfu6s3189HBwpUMVa6KXvZA0SlOPB2tehtme7Ra9ugSFH
k8qga4nNxT8JnNh3ldhA45ZHFnoW4bvhpwkdOju+4mclMk/L0VAMv2FlOv/uvYsxEqaP9oELrGUF
4fEq5JKdKFqWT6D+sPDy8maK5kUD99TvsT4KYkPyM6pdSJRweSWYJUXy2C50GNv/uuXXL3DxxvFz
40gInVOumpZ//aq9VYZdfCeS9BjGh8kEFXBVOxQ8ZDGr/g1XCve0QBzNT0GK9YD7wSM8OWpsbXjY
kztrCTfUVA1t+tHoSmoJYn71VqApjTqsSlj8obtnkijwVEY9PCd9LUFN4CP08//ZBv07li3Hmthv
MAYGC466PxnW+KUE9QKbt6Nj1Ca4k1dut8KPMh5TLNyp7zsKTC5G7vmxII5O1gZ6uVCeKLpE1xat
c/pSKBTdTDH3fRvIkj4Ab4V+2Uvr+Raiq1OVJKY8ZbyIqShqHm1FQIKfxjOd97bn0D89crzR4W41
Bkgd07Z1C7xMAfLd0FOQLur5wE5mnWI/wgxkuata7/JyJ945EWb8T6us7o5OdtIdaKU+9EZwuRl0
KKavB8vVP62Aa3WHg1UnN/cO5EoP8ms94xSNYI7+PFIHfgVMon8I4U9pNWQhSC8D2YARX2Z4s3Qt
IOVrczcoKoLuXoWU4EjmIpuhBovoTwqljVFfaVY/8ON2twAFwK9FrZ9x8wxHHwEFCYconEcxJA4f
SNtR8o/ZuK7FJvshSas3AX8dMUoGMneCOzaio64ow6q7sS1r57pukdu32FEcbtbWL3MUNtM9VJ4r
owtj2iTEn3Jx77pYG7iglsznPwesdUxHbP5y9FGr/Sg6qVWRk32OiM/XXiRoYi8sRe/cWvCy3Y7N
eVLXxHCQkeLC1oYdCY9iA211uk1kWY3+yKxxzzeHTppJ6dky5WUPoZVJEigw0fOUlnGPA2jjhxaZ
tUiTvJ2rJLThz+fL8IokY0wY1eI0MAQuKrJjHxRlh8CAeS7hlp05xXEvlZUQGE02pX34mIdMnpiY
gGv2DPFEm0sCDcL+xEMXHkbcH511JFqQagvrypsQeoz9sHfx1yHx2ePC9g+bh/PbG2KnziZD2r4I
iX1yAeVyZd+T/P1hRVzKSTu2KCinnqOZA7JgjxaRuem6XMbwt/E8tAloHwXB0mS4I9EgB0rzoJiz
XSOzrNfL7pZsyo3AutMBZFxFJ4YXyl/PDQn9qSEmljxshabVE1haMz1UCfCASVAPRiwqXQGcg+tI
pzhnfS/X7zTMENNo1DEpi7IoxQyNgLHuu6h5zZFtb5t1ejwhu9OUC0gqLv+bDcrrUCLo6cdE86Rf
W/trt71utooNSAXPJilkXCm+IS+U929FlP7ZqVvhQbiC7V2iuAAY4FqcAYafNmIYai1M5Ic1GL74
sRtU/REvfQcpL6P96/bdc6bzK/OkhtlghDqAXodpFDo1LX1QtyIt5nV3i9oCKEen8jKXRPsrta/Z
LiGzMBTpiv4YaDlWE1eVsDp1wNsvNvV7oqNvDEnk8iDQVPaMlRRIUz+BDAAmjydWYrg+FT1l6fXT
X46FIaDgWl3HETv/waTKZdQqXKcyxgUt6GtVCyY52TUfKoqW1OKagvrQth3hbNSJLZMjEV9G9jeA
L+fd/mNNbF9XEq2G3ySKLcG9WyoQRpLYFHQShiij9AAgrhVQPtwimC6YYyO5wBmW72LBIjWf927K
2/jFVUYb1veaUY0OyVYwBcbAwsx+x8AtksrbS94zHHCHv8ZtB7pZZkjRhvoSTpYEQAqugqRllglC
7PSLHY+8fBuR3eSgZnFgsJAGvdnQrFHe3e1JAOmG+LTBM5mWi+4UBYzEs6o/mo6Z8MiAMkGph72f
JiGw8hGZfqzew5ysOOHddsCGbtR766xmMS0i82+NDF1F21ZGzz4oZlYpxwXoIb4Rk9z0P60hi4Uu
3bgLTpTjPjIN6ybLZKQtQmzHsTAhnWQb0+8VwWdeewOmGJMzyPrfVVaDKqgejxv/Kl9irbBSAr50
vKDlAJADjOy8BH99XwdKLdj7du+XnZWeU4sybxuhD5o6TwfoNRXqKQWohSKdmpmH7FWj80/2tiaD
67qr48eCLXKZuiaKjCYW5FD9eXkb+Kbhd8vwRqX8OaBTmF+Sa/i5ptDd5HdH1fkSWExMroy7w1O9
lyS/PJC67laP4E2cmQ0aSdkDgBfIGiPTJHCqSvPtmrehDglMRdUZ9tDZiZYpFweLuXQdSL/9gn9b
v9kKKl9cEvSxn1P4ERUUWEK3inhp0w2BuI2USYiPZIwDwBv1DYZn+fzHGY1SwCAZvCWMiD8DU6GF
HlwLXiC2g3Fk3+aOc7ixMOwURZGTb9/basLUA+Cpd0NWPH7d9vcLwwRfuzKUwYphQQNxywXiwqck
zQAuJyZmSVk/j8lNxWMNpwyX7v5wl5QMDnIrSF9r4uv+U3YYm2EsJJsKZuPTYWKx58X26IWRxpu5
xfzn1c6zvN6+5sZ7Bj2/lvuFeUMM6OD/Et/kulgN8JiNxxZLEHkgeGn1g4utdi5etc5Lbfe7v7Xe
UEHy961h33YkCBjXn5vSyjpJkEqeudHRG7fIsWAKXbQ7flhvV3EWTA33D3YTS2sDrGPjIi1yzMnr
+s7cnHJapvvVpjDjoygBV9zUFxZGIF4RNDR/5EHmdm8JiJ6SU4qgXOZ6bfj9EG8PHbhEyH0pXfSV
rv7BdmOr54sCjaXPtBh5LgMJwTOzi8vCxEFQpy8H9+1j6rmERodiQtIpTfMRuibIj8UQfmesFMtE
Ny6HZ47gsrbvGRIrA9ECoqHDSYiDau6Z+lcfEMnU9JgavraIztA+jLe8ykRMoYzzJ4kusKt8a1/4
33oxdF/VIbh47c6LWkf4tDctchwleAUGTmLMpEfKtyx1EPdMGWHXiMDwao9dJa9pcOeG4ymxSS0H
YUWU4hMlOvik/ayAhCRFIzoop6dCExEivwdZbvvOn/23URXo2VX2IPKkAWZkSpEpP7ODyqyST0EJ
bf6MVfTxBYRpCDKKsjf8FtcYsG9RMRxzP9J15KgEEBtgmVHdz5Hw55D6WDz2lWlYFbjheuDtN3L1
HHxyF0f9954PM6+E5g0m3KletnAMQc3zaV9nLy+6Y6kJrlRzBCFkZLlTBGpDYB/gtib1pQ77Q6e5
VgberbEZHDjouL4UwqeVosMSArgUpoP7QT/QE0i5SjQ6LiEIy+CZZEIiNS7uE7tbyX17Hb5AFkm7
g8uWU/PGcFCOMhcRNMeTAMynMj3kZ/ZyxRFG2BsokDRpP2DLKdH4GkEsoZXLeI+xUAO8Ome6Ncdn
NF8sqiCbXNwByBswAcPY6vREfjlAaaO2GZFU0cAc/STeEljzQXxBetyE0TbakL6tl2Y4pRwpfgz8
c2yQI7HqRvrYJLL6N2+NXzD+Z1DI6d6M3d5145HxtVux4SReOf9w3zuCo1m/2l3kQNnzr4B/eNaT
RZPEot7IhC+4PbZTpkE5mJEKkLSHvCAMDk39GefUHysJ3Mn1ifZ7HZWmstFPFi8IALlmvhOOqdDl
1014d3ES+CQyH3RhtrBi2Uw9OzGfA33tCqiVDdr5bKwIvIQYsc7t75Z0sZxZPSAGgNKI25k8MAzZ
SiVe+GeOrj3vuPCdC+v04nGTr1spoNbbQTSJj7QuiMxeITyCAvB2EyA3OA7NVclJMkRHBkl82KNp
vv96CBttfOycGhWJ4q0Sp1riWtPUXh3yCjIF6O8o4xZF5/xULUBfrFgAxzMNUyzi29yambkA7a7l
zFKvbZi0D1V64zxr1+WFB5rQJ9V4d3Pb6iufKwGMAKk8DbWLklAQBbeoHv9iZRHWpRE3hp69zhms
/dA0dzqj4ou1QLok9T76DfcWtIIAzyho1zJf44LtaFjK/uwEskqvp9I+oRLQsQOjPozrXS6ebOAz
mXIWTowjMi89IF9mSV+C7BxXZAxK4AnZZWh7csrDJoTmEm0HYVKRc0s3oFYzm6+EoY7UEG0o++md
s4sZnO/QV/2VMyDsNX9kBJGjMX1Uk9gkCYROwuc1zMiLPL7CaHtQ3chFyrplY2os06hChL676bGO
/aA3jZj3Jcff/v7H8Q5c9nl3EwUwF85eu1/Kb7NT7GeKzRJjNOwr7KBb17pCdKkC/SMYEPTDeSH3
gAgShdR7XlB+zQ05YxU62CteXdUos9pnAJRm5VjCJBQa2CaoYs9dCV38JJnrUQs9/daDzkdQAvOr
pPqDEH78xMFe/Wmis/Vo9Yldnb/+fIzfzqM7SjkhWyC/1vGUpct7IzrF3Ci98lnjPMFFMb6CjVWC
XvZSNBdscinmmC2CI9b9EGTlk4xMfWBJwzHN4QA1OxjM6CCqp8yZ4Lx/9GfGt3EmqombX/gYQrmF
6E2P81U2e1Bx7YPycR7NoRKKOW3pfYNvNOEAXjlFp1t4O3ZUVRfepf6y7x2J+QhU+Vrtp/9/2b++
7wf9AjKe2Afh9GQyUeKCND7QIkur8Fv6aMQUcJ65D190ul7Fq+74tEkfIb7gPtrPgS4hP8ljomKX
QSt2AbK1V1Bx8BkUekxpYx3M3VK6Jk09aCx0LFSvdInS4A2gN/KV1tF5Gsmfds/p/G6QKO70AWnu
QAL+T74mnuSb8gZJQKZ8DZDnSgDwui35fjZw0oBgqBcfksnHwXKsGvTf4CtCPGNQXDU5eOX4wcWB
oPQ0oqHGZ9AbAICGPI/tClQKMBvtMsJ3eIIQycqo0f1iDcaxHE7yJJbWwL198Wnh++MU3VnsmL8v
yZMvk/BTX0ltOsiw2zPzr8U2bPKLIO7Ck42kL/curGWQuv8VvJEePY0iY4vhoPlLRZTxCr/6jstH
3XNTFAoZPwm7SH6y01rhcDNnl1RqQB6dXR9UUgdYMLj9qNJSztKjzaHx89Nk0dBSSdtZToh/TZLQ
hhrXwSbPEwE3UwgeMShxdDYkeG+P7qkLUnXuinC8zfp1gQRhui20ZHL6GYTiw21PgwfYUiJZlGYI
QCRJNUXefcbtc37Vyh7ElOkCMx7hCAE1HM8nqTlmqm0xFfBRcrV3C2uVCLsS1SYXmWkuzeLWi+qW
0JfPgUszV16Ww7xvgy24HGD/het+Y5cm8jF+IA87S8kjc93Nt9PPMlAL3aMgYs0zVzltQ1teE0L7
i4rB/ouc3Z6ITjwV1MTiSaC28bhCCUnM9Iz6d8Ph2dOGXOvPyRAME0ai+kYGuNurrV/uu5Z7kMOw
PY5YGXRQhjomFnz21okNI1MeweO3DtCMK24jIvvYmq+InPMS5zfz+uJr/rkzlKfEKrKiAPjgzyfF
McadiAWCnXRta4rhSdCRiMIBH0agquigtpP8Nk/jXNwg1b0tSNMcY0ql2MuWfOCpkwmvbdymG4ci
pE+w7aEEB8XzR8F6ZYLtNaOXq19ltpfwOxv2mB4FTMja4p7pY2Ia7U3eZohyeyHIw4dZ3C5T/tnV
8iTbMqKfaI/AqJZ4EaJ07oT21S20Y54gF5d9A8h5Z/QVGdvj7XEnn+ZmIEpVuRjXTlLVvUmtQaCq
y/ZeIyPL1may8mdO2BpPNHVk6IsK09qS+mfUQSGaHIAt4rixt/CPUKaLGEl51m0B8FnsoOoCzx8N
te7Ov6W900C+Rq0d0+7J0HVwYGtzLECzwX7gn4hEC5cEK+z+aUmeep/6IeGMTlsb36dzSPRxQUt6
oYtKAMzuRockZzNTt2H1OAUj/8IcIFFEwFeOWia/vCN1HYCIyyWNszoLAK9FP4Iv7Dk9glORzX5V
0VK8z6t01cVP3f6jJJrYUHuOom837/1TfQz7NIJX9wiWUXSVfe/3BTcEk1eFvkI16/AOF2lZ7dbo
0WL1HbPNMxWSnFscL7kz26pKLb2CNfHQCiDCxHcFnUDOi8cg2IDyfDe0xQi3Rzksa7awjG6Y9QAe
uLSgl1YqoN4Y0ucfIGdGZD9gnpsE5kGPJ0GbdknjkDcLZURr0/vOLLpBLeCBdtHNMtrBpj4Nf4mT
jJg9hv+N0DegqzZIhJaIm3TRDtvu2xyD7AAQdIMulWdMPdEmjqYDAi8OhxphKk03VCg3PY3Fx/87
HzDWWqX5qoRQx5O8cfTWLiOam9ixDKnqGcgKlJgnNEuRxcoQ7hXbKhinli93IUTJCBRNBFVjLD+Y
Md83+tCH83zzlf3mURjSXF38I/msnPbi8aZjVvW/ebm6L5REeh504de60liEdxYoh5VVQHgxPhAk
ysomdC1SNhLMR4fQRLwBlqpmHHC4hLWqFz5ebjj0YbQojbRFJV2YR9s3DVWclf+c6f0q3bpajwyq
AdEQYjdBiZZCda6bf/8jlMJNIKreoVhj61tvyqlr3HyCSVfPu/jeKtnxH+GqrrbrE1koqSjiVAg+
DjDcfbu1I8Z9odcSvLpbiq0Y40+toVBvFQbxWFBld5u1QYYcOokxkiEsRbbbUlB26CCfr+e2MKjw
CERJp5UARaH7HD5zLtQoS8luFnuYaWsy2Y25P9f8nv9F2v31Xf9S14v7FP/Y4MzxR4WtAxjjxF80
peqBKbUjSlc0lwtIq+8id3O99a3EjgiEhj19EwA4LVbEGP3wmZHVnAcjrR5wLoOqrchY4dBFDdlN
gjjtj7OYsLACK/gK9WqiB9OKMrD1a7MR2RGr7KmIQwtnxmGqXzsbo+kTRv3s/cOE2sg9/2vVpD6Z
AY1rmqRrKCAgtqWGu++zGmHDSM513msQlYv68jiD9z9G/z0UszVj5AnhpmME3OuPnTs1Cfuug1Rr
LbY+2AsUUHHJEAMBhO72mh15FXxEDCJeZmGhcQ+IBKKXl8NCtl/7T2zeg0n+xLHdo6iqVadJ9fG2
FeRFGs7P4Q1pR6o8583J8BkSpk54iL76Ytw+ytFOEf7GhbGZ8zTKBzqEURYi+Rkq4HNBEmS2Nboz
vyA0wPAsDivI1ZpUNX6fF06ULPIrTLIqbM7b0bHhcyr/42UP2UAziEF5HoyjiSa+ZNtntq1DQM26
Iz2mUqdJCqwwX3yNNEN2ACQwu/EddyjYl0OBG+Q8zyBoUDe3BneuILodmUNumXa6I0rXKajYcvkx
OOjstR6binDqHl3aoe1ndkaMQTCLDjQT5CB0fUM8fgGmKtCZUbaBLGevB1lkku/HF2bStxgoNqtZ
c6CGMgGgdS23aZWPN2xeIRV+ZiQOqB/UUVBQThhwQOdJZEoKXowrcM3e8DZTn/DNUcBbrnY5vPYx
gBjZ+m9f3DOWcpGf8T3XyDwmDTO1qQBRWbhY96U9SLc9xE7GTo7bdvAlJQGxKM5N/T5RbWeK6vMU
rs3pY6BnGrQIPeIIlpUg6noEhqV/hLpWU/qZhj6VDRZesm3UUj66RFlY+huH0mLHqWn63zpriLfy
hagO5tgMYh5hJBbwrJN2Z3v/jlGAHlwgBvCRkbbnVgi7SZKYkif6D+vWWKbtx5Lo1nbAxDKJJU89
gI84kDMxR61yr0cG7oKiVbJ2RHwGtW38qJa9VP5L0+KLcN4C2g1NR7DAGUsqRIGtI5e/214l3ozK
mf9562PkZ3/9wVDi0m8EOnZ4IFomHwVJRdEnb5rxwp/XMWvtqskPEdBjB/QhIdEWsq56Ul4VwNAF
HTBEPJlsbmsdwv9SgKETLF5Ouw1N7RBC5hGdEdhQdUcD3S19464fR8mq9Q/dPHVi8rAMIm53lu8l
gOybpGHODIN6IETmpefnShBkFbr3QX3SJ2vSs+ukUcjURJ+F1nrLfvEGNyZQuVBg/Qjk8jGV8Pvu
p7lu4j/oEczKrR/+YiFjsiroDmi1ayEsKa+xKD28/W/+nct/ZZ1Pp5TzUg+Ncd1h80LGVLBPQ7TI
3HJVw6PRJvEEEXl2CvnJ8na3iuofaX+ZdSVaXAZiijm0GP8ewwLnUU6Gm83ONAVKo+ShdJB9zoEJ
KnfvgJSWAqAYstSn3MOEVXwATIducCN4o18gDlLqHtgmOZhiUCCgcdQU4idcm7JEQS7MAAEw6ELF
n5YZaYJIVar8J0SkdVYwy/hY69LFe8Awv2a93MpBt+5JtOeB4VPrs1uDfiOBS+pPBa9v81q1GTxG
otgokoqRRxyC7eecDgCPBOdCAPQvFqCwjVkk2lRVH+dtuksJ0nTF8RIXw/1AmO7DzZLr63gtKkh7
+YIp4SxpQknKPH1nHpO0NIgtu6hljRnQOReHeoEIZfWxoAMFvbIKmLdezfYkNt5yxRcZ1rNk4AmK
XDqRXsJZX1TZj6EnmpfWxwBA50/U92Ba02IiCE6mgbo7g0svOsXl0DNLKYk/w7Ae+LLO3bi3wvME
G0gGeioWLcKKeOv6+QTVRat5jrZL3h2l7EMpja5IhoVKOiQaP3Jn4BeBVNcjz/D7JOV5leBj9zsp
hPhvVSGrdhe0CBnUBQs94qqr44VqYAvSL1///bT82GbvxYAOW5rH0D31QTmGGKn09tpQjGqaoOlb
g9Sb2bK3dmNOmzRxIHTQgjJp8lSuaL6B8ablnkGqU63AlAk+xbfYLYpKLqkT2Fbvg4l3f+JmY8+7
SyboRMgmfI6OrEAfjVu4yKKjRuzHdn8FjlruXNkCxhMiLRtr1zZy/rn30Yi1xRix7oUcIHkNvzW7
INGGQTrFRfPCkNQJsEqvKl1ahoLQaWpLXRX+jKjNRT8fVeBbwHYjLqrDauQUJgE4vPNjywmKjvpZ
I5n4vzKJvpT9cKDXfBGAm0e5GZDp2x71fVsPGBgbiMC35sQtc8EQra2GpdY8pnwVJBrskKEWNWBv
//HuCOwE8IxU0R3iSLpKbm9EBKUGuwgaJ+HS9B1PilrnToNIt3yB/shTGv6+aNlK5q4kqWb9MsZ+
+NT7qjmPpVnZ6tTIgZCDKOD4oDAfSJ1M0OKYwi6xVHdAqvlcFdwe2aQBBXHzjtHGvqpgOhzKf5iM
H+7dub7Mj/FCH2HCL+TkBOWwzrKj2NsLooSqpz63+GwiHFARB0+c1mTB9a0H0vztc7ZydjpozBlp
eMslbXXeFNW6J/m7jUuCTDEfFWp3XU9l4WXRGWQMyM1/5IMAqwBpLXDNA0RGrTC69VlPhN1P5d8H
cKhzlluhsblbdskw2pknz7jHt8pULj8oBhdX3DUWHmFRODU0s7Fc4v3a+ClKfNoqYXpkCoEjHLwU
Sst7qk1+mlMUViLpV34fMhgsTQCh9TXji8P/hgv04yl/ptOF141Brx07lBSIj31NLh8nNeKZeqAU
xHad9j46MYBxjOqB+zzQycUyUDjDN+vYoXRu8g0TmDrj0h2Z0Xa20MnXE3ZrGC0vNcRASBPCyIXl
wCWWltKMc3pJatKCZS/wZrNpwCteiQlAEZNJ5KG98a9rxhXN/e0ClXqXUfFvvTYWnP4nHaBzhKXv
/jlT6x680YbdL3bbTIb2kAYrwfwLzaHa1y7lU0znoLVMpa/2uOyXaLbifLlgLGy6btfS95i04B/s
fOjL44AqQCIVdQBc0NUb2nul8h2zgKgLFPtkgCHY2ZRC4/zbvqjFgertLxdbVBCUfMNO9YIr9BQB
cUpVcH3gL3dRKv7A3IG1JC/68Ao1EqIBFDwrk6TNSVWPapONf4e57X4BLNQ+YHHv4+booAK4kdgr
s2AOUCz62mNtqdXDZ7j3geHUeTpommQmq3f8RAGhJVYswx26rY+QJ4S1JC8ed3DXZC6jM1xH5cf/
6q3jOk+8M/7UsiiiRmAa5EQ/94Lbd+NTyc6P2FwSRM1M7HbTW8D62d9Y5b4TMTrSfjYGuO+xMUXE
M0+MQ4BT1AjqFW9R7Omnu5blAP1qka3TLslNxSgC410zMA+UNav2OEs1Bvt4Y3uNrSjahCjDtMhV
PVnGxXX1icieR4qk+KEDnX3/owaX4tvj9gk1bLPncN0m1WeXZjxdiEiDtmHubrQ6NmPvbkwrKQ4R
8nQnnDZTm8axZp64AxlSOfQ+XPhhnvDe0D8bF2L43HL7nKB2Z/NFcTH/lsH+rhkc7QEUDesv/73G
YBq6vOgjhLqoVdMejL88X/PB4DSqY6fzKQSd+qcVJvL6ZW5mtYhzrLGhJUjeMLnRQ2NxXVUL6XoR
CLsv0Sd/Z07tK6MF0QylJKrJItVr2ZrSVykpp8vGo8D7fZI3gfX+NgZW3gJN12f9vEk9S+nb918+
HpSEPJyvzNiC85MzQX94mkN2O6bxEmsckqL5Ac6MQLM6k11Pft3xho8j2js+Q3KWrGM5bmucBB6n
v9z+/aJfP4dlA2cJB7t4JUx9lKc+KYP+5gapQVIAdm8hS8+idzxNNQmyPiZarz7tszKp8f3NJQuf
1tDjQPfPyGZ+2mJ7Ywh57xtFqGcSSXET0ley8W0Yc2weO30/doznhdTeqZIcxQKcbM/QuDD8FJ1n
lZdhDxLNB0ehCFJQVH/T6MoW6HoadXh6l8CtKNjGZULSBAsnFB4TbLjngZzcd1qvoIHwyA1Hpnq7
J4P7GhhwCG7ynO17ULjgcigaZm1temxFF7g4MXaCA2D+eqKZwKHW9E74T3pB80LCcXzP/8McEnuJ
0np/r6qvTs4X9xfdQFZW55o2JPAgURls76fUeZkgqMGjRTxWEX9MhFHEPGlxZkEj8PJBstN09fAz
X5DIsbKmbOUm+4tMYqRGcrxXZr6kuLmf0VzCCg7D43jF5YIQg5Z8Ytbon+ArginIK36MSryS9nkI
EOg26szNYY3pCtlNuTkaLzgoDxad8GX3moyvB2Olokx8WYGiyem/k6bzi8RuNRmV5cW9vACIoj9f
8EDtWoeY+ndZ1VHA81eMoF8xouv749IasfW5vV5wPViB4x0Ebj6OA6jPd/8cu7r6vW201eWlnR3y
P44mYNquNAt+7t7ZH7yBhMhDs6Omg7yhMEgfW9vk71m+L24jFW1GPG9eIEMZHZWOGX6NZ1bf3Mvt
ZbTq4rlNVsRS85lL/dboZ35oE8zU8qYMo7AF0VMER/LvwtWKsUIm6qQTozpj0YAXtVdU4NN5CT9M
gQ3z7LK5ilvHGU4v3AhZQaLxBjnsb4f71Y4LyND3dwfbvkKQ1yMnwy2Qu0FUxLMqgHgF+H4ToINB
b+HdOg5e8TzLz8Hz1RwJACEjXNfVzo2bMpBLdDSyoJs4scfVgjH5m4MmLTV36+26AUp18tvx6ULs
uVf7YmQu6I5nxyOQkPUGTzZT4wiigNbqs3YeiXbt1RKPZZqkrprwvZnYSFeoBczBKGQVVBqjB25X
2NqXq16OggB1yNWYzOy6cYorlCZ7+ddtIbWb+FvBBOj+t2FEYF6Hr1bI9NwFsJtFHfQAzciXPS33
YtUfw9SovU7gcV6JqwRyg5oaQ+x2AFooCfO/Q1pd6mYNGzIMf9+qOYZxtv5Lb2gD3ezol6SzBEEg
u6gMKLNKGfdSjoGZUZ86zUwrTugOCpVL0NneG2AjYYFhyYL7ZkKgfFJL/KfyE6hGmLW4ZP+eINcA
lFUEdPGrQe3psne3B1OtnsFeZg3w83RGWrHgUZeBJ/F2iDdf2EPajSWb2Dnf6E67o+wtQOvZxrfk
cqIFjSVJxt8DMjq2uIrsY/30tYx1PjCAt0nMX2fCWUm2B6APAOCyAJuKG5SaTL2kqGMJHeRfCOwv
2MK/OLggC+N7LTJxfi+91pJCnLoRJi292wktahKolQVgwrcHzcdVJxdk+9g2N7BKUV+guvYGyZfv
g6c3YwDivwuLMhZzHjV1k/583wov9uCc7qaoAhhs5vfsKSAn/HBBttjHcSgYIyqAmcwkZMLddtaT
CZIRD/S5qBF5sslRLcmZ8O/xMD9OqbGeDM/MGUH414BFtrWKeSJ5sMZrAbBUjf6H9dmTvZomrwN8
XhKNwZxA0tcK69PPi86cGYd0P0wi6LOh6HUo8EyBaIiR+0cjIxyTszvyFolNdl3QCnI/TmVny//i
ca/bKDs14LtvFzwIXIp02w6grc4rwjhjBvatzeO/gP9dSBOfyDqP2rSPfaqVDYXVT0GsgvXn9TA3
ZGZUEsuoGL841a5mriy3zTBPOo2CZXYakC2xmFbT67oncHjS/dRU91ZuoT9K1Og6UaG7PmJNTFrL
U999ce1WM6tjgkV8Gl8dathGAFwplLng4XMbrzsUs8AzZQMPC4j9NwlO3onJsbl0qYwoRS8punjm
W94eYGiB5e9srtFxVJGHtRiRi8lbGvtrO+43Ee2mmOr+H7UBzpY8Rhq74ml72C4pHjhLLf5z/kpZ
0mzFnFe+XXY1AUVXKSW6dk0Suo3NIHRM//R4RCK3gFcv+bV0kLm2WFnAoqyuQDR51untBYHGINL6
Ht+aVkT0IRvG2FX3+avJswp1u88zqR+qbPOAJSYtqisbAckMr27Ktq4wka2c1mNtMsCha5lcZbdH
+656c4LfHe3O1b1j6K7e/HxVUUA89pBE9/Dvmm+Jm7QB3WLnwXs5JRybwW3i2gPCaWehxoF4f5Ej
yG8jo8mrOTLoKeUNd44sTycnUv2vGKjyt5ciNKTLd6wbE/3jMZSB3fU+r2Mn7q4Qbx3vhKI7Zo2R
UFuj8bnoaj4lqaRUrAPy8G8Z284aEM85fbBOH3vdUidv/BZmXPm/2WkzANph7hWN+6FP1QkC7DDx
akT42YQv6FoDkkb4dmm0YUyNvxFQ8/XVmsP/5p4nWv/toaS+cb8O4LV+J0OrL9ry/13pYowc7E9G
NA90CPPXhdQ/a7YkRrPwrHOmXgoWes21QLZ7nqvRrirp7NgaOehdGb0rBYVY7B4UP+vAlwo6nVLw
dqRpnyYoFu/822MaBVLKuB4+dLl/bKVG3anAaQ2ki3/6x0N3gfuCXKz89WrpVVwHX0+mVNSWK7nd
NgEKf2SU5gH2EWQP3/acvGdiTKlw0KCDxS4DFbGendUSCOZxqR0gB9sBeisDW2shuHbezWHELRmD
nVfW3jdekR1cyhI57qbeTYgrJqC/U5HscG0Dcf+wNePGzL53TCcpVK/fhicE33BK0hEsP7B1POBR
19Uaf1n7H413C3VNOR2GvAWgAIDssJL6/y85CEEuUoCHrQzdwTJvQZ5e81oKqecQlIdInybU1vrr
YRpluiX+3v3udmc4lmH/3yCC3t2M83nd6xrCFMprMVUfRg2j6kZE6d2u8djzMUH6hHQeJdJ8bagq
iEg76BuPoA12mcAmKMejuQFMVts6h+ZE2w7Iz/LMLeEVfuXqSsnqPmawJPrQJTb6nuntuRbtKYiC
A5/7OnGnhPrnyQLjLX5SHkh9xjBPWjaf9i5oOUbUn5wCQW1mKHyWtmRrHzPDZPsuBIHI8LKZbXCB
EK3loO9GOVCT3EgCDQO0RhdwSpA7CrzzFMh9hk+BKKX7F6O7Tbj5gcnvE9AKG5R5MUmcZS+UAtlA
/gNTYxa0kzB3IRW4ESLCWHojO8DT6zEFs00GuFswzRfAZ1I6zv7ZB4+Nc7JHG5fg8s82O+cxXfim
+fVGcvfBN5tlAAOrP4jI6cmbsMkDJcKLFFXqOheGWzcsgqvm6eQ3Ex+uCgISTRsb803lcioIy9PS
V6dBhQ2eF8wd7ApObe0TgJrQE3JPaZ5I5ynaOA2WY13wxU3seGQHEh2GJdX8+JnZ6wHmK2YMOfiZ
cZkDOYMPsJyT0wu+Xe2ayaSmBnqctVgZwLBsxYdBe8IZj4emF713+SKKcnkxm1n+acKcJ2MTBRbM
2omgwE8k4nvF/tIo2tBbWGFIf1+lul2UcjXT03uZ5u6kQ++TXOyoNHdJgbnd4OgpfHx7I4lIhlzh
bNrLAR1LtNe7KCiMuK0Ec1ghyDMbDM+lxCsxPq5esxs/LwfvmfLXjP6LZWGqnCjzvIl0dhfKgt7J
FwfvoWcep9dLhu4pvLd1Hlck4Kor/Ax0/dZ8FjoDmIs9r0PRjVvuHSiPN4wwRC42bssf47/kV/Z9
gZSkE8SYZC7X3VenXgnNW//K3oof37z0EKSne10Cl8nUtz7kBSed3zCWJoE+udKB+SopYtnuUDsl
7q5vsrZ4Ld14Uhcsu8hnrbjhainCtCkGWqjoPsc6xdImMuhNKeC219KhcmIUvD04JGYP5g15wwNs
gp/48hwvybEYVSlLdxRhx3fKK3V5diFi7ZQZjSfp5CKnAG3OCFysrbqsI2XMio7aqjhmqi77K0iF
UmMnexvOHLPBJSckdjNyhxBvmtARuZfaD2aeLz/ErbqQB2P78Taow5+usDHJAXC4iHA2+TR/1JPf
pvlI7T1M9cfGAKpFDyxLZf+gr730IbZElQD7b9qXQGbUKU5r93vaNwXBnQbBoC7fBX7o/ILl8ZQ5
g9Vs5ruChpoDA/wVPS62lV8OO4ILn0aOYVa/7PafNmN09Qg6VaqNarpxRfeEYt8pOEhVUhhGnj+x
2eeF3c8o0frENBT7+avmHgJzZZIVIK8luxiluzcVBBVOHm/cRu7KR5PCJbA+k2DyzlYvMlR6743u
V/h3hk5mH725Btjwb4/7kX99sN7y0B36HLCSTdJdBkmNwZXk+4BEnU8hU4D7Jgp3go0crvZzn2tZ
YjrXPRTtAztZMc6Ku+6N+hanx1v8Dm4ski2sdnFLV6eJNRhxNubUqC9LyNSt0xJ9dPfQenBKhtfQ
AQVwnuvXFTPpTq/rbB842LyPGPE8H23dW0leYkwBR1oym7oRHHu/+6F5t6jKDQfrgcJ57wRIFwne
+mU9abhPKgGqxTMxA9fO2EDysqVEY8dOORDHtcX2Wiin8jQHMbjJLsx3ifRBYtev5NsO/YGmY8iS
M1T2cEODCYcnz5aHeF9NyoBccy+uSOevNj6yqqCVtZ37lWl6S/dG8iQJmvVApgiLdzEqOrype/e+
OIDllSBUQT6WfoxYy3P98L+opClAZjadRkllokJyz5E9DLMrPIA9x4dU7UWTEnu0zSbp2LSR7/Kn
ng1fV7EQLHxtoiWnZFLXgqFHN1/JStiOJL7dYYTUe1RgNN2s/xEnTFPJhAaAKLq2Ppxyla1hELJv
8NTYTTlXxivc1aBp4Ye68t2NqrIOWa2IFwh7PQChFeE3Uuk5WOlzZbs3CVnFwSv2418SX3yj6bqm
Sf3EN83aYgUA4mAT9LeonWm7Z9+ZA1Qjao38zlZJRl8QLZttH6dgoFQQ4OFHCjhvQCq21FbrB+9/
rxAvI2iLt8mERDhEi4o9I1zOcgqFLdHr5QePKTaQCjGSOy7jsmmlFWcKOozXLVjG2MD8teKAQF4l
lCjglbwNdg4vqhXoUyrFotXmTLdfDhW82cgyrmgaUin3ecWj6FQF4WtiJpow4WPGVn1v45ZBHz/x
I6tI8DqtE7FA0aTkXcmMvWi4vdi3Kw9nfChmQPKS3tmqscgtuskYBo3kK2F50yluXngJgHImKdRn
Ne4ilWoyfJvU30pLp7fRNl02GsG3eag/qva6dIpEL1f6BqmHSZDJ9olufwy3FpnpVr8/6c9BOzyc
OTc8C6K0Z/Eh/H9IRWwuXEPFEcpUK7ouizwvPC8Pf0w/6j/TA2aVq0RttYhkmB1/NPbu2FG+wMHr
TmOoPvv05NG14pQmhaX60a5XQo+iUJxBhnTV/esLylalgBL79FN+ieXFyfAgUeSF/dOfDnljZ050
Fs4GBiwnFZmUSX8fJuryJEIoJ5ph9XaKlyvyEwlCevsjzsHa9Gs8IqiD/dscbjoqypplaCH9PULv
r6uBYyiudKn7aJzR/Rau7v269/fLLD+wCkJlZpHSseT07cUxAPeYqxlaScDs7de5hJayBU+LQePd
39Mp4IanSVNusBu2PNFVvi2loFUHzYe536tWsHZhqudGUdjtmtyaUen1k6ZgbttIEV6A8Jqh5pa+
ODxeLe6+c4eB70lZ6I48A6QriCrY49SaU0HHfr4+ZGvXzVgajIYqDXCpilSUpFkChMdrEQeCWcoS
hsO0qjEgF3TY+yWXpDD/B9h8bgDJLDrsS+yKd3XjjTW7CvI/SObBcSbqdXn7NFPmQqjoY/f3jnwa
4Rg45BT4T1H4eKW19onoj2BXn8beAlDiDJ/AR83mWd7WICkr52sOFpYsD49dKdYJl2F6+3ou3WE9
YpkxqehQD45PW4/lwZo6Mov+vA1D9QC+CTMY9QEIQ12jmghs8+LAZxDVRay343gD2u7Q2EUNZlkb
J0bUEoJewh8pHgh6IxLNA5sQlbUTZqQL3QTH7bkUgDafxnBYiPlsktfYliHNaZWewZhHtrdymM0/
2ZXXGqinkjFYd1djj541Hvh7N1x1UccJhCsZQhv/LrCzq3cPac0H06Ctcr1wtReftzesNt+kx0Op
uRY0fNQ3+pP8TnVXYw4qI4mHehYlqu+VjSzeG+ktKLHhvuaiKWiXSzKEEdOtpl/GGDYDznWJjUzs
6/Q+JA4KyEX7tlOoHREYuy3bqY8dov6wfVbuakEnxUv0xojQe922Cpma4YuHzhYE3Syz7DTQwaDK
2P6Fv8lRuire7NNuf+01l/O8Xq7yLZYwi+RQoaAiPqK/0HfoGXdryU7HL1V1YzUEpuSWpPVL7BrK
TzZSwABY4imNUb0EFxAJuuuSC90pNzZP1dNKIDb2YZdjzHHY3Et5tWVcoakYLaITHOKE9MdKj3Kt
XlZnyX6OMj3Teoai00LFq5u5P6FCAYKBUh9ZC9ekan3O8gcl6nh3myBa2nq3YQuXnUSfgV+K2QPp
egV5ftGfPpTP7OYaJX4A6U0wd3fG1UHEu77YNr26R4rE5AdYHtXDOZzU+pp3vDU2d4k07Ki9UxDx
56VpaZxaKS03EEmU/jkcJA44qNrk0wnru8PLJFPk3reGsspd+WMPJs1+pXFE4qr4NtriXNr9If3y
A2ODuuv6IxnGXYqGG/B503BExg89s8lqsY+6PAeb+kukRO3FoTP9+w7BGGIUzmMSY+uzjKOfDdjJ
toMLY6JvG5BUdX/LcB8fCp4bPg/QODO1EIK+9js87XZ66scWP2Or8VcNfOBX2A1kEZ2BBkpB3H9A
+KDgGw71cbTj3rxoNZduNJ2fqdRSBec5MOPzqQ82d3KlQzbcyKPpfkzFn4E4VLObpwrhgOmidwtx
Pf91pjydf5idwdxZ5dHFXFrEwWfA9OWlP35PY18LpxDwaaBU5wBfEgnVdSfchObZT19ed6caDgXX
FxszQbl0plmxlrgfz45a6ZBK6SxZRGYIHXEz06EOvI+5JD8zHvSuQzXFEdZ9Pzp97GMEXkRLggqx
rt+zznOfoFh3yIa2EuldDgLgzYqheKh9BlXucUyE5vmg/K3wJa84P/KyJl7etY3pCGohvcOAbVYk
yKCPVmSaXUqIdb7IIwChGvC1DG+uLNkQwAu1i8caIhA+H9d18LYQQ6JU4es6IoQ+zXGMHfYOx3jL
eBjGdbRQdKtPb1qioSuV5FJASoTGQEsoJzHQmFspAzmPdEOnZTMRrLOEql9q8hLHWGrdeb9TYf0A
swARbwj0baZuUOmc1sNaK0Twdeuu0wQp8IHzRTIU0AUzg+PfeJEt0/Sd5HoVkg6pro6PseR+nUPK
XNCawHVH7yX76rKcMrkZ7Zargp8141mc9WdMNU0k/0Z+Dp+xpb5UDHvwyDvfi9gHvLG6MBZ3c1iW
3Cw/p6roEPzvZcBNQmAtJtD6Gqk7bFtHEM8ZGBJk4zZRlDjSYbmX5uP6uip4kC+t3kwLsGX6bHUX
60nGd3uHkouh3q8xyOV7EX22fnJeTok+WRIzeDZJ84bs1NI4quP54vsrGjqL1JW6qV2rlLjJczPl
ahzhKf5uTkH/MA8PXybw5Ic4QctUSI4GBdrJqCKjtnE3n2jNQ9PvaTxeNHqtZMQXJ3YU7rwzcwbE
hPE1Abq7Fk9Ng7VYaCuUdsAAb34hKBm8HVlDKFT1/7ETmW2rhjOODp9gV4BW1oSct0wzszI3MqkG
zG8G7Cbo4YDlGy9hTgE+koSTzDL6zNJTN40U1I3J1Je3dObBp1d4XNc0p1H9T8VA/OBeD2vHdEBG
sZhStQTFZMWAV0jNzLUvI8UR2bQUxtogMSwUXizvb27f6OilDuZTbkmwFvuwjSd6aCxH+stskOIW
uV4frn1wFcCWGdX86fLGh1LrhKxR9J/RydNNjuJS+HfF7QLMKgbYaDoMMnrP4oFF4Bbq572tl5td
yVeIlQb6Cay703xYw6ufl3ploD3d8qDQ4V1mEBsymoQ05yt4Lca71xR6YDOUBYiyvp8mxX8dIqNf
sQ43iNricIuv8P7DqcN+k0OXWL0e7MndFARmOejzBOjMWp8+V6WckSN9pvrUhVWIwpGFS7jtzxis
emGU2TF2XHiuk/llnRvd4whbNckNoT+0VKBSWhhcP0xrFJOZs3calLwwS/QzgsO2372WaixxNQ+v
FXZt+SQkb3KKL50B/oHYhFyLXApenuAQ1dt1pw/MmY2dcHWjX5QSkOb5kArBHRlqTWlMZK1qh20u
W3UWBSP+6wkiMca8inC/BBfQ9pGEuij4M2nW7m5pv1b80G1CUik+1dzSbkjEdJNbFAQDQpqWKcbb
/RYq1bcJWx8vJDeWyHBxWToKlLZSLXyjlaLxgmsRt3Yir1wVtw0GVI7QYEzeE0WVbHTyU6dH4jT1
aw4yWDvLuYs9GasYsIbSTrzq2pOSpP/VYbOOq+VHqnzsyOCvaV1i8mprDyfNuWxQtMYHUtmRSVbU
GpzV62F18JmKjn4AbcYyUZR6iD/t9itdvLDHVtOBhlDejhWGZC1GkasrdJJ2JITflh2GbL0q+kUs
ars7I65RUnTi0lB4mdUa08PtHHVcxTOv2I+/Yrfh49/dVBsWmgwwOkJcUv3V1YTmzfg0xDqYFmNU
7H7RwshQOTlpKlPB/mK2piAnM9d4OkMGkv2Xi8Z7COaMkN9+q73nOy9uSN88MbCMt1O1PZS4mEnF
djKCByzOqjL1h8epFc2r4eg2TZ9yE4qW3QWmjn5/V43swxoZwEs6dBmywJnhuma8yGbKazh895O7
+q+jbJ7/8Vb4MKmoM6ggWkRDJJK6wSHTI9Tc/apTAYrGb0+ttqOSUwXSmOACeP2+wHEoewNmT/0O
Twb77vgAG6PTB+ITG1IhoDjKJfBbZ5HrhCHvhJ7Tl32dQxj6JoYZAdNVDmINrI/m9SiAq4RZcr9P
+23kZTfvDPY0KuqmAQTfqwsyalHi0Xkcb1shU12vhUl2QapXj1ln1pU5oHYTEYFj970ntgpmLGr3
MU/S3/pjtYDcU+KfKstMOX6xuFE3Fr5CcHXuLwbd8IFR/Wc4LfnvXDh/RkMmVRpOASm1yczIjQUG
kqKjz1Puq7B+k1RJ7fnOCuGXBka7ON9M3kvBeN6+OpA0CFSQ29Q1tX39P1LfV3LkkPI4db2xmtw5
h1W7+lrb7LAcep4VBI23RHbguTq8ydFIM/Bo6T7R0XFXAy95ClBeeuuEwjLMAPu6Mor5mwqITvT7
EdQU2wv0soyPhB6byHDx/a9Pl/wb1Nvwv0al1p60i3d9NtZ8a7DyszXxoFGNRSfE0MOYSft/Rmbg
YlvsVDqptZRDiXtnMY3PWaexp703GjNVOZOyYoDAgVLoxCYjSXInWU7qO5hGCPZp4cM/pXdCuFHm
rfbJacSIf6Cgyp9e1F9N8Hy9p+up6VWLokdN+azanUItTZkTMxyJx5zRSEVmrEa7GWy7wnFsc87d
LgOR52FO2Sx9ITHhqwnJ7LCuDvjqvzSNHVhkGaAOH/PfMun3BVdr9O/yVtYls2Vzm44+L0nNhEKO
CWK5X/Kk+w5TMxNC17WP7+vYGkqAKc3rLXdc3c+LHwa06GvvJcV394ysYcGI/nM7hGHdZFdi/hUr
XEmjYAjTZdmU7x3ge8D2VyYBZetf3z/wUeSb9Ml5v5AuXIz3gyHzeekefpZjZrYkrDRLk7r/U+xU
VaXk8yjVUVImEIajv3WUche3N7GLPOJkTdZZ96sn6aNhseaaVXZA4ZmUX4i/ynRwpX7sxif9yvlY
0mUOIpGX4DZS37B61HwmQgTEDPxh6dIeXQ6Seu0OQAdVs/074mqZx7Uf5rETYO3DHPKv1G/Sn00S
EfDxR9mZj5rjwQeF7rLA/ZiWmT3ZRpWkpJwAt0i1KsgtZJ8BrPAB5SEFR+TH3L+wPnIp45sJlc0f
rJojvMYqx8tpse/rVzdkDh+rpeifOHpYD+L51rApMbkBoIo9XmkFGnuUQr7ovgMTt/bqMMqU6Yd7
0N8u4+drnNU6qeAWMFTYAhpzohM8+24SKxzR+ZH7oCGx6vDLxxBXmaSnmuPAznk0PoKjNbsNzmA+
oG5ajjcZ9/Ar4MjXX3vgPOM9jB2L19GB4KadJcjxpfbV3tsI1I8fgP7/633tjm3MMny7+8/77GrM
S9d597TwRiIYnC8F1oxOWkvuSqFlCwdiqsfR8MlCYvKgKto9FxteeyEdjH5QiYLJu/670fLSSYTg
JIVfzHxm6KNYhcTskP+gWEbinu4CdnG853ojV9pT+rngHOUFKxzkv7p5V8CDTcXdUQdYMFm2bXDv
XZxMgdWC8yNzJm/UcRTiJwI2Q40Fwcf07HUaZl9DX8uVdUVBWi9czcOitM1Ny2VUdN53QelDaawD
IjuO/icaC4Hn2h6dqJxbIdnKw3oECQ8l5YILOK85acFC4Rd/qXb5fWfzSpwItWFBs39zFLqGlgx/
KuFV5hCFETLOo+oQxM+vDi2c8pVpD7orb5Gqd+pUJwtBTQ8+sCfEWBxVCoxIgSxA3n8r/AZVbi5d
tqrbgkyV4+YIEUfUnwURERQ8uEETBTA4e46uZfORcgxyrsrJElVqTYMTZKHTVJcfGm9YuHXcH42p
xnCQ4jIY72rv6fZucHgFRnVVNPaFtVz+D496yOQzRtvkvUOJSzP3YTRFJuIAhrQSqtIlP4mnuFWS
fUEyswBaIgNz2jjq8bvLq0RIU39nAbWOmCebNf3UvXFQR8e976bZ+WfUdLWf4V6XWzu9am8SkS5Q
qI6FZaF/1cMDtOS+A2pF50xC30Ewwfmi3r5s+Pyydb/EcFsTAPfYeX7yid4xDz1T781exuvs3+VW
N/h5NB3YYLAIahQvkfFhV+Q9dwbEAumXHbnUDnJcsJSiv/gKaUG4PAZaL010eZZ8kXGb2CGioWex
AYGMM1YCqKyz16oQTSxGKd8JKUIYBEh84+cx6xuL1stcrV68iSnlfV392rE7bLn6KqTn7hiV9VF2
3SKpUu2SSLK1PBs3U7mWyaYrDFDiQl1HwWwvIJPSMTI4eds0wnfnMJgOknnhD8IHwZH/TkGJ/xfv
LZyiS2HhmnlL1eqWsNLX04UcUwZ90xGnwmVCs8LAHi2x4dmCUZoj087VEyc95A5WFK4fvRuEt9Ko
NiYwxkPZD/qhOYcewAa9zHo3yCppIHZKQOp58YuppGUpa6iTVCOuZCOFDlGNnuBJIgU06My5NubF
Dma3Xw0yN1zC2R5RymEpNkI2LyieaTozuxkqBQQ1PqRIQNvZLydZccMJnnT2CT8JTGTGkPbyvxk9
NV5ypKrj+Ap7ZB7nGCQOm+FSCw4c+km/BeHLMBEswtx9GvPPWcN00nktdNEz5k7rTvq1cx+HhaUj
Hw1lvOZfC7M6s+OeukKPHlimpEjAww3zIr8K0NDGxK/og/3uNtRWfHLVF1tnOXDTd5jRywJG0Ti6
0J817uQsdyf8zHHjsXITPfItP/lYtdPnWvpc67Hhx14c85SqisMR8h/GjzsblKbOKz9hd7vvm7dp
Nkerq9UXL22yRXmnx/O0jKEP/EbVYUkyhb+3NqLTQ/AExnBMZ129AoNvlyGvdUWeVoJsudr8rzOj
WG0EHKcWdVMlreDy8p8FYpDy8IeX+yYfh8WxLiWrRbZskWmDLc0D8CryY2ZDfbHElrw0NX2nMW9s
CLTkmkFYCsQDP7nce7GoKAfsgf5BxR3mZHV28081pb003J5Xxs5GchZedm6IDITTmKK5qZ0Yjb14
a2Q3gYAV0NJ6X0E80JtiUrPbrS7bKJikatKHaZyDh4Bh9YTu8moTaM7mJz1tJXCiSMBxFr2zSuue
nL/UrxSkuo32l5ofRRou1n6nrbCnN0EX7gAO8FTO1BEVU0WmSDrU/zXYe0UPJgF5rTLxPjc22WfE
2viSf48Kq3NB+t59Om0nq7d/IR8AIPY9tiU/ENDG3I6GUSFp/K7hHMmn4y6Lnj4a0qdfTHfDZ+vT
GaZnsAjNg2iG+A/mPpka1llTrEGw5x6nv5HcRSlGDj/jHCR1vtCGa8HCf5A41aDe6wiDANMsSYpy
qjvMuM5i7XApj0nzCeivCdFSlKTCZtP1NWnRlXw+E7OYTwlWKV6qzQPWDEKR9JUYhMG0xSHQF39O
S5NyI1T12Xy1EfpeWzmQSfDU2kyvOpCvxScb+mZfrAYZlfPO/igQh8+cd+hpFpi0SDzyLaYFx9S9
FJxY9+BJNamBqniThKX62lFJwaYAkTyX3A/h6kIpGU+Yw3cwUAqYTT0bphpi/7GBA0qoOl52NnfO
8hCV9ny8A/n19nEr2SMvZz+kbiEGF15E4IBB2MgeZSzlnZvuzPkhIFKlFuAUsOp6d5B2fPf9MYT0
XoKGpXal9cGCyrWsyFRr8qI0HlpdplCRl6KWYIls8TE4g5lFX6UwghQfxO/UhNzpplTA7xWzXHJl
wyHg8YfQV3wzTdY0YICNp9BCVWhIXzVqBx/QRedGDO4eabuO4Wk+tpi5JAnEZuRt6hYkHZLnCw3N
Pg5sM9xZE0WUVCInDNqczAK3hbg9Or0C731sa82Fuq6CeHUDLAfiqtdmqFU+f7egFRvx1CLe6F9A
aed29lbterjfh48FeAzqAXDh8oZ1iGztVww/g88LHZ8qc1vlRdHd5EFGlZpEf2FMW6ke7Z5w+ytQ
9TIi/JxrjlMEFCYkTe8+Rc8xmiym446aemQA5AeV562Gl3vF0hJLvBfHrcWDUyJu/o7whKV7l2hm
IxJRDjqaIgrtZRjljfMn9rreG2pa5rDHq5HEvSaDX8ayHpl2BHTM/7y+H8nW/p7kmDM5GHDN5CqP
WGUCFhlvNEqOZr9GPVWTYLNVFNlh4IA9tCak5CSMHMBw1LhME9oKUFiHjHDQsmrZWPYI7DsZ4bKW
v8FjfRToOLMOK8//XJYmjbsaiTllOwFPYJPzuaf6hOaddegGt3qayn6DmpmDMlXNseoNqQPyQYbc
KeAuxjkKEyLVBq31YQXRGFezFzMHD8QV6qN2GtGZWvRB7PrWcJ5b+lv4mOARj5CiKMa2bg9izt9e
za5oi0749ertNh7gBpn2XlrTB1/0pSPIi1n020I/YvwVPp4ahkwx7pGsRikFWwcWiqR0TmZgtf/E
+wT6c99Qxmi4kwNIDIsgP1wjBaAl1EiUjwHS4gElqWiT3wgBTeF+ogTevB5MEjZDTOwW9OMWIVoV
3AT7qR3E+iECn36alft15cCVVH4RBGuUyrtxdhYFwdHNQ1hsmNvG0UachH4Gfw/ZkWHxIqD/NRp8
+7MHX6FMixSDh9xoPkjVtkIFuDfaHR3h+80Z929vUEhvdTjRlZzRp11JqqhHG/Hkcnpzj/C528Pz
AC86SvgNEA1mgR7jsfM6bGjlPDmjB/3s+9uoaNdMHhY9qmShXMVBPOjoWLJZeSmwL4WFJhLR5u0u
yUptSlZ31SKDK3DPa2nBFskODqG6u8FQ/gtFEinh69ATQcnn38N7T6zvPYHVZezgkalDZXCo0li8
eYGyVFZSF6ZPsmpLjfY6WIFYfwRCdEmf+r0cZT4O5zNOB+owH0CBhnJ3zpi+lTTuWvIbDDVk4yz8
DiA4z8TWVJ5u3MQc3BkITMMPuv1VJ1370eN8zcv06Z6If3bTM+ax/BfjCkBCuE0DST9dokWwXtvX
aZz5SKnjrxU9J/C3OA8w8okb2M/Hr/bw9kSvQcGtrHQZy+ctJNVdZ0ktn02ifZ4G3AKjpwoeltdn
Zb8kcoEjbAKln7f9LjkBjERRuWr02qpbnnUEe0iVO6CL2n+qnU1UNV+BhAw07jPf2Ru1DS0uE9OX
oZZ6TlDtV4B6lBsEbz8Zbx6C6WFatPKgHxfURhPuB2B7cXyfYYn+XOvraxY8gggR59hlGHRNEidz
ERy2YNaDuGoXF+4U1l3Np4QjHiDXofwxNHto7aZELW4WPDF417zgOotxHs8vITpmdGdBXIYukDl7
BH87JTKJrLR6OOF3jAG62cs5VARcBMqYRzaWkyrL4Q7O05gh4wKyAo5gVO5KEKvtWtMT+yQR4vHf
fA2/zkYFHseRrCAbHSbcOjE6AHOnNSf1ahq2QdYTeMI8/hWcGV10Lu3vacUSrrlxeZv/E7bjZqwa
1iKU1RxpA7Ge/Vi6gU1kS0Jcg1uTJUCTJfMCCzHHtU2kqhDAl/xyKVJgI+S/rLSAvmzP35F1fkJc
i4KJwEevYEKeMry0gPN3Wa53f2P3pVcdexuI3HHlnowq63Ka6MoiOQzugASLz5uc38IJpA1/zt3G
MS150+899Ps6vqmObZMbgA53krq6W1eW/j7yKU3+qvnAF7lHXMTWL8lQ3k144Po3Iuif9lFOpa2p
dg0NzXoKoI8eb6fPwJ1hQYvmZn4uZ5a/seEKqdt+BLbOJfYTcHIeetjObiG7D/bnSzmtst+G/YGt
qtkqNt8hICYtgb2sHpZfZ60Jc/q65XSL3OfbqGNdY64mqXaF0XYnHgZqF04rq76Ixm1Pz3kjbcYz
LqEPwhTzXV1riC4oD7tRpRd5m+D+HFBLKVu90oYhgpmHVug0+EKDB5o0X86ssbOLpT5Ca0zvSfjJ
S53m1QOHDLzEo0dj95PQZBPId45CDBbdlhBjVKKkU8lJGfsnUVQRrKibk21JjuX3XUp0JjkzWM8h
9ZPDiwmigBEdLUmdscDkuKOLe+GWkKHBe16NIPI4czQspHpPKuF3h27WA3eb9NbY6Wge/wwhoDtR
ULMvVmuVTLWLWoKhYrINmSh85sSO2HJjmIfpsIc+W86hCzRL129MGm7hlFJsNeMgI9XHadCI2Avl
zuiGIn5PjLLpyZYXDErOgXQqaH2YkyE5yNFMORJFZ89oWCzGsLi2wvHufzT4itADACu8JkVVPf3i
HUmSQfL99WKbmleSEkyLzl+ocNf/FnQHPQvZTQ64HjVv0Kxr2NfC4Wx8O2DQdrY0jggSH+zyYfrr
RT65brKvzMKY0+8dLipCNilkAYsd3lT+CEd2hQPKkYBaSFFrthGWu1t62nIpgO6/nUclNqZ6DOiX
I0cKhpvyW2H3g9gWs+ZoKqTiZ920q4ddcw+F5p1FcL1OUV/WWkKfRruBhlUsiE1O3CbgV6+u/JU+
Wa7C9X3YlyuZQKmDLzfyxbabNeZeELRCl4ARR4qlXZRXXy2w8hAkGmaRT37/W8bm4T82e1OcbrXf
pCBHq/FQBaXzID2PwvzXb8yActGNvTd9KOQCvdAJspmpo0qQtwfZH9o5HUa6BhDeXRVl6jG5Uch8
M+4d8DTDytEkv0i8JEhJuUuvGNOYZReiIviEerl5vSxWYKRRRQlVbEzYHYc3Jf9Sj6n0bpzNO7ZV
Uz1pI6mP27yp99zwwpKzas229LZqSRJFfCdz79CfHCdzjKVDjOh7+6J4g159fKRrVcWFjwc8O0m3
j+JLWrTu9zJW4ZLJNi0d8Eikt5PPQ84diIYaEsYHTT6iOgqVabR4EEzUq+xpmr0DBz+gSVnp9/hZ
Vap+N3Y/WAEE/JGVee9NhsdADCBUlYO/IMl7AASrkdhjuDygOi4KBO3aczVDWHwagPpWtZ/bkl/K
uJJuP2egEYUug9eGBy1KgJBRFZZLD03pptSKzGNjOC+ba56G+ZSNyLShply30p+bqdj9kRMhVyUE
hJUfPxTCC42Aawpcy8kNmsb58YjznK1tlhLwWtxkpufzCZFjdm+GCuy8edgHexCzhxPIm4OxXw/G
9WCWREXP0Y5AyFYvP+mEnsL77YNBSvJjl0ENBkSCsJ6kw432SHgFsy09Q+YrYVuBlI26q8G7u/yh
ltHiwnCBeW14DoVH/dspFjAbYdoFXQzIOcDNSoGUjt+VQJLxJ5No7xtkIsCMCCFjSyZ+Bwu5nhbi
POfPMOffVHrMU1rF1ytUjvnCNDlx9IU5IgLgTldzn5hC3nOG0mZpJFTpt63ckfA9Oc8sF+fERxs7
wNImrpacQXCpdMhbz4ZTD940jREHoVslggZa0QAdFvmHuR787I4CyEV1G9JOW/4GEA0fVk7339NH
tSSQvi+F509HZrHfeV+bi8d0Q10+RChPhpOArKCOJ8P6cCQ4gyHDdWnfheRPlseWtmv0paZbWPJq
46Q01jXyHe8s+mne71RyoqD/PKSAQn0Y8inhJ4fplbUyMe02bhpT3Ihl1fD2a9a27gQE+wVmAtdM
QR2kqIiPvWRmdF2SyitjJlqe8RUOly7Yt22RvEaif/nVJYC674hIG4gY9ZpcEPpGViKJOSjQEuEx
/rpQrzD3nsfCho3sJ9uauMJKSWeLqMBmexR8Hd0hzefQuzLqkf3eKcUPEsy2nyySrnT1nsNsQAr7
WPgtrT1c47/HhFlPWWtg6V/bgC59Un/g8KHyvVv/hSMXcCOSeB/3peMEoTF8kXcKVGnRqAJk5y6l
eDDY4w3sH/293F37ga07LApHgZzEDA+fOSs5Nn3AP7cRDtXnKLdlDTUuGKqwKfBxCyuJaJVH9ZcY
wbHHQGvkFr+245O3TmtuHFn/BIqK3nGtLmNSTIK79/BViuAQTMUv1EvsBBiiXbIH7LOkdejv6L0V
E2eWZE8yUgtPZdaXCGP/kqIcIvBUzPKwEo5Us/rgojql+8SC3alap60bP0roelQwAXM4s9tmMfTM
5UbAr5CKRCIW5QX/4R9Goy/LUYYQIPY/JnRyT2QgPcz0Q1n3xdkjMKJZHv+Dlv+rcxLNEo1WYAHX
/Z2rXFaAAjzFXHzpEVw2xIf6EHNo03SJDLyMNyl3MqMlVftvCqtXJ7R6DTNqTFTpyZmDFitqdhHN
wCy6k71dAv8+NNyBta7xVM030qlk4jghrkfI6X7tlMmiSrvo7gUJib4411QINd1CbMIMCDeG6SJ8
SjZluwKxEbQFeAmVXhsYAj2cH/rZ8YtX8jcdmvhd6aEhHjQl9iNFXD5UVZLuAX/JiQ/rQoXKqnU7
m1XInmDYF53fagMTbqSM1qOjzEu/C1xCs6m9ONTeUvAOB9WgZRd8E6DGJrS4/yuiLt0SS88yevyX
/sgDdRcgmlxHJlHY5hdoZ0YaE+7+9rrEUGaWcgTf5JCrv+V92XAWlEAmet0v/QQjTiXdp6+Wc8f7
foX2MvFLxMYWxwsqgozQdqWDgXuyfL4EwmvklPtuK6eVlabMT7PzkpEyJ+hpdXRkxJcyxc5IUxD0
64y3Sz6rtR46nxpDd7TX5j8zwiTsCt6nzORxh3v5du5PffQ0gFFX/uRnhAuUfeRruO6eUG8uvqyp
HFqAM6M9RkZiA5DBQ098ChnGcaVJwujbMLbzIEEVrWShjEtT0EJ2+YPj7ylrt2S+naUxB3g9txCD
OjKSFnfEo6YgBkeLiLSfJ9kx6zZsiVaiLROvC9zFAHwcuZwL7xOwPfCAWtVOzSzIrd3+G5NF+asv
J7rzs+sNSEMQ5hnqcJp2h4UoQgqr8Jj8MQBbkc3upXIRpW+02CzJ0lmtXyyRKgdIbCK+FfssHVNO
AVOdQ3uo/fFeBDEizKH0/GvmfdbEupYiauM+NHRrRqptzvEcPC4684rgSEakwYI8ZlvFbiT+dnTr
Nk7yE9N0PZc09LYhxu5aEEBOHlcQcbqT1F5kadz6HJsRwgQuPrWBVvqq/D3OLE1IIQgodcW5u+Dx
wCaTBfCy7fu0BESVolbjb5ifVaEmjrG0Nem2F1TYPdT/6VituuRj5761a4Vx4/PgCC7+xGqXKowZ
ysbCk8cv8FUaWa+KfWTGfQ9OJ7WJZe3JMPdGLFqXbg+dStq1v2fJlBOkes7scJGgjHlen6nV0k6H
zgKTEsSbX6/Di3u2FbUH0rXWYQxQ5qR/EjFX75kaJP8TJTkiX1tIsvavN8jjIPBOsacutTk3PXqi
JkSWQ1wshiaVVoco050wyt+N5hv4OZRonSQ1vGZ+5i91fx/WEFG2s5uP+lsZA6vm57rLLL00NNcu
5Jz+KnDyNOmX6dqvFI/1XCS2ogzS2BZUkFhSYpVRzYGg3JRJN7cpekBCRg7S9/XSEW3x5MLVl/Q7
9oR926ITAVXHONQUS7DUiSetG8U2Bj8xf9j5hKwbBsYFofUuwwsG+uCy4OnWSY8g6xGXFWId/Ya2
kBkGGaoOc/rRl+70AJFogBQrvWrl7Cj6in9Kw/6II/Qz0dN+Z/nl34FW3lOIZQklsER/GgJAWZkk
XjhhIt9P8dcVNfdZikT5eF2YcH2/8IS5m6lOTqDxVIKI6CXoKWGxQb0qttMVTbPX0PKC+Oc8nKeU
Ml0xZ+ZuXInFouCpqb1RLqNikn+FO6Nc7emY+Zvw6czV30rfRAdbo+PFFfLxoS0Muu0Kp5jrEo0M
CHWzaUnNAh3MhdKhskpM8SnQCwdPXiyOhCMbZzkf8EjgfQYYQBksviID4XjNb++JwC2XFhHas00t
v7aNIylDToFOM25R11fOOjUCw550vaLb8A72oSkHkaYuiE72Uc1RVl396fPYWMfjWxX6jqxm1X6x
uxB2waZPhQdOvlbePIB7NuUUbDxA9pOxy6BzytzItDgVy3Hz62l9eiyBAm8BVMurOINHQ10KAxdL
OXEAsHq05LqvHHQgaBHax5hGgg0gbB7Yy9K11C8nDy6+eWN1ahMpvdkQZGcvbeEw7cly4z6LYDkJ
aKmmrO49BH+q20Jb9tXXxKOBS/WWhWEk9xeHK+2tO6aE8rzxccYHh2ceEKAoavpYSeiStE5VJrMy
6414zTT5pgzfOzppdHhIxQK7ecX1VYbVv/QRPFuIUwazVGOcciOmLsbCF/JrV58wBE8uMcVAZCtG
xboP6Xbphzmn/fJ/lDSHjofRQsSSIW7KKTNhOSNrdlbi8cCDegZaUmZyYCGiNTNv2Mu9yZ2PXC5S
BZ8I6Me0+42DauiksOEAvA0HwrohvGziMiV420Ux0Cst4wd/kOLK+7yPd3j5wDCbD3l+B+WGAT5P
JQaad5GyL+pgEa0YzAPRWyD02GElCD1xFo0t4GtHPrktjbXgnxyUqMmcVyLJnfSXNqy65UFjU8dn
4tUk0qYvYmiBTSinAZCWW9ATPVERb3QzP8bDUpAvwf0vmLeJwVOQ4Hx4oWOjmHZ3Ch2rkvx0MFad
0gX0cv2QrrgcUeovDMK4aKTTrLEdNM5YpOJqqUka9bKW5jmESLKPw07Hu9DKkMAKAuzYOQnlxjoI
OTs1C+eQ/OG6R7yEKofvnarJzri8E+h8U5FTwQJU66f0e+3kk/UYX+12rAPWUDH6i5AY/kaERuNS
nn3fSQxPYNLmBtANbnYFoemvmgojUy2F2y2Hi3/xX8dpie5XVjmi2eLs+vuSaxQtT+JUE9bp6tY3
p/qBzJkAUnEyGp6+5gTTnX3lK/rK85//sYD4u8NWJWpEXqqXGlXjf4VMaI80OU7LXyCqFxer04OA
4hmW0cvXai+MZm+PvFBKobbr8k6KaK4wFZnuhiIYdkuhguwojpTjPrb+p2B27L0RR1fnd7zy8VOc
w22tG0losP7HnyuKUlPHfiBCJ3oRKveiM57xU0oO1DtV4TiMMGkLs8JYlJqZ5WDgjEA4atBcDiKN
1nZazgdMpy8FDZuipAmmZEZijXbn/XPcz8U6NkWZ87mvAe2/CbTj8EfGU3NIgP92dWwV3zQbXZRs
7V+KmeEQ8TXLeEOzLg3KGuB0Zt9B8hhPFWtXJmJlB1CA9EbMNA5Ti8YFvD2NRoH1fa0bq6QG3C5K
y9qB6CCrn63chZAmaSyKVEhNYB9/oxg3/4V0Y3q4mpevwAeQxpCcLTtqoqXKEg3M1GVvyrcbPH6K
NKR8XIh3wq599tkimLcod5zggP3TNzGsBlgRjMx6zwa0fCUtEtqyEBVEYAdUQ0xcPghDFXgZxl/h
KvDtZu669Ulx4K0oMAsR6o8elgFz9RKMyHDO7x7o+p2oY+ER3/f76BVmqPI8cHdW8TLAKKH6aQqU
zPCS3VF7/aq+Thj695cw82YMOyedg1yU7ZDyoA7A7tsIawwlYhP25CTIUyzoeHKN5h4EyCkkhYWB
l5NYIoinLpWv6buIvSTo25vJBxtvbCf7TxQf1mLOykteey1K+HaIzLU0CcXM96bYUa+bJqfVnB3q
hnqSm3BMTUFZrI3g0ssKjdbUtqogbVXG0K/s00QpdpJf1g+OpIfWqYGUlgCcWXDshwcuF7inTXnk
Z7d8k+1dXPlj/XzsJxc4t/USW09PpwwQddWPWb3vKs0NkIX9OJB/5EUShZHW+gfV1sehKHACPDV1
PMK4TO1ozdqSlNUEPCcdiGcTtPZaXCxo3zFHs1uP4XcMLHau7pJ8h8mwK92Y/hwGXKbPgfUWMgoE
Kq5ofBCOXsrpGDFhvhxqACDMTVonNejUI23fHC/PaFJ6ZSuyfHQeLquVuP67EdhaVszjyRMgiOjp
MmlU3NbW6WlGcediAnhNTVb1wfhYGnBo3ROfMCFiDVGeoZii60JRjVDWfHLkdTMR5g9utOVyVf1y
ubuG7lr5yBRuZPDyRwFCulj18RnZO+htcZaDqg4uluJnZRKEkk6/1WF+Ftjh6jWe1CIbk96obglE
x0lraQrbFv3uFHQoPR15FPxD4qKgee4d5DlufpDb5hhpYLYBhGxvMyDA90pjKHc6v8wj8ikEAHHL
fB9fT4kmRv9hLm5nW873x4AdGXx38G9ihoUnPkCMioYf3WzGNpXAE0Wp/DIb/DJxHixykzLAQmrp
5W9f0ObvHuDny8O23ke01bpzo6SFKzr7ZilQ/kkKfJ68lcpVswPZ3C4c7YEc94hafP7u2eItT8Sg
UmhrymGuIpGXBjaxVQHBAQgjHrip3Q66Ig8mfx5pu0/WoN40jzIHTjKOZCHm4UuIomEzCZfr1raZ
VKvFGldjtkV/S57ZS+QWOXWyPTRVa9nO6IC9q96aTJGtiXEl//4wc/cffN5edlJpPMJdv9BHaAck
S6pOozXhKgkDi3hFIwqmS+HbI8n7plicglWwm90Hmo4r5i2BYp50feVK7DTsh6fmK7iT2XYyRc1t
ERwEiIJSCz7I5+c/0oKhRea8Q6Zg2n0skL+DH2ar8t0+t/J4HtFzPetH3jFn2okAqYpssPfkIvtM
E8p4e/i1Tqzy/C/0D+D+2oQhJlKPdO1AEaPx7ILzcVzxxB9wTr/qN5NfJ170WWAphvOUP0SW0uX+
hvE/gEeL2/SYgCBQvwgrcGfGfcjAAiTkqjoSseJiRsUHQaWmWz8as/TcJqM0vJoiH3q7nb680D7N
vgb0AVa/jbbTLlsfV0p0ZlVkTrk4IfMzP6JBPOuQtNYqa/PqsQVPobg6x3qz4N4u6nczoTF7zUWY
ZYUdrQZU8NYZp7J5p9vrB7/tYJytftylmi9hhkseMeX+cecsyBesdAdbLsyqJ+MVdgozj1OcfSaQ
kvTo7vLVL4yXRfJhQD3LD9ctseVruvT5vcPHZvmLdnirdamvy8/s1iH4PuwY7+pvpMv3Tuup88ef
uQZ3GTiY6I6kZJPK/8kAPPLNxY20w3GEU72AJl6fEiKMEIFGQt9dm9oux86OSOjN3UBfg8/Wxshw
APuXrLF/7SppmfiMDk0SSYAe+JnfyepcH3H8NPSRlgm0qQlULRoBKwcv9+lrCNBAet9sCqzcDnsz
pZzdVtoGq7pqnmwrpiu/2/7paQYALu0AjjIa+7UrNolr51GJoZkRPtxUmwGReOZEvwd5RCHTvxhn
++b4vTyzPocOYEuBTxlpqbW/PRFj/i5Fcix06wxrImQQlnk4NIn5j7KH028LVCYa4lc2sr+jMI8t
PPuIg38NJeyaI/qHq9G4wXNOxn8nIk0h0DQugok5SGA3V1A+z8RH/Y8xCc29B9RF9SE1wud7GdtG
GnugF1cSW57DuQr3BlZeqpZWPO2dwwd5+NV6GXbMnESqe+H/eKnog0BD3Gzyk8OlN8GyxotHhS9h
rQhDxei+sG69XMyYpY40BcU3hmt9yLREN5yFf0rSVwa8a9OUsDXd8E2eQTNDXDKnTyFka8yHIxx+
vx8GBxAAqII4EqdNyfb5yt//UXZ0ToYGylwCgrenwrw4GQKrU1BGtPp5lLnei4r/hPlQTAQPn2/+
pd+x5Trqbo3tAFvvZp/yr6+INhHPTppEgxk9hSAxj1Dh6FoRcd9Tz7cBY0Cxb+H7PUrWa7xn36PZ
p33IS85lLuiIpB7nGfYN/xoHxpuFenxacwtqA/gG0MSDhJnH+VIFEW3EaL8xrpva/UzeMlNQ5R/r
vMej8Zjj4RQ9nZhv39tlVvpZ/lHUi3U4wdiqYzsN0Twr7l6vX3fco7h8KCOvfJp006tTGhdSh9g7
Pt1blTkNxqg3gmNfRzhBvFjtj3NbUgsC3xpIt/XJDgmm2/GXdeRlYYmw6/8nxMK7wYslLJeFaIqD
5MOS/+ZrCmx8gJSPGdj+tHkb+V1kyT8gueC2nk0aX01Dy2cybBMP/Vo+RdyrOwcXwDUoBzJwiRor
J45X5QgrmPZcF/4IMxJTeRz1bHlLxrme+ZE2iVjfe29OisXczmErzzXRjDl0a2SOmNM3oFdC9JKF
QfS5VrlRRexymJd8jFhE+u9Aj94sJ+a3aA+z2PGBO5uSX+hJGy+wN1feJT3iME11iHGtqOFxW6Kf
ynMDF+r57k8OCvYnK6zSTo5NThhW/0vvCjU+RqH7ELBUdII1Rsg3f4g/UrWFDKeZ8KfHRqA0qpct
U19BP14p4yKrsbpTRFMI4jnTahL783XoMiM24nkketWsQqWda0SHGipis2FFV9NP4dLkKXhPyRzN
kM+UeI2XM/2uBP5dK/IV754q1Qat1imG6cGR5qEAXLrCIVC2byrqpUkeiH2Gx4v4lFYdEI/GE8oO
qShtKNKdxaw/4EKWZ6E/3CYXvbAmyI29M39qQ07ICpDI7ixAkjFLoehKhb3zw1sEgLN7HPz3DGwT
tFmFLQZ9MnvSwcmpFzmC2Tf7JQMWmThqPMpJs57KMRth/A8QPGJ1PrB3wy6G4g8wql2UunLaDy8p
8NEePIzCOgmJghMPYyRxO1o4I6pqOhd2cRdrDXvrmvX8sTqFvFADOfD1oGeNRD+fUIQcK8Of0CY5
yssM6+leGE1RGILhz06IlypFs0goLrzLkx3XV8ovlvUnTxdBHtnKNQlwhW6aD5K4hkugo+z92/NN
KDOxbuIgKCRSiW5n4Uk0aI8yuCMOWkg3pc9qWu8JPUm2Atfz4c/6KTtXUplxolmCrQdpe/YWds6a
kWFby82vngCY4bqx3iV9EAE9y5HTpRqg3NrBDNYdAoLjihGyW07YcmxwhK2nfNFIlLgcLGOABdco
CIQXxTiYn8AMJYeIF/md8c36B+3bU81EGxvtujFzWYNGAyhcdTNCjCQOKh/IgxYNgwT/CTOKbihe
LpJBnseTET7lrhuoa5oegqNQyHJQwoNSJpp0YBh1scF2ZP/o0tx52to/zrsGiVEjnJTNvkN8UWKT
TUkVH8uxOQQA1mbQwAbJnqNaJUXJHFxhyPrgYdq8s1yy/LXonL0aTArdX2/+kYZ6fTuXbBNWmM/7
u+60iQvU5JmCg5TiPsq9wJ4JeNIuMcJimHdWNuAE4xRLC5G5dp0Jn/xCRKSkTNUYKaNez8Jr31gG
aE/14a8O49/+69Ee5Xm/BbYVOiNa4xnEJRsZA/cyrCR7hBtD27a6OOr3328kNPVoSNx9B0XbfSR4
BmgUkA2MkZGpuf4YnJUG44OKF5UOT1Y9Uf0dpTPk6qgJvVLi7Q+VI3qPCFmw5oEy49RWLNr7tvvU
m6o9s+wNX/JxEtUdMHcY2450/TE8dr3PqtMH/5POya9tlWVJ19NVldY/6qvc7p57Eb+wUAHGf0jW
YdYAg2gXQfmD0yTwdcqKTpGGhVxRsxHggyMYi/MkH4klqorwSZSe/CaF9qJyqKb235ckrVW++h+s
Zfju6rkMUorMvU8asPlOBB8FyAvVGokdgeGUer+qBTm+ttBKmh6DF+Gebq+fvfhyqIZKyahnByOb
C8rqJrfGPHZf7y3IiaRjp4epTAKsJzmYltYN6ysu4+9EBacG0OenmCrkuZSy+Yfo8WqWex1xSlUP
PhWabDr3WCHq8EpoWgo43Ey5bJ1TO/wtIrDpA292TAS3HwYEMsJQboSVOE2yiUAO3qhnmyNElYqZ
HzCgggfwCbJ6knV8mc5IinHoR/fUCd4mOzy1+ImBi/HiPc+sC1EkABMbhxUeQkPWQtRTIOVkWaFP
4Ere1QoAXe5mTYqj+OZ7IL+ClQ3/GKcguD8WOr/wDQMMTfT8MJuzYhRmrU/ZoWaIAHFh3h1Q2084
tTsXefxIlics1w+u9/rBXCv7KB2FRuxl0SoC4VJMILfdf4DPSa92wTuIgiM1ezX88nzi01Wb7kb2
1gE0O2LvzIL3cylRpUTdn2Dfr3uZADUu/8UmyOoQ2xb4opbS+Ryh5PqSz9z4D5KDnFRJtI/MMYML
p7CPYQ8Q306y92O6y/p7mNM3VoUJZwKzGzvTBOqN5+pTntwmo6ild0Z9gBMsmZmIZNriew6BZ+fs
/qTDw7V0Il6fgGTgTeJieSA5Tb223ZdFqmrcuboIBA+E6mKlj84D4kx7Tt1JYbOSDTMBr/SG7mzC
gBCV8r8kkNCH6eO70mo/sPD9LminV71Y5LCoFRAq6GlLvgkcU8x7kqnv63K2B1ErwFjoGmOz+oYE
pqRFQD7GQ+1OuKdQcnJ55qE+KISLlWvPNTn6bzHlZMv2+2SBgvACXv5M7vmiwqdOWujAUpA8rpzs
8x4BBZGuoxwfpXYCWl+4J9WUcaPv8ff6KJ/fGovewKtnY3HNeIxawtTNIBIk7qs9vLNIXYXFQWmf
AxAH2RM/o/sjkF7pR+0j1+U1xVMtOXoHA/nd6NzMuipKnZu0yDaM/beRmLN2L2LxCZk2cn25B3LE
9azTxDKiNeXzogv4shm1xu7JD9QLMh4biK6ItWJjpuDBs09dG4DoMnkNU4Mc0/REnBVb3DeeCe93
4JXSzRgivdMMQVbF9kys46GdTi+wqBR28H/UYp5Pa2MHf2XFKGFge/gpvodugSu3W6ponCzKxzrx
qYyI/Do1qYVPzBbFvB287XzYZNtgAVA+C2SnEP6tocctTz1zdMHMBGCMYkXidT+WCoYxNlr/ICgg
GyXU5AdywqiNWzJ4STJiP8ZQIR6GnIGLK8/gE+6tsh8xVMyGbHW/oHSGajSTl0BDz/WlyYr3mDGf
qveG/OYRJ9mTG+qXpWKmR2q8w2bh5522GlgV/gYlyUbksXzojP9lDjOn9ymHv0eXrfHbG2C0bVc5
9mFoQLZYVclCWaXjDWTcHq5MSJ+0rVPq78a/LeBYW46EgLw/j4xGktNk7yQTGbBxfWxLV5Y1d0QJ
mhkkrbxcJHEJ9PSqM1nDSAA5HFgzXwFY0qBkSN9qVJyAOuiHKqKfYXMcTOMqdolSD7sKFwiacDDS
QTFIlmeqE7bjoGmaqp/jkhyYQQKgnlW+N/rQGR73+zHEo27hIEsXVQZqNdZFFE/6Rx9GECOJEy1B
DHvTwdBnmNiIuK0I8RD5b1PnZSHWvw6bbX5QkXnB1wFlYzJ0hhA/fK/RIcDnzqB39iuN37HOVI6F
fB7H1OztlnCZspcMzW129Fb/RA/gCWMC2m6/EZt3VrWbjHEqTsfF0JYzADLJdiP1gTmByI9igyuG
ipT1Ptf7Fk5H7ryHT5OmXkllDekRy+TO7q0X8pGuJE98/RX0USo/1u2tvk5Ga0Gs6zviMG8I/gve
KNIFgVZ9tmavlH8OgXhANTZvRW+74vDCK413OupIxa1IxXGYP2x+RuLSz7TpnacmfxE/vNX3oy1a
f9mOipGRPJXHdvIgxTJqs0IIh4kYrEqj41yrPWOzxUEGFvIm85qW9Dxt7krp6+e68Pa7DgKSQ8JE
te7I9XbYoXxUHOHpHTFH8vPunOKQwyuwAXgQr66OZXqtlLqVLgPN/5Ho3iavWq/kHNf+ZHckBXf5
41NxcnDbq72jOpcbk33NIk+lRlh8hYIshVAB1lrINHgaj1bOtdIVONq7BKLDrKAbBMa//N/goFK7
gDLiYv+t3+E4S4p89Hyj1y5ZJM13H6sHyggKIDfm4UrWsPaFooikkc4kmoJwf+vdoZ0Pgd7EZk+a
c770HnKtQeMYrjfb0S+lXQY4sOzpAD0DnFhBa5zKjC/n07cmXte/wQMG1NM5JfSfWPlr9njXW74m
OohofuMy7TgGKvPrbIM+9S+9t6Yfk3VI20S1UgdSYbFGuajdXDG/0oSKm6kYtSn83knTRmp0j7il
gYy7IzH3lvc/7auTDaBL5S/a7NbCT3inNLO4Efu03jSJP4tj2/a47ATPUcwDAqXnKv5BlxIIjUhO
hM30cRwxc8KTTUQAZspq2+qNH5NTR7K/EyEpPrd+md3LNWPQFTXoiko1uxAKQwDcOAVnWnPP8GiW
01cMYvI1acGJAtRspfuND9TWzpOmzy7RZ6BWJYOLw8TogKWK/MBufLFHe8WsdM4g0SibaUfY+mS+
9pLY6LhriLZL1VPUy+rZuk93upf68uIY64gljDWDTX1ZSW8jhX7iQOtQ/t9d87OyM5UGznv6FOTl
TohOtmuWEgkcgbhHbHVNRu/HEdl2hY1IgeP+zHB9jthHfaV0UYLVPpx5G2317TwSFIAVATNueoh4
Bwl++yMIE+8CbL151xvqrmYylEzryVpUuswHsmjuAtC7LqYaSU7hiWnNqaflcEObce8urZWFFtF3
Bs5OlgM72Ib7YObOj92qWaN1cNug10qGGMv7iE2SMjjdZygdXHhha2SY+SkKY2829w2qHB1WoyeT
EvjLtdI9MkM31lI7M3Bwh4VDC5KfVjY3jiUx2mVF0AXfDEuHoawXduhtxn8Kw7sYRqHtv4POXB+s
PcH1RFua6lHpiLZsuJwdusvb3yVI2kISb7Lv7jNn+KxXzawRRxmh9LsQYqr6qD/Y2qspqz0GOkt4
/hR8DoHISPKdVKHdmrVnyI2+zeWwDsd0uo9EA+C4G4E1u7h01Hid4cjwAYEHQSM+k0tZKOU2bpDJ
h/2nRkTNBn97S9rPEa8+/08ng4lYjhFE5N04luRUMx+Rw/xesxfop64ojnK8TUse1zhu4Ip6r6PA
V426AwLtyPlh/EL3IH+ZQVxlAh/suhnEtFi0AkeXTZOtWveKL3q3cvXETmBcMXzbnFUwLbYvUv4g
Ufz4xHY027O85z0gcT0u386mfBD1j9vnoNvlre/JgNIxAkonqrA5IreCzHRsAIJYqy9mbCmBYQle
LRGneTjMx3jco/+6ENY//GQ3ZIlfeK3sMBN1yU80IRmZo7dw12/1ipHfeCyBA00aw8rDBx/wwP9o
kjTR9sQv/r9LYNygH02fPdZlZFCP8E9G37IYAk3QtIDEDocEQ3sLEt2P5oFVLlpyJT6fPKqghyav
dTT4r4CICW5Z10ERRb247WOCPs9OyqXzuoZe2CQ7lIEeI6tQO0oaQuoDnTIHE1cyjVLC0NRrXGJ5
bq09gOlbAIHuCihQTUQ6Y0xjpkxBY0FOeuBnIsvOsE5YzkkcK0aIstD/E3f19rfKuGwFFOAXTX+A
fxGm7bUo/pkm3WPXoJ3Go/WY0L7lGSr/r3/f35m2Eo9wKuH5B/kuuz7v2RqNMi/gKIyB3+GOIgeQ
3AiXvLBHnlzCTpO4KJF0jQowsj2aB9hkms3CRX0BtiIuOu7QjOFNF/3YdRGQAo1W1sYEEFoNu4sC
df+NMUYdSWH/4MTmD96TQNOlb8FyIcapV+qPEmHZLE74e7lyVpNODBGcNeZanLaWAkRexEM6DMDf
UWdIEpx6CslUnhJOKjE0lXk48graZgvoM7P9al5ckc2SZU1EkBJ8LGWXMcML3Cl4UogojPa/XAQ9
n28uxEW+YesQRkxQ+fCE+3NpuRzMsYDkMUplbTwxpaV4ILTlvegMA5GgNs2MKvbMgKXxakYtxWt8
+6aFxWNRh37CL7FtOw3oAMiWqCbFAHS9KXfzEAb2BuWKTrA2Gb3/tgyQlvvpNPlSs/cdQaMhCyyl
Sc2h7pDUjeuTnvJY+xUvCOyBrVDB7SWOiqcWzIQTpawqUoeeG2g6a5SCfseLegceB0TQhZFnCXSc
yiaVJNWiN5Ra+ASm6w3EmpVv4K07nVvTMy8TdAJm37t7OXIBrpnBWm61argFyjhGUZRIjxymTHOM
TgoIQP8j0gjpMhY98lYyGj86cxft6c9+HPoqeKbBmgDAAGM9wSTIs8OVEyayC0hmcsnAWCeflro4
8LYNyOJxf84xBb45u5JfkjQ4bUT2tCXrCUlPD0Z+Uq3rwLV4WKcwIwGQm7STBMwSLwaWexaSh1Wp
KAUdkQGYHLtNIQv0rp/vTW0BDBhi73W0bzLeX+bKUFRx8POZeHasNUAnK7qLIvE8xtDazcmhNpx/
U7fa7l0/RDiwzaXmTB/sM2JUPDaA98ICzbCinjhH8EYHL5EdcRggeVttWi6Zoy3fn+VaHcZQ7xXv
ru6xxfbLUK9cFPb6mge1xIITlsphIvrcGLGAq9QnjSqQKRpFtQfJRw9oOQyzX6nINEsNhzB9tvp2
i+y0zVY4ETc8XN2+5vhbbReQZvkBaWR8pBfszRZJkBTUKgcvYSLsNB5FPFdzZYsjeQahdYyeffs0
GasMyOWeM8EN8MHMKXOWRgm/V1BBFm0fw3BuEeDLS8vAP4p6/ECviZdtQr50Ilv/VaNLLuLWrTEJ
VqUyAfinz/lI0R5v4mRFEcfC2qAsNad4xdWENUlPF4/Y7AUpUZeFoYJcggkPziW/jiRvecrTls1u
16Z11c+cjtWoFOQisMhxP1FzkVuhwqwgiIpZBVbjyg8kJK/mlpKzItOnnKpqQ2OsGgIZAT1tdNND
og48etc1LO+ZcJ2lgvA6Mg2fAG+9e6B9ho5T18c2DyRHFMXcrblz1/W4zs1bi2md9aua5GAOt2fE
J61wLUgrgCfXGRDq57795i1eByakaV6Nrz7sXvp0nuR327m35hkan3wpFZupuJ0YcgVikj7RjdaI
rxnhXI/AaOQOoGI54BS65KHv04ukwHPgpC2dPefkoDVu2UnX2kOssv6JH8pgwLbXcg5h3JZa5n3q
6NRMlHW+j+OGA1PciMJuRABWRoQKPqHhXP7UPLmAeeAkJ08THCLRZTBmNmyqiR9TnYujSrt5K4nP
NHY0ir4KIPq+3qkOyBvMFALds5byIX8jn0lZ2Ir6sPxrVcUSHuIeSx2+jLUeZqdAbFy77v8Y8C0f
IGJWYKdItfYs1ovqGMBs32wsWYXfRgT3v8jG6x3RbxduzBRCZO80EQmD2kcU7JFo3vaM2w2kFYDS
KGqbIcdbDfnjCVMj6z3q1j8h6XZkum8OQJMjEbJHggNgTkZnwoy1oULvSIcIL7j25wCA1scKDdgT
c/V9u5IKfd9cl/XlOXmPcqJ+23uYyfpfV66uwavmova62TJWZp2BQzHOrTyIKS/Ts+ZeQPpM2Wa1
zHxK2N3N/QAto9VIFhFT3CD1OygVqst/yjIKZGP0fVfZo5b3gaxxNBvAvYvF1sryII9d/NEtkUCm
PSt4OTRKAc7zZsRzjP1AntqM7v7q4LXJ6dI8mpAVmhwOlIKDiOHC9yr3N/o5Qp5Z1+KS3tGSJNS+
n9+hAXLZ8q2R1cK6CIR/esP0UDK2mW9BY00r6BVTWkHRUFdvfYLaHj/rykQljLKG4cRNYibUaBwB
ddTuuo3OhUNlJXGm4ueg1ucmx2JJVxrvl1iSRsA8pnkWhL4Qgr1UF4T5HUnJr/hSaNcMxVcgg8AR
u0RJgt510dQNUggDqNfzmrYmRZMIj9DksjUHEILgeRURcUZLpkqtktgAsPoJakx3YeZ/Qt4RMkZb
mpiOaq9rcWue6EOmjpwa3XC1BZj+4GyH+cw/w/7k3vdl/KAe/n20GXCbf+KiSGd9ElWdRJG/+Cyy
7AkeKeK/ZcV/HaQNK57DiroxzkNHzBCmiluz9a8LqsN5DZTzRaNd3PLc6UEA7CfKCyUIJAG5/0Fh
Q7GXn87M94GM1wle4CIEJz+YtQWQ8JHPYlD3DDrNyZIpAcskHmnfXkKysShMhS6ogH+c6pxhcpX7
LUn/9iFe4JcTw5J+P8G6YjXfjA0fN+gUdN+ZUIZr2HB4g1lX2Trf2S9aow7bZg1Xyjmlo4e2iBUG
5THAC6qtZwTYl50bUpuN17BUmp/sPXBfo4CU3Bk9M+mbWO7gJ+HwSP4fgNmbLQhHL1fXdKa/MCD5
RijEeGWt/S7XhlMlJLKy/DnelxuVx5vPZpc0l90tfAMUZWwLd2NYTAzQTRqk8SRgCDzl0aNT0bWY
TGzoj7SMxQLQr9Ah0nJxUeBNQr47LPX+Trqd/aWUEg+B24JVM9SjGH7foAPI1B3Cp0GM5+tMRiNI
8zUXSX7eVp8qa2HIukEGnQRnGwmYdJ9k00PrrRAKTg5JhNEpbyEa/BON0ybcHHEYSABk0ooqxb5Q
u+yjWf1aA2tHmbwLAKZC3awMhEu8q3RbsHjWv3eqzyOiYBsrSK5aefN7mRaovLnbVcS3l8aQTOZL
LUv68haX0cRAVzZeD/lvNODxmP2UPNiF/xglfOy1ca+HTgPQN6BLD2JvwO2YbfD6fxJg6A/SgRO7
gQAoUSE0SavzYf3IKRe8iyBgmKSmnHVvXkA7/8Cwh83IhyY5FLwD4YGv/6I9hgAymDcAGnLGKly+
/V5NrRodva41XaA7+2qEo1z6fBp2iLrpss9YYJuV4vzZKP+wquGaa8ghXg8R3Sf8MSSk3S+ibRoI
tCmj7GbFzM9gxXOndQ5sqjTuGX84wRpt5QrTFBtL04bmWbJdcC7xsg+PiDmcMsBiM2hpho8LMZ7x
1d6+0xKs1Tm8Eex+bhUR9+Nsp67gDlkXbd7wXiPzmNDXFC/K8dV/gmRPxX3SvIw5cwiBf89FR8W0
0kPAwwCjhBsPAVAD+0ZYVWslS7Xh1fcKA8KE3Vx5M9WLCS5JfifIw16NjqqkNMLa/fyNA4wrEF4h
n0E6XlsIBJt59MNxgMOvVbWIxIFMtzskjKPgX0Izi6jDEtdTEUnJzcZr90fyr1SSkaLNXY/la4KH
ND9KlfsNodH239UBcBSdvNWBOHlsGEc2FM+EEs0eqIriEb1rOAHglpx6xDlfFi2itUi/4ueFzyXF
E3YlhOn/f3Ma56bYrHxSjEDmOfcuykKJh3utHdMQ2zfXc+hRBYyQmacGH/Jj+tKZf91OflE5dcpd
u/EyAr8vi7anC4QHIgIyTVbkKckQPgArFzJ0OwuVDnJG0ROFgN+NToIIW0BYzjA1+uZvGpxUsN1Q
4K8Gp5kk0JD6MIZBVT7OL172ThKNt/P5KuIky9MwbZkJJ1/nHKmAZjbn8gr6SODnx6PU39DTThtN
i5R4Al7AS1UW8RsUadPU5OhBNj0ghIvQWfoRxTg7clGp6KaKvf5XuhJ2T8KxYTMLvRK2TjM/vXiI
hmBZXxR9VYn7XNmkNlNM+RG6LCL6KBnRcadG32oQsUFrL4gZoCZb4ING0YzLNynNyLSbRJ+qqBFD
Bf11wyi8krBEEm3bZh8gPXsYzFgBd9cKmuNmnDvVP+kxL3tJVmNISf5ZGV6WcgFVMb2k0NsM13Z2
fODLbfhpvSq0bKM90NU4B+qAyOGYetH4yaLW9ZvXlATm53YrhV7q1q7ooYcq0AzP4tA3Z57mHGet
C+OVoI8xpYDowFNiDOvv2aFcwu6JuiGlDnAJeX6SGAsWdgfX1wX/SErAgfMX6/QaqX3atkiD6JFa
nEoQLeIQbZX5Hpw8BVpZl6m9a9dCdMDf6GO2anYPsX1zaHFMFDhstxotLqJp97KgkDQ0VQTzq9g2
vSNU7JJLDKBKQu7LIZysaViLDqwgbFlfvirSqoIdy4QIJ3H1jvjC5GGpuZLkhI+5+cPlQlHptXmY
WGYgnUodpGi3M2HutXhVXqTKumSpe2THaourm1c5hgpkcBVPoFEQlb5Gp1YjjB/DDRTU1dsBzHjr
plQZm/iINLbeJ3ZEEAhHIHadqcqeySHbYGS7Yuv6dlJ1uDSNCOCRPUW/Vm1h9+H/R+1bHiGh3zYK
ItVBmfV+Lsg22bZPWOQP62ChO1W9REq4YPOJ9gUyCYRF94hBaG29I+LbWNhbiqEl3C0fsk2UJqH/
xDM4WdJuCLjqayjVLLHHzywjEAf1zH9n+lbZhbcVGbWyNOM2I71UKiwPVCSPS0l7BGiKroIfNSHm
3qbNyVBoTxynkWeN+tGdtfmloIoqdWgPG5cZOrX+XCg4T34duxPo6/b/wO3H84MnUA9R2Pm8i8R8
FKYkj77uiyjzT7zFebljepXipNtD+YRlLwVMdzJoi2Z5zvrwcGLmEdJm6k6iZKDvQEYckfrOBOxa
SxE8kL67l8u74fanz+WlCZ5oGmmYcgeb5PYV4X+s+fbaK9obh1pzLlTlosYN4+bzFTamgFeRaehL
rgQ/EBgbjEZFZE3hXixpYFsHOXFgRxnMQMeDaermTeeAx4xo4wHWDsW12/l59ovSpB/kuEixDpf9
JLbaUmUU1CizYjo737V9vzjJaJlGbN2eJXQzD/ofXyhvBn43Bb6XAyuKH3cCfwYPZ5rjCfplm7sf
oibaQ5yT4yNU7KmO7vQuL2fEPjnoXsn1syx50/LKTw/yj4qH6t20FuJURFIFNnZR/VbV2CdSpIen
mnUrPPuNXKKM//tuLNxIC0I051EJ0xGrkW4ZrFytR/4/hWtyYc3IVjJnXRtcdlhklEsSbBjEzh7W
HoXQDtoLjV3SvtU+xLkEgU/NjD4hqbPq6u3JZqKvDZAooOCaTUyapETQduxtDhnfFjz8KPKkrKUC
ur5ZnZyCiQk/OiU8T5bLvcML3/aezp/0OZkWdi/dLXnDZenZhga7VpOsCdtNbrC9XhYW24dVW1Sj
zArMWM4kEU+ydH6r8g0gqojiSW0HH+Jw2wMGWnSFxZ4Z/STaBu2FnSM9xNRbkK5yE0cJCOvnmwKN
+26rdAJXIVy2Gx74A0KSIaxZ7kQbJWiCf7eaF+dGPx9u2op9YtiB1TOc0hhGf2tpNWG2yDPgLeiv
rXFc+5vyL6y4OuClMfbBLTqK4VRUgtmUKMfwIlJ+wA+2V2fOjBgjbIBx6qByc4rjgerK0UJUy0jr
ejU3N98h3ERJuaaOMuXyCiEuSKAd0RRerYE/g5A+2GGf0t+lVFlSWKAQHdxSoMXUHq5Lp/3TWvXD
Ih0nPcg3SdzPvxxvi/j4JHL7zi9Ekz7Bi1CCG7HFZitC6UE1/Zj2/L77uH3l/W8P6Gx6AtLJt9Zg
r9Lul/0JdSNc8cCIUm62Gpv1nKQSycWbJIId/2qMqvPg4riMpEAOa2cHmvAfUSNUmSPzQVC4Nda9
zOPkG8LAtRizepk0JNgzUX0iTX0CM3ia+M8LwtqxFVRf0RuxiIyMJBNFQlKY1RcqFYO1j/zziPXb
SNjf35FtByuKiNoRHZREex9uG8Cy7FAtb7pi/gFUssWJmiK0Mg4z+UImTwJm6eZpjYUKEYTq/b9O
Zq1KH1vUPOYgus/HAFmeLZ8N6OOdu44SiNJ6k6QCth+qG03wB+wMay4Q7CtgeNmiN7HGG/o6kldf
KaHusO3fl/uosSXsDU/Cpm6oDxR46HrTuSmKt5ufMupYv9gdPTztJ2NFxQk1ubTElTNA95sJc+qm
JFylwFR0hxUrM28FZsOFjbQfF8Z63J2ycxD34c7FTTPxkmkL01RpC49L0YUcT8QM9SKJpkGJ1+FJ
r2wZ07hSwr7CdcsW3Bi56QHvGEZ7KGKKjDNBWLUiNghp3PoARi4YcmE7zQWv8MVxdQqD6LYPi00x
NRRkaiCFtiM/bbLRfVgcG13m+6VzoJTLwKE59jwKy3gZ8LidP+J+7cgX0DXUE2DzsKfL9AFr83Wf
ZRRzrkdcGX95kSdGv2VdljXQdCblf3TfFjcdQEKT85QDijjsvqW/N1unlTbaylVg0J1g9ev7uFdV
y6MknPTlBGR3AnyhZxRsUQImirhv7Cx+i8Ztq9BPRbn0ucQl+6bXASowbERcXGzVqrPGSA3pVWcz
2bZ9/F5hHmmlSx1l80fxDJwr/cOEO+AI4qpIZEygfqQyhT5PO62sHzceafRsgE0frhShRAELC3or
hK+KFbwLerLXm9hNfutykWxNGk2ioAXr/TADvPhzH9Hy0vZqRs1fVLIbouTI7ZTC4OvudNzO8xYk
GuvaWY3quDWEODAQq6GpgoUr+LiDMS4PFRKQpIYFQ05/FScjGUKAGUSxaO1mdJ2edn52J7szkNSl
Zs54oqbCk6YI6jN04/22GwBTtQn/EqwBtLUBAnx+HuN2O1vRbqamLFAa/ZHfOr0KpVLTaJ8v3ObA
FrunNRzd4x2dI+6MTbELdYouUyIKhfNhU0FVLpfnAYhMqMvmhIStWvQZuhyn0iUItbUWuv8GUv2l
l4dHbF+Yoy3AnRADWHXAJeT6GuEc4WXiF+eutJGiFYxp0pL0dm2E0pT3lmV6QokYZ4o47zVwzncS
aRivPL5XBZS1DHtPki5s8sr07DPGVGRYkjFhYQStqP+n/wDXxnBsl9Jya9BvCldtexeaM5JuP2I1
INJifI7DR8DVOIdjTj9PSPVPAUzfWcJcrr/G5JDdL3T9/d1fq1lufObAwtyjc8HbAq5vGuyfnCpN
r+8tCAehZ7DsZdZ5Dl51dj2WjggENfubBkwX3fQnFSCI3g2GroXYjfh+ocnkqxuCdZt/XAp93RC+
g1x6aXSqLQ9zOh7z9yw5j5jV1gE8vBkoNS9lm1+adBtg/ppkOXruYJSytP0wsoo/jrFCXe3XmvQt
zWFlIcTWP0ryNIbVuSIMq1kLRyA2OUm1QC8gKbNiT3NcHJoZi7kbx+F9Hd4OoOAqjFsoerovs+6i
eNaZVvjcdmuZv+NXWWHgh0qEeKn4C7u7yegbZBBZUKYtNsNj8tjgBVRKUfuB+MaY1gewMZ5rceW1
lvfshgMxJbtMLl1rDs4K41w5aJc9qjxu1ijjNvwEMttYECOkB8m3vSSGjrgUauwIQdVXU3HjduLa
NSIUAqnAezR5mvsyCGSDKqoov9ew91QB9FnNFbtsfHslhLwXGGMdxeIhHursg3MCm7VB40FYH9Sn
LhEVFyV3vVIBN+B2PRD60P9z1MpP4w1I5MB1IUIbTyX5hLxbK42Q306AEQ8NDh6E9rYhCuEPPmbN
BRo7JneXOFozb3igFD5qRSV2+ZXqeJgtJAsgLKcwdGEUZlNXe5rtDFQl2A2wYvkpEJRSWAaw9olD
PkJV2pfEy4EWdy+oJmIr7Mi/+yGPMcMRvHshu7LP1ivOc30a8hQ72qo9cxxijDbHxRe5VQomkwGB
0yMhLw/KxXlSmGH+gSi1171DrdcLQ39ZVrlLyKLu82tUcOmP18PkZdmDCIIf4gh5oyPpH6k9RNJH
/YH8mud2zpKCTpUiZ43d5QnSOCqiy7CDSvWK8flOwM6/ezkZRK0Ld66rWpZfRjk8MPMih0Nf2aGt
S9zEbhBRFFlIiUquaGBfjxnG6cIV4oqOptHFvs9WaVF4HXV9QwcjoQ8EOgJiOv5m2wKtQq/iwfo7
zC7+XgmBJ3KBcL8ZM8PWE9g7LTT0hITzEFtPVy+rFu3Go87ZXlJjXYwtS4AkQHdAzSlcx8Cd8yZu
9PZDKKaUxxLWEi0fzl0GKcEM/lWuCtR5Xglf65AyFZYEMdcTGasHM8mYb2Vyv5paww9G/eN+yvIw
zxAbIzZCNnXhL9JwW0UkLX3EBuMgbENZ8tOirqu1mYPpqIenKuKBUxeUqWIs0FrXx/PEgtODLI/I
28aPUimRQK0aFzysDlFP22VghgC2M2PN64kepWt1ERinkHCHcmjJ+XGcqyfqS4GtILcbuBXTGgM9
aB3LaQ0okVKz54eiXUM2b6CMnI1ta1gYryPcD8sPsSH/+4EEst/7j4MOC0SX2GPLrzIWxi4ZFxMc
AQ01HKFzJvPWO5d4RVNigVCKRvYlbvoenR+Ek9JpRbT1SXqUtxHCTLLADXoW6ZOzRwXwMeVf9epC
mpB3CAwm0w+vaEsLgetV1Qp+079z0uQPzQXDLctVPUlaL4NZ1s9AiHu3zwGfIP+Ye4Gdkdk2IsGs
h/MFDVFsA/6VAzf6sqB8ltPVTwn/vBZylemDi3otnENnwrbpYekG+DD8UqNQExOI2jduM6cFVIkp
UndC5o6Qh2SNiF19m+Q1g42rRY84zX2H8tUvNJ7o0rtNt1Veoc6RlvtWhQuZsjxW9zqIxgtk2clt
y0T4gJznaaGaNkbQ4HiyEgz5N6jwjfhaUSz5kd/320y2ARo0eUCQcGwq6AiWpD9sSP7gn2JyPcOJ
Zid6biETUjKp5n3gzCPWdq3zorqzlePJ9c1OYaNsKcgXmK3cg2fpMRlfjdEzrC0RbCzTASpCbGlH
Fp0919vi4La5RgOlY8K4/1BysomvfNMLNBdtvj4Xq4i1HD/lRycpmYVPdYlXROlG/z8fPDG5ZM7E
dPiCWSo66x0fp00AKrwI5Kxrs3i8GDdO7ca1kcs/1/bEqaLId9kNPdEtDSnuRrRANdQ2ALqU5Xzt
k6NSEnt7hW8dyXLqcwYK8nOUOAsotzI+qIGIe2LhKJCQljAnvY2AuaEkKn2QIU+O4PsGJtjdiNOb
PB+Yz1PDmrfHYqsimwvpinM4sHhW/lCQch9jraENlzpP0iGBksVzsAYcYWMcktnvVeAWYbRzVPpn
B9Ytio81rlry9hVaqp7mFzxheqbr7tIr72HgK+ubYJsD17jQfGav+uyey/FeLDh334nTnYzqlwGm
0+HWR1eZaupFoiTjTzhKMbOQDZWrYRdtsFNWW7jIFoGFnhCPgk3X5LoZc6HDJhdn+qS4bdnFatrf
Wi2cm/QwUCoCgUzgWz83xezYweVHpitRs6eWGHjuTgI8oIiFtF87bHXno3ie/yeH+c396XPYs3Ps
v6N0lWPoLSD7MJHW96AIMMlTNdJQLYFZzge61x416tHUheqEv6FLlhpEfZP3PRAOoOXunx++gY3m
+74Z4u8miGdqrF1ur3mDbulDlrMZ94RR0Mfg4mY7xxlukYs9zBYdnsCFT+VVsA/Vd7Dlylmjpj2v
IXmncZB4gnBXiqH5GEp6ZL0FRGm4LkNDy7efoqKPubsNEXU9m6AygV0cw51ewrp0aif4T6buIMik
Dfh08mUSK/nSGeKf8hyJhBhL33oCJv47750WZ8FJyPfxxD0E0wawOAmPj0dO7cMbcuKJd5JZuDVz
lyGSRmWCOufhsrL4jRozPtLd4dWKIh5CmWd/HleVjN3Wv/C1yepabj2R9+VHoV9LVdQ4WsJNqyla
vTwA/JMCIix5rniij8KOuFr1eW4Y7Pvdavbedbj69quWb52L5psFzicYU7c8w0nybQgpEnoG+Sub
b4/OE5gVWvZUUJHXhXGAMAdTkTJdXQXambgjwCV+R5UFabaTCXu0m3MHdRwG6eZjeBzIYbvB5rCr
H0oyULImyghRylrUqXaEfDgyS7hjxVE+GBOod4MvIxqT+SGKJKk250YPv/kioBjfJ9N72PgoPW16
//UkuqtQ2nmVIlYgIY33YHAh8TpyfNETIuYrzdh7amnIGuYbFy2bN48DFSliDbgRxpjGhkZcUUzA
shDssRmjjvBpcLi1rwOrvvZdCn9gnjxvZs3aPLB6C4l9bsp5ElaC5D23B3LQ1av+TTe8M0nPNVm9
3jzb7DR+t5IlVk8lWEXxuHhSjNYN/WIixQOWSkkUUuYITkx/GPp2bImcQCddyvQXgfOUH++WMPeY
Db5gpG9lY1i2CdW/jnH8L0brh43/1FBkjLIvBH/9vjhri7yZ3nEZr0d/dz2jyNwmfYlEFb49kGh1
7XpAN1h0b0kh+yfyY93/JX7oj7Q8PKFeaTottYlM3qvL/Q5FEHHTuJSvJaXKSuu22/43JVeiUdv9
bW4lBOrHqXnfAFAhL/fIjIgsaPmdxDX8QZ0WxGfmAOs5zqcXJjU2ycSAEJLn58sSTc2dk52aBC7M
WM42oW+OND0gP6GbJyfGorp9Dt04frhTRsCxDP1tA6qvaEu12LwDvMmMz4375crd8VVZUAdhfB3i
mwS2PimClRytF3ngCh3MFIfUeg1dkmWExpM4LU8KyHReo5E3i5s+qQB3bDQsOBpE/CZI8gN+CJyL
pH9Rq0+SquwpxX92GvZ9ByVx19wLPpbYavteeBuBMEdxoy90sHfhSCuHS9AB4DfTM7tBUWIDGxj6
noNpIkonhh4inZZ8FVtCcoVcofg+qHUXI3TzNierBEy/vw7QEVtLZUQFTOzm7GY/4dWpj5uwlfk6
WDTdbu/kUZym1fVDAiwhg5ps4w8thIW3uq8XVp9MHf1yDL3Ufw7X34ML51j1dQKfx0UyHXP64fp2
dgDbnE2CC55iU8os3psQDCrXNF/e/0x1dg6iaKKf1Mhtizx6UW8TxQb3uOKvQvBupyq3nPx0nfZz
FV/PtPigmFSsXRyg4cW8RplPee1hBTTd6v1WzgNWtzTggZJPXPJF33fwwSGN/Fv7Q2F27ULDFXwK
jaSboQs7pYty2My9GXf9B2N4s0klLHwNsdBsAKdhyvg1mnAhjI9n2mgybLrWg148UuEbHaDNL2XX
hHXahImjOIup/kbfmsOC8vb3wpiTd0wbLl63nwtzNTsTwvAbGP5oJbxjfWrPS5f56MW49tBx6++D
jmWRiTEBa+XKI4dIGlMimcAM17gbWtgTZ8s/WknwRGmUAdeUXFLvEvYz2IBBc//VyzXfJRztiQC8
aXK5Uo3gleW1rjqw+Gonl1Y50hcZOSrsvtIgGycF/j1PRJTSeuW8yINs4BtDN8Yrl/RVHBbv6IwJ
AqZ4HvtcQnuI5j4uYYZCSj84VT/wfk3Kf09UFx67FzhwQ9mtqBkYwhKpaW8lJzu2Qw7E4B1t2w4+
L7xS3cbYYG59RIIna9b7rrZpzPmEvV6fgSnL6tXhzJCUrUBwnFHTRnzepKwMIRpwXB7e3StcivAH
nQWx6qrBfPWsiXEY/JXRjYVNulUMdnydKMFqZJ6+DAilMCCFOVHwBMfdehDNcB+lNZc/n1DLxi71
UAe+z2u/9XiCN8VG8TBihrjnrqBDywiCqHQb29oZAEgtjTvAh9osCEDFcVCtro/w40ojkAAm7/Vw
LXo0HMxLrgyMPfKxteWuMjITyfO/Lb/h0PtyMblN8nkod71dIpehVjYFnt4VPC/Tc7l2BNLoXjsV
nHvIFqfP4uXsZ+L4GJEAPy6NNgiQlZ7KMCGnWKuENM6DALOx1/cy+FvJHqNnRNEHQo4zPHxbPLVE
lg2G5h0NC2SyCNFHEEGon6DFy+qCGHUazTX6RUegOUUkVQ3+Ih7mud8tUhPxe9SuofFk/Wl/QSsq
SLJmTr3hoL4yd0upV3M4mCzAHyA+v9AVFLgCLanBtj2dTDCEI3b/lMYfcQW1xRkXPI2j2mrx9D7N
39MapP0x0CDV/lyGx/q4NRJPkNBUp3qz2eMUNvky2e5zO6Beif69GFZJEsMdNxYvqiz5zz82aZy1
fgD//ii0sAaA3M6zJHeakH7cIPt+TuRrbHierk9cuLN9ZQbBHvLT0Qihe6L8AJqM2zVYlDUuoEjl
aQx0hLdJw7LNw5cblWmqQfiiqu2u4J5rf4XMzxnLUx27iREThH0BbnRH9ULpZS/oCyUp/vX/v5NG
yH6BN+/+P13LME01IIHyg9BHVYjJAIX+6lz/fPuFaynYbrVd/dMN0GPrJOIyF0TpLwZz/BRudXo9
4gwE65WWCtRzSWnpHL+WFfB5KyFNwTmLyLPeEw/xhRdI393yQQne5o91LvcCrHfesDdd3v3L3WBb
bjhw+c94mBVdbEjxZpL1LyKYbEmnFgwq1rzLeLkDCvP49mmxbTjiKNnp5fmRLd7wooD8mJx0d3Pg
0F/vuWD9RLYTpLc12lVPINjRR0IP0Xda2UuOjSiBZoRFQOQGCuwlnPue/OJHPLbXRYAC68cojkHT
W5BfDMKFQEZXmixpPHkBBuN1HOgSETJNKvHpOWNIwxM67WVZA+dsk+8FU96DcHURPLJbv4PuCgfV
7WFH8AKhLdviAzeddsvViB4bfrnhL1fP748Pz+wiT3BRtr8ugs0LIHGgfjl4XKyAp7f5SZSXNy+u
1A63l/bdCuaQr0Os4ojpLkFDuX/t9qBTEfJJrbkRfk6DE27j8Xn++3qtj/lja3XYa1bIlzVBFh9U
wZ3qf9q0/+ai5ecjHSvrNkynDJuhczlonpN+zUSdxSsAxKy9nHRpPhyLu7gDvrmN2nWf8lXU6FAa
Gdjt8wqpuxQptle/lQFO/+ua+q/vpXKGsT+mhcJK8ocNkmxQVIba80cFtuFj5uxq6GxtUPkFzvfQ
nihPayhNz1uPtfU4VDV9QY6iVrHgViriF3eVLka0KTvEDK35EzjUwhyXbcsKfhmRg8c2mI0DV+uI
YpW8w/99GDesJKo9kBvAw+lrg1t9AUWuNfg0//9GB6IEB6qliW0lz0xlHuabcJZKPTYVyY3FFXI0
S6XqDxdhQp/Mr9LnThix6j1yzenIx0Fk3f5NlncZhBP2GBbCVy8944/dO9zUN/xAHVo3UudgwmOa
+Dw1rQHD7r0TaGOM/D3KzK1g81BaoRJY6Gzu8v4q6P/pyfFE8nHIxYtgoy4NCXqxpIJlt3qR7Nfi
oe6uX6KZsXlu5iLkOzSsHwHyKExdTSwcq1dlyEq+uF5rz5Lz6MG0BW7hUo6nkvYai2rY1fWPKKDH
1HmZm9N5guavF53V6PgMAg0ZlQkcRhv4rr0XPNcTQbeYP8hr+QaS/combidQP8XEf3uVpXy6FL7U
HFOf74q6UeHnpZ6R1hxq7Ua5LjGCol7MwebY5WPXiel9H6DeohIGR8yZhGYVXu+mApWQeHONS+kC
YUYNy8KKKkRz6KZduxj9rVJ3J0lG7PexG547L++ZswWasG/FeOD4DyyR2N3GIUySDpzf3/t+6lM5
V1ftGthMJGywdkiUtitezGBKxEZ7ZBlMyDEa29B59zpER2T3GvkKJyq65hB5JOML7ilv/JsYyBKN
o/Mewdg77x/dk/0DyCfv+Y+urE3lpOfDdFEu2TRy+D6pVeCLJ/XSvf3I6wlvxCjiQrr8FP4QPTC5
XW7OCAmUHfBv8oyJs3hhUOrH6QhH5bOdjZdBiUOkwrLrY84MJILNv8QAlYzhiqotnK2M5qf1QO7y
d6UTHBIItNqHUPEiLZ1XhQvqPzzY0RX63dcMgeE/toOkAsGdD955tuxrqF8MX6qKfXJIPWvcljKg
w6jM3S1mkRp/Z1a/nCSHxyFFpPlCKtZv+BLMgHiq/30g4qnUElPewcu53JPTkjZdH9yAJ3H9xbjc
nMQQUa9SuBEtjgE9LgjxtYa9hidKuVdbHOdjThM1GmGdk/annv4ZdLBVBxcFFgwSRt/pO5Rgu2VL
/T7hON4adDjjN0lD3G8N4yuXnAK8qG1Gvcz8qzrJBT1rQVrdSTe+MssMKSZVbUwyN300CSsy4bct
+S7ycZG/wgffP5AcX+F8MuCblC+7z12sUH9BlI92RtfofAriBclg7335xYZNhF+jO3A9Xw7VcHYs
jXyyq8mdLx7kPbECz5hJqNDoGn5sbzTVI8rUx/FZIm4gFs/xVySnLE7OevsjifLXLDhGvZqmkVwD
m+LIRalR6H5PNx8kQJ/0HTP30zEhGdSpcFoLThyVH2SgC7iiJcO17CVZ3fI+atMuF2idOHPP/K2y
JaZM6PL41Y4+WRKH5LYhNa7KeuClEFz8OXpPId72sunO1DJgeO6pgH1oH2zAxO81dejas7hjhLZn
w1lPVrUZUmaRHtioS0VP9oT7ZLyY0Ml3t+A0kV1fwUQvIRD39xbky0hDmPyr+UTSO5eocsqFM3qJ
5Pg5PenNcFC2VsWeaHIeucexBiMqrt5FmMdbAjNAjyEDfb19FrF9/oOUyaXRsLFM3ZvZQ/J3/+Pc
0jp0XuXccLxB+O+frd2178YDQeAPdP3HvF7oJP6VU9wBYxgVUmx1YsSyYVdZdnTNFIpdvEA/PKsO
WRusV2XhYSPmixcFmfb8afTSziPeKZqFdjd2hA5G9GzCbJDX23a5tFH+v6ORdfjKHlk0DmwNeVTH
pT/Qjv1lm/NH2Vd58z4s6W3sHavH0iGnnH6EdhfbvbNx6tn8ED/ANAdKLpjyqwaeJvNw/gWdFjoD
7tuF7dTek4oKqGk6CMEVjG+4m5BWO6Bny+iXPkS6iEdM1P1PP44y4YER1ffRWMR7fKHmbBJ3zR2i
EhJVDBxmMIvJzu0scWx8knr0F5vypRPRoYNSbk0j6STLs5DmThbPBZbsz0h0vyzZiJ8Fq5/PzV45
SVHmHsIeQMyWYSiKzd4pNRZthInRM4XxZ+25qO3VX5sOl0yp49GRwL71C/tbOBlfDLak7le+xkpS
aVlFRFEKXh0XClCirsEAf5NsscdeiXzbSL7DmXY7uJDJps0Zwnj9YCDoVwfvHGtkILIzJzAi/wAI
ZVGhlP3BEZtxZC7N7/4XNagF6CvIq0EwlKHcZqkP3u7TFpaEYQRSNNNaqRfuWih6LYQC+dV2nFTX
CQKWiHb1QxJsy7GmDDuK2Dto0Xh56DJ1ZP82031+RxIko8bm832jidDuF9qf7/x+G6yH/3S3UhGO
xF7GGp/giZDSdX9bw9YaS1GKnT+dUZJ5nv/E8UOr/QMorg4ktHflI+h27QUXRmZrw9AHOsTQZY5x
2psQhNqIYyJ9PuHopPz/00aXZZ8vdCHcQi21Bc4Evve1WnI9w0KRSurIDyaNPnHa9FaioxMV8QAO
YGcAP/GmltQriamAiQ0I/1MBjBoChy9HGHm+x4sdi2q1S2wHBm7vV76YEh9PiMvEnlaKVKkNT6uc
LCWVaK9NEPR6v/batMcN/t6dV0K05j1Ex4KAS2EqRxlQy0GgaAiQUGVEwrakeaENiuUJsc4mfeDC
01hfIos0MY3J+RiJVvb6peJbELiausZs7T7al8IKq27Lt91KEYCONCANSMgqrwzFJpaXAxgL3j3d
+c4OydG34OqBv/ErKTskVoTFXQv/oC+9Fu3z7jNYSkL+ND3HpXy1JuXCTU39co41ww6o5RLWHT5J
GusLphCyrTvfQXtnWj3jAOpvkmi7vPThAZrqhGyhHWfKbN/jayR07SiM+ose8602NxBMv6hGwrqa
+3GjX4OU/O+3yky1+Z8Wo6NB4bc508qa2Nl54iXOjNe2M9wmtJ6fdPm8/c+ffGXnl1CqwG3SW0np
FzlprmjUiQbGYdIEyphToN1BQofZzRQwDzXtnS04AyP06s/q6rLWO1em8JCOyt3bk5vYXD5nTcta
J13s249aeNMFPfQqkxh6HbEqGC8TCszJWbfDY0C5AQd7HLX2Ta6kFPRl0XDaqAxpNPrMTMEpSRJB
ouLT6hyUvL2L+St5ovuqOI0lnBg9g7v8OoX+rCFMAhAEWz0Oiw8JVqCFJE91GTsE8Qx5pzclLI5M
xq5mgf00NDyvbGUom4PFJG9mfs+ULkHlIGT7Q2zsEs/JFH1QqrUm2gnx8KtaLKoAzfLux6tuJiwr
QttTct0YLX69Wm2eVMXM0ennZH7BPXlahJxjDjMS2nB5C9eXm++LT6kE8Z/+QxwGzvSn2981/UkW
la6sC7TBc3uvDvrd2Fx4RhBkC/bmRdG2sXCKk7b7G0ISDF5ZrgcI8fXx8jKI9Rdp4sg+NWEsJgHR
XPbpk7x3SnI7fIXEK82MSTvu/vofpCVKJdmdRffUCUhlLa8MwCxOV44OZyeK86AOt9WucZtBrdZq
rZTflKrFomKUzC1cGQMCMa5j2FZilf4vV12eLrQkQ8zLCk7GwfhN1+/BUv35qbkps5umdBBUtOJA
yCujUmbPFWDbFP9CKZDMjx+xuBb/2cMw5gvQiXAk43bAUuLhNYuwR22MZj9Z77atCYiXP6ds2Zx9
JmifQxGevh/SC6z9BGS9RFe6vKMc4zaFWoFrNjwNiF7MDJlcFciUaSwc8XB/W9YuViG5pbQfpc5H
xKbopZLkHhtgIN6PrG3ksRRQDqP1VgTqKma60lChdegbDqv3l+c7ydUV31Rwg7IDQRxEflFJKkEG
FTMiTZiZbfjtcbjidkkEdkqdh6kBo7g41tH4oe/OpKTWxZTYW/U5yf/OYf1aHJ68N/JhuSJwuDd/
Kvd4Bpi2t4Zm/NIbz78f/aWB3jgBiqgSWtqrTEFQEtMoBS50+R+BvLD9qOlZoLeSvf2u9JnCGmpe
v7VpA9bp2l0x5H+D6wuIKsl24vLkCXVdwc2K+6X5EQMDFzJp1ZFq5c9H9Y2+BcAlAkyRVGHvbuyv
gRftVfkyI3YG9HuoMDd7i1u9sqdMV7Mbb6SbJWgdyfkG+hR6x1Ajba2O5SYacuxoe4//9naQFySx
beNH0CkJadMt5xLeV4prennQZ3vKM0uR39jyp6EBURcKkg4YCtANDDVhKHbFFaAoIEuEeocrNqgG
LQeWKd08tUJ1ITBs9oGPMJaTxseJqwfPtsiBZCPSCvefuxsiptHhrU4OcndUN6HWvq9WiFvQr+O3
Zdl0l3oFSQ+3o5ftuDbPleBFAdkzg7DOkUrVyh1/9f3TonbdPEGnFBZJUcVFtIxtW/vXVmiuEqO+
v6zODK2pav/jD30fwL8Up30AlBMZ0VgoLu0n5pWMvAKx4lzkTa87oEBZhIQzaJSPyfxYLmO0rvQX
tBC379XfXjSxil0kAjKObSVD3cdClT+ei/k8fYR+D24L9yJSQdP0EusdQSiU4sUZ1bVT6Ape2okg
Hz/RnAv/0u9XgR9R4QMjJUerWFKs+XHoPOpKnsSxgnJQZxUgACKoDAGCeEdN/saerhO6dRpmqReF
rZu9lUbJ7MKnGpPANFqingvtZbeBT/ZUpVXHCt5ByQfXCTbaOdezCd6wbCZgFWn88fXf3dE2nht8
z5W9uFIQcSkG2/rEUQRS+FDUTd6gIDZxNORAi3hO0+Z5f08eU8oYIyaT96gIaSPQ0swkaTzVhtBV
njbU9vUveXqw/dr5XNX6Uq3mMeODg/+UjY3RiGmh4R5b3oKW49ZpddDlRIIFTDHKYx1b1eRaJUt0
WePAJhZf2isq5nN0zv8iL06ah3UTmfzZmQ/si3RC8m4HBVWc4bT/lgf1pvLVVCesDljW0Lmma0gr
zVQY51dcHrrAIh06uO+1fuTee2XbdMvO5bqwhV89/0K154CIVP9rdQceJBae9T0ci1aEUI5Wta5c
XutnOnJRefKhsrvIrwwCJVZB9UaWI78mu3p8vQeBVvaeEGCH4BUG1qjmCY8FoqV440fM5LhrJDeg
wUBIaw3MVgvRXElrIcns63omgp9v+ptVkGuOZNK4b+CoQVprzbjZQU0cNInEdjGS75L+nLDnYOPV
lAw1mgBDvOE67uppzHosmIVSjcMkba8kJvd9ao9mY/32RJko0aWiunGzIGiNaT88CEprRnn7jvSr
vUvb4ZWGP/XOjPdwNOxL5DsrIF16VC6/mulnQSAaN2wjFTpqPU/XPpTRADmfV6y/HrOmyFoPikbk
t96lyr5lFrDWo1LOgQ0NH8b5ymvoMDYo+x6Jmng9203+G4anP0S1kE/tvNyosqvQYtT8igZGbwtq
uQRnDtXpA9DlnJHAX6iY13rbPVn+wFC/wrgz8sLe+4Gx5shh82eaJyRpRuaajQVGDUQ69e/i0oXM
FZ9JNkF6nBRYq/BO3UMmR1nnWqLosTe7KW3l5aYouWbZiKGpBvHBioU4QurZqHinCmXX3t1L2UWi
2EDNTLV8k8EsJZjRTk/5qR71nSuoGSpWcMVVxr4mndMYdKmWXKs5xw9W9hCIocv7HPVENv/Df/9H
oD3YKF19uoEvtt1fQM1usQ2xXx2q1OlcCtZB3yDmQWJPX70aMZppL2kgo4I22fLdvLDtRDc8WFjU
FrppLcgpadGmbHqXt7MqCPus3ZMtYmnD9l11/yl1cxqTiLN1qXlOTyrtUgFTUplMnPc9hwYhoJ8f
DZSYDgL5BVcBt8EQo+v4iYNsCxk1wS13NgDb/81QS5i8fB5o4LyTu1tkgSReMcgmmvUKlDq1F//6
iaOAq5sAOgNH62tHeYsp9LKgHc1EXtvWJTBQKk6uoPJx+tIMattpciOnpFe49H748ovkwuLDs/VZ
2c+fcEdq5dRkJ4Z1gmlQYqdShHVEP65JJPDBmS0rLe39soKYnxaC8nPzjwp4CQImt7pH7UlYGCWn
Hy301edpfnrKhJJXgf0KeYxTwXGOrsrU23BUPOVRTXit33vs1T8RfD87FOCbFj4CZ4528zdcunz7
UxLohjLIAq/5bLe6PP1ykw9Sl3Zf2Arp8NiY1Jlu7/KM/01QforPYm9nHYa0Us0AD2UY2FOhvz4n
i5bbpihtA6PZfVGYplDg9QkG264TC8puzleCgHheJ9pyKM9AN0F7sch2vP9mAZZouw45gV50Ikvf
V59UqbQm6PBjM9C3YwbXpoUHEFCPaPvcMBXGuPUbRGus7fdZsJ20nsJgwpHCqVH8m5f53M2f5+eO
e4zr6RnI1QI5yQpw+16uqrxVPXRukqHvz3yVeWCj0H4V4xwlpA560m4xJki6XZOsrnrZgEa73aOK
n3mXO9J5e4Rn1g8OwbVpDQNJL+fHUIEsFq39PN9YFEHsH6lR0TTx/Loz/k7m55iLvAeRw/hzB5dA
h3X7JtfOTx3KinpWtpdzwHH/jDp1iAmkA50yKUJXjuK/6Cx6w4K2pRB1+Id0mgthL5g+tvOsC0IY
glVVyfitlSWdEVWV7nm6YJIlxjyRBwSmZMzBiVFTWoInOOnPBKZkYnjGqxtYludcezCni8AjlJRn
8RCulJl+UIULsC9Jl7OuzpNMKY2+nMSLh5gbpB33LssNCR/0J8abShhvDRpifN7B+m4pduL6jLvf
pkd52Bo7Jg1V+JRhXVbxe4lbfwDZh3jG0DblHxZ7ymw0Sza0zIYtPOnFd/oSGI3noYocwFHblJtb
2fgF+i6mRTyhEd36OGltZFix7bFo5BaMd4PuUKpbNy+iZ/S31yhA3NGSmHcReW8cd/kL9DdhZbP6
LyQh5LuIF0LWk4qa4QF8Aer2w/0dAkVEjD9JjZZKSOCCaVStggWaPDFbAS/ntOzZmxQYUnfJmPGg
ZB1u0Epr4oEyX2QiHHfJ+jHujqvnOQlYlww8PlheK6JL7EeKHyu90I7SbygJGzYEY/p8J61XNXPm
5Dj/XNExGaFmbKCmFWvT+h3kAFGegtz44uIs/JERvUuc2N9vg76x9lIlzjEwPprTBHRngUePatuA
9YTQCFtySMorCA3qwSYvaP6nQz2KabWnE6NSe5yeEnYbr8XsO2kZrKD49YdxYIe6DiSfexk4SIYD
TyvvSyW0fwmYXr92tBSL/6CH+csi2ddREae6YtMpsv9ahqWeF/ac0y7admVQsKd4bDZ7gziTNJDZ
e+74FtqLP+IX6gEWBPsouegnqIskcpBqn7Qxn5VMDAhSNQlvJ6MMvRvRON2G+UqFZP2Mqx8CdF0X
TbNTszFG6wlf0K2apTow5tAhtTvbQPZzmsKdzjRdKC3md3VKyzQ2VtTkzUvdPqoU11YTIwsAnYPj
hGmlBhUgHfmabfktNeZIz8wAttAegsa6tHzkWe3/TFBDn2WwMwTsAIYBC8NT6Rw/n6qcpI7hwp22
R8WSawHVNmoSzKJ2u1TkqN7xIVJuO677nJI8DFX8tIMD/2nS0xMOk+3moaX2nNcKlp9FEFcRSCtx
W8FnCWH6q7F330nLzCI03fVe9VJG4NXqel1RHjKzYp3ek7REhccd62j+Mi/inb8fsxmYYFQCtymz
8wr/+yCbqjV+SHi7tv4gP/4l+Sk+fy0IPnvUpXHUSECX3REYNi3GcK5d+2hyk0IemE/DBwOCgJn5
SDbIULO/Rn/ZzaNAm1+SvzAZtexVHcNrXzp/70TYD2dhYg1F8olGrMBzM/8w01ZE6jWchl7hdH54
pEqSUrTanopQ5YhjEh5Udnj8fLNl00V+171nITSRinWDH7fPiMis8ywY9q7+CZCgZ+flegDfK7D0
XwXronY71tEmZv6Vem5Mi/7+dYaACKDBpSYghdIMB6bQ8PmVRBsdIoOSjoUun1yhTVt2eQP4MjW4
PDUjft8r1T+rKJOFBBfEa3Vr2TbxlIx31nLnj+ewfy52pvTD820iw6UeJXxD7N9v2pd6MMsfmDg2
OQVGOpD/CxoH0fBYYKXbpTuOhRu7Lv3wRfQD0jo3ATOFoaghumtdUzkHT3hucDrZ+qZqTnceA6+X
zIHemENR2/noSl6o42q929shpgfpifur6GW5DqtujubnQnQkRYp2BWyIdu1PYI6SfGDLNLr/JDVv
ezT+LyBnaMoUcd7JEi1iMrrq7/w4gGI7FS98ojXyzbNS/qzp4d3/flCOjzTfcXfpced1xYa0xuSe
Ja3pZKP3gkudhwwhoC3tKjk4zRA7dLh0r4KjShLfLKOoLAdgDQ0iOHbiglDbDrSjo3jlJ3WHP/hd
LNBG3Ksg6NwtsQOkuP/OzybDCXGKqAgSJqjLQkD6aPf4eNX7zx93bgQYUu1+e8Af590i1TV7e6R9
VV3G6FNEXi/7n+6Btp4J/04NqFQ1ztK3Bf+XI8+H/TCwdhspDQpKRPH5+mdoqdVqZmmIuTp+TY9L
oIKUHAGgUZYn6LvAHkqKzjv2099Ptu1+RYIFOFWqlZKamMWUXoupr8aw6Kqx/rqKj9xZ78vun8ot
rqM0OZ6TiQmk1BAI6DnKZxXdTOoVYt5AzpkIhUQ2AngAOHexOkmrEMzpo+Zu54Xsp4HaRGjCdE0K
us4QX4i+/Iz/7zH12dbRXp28/WSeCVEJMvI+52JJjDcOUKO5gxUONf76Ng9tvGuq7lfLo+sfQ2ta
W6Yg5z9VOJZE12F1/09xWdY7a3GfAHqBZXTwaChQU0Wbo6Dxp7ZYDqvQdzm+dlZp2vLdtn1Cm4WQ
lzfoiBhVU/5iYUtQRreBvebZQmytmdxaXX20+I5hgTDk80TfrkjAZRxkH8UmVu+/bO/uvqyE3r3O
BBB3HU6z8HVDDJBtaBegX8quG3DiR53Ls0CvsXd6/Wfks20TSHP6NmEvAfNiAAulbsi3k3KUsr+1
/DghaxNALGY5liAMCfFQ6PeP/pyQZ1R62EtVDWKCPOZJKEQ3yzprzo7i2Ztl9Da3YIdLKftxKD8/
mANGxVeORMnHS4sA8dn1RAtSzQT2a1TVJx9Bx7AAIcHIthTbe9W2wb6lwWSjs9y+NaP7PaUJSAuO
ZZa0GOa1I58KuV1RpvQRdiL6k9MRb1IoVPWgKdRHBfPCjOvrGpx4waa25E2G0/2qZzLuRbqINQ1A
J3nKWh/fLH/gwNSvuFF9Q9gKmZ+M+9kx0jq/m+5ME6P/2qqvWFVlu36dKsVrF5ZB4eVdyYLpyX8H
jbHu0tdqjgcF7iGJNTNDTiVbKI8w5bqLuq8DzALNc9IYImvdnWb6ii0qxIoHsmDLFjMLZKHi4h0N
AZgZ3Hg4bEADZ30YcRnu4qLKLU20+Typjrax+DJD71KfcGq95WBYoTSHOxzp9eiZnSgu6hDAKfiF
2Mvr1lagd9kVSvR2ucK2V8DEXT7PJfBsO3hkrAltgEzmrIghiCLHtHAAeGFbWNFEBHnewe5RUrcP
cRpde3E5+KFmIp3eOu71cjOQwU3tDUtmPgg+1c85r4+CS2q+4H011IcXVNmSZlZ959rEFYl4+RCp
0Nz1qvEa9QTjANXzj0gSeLiN079s4ZHtIOOyDUhlnifGafk+AxM3xi4eqGjiEq0yA893KlsCA6hD
f00MJaV22oabWj7cKZfFUjqU+tIy6l3/L5Vk/ld4QEBLNqPKWIkLUeNf1BFQJCb1IBe8OOne/x0q
NAkeqtjxhqQRHqiUoIxpjOS7LYcuambbhNdrhlFCa1+Ele5vT0c103EkOxjDpe3ywtPpKFszfMOO
Ks/5HUCG6knZ9WmAuM9CjWpYsNa9VXpQmtUa7hUHZYqWuO3WwNakAneRO/Q59F5wNtx9p5sRRASu
Lg5VYoqwMJQcUg0+qUHVIdhaBjpSmYmFiYFt9JvaWdyy8Pz9yZUay3Tm+S1LA2Qi5+GVxFyky6Q+
NnjvcLxY+rL7RKbhdwmuETQP+BejO741GMUXO+wja4SQV/tDd8xjQIlJOV9mocYO0sN0oeX+hUOm
VRuz3H85kkcLTrR0vTfMVWoolizrBx9pnSBSAqzK4G6wNU0psqaSpI604EgGvjsK6VjKrfpHETpu
+33kvNKRZeXKGFuQ1SbUnMuKGRhRsDGzZes5EBXhtzU752cg32VB0nVDR8V1/kjZBONZtEdnAvzU
UBa9eCcUMy8eVQTx0esfSpHuhzLAXAu1V0FYvcpYYRglEiC3NrEgH0ojFyXS1yvgvgq7KZLQNJQX
FT6zeeXNgvGdwmuvTJzQixYeraM40pZ00hvNyA87FPItFXdniwjrOI/LHYPZ24Vv4q6hBDx3bSM3
KgR6ZqSRFaZbqicebphvhvbJaMEOC/kDjrBynfjow8T2hzyW1zsGmL5lED4YWpeKKl4NhJoBm+qx
4EsTJehSgNROQoI5CAFIL1qdPwy+oIPULKWJvenq8HoNkRkW9omDFwPtMoUElyNjlVfrL1Vd3DxD
eQfWKAFQoTiFI7GiZkLMxJFZMQFYieyHQ4m3XdicBOPdkc0gymiMF3fs7IkH0WqfBNgHyHN8tSZE
WfCdgT5ZpAFhMUd+Smyus1Xbh7l6Nc7p9/0KpXIIUNzKsqmRY33VHuVCeK81jEr3XpXsmCWwiA+n
Q1gkllGrcOV9rCUsR0vR0jtZCFCOEnsLsQ95y6AxuZIUSLpuWEJCXma0Io0n6NDSqT2vayxC5JDd
zs5lVAxR+TtQFr0KHtV5zBM7nqMKgqD5Y/lKak5yygPHWSQ4/b+aAH5OTXYiNsJU5Um9Tndwa5Dd
2z37qTGU41rwb7EsaXc4aj+OQqr2/IxsL66wb7s0E39QHUxglMsVYZkr3RxlCMWl/gCIsgsY0osi
kr90bF5kYF+hvjR+MiBpbmpx3pAwkou1PFXH01jjC1XqeNqxen2MYSP+bXEqGztETw9t5E40pcfI
amx7jb/dPPQSUgi5td18JD6a5TEzwuJ2EqqbMp4z8bD0RRQ5m+wMi1f3paVWosgX2d115FVujQUK
AD7TNVWBoByHBBGNi74Iq+oSsGfprjmVtlR04X//Z4gOddzRHU/zZxwZRyQ90zhaN7HoNV41OQT0
Ca/o6UMA2r+uD+AYz54/YuPqNiNpgFDdh7U2N0t4Eir9AbYRMG+v9wvPvTMjcqK1KCWdN3RXhyJa
uV0G+jefx7wK9ELHBQZkvnin+sMVV3bUfHpVVtsxZOIO9/crdpEo+uFBuUnX2sujLZmyBKNXnOZA
MiUpkj8e5E/Y4NCN5yvvcBrP3XBnO7V+73QiuTLraQmz+rT1BIswpis0W6qMIO4zBXjfST/7CjAk
2YAxSuilMNp6MaMGpnV+HajWljFa+QuEgyN8Ltu16cDBqDSTOYnplX+U35ekxkpC695G2eICPryb
SiNpnwmb69n/EVYi8lWoz9hN6u0BVbnHqFTa91G7Sp39A2U6PlaobQdQ1jcCxy7X4TVpPNKAFzDi
bcH2F6g5O8tSQ1FsDxkLvJ9kotNt4L9NWFLFCYXkG5tfkFmgW3P0deUgW6+iaw0b79wS2mNSxJ5l
9ay4hF/VWauH0MsJPZdb8ArIGJg5BuvU4A5g/RTGeNzZGLRBI0Fh76K7W7TXYWQuMNleiwo2moZf
I7QFvZpIJLA+OMOS+pBvG3bZed3j6wzhk1NzqiKhmwhBbK570zokE67Axa7QlQpjATE4qnsu/HOB
I80sXYtjr8NfwJWqysHhBhmQbSKlWd1U9PZIl94jxh3wcjRIwrP0QsQXAD5KKM+EzuVek8brGoVM
SxpXP+bh6o8ykJQOdlAewwK5ViUEIz8Ez70IKuKKYNddJ4stp95lGdN5QSsjHU/ucUjhqxSyMQ7m
97YB2hsilDlM4vGUsUPmq4s5BQ8keiFpmS9ViHAlnW9nk3DqV0Mf6tBzIMatlDeuuLCcxqUzUW3/
ikIpTCAym2PUekZj4i+PsXClunNAfcI2Ys1uKO1Tq+mnelfHcsOAhQepVLeF7e5+c76e8lgAXchr
ueNLdE9WOLkzTxMQPaf/mZQ3Qr43LCGEAeUPLJKeXte0NajB+gGMxlV+B4BJErCCat6W/Ffyi4I1
q7356H+wKYG6wEdVxdbRqIThtmArCfdHd35VdzSykTtDIKucY8MaNHuANiC5B8/fZfVtOVYvZOk4
lEg2lJJREhIXgDofTQ0CpwQGEItiHlzCUvZGAGYb5kZF+tc0kWuRMETFVgXk8BshTTsgkjukqLca
+icOStqDflnel3FjdWc252fLX4mWkmQ5cW7PUyPytBtvVMkzVmwRLSMbooiUz0XUxNt0+FmSvRBC
qI/suOcvj0mE6ZoUKZuSos4KKHIFrZutr75xePPv+Mone2evxZ4MXXGjFjud6My0v+2eCyvUAJSJ
ItVNc808p25SEGs9Or9yxHr2hDm0h6yszgHu7mhiy/YnWu+KE8zoopj7J95hHigUu+VmrazpwfOZ
Gnkd4sAFBikqaG6VE7Qnq8x2lKiOZaS8e220EluWQIqPnUUNgAtCI2/vA27W/evcSknziG+2+w8k
RZhxR87RPYx71e5NhZ9iVCshd9eae0JckjkQusfWNkE7E5ZDe5X+oqsIcof5DtYRrlpxXFKGExkh
ubru7mLog/8GWnvBCVWNT7zQati+gXU5vEhrG8LxERA8PyNJh0n1WfwIae3Ygs5Rpa06U+VTrFkU
VIGVUkjLmeWgFCdlrPEiRR6ulLXZKmxZFgYAec6iVtJrS29xEVWxvBF+FBThzqE5BENXr7UTaKZ9
JCdnx8t3oJmhiQKimkedM6hJ5RPnn2J1sBAJOUYkofWuUnL72R3hbJwxhRprE6k2iwB0lkAsJkTL
u6EdxRyNE1voYh57mQCaRkCB84l1ibCiZ86o15D3i6SfjdtGqcddutKLd7AlbsqvnW93d5sfgT01
aT7Bots8jviFMr8sZSVLOe0Zzr35rmNqQBwLB+i2T4FcnPeBTPWXrhCxAaiHh3RbSRPeedCgJ0DA
F3rEBIwPqeOM76SAEddzniLrjMcP5WfpYJ/VnYjrAAtvTWtZWgSjbrDUtYtg6CuzGBRWawH0zf3W
QVN6DJCFciVpfMoKKzEPw4MLpVW2tZpyYlCsS/jVbairjuVIvL6bSz/7q8sAydHZR4v+gcEv5442
0q0I98s0xIEGsBDJRbFybFAPxvkvQ470nwZ1uP+pzUCb1Qa6a15wPymbedsfcQjrqWPO36AP5TAk
DpC/16ySboLPwsjZAoD4dttbxXwfNmk9W/U+ND3hl0Pa7xb6LyOeLxwknc3aHk1uo6yW4Ur37FGH
fpLAfclysRotytJ7c0In5gslspm904qGKDrHhgCGgo5uAi96+plVPW8a6OY5L2frlAgpYmY/FoOu
TVeqm2OI0/ppePSzOzW8I6k9z7bbNN5LN94+ngvWzbHcix5YCC3u8DBjhE3/kZW3oKjaThtmtHkB
CQUNfMiU8106V0YUhM3uH5xhq4SIoecR7qAaX/da5Dj5nHuyx5VUDoku2Eh4iVgSBzlHKCBluqob
v4pxVplmaCwrPkQ+c9Y4hbCzFuZ8tygbklZ8u96COm2sXk8/KtNCbd4C7l6Jm41xJhUwnen7fNPQ
R6gyErsj9EiSwEN0LwBlomRPEYyGKaqRWGQ7K8l087+Fl5dCDiTUykImY3MmZvFu9fm3e5NuXdyq
IH/HD1WW/LhNohei7NgYPw9LX9KfgnZyWeCLKC6UUczZ1EZeSkCoBJVWh41fpBRYwEBKFSS1tVAV
mD7jZa2T6fWcT0+tTuMOcY1h8RpFRY7OB2QIFmpKDPYB4iMy/nUx9St3nC9LIm1gChIzkN90tx6K
9fZOJkrXL6V72NNbynjJmOv7c8ih7USub8GoV7prdu1J/yzh4sMHe0Wu0dDIzwbXaO2wXo6l38Hy
aQwCgAwEOPaYHzDpSho5mL61RV09vz4hc3rx/rxXsrUz7y88FJFs6ZesuIvzTONbMQ7Slg75vZ7J
BAxwJB4dKOYeQ15LsUF5m+Xrn/1xn7l6Mia9MpipyMsruHQLSUw+kXxQxOwB1Kdgsix8z40CWmey
XPGvnKpuWE6b8giNDxbsQjA2wnHij27q8APDjxg00M5nSrZPdlsDkGrxVRT9qQzw155ZlxsrolJu
kyAtHcsX16x3Msn8oCgwyGdyxS4v0uGDMuaI1IV28lHZYpyuE3HadvP/dUPcphg64NTID6scRKc2
/MMm9Qeeds9RE6jcMGk3col1gJp0n/wkxbEKk16VqWjrgpGO7l8L2jCMTOggqNwW4mU2EypB0MHD
K6S5pvqyVSdEG6IwRkU3F1RXDdJhv0PIkx9aZNYs5RrTKzcNNccvm9jUM4tvru2VcKNfC5SUJVQd
Ldq703rezlhtk35jXMx6D9C2Fyi0EWG8Q07j18kYWi/NPsZ+fXVkMy7mgmKiQu0anHzbBxBvs/EZ
X3EVqkMMf0TPxWZlE1CyiVT3l5F3a6XHQNXJfHboGgBmrtvdDht8KX7tpcVzMxtbATPtz68Rt2Ej
ONzMcoNPt6sXCN9MOMhi+nsNxh/9IuKW9coeALDk/9j32M/o/vk6KPbZwC8l7lEouI0a+c/rwbzl
V0BZ4RmaVctGDTmgYSN7AMWgdwdlaoKhVhbTqBMAxviWAMGizCTqxzGH+1nxqCdJiwNChOCht2L3
M0AjuuPnJcgMIAcBsTLPfgRDXlJXM/48pS68N3CpBWKLMUjo5atuYJZ6sn3IuQR0tAPZse6cdcAo
bnWzAe8Jbu5LIFlw7b+lpeZftZbGuDdjss35nq9dzpxPEfCiqJTVJhVNupoj5Dh4vm4ArMkqgJZP
iaZ4qVrRODl+9EGtoDeavL7W8VW+M5dBQwDkRY21R+Wk/wPhHCcyjZjxIhOwVI4UyvhItqy+uvYY
DhFbd2iG11Qq/M2g72CCsW9IYNHyA94SXdBuI+QmtEKwcBJWpLGB66c/w69X/9lgZ24+34kfaI2f
F41JXuyXv+8ZKv5gAv8FFCs/c/jb8frQC2BqmO7WazxP4lT0Dp+ZBJA/MzMMzU+fQmP/JUA5vQKX
T1cwjdeNEXqr3+hbcvHbornDjN56KPg+O07GkAfTBvRY4T+iw5TRjJUo3B3wr2Dp6NgSxb1BKRmD
uYzJ4IkVKm22Ud4OHZOY8xn1cwsKpOp8rwOVNxosXCizUk/chGRXsu1od2tLKIJkcSzfvwqcZXOJ
tUYZfTtXT0FjqA9l0bN96VFxP7p2Ylm/BTr6HF64bKQODvS7sHm/YCTCbpxv0HIlXniNxzY34l0o
AsenzvjsMyYZyl1sl0d7XtX1+ZPzXDI8KyxFsP5vjy8CeR9lCBYtlrTNx+ETnMO1nal8pIIePbrj
nHPqBqp0QqmLDDy5paC/4HXOXf14RCIMSF0K6aIL9TfgnsLbJV8b9gq68lUeXdOnI6lVSRwXllen
NVB2Da4aizVInrrqsOU6harJm5WWu7k+Jr757paWkZgPKB7RW4DEEJq8vG4G1BXKUORmO0LdhjRE
Iq1V828R8N4vXV/x9gw6ART2+27+N2QH93AvMhkgPy7hc+u0Y90U2Oaj1qpSUNMOh/WkdkTuYdMZ
B2M2UXBKk+UNsh5nf1BYl+14+NRi7HeDHGZ14wony4uReDUgDya12R20ZgAg90jMvBksvW5NNERt
/1BM65fgyTyQsJgGm5/hVx77889eYF18VU6gzsjRcFEpddu917yXQOxcA6MeuIxfmTZriGUoAm8N
bAex5428QFs3ADi8iRLG9em3tDH7RfjmByopSGDIo2Jsymh/4g7w8tow1AbWty/jcBZRtUjc6rPi
SfYv6Qj3O7LAcmjg6IyF6LQyZ73AMaAfW4cDOzQIvfKSxvzWqu1WO/fdGlxX1cTmw2NpSfO1UXuc
avPqeqdhqYLMh7x6sY6Im5hXJ9x8ljbalOGNDWu6JprkZ2KA+o2t+kynG/gPXr31c1wro3iRtH9A
jTeUvPM2UQwqg3F6eoV1O5jsC0GB055PDNrWoRZ/zA8alyb2yTQPC2Ui0T3FrYfh3iubBhi6YaCM
1BSj1IRP8ZDo1BQbPJCfwzGASF2JuvAr5el49iFmhXZ7ZOFzIHJwnMC6A7SBVfXfgzh8bX5a80Cf
qDZWOs6r/aOjJF22bObQcfTx+wHDU8aTn1mqU3Hw+6wwatcbEExQyuR3Ps8Qh0USbspbVQojb2At
xlRsvaeY3iYyKlMzBcTsVceg5eoEHK4oo0eBBSYEmEXaHY3QtWnqLkLDVUwoe0fiakp7U4Rn0vBT
MIJSEoj7Wa5cH8H5Sl7XxjkBZcAlWoi6xsqz8Fiwa3SLS92tiQ2n0xSP4yt13528KiT/gWYreePS
jcJdWcgb1fHYjXC5tuObvxmQ79/hL+VyG3/ETNNDcIUAwkijrZYZMfNbncVeV8FxGdX8vaQl+Xqm
iR1hcJJGKqj6J6aetKuK2P2M3egdw90XuujUfjHjocePJWrZuMjLUkAW7hV6Uu+g8ssG2LcXT/FB
j08JvjX9mnivTtZD0tB8GmsGYZ70rSolXe4S4nn/uuaMrWQT2zYQoFuFX2i03KxeNcKP/TkrU9eF
LdOSBvc2D0T5RnbA3YI82wAcyOTZbKDfl+JI6GR6NJJPvrboFgBzji4s3JVICIafGt1uRD/b0Jvk
WlF9djgtkV4KyUAZcY9Cosw2ZMvtUkzwbQpoVOpzJZAqPwdrH3WYfjWeOtgl40lej4b6K5cLYudo
A7unREy++rTgoIVz16CbnLZ46mQhjQGh7F+UuFDtAb0zlhZsOvwf0no0a+oQFSV9BVVM/8SNOeLC
US2K91jGp38y1IlE49f5TXySWoWuVQySpVyL7/iIj1t1fEWxNauWPPKcKmu2kSPUmK2/+ak/R4NS
Lb4eaKpPzWCI/KdeJpol8T1Nf+tXX7jB6bmSHyTm7DntV0an5GGbKWc7mFaPwt+IHxnlS2BYU5u8
2Mdgw55BsZftmf76nZugvHMs/vAuEXmtdobpkrKQ/4C2d6WYFueko0UUPQSxmB4jdi0c5+TSDhjy
0UW/nUn5EDkZz1xKSngWpfEobq88Ip54QYOIknx7k/zcaM/iSEEY2r3ATcAMHRhXfPzBpWOS0arU
IZDeqC+AUKp67c96TA3wIP7ejrpq7jl1o5cMVg4Tfg52DBSyBN1zlbBFn6Qh/ZX/bnAZlH/FUkb4
9T80kewBVtvMKRje6ZM90rVJJWuSQx8IRZtD/1lONmzqJTOiWXp/gHz3iUaWikkFr64+Q5Z8nq75
ZKGMKqEHWgCBJQ0qyQ86oFK8U94HwDZgc7C0NNMTOSfBP5nDRVCAwJviZcxQpps9yECfyeIbdoiv
nRb6Qyyhb0CRyyL5NPo4DzLE9B/tN7ONouKVgMpvdmLebE8TF9j39eC21pgl8Y4PSBUlLndQg4QO
p5+q3xqeu0zP3mcz/GfdJlFUXZAadhQ/oOcAJyvsYfDTilyh8U8C1fqmF/geNo62B8pyhBzmKjvQ
9RnvapGx3MXrzhm3mZSEtq46MDa1D0ZY7Mj/83KJsXDB7ZypzKy+RNqC1pG/7GuRugpOyetNcc2W
sjRAeQH1TD9LR2sVluoMifh09HqRaFgeR1La4MVIvwEMujTnotjQjzPy1JNzFv60wlQhWNg+iKx4
Jz2tOgTlmMYyrQqYU1YP7u8jyGJuYkaB1shnzA5wVINRdJrS5QsYVysuc1iL4zgfVaj3Q+3Zw3eH
aXNNIMQx9pX9X2ucCQRxowBLGooKuRFJ6sA61LutwXGJzKOgeiPuG7wWki02qqZs8oGYyCs6Vodl
HhbUpCpdgpyLJ6DGBeEgDiwgf5+CvN+uVQOwf+eq+JYc3bpwcKBjJF8J//d5sRwjms7Kf5TzDzmw
zcxvSD0xuT9BudwZT9IqsQ9SrVKkQY38x6KuYtvYKf2uyHj9eGQ+p4PjpYkMolhrr9sUgJlJk2pP
wZwS/HpXILR16qM3bBZp4MBT0oWOCcBqcwDQpFmipkT1YhFnm6E2hW9I65wLhMydw+d1891yq/Cs
MRvialeuy+9XhHnSW80QazfCI6wsiLwKxpe5/aVZf9TOHjYUKvhKSu25wjYG32YdcUI7EPtY5fq1
NHSC+anR53pVKxJ+moymqEf+RPrWLteyUNDz4kB9ue9/PrjD0Isb3SZAmnL1xmWh7ACxJiakU7P7
IfVlE/YS8QmQucmO50Ws/CDBLr0LZM6+np7i3CDsmTkUpyZ/8QOVVZXQBLw21sJt4o+qo4lEJoVP
ZGqVsjKVtVGjhopm7HS/NrEzYs8wftVOhwcypGZeZfZrIg/F5sWGnybhU8KtGjOXOJTjCC5ZhKez
OXOOdRhuTAzm0aU2W9sLQpb8tH5CU9PRuEDRIReWsuiW3TeuCkom88vrZnqrswD0ZVq6e0dHSpon
HKOimmnAzYdssv2e0XUGk3dtrp2aBRHZaAYz+xT56Kob2X0P26cWLDC6kkD77wkLiDkqj+Jw1Tsd
pFX3kZmy3a+pJJLNI1kSp0efZIux2ceLfyhNCpO0F3NHBAbcdmLseM6ZxXMGjTCHKI987g0n/uzN
N0I5aCkjwSFBoOf/3WkGubpIDGf7FNdsNi87lT3orQdReEvk/25YDXELcMYEHh1r/rUZ7SWlnW4c
eDYHXSuiMQeewEiA62eKYuv/RtdRrcoJkYKIXnTxTiDPmVKZp+9KFY7qGzNESwG0dkvexaIkepA+
QOve37Vx1L0/Cv8J0qGtJp0FhVLJD+3Hcq8mngsBocAvLqwbHtoGSMqUDB5KB/hVuAUU1bdMZtEj
SQN89xeF67kkiaEa9dMX4rcbdLhrXZrA+RaFDgSm5POM8SN9D5NWU2ugekVIVLOVeFJnjL8h3e6f
Zfs9nWkC/mFi+ErAP8p+GinZ548PuK/bGSGJ87w+FiNuBXVdqIJX0WmQ1dinEMYTYW4E7JBJvpmS
EoD5qX2OT35M3/M2vrkhAAEivWP0Duacq2LesS5cQxAlTfMG2uLEZ6e3k83JNESOBJKdcWaTMHpM
kRwyyhmtyFr5wvrGp8aN98kYFGY5JE4QQNJQhKiZQyaqo8RTFo4eso0gP/im0jyORMzNlhnWM+4k
rD0IheYWUdJb8Dr7ycCL8GMnbxMoh4UQ9vyISa+k2HX7CGFy8wnG0ohSwKRcB4j+yCMkb/OgnH36
YJeiuY4rOsQWDk5eU87aSXFDwybJhtpeco1nQ3yGwachaDVg1VxTbIRvB7iFOY0PGyRJBL7gKN6I
44+TsvTzq1mfD7VyFDMNf4ZpXk0WvTF5LjuwWEWORrWr1FO9L5H+2sG3sAAbK25AwNogfk8Nwsv4
kNLlaiR1Zx4wK0xWW2XUoEMh98yqwUQ7O2VHclZBPC0VzoAl0hq0H9Tpe3xJHobrZ1OrNmQKyHPp
mvlA90hY0B6thMCgMsFMZEvJF4hbUgXv/LfXia5ZFG7/SBFsaT972s80XrqfoKFgIP31O/A3xVxJ
K0V9+yjDJxMk3rMMOPnHPNgveSGG7RNgbNFXS2elb/4nSid3B3G6Vte0c2xHLrLDIMqIsMKSGMpq
hOHwHR2PknZqGU5mDQbNmnBel/zmTS8R7eP2lgpuOqeLqAMpN/3MYM7ZsRzeF6jsVksuW3/ornQn
FRU1uAiNlQP5FGeV992jmO48cJQ5GSK1aDHf853qZ0ba0v/Bqf1xJpFC/HrYuBY1G+iA1VC+O7zJ
u1MduHogY4qf5w9avKXS+0OyjzaYLP56jHxNOtEWr+B4ooXgJQSklZcbpA962u/1LfSaRURm/+mb
RywJ7f006MwuAQaBJ0Czz55RsD1Cz7TYRAtyATtj4aOWEdp52tUavekLU2AHOZMYjQ4Yr1g3p/dU
tULD5fvj3UMEWCSE3o+bxSOs3zyVkMBH50ir9eL7mVj2QnJIDP/cFaHPGjH08f/9YlikkAudX5rp
bccRhB2d/EAbgQMFbcVpd1g69zOG67G3cLRd4Fm/DayU5E3Vy3qm5PrI96qpPPEkPWCku0GLDJXF
NJhdmgdDVF1bhaOBX2AVrI6NYk6ffp0vNvgAufNuJbN8oPMi/2tAOtflptZoND9HmzzO82mnu/H7
vIiRDHbaPQ+g+FWOn4nWlJkNIqxrEclU4R7gUkRYPZGOwN/4ToaUjfORav61FaqfSLaZDuc7ijq8
kSSYZviaGH0an6bI1FSDFne9tFqfTLh7p6D9gHFHezOll6uakZFJ8qsBtqKnVv6G91gt6Sco3RIO
vWu2GjbSKh/up9oyzw4p7GQhhjvAXvGGgnd10m38cd+Z8c7bwqyngQfyomcmhiPJVyJPwBcHSLce
eORguZGXsFpCST3mWZ/Y5B6k9aISnpvhN4GmfZywcLCIicQ0jIV8lEFdESf68zEuG5QAZYx0BNJT
ynVzxeZlMW+kz+f21g7JJa7Aa8ODev2TUonhGQOE0IeAfbBkF8BFDJTMCSvQ5us59KHzLvos953Q
R4NZBbuspu4+kH6zMxLSX7EgrctRD6fKPPzPLiupaAf43NPPxvtQTuE3M6Tj2kxEZs7MNxqPytt0
0mS4ec5gCIfMy2LkOfO+ujWX3axiMAPKCCzgmOW/o8JFm7olokXsIri7HcIWYnVWVBcC84SRnY92
UX4lX5QSxNt+y8p8acTaWQEJLCMSJF7R3RUd6yP8oLAZVon8GM7AuF0LPgPXSVMMdOJ/h2uWYrN1
2SBMpv3CT42y4aRu8jg/u6P6kkrzACmWK5rzRN+y0ysyNZkWLqJwri5+AGwce3BV5BVbs0EPkqw1
L617zN+OBdcaO81HB1Q9hT6iJR1tsnsc/13NfZii3gxUUn43IlyJZ5e6x9/dqaxsRpVt5HUvw3Id
zp7HCL94+WkHxHN+PxlsNuuYi95SwhKu8gBV4YxG/s6PJkW1kSMfLpvArgPE0nF64L1Y9mT5ihqh
YFaawcKKOsEaz/MLGjTLrZY42DkObZqxnhjq4Nqi8kMdZAGotMafCMyMcpp7TrT00T/dQnMddwpm
eOrmgpbcvQ6ZDGBc7q1oQdzGWB6tt/Pyjpecov6lu2pC9fbN4PpNVGUmNWn+KwA2ju6ehPpnB6kh
iiqGVElezaqM+JP8qUEzmqO/20eNmjm5yZybeBHkvtUd9LESktQt5/1qz7iu/GYywGuRdR4uh8IB
rU1sw1CPMShpcRkyzhGU/hj9iXuBrvoJceGTUoyQpeQ6uP2vG3RW6bmMGMOQdcTzJ/hhEgCj2bLP
8mBuhu455ZvMEpjOdKU4NCPi6/Q4OlBKYT3k6CnWxlKqfspDoLIpA1hWsYa6PFDk0IAT9ums2hps
AcaUcLnJW5pIh8UJTNav3kE6QSpgR6QBpujnWAJ7dM54+PwM/UgW4obYrQxAsX89NPaKzCpP/H/h
VL+l6+roOZXt+1blpKB2qkj3ByyP1IrS2e7nZYzwqpfT/qW0mXJRSddLktfob6IOa7RdU5i50D1C
jY/ptbayGko6b7rZLahZWjF4MRDpxig6cHnas5+gaE3F64uczPHQlf4oYvjtsY6cqQhtpSsMShAH
gTGVuHGLCUMNPDNs1ACxazCgPDLDy28naWu31mdfUhPT+wSijdPsHLRqzLlrolt2CrIx9YT9VxFp
PoVUupKrQ/gdahqYMLPRH78WaCIPqGIfL/nhYKz4YajnLh7GX4AvTr6WuTLpKuZePrU9xWvXVmOO
ofN3bWhJZjjH+nHKF6T9ohcPJG18SUkonRjkI6TXRf18W5rd7K1tZ+mumFAeDG7INJoH7rYIMmIn
a2xTCrFyl1a38vZRMFxl1GTHcKpyoLk4cY6y7hUqSztkVOs4cT8z79B+mmrPrUW6LvUBGqK3NkV7
zVzPOzAphmNvQh3j/jcL23Qz1C5cmCPNQXPdf5L1kVhu532MWw9nJcsygO0F4AugWtFI+LrSqo3t
bhC8ypwmWqhmFTqETkmcRCcFemk+GqAE2DXbVyGtSaBTIn7eL3b/xudmGM/+eFUCrQDbMQRSPzne
ATOm85TmI45m4ePD0RutYyf/enP+xaqzpfs8mQuShf5dlTw5iK1Ht/nK2EtmgMZ4iDriuMJYk7EC
4jKE1JSRMPvB9BJOYr774+mJdCvt+va3l5kpjT9gx8tndkaTS30+qIMU3wkLHSq9TlT4hVH7o1LU
RyXQtvtfbr3o3hWV4WcYwFMULSQuyE7oH8WKyY3lo4Uu0wIQGaAZFoSuy9i24968sqAGUcC8bttc
+z2hXE4B8KVg9vov8z/KC9oPUk5kACV7JLxDHAfOByWU+QPo6fkidsZJMhv3rxgjk5v6YebieNIp
Gkm0jWdZxfFV781Uif5qSUh8PqH0F3vrOP/xNTsRErrAecTPVLPnxhYVJtfyUjpTunNxztjZbILi
mJpq9VTboU4ael3LSWx5jhmid9kKFZLYNXsSBaePmESgYvEKQBUMhEra5E3EndDcM7hxqORrfIKc
O8HdQ2dCWZ0xFULiDCeM/ksF/u/d0N1sZufmXULGXwI/WYVx7/C7HeTkLVqLUvbCb/jWF6XV/O5r
qsWIvNwFxIxsXprA5e0mMh1KOAtKrzwZD6tXYDAZjwvPyp9xhUp4w58xtoCvCpjdDgzhUT9FIJPE
GRFD1NLMP825d3lAATAwPucfAD1ks9r+/2ZBfJB+LwWUiwWOiszZ6b9pCqybw1bxVvaLmfLId7UK
CQcmNkkdO2IDnOTb/lkbqa7AkW/W/tr5cp8knpCOY9K3Qb0bmidyPk+ZqPDA/RDX5TBHqVBfp2Xa
FpaumuSpYA5pC+LppvL3JO6asQ+/CnboEJmRH/2RwLK065tsfe37SvHUKu44G9UgDl9L46xUdNgP
DbfI3Eo7Y/A1lSS1pehO+T2e4AxD73PloW9Tn9PEhhu2d5gz+LkVczSOmieMsQhIz4ilmtvD7VV4
678mfT4Kt8dqcXsEanm5tX03PcU/LOtcrCGizhzJ3LnqXBvtJucVAVUhpKIAIyX24GLt3TJ/26Co
sLGXLVv10tPK0cB9aGVP4a4UihSQm5o6AQjtaZljn25FiEACSxoOYLdCP7YS7Bw6qAzW7s5rz47t
s7aRW7GtCj0yJsXLvLOhhO6/dN/HorE5ae08TuS5EGb5O68mThY4P/+LQq3SQFuXkPbRyKj2c5iQ
w4tYsncLBpxdE3AV6XmKCR8kKrPbpe7By8pg/L7TTYpdZpK4d2dsPM5eKJBHHWkcSE4fOaT8gb7p
4j8R+sasJ0X6okKgigH3+TDHA/NsX/iU5wEqV3pZe3qZYLJwQDM4EL3aX1HK8az4EpBVqcG3N4Fl
UGeI2pP28SQ1kUnxQXG/5qPBJyjAHlN047eW63gRQvcNfwzjGqRr37adDQe7/h2Ffizvjp0190mP
qrQCv+biYUJDuDLQLcgr8Rv5CAW76TYzW9a2ygD9c2vHMKOZn92R050VFMPu+BQAJgP34bgWyJPh
SUWRdbZqz77EBLwAOzn+cOBOcym8fco+fMtU7JfSXBAzW67vwh3KZ8uGCX90mD+EOI+Kbc27rbZG
y4gE91sFYDVRgioLQiaFxZx3xlgKDJPcd896z24E/6WetoJyYn466sHXtRh7mZJsVMZDeb3+oJ2L
6oLA5+T/UV62XFyLzCVvq2KmDxUMN9C8LhwBl/qRMGRlyVT6M2MXxBVdNPBI2655htsh8rU4ZSVU
2RgIKoPFrt6iNigoYM4lYTVaj4F4JJYq2hlnB3LWWXTrXTum1DhxsZymJd7p9exEunngqUd+lOq9
tYDthMd3T7kkWLIwy1mGZaQT28KnfoRqs/Az30fmaAyNkN6v+OV4/A5+mXOYMNfUQg7LJ13AjvuB
ocGZfRP5HeDM8afsaQZpocucsyDpn4NE/l/y6VGJ5BBY7j9ksuzGnmLxm2WmbX+oxi2ncmPL4XeU
IIuTQSV7gkLR6ZShTwv6Mr12NvkAml6j2AVUySm5tvUaiT+KYObdvUZbYDi3pSGC3Sg/Eklo6g1r
gmaDktIRD2BT8oFkUCX/7RDmgc+KZvjadFTfgOXzOhtQZ2fUDfCKV3iYTxTjI00VUxhVun8XMGuG
se4YdhG40T88FbBGobslZ4YJRIz6NYDkqpLjtgJ+sSToZf/xQ7ldXslL7JVbqpwCkihw0sNf1MCH
miFHXWhmnvUaCV7F/PvCy3HBF578J9v6/k0Pms1H16yEgtaQsiDAEyfSzvAvuZWDOZGorqldvW+Y
EkkHjcCpvzQKuA25h+EhuvvOi4ArXRUjd5f/DaqTK9YnnXS5aEh50psf1QB9V0/KVHAp1StPmy54
Q9ZVaGMelR0+qt6exPrHX574vJuTzK8bhz8Wa+zH3jYYAY+91byNNlRnFRvSzEA8xvSvCOxrORWB
D+X7taG40wDVkycMDZcELWHRJJn4tLf98lJoFtJ/5jIiTkB5IBHL4ilTeBURIl1m15PCRbv/ZELp
rLu13S5bJKgbSYwqHNb7/gYIM0dhwI1fBArgPaeEd4+wbOsg6xNUZ83QUTKdvGEJ1hqQar64wLku
rI0/h6BrVd8rTVZSJMXNdvpMO7fPaC1IQ3nsbEBvPIU+fTXpKiaEMbHL7VABg0A5XzAwJTpzz0pE
V2SjjM+adtfkI9EOwaFZjipE5umE7VEbcNnEch8vxkFwg8ErUkRlzRxmmQr6odBw3axncUssKZJG
yQZxE8O3n9YaumFimKKrSpsd/aE3/VmjGrkhTuaCp+aNusPrpd3g6l/jXQ2ljh4giLCaLP9+24oP
Py2ua3SCypxvSvCDeK6Els63slNf2J1iZX/lU2wyEHqVxHYUnR+vrzZHD4AE3D/ajDUspKtdOLZ4
KLpSXVsU60i376zlBjnGnAcrFLPSo4+ITpP0qqm6E9kNif/1g2My/yNaN2od0fGJhKCgnzq3XG5U
PhZcQ19faG6fi7QPg4IbKRO1o4HKGx8yQznWgO3MPBvIaz7dXzCsvTBaKKCG4yW4cS41H+luleeD
QIRVrx3qXezwg/BAuovcLsGkKqkUOmzCVACfyKmVYO6K2XU/2XGfo7EtcY8mxrzHWX4ontpoXG+J
+rdIQPZcpFvR4JmbpY+LNWHK+PFZnxsPqVFzzYLK5LXXwyWeunHg0PlMOcIeb1kLwMf3y6eAEaXc
9l2wfYxkaR7c/ufoOgTcik7RjHp31v48vW/1GZqr3SD7TWzHMQUYRVXQIrjGHtEZIbg0xdQ3InPy
IrJmHjd2anPGP6LZtfSMEugXXjQUWQJdKyry6nQsoUHcSpEyhP0Z3wgBbzBAtfXtPER4gX7nMXGQ
wgCsENGbMaDdy0BeNjZ6FA/TW+gB0Zf7vdRLMewC3SfeLfuqug/FNxYD6iKFz+a/g95JHq62qK7d
wro0kbluUWZdxeruic8bFae4I1U6YOwJp21iLmy6W829xrRz2kTJvPahTxd9+uKx3JtHV8fpqWbI
8QfFH3WWtXbrvILqkosNagD+VuGryvViC/CEX6FvqNNcAPn4kaET/ZxUU+vGlJAAHQb1MSFi0ufu
Bc3ZMo3UWutpibKYc6NKCm75zjnhzuMgbdJ5opdt5RGWmgEyaDaEPLozhNV2pofQ3HDdBvvsEr52
tMX7CMImbfKiMTdZWV39nd/R1lwhK20fB6aEdSYk0fLjTZQ2kC6OumAMNRBkgR3QUP2jGyF9Rwab
HkhDTQvCVI6wVhwryZl2LTqV8R3e6dKSig7TDloofRHC4/OANw/EWMkrKXFrNxvwPS1soLEyjMHP
Jy36oEepsWmXB+We/rmqZgAYxAfM9O7FKhN1giIhAETpwVeM1P26NFtLYmfGPiOVvd0kvYexJL2i
iWMBA6oEEIG6PImUJwoVvrMdDadc2B7H1xbIYG6BwJVYPukyfm0fEbRX3Wp+UG9eSFpSi+7Wh4gF
CJi3qf7k0Jv1E0ZiBZXJky9E7iAtxkaukRRCcRlUPoSef2Li1ok33u23/14UjwVX2tQvOzwVZnI4
uPuk6Mfh0J9+Ssm3PZT51jfdAA+DJ+zFX3wLIjqRiFECJppLhRWWbZfRAlvyGnqZhZRy0qkM16wg
DoKyGGYdNZdHVWUSPcxqtZ4QoME69g/Yr9+rcnzT/m0WyfnrQj0WRnB7HPyd7PgA0eMYWi6PRL3r
Wpc4QrygQyAbJEnVinjcQTcly8nVYEbjMFNnNm4qt0dTtHcC7ZXmg1HGdtIyFdTTPfhlMDJxrNzT
1ztmSYb6wl62dShIYd0vpFIHHgHIw8skb7eWCkszKVp0r/1XL1xul249oTSJKtyn8HonLoaPZkdQ
kS2xkqUcgU+wOHbkgrOuZHqJ/IWGG5xMx9siLQaw8MC15jXpm9O+Hzq+csCazOPyrE1BkOpuWfhD
oDnGGxwVysPDNFhDNs3eT1P2Ah9rWoAmQheAPzUL8OzO1wSYD5+SO8cGM/l+BWSnPSzBTooGVQPs
Ugh+CEJhnois0y2xeB+41ojtI8MkVSbN3qZtae+3/eC7ID+1SUg2cMNGz4ftz2uhDID7eiVjjGtl
KSt7VnuL6GKIkhVwj6uDM4hP0h/0rnLuNzSSp2uE0NpIPWoVzvp69BVcxmtSrIBXRpq8Rk69XzPS
fAiG5rxVG2bO5eZjlxL8iayPko0YskUuXOGDIOocA+iJx1vuaah8aJjtN2QUjoOfH5N4bQ+ZYQwP
T+l7ttJlAQzwcw6YQqwdWYX6Fx0+llOd7zuTWSliVqJtEQEDtMg+wW1gOo2onTxarpc41taxGgPF
j1RE0u9U7tdCgHwAxPbIomb5FLBEmrSqOUKKA5XtLusncydeDKI2XxdR+yZvQ2yhEKXOSeBitpqe
Mss0gHtAlaw2ZefrDDh5J17Xr0VaKHDRqoUtoJbANke2OSJu+Nv4GSa2T2svp6cTQI1s3KtmIgBS
sXHEm/xYgsPPB2oEJkhSQVqXrJR752T1LN6Th4K/oNlkvJRCxpR6qfFBjWMoZZ6dp+7wVjaV7qV3
/N/qxbXsCZLvSzErXhKz69Gz7sRgExuW7fhITOWwqVWGBG4e39dXe3GSOPTFvhagfn5KzjvvDx2+
jR/e01so6YVgnqBoPJzBCkUWCaBV2kxBMvVJAUNulJyJOa+0kFUKVkgdy5HAoSQGpHF1lLb27R2d
eHNTVofPs01KB0QHDd5Ub3UsP2ZyFhINYgKWw6VrORetwnIE2tOcjZsfIOqOqdo5D7H00/R12DLH
zKA/Ged9Iy7aXXdC+8oKaq08ESdaRbSK50JTRRqxvKv+tFs+UNUR/stYZL6/qJ+rdjfosQbcO/Bu
Jy2sGiv87SHsUqsBu66IjUeCm4gbK4MnWKl5lShZ94MzKVd7hIlOw/tS+5A+d1W5KCNekHZTsZLZ
pAyUetZPJCkijV71di1v/CGFGm6Vz7rF5T/qAENEjxGmg/0fSureq8Cfq3YVb6zH1JC5wMr1Mq6P
UCDMAwPBZ/R9Y24SSQkCOeyTY/wNrA4UAR8c3pi6gZnWHLdSm8Rp/toXXnEXd94kajTQVMZpWuFF
+blJYMqrpoQMKSQmbgkrPAd7uwfdnOYoPugk7NhDjP7fZiV4CHkcBa+9pRVIaokoRY81cM/K9YUH
X8JnqFub7DyBjdhFwLY8wq+mnZN0C/PU5UtJynSrad8i39TLnSTe3b7r46mni28M0mWeiY1xqPzn
K7Vjtx6g7mc6DRhp2z1da2Ya+2Z5dhkWkjiwMHF3T/fd0cKZwNpjm8opSNxQBz30KqmjUwNYY8uU
ikPvYfWpYQhNYJuPkdu1d6RnEsIc90UwQysouun6YwCOTbKyS1MaS2gPW4lnvd9cLPfAXvYc8A8M
PNBcKhQOw8Wanuzp5KRIoTqQU4GYoiur4sL8tlON/057W1kmGphj+36+KzTCdZYPZ951HdQUgs7O
hRCuJkP3fT+mksBdZTPjOObvxBbiHtat3E99QWiyMA1UZKnW8TZc9eho+2ETd/Ya5hBK9DtzZQ88
LSWAgWgEP4KUcQhAHf2kj79ViIfW7ajd1FFpnNB1KkWBdshbhGSwnorOpQ48SDf9R6Vof2G6YRSS
7pGSRi4Gy/X0M7Wn8SQqm3PvkyceR2lZpHyvs3dlxxdMAwBLQz2yqxVaczUHrfdgGSjsjTvy+iYH
ElacoFbCgZ8hHK4XJJxkxGJFG2/Bzz/s7wz4z6xvX/iGDI1iyWABAAG95IT3knBG10JcC8J+tlRy
P+sOpU3OKfBbxD83j3wfcs0yp5gN97nUUMi2oY13cPkTwbjzFsv+l6PGIEtdxgttVF9agwklftsC
sVWjo1lR9O5AawknNISlh7hBSt7dnzqAbADMqZFcZuY4mIrMvJ8e6BWOE2WqmYO/3lZt2PeUTKx5
fwFHYWmuqreQ/DAic92qeV/PgrwqRXU6qIJwrpVew/zddEKx/tHdBZHV15TkwIZsxZ9qJwUerRQQ
cSWZ2qWJDzi3IaBGseWY6jYdlxiE5tCmLlV0hcVzcT6yV8vCdp/71Y9qmnP8jrObsROXNXQtioS8
hN9PR4wzM7aD6VMmcbgtIcACiMnHx8zrC4BbfxhUDnR7yL8hLiuJsAJwptwYgssDy2s/+NJ+vAvv
C4PPCp1e9bq1FoF3ec9biLp7szz0zP/A+a8kXy86I5+8nfj84LRWslrWEJABFqBFwbV+6fuqZwLj
wdvMPQM3X53Vkbr5TBU84TEUMSWsdAzeUQI5xr8kbvePPjlmcjvLELFX67p8sKWX0QkwKpZ1ddqg
eS8XScvmZtS1oYzgfVz1tbfhMTepi2EVgbaaBF2nLowhioSqIcvbkibBe7Uy5WnvODAl2L7Cv1lq
4vqwo/rQ2VC3eZUT/lfUhKNvkE6eaD8oUJHzEEBfcWjx8a4ql+Otkq6TUFoTrGHQ6arA/LUA0DnT
FW+/qIZX++f8CM2daI1RHvAszGwlU7UJXdfRR2ITYRx4JNbli6RmhxXjHZQz0DwdhOBPdA2YRMtx
AP/8XZuWuOoOmH+xD1h5Fiep1RqOIOLkeJhpKbjhM/SpCYQ90yS3zrvrv8IaBMQ8Fe9l+20vw6U+
h7KgD5TGKkNjUmxU6k4gwnvBv9jvak4KexBNsNonAuxeuo1QazKPDWmLPCgbnjMuMFJIcgINhVRK
pOQQ0qEZIdLVUgBNCvCZQLs7OMlhR0Oyzx2us/xo9/FSDurotax2pI+UApWC6EfDxkjQb5JETyCc
GF1YV75rYrCEakugRd9bS4tuzaJrZJEo13fpUbdUsQ+kler4UGb31NG4UR1t+4fy+SUoPvNeP8j7
3QEoV8RVLVZc83rreYcTPCoTBHCuYQXZHz3Ny/1Y7ryt5NkhJkyNJ6qhJmzFF6CSmLMxbdi7JvjQ
o3WC++dkXnUTNmp3wxMJl98y4eB/dODFzCQ5VnXlgPpExLcnOJdzz2jt3oH/QlhG2lRS9fYrrWQO
fLDYRQhl88qyRkv5YJ2sGk8BGv9eyNjKnSctVmpoVk+CR3LlPMbEU3UTAuorFkdGPY09BihmEL0H
+0pcI3UxrAYAjGa3KkaMqyFjtCpMQDZDABL6PuyvD832YPNlNe0ubc2eKaQITqcF6sDf8SvD0T7D
b0Hof9LAw22NXPqSHDo/CULT05mL8DgxD1aJ1zi6Q9DCFV8pC5fLSBHlUG3XoVT5JEdXM1BNA15g
DqLoZdhu9/T1gj4RKj+DjMzJ3bW8pjDCFfQyL2jc8Rv9a9cgFLkLigo8NkQzOK1QPysdljCv8zAA
976x6lBOFFJxM9XJSRKlSHnFawkxlkdKScQ9WCTBK7v0a13APg/6oxCPslwTKwdZ5iL2wxWvYx/+
w1DPZ2/Q21eJyLTmLccducOO4F5o4biMK95jbvVYlj26k+tbBaB/k47VRBXe0pUDJ/3VbhDRfiJG
KIX5MsW2V4egmT3OoB9vwYQdUhSKGJfZHqYW2+ukA6SvrWhov8ElMSizG762KD59wwpEhi6Vy3a2
NwECb1G5udvi8XHu3wdA/712qO56uFlUCsOFvcoZHsD7+FvdUr9pnvvBVmXor0tc4acAuD7R9/zW
KYEdYG98D0K4PykdJWv3NnSzxpwXf+PMhyti05MRPwkNAXXYG3Mu+Hyo4kaptcAErgIzyK+l/1BP
CdnATozUNfdgBt+AP3Bvn1XudoIUezFa/tO0nIb2ZHysdjJcEAQrNPK75Dryy5WvEIbiaz5JhjtX
EBu+gr/dJhmitN5rA6/E5lTdSRxW7+m8QW3ofQOBrZtZat1n3hm56okIDB8TyUvcOeD1YcXCTD/L
AUERiuy0/wyNnVrFJwpYAimxH2ZwXuHfJHQxSrcQVaac+RaLDwBYOqI6WB+4fZYYngDV6jXlKorY
ujpmsf/xuEAPavnG7Ne4mRtUpHiihjs7RZ6LjdSCsnigUZFjlwGB07kkYaBdK5/EGB9hxPnOH77W
NOcanaiCzn6WUEudXpzlZE23ZRizPLG9t63bq9hACXNOvnz2kWLg55qtSfbTjIj3DGzb7SwoMpS8
6rZ+2SetcC3zTXVLS6a8FVTip7Rbi6L9t2pI9mt8AbG7Q2ScjINYM1ZtvWcZpmnB6g0ITEvtELfa
iCS5DbtxmLgbGCFxi5/bCg9qdKMKvB+WRlrMDvsxqco45mjKc3O25OhVw4C1cHthW5s7M5Ad6sUF
aG13u/mlwq1ZQIr+GVZ7dXvXo3eUerQ2ZOESfiMNGu2P04rLW/0EJV6HiiPP4qxmqQvWXC4mGvTb
sG/ry2qoON73ysH2amZapX2UzQ9HJ8/ysfWghe2ZcPP0r//+8LHxTBBVtY1qPukJpoazBJJVz7go
K4EHasbSCYfb+rCO5dgpW+U3wG4Wi5ePC+d4ANlHM2BqQjOhSYxvPYJwDW8hxgu9B0qRdPQ1WBqo
1zB9lk+pWe9khCxoiKtPK5S1VsQrbKjPWIf1LpWf0bdvDjMTjgfOKNnJ8JfCYSjfiojwKqZYwVQO
ozQJ5W9vmT2OHU+ABJiZoOFob0NNsyBs5b3MXElV0NHBhzFNLOQ5V4wv2y9bBoH6oazkK0lh2iUl
YVJZRo7KQdZ7WVIu8VE+R/4HyoG0z+mi84ZOW5rp1msCQGl4yhjNhvmsdroANC0Ox1Uv+dPHe1QD
zVlW5bwMA5O0UYJ14jWWjetU3dzk5y3GWHnOoTTH4KyVKnGPVVOTZc2rcV0MC/nfUKfWK4lCmLsw
pGzjjivAqCfHVQ9T6rK9IibVGIDRMjTMtmVYW8MyK81C05XY4xeOLUt/GKBzrvGGXTfBhDDPi9ot
U7rtQI+bgUJ5vSz0H5vNG7bsCyn6YMGBg3sXM/2z11QSA0LwqmeBOitQJZiMh1moQekwPLTBzLWj
3GNqu55AfeCr8/S2tzKsy356iTrG5ZgHxK9W2bC+hnioHnX0EtXaFTVNrol7mIGnTDTWrGy3Db7Y
a/F4G8OjU1Mn3RDjLKZjgm2Q8WEdjDOPGfaG1X6cwHVoBtJNN/F73qdD8qwFjzBesAgAeKOLHpPw
y5ylGXOXzKYh24DDHjT/D5VBwlgtBw9tUX/5t6AnEzP2NnSKeR65zvoPpAx0t48j4fuku74nRO2m
s1cFXV6qCG1NbGKtk+roWFeCIQLP83w2yXzbR9WdJsWehBWfv0n7OOyvHvZSX+qQDP1WUdStaOf/
amrtgzB7doXTKtfaitX1LOSq617/48kbPXKVoemRkgklOoYNJeXiZo+JmFyMPveoW4199gjaDue8
K08pA9fq3hIDOg5BCPSMkYaDVDTIll6iYwooRIW/c26KCeGPKNOh+lV+tfA37Y1Q3mD1wjJgSJeJ
kTyaCeAZqcw6dDSx8x4norvuKEHUtW7WpNohfF1j01zkT+VxublaWuPUXsXcjvDrmKkREJWos8+m
RenYr2o4ogiFB9WJdIqMW8jVK5sBQsDVB5wZXmJFO0xrQu1lzp1GQTpJS+n+3q8w7tnAreZ2ikhY
zUA1jFGoY8m74PIDowdCh0HXraPdcPfnEoV3bfKOhU/s6BPCY1Z6hPR0WjC98ouFDEiNhPQAMesm
TymQsYgKlI3EoNNdckSDsJ9AMpFnTq0gdymLSOt735Jiwl2M03wwAVf60XvrAO7e1l8JegLzEcgi
v/7tCTmX9j2Us/Vee3HPiME28XZh4DvciXcy7r2cgdr1aYNfUDeE35N4ur1GYhS44YLIHR5nQyRb
7y34nyTP0VgKlfO8GexxqKhWJuj/MkU11mYzZPEl36036b4wTRIszQdNVr/2ZHJukYoWrjq2SPeb
wo+BJSi+IY3By0CbobWHh+yp9VLF3708GEmvUE2CdQ2O6Mlomf9q7vlU0i2A54CTPtIGrX0CURSg
s4uozJsNEcVlKQvIT+b4G43PhWZ9vTGlBNKMJNgHNiVVKYe9IEoQlnSnMYYnTaZUKKr26vjsJdrP
pWuqKIT6M5jgffRrahLj86BElRgxv0zVprOMvdWc/NimKTV501PNZdCk25kkd8bjy2ZwL6hx3cdg
vle06sJ1/CIBL2IlBQpeJ2dP3/SwC5aL+ubb8yFIY3zbCZZEh6F7fPeB6W0Guf4GtqO3MUdgySlr
r/oUP0W+TCxpm1QtD5tQT7MpG8OgcWlU1c683g3tyPzzwJaFFgXRizDqoIQw06G7OmPVunulClCx
Ab6Nw11Xr1yYVMm9sM6ATJOaornQwBxmDRePekGOErsv3a9LHvxnNtNoTkDZzgOhUENu2GgWZbEn
wrCJYQIE+9vKZTMwB/gyQcrXdGPokLHWlHubYMG45oaUKrG5X7LRHxlPKPDdu279Uw9fiknRAHU4
NhkIgM5NwgBqTo+9y/29D8nwfsBC4EmGB/k9wrsWwfUfitNA0g6l+nhqKw5K83XX/vV0DLCMVguz
FeV4F//CfjBctiy+De+buEjkGzBXTsnqdi4YcRmX8UlytO5k24mbq+qjPTSseYqfBgv5m/g3DimB
p2TsGeXTrkVSxUdz8GOF/G92jL2DJaE/7Thcs+2Rluo8GtrHD6BHCzmIMr1KqR4YaYQ2CuogNKYS
vNS2ZvtFSyg6AnV/Pr3/M3xWfFqMyNc3/EKIA4Y0Zt04FFlj1q28CTsJ/5hJDldZYnqClPO0MH/k
WKRpuZRrmvtAaAa4k0GLO76BMWXIzm4qDaV7MipG75VMcA6N/Boop0sj+Oy8NC+rY9jFPGRdPagp
SMUIBcv//yP7qJeHqazEypHlTQtf16sdZq+IKZ+RZ3r/d2FohQF9jdULKD0LPsJ+wEjkvUQrb6X0
37afxbWTxgUoDGPvq47gNN7UaG65X042ig13swy0NBQRSVRZZZnchPTi/qtwJlTOQkLkorElepuK
JvznkMOqzKzm3F1mOooOV7jkXKF4xdxF7M3soUPj3eXe7H/lzS6GG1eMY0XXNnSWrgJkXgl6c1NN
swe6/p1IreDL8+3MmVX/c0Obpr1OrZQnXt9mGa+I6EUZkNi2fEfV4X7mYohTm1vtSKHbRmTKkD10
IzW5DL31GCcz3NzI4aMC884zC35QMlv/3a3tgmvmJAwjkXsR4z4QmUPFWUEca8WtEzvZu1v44H4m
6K8M6TBYAuDSPvEUPjc0RCk3uGb9mCQDn5LEL5HZrDtw80RnKc79+5NBQt8QNq98JbKVdPAC861u
R2OS3wkG78sO+gptG9aQOzoRdYwdloD+sd8BLgCINTOdd9BZZu8SkJL1S/ZTr16+qvawm5zMyDmH
YKnHzKSEyWVSjd7tLZNUlXBJkQv//j9/qQkuUVA6SMLQNaTCDtK/COY2qGwDcvQaM1WElHYAoTQT
fsT69HZBrB9VhRs29/rkpgNOD4iHByGF2upqYXuFQNH65vZGdnINFCb6frCXDz2cUNVQqeYvQzdz
bV9uNrdnQhY5xkMVNd1Uma6S0fNMab3VCC4XcrwVSfhEsZPn7sz98jS/7LtbrH2Mopo05EXy5TIf
AGDErR0bJodBvNy2QzFFBjSOkFbP5AAS8h8EhRvfp6ud3U19HOvu0U3fbXHrzFB18knFtxmM/ydy
C73wwQOH967ygk8F6NmnHcGCPcicg9dQu2J4+8HW4zwUi2xwn+/BA5AiCTy9DSSCRpo/nCvsD6qe
x1V+3SVSL6GXibWV9QxL4XtKYfxjcYHWweKLIA21RqFWBa0kcG/nUqJ4vI7Mg5OfGs/LMAtXBqOH
9QvEhrS1RJSZwiXSF5cDRxj86+6Z6B+zD3YVpDUxIGUR+C0GVnolUowQ9vsYhj+0Wlm0DaSR8k8T
YjzG8e+tt3ms9Io6h8mqg12XbhU3lcHkO0JETo9pAGXPI4nT194FkmofKx3sFdcbDy8bu2aNQXDS
xVfeT9I1zHZ30o8TF+0jOPY65uLeyxQM/WH01V/XzV4iFMGnawqT5TxcYpRMLO1VnW7XSYOl0aJo
ta9GLwup44CWA8BB1Jrc444gUZlZPfpJXSmseojXVTc4Y5XudFInY0T6ICKQCj7LQmtwlsMPAXw7
w4rJsVBL2P9YLV9Kbm8u1omTuaAUWqmEbI/45R42NDjVzLnCfmSwOG0odiPpbz5LFgxCMt2pNdVy
PwT76b2uH7hBV0+6Y8LL25k7Wm6HpThYXxHHZRSLNRaCyPFG+z9qaMXz0Z//Ug6D/HtAOcfXYrwr
Rd1d6V1fh01C2IR8NBivRUwhM5CBsMDSW07aCLKFO16pFY/+WsIoFsbB3wMvnokOJvzonnDthj3s
GwWuZ3n9XuaXqbu7zh1G4axHdRE+sPeN/Wh9r3tLEiO3NhvlhbbDSaXdzWQxccc1IBGeZin39KDQ
jCAhsiGZfh/FUjej1ZV8aTiL6okh7njMr6G8CsRxfX18XFk2UuuRoy+MZ3IDY10KlPFkHyC/36uw
8t1+YKWgb81IrQatlNFoW50f+HApFj5MRO9UQBBHNUcUOmLZHLFxzW7LxHm+SMlTBFwTqyN0rSGM
gFwhScxR+SUBLPAjk+haZa78gIUgobf397vVpLJWTZXD7BiSGjkcSeS1y50pxofY7SwQowLDGpem
HC5b7XHnPESNmeagXt094RfC2f1bgOn0fDvYaIaNHEiAKobQsYOPtyR0HiPAtuI/kwSnASq8nyEW
MraBXPYSiJssE2IJn0GirnJK+WMhvBdIXl1pfAByXLPmNPZRI9WWTgSyODp7l2hYu7taK9TGtAuY
h1GRjTBBbFXlV0HtNO3UnEcdu6y/Xd9dkjivse4vF8apSkypxWT7SX/7DSscj4RBRIwhC/d9GdCC
J39PdauTUPbsSzUaPQBuXr3EJlEfjaJVaqk+X+CTzi7sAepsBZ4ltSNn+CJZgajt0ZITVDQ0Uo2f
FrkzrE5qC2/747sLUb5PbUlDYMkpenxSDxyhd2Q46yqWTAvNIR0kiDAuV/beF3XRFgvGhD2elYip
+lylIBVZPTRMHLeT+MJecpydqeX42BefdlY8cOAtkEQLyHoZ8ouPcCYBv05D1S0yqYGtfD2GAbaB
Sb4tkMbs8RdyRbbGsfLBisYo+RXVy1ZGLopk90pg3F/u9xbSReKE7So6cSsnVsDfbKW70yTTEjL9
5wgsBmhWjOY7rghTeIwqFD8ZtpeGQnvsYcc/klusOY4bN8aq0IvkxTPbTMCE+gxdH0d/LxyddZAN
+xsewjvOaxboqhrerDu5L5w2+zoWwV7SsgFIFqaRtL75sgqUA+XHff5RtJyDL2uADqE5ZeuLABfX
8Fh/yJxNn8Uo/lJE/FdMtINY/oRX3BlSOoz6eD7tvQsSjNVR9/cudZrQalLuOJ/zvzNNa6Yw58L7
bPh1BTnGk0MX4zlowvdSqarDeH6VXvRMcWHh5fboG6YqqnF1gfFRGuMc7kmYTQzrteaxg4b+eCd2
gWKmacS7E22tYrjWzejDert7s0B8YFHXz8unMx1qUbDXrGjT8j7+O5ZI3rLLFOzEIrLh2iD+2vhJ
dWnRshh1qq5xrT3L6z5yDaFbW1Dp2o+fZtqEX2ZOnePGAwV9tElaCTj7/QtuvqBRa0omwfQKaeWD
AAuvBdjGP742G1G8hIzvO0DRUcg5l62BHwtAD+XieOq/0o9+HfMgYBTmVm/u4cn1bs1M6WWCJrjA
Ni7aTNCA24x94qJ+2Uk48lCWzSOGCaviL+vlTXnUjj14T6WbHTy8XWnZErM7WOX83foUVSRfSIiO
p2mvRF70C3t0agdf101UbEg3gc4/MTiWmnE0pOnKR3QQD3j97IOvL1T5yCaN9e9cj2Shl1GAKLEt
bwyZp8wVkZOxwPksMMJm4dC62PkybE58tNvtyRc5qiNMEmvpWsoYq6gtQ0hMWowLPrMktMbaI+BH
LNSo4n/ZDvevBswLj9uQzmCFzC+uFNMayS67cXuliuof5Smp6ElieIL4BlAtF5mN3Olr8emM+k91
9BqJ3/A4etfyjSyv6XP0V9X1dLx2nEjk7h1bpWSCxf5f0Paj4IQeZzCj/Z1xYKj9lYk6LMa8nj24
FXYQBXDwe15TIxTX+uyvLg1fxzJpuwbybSOG8ohZqYLx3D9h6l1Z7OC2pEy5ctRLtGYV0wFASDdC
XAwRtEkW9Te2XgioGvflMVw1jaW4CQoP3yn90Dgn3ZSuEl3aA3MZfgZEzDNMiIKZjuAI7lsun7dn
lrYG91JcwoyAC5CkGd3fjq+lYV9dxa4cAWJxFc5LPZGpfMtcqWE0PsnaHLnKV7cBZonfyg0bno/m
mrC5wXXdrFDlswx2wdO6OFOjLTIyc8uEEh9mBpRz/mrMsGdFaeCl8PM/AnLrwvoWjUtCpvkB4PEa
9jJ5aL+Je7ydoFbs8Iyf3mMUA4HtkCkdJtaXVpYl0m3WNoJamIQaeTrPQRAvo1Y15YUTr8lK8gIK
LPh5RJW5eCqqLlmrY6RHa9I7u/kDmFlaC59o8KnAcZyWlzbexiU0mhZD03+0ISF7OXjlLGq5yly3
JQo2eOao6xqG/PeD1njPuziXZRvEQT944ofZsES0s1tc2i+/72acR/har1BcQg1d4xYJbs4a/QVc
ovx1mQVBccPz22JV+OFmZtQRITiEFq/qhepMVUTgiiFEtY4mQCpjBG2clONfi3I3nV7CAN7rPjEP
Eo7H2Ur7vHNgVzUZ66VD2NtTS4h3vUxi5HbSPGnIFnc3ozzXOZlGlCXlElHezxlffafHuxEO+8lr
BeBBEPmSGQjtloSd+7Ull9ELvIC7L4Lxr6MztM5MsuhtI9l5fD4FZBAUH7QWYIVL0WyH4Y8zUi7K
zQPZkFkGHVbElgJeBLDhhn4jql9dJcajje3vYGhy0GYo4Zy0dgl7AoWhfmLKVy9Orm8RlxebadrJ
rIhqMqG4kM7EDCUwYD3o2N+rP52epnm7QIIMaDnE0Fz1c07q8IBsD87FO78YYYDwk+etgfeiuG6h
W0bhXXdFjoWOx97dafmm2DyQS5HCWQJ0dzyTy+sjBZlbudrzCc/evO/oZU6oa+sexgkAKDshnJtT
jcNNtTeJEvjRl6pdX1nWP3OJMXZY8+1E1k4z6CPEE8aIdAdp1XTtuYpMD/OrDIdLC4tR9Qp/nqMR
Zp6SIPuC5FZvc3Ae8bbMVuM9zmxzypmwayGK32mQit1S50sxqaRVo02yVeFIKz+W3NE/yNR99TiW
jaS3RKRx4OoQsq6NrOnu9CtS766cDiSeOvxUH/ETUeaRH7Ge1OQW/VjlrY37uIyl30ByDdRpQQSk
FRAahT/3Y65Jl/MAMuBx7ZBkkFqX7ycNPYTITp4/pubXKLpNBUVtpyjv1lXbqsziWsvF4E6/D1xb
QSIWrhKJ2YKJhGN5LNlvZzA7jgxndrxZy4LTitlBwKrC0dGU5o9j2uApGYy5zjA+YxTiPvU3v78U
U+lUfvlTJbM8ynja12aHMrrZM6oMCfZuQk/PrdGOIX7OYaVoSRA2pIujJW2J0EidX94wdkSXkocY
PuaoTYtCwlSoVKAKmywQ8swGn3QTCSPS86NXIFrnQCITApCeEuqNa1v6Rh8sWRcKjRD2YpWQaToi
wn6IPD8IlKSghcWIZkVsy+E++VHjAqlPJLNB8slkvKrA++Ztkv9pelkHmsZi/G3P3DKPCVBGA/YP
kC/cEN/wl4Kn3H2s7xeS8f2SLCtJadALQAk36ELdPfuv26lQlnWHqbt1P9gp9yUGZ1QNeyYdr3rh
n4HblrCn5yH0ZqKTlUei3uTgT7PRL18zGkrgXIVpuqhuAhmVIC3tzQo4llG4uaHJHm3qY9H3kYFZ
GwxecITb5Iz74acrKWLInGMfq3EH5PJoB/3Ji1gfOj/rXZj9Ulmv827aPXLJUeKrUa9e8kyDrzeT
nXJAYP48iVaKb68l638rOzhKdyqe7CGlniufw6zmM5wFFOT7Dxvyn8qv5SCZnw575acOQBWmoylc
8MvYZnN8+G76WMKcjujbLp++oo21Te6ycOrHHepeXnUlrbdnaaMfMAczwoyikfhqNiMPJ9TmfHYa
OIiD2KpdGR77XUPvcXzsm52EeK7KQtDwKk863daFlWoWnlMJrbT/XxB9AZmMvR/KucmLa7YuKvt7
E5Zh9TIjpdit6+KkseX1f4FD3lnkUAS88UunKeMPZpcHqEaMoNdozuYweQo8pbn/ukePwgdUkhpc
pplvTsIQAECdpYvmSLjOBe2FRKpakezXxttIjL3kpG9h6CcV+AhUQwSJhV7mJ0DiWCH2w3TwdQ3C
XJrbjZKIF4XYFjWs11KMGsly/ZxcDTaj3ug33ey0pTZc7uILnQ2qNPtfvSlbFs5GB8o64nWGrhME
yuLv1etXIRiMuehlTJgUTOs5GWp5Ac8syYFETYWMMu/pzmRkxN9oSXBduVHG7FNbxsFy1AEUrRJa
4rLklLTtci0Be8OMudcFIncx0NN58XDTQ5C3viUHP9bx+zK9jDuzbpFSvTjJ1+Yy9qPYJs/qude+
Krrk4PcDTKCcaQnPGxswjf7O9fMq+uEj0vcz2pZ3PdVJGz/uDK3VeodcgT7Cg87Zg0Wd4a23Bum3
XFjCsdUMG+PYFshCIaTRnZ1gECFRlFmU7E69AJHw7njpWv2Inc4aNe6jMW10JosLpe0vyDVmRHV1
GrZ3u8nbs5y1ZNMH6etpAakNr5NwdlInGEhBNChyrUSIEDmB2R+VljwCNIjLx3HbFmXgegtPb9sV
z5o2/Vu3bRGQgNs5/fsSImAeSrRH0ddZjV/Zv8Eqw6CGxk7kVbqy5UfIVVghHufbpW9XwCSMDVXv
TCpxqogRNFmaK0d6hHuKHSs45bBY0XXtU38ITs6FDSCVSuzI0cHIEx7IJD6aprobAKC3sNcDnROo
rwnLtih2HWJ//FXgzDgyDVq/aQjoXzxl6rPEoemSO+Pm491ZD1eoTTFNluVa+CovypUxRiQu8mWm
PGBLRGZ9me7i3CqYZw5FCKg63CPk04D7+GaEjtJPnBv04TuzJ47OMOC1qdAZm13rtPz4w6RHhugq
fyZg6utYszmbhE2/ejoiEhutCY6J11shtcvtMGwgnXqMJCyQzm8UlO3A+RafZXktcr8ZAWDftyv3
cbvos+QI9lp8uKDDNyllX2A7RpWlAfhoJavcLhRpOOJZWkznW1kCO+6HnFTT1ZaTOeDqLdWbP4O1
c1D5XFqvdcZEVk3ZwtamzH3aHdkU+4lSRs5AYp1L3J6qopMCVsbeYwrIn/LtJ/JLqAT7xrXNeNH2
iLpejVo+vyQgKk3mFmHuIQKLQ81hPA61k2jJf0YVE986jOe1FQIH32N4k8SQNCeutGi1yE7Vdn/Z
0EEKpqq6N/t5BgYrKKovQbyXZCX9J1uNBRnoJ3jY8KQFPBqrsCSWQ4m/+jG0xMesMKXRL1E9prTF
MSpx5SiaE+JXwEgNpozY9Hf0LDRwMQA6zT3gP8OsoK+Y+T8WqFmRHYR+YEhMGz9Otq1g2lzCuOVI
ZKOpPihN7y1ik4+G4fRHybnNu8bCQonqweV7OGFBqvsNkgA8U8/PF0YLFNnG7I5Y6kaH3E2sUyiy
X0CFW2IL2QmAs9VO/65geHN1cWfkzVpgKMrYYG2Os1HwENE+gwEsCYazD/IBufOpJwws/IiTdXFL
fSttKjy5g5ZFpKrgx5KGzdex6XXfJIVUiHkg5SmDrAd6kSrXh1G5tWvnTVOcl6cPZK+DrYqI36si
8Sph5YVYPgTQqcEvkuKd3NMhUWzpTw814LIJFNahAySUvsx9lBJL89AV+c9hJ9QYYszsoSyHN+OI
gry+qyVtjUL2Eff2YBNLewfT00mBWAsBzAWORhh0i5jGaqvfJhPgzD6/HRfCdagJAvtWz2S7Ic1q
G+sFBo73AYWZycNqQBYU7/ckdo6GnO/8L5lz3zpTck5F+6LgGT4nds0X2Y/klqcqp8Tg58VghuII
9OUp5MYFFuWR5rmJh2Mf29Y+9HkrDXH0qh29cLFta7s0ah5Ac9g+FmzNtjDOH0/uYYCHOf4U3OeB
kV7aEv3k+x3b7X0xXCqyUEXYyywVT5RgOao6rMQNsxE72BUm02s49K7NquwwZzwKXw2cVUN0FCi4
ZddDyTMA5zb6DlEHEL724CcLu/DLmBkTkL6drfp5YAvWQ1cbJZ3m+g5pC5JOxXvI+/OvBbJkD7um
BA7AhzuqeTvzkqp+jGmUxr6b7OwhCsAkj2kJynqBfGv/0LBj/0TlcPCN5WSsHhPtRAIkVC9enhm2
ZnDnCGFXrAXEbypDV6AdS4YaJI1dJaEcVzHXUI4YEGuFKFsTEV5+CaYNyTbnMnUTMuPe//LGBROD
7OEKdMmR58omu4ppeqmWZ/GH+621SksNOXR6Gw5B9OiVyTpHGUTKI4j2Y6t06tF+TFf+tVsFQWOF
w3Kh2kMpjgnJEYmdPq8dD5U5TQHFu7sAZ0m0D7ea8YTam8N4lwoLvKSXaJPBWuZQBLN4Y3lKCxYv
yZxx7fRy/lTujs557xadNh5922pPyD1onfavuQvTkj/5qe317NdnlCc35O6v2zuwOLsYpZWMyUgq
8pL7VTO0tooQKGnooBV1WtqsaesDFoP9d6uFH/yZ5vZpZMA8uqFxmMkInRxbRSMrs+2VjRwjJIgV
F6dEB6vUzh6Buzpu8ngiyoFUEtzmBtvqx3KPn8PfYQ1dRJdhlUCFAKclofjprvNU/bhG71Ms/9IZ
+TSauOuty4Mqvwq753SipgOnzkoVDIMpgkCBFr7fEwnO5ey0E9/JGUbx3jVPbHGIbzRRIThooMhq
momzUsSPFq3EAJe7t06qO5pdQ5fOv+0E68XB4isVBDbr/Tl103jDdTw3yB869o1HTHE3jvZ/8teR
/DSXnD70AxHq1hfNvjmLRG/t0EmfuXe5UVXHAkIQcMFB8zj89zuhDfE599v4RVM1KPUNC0hu7YRT
eRyiHr7w3hAzEur2x9/TwyGUt41c265cEe7feAFQwvpS56qnGKcf4d5k6Mbp/1BWC2nEt2ZwrqcD
3W/IXUzmQ889z7uqLqmaZ5R4V0eBJ/iPq1mjyFuYXxH8MCARspV7c3uTmNAVDrm/Gju8atmovE6S
anWZuG3pslgc/X7hSjbaeqwUrRu5dsSeHMrcAl5Panp0yKoaihC+x3gwbNPBB1fUPm+l3HmhWpvn
TDOvfnPF5istsJPRApIB24SbRDF4v7T4jxWP9fvzTT4Ysg+Sq5KXyqh3KVb81EcOaoWwl2mXSU2m
jBiLGKvDCCUdD0kgZxtjfLDTjYRRnQnTSOTJTHGecZVzTsfVIzlO2E+soW1OOtP9StW1xiEkg7Oz
eioG3soLq8m9cH92XSdOXUhh7eUSqvApAHWZKu76Pn0d8j3y8JXrbMIh5UcqJuyaaxB4w0Ie6Lu7
wW8DmpYpAJ6tuDmiewXyFXF+n5gN0pTWrKxG+LXk9TyTV1PBmuNwHfr0rNbz2TcERWytg39luWiP
STXz/lCHtRlLwVm6Q1F4RH8JT/nA64zTz24JEa+ODscxBPqDpU+CXDxBHYs0rnrvKvbiN6sMxeau
2T3e3X009eoLcjLBvjdRJhgIR2stWzLd8TG7EsbUBDk2dJRB9bzI1qpnlL/t6LaBJbw7Ya3rbuMl
ZJZ65PhCBTxx4G7tefgvKNDs/A0z3pZvALGv0l4MpVaewAqTBHoWLbomDC1gYcNeNLmA4LFf3oUt
tJih+/GqC7OWOag1Ge9y64vCJ511EO76aUbH11bdivRxLWXG54dKOYi/vUb+zcJw3yYVGxiKsSox
7sH5p2gslvykteXdB1XhIgNoUNeU7kr8JUz97pSvkF4/3oPyHBlqL3JPsPvZmwLHpx+10D4xv6F9
JZEGgpotRt5wVq68l2Kf2BWAp5XDqIGFA6+yGolA+zdX1Vy1PBMuKCrbzeAKHoYnd4K/1TApPEtL
cguyXVgvZRSAIR8n+mCU4nhPhDfQlhUgR22u3hfxW1ZcqyirDAUVaFw/rNIIM3LP07hLC8+F/XWo
9BvT5JF7sJoifJxYTlRzBKtlXU+7RUnmlcOZOC3ZCFF5vKOBhdCDqR70g8EAjeBG4fw15Ato5Mla
6FU96lmKCi8TC4RTujIj6Ip1ah5lcwJuX0cpjZuJYmyEJTmup9U3w7fGS9fYwl3MHxgEwk4j4l1p
1uUbvbzcRE3eHk69urZ1EI4J6bThEdpBi4FXd904l9FZOvgutCyoSuaax0HiqB2rCGpTB1H91ZrZ
/BC2s9aIUk8+CGVM6fuMpLzcuGmPoh/ZOfAu/4FULasN27IQ7K7IFXfAafupYQPgf/iP2wBDnbE6
UYJzUy7JeOYeSUeXuurvLXXkprmYnx5KpNZR0Gx7AkPfFqXGalpVOl6Qo7p1ogoTbPobVN7jfG7u
4eIvZGiP/5e3xLCrWm6y0vWp7+7tmgeRnp89WTRSWEWWBVw58gmoc9bzMEF7kdhSZWJbbR6Wahyx
ojWOwcpdN+4HjRdHV1xyGNUt0/YV7rIPBSPD8ylHllvwQqjH+ykXbnouPnDxc9o0p55Jwul5vs+S
E+es+lJzIW3H/yebxQ9hKW1srWo1gZmdaBMwWlNz/Qo0iL/dcXU8ACjYgJDo1URLw/va+8dlBhhn
GEev3WCNEK3l8zhVDEZANYxg/95M3UkCaMn1rWqNxNxb0mpRi02cT2fprQhow2UWFrmFR/bxVUJu
9e816gJYPtr+DrOsUEYzjiGRn+z/cR9Ss+BAESwsIuJts0OICGthgvHUqcMWQ88f6kgzMGgdsnDs
wtDLJY+O8i9uMH/GoCH/Uv+a9Bru1zm9rTXJIhiaez+0dISnhG+4ny3qBwpFu4/eFfCX9WkSzJTb
Qzyl2oKeG2PzfYFQngAT6v2NILjv2o5rO766UfELeKyLxnNBSnZjyGNlQSk2j1a5jNjRFJgqV/S+
tRPMfCW7+y3tJSCWSOlXcBpp5pNqiBJq8JlXDHlBGu3giosWjKNVPXpVRbZmaB3KX0y+mevybGAV
cLQtej5ApGLtSgC6lwvHQCzufmvJRkL0mMUN7C9LPDY3Sw7w1o1Rf0m3GO2q03UzCbZU1wR7Xyxj
ss6deJh2v0qTFxVBnqBRPDfucZh3EZHGT854Mfpov2Q7K/bA85xg0vN7WPBrd8IlufHnwsF89R9b
fbk7a7t5Kckinm7BZsnw2eADjVrFi5xYwmRMrAnynUpauqEDDeh/2DcinMPkX882sZOm+Kg5jHyp
d8qUJV2MLrjOA4hpzVSDV1Pdx+4SgbXU1eDXSP6ZUERipjs18lP3P+hwaITYXIjXnJgmc1+IWegB
kZm+f0pawacVxQWhF6eXQaA/a+1Q0uGn2PEh5xJydkt/eSTPt9CQmcnEi6J+hndk8iTFvzPLoMpf
R+ta6Sx52wEa97RGExjeqPDVvnyEcMUBQ6MT5bG8XbWLqQQ87i3R+de8f6aaX8D9efXmAFI4yT7j
bQdEmses53gl9bNi3AkgwRTUijzlneoDY2e8TAsO9tcrcggMdvdhs6h4wzDck7Jdf7IvGCKMLqgR
moJtmd4DhLgcLj+W8TVNJWK4ayXr0nRycpUZppkTFm8TTsOcN9N2kazMQcla3dPMCmF+r2GB0v9G
DS+FLXcVRQzEB1q5wekO+9la47WGWo0ooUtY4hMXKdsyI9jgSFpB3qEl0aw/+oLV2nPszL/iYToB
rLqH7xyENoB7aFc9+PfOGxUKZk/MGwXCb0NBwDoSwwzBIfG/ekdsxsjq9UGn0oAVRrVCe/hMrao6
0dqsSjvu9TDUlRbuR8D+2G6dV5bBgyfIxGherRs1uFgqYgbvDWXjc6UObc85QfK9B6p0rAIhRdRf
Wwn/ZGFEylXqCcWD0/uzKBIiKu89+BJLkzn+ZV+l4KWGkmkhMY80GFuQw4DgLu1AAKjvu3YCYkkN
yRDWW+uw/rbdiUxjrnmcvT1Pq4DlHL8guUEMwiigy2AP7XJa+R4qUsYHP5aSVyGvIDbIES17YTUN
dpywkxLqY9hyrkNHXBBKW48u+ZLuHfCjqRmgtEuz+BqvnN3TXviVXXNwbCKwd8Syw+OZsHUek30d
CZ1gYIJRaRQdXGUj2Ntk9fIzTFFBlSJso21uMJE6cL6BC1HUZad+hqYFNnEL/cF6XRLGDwJ/crJo
Uo8rlA28caFy9k71eVr6IlO4JGN8hEes5LwIeB6a/CEjZDek6OF/n+tl5Z70aXvISxQ4FT1XDZK6
Ldi40eFxA2voCGsXti5ysiMJ18XafgsKXz5lRRTrzEMsT+ht5ftrf/uBhmKE5pNkPbP4ACQFKe1v
O0pwoqwd9DjOgt1vhX6D+C7Q/YOyk9PSeWMcvACv1JyPv0fVH4bCxqcc83ag5iDOIQU0QC61oWqw
Vn0jdiWXcw4ZHqzk7vPMHhcfeMOMpaR0FyKR2ZFRgg0dgIwbhqgObrtsDm0+WlEoowKHdCp6BB0r
G9xNy1ZcD/Qtaupz/bhwuOl9juHcOk1UKuBnzOuPipkcFJ+mmqXjiEhY1bLoAT9LEGhUF5Wh4HAR
OmXRrsV94rV0O619NW7P3Omvs1p+/dWeHa45WP54MAWHlIUh77b2fsUbsy9D/pi6cEoG7mXEgkYF
OGpdSaFNZFoMlOVQ+NVK6qSiN1LFLR0Bqvb9yoCikECtC7+FAqHwGnb+cGUow2Qtgw+mCBrOOuws
FdtVgjKHkja33LD3dAAarljyswnkDOGUzlP2oXQJFQu28E2bAhsV+058swr1ARvWN5xcpZpYe5pf
UMjMs+Cdk2tst/PP4uUkmgHJyu/hKgWH6h59wkm2K+y4K/u7Q9YnkNk1/n43iHAjC5/6m0//NJt4
AtIKyB+XwGz2Ll9xI7tYLgNxFJ0TxuweQfIeb+JgVgb2cPxlyQ13czETOXdx0iByMgZDupiwGq2l
ZSvKoNXWdNnWPlvickoGdRv1XrmRlrt9pS1jiyMOg5XaNNUeglxzI4bQknRxpEwCpPvhwwh8EAnx
S5M0Kv5zKiu9taBDrrFoM3rtaz/0d04X7I66oca3UKWyZHwBJp+ek2DcIJ2GX7kkoSQ6EAYRbHjq
b3s2PhBhYmYdrqs/lkpBcNgEv+0Y361FdWXWcD7vWkk6MRmYZj1uvZ8g0YDG6LbiRkXxNEelugTX
w/lt1rVwEY1dgsjufSiV1MpOj3PwNoMaM2zitD0uTggfammeSXjyi/gam2R+eyUE66Dqq59/OYAP
BFmLS7Z/UvAjRCekxsrw5SKHx+gFsdqImPIBC//otIzW5t1ByCCOrJF7TDw+7ucH8r3un7kb9k4S
DNImY/gWxo7jYjZGUkYf9SZjgimX2OtqNJXmh/apVRY0FFB+xArBiaG6uqlMwjQAIxrg5Jup1SRe
gKOYU0DGT0OMnl+5rAIk0iAVhPwFkY8pbP7l8ghz/GfFt/tTrOwYr2v8cN7ri7565/Nvfarw4nkn
3PDFJl/WDisuzkuW3+DbegaOdB3KwI4jnuOa4HWbnwejGLLm3GdNp5wDUYr3otv+l8NpOIGr46oM
Me/S3lXNhDDO0B5YRk5T8Xpge1oaY91u6umA08GmjiMn0R+m/kItoG58r3yBgBJr4gwC6/AxOccI
4h6afYCAN6o7SxnCc6qJyigzpPz8+jT3e8ib8j/elUTfxtTOSqx+46mUgBu5KsZ0zhiAkdxzCK/S
quFGVozoNPJj9j2UcJ4maf0Jz6ViyjjLJ+ezYrrC/WrTkWAeXu3IvExkJuIuHtbwEvZlY79Klvsi
p9OR14WzqhZaD9H5qN2lgzHz7zFTm7oKIL+JzNngTD5rYodHun+ayI0UzsnLso9AurNgtRKQBMxd
nUdptCfJ3mfipQSLgINuq0X2fPXj6DxB+9KULNxJHs6RUbfouIQ661uBMgMNaBz3DAEtFUpIvqU0
I7DdSxqwAk2TTz3TUOcLHpiCNlu3++v0ub9kcjW4dZ3naIsIY4OfhpfFMIYOaMIz32YCsG+MSqMQ
AeGyfI5qEtrXh6WjFXqhthNABG8IriEohC1wDMq7nk3cgPFZ/yKU/zzlu/VItFi9E/Sp0fAXK9gX
4KFpQ4n07vkXFR0zzHGDMEjFk4FQ4a6LjAKjvliickZelv7nKjPUJLop9KjOmWcJhuV9/xYQluld
AN6yAylpJqU9FpybCbW0sKS7WWnU9zT1J7YzDKar3F8GSjmm0WUnjrRQl/cE7cNoA/2bw1x+kvie
Iv49mPp/9Y758wfRTz9QkjKRqynduhRIPWFYG5Pj9ciDFrpi+LZYERHnAs397w9Nod3RPqjGJyI7
scuPQiagh/qtwBDz3wjOUYeNCm7nmF8sSlZ5kmkfTN4lwtwxyEG4+antcIcK4PFS94YsXA9as/cW
mIP8eopY9ALhBsZgyz4EvN+thIykw9Q2xFThdH6ZdMGAkihy6siqpYYIzdrkiTMPX4+cXAjXxZoC
iCO7BYnIuwFVykCUKVq2qebx0h9ljIV7hgOSxAahY11lkrLehUGrQ8bM5yeeS2+vV7KIcq0JEsrK
eMRGo8Y7viSin0+1m09IokmVfme2lhld8XfEcHLW8V55tr517iELwtFejQe+bGUjp1bSw/1vSMDD
az1dlzGLO65NWRTTcKod3vVfVwtpA3AFyoIPla2rr4+ndoCwTmhy/heWygLs0CDszn9FFTsNWu14
547iJy2qXNZDPAhhdRMokZmmj2tNrTaQjArLPoaB1TrXLC9Qtd8KPApREi4+1M5Yl6iR87IsngMQ
w7oywZltcokFyzbvmJoue2JcXbJrXa7zcL+vtqNDz7IyUnIDcqdP+O4DaGPChVnwRJSyzMRRyXU0
UIrAxFTsiTtM+TrmcJi/F7zVjHQsfITi5lLtvlHhQTeTiY85Nh4dq3A0raHfqj5crpn/q3jD+3me
a3eJ992rikb3scG5Q6VrU1GXkwmthwwJ3OFnZMDv7Th4a4EAJJIMpCuIhx8aXi7WKM3LOr/5+iq5
wA3W1b3qgsXpY+z09p68WQetXAPNU1ki6k0WAvtnIZO0i7cOK86eIjzv2D3CGzBuzMLWQJNm5Og7
hXjAobzosnUPS34wXaIv4neG+Cbwq3sMj+QmZ2pGZ/h14k0bs879O62EKPKMFCrRUGwv3m3MAqQq
4FB4NzXJhoGW97QozYxm+sMbq0ViSm8Qrnyvas6motHwlsk2xRQwhCLCU+Y/juBbq/lE/+2Nq0rA
8TZNySS6Vyn8e9mMilR5PMTxD5l1bx4V2ncKelhEdzZsu8iIUEav/EEIRGJWFJ4cC270rKwr5O1h
U1VDW23Edtabc8PIyc2znEFpOIkzmahxdj83iKKtJSPli57se2/SNsxo7E3UeBlEXSb3HHShVuri
VW8H29AOlpAvgdWfdXzIO/JP+JlqvLm/xpllF5pZ0xnvVnsxGU8aTZsDX9mVbmZheOeRU+twyZFD
W1WcSBmQ6QaCu7hbHLozs3YuzVZU6jOsSaBnbVPlKgbeypmQUxrA/lJLeu0l9jV0qegL0Gqe/GZ0
qzKTsBHP6CMmkEouOxbLzQsM64WUFmEDzPVur3VGSt3ehyl18JXDNj/pGcxPBFHlWe16GCAFEt95
7R4WX8NDpdFpPSns9jnzzgqvmyeK9K7lewlx0zjDrDVpjkpEpe1qFb9b75ancsgX0XgC5ULyYYeG
0S9DgiSIGxiK91vaWbQNnPYcJO1JTHdFaaxImOgsBQtrbzrhkFip8PxuV14syyHb4lw2No+LO2ze
jeLTKe929o8GGTIrfO/YeTjD2NbibCQ1jeCpImEbuwdEfqeu/GgpJNws0aUsO4l8y9AO/2X4gBBB
6/7JgDEXXEdU5N/CtfDQ+6w+byGU4fG4thvWdQSILwmieFYJt16qDZa/7nQdpYj8eD3bEbCyM3CB
WfzTiAeucSz7jSqLUAIHo16YNEgqfPaRv8IE7b8t0fOHOGx27B10tg2Td9LStEr0DgygOEvRS4CA
JxOTPsjfRmv1KWNTBksqxfUWbmsxejvpzyrTRJlFAPa+I+vfDXdXp1HucusWh8z7wHRzj4UNZ77C
iDvXFUnNYQWgYC5Gpwaaxo+/2QFRfve1Syt2jIoROwkpWisCdyrdgptBSq0yr8IoGEhQzpNvW5Gu
/eZGL3xv6iP1eJeOfoLSMge74u3YCD1nBIy4/Y0rLeBLnJZuJudrxRROxhgt+1dlSvhla1X4kdbV
HafNs9eSb/mrvb1a6YCpwHflMETNlCIOAolqpjoOWXVEFsUpPfhMAVuYhgKZrNLQEBa/4/ucHmzL
4o8QA1DueAz+OO+JUFY5QJeKhXx1BrwpD8R2e5yl+MLrdVfFLGUfPfza4tHRsW2xpDPWt8xUzgsU
wH/PCnrCZoERdfYBAaMfc+a03TGzCTbok2CJuwCzshk71hKuVwb8n94YAwCjp/LzspOToSmGlLs7
ZGdajHZV2HnDbdZLHrY3kBkXh6wnUz66S0nqYIwj/IaS9d55YqlUFqdmG036zY3FH0mgHy4M3GHg
bRPbthGmCJfGV5TPhG8bMcmAtdVXZAXGKsMMxaYBRy0VALHSw/NtgwCgwU89/Bbw9IpULe4hprFo
1MrClx7gGDGZlb671Pu3QZamnxjijAmoDglDKs8iDDwWlN8FiEJvMjiAJ22aPHc7T9SeMtjuiaZ2
LMoMg4bsXKq1qcVQMUKp1PCyl4sBzeXavLUT0nTjFdRM+L2Oo/qo3WUlDhy3MzSlTKgSFMpGEES8
xW1IuzgOgkN/+ScY/YTfPHvAPtDRNKzK9YUH5b7mwydvc68UTVC321yLXOY4kv/VOal9UeR9ns7F
qMSuJGJfpOxQEDzMi+cz/C1Kwgfje851q+FhBHF+eH1oZjzeO0RyB97yH5Mwc6sOr7CRDMTi/0gf
zdSusGu5jZKstPf3Ry7LGgOPDfnxHrpLH/5XZBd0OTkGnC3M3yCOv4DNVi0pp/bFbTytXNTelIKs
g0u7wunYzPbh7HdkgdcZ/5kOkxirXk9HvsSeGCOEJ+VexHq1IKy+eQED9wBcXrUqhP4HC7wJT6DU
miHlwjpL51VPCWj/XIxGOBuuz1WVNhIZ39S7q6lE0oaK3iJHf0cnJy0Y/DBj0K6nGq2QP/jWdj1Y
EFcTmt4loAtI6sfmp4Um3sdtTHoSOBQg5XdGIIo0z7yvyLvbYy5epMpnqte0XvEy/XDoQ58K4dOp
nXvsIEXRDjOqTgU3eOBbm2br4OGxXfRvcHUR+sZIAmpDgj3YOHolzhKVb8CFDla07bi22rt1SLEy
nXphyFNfAHCp9c9XvVaAJXfYEjBoYd6Mc51JBt2WFi/7jDQKFJEN5uEGntO5ReQFhGoUZXpRO9sx
oKbv40kM9h5UOltzEGGxekKUQXlHG6V8igvL0iBo4q6aEbcNAHSpdxnUqEyxa5r117YKylzX50v6
pC4DsOo5BGZcWS3E7GAmSMkfwWNduP2DTwW+ZKY/6x0xmy189V+oMdqUe1F+9mGAaAtsAHhoGddB
Q6+UyFJmiLnh5JRy9GFgW4OSIjeRZBXqbdyxs44vdf7OuE+fDCtMwz4jeJc/a9n8fhIVdyfdFlHS
sf4XJ+H9s/XORPQw/Z4cPa0+/IVdH3fZt/nMxC8ihwe1J656f83ADLy2J2Op6ZhL9gWUDsoA87j9
SEvOTW9nVSg4ZPQfoQgw0JcWvWXckt+LI6wv52x3g3yGtyAlNoNCZ4sybxSyvJoNd4khTWASkZBD
y+ST6bAoJcHL09gvQkDU/sj/BOFUhiwHr5WXKE4cA/S6l/3ga9rkCNahnmvIiy2/DDB2dXMbM2wW
vndC6Ocg2VjyUaAJpoIwDbsfVj/Jma74+8f9FgXkeBSVaD702tpZy8lxXmfRMuyTBRvQ3NlXpXcn
DL20AI0/bWZesh8uSnqo6+iWVTwDYqob2ps2fw5qkEef1d8hFlbuifW4i8nnjvTxEksIM0RklzAd
z2c3VTjypsWHMdg7bitANK7Do5L5KLMUOQdsqF9zzjM2RpX5DjEZfXHH4+Uw1xyJNFKgVW4nHB0N
VXOOctUE6Wtwf0kVtJuXHcHzNfmnl+XLpDqKN8aMAsZwZ8nzYbDMCzUh4VCZVhwLD+Qk3WBzLk+W
bNSIneKvwtnC2MZAQtQB/kSTlkVQAQHseKVdFXgubEH58kqJyH/xmv2x7o8UMLD6t6qCRFqySyBw
OXdn1fY7Ft6kUwxMrif37UJE1qdTuCI38EOizydAUg3W5SMx96cViYPhWv99ag9BRZRfiF286UMn
ADPhLB+KYzLpgcTJVW5t0MeqJAkth+b26JSbfniUPACWq0iNeWH9tie52u5GkX9YzDKzXEcr4lK+
AkPoG4DB9P53vVL4qhThGws954v3UIjldo5Vh3VMopydxWKflqqllis5fS8QWiKWaB8S3wFhFKo2
ZTyt25LZ6sfJGydjL83Q0bbzMAXFH6n72U0JDkPHJmgGKXkgRf2gx+4Qpj11NXTXJxLUEQsyhGo3
3zsUTjCHY7PgL2hvaM38o3C0EhziPV/5xudCcle6azga6vSayxm0NTZVEloSOxC/dvLhN4S67mbS
0MtMmhGSTR1QEfj8i22jUf3kwNbRJnurQRMrToFkU0BxI7jTSK16AU9sQ3RUYAlsJjATO4kvJBq4
QVYLOhTXAYTC0dTYe94Ni7ZY3hC1k06tAthSKXOzSxBNtZ+w6UJVmO7u0r1wipzBCYuyzuB9o/8b
15HvMQbWfZHhMs/h4sjCfjeBPqunQZuhYIesTurJg0qNvHT+vRP0odM/wu+QXTQECvcg1HKxpvRt
pdulvUBAMe26NLsXGVaHA7UeHyLnO2v7kE5ChUL0pyDd3Q4rCxrMZVk0rZs7BVA2O36JzjwvNsnO
R0dvPkT9JDmGnHsyo66ESnMACijlk0nULR00U6ep/rfvA3Job7qFeiR88LiN2QFPCMx6ersTIIsI
lZkyaX8nIUxNi+q/L5BHEEyRtYX28Xzed2r97dI+Lnyq+UDX9g1zv2KL582Az0YAgVuaP9xiRMRd
88wdXe5U4FnFkVIE2Ce9eNJYLUR6VOie6T68r5dMMbMetFHII8oJK4mU8155L86qpzjlBhI7fV18
B6/ksPlbq3LIWWvAB63pIPXSqyUYN1y85GrldhPzXGJIpMz0h7y1jem4wtc56w5tWmykJOoUB/6R
PWaATtTEXGf1UGn5aS6ekVnpvCQ1fG9BAgEYh8Kpzg8/jmFSl0h4vv6P3E9ZRQXZz34Xq42zaX+m
M8PPErq1GFluPSCstC/dmRpFsP4tx6L427n2eBAzogIsBxbrzaN2VYCiUEhNnysK1ymTsn2eMmFg
y5VjoLn2hU1WQzDRQ0r+MQDyX33GdN70dXZgouequwiDU0Qu+B+qXrAe8attNaEfbvDYwvKQI5GS
fiA27n0rCEuVtF0xh8bJyzcmAmhlrNOyV8+Sy/3sPXjqv/mOWvqw35lb8/LBojffiuW4vY1s2YSv
aeHladoxLzdVd67REZCwC1ZJgM9JklVZu2VRTNKeno5fYncjIQh+yINUX1tQnxlAW6TPAMysbitL
cI6eUoBYwTvYRICRBbelukEzRCZ2WcEr+Alswr+Pc9k3W8JMCC82YsacZDTdl86s+bx2hyMKxMeK
J6ETjLNOg/kPZHp07WRabmyIn+B3OJifInPzkgBuSnhC52YYIgUvPoFHi7I4/tBZf10CzLE6XYct
Vnf1/UmYHrIaz7l8dYWfKnzgKyKiSQ8SJLmawuirKXamQH6JQ/e78szPnq6ZNcykU2SFwQANrY5R
yD5Dsvh2eQZ9alZBkAhAau8x2ZPlIu0GSKhyIZubgh1ZtDjYzcgpO83Um0CTLJ+GvOKTN/s1aBml
pHGYcApuRZOV64cVODh53J0Agy+NEKFC8e2nISveo6/5Q4x4fYsV5/PWZnne31eJljdi104bc5TI
NxLVBo5M1eHaavu7zBcYMbJUdGQ3oPSGtNh6Ad+GemkYtrZgepjaG4NgvewrupqKf/CUK5GsQOAt
jt0RHGJ9TNASabu9XGjibZ6zBnrCZJHNVftxwMvhCu8cRLBl6yQwA0BNUm7bpk3UXBKcvNrHtFxV
tYZUpimDhgw0MfmtkrWMhAZCcWNffPPvB9xzwBhpKrMG/zwDm5OPg4hj17eaNcWmUN+rGM90YP32
rWVolJ9JZTswUjY1UXEDC06+4f9JPMKIVGAOPztl3Lntwr1S+x/28wQ/9ngPt5ypIh3REcoVqTYI
rM9I8ykGrpxvFsS2tapwqeWGNhO0ctc1wMyBiEctpBlvSR4+23R7ZvHOlDZxMT0ocB1+/QyMaO9G
xImNg5HZTrx8YEZvA13bMW5zgH71sjTyhYAhkhFBH74VislWpb1O+b1DjRhjoJ1ZtHd1c+c7TLpN
gSrcZPWjRgY7Ie6jv2FoL7BZIhDfsJXt8BWJypUAF5R0j5Wqnk3T/7lmGnW9XtbXGGeQbJOWidYt
bqFM22O0ZJ4mtI/w4rQw8un2B2FQQ2LjSXQExxid5P6VXZaaV72xosVvhUT2PVLnbo74i56O87MR
m2i4WCyDfUjmbX9CtCY4GcOor5VjiNsCACYZ70DAC8N+ANeIdCw+o1RmO9czQWnphn6XRJv4Rf+3
8lTf8PsrJUf2KvyyjNhuN2VGALeW4RXTaGqKP/r3YjfEJA1e5PtoUqfjWQgsvDVIfXjzjhNLOjC2
VPanuitGEYYkMEKmW812g5gEBT51mP05engJy1oxzMrSEpI/3EVejLmErbj4MpgUOcuzhLbOmu05
wbLDDy/m3fFsDbzIRraFxMBZBFjO0fz0//FgX1x3LRii2eEoHQJKXT41NTc25hvojsIWVHbthoV5
lAt+zedE2/76QQ1EQUst+HDPiwiBe6jb1It6xybghDl9c7cXaHK6N45+iS0+ObLrV/oi7M4HrPkb
oNh5yUJedh71cEJW/IiC1w5lSVkhNVZ1OZgdMItQCA4/k9jV2xSIPz8pHXjZI/vkFDtVhKLveMxq
1dAMeykAcUjFb8UGGjvRPlRaDZXZ14WRLOUZX6cByeo5Q90AAs1bOvm0JXtxGM/aHE6wfuNHlhSo
VzeD9T769zfd3vHh0OAiVZUdLAMpovux1SJR/ih6nsd1UAlv8MkaJhVIwYd9KGwiiyCSD6iy3XPK
vUMjeqBvX+JNB+dUdeK3mIfB9J5VMulJSjIc/gGFsPnAUsaA58HCcG4tpxohAScQ81AgqbbsrGwu
BMki86piNvZSNBNySI4jN+SkElC7ola+3PJ/u0+jdQyizHxBRvx4P7QNy6xBgdreWjs6w3112oP6
zUy3T3iu4qf0IDJzKCVmeG+vL9lZkuwen9oWyKazw4i1RtrzLbJpJQ50uyZeVG0lpXnaQDtsdoaV
E1N+brSwjjv0Ax0lFpgwVlgcJAQ6KjwrYKXdYnxcm03bysg2ZFHYFoY9h/tqfcXVkO15ggiOJn49
CCETwZz4et2b8LSdZwntCp0kPRn7ZxpSYldzK25SdImxjEFrVPc2sBFn+VbZIf5709/+Lr3dysor
kkLxyc2baslJS/DOnaL+6VdVa21Ea1EytXFyWeVCXB3aYmfrfWRNcNlHVZvWph8U1vP+9A7WbHMu
3D17fnFtlMNVbvzNe2465nONL/hf5Br6W4pYeHrZQQcJrVrjul/YPegGN1Gz3wUBWQrEhdsomJye
mj+DCQf8iAZPvp/MeJSNgCl57oO9vMrjzvBQU8wivLXfCK5eW5rueLd79UiPksJnvab9q2idvQpY
PMzECpNqK30BKGGPqJ8Rce2A+g1cjmzecktaVm4dN6pgfUH3Sbuwz5x8EhFUDtrP0MKWAnMVduRo
/elsTbDzmNJqFU7gieFKtBX8hoySwu73yOEfejxYrJBoHn0DpXL+iN/BUl+EtKM/4HlB4S403dVw
VtssYnCcbUywckfOpxdHzYW5439O0be8sbUlDZJieflll0SMtdgCUoDDIs50i2RPbxtgg7IO20xU
bcSVjMCJh0hFw8Eyp/QOiggnjvfl+Apj3L7phe6JnUBLCp0jYcJR1DN3QDrGflpE39wQ7xPLZUsz
1PWO3ASC8s/JiYkIwTmkbmJWXaL/JopBoxTuwgQo1Ve7s/p6Fkz+F8oU99z/UXTNUlSZjutuPDtp
/rHuJ20+7eVZIqJ/t1tvGxSLmm9NrOVRhMkfHCrMTjoAJbsuGL38EqMvoMm95npJDCkgzpG4YTpK
oarDgwCuZV+NGjVrkf2AEsFrnKFq96enLoDWKeR29McKdOQpRpJr4pJ8tFjtIjo+yoKXuOIqeQ5U
IdvFToR/q3Uhz/Ce4rEfFsGFmoUD8rNB7SF+vSIOSaI/87OdHYfdsSvdBUvabHYpyxYUDwL5612w
ZTkvR80546yUwn7dFf7Za1KBnmZB7L64r3Fscxf0Gmr/7Wgr+uqzjP2kkernHL9dKgtdLlPotSEc
wes6mEJY/gwIlFToD1sebVDyKjO6i3FohTK854tN9iJn73GvsL80Bmpdx2NyeEql6HW3UJZMM0IM
twUljEzE4kaNsh9o5OH9k5URvfb4pw0a4VENY+GLicN2n+8333nxpXTUrktiDrBaQ/W3y+2BZKBd
4cyoCRLfP1atauJ/DN+uRsP9ayeYWdWYGXKSYZeZMr7/joiAqHTE42mUJz2d+V7gyYx17nfK3aza
oGgioiH0wB/BNtxzEzku8SVvG+xbQ6mBgNIvFpDw1sqLu/MHGjrW/hS7JG6Vu5j6KC4m4JDI7Odq
v+lw0M2MYe1BGYgv67Ktw7ANn2obRlisTqPudUzzBbM3t2diBGEbHMYAf+7D48GcCyI3Tg6iDQ0h
ZpfZvN8zTgZVF8KeKogYyW9lfk7JM3I6iNjMnokHBiXmSbJJ8domFKfvV7dQOMfBVOTRo4rCDU+q
r685v1WfTMKCZAEPXdR9ksPzctxcBgGr0ftNhnOcE4Ab/lpmrXA8nA1uHR5TeAJWf34NIhpjz9C2
e0Pecrr7YJPesOpp/1RxwwwBlKIUaCXrb10q3C7XkuWnAYziTcwhF+BZcjYRZtquc6sEAZ7fE1iq
AD3iJHzmIQFXTHuQrm1mMh1rTxUKCCXjpa2w5VwiKbQSMaHwOIb+n6Ez3d9uDERMMC/WxLprjJXp
T7kQVH/eMLdI1aPORAGqIC+hOiyveUivDuAxP3CTSD3jq8wF0820zdAlvfA912Xe+2sbeNKuM+O4
AI64sT9XazvO/VeE0MVdnMgvd5rdy1+KsbBzRxT7qkI2T34v43aTlc2jwu/NSFGazxe8W4Afy13o
anM3rfZGitkNipCHpNzIj+i+Ezip2LC2RXJxCijSP+roCnAyM0wsCKH5lE5VC0MntKWzucqQEi/e
RArDOMSqUmDxjlFnxN8Z2cLR7/uHS39GDRnn8vB4OSOAonrCb0vmz39xnf8agilKEoFYZIGRF25H
CH0iOq+Jp43AvO+klWE+ZS+G8P23NtCHLkDP1vMJK5VXZSDpqMJTGdZ+VBLsE5cVgWkUNT1G+dvx
Js4BiERpAdjyTLC+RdwDeFU45qljH+0CLugFJ7aqRs8mwKWlbnB8NmiFSxcTlKmmCT/UXxmZ8NnW
XqM/nMZNdEBae6b0glAFUjWxSn5IM+aL0XEVRrm6bEYVbilM8undGphCO65VZRL3FIGnk2TWQnoV
T9ImeTj7lE9aXTzDObImTU7PDBI0R7Kf0jpEkJgHV6iZVNiBEz0vq8qsOvyx/dwfUDdsXFiSGJyk
uwB8kinsQxLecVYZrqYc4jr0WamNHIQcKoEfby00XyOKf5rnvHFy7G7elsg9EcfZ1JNfskUi/pjf
6T9PLmt3ui8kRCZLVvpoMqXa59u7G3p2vbamHSmFI+1f/xC5+TlmMVjtByrOuQprvFpwoUtMFSp3
Kfio0mXfHPdV7XpykZHQF2Efrrz0mtpbI1mkqJQWB+727bjKVD2lJYJDtFJoxRzIwW7WllXPQUgx
vxLcSDbnTG82OXWL4mUIbwUe56tgUut5/s35+EYgivTTKMUswnOBSWKQTiugnndxjjDJ92+jX/5q
qSzqAGOkiDEzr3jiplBI2Xj0qS1lt9BpXxxyW3h1aC9bWaTp9c2uocCg9OoxeWS3WJ/c2GNpor6z
e6RGLfG2ys82tCoJ2y1ZA8CViKmJmXjRIpyC4SfKaoMmil+EJEmCyjwMMJTzB62mHEkxc205PAcA
WrH5LQ3/Q3Hb8/aL3tKtfmjPYty81QIyRKSQQFqY3H2WNBumIx2wu8VJqt2DNNX24aPvgq4wvaYb
yntIWEuTIX/NTdpB1z5lU6lAXWoQwHYRDlJtvodUzgsEMNTyMaWPkEtpQAkiPEGSylMiM0Bg555a
XhjmQ738eS3ox4/kB/pjMMyWuDxV6hBPZXRPWvRIeIE7wIjzvMPZnFYHYkCWJTuxtqPhGIY8OSqt
/KF/q5WGFBQvUlzX8dOCCdPzFlrO4A5KUZ2lNk5wJV92Llvfr9//c9uWClSKc65fzuwuVNiEl/SF
Z5nm4OhJVvv/BDu5QgSAiR+BCbj26WhECTThBPXXd6MHlBVlznYoeqDjHvtDkdZ8Yfx3Gp+SAjlm
fGwT6pvMNTXMm/cNHf4uzlY9cfDz6qX4+fXaxp1eEuvWKix/473JmD/ghF5FDJuI8ZGZlc/DmhVq
5RViGUoNsxFIyaO44G86uYm5O1MbfN/ykIl4IcVBdfdRB3I7r8TKxkxdUEyBB5TT9+VGUj3+4Bm5
7Pl6LpednNdmR9/EyjIq9+rWxfHfpi3FSniXfG8hYtdyKx4T0cFqkj0ireDqRsJOxumIswHTW3lP
aF88O4Zgtrq2uSDfVCWX210dkURC5XoWXcwgpqyJqV7sXxvHrorGdMP/LffIDoOFkLmrVRR1Y1Fe
z9wl6RxHzOEWFuz3sOC6N23eeJoJOq26n5KnBv1Z6pqFatm64Kw0PBKUqe30eB2Zx/b29CU5Vg+6
aa92DYXGJy4SVv4qVzmmgOtVKvKM2SE28X6w4kpG+XBqffnEhUaUzo4tvKMN2z9AZthTArOnnEho
1uJkefZRVpHUyDLsiMOkTeZHn2OGxu2IC+cTFm4cwPRINFBE+pqBqUIK/GLxHJLako5BO3TuHXAn
OJLF3fQ820AagosxTX8Yk5mkkA6NrdJwUOxeOauNlkc5znmN6OauvhG9N6MmPLAlbed2p8aYjQE6
K302Q4lVLS0jMuc4aRbbYHGLFMP8AhSWw61b1Cu3ZX4Pd5NszkF3hxeZjL22t0BtHFn0EtgUix2T
M7o82I9kJa7TMAaEcwk5M99IYDfb9uWQlGcXtuOidjfRryz01EXp3F2m7CabbrhccCZvLnW5BZf6
1sYBMqA+3No0R9Dl9bvrCI79ZfV0vwyM8rPL7wyi7XZQZ5AuS10fmp/BzF0eIkFRXg/fGSDpVWJA
dDs+0KGfWlU6CYT+LaDR15IMSEDM64lJ/RZg0eTKjylZCpnocYp6pXWC5nkJG7IVdbjc8KXv/HRe
tLhWtAeigccRuS3WSf9/Wt4bDOkXcMD1OekYTLqC0Us2GdnJo9GwG23GNOI6e8WUE5bVf9Djvd3C
MLCGmjBRTiSoBmKZ6YkNiBgVHElqX4ZMNvifNAuoHxPTu9UmZTurIKW6pkgn2O8ABezTvBe0Nj9a
JvuspEmAfp+T1iC9heNeqIA8qyscBhxeu4eFz3oGJZXdohUz+grb/iI8l1s+geDqKmxU1Lbci8bu
VwF9M9I4LJCYT2n1wmkaroNXMbrUFRW6TxXNCujG3CwjDm//KlVnSkCqUTAfFVuuibFFVOtJBhG0
VDRK0SxBVNnsNOlDqDE+/LI+1KlEnMmMv8pHKoh0Byy8P27v4GgulqD+XzyYZu50ChSXe3qeWCP6
HpTqP32jeSgQwMxqXOYASCzCGVGT2WD5TOEVd+jhkmqvlpzSmKExhKENo3CAsGPkZlPJv7pJfUC1
8n0Ba01d8dg3017o61jMuxeVHS8LoaTMiJPMLo0dSZG8f5oAzR2DOpAFakqZZLwbPm4uWlWsgPTo
ypa3FrPT9HaCfdB8AhJlMyOu0j8W8Ufm57rLuhHGlxl6Nl0xHhJKEZG/gQgbsqyegfLr76K3xkIQ
QIA3LM4ymJVpXS9Q5+PgbVx+ymzeMdush8xtDuwlWwoEj6gey/3B4bG1iK5nyM7c4FglM0Pvfnm1
pnWCvE20aYQRfN47NaxeO8YIfzjbPLcgontI3a5k1u7vPcKeNVqEwLR3Rp2mXriqtqANxZSjinF3
nMAZthm5fpLPkl3sVfqG2GUleOYYCQOBZb41mdB8H6WnpuTM0u7idAyXLBqnQP5EYilr8haknUCF
Zut88UYNJMJCgAt6Y2LpnHBiGJy+PhqYK+r/fAhPBjl70g/J3blONR1EiL2CFIJd76Qzu9dseLg9
vw436V0o433NUqNpnT+JVzKuO7Te3SS9f/zFMlHtYirdXoNHacNOHtxg/DbiHjB2mQqBsc+YUODb
ciWBHmFTRFjgFMntwfXgiAbaUDPlctk8kE3zqaucHEEjraxQhd8WV01r/zcz9GObIaKwpOgEd79a
Npg4lm/zCA0/dHwSYP721a3nrN8Sf/nA+B7gTyVFyoEtY+GEf7ar8KrgxRxlQkbhMqO/WO2lcsWc
y/vbcTkdu3nUUuRI213lHory7RT6myc6GdI1coegLOBAHaizQS+hxTWDAHpgk4Y+l6GfLWm02EgS
QG1FiUb/BpchTb8MbqbwwgEmDuUD6jQYD5VRsSCLdX104nBahYGNPnvMCTOJw6K37+tW8QbTlsJU
7saFFQI2aXkoceWiBH3IwAEm5oWrbgXCN7VfwbYuDZoYeZJrxsp5ak59/J5qi/KpIb4UfUgQogzJ
XIxaTxgdPhqzJCKKSlxKwSBgffiNfbX0C4+7a1tAx1DNiEcKtvTg6+8qgm1bDdcesQqjhcZsWJeY
U9kQYhklfJHGxdUb4WHg45JjvGrPewgCNMkuQ6AsVAK2cufeJfD1cS/EgnQVT8hjn/dzLtjg2+Th
U2FzJdhii4wfPvCBzcz/M/KnFzftAN6soCtnAfiFyLIwHJIkgJt8CMShiKiLpNiEfV3M2kMvMluJ
K8RhjEZ9XjxkKfMCsrSnM5C0o7qHd23/3KHohk38uQ/3In+PG/kltNLDMB4c/gM9RJdiMuj7PRaP
wvVPzmJVKCK8D31HNBAjta/doUxdfezOg4OiaBHD7XuSuiyL7tTWhirD8vxTlv92AR8OuHmYbj9B
Jb1jZCQ6JiJhK8K/ybr3RjEFdeo418x+iVEDye/bdX0VqD2ZkjcQm2R0kamDdTJTYqTx255KfNzB
5cfqH7o48sgSY9oTw4mbovFCEpLTPfqO8ZU6mj42/ZHQQdSWUpEeSaZLyB3s8gJ11XHKoRUvhNrf
KdH+11L0VDEi/eqslerVZ4dNHZ9eHD5h700x+hPU0fYX7Gc8O9e21Ti1+cmd1jES58fUFCFP3Gct
u9sthC9N5aaoy+eQKFPnQLj8Tok2TxVekAuJ6nVij6QK7FpxxY2G03p1K+F67NaRV7byEJf1xdtP
z0xhnj3Ucar5TaNT6i6YbOIfTjTtSLRgOHmgaWDxfuoveQ1EmQw4yMfI2U0zV3VRac0gnVwRE5aA
NqoV/kZUBv3g5+ycSpvG80hS3vkW5l9GlSa3tPbbSunAPkH1Q5Pg10uVcOqL6SC0gVSJeZblseGG
IjMD5kQWkA+9h81GIaUFw/6Zdi13qavX8GtyO6BWiq4o0iZcZbKu4W1MMFtBjfbUrUrzc3LVlUdt
Oo6UgY4ONG/5wQvdlMAtAs2jSXgkHGF200ne0BLXrcu8t8JDgCR69nhIhjxTF43xIBFYX5IVqGYz
2Kz66tZZPLwoRGbe4rRIE8lNLMtfQzrlFkTMt2epLL3Dvj44XFrZ/E+rqN4aC+7DZf0V43Sk18UT
2OvfrC5vE1J43aJYR248/nzPo+H1oBVZXI2PihacRM6IjVxYf9PwCfW31U/6ZqlU0SyrQG44DxMN
UY+LhydUENULHMFCjWcSarH4qrj6vMrN4VERVqaohGADuYbVLDJgvLRNVWb3vuOuFQ8dGT1D6MVm
Lk2mLnInmY+7STGGLKvLq43jlOuj4/jEE9A5hPXlq98bTzC0sPNpz2aAqrPnwNub/35JWi1PSFuN
pcB8cmbJoYOVL/GOpzMOWxUEoHnMTXBv/MGbvCzST0vTWN3JRhUzwwsRHwjTL8Uzr2ZDK0S9rATT
twTOVcJmzDjMfnBcdCox/3UgNronfGsiSOIdG8Lukr2H1SEgGh01r+83EmyIiGemQzhPa9iaV135
UP8rxpJdRbaLxTV/oouuGNB7ST5FvJZyq3Ir3QBL3CGXGbSD/eeGBnCh0idZPqEcvzXLm1Ulzj3t
NjTrF+bE64HXAGJXXd+241WyBF9WXR7Hf4FlL/+p3imlWzuraIV7pjs3FGd/lk/7kc1ZOynXj127
s2UzWD20pE95l+fTvonW6+/La6lORySi/f74y9/ribiFsN1vYS2Aa5H4ag1PLau3pDhb3WSRNxpR
sOcSqHTzV+eeyj7KCugAXtNqbEvef8ycgHmoUCwr8r+upwE63/j0NMi2YAentZOucFBPK8vMVPui
+XKL+fWjJfMRf5ANXQPLRuqg04V8xrOIMI3v9h9TiBBnVX2x2udb72ayuzEVN/UMOH9rMMQTBk2o
jBQV1tf7kkvX1cxuhz2qHyjySnpFQ+wgKKSeXg4EjHfkQxWzN10mNecsSWQmHTnZqK7aCLTa/jxg
C3x2mF1qSdGUnGX5taXeJcqSkmg6k7/iSr+AaqEs3N4qoqzfs+kLVSE4NNCXtEH0gH5pxdwjw76i
rW0ilwaviglbzNVOMd4QxE/IVRfnUcAUFMEk+zppWCc4uBnC3CdwsoD74cNyHwuc9vmYHSriulqv
a2Ulq8h83btVGbfZaVcV7/MJzufM/vpT0kkSSdDmCjlKCEhMYOCCSzXiWySSEDllLgSVaWEb2WuN
34GEpMmYQF7bNGMq81TuutXL9jgCpxaeJ/61J773RIFdXovf0SZbK7QKsAYGnYsI0FU5P9hDYTD7
k4+eL/WVl0KdkbmYRZ7hpbRmHt1pwrm5s5AKAfLzHAKxNWYTqHk7U+u08EtaI6l7ZlBxVnOJAZl4
Tb7OtY4D73cgoI05rdfc7us4ypAknIoUeIt7p7pzRFi3aPMOA09/gqXe9e3YDT68tAdiqOA+kUft
3jm5nqAiun+IETzz+PULtjhe3VkKroh/4mEVeBz/4g0mNWG5qLK60bY6E2j4S6Whf5XnLNs/7Hkc
p1DOmIrwzOGZCPQoD89jn50npvJjK8t80u6jVb85f9uUdkxjCqoDDeZAlQ3cOTKD6QkUEP6AnmWC
DeL7GGNVOrfG8Q+7xbKvKQvIhmhjXntujMax7lg+iqg5sAw1aoEEiSi76janKi3puQ9D0lE//wcc
Mv1tUmP1d+76RnWA4zxw6EV4cxEOQacmh7dn4QMymxk0+Fyc4M8wPUJ4Aqy3hYiSfI1wjgSB++T8
r2bVN3vJX+KccjqOMaqkuP96chcU3NqT3m/ZLuANZSI47JgMucFGYpa4kRaREjDAlCvoVn4xWFsw
7S69TGljNpCZDOmbOURgcrJo8yh1ZlvgiiS5/PygvCaZy6sclQz2doZjtACHMt2QpA+kQAe5GZeu
OJ8jB33974R5+lqeYvDX3Dm4L+Qkd05fIITUx2z+xskyN+hhUoVF8ouoJWzU58eaJ6HlDFF9UufZ
pTQ8mDqOkakFxGobtfDi0oKRIxIeFUXAYj1j4ynB2G4hIJOpDiuoHSd2x8IMOaLhxAfh54FPfuYs
nN8Vh1XfCi6CMZSNASPSo86WEl0jrJGdbol6rNk5D1d/ih8okZJsrTicARiS786wKHHVMqkpahdz
OiQaG0fFdyUnF2aAMN88CDVvJZEtbhWM77kQgwucYNwVVK8jcA724++fmux/PT8vui8m8oT02T2j
y7Hb1Mx0jJCDTHZmakKKl9TjGE/dAxKNF4E7h8zLgCORUS9O+1BqEQd4GqpwhPtkq5h+IWfhgtmB
3dgF1BkP8xPZFeuJOSACnGDD1E2ZeSLnceg7fEAbI/2fsQEMBcFDLcXUwTLfHnfkKuSsfujRjIXD
dkVZv0dSjBR0vHak5m2wC4DW+tFkTGUU+1+yK72y32By1X6aD0hh0js3IgIeTtesfSDaEAl7B163
bHMimhQ/zVIZOORPtqBP4oMGXQUe84IjuGcM0UcGxAeADyMip10t2ukhFedxKc1U3nGMJPH+C7QW
+oa7H7JNbsaZjKBW840I3gACAQ/Oi8aoqmybJVxKAHxin00k2sskNBG8c8SJjMiyGvVeSIQLzFg3
+ntNMaVJbmMEwnT84DjorIJBmWW+db5jgEe0XaIffMq9lcXFYTSacvTPooBTR49iQ/jNZDwwjRft
0dtDRyBc3EbhDBCkanUk7ifxhYFSGLyIzvPc/7KEFla9sLVreIc39xtDWBEp9BCzJFnL8Mx9ck5e
j4hurQF2SB0pnzKqA6FHbikk7GvhTY14yKpVB/AmxSjbLRXlC6j4XOkxkqj/kIQnJOGeMp58oheV
Ms0nXRYFJoAKozFgUcsom9Sc/qvvWlyRnY9ViYwDYoQR0MHGK8EeFivJEvgyXasVh0sUB6hgZGfJ
JQCN8LcSnQlE5wgvtX9iQxyGWnU3QEzpc/9BBZQ10daqzJNYkq8d4Dwr1f3QNuqE+sRYqf9GBOum
tumn9BfQttZv96CUsXshgf9LM44KvuQQXOpXTCZwuP585ihZ9jzlgtUVOF53oMGYFwydrUUxIDBD
/iHHKBbDVbq5SEmpvjWzz/+DF6NE5bOTabg/Ewy6ihagGIgwN0I2jIxQtRo+bMni6Zm856GkKu3M
0xt7MZkkBK0pUV28Y2pzdnaKcfxA2X5gvgfsEDYnQsuj01JNSElIbhlVr4iLw3YQ6TgzoOOQjhBj
lDhy8a//a9oMxB2X+pZbOJMGTJMXdl1EjrjhPPoXxWdFrB2YyjG8grxPY7NzIZC+WzDAZ7bVGI9J
OGuy0GhpWFpkzNnzZNTrftLi6ILeDlqHtUmrXVZtBqI7DxfiCS2mvSYXgcu4EjMlZHir9YRq2bI3
8SRXlmkt4fY9efYpVVFwKqFtns01cY0G6firewaCiy+Hj6C/CTCx7wJCmrVUQrknh4w7dh5uGbd8
7zYCnY2idh7oNW3F4x7RMXHGzwYHWfBosPpJMy3OdCUO4/SAVwmdgwwsxdKYVvuVUNVUyFQ0Mxyj
9iqA/f7Q1tg9P6wq+pEo8LpOX7e1ew46XBDNhqPV0yb56mLgeduq9WkienUrLgwkscIjsVNmEb+X
RvYOG26BMIHpdHRkHgJcSsFzR6g9cwKNcn6LoUjUZPsY84ubSzWyHRXcxm6/gprIYY/kvLxJ7NT8
l/+v0nmHyH1yg3oqhU6xXnJ92izp8OSowElKaVHLL17nWjYK7WRUMs834mfg036PJeXjtMn9mEtu
id3cPuKqeujKyvbnckxdcJxRywdvArPDuaRuYaXvopHOqhte1TRTTbG0uAudP6GjzU7FFeu1Wbmz
+gfNm5C4300pfwnlxUPeSIANx/oS2q4NUuXUIC9D2Ms8Tj7qnW9cYqsy/YUQS+fCiRQUSEYhJiQF
nbc0N4yDlEx0gFOorB61t6KWhfQGl9JE3H8V83OGmSvjIS7s6EJbtIYHpzixBddl1iFX/gKtITB1
VaVmTEZDcFUv1EBR4C4Ac6L0xlQG/jwBxXpsLQGgZ0hXfp9YqOqSpLR+4BgLdZOsHXd/yhCdMOli
BlzmjYezlbxOjRbHde4iZl4LdncCqFmqhFsTbWM+E9WKXoi5Nh21udkbAh9LH/FBPL9tdKsdjlm3
TadifRlNuhNOINNG6pWvz5Ejy+g8gsl6q+wMTY1OXNAcQ8PrJ+8KOAeCUjBA+KHDzhJYmuYL8vwx
HG4SU9K38FRHvqMd0sFOc545FxXETk7q6JVu+2snHWOFz6n+/nmhDrssFth9Pg3VjPy5pbooLqr7
nXMp6r1kG8lGIEmIkFQM1MII689LOzMb2/N5Zn0InBhHv3sU/sfB8XNRSV80VOouFD1+2fGfhCyj
cjRTZqKZkeal25b1Mq5IaUyXhopEyC2F0zcX5A/aG3xlzt5zZ54I+gJVhGdHqh4zQLiNuAip887X
+OcSGG9+6NI/geB4U2fxBAdDUXC47PbJN29mhyVcsESvDcOq9rARDtWmtx+8iytW99vxRDiJybhY
PxTLMIR2sXbnQkOPT+1ysaMgTL07f6cyahiW1J5bPQU5jtLTOMjVRHHUBikW9Ltp/arhTlQKCPH1
e/f4fuuU7CSJe20X2FuVAK1u5nvIcKhKfizFce4Mf9xsUFyJMAcYRbIIPUps0iRvHvgC9M5cbWG6
kkFYmx8S3ooX2J9eIqGDYQs4cMVOuXWy57HhQmNzukHhdIN4g1yVRCPtY810C5pNE+TdeS7eMcPk
mV2yK8DLSsR6faIMqNTDU9F6cIRfYPS9g/xuXgyLT9eZyFeVKqramAFWDbsOrrlHN3OGPJT/vj1s
+p20d7fCz08qsda7LDuGHK4nZJjkee6muxKSdDMMAlOGSOO5sGjRjwz08z7pjx0sMYmeMYJTCqNz
T/ufrdJ1DuB/Q3GSnUMeUdkI2Q3R47tkCTfyJFYBEZxrQYZhbaTEGfs3wSEaLyFIv0mYO/3xI/TZ
W/0hVa3RAKqSxVmkOopTUyxrv/glwlCGnxVtVKUiioxT8DCjpF+WrVWAZMRpKfatKLChV4xgA9b6
rgxN5nEE0Sfoa7QNAi8WeCn8J2M58vdGT0ycY7bzNy4gx2HlUgv1AZVDfY1sXkVYDXEyJYMuJrpd
DZBGY3TzwQXQ71Li6Tt6O34JcwNvgURoaKlrAbgEMA0cUAb19TFJ8cAA5gItGGcumy9YCjIEPzP1
+4VBM90RsQwW3bVxHmwTn4ycUA/QVTlxvyr50c3M479sylyqYaTmC460SkQWi2oJEUEZ+E3ehFZW
cPZYFYDbdIsjElnt1XZT+hEp+rCYdTu0pWOhQYJfeUKkP/NuLSuaK+MeLlvXMPwQtvIGZMBp0Gkv
iQx7KhjjEuqDTlVZILXdayBdJnIYtJsxmoTy+6YBMF9GI/jYCpIOchWv19Zm78uDe9du5gcxvha5
CMs1uyHJFqW7CvnnTv1axGcCcUtMWH5pl5cRU87dcoM2PNPh/hfcvE0ac6RJUDl3oqi7CkYXoOUN
+/n5VxTPB2xAjHimzLCUoY9TX/2Spth40ArIerfa+y0gtQw1bTF+gHHCP4v26jtlS6drqSBNKlAa
/wsxYlHcLBxhXyvmqfpGe1b1uEhrvRFYGSd9ppSAbRjTX2bt/cjfeUUsM/wtbir1mcLB0DACqWOU
fd/Tuv/iPNrW8LWycmIjDfOoqB2w6nfomCMygYWGBlJnPGxMRGiyb1dk3CEnOyErf8jXkc+Yw3Io
gmy/WWk/H007K3sJsgDpHTNUDdOEJk09OX/J36X6Xl5TTMWDQpbJpiH5UWEuFKxrdqfKRX5JVYIh
VwjRLOd8Ch8kRo4Ics6Wy+lhPFXe/7S9ErTFgqVGSCawFVbBXkafUP9l9VT3lWiUZD7TdklDgNmM
3U9ayxtwWUIIBN1rMPfVNE87+ZMkWSR5sz2qrv31LMUTj6N4cVkm9Eug+GjY6EAsDMpnzKqe6Qj7
5PY8aynnbrPN4oh92iUzTgxFS3k8GKzODA5zrJPfoXno2KL9h7Edixjh88S2TzaPaoj1tlY7kPPR
x70y2SUTIm8IfMgLdclWL8UbNjyeQm+1edCIaWFU2F2lE/sOyGbRrBMDqnd/4giuN4LYgHT6OTYm
6UkACYBmS0FuFZrIzBhfJTzZDI3RAmeEYDaDSr+Rry1FHTfeAQ4zhuMGqAx9OqgFTsqI7EyotZ7r
Myww7MHNWK+9LZQPEKmmC24M4b1Z4FxYuoc1H5ukC3Z0/c2xVozeZxibs8W+8ppGVsXgXg9+/wLy
AcDph1Eo8Ul/1Lp3148q12EWIM2jEAjdCy9d56YCRnFGl3J7UbZlI+8x4qtV7trn6AGBvMDVI5HX
STz8az0a6qZwikmp6xPGiNXQiVKzwjrUVJzpvAY9pUioE/vusVeXLpZQUQZJZ/+cGBQ/WSjCXJ/8
5jwocN0CCpVMdWEWkwqmyZAo0R2jKJoOlEcg9DP/Dr0iN1EEu6HYkem3MgvEIG46ozxF7DSoDBL9
N9L4t7DW67KMagFJIKebQDVQ9iPnJWIT2cUAyAlwrBBhRwBJo5qzJKYbepeOgkBBFQ88sjnJKHhf
jUIRU3wAw3lhQmyPGv2uyy1vVYTsX2rD/AB/xJyLHTA6DAzF35dPxELIpOijnCfIyo4ojPkjcoVo
7zrgaUWjlTb/U+TJvldoc55CJHDRkXB3kKjz0LAHNO2lmAYmXdu4M/RDJSXPdKoBBTjy/UMkIYPy
q/DH7fRSIAKiaQbnlZ9bW5IGET4200qRXlO/Xm1gP5DsOied76T8i/5Vs2Kao+g/wnX74HtgZIYO
r3MpZ2gs983tOCK9S/kmQZ0J1knx7qXfNB+v3wB4zHbAnoC9smEd1a3ilriyjIfvcs1TrR6aP7Jw
XPYyjEovZipd5yaG9XK7OXi06gCCgmzJXYa1ZVoD501j979a9AW38n9Zhv3OuCyU88VEb6/TrIWz
QejQoQhhguYNQBtGUtGi4XPVe9Kwm01WSfEevxQ5vs8s5wl6sErtgnPrH8lFtq5yH5HIXydz49ld
sIMCzMH3LcEMpiCxzFvo29x5AOm0MI05TrzkgQNBXRSXs+OitFZe7WinxyW9ixwvYuLKhpX1P2qr
ZtbssCFNaTQ89FgzQuZv6dm0vWDAurDdzajC5Batlg05zgNIBl8G+RArTErf27Q+X3UxujA8Q0nK
aoV8CHnkdPTC/2TSZAm/uHmZ7Vnj2aUSi3EWYU+Hp4n0iYUNW8/FQEhpyIEpZU0E389qn+MYwrbi
haVfvRYh2ua/Xyr+zTmTDB8NcHIjBvz3qUhYr2IpgMyk9VqO0XaC/IQZ1DMS2rAXKnfUSE9KdUf1
EihplinzjWjlZkWodY+ZhXYs1Ct1m2zMYNwHY1bM5E6e5DL52QnTJ9BPE5EfDhH3bmiCV3WYEYg1
HkNz2vPbR1i06N3pU/Gx6fnVzIiqoc5yxTxV2PlLtdW5yX1oKiGdCoDdF6y8Ma59fEhgtpEE59Y6
oIUi5kid651DPnLl7uBUL3JNutxG4Q+HNuWNXA8dIFuX7c4vdvzreEUDxbbL4ZAUBhgW7blf8INJ
QoyDFyVF4qExIlteFzNQZbRSe2rvBITJoT7g6n23HnlQm2G0zPL8m9tz5/+m9z1RDpjGA02ehXAk
LZYVGen9dYTvMXPnu/3b2yrGpXYqx9C6JESq5b8XrjMdB7a+e8FID/qMhJIMH7F4dmp0DBLaWh2R
terLKOjdbNmz1k39AFnzS12N0TRcfB4yua0x7QN5EqC5+z/28SjnKO4QTgVtdVE/G8h2Luqwo0VM
7fX/pX9OWoiMo3u5oE2ZEgFnIlwA9I/eturqxtuzo6MEjWCI8IY8AkTUzoTVssQ53SMx/NE4n17+
kqU4eZP3tgk8xfA7dLFmJ0BRF2Y+WD6z44Jm+G5I2Ds9x3B/roxMj7ze442BtiPd6fqjwFrmK6CB
BowaJrtegVzp+v1GswiuM6zPBZ4jDV17vzdxervbmZjL3EBYNgMeP1HG7zIKXpQbMqYAshVb/pLW
brZI+l0QuaQ+1kQswXxaNm+Aewc9FXAWzDN21Cjgka593vJNwedpv8kVNNmtJCzhQuLSW2DKF18/
ii50od56cEUBxZjA1wLVIg/Xxy7wfs0w8AgyrakuV7U7OO7BXBVHcQhWcGjR9gpaM5BSNmmtakWT
sdSfWFloVnyCpFlOsq+qj8eqNRk6pcx5GIfTHBvODTsswG62Kj5G9sl0vdt6aC2B/qMqYPm6B92f
Lz1TIOZGyjC6Xhi77EM49GUByFr2P67M2038QbixmVAODDXolPL5klQfiUlMrHIxFHcPSDRScg8n
YSuMBdsX4uqf9XZgDG5QIHQ7Oa8rt8U7ukbPP14xaRRewKwzJMXgXbjJej+p6zcZXqtGkV5hpPy0
qHFM+Gen/vrzhSyPpsQEI2nHMBScJNDNVuL/GvojozMzUxnlH4RTVlsINShGfDenWLt5ZqO0Rupa
9umsoNdvhWgSzc/qiOBQ1Dk3Ak+Jp3S2xSUMXikOg3hSOWJJmp89EbLH8JCaLHB84But8ekjQAVl
oUKTOnVXcXfu3S5S5jJAJLiM+vDontcspVsoF/doqFW/oTM02LRaeZn9U/TDOWh+t0SjEk11w/vJ
mvGnXW+fpz0Es5SzHXgEgl6PT1lfkSe8Vc5uPCrTCB53LJf0o1idOTyN92FVyJ/TXvoL6xgBMWjS
jh/YwLzrkCaeEg3GVgQT6uf1DhtRId9GfJOhwoMAdDAclDNU9s4AL738q3ZjptCs4eT1TxgWTnJ+
gVy96q6vNGDi+i7rtSpVbRRg/e9PwJAxq2V6X4fEA5fBMQhLFssCCQg0iviAXXMY39J+YkJIQzD7
OtRy+yHnl2EyCZHFflEWmL1ess5YJM9viQrkEKcLjyJXe521PzfIZvb7cbi5Tqi8j8p7thTkwfXQ
NYYS8/NrDECzuWFSKSvycYbBa30g1MH+3Ipygx+J43mDruGKnjrdJ3Wz7tjBxJZF+m1vBGVqk6PK
Df87kB+2EunpFwbZd9t7V82BalFOxdNODNgfPbMpSL8ICDG7LLomYY1fnGGT1nijZaA8D2t1nzkk
M8OnodHS8XJ7mWVuMd+d91tBdVVitB01g/n+q5+4WryD8/yqswx1vmhCIX13shifQWpm3CyCXiqh
RUesBj2PkC/vviDS0sbCovtJnqaQQJU1a5D/PTqqJx95hZ8nL1SURpfOOu8nCn98XtIiRxOjB/Xh
hKvgXDy4IQ91i97HD/80jLAwnk6GV+iHsNw7OEEb/KoMvW1UwNda/Csfw4XPan1/JwMkXCHxR6Vv
j0ETTPMuYWAFO2k1esSfb8hCGkW5OUQdmICZtuJ27vptSULAvWkDkUD1eoEPaubRfgF/vNoxwYGn
fmU+vdm6jcs1aEAr93g1fqfnoGAZaUD9vLQJnuc8S2XjoBifdOTuefMQMJNYQ8sL6BBFcJn9vRms
5advkuuNWhA/ZJ2snxyK/jZfdV2Iwxe0IZ3kBFN01+ymS5tbrB2c4WDdinU9V2I+vyOWkuzgl4A7
4eU8lDOouvC5rWnqPZOosHW4CnOn8zufs6t8WHVzP67dPcx1i5Dlfsx7nMfKklsJbLdk5fKBvqOx
Nup1e1sij+vSI2KPG+/J+b8WSEyW71miXAFD93pbUAQShm2OrkbPKA9xxAjBkSljjEoAIcluMd9U
yQlPn7ajKXnm65z/HQmvVVzWTrnBhoXw4i87eDfHxFXkk4utkqj1yYTMrQP0n+AqBkV5bVuKDz6d
TTq/+3QDZRmTdAjqWapJ9/rbLlxD54Y1g6w2id8F9kh75HArO/RNFqBtdYEaumRq6kOfDGy3tOCU
CfMTg/h6OctCF/O41u+Q7dHNyVSFvID4m3CcILpgkGDmHXmMXoB3aio3CQZX+2QucNA6eGKgFZTO
jSPCxoOB69nYi7Vdnbo18Yup6IyMis1mrFab5yAqLDzeKnQWOdpd2Pmz4gFfHIa83xs++yOnXKpY
LzK5OX/1VNCNwlLh2TUN7XzJJ+/dM2D2jcQuLzFKeTVcDp5uaE5RK1ZihkHw3lqur3X0dZEr7d+/
XrxpQFJpvc79PwEulfp/9pfNj4N/ko0rQ/HH0iJ9WSjIQZm2et4hwu5PBdJHe7DmQQklK5haMwQZ
nUoi376lZTqTbZkWCzGE67Kk+0upKFiiFOMo7XFPlqx/UUDGfA//GmXWjRX4mB1eh2iR+dU2vCIr
70PZciumSU0lrYn5eZCcHJG88mj8eHCW5dM/I4fVX3tv2k+vjUb77l4scb2HqGafD9bJNiMGoaQG
yj+owkrRIfmBxDRw+0tO6Jpml4Xa3RQHIv9bWFDeJzmfebUZMrDr/haTPJs8r0KyI3dmSyn/O5HS
UcVa23Xmuo387hHaGk8qEzQXfsXbByUFAXk1w/Jru6+su5I5e8nR6a3tz/5+yNeupcKOCnIbNkBb
hq7Av3zwHpYUZWSR7E5tVyqaL2UOA00f/4tKq4oirvW0XGSwDpW30NUMH50ZCP2oKo9IUoOGlfHo
jJk5d/NVhh8YyGgtY7dXfykJlonSYG8VQuDTsIKj3lDoqPzQG9rfxPKf2uIKjOmMK1neDgLQ+xPD
Bx/gT2+S1QgFUVsmUs/etTJM8P6ZB42eDHXifndl3oCYN11NJBu8FnbIP13quZITDMAZGk2GMF2r
MlxdUvtCDjumzf0mC00epty4r/ra/eDVGH/eX4/TKwylogG5Dnmg+cfbNlZFnTwR3jDLbHW/7PxY
Ih4fSyU6pz9T2cem+6iayWfSRsaN8Ebxua+TPaO+CNfUwaSQANT6pdIL0xRxSoSsq83Fnh9PX+u6
s7hOZ3nhrucBUPdXP7/ux34K6+sF0Z7EeQSFcwGCN7vDaahhOIStDHTLvVa5S1MSikUR4NKnlmQ9
+7Sui32cFhb9MfBd9lPyRVrvgizS4wJuUxZUiq4OM3rWOqRMQi4dSq8DqyjSjRVsZ6MH3+uEDaht
WA23gkqZz1AQ8p0ED/zXXN9Q0Cm+hicwkFoSBS7p8Acz9s7xUB3mljGl/sQ+7/140DuAc2lK6zkF
9bm/L5ri14qBdZh9J9FwEJOiprKgTdc3mWNH4EW8YKYifGf1QMK9+5lasvl2aPUe5vy5kt4049EF
QihX60wHLZ6K8h9av1KXtlFc/vnv9OjpPwJ+1klu6kvQv4cPwE1QPCWvARvdZ/MpQsOgFVTr/ypC
onLwBjZVtOX3L/+r8nLUKUqmIhE9XC93TcTA0ywWVNBe1/PcGW34HombX3S/qSpEpcxyImBrlTEA
OlaoDGMSh3quNSNGkhGu2I5al58y8SUZjECEU7jh2EI7ZC6uKWlQNciOjAMM+bKdOV2O/5/lUOpD
k6BwvUYi4jvETOH0C/sQ2YDxrg0VL+RRX+1mIvpfG8Lmf1FRGgbSayiC3rm1g/cZ8QOzhOhnv7NH
ISKPYUpkmLeSgZWOvmtQBOAuE+jNrH7G59CIVk/EjLXjgS88SPg2Asp60dPXNKBhlNYQvvSeaUIi
vyvE/2hspBUkjyO7LMQRcCFAhJryGpBmMJDxTJBtY/fm1K3sZQ/u5sT/x9SjMs/99TwuFOz4gc+p
jq8/05TE4ugK/3/ENaea41XL/cKG1qNz/Ixz6Oqap7HbMEP+ToUuHhwtMeVLMel4oyMlGLKUZ1Ko
OL0LNzZWc1czGwgpXlLjBMYuRgnaQxy+r+HLJRpfWRoTSd1b8HzmbH9Dp6bH188O0QxKrkZZQBKX
NaMnRrVJXFgnU5DV3PEd5Yqext5V8vQYQ6wqc36YrNeRPx93/wgypZgU85w0hkpNU2IOR4iBg96J
wxyBwwXwliD0xe00DwMstYhERukvA5AE+FVNY3+VlZcaN/XyK2XeZVjMhF+ne59GQ3nbSXC8neAm
oz2OkqwFtQ3yHrRogmUnRgnMYGz9V9229Vnh+L7XasrcK8u0/JrFDNK6Zl59upNraYJdNtPDEzxD
c3PYNIB3E6Nrhqkz7VzFLlUekm9mdc+1dc8Zs+Iglhw6cJlAyVE8QTqIuImgEO95bxZ7c07jjgEd
Mfx15Tjlu5wdnCDj8SmnDK7zsDMTPAhVBYTVGU1RPCPIIpSJ2QlkbLLWxKj6uBjfy/lNos37/b6K
WA5AjGb8OJhejmfMPA8RcYaUq1gGVe9mMs2UWGls4Ien4/dUS8FsEWA04SYKqt1+B05C+UZzeq9a
HXn/uph8YW3WiEpHn8zZ4+jk4ATTEiYqAfFYHc11v7dm/Ury+upGsXDSbIB+Ah7V5MDKF2F/Wxjy
CYfeRwrjhYav4Eaux1KTjRSgC9hmJJ5XYxjdVY3/xoi5blWuYjvwYlCn8hHVieZj8Ovh8wP+ifq9
JuT/wmPKp//lBPhoASaxLC6wD7V2TgNOVgCUATNsqwROTqaZwYvvWjOW+lIMDxZ1T7DED0W5d+As
cg3O+iiCnfV2Rh25rkMfwIyqxleMj+g2IznERpfO3tadZdZ924NzclKrU3lP3/3ZG7Ng+9LWQ+r2
F70HPcizAATLzc6KXBtXB+PtEFLb4750Skj2m+/Be8Wu1ntHI+G+OmBHo0fgJOxLAdYzBuU0+RCG
FoN1RgAE7SN+gLPSiDnjHfmox+jw3RtQM2HNcukHp/Ft1pPyNv3rPEU0hs5UIeZd+CHwUI2aD59d
O847Kd/883eXp6OECXjwjJbDVx+vWDnXeGAJJQzpOrur8UQ941xQcCCChaJ/kVfOPn/GrfaJkqGc
zcEksxBaH6F5nv9TwLD8O54HHOpv8gTkibzrIehrXZpNYVLl2TkRD1gZ3iemGf/fSVP370c0kiFN
ghKWgQbOQFQjRsk4rRZ7PGwwR6+D8ck2ku5o2yM+HWqvR2HNjlO69oK5C11tcuBs2adTs3w3o5q5
1nOVZy7RwrWiJJwlCnPbDmKUZGMiMqNPc0DMI0CnEMVgOC/r95YX27NuYAG+dmnB0Kd9x3OqCX7M
hYFcDOzm5D+KRSotYTc9Lk9+Z2ZRvmP13p5FS3buNcgx1XGfXhq12QcRVI/stQHfp6Xc2AV3of5+
jBkCzymhZDc68KQDE6ooBwnci0mgssmyuUwPUBbPg23gY8gyigIuAyN3JRZvjUV4srjUGAPsuCuF
Lw+OSaDlEq3YGMkr2kbRMoAL3sIsaE531jao79DPLwqNLHeFgQjiWheiu1Z39B+0L+MT7JBNA7Fi
/8XFzaQKQDP0JLFgqQ6wrYm/oKS3e1uIiUeIL1RGryhxcYS2mPQNjDsLCME+t2pLgt3JEDrDLUxv
StXphZsiLX+ep/EKSQIxGOAIOGDtUjsrQCfjzQ3roJNcauU+b1lzW5fE/tFeF8BemapzG/ISwbbK
Awzr+VnfCIayFMYeiR2hwpoi2TBVk4ma4jBMNWEhxHKUZ4rUUm+1fNTDfpj5IzzCmYzcPCaHseWc
2mwjb7wqqNkn6RjDhG6DuxvTN7ZXuIb2cLFMW7WDShWSZOWUA6QxtGRHe16zVvL1m4AA8uv3yYK7
pMzVxfxwcxR35ZmKGx1sfZDzW4N9X4pytNNzZx239GErPEFzMTnuafl2dum3f4yL+ykAV/z9tXnf
JZqu3S9i1YRlZ6JnyYg3Ot7inrbbLmqz8CQW36lmbpEGpMasuXlzOAwISsQU+wYZBCKM5NKzrf/b
46WparBrZEigRgg1QBvdxaQ0eiB9rvyHp+DnqgzFNpwHH2pGfD1B1taWkF3LN+e7LYUfKuQLAO/K
oHPfemfWI+ML1lEj3J9naNu2G5w3Yem/0E6HzbEUgv173tC5APgGJrgFCuW//SohXxZjmbB8aQbo
4bJ0FnCbXhXARf9R5qScSWgCnadoyJnMZ2EO2aYQd/lV7b1cQvZKgbxku17TzfPF0peEMTnApisS
/igeuCdpE039Wd5XsWrB3GeYslDu6vDqwCVHzRjwPp4bcmM//MkwNS68c2ZqJTN9FUo4hfm79VAf
/qpO/gcwji2pvtRlv7AHgkPzT/SVDTeR/JgBHIX6DmSkjKqyp/9kl78u83JFmmAJJso3rtCEbc1L
V5eZ5GkxKY5Kc5WEg+RtMeGRkFsdq0ztJ0SsmNtpurgY7k5tGCsBYCCvVw0L8sY3U2HZ4vb6b4NJ
QkWZN3dcodNA5GAdKez0Oq81SjcOeliVyLthIa/15SuQDBmSP/DHo2PPrGtORQc69JgjVCKNnPkT
YtTxyEcDcGXHc8sjePBUJ5/S3j81WOwsvsCLlW4HXgBr0qmtmcFgbSG5DYjDBgWWjy6ERhmBrnIK
Xnxomt2dwrAZHBeqtjuXDKvp+R35cwWDsoIr6pDItHWqMSWmqZvEF8XcMxzf65+cPRZ771PSkqEi
I7R6GSrsxMVKQlSRjHeOVVo9+h8Y2drfAtXKKjFYV5wSbLN2UVC3Nvva1gHyKEAco0Q7Y6L4C24l
0g5uIJKCjcIgCAvHXXrP8Nc4RD+NIVB+GUCNcrQzfiLspb0GQiu9mIN8rMkofxMumrosgYmodNdL
YLbrHkzs3IY6/tZyBZQN2RMJh3ic0AYf1FyY1Ft3KAWKSpGTyYHHV6Lj2YZWOPV1wJ7FouDESq0m
j1nETQY2prJ+LrzGvfY7yJNysavH0EHPPcW1QNnWgK94xgff3EfGLk+lK2gaJxZbhA6NTI/hW79K
RTLxAhS+JWoWD9guECtja+M7vA9PKceSophC3FoHDlsqRiWlxeaGk5NGpt0koP5tzoaJ9+H4E9Vq
4hdzR5BCEM3o4L3f8ZasTqFN/p6PNE4JnK0iUgIQnOFXAudH4dOxtaA1xHdba5AY7XaCn2NK8xv3
1zI3v5eeuXoIgtOhF1t3PMGa1WFT7LOISCDfwiAQnPNKsPm6K12sIKiGmYmpYQs82W8mSOoeBZAW
CXYPPpRLIV16xT4hwwtz+b3WCdznGrOMNQkFeqZV3n47MKUlcMscqHeWx04261O+ldRpGOA65+9E
162Xg+JVI/aKG44IPpo+sp1ZfOhTn++rCDwFn+cT5NM/568CqD3etnB6DMtbr38eYUkD45bzDLmy
skqMeDgDycsuLxcMxUSXrYwJhZ6NGPzSSyknHjM6prYN5HogZy5D8mjo08vKfS0xUdFmMX+ST9LV
5zcLQlkejiD3ZtFH2vCTFXUYlKtfa45z1MA+xZL5jK0oET1PSkzRRfIlRVH0DJv30B+HH3rN0Sgp
oox48cCp97Vn7A+TNGGw798PnPOgCGKR5mJYtTjwjJ0ZAwnorkS+Y8n+nipy+HVxQ9xHyxQuD0mb
XODWxaAryqTIwXpNjCULlSIpjBEKCJCwHYDovHBzd1uHaJeGoYV2KsjwNCXIy1OpzmO/XOrNxwkg
Sv2JqB5UKTXzmlUu7HYbqXjM6T2NG2c9IgwYcwwXxOZ2JrpdqsBn/PKvK+qqVr1JCcub3EKTOcO1
dDL64lvkQqBmAZuY1YmQPzR5+Yihv1Jd2SvQO83w8O5UahEXT3/3fEHaOvoI3FNqFI3Lrl+LebWB
5hFIg1mPvbJaGpQdot1dARQSy/BGO+edFFtzTZJCy1MparkZa34xemhPNr1kcmPoIkNQkVglVlxD
q3lgI8A8tQRzaVeJPJq4wGFLCJ0oUI5ApqVj8TYAAel2sFtISr4pOqUV+3OmceSEDFylMd3VmmVv
bz1eq0o8afbSmKvq8guMxVaadyiJGwvb7LHX+9gOJrAv5oUkrWTiddbsCS4QnlVWoRJnktG8duxH
noyVlymcyFy4CakhVeN/lP+k5u+au/sizLVZsXeb5j8qCaynwQd5qFley5h0N4Vwg/0Q4sit2AAE
QaKR4/DJpVNIuXxNSsojY8+ssOMCsLTuEPizEadCCPeT2uGFYg17nz/O4hVWLQ1RftN5pjFpHZ9G
9BA2k+xJtsHB+mT7ldEf1Ud5F0YRurz3a4+s0UOgxAY5JgUHGKTYyiUceinKB9QRkUE7Qh2xozTc
pyIve+zTIDOF+2rAZj9mOSuc+BtoCUr74/Q30aZBI35eavFJvxxegFA5ZJCfMQrEG6oadpfNOzz4
HYqkjw/9g5DOBcVx0fZspJZESZEzH5R/RYJo44Jx8oZi3IxJNTtJXSteGG7EDw0xjDpsa8eWvO1O
qSYeInYWIn+wXwObfmJiwvz+Ocx8f53+eiUGaMBsE5UU/xArJmbcoL/1OOqkOmdwS86o3lLAtRxC
XV9v+mj4jNgVdJjQuvWO2zKOB3Xa5GeGScETsq4I4/WQqdFj+6c1vjxLtNaL8lDHZ66ZCUTKSa9M
k8yh6GQ8OhvE1UyeAuW5Pk+Odsnj08Kodk9PHqgcdOQMzIxKAEnAmdqyT3H5uGRrGJk4qt0V85ec
ejpnvVSpQZ8JfDsU76eD24hXh39uIs9wbyqRafuZSIV52Zd6r0fnWElj27C8vuBNOiwpy06xSBin
8rbg5XTv0VdTi1K1H2H+xEDvVDkmeByeTg9zYBPG9wh8n6x/Ww87mKFxj+6mhXQ479izO3+gbk+V
BVjk5XSZaxB0Wnvf7bfE6IN00u7Q7/LPa2ihdBJUZoNy/PsC+nW0cvGlhqS5loO/xZ9kyJ2iFlg5
8qRTNT5rlyulnmD6pjx6kfITXRpSz5jrnEtaRS/uQ92Jn7pGTgslEspVNG/wk20+JYPfhgDMM4xD
TlT2w0Nsff0eObM2rVxxqpipW51B/IaKDqIMUfEZsBk/PqeuwbINIQpswkGVh5PsJizcfSFqbzl9
DRf6Tp8cprbWhuGbrBbO75qAiI24HeQZpsGrOv94wgpONww7/oAAnEf1KSP/DrCuey/P1f9EDat+
5YixgqvipHeT0KMAv1xp4G0mqaxIFytXBVQINrW5maPXQ9/xht4QdYDqTWnUziIB35fcSfMvVboq
9ikOiWo3e/k0J1Re0gjbnBFaoODh11dyPvZH5me+Sxne57KulqMTgNWHrpa7r8de03zXHh11UATG
XX4yPcs1hl37HBPMLQxOdGNiqQ2mwFBOjn1284zNNJCUTKEMV/cToqQOa5AklQY+qDxo28W64lgF
V+ZAYzjatDQObSUNBcUm4GyZ4eVgmK8mr0K3z4hFeMI5oHVkCG/Yz6+0MjWSQT4zOaO/wnbOSDsg
edOAaHXbAZt8ogrQty1fLdT5AwXOmYZD4ZuDSJitrh1HVH2HGWneGoXp+uFMC6Mixn3hLWtEZpCg
hTpy6r++EIj+kM/WTWElv6xThCg+0XvyXPIou0nS4xX5O8ee4RKHg1bCZB6yqH/TnCasLaIpBj+q
fM7I6BiV58psO7X4f/dNWAC/rX8wByjOn9jyapw5QNHFQytzsPprQjCwNo77NQ1qvXhSVzAUDVxV
Lih5NOkw05VjPOemQnNBeimTvoc6eEoS+H1S52UcKcqYkdRoilHEX31650K/iNhnDBA6tOXFj3Q2
h+WTQ1Ej5/gAG/wT/Z8PrXTnmqZaNoBxr69Cvpf/kXAfjNXm/qKT4TmhETucUX960YDxd3e13k94
mL140gBirf6XcVc8brhwqzw0SCQx5Ap+oWjjESZWJ22+MC6feke7Tr6bCnq7SgWyOkcarxZn3vK3
K5CmPIyyq85eP+DG6oPwyrY7Ahd+Sj2x9JD0rAf3Th/JHszfd7OWdi22psQ324/uqYg8JohLMhYI
rg6YDEc0hOb9nPm6RAvkf9xeT7+xB9gJoJ7OqIRPmEYcnXrLsDE10+fOPFs9NlqW5S2KRvhao86R
Vjv0NG/t6gK/1Z0gdNDBuUEaFvTE8DpNL/RYM+iojp4E7TZkaBmsLpaUqWqb91AMu0TonSeNc0xi
/fLxGf8wNhnju9aFQgbUPfioseO4PiMwN2eJSPoIPapgn4EixOxC+f5Pu33BI20vCedynmONszot
fzeEGhFY4Jx3lOOignR6FdsFYVXwiPyxiuVtbHPTiD0AWG3scIlYjy6UOQugGDCkjY3t6FbVIdHX
RLxvecgNsNMRUSUviAJmMMaQ1nGG8rzgiJXHZj1WaTZ95vJjWVSIdGO6fxmN+epP2mpLPpwrfWvH
+f8n2QnIoExpD55snmmHFlvil6b3jJZml1RJgmwfz/5GVgM18nyARt+2W7Ff3RMkSmy44JDXUkdC
CS0G+YEj1PXtRZ1ZAZZr8VMLJbPqKJEniLkTvjaCYSlcmDxR6HvqC9K+pAy19vTeV+p0iZuDNeYW
CndpaL9lE/NXFpv89JK5AB5XhLAz/s3KJh3g7BHopXoq6mVzM15JLGTaNKFswE0koMwt60xSwbp1
ohn45nGclO1QPYtnPpuBSLXtdqS1sgQ5ILUXzQrJx1IZMIp+I58JxoHlsSd2hspl9lEpvOdNddI6
4xKbky/4qtrvdHr+xyooDChVxJVLx4l5LGphPz4bZX6s4RtZaYdh9t0hcaX/84o283jRb/j6tz++
+Q61MKxQRjfsfHx3X9HRk76DlBluGplYI5phBDINDs3jeQcds2ZGXE2J6koiQSxu3ympVXztngaS
PwwcHrQU+cWJAlM4tAgrkm9sc41K1jCe2nWf21HvZtduLTEqX4KXxtl+ag4aQkGecMX+FNTTryJy
CAEKAsdhxfXBII/J8iL3be+NKYYt34Vl/zWSXdg7Ti8fMVMhQNP/oTukf9CJJ9ZzAQIX01FmCbi1
mxQlNR9QCiCNAXHEqj+H9IfZURYcj1RV98sV3cY7ZdtHIW6xQ/T8M+Yg4EF4v/Ri9vKspsDmOxsN
IV/UGhZ7ojMiK9Oh92vcZFyTgpe1hnA1s94vPPZo7p66jXtK/vXvq347l4Uu0B7Yf5Wm3qrFvUfq
03ESHMNu0Sf6YFL+PsvabS0T/0PC5PZFnvt2PEIN77nNqyjvkKtKblLEsZOSv64J0UxDb9Ym5DhH
oj5lXlW65mlMKdzfJcDwZkl1obgw6Hh7Wmc/nZxYdad7u25Vs53uWegfA+jTZFpq0KTQnrSkv1iX
JQPhhh5Hmg+OXGoPr0nqhrjb1jwjK+noiE7VwiFKWF6qyfzsl+FVuL6xF7lXxs2ux/RfhOy+REcD
hkoJE1tKgpJ9rDqEC0F+siALjwx2yZLyeeuRLABhN7RNXKRnkwJD2HkU1NXk2OJEuQ7UOTtA0QyS
22vdcTphgglo8rPxMZzih9XGEYIzexvDVwSYA6CuA2ENsvxphfzKbZLFGXFgkKnAb5HsEbBDmAAx
O4ZLgfvBJ502VsA2Nuio9TF96rIkrgQA5T/nvpeFywYPlc7/ONuCCdJHDcy91G+ERyntQkMAK5zd
gp/O94528DphaqTgM4ljhywTyP/baN4LR37SJPx66UypLDuuCjI1Nyj440woLsxYYPsbM9PowODe
t43lHgg5iSpEBN27ON7IT7xi7JiQr9RqFG6iVeFQ9z1G9GZQI9WzRXPv9Rf8V1K6NasQhB2UQaw5
xOXf1Zdlt09r/60IxEl8IVxX/HaNvdaPnwSZg0s8MMh0sjCVMTvyV5f7osj9uRzcCtwluNPUVB46
A1z9CE9NPT/aop1iq6ah8bzeOS5OQf3TVw++tgnOCDftULQmm9TII88dKl5OhOEQBGZduEAgp288
Z90bdFwW1DpevA1IkpN+hh92NLCeqF5ZiqLF0/ZnSLackIgDFxoO5a00RPo8n6LGvT4sdRSBktLz
mXxDvtT99Pt6ugS0B7VtLUNVD+HAmyxt0OQFepCUrCjMLR9PrmZRcChbO72huRGmBf5Wf+CnIMkq
aQgrvOuFzIxu/VZgRK6Q2eBstT+saL+FNXrFHQSOURPCVl0hlSBkx9Xly628GWJW62oP6oVPKGXf
rKQCYShvAuMOkubNm4MmQ0V9EHm/+8vr8wmNz2i8PZHa9KKTl2l71mbM2a3sz7sZuFW+OpJe28Mn
wr1u4OL09J5zisossrQznGq8FtCCD/lgb7bXaR9QpmADRrieGlTrjjTiD0dOdY5B0ePPWuu5Le43
9RJOFqmAfay0ct3IkOTCQhx+zDcfAV6dZT3VZyr1wiRdLrvd7pOkGUw1iSgcV5Wkoac/LAZli35I
KE3qLVvQHHAeeOi9BGwa1y8zwkSRxdRsfqkXenqitq0PV/cH3J1SnzlvqNQdwk6rg0N5waE7m6wz
SJGoXbgU6/T1aFaQ7l4XDGduqOGrxUTXj1rLwNbMPf55fBeqbcsawSQBjkcNzj2Fnoz7ttihUwEL
7317Fi+fHWe65+lG9Saow21AsiARdWSx3n1ykv5VztHH3N0igBHuIROoqMlLxzNREwK+oQT8YnAW
NcWKP/1wzj3O9sIP1iMQURt8P6JuusFkoTRxsvoM69gv4JH7jBcQYRFRSS+C5fybsMaDG4HofAva
NUokwTeIhTgBIlIMYSaCjlSquXIwl5anRRXpUVORy7YTFGMWSzYlAn/siJgpj9Az/wvL+mDILuDA
kEYdkjx1Dt54a3NKpKBwJWOBXn2DGMshMaDr91PvizDXa+igXtA5MH32HvFJNMBvio3rV7T3rPRt
F6Zbyo06ulqwXjsS0OU8K2WtvWY9JmqpaJY0n5BbhhVlLJ5Cr7Wrok0vE6o0/W4dUi6aq5qJEQZ2
bvjCDuXSYh2JlNtdmp71Na3ZbWVCryE/ZbPZZxlRzMWV9kbmrsGn8XeQpJVTGQiYDU6kaV/sLoVZ
gX5rsHJgqT80yzXHjg6nDfoUssCCwWmuxf8XC10OwgAPLgOF14BuffM6e6oLVe60QQGF8YKz35Gi
wIy9fnrilQoH3iUuynhg1dDdYwnNU+nG+eTZMJw2fx509r5PQNcT2tOZlfFOc3acFpVMiYDTgT0O
718G+Z8v9V63GC0mc+czrGs9I7994SKLYpkjhFzPzdvx3tLHv07IqH2YliKnFNVqhkGiTh1DyB7z
S2zGkyYoUSA1pVEekS7K9SejfH0FzzLqIG5aYXCBeWr0Dg815VdtBdPoXTMP+OSv+Mw+s3D9TuuH
qs8G5NgfxtDtldH1kdpi5U4/dOVTSdfQm/d+kjnqK31XXT3v4SQCZ+NuttIWCoKCINHjcBJ5KILy
kz+FHQMZEYTPbo6nXlkkpwPwhmtbRIT83+WAAm2pnTaIlZi4T4ic4+snXg5laqOqJ16kIG3KnVSs
ojOZ0bXs/u8xI/bxwEoS8uWnkt6nbuFExtvl8bHbek8X7HU/cYRFcVLdpCkm0Uvr/ZlD3ZLr93XZ
h91oMRctT1psKCw/0kNEQyG74IzEUdqriY5cmKZBFXSvEELuyOZfFK+ZD5hKscp4TbmiB1SGwAje
xvF2w+67U5frw1xze+x6fVGUvxDk+gFxI1V2E02gJweKR0ZPNItvha2LrJvsbICVVJlp0C0ZiBbF
V+54SmSjBBzM9xXQFzEhPD68CwhBjto8tR+b6Ys8QUm5c/Rev2Y8+3oz2JnBra4QVpZAeJTl9YBQ
7YMikZNt+YBRtLAAlOWiw94P0/wd7tVLWI/xGDeIfMjsz/tiHR1+TXMhmfWNkHzoJ5ixVeLwkO+D
D+w4xgPqfu2mdReTIYmoYECXF3UbkQHgqbqWJEaKedXzsORQt/0EvvSrucwRCdEUC3lVNIOkDNav
FxNaH3KVz63XO4mtPZsPwLwYT3PiSev4KXZSDLGaFSJZc5s/AuWwFAoGBq2xGO5rfWheMWOPAyh0
HVl4vUUJW0UjvH5io0ehs90jj+aL65HZt3D0pOtaJi9m0WtwFXneXJK4p/XyKfP3rgitxjtT/T8e
Pt2NkycriBmOfa2DopZbqRDiQRhJuhU78Ida7nT2DFDLaVnhsP6QXDba7yCdO3cNemBDWv+S/iOR
UgfwxTW9EZVDN/NlnJxlyR92IWhQgWQP4l4f+Jaki32m+98klz0StL4kbJAIqM+3KhTl6PAIeLLg
k/7zVExnwXtXqMTzfuLV/HB19DFVUJOw4ANZbjUKHhBjIXzm5QRijKUegveJun9/o//7k108Y08k
OosT2qc4C6n7FO6DB+9Gs4sE05Pdv8y+zTCDM63d+2OjdtXFq0O57xgEHn4gV0w7WBquJ+POsQAw
Zv880x5P8uMN3iFqQBAeHjC5d/San2tm6W235Qu/ckbMnT342a24OppBuDBzT8+kdxBak+ExS80p
flOzrbKVvcOQqUsnIo0wXsNdKcr+oyNb/UwvagL4EM9aUzLR/JtwpTS48h4m01Kp8Ie5orBmKNQz
1UVzZu4zmhs9dc7Q/1WXnUqSsKkPVNSxAFR/jFQD087d6gYHQD/mpDAkwPp6rLaAhnvyHjXCt66C
UN2Dei0yyuJsyUQ69wNINbH99CnPZveBAP0pYFm/Zz6FBtxkuHK2eJ4rWcfE3+h9S2PqYLZ22Ufz
qlT9xD6AJEfl3zSMHjeynGNCPK9JefSIR7u3suKMwQoRRQInthRFd8UGlVKrHhlAljTDdB6/bREi
UZ35hSyIFmenXs0oiw387Lm3K/YJIPBYipCVJLch5FTBaRLHtlIW28P/oSpD7hR31tCNKsSTYWUu
BoVcJBZ7DBUoK09nHzBisU1QzrkddCdb1BmVOU2Lh9WD9ii6oGj8Dy+58qEbkQPLbVj3bYow48yL
sO5/pnVjX/CgxuIpa8Apg00FBzAsCzDfRaiXgb9QtIQs7j8SeiXrrFWXyxVQVEwwgCyqbffurxrg
zb2ehi18/i+dzWrMx/hm95UoH2ksqWdNnjz/G6oWcWfCgURelxxXlaY6+L4pcSOif8gaHHWYBo6h
vU2A/fWWVkx8hfW2kGKnFeI7Uf2MwHxgDkJfi6YvC1Q/TBm9iWIFZAzJYwZZ9u0o0QnuZaZ6njNL
ZvFqoLllBsgxakfKVz2m2u5aidY8QjnJBx5cQ0U7vbwFb2ZU58ylE1dFUwbGLdVkPjFDSMhLgrM3
csBYTfPLj9muzfup1UclqZCyviUJbGPSpF4OusHYj0/wLh9DBXEL5mXBGyHfpA7PA+m/B2IHXWZ5
IxZIGlJ4UeblhkreZqYhbXFOYVTWQ58X602ftW4qpVeZNPtyAqcu+igVl7EWdrSeOn6+bbzNcKav
0qN6mZQNtMrTavCp+PHOOcH9jA0yXEI3zwOhQ5PtqchDxp9gNgNC8QjLs77H3pkRYO7+eEwb477f
9shuXYoWr3Hy4uy50I1CvraMvS0ikQlW6DjO/xoxvoPfyWgIUzHd1+5tWr/FhtSif5WUpnGw6wQ0
1IESO3pyHzqvFahAvDK2xcVJ9dut64DMBGx+z/J1eib0NcQuVsPZgkOSSvbPCb71C5O1XyGFGcDG
q+lxsKYJ3IOxbcqIXNTfvSUYY69L4VAQahcxTJSjPkWlQKHLtqF2DaCrnye1Jhf71r/5ACXJTgSB
Px86EP/CizT9Z3H9LyTLs9PPxbVXEy49M7xDFho/GzCmWy+yz3FOUHJ8KKsz6QB8pFQbgF8BInzF
3HPWvlrzikcy0/K2pXj2OfDEgCNDOAsvc95kB1c+2oq4GOnvGzHxwokUEIBE8Ex1SvI2k8ux4U+z
Oq/7J4que/qv6cYBmXWD8ocSYIBfASL/vVaN9aQGgOwlT4ECxrdTKjKbhQWhYY8PeWxJWkstflhm
1BznFi0I49QYZP/QSAnBWDVzrOk6RdigUhEvGzmxWrJTripYFDNGmlfTLt6pWhNgyB3JN/8pAve9
iLN5i5tKTKTrobz1ZzxDFo8rNUO2T+NdkiwpF5SYCSGBgSy7Qxw9gOR6r8VQlsROvePaSdbeLP7r
xTKwnqgdd78QD00n37kP7db2pG2Bb8wc9vXj0+eYSkiF41Nw3rwrpsI8HRAgTiKW+rvKTihEnOFE
torBIOXUaxtCMh89OZN9eOAU1t5YgPzfJIhfDoBNj7mtZSkeeVElPHM68oqE/MJ6+ZHwfaoimtxD
5XAKm0e8LwzniVRUyl0ITH/xbRXYfDk4/Q1G6hRjkFAvAnBT95wV9Zxp1DOHZ96NbQ/jOexMwtl3
zqvmusI3EOm4WgfMey0Lm/VV0QxNXisWUI6A7Huwn1EoWeVlY/9L+/Vc3SkyFnCju6461yvdN5Zb
V6ZJThpc0RoilXTEGBD1RNCHQ8gK2gUBD71nX6zSF91yk5whFeWnTBBbvRZBVnBTtCKbgkecSfc1
OX+IzDWO41IkL7MtaY25j1nVct68tKMgpBXFmImhJB+Bzopt1zZGtoeYuyK73/g5jpjKfJA+k/PJ
/rasJmDQ4if6+NGW4FFzZEyYWRoI0gdin91HFI/rOhQpvdgjCuvZCQeHGiGQcJQr8bzxA41hCVCO
ivrkGIEfB62wi4xm/j775dEujip8wuC65YVdHmBgBQovDBc+dfvc4W6Sd8xUsKDFZDe07J050NBD
ms2sO5V8D5uNVhrq/0DmnmIyxXb38tRi4yUQRUM/UGWOMfMhh25ZQxpFqz98ktOvRU1I4hgLpK+k
XQKpkxRAXr/Jra3wKi5Ggnn0ctiZt/sx273SrXeF/9E7kt+J6WicwdKhhTCBwpDA1LVfHtGguBxU
mnZpz1wu/8Am9dETf3klcycgicjCOma98m0cpqmll7DNcOzVCsq0BAJ7bM5S07b8CRhgQT8z6DIj
1HBaXZ45gFGtiWpFF4ZdrAy9zE1sMFZrPUDpUswxtSpWxErcQsmQZ0ADhA/9X/YpeJygH9OBGfH2
ErGJNdtzDFoAT28ISYwW0JB7EfoJy5ssvPM0MOz2ihJnlpHFdcK/qMj/9pVJ3/6N69i8wrxNkz3S
2OeJkwNRr4rgziNRvNDryYD8kJnb41nL+++WUhkK9+82UK9/IaCKng68cM/iqMlmbspBpYfQJ6Lj
2KcBUDGQLrTJJF6+fIcY53Vc0AiIIhmqSqcVwdzX7db37S8MRNl62KEKZoB2apB+R/xiOZDundwD
FrTBAo4/3MQuZyjsdG2f9Bfk1slVNpK0sVwxxKB1WOUChHTwQzpqeQqyTXjEJSXf1hvcAANpFXCL
Aee8+nKlFGUvl68czrx3XLIP886qeLwlnKpkfZFAOtFv0HKOwKK6P8bDVzNPex5+JYoAIZlT2Uzu
jR92foQaU5tzOEFJfUIg4L67B3hmWHOsXIDPBibNRwJy/T88PDz91u0P+wmNfV6qs2drcJI1dA0D
YFs2DfwdTHmUCctTWpQCg5T+qFN6dq79SFB6qUYZR6pbB4E40WUMeBqkulKXtL/6EYDA0GiLNAg8
SmaHGAz9ia4J3LCcF1P040CX6LjwpX7aiVU7jZrzjMJ6TzY1gtTh2fKdhosBumkfKc7ovP2K2tfo
Yf7OvvLmLGRTc2AIT8xKuOlGgM/AFuP2+kIvdE8/EvceLTY0L06HglR+JbtsZrcvqgs1I9KXuVIc
f52rfyYHyozCsMLuMtBdUFUSSA02Xo1bMqJUAvTfk/cOPVGfpVckDcCTwaCVe7H8VySZewF4kfzY
+FbmkcMxxKtNtWXByks8NOtrP96CXyYhkFFflY39UrvywUop54C4T+NkkMNc8PZoYF8LvEdu8AnG
6SFJl2Ocarps/UyADhBdzsRRQUAcdVLGXmRnPHvkYNjeL70b/JO6kExheCH478mLQ6zvWp5pg0Yr
rPTMazcP1ye3XfMaLMWsvCTnLzI0589YW8AYskGeUaTxWUkHmtb+aiCpmeHoorB5aYmgPuE96BNu
EnRgxzBPQDMEL+Ci2CWa7c3R3tphqFKMciYVyKsPDOmWACrUHJMtWbSJwlBUuI2HZgGQ/j9yKbvQ
Ua8ZC3H9DUAVu/brI3tWCdp623k+hWi8AzsafQF9D6pfp6QMJcHLXKFkX73Cgh4xytbGZMpvqC7z
EStErT+7wEDsyItqpzNvrPCkSTRdYX67VcCB3KZo4zbVPtUkSwvYRU9rkYb6O3msXBh1sKnuPyz2
fVGwe0vvgaS5ym0YGTKDxxzdmel9/mTaIUl2ZO99e2czO51RTm3Q69wy0by0yjXPKeztckjIy+zh
wcpNEAxEinMNtBI9hpbLsvMbMHmwA0OkZKzaKRYdK7rKIDhVjUXqpcDZRMjMQp6exq27w5daZVwz
612j6nTnYBKW9jiQ3txPUXoTzKKZBwxEj4dUUBmrdS2wTmz5XdiYkaxO2fqNrpI53eSX4RAtzx95
BAVWS9yI8KQ/m3Bo/KKbbPqfJirl3DHNgFDXCxp6UEd2qp48SruoC860prZX12kqsYaDAxJHmtJQ
HDfpUCm5Q88ku5e8m8Unw5h4TUfnGUUTi4HP5ASBioGexRHrU25tlQWONjYsx27zPLV0hCKn9ibs
SVfktXUDTa2vKjgjYXnkNQ5xnB63qsbGYH0cmZ+GEDxRJeP3JZFkgv1+85utOXBZNmpX3SP4NgXx
4CpHJtxNoqxTucQoMPRRD/FIaw14RLlPP52GFHll3yMc1aBXvby/Dz6FhxKli5OOYFKS6yTo1YO8
6jP7c5A126s14+DXTAFAaWJslAwxb7kffRT4y+TdKu2/DIIp6rVotw4MqNvGQL6rJcuVh2d1ga6h
/9TL8r5qnfuhvOpSpwgVMsqQuvB49TUSrz5/mQaITGgO1ZHXrdqv8NYneo2m58s1HVbNXu5o0UTR
rom0g9u9Km30rNpX5GbJpLr+/SktusK8xhNpXn68v4ZBpKY+OwP9QIDkc6gCMSSiF5TdNCws1otU
kycNh8qmVeCPxAkmQ/2oZtifpHu1p4ZJPFwJphlDHYnETZFMqHxiIsJi+RbybfB4sny9k9YUfps+
7YBTePd8NwLcSMkBMglISlYgdMYxra0mo1bZVgDY3U27Q/b7tHOD0sFWpKhrfbILnyDK2OKDTv5a
x/6EY3z289MGPGyEbdZYW3bHKpWeDImcGVBvzGn0gwsDBgIIRbUAvUJZbDEy2Mnp9KJ7NsaD++20
9iSr6DX4mA9PkmhcIx9n5Lrl/hyjGkMdm+x4vW1kMiXqyJ3G6rVcbBBvhkb1HoGTRXhyhg8wcf9H
VDznzH+65CmU8BLz9HlpbxM8JcnyXECgAbH2OQnhLU6xjTlNUcq07rrQp5E0AWezuUADS3XJXnpQ
UYSXHdXLvnpR5uWJeEFFjNP7DL55Z41yhwA06u6s7dzCq8oUHg280u9clV2NvEIM7tk0LvgD7yRg
4kxr3OXFOzrrCdiq/dt9Wt/foSYPGttKD+FDhH23Fqw50/aojBPMvE1xdwGQAuvrf1msMYzIX0wN
XEXpzW5QPa3vIVeQEUMFFKBFYG+1FwlSoq4aqnnH4wrGEDeap/5oW/76AlxYBZdIYcSKTzeQDQbB
qfzYwxnBbiXrAK/geGWZmgnRHY26UNO/U2uBMwhxo/9dM2qEnjfM3GM/0p/SV6+w81v+fwSeazpD
BT+ow3ggUoBSHdbnIBTPJefwCwUfBajeVrHk75dAZwQ4ltq/oGb2i5Vw87gI94oMNJ6Fc/5rpRLY
lPqnZ1oMHpp1vac2yQKk0VObyo8b4adHwJ9RFs+i8YzAWr1k+TgExE5zNztllYteqrF9kwo4wok1
AKSwU9rTMNJS7Z0jdHVg2fHAgQvgeEJf3kMnX5qLH0zqCPvYBPP1FiREttaa5YCTOKT4NvcatlOW
lfnJNmZqaU43i0hXq9xNe5oFA492/y8cVD0QklrCbIuj1WWixUxYlk90Lr94nCkrt7hQZWKAvYAg
JguHcpzEXm23TOho1mIhLyKJtnOaT23kufcRIpczVKmm+f9jL57ykMCTMGAnEf5lPYaTA41p+wL2
gCelwzUcW8/sUF65WiOcQ42hC7sNnlv9uNK5GPJiKlY+93BzXwnbnfSwUjW2zgYU8QN+dPQfIRP8
y5tyTHIqKfsLrwct/lUJWVcRZ5f084uoC6P91j2sUNK6fgolwSoRdSpkR5DXLEt+KuT5/Z7epNy4
C3jje4ZMR15h1ynPR+DsteiACEBuCWWLNwV7pWxGA5sPGVlRN7+wEiNg33Ypb9vDikOoMz5at8p3
s8Rwe6E8+GN6JMQAWp1xAcF2vPJ6kDReDH2hNwC29sE8x7QJ7tRTZueUe8wmVuIj/S6v0to1jPEY
IkCrmpDf36xm84G0EAivx01FGZVQN+D0G+6y9iRG+xC5BmtXRKTmemjeY8ta8pP458bXXINhZ814
IcVl0ai80mko1HK2ql0VGpG/kmq40LYF729Dp2L4Kflb84FS+gWiFbiD9yWykidNYYL2+E2U7cAa
fSb93lua377Pz1zRaRp05IcirIIJL1QAJ4MWOArGBqZ8b69LydYJeUsNYS2/ncWSCWDEoCPhR1/i
wb43nl9Z/p3MvicLJy1RKFE4ZbVk8ZtZArW0bevzPPkpI4BOSmz4+9KurVoyT+MzY9ux4k/1Grqj
v4+2ZPMHybwJtsDBcccj9VhCzPRIDq87eYnH0T6e4w8IvWOYGvov6t4T5KDoKTq3Njez0uwow5N/
mOhWGvJ+qKsuda+bYYd+yfkPK/6c6DmR54U4gaHChME9ehz7i2Vk3OtcdhENagokA6OuYxcUtkFl
0JFL6YVDpQA7o2tG7IqN7kS1qFUHUgk0hxulN27ZONvw1He/Aqi0IuodxvdwfUo8FgGh5x5QWuTh
msp4EGGlUnUCiJY1N3LJE2kRLXbRgGFTkJgFPxZSKvc42mI4qUr/XcczM6fooKXc2V1mvsNUaXUy
jCI2yYyVncrQDLUVKj3qYhf2Gpm3vSy4ISiyaYKrW9aDkH7kCZGI+7FVbfWvpjm1/5knkWuTm8HS
OZ42xpthrQmdgBr4BdzNl/EFgJxJ6mkpQBwFQ1tar6SBXXZAkZzdF5uqCkpOlEs56aK1uk7venBy
mYQNj5j0PKFYOSK17B1iSB0D35ybuTvXnE2opvZeIi2IL46owojtdWjQz6HgRAHKWf3wDltVgg6M
Eb4KI0LoTwU50GDAeO86cXJULCgjbHGGA5NCkU2AfuJCMExzUMba/btL5Zq96a8Nv4wtQXcCxRoc
5GZmZsoifcwNuGf0YsDO9pzh8kcqvqruVRuffyvjDv3EOlfYO0QYp1CESBBjRIBSEhhh3+6m2soz
wSjuL8UnUo3Uz0cf498q4z4o7khO5AIliOC78BazPyk4tK+qsnPFkQZHxb3GMLxyx0nUiU38g2Vk
eIRakwJHRr4tHbHHG5R8AM1X1txxhdDxDGFlHTP+OVB3/a/LDRvCs7ZTCq3UKy/2G4fsYIO1me9u
0Hp5O5TT8ta0MvAmQLwPDUzUiuEVPTHXIbyyabLLj35SHfPdOhxD0JBFwLyuaaImohcDnGVl+MWb
oXj7t/k5Wm+gq5Yv+jYj/Vgsp4Vb14szx3iBht7WVZzkjO9QN+dtaNJTKLfepLhT5Z/cXKxh8K21
42f9d8p0oCc4YRgRl3jfw4JHJqgwCYJlXleK38Mi3NiX1A0DCAEJ4z8uceG8nL6V4wiGmmjEkEpd
i/KBV+GvYyO5lUfyfrL2E1MiuLAVrBgqyBnGyF1xU6zeb33pdPH+3ZBeC3CHZG553L1R5fw0JQxy
fjGcyqvp6VRyPz2+qj2sAltRccR3Tuy53O55zy93eETUPCsfG33ddr2UgfYrleXzglATNn9cbnh2
5hGf74nhstA+9++pYIBtKspgwL+yHBAAeEeR8k1biJnonh2Zs7gVt3C5q7Fbg7g3/r4KgyfGqvLq
oluQpVyTbeo3H52TfqOzeMAdGQc/MyK0TjjEQtORJaqra7aCwZwwC+X+hfmmqZnzTqrpVUIX58R8
6RcG6zx7VjhnEbbeCsw99lpqKwiYILXM0Clmlxsj07nTq3mGDOSLUeqp8RxhquNOdELiabJr17fh
ZLVbYqFIN6N9f7adMcBy4I8yxuVeGEj6ZOuCSYzkiwZQKVKXqHpmi3I74QYzqx5uRi99cbhyTgtb
yn5Ch1VbTjG3ynCoRDb+PeuSagJkWmc+MznK2mxdfIJ2rujQtR6MieKHrLN8jWh2CrEOWj8rR/1z
WETGl+tg8ih915n//i6zfL46FDBxBIeWO6r5poUiCRES0SfjbrJLfNyP+RYBAzFd4tCTKFHVk9j4
2q7dsFrbsVrg4Lv0q7rHhlLyuM5XYQMCjnjiljl1AuiJkldVnRDlJ8qNESUtxagA/uCCDUq08NYj
8fF5tCH5rhMVLC8Slwmho8RJoHVZEZvrBATR1jedsckhuS7z50nlbrsv7MQdLQxPxp2Y11dee7AO
mZNsh9sLBZRyAx8JokD7orCZdCaOv+yYFdHmm58H3fvPPXit1D9b5khLAcHChOe0ORBcPKeWkJfy
MtcvNbWj4C/OpbNyELpkmtP9zqH4c3eXreFGinXCulGwvuLAv/OmbLns9DXoe0KxVcD+nb/TnAru
KzbOESPuuMzxZUyDe18cvg4egy5spvrfNFWFtR7f+UgvIPMl7QA8MFDyuB1KIjo571GdWIa0qWEg
aVnHxiX+1PQGeBFKYI/T+l8FtpYGCh92OtUaBf5rYiJk9mryMffhgC4omJwp0nTlxRLEJXqY26if
ybKjYwk/63JTuObiHQOgTSR5IvEA9gYMzKSsQRjxQ2h0BF7FOTrj8pEsB7QbW+2ERCfgU2jGCVVz
WsI3Xhyl4K0hX6VQjvTSBkkjoumCQIlMaRa6xBf4ag3OIpHs3pqkbitsc5aCbhtfar8VDhVWsrpf
Na6WbzVLqOvTPSq+dDN9GiZ7Op1civNWBI30Z/i3EpehTevOkFK4XEIyyqJHVUIdmoJ05WQXRIz7
3wCQtDPhbP9eghbunBU43VxXYxEG57l+1UbYYICRb4i9yo3yzN8AVLm3TfVQe8T6XlT/HQPpCV7j
q74VYPrxQ41YoL8KaaPPA05brSqADtGeOkSnza+RCz1PhD4ZsyxCN7+l2N4Tf7Mzn72fIEakJtGc
c1OIAvL38YYpNaoV+LGUNnkW9TK4O05iz2Y8Jfam1B6dqHxxEYohziwJWqjP2EgmvUdfBijWe4ag
E+JUxvtlDrdWWplIGixfmAQdJjDQ7NQC9L/YuyCKVXqQ5lZNasFTHykggIPINlHa729R+W8RdKni
iSF2Wqprofcu8IJPOSAG46hP6jTp9SF/3hSjb9nkH1JwoKTJF/2nvouZEAIzADtlWo+H6pkj8LCT
+M8X3VCb9jaSBorMoeyI0+uVa+TgcwrUFwz575QqGx+hx7aSuXMdDCt2iNh96n/wbHDPu5HIzzVm
ckgtdp+Y0hb1Jwxd/RDy5blgYqZoPZD165NcP/70A0BfbQUKWLZwuHKVHNcmaurAiylS2ML9NM5H
rOWIPxtZM4i4/DKn7GyHY58RBHkINXmmtWd1Csf172+Ppx2ExNfTMy0o7d6G+xo7DGnWT2LikCrg
tfoRdDNIF4ZIzIjHSQZFhXHV70xZw7bcbKYZP/JKLx3JDufDOLLaUwpTdXP2SRXODXVI3tOj1Ayy
lFbm96w506PAvCk3rhf2MZkJSlISc9I+iAo6YdaO/goic+KfMwAE9WEkYwduvXICflv0AgMCMGIF
nyFidZBeWJuwubRqTRy9uTVktpyABwujEqedp2tRgYGdqzW+lAyzlI+TtXf6kIZi61+KmwbkjSyL
hpp6N8fQCvLld7MZ4YHZ/6eZqhedY9CWCqbPfxZT1N/jjZJOTUPxoDFDxx5t6EnX/JhDJzSP6MBS
XugTv7BLlvWNO1p+xLW8H2MZOZDtPKLViWxMzbrmEuISDRW0AaegoGd5ZMV7KnhTUQOKNViwNtwF
WiVvvk76nCP4aRetY9HB/gqPMT50y2rygoPBKuvnXIGpZlyjvjGCwJJRMOE02wn3ajItmSUrbEQP
Rg6NUwLFN2z2HpDvMHqq6qIvJeeR/TpbJT1+ZaxFrMGG2hS5PJlt05xFTE7rWMFJyerbML6gItx0
TqJVqkcitmRWSj51BVfAcrk5O+DhA0Waqt6X+pXi9yb66X1VLNFfBlHOqxd3Wr8CgvndbQU1QYgj
yeTyHzt4bETUOe4q/XjWUpY2/g9DfZ8mKK+Ngn+u2rNDU6DAXPBUQK/fh2oqMv5npS1u6+MhFvaT
nY1NryWsNMB+oBIRLDHIXjX9p9CxGO8pADqAMhBdAKCVhqW7fg1gQ+Ng4dtFxrdnugV9i6RK9tkx
YdaxK4dAM8XrQs+FaAjsakbiNsSC4o6/fL5vpYdXk99kUAwdVtNtPkz0VM+yxdvL6HsaOzvBHYWZ
b9M4/7eORETGSvERhP6DF0KmsTyvYHk2cRvsxbHsjMaAyp3Z1XuD5FgT8OVUpUPnrC58HocVEnws
1TwMpg3yn7RDRX9UPBHJHefUPOBxCzmhyAfJqyyC1YOU/OHvoZRsYt5F75Kyyuzb8GiBBqhg9ooN
c/FpTA7jOCJzZxKD/SsFqGH1F0qAHmE2DKPXsSqyzI10AycU5dP4a7JZwMJnOFPVgeiHjfpb7I2X
rMvqlqjz78Fimm22/Q++WlnNsns9LdNvuAMtwCinPpCmqEaTUxkPhOBMbBhx7JEVzFvY4Yfj5ht2
7aqATmzvJJ6QaFzQAysrQ0SsvHzfyPz4hjK1VWAhZDLLiWYv8fRSc/WWtiUI0MAbNlLZ8HGOs97a
yyl7VzF62u+Ae9J8c3OhSkIfDBrNRnDtcQnHwsctHjGwIzBDQ6UoT46YZke32bVAiy2kXCDj3H4r
xEFKYtxGFAlcOepa/NHNeg00XvCxX6gqj9mTsjcIphyaawkvTyoBQJKQ/y5FnpmruRCk2TgkU5JN
qXG4ek2i1WJapg7Or8mXrUlSDCs7oNjU1ID8VHxAjUhnNppBJCZE6Sw3NiBbBRfaLaEd5iCf7GEe
CAXIWVV8KQ0kzj6XgFW8LPzttEgwAAulYFm3lfNnIRmfF+FnGDrnVkQbkRWAxM0kixPsj5g7U2J9
ONd08dBU7m/TcNqNA2oOH1uk8+ZSzjvrtny+h2guzZNwgntwP48TeKXT9DDlP5J7rGE3c1E1w6Mj
iFbIlL+jgKaARbw35c+/ChfmHj6bU9qKMh1emPbGPry12zWoyV9+XK2JBsJfyIgJFa6rUCu8ftgP
Z3OTMCk0hjfpQb9yozv2akO3AsToXWJsOY3Mt2LWAPBH0Gr0LAXtkv38nzxH77sx6FS6eoyUsjy/
Vy2BQwQrVEWCSNNuZBhhuCVm4E5+mPkRUvaKsl5PcJNd+JraapixFexiXSwSTovhogOo7Mqtu8sY
pPAx4VRB6+3Pa4+xzsjEf39kIcVaIhfWukAQBV0DFyXCk5R2l9Ratd9xUIGFUA+XTz+O3MsfEWau
nTEBvLm9q9k/ocOBhIX9RVakseq1NPcFlnR5EIxhiCk8vpl9ttcgX5zw5mb81m2O1FSCBg4Xqenb
9VdvWmgbpnoSC2RJRVDW+yCMOz60MAISUaSWqJgQrH7Mv9GtiE68H5vtP46R8q+T6S0tCyR5tsK+
ZDz+YzoVI8zm4o/8OGjuxNEDnY6yu1GCkB18nI4tDR6F2mX0/NasCvyE4cIXkqwaeF4unJT3xWQP
AYyo/goaquKHg4lsFeZ2ogQQBOetmBfwCmy1aWxZuLZ4bBt/X5qdgQ3vmXAkhJTlRdpn3fnVDFVw
1yf+8wYHflPlNgCynrbjIjG17iGlVn5kJgPxSZuIplWkdU+E/oPkC0DV+t7h5yWozuUPxdoLbxkQ
GX10Vx/L+iHwPeAYXhlURkbuMvQQYUQmEK0WB+x21st/mSU781oZZRaNub6Ey4iMi18bcNpJeOVJ
96p3MvczWxgL6ALCW76bY1PwE0QbWyE4IhP7By19wEpGQB+SPdGs8iXMtOm1hA5ii8addjfSpz7c
6tTt4eF7w1E646ADZJzwmZ5ZrbUZvUEeOwhURIlV/rOImCmNlSOQmVt9rFOEATNR2n/WWymLI5po
SCrW5UsLj/37kIZyj0Kn1oNhg43ZOQVk0/ByngpSNkcMZ9xdJecgMaZONtUkB6HrtxbRFw8YrtRL
QwRafRTV/dH3N+GzhIZambYf7HQFop0EaF+NLvDPTEl507BDfXrJIEb9HPMYKCEeOFv79AFK2jEe
r53G0Tb7HnwvAX0ee5KUobxMiJvrhswL6c1TQu+NNloptKIw/mLNZ/FzoNLkX0NrQC+LR+uBVNao
mfDJjvfPaAVHx6BaejGrnZnvy+lw1Wm/2JqlvTTKzusDFV8R8x4ZVpdhapvC4B36ujOT0Q484oCe
dwXT0k5NXDAYOcUEBroKXnxjg/4VLJI6R4/33v3LEj9eOPt6nrZVo/2KwmNS8WJ+mQ1FMT2vzcw2
YXg6ZZwjYDvDeYAdmHb2XNpDmRfapeTxqEbfCeBGfeSO/Tl8VY7HhrEx0cefZ9Xynq9veB/0w2NH
Sgp6LyMQC18y91OBDHOsG5iRgNhqFZKrFmKCL8/N6CpZf9diAkm+uafTCqzUWHNaarv6diOo/AyF
uWK/SzZKV4ssdwsOGWSJLQJPi2I2x3mDuy3qtaUGyqd7lIKCw1ye9MuNKK8hjGKMw2pQ5Z0KzeQC
7qFBZ6xE4GKtG1w2xPTL9BXmUSLA+H1vKXT9ddi08XHiVaud9rmcIeQq3FryWLSZXScXEUHYehfp
zxRS0Yf0hcJLXpvjkhltuDy3Jj/dCGn7a5JjifgosqjUeFHbAi8nwzziUEdqwY8mUS4Iuy8+G1K8
KsbBTAoXxI3ineTk7WfYcxk6H5Qnxvg/9S/86l4uNWVnWG7inBbTC4EjBTDLFO0ORtQblJH71f0z
3thZ/Z2WPuM9D2/HE4u8X3Ld6CxBAtdQA5sNH2W0hxlA4Yjn1N5DQ4xYC0m73tttyO7hBokHmxYr
04JRqhTcqIp5jEy+JRPlxPInVrOP2NfdgL/wDUWQAP2masnwZVLm3euzTMkrgiZQsOTsksANq0nt
qs+s4K7zKk0n87vlFRMvv8lIEOhzI+6BbvdGrrp0K3kQcS0WHA120THSLIIl9VAxo/t6q6eBseLb
VXzvhyfNBWo/QyVgVS8GE+965cLkRYHkl4xGg1E70oF+VcJjWWjs4eqDNvlF4jfFcxcZUt2WWoL8
tSJ/9i2+lIfBuiXsod6wjH8vIP2sxVOAduF5XGus3bmyn4CWcmvBuEAhWlxcCHH6wdKliltWLXs2
6o6B5DiY4uOUOhecbdWL5+TIhUaEjKR+JYUXZ/wCoZhxi9rJVlQoebrwIxuTSciRgni9EUQ5Wa8a
Ii8JT2uFqSShYQllEisZtDMXFAaX3qwerfmhT12wMvSh/Hy1S601Oob8/XblOuT8x01tdQVGmXKf
7qs31c768j3qI25BDNuUVZS4gyKGRwCeVjdqHplnyS5VK8vxCTsUUaQUFB+15WvqNOG2CkY2/qyS
2vbMy9uVUYKKfEv++UHZWUqKekaBHiyTFfYxocDmCcdtuoevnlJo/Vitk6PLJ0/4+UOvZ4ZMonA/
Ra7lLHYrX5phE3uZumkw5+KLXQAxibMxg0p0wlfvq+k6FaYMnte4d/ttRZFOu7zEdNOH49azyqk6
xE9pPLM2HrUxM7Cr/PjxFRTV51Sxp0v6pUXvU8H/a9W1PFOA7AiKQVZlqkxuNgC+4SkPiCDHFIZu
Yz6i2QijYCTRAIUO5FXIWlb3KztbhMmB+08pClgooptRWMtRmDzNHPVpBOs1J38OHWrrLvDMwF19
URRidsi6WC0BNziMTBhTbAUIAjkWeT1Hwk4CsnOCpuxM1z06rjWOoh1I0mUpc3AGh9c3P0jG7B/g
zAIyRHuWbx3BGDr22MKcax7PzeHt1392PDveQSxr6j23UstmTR456n9CPxwdbKeOlhm7qWUNZ+bB
dwe3vmX16aQ7bNmScdwZ+HdHc3hbwA78lttnaYawk7WX+vVQdawfDFEYoVRmkIS8lQJH3LTKmvHt
A3vsFW1VoFxFjrsBE7OiDDBlEE0wsWo44T7Uv740c806aCIQvfwQHEi4MSGpHi3YsdpL2+mn/nb4
IN3tgyfUId9DFvrXexG+Xedhhfw2bDg+Ycpvw8DlqyJL2cOnRrqX7+llP4gELBmCMxyNL1ZrWgtX
A0aM1NfWKayOyA/3v+k6d60Zpu9Mz9aOunKdEVuobCJdGXewMea5GvMFQ/cPxXNEeNU3p/Mr3G8k
JnclTI90RqjSto3ULn85/AHSFPYLwuLE9M3l0GGoUvEnjxoPzf5KeAYItspixwT7K0wVVOP+SLz3
aAev/xhuGT2YTrYa4NWHpeXFk98pUbTK0UTHXsbxkdTIQIbivigsl1VIzvi/GBRX5CuqWxICO/+B
I1hH3Rnj7c+beui+KObd5WLBjLyuEI+5jcOfS8jtfIeKOHAiQVm63nRgMAE+mjPhcTXWRu+f/qku
nd7BnhS/SCy4yUg8DcVgqQZO1cQGsqrK1hNyY88R2zlRfXF4cPwdpwcrIwYCf9lGklhdykGzRNS6
afvbKQe0KD1jaKmMrkHrGDb8KswUVWJRMsag/OEcCh770DN9Ry4PYsbIZtxJPSL42XV2GBDIlfoD
5xMnMb2kRnMLzaxZoojJ4ws9ogaoGW7jhVW2Av5Xjk1sMjCtj+rzbfs4gV9ezPaU+GMURTHwFPD3
Atgkz/4BTscFCShmva/on8ewXkviC5m5R7MpMOiMwx4K3xfeR9ESWD3DFzBUZ2SQqYtEijny3rG0
2PI7YlPTEplRWj/BBe29iljmYWJ7VsQEG2mQOirZ/KznHTtZyTgFP9d4FoL0QFLip9iJqnEL5KsV
L+SpPH4gh4vxITRz0SBgHbqV3PWAoNDR2t+SqNuBlOsU+lQ7aoKAQ81h+JerrRdwiaDSpE9QBPFA
VK2gvAgqF4KEXxSP7PgRMwO8/DSQGrL9FRfi5/nUD69VXb7AseZ8AupsABgnZ2zbBS/Cy5gjQ142
/Bepz9d97i9uu4QJ5t+PT7D/fezQ9+6szC0iw8JEM0rIK8kHcsUe3yaRxBXyJcAMbWjzc0NAunqu
M8d2qJpbBJdWtxUaW04uxXeGcjo0+ykIFFbLNF7pO+FaD+yDNx5E9djdOHidYJTDXxEubKZz4ULa
EiE6XAcd9GaGbaBqRsu2/vEm6+NPjAZyprC4cR64U7KLbm4+GsFxBv/UMXTielnxnqE8/ZUKbkgJ
CwD2zGf7MdQ8fhWHM+vSBFLGvOUzKD6QP2ovQmIy+IO/LWbIIj8jV6j0kezWBhCk6Qo9bsDyFC2T
jaoH1wQRNshDSfIS4dB6LZZ8GHZIBNctVxvDhLHPPozDPWGAFaMtxCwk4b/Es/llPGiO7Lyzvpho
PIVF7GIfru5p/pQ/MacQ+YuUICuHfyor1hCW7x3/WtmXPbFhNX8AYsa2QqqQv6X8wzUVOJzuoJeS
SU+G61/TP7YctdEWPGVfXZQIUU0Zql8KcEFcvKioRQLeNBz3+EoCUri4OeX1plxMjMDl4TJv4eRE
dS0VxNHyjRq92D5j5nqRsne7YgLcSJ9KEXiqMjOhhzOk6OFn6fJljIaX1yCC7sn2vllyIQiWlzmy
xgi1gCER5arODii5OFeiVMFbThEz6Viu5b/h4WW4uXLhNoharwy253XrkR99oNyvCrDfVHOXTK55
1wnr55f9U/OkStp/KJsmx+lkkCDs3Dk+W81177kJByPlr09mxfym2+uOmfF2FfkovJXGbp+ZopdD
VDVsznYffCURg+kxY9xvAwbghugmGEQX8Ps4jkBtQqFG5bgWIG3a0wqLt24PpJl+IoRCuPnaxMsn
gyJwi0WiPb7kNEZdHgB+0ZGl8XqL6+TDZgqdQ3f3YBj960AC22B29/IRgNtI/7F2V4LP3OMmsLSO
FUy3LF4gbBe/qDcyfK5N62GJG/+DtlQtmzLcjrxO230/23TKbgzZezAlqyz39vlHOO6wrF5vIFpN
MGQeMgfkfQa1vY67SfcoNjoc1DhuK2cfR8s0hJ4f7+S/jsQt3dbZi1DOZyBwgSA9NzJ0WfUX6G5R
F3EOOzZcmBxsrzOEUWe19xO6mKVZeHnxiN8Nfn48rWZbJ/YSfuIXxIZm6brFNPbM/o0YmWFjETuX
8Ra/TJFuktuHYO7ocAezfmDNq7fEt4oXYoCvO66G9tyqWxmRdmOmvF1DwwF9Vy8TZTHMIYRDODQN
EQC9pm+rDQsfSlTcorOLKYHk20v3yxVc4E/9zs6XqSDVADw6l2v9BEC4v1Z9I/7eDbY3XhlhlsL5
IJdubZBm3jN+aFAE3HqAoMfCd+1lNDslIvxd2cpVTPaKsdHcqqeVCiXnaqrRR9fHwPaYX+J6TVLy
3w/gzY9jOSFVwTCAdmM3bx/+uRtKHsT67WmclqnXl0NdiCQ2kawkK0nR+btcC2km+nE5PjENpY22
+ymG/w7VEKqWG/sgfEMNnZAD2x/aEG51K9829q7tv0fn79O4YW4//QeZVY0L+2xDP9rFlF8yEpZ0
M1o+IFqLFLvGPVR5p32S0tOBtleDFeQTMcFOMt1NutE1ioY9bu58gOkmA8BoOFUrCk0ZxLB9A8zA
BEZOEj+qH8SFJ5XxUSvd4uscCk5dFfQgEWL+0RkHqB0WGK4uPsmFbon3M+eUuFHdankNCc64Ndbt
wmE7XOjJ/3vK4RHxswagKjdk9JxfWGM7w+IYEMcDJh2JnHPYd3xCaN9mmdrvshiBxzNHwC3YScM8
dkug0/mvQA4uDnVt6N8y4t2YE7xqO+L6oM4EqkYleubDmK+GrB2f7LUiVyupjFVAR9Ak1z5MGDng
KmUVTlr6ARRFvVE166Ytk9Dh1seVswoId2FpcLGn9SUftWOpoaz6VZUCXadXVhqiezODzRusLYVG
s1GHZaIB8u41fgwIW+s2FqrdAztMQBeJVRu7aKIrUbSemaIpO5PJczDL2Fp6iy+zpvstDlGXl0Wv
BZV7Kmb/C9WZxBtoVOR1yj6Li43E73aZqSBFvhnuR086CukndByX0PDYcxeqtIR5vbceMPQSj7fo
f03bS6BDvhkpiOR2Yhe1irN3LYpSLdSMdroOmqsO7lFBDFeQA8Cv6gXpU15kFtHs07+zVsRC9yVa
1pZc/JYodIe1JsbnKuS8EEY9EX5+A1/cJJ0YpavnH2UuJIpRiq+Gdw7+xSaGaz+zp01hLkM1IXwM
kDM4zo6AJOSYbMrH/0IBF4uDyFKbv/86Gta8XYH0bqWX1XDSgR80psBYRrTpXgvtTlLLwQbzAbsU
qaefNTpI78j4cqgplOyVgLcwLi7tU5wvk81OKeFkdS9rhg+L0B0JWNKgal24CjZ+u2mt3z4iKSkK
h30AdzKHfS3/n50uX1oZzkEaBeYW69DOtIUcgZZpr9K2yiF7YmpFRC4a61Ez+iuX4pRzgwV+q9wi
hLpQWsMtSe+P0n9EK4BimpwJm4NUXVkaNexbRvwjrAPF0SFRM+qUcYNvZcZm8Q2N48vF9hhiTn6E
MiVra9vV1rFyjIIkho4OyRFPbqMzHj3NIU0A+WI97sBnOMfeDRJuypeD88mpsOYwzLBHJAZ0Qiqi
j1Xaa17jcL4zD2+YUYeoy2KN6M5UNLQjkiZRKLSfnejIPU2/mVUGQYnb9AeNU9+Yd0BeVg68WCWe
1um6rLE8vD0p/qVKETp6Z47w4lloQn89aNm4JvrApWGKeyrECYoD+dOkOYcL2xDz3Rtd5TXjw2PE
Qyer46vWvxupp60y6KHc+D8Z7J5Lf6o22UlyOrTAp0NJYXSMCniJgC4nuPLrwY49YyLD/jCkG5IO
hq8vQafN/eKa4L8I7S/fqLy1z6yJ9vxxsiGV0qrO9w3g6o4OBsFbU45+zks3YuoAgvobjis17l/E
05i6CfVk+QvBv43tD4Kq43CiBiMxabykB3jd/iP0d5I3hgW+ACcVJBCwd+Y7TFXDXygfuWaBbXKi
eRDov7wN6eFglkSg4COAmFzvf6EzcR5lIlCwd5NCkvh/b47X2VloudxWFrJujd5zLbtvprceS0yv
1jNBj1TQt47vnsiMOlzcPXK2Y4OYP2zh4qIagJstaUnht0LcQFj1dx8QluTSlJ+4aIzzZieSmN4s
k212tH7MNBfbgppdXzoOfIrySixp4YDMiXj2SXQB7ddHnbdogpJUhu1ndkA7WEdfP2F+bzbPJZhb
sDfynENQow/Q84W7iYmOISyXQw3OYzkQt4NTgdD60dPXKpnQ2/W8phhHTDeDC4BDQ1YdkcDTmqyy
alOjsNW8QZFl/AjOh3wB3QeeXPKTcKYErdwcM8sGYnAZXG4rj4X0cX6ydj9iCZmGQFnDnBKunKp0
fVSrEDeC0OR1kfYYSdVXkrhmr0p7EXVvdBDHITQEvbJWNgDZEuATGGdKuf/uaa1n7MqkrDbSJxHf
mmNYALSoJdrTPI5VvDShgh/e5WEXsPYh0xDTx3eCpL8fnkr3TeywyhjS4UKxuPo6YHinG8ctuyG5
d0WKMxyQuqvdhyejQAmEPq+UKObGJmcLD64WX7DHICnmIoENJSSNMobuye5tCc86g6wzt50AYfJp
T+fOZEnHWe1QYslZXS19bj7rVXSj90f2f+zpSIo1yFMWDrLzZ9JxRc3j2OHM4JM3b+MRn2dc5amV
LH/QS/tCWOeBcc0b9SJ/4z3oDc/z81hGFwOtZwmHO806d9761rDtRZ2RVBcI6eVS+gax8HKUSHH9
UqEonPfL41jmqK5IqgqFjXdRSRX4lEq8rjUwAUUlNWnl8KbFLG/w3NuSfSpWos2IFPVtlj9QaueF
OxRr/mnTTWF/cBTb54w5yOVzv8Ok03GfxnW7TKGk4HSKfn1R95CDFVWvIDMu00ymh+LfEBC1qlqA
6brPNoUD8vizYHLi2oBAW/OZqK09gksqLjHNsyHwblqXGkTF7Uys8+HYPFWZv9daAG4q3rIMGSa+
NXzjoRn9O/ZlMmPqd2mtuCIR2OEp0T0A0MChIuUKOy8aHJvegaEDLAznHDZgmWFuWdMmMs8PJVew
I4KzrgvB5WwJJKKZTqqf0Jjwqk86/rPfIQ92Je4GzmPWDaEycUjbh0FMH+xoXo9rSC2SufY0v1RO
KkIShO4wIDRxVdilqMNWYQJztCCI0hGrrxEp0F2xYdPcAVOQFhV7GBCuMB9f51f4mfMngrg5iCnz
rxsgezkMMK6HEmEl4JQ6+2kaikXgpXlJ2mHAGRU/4HQt6kmfaw6x6rB3+8OasJVGXgdDL/SG98bM
pzDQqcaTwKaj6RjYnpuoTdHUMswNrTPdn7ztjHQ9MqC36F903+wsPLPhANQxXtgwc1wSvBtvb0BL
Io4Qzesrx6vHNoxT3sdOApHcR5SDbwd4jv7zYENY7WiixoUbrl5ElhSFSpWwjp2M+8fNElnLlNrf
iJuWpS1wthWWXDMfovKS5QsPqgNB30ez/1aEXw9WMCHpyxSQJBAZ5bMQc9Be/CaZh9csSquZTH7Z
TxoV1FP+piMlCWr80f5jDkbQSZjJWjWA0Mo2zMf50PHi+fVAkRk/PYiWgSJrY4xW1roGxTorKAGu
tA0HGoJF9lZwB76/vfLHVAiWPLkQF2cOnl9MVVNf/lReVgAs9KYBrJlXA1igXFyR3RWLLtAszuar
JqEv9yPw7Ypf6nduCvwkoawlCnYD3RdYS6ZGU/cmM67TMPJBAOJ7oftT2aNCBgJRcNJHmOU02h+H
ylY9auotvwo7sLRt3wrlOZ62/oYrqWjbosc0HcdMQ5etcztrwu4qmHZBX1/aXrF8hc765aUksUnT
HaZiJFoH/sInbwkAi7bKhujSQulXWYPHkSpfnK9irZN8KYAXMw4Zw2kO0Hzto64O2sRYdqZZGTkf
xz1k10o75zW6Vq9r5rXvqdL+wCiO0nb/E6wBLBWUM5nNnxboDJDMYwgdXqlteFefNA+/v1fTTVf6
loulv079NlwgIsJZIDQUOfNeXAXnSnbtNeQV4Ht5KKZ8Qvn/nbr5JIXA0sJzVPWFfrQDbIjWCECM
ZS/pnibgXvyf/K117rNwN+gtcIEngI+13/ky2f76oTgJ5KpaZp3WJOI22j93A8+8fgrzKVYgid9F
SORpFge8Irtvdr6k27oFBg8oWQI3hlKXw98SotYl/NbkMtsUZrnnW6CGlCz2Y1Jw4xvCrgF9ZrLX
cBCRnies3wWF+yqEv1WgoC//vxblmUoUtSTyaE54ynnresjNQq8kA3jvLAuY9Xph8oHpMB34on08
jdiw8iH0eeL4BLDbFISyAKo4p0wUpV6QuVcDQwJIgYnzlw8J1EREdt6MzoNCB7iuF6gCisAscdUC
2op02XUEB64XMG/pC+ijVRiNYr/RAeFpF0LcAvuudaQD9tVkm58Z1ps1zc1OPtbxjs/jHJ2pakTh
91nJE3xGrtwWKgHjSukGQvYXQPDz6kk1MKw9wtl01DsZ3hNQygGOX7n4N1++J0B3r0La4Sr/DqSW
WSl3x9IyoCAhhNvyZ150eHoMfbnBSn+NnjCudHbSPhYXgTFz64MeDz89pPxgZwXTezS1Y69XZxQW
YW81SIMrZ1sKMpHO3DkQu6NpusBRMme/dgqt6hCjh7Ne2Rmrt7FdN8eVqqgJd0x2a/UrdqG9w3s0
jXT8ybzGxPPc0FGpxH0hBGXHV8EpV1Rhq6vm3dyl0eMW4TSHWw7AuABHBlD9I+u6NKBMZLfkZ9zc
H2G9BnQjxt/I2HWzNgNB6bmW7pp6ShQj9V53dVJH/DwcB61blM8/rMm7TXpgJge1OIo0zFTSlaiL
bI+rc/qlCUQKcOmjOi413oClHGR9wvyeEZtAK5QV4oFaxYH/lhmeD2dQmiaXhxKp6orrGMHWzoSU
E5Hjgr89QQVGBli/ir0KOLjtwngfvGAN4inyY9veTVczUb2yZ8ji1NeNhuuXO8YnJF6vAOp02FmT
ao1MFx7JOTWIiFAoKWhrcAFlMkIv7hlcBvpjAFiyAkZDSWxMyhDzo7H/vxekpPm4f2yHEV4BMKY/
0FqU0fXVlf7m92JUBniJbNlcg34RA6ZhqJdbD7+Eo/0pY/+MCmern2JRF6odX0VYIMgtfve3pxYA
w7DHWIA5Vr2hGW9xHs5qFzp7xVONmSeE3Lgo6npi8S52v6KADeWBHI8LHcEKof0nuwuO0XiJ9s9b
FeQoDm+6JSV3jKpdHAAf/qGR0e2997KQNVToKu0XvsTo/f3epSp6TNrYn9Qaw2Pr325Pd+WeYyud
xLJaQlWUMz6I5hYdFosiuHHiUr3rmUkYdBcaFFK8oV+UwUN/3i2o/SQKfzWRc6gOKt6LUCMgC/4L
Rr4RSyRTpmhnbKORT4tYPKmXwMkpOaJlgHy/ZGXKAMdwavpd+bJ5osdwFZ/ct3/DcrxXL0DmgZ1S
XPtnQk/o2UTGj1eYQnJ/XsvzrUST5l5qoTs18srGFb183ta7K/WI57w12j5mWL+K/3P6nia+w3aL
TdBD+WeOb/0jLBibwiTVGE8GECvOzBuoId2Qia3GM11BQhaE5XouAQw9jJ+i9d067uk7IXFzZqP5
AVLbjveKlrajeN0SaqxCTO6U0JUok2X7ZjxUeU2UtlZMyZb7SQv3oApw5zfX5idzy321Ndcpn1R/
mxQS/1TZurvME23VXEaJUYGhR6Iw2eczfSV8iwc1Cvv9VFoy5c/b8StCLlJXuYx0PZnLQ2uZNfjX
7AxfXasVD8Vksj9fQLak6KWHFBrMVi74t9qrngkZnkaiFJKYizDRu9trL/06BX6JaVJbE03eUwSa
JfOl6aZLlQ63DO5dw+dPZsoXI6k+7mozk8FyAKkFjme0Q/DOOgah7M9zZRFBrCdioXC+G9Io9/NL
fSHqTjiNyK0eCNhAWYXJc0cE4XAwHcQlDnkfmLUEM7ksZyLlMsH6JJ+IzZynVhdljHsW7AhQZbwo
0T7MLGTF7zn78FLWdGfsGAvbA90KIdggVaVbETJuHmndx+rRFsYe6mcbC7VRgSWlBWjd2PKPb2FN
/Xarl3HHFBRaroF43N0/xcxiEev0yXRjlgEhVwLkL1HcpRK6vzItbb0mhSybrnb1zrInFyC5VVEj
jmRbfrgYgJQqJkx9N3flOMJTCwOOkiCkI/AyaoOmx4FKigmVYimho9HMgLImAI5s54XY62bYgPft
GR5WnmEXlF4gJoPkXOz/pcevh5kzo/27oAejKxP3FcRXejnFod7A0t97SgHVeDs1eF1D3CkjLoyl
OKWpze1BJrnJk7mucqUTlWeNhKJW+lVfgRZqsBQ+joyVGleUpXweJgtLcYQhxlnK9b7llpO22583
Cjv0vQ7vleHOwU0Rn9MLwQCfEJlaqShv0KtxgHVhUhZNbi16GbZAHodHCQCPph7CpUEE2/JSABym
bmq36IxxxOrBWJjVmLD15DV+JEYSbJ92k+Yc+uL8zIQdjtY7/au2aLlkbNlgwBu956qi2VMqK5sX
FcjvdKZ2RkVesymc6zs9T7eKS2utQVxdGl4J3wGeIWTa+RNCrCfCTkH3dzr86UQFJSEhTyBJzvuR
A/vKCs3AkJj+o1AJFZCWKXsg5PppA7tnLlyKM/gQIMa3y6CaqM6LOYwbvHqNLr4J8O8FSoX/shoo
PwEIu2sUNaZ4pzksqgHsvLlozImJpCYFWHUGACF7yW6l1glmnPGuqeKP2Xf5hd80XYFkAJVoqrPS
mHRGZfkgF3jt5JjI65aiekQKLSe2NLjClwZlJDvZC3Js4CpyNxrfKcxKy7NZy4fbbS/MPU6PsZhY
UCKWGgSIDYc38W6v6KJqYOvWPUA8CvBxdTL82gaNwfAm3dHtJ/dx2zQNBvD4T7k9/T10uL/cplnx
OaIHDCTL0BGoh6gLM/jdpJpZqi0pcIsc7Ik/UJZzewCPK584RclGIuoq+jTlfxzCe9yxSSxjeeM7
eoREg4QFQzWIToRbFVZiUt3eDLfzHrDA2gFbuzIqgh9mkr30v33TsoXesOf+Lb90qE3TRXnnRRdj
6F6T1C086OqaAeX6qEykEqg4BadQM73zCoN86P3E044jtRZ3S2Hu/YK/HzwmETy7RzZDAu7lE5if
usoWFrDPtc5Z+3cfHU9oc20/iZKXW1lbfZOifN+xI9EH1DrRxRMlLkuhfQ9fGujvD+3ZK64QcOQT
tdKqmdZtrlbhCNR0gsaPKA8SSOG7RiT9zinxOvdOeLVAuz0Q/K8HhXAPgAL0zm/vrZvHDgeyFq7v
adyEtUzyWhs6ZdMJ5o8V6lmlITYh/6wOqTeakYJsBXngoJZFqX+BmeeZJ9qRW/P1vVVrV+M+IvZb
ZXDtKcXKzb7lLjaqlAiaPmZ7e0xbbs3WNC69bWYX9M0W5NB8S1UMiK0cRLpBJcKamI7MoXVpsnLh
JPNnt6T/73XOT7Vr7htXuno8wSwi0b6Nkv2PpjBLnbWlwd+8mVPjeCGYZxXLtV6QsvUXuoQjB/lF
3DV2ysqH427uMAlL8pQNvqt2zEgob3YItezOJ0U92cNkti42GcGQgTbq27zkJJE6kvGZFV32OO67
IQL977LVKJSNHIW/R+ngD5D1fHuTi8ONO9DHNYS6E6fX76NQgPPSIlW1EtrnyAsrHDeKRsKc1A6t
SODkjzA9iep3R6jZA/gZS5cx1A5MWHCfJUtFwbLJRAR5AxoGBnd2ijj7izI40NU9ja96XP0VNYMy
3ySPZ84YeQ3aMghlG8FPXqw7InrhaR2XredF/ppYlX34rdveXn4dE0YiIT6ZwbDAonDwARRQy6e3
nOFVNJ16Y3SyEaF95kQXhpMF38dXZbVGmsK24yv5+2oSCeEeULhB6l1GuoxkfTPYg9+9ncR9Qy19
ibdz0I0XJkdAqyTEnpm7Xld80IZOZnRElhMFfNzofOYq2dWaPChSrsCAFOI6nlwBM6nVXlEW7Ijg
k0KtIycoisGpcqVSJBQpOq7MMnCmY6+ACJ+WyIz5ADXpx88d3by99wSGCIDsstmzqX9sV85qVqGL
bH1N0cz4FqSK6LMgP3uTbGTjDR1SmT6UXFR2iLJ6RtW1yHJt1UN0bKQMFjPr1tELR0El5rakHvrm
tv7RyM03MdcP4bVJxnFC4s6gbQB8XMr2mkVJUJjszcAtWGc7O1DRhOmKK72y7rC9oETU6UW1BjR2
wzjgOwhclCw89X6jnaOJ2yKO4L0/Bbg7lvrraEUkBMtcWE1zwDuXSAvh2e7OBNYn4E/hYFUqrBZJ
u+l8+KsjZwSJwRwaszn1teCCepb4Id/dL/+5UwHCJVmb2oAyGVoG3ZNb4IxTlTkQNyWGw7Ftv9bu
RWRj5wOjOW8+LGoT2/7djQUE2VHPHOB38LymDUGSfxsfce7UfHeGEy2duwEVpBcgCipah6PxK/X1
dCTmefif8Uc7Vo1xAqWGetkP9ISZlQGKnkG57nHL7KQjYp7ZihvNUNrvWXv/A4t6F+/bQWU6GBCo
uocyznEINxKSxkqI/n6nlzUU9TyGArCqbyZewDPmDjaqat7kw/1Btf6J4eL+/h2xrKTcPxOIni0/
EGNF5qZl8wo4IN2pJj9FuyLSDBdg96qw8wQwX5AdwFudZsJ4WGyyBLUmhIzXBcrf7gN5B/p65D2k
vuuyqjwnBB99SvoC9R92XMVHX7SrQJr0HG6J0NsnznJGbT7eR9HItpGtOqIEv/+gJ0qzagn0qACl
ttFGYqrj34o9FvY3UkpTmZHLJY5/CIebKenxxOvxTBNxE8hoyHJv69vfEFkJgVIZBvqT+fhKxmeU
csHFcGBLsZ8ce5st0amH4Vt3D9fBmNn524ypqy20pG5yWUoK+mXrovz3EfZA+BbB5+RGkmqoSm5s
CbvCJB2z+hyVF2PSq59K4gj8prMN+G3Rhw/fD81ynCU7zMcQO82GxG4B7Gtuq3k30tEEbOkwRTpk
gtn/Y6xSAMkgQOx1pe+3wijkUjoFHBLgYkOtAUsbuJ7CDtbd5StJ/IvTbbikWVPrD7kdUvofuiBW
XQRn5UjXBQ4uFkpYnYtxoCYXfybNVrojcPZKuqZkyaBCJabQUXhRezlmzdBN9g6CK6FzJNBZvu5g
klGOWZjvh8Qe8D6VUOe8i+C8qOmBzIJgnDzflYlHYjTCzF3mlLaA8elXMfTemc3Gcywphn3KxkSD
ER93q0bPARJCAwdVEAr9sNxdv+8nWn7L5c7u3OrYcj8dCGtXW8TWzVEUIeyA2CUnaVrArtVHBEgx
B1MZ4exPmdVyzupbpFU6lcB6Sm1BWRgeqo6v0v7DgXn9WvumtHN269DmuxvOnWeA59jsKA0PqOVv
gisRxSQVaBx+AgyeCVVIWR31R+KtLmHLNzYXnosdKzaM8aSCkM4f5L98Q1wjJzljBbh6K38VHzsY
9djjqVeV7b4cr0nFjaB+3Xnk+Kp8LXheKScz4hipX5do3eOe7yvx/qCS1173ivLtlvcMqj1IrD6V
j8DtuBMephFxqfHcRCphESpC+d7RVEilBZBmOdWor33Qb4Hm6jiAbNPJOztS6W2IKS6jufN2ZgTu
X8v9uWlnONtoy7qTt783/Zf4Xl2OCIP8zbC2A/XB0TozIGr0dR9OGh0BMiCxmi2PtPVYa/bKalf2
xh3PZvb7N5k7FWwrcxtZWZhW8NSwC0tG3uj4Ma2ugeQ7m7GWTK3enbk1c00s7kv377S2+158Y6Os
O7Cc+cF8Su/jDGeRZcMpDeWK2oO63Fk16p3u5qRvVgifM4Y51M7yCgvrMZT2AF17LR/Wl86V1bvf
OtNgF8B/whAjNlpWXmEVkm/FkwLYkJ7C3dwgcjp78phwwAIPejuI3G8HvTXN0tMlQADGCBWT+j8z
ZwTL6YeGlIinR+nnU064nyT0WlMOs2YssRPomkbAdkgokUGGxIPnsw8u/wJ+aVx01vAsyiaittIy
g/LuaRp5fBo1u5p4BYVRAlCqiXX7afcN4tJ4pmaGTZYnBdB2gwersTlAj7gwCz0RlxlpFkx/88yX
+UY5CQT7MiDYQqB0INL+7df3anG725a1VlqyQt9zEWeJHjJuv8x6i8a/l4yO0fk5aOCFz3AtHrvb
or93PW/rN844FvpkX1f+zplXKXn14iRK3KWwuW5UOa2A7m1Susv6GHNN4ieGBlAJi1upP2VzYSkB
/4NllBa+elFhyK/23KB5JOQkFsE/6jeFSvqsYr102jvi0AFWV3Q3mFGCo/8hz0ar1YymsL08CvTY
iRyxM5R7QVWVhMXt98HDgZla5dgmbLV//xBAZGN5bFknu6P/qIZUN9PQyiOGBTeiY8M4UDxqO49Q
mCVoNlpQGxOEKvK/YcyDoHufp6VxQf69wqwpPMVPaGJsMVQlE1PAhAGqJTQtUZajEvyGaP473914
NjnLrt8tReHV90X7cck8rKmmd/srQtlwBKaMMs+irO3nckX4cTTSrN9hnofSJI60gqwiErBaiS9x
caNSkK8cOeYdMLKFpb5oRvEtYlBsM9XqufsQQt+a+Cwso49IiGuRUruKf1YB3z04sw71xKuv/+q5
XyH5eV5ntg99GMSque3ebFBzhRrM3Wj2sXMEOnhtbQTu0mbRQPr1342UqneouayTye05S2C/jnh3
UuUFW9a254tkFYDL9jcznG7ST1qiNw1TLVtIzv6yu4QQyrWgN/xKuX+xYXCtyhENswmRBvDxiI56
HWC8XC+0Gd6yI8xoHOLbIpKpcnsUWsZZe2LqWTtyzKEZ1g+g6jC96MUQPlGnKn1L4idnPyOFIXpr
Zvj7bKhn/bWPWpsxCCAlvX/7nMVEL6KyzVbpS5F6c2XmREUPmCFg+N60etLZ8BP75uwhEnsKn4IO
vwhQjSGEWqEg4TV2Vxg84b/GrgcYPTGBXY+gjl/3OBxx9u7a9wRt0GRXCzf0sQbq9ACzNHXZ6YoF
DyeLXsNUAPYYjSwZgEKULg3wxoBgI1wiWPAXDhFrr0VynTi0N4EGmjTp1/iA4XPWqAAnX/94im/t
od0aYy78lQ0kyHBg0bATxePIhVni+imJQpl66IrL0V0twbDKk2gjUevs67sE3QQl7o866qduxvMO
MDLbbvNM0Z+OI/mpthiZTZ7oRERNP6m6dq0UfvNjb6Wdt/2C7dNSsk94YZphgSVhDrHJFX7IpjdI
qG2p9R5lpHgOSFhH15mTbtDYoHVZ3ihnNGyqm0rtmrgDAdW1GrO4VDh56LaF0TQ2z2uvcUhANney
XYaHNt9YsVGAe7lcnK39/t8wSmNWjGuaf0+NXOiQltsY885H9y9mBbO9L8Fp0GP4IVGD9Y/HPAcH
PXbH8r5BoT2Rk7SYXjpT5X5JOui3njrPUF0hjn4H7j9WvE8sk86WascMAvR1Pam25djDkDuIVJV5
v9b148Ielw8VQQinvKpCS8KiF1Le4HeVdwr+0rGBQUWXVLtoCyiPhjFf2HQ1wTDmC+czjf++8wmt
k/V8SQn8wTu+0+zxF63kQyo9+3gZ7sqoUAPaj5rLf5Y1x2OBgNvNvG0yWm+0Q4J1evO0YXTOiICW
jC1ohCz2b1/jM1zSt4f7Xetqm2/6bdx0He+EVSI5ssSYEVkpDuHs4or+22UbRKJOaS9kwUuLNkkN
a9KPBKLGK4vOlbgjYG09rUouB23zsxRcOpLbi2GLBlgoM+ZYRF+mhM/ALoW4HJ2xfHSppkjq5Lt5
OlPMRbIO0OK09C8CSH0DxSVpeHp4BlSzDEZ5Oo1pVcfya7tOeq4icRJtb0o+6fd1GAqty90uZqA0
rwyMHS1zyeIVqzioquDWeuYqQ+YU4e0tVGqw8Yy+edqG+9nB8eTLutc0DuTPKy6Q9JazQeE0TwIu
OmGsQpwmrFP0LZ4M2LEUXQmq/SGSIeroOeuyGjioS9XYBPitR5SSENgpUAoUgkhU1502s3uIYn4P
9iG1uS0QA6OvcwCGlNW1OHiZ/GP8IAq5738lYNt3PSsWesFy2g+ghjtyOt85heL15nIsyF9kgUqB
X92SB7Hpej40g638K8vFA3Syptf1h/Avwvf5+n3PvnXF5gZ1hn7uJOl3HoCm1BMTsUPHL1cRIJ5G
oIPjmkgSUlhZDw7S0CC57Y2+6gKIMLcPdb9bj4936RRWSGKJ+Z2hsykQkemWiNaM8eLXq+281jnf
pqKMvwnw0nEo2aPGkNMu3nW4CPdpwe+V7Og6mWdCZ576H5bAOgmmVP46Zn01keurHaGU0GaHlSJm
FI6RShqhnghPaVcrnkUKHW66P3cmzhjx02Q27rFsVcNkjDRHggGzkio9gJksFCELigHvjwortMZs
RfrbwUmbJSzIbJol/8ddrS+lo6rdqgmar3IhhMuFInON6ECvfmqsebIMPa5eTy0JteF6wEiMZVe3
JqhtS0JwLXoK5oh1H8tlaczkBcprFyoLi0JvIxYiDmrcyJxiWPh5SdDxHjbCGBACFYyDicEMqsyT
1VhI9XiJ3FpT6dL7M56xXEimhVBPKO73jqdRsH4PX9a5RMY/pM1Q+u+7dqzZBT4uhjAqT5fFu03y
XnJdmKY6M6Ynyq9u1Jn0NI/ZMhSCmWnA7VFjIQfCLAW95zJ5Mh+JyV67zQ9GFeNg3KPK9buJQpTh
ZiuTtAdKs6qEJDwcG56rlhUiBHh/cB01CwU7bvU2a+hF99ENmQGmALXCeqPuBO31ymaDDo2AaUBI
qs/6w+tJM7aWHP7bqXq+AdY3JA1AsyKgi8MiwCjof4imdXXYMfsW3FYmYVpahlcRn9G+LonNmgxb
0bI2ma9zLGKKT4fpnXm7CpzYg0yi4FphxKkTJ0u74ljnkwmz6vjLCtcUxbNd0u4QzrPUbfa5iqT0
EIQWLHPSqwut/LU8+FlXt0VHwJegpQrcVYT8MseVitBAUcPXL/3NYdNtcLXD1owjLcb4l3C+nh8I
K8LbpNujlqiFXEzL2yLG7Z8ayUOp5mKT69D5UmQKKqYj2wwnx4/77zKoW/TeNgG79AYDUH0yuoCS
LnY8wt5gCu4NAERPmGkK0lkLAdpT8n4nqc6oRcOOQqRvwgyoN4E0z2B22rKrY1mWw2hPJNSsEn0Y
L1FeglPTuuigMkgXy/6e5f8f4r17CCZYn+qenZ6FSlTMtiHg4FJd/dzydPwnkrjrwwtJ3bQ+oisT
jUnp+rhi9adSfixJEXqglwGoTQ7Yuu1mAhGUa+Zr1xZQmyPPJwpK3iPa10sGE0WtGiRYawk/Gajt
LuqqQVNKKYz2QtBtWP6CMjvdhKNGHYV/BNBBHvCp17lF5DeCg/e0cz/XEXH1g5wE8zHutEZ7QUw2
3vz7x3Xql6pwvSD5UB+nHCMY8JzdcDKKJyLZB6kXHCZb7wYUW204L0p9KDLuChtZ6M7qx67WADJP
sQo+5gR4CqhsZLpOazrMEjyHz7YeHe6bzqGJsLy/YzIZa/YTBgNBncuAm4C9Ukk5xz+a7MZ8k72w
8aFIf4sG0qGCfKh29NkC1gHaM5uePWMZ93AD2AthoDmXk6O+FkrEwtWUhnole73heL/jnR3KB9EG
itL0wMh+F6Q1B0MQhRXo4fXX4x2b4bTjf7LTReAQtubU7HsgewrjJTifLFuhBpHshJR5Krkg5H8S
wsdMR9CYaIdjlZrzYJizKVBQR6U8XwNr1eDB2qsK1q96LW+9V0IVDuwOFpGP4Xl/3UbyMFa8julB
GbslMpaXLC2P7M30bopBAjg+YgT0QKxgi+c2dVo5PZAnXRvLPxYmhyp8HF7vIDOg6coB54PzH6Yx
Z/sYRerG31XcVqRcZT2mOBQ7EKJ2JWSONGj0jwkglvn07s/lAWVamd2pZowJFO6+EZHMCu+jqkJB
QhHyoxiTUDm/gHG5FsmZAPBrORwngmtplZRdWE05al0Tl9NCKJklWZgnZ1YRvHb1tBCv8IhTVYU6
idVIbsiUYj9FTIg6MjYgQ19XteovlxqI+1fBmvXXTJCZf0tq9/M2vAtbHZM/cTT6sYECey9ezTF8
2NyQXeEzhnoAfS5spY/XmrTCVQeT3ZAnRUmIT4/bXLTw8XxEDrhHoa1MmOcKxgELPtSi54BROxNH
WpCxSeNODcTqFuH8tvvuzKzQXAC97S15yzGe2kuMHvW1JwiY23YG3BDpxko/lxR7d8V23xmP5/uQ
VOYIYl9MXahiK4OG996apM+6XTPpdPvV+8Z6I+LIGrVHbpsnSZWhIcQrrn83/8UB/9sQaalol/oK
7fi34r7yOAyDiQah9hEfY8O3LvDyEAJZTDs7KC2bxgt6Nb1siMeK2ylX9VCSK2Y82vkZlraN43i6
rZ1g22FJWq18RE3LR+G6Pce2/ANySMrN0RRptPTjOS3aLCw8h9FA4XbwqW+Ih8/K86blm+LCZhM4
q+lHOjCtzIEXx2WHcphXo7AvnIIcaFRhY2uUsDP6pz6NfmtqESF1Bi41jki0wQbDGlExt2naZdRF
BkOYJmcbDN+tg9/uH+0nCkmi7S6H1j3NoqfxE1WWwXc3s+8NNIwcZwFBJj9F8n2N20aIDdwQrYxK
YIYovgIYvRJJ+8wkmk9aWCQgykNpzDKa90vG77uSVnzF9PBv9+tzIAKHwwF3tvtozjoSqoQ9EUEN
gviuXu+iB2ZpsCJG950kVV5CM4TDEGcFhmjbnGRyhsTHl7ASgiUOEJj+ugV0ZC5E/Tb3lZ/niiqf
4t1567K4MMy5QbbTFRHazuT+GsP6P+hHtEgMk+gJ0kKzyDIRwqxfsFQF3GsDI8I6pXTf14TDDAIB
OIHhQXBjgPCt9K/yWZEIUZAfFFpozm2A1FnNDthNUQAodOjQmNr26a4PaxARbhCmVnlyWtJWINIG
UVH4nAi//oDzqbqM9q4blRj+N8KWiIK8VAryIASsfHZ6XhsL5cT0ZELCgJeSvbyQiCAqqX0l7H5B
vIeMuCXmtBtK2d9APCW+k6p1Ko4IWPeAVCVS2xUcwTmzhiDZt/Y/V6/Dy0fWUGx6jIDQFMI69C/p
7BzicfKtNQ0O3lmPYwhY7W1BxkhVrt+Yeja0cNE8sOkWLMCXbxVkPDTyUCP9CXx0RnmFeWHQbDTS
7C/bh49wIuO9ZukYZJuw8wB3H6V07QTDKpgWm9HZnmJa3tlwCmF9xBej/NaUt5NPrXUPq3kJ0/wm
cKIo5TMGXcdELyyHB4/vAQmoJ4oq11E3ZX725XdfS3Lxo2CNEDISqvA/W7OJRErxYoCuop806t06
qlyX27Puif78bp2XboNtPPsUjCheVYpqhg8asK/Ndgmkv7o9XtLKu2MwqySloUpViRCXQJvdpOGI
n/7Y5/gQ9ZH7Fe5crfBbAUII7yQcPtvSa6SK3gY1VILHU19+bZvFyeCyaoDxIpe4K2FFjJ/CrMbA
GH43X2XGtmG9hJCvslpX5MLF3PAKsHRYz7LKxJXLAu5uWb8MbhiCQEDLUsXsff7JG52MLvgnfEzn
Qz9ljLCIQsQHSuU0hVi1WU8F/3SgmOMedRfQcmj0kanS3xWPIPaYO1Ec+msTegMvt5vjX55GoP+W
h9Zit1oXoJLVY9Yq7HEBM9hnasKdQNReJEzryhN4skHrMhmQeR1zygQL0ZF+9re8hiIorfDm8fuT
T+R8/nitI+jJuOqEjC6/VKPWoaDRnoNRxShmWVqz4sYNSS1MMlx1BxKoPKt1V+0/uXfBG2su8AZx
4+bv/B+SmMDaaQjULIf7fT+hYLFP6OMcyinBVdShCLVfTST3Q4HvdOwFK/yzPWqHz8ljdNrCPwIB
Lk0itqm9u0vpO4gO+lwkR+ce5kmijEh4QIvDb49pQT8oIkjF4odDk29qvH38jUx1ibcUva6Z4lsf
aORmNKKVrF+wd/h1UYc0PaxREHNDv/dzHNnivWFrvYRL7mWIiBOoc3NrYMChvWLChmsWJknt3rKM
KCIQ7Sxl5FKWZyIAh7hPD389P68LOtJxbXlJxisVtXuBIRNRqEGjBuGk9tMgyaXAnFWB6PPqPRlD
1iNuY2ytFXW+IVjf1Gg3Ni3jCTwvK6etkZ0eH1kdOu7ukBD14D4UyU5eCiuIWBCOSxF1NKOTlNKP
gWV8/IaFo5HRjYXmlFQRztiOUy3j7YaU4z+aoeh/IaHf17wzHOqaf1qWcZSd7/11+R5QaLxYt0Q3
Vn56VZu9TOSjaOvKHEKMZPRwbrB9oUSwiY/Ycgj9Fx6rpQF8j56imoZt3KlY8whq2u+p8rWoZuxY
6OS2R136BmS+ywMy0T5aMpvl+oPtyAkVv2JFMyfggvWG/LaH3nMVOQL6sv1NPaImzZ4QOpUXvRa/
DDTK45SpKrb2MBDSZStQWw3hqvGao0U5Bp2ygfG3+MIEkhUoadGEf9jqdICxKc3lmm5dVFLLTORJ
JsX6xjcE+rvwm6LkZIBmGHuH90Jvo2kLdokiv38wN5qV5PWajnAOlyF9naq1hGaNe5fpD0VmDZBy
HsaDIGl/gJla19tP4H3AfQvt2tX4Wo9nswWg9NE3un2UuUUTB/ThXlgVKj2WM7gSf8Lt3liyP8g6
dEGrccelOoDy7fv7K002J77hvc6KNLMuignsLIv7OV6zumim/1VdPDXW1x0N1HgxyZ5f01c3sc0K
Egv9sVPmxe3KSPbI24ulliBdYhy/93bNbwMH2Pq8sQgPb5NL3JwW+bNsAlkMGOkhkyLOgSaba4lv
qGTIZ29sLOC/P6vACUdpRWmHpyF7zrE2ou6C85wtVNotQLTipksVFTB+toTQ36HZTb783xd+lt9b
lgh284BKyIPVisWg6BVCrfgwSB/T+rTncHuwP1x5oByurZ1dcf+MxXPDCUzOZ90hufWyN88iUspG
lckLdk+1ILBt7KX7lO+8SHgCX0DhuB3lzT6fbUoK46mVtGQhCJeqtlluLW+APmiysxjHiPzbGNi/
UPnwFuMguhOBnzH5Usi80TSPaY9FSuiKHwBeFTOz5y3/+qh4NuYtsFbfy8x8R5SIJis1eQMhkKfF
73yFp1pc67L9roo/OwI5ypHkxXYQjoAR4Ay5g5ky5g6eFU9KGysdGjMQRT9gGZWDIpmFyimZTjhH
FrRdxlO5qEh1M2lF58yDuTp+SGjn6GGQb4QHz5/OKJtux1ZTUNlr3kA83rJ+2LnUmY7sf2UhZs+6
ISVj7wRUlYLgKnOLgQ0amUvksTnRBw5aXWOxW/upE/i+C2dDEttIrv/yXj0oKMSSnE+yG9LsSy4O
cfTMovoa1ypxpcNs/YG97eDzM3X9WYkNcVatLDj+6dvx59vgY/J0/Q5ieodYcytoGKCutWvemsT9
uR/boYnro/N3tD44IZyKsuT6s93nsWnD6i3k+d+d7iNJjnivN3k4hJPQaDsq1XVnbGBALiU6BvCy
Cu8lBk+Eb7MPPsR/eoGRXjgpl+8YhEYAl1ie0fesQnAQtR12e3BQBL6zLKThbwhoWNawPoD/OuiF
hyqSexGaDgP4Sk/yCtkRQqliYaLiPRQWwdCizQTOl13tGp8Wj5VG4El5bJHPLdKnqwOPOn6D7Wu7
k4Ph96/+D6j7wvU+eTbWHbw75Wig3FOV1q9lmbBSDZYgzoUWUbGjZ+i8tG5N/xDjRi2kmLOW1Xmy
/gF5sdheg1DYicx3peKde4kk8+JvkajE+75q2kgv2eZmF4eX9gtbLhlHsczOVlRWBsOe2u4j34o6
dKJPidThk0uJh+y0wnwo0+0lQAMa2nO9IgO+AkvEwCsdwDC3V/xF80RpN3mz6WbgoVDmPcTMRZkz
lg50SDQs7BSaltup75ON51b722NGA+hmKWVOhi8ZqzPbtFipu3v7aqrSpY04VLZeLEY98WHXAp7K
2sNYlgv+4bKF4s5XrYQEiLotZ5mvHHaETsiHdduCKPCYQkoteSOgQZjED4BEATISVu+SqKZjOm3I
BjBCigylWB9jGldTbd6PkBAFb+cBIHJHXFDQ6y8FH9hEMIsG+dRLqF91duJqqbbJACcA6RugpuOJ
LMNbYHD/5ZYQDoTWSMg7qNEIdKCMxxwLerBfYQpRt7SPaDHtWoAuv1TG20i+PL60wSoBZOET5H8w
dYnVsDCsZvwlmK0o8QfkGdssoJFB669vZwOWigK0Pn9c0FEN2cRcE6AaAfNgtArbyNbmxW2ILeuY
WQLc/eHTBinBmT41x7tNUdWCKW36JXVQErV/e6sU7EW5R+tG56rjILLEJ5IMrGG0KDtnJyfKQhUu
MEiaMEdjV585UsEakDgBt6Xcbamlyzpvhf/uxtYadz5R9pW2g/7+K5sXusJWpMI0lHiN2x+vpJgs
kiwO/SVf/9GpYHwZnRoy7KTQesD9ygNk29POif/kS0mNG0/7SDSC73mWEvlngx/STsFY2ZABEZJu
89Jcd6A3iFOBN8Es8hnn8/8Mb7vkcW863jDY3ZRwoRu8DwJXa7HTp6rBZOdsN09GeXqTMv3WZ0/R
pZgOIYRvw6ZbdJ4ZcLeazWcs0V6W3mLTcPVJjd7F/82Bv7jZvscMpXMy/WuvSIKtUiMJyanEzeYY
K3nzdpiW56MZQtdbiP/ChaGHzLnHp7bEE0l2J8CF58+gKU6YQmSoAti+69DfHQbERVnzn+71ueSN
fo38uesBD+ZKveHwXd6/WZ0revb+IsLN5jYW2e++ykBh93kuy44yKOj7dWL1p3It0JlthzJztE3w
yWEoP0nyiHwhVD4SeBMYQh77bAMJ7qOZCIIHouNnDiIjPbDgJZ6/qCJSRAYz84AUhkzMC+HKhoc+
o9FbhSWX4srJXAaQ/SP/X7hqt2DLoG72/9Ix24aN6knAs2C6amXVyC5mKdJi5pc2Addpi9FQoOBT
o2EBCzYmio2z5e+dNf30tS4zXgVdLze+qEtwcCnZ4NydmmguSGFMz6tKJIhkXYxnywrVzUxC2Ajh
VD5VsmMB411iMrFf1OJ44JWI0YfTkI75S8XxcIQ6Qd8a0aeMDYa5VoTqU9JQSkm9D11xsqxIpk4p
fvZK9/i1YN8G92G9bMbTSFgM6ebbecpn3+qrkHiwFOsbyQqoK45VSqFW958jAQmXS84LhovVWPiS
8dm4ZCwN0jPubV4Hj9A8F/FLV1Pw53f3Ex3DLr4yRLdqE6F6zfZyOeY9rTRB1BRJb5fT2L7PJhNN
sQbe5C/3vl0Qbcm+mxKAtrt4uR3f/YmyVUsS8Qn0O0j31Aeeg0fAYDEDBXsnBwrvBv0YokrA/Kvo
Ir12mIdabVkOrJKHjUOiOYn65PCTvoHYHuRFUahtAbGOwbmPymW292FdHY0+SRqc+cp2QdcK+QXH
fdFfFEWi09vzXFnbpCzfXw8t60oLYAZY6scxQPhZhuSaD8Q8JcKv0q/UUrQkJQpULeXWzODURTCj
DffzvoTV01oMZztlKVR0XM/HzzcXxqsQXqoOhpI7KTI7G7f9Loxv7v2Uoh6A835oxxcMSpC3IF4G
BecoSKuZ0Lat+7irfU7nCabqQ4F0c8BoPxuYxcrqP62/v2OUepP+AaITVPVYxLdJTa2A+oUWmIH/
KYpW72FkDwPReVPV17moK2UTHIU7/GXnpJxHN/bei9Aye2NV88A7oG6IZbEzIXZuYBKATkmj304U
lqAY86TW8mwof7oeKvwhtFbWNPf7SmKbOgEGHUg43igaSjvkyi2KlSJpbroxV85gS1Quk23DQqo0
mvKt3mYX4sVIntTTYyM8Hu1/5epiehTYk8OPHbRQ64uBqJ5Yga1jE23r52Fxt9IR24fxVY8kaSL6
dUyuVLAfFIxZYJtfwxQzSuwnIr7CwZUIbd4H/JxWYgxjO9pa1b0Ri6BOOuhIVC9bFRN1qwsZMIhX
tw7qnpcbrqiqR2VF8cRTrKeo7LvDf2OJsqLgoDcZQwQw0Um4nMWdKTkjALLBSrwxxhfCl+sjdETr
+/ywyIThwDkPGn26JoiZ8SLGVXilKwCK/tuXX9kYWAEFafBvZbTaCHWYgubk0tvf6i62wdrdncEc
ImTGpzyrXzJ2Y7piLRMyaP+0U1LjR+BWUYD6Yywd6JhIyoHMwCYT/7I3KjGpu+tyoAl/S+OzP9/1
vPL765ECcO7BZTMxh98nG7upUwzdESEj6pgGVEQclUMOC9ap7d3hzimUWI2pvPr+XG4Vsyr2DTrj
LY0bDy7E6gVqaxnyz1z/Kahv1hfFcpLIB6LMdp0yYNFY9Bfe/WBaC+QTL3JpSutDyeBL2Om6cE6w
xJEVv+1cHkSOJ9D6W5vHiUVTE49YPcQ4HEiKASWqYaUST6A5azJRG95K/b6c3rjiXrjujNHEX8fH
i5IHnuDuo7l7ustsxpQVxesjOLVvn6YavApxXr9Eo/Wdne2RwAGOHvkAbkZvfSpI1cNhIht7bJkn
kuxIfsWeICBWlzwkTOdZV1RHbgHfGdyWzb1u1OQ1mnxSsDYB+2IkfKbmqOpl7j83v3yH1LXb0d/1
Y9b3I0GKOzjx9W0N2JsyzzSaxqqg7hp+QntmC+X5SWxYjAcZRUAGuFsLIjLNKuD2GwX6fltkP96v
vUa/GQWQQiFEQ04VNGHymMWB6PQpTXdnfGJALyPzQk6J0UZiUj8en7YnrV2fvFdjX4WTLtF72ZNt
tfZhovX9bOnQ/uFFuYz7cENFo8imW1BcrCPJRerxIBN8rWjDtZ7UyMl9AWyGvoznUtL/1QzSJ+ML
eMPF61Thbv8Ct+aAmQxKRLGPpq2sJdMIpFT+B6L7vaUcC+6QHetLqITKCOLSAR0OjzUD4+55l7Do
3qxw2+1xIuT0Dicd0dLXMwO8i06ExeLWcnq1AeBBY73h+2IZHqhPJCxB4V89/ZXOze3LNT6Heaaj
0gyorAWA0HHa6IxEcOw2gcSX9JunnpkbwRXyGUIlY4a9ZX8tOt+WsMX3mqq/mLLroKbu8ddET1Kd
YxC7a35A8ykYw2QVepvK9xTmWQHMTqoGDQ2TKrwC5zrzzMcRNPZJBcRThe0VVKcnrRLfFHTCNTyI
PSeLY8hSAXjyMSmjNu8sxMJu9zUXZDbDzkSyadCL4ww6gl25MsZZmjUjE6WIRU4KOUTlV5DoQ2IM
m8BVTgxIbOcjtn2EpijF0vJqZ71upwzWjjSutUPoH/UW4JOy/6O1E8Sza7PQ+6+NvelCe76ECyDN
X9KMsoNELHucw9+Iy/n4zC9QY409u1gKAQtSInDdQfAp8iTs8i1jl5QlGAsA2jky0sWtJUhPYvdw
nDhqma4Sux+UHoheOQnxjlOidfPRl056bh3/7zO/jiwJAq7Ewr1LQHry3VViaWTywzRfZ1Ir1QM6
zdjpy2ofcxjPQ8h35X1FL7PfGdYj6B/sOKFEPGQZqDPBGO3U8iJVKKivsBAjlHYYeb701NjerBm0
IxoNSGRru6eYk3IQ8hVTyzGdPlbeZtC9M/jv+1qUp/2UVHO/x9wupi0DemwuF6DksIHApnsxKzFI
BC0esfPs2ZH17xVv1zE91FIvA2MvohW7rbAaykELYhsmULgdO9YCzKdtimfTnxVxNqVFIUUZPF5F
iUe6kmbIJdQWsYXDY88QjY5o0n88YfVSLRUZo8eAIMhluYl4y1azd2OElcpCpdIg7UfUS/0D+meX
gSwareCviRv6WY3sgH0+BJgJ5QlsCpjoFkZCClUniv45MpG7EUsoO8LcwS+sELXQmMCwWYCaOJWu
RN+N0WRGg8j9Cqgys1/pTMCM7qT5oxcLWVrMCMOqFj8/eWDawmvgS+NHRRHq6G0u56EAJCv9G7Ix
f93L/JHBX9VjjvgmMVqGiZ84UlUJQ+0+uKXwN27H8UlyxXHFX6R8pl6OkYU9y7Kb6Z7IKrXwD9oS
U6zs2x9NEELEftqYQrpXjHm4xPzFVbI2hVCEq14imyzASZMs10tKzU6mVwvTpQYnYoGb/TWFpkXN
mO8Lll8Qnxw7qxJUS1E9PwZWixGyCQI7HE3Nxf90V+z6qbc8d0UkdJLOelwDbXX4TyulUG9dwFLk
KVxYrwc6461UUAfM/8nARe72dLvWI3QFSa7Oq5e+T1sD8k6wlJgC2chQIVLoRRmVJGp8YW3LGGFQ
6IFEVDlC7Ib+pqQHWxeLn3aEMbwsPu/T15ywJECb2XprhT/AVtKE9/nSnRETZZZeEsp4eL9czVrl
YwLmosNc/lp3g4QqOTPbEhzUubSEfDJd30i1TxrGSqnKbGqZYlPnoJGYceRfiOdoCecTDDlk8Kif
9Zby+L7Kdw5kjQg8UM6xuUIYSueqA+NIwt4AIN5MwQ1pWKj/z/+3UKCeVMz41nGX4HuFG5ax+Kbm
RvQzSo4IpMT1czqezGYj5xcebBqtttUDyIF9F+5EBfbGnaulRq7eyI3tTV1PhPqFQF6RBQFPyuy/
/Um42uNo46WZ3jEP8zG5aOEXtn2W3eAtjR6J7QzXZtMCL4LRtSPn3WP6RlNtPS3r1tsiGeqTwwnb
DpIJzbdZb1muK1BWkdMpb54B/+OKlpD18LsPwxOXAb3Ri/5K9IVWBkH1F/IdFFDKyPQf8RtXxcoI
IH9jCNoIesoYQRn50mR6FcD/07vSYyHVsyINrbVYIHPYhv8yfuR9nB+G+bs3WwCDZfWR7fCDo3QJ
ZmgcxPJVfntXNG/R+0jnRsRnmTzg3wA8ObnyzSHE5qZOUnYWBNo54XfPy0yI+GRQ/OAF5XkMcRLz
fakq0B04g+S5AfRBnmE1V9BDM5kgueX53GrLzu43dYDSmJ3zQpjjvukFrZA609wLYYNCCBmZWFFk
IKyAlhMj4v6xVVJlYi9bliGTi4u+y/WbEuNcHOBQo+AIWqwAwMokM3t7hDK8vvnpo+AWsZEg4mRJ
GbBaiJOA0isOFlRKxDeYlp8B0eOcbfFmpIRsw1TnQiR3CXT7+Sqfg2R9UvUNwydPG3XsKgy7OHcn
tE4/inEAsO7zK4TnhD7oIxes4c7cae3MLj/+92EyFYmnnen2XOiJxwNk2+CTtjrTUvdRHHmsfyH1
bO7rCsgOZT6vdscPD0WVwfpLw4MVWXDjDpXdoqjBDwVBZvUUpAQAfV1T1VkBFi/VtCMWsbd92Jf2
kjOEvES9k64QzbG76WngA3qVr5yLlygjK552gV3z8QEttB/Ql0D6myVWNRd5Sf+t3FRMxnYhRFmn
9MHUgnTDFQ92vQY2ppf7OuCk5sdaSy33U5gGbh34vGTk99YcUq4P+ltlBfMGrqF3GKZ0xocZprjr
7Zxu+mZfEWqmIg1BgKdBhFat7wR5k+GAQejoNfrCNr2No8NiDofQ7xR9k+ObvltORx5NDfs3V7NG
cQ1pYK2o702uc6nokGF/eu0G/Iyj4C5OP0cmi797gVkes/NxyNnz/TWVPpWHNHx4WKn3Y4G0Bm5R
mdO8qHE1qiYkgNpjsC6fRZ40iUhcygeFhsRuCvVEPR2RjL4MK9UcMEc5c6JbE50dfA2PopcsQI5j
PZqlSEqtN6kze89tFDU0GIsxeKmrBd9nfEcnoBIiISDZCLMOstSn/jQnLk679M/nEC78ntnLaXaW
L3yq0Dh3TfZzbiJXfuL5h4IvgcS8yB5muyLjXu+Vgzt7NvnlBepDdlt+BchSxpCWBCDG+J2IbiEu
lS+CGgyqBeQJ+OAbsLGDi2Pf+3wfW2dzg0SqkBp5aqQsDOy54WMOatVheMvyZaPX8FgLa3zgb/pa
KOjwYMoweviYdn+bLjUN2A9oG8wuTPXQoTQ1Xh671AFTU45BgnxLehOxSeF+9ceITKPLXLrCD4rx
Fzd/1oHBLBmHadEZzswNCmb/5JYEak1hzvesCgJGheuYUSrxYwMVj0q1YLe5I6ruPMwnydj/ezCg
iqak2FnfWXTXx3YngCchaFqPLNO9rO/JUmbuueqbVKy2XWcgQoIUNlH+fULkywjU+4Xxg6u/EDAV
cwzZJiUrKLqv+aVApmbJm53+wytiWH1V36x7H2OU4RLRRIBk6khXn5eLf/hMVcMDo24s1dWnxYuH
WT8MwpUviEh2X39JonZTM2m18lTrW4Rec/6UeauJ26qgsu850QslGIwN2Z+gOd6n7EdT1MirSZsU
szYIpdsy608sxlJdocBoURSAXmTjBAwnM0ztuA6BP4gYCLwcFVndUZwhKe4P7M8t9j9KqpXVik+B
UyuL81ZC/RRKT3cUHttRfNWd1J4MH/+uihpaiLsZI7ZRnr3howlKxETosFLs5f1V55+FW+OvKcKW
hfLhlNyWWmhZcvOMi50/4vyRyb7CcrtsdGzlnMeKEriC4iBnLfhKqkPCLnmaddZmTt5NuInDPmmt
WHavoyXkYWoLuguod8cvdJmhPbwAzrG2puzu9BQijlICtPXjvrKXZXTF6PsFykC7d1+aSI5qJGf+
0VrsSqJonmJAoIMdQuSNRW1EceyFq9Q4xYDpUMcNaEt7fP6E2DciZvTrPr5GLnV4YAKkFcNgxORO
yWpFuGQhtOWSs3hBJOnFGfsfQU3MlvR3NooIRseGl95E0k5cGzPUqewlBWPCgueKqA2zVr4WzhIf
lxg3toNgW2JY0Wv6bxeCU6YCOoghi5iHKXK33dZRRw3mjIOziZDOs+xnCupmnoMNwg1J7BIVtcjF
Uz1FuxRwOtNFx0yoojwc9bwF9CxeGslVvUegypHfcNbvcpakb42BEPm6bWA80ncSzk7HCcuW+0wf
A3h8zDhIcsJlA+J8VCpOFCiL/3U7X1hzB8ncMiMVy8MukjHu8KOFt+LYjFOSmLXn25G3CNuVQQDi
gaT13PEYQTIGmm/8AmsoOv6vlG/MUKL6KJ4TH/TGPTg5qqCO5CsplydIo78zr1qaE0m8vhNHihqg
7gV8nxqD6C9AFkyI97EgfCY/JBK8jegEMox3vcGHqUzW8gzluxJCAHuC+VceeaqlV/XsoOzexRVW
uom/tI+UHYOhauu6GrbwGPJqdNKj6lhvr1S3EGpmiocElVWV23eVd7/MX2lLz4KExwsvdFkgq0mQ
pqZcaS/6n4QLpJdfMFEuuBcdjHRZqXEYPdUX8imC0ctqC4mJ1ErJjZ8AnScVNguwgPSy9oe9nFAx
lDlOgrq4dJ4FmX6EDwMTzqR6IUSB1wcMb+VJVrmnW67TUNxD6Yu2F7XG38IBa8y+boZ72ah1RFEU
YXbkZWTK5zjcNKFs7bfJs00zr6VD1FOj8327Hph/QTWDxcKxnzgy+IfDVX/Y0xawoSbGD3GhhWwW
cIvLKGZDkpFpGdjHeLI66A1j7GxphDMZDsyJ5Ynq9rdb1JRxgaaOl3/wsJTioNNaB9wPOGzBHCrk
kTZRyazwVB+Iq0rHEPBdWi71p0umTXCyQ14Cn2R6ZvcKYPoV8b5ZRTBXjhHTBPvEayIKWok2jagu
UxOe0SVZTvFnT8i3klmNdmsrWxiLnNFakxctYFAgMfOCgehidqVdTehpXoLtFUmht1qkxDqYaAmL
uoAmd/Cxbd1OkUGQIEVyrAnAziyvDOqd0r22M9cEcbzLag3GyVzq8Sz4H41wpr7b5zTx0oRAkbKJ
smdq8Mbh5OrtfrztjjBRj8Wws0LeaV4Wno93b7oMsyJm/F1JJzNvIEJJFi+ITfjok8QfC2bqFkbJ
TjuSpxXTNvholNAVJvyxi/RBQ4o+RDRaXK/t6WY1I6YQg/4FGAKNLojI1Eprd93N16/ImatMG5qb
LkjzkpmpsejzTuERB8hDVjo2aXZYH7LO3/zivODEeQ2igRXdmNuI5hvajDXM88GGvUtpQt8fg0Ik
0tI8/EhUVChxX6p6w19KQkB8eUrOL9UY0YEh34xpXWQyekdyGEEB//I3GIRq2C3WVsCAl2dozK4c
ubAHUuAgd/HV2UTqspg7f2tysB1vh/48bFN+H/FcyfCPuppH5dtC09YAjpFkgEvQtQVO9q4GrqHW
qxRAnFVomKl216zeoiaaq/1WKxroEqsyRcANR5KDWTh22G/rrFANMV21rVmbeN+NNi0E6s2JldVk
0Lsjbnx11p2IrzIZOAVQVtC95TmXZj4EAoRkoswpBhZJACHrT7+6vhcE3EtMY/hKPZPauBm1QCmN
nrhIiHYVkwIU1e0yCr/FQs02CDchqGk/k4ppqtkFoIyir6DdAiLAjsO5a38r98fzwfKTpu4a0Sgb
qxfuiQGHys+bfPsSzbPXOYMjmWyw3dKGgJoqkqV5mqu2vR2WZ2noSw65K7CWpPiJb5GkHkOWA0d3
HPoBUMPvxlY/lKY50qRrzhv7tDJ49XnR1mVERRMumQfBR/HJwNRP/p33LGyZRozW/T1WDXpNHxQH
mwYLvEUSzA/QQyaHtiX5f7LceEN6+KIYtPCd/nCSU7DjAqf1Spw6TURu6EDmcV2pJZQ2Mf+xHO7p
mim5Riw8Fyh3qFgscuNLZTaenJw0YmVmGMIiE2aWq0+4q6QHReotbSTGi9+Kc4CglUt1gYhZlWwL
tA+FqJRYJAJX9rLZF3XHTm/4ZCideZ0onO1lKddjj2yInPFjRlv7tDlFyNk8GEfJHp1d8WDlOKKp
dnZ4v27/Q8ezVLta182uUm41y9ZpT469ifXMLEjPmjIcbqyb6Mj3r9v9HEbJxDZpFIHkBL62mawd
CPFTyaWvSi5/rilHHDRsoCtF4cdLINMP6rZFKTezpF6EmfKdUnc2mYbhF0xhrXEkUcgUA/0czMD5
es6BthOooQCB6g9Wp2xzz+oFtcFRh2XxFwR9Go/3nKHVnH3uL/WCr1DHPQikMMQYhRqJmsp4gznI
P5nxyjRbiwfYlufI5ClMvCaFyZZm5xlSylTK90uCh5cs+7CM/9XUOYTUPNP2IWA3ZdbKa4sNQxVa
33uHijPQo+q74GsneMBkvlPBGBZb+u0HyU7g7CHWemH/RJAAS1MFZy/X5Vq6UfkAp0Lh0DlPmHog
3i9WpMarjdDxJgEpoGiESWAyvGP08p7mVTEVAb3fE7Ck9RgMJKYP2WDjHlnkfP+Pwj3GaxKIOYj6
/zPsZPj+m5/iAt7kRP6bqjc5fs0y0bSUmLUQB2mDYpZtatQCZWPYASKR++/q+7eazOi9aNQnFsdq
N56yBDNY6bbABbvSZjZLqw7RlSUPVjJbRwufR75iQZuDr8LI7NGRglC6kJ+3ps8np201dBgeW/T6
1Jv3tH21Zku5SHvQsMP5Q4NXRGfHq4u0kOhsto/4F9wjNCr1rV7unFbujlhBXnz58uNncwbcRchP
mIl15elUbShW02ywnIB2Uett2EB/frL80gO0eh7D8nx/h8D0wCwLiTBxETboonU+DRF4fKeyZFok
ckJK38sJb+UjHIKJdHtg9WZt4FY5MpUIMX9T4Wcrbn4N22P0xn/vWbsQTrlykpGnO14rM+fH+mpP
p8jlo8zUAbrjTL5H2V2EL/oRQSwKToeDGHjBLmz4e3LPU7maAgqu6IXQzKwZ7P7w+0P247ttTw4l
xwnF75BCvm3rFw5XJqCCZy+BkBDqxVD/lYY2yFCIWqoppjO6vg6Yr85JkAiMXwROZFenknrPIHUn
C24jEiBmcTkOthbUyvJNWRinFwhHSGIu0iEFt/7DnDQ6FjzGZEWDnPnQn3TZFs/PTtNuMZKIqApx
0kbPUa6P/4XlSbohsYeydSpABkxdpENjOLFQ3YGSoQyvja+nm38XDjqY18SIKqcZJ2Hnij59XrLE
1bDQfmEUbgY5VWnHNUeHVBaK3GZyYv8HjYrLGQfU5RUWv28DEnCu+hv7tx41NSNUqNC8BZRXecyF
JSeoBiP9LgapNuIMS/6oBo3XyB+wlv4fVWI4vSK2lF+WlBrf4roI+Leso2ewOBulLnF2fYTcHTt4
SvxA3NtuAe7RE8+3oQV/DHbb31umX5+LhIFkcGkpbFzelGzFDgI9vFJYw6NylEPhZy+IEIh8OHwR
noFl1GWz7sN4ZFgH30G7GaHr2ew5li10RYgTueQoQWEe6OW7+Qo44MM9hyzQukTO01fHtXz9YW8d
weuTIiSOYwM1NtrU9T0F5jaSb2rgiJz0YewhuUj9qcdZREaLw9MgnEdg7Vexu0DONr3x/Nq0Zemh
pllq+nmtQyRPgSJw/WAbmhnavB4VnrR0+9MMeLNr0Eium0Pq6rWZsHbmLwiXNVEU5vqbRc5+vwD7
m/TwqQev1HQUxSC3LIDpXb5BG6ntTAj/XG0xE+xzQCNvXPxrsXrPBF1y7czHAYguBhhWfq7K2TQf
K/fE6ozZKww8wSPCVw0jxTfl39eyM90cEkqHgocdJLpJVHFdN+ClCvZNPQUBcidYSMWwOAMLDL10
LuOQ7eoEkwHVXDh6u4FuDnQBc8qkSxDo+MA9nfTDvR19eGSwMkkVZV9Ncus/pLw0A/aFfWwiZTQq
j2x06zDYFtCgm1ukoc0x9MJrk03ObZpTC8PBTGD6teY7Pdi0kT6TOrsp85gNdYX302PQz0m4LgoY
xTlqEdbO6zhnQZt6hwTbzJOHgtgZ648ir942TP5YMIrCWpzqzXCeTsd/c8utnuH1oz10OLmqmrBr
+wYbaf1MDEbmTQrP/M9mm2oLm9f/7P4XwIkumG8hj+APq+xn9REUNMc/rO8mDt+g2Th7HYrMyo0e
v3VoQJTjZVS0oDVAlTXNifqsLFnFKwvotLWKsMXm9/y1FhSt4XK6q4mzu2nClZzNIA2L1MYdaPO4
l7EZEZcomdlCF5oO6me22lfDdbAewbIKNq/k9u4FekHV0ja80lzQnDVGoz8A1On7ffjAwqA100uf
z2l6MQhy58wy+KMwSuYWU3cvGWTolN4V37WJUg0tE2UG1vUaSxKjkxPlFFeWrfuKSjCCDpv/a0UJ
jpiZCZT5gb9ZO6FXq1/W6D8xSrT4vnFp5Au2Gr7DzIVkuKHvhy3YoPFUqVzYz2mIZ+Bj2A6xI321
M7XDe0Lj6xay13yE4R3RmhgjVq4tK1BdvAV8GKWL3HMH7W7x9bDiyQ5WtfxK8zIu6VpE0cBROuvg
p1JayTJdQam/nxk+3vUjMVMwOfVE5Txcqnj4726i8vXx+aj/5qpy75KrU/FFesFs5jxEE6ePT4JV
nTWeUNf1JWb5Frb0prmO4tQqcdXdm+fMA564EPUWQ7ro9Y4HHaGmm4j74HWhkrX9lvcLQIYqPRBC
P3JdSMEyjelYFIM6HjxQDeIdsyKKUFmsIBebOGxBDI9lsiQSW9H2YhtAKAIO7XrbWNuCaiIG1ZsS
6q8/jyalC0wKz9qb1kH10ijX6Tov+LmgXmKe7WLu069c1neA6KU4Rkh9uz97p7Cg55vwlf1vZI9H
q0S4pL7zNmog5cfRzPmptPz1NF0vO1SS++i9frSXaVjrd1Yj6Uyo7WZkFbGVRan+LIchMzPgZYLD
3A1mYAVkRl2oCBt92kPWYkafafUCaBTYztbYk6Sc1byY77/g7GtmOpKcrDspwu4Y2lcjblTs8hpy
KhSGvF+q5Z5zr7Im3Ol48PyxsaHk751Ni9lM04ZgDhpeA/AXqJrP72Two8lGiDBH9Ze19UuFTnns
A3cy7WNE+7RnFoug9Kl3oVG4u7KWkbu+95DEWbdEtdyDVGGyq7QN4b2G6p0BXbY6UAgodWS91Oo1
Dx5ms1pBtTsjQc2hqc0Zb2XJYRVHF95C3vNwnCFFeQ2QKVJcwNr18tZ8l6qZqgaNJ9KVzQ05xRX6
pkkqfumjegyQvJV6MN2+e/YdZjMKMJvF8+Qg8pyzXX/iNYFRkUPv349GlhxYw+fJDCFSOlmvxj4Z
HjdhVF+9tuPXipeK5g9OpR/vaNQ1t6M8X2iiieZ/qJOzpShpOxWbOqaDNi7sj8vq5z2GEg6lIkEX
egcDIlWbo8filtZDQq8TUNmjaEF2+T+HXgBX9VmfMZ9Ubx5lNeFD5J52BZvwpPL37KsUwvhJsrjz
CdDWuZ9g+29HOZ5kNxO99I/0VhOzQ2RF4CL/TqroABPF1ur3NPLAX3XVOVOH4tktxU6++xlN6bTR
U0vV8lvBIE5zCjjWVufcjFj1236YPdly5yQAej+SZ/5rYBnGuamA9Ak1wh+VpRIzWPfzrt79ZBh8
feTCRe1HtqxWLrdZMQrg4wLRYbTd+yJFRwygprPxWz/GRxySuQgDUBw00l3Itg9U3rNiU5MwSm/B
bomqAFA/C+GnwFoKj7S2Q5UOolERO8PbTco49pHadyOmGJ7Np/1m2AxzPdgNpRdkQ1/j0u82F9Pb
IzuvAseLAZEYWD3Ms9jCC8Rh//uIyd01a25d6lW0NjGWnaPHXsfu4heZUbg/7vzi3JJAiC1TFdED
15K1AguN982Yr6m+tVjR0Zfa1PuI3tC8DlHZ3FcDV5SDor0EPqmHRS50LypFUY/Up1EJ9iurDneJ
2pGx9spSV0EFB6OdZiUu9G0CFjCjoe2jwKhhs/JwuVRdFQLbSz+FpOSxtieYSMFMr531eq3NH5Nc
NVwabmtKRisZJVYrmEN1PRzDrn1s+1u04+YnnZjenrmbT2PsmfMx/d7X4L1RolG95YQbmTtav66L
wd+I8gcynA114MUvjTz7EMFukiZ2tYJYAZte2CxOtsgt3BwYso+yvj9F1OvKVp9yux+T5R7Ja+Qw
7WT/7ZWfI2sSNzpM75gIK+uu3s1FN2h0icTI5rzPkCuxTvBoOuXui8Hsmr1IjPV8RAxM1x+6laUk
OFpPNFiUkqldm4T4uhx3bQwF06i+KIX8QnCGihArKbvYUnhyszcKThUGUb6ZyvrCAFCaSxIOwsA2
MwoyAS97SU9Xzdkk125GpMrfCLtUGU2CMuVjQQeb6yyjVsUph+UufrMpt9SCV4kRCQHDnFHwBfk1
3Wxxlmmt5daIwZ7VEC3wLHIAZMvB1Wt/Hym3GYV9OO/y8wdi6RaIGUan9BmpwQ2obo+m836X76P+
EA7aNtkC1uWVOgrQhIJxZundzvV5uDRnDNi1wEabhqOEbo16bnb1Si0AP2ZwlG6+XxjYvcK6r89T
K6t6REl3YR/sIwZpugasHtZIsuW3OHDGnTITADNYijLL9+xl3FSc4QX9X5aAHedsnE0zomKWzySm
PpeH5tharFbmkeK4OKPKFxBa5XvAuEMsccAy5CW7IzER6NiXRhGwnTCdiGN2pgtDzxycbJUMd3i+
hG78lm6WHC5pPtW0/KHWFG+WFCibFrT7G6WEFrmmcXkDjbfZBjHxU/XdHexvi40De8coa83DoTLy
svNm+MkI7D8a6KZkxib89SjSglqNs1b7kqWtCCRhXP582PnXq/Y9DGNpGk7Bm34f19yxZhf2HsJg
ucesJO/OegbwRMIF6r0LcAZZLEbZhQeFrXwie2DSU4Blb4Q4rl9wu54t/OpuC691+z0JCPufjrs1
FcWoZ9Dpeh0aXAhSIaci1QLZ6gBlgebqPOSiHm4euu8zx9m72IoaJPhC3LB+D8hVsbRHSH29197c
Q4+geSWUsghOagLIFJvsDixLG995fs9P3YumqvXZYYuCnT/DpQsaemlA7eurhkIm9MyG/DndcNjC
A0Z/G74Dt5guWip4QfvvYwm2hf8pDVPstRF5+z3ZmTGRUShpzBOsFAKgPtR7woaH55/UGY9mQpOh
5r8F7M3kIzeVuTQDBABDnwnvlcPPidFu8gFOtTXbAm3rlsAyhbp5Iu/OgdP00S+C1iS5yFdoowZ3
ZcRgP7Vz+XcBpZOsc4MMQ/Ul09vEWu+/12zm10yuAjWxiP8/cZFv75IknC3tFFdNCDJCHbdB6hkh
em8wZXlr929C4UmrGrI/Hk7DJXrUJkgz8PISaDD68kmcSzcC9yjU2q9UFru0uAC3puG1453RnC7M
uzAhU15OV/NuP7ehwAfMzvbmL8saCW+9BlS25v62GL3q/EHe36VjYao1d6RoWfh74fnzcR+U4P4h
tlOnhj2NIu/SX4qY3HMPw1Flk+lE8SvnhJ7tKu1p0EKfPFiVRahwoWyNAm5a0TYvbJ4r/9MeL+VM
qctEBIazPo5nyhlhWrgYysuJuknTvY3NXPZVS90+ofgSZWVtIyXqhG0rDHGfuY4unBKzKgMNVd2C
bqHxoa1x/7cGSXfvbsCp44+LPLeuBeuNX5bZtsOtHqa7i/AYaEc29ERwAQhksxfnn7vucX8RKcTg
7VVy6GLheWZjhBFagSbmhmG25iM0/YRgsRpU/MiLRt0OvftQJWUZRHWeIP0JdfQSJrDiK0PJcUXu
95MZJSBgBlcBaOhVKYjy+n25/r6sH9xiT9v1txP/0P1pZ+9/rCAwafIr9DhTalFFPH1OVVmQI4NH
XI7mKweW4BB7wIS+LfMX5JHQKZqTdpA9WVitDUFPHTxgifn8L4O+elPNOFDYqQ3hxQVvnuxkBWmJ
S+qtL/z/Hj/rbUtkrJtNWSPK/V0ji3opA3MYRmFdvD3UvdDV3P28s7Kz2MczeRaofRXQqCBq6zil
xztD1zUSRSUhUvJXM2K36jeiBk/QiwB0oJAR/voPfmYIRSl/MV7BkI1jffA6PO+UKvMywWYE8HRg
4i9bGBHoidGmrBIGSAe6Gziu+VOh+gfmfoREIhPQN3DxWW8SVsfE/UKcKIJnVNYJjIJTwP9LkhhS
wJcu8rBKMGHPkNUuVzZ1pMC8v08dLylqWdnjvq69cmgzXcLsfTiXwk2j4BQwh473nxlWFIFqgcka
3l1Fi6MZFKzrR60TF7ZPDlGyq1795EwTjgmM4xPRm/gPmSdIpmfju1TDMVnTjhLNyY2CnMAXjSLZ
Vq9mr0Vho+Uy5Orza+Vjq1RydY3p8sCOAV+vkkEsTn9bZsFvtklT6K6w/yZjVdNzOQJtv7QdNCPX
ULYF5mWaC36twzrX9pHbJAQHamS+BH4G0Ll51TJwdaIIMNUn8O/AKBUA6YgsCX4pwXPWIoYD+BMK
LxY7oBzW3vxXLjHV1FX0kFPigwSmJWBVgdevG5BmAzEJ9IHdzwgw4P5/JcWhdYal5pOlOu3wwpB3
d3lfPMo719798m1ZB20Xywxkwd41SbfDo3kqVMnFI4IvdHX12keTzmwNVnYTxmN1utHlzEmq094o
NAhbJ+OH4wVwasFRWM1lcf2oJ5/xSD2/3Prr9bgl4cIIev/CO9nwmP9NhhbEDu8IohelwdxSMB26
E5jAnedMQxrUUzJK5cuodCogKZDXQjnniN8k/z7kgMSkPYal5yJ22kWshx62eLhQ5X/4kCwqe8Uo
7k9PLQHRBVXxFnZWLw5HK54GsiPjApVHBl9YdFggzgTGuLsfM6U8S+AvQO95epZppst5kqVllbw3
vSw6Bp1iBn4eMf4GL+nRmP9JKOH9ZyS3dGk8At2TsHVBbQ6oC5TMlHIsv4qzW9k29TaZG/av6s3u
5+Ceew17hXMYB4IPkyhslgsxCGKVSrz9znSnfsKS26OeMQjgge3Onias3cYU8r2WeB6W9d2auRj5
asqstnkcy8xjB/JpncUYc31pAx6VfMR1LuVSlhFW2M28U07g+UyOzUOpQDx2g1hWQjh5YOoxaWSF
FwI4M8x8mVEyDIRI3gYRZE1ZGvx5RrteCPP9lMgwFXqkEei19Zc/khLavnHX/P9bvhWRL49qikz6
Kjp/jal6q1HgeF45x4hfz7gmxIIQ4myNZW0urgxsufvB5ybfKthu/dZC1pZ7KPcKZ6nrXXwmxWkR
X3v5j81rBfY14zGZXoMyJRTYBVzjoKvkurCAqpSQvUZzxVrCGPdOYSmJwkoBuYXo+Yt1pZpUK6aM
KNSa7e/kY54Pc6aUGyzSpeqO9twccwN6NTt+zzOO4Zq909ujYAGNpJ/MOpdmL6NOF4eHfjSj0Czl
45YzJv6ov9IxUZ4iHJGUk0wyCiAsOokfAmwcXqrvs12EHpBzAsCZ1pFEV1TbLKtRywTrVS+qfnLp
lEGfB5U/SGdtN9ALO2bOg2FIRNSQPOH8LG+n6dMbOLXt/0FDP1t+vXbp8DmcFdfXL53tDJkOqw5B
8XbmxRUOBHukJvyrSjtL1u1CWNO8Gh4Hj2tFN8jgYVHJsJcCylQdlqFBNI1EqcB7CXvbj3/wp90n
X2qL03OdE3HzWsi/gENZSX67b+vJvY+h7T3OYK52SLUMudStAO9MK9pxeFmZcr5dCVfX75DuXUVs
Q7t1xGkucDT8TrkU1nBBMSm0I4fKWhJi1h2pBJIeKxUtY0wj059MsSXPlWwC1uoWQeRzDVBNtNv9
sqmUYQh4Elc/QdagdKGLlbV7yT4UiGcVco7RxfN/qY4Cmct1Pc/Ez1UfF9+/UREUqkynzWXuEjBL
2m889SN0q1inQ19aY4Ps2UxI4PZoxllMBkcorXHOToGp3c+oDm2UzvmDK5X4ZgTcVtOlB3HIgkUm
uHaEiBfjOmZ336a5kRYRRW4aLbd4tmJoQODOcWUYJUnQ6nYvrQ9W+yhbJdFp6uEqeKGAiN+ts6Ng
mpkZqcstZnJNI3CFD+8qMs589IK3T7Ehr6h2PNnqypCPpH5bzlnystvDFNHhsKutUslazSvzp21h
VUdWaC3tuBloLYIe+J4TUKSiudAEV0zPLNcORQRnBV/KTEnXLYGszcUhiuXSGFSK9718fpz7u6ZF
VXxVEVWe8VuV/VkA8w+AdIaEKqLuWunNUVtlY6lz27vNSO0MOSJTPk7SEwyny80U5DvV72EJ2DCu
wR/qyLlES5NWffU0wq+64uEM/V2v118FkC/rsLisZKUtVTIujINfJnZ7yFjh46uqVf64LL1Gg9M2
3mCbehiBnlR5+/sc4jtacfE8SHLvbgeqyExg1nPzbh5LyBO4C78hDsU6BZXk+qt3VYb1WVCscB//
DqFJmePt9lInc0BP4djNH3g1KUIuwXQTGaGPXcxsPw670frY6YPI2fX5GPXoB24pg796wBuCoeac
ca//uP1yIdq3fSXPeoG59hLt7w+6v55jMdZG57imw+XyT8y4HzvG9pNzwI9ko9Fte61Wq433GQwg
vF9bX19Cvs3VnDg3TRSwq0anTHP+0lNWwASuG0gj+LzTrbySb2Vo7A2yIAob5dhemrrcjVDBl+Hs
YMZm/NoIZaoZEAmSqNa54umqRUonhSE6i1xi8y9Pgve9+R+OVfsNVO5uE6zbh8EPDtJO6l0p1q7u
XHGTM0L45F61SmevkWNIW7vKqHFHXh3jUo9bQ3gvdQWrhJvEPdb1Vs8gtoOEnjkdujzdS1JMqZDu
SXs13thlOCYQACGRTwm5u4FhOyVnT1//WrZUBJ4B9jrTSij7mQuVoiKGwjtwf5ltB2HfzEsb2vIp
SJ76jkfh7+eC1g6RePK8NnVCm4PRjQ749J1gEMPR05SZ8DOlYYCbqBTwG74OUKGlWVSmmCe6Q20R
cN9usQ3Q+jGh/LVAb+YNKYvVEnUFfdiLWAjtKJuGZQZoeUdzU5Z4qfhlX+m2sKE4WGePlmGQrE1M
OYy0MJhaxgZWDygHJEu5ffVcabr8tg8W3hBRlOD3V0WcdiBcyST9TOQ3b6oXUFD9Vwrd9mKVod3O
ElGh6YfB3p7cNUFp2+g6Jd2Yz/vCFm+H+APP1PcVw3GecZed/s9vKu04jz+5bl2U/03f2sspIQb6
5TFUyh5NxIXMPvfIXo5HaddJ1uPCpYA+wXGwDf2OAvZ8n7K+tbhEfrJtnyQySpABG0kiygDpjOyX
5dWS+p2xfzjxo10o4SpQ+08LV3zGGFm33N6VTdFPdW8suGZjf72ZtRBRqXAc7X56lcaIhWY0amVy
f8TDiaSdAlvrLe2BaBjireiEUmuXsTD/fUteJtn8UmgfpjRzmtIucMs8W17KjpGbjPJgLCshp06y
YBaTTsNgzHkHnSW1wZ2vHahXHLohJBGr8TOmGF2AfVeFISEVdZJUkw7CNaPKbz8AckXBTGogrbC3
R6MGWloKRj4PWR0BZ864Kdtqo5o5bKDzA28IQsExDGd+9db36YlpA2DO/icUNn9FeDD55r33H/H/
EcV7ZteUmr+EUNJ09ZvkHvnJClgL+/nlgGJBLb2qkl1N3hEozB4XV2hlungzCykeM5V496WcnsKA
B+6OuIYga+JWt35/S+VIR9s7z6W6vk+Gw7edpBPz2MiexhYdsdyiBgdOOfJy84KtvHt5LK3bkoYP
L9kn5evm555Z0u+/Nd4GfLvuM05LzF7VYJyhN5rLqJPHHAGo232q9Am1wbm4JdcPKvAz1R9Cu8NB
38WhI12006QDp26+qXCpln9Zr8fYc14REWhp6wxaO0nn6QVy7mhVd22OE/ZP0JtCZ8DoF+hvW5vN
LKmNDaB0BUvE8eJ862jqdx7ylkmSzigeKyE4pGo0exbOFhmwnEOWT0LLs50y7jIwhVQOkpHjYF6E
gljryIA78ICECSedfg1futZpvZHii6iRb9O9z/MImT7ucuQX0EG13zm4kTMpskFZSGlDvPqWFLdL
CpCHExD+RsvnvFICTmn/bDgseT+5B5X5jEFSjfPJFcyvWmO2lvQ2gnKfOWEGHSugTwr9ttq9nQp4
/jetMxPxhJY+DDYNqdOpB1fRYfR4tCWGeq+2+5pvIfPMiiOtxborUaUDfGpnpf+khq6FwXLs6GBQ
i61AxoEUfNqmRcjkYQY7lAPf4pVXq5twaSFpDwrLqEVlZSE7xrv1wfx+vcLFTAhu0fyo8HR8dxrn
BayGtC8NYY8rGmIzpGz9Oi89biVea57QAJV/sjA1bZDOJBMActlmyBtBSRrC1OPIliwaRF8NYBEe
al8qzTCt1C7WcsKXCwDU/8FXbwEHhpvQQaq0uqzL8iu0ozil7URAQLC/MNEdAayepSLCHMZor0Uh
cY3Wax2QS4p1HzQZF63j/68X8CTCYkypBcF8RpdQEPm5VzqIHLfu4QjZ7ay8Gx9Au9sJ9EkiQ5Mz
iMzkZsVD51l4b02gEd4lgrODxRNrA5XhZjjgStK8VjRU2gaufhGBo1Ju0F42lmFQch1NjebcPgok
TV7AMx2iVaeCzvuBjSsASq2bfuVt4AQnxOVEK0iUYHchkXZsNMqCQoNj3ZfPtK3KtezJ2QdoZb60
9ML3KlgO6ctnwE6miJ2NDkyA9u1grYqNcM1wJbR7Etq1DCYM/ZKc2rH2KmyesOSPlVHLcdmtWs5I
W1XfDTijlS6XT0t2XOzSzSCFrP8/mV7CjgWhkPxhus8yROhUB7mrayr9RKNvFQRRWBab5SUV+9yS
NDq784IECeLh4IuHtwEWdrE1WlaV5AA7+SQmSv96uE/Bk2dWKMT95s9ad4gKSLoF4xWp7E3RrU5Y
RBwILf+rskKESnlIxqdHmmRbEOcB7ljYMI27aIy+6yNriBRh7/XbwYKGa8+MAkV6z0lstR4LBjVb
pxyiHaV/UFqCx9HNg/PeVZQqV43B+c2Z1c8u/Jvdi+FKm/xAJSUPZispZSE0lkVZ9pyaW1uMC3lL
hl6jrz5nA6hsRFlG/4+7yAAabDOb0g8IwiVnrdKVl/3ohM40VHNxi1oWH1gTTFFVAGygI7xK7PkK
QN4C3SRtGxGXG515F+uh1REJZHFaGbrgiRHmUz6KVjHcayH7wCTkytS9Aimhw/xpkoJ9N3ET4D3c
ZGmpD377NJSsbNasHXXHE8mliz/VQ2VP6+P+jIHB4zeAw9hxZOoCwNVBU2nSYzRSE3vaNQ6cY5JZ
yLgyU2GE4GW76L4j1A9SoaSYzGDJSgyy2bvn84V0G23XXBTfIQg23UQC6wXna5W4qDM37eDBQDlp
jiPYAG+eU/7oe7ZmSILsqDIiy4JpYXhfzW59Q91Wm2FhvL7CQCa++3AhZPwImy2sX9oMkuEjcn6I
m9wKG6tSTAsr2pJ6AIWwvdQ3TDW1n4fkblEUAtdcV0tbZF/ewGNT6DOKt68DTv9HhPv7uvTWC8/q
77tFlLpUWanmHpc/rHb84kCBNnwJYwVb9f9wLJID5pVYSuyk8xDyes4nStjp7qhLD0nBh+x/ziee
XNQmsGfBawBvpw2VCjovZeZ82HXW4+4Eds9ogyEbxXf69Q9GQ5ZB/H8J1lTsQX8pFRn+uGNT0rIs
o3I2dziskRBgUIdG0ZBu0rXCCmi7pOmC7Fo9VeqhUfp3oV4Dx9K6L02viCEkFbXDvIW81r6fruBX
amRtLbo/cFBH8J0gOP1s/rPNBj8FHJQMa6sXKMde3EieX4pcMcxd8htSn8fxjzSDj27NpWPlw1Kv
RaUjtztbbtmgqyeoAAvg3jIvDlNpPZxALyx3g8GoKSGMaSXgyzA1ZdL20NCYBhIFnIiYjkH+lFnW
IpxhDR14glMoTwSxbQZl6L7mwuzdAKU4dir6w0poIyUY40YWgTMRTLbWaVRP63LSJl64lD2owwUM
Paqg/Yj7AErox474QovJ3q9cyuTwFCDwTZDjsWx7LPgAamI57klUsvLimTy8ZNPELdMISOnXK7NZ
FjGwulkhfTE9rnG+MguAn8KJ3F05z+HxfX9zQX8vHZi/9yMHSQt3fEGPSkDwrhJKjRHeEi41YfxL
Sz93gJWYe+KFd7DH5n5t2opZ09WseR+pMTVUBrZbwrXMWG7PLYgK6XHdCNCOWkvKUXaSTygphBm/
gbQLFBjdT275my9wuzLgQ5NRIPZlwyRMSzvRcVyq2ZmWa+QMeNXOK5C+vkqZJgS46LSF2nsqPISm
6eRB9mczdiGfkQ/BQSg7LCwa5yE9Al1YbGakBJlaiaWkEbD57kT5BgRqz1N/qaAp1cwJtVGVgzBP
M+WXCNy8xLIGtu/bqKRQxkZvvcVGqBVafXMnOlbchKIiLP4kb43r33tth1cQZZipYOAq+hXggQ+p
ER7T/mKIk3xT7d0NImEjC+pPR4Nixpf0vNq7GUwLn6B8+ze44Z/ILbOpGtvpvElxACXKpDsb+PIf
SPtEsI1w05C1oypsx+r+UDhZ0tWce6+Feciuq7pxrlFo2jiQ2h5PXqqiEtniJPuSQroRMcsU0DKp
kZeT70yjLGYtZlupxgDEqR+np+vrRDUJXRwlGgWG17ytp/zVnZfLD56XyLW3rYIurFFYoL3i2ao2
OmqJtUVNsk+mwKSpuzA0VGMGRASxYgzWjmzjJ9ty2KtO3gHZ1TuDFS67ya2pJm95yzDQHj1pZHjI
wJKlfX5GU4Xxd5++/vHCx1C+AGAHzoZUWMoHwHi9kkU935NnYv+JYYufvpfURQQCPF27sAf0Lp9S
wn0CeF0NSz2aOttSMaW+QW6xTZvb90k183KD+mmBkSdJg9G1cmx6CLEQ0d5qT0jeuD5tPW2M5u+A
zbDttvD+AeFAAYaH/wZQJ9SUQIJca6JqLhIUXdF9zrHz1r0wcq31vS0uVupSu+PBEgsW5Fn+hSUF
zR9P607hSWnlHbW+MF9+Rk9+sl9UEHcXKPlTUvcGyHLH0Qg16S6rZm5+VvCYEMpsrgFcU/fgsIv6
GaPaztJhPCNESrjPnsSql8sE6ipaCfUZevHsCUD8aYmXwSvpkBmtd2+eJ0Ru4o5K2rMsCoso1RMh
kCQC/vH6fBRl8s/RR5JlNM38PjN5RhfGmqi41oyD+coY/DUOM0Uy1ICSgp0sf+Q9lEPhFqABgvZo
3+RdbeV+1rUZcMN+Hh8Asvn6ON9inBEDsAByrZ0XDsgSEURXfpe6BEraLEj3huuefxA04TBVrDuW
SlRSfxJbO8ZJkbPgwwyjFgwTSKRJO9WEeQLJS6IZhleNQMcAaW7D+FS6/Fr0Siq9z1Gbch7m8/t/
/yEgQxcmOWgqxabvaSNrH2OxDduQlmNA1ADEjsJQh2NOBCwRxT9W95dn674l7alZJb8gjf6ArokT
pXOIG38StfDn/NGbMA9dlJiDqasrD8Q/hLP/4wi3xrBwokA2aE4wowQa1S3zzyQCxZVaM00otFF8
saKHHiJWbVcQ3PsJeSSe0YINOF+woy6KC94irr8Sl1OQW0Uo7zAja06i4kUCbJ0DL5VC1BJXzDaw
ZAz7cxTxc+hzMECUqJf9FHVbHnf2HKbmowMnmGf1tB+1XCJgDFZ+OJlNuE/NYfYGoivZd0oPQ/a1
qsuqkV+kItnZ9D13DbHGTqQz/HQANaEUGRMRPg9ncDC3LYpeq3g5XdTDXj5h4p2w+8Xh8mzcYMPN
3QgeLtmjn9Y4Q13FabSx/BxIz+V0Qiki0TR8INcc4IkaM80aiE7eWf92L3OMs6J5WhRBfOEFF2JO
DdPiHipgczOEdwbIcuY+gVGoz1eycUquIbI65fOlIt8Poj/kX2VB7nx+fjgrzbyfkoen73/J2Zp/
nA6CyJ0H2hllRLErvphvuU96pqF1UpDR6Bz/K/xTbBxVF2bJNdrdIXiEF9u/oRIMaRZeqpmRGIKU
f59HFzJaUabeurRdeGvREOHO/fHa5uzh7w7JkCxaB8FFs7CRWe1DXc0QUmo73F0VQymQo+TV9D7t
bASo5BCqNO5j9YrnWZbCQy2LntEzLlfXVkzCQHyW61P0dCSAUEeNW4OeGW3pNf0AC7lrYUtq3UFI
gYAxJD6X3uCmRH0PpNCIJz/16aAo8GIWK96mvgZ2VRBNqZm9wMqoZ3gG2FVFeHzviPM8ni+wkH+E
vkX1M9v11JLfxhxU+kaRoizGHDRgFuWh47TiP6s8naNch60P8hilkKIwc7N+7uKg+FdZQjw43cK+
crUv4DCOPQrdiJ6vBRaZBrLgvXXAhVhrNwCEXzdibK3yG6Wp7T2ptdteOfyyhAPGBnJoZKCqPbxD
2fe0pUvnbBnpps1zLSY+z2hLe9n0oLXoBhyoiyyryXWDMOdm4BlWGZ5xJk4H+h4TZ8lxJtjLVxkw
BVmNNYr6NdnMqPGUffUVu/mO2vJKb+daLbFyKa9TeBQ3QmELhBS/sOKdEVSMeqRC3kB+qwOjx/K6
bz62sqm2lXs6+zk6BmK5R30MxvxaoDOKvYNRiJ5MJ5ZGnJdB5fH0ewheCgtPaUea1QG9KO9kvWwD
9Nhuz3A6RM78tSwFRAKFLUbJEEDnI80u4eXrIsTuClQOVjkEM27mbAEeIc3YqI/0ErGRrWjtC7fr
3rQ+eDy5Tfh4XpMc08oQQ4ZISgIfCHhqfQnMxcwuJLDTGuizNm0HxOEvDuue23M6471WrD2+joCg
+6SpMm1RUxg16wfyC+PQtctGIy1exjp4dUuQ7k/fBTLHGREkjpwrvoFFym+LWmhSoyr5qlXaGewo
KbiwWQy/p2ccK1c16s0dmNCaCdFm90HTQ0YIjMErSnfg86zrLcnTvMSAgJOB0T19Izv7cgvq/e0M
U79yH9teDj11slWi9vLRkJqZtETaI+2Z/cvMjs1vhnV+kISs9LL4nVge5nMeRWmnEi3G2trA4lsm
kLkn+/iBvSZWmmV6aABDlOCsuUUu9YzsduhJrCq2pzQqnk9VOIPpOc0nMPG9uANqehoz2QcOicy7
LCr0rlo4ktBRBgjOiWAX4xZ2LZxQ7KEsZyLbHhVZiH2Ot3AyqP1ImrM5i2bvGH8+z3VQYk5e3rDO
hlvQBo/cAJcJhO18HFgaFyaPvYcsUPvR9Su8k/uguwxF6W5zbBUEAIOUXvMqYjvmnDpg/ksx7jYD
mkbrw+4f4haM1n36atGl6220nO/KkcgL0GNYTVMUPmMv66dEYwVNhUUcMdHEAwMTosnnp5U8WyPu
l2HQPDHmuPOWQ4K8UxlzbG7mMI1caGFwj5KAI2lL3+XmoNiNX2hHFT4H4Hy/vOlN2XmK19fNScz3
yim+SeYjZJCc5d20zBF9v3UkLpmMtEDqpN9ViYp1/O4IagMkGozHTAEOV2VvooSj1+Wi6h/cDIQf
uNBjCv2lPxW1BPllQjznUFjUd6wSS4N/1BuOC1Sgw8nALDsj7/kfESq+5G/Jbs+90cYWSCpRORAV
EVHHfcmYRjYlcQzR9C8qwmirbkHHEZdGMfBoi2xZTU4Hf6tLBV8wTgsnTS+sCIc9iIbnrzDI2oNZ
p/Rca4jXTH5MPokXIg5Y5TrQyCB7eUUfagkDmD678tkv6f/mSBe9rc3MAHZUuh/RHDbMAtxLP3U4
wJWtDaT5WITeYbfAT+7B7s3KR9/lFHS+kzUC/qPx9fI37tJR+oPHNwfMXmh9JU6S7BTHZHepCmDf
UEgVkpPp0UmHWQV6BZGLHCmiIq2S2hE6UOkLvktNbwS6MIHayNwo8J/87hn7Q4a0JJlFpotdo+uO
gQ1nOFsQKoIeYD1PszB8uQQMEKr9HJy070RCx7jI6O3ANsn0CpeH8g/lG5nLRltmAV5eNd4ML/B0
g90ThrMrwj9PMgmS4SIPQSAJA+gGg4MS8n+1kgsL415IAGUyXs2iJzlcziOYbkBkZoG4jx8ACkzj
OaqMnsJpbAQBXN9C5G+9j/hU2O6ngAmFvXmdJiJ1R5u5Bub9IsuQlJXFjsFr/j96V8o/gHYAjvPo
d218ecjgfdK9m+DCo6wTLDvT6w1tVR3SfX8HVYP3sFd5bV5YzXSLNGF/Bzf8mBEs0vALUg7ee+ce
Pg7J+5tl/ESPGPgRxcNFlEQL0RjwVoohDK/9EydOzfctF2lH47D1Cjp7+IJ8BQBQmVKR6d9hq4AX
XF8Qf6Qs0/BLUsXUQ4u0y8d9Ar6S5h6TBckUbSE1ddbhAlzPa0/WNwkt29if0A3T+6e3uo7Y2Ku5
OUaLeqgOVD8tTWHGb6qtMLgXsWrb8FsbofD2WHaHgPhQeUTawhBENHtxX2goMjWrRr2tDY9zICnf
4mkUYNy5ZD+PV5Q0MZUcH6HHNi5wHgP82C49U6+d4UXci1JulcO9NNEAA+ftnK/+iyxUAnlrLxS4
g3/nKMLYNhw/UhTzle52G9HmQMuoxLgjxUkk0k1nzssbrpq7vq+53T73cJicBw9ssVnh5jsLXCJi
xhNzRCR6sdH9jgzVy8USlcd8vfZNgmQD+EZ6aykEpcuj9TvyNOm0qgbIDLngjlSsYfFfjMCzd/mc
ZUcz7z2NjX/wz9Md1DFSus0WID4gowi8KdAfhLjxksRhh/WE0PdR7SwUsMcx9XcVWqxGCJHdRiXe
NxSis+0VKvCRQFS/7KRCr89v6gaae57Gmue97AFpd+UYNhN+nzANhe8jY5ULQtCiGDLzmLlvbTH8
V6hxKq/FpQ07TxHtU1ipowFYffPkP/iFV/KNhsslFgtRyg4AV/5j6pFCRUY4niBgMVlBKUK8rLa1
5/X391uj6N/GWWkeYMhS2URaGAB2cXCtqSI9BnLeWtTE7O2D3JwhmYzywrJ/r94JwfrpH0D6OZEK
vMM23JnXAzRs9WuH/bZWmBug3XX+zyhJvC759abC/Z0u3PeSpEt/BRniWNVOc4unbp1E4CurD5fT
BZk1abQ3t6pP4tQDK+4uH+oNeSUDGLZUcN3M/EuLFJ0SsQJnU4nwRnFxsVNm441q+JOWLka6FczC
4Pdb3dM+vSSvbVeTNfIAq7gxUd9b6nIxWeBdQWg5gM/OGb3BBkZlysZbwdswTggv05FOs/XksJrl
41N8TA6mb2aDllwmWw4GY8ZoKGCADDwIf2qGLi9IfbyD+eeb9JI8tQJJd4zxPTh32c1d/RQlwZE6
IhuQ12FKOlpF2rsQH4xnIYlQ+yUF+xZ5cjHku/mHC91Nv4mrS/1XNSmiryQADfJPUn2kwWX0ZbDQ
HN0q9pCqADdh6E/KLpHkkeUaGe80Hi9lkLBBvGFT0TeFn/1bFH5cjLSctULq70gc4NAXp5FpbGGD
gBinUvJnl6LZ9WpksdzpNa1QbEV73XNuNGmny9XTSH1D2jm54YSJ2kYEIxOROJOTQln3v/iYPHaW
JPCJRzV4DvVlwb9ZZXT/JvZxLJcxYH76I7Qaav/HPxX/eo8lsDkmBtHDHPu8QBnKv7L/qVhCn9tN
KxyV7ZjN9w05kVbC9wsNH4ICEl5mA+0zopAKtG+kgbB0hujMl+f8+zb+Om5SsGvF00blVJENwOpA
s2Dnh8dsyqB5+ZDrO1toxcmuiabMyrXHN43CZ43ejHaHXW17ferLbo9TBItq8Ub7cDswto/YOn75
+CCU/3RB82mvki3xA0FGLeJM6pgaxhosccDpzNxVZqw0Ag6KjD2QKju2rxsI45x1s1amJSdybFkz
8rYatZhnX4QcP0p+gblrVv+aQYQjJwpcnIhubEClc/d85dq+EhVI7pJPNgeSEXrMzmvxuzbOHLOK
2FhT2FcYtEdafj6h5X87bM6qZC7UQJk0WIZEUKxAujewK/Bgomx3obIk95pzdtKacLQ8VF4kNJjl
lVyNjTpuN/1FpDuABD0Syv7zLeuMe75TojuashHDNWpCfy3ZcyrMsVSj9mQgRzk7Zu+aonmZYR2I
GAjx4tdrAFYJss5NYOjFy9/fUDAQ4xWe0q8liaUA+dp686BUWIxw9Yq3aUpTW1bqtNbkhaLAUQsI
sRZ0JxNrV1TlDrQhW4O52uzjx7P7jT1EOZEe/M5cNpXbtY1jWrf3PpIwwGl2ySwy5FrvJ1ysPTdU
3U3/w6aNXV+Ss7iApD7i/BY/j3Emmf5VTiWfH2QnhsIiw4C/6TpyLgnwrIKnyJ46LYyQOo8SiHkI
Kw1PfesQGYihRLo5gjEDrHxfX9vFDT3N1YHm8CcoyioZoZ7gauPW8wxgQTVuouOD/+6gIB+DW3uH
lE5h33oB44CzKrcq/NAKxKk8F94YLDYbgvAXUTQj6vcX6SSkAzxpqklZUf+0Bek8e+NmY5GRoVIF
hFjS/0Rqx7OXbueOLjrTqgFCf/NWxQQ0w0ghDBx+QqGCxKGgVTWzuu7UYHq2YK3YmpdA3wFlqNcX
0tHDtKIsssQUzdXtTjHUBb+st/sCI+T8CoFRNTD5TlXrXlR3ehOmSJr0PiPby88GC/6+S5G8WpG4
xmllTwolNp8OTATGBYj9FSUc5p/saykTAI0zZpbDxW8hptSozysaaFLl0YcHOlWXnFWl6YGaGjiT
i8jJ7kAEUUljhhBX5oBI6Gb4Eed7qPmyE/DO5awzswUI0f9Fc1wdjhF6O/4MIqn3ce0kD4Oyp2El
ncyj7JcUBip6zMbRKL3uMhXXKprN8Zhelu1czj/epuOfQ34+nwt2eenMnkb2/4zAZP4os/KjcSdb
sg2bVZf1tpd3pLhmGj+rrVXD8V/Dh7yooJyyrYRiYb6Vp6h1wOFGSFSc039CyUGB63qIi0DIvvZ9
aX763Z+s8qgqU6PzsYPuPKDGKXXOnScEd81fkDyp85uuZT3gG6mgDipQSnQDCakEApdV+AbsWQfl
6fvQ5kPfXivLFf+D07aTkCmGZ3rf42RHWhmQ2HkDy2kTku3t/fumRrfiAKnjxfXKy15tzgcvD5NN
0QduqjvJCA86FALA52/nO3AwhoboJ4sQFgcl9zkSawb934+X0ZedlO/ntLUfoQgXS7ec+4ZK0Vlf
PMV5CNxsTF7Dqm19Tm91Z+R0AGDIrIP69Qzzo+eFofEBwallRZ5kkCZs2sijFx7cJkrSy7Pxvv10
oCAjxUxgoE4vjF624CZCUoUjipErx9Ee/BGlxvFwZys7JHF65JsoLRGF6BexQ/NQiiHp6c6bIazm
zFy3fTI6drFgW3YYAGntN+DKLZ6QQy0UBBykLbb/eryImHTHpkwt8NCd6Kutfkb7EJpEhaskrCuS
/iiPgJBTnfK2KE8btBjUFFlYUSh7+k6xh1i7kH+pR7tKU54W3SoCfpgXGsCiH20tSu3h3BknbeZG
Mq5oKlibd4djuv5bsKeRe1gtwJcfXPvNQgv77+ECDEf3WM2eCu5luUDK4tE32va44LwvjqMYLrMl
e+9v//PHlwyrHMeEUQIKgNcw0G8Bag4Wjlu8X14WviLeKcR4kbkA1X+aTMTo4YzMB1N/ue3YAvj2
YAO+6/HA2rnJZfa8at/RwvVsxFp24vGT0kqEXse8HgqRcrVXQoKEGuJJr9Oz5+um8ekYAsmE5N3x
69UYxny4Ul5WNOPQjhV8wgtTd88+s+IyHG8ldEa6Uj+NCCpjK0So5d4uNNiN1tk/8tenX2t633CA
gXKuwPQeSQjkcrsSrAFkPQ3drQMqQ1XDvDeMsnnlrACjNZKZMg12fqmi3nfZtaKambT7LGS1dOK5
tv6MCT4sKSUyVj/c1IIaApqrHxwl+GeDJ/1+9EF+JgU2hguUuHnuN7nDXI4xA5P5fdd4/AMZ3dud
xcq/2WWecz+lVLhuYu6mAJ8XbKijczvUaFvJoKvs7mDxiVtswz94RKpDoruwNkAmZVkOmGjCtWY0
jrPvB068vt5MYj8I5aYeMvMo4LuPOvwNix0NH+meIGj3DqTDL4ueODcRGCwia9i6XRTICD8ufQDO
V6y0plS2ZengGHAmn9txgsLJWUlhhKaBqkIY6NvqYhjGhzak7uAkv4u8x0MrX0iIgcrNlm8R/U2o
VMPqhW149iDsjuEhwcrkMQbcGV6mpMSX2AmIxk+67LTvCwjVK0T1QQqiuEAb/Aa1LOTGSE10ejPV
IClJLOBJ9tN3REWlzTmYWXw97JTa1I4NJrf0v9AYA2deyuAE5wKIsbST6SZt1XviLpShCiIR/N8d
GIoFM0iA6urx69qaaCXjICIrlP759nMGQFK05FzOJ1ERGtMid2aNROml2RMFJkpG7qYfNhrdWHuo
D9HydCryZGQOJIhSsXs90z1E1pHeB+J5fboE7reqathXl1tWpfJgEck+V17BlqSg5IpquoiWvFmg
jpkQJhL2Jlx6iJe5mvJcWkTLCVMLUr/b0cPD0joK/cWg2BuRyAz7AWtO/WKOKpAfxaZrePBLLDl+
uIcZXIAglKPMq7oB0WXLlSyb0RwUEpbI5GQGV8XsM7GpUil/IBx5BKd8N3x8FJYqd0nUEvMBEHaS
UaHjpX4QA+OapdwafKrCz0ePTgvVhMmM4ABfTOYLYkV/Ck3BOTKroXYN6x9YUtaRTlHMLW152XyW
sK0AM8g0wFJKyftohrzwDQfOu3q8G06NnN8zN5zGnvzZAVfb2aWZbRH8bREel610UVW7xYbxT9/t
CzmVaV4GvU7Zc98BQ+AFOpbr7x9Mv7bku7GgGoyxWW4id0VMlATpIfl/18JmlepBYEbJ/bZrU7Yc
cywRGIN7yUib7JkYFvJEIjcW7FgBKQk02mTR+6KHXFYGFbyXz3rCpbESqPrZW9AH1F8qPi8ySxgw
EUYPXS8wwF/dob0FZlghkdZkfPDJcKZG+Jrm9deOY8fRQ/5GISdrhhg+SHSgU1+wIUwpTAp5VeEf
wj23VH9Hs27qRKi/bVMyWPLxDW0jLnvO7svZ166SPouyXsDhAefwXR+t60NVZIuLvXAkJA1UxNZX
jrxL2fXAs3WJOaAZiGWpNyckqrnC1PQdJkrGDJLI/cKdALJ6H4eQMuzsxfSkC81W6/EE171WcQLN
riv0+VLlvk+AJpC6RXobm8d7f9CHUsdZYYHRrEYMaL64jZvL36naqb5lUyuR5zQHf3neHOVJT0Wt
ZL9hmLpFv0iv2XOKmvVt9wF9nFBZ1tIYFVnzBTixbN/Z1P2jUaSvuosuXbVwjgV0wWIoFNzKwVb+
njvPxZ6DJglBsr7sItD6woD2iVRTcaPnoSEGuoP2LwIauYhr9+TDnEJzdw3/S4hELQwV/WhBl9I2
Nrtyxw6SCGhXv0BbXAeiZRUS/jbe/RJqKfniriM+/tDAXSvAX3xkSd0Lg6C/yZ0esmzgrnzWmYM/
SGVTI/Pm4tSlg4LX7sbsze6VrWY9a7hFQAmpU+JlR0EdWBgHxzCla7MB9qDsekUmtnC/naIXewWG
8aJXJA5XPtgc3nN8rv5ZHJGPcoh3TzgxnYcZTyCBbwDXESg+hhGEQ993TfOj6rFMQQnSBaY9hH6Y
uf9B7IUEyegwRvi0kqmuAIuAhZpR8HP1RGTBmFn5McIma/2wRREGIxb+SRKlShHYXrcmMeXRb0Xo
ZoPjaJ43np4rM6GMg4RxSLxSIfE0u7j1W5ioYnxfG9JNN+wCdnkU4cbiHHyIx+wmQwc5bKdC4gkm
KHE7wd3VLgBzzpejhbAqjv+SHxdQMOuM2Weuz6ZFx/jghsU9XRdEKiqkpauXU8ZClf/4VC9FmttE
/bFa2aoHQVaBq0czlDaMG1B3huz1TTjs3I6H9XAQD08A9YnprLl+MSWovAkqpR1p/YNSl+xU/4GS
MC6+tv7dtRFko2RNENnbytdjpo2w3JKtf9T7XTXpauWBivyfdCjwhv01zFd6NSj46Sj32loVzzum
kTrBsIuod26NqjkLbC45c4ub6NTuK358exieAipg0niqWUmXWpyzwIuUb1I5GleH3GsPWCJ3E/uW
+X593eTlxf7tGnoBzYgXJqgrKNNsrHD/ePKBxOFhkN7oFsLFo7htWFLgj6el7zzJBaaxJeiYswae
qdaI2HFOouhYUz3bYJ7p09e1t1ouRTwDVvsy4J/Vr70wUtRtPFMrGft0D+QfxvZkXF/tdEe8QuPa
Ej6nP6JT5n8J9ohC6kEj7MZLaWx3cH1i8xnOg8++LRMFM7w/VRqY5kS+oRAky3tbp48iPfCnYrpH
nHRWas6Xpy8G9JClleZPCkijUGNWJlirrkrcSS4rWfs3FzhvHto5FieGhzsmS/n6O2mb8JeHo8kk
YVic/Ptc+nLHj+N+Z3j6y7X9TbTqc8Tj6xUmMycPIz1RPYX/igaIHxeuj1FNl3TnbTbb8XeR3mBw
UQ/v8B1w52p/vaDrtV+F0hslVqnB1kTI08s1kb8rndZxLDySnZqg7TAV46ZG1vZhgVnY5HmLP3TT
82rhQ862pfYcGdYj2mHnAedFq8oPyUsyo00USO53WG+1xcBDFVbwT36rWXWZ8OoLKGpNdj+/p2YC
yHlH+5eABPlrgkgUI170gcqbvEyKDrGc09pUaLX5btQcYDXLbDJ1gqaq/zKqSkBAx3mjnpULYvTh
NZypGCZYWtdP9CBBVoJD1YwvfqIeU17VT6zMHQVEBQ9G5P/0mvKYKmok+kkjxMcNVicLnky03oOM
X4wvT+PeT6zxADA5BSoirsQZwqQp/stdn0E0s+69OT2f6X8wCA9UGCPTtjY6VLtm+lpSodAh8pA4
/UakYVHcEtEmyclibiHqNXSce0FzvxNfj84+LHSMi9gm6rx+ZxE+3x/AkX1MExZEgfDPjebZL2DU
wQgI8MQSjE7gwUs8/+QCjQWRBhN7kvbJJOUU3qrsPHlRLmUci4/zTWt/gr1K/D/1L43oiMqFRSG7
RuULAmLzDV+oKpfQKde5e0jKgM26YJWt6RJ4IIClN0VNiLOwLoYs+5N7HVCvZg2KysirYczWCpGG
PAh3q3CUa8rgBbYX5uyKDqvlOAw08oAw6xH+ZEM51QMRz/21SEqAuAxGnB9QNCg5edjhAX2JBAcv
1oLl1P2jDBjojXeY9PECDxOZsXQIDJoG15Ok2oxZrFFdVI2ByoRa3sL4zl5ilSJERgag/VgITBEl
1TWjG8Gq3VDkS3fwW58HgyO13GoeZs4Vt4W5H2nJPPkZ6Rgm91yiyMABrWEhDTZMrzGI7AnsdONh
VP+3EClkYwE/t/+qWGOeN3GwrDRcBz2hOggfAUpHoCiEhWYcmnlDl18MsCM5LyT9o2SnmMZZCdJ1
FLEZBu7eSmNyKZUPY076f0AhbDhBiQXbrH0CtsbWAD4xMH2Zgttcv/XQ3S7NgEYbFz6nBeZRxfnt
XQ36ELQUdzZNQ8Mw554pt0cHh2VjWcI2dlOOX86YoVpzQFdaZFitxx3JJId1KQHqmN2BJzqq7lAe
HO3mWbpL4+K0rgMLqXGD4iuIw5SomonrncGh4v38rmA2VXM7nxbTrn+3fRFQKf/b7F6CQbhaLfQS
dYwoiAgdBeUq5NT/vh0PKtdArugh2BJKrNWgjBShSxLhjrrW+ODyPgEoM8vZR34yq4Qv7GJxIE2n
MKuG9Wl5LH7NXGxYatjY8Yy64qKj2jAEDqE4bksZtOK7qc97ZeLlnCOKx/JZRyGrkiWRLRTLUin+
PIBX7kADFZKJ1/pn82aeQaAnWQwspu2mScI3Bl3A7Ix/il357pC5m8y7OLzhCJl8FmDjIyMgGiAl
kRBjddCHGB+37P0PFJ+/0fI8D3H0r32VOwk1XHHu4oZpyXXwR7U5p62FKcvolypwW4z86oqyKm3K
8O8MrBfX50s3ApcPHbIJ7juWWIlPR7F1yHJ7wvrbdTTJPePWbtDcwZL7p7G8fXatC5u2vtcay3uY
Ucwdj2VDEProhNMAhZ1Nw//PuTJgyVBg/HwPiOSqAtVGn24ViS/f1btHUAreA/eyAXT2Nq4yQnNI
jF7jV0N8te11pzFpXOM4QkbNzJFyGezjpMX6lXSEE46WTw439POjsL3Vvf+DBJAurVf5hfg1f61f
lzFNDGVAQnOIeC8wdFc2yQGaK5gDBiGY4bCfPmwWUqIf0x1stCH4YMJb4g0Ys+EAUgmbwuDycR8V
/T4+kg7PHgi+cNhGSRrAaQpy2K8qRt5i/arh1nbeM17lYyBMwkf7j3/cIuQvly5IK5lGIyf/uk/d
4YHofIiKm0locR2sgoH3k+6UYO/Y2D6UgZooxwksuekp/ksOc5VZg8cvKklz9F42hbuGigw7XEe+
BCQ8wihz8Q1lskw5NDVISuC/y6Lg5sGJvV0yN1Mi8RJkcss4Gypk7VSW2m9z9mkSne9Kv08yNO4y
5Q65+mHKtnk6auQASVTuuz5Lwm7pfSjl9zP4tStlOz87w2IArUEoMeSAfMviGdWD25p5GHtXwMYG
i+BYsZZSgZL+uE/lHB/FdiyGLoYoOewBxiBQFXlPRA/u1suLk6UwHkE9chwX4MVSs9sYJptoU294
7c0iem0pDOcz8aC7YTWK0UNrr4Ye4bDnNlT8fLcWeGXaa3G0jYk8CtkgCrFX+BwaDlIG1kqIHjS1
paGmG0QvhRFu2yJ0OTvmRUHunrToaquS9dgsymLSvXshg5bsNnk7CSvKgjuNM2RkrrpU09tmiIy1
lIbTLvhY4MMlnXSlOTJG6Z55g78N2PG+1QubW3AQqMt8Ts2is2Pdj7Ij3JPaG4QoeHqF7eCA8N60
DP2q/cNrw9TnBkS0nQklVW8F4/C+fOAYTeA+sDwMnc/BwFrDlIGqF6NlF2m3UTcVMd83z9YEpoB0
9UtqmwmrpYfM382IeJgnM+VLstUNrlTNMSAOngd6tezUG3wsGs+NJ2tACEAE1qYvnDmX+jovT66Q
rDgms+FE8H3oSigXmK23Jyp95XVGVmuCgbmJENYIr2bmdaeQPDNQ/Bv1kxly1A6a3bNhBNZJt5RH
UU/602R4DE1xDzfNAXPKVz7v1YWPDCSHRhTuBOvzYzYhykZbk3z4VQcONIHzLKtY3rUM2bU90crG
Rn/nKLATGkob9LqTJfAnbRXq0S+/OQWKumew+AmIfAf9BIgMTBPxqvcG3nU7WQCc56v6KZw4RmUF
z+JtWO6x9Hj/roOP4qCZcUKapwK7ANHL9sT+kzjUEIC/2geLDsRcTUydFMZo/lbp7VW/bhE1QU7u
Hw1U4XbyE5Vy6d8ybXD/Ip1vxn88ENiZcQti0P219skNHNHcMOOqKFcMFQWk/yxWm487gN1vFsT7
LzlipsA4TsDaBC0iqEEjx6lcgNdLzJ36fsjYz7En2ZOWeQdilvzDXZFbgCLNBx7ZWSaDf2OJqsIb
kZ+frFSOKFl4XE7eMoOHAfEngbPeU6mfcE4d1tDfsdwoWvxkKUbB0CxFwmzQd39F26+bAVdZmKgh
KF/JWwveBIJkigBFylRhQlo5AZVpNQPndBx5L+mqjAMPBZaSVJvIl+zXupar0Dv5oHneYOzTgdoV
l3rDE6fTYo4AaUL/pt68OHefsNQ3CFvGEjNxQjt6A+r9bDtqnVFShYWCrOrQ4tQaNerediuT9wwk
hC/WXFahGAevAt0WokCEg0+wNBNSPbFtHutRGfgSM7jWQyxGElCNI95xfJXQelslvZnE4AWpEOkg
dpBKTLAl6uxpvNhPfvmAHKnJ8/GYc3yKk1PO5uYNfcfa+edMlAlDubXCMdEoWIfZI6n04jG2dfEi
eqqsTK/NMn8Os0vS7I7FslIcZ4AtJitDEONYPjKhWpRj7r6GYw1vY5kEqOQc0txAFgZOGkmu7sId
QZGt6xGDYi2X8rQR91jHCu7ZhUAhiNP6DPQM66dl9hL7bImrzVh7GcU+lVL6AXP6Ynkm7HVpFHfY
76Mmv3Gm/tj1+sOWtJXeGBbCYwpbLmfz3IBkf2cd1N8maquj8jf6UWxeKg3t9rN4ma93xanrM73o
Jpfq8EyRR9E5h871yQMc7YS3ps5hc/NBAKZ6WBw2qA2gCAlBOTYwNTSBZ7KvlW2DRHsqas+qkH2W
b8DLBlmUDqxKHHNOeE1ibsYNBOM1rfyfJzshRjrTKNjoujTiS1G72swUcaPwVXCj0zp135A7z8+i
eu1HQuH0LkLOR/zX8zX7q0llxQwsQesli9OquVLTYzSOua/MiLe7oC0ltPGcpsV6GnFz8COtHQrV
hVU3Qwa3X3WYmmNqRhA/uAw+oDpuJtZV8UW2RqJgD+b+a2S/frPLZJF8AqQcpU62HidNEY+HnVHi
n+iJXPVJpvx7dgCohtb2gdJ6OqdQEP/33l/ntQLBmbEwU2N+hKQY26Ac8d5wqWajAC8ufLH99J2R
Y3VK2NMiV/OwZNome3AbTXyL4Q7hluzSpiPJiaitUoRnfZnglcEzDhs9cFbnJLv6k7p1dYZG6Zp3
yorMcVP5LEoFZcbh1gwPky55GOjmkGYLOWQKuHwR4Pa6Pm3HWos5/Pob++C9VZIhl/czCvXug3TT
VuZQlv/+9GGjEoh72FXlsE8nWutnyIpmvKmPbkccxTSWwUV5PGhilYcR4mfmlv3C9MvJz4+y9A/A
u8MxgtEGjHH44eCBUH561PCZ3b/lL/HLxRFcaZTQZ5Ff+lDJzKjo+dYSVWb/T8f31NXOy0Ert0yO
Ef7mGfejkNzpSrXlE2UQYkaFNPeBlcnBFgP8S1/7G8IBfd7/GlqNDOm9YpLIUoKzefFROA3bDjIY
1V9Pe7keYRfkzJxD0buyrmopVwylKu53WbwR2ZS5k+g0Mt4GuhZ4xuAgBsbywrfD8WB0+OqqYGCP
z8L2Rm0voouaHn5sh7WKAZF0Hwo0joAnHuMXWo9Bp2qr51rEJsqPTXIYH8h1TR7sIxaX7b9Fqt/b
9VSLuVbMNC5e/QSFcMH2P9vTYWPIk6jeLm02I6t3y3uksDa8yjCClqgGs2L31e7tauikYXAtrlh1
t6Af/r1/cqagIdWm/x5Btw+x3LY6RPdqj5ggSqUu9V2MzAFjc3JOv5AEYkIxd/fP/yqSUFZa7QnN
PVm9qxyywe8UC6XT0kIHyzUe0cFAp8lvIndadKPrJhjhXY8zAQOQBVN+KqbsmaRZhHP5Pw/IKPkP
KCjHpWpnr1dx3HJjICBl5VscZfPOH7KZyycdlP5WrV/B+7tMVrBUwmQ13NNyUtysIN+6GIqGYIZU
KoIYBRS+LhTvHrA6vohB9OfzzP40mU3eEjHEdWETIW+PMZ03O9PFAMiBSo0KmuzStZHG2U6WKLd8
2gIIhJTYoNKNDCPo1Ubvm6D/btRVN+oflgJyEG2xDqkuyACzzT5op0dribQ1YRlyh9ru73H3Nk5U
dwn5HvtfkraiNo/lxGhoWVRVLMZM5U8ISnfscjquZ3pTKjUzAravu1cySsq7mw7mlj6gWt/35y0g
dG8LMi+2ctGrV9yLUVp0nyjGLGHhPcNfuHurJ293eGZDMnvD4v6aF+Tr6e9VGWsOOPWNT9p5HPnR
RHc8X9KEAdIDP0xLECkGrCzAgQdest46dFT/78WspYmK7SrLPf5rwhzdm5uzZhhHhnSOuFapeOqf
MbXTDuM08O4h1ctvH1dwHCYvhW2cksJy5SR8jJSBY43xAwr5vEnAybYeX39rhmTkzOcfaZHu+ONt
nGuh/kp4W8fxFdCs2gCDmLJH4OmKzDXKoWVNmzbZR2FukZ618sFJxAu80VvxZZt19dy9+edvylbv
pdYdZlQYzaXrQGJSAUvSogHCU68LZqUnQq1OICleMov+U5nt6JxWIrkFGZpHOOYBifU32MOBX7z8
tri2d73t9e8vN+Zn5DmJFqKAZ99QQKMRGXsoMb41WC30cgaDQvsY59NCv4dM3fzK7HLGb4Y3LN5S
ytineI5UEgRxHoxrmD/UhquEInaQ5u0DXoilqiUAJBzvnlINL1UJwy5XH2q4JWgkdmLRH6vVUUZM
JvwNzMA3IA9Vtf4y+1p/vv38q+PrLjGOei9s9yQukuL6rpNbu5MnHfpsEK7QGd3jkvzPthxulC0M
qENikkeWSjgZI4TWDHbEnvv3OMg+0Tl2ZJ5fr8/5HPwO+7LOn7O4rAAXTqhbo685F3HCCZbBzH06
nnoYg7ZqnA4zhc243j4EBy0HLBZ15LfHtqTPO52LA71nZvttdZU0foRBihVHT9ypqrknziAWTOYF
6sqjIQwtuAPPq1TR8Xjlucb3/JzXYvUU6GPCjkrOxZyc/7l57vVBmEKMLF7kLkLqr9N4MPQ9yuti
JGltqu7Jq+cb6TA82OcNM66IQ793Kfh+OdhOV0HzHStHCXW7TJPilWmqs7LjGdT+jg+Q92/HMMPI
m2d0uyaFTjIjzLDEOhBL0IxO6tThz2prsT3FZxSu4W8EnhTfbZVSIO1QFeWaudUqz/635S4DGovc
50a6BFQ69WHk97GiUDt+ZY1NqDV2Dc2afWoNx7P/WuXHhdP/9JWN3+jbuwThecotTno26igjzP6a
PdkQe6notU5f+pO52oNHH4f9ZBo9f8ZOpl4L7/PyMIMCWkCTgAVcm9pbWYahe+bLYhKRX5k8rSxn
6whlqrTXfFGEp9nptxa61hpUDD11ptKF4fARXFNfnhjpc5g1GT/T70fP0/vHcf37Cx6YlWY8cuhE
D2aUSbq5oExaeunBnOVz2aDfeG57SPGPjlcETBjNdUrRU7hdB3yKwMr9t5ECso3ldkT26xi6nqrm
PzWgfeGYIZ8QdRJ88w5jZrmi18BlhKCVSs5LnvL3VA8zE4B8YUA50jJY+3dFp5RtA19GUCcbdqZt
Gy6SqiYohMzVRJelqKPekm+sEYhcawwyTXonqKRXd1Z3bYS2rleBkkyu9mTBfBabRu0L+yWMNpoo
o/+WetPI43lBOYJo6zFZxkmv6F/PD5D5pUPsczzKfSf6wYjkG24DoVVIQa9dqbBcJj7NVg7vlOuh
FQAGu/3H1Qp8lkvft3G03zbCvVAONpElTeJrhGqYiltptIM38Uf9su+NKbfodJk5sNKog2RyDs5A
sRyLiQfNQ1wPxD1jw73TpL7OjrmE/G3NCF8x+bf1tr33K8khnkaiE2NkJdwuco/SyCRn6qQVEgqo
6eW1cytaz3Dv253QPtw4atvBam6lWh2Lhtef1xSRr/xR77rXINBsdUVbTfCg24/TD5UTE5pjYZh1
GYUey7ZMgFT68JCwwvGeWID0L14C+T460mFsqFd/m2B3XxQAj157JDic26fgTUqkM4NL9WuOu6DA
ZNW4Az8FNcanq4TiM80rwli+2wRAhbSrdFUM5rRfQZqOE9FREHtzVpAVwMcVk2y1bNBU8WKn1Uzs
u2QM7BQuojWrM0fMI9N2Ml89bMqTkQ6o3dzWLnVbIMO55STKhN6NtF9N078wmjzjFLch+fJ5N7Jx
Ka6thA4xwjbcG+IPfVzWTwVAID8sfW2bHwm3k8Vcor2HC5Ti8XfbJ01FBz0e+dmAbgT2EJAj4JzA
TmYIr6YpsbB1Cws5zjrHBSJTS0etXPWyP84eck89HJslxlsFXizMa+sDpPjQnkmaoydjFzDW9R+m
mQdfQh2b+PKHPQAb1+EtrNEB0g6WrV4+TlyGsiy1QMys8xJsyoPeYcU2x+9s2zLkma73RwIHQIcs
q2m4tWJNESXJhBMt0N3PY92ixJxBd6fiXNMbl2Kf8+eD1Fd3mkCh9sC8mvEKKgp2dxc/r5NaKnH7
zsZrxoMtJ3wewWe8l+dCSqcnqoXGkRvnesz+61GCMVyNsYRAqlf9n8ME0pUSrppZNaJsR/9XPx1q
zpk41/41xaWW5UQGYXFlhIcIZ+DAIinDMMxc5H2SVuUoSy2lstuQSGEzdyVFqmTP1aG9DhN2wbej
i3ev0i7f3er9G+QjyOa0CVJcuqHfggJc6CTkfRIJ/pqCSc22+4JLDwDmvU4hX8V8my1Ri7IrqUNj
QyM3fd7iie9tm6+E6ycQwAXBHXnvtfYOm/WlvY3M5cDFkUCv7zyJbKkMn1TOCY5gbzgBTOlEnIQf
0W7BbZXbzAaaKARPdrwWYiIdOGVWXdg4+yu4tRWB0Y1SkeUNsRvgN/t6N7kWYTHEfc6hsjfCW6FD
wwlzqT82C0ReM7ZWRi5ss1SVViOSenR9W1/3Oo6E1vOwDV6ObewZkY0SRTfPwYLUmRV+Bnw88fdB
yGp8BWBpI6wxNQz5f+nG5r6AHrHfeqeqEi22aSrpcRs3H0LHhF1Jv1u1J3W1kRj1W8UYSM1VbAlV
fqlb194jUzHwqieXJzPlaFQOyu/tV+RM2Ruvd9xclJSigUEfLkf3Y5QeqvVVBSEcBDJqe7p00li0
GbgD0QKFfIKt/7cWwUWZNGTUwa2W80d6zm0C6yP2yDDSrxGjj/Hc86E9H9io1rOkanIZcXA+/Nfm
HbGhXbdpfhXmMezUax0jWGcrQw40eXD+AWG0MhFFuOX4MiuK35yiHVYTT+WSDjbdpObdWILvcwAB
W9w8doQ863UnZzrejMem1Be4mGXHtrVGhuC9vb6tfTy1iaU5+KZvIVKjcLoXjbOFiOXmO0SECVwi
zxUZCDoPJ0+mVP/Za+bPJN+f1heImRpEPo6DfLLzZQuhhhGbdYuxzJD4S9Di5o0YBm5I3F3c+3Rc
vQ1Flo1Hn9d6nDgL74/b1qQTT/H/zdLU0Xdc7dFsoJJUp6Q2bO8VdrxWy0ikADWsORuM/D0DfSa/
dmR6GzjTf/H8FLEs/EfphkIqflEiR802V3zl3vMdT+uysjuIAdE9yKU/kLOBkGjV0PMS/jV/cir8
C0DCMJtxWcVKbR0WQ4qGQRNG+8WqLpjH2gfOgVNUJh9SzxCcAfia2qcasOKcy+/+bJK8kK67BHYd
7NSuADAhTAena55Dj3Ru4NQTtP03F/rv607OF56+5uaLB+NbWvp9sAU/n3dcEijn6bBDn+xe1btw
4eIJVII7E2Oul8i21cD8GqD4gTVXe4Eq2K7zvSaRAaU72p8tWT8s1d65leNHxX/GJTMSi4GDoP4E
tYVb5oOn0KHp8hlt8zKNpI33MHAq0P5p4Q6fSVV4LI87qeRZT4OtJfZtYeUqaU29E1gS7zoy1hTF
2MsHVI+Wn7yoMwgh8ys6aVkcN5JxTXnbUzbtqq5rTfiHI1PMr620Sge+E557PFA7Lu7GYmIgs1Dg
9iigVz6LK54jjFq3Unbw176cMgRRH1EdlAvKWs6fUMEghmRzVwAN0V+vvOnxpL/g7666GM22MVOr
utjO1F/fyT2nlOUU4cbPuMLh6STO47MhIb+cOIymZJHTRMQUOsOqkXf5nsiFp0B5U122zqYjYqgQ
DVMw4jsg+oT6H87IzzCQHNNB9KAoV+cm78JujcFwqYGHsSWRlC9H0+VR8NIKCjz2Rl+/63YXUE+z
bnoEK7QYPVmwPXZiIt39nMtN1ID2uC31kHmJOqibHG9A6rjYGEdj8kKfb9QZZzfRwV1rP1yBiqt/
dTbaMLD3ihDVC5NlEwM8CcTZtAqbupJyLL6x6cSqj16tYtqCi/hq/rRojqeTF2kXKke67N88dLIv
/khEUf1+gCwC28qfwIsP97lTsG7ZP6YHX0fG9Yjf6k995L3ecawd8sn+6pXkP9m2yqpisL+538lH
+GMzItKfxDwQqCuO0EHZ9XNzur+rH13ynsYC3r59XZTA1lkXL1ZECyvccWHTk5FbL0R9j55fxCyJ
pIacZJ3Lw1v9DRnMMW8hHyZMr4wVdJJI10fnYrB2dCqueZUIcfyzWaQXw3FMzE8ELLGz/hWr8X+u
uPglEJS+61kh7FuKotiX+NlrcfOFCKJlpqmcIs6D+Nd7bOEJZqHGC7X06qZefFHmwNlZ3vp5c9p4
jxjZEOLIBk8zEE2TLiB+J/16N/8TO8D53jZW7VaXV8P4DwlvtOVSCDzwVt9iiqQvnXah7rJQC9o+
nAsvwJhkLxDiKeEgjG+CYVJbdIC2csbRDyeaxHjVA1gJxWeK4qXMxgwFHD1CRTDwQ3mTjE1TRflA
5ptn5JokGhOVJSMeTRe5aKoo2v55y7aTvI7PwqUJ388a4e1i7IfRU7N1RN0mCTd3W1q2INsvFqVP
+0Wcm4qTmCLDajEU0G0imHaMYVijnBQ6aklkMN7+gACyZZ3uE/6cf103AOXSmTqsq5b7zhPZT+2K
UE7KhWv0mACVn8S+qitUE5uvnLXHGURFt+oOtBkoEnkRJGu1/h77jW0gT/L6+WVnmK9SCudei9Cx
j1XsvOEK0i/5fCoVRfPK7zuw53HrL8lsKKKB+BzCE38V5JFhh7GF8Yn7JIhzk9zhAkUtI+/Fxk+l
XlyqTTsGZxUpnbboN/T0JJ+RuFqmC0o+p6b2+M6vPN+ewsNc1GJVBKSYdw+Re01vRwiURiMmIw9d
uy3K5LEAQdtaO+hkJl1Y4KIpyTu+b6jodbyhIerT9MNrPnlQF2LWBHDafbCTDhIWqa3Bt6QloJxs
sT0XN2HLHx0YmejGF2hvqyYk2kHEI/sVgkpc8LonkZQKsGXKBde8uMsfC4bp6kNss+RgOkQzYSuW
qVw/K5ZhqZWCetWyVdncjjIY7fwkwaLWudp89wpLtSmnW9b+Mak6Lw0/m1QlO4MCkR8HtFtIlCQK
tiEaJat+CBQbNsxM+ST71aw7d2iEXU/gkRWg4xGvKOGDIv26pAsUVtM2smXO/whw8aNvpOnaaNjS
/4BNHaVuMPbCZVs95EBQbbzNksYGKa3hn0AFjMXmVSAmZaeKmDHGz3vLJboJQWx++YE2Mqf4Zi7U
Qid6VVt6zm80E577Xr1S/zrRqTpJ7tYpG3v988TKz3mfcsus+PMAMweRYG6dc7lvwG+1u1Uhnbxl
/6hiyfr7G4HKRN4JjK26GUVfS9f+aOmN5fTOKJSAU75/pKgSVyyYq1UyrHnJ6iNiuO5ZjGxL2OTk
a8orqi+PiBqwW063KTTEn9v6O9VAFgw0EspLnPWqFGpsXyfiDxjDqDlc1mxvLn5zyeXHf3e0aWeu
HtB6maCb0leRuOO/jD9t4dAVKDh/GMEPw+Jk3YqBFJ/hV9AKYs1C03faAmNf+1bv8e6ez63oJkB/
dfP42t3tYB7vWQgn0eLPwdUm1E1x+7zho9aEAitU2q5+rY5gIp2ir+YAyFkoJVGY0NW5BV2JuMiL
qeBKOybjQUqFWHojbinGRL3jxzaebLmDyF8w7ZvRvlemI+MerPIeLXTPLTLq+9WGilH5LClBJmgT
01Stht5vWk00ZYWe8Dyl0uHXsN4jnv1UtxK7T9bxl8Rn0/uW0swhzwOAV8+sTgAzEpR7bWhz5+xx
eOpoj6r0t1chNOzkjjboTx/CptF6V5AAwM2AgdxNSUFDc15M3Zpic++qKgqMsRO0YAqDL6Ns3wrC
R+4H+Ylnhkf96oc6H7sHqRLodvZDLn66Fh4HDVtDaKZmPClloVRfl6S8GrjCRDBI1LG1+GVhc3sH
ysJL+wc2KWyPPRe5DwY+A7SLdzJDqc4gC4LgSc1k6NVtmv5mqAfyskd5jN5UuZl4Md5LUwQcr44O
jqwK7fP4kbmfbrNu9oRMcm+eGPBhjojvL3gxSMmGKx2TqEqEh33jgvTCN2GQzsMSJgOU434use5F
FCbQ6xaXYXk/x0n45rChHTvuPb+HqgcbBiCefEk+VOIlW71lnZtc1UZjK8LnDSgZzowvo2xIBUoE
75IIzg1cCPzZVNO9nWRlwAkR+ETh1Hny9I9BDponvgpJOE2KYNwCRSdYLMewgJJ86hEijYGKa+n2
DSuAXLqY+FbdBSiOwJCBfbo0X+WOdGfoHScJKYwypwzy81+l9veM4v9BtZ0Va11FvuCfuXf9RVgg
NhS82SBUAQEPlecigaTTOz0p5BXY5yDG5np3pBBO9VMIuUyp1YehwPPpkbf91D8wiXG8fXawbMDO
xpFNOA3/OXOchaZ2np10SafW5R7JD73DU1EroQhBFkrwkYKx5PaXGlQ79THDI35sD+xIQipux+of
ExF7CIh1kkZZaixPreIRkRsbi4OsZQu7g8HQ8k57WJBloM/schScAM7fG1rVkdxvsL8SY42oThoz
xpmBgxce55UtWe6ZsRceYxf+PzxoPAsY45dMzP0U5ZNUAw9OKwDyoUzAoDz6/Tkmvmc+tEjmeorw
4fMo+souqkU2TQR+em0xgVEhAJj50ulpSMV6W6O7Znqw1T3KHrHxKpTArKxoxQA4Ja7zjl5BZGbe
EZujFyxPRF2xbkQ/D6LmPF+fy3jJB3IgY7hTtLo+Goq3kpIhoic/b1HTDgf4pjKXM2d4U3Or/9G8
iIsf8oP+7dMkPODy5yXQ/XIR3mq6cQpUUfTKoYef996MMBdJH6tDs8jeZXrpEHOH6ZGI4kqSP4tr
NzxLwZ6aMcgwq1NRIQcMfL3BrANtZVL+qHswKfPlrU/eHccJMFyEz1RFFDDWTdRZlN3AFoE/LSWl
IKIjWeJ4TAXYXAsEY1DoVVFZnJOtWhr0wiScYy725M4i1GZT53UksLrH82jatIdgz+QWVA6YmeLk
JR/F7yAoWwR7VKr7Fxt013W5H8BHhd3gGmK3NH/RKpV5zFshyRgea5gTJ7PA3ajhva9tRDB/lzYj
dxuONal7+LLN5ts9zAbn9UJPuRO600tKWVvQbBrn/xzJZ+ewdQph+QvUHaTnG6CVvONLKCdWICvW
d0i6SxzbZbjQlHe+edjvh93jbABgkvj/UnSZiOxmkl1PugObiJ+jKuvldqdXRKbQMVlyRRXuM1gb
i7dbGlwJJduu3lDnoQFoDk6pF8vVQdknjNOcIsQp+uNJVS0NuDpslx37nGxjSD8aLInCukACsqSr
SJ5uvn/75jl+Pvd0lfXPGSPsAjdHRzu+DW8ri2lu21tVszC3R7+v8q1uRMlXjKBuBHo/Yg6LUo/A
6fBwJzoz02Sd5AkKC1GjgflBxh/byTDjT1zHl5IUsnS9lyJnHUel37zhhhm+tMVcIgOOmIXSelwr
oussz9jU2CG5ELSgNuGMbUv4EnK/sZxFKb3WHPlmrtKfNhHTKidZtuYFlEpm9fOX71W3M+ymiqSf
tW1K0mzn67HM1BxWCdlAygygq8c6VivCT0fgiFPcJL0Wtv4aUtdmDo6g/uy/RCRORbmxm08Ts1sP
CRUk+Qap/OsqQUlpPmza1eyaV0quDdV3HgpsfN18V1g7Jo26NWk8yIdYYPzAYdMpE9nBeEntTHp+
QPSruKUUu1IgNm4v7g1N+v+M61TKUogiOYbxwMZ3AQG51rm3NqAOqQr2ST0LKfhFBna4irdBoG0b
Cuh/qxLYcODC4NX/VpGVsHSBbFDYrqUUiLuccmtdHlTJJY6giMwRfTPsvBxzMZpgiDnopo2061K2
qIwI8ajLKTzIfVpnCEzKADzImGiUtOVm02Iuch4HfYYmw0PAplUk8ht/WUV0c/W0hlcrLfiJi5U0
e4hSWbHThvUEnhi1Jy80wW9a2YMd5J+OoQoWqro+8CtA9/nyF8W1rzgdTECyNQBXpOx15oiG1W5G
lN9LxrOBI51u1nrUtM2hcjAmLyLCshT7hvkPOuuQmPCji8+W+3MdCY3xXgiMadyj/kZEm9E7ziN+
WmDrfZ6sIflVvuCXRNqht6tkqxdZZb67mZW06HWGMa84p0QFWEbE7YNiGeU/YjGHbZnAhM42UoGB
GRfOGigwGKgOZBf2XtfuZCT5CJI+yPl3cls+rkQVX0luLi2+ODuwkTqY4w1SfO1GkgXJhRogjM3/
50AcTE4xJsJba5k5E0ULfb2q72WK2qH+pB+qmNV+hPaChwR2fVX5Xwznav+Ry04CgIa0ayFCW5uF
I6X5THw+JhyH49/pw5i+Js2yt5ZcJdTAcgd0sK/ZwFmGjP9r+35ZoHCATIgBc9k7dWj419CquHAD
81kXvbZTqoCdp3DrkBxwOTPufYAw0lwZZtb66pr6QKmRXxPn2Rq52y6RME+ejKjLInS+neCQdFSl
E61gHST/Tv87TS+BsY9qUKAwxCy8LOnLfVC2XgxktGJlRozqYPDpLIYKpIXCYAFLm9t2cIccx1Pk
oWKEdnaSejbDoHBkescU8F2qPh5IifKdy8vPI2B2MNalNzwxriAuarnEt7iU27/JFnxB4UVZaqN7
22l+tXtmeIjb3TTcKvTogAiZuhTDEmwLFsRqGF0mFts7UZsh3VI+Qv6C37HLsKxX8M1noA0UHYXJ
9FSsi6cQIbbgSBwTDLzF2WxuzHyKIYUkon0ZhzI1kbO1DxLn8dM4yoVfpqUIq2MbpmrsSKughumy
g2IaGeqizGagSahKVwsGUNrW8FvviUmmTd29Ub1XIQAugAqrCXkT8iWjrPftNCD6HzQ2iXo1sowL
yo/viCiJ+xe+OKng1dbUIjJwyZl25r1rdUTBdQ4HhohExv33Ow3Q7LQ/PDOoY/poniteSJIL1+/t
lmp7CsClauJiKgWjoQc+06GrcL0jSqzwzBt6tO7UhmrOSVIGIzgspm3lZpRGVJ54sfd+5dAfhpxT
MErjZuQF/Es3MJhSiIwosRVpkB1g18tGMLNsbzCCU/Sy+bkaUGcyIhA8b+3QIWrX5eMMBCzLh/FQ
5cplHeRFQTRaQiOptEd/v0GxnWH0s4etsiOtd1YPWyCltzb2i/4qgsUAD7b/wXMxN2iX6Le0zoMr
K6Fv4cNQzM0bvlVtKTkgINciTfg2lXruQI7dWRRVqdXrDQzn3ekmZ8LHYZGWpcZwv4G/7x6kgtA4
WRam9xzSKgKHHdkaiLhh/9i0kgUdC3N8s+VYR9z+O5iL7mUDKogvEvBaUrlL4DoYiA836Zq5mOUf
8zu1dgf1Xhks6aPMLlJrIK6VW3C++7iXE84+HElhFO3A4BCWbdkqRETIFNKt3IduYXzStQ98fMi8
NtuRZX02PYwxDXCe6sbP8Uv2WCTrSpsJrR9NaTXRmHbFYD0fzXWjlkDw9e1yb12GUGdffdjp7YbX
XYUBd0RXOd7aQAU9gTcdEMXBLHQXw5l3Ju6CQckQLUVxxUjiQsPF2JtMWG9Z453Z2Ni/68BCpaBL
KRTVwANy0UwwVXZNeTh1BI/jMr2fL+7ElXGeRwiBZxt8VOEEekUGkhZWcUbGXM9CIxCWDQ42EGQb
WNpmJqUWZ61u0JDSbKw+5ft21OanFon5KSiN06bZXLkQDgN2vgCWbrk/SrBpnk4f/RX23jIDqy6o
KgCk4TZRGKGuT90Q2nBlCRefG1C+xUdKvDKcHg2sc6Cz1xzCFxXLaYfC8yTJsdd3oMSUcDgx9i6x
5As3g5y5S9t1p+udgVK0pqJ3ZNJN+jyEWpK8X2QCFxBuy8BSk0SyFqJLSuiv5ugWEpe+QqK1mHJa
+qKQE7MqpRE/e9OGXne2GhaKYO88xBBrJ3f8T1czGfH18i6qIC+f1Zv1FKBPqzOzOuPO68QgDz3G
gXtvtUW7wJHvBwrwSNPQY0m2HzSsCpGvPMyslK6kxApn9hMGjxLps+tvgh0CC0TZIDrDCkAZmJUn
5LPe9MD6FBtTatyHbun++/zkAWjP4RbGq6OHKLMzs420qF3eXUSB7SSgPGVLkZtaK6cs/+S6FxQk
59c25FqWZIDXHIwxJL2VEvgnqiebGRPDlDC05iYL0Z+7RosMu1RUSTqM0Ocd7XShU5vGuwj+0Ka/
wOrBfu1OEqBmVLLwETb6R+pZKBrnr2td1riN5Dp6EC1xxEtoGUmklKW401G7icLMKtdCWub8v7iT
u2t3Wnr8ojpn1aI3RWVZo3MH8VO69Y/2ipFOzFteo5UdioWG0M62PPrcV5oFdouqF7sbmBNqWhId
66PNshlroEWzEm3/ZBc2yyB6ugx62Ys2vq2RO8XSM7FcAN8GuxbgaQoDSOSNRceAmYsk3z7OVvl9
+3uH/Fdp+bOa8sgAGJExd+wAJZIsPViIa+rrLp3vs1ERDaUNdb5NJKRbP09bcUzBXP1xWq167hGP
74zyXXEWk/K1ZqazuJKufxiN4LjZ90iAkJu2ySpiTQYkp+7KMo5B6jlbktPpBD3ZyrylZqh4lzd1
zvOgcP5I0eToKpuAPoyov9IAqggOQ6DJeH+BN7Gv9euayShWdUQAoMrvtFn2BxUTiyQQaaUM1HXg
yybM55MqszrEVSEQpnVqV7M8SKT45mi3TUoktnCsc0vlGZEtYAujIl3giPBbcexE4UQGsjgirZfW
oIoPXpIltT7s6U4QWu7Xf0Dj1dEoPMnCRuK+pG0FpByy+D93Fq2IQXCnVGpiW9eXgtJTuk4PjI7/
daZd8+24D5FJULpWLrA57j7J5PnB9mSoXPfUoZl6NdE9VBh9tmcM3Peu4h+l6mNSoJKVzKBvVb0b
J0H4mI+DawSnrgjKgk8XthD2t0b5doWp1nvbISk6F32re1ioelpp6Zxro7bF6PLgg7DltjonbgyO
U0eddx28IqPe+Uh9R1zcPRpAez/YFgYHaBiHAr+2CVce7f8vswkxE0UgUum9RN/YUtTldulAZDAw
/v9mbn1R8C9SttFR56Y/J+kRqqvJ8xCdcxE1ejp0it8m2B5KyPtsHxz7DjNV6yJkZpJhZZrwSmhj
6eaEiXGGhiah/3SuusLKUnSlmL5vLrDd8yVw0rsIqr2VPmFiH8BMHCPjRckiQ8pos5x8oNeD5c1G
e19YphIgiAXwFPx7Z9pe0+2jCGuF5GzjnRHMxvNf58J1X6GcOEsGQCZw9vS/NT5wF3S1ljjD/jeO
jfXmg9KfH9BmT972yKMR3/cm7eCiCfGwW6QvcZ+UFgN6prwrcmCy6jTYF32vMYVhaivBUFgQY/Yf
mJU+v9zRBts3dd4wJ2LUpR232zTUN1U4bPVOFsl6MxPERHqYO3NB4NTnG+QHehsSTzKcDoX2tfy/
8lzeeeojddavrzMhnBGxa9+aAa/cBrGwMcwBhvkHmuOCcPeWzZ3ad4lLZAj+OLkEZ7jBN+PXlpr2
Kyr1nhvvO1IDKl6YqbXgu3NeAUG4/iIYHBpo0bpCW3cfVs1AmxNTJ2t9EcRPt0lCVvcltDQXh0dS
d0e/NpdZ5QCk2L/ll8JApA3etlhkzR50XCTpvF3tL78kGngEBuKvlheFndiUrYSBQ5OdOI58okNp
oRJQG4QIsvIrho/569UAntNx30uv5agiLf5ESCMj9f6Tqt9Cj4rUzWjFPFX26bL7ZdBTXd0MZxOp
/TN28QJpCcrLxGCEWIdE19rH3TRvG4PIm7KyoIuyeQNI/JeVUxZYDWI3NsRG7EVWQHXhdZJysOwy
GQgcnmUk6kHubk3ZtMSjrbOeedpTv6zK36EvcBlJ61gTsO4b031swiRTXdbvoBzXekXlYop8QzJ8
S9voeFDmcnxEOd2ZdsvRN5pbMXDtFADz6cAq1WYDu33LzQDOR3bqEYhvMo7wD6GQOE1Hl5dxJdTQ
Mb92zpI4mm0SZeTMOwH8R3ydOnAdqFD72jdyXKa86qhUR72mmrwZelsKLKGwFYLpXBC+oPygs7f4
8kfLfQyYnOjJTAdtznzVZlGgc7KrV2VNyugZGls7kX6tJqYfyIhbswJKnUnME73A+bhQc76tITM6
yB77iraY4PRBRn1DlMAhNYF7sC9cDstJh0fMIa6xjzcJK2dA3U9HvzF43m+S0GqmvxebZUjjxR4B
2TeEF3Auy9QVyy+QDJ9e74oIaKJ36Tow7jlmnWC1fO/qh0H0qzVMITrD8b7XzvVa38jg20lNHdMP
VQh1XditqSdtKro0SyUzb0b2MYcejNtBB4v8MJg9SitCsmxHnDH6nrc+VIV6kYfXVO/W2+3n1/xP
9gvulLhBkc/xovOEOBcrwAPa6AdGCJI6DRIs48uNgtwuJ0TMSNxRfKn0Os8SbNrwkN03916fZrJQ
TUOwY+70oUOkR+YbOOOKM3NhhDGkCVKbGkZzb+7hu8tSFhLpLSlvX3n5YcGLZ2wmmG8kQx/r7brc
3epqPoC7jjQRU5yCkn74qjCZrtW3RB3qW+FpO3pSimb0cH7Be6oQ+KkwXNa6u+wwEUcwfWP85juM
XBzz4kBtkkySYGwSfh5kdCdOabqr4dT6QHvWLZm2osNRVFeix0F60kIjvSnTwei9mV/MYS5oxK2M
DH7Xucep/UvGZ/hTyptfuMtLifZRhFHHUXW4E62jsmRF117csvIr3t/CtDO42dkNBaKou+jS6ncH
jAY7YZWPk4aMONSkNKdwiSQTuEtt/DapZxpmtdP6T94f7ZWyOJrCz4CAx2v+tw8VtNCZShFno2LG
oYglNBMT8wVMPg5J3H+UsopQRmAfwphEkLAZjRsptP7BXH5bqCCpM8equsVTj8VPGSKlz/y/9nnz
YTUwVY4W8tZjOohcvcUvLKumM2NXOHlQiboCvQH+I0rT9x7MoQ8mHW+pSDLtXx2RkYccLlhUEC9l
D3c9SZUVcitHi7YysLBhFfkMfet57Ayb6klsfe9FK9SPAFA2UuCS8uwt7ksbrrv91e8RG4utI2Em
KYqdfCvTQO+3kyB/eh3WoIr8sJi3QIwd5QATdQGWRgzZjsAEmT2GI11QyD+4y4b1o5wMWmBUHilW
u2G136M/XtJHzw6SykhFr0Rcxr1jhYc/0/ZtArbX7F0Ja+RzlQ22K+fy55n/is9SxcKCKap64xzS
M6dIllfZeYp6wIirYH2clfDh/76vlK250BKS0e1SJ2rSV7RXDcqaYVpKEWDW9QA89NdPr4JgGFoh
UAkLDb/qRyuFl5WDi51cMattbDGCM0vLvB+nCiks3I8W8QLq/Ee/AF3Q47o+Qm6WZs2+M9qirVta
mB5ySxlEe3WHInIcn+/xZMrlu9NqNi3riCuVxZG4FIQWGLS7ZH09mX8BPlKufR7pNXlfD0QPp6d0
QsEL22Gm5KNmXzmGwGU0jyJeCAS8DQd3hcRCS4UV3omMMjr3vcLqmf8IO9Gs2p40pQ+qEXVOc0Zv
/tL1SY+3BNFS6GQGjWWWJENCzeczGSRBf86R4thpG/CKRIzChXO7jQaKYFRN1wDECRLNkjwi6FGx
I6g7dM1x9nVpzTWIXpyMHLUTZ05vSpb7K4i0qxEpfcc909UtPPBBkBoGASnP/p3fVPJlmrEIKjvu
gHt31MWh+4GKmJkxxyUyySHDeJW/A7gH3dt9t5x+ePEj0R8/f1aITYBmdWRkxbj44/YeAai9E+BZ
MvYzcM4itcay1iLAWAz+jtiC5kpaMJ8RWq0WTdyTZhqUVIM+e3FiteakeVAOyzsfDnht3ubXpcdP
/uQMAfHnQx97UlXBJHcJLGCvax7PHTkndjXGrTGZcGvmLXnMqIA5lAiSZs9ns5HVJ7wyhZDpxNVV
hLeexo6S65umAg0GGAXewIl2JHzJMVk4PMyC4NYLRQYihRZ9bRXKnWcVv3wFWuI/UGU4XbqPXf7G
hwUEEpdOulLF1QUyfHEc7AKQ2tqBcZdTbFKUOHTV/Yi8Y2a70eQE1gGDeN65r3MYArINY/xzmrFD
GkQl+JF/ZS+Ri9bkoiJ/75GUiFdy4FE3n0DXfDGA5z4dUMFagNMXW9LMNhpWa1JsoghyhrLu36tM
1OUiyskv6SzIIxK/8T8S2b8t3DQhYg7j0vaQZkLFpdN3ELGwpfDz7v7OxcWOvSz1lcOhsdpJnaGI
5fQQhTlCRNcmpbg7d4pSIX77CQItS8vcjiU1sjWGmU2XDjwRNSn1/3gK1xYqJuxdT00jD2VzspEM
iL22I7sxzgmvuADQhRNEescoO0sTJj1CI1SjJPQ96zUR1actHo1nuGkMtvcX/tT3Uy/2rO2CGvDS
6Si1hHLR7VmbF3pk848HkI4lRmNs1B23KkQi6rr4LBcn0HApa99vSDEAfWzgodAL78AM7eJ0Wu/z
GkqXQSx2pzOMVZNyGgRz4+Dq4YWnWngRfeqb3JIjN/Ib7RzSvQGlqYot0GC2GJuAlQlp5SfcPU5U
IHBnyfqt2qqqpl9i0OeUJAOVLHxvZ1fKisE425VsUCj+7+ugtVMImWZLYbjSES/gF30B7ZRdOu6g
udUxo+Ld0baOWoHOvSQcXIUvtd++lC/wf5EzKzxRDHTdsV5vus8ByhubfBhWjYzYhEH5DsdmuOfG
Pl7eOUVmKbt8ZzkOuwe6nxD04jc7Nj5ApEQ5w0ysrH3B+CBagdGnga9PRXOJfuMePIF5HwdAgZYf
6Y/j8eZKLIUyePDlhcZTY5wq/Zg+7an7GklxadeZScnqPJmJG2d29HDcuLKFZiY6xraEFkad2X1K
tesBYZhYGslpYFnQ9YdVFRYiVXkUby95cVUURULsfWCncoekn1eUFbJ894Uxxy4j9D8XDtV0xBqv
cwxjCFI5qODAuo9V4aMGdKzMj2U5MrV+cIn5HT5CriB0xCd7iNRa69+MARAGqe/tg0O4DLyEJzEh
KPfl0BWGnOkHBm+yVBzpMQfjyNL8vvFOZv2mtbTMT6GK8M8vsKDfU0BuvkWFhm38dGrUef8nLizO
HouTQsP6GCV9O9MvcQOKyHjYuKhXuit2semlmD+TXgAT8Dlz5eK0rSFsxPvoRMYa+vJwCpeGBc+1
Ym1i7edEspbXhFoK8MB4R+3WPgfWZvs3zgU2pEu+HfQMZ2fQvfMdh9PdFOKSIiiC1SyzSjUUKhMI
loZJdjm5zb+tyD4kppW2HRuxaTK3RvOcVuA3b1qMnVXER4e7sbU0js/pLA3AnvIwRLzrhKyt1p23
g2sF7pmuzyi+SClN2XDIAsd2lbL+xqPFGyTsXSrmuR35vJNbufifsvSepB4wSKBRDE29N+fqodZk
bczm2lf1nFQvxdRJkTH3z1S81F7/AKrg4XWynyRQ0qjojEqHjLRAXS1tD5rQHI8FIAKpjglyU71Q
HOvF3MQQhvmJH9XxIEiBpPW1+lHJmwcwZaoV3tVGwO6Sd0CtSABaN3t/qm6mVM2HyZyxvkw2XWi4
I4jmNSiTEP1JguoO+RX6xs2m7cg9n0XFJ4HYOMUn9kppyNAvkPVxvvgJINM189oSghgosneheKkS
gO4/I2lI+fPbga9yNWWSegwJiGT7ennnIVa1/EA1rSzVAQexbJPdRbDC4FyyK7giqgJsOaUZ+gzH
X00tz2w3aCzfj5s//+uJVcewfxfeXxvfkkEvRi7iBwhd3BjXleb0H+a18Gru7Yqxwg5Jt9SHQEHx
TjWtmauXG4bZ27+QWTmy1DleozCtXSJBBO9XE9OGFEn2Z6uMTqidY1iSQ05DDWH91CifxI13olqm
b5IGZQDoCAWoxfWV3tPSzdlZrI4kYNaWeT5+81BeMS388rfMYCZDA0IDZWCW8h5lDf3V2f12x8YA
yUulGsFxvp/k369TkyerVsZY35tXmJbDaIKk0VcrniQ0TDhpNxb+8Xe7yLTdDeeGJDOb588TOYPw
Ev3p/6DiAsyxVx9PZRbJIraIq1ZhLp8P1eRZmASi1LHMOnGRPKJ78Op3KR45dLci+c0n+pyA3+KK
HZLksXhAzplGR4Q/+4oMA50WdtfnwXF4zq9C/OGcHiUm8okj6nYRKx2BKicNkDZpRXB1RM+PfXY5
WsfXw7jjQu+nVKGGLi2wshdQ6C0aNwID2zaWKRbsLMojjlLkHADKDgB5nnk1/Bt4IJHUTxCA4ESE
57av7TVN+GUHGS0KMUI4HSxJ+gGIvoMOIJiGjXz8pVhzjar7AlKBul39Mrh/77TWQSqt3rHGee9O
V7DzNGm+Klfnnxc2JGCPT4gkkZOHbTzrAA02VAQzwF+Qy8XipAKQeVncxbuRlKLHIwFvLVK46oxZ
ekgjDMJ+oHCM/PKITSzf16N6rPe4AY/jkFKXQyqNH5UFBnuQY6gQWW+bLr61x7xWePX/QDIXjcIo
3HRbt6ykn8gTjzB2xav8vfgGp0a3gPVPun6l7e31r9du+kO9nTG4C2fbtlShXAaU1bApJKY7dU5R
hl67Wdi49V40DALVH1LIHVqz0zTe1DslAifo+nX/RzNjgTOp0hICxGpLhOTYBG1e8HcjUNgPGfgu
Mjhiu9l1CGFm+m355k4r8V9TfgptTSVi5Sqj0F08PGg0FI21CIcPdbi8M3ryARQP+XHjKh47x8Kl
JuBz0GstfnsQM4Le1/pPZxMF6B6GI2xWktdgt5lR3K58E2rccNuoSufh0I3JNml9Hf3qH19wjNnk
T/EZHErrPyxCdMqkFFsg99S9QUOrk/FZqEZdK/iHaP8pQ8bLFmi9KnUL3o2IcPaneHDKG8GKA8d/
0so13ROs/oZPsqjxPvoeJkgEzWdx3f8xQp3Tx01b1FoBoXf7fRBDbjrtzt7C253l4FgGW+0POa2X
RMZymXl/MHfA5cjalsninNBeWrSi7Lj2CE9sg74NVgh9n5sCZxxjqcolmRLpRN5f7xeBu68uItlz
BKM5ojsGbgE3MESmfLtuOM4RnweLg16xrqJARHWRwtOCFI7uFR3FpfmzXPpAQydfadhVBrwIQcRj
AF7W+Ah7g3RSl58m/4zwwPb/MB4aZtPgo//6IfnDo+D0krVsjH56VyqStMTm4SUcFkAa2jt6VRVM
xcJXtGFpNDR84/3pIX1j1LwpG5mnbCe65fKcsB4agCtA9wPDNCSuSHShy06fvv+x1XgePF/kGXnY
FdM87BS7nG627aU4jE5WzcLN8brLlDpOl+73AuDlX5Q5zmPixpIt1yoLxebxZemE0MlmX0P+oDS+
GXQ4Egw6PCZ/mqLJGYiDmudgRIIeBXXE80FaOrBeeHWUCskypRb/TfgTxgpc6Y63brp8Qvfcg9vN
zRx1J0Bv0+Mzvw/U1keUlHXfZj1wboP90cXpgR0jW3KVHq6Y7YW0cpmj7hEOnYpOyOxo9F8+2ka/
oOM8uB5niOoV4knMaJd4GxaLH7sLEPsS5PHuvPfw7FLv/DE8BHOlYECcY7n9HrDyKNDPZoJTdgZU
Y0xYw1V8hML81W5KDQ455A476iNsYbcGgAgdub4RO0k+/966BV7I7wEHLdjJrLttwu5OD/X0iDw1
1dkgijd1GbBjfPkPylHNWEW1woSJVyN8anmvU1X9ZrLtxt/t+cpfIzBWAPcumJ5LWsO3U8JWppeT
LnDjN3Qk4iPvYwCEyHLKOFaBTQ+zdNfrwAlIdYvQEq+iOY4S/zPh+7rtT/Ypz1xncYiGcYO+GEEo
XnN/Ks+/rv1nGnE745qmyJDFmLiOR0M+F0kRepr1R/JVi9gbJHQUrVgvrLTwLLrgi4mVScu4c+93
+DG60dWO+2T98zepJLamGdHchzcUVvmiGzGqcfn4/IL780k6UT0cJfuyki41E2AH0ttB+rm8BeGg
LA1BXFBuzOx5ZTAFHk6exMK//ANbk8yR3b+bPGbcDcHtPeRdd3aPFNt4RW5dE1aqWTZT9hO91xNs
G7/NhSv2W6rDX/z6zSZVFC8q9bkSbo2ftTK5rkAHb3QnIhvu47Fxj7DTedBRhahg7dJoj90E9a3x
UwCQxafCjgJ+5L2qlOPNLA5d1I0FUSRqcHduWJkMNpHWiFVeAKQnOdryiHe9voWg2d1p+DpInWQ8
R7lrCLH4FydkCVPy58pXQrKhghgPW3LfzcVI9Gt8Vf5/96govFs9XyHUvrKHz+Rd5FR8mBbVUmz2
wqk8uOeCSmo3uOVJHFJpQ+pjY/BtBKB5I7HNx3DN6uIlKLenuQBiC/q+7T52SMnLicka+QjjMfI2
v5SdFxQhIUj+8Yh5BaqUVRmRow7nqXecsMrCfUy3vSAHMTvkSqDoj1U5Z3GY5/oYeO6vWO7/PLTj
oeFXdRsDeSVXoHadAx/j0Ttiodik4cSbbVSdyKBGhu5ssdPVHih6WAr8baph01aAo1BLcpHS0pC1
snY+0aKJx7+w0OKyvmb32J2R+BFI5GdUPaTADeto3bzjlHUn5FKEfzv8bx6i8BKtVPhPtW7JbuzG
ntSS/8DzEicTmHxzWU0w7nbw9UoJLKQ+OTpQyns8iSdGik/VWxB7yMYv6hOMyt4VYDYkYTxNFVrB
zDqeBtevBfyRJN/gpa7h21mFfWYbOwnsyvhXVT+XuCRv4mbICQxRpRIhmx+tljCuogVp0zog1QdC
N+rEdNheXoMnB7WQlbjYSMTo1nSwny0nAfhGZiTN4r8PspwkHkpBsjOBT704GC8w2qBX0Gu2H8D4
eJ/kckAXC9crDBvXLTF4Z+S8ml+hZj63VUYzt6/AHVgVb7JKuwvD8TdFS3Scw6oXzEhSYRORCcMd
kWHlLxtLfQ4vbqovQQKlUgUkTE6JRwp8nrujrYMfw3OEYYOTSXOYdasrutUF65F0PYaPhvPPXqtS
8PZuIdbuDo+xPlfth3PYI5utQ3SyHQ8A1mVWgVn3GCWOZlxBmIFcxt17VWDm0Mo84F/IzKyxHCmr
6tP/Q1ZiCKywCSb9B3D+8GJGI8KwcL8qPGu5ZEb9AhRYnPgh9xJFTiaQvvQY693vQRdorTR0H7Rv
/r0zaEd2hnlsE4BKvHF+buDUx7IpyKyQsWGQs54aaBclPAqHSrLtEXBQ+OavbFRA1rGSO5SSt22u
GMCYq7FaX18nEI2qoEzJUJrHphHZQLLZiFvdTHAgVIKTVjSNv8PrTAhgApQFryJOHy6SoNej+y9r
J+xgoIwkhRW0l5xz28YzPrtGcMd2CQALe9GomOXy+pZ/pDNN3nzb1KG5Ir62svcsEhpOxJ1a01i/
an3V7OBX8RW0oSuTA3qW8J3rkFSqItifSrhsu7sn3mZSZTYak4ZuPJ7hWKJ+7hDO9q/L/sYPk44m
raHgJ4ELYLRj3YdLhDJp3AJKwFcD3Pi14BQTue+Yj7ZKhP5/osS8zDmF1WB+cgCNGYZredGETh6R
gA+eV7aQ5sENJvBdXcHkQTR51Bk3meFzAzfT52SpQpNzICT2V7mjoSV+ctd6x2SzaqeTuQviGOQ1
ECheomJucSE6rX7iHFG+nbeyYYakS8R6aMKlFnEhkgN4nt2B8z3Y2DDr2Z5Gcsee6FKHOdkT1F0b
LAey/Dvk+WUNR/oFuWOW9xeJ01OrmiBJM4XXKpFliJjQKk6G0WoMOzogtV9n3XJs5MrWRxQXgteQ
mgPtwNBWKCixM5d8MkNK0aaWgqtYazQ4ONVn6QucZDRw5iq1AX4sBdY6Zj/Hib2NzcwKJapl4P9N
au+ySnXxFswzmol4h8WqyVfwQOVZbgw1tQkcIhObec9LUFgqB396bdlHUnkGt7lg4yA3lNPJeTkn
+BmFWNWZ/zHorKAQCMacY2Ab5PT2bBfxGOGO4UBXYj3A3CGGD9o8H1FUCz/hK5/I6GjcdxYORNjs
A6ehLDzgNF7TVsZTJuLlqnJE3w0guHtJKMDL54DkztM3256Vs9lyOvaFliEzUgNiZ3oIwJKhE8Uh
zPmmju3LKy1lTNPeQ16dlnEUDUsj0fci71R+tFNcNetStQL+WXwXuXLz2QJWuxXCEaphk06Lu+Ny
arjWQIIhS1BRjB6JK9M39bfwgV/Mo4wpH6AhbzVB/pu8iLUbB6eh91Y8FewZeUHddbX4meUWdrpz
6X04TVF+LJ8dnwDkN7MVg/gNcrx8M4+8/JKDkwtL3day7/rn3SAzp63e1FoC1ya7vgp3gi3uwxKL
UKhWnLBhISW59I4dnX8wEc43CNvNTHe1nrXelm7OaaoLrKbRfHitSBSOmCq+w+AZCPIBcQgO1lsu
2+lzY9VCf+nQ+BvAfjPZGBOemZfWJGExCUhB66LPXGf2Ebomdm16dKCUjVP7vQU0t8mVjiXZg0Zm
b9PjtBNcRM5JRBVEcWRm1E5RQdYlQAKu4tPCRk2DzgpBMT8CAYe2cYLBP1oLmXp3/vgTYAuoWcwm
Ynxw+qlRwVparY8CfelBLqy3kzu5703LtRvyovUeUQqWRMrgEBXvAlB6+L51UyRLuwgjYXXOMZTU
/7bl4jYWbNqX1fpeCswael7e9UmxxlLPNNJxAGKjQBkJPDA94yHP9HhKwLOmew8nnt7SEogB0Axe
qUrZ8cdQon/GpR+go5f9eVm0StxAxhcBEbboD7osGnMXCXlduCViTW4ELyiUgIF4H4U5eqSaMAdf
pwbVPrdejqrWMS4unCzK7XhTzt1Tu8K8ibPzxh6vXo7KR0bE/8UBhxiesXh7BBb5cWNrOEnq7gGF
xlfXg55xELqJw2IZo7X7nzpypljUs9WgZk+MLBD7o8B4f6EX9d0B/uEN3mRu30WUc6m6S6kLxtkq
E3jNB1HGodPZOOpOGfy8NVadWkz+7SXjhE7tnJ7dj1+6aVYNCJt5zVHB6HAKnJxkH3kl8GGCtsvV
hjaezC1jUkw5B82QY7uSkNYJ5pQXgOQOXXGOo1vExxf1WP//jEnBHKLpuDwjNPOUdyocvfzaT4/v
t3RMuw0pPLqWfsdhiCRWoCfPa5gl2ucKTDeZBVxacJwuqW+ZZZIMuuT/YNvnntN+wlmiy630IxCg
XpA/v8vou5nRS+2GgY5Ewm+7kGNc6FYrVJYHRAkdo+bLP2qduHse0RxZWmghuPVSpHcIb5qazahx
saVbJxqyIRru0Io6O6fS5pZWphemLGNkGM5f0/JwNxQoykLHhPB9euwvqRvFDk4yyDeGltVeY6zZ
tUI4iKzGAkXxZ+lKpMrmlKdaGNMbUD8OEW4rKg/T3KZSpyGoIYo+yKjzoMbmV8QTCpeTaHNWi/o0
c5MeMAJT7J61ZmpcaDnh/RRIkXS3tr/PXg3vKSr245necBTCbcXaFF9xd1UCaZzqAaeEOIFCwQKi
4U0jbSchRMU4rQgWktSTUBTEBxBNlnjK2RLhokJaEyWXW4rkTxF1Lr//2A8WKSvBD/X/oVlqNlyA
bVfPsjyr5hMy/0tyAhbK4ch1xFa4MFxz0b0YsVrLLhWTp7he4vXfoTdUZL3uEgDLLiHxcbsivyTc
7GWdMBx37L2SUBAxHCJgtICbm4BUp/Ibk+zQj8mN0nQXNY4pVsFY7r5FF+Kt5Q+Z5AlAWYcxzRsG
qbUonGHqtq10PI6yN0gHTuBW6f3SBmuwk7+nB0oV24sLJk53WbeucF/e94EqC4ZBYxSdVnAe8lMx
TByaaIfctermGbnSqNVGhgO4Jttr/0E16ivtl/RZGvc/BbU1Xx3xBCSnGRpxR5eJDYeTumis8dVG
NNZP2WtcNWU8IcU0ybUAE98TIPwADuuw1nfoEDPrZnqe9+zjoaMGK4HgeGkWkVTkMJ0evp82XGKf
y0ysv7tXnPHS/Cdc+/0PPHvrx8u5igHR2HDsDt0umKP8TS2rK/zngcR07QAlqfP8JSVE/k54oRyc
D3HZmhj269zS0ZV+aFo1Ttjt7xxTNYu9lwxMzp2Mll1RkvNIVToxFcZY3PSMiapHaH2i/755VdcG
F38uHTOl5QMnuf7VaXy/jhKKf5EWRU4ky+500TwCfC1PTv2AiJp/psxYi0pzieRU8hODjew8mOzf
PKPUWySvLktX6e1KH5E90UXgGXRkmf+R0HL0cWRvQalne7vfYEpoMvjANquRLGlav+oX3262OuEr
GYUlRBtfeauZNgdJYsXOGiKT1hq8c2zHrU0GMC6a5ofSvdd+qu2JsiN9dqyWmJLGA1YYjbtC7xxf
/dI+u8GWqFJBOP+svvMS4E7KV4SL3tjmwxUHjakF1zC+xIe1kCBeoRbjNVOaoUzRcSIcJgE4wqRm
gF/NZSUCGXq+yN+2GPHVKjwVOEfMfV5QLmSFrki9GpsCGrHTDpJCS6rZI/BhIhDL+VP4iKLf2nra
Jtcqpld3QU/bU6PYp81bFDU6/6vwbsQ/LgkOl4Qz8H3ZDRRxCvWQNH6nwZaPof/ZA+P2K+x5dx6U
9wU2RbmfG00B9bMoKpClhJDnvNKX5Q6iKjfMqSkSSVw8PoqONhzlDZHzkIz/qtVWugd9JzSuzvjl
QTPax7dsYRCcxCgkQ8kTzaq2mnaWXx8N5zr1ojLWb0oZAIk+Wwy7p1PULYUfTuEN81RuMUzYm4dd
CvCUTWbEha/6bZK2bLF+wP1pavZao31EbPNtKMPHFPIjnEC7W7e8OTT/5P4IZ/wCME9zApp+XJ40
AJgIWB7kOaHIoZeCej/Ubh5N4OYpd5IP8Hvs2d6P2pTuuXoIAKZXwpkOvGnCQjIb9GeIgJwzX2ET
wyTI2CqP0oN4ztAPaf5AK5TCZdNy5U95G+J6YvE4fLuIqkqBsSwOfV/ViShPpx0iDw0Qc5kVToUk
4EYxmtdZhjmP1VrIBynsXf7hoxxmreg978g5t5rBGA8QCjjqdgF0cziW9X+9FzQzA3gLEo5ZutUj
hvmN8BAjQG9ECwxEycYWY4c0H6mo7CWibK8f3dz4wpvr2dE+FI5q0iULhQURdPCgnYAf/oKo5/uZ
KWwRT+uPH9KSZDYmfclM42wy+BOeSaSnP5h4H5tRwzZbzadrkbfsoccEa/UbxhIJkO6nD/eSRIwg
8NhFC6zSKYYRKBKT937UEillZh+iCDJJgA/lB+GTHGUJ5buDyGoZN+w+9giugwy+2iSFgC8nfeT3
qbBJY7cYjpaJ25/hbk7HeLsiDg4wBRpBXkN1Bw8rjKUcNmbLWVhRrGkEQFr/DaamRdyZxa7uYNVB
aQuWyL+DHGdNiZx5X/LXI2jxCQd83A5H/7KqhJoskfRwwkdfPihZntGbnsR6Ea4K8PCKEnnmtatA
9F020SRfrl6dZS3Spz091Rmmik/MoUO9OBsL0wvADaaHlJ1zRAZ8u9CGwe1NQ571GEUEoiNvb9vh
LrsHBkegwhgpEvb3P43X4MdvuvzTwKcmQtfCewsb1bXFXVrVx899v09/jfIn3rA9ifpbmmmSv3mJ
/Z7xw+dqkQgpcgFAhqHdmQ6lS1c98tLQ6Ct5+MkyoECi71DvSAQh7prBfyQA4yzxc0g8yopX3XRm
a7pYJoUWrH5+2YiDyMWWwsl/j+H++PNi6AUZ3t41JsatYEQPhkeO2zii8BuyT2a+Zapf6KN023T+
cKT/b1CxjE+Z2YQNXGXFBgVPDyd9d2qQAiBbXxEmkY96KqvE8+SNPiKP3AD3PXvgPl3NOgqu1nbV
C2VoB1hsijzR/66WPy39Qn1nohdqC0r7b+Rco/C//UTe3TFHtU4bxnW7pESocVvYRMdApL8EPv3g
CBYFPlKSQd7DjBZF3wW3ZJ9EP47Dwl8tmFlLep7AAZkZor3tplPM5AhNzuQpBOEpdDOaNSl8c0RF
AGjK8RbOFy/J+ayGNsvbg9STvLcgVzaZo66E94Py7o3qySE7eoP+dMeQ7nc4nrtYFic/PEEVSevi
QOJGtsOAaWB0umkYUy2xCDi1eOPiZ4qA2ocgwxOK+L9itYcxttclQF6xmK3WtqO2Fm/T8Ccs4SdZ
P6wK9HV6x8UrygdfwipZkisgnTwL16DMMi6VlyXXLo1D+IOjRwQlyHBzh+YGqmkEHQG8pFcnirHR
/kzKa6Th6s8nja/Ob4sAwTXJzpQWV7f8xyOENiNqhmZivjFK18TFN2ZiHRRRRBiS9sXdk1Ofy7CI
2224AiKMpS5xv1gp+WBwjjFOqvQiNEdEwaYIxoOqPv4gHUC0Xy1hi8PWmhCFmJoZpigWGugEFW+T
2NWrmbPoC5YG1QrsKWEUKJnafuotg1sWvPSOgI+y8pyi2x8cjt1/Max2fXueLZGeQUMhaC9WQtEm
TwnSwNw3OwMTvw2/tLvGDz7DxEKaq4aCrv2pJoTC6GlE6YY0SLi/MPYpCY1sH9ZOU+5EZ/L9hY4C
kbKojqkrdy5jjzD6TX2r6wvJKqkid63Rxz9698IdmIoc1pKdqjywAaCVEKPDIZbO5+gNfYHVwE6w
BXY+Rz1h+L8DG3rDvypr1Q2uZ6fqhE5vZF98axmh4ygi3VTp7XX+m9WivbSdYYCVMPC+f99RaiAD
z8zfroVMdst7VmTmOsDBd52HIDOc9PFvWirhZwGqAb4wRYWlNLeGRCcUKkzdOqzERDOd6WsSJkXQ
2TZHG2czYlQyPNJeF0bKcvvBRbZIdMHtjSQlnPfIP3nFp43FdqWoU253QCMxZeIqafQ+xBC41dc+
v5yrKpotHqdDQH+VIoz6F+RV0xPaY9TYJSQH5+kA6kWJ/ItOrRajtUruaf7Y6lwSB8G+VdvplywR
imkVZKrZisr1EAAoM6f1VBPe9mmwsxb//mcdSc/gKBmhIm+y0eHT8BtSlIVgL+QGw5nUxbY9DTGf
ZSJtSYp5pqIP9Cg6oe/caftZNFMjmscwEbRS/H986j+LAi6OLl6zkXUgTz21TcabOsjjAfVKaftQ
i0FWTRZ43zmeiFpC0VGPya15r7an9sUFgPrcjPvHhofMiD0/eoYTm/dmUnEP1LP43sxPqe+VXnva
tXiIpd1zwIzy/oWeSuo8qWNv4tjRnDWRM7ZaVhBuPokIsXEUghMu4hrgNbPyBYyBaaAIlhOydfrN
XvM02BDYpAeCuRHEK2qSqdH/yGtFiDgpOFh3v+zMaVWQuIOpcffkpvw0OR+6PKN2QJVG9xNay5Yh
2qyegsjWqW1P6aoWP+XMFJFiSm9SEtANw8uiB5Ef6+58XrhlqCbFRtoc2Ks9GjqZ49PoJ+qS7I0K
OXyCxWxfgq5nVaotxsEuddCYzJShOMBwhfqsz+yO4s+v548KERgsvuCRcfdf5JgTxIB1yjoqNQCy
OZhxycUFlO3lyeHKUDCDT4yPhOUlPXYPPQ+xc5Gio7XgUSwFiXP3Lo1kiFEvriZHWUnEBN78LNk0
DoGyfXDZlVL2lluq0LcEnHZBAnL434uboggMhcI/R7YWsKBP/Yq6IuTUx5YTdg530Izj8tqPedZB
0R5ZYmlOyprZutsplvb1j7bT/8M2q/pdZxoJHQuL9/xh4OF+U1XaRi9uATQsxBdkwq67W0GbMNhH
cUX//B9le046CkksC6RNis9HcDnnVpkgpeJcLIrHWcloROLYP90yrq5B6qeUMTrWveDCjas1yZOz
YU/Cz7w0EcuE95ovu2hzTjFty6dHQWYAg7axnWQPb/BuSMyMyNqD1wvvuRk59xQBDMly6lckWs+j
TloZSU3pM3XuJIwfgd2ZLsQfrOWZc6qxE0ilfb40JYfHBx+hIOsJH5MpsEz4LXfmPzL5JYtwuvm4
QJm3s6WmYAFhNRRHdOiI/FF3UDNTJdomtIgNIbSHVste6obyQQDYj7/sXKDfsX6985vDC8Rpm0xP
pugmLZalRf1EEKxQHDbSfAW44Ob7VDqDXEj4o228ZaipdPZeIbO5CWJ81EgKeXCjydlDQmbdmuhZ
Ljuu8E7d1Ii9oRowYO1GYOnSRRcLNmObyZq6Ycc/bgR8mlc0LPTPZeahbzIApmo3cGl49TYFJT02
zbsSCB6kgbqrBNuNcB4A6vZbAXJP4+k2Nhj5xFGaOS/9e7KYD0UmMIm2gDAh84LmOXP/nHFmfM7A
It4oPtDh2vG/vRmKeu4KkEjsTm0ywgsHTTcdE/S4W84xWtd89OpOxjgitIm4pzWNjLBZRRfWzbGz
lMF0Cra4JwdHTIEyEf6HRINbmY7GEUF29qo+CrcSGM0BxeEVXF+mLN43chzBXEBKk6nwCmTFqDg6
Hkb0Iam43C7kfXT86yLPdGztg5vgCim9o+XeVUpJnzIv5IVqsZYMgewByTbmpj1h/hGsGmRFjlNy
jV/ElyzpfF6Z9d3KxDsInXBk/KRDiQlSsXv9Lf6YGkZvaxdBvZ+FjpU6Itn5VsL0tfT/B3hM4WPd
yZqOmskhJOTXqoVSxk/pfJa2r71GMAD2x3xk7TAbzMB2zTrJedf3PqPJMKr2cBF1oIFjHj3lqpMt
J6mj9OZ5zOYLEFAAApvgt/dBc1eMn6w6igKWE97Zt3eeaNdH05933zGCfgVI07Tdj4DjHuvyLF9y
dlyuVlsNueNHfUwo4FjlsShSbFZDMUzyJHn94+b/k/e3OXsC+ZJiPI7QOaHUa5wt16UQk5wvNDVY
RuGLs/irSaJFnCOkv8eCZdcRu2K4JhlGP33wuTX8B7k/RMpVQhNVpr4IU8aKo/KpPm4PhI9GcE3m
QUvoFAmQfQDEKjgC1t+ndmp0RVipEX3/vNlUf+3uj24lBh28EgP36q1+MjaVFNzE55rAQN5ADHlG
WMMtUOggaXtK3HarYBaCTj/L4Eop42vH3P3E4/bsl67FEO1DiSXL8oCVw3KzK+9J0sWqWfU/YOdw
xODRub25Za+6RygOVtmibxNS0NXrE92SgeUL63Sh2zXJIT1AtJoIbrFf2oDyE6+jiq4AUH2+1D8o
IugMtb5xu6OVQwVVfSvyzNNZW9UiwvdVMh/qokvLKK67VGRteLYsjxOxqlYB4IZKwZ/3tVNwRrTy
MWQT4sQNDcnDnU7rfYXT0siTLGV6LJThMj+pKybdmowyoGnSMjSv9MfW0Bnq8SMJ6y4nY48EmON/
xDC5EqbK1+Wz5NW167a7+uFoP2mfGLkli8UUWfj+pDpncyUsN6EdopUWxGSBy3W2Km4A9CGF/i3l
IFq1qvPIgnbGdSCc9MzdhiSq78DGmqhOKAEM+9kcu2vLWFkNit/bGFDVHjtRH1yGnLsECqoLeKV5
jaaoMFKt3smohdRQWAf5U1sLjP+uRuW7/XuQm5hc20RIHvwJaZ/Vqq6y0WGQAJJVym2Jbs4A4hsy
tR/8TfrUCdWV4lHT83W8m81pA0ri4r5tWwbNCBAJVYbSzZ+qKaxyYOcMR6CZxVYga5AUIACl31lS
QuvDAY9cz06wRsFzatGxMxkZx+Q3Ba+QULSmtKp1UFA/9t7tGjp0jeDXGz/FlczxlNOPzqQ6rLyE
3am6z9RpMfwBY+3ljl0FpeWf6F0LcCHmFOHr+uuCHzjVu1xP8Fc3jor2F1H/My09xZpZJSC6X3lD
FOZA/eBH6OWOJn06aQVXHMYz8CQeAkr4Hl1nrx77hDmYSuFfzOtAeLh6rptw+knOufU8R8mzYITl
HD1FoePxqomlhhW1Ru2V6xGeoYEthT1I6Yh/i4gGYoBYBPzXjr6YFiUAzEMnW8k9RBbuItu6vdBG
gcfV0qusNXFmbAa63uMcWT9UTwQIXKkST7Yu1ZD3S0LEltTAePR2AB8Ayyk1QcQJTxns6lIyYqg8
BmQu+qQ6Ww16rKcS6hvb1zEIr42UWmqFuMOE++g7bQQpNueLzBQYaLNoV9d2oA9mgy034SgwQIrr
3PxOBbAKoy0OsZ5bg0NH52oQK9Es1NQ5YcMJUA84ArjLR3BuiwdoewX24SbZSLJwJnYGBxtuJng7
COXy+TpaLuzhYaAClBhmuS+G6jy3I6J16lndcpLpNgoWLlbRsXx1+JOVxFMz//YbjexGXhxsLRAf
YrztSs+466SxYsNkNi2mXmu1R8VOd/++lFVUmP+At2eh9ROJca9loh9Gp2LPDexHAlahLpA1JIhI
4B7XZIwZR/3mWS2NTorBUJMQmBAYePTbU72/YPsylldA8S6EPLzopsCrfluEW614vDY40A4ADzU0
MFSH23pfFZkky6FQoiNiWik4ILgXra3SbAKY7Ix7Af+Yk8ytplakjSANAD1hBiNEIiXQA0JZPr9q
lqlaolr0ue9bgzgjZR1JUNGQG/WQ3/Awqr2Qe1UU95fSipa8CiRUCTw4hCJoPEqlN6q+hgFpdWOw
CDsiknXW2kQDbNqnXwMPj1vrouFgtuIfvH7o1NvAMLYEPnMwW+bRoWtl82bW8GMdgADdBb5Hf4sx
KJqnHjDlphCI/CCKHLDqv9IZ7A1Tf8k0UOGd+EFEmbVQHHCdZ5649hKFX46GkaMg3aj75Na+hpOU
uC1kF2CWW/dy1ENdrjapsI4qhthES6SM134gIzaIoUfbjn/diRYFDR4VNfxW+bECJcD73+qAl+L+
w7VUprdhq00fqlmHnbDwmBNKiJhORbivWsuav0Gh6VMtb7lrqhtm6ijjPg3CVUpmPYl+ShXwdVPA
j8JR3uN+f0fkhNSXgu8vKv5LVV/DrHKExK98+hNtYicQoury/D0wLQ/eD0gQp2791S0oEc95D+2W
XkGuLn4uZ6VsgRWQHzOV13G+aOHJquZrNyoE2M1in7WZ5x/k2t1Pto11/zACc912myGrwYBH6K5N
PuujRI4pycqqgUz5dA83ucOqlvWRqpwgYNbwMm0OsIp31HSrkSyBY+afjBIJEQyeEOaUUtRx34Kp
69LfUshtxsfwDinPdbJ6uOEMZjGPkWdykSW0oim4TOl37TBdvGevA1nBgYoM2XTlrkUE/wCtGPhN
He9Tr/q9IFMvZgscVZF1SECq5IFSIXLuFUfkRucpOKWFInRLr2MPwNqJJytWPM1jQ2dX75WJY31H
7jQeueA/bKrU+li3FXs6E3YIrg5aITZBiMD300IENVT1q0f8YovGeeCnEHg0kYdkTu6WIkLQbjho
ULWVAb0M08fYZn380TgCk3F7FUhHBdloGv2hWC5Ga2mtftRitpP1NkQFYDMYlztqFOUo83chftXp
pMSJ0vx5YtbPUGTgrrHPnYsHbigp8dmjOvlkg8eHP+LcnwcY/njNPhkXzMN5aNDLioTufMYYVZZz
xnLny9djB1w7ABrp/Sr0LsI7IucUJNtYcQVENpdD7xf15ykG6p4GeL8ueeLhcSr8+STTpeXtS+gm
LKI1CvmISbywgYaYyAvM3tttuHHr9Jo/tEpzYkd0yP8b0kLc6PJRBy3jO8KF25MnypSpz2Joimxq
I0rQW0S9VY6GNLRnoZfCf2YHjcxojFxRPmdxJNvAFCotD7qPXhS11KZWXi3M7H7vsE5a8ISf1avP
P1dnGv7xNie4LCawUna3lAHX4IWRjR5CCSwIONJlUXg5URatg7F+3sZvBvwuh9GK+/04F28rjdgT
sUhflAtd+OPdq+m0OmFsvOD2+iKKa8eoq3BcxGE7Qn852qCT07aOraTgocbb6VyjVpeyHbQSqf+e
zQpci/550PBTdTtn7s0uYsqOvAikn1WGjmhy6Oz/Z1aYyO4cZ9SFk1PJqbmiIstGDpit3CxLSRBZ
/rLftHXTSRbuEalhkid59o6DFnEneMVsIuZXbOQvRuUt7baBaoa+jWPpn/Nsu1tPsSnwqitMLJvL
5VZ9Ms2AV8oKIKqjoa+M0p/9QeTM8c1Ou5zX18LlBhNHWfQawcphDhijafB9Xq4LCtQwIzEvHLIz
As0gifTydkMhVz5+A42He9AVff5YIRjttqOeOE5Gn5i+6LwPjQ0A8DFqYrICyAudXdheAJe+A7iT
bk0NPspBTrXynsvnhexKoEqof5RuDSrIPP4H9LYUkLKTrTxp/k68MDp56fZ8j+SXyePYTdHw5nzU
a4xGn2yjTeF36PZDPoJuHJnAxNuo1JRB1Bky6S5We1ngBDC5JFkBm+v32G1uoqtdasuSff0eLfS+
BFD5K4RF9dx6VERmMnIl2o+1bhDEXo2y1xBxVpe1wuGFjv2Dr4UUEhe0FmHEm0h/OQVs+sGkQt0b
hp7fMrHwwsW3Q1Dq84TSGKjEamWhHVTlDEs6oobmrjoao+LLmPKwLI3Ux6s8lyz01sfQpEVPrvp+
URJ0ZwTW9Exhu3g2lGCG4cEtoFWbsm1AaD/VO+pU1VeBkp25WxOvAJ6Vy++Mf61aUxdShDFnP+79
BcWjsPiCAgkYvf/x3fLnTv9/AoE8SINp6HyBjLqVC+fhpaUdAz/viScmkKOteAo2IIWzmKbmxLXq
9xzJL3MkVfUPg2La8PXYbhwuyytuVkTI3WK/3wWrSKwMBjf+jmi4iOaUmMaWCWO8bj1IIDbRrz/I
c0PDRMpyeoQZd48J/MxBC+uHwMdkYRxtpmsQiGUxuqgFkk2GT1I3XdvvLa+LkjKrx26mi/Heej6C
uisn3gMF+dIEQ5edHq6myrq/J5aWk1SppH+DmxG4lZo99xDaLE8HkuF+McPpIm0mOXG991MVtqyC
72P68a3I4pISvijewUdC9Szne4yRFEq3Tdd81AWrA5SvEe3xD8ncNekxgGB8EWWWcBzZpv2s4B50
4HZznyl2FF+pG3GeOhkyU6h2Zc2gtHqvLwyor5v57gsq0pvDw4GE/5ofYw0YzCJCWAAW927kEuBR
lfSq+7HC5nh80IeblnEdZ0rXCmB8DUICVtalfNYK544ZNhWE3l8+mmcc2q7taIPD/3eweeYnSbQM
gcq8Ur0bZGuaOgdXNPEJoIHEUFsFcDJr1TnLIFrXmxjBDmL6IW+ibZxcQcKl3IVWFB+Edtp23dFe
GSZ6VqMQUnPqhHSZpoPDEYZBcmPVvdoQvL9eZZKLENOIQpjDrhEFZyfRXenHVf2RUql357ni9vrR
l1O2v4J28iEW613uFnckbvzlX1p6DePWy/UHiHYUJdn5petFJWBz9h1Qs3GetNzajzYXlw84u4+b
3A+zubKYlXwQmD574pIeqaoTe2PEHn4enruYtOLETtRV5HK6tDPgMu7vQpPLMDapNrUvkx5LI4vT
HPUVYFIg9132Tu2N3uZ4EQGXa8GR1N5iLBjbtO+GaPJBgOr5Bcgw/R9Asnq/sH1acF2rwFWnlaNB
cFJJGSFzdu2OSYGH374YMvnF4NcqPz2dp/1zUD/VI/LOkFS+8664zXp+SnvCma15UnXahFFyDX6Z
0bOsba4xPzhKZqGmP5tgDsHpVUuTo0YpE6nGMN0aJZYCJM7HEJwASSHXmQjmVtgOyUVmZaK37PWQ
WkNgIbIbF0/EEwV9Latwz339jpNj5Gnttr+IxGp4Ka6/J0UYNgvuJ9y49GTeCLxgfjpZwo4i8okX
6pA4N1x3V8AaBfgkJNsdS14IyaZseS48/IV0D0W0FrY8OGUCrMdVFaLBY4wYo84xcIYvxYTVEUbV
yL6TXykeHGpAeKM2Ue82bfewXoHm32tLaUJH/+VFP0YO2IMAVLA2XJYtCpZKfCJ3z7ZzC+A5H4G9
6t5PzOWwUen3LLFYWObFODhZjB95FQZgKPhXVQZDqQX/RjotaO3vLC4vOhB9BbUSSkNMaiotv71f
g30WSnsprP4t+kwIPpY6piuZ2SB2JZ7v/hGrYm+JxhOHXAe27lOFTkXxVM2uObnhv0DwP+8ii8mg
8wjetXf4nTbShdoLMMCxaRiPtFaL3HXV1ZV5YCw1Z2YZJaETh6Y9k3mxbTT+W8zgAAq7XZZmRlNe
2B9MPnEy3AF9wFlfEmPIjrBaL+tputc/UI/N5Ysef1iwEqQ1xP4x0mx4/cN0IEw57ZPO1E8vs6oW
bVImjPGYIygmOXois4BMJUBvPEd+yM0XnXySiEDKS9XVbUYrM4xZZEQq40bgikC8y+zDqeJ2o0Uo
nXxTwjsoCgL1ENxwHdKyrxWd5HfVeVNqZVCwjnpkSI/jYOc91iRwXiOVe6VmwGIyF+o14xWtpc3E
YEr84SYR8JzYnqpZlfKg1G5nKc65noMRglCoRhW0G7GVZ/pHnt2RBf/b0xDVyP00lLXp7fUvHp/h
I7ble4V9vnhi9SsGfnnpmAs/+j5YObTfMzS4m6uVIKf/OK4XBoI3RnZ4TLJF+JL6PQUi9boj6c4Y
f5VhZi2str22rlc5dBIbkEC0RmSzy5SwZbaBSHPdn0ELu2Z6PDjtk4sifybqRch5gS3CucFzAnld
a7cuYjM8RiiZNlWcRMEOw8I+SrFhaqS5TxYbvIi7vw9sK9IB9b/1Kt2HQ8fJ0BuNxXtDonaOlCf+
PjyXRecoDpvZtJ6Ei/+77U8e33rw8RS37+NM/zC5pY75kPL58nAc0I2Mp5i+6lNavJmD/U4tmVUF
x0CeUT3GnwJe5GSl8ycNNr6JfkD2HmQGuPyZ2hS0mo/SMo66yUAEhC0isDsY2tIKshkJuobeXkp+
QPwdC7B2t6anDdUUatB9aCzRCc+EjRTFING09FQlUwayvpp8XRQ4KJ/PGBlkoXVzk03rzMS2XSxd
5jICRMhsmFxCnevOH1ef/eiDX414lEw5KO42CxvzJZovVi04tv+87Sj5w/+A0XohzOYUjx/6obrv
RDG++B57JEHR8Z3/c4221Gswa2D0Ty8nj8Ora+Fm8iBppFaVmuCB91o4P8Clfm8FkZCuo/YMGMBz
7nLge6TJj/rWEtJ4C0vNoqeJzKVruEEqh3Id8r2nQRxGq4K68qCD2PCJSJwj/HsF9XCsdJK6DfYf
+1585VSQq4FQ5mtpA8Q3o4oojN4aMxxpPsetwCiZeN3bMGzDL8WX2HVQmuimAaOxdnblCfoDUflT
+rIEVG7YMOtKRjK2dceGMnaMDqxUpL2+qNVK1lvd7jjfbrTQIgKOtevLrGS3q/1bcPcO3KSbtAtI
y3ur6O+RLGfLuoR0A6C5hlTAJ4F3iwAFL71OdTtqKiRGEpkNuiEKC0atF2+yALBJ0t0yTR3+kXiX
4HodnXodUAIX24ytfB0/IVWZr+rXIMWbluvNeF9/uVoT6/LH3J7NyfxtTHxsoSgy4nDjLtgoT14D
PLpeRP/Sr/nh3aPItbIuMxwmVo3vDPIFlnzpndzvGeoZ/H/zmopI043d0qhKLkiSd4vojNEWu8+U
xuxxGsif3qpyYk3nTdSpeKnaW5/WGq1UBumFbaD2luih9uo9byOTSQEg/2uXIimvCfl16T3rSGUw
jxTddI1BR4vGnPQWvradjuRwKdrdYeihKP+Mgtf28DIHR4a00f05OjQJYxHsE5S5kamOW03M3YfX
KKn8Tp9hZ/SLnzVsKrGIw+QNGfYGp8+0OMzFz+TPJaEeaJOS8ACDJ/FGkWKavP2ZzaximOhQz++u
EDBIis2Zwb7HScmBptWtPdFMSK+EfKE6nrNr18aJNN/6nJmLev/y12uMkY8relff0nCPm0JxyzAr
Hpf5FLgaL8LYLlF2mQVpSyK0nFuPWHUZiZ18wQBtTTEMXbbWdAbH7T9oljJQijv+X0nAiLe9EusI
ZvWMhGCbwTf4nDmvgGZ6r6+o/uMX5LDS9f9XF8aUp1lVCA7d47sX9TpgQepnI3YV2RGxSB6bOlcT
YYmli+UOEI85UfNy4Fw7e//kS98ZmpQjTao6xqeTd5eqOlalnrIPGMrmZzN/NMY+ARN9+62yqj2m
WfPc0VU9ng4YVKMdP4J9EyWA2hZw87WZOiS1+uk5vObAdyQO5HacPBRHvHhuqdXRyOCvi5hgJkCh
qnecRY7IPMzWfi7MrAnCLwQnOyy7qU4fCdu8rh92WKkwoRnoHcFIS4gAwE88uO1sdrfQ/PDNvIY8
n6Q1cjQ8xDwoaQy7ei+EUsPeEN5COLyFOOMYhbiHTDgOeUCuTJhRHtvVL8gsikza8ShR8MCDKyKZ
Y9l+g+FBO+BY8yUz0QINoY0ptj9GYwJToFR0OKsp2wljrUiEM45TRg0aF/9X11tZDV2CboJOjDty
jXavxR9VFZKpQx05FilzN1188BQRvSrbE2WUSh9WxZdV3k3bVP9ohy9not4j6+1hMlIet1Y8dwj5
kwq6/zuj9s/Mx7fn3pFYZQssC8FpPBGinkBsjva7E4MPUiYAIVlZs5jrkZZgVjboPHNn7dkCh41p
oxwKeUIHWjt2h30d66E0t6f5zlA0OHS/zk2vYIal10L3J8+Ov/FY33KY9XvwzO9l0pcsGDqTtTaj
HcFwD4XoFJ2qKs4eHzu5INPhvuhB9J8VL5//JAKwY0uYTHzVQ6QhHq/Eqk3YCpo68z5ldscY7qE7
FeGx1oHX6C5nc+aJ4Y5uCaX+uQMjhqFdwdai+O0flXh8ZU01tpPLEDkvEVtbL2nwYiYeyVJ/e6CP
dLDzEhuB3EPhtjQ++VpYuvWWH8053/EwZnTUdvWv6AiPhBRKO1mo7o1cSL06lHDCmZ9ZRC8gvbRj
k3j/aQl+TqVHcE8I05MCq7/gmmzLLLW6aO6M871vvXCcxOI/IxLRVvFDemEF09KJrQo3ysdBHm4H
UvLAx2UevkaA5GNiaRqZHapn+kLcunJo41w5VZOsHQldd2Rx0vJVTwFSdkG847+V6GQBfgYKYSoH
2NHW22ZzbLekRmoQ2y/tBmLh/gxtVTxjVnPIyp54oQjOwwlQZE1XYsBfuRQ+lRXNJ1RwYPjK4sNo
SzHzVcqy3xnhT/vKsA3Z9fYakKYQv4FvXK7El2l9T3NLLACLjzOQSQba/jvexXZdAaqgSkzZJHJL
FyVQE9zzSR9hiThW0X51xtOhMfG/TPYALys7sNbWxzUio+HVQob8DnsuzMY7uPLfZVc6pLHiZrns
Ihbh4/ugnizhB7lGBTD9ORZv4XRQdSpIDcna+2xX290nRZHoKpGFEBiVqffzacksQMqNUarakCw8
6xjCv2Uspb5oh64KUeSWEWVbJSgMCNFdAIoCbBAXosFTdH5YAYXtfFqMpoKmgBpRefKD57xuGgkN
GETiGCNbmlAGHW+WobFPBEkxMW0DIkBnoqaAshJFHuI3kO3dei7JknDsquWjNNSh+3KeNdteUISr
OYjai/wXGxHTgU1VesqLrS/b/cdBlFgWgcB2nPKBfwhjPWpPLnJDxTxTVGUILl+xuKoa8Wy1wCJn
pVISrXwqZGDOJGlvEFPpdF+71bOGPrhNZyfMnMtBH9ZiZFP189/e6ohwGVs5zoTjlE/8LbOvb7a6
y4C/9gO1ECthf7CS8Q6xYcw8WQ+YpaNuC5wht5jGRf/BUf3wwqsPuD88O2MpUlyvPsJWbGtmO0xy
7Dia2U0JP4usrtvky/CDdhWfOL5hNOHrEQ0YFL0J2TabkWyRmsnbAD/RkIvmofwdirstidYBlVPg
AYzkprMoprsd9jIllrtA7KbP7zaXzbZESSBgX5FrmXIBtjmK5iQtIDf1EN97Pbu4fvcemvlaz9B9
0SgXjbSiivHrLVpYlhCmT/GrGe532eY+TGaP+OoDRw0u5jxy0zs0/ABdhZ82gQR5MauRrzMtBYic
RpMHIyRPWAV2arIvDH625swK4hBh50MYfkupytOqW41IiRdhQMfAeefPaJvBlEvYHfVxuZFYfDSU
1plcPKwMT0QbqA3TDP4Tq2x92ekGKf/wDCt7m0GNbl6LtuFsj2N3yXQoxdqtstXcgAQCNZsj96Ov
IKR88ReAJbUqDqoeRjbvoPvJ2/ZUsDV3jrZMf9mqxEodN0zTntAwV1KHrPWkNC6tRjemqbFUe8ih
VGa4Rldd+RyzH0ilrw4zoryPswwLGO+xP8siSgy5ohEv4kJrdX/fBZkfAzseflXyii0tY8V4mLRv
fvCS7pgvcj8XxMxrBykuCVIYSvUIQ497mpA2YVv36FwTMmZ1RC9oGivut30v/uA30FrrqGYArLZK
jWlgXKhAxkOwqukzKP2CSOGW9WgtYeD4cnxy/QxJHZkM9uBKwom3KdKpahSD3RI6XwsvLl9ZOav+
HCh8W6/n2Ar1BW4oeHEByDQjarY5247XSGlVIGrM5AMxS/NV47EJ+eK6jAel+Adh5ka5/U2MQL4d
0mgd8aFLy/6XmY/oTMMuNuFe/QRP0nS2Y5u1h0HrBQzhWujFyZ70LhFrSvBNQKuKKHzPoChlTCHo
p4ib9LRVvD/BMx9IFP1vh0pxv6WjyRW587NQNNf8rn9MppGWhPKsmEs/OCKxmyw0yMOLjF10RuG0
/e83FwQFSYLNeLXZOSJIPxZ+YeXwp5q7aGPAoVc/UG8ANd+FOdLv99qTwgqXsmoJv/SWE6xEMZs2
+C2BZye97UP+nMp9lbCylD4b9yIDfpWffJhlpcTtWYpUCnKwG3GgnvqE+VozVIfacnLdFAIbUIqY
msGw1DrUSJcSQUIPjgAAeoSmL2/J7BOALWKhj7mQqEji9yR7NgrTvwPqDpL7Wx2UHlH/OI+cy4K8
byMGiPyygrcpODV5h2GQ5Iy+gM+fVV+HPxVlOC7yO5lAF8WQrOQQZfhGrpiwwTSaCnlUu04ZkcNF
9WQLH34sM5FnaeYnSf4dqnXq+N+kJ49C4bV20Jo7uChmVrQPR5Uugf7ps1AMBoyI16/OwWytLonR
PdBda4kWP2ubUfI7WQjY5Itas4myvY/XkwpI4PtgcVhvCLvjNEeqQ9dfT8pctgvQoe89dNYceXRv
gYuorG/26eHOI8i2JiL19+iU/oTj3R7vAUwdz+KMr/8rh2HhVuHESyWIRc3BduLyEYYjnAGc+8U5
oDUseMzLB78oZCiZZzoJngZerSZnXpLGxV6wL+QdmbQ/KY0e0n5z2kaZcz52kZRyl2jSQk6sxJvT
f8MIY8Mzxx9nEe6VGcvQ3IN7oW1saWjgxTI6rnEoCpUcw4zmiYxLDJeK7rfxU20QF9bGIb5d48tj
oGowzbVlwIHaEN9Iqe91FRo03gpcsRVkNao7T+6r4YxU1VXZC3QfQg2DL0fOWlGjeGKQvHnYKnOV
oe3q1rYd9hDdoXmxBMFGVY5rvznKMssZRHNm/0qsrqNPQIJis1gK31bRTuK+9YluNJxXYTpu1A7J
e2cMNagIyxoyLsQN4BN389qrp/Q3Ojx7fqh7tVcZ6ZfxystHOVTViWSxBJiRDSr1mPpXGforjta6
x7cCat6vpHTWYEP0hX2g9wWTlXZRg6uDsFA9G0LlDV+N/mK3Rp6yL8d8Ipc4gRL89RsYMA6jU5Mw
BTtrkMzONeuhqoSJ6vyN3cfvgBWObT0LeQZCBWU1OepadiwjzGvFqJY+LUhcxOvRh3KebB2S6KGG
tviOiE876hlGsT06+fzcS7+RYyxG0MisuUx5y4341a541O2+Eirs1EKKkGa8Fmkqyhg+Z0NO8GQc
e34H/DAQLe3aaTVZT1ZkKixx25yHTiMGBuSt2/+OJbckiUltaNFSK+ZVC247jUlygRQvc/MpoCY6
E6myZCc0VKAfjY1xskqpIP9FFTyTH1YwEwLoq/P3xAGTHgHq/YL7nex/TlFXGnzQ7bPAUkUlZyPR
8DBvpQY6NYpvbNhz8f+kxxh2qXvNw8RmfauElTyom+yv8RBQMSvFtid75IfW9dbb2cugpAQfiuzq
PN/WL3lS8PjRdaXdgmpXLn0HR2LdKdYB2i5qccwa0tgGvxo9CQj7codYNkYcevqqqC3GctXY7sJZ
CvGUAATAO6fVrriRTEgej1pKSG3/04289S3NVJy2eirPhLVUTIK0TJsRsp0+3aiu6BRzW6EiqmBy
hLIuFEYQbpZfEB2SZy4UNgZ0EmhDJa4oBpiukbbpjZ5BhGQmjERaD8n/1hqQ4poj8hZhwLxJp6N3
OyaJXLis8h8dB2VOuIMfwGmWS/Wu8yT7a0AHKbG+nL+VyEJvaVX0eVIlWRAw1+ufqa/Dfv49PB1z
tZZ4u8IVz1PwFm/9gXC5/StaU46CRja42vcXV/46qkuqtjRH4M7vV06nnojoSFxNmKwdRCyNSkwm
sZXtL32BbNtrwz6LufcnO0/3lNWHmtw9wEFmxEyacVtSwZdgggmgX84r+PwchVz1dBmf0NlwXM8i
047duWdD2hdYc7FUD5lU+HGKmxbFuQqICh+r+EXVD+hgeV1q+52yrwLgQRdgXawk+H4UHMhH5Bzj
KTrnYSsK2Cx03/FMlRUgy9y5N1HqCCj1sDbZps9srzGytumzHBjsFQBHdjCiPINIYvehhjwkVqn2
gEfSAu/H5FJwMAvylsWfBeOkc30e/LEB5SD7T7vfRqy7/o9n6lqVwJFRm9km3QLmL1NatfLOMFk7
8sgEhuzTlVBfciaVv+kwFlL0IMhjdbaCIXA2mZ9Ywo4zw2IwayiRwk8VWtpYMoK40QjeGboqCRG1
61MWboULhOJlw46xG+V0HGwxVOzqsRE3vN4K/+T2Ni0NB9UhlrtgkRfhOk4rFgzR1pOA9U9xno57
8/Ytk5jOTwTV7UOsxpBbn5aBGR14k4E/poh243nQUjnYa44o3nhK5mGO+z/qoRFmEhldrYsdjqNY
NaXoM3tEKRK6Ffg1FTvGtBYAmpuwDU/RLu25C4j3mVsNSw1aj+BbWMLDUn6wqbV4HfLwXZqnHa3h
mZXWidKWIXJtLugZyu3QmsTmGP8iaFYm0teFo1yS2YSj0pvm8wVCgcj9R1mhhFGA18yWNVpf8jAE
1oHmSCiXq7Dvyi2AjsYmRDLyiauyo9zPDVlO+FIXKnks9RyiUouaaymwH4ArOTvCoBBTNvgn8Vvd
oMuVV450AZVkxNnUs4VBB/F40XvPEWZnosyP4arX5x1VZig8Wmjvh1+IylAMkP3+RCSBUvdeizLg
uqPo9YoxQS8eFh8cXcOVGDwiXkhoAzcGvUDN3RL2qkz9mCCkZAuteMWetnSETTs8UllgH2434Myk
2Je5LDlw1uBUHHZynn8+wDeP83phrgXLc061mAjDFg2Q4/wpoc+friF6cScvS+vfD4EI+w+777Js
PiYEM/p2RZSvcrZ+Tz+7dsuMvV0CRUDoD7LOST6/Ych0xZy8RXQfdz48KdpF02n338h9Zl9KWW+s
hvqfu6MrDtTpu4Gp/pmmkEWeQ0DJYSj7cHGXd2mMWiqnxsdxVjMipbMLzbOJEku/Ae7qR1HD2wzX
LqmQkQu8wG3jO0Nx49iOgD6lo+kub/0hbFwaNZPeUa1U69enVf3NltucpadzNDOtxje8LwMVjWu4
OVX2K4yEs9JBZrCWzQOUclUWUU/jRANVmeiH0DcB2q8X4gWN3LBmd99rQTg3PKQcWC5vUcb/s/i9
Qj9HSKc3MZeM/87nPyYLpnWDIeTD5uYag+O9loaEwfj346dHEDYo0td1OP8Oz0gwsgClBf8gNLYN
zBaWXewBqp8RqdZny+qpkcCWKd3pV9I7IBxlwD+Ny8dx+8iy6jeMNCB2PfL+PQ3Rm6ExKMcKb5jM
BnORAz+qmQXdzjWRzU/k9vul0c6h2vvvwpCw9CWPmAreI188OgJRXUmOiz2Jqw3bJJO1MkLGCek2
1Sui56x3MrrG+Ut2BtVV+i4GMvQbNU7/KgqHN1oKNM87WCBtGYn/f4Ka7f4YZl3WON8Uh/xeyG86
Ca07RL+u1/W+TTN4q8RJkUsHGflon5CeL1l0lwMEaqUZrWTXEDOhkzkL/8njI+f60ulF/LGAOxjb
2TAk7N+o69tJycmGDwrN4UZxINIk/WWYDZYgilbbFl4drVEnzZunGqL/f/qm1RmO3NlQCSH0FVCO
hVIvjxLwTW/olb3XQJ1y5MMTy/YgpvTLR8jRPJNGLMrEHn7Jj0efEhJer9fbUBKKbVJ6Y1aTQkxd
6lGfzMdddkcdBXCV0022rbhJc/FSkvUrCcV0oIhdrfEE2uUiwOHfrjfN6rCdYyT1vGECfHP3D0Vh
WNYSWXvMAFkTuohXCf0/fra6KZFD5eaLXhhFbygcHfpVs280v2C+vrkdnuI1+eQEg3CIeERb49eP
Hd8KKrLSUL29qoz9r0ltK09kPVC35Mhz+kFi0yq8sO22AlMTUhCrf5a7fmDhVCrHLcVJlJ0Gk2vN
RSQUL180+RZaOwQpfWhW7HkB4jIHUvYwUWp/bF6IxOwd3A4tBxMbR1OqTWmkOhWygS3dbyromYwZ
iM0GDs9/LCJCcuz/C9ApvpQJM9rBeRGRgoMQNcfQtVasshpJ7nkVL1yqHbzIP3VzyWqB7ibPGEH/
77lqE0SSiy2jXyrPxjinEQyCAfNv3EuVCwbr+iIJlobi29BgoIe/P67f6H/89OO/cfm+bJ5rp9c3
ZjL0e2/THq5LbOGgxaavpCTjFqQW1Zo/9Xy4GcxFITmKP5CAQYGteXkwr2s5Ba3i8/2rQCilL2rH
MWvPDvfMabEbXWuU3emtviL329vFErsS0G/DUtmVD/fvYEIKQoeg1DCdPvFiD06wafj8NptQ1e+D
j61j1sbrLXgY86GzM5OAdN/jLFUCenOAr82Z/lB8L3a3nyAjKkNuPi5eU/it7Vuk9o9vz3RuzsaR
CtTEz5dadQJn5O4rViizxBcDjBTMOaPPn7HRgjh2RHSiqgmnULScSe8fFb7hdPdQiGNmtqQrBEIl
rb7W1DMwo/FnotHd626A/wIwFxsocdLoyKzJEVRD2SDAhFDClOLdYA7uEBH3IfnWZsh5lauDVlZk
zZabn3SjX64bfJc00XQf7YOEKqnNNwiBdkrQ/54cEeuUh4xcPA+8L3puYMYYQU17/y/mFQFNjhYY
8Y6/il4IzD/qhS00FxeLxQfzuVK22ulcn9/DpPcZzMvAFAPRuqP690aTjIY45BWNWPGR52ImyW7h
o6JEE45Jtjv6YZrE/qhbNfvIxBm0NO/GkIRSR8XNOFFNHSvCSyOWqHwy4aaeK6sqDAw8RT6+c2WF
jJnrDyoR73D1ZWg/YiwpX4bA7eg42NYL21rR8hBzxrHSKXoVAHspHm+VHrs9mAzvGfvaYWUxGVbR
xEKo8og9mAvHIsZb30D4fy8k4EbuE7Jn1jz7ZLW1kKtZke15H96BTSdxqM2IxN247iyVwb2rTynC
dHendGtmvpgbxvW6L2QH4yJputETUw9hlA8k4JmmlSnc6Ghmwj/cP123LM0Taau8b5B7QwMvlza/
g4Vn8hhe6b000HY5NnzqO+xuRcJcLVeZhcbKmBLA42ZOdgwDPOpxDncfRww+rDFc+n7payubN57n
/VJl5E1HnYeL9EFTM0qlPaEk/tNMnDQ50iFZ/x4SGkfsJl+AmWiJPIJQNUWvj4Go3AnH7jKI/1zY
EbkZShXztzNSlTy4OQUABnkzA/2ykfArX3hm/FMMpT7Q7ZUm4QQg38HZaPgyCUm4jl66Qs9tkYYy
jOE8sbuB7wPC5FX8iV5em3qpswfRG1KDlgYU7jJV5Nr5KPPQx4aVmFPCtF5wP9t4iKZ703S13a0j
QAM/gN1ImQgQYdcgvRIGSN4NJBjKrASFRNvXk4a9N67vVNRdeIodvSr/sSH5s92YmyWpTEzAXRPR
GtYE4Tvos1wytHRM05Pi1eyetqxRrFkBV6mcywW2TVacRwAzhq9WK9xWgepAEo4zdYtC+liKyfBb
1gmk1cUE5YMm3xYaLQZo8hkaM9beRiqWVGLfvNqJ1ZIGZSgpkruN8C9+UVCsHbWBCmRHLxG9TPd9
Ae1+INH/69ud5QX22CjaMS8/7CjjBr4bMxUnyR/AKgZTCbjSVroZTykzXgM6LD4E/erzZ6C8b93Y
JItj3+VdJ2Yv0+4IVFe972HzC36J9yechOsSGVYU7HQlsjY1fc8YAGjupZtKQFTZwLJU94gdB+2r
srAqkhwAxGSAgPuLYpp0VBYZEJnJWRIW+dcmvI94VufjYNMEWSAly2ASBIVQbBM8zWA01bFaD7x8
XNS09WyMSC5/V6Huvka8vmfPrQLEQDmLfsKz+GXn0bBEYaCZ+/M4WgZDyUVS19l3zgl/9Z87frX3
ayjJJ/mCcc5/VQWeiHcHyGw7rzRSOTAb5yDLFgQ7EOO9j8CxReEI4Cu4FtZWFB59xTs24XiyjXDW
Bq7HWo8dyiR0MesKgeV8vk2cyZpu2PwOxEb+qyuu7civ+/9qt4iVOajLqJ6LbzofCrEeGixNbbUq
hhdzZWIGScDse8b7TCDstvVlUt0knXYpcgCMskUy7vvyFYrw5dQ6O5ftjv06P4IlYwtKdu7BRVjo
GAkONNevokvWTdij7hmZ7H0xnHZUuAn2n4Q2e9n3eGQUds+wvO11+km+mV45viu8w6Dy/0b8l+gW
1taNSojs/I5KAjZDJ8T39ad3IGjz85JlPUhJI5vTtuVVHDdEayLKd0hjTQxVzn/Dh1jdJyDCh1Xs
zL/K66Dlx2l+d8Xu755VBmHD/Dx/7N2FwG9RMJz+zVPOAu4HOj6rMgWF9I5N9LWky8n9tMqImMXC
FP12NLnXjKH8Fyn8lb/3jUoGcrMNUoudfE/Z+zh472yXs5zH0qHnu/AS6WTSWA3rG7KYsAUYRiB0
HUxfURZz5yAnLpOy5jxhVJjXRUVw3EdeAVDlPtel2T6ycS2lM6t8a759aSznk3Me6fHqETDJSrvl
kCOWCQAHuxig8yRNIrBuq82u+kKsRaUi34mLnY0+Pst2nkhENtB+6RhIdMsiMh68ltBOg9olBdCk
LzmEKdw/OXfEchjyNUCHP+dRVsLzGaAHvXjSn1wVtGqIEAwvClhsxlruXhdfj1SmgmR4tpzn9VXO
/JMtLLobAObWAtdLX3aLKhOoOfB+hUgfGJZ21XKqBKfvmZ79VxsmVT+pGX9jVKRj4PUcSixfsjH9
w0NJhF/nM53U7PTvMT71ReEPMI/Lydz7WWv7lXIvqz2QwktCtmqbQq5Lq4SFpMmVmRjB8Pce2k96
Ifxe7okP4pL+pDIUvTDZxyhDra7xER89Yqy70Rl37qBithftNHAI9h8c6xBB3ky4TMyuXSFgpJnc
gGY0SuK2zebSV9ruqLrovSvLZir1FPLDFq/gugFXCt7hlNnUeIZvZIUl15J7NUC+vp/wP5DC3c2n
b6NFbDTT2sAcwhq26wnVCS+nnxEQEO63VTEO8q5mNZkUMIIE5lWnKSM8kCT5D+rP3UF1z+xD2YaM
5mBbwYImEHq0ICCclR2CPJyDZNR8d7Ij23L9tX84LASPOfILK/yPJ2sN06RWaaRa7LtfBZIl9MQS
djB0AF4aWM5xqedD+UsjC3cnyFuYWRwpXcgVHV51KFL33Io3GJQKbtOpNE2KlJKMHobAjbsIrw/9
5W5KLXLcZSI7wd7FM/Wh80jNd1e/8zg7wBh6A2gdH8iuTsIWhAxOeivDLE3NGS1H9ljqwEf333KJ
xjhUi6+MJ8WKcqEjcA+qbgQUzhypTMVF/Pa8Yzyo4q7DgTOyZzkm1m1AcedPNvAHqrJ07c321zd3
pcxiewuWzhHxlUEEZ6d90tKk5Kq8MPpwUYncag01ZEdxwvu845brUuArwCdKUkhTx4i1M0DITcPd
vmjJzFUci3Vxsp3qBauuSjUluB6jLQsaxsXVYIbG5xRWVS8goSKU67UJ9vps6ABiPl76DND10jgc
xE6De1MvI7aUhixlEFfYng4Moj1iKU4V5378oaw+rZmUWlO3Bzggbgv0xTh4/7MgKTuM80R7TO0g
qqKB0qg1+360quNfVas14UBl/TbWcWVDVuoP2AAlyebT5yI7ovbv7lrZswflBCpfaubNkiT6RXHg
nNvLOOf2SnUmuKwyNve1d4xO/ZESRJl3n3j0+KsFcx4O5IWQf6Cj+ldYQoNVi/Y01jYilOEQodf5
jWD3pjJZAdeKRRtR7erc3OPzP3DsS7ydRHw03yxPeKK3Dd1Jfr3bF+TF9Z5DB8imx8lRe7/jJLb/
iGW7xd7jaKdVJUP2RR8HUUh2zR6SC6ZX51l1E9o6YD/BpHOptojpmzF5Zy2Pnfid1VK5Jq5d+Ht8
AoI7isrRpqZV6AM74Tg/qnMe1zCErZWd+HLNqWe8zml9jO5QMhZMuaHmpSMNhG+EIfagthP0dPw9
rdNrz5n+UKX57yb8sJnlptJga7ysJZ7wByHZSZvah4MfPIpwGZ5b5Ie8yv0lQaBTmrPqgmkOnGuM
sQNbHZzJfZlgvQ7ARZoMHYVrxC94DYrqi4wCBULVXLXaW8PfUnz7Z0tzX4ypR70fE6QWfNU2lHCm
6D33jZZTzbr8wt7w3bfYebZeADn1kFVxEA9H1wUkWMyETd+FLAXVj5uHyZcg5gTunDwXTo8VKCHD
ght/yXTlIKVC1Rn+WWNad+j/EMt52hS2KTL4hOtHXZL3vbWR6Stj1fLWKKkGu/kIWMRdQ9NT0zlS
LgRNMLjW/fjLq6yCwMwkh677XoT9uHpixF/K+iQxV7C2V/f6JdwhTpHDVQNAR/E6ClocCBAkCJd/
ix4KTjmegHSYjM9u0Z9IckE3ufYeHX6s7rzCXWizd9B6UwHZHTjmc3mGYu8gQseicdZmeIT/kKvG
A5pELziEclDRgDhRs1pCeZMD8+5B0ob8j0NyNYN00cAk/eERUg87VsQYYIe8Yd17l3l4I/Yq5OAY
ZXxkrjXhcI6gkGnHfGjM4RLssTh2qhQZfzM9ZWGvtVbCFyEiyzT+P/NnZsAJxh/eQ24+BoxqSqdG
sConGUhAveoN8ewGRPKTH3RfGta5Ie/dHeFEFDFSDSSKr3goRzT+P6oqU3rYOxeZN3vyfjP6pFSg
vMTS4nC9QOw+nP3wydTBI5u9p0OM9zGVxQwGZ/gtSGi5rbyq4khbQWxHGv6u/DxCXzoYTVHSZczh
PRxi9/yDP6ltjAD8A912uY4L2f5iyCIAXhuVsuYdDmHG6rElzYCCG2wc+7ltGv44naMO2nq5qfjC
x3PDdN/gR2R14ccjBPbCDIJGSCccTRTcEbpROOuJjdk9B4s5OXAD9pdt8CYQeLpEXJVo2hBkW6Z/
oLc6Vx16QFhlF3rmVpZAlocEHBowAyTP9rRGpRX5+xb7f8uEF0uj1AffKn5kYPUz6M6TkuXExF14
k+oXFYgDfrebk+R+WKjrY9cJwUkli3eI0eCQXSU88e6apbm2MamAPCCoKn5K9ViIUq0dGuBtYPW/
WWU3meg8/yIQmcoaSytBwKob3ZSa+ivyNRBtSBfJEINcR07zI+3kUPclm9OhqkQpzQCLED2BDzOL
zxBUuUGIM1YLBMEeVDR5xFGnmjQswq4oap48CLJyivwzL7J3M4zb/+XnEFyoparebDTcAvTJrlsy
Y1uWCdF+Qn4f9MH1JWeQdp9xIU9R8uuW7WcSBExD7/w+TBEXrEIInzjXHRuLYdDEhfPII73PArVo
kqWXW9y2t2iv3qrwHLZw7kNPwW2tMHfwYpuvQdeQQ4qHx9viBxr+hfMuZ30gkp7/YGGGCAK3jBy5
S8X29BomknQId2AXef5LIMFPdemaCAOhBQDDXFYTla/XCrBByd0jXP9U2leQOKGjEytppe3c+dyt
3kp3V/QIPWvdvLJklpejyqqnqfwOrgSrOYnoersY4/6KT6UnmsjW76+iitLkJBAvfKOT+xI4bvRG
roo0Id+EQlgNwzDKhGuTKJsTVc1Sc5Ggj8Q8b0GmQIoY2mw1/PLJPKf8dx/h0U67+x9kfiyDmrqn
I98wEbP69Zlg3eycUsJur5Gbj8TP65+ItNNQfDNtMPdDr9UCkd6Is0eu+fLOhD9rhC8ZEPa9zdZ7
88Kebu/coeMXWg2dg9WTm6kUwFVQr+3tKmqXV+tC6+/zAONAwEzrHh2zOUz4TH5JwQxum/zGQgMH
sQO5jVaiqxJEQv7CExM2Zuptry/9fLinKHth5P17Xy+ZHf8KWlWa4a5MDZhH2yurDWfkMW/L4Ci/
qDBREEZNuUhYFixzBnQDmuYzaI1UV8sZlOFskwKvZarIJu9lKBc8a6fq1VtmuCyM7mdZmC8GYYIo
GoRO84qMv/0GJHUjaJb+xpS7rrqu1Dc7DJ7lU4ujV7OegzGH3NFu1JH8neU/9u3BL8RGKPkgjqdp
Z2jv/PzZi+Cp30Fn3unu4irhmd2+XCqPommQnd+VXx8cBqZyAvqh1anqeVyOJmfm8CtW016I3Sa7
DYsUIY+yjNB66geeUL3rKJdiJxpgXg43vpoJj1VvRA64v2lw9h+LVa0PAR5nseniTYkRivOuBaQw
BglVwHb+u+XGMVXIMzMPKNCkIg8n48sbGiolZJ12SsHutqnmId64GwxkfiO3nJs0seq16naZceX0
CUW5olEc7g1e4dVGbCw7HLdDY93lxKnmIrMJq5N0Q+J+NhilF8+Lp145JIplqTM8qauhR0ydKcVB
OEH66/fHTmUQhnHUF3DJA/8Tkb2RB8SqBJLXxaFiGT6YhujNoEN3bdLWW5UufvcF0ctkly8ySqED
GQ9EXngQy3ZMxNpo5acZMAOeZClPpp0Uc2XKk8Sivg12oK0v4TDfuiXqlxzxKqUNpOurjIoKRoD4
3gSL74DAPXlkckD8fOO2Xcv4zuyEQz5w1Sf/4co/FehbKtUAC48AZ3MkVrthQKjrbkFCYxHKv7di
pQNgjDjm/WOgjHJLwrwCu+l9aAsEZaigHGk67pqGFsH38irm0MovvGCDqYbBWQTWNs+jWypNnVYg
Uh1kJp899+WvQ24cTDgeCMSQBu5+0uvDIzWsaIFaPZVbJuYN8g0FeI/rMtPeNm4p35WjJtDzUrzw
XFezsl8E252Jfu1nsXR7vXYHQwuE++DwdAYsCn5gxsNAVc2t4qMi3XQ05+tZjN0tLqYL6dK3/kyr
ZFLU6+V+rj1aVhus9KFdI2V0e58LEQ+j6F5CdImZ1PXHM5JvP5EV2niBn3hHf4Um4QWv5ZXfiS9+
mHonPMOs/Ewc9IyxKv/A6StkqxaovmaCrE8ZuXlQsEceS5ft83hwee/njeYHQFiYTHH8xiXYXVXi
eTW5r0QwHZePPs8qDUtkSpPwVtK6QEAYN2gzk11l6KDTnV8LkP8t30i9FR0EhJ+uprmx3ZetJlow
tO50T3BcdAPZRXEsgIRX4t+BamtZnh2ZUig0rWBvWEc9y0kI9anslS+HLo1c9rBXELd+uq8ztWDt
6xXSWbgWxB7ul0u1jf7riNNTuODOQbYsjQTo6Diw7/5Rgw/oZT+nNiP27FQWKUamx1nKvbj++P9Q
V4f6tTOFtOqOxghPnEwF/lNFDVlZLwQlEQEnlraJ5m9nJHaOsD3ZBEcmlNDdq/o+vHXF+WyDgAX1
Cr+e+Dz+NcwgiAHA1/5Id9CYxg9i/y4oYk5ELkQMJ/4YacV6PPDPQk4ub7v1fc1HwQcFvLtyCZPb
fj8ZXRl0+8+rorAZlgRn0k38TKU86c93qy/9x1Q6Ds9/cs/pEjdx/QS5FYVDsuUV1CMJe7sZ1Xcf
1C0AsKGrqxX32OGOAd2AmC8KGrNBuUm9gfaut7kjDDdBmHqKkmTcy5QewkIUET+AxqKF+x8Xz6gO
FmUi6cDNiYzSqAL1VLmyoIuzTB7Zzh8+M5pPA9VW23Zysd0BAKNTegGBZC5O4jGAsJVj9yPBXBxJ
T66eG7X8nKAhKiakOP8qt0fWHjUVC2TIjdgGKDyKsah3YIRJhM9TRc3uwW9vbv/UVmfqFblsYbdg
2YRcAhH4w3jRkbfCR8e1CbHdMOffme1Ir7RvOPKpQ7hSpr71pn46kGZcQTNZeyzr9mDSOucpzzpa
gnkgNQgF8JuTEiQWFwGjVC92r3NsrXDzP3V8Mq8lYt012Mk7RiS+gP6RWdPydrgBRxa1jz88ul4D
1KWY0jzwxjJ5jo6bShdo6TTx2MxJIaJhBeBDgui0ne9qFLutppbLw4+cbUPlTD++kLUg9Cnn/Mlq
LSzC8DxAyC3PolklCmnpVtrlbehvcaCx6kC+Rj1FUdFw+GFUXu8PTounbmA0m3BvZueCq6/9IiDq
NYtO+FhZDmsvxdhG5vk1AKYMkqZEuZjuMfJFWVdpUWA+UQNdXp1r/2VlqgAPuJyfniiq+Mj5hqkk
Ie2/JMnAIhPwd3mokbA1/VqiKcThKiOrqru+dUga1IJvtsoPk5EwL7yitV2XE02K9Jp5xCv0ekeW
n65o7mPf77TB+TXlfLaBZNU23mQma4lErf0SlE8psrgxXAe0m2MmE6lRKktsFxCGMBvsS87EKcpy
ZVGAjRW3tKjUGd2NWZ8l56dJho7BPHe+5JTXu5sYVqlChsL5Ld+x1Az4e/o689XwmmtdPuwbahIX
hfgQUiW08dI0mJNMSPa4pP24plfr1Gy05hwxoQExIfY+GnCer+hNLMaA/pEpf2PEgh9jMVI7eIy0
F9+d36faz5/6ShWgvOTbSP3rKk3M0e1CijFMD1djknFtpeXDGD78j7CqEhFmH+jX9R6uWMxggFnF
u4qRXDgmZSJR0hccr32XW+hULiGls2mKYUo3KF8EiF+qVAp5YmPb+YJfIev5BxsK1wC+7sb3u+JX
ZzuOP4pVj65bqsKb5IDwo1SRC2gUvc5BnGR4Bu12f0Nsi5wpT+AWqjJ3nlqDI0KBoSGdxlXa25l0
OrTNxBI8/7tm37ZuuBSreorLInE/aYBdi+0l61y7wg58XDvztqKBCsFfFO+Oj+ubkZdHAWOMyzKX
2PeNF9RN2ajdyWKT/GsdWLtQ+eT5ZyFZ/Tv16lUMuOCVBPPIxa4x8w3fMFcGoSQJdD84eL3hVUK9
9SMWfi7ugXbaC99mFn9NETB9hy5y6LvHsAYUyuyQZW/EIPq3xZZPcANOkWE+pvMmyAHYX1IJZ7yX
vl2lqdJQZEdd2D+z2SnKYQ1mbXbkT+lbCQQek7KbJf5OCByrRJbzpv7Mj5PTgA7IbVESRqDZOjph
Zy+K3W+e6AYZb+SIiLxSAi9R9Faohrf4mg7Siu/qhFMe3Gv3vBVj4gWq2ZBRTdf2LjaUEniDO0I1
89OJ09WWg0jphSyDJhu54WqSEiEMSfyALt8yZP3oafu/wZr74B0Z+tp8aKw3Dth2xx7vj4DuJWN5
syMysANbHOzW+l5pk0ACSdCB1BuuZxacCZRCh0398RdpgEUgknHlbxcNc4SxxjfvAKzlgX/huS4b
seTycWshRfBxLdIUwF9DuoqSPluqPZ4p3keB8Ysgdkgx9lk5uS95vYi3YO9UFD6MsVdRszouYwtu
TH3Ii2L6Go84HJIgxuKWtjZUCSgzwPXBAx1bhirDog67RBO2tNzlqQ7w9G4ibj5dWmwHPdcw257+
x9Q9uY/nUcxXodCEpLYo3sJT95grQ9s/59uhhj/T8c4zzq3uJNX1or2NjjFQmNZ9MjjbfALAC47Q
JI5Uyn0gPfMM3H0mnxb+1WqNUgfgFg8tCZAZhTyAHxAUgv9TBTm4q1mCCoTE4BS7tjaIZKB32bd9
c/hCMrOPk69/wOfjsuZ7OjrV8IemWwhAsn4WoNS32zPVbK8PjY/lpYSzEBNey212i+iHBhB7LNJC
9lRt7IZKvWGKl7hm5C38vl3h0X8KmHeTA0TpN9P4GvfJybm4lsy7ZxRFdgltDXprY+TeHkpVX15K
ivMGYMM84TyP5tDZvxZXiV3dvZMVtZRStL4S/wKEXESDaPUB3HTehMiyBxb1n7AGt8rxdS3FR16f
4k2eH5VnWrZcrgCIL+jI+VXZZTgngiN4EKERGRLNol+lJTwxVJm9zLLuiXq0y/1tp+v8dF9q/44e
09rClVJq/lwW8k5RrrGtYvhfUIgK5fpbl6HVvTBWWBZFYpw0vc8vEcNfsnUVW0xb8n/OFHy0lt+H
+0dd4MpHuOMmLaG40uXgDwtSBb61Ysa/nUw3RLK+bsRy7fdotIkEee2pUnm3xJG1+5Wk8leVycRV
Y/YgNhprFmuTv1SYT1QqUwaeT6ps1a4ZnhfKn9A26K947ztUXTpiTlcNOIo5BL306QNxtOMDRyV5
3hdY17G39DAq+KZ2ht994TsofFyhsciU0FCJ26vOxrEmWmmciHSeBHv1Z1auJBSs9s3sANutdoTJ
z0fkwgdLZ1uMImEbmdBiHNMSEU6R3SykEgElg4NAB+URi857M112+cr7BWYu0S76hP1oxugyASZn
us25jpz2v3xNm42DiJioD3k0PuMDSdTfWfx2Dtwiz/HdEoHpJCVjNFfnSPLtRoRcaD9hOf1db8Lk
RYIhWzfxS5ZhEjOBg4bkeFeBw2OxiPY9AfBj1xtNZGprk3K3NemcCPKkHWsc2qgPrcHHfgWTSxlC
BGNtpQlB0Iyl6UgILD3ExJJkHRkTjwaxix4vBv19Y6JwTjJI81igcG8Tj9iYktf6jwsS/YkFrhtt
3ZSWPEPst4QSbbOAuFUGLmPm4PlI+71EsuVOfxCcIZiTs6O6KfxRlgbfDzGC1s3RLE4btgVfVHrH
Mx3vchD8/YsRbBNORHRvKY99agVb0X6jdJ4fk2dheZIiQMkAgEmfLNzbN2rBIa5c30gK9DQV+BnP
Yv19/7tmU4h8FE1kuMO3IipJZbFOo2TwvVpFG82WpcfJ2z1B3ve6WjNtX7w/PVjCFc491fiI2roz
gwxxOr/mXWE8Z8C4Xk8GncjD3UnpdZbeZJlpmrICvSTkja1CMMfVQm9S6FeylZQBTt2Q/4NvTX3D
AjxgefH50gN1t6c6UHfpkvkwcciqt4OrG09JBvModYO5T53THm/CHq/IL83Y+hDOvSxHksz3kYti
lwMYL+Y0ecI1VRPJD2heh5ymjO7SeGUxkzWD+JdgigE1QarTNAfiC3VP3MX3tJuNpbGvldEQk7hG
iCmH9X1PsGPJukJD8po2fEFSTdWIZ17ovjRL3JcTB4m2y9gHjJ4vjPkvyS6R6kBG4VflwUceMmGZ
tPWqB09RIAFlDt9bkOSYYNXl7AQE2h21lhbGvgSXdO+gq6GA04t3/9wG3Toi1FHGw4CBXmVKrgYN
AxrobUi4jBPJXytDrlGKYAC1ZWgIRuZF92vU5siwm2hgi5DzDuzGtF7wBifQGUxYA87FSpA8JvGA
BlX9AjqrhSTuxKNAqGnnvw9P3xauZruZlOhHOrjHnIFjTHcqtiM8eoLynfkhrkQeCyu9tW75WjxT
ELzWcSsFmUkwKI0dotmxLwRM6/fNHzCo0Yp+gOkStZKQEKsjLn7NnB+mR+hlSUFGliPpt7CbgSim
cqCnl2W4QCqF33Nb3D/qmqRjkbyvW//jxFFbyTsvqz/Q8UGnyDGEwzAq8iNugUSTny+mbyvvdyud
vw/y/vBIHfMG3rtAdgWMdjevMAS/lsertzPaB7xbT8BlRd1lN8A3izxN7bOHnU5IbdCYb8mcShwn
77nhslVtKltfsBIVsN8YYqdOXifz0dHxYAz8RWxhYDU/5AkKB0XLQb9LxyhSarqYIM3wTPowWg1B
CXKb8PGhUgCU2XvMGfspBMtQK3fi52uhLwQFANy+fhfIbunf6ys1dI/+yDBYvhdh+N+eJ+/3hTel
SmGmbAKSTEzS+3Oijj9HDxFmcYsj43M76n81bCQ7LTpPCz2WOInfVoqvvsygqtdTFrseRFckYUoT
ATNo8RUH3QDWeXOcxl1Ud7amX7BHP5LM4jzAuyI8mybnKRFVg/YU+w64gmnqm5ZxhC/fbVMo9Ozh
l2S9vRnew1M3hgI9LfxjSUqM3JGG+BnCyhQTQG6IGu/HiGO4dT6FdrVdzum9Nlu7bfja3sLV/V+F
jxK1G9/7915hNyotBsIzc02GRk8drqoMLwIMl/iwrQbWOY9vX796Uw4T7hS42DRzBKJUH4rw9Mjj
BizZT3LbBLTuPp0vewlQWrBOsc2x4xt8FmCZxuyGpthp2C46LBrSMd3dOfBT5YrlQWxGT+7Al+iZ
K/xnBHCLL8vKo2NaUobcpamh3uAdnvcO3guSkDti693AiUB1qslXtiNheePA2S8bTEMkFv6mXU+n
xXu+4j5p6eejYwLry/5jPg/D9gqTZaVi99hE3gyNN/IQs9F6A3uZoVEb1SRqb5ZwhGcG9GgvkgY8
QMbZLkpZZAkSZUYLiVH6/NcEuivZ47Iq96BH6OaqshNEcDJTmtz8BXN/15ipIskRZxVEItrB4Ut1
6VwfU3fPd7yF7xOMceCjwAzPipAZYLsxTqkQ5rAYfGSLOcxt21VitdCJo85mZOgTPHFyeDIGRg85
qt7Pr8XT/2HZH+D353xx8rshYHidvg9AszYZ18WdeYtogm7m6BhXm1arh1c1TfGCapCZhbFjh1e7
BWIcVuYfru8SzHsepr/HKPORJ1lkvMO1zNcqgUOrS9hkuq1DOmWoiU6X/0J2m6RRiEvwzGkwYLuG
wFt9sjKF1TUbQRMkiXmIpScWVvftTmkjaRSAM27Q/pt11YbiqfAcqbl8fd8yOGEtY0gddo9XOldb
VFWvg5p6GwmB+NWkpTbR9Cehvz59IXKz6PyrNl/QZDcT/O4xmmQjw6LjOVZprZXscXqis+VlQfCw
SscUsGdnB7ezbF4zQc/fDS0c/Xud2P4WcPZXppK1crgiW7m8kmWSMf+JJMDrjmuzIUKCNdREsajL
aNRdpzu0M02NP2W38QNM4GQYh2k7aMIc8qtucDtcrUZBMmobyKLt8h6H4T5KvFOOgoUnim44FGun
TvIfz/i61CKeZln8J+v10rcWud8M5sTSZjnKV84Ro2J9FrMRBCK6CBkz9a6TLSkM2esEf8atWMJZ
0Gq8DNQpqmllkklyr3yzFSdEWbWpkwAuQQKg2tbWb8E5Knuc7YMUIsoU6lHZcPB2s51PYgSfb2d0
FDps6mIvV0A2E2Y/uv3mSXyolh1jA3uLHSCRM+qtF6S8+j4kHQrW71iqIjiBsaR/d3Qx6tk5ZJOy
Nu247x6tOlyyrd65331fuj95qTOiqgBbYo0iy2pT+6Sviz/O28cZ6wwEKMuY/Af5HuNt2hlcrSMp
TBQUY8DQKYdJfTTQiVjwrBZBy543y8qfBJ9NxIYd5BwSQWrKvOpdULn51/i6dxFpywi/T8VpGhbj
PDjtPi+5j6hgigYNY//dFgTcBrt/Ufirosxm+u6f3e0pcZNWFZdTWbwijYKdofRrU609Y8RAoR8A
X9gBtyFRQPL24HMfGrNTT7EfUH7mkDVK0c7JCfQrG1J2o8xZn3bpRSn4C9z3WH0U13JAVk/FPh7x
vVgugm3gR43lHNFQ2IrrVuo3m2p4rBNjoWYtP+OaM422xVY0bEie0iaSNp0EXeEx85YUGeaQEj3r
Q36jr24az/v2+4D5bTxqIim+yk1TxuwLhaf1oIQBDpH11pkOOAQf4ZE9KzfsEeu7OcBzPmHTHHoT
7q7CSKVF4LRekjmgY5f+4O3bfEd+Gzy72dyDN83RJKZyrF4yecp/5k8GCfMFfuKgWUvIsYxHNdAN
wLRV0PIlQ3goj4WvScZ8MrZq29fRFr7i0HBJbw/sGOOPKiLLBsYOTisafYDLBi1Zrcd3UsK05nPU
I6kmg3U8UnfZGJll8+c+fPp97IPbeMVAYDhST0YkihExcG9/OH5DXyEzjT3OHqeOPfu4/O5ti5iZ
E8eUPwDQKtVBt0LRgHAf32nFmfySTvopizT1mJkNUUka9ldqHNGqyLGwB05uAvPgQAHS/jNe8cad
/kmqMCPIFrw8ZiucjC3UPAAE43Fik6y+aSllrbE0VUTO36wgbc0PRwDFPT02BX2B8EX8HTBLfxiB
AyBZwZtF8bXX/ASmQSHpXwrtv5oKeoQfJRFwzB5rfNqKJjU5BSYm5GQ03e7F+PHD2Rwjx5MY0ljJ
4peKHRgkXum8jIXYVCGyOi+/8xmA11b5xMWNhqOv+p7bReuBrF7KQvXroTQWucBwVKJEL4IuE4Ua
M3xTe7E9fM+vTvxiumW2aEe/9L5AzpwaeJbK+OuDNZ9yJh5aLkHJso2MnRwPKTBz3V5wSCc1PWi9
ZJpZP0QsjEbX4ctd/EmePLzUY88fiUOMTSXV7uoRnoc2UEgX074AE1UbRYGMdsoO9N11wybLkgL6
pw7RItcnpLDPf4UxDyWkLglbHeUm0HYi38aRyDSXb25Vti425uwS46tkopgK9DAC8QAQF4x+Ib2f
r+lXUlGi1cC90LqAmaZ5h8ixeBePbFE0hygtm4McbUuGniNOQHhzForiSNZudxfi7R89mKDxAoop
EGUnkG7sPL9qY7IPaUGiCmld9tPvdeYN2zX6CsO8Y8jv8k7fF7W7rl5NgMsvfrTk6KSLf2PaU5ti
cKwXs+gn2J/QeI5lr7PlK/60YkW443WEzCWLlleaPWPfzGhVfdanx8xfYrLK6nJv+zrZAsy/RnW+
wIF7Unv+5/nRI053XmXsAaZI7l96apuSuKm0xyCg33joF1atXuvGB13pZy0Ld86mP1Qjf9ZzJ8XW
LGuDcX3AB3grRTwz9gYS6BuamDGUnUxjj4nslX0Qa/ned6MLHzYp5avWBctENX8d9o4uZre4hIU+
bFGIla6GVnRhwWOvt2L/iFZkNFNLDrjzCQFw0YBH1VYHTTpQA/4gA78qgOhnChxxzJSdDr11/j5W
k706kYeVSVX51zGGYwnJ57Sm/sWIDzyheryYvX+SZjQ8jtccr9c+Qw/iftKH8nzRHL34Zy90j17a
U9MiHaxkpCA2l8Cr3eBo9qjByfBnu86YAEMGGYiF/Umfx3ST5egYMHei3aEYpFCrqJh+oMsir0oA
ph5e+ioNIwcn4lhkTaXMx9jm2RvlCiMblFE2c9K5Bb0vKwSX7x7tkf0ddVa+7mqv3WD5BEoG9PUr
a1PKypo1EiYkcroAYe8oo5BDytk8/HnsbnjQekhMpZgKSkvDIHOxYQJnoBgpY37htH7TzWRrcdbC
8fRsfusH6tD36o1A8Ff3yFS8FUSfBeZUTUTJsVKVMbstElzqVVtuM3GZvR7mlN6w731lvBtbsAjl
/ZKTbZ1c4CrFfFU/QO1lAaW5p0bvpKW//gGkSzDj2m/aQWbSEyEg9AKR356Z0YKNBwQe9NMRnD6a
sb/LP4QwJ5qtq1LTGoagXTqq8Ihu/QzKYz1Asw7nvDShB0TB+DONrT0VNI0tMZv8BVkdbHp3KNNw
ai2ZoimlcN34Oo2E9x2LpuNPmVcBpTBFJgCarsgLYv4o/sanVxaVsvO5KKEsBJ2pRKonj/8T6omR
JwGSsbpXCXWDp0/kc19njhbx4dUM0mNy7Kts+XqeqK9r/xMgiBmRBH8eCnXFxknPPLdDmYPAXsmd
Kw5rnN56eDuLryBPoECuXfnpVaks5ZBfjVx8EilcPERvXKxp6auf7pkOKeI4iX53iHEc9aS4tjdU
PLfpcXSC0RC8m8+W2P+P5E4k8mllv9jF/z5xwDn7a0qRqikCXp4wDfqfpxMSoMG1MFEFTwbeEGdY
3Kjtx11RoYYQr0tHkNzp1hoAocdc+GkN1V9FEo5ezNxmOVjBL9DUG4w1Gx2Z2Syid1663VIw5I+E
+aC2uztc+lM7rd7GRv1WLB79vnjmdfwvHa9wLHCJpJWlmYdwjnTcYMaVZx8t+Hrk6pHu5XuqdEcz
I5GYIrWXs7kKOycGjzj9KrQ0sqkxVD3SJ2EvcbzH9IS9J/l82+/x+qA7RLyCG4nSTKhbdHmKYEsr
8OOjQKFyT9GL4hY8BSfxkiLXrcxKwBwD9vfSzsBzFj95bipQifT/3UYzomW0f1QCFE9W1lqM5Erd
0X8aGe/bV1a3RtoIcKDMyp4iyC9rLsO7J3cQgadXmZeeNEk2w8m8x3T4gQfRWdSjNgaVQz3pXqRb
rPgWwigeNgVods4H6eT6SniLXrmjunDQnhAdkW61R+8frSEoUAgFza8mYdKoDI1V2cYkHoXmUAri
I7chu6hB4hWiD4NOIJfOgPYeJW25JDCcD5UqA23vyABBuD00gw3J/WoM+xlPaS4Sutl2miCh2YDN
4xllOQ5POrPqJ4rbgvZbNLk3TdPS4SVSmrV1ZbrGANu1cx+S9OuXRKQitMtlaW+J/+8lzOI1yHv8
MqmqBK1PY+3yDdLkAriGL3+MMXMb6G9R4Ydub57PKbSo0aWZX3KRn6MC8tY5gLwtp9W4iGLAOb3V
pvG3M6vthTa64QpmeTp5BFZrcYIRm7J053ou2egognA2gJzBY+JlJpGsZD4gdCZpU8RfhlnJTk7N
5UDG2rDnDQhKRif6GGS24JI4Y0n3Ba47tXtXoB+SidRnLfQ2Dk5lewYTdKdBWAqSMI/Wu0klkmRm
3DaOefXILfruIuT6suLGfrfBKo1Lar1RFZvXRFnWhk5nJ6J6URdLZXOz8oq9vmlm8ypEX99B3Ei8
HKG3nf24yYiN8Udd9EXEvmdG11Ugt5Ydouq74IJ8CrGbpa0jrWurZSfljRuVjd/FarcALnGTH3iU
2gGSLSB38cTBCbmrTxQeQFMQpPKeVHYipAQk0RMUmWTn7NJUZZwUM3fFWqSkqlCv+MvJCC8sTmTw
ZSOQfSLe5rGXkfR8gPfnnXRXqaAcfJ72mG+nIV/oXaOZHaZYW27+C98zArejR3f10d9fNBdWXAW+
Ydd/EPxiITcsGCKmp8wwTkY/ktHXV1wAIfJCiNOEbqTuYRbg/dD3C99RVmFqyVq7BQsQ4u2A/ZTn
2s3xg8sNzlVtBDlH39/xzN6RXCAvHylpeDHCFizZvh5jYFUAm7jATprrCo6Tm/oNNqvvBxaxMvlr
C4XriYujzbyDgG3g4tcAIFKeJSbm+3FDY93oRluofhqZH+uAZaqn3Mu5ZQdJ5Y+FEVYJvLxWBsij
Sen2WSHRb6OxMn02NEiVweWGoseGIesS0HPT37UeV30O5V06WMeP5kQOD3xHgLWzfef4WXkoHPoz
Lfo++muEZYga7KbVpDlVB4brWMTdKy5kFjbdxIWl7yJlmT4gOkkIgM3dG5xr4zQLLEH34RVQEjbe
px9WRju8zfxEmsY2KUloaIPpca3Tl7vHZisD2jqBs+D6b7oMV616011gFNuSjrCFoSRd+MVbdovq
ev2EIF+eHxfyMv+CDkA07Kov+MGABp8CPtsWORSvkCR/uPjMUK36n3CJTwh7eIu9clRcvftux7es
Bo4oS7lT//xaQ8fFPSGHUVBcngVtHLB5qPS5J+yNGC0GvYE6AaWUCF6vh0unMquJP6Q6aV6Q6JFt
dOomSQwYfbdgdFi66VVKawxfpI2zHBhgM1UgkRKsJJTvE+ejbWc6+st1e4dXnv+aT8Amke1vPs3W
piIv2r2prdcNtJa7DoCjfPY+ILdvolCZ7WGJ+DiebRdlObIsWerngl0NM3bT3Ov9pLjT25wPUk7l
uEruQjiYsjYEj1hx5KtADz5Z7AH96ZBSX2wyh4Y23RfTk1PbTcyGktLaIDgPedOwyeA5RJUIiDdH
vhenIAh01hyT1g9PoB8pRKG7j9SSHu56HGERD2E8faTU1/X2l7saNP+/zDWjTPf1yPLERb5F75Fp
hkTiGv5Jqxr9RsFg2JMPaxTqRwCwb0ToUGKRq2KKQgtep010bUmMfJxqMvF43j5WGcJN3iDqt68S
oqdpgiY3hSpozprDX7BqSv6JVRTlFQkDcCYZjai9lVZRA8XXx6xdjJMEVVgaPIPFEn9OM7e9YFd4
H4SHTSU2F6EdlqntFICY/OoBmu/SAJLBTfmsg8mgAxx188RNPpkgmSkiNxO+5/28tzkSAUNmhiXK
qkABebeSuuVnXSNTN2de2wPWdcJk+D80tAp5GJDEDn4oob6IxAn5X47cvQ6H6MMCsLnKXGqHzOkP
hjVkxHHu/xopv4Os5d4454cG/jcDuv8ePcTX9j9ykbcCp2ifR7t224D0GY8yciuif/DqSX1AUeLU
0GMM1zzyx3BLaBcX1ce0byCsig10ADWUIonGV6SjXBdF/CuE+MOo6RyhbeO7xuTmgAsJEZ1hI7if
lZAmI8PAdWbiTkYMBg2qGKd/XNQHzx6c6MsxaGt3LOlcbBfjXqx8satXbqTB18Pm0xjiU3qe+SNU
e4MTaKnOddYzOmmpRhpHdcNwv+e3Cj3UOjFq7QFsDduT6xfHKMhVYi0V9i+xD7r0tcH4MMKOqqLF
3RQSeW0Sk57c8ZaJZs/4XLhGtHVUixGseIyBPB16ZZTBfuJE4vs3OX67OSCbTBi3+PfuotyRCkjs
9Ju+B5fzz44VHTCAobB2s8e3vRJIhzEkfwv1U+9JGltedXq7CSoyNsO02s/BpUYD4EggDkRKud8P
0MRUnMHdEThM3riRkqw2xOEY8GkJ2FPAm3SRvpoqvipQS3mR5HV6fq49DKuqAWi9gciiEZnjIzTr
u8Z904yKp+V/eK22CWUdizqykj4a3BfRhsm2N0c1ML47KHHgDcZ2xWCeAalnvndiSBOTjS4hW942
CCpGixdQh5ZlsFbRqkbw2efPtoT/3pxmHRrJPwiR6uMnlBkt6UFUaQAkwy1AW9XRsR/qUKKNt+Uv
Vk3WmL0/Rwk1jctrKsNKu5HF+RnLPXJEaMUFgQ6Db2oUkCp7NvvS+Bq9nYHJGTt4yQhDElBiLYNG
kAZblnDDx/+RgxKDVDC/k1Ys5pf9r+so4tg4UMrzpffEdhY09Hl1rbpoXu2yjjQOtErEQ0a4STac
y8vN5Kj49MYfbgi/1LERwik1IzTfetaWcCuiJ1kL7DOxi70Nk6oFxc546st8+QEbxEyEbkn4+z32
xOAtLNXw1fQQtoulpCefHql7qq8mqbZiX/2iqrmbJIe19d5a5obwBhDrwUDTaVFJ0ThAy+z646rr
qFGPgKGyU8YILu6tuyaQHwvlE04uYmx9QQ/d2FTiHostT6cgZ+wH36fPsIXP6MS0AC0+1F0KH/Q+
grnKAMKCy5/jLINx1oxNsPAHx2KYPuDC4wXCgd7kI1OtZFEPpD+6qKMd9p1GiidEpMNImXGKAuFD
x3MWV3cGl8nb42ZwukxaBXcEQesTWaO9oCxnUEEdiGsJZeOs5oUYRrJp8w/72vHwQOKzgZO8W4nH
G/DHvAPyBAtO7TZlfSyRYw5y6f1hWi6q2Bu45R4KBOc9rV8QQiioLMI7+63Bk0Tv68jSdDsP5Vft
k31Tqt2T1S86eZHoZ8dd8Vwnw0FsqzBY+tSJglnPxq+2aW+QnSPrnx7WeJEu4MIKjFdynJGrk9+X
bYZfFX33yWBBUjZdfYZ1WV6Ml2+0Lg9KM0U5Eczc4OpEI1WRkMvk5Ua1EwO3a1SVrCH7QOTub+Lo
/O/XgqWnmRLmf3bW9+IOhx9t3fm9PwfzMOUpnN9OBe/uz/PjFV85lssM8cl8ldA3SFf+u+gHxXT/
LlUbm8pN7vbC+5FRJtpTPk+HuF3NaKKVYfIG+lH0zLpAi85gIk7Jz3tU6fw2nogaay+gYqSHcyJh
/uObQKaSaADuLgQotsBmj7CHPqnSurwu+Gc/2p0RYHl/nRQpspbSP2hxpO519KNIbdKknUBCxH2A
xDPQkgqt21bSWt8Yo/MpkmPF8HcJkeG6FDB85Jx0H346B7+p7JgpOkXFkNzzdoU9tEDBE/A8HWDl
woerroZ7ZmYxnhS96LaPINH9xh9BVxPDfBiPthDUj3/MdZuYZlr8SKElVqx6azRoVDy5LAjA8FcK
6xK5qzq609mwuJ9FWpyimrxpqO0w0h9UaKgcSbZ2Ky2n2Cgtn0ZDhhYtudsNDuPzO9pWZnR9unl0
kEVlMiIqY+mZyWEeLcM92vTa/Beuxm4uXd179bIWTO3kwfJCW7yhwZsS39GO52/WS9OYkhOocrtz
8+tzpySrkElwRzU1eAYW2+WfwF4KTzoplDQH2lzt+U12Vij4mH2M3SQtc23herBHXcFM15lmrHDG
aGbyUQptG6UEZC2BwZV/a/FTZP31lmfzxwaNmg5YrAeRdrFLjBXrbKHyzsnklmQIVBfX+MkR1AnU
6LjfCmf3+MsfDGts/COpgn7lu3mRe+3VFmUpSDgaDFBq/FHCY4Lf8Rf4qkXO6JOvKO7xFYa+SlKC
R2ceo1CvoAY/sFfn2xAm94tBXCaKMG/Qw/LU+9FhVx9mSZJRQtBxn38xpSjruro9gUfkKQhO3sEd
Jg+6aGlsp0fTrmaUrYnioU8reddZJ9iko2UiyYU2lT28X8NwrBNyurkWd4ieyPBQOUXWTG6cHYDF
QQ79YMg0m2aSOXwFlfGLkndMkg69AEN1V4bNFpjEt8N/AKsYZwg17s6yAVmf3XwvxYbG/l856wWc
j6dgzhnOefmP3zhPIc7dlh1iR8iX2bnhxPJnzXv9XIWhe+w6pGEhv307DQXHCrkl8G6zrJJ5iWFy
UFrQu8/xQMpn/s7tVu8CWc2T58KmcjUyZUDEskT9M8HMU+3lYpI+qzxrFLcJLxhDzL72zDDjcERK
t4kOovc9ExzPt6WNOWLVtPvQi1geN5LOT4qEw9yIMmGGhHjt/ARQsXm5WSXHeixix94AtMu97tvh
95ufNWGu2mK+cv5t9rYmOitrqgJXSkU7SarmIXpS0XrnwYbZAdt45AlUhOe0QGO/Z7/l4a0zL/BW
JWats3XDaFz8qmwF8PHXTmCfIbD3+MwUubLKxI3lRnw9bfR5ntxUauvdo6GegRzvLKP9dvrTWtZF
KpsG/g+br1t60J+0TkGQD7RXWpsenILWtfyU7y9AkH0O+A+Twng8HmHeHjICslJpnEVK1aQUHohM
iFRS38ShkOOq42hpwPHYpURnnXhFSo6eIfWovm1ZwJOw1f6QU0h2yjOrbfGz0wm7UJ5ZcM/A4ai9
WYa1n6g3OfrG1FYEd3EDD/A7FnpIzE8/l9Mdd/0EYLCOdlDvWqxaAo0MrzjZkA70YvGJVPe0dre8
5a5mOq+KA89Hc5ehbWlakEuMKipzQYrEFa8/TdnB/E78ckCoR+27fJwdDHUXjMdxFWcfQ+KvmkUU
/Kxj6VOXsf+ROSIaYAxPvtYyeynNLgyMc3URnITxQj91BooWk0saTxj5Mp00RbCR8+6jOV5iIJVr
3Sf1PcOehxS1/mFhx+stJsfeHRfTyYULzfpJm0fYCimBSxRSYnOk2OlRrc6zdoGpP0QndOIRgTE7
WzK0KpA3/WUcd5UBW2MHwFF75JlufhYOLLm5HG/lO7CRUC8q6gabwpg2N4KGgXao43xH0Gl+pf+k
7HxLf0p5RnPFeafswpehJq/j2ZoAYslcqwgSoFVbl3y+OFQR8iIqmnUMuLAHkWxhGW9oPA/7qWho
VeKSHxezrbKGO42HwrYNExwpB6hzubH2tMw0nMXBVdmkusRaC3Nu+l4Z35cBuCZPvW6XyIXICBJT
lTYIEE4Dhnhb22R1PWK90RN4966zqRorCE4U7qNi+gqGeSVV5U9rEvCke1kwNwLPVTC1RQZB/tkt
SnUpr2pz4ozy2i2i1RE7XsHFjL6BW73eUOlz9mRCjkUxf90LhMTPoGZhu2Wz5b7tdJYHPuOb9E/F
z5qKpfC7M4LMDSjV5ztVcCswYbV40YvDK5swEt+ZdrRpT0fyrFh1e1LB43kvTTtK0HiK/kMx7A5F
8rfnM6C7LykRS+AzZ9cBjZ8S5d+4G1FsfKJAtS4ka3HpqIoEzpMR51LG0F9FVS4HonzHQ7k2/fS6
OH0aZ9qT9y2d0Na0BvUBf5XKHp0D0GcJyeD2B6QkmitJdcxRYEzb0femXtPd0GTDRTgSVuM4Bst6
k1StfazlVPLeIvCDl7K/H1ywGDC+SaxFbk5F7DHkS1FsUUOGEXFvzB/xkDa7BW5fNh03lDucgpka
wuqSc8TEfR386cI/VoVC5K7OndDqvKy3XQlPumwmW2qwv5Ae8HQXGmk12INPfhWJNs9tQ8X3e03j
LVpcnLKtPrVyfmkk90MiZe8OYOcxp/8/O5RN/GeDnvx69/ZkgY+/otszz6a+/rXISXS6TuIaf5hG
uQFPzcfM/404KKL9jsuryuDsOOpSxdbxQEfyMQ/duF2uAm866iMUEVH8BtVGWM8O+872oo0dL6pK
dVhi3buVuajjnN7YIIFNN2O6+YpOYYBJcZ6YWsb6PTCMu1tvPasJp4JTr7XDRPH0IXWrLAB2k5l8
fwiPVi7cdMwjUw8xS36qKuUuYz1T06wAybA4jWAYemBRYu2pmQtJ4AywLme4CMTUQZ9L2jDgVzSZ
K97yNPcr/XRSogLEEsR9usbFXesm+v9iZiKDYloBUu5bQfWXEGLS63E/RIKGWSFBvN0A2lV1YXyS
v97IgKI8fX6XY2J631nzMebjhu289lKl9uP5I3dc5bal5iKQd5/9HAeullSAB1KDWmF5wqzFMTY6
kETXcvtqpjHD9vb2sY80yFjUlam78TafA3rWgojeDgONWhT3WO8CDzkqMSfYtYv0OCSvyaEeR6bI
W/oKEu9vcxzniOTRc7dYtXYmptpyNUotEIz4PSBnCi8/CYbnljxwjPPahIuoDsnbFfKF9lCqZIGp
aKwL+OTY+hSOeCbGggkTLo8v4ZXsSnV2Oi0qyVCZmvpY/W6WOBCEArm0jXc+Dfc2DZ3KX48M4OwO
pPZtKS0yUaw495o39FCtLPRtY92BWXL9U77nfqOq2NNwRB5/GdlHkapjrkLBcEFaTQEQr8+QdFl3
RQjOUYHvo3LwlKJBLey2DNFv626junKT0ndEMqFEVfIu8lYxutSlq5mwH1WX9+UTYURpz/FIuSud
avZXS5nYbzuz+PmsxJEm+m2zzDqzZum8evMGqvWx9yHsxHlYRMhs3W3l1n6ZsrPKsSyUsXNaBJJK
+2Dho7O3MYPlc5O8El6HnDD43C743pE8FjbB7jDx7knWrAmaeu2umf1pIsVqKAVzPmQycThCA4Wv
huCy2+Wd/9eWo5L4jjOszlQoMQivUnJ0QoaY7ji8oAptPiEtmvuvFubQy9YMTTGVNJ7lfx52GdU+
vjk6XvRd1iFj516UgXTh0CsXVMOrdNA4r84b9VuNsCfTrxq7O41P34pCrz8Kam7WVk23A2rmL3NN
WDcWw0ZI78/Pa/x7D1uh5cEbzy9fSlJTG67/e82BT63yd0PUIap9dsPAF5dQm9tTXZM3fFhmRaaP
1A3r1/Ay7nS/PVqX1RvgnTAnAl5rFdr58XaieFv6HE6o8zI5FXRxJzzGcGXa+nmnm8axw58jTYTJ
QNCmGQySOqVUVHJsPOWJQf76wWpAWxoECqA3JnKp4dESOlwUkFeVmbkRBlTh+b7bGBfNvqEk9cSc
zWQNPNFUeOMVcspxepA8wTkTJaD6okm97m5cCed8WBY/Ti6wEYUfNcMLgruGYBcV4/Zoi/MxFrjp
hjTF8TkY1kdiH0mTW+1Nm6u2doYMmI9Nw1Q2UqtGVf0P1bLiybMfWPuCD7PxQuHAKvS/FgameEDy
s8WEqjHhH5uyL2WSRsezAsYVZTX9xKDhJsT/hTF3c07aQCxDk+Lyee6qOTuWf35cXaE65ceIH1Md
HCd06jwOfG0j++hH21mzMrbB5Y/8piSmYx/t2BnMVktL6KBJfGQ2FvYJWcVHZagA4OxTfiuwgpWt
V/XkXG7mLxA+bE4E5dMvGWezB/rXu2KizNF8rSWF++WeWMYrrkgsTOrYiWn9zUqXg+M1jhyAOwRb
lZQ56s/cBLEmn/2ajxtl//nZkY/K2JaL5LR9QwPRhxSnBn4E4/QzM4zaw+oMFOEPapNh38MC4ZSH
8sXCBTRlOUjA1UILFl/es1ZD17l9/srs8LLRUnDlgT8M4utUUhK2GiRrRJhsHMHCTnfNQuobxzkq
YNfxbiOHp6R+8vRUoseAUxGMCz64HQ8cIzaer8ChCu20UItTGMaCx3M/git+eaJGt+gHTsyso0S7
mruuM0PyCRokbWnbO2Lkv0PrNnSRq5PVRzIYrEAYXxfAc486Un6QBwRhFqy/713RfzDB9b6D2cF+
+0s2NoyEX47PCNPJUjrZVhdOW5R4TntuLwhH2+5g/PtAg7x+PlsDy4mlLAfzpuKrvHwOzFSV2YK9
7HEMSnl3/A0xaIVkG0zyMD1ITTI6idppNcGyh5ZvPasPHvcpPL4VwFq7zkRbYyYiTzG/x9psGHcw
SITtUNKHXlXxX6FYnzz2NeY95UNmSnAD8c5WXCzbKXBEvglJezrh7fMwEWj5CfeJEtYZzp2yTwxj
Si8t8NSFhu9t4KRtjixf1ADTMLSCOhWbgoGCzyl4kXXe3pVax6pMQAy54LZMOn02hzJWtwr7gywR
z266TO+n1bW6XDirCzKzoR/HxrctC1tOTLzDHazUWQwk4klPEeA4wheFkmdztque0ZoqGAakcmRv
UwhsuYS8kXyCFf4agqyF2XdKlYq5R4E+H8vIii6iVrVT8rJQS5l3q+4dTbi+Z94M8bOLra2YlVaa
XWzN9WnkpAEZxH27ztbE863R+rBZb7oUZciRdP6OTwHL0NaANlhXVjYYULUBkkG5f6eUeqKOLUrU
oEg4iNnNWj7VYNqJRQ6zci7nZSS7NgGEQGSo78VfQk9639VQjQlhWdCknMHSy1VznmxTZZNs0wWS
IVSKFHRlpr3mgeCLutDoOh6E+BUYyfyVcF8+8x02IHeplD9/fh5eb/Vf4x4dxnr3Mw67DzauUvmi
rI33RZA2ROQkCXbWsMVcU3132mIJE3FYGlaiqf+5zwRtQkFGsicuxKDrPnIMwGCXOb6XmhQRRFkY
Iy+Veiygd/JzL4UKEyZ0VcaWjj+ZfSy0nL1FwVG92PMPdA9zKCPqc43LgHEYnflIp8HC91Mb75IS
4SFf+aRzA3u0gZyt/a2njYRjbi2nIlZ2VQ+OM1vP6BdzSdC4FmQFjKaSA3rTU4FkblB47SRFB4FL
Yz3zf4LCHmKxcV9mS0HkkRiLZidbNKhkkQKHenovzgngC70PACnCwWfe8Lnf27OMy9W/S+gq3VeU
XMbf0nOxgI1WE0aDSrPtK9PA5cyf9WWwAIpq3dha60VE3PzvEezxPfs15uVWMjlHncqoP+U0ttFJ
eOUvp6QT+i7p3TcWi/lDdJOu7PUcRPTFwQ6gFfN/YkIEgYFJF6sG48Sfz8AAJRUrJeTP8X7Qj+K4
4axIeKyPmm4lPjucspoeAM8xLVD0U+PCt1RNnmS7rmd14JqUXQpKDNryB07BOlNMGH9IdBq8mzpZ
2WJfVKEamqOz4+quplrSk/rjs1kPooOxmpfJQWg1srtc6Wg2dU12QN5pPUU7vX5nLHBGXbo3LFKL
DdAwnm5yGS3uJ+iGq9AknRfMIG7ic0jJNO9tWJIE13FSPKohGKRzTMgDZE+eNCpVXbmTiN/TueUl
muF6A47J1d1eeyapsB71suXZjRKO6t30bAXVwkGP7fwUMwY3i8P8Bipx0vDs7lZn0lyRaIwubu9p
hHoKrMnbuPcwz93XPgXgpV6en660ZCLGp+8DfJsQhLpPaCKec7NTHBmCpzovdr9ZOjcdfD53IDb8
6e8FjK22Vyfa6w8MFi44OiVFJ8tXZXrpO4Nog6u2UQGsRZt71Dm/K3GyqEs7cl/V/LmSbkbB2AXa
mThHgycIlgfJdJ/ndJYvQS2V2ZSpa2iLyP/IUdJ+xIyXGTUGgeE1+b2oH80dVEMrH3DGQ5vx6SKZ
glk4q/HWuqWnYyXyCse9H+u9Eqr8Kc3AKT2Y6farUpKXRAJyY4RXlQqBEpazJmjKyh59vRviREQi
uFAGmOBKF9jX1eCvVeQjthu0+coscQqH7IeZ7dYxpI+Ys21Ls5hohflqsQ/7a8OY6yLW+qc+m24h
8LS/meVkNkDUE6lj2Cjim/qzUztJJRdr9Xd7p4yaHzS4yXw+EZIjAmf1XJ5I9xgjd3Zrao+KyolS
Q01JECK3QlAemA57vhxblZzQLbR0Ib7jhq/O1xJRvBmjF3uCeeM18eo2mlB9lkE7v7+0TSRTAtH/
vJG97QRC8n/99mrNwYSBfQutw9UKbHQV3BqOk+NFic4l7YZKwBByf+DyqfY6bUQydoYcv17YaK6q
as7gwb/Tkeopm6LemJ3m/CY90YAD4kdSJF3jXvpSuWfOV/00xVbk1FZOKloAX98b1ujK5E7TCggS
4NKaeDCBwGKGgyTBrsBXktxVUVESqEWOuoiV1OiU7H2hHgSiG62fWOGAs1ECusKfI46EBhP+LIUd
11szXmkNWqRpaNpAZCNTBoUD8DLSfG6x3EEJNJSmTShQ9FieTE9KxuoY4sVu8l0EeqagHIJV1CXC
BZ646B5sMF4AyiEcxHsusZITtSp7WXz+Did3HjjC5M6NWA/wCrowpdqQ99DfGEkilAtefrZ1/1HF
CZMfGi8g5Q35JsPr8K3rjGDx5yo1FHHJeHOgdXDTNIn/WaI8uqJWzcF+7MYGIVt7QhmV47DKUSdO
1k0HfWzfh7ZLZjrDLruwGf9ucah+/663ZKbuQ754WxiE/L//Ub//5QFut8UNh+ejY2ix5+bXxetU
k+qNZWBQZUh6Q36ks0vkBdeAE69UtkxstWPS3buwaExMyaRfnIB899Hqt04rTo/O/CgOBUSR2mI+
ujz0IK/1R4ohBq+vSXW5I5gji9qndPDJ75+jYIpzKaIdGJosKtWZLv/peh20NChghb3BG2OpA0K2
uD4w2jZtgkU/zdtmru83sam0xot2syIpFV/Ufvy35320OMEZGxPZ4L/LiCvOTPpMwPbfvPn7sHm0
3RvXWJ9DioGIjGJrO06BkfSgf/+99IRrTHWa4UvpmWswC/LAF2BUIfmGb4vsloDN+aU42dS9ZFLE
zzmF9XhN8zpEOqyzFFY974RTZ0nAOShH9+OXCKrbdz/jaFkL468VU2SO82u0VMphMgRwBorkfLUK
xk212Ox/1xCCRZn1S0RY8MX1PBpkO8lwxx8I0OrynQsxUwaekonJxeG54Ho/bPwIkoPrFwtfrofv
JTguPpqpJ+SqHLzpxMYHXQnda/0d/qnPhJvJMcnw93W7fMZwirabGLwwxmk4yBXYvkknids+HIqP
DbfWc5Ns9kT7mXgPgOcXmFiYWaGdT7rhOtF+8l+wGBWbjLuNqGYpw5fnGiPTeVO/5ee98OZRUt59
KItiRQA6wbLYXPq4x+04K/EUEu8MmLDWftEA1YD4LtCzc2+dOh2WAGtX4XO+GkM8JoOlbPOEa84S
2EgaUvTPL/5PTUsGnTDCdsTwxgHlL1xsLaFTCUG8GYIqu0jKg3R5hvCJNbWHL6EjouYmfyATBkmY
/5Lk5mZEHSzetcWESWsPhLTav3fK/jEHNxpMSpYfwxzWrhUxrAshsa4hWvIaKp2gurBmxeFcuG9o
V34bntQe2Acme5q8Fdz3zcihZNnP+adI+Aca6A15Ref+PFNiIEB23wfbKvj3rQsrcgT/k/CrSyS1
kMMvAkIbENWzeRWaO+Wq7GEN6Yt+r35BvEHva62Wzx0rb6W2NySGfRQxmXAIv/oAoDXQWJQJHKHV
dlomP3Hg2zHnzz5BNQu2mod4v8KVY3WvuzqnQma/9pXiDxRC5Pd3kQwEp49z+69N9jTFCqn27KCB
m9Cmslq1CrKyrfdlCPT6OkuqUeOpBUtvmxfriOY6wnxAh2lPkWY4N/8qCd7YZbELZ294Nl8stW1Q
AjECTt13qwyMVuKfytSEWkZT2qXJ2mfO5LNnhu947nfMgZDZyPVDwfwGLCucwSsFPYjuu3XJh5Mp
m9Ys+jHfRQ7aB4cSpUaYQj89hY7UfkVoCpkyF88ITi8k3AmWcsJjnSnITtXqvpmAf7MYX1oiWi0w
JY1vFCpBn0QfVxG+Fm0hOKiF9H/qVNWEjP74wgop2CvM4AtU0RnZOd1mnjjTynA/AtjzNpJAEfaP
yOawo5Hxs7Ah79r6XT7ScqPq3Z51N8E4r0mK9GfsZDDedAxM6H6knDGbRcnfuwZ+H09OS9TGQ/ff
tlbsOHVZPEBTz9MVkQn3gjsC/de0DtQdLcZ0KbrB2oAPCufShhNzcsicqmWS6wK9juLcElhfJ5Sd
i5qxhBuLmH8rhbOlhG2l2RvlXbVaF2VsbcukEadRDBp2/T/6esx7GjLbxExONIZWQBjJS8TTxk97
STtkaR+al63eycy5mm5UgBgJAJ1rYt6s0LKLmqg85UESSy7MvozY4Nro6I0bvI+va92FWv0LCoUF
bForDqxodz5vVP4Hn6eKO8pP0sX92bA4InkFZicgK407zz3fsjRyc6OJ6cVlCsBP0sQepKMacFTh
rwIEk7vlqcgxN77txsU3jlOYS9CzRXO2mqBP37F0pSiH3IEk3HgwMz6KvuBA4vyGXr2gfeKtClV2
bK17SGr3jcZJ7Lhtaicphrs0/B8pI3fqDyePFGfBdILoLqtyHA9r36Ouh9I8ojDKPv/ueDNVzhvZ
Swj4/a/3gTAFcKzZDeEix86VziahijUA4G0e6gpudGpgs+CuwPJSnbU8euYqGt86d5AkB3Gmt9hl
/Ix4SRJc/Knpy7KAPUnscgZ0yexgqBuzN7pk0Yykz8bDxpoTAqB9hc0qzdHlinrPh7Ora6nwwRp/
N4jvwjpt1teDNLZGJ4sHMsaN7K+zIFT2ZHuupM4qNaj0OLIdpt6TIs6YESyoMEycM4XQa8cF35cT
d9rwgpiKaLmVtDfwMIP2OHLD6lPqP9TJC5Sgrlb6Spsfhm1nIQc6nN1XVRCr/sht/vjImjGt5ghF
b5QAw7yZe4CYDsXwpkFlSTAVQhcQRP+HKXa6CsVbyEj7JqBLpolUfPhcEouveQbAkAtScrpZQMcu
RFYltGVlTolGdRBlLwaca8lR/dfoXpU6tUVVdtrhK/gl/2+ROXoXcusbfO1H5ufJ0euMLrJrCs8h
6KY9139PWAiksWggsedLPUqHSRaz/QudpBp4e+Z9cR6/R26BzvZYIFjgcR0bzXITc27Vdm990sF8
jaowOHILa33EDu0SHRamv70L7DnxEitmcTsJBbcW4o7q4bj+QvN//I0esU9OPvEwJ0O2f0KjH+Q5
RqDhGEqgMaJJMhMywy704HrxZtuswyLn/OmJOvoXP7cqwTY1fEhhRMNnmrOCEKbzLGJsVzyntD50
+ey9NwovIN/1yFiWByWzXjRGqDZ1ACbKKO/7sQQZZFmgM18JBuQqu74tUEfNSKaPWQL7x6N5PIPH
k+jsn7ZunWAJMM1wCh7HnZl1Cei3LdGlFxYfNzPgC5nfF4pavWj215nwICA7VbS4RG3vzz01KdZd
qMDilWYvjBqUgjBjXg3JbcdhzGT3IyrnXVihRahWh7GWDrWBt2yIvj0grJHFy3Jd3kaWHb4VHcYK
IRd91UMbSd5NgcBE4KjeTjbXz/5HkELyD6utqL82vMFH1IGLSMnXoPqaq6xSbwsLzKyhN+pRZ3Be
PBLJpU+k3rvfCdbkCNXqzGYlh8iAzABYdtsj4/eUIxxvgQ7lMQGDhawaXkPj9z4XjFkcxz+7tVfk
vAdTU2kZkFW4WGYBOTPZUeUKIhyrK8NqDefXh+0P/9JKS1rIz8JwOTwYRiebOh/RJ7pmhi2JL/Gh
pqTwlVA0ptR+D5XyGrucnq6Ft0Mwn73qnkgWZvhKldz51251gPf2fJ4V9la6j8Fje75TxoOlELM4
p56j32Q2PN1R0fEZROyCoFBqEt8bXShKvX3HmQ8VpRjFsO5C48XXBOWZkNsAIZ1LUAjiCFXeQ5lH
PgFxU72FCKceAAP9YUnNtlthjtGjohrcvX8izanm8xd1TBe8El/HTECnSfSSKghyCbm4kRiluGPy
UgQcli9escTf4G2ZNkTvbBtg+TGa3HwTWvnOrVPi1O8AAYMMYTdAoZ1CqdLdkGlwJNmGIJkbkjkg
EImiOuYogeU3jv4kXsNhRrmIGz0XrihadT6P4x6WGF1UpQetMZ9sVjXNVjzGcdfRp08/SWQdzH4n
IpI/gDwheBmyy72BcEJWIlUk3meP/jxraLDno2t9htEnXeILLtBCNj5SAtoPbnQB5W9h1qYIApQn
RGOCdPpQWTubx3+MTPpI1OZ7kerKcfek5Ua6LxYXYqLkZnlCHmqR+PxOh/yfgN1kmwy5vYYBiT1t
G3QUIH92v7muHB2vRNWUTbYFuCFvCm6qSEcRYUijH22pSd3fRYP97savrXOqRIMCsV/tBhuOrLLM
CUOcL/btbNPsns7/L/UFVO7E3rH7V2xldM2bpYIb3dh/xTORjh5TeR9iGwWSujvkDl3qq5Kig+XY
eaJPrGN3JbI8/R2fPN3Wb1xVDFx7zXtuWomEfPtIPd1gRGvDoXL9ysLIpVFN0/R+EIn/RdHWdr3z
Hc7hYNOThd2tsE1IaUaMOocaqNN4c8+ni5ok3GhURsh+w5oa9hV42zPQeE9xIuZ0jpRe7yhU/2F4
3642Suc56Y/Y4wPBUTYAEtO8YAaxi06UE+sGTkeVrbY8M7/uDnxGLS/WbgD7FW0+RVb3R0DglsaG
EQSNHRp0eJ2Tuoqamx7s4lqdpnSxVVEtyjR5lxkSsNFDpsQaHxZiLrQPUp92v2XbOq/BO8eEv+OX
Fq/SbNascp5GYBG6jBNWxWPlV0PO4RLsXMWgecEnkU6cPPasCq4hq6FumFcgnTmLcgCPjOhF3Tx3
1bKR0OVqbNVf4Df/v+pP0zfaPaqfLVuHNOvxR55jm0mFLA5/LV4IuxorOmkJhWQYOJ22q2SeKAcM
AD7AIncxvL8JUqyoJ8DIW+kDe38/LmjFYRJAB00DCCmubctJerTf+UjAdwha4pgdWDQdnJwgJRqB
4C3mysR6KknVT1clYBUOCEfUd5lEaJ1j+YgNlWM19WO/tr3wz3+q26qTxDuhwl5z04iw6FYFSFz3
dxeS9cF+cmYtngAazf93BPTnf/iRi6+zy1eFVBDVUNloQlCii0uJgQh672T8d6ChpxFj64PxHaV7
uKex4Is8LcKFyomv3IMrMiLLpj1Zj6ON1ipXQ3avrzVVaG47gCShm7urABlfS7L30YhAv4tt/56m
fPfRNL3YRkfmDbEhlBSvXSko4tUo2O8cdv+J5rMxrOe+EfWLKMPMaDJX/0KiNLqa9bWW8d1T5dJP
p9JEwugAEPwV0G9Z/IC5SnZSPYYWBrkv/xZTUtuq0cwz8jY2apX+XZD1kzSe8VZPRx+HO9a0TR6j
yzlEoMR6yweoYnxaE9vxJjoza03SifieaU1pTbH4QGY+IpUZi+mPBxSgCYb5t7Gjf76Wzxn+wPwn
JTbQGy4ZT8UVqm29w/Y8evc/kXWBLnQb30hUZPLChjxwMnk9ASh1Rc725rjyzFCQY0nr9dhXio2g
89ffbV3xXkSHarbIW+CQB4sRpBElFLRQAaVMDyM11JVs5NM0iP1Rn5cokf7A4tCMpxdsUshhouQq
oJCVq91OsAakCXs8V3bIsFn4pbr18lNfxx9OB5ynPtBa0Z9+Ui81quEqhq96oJaPe7wyw9BtIa4B
10KFxcZf80qdfbFZlnxaU387yeU+ols8zuj6S28uXpx8Vhu9b9kCM/+SjdUFp491lts9knQwT1Uu
Or1fYJb9mKju6j7lvu0uv0I2mPc0O+DEOsBAfUpRZ7QhMuGsrNnMh9lBW3/kNkmtXwFTvzXVsF5L
qaC4suIUuJv/clJonvK5LD/e8iXD8RSnUc8h9EWDMNUvpgj/wubr+K79oJu+iiy/wpFn9Bw9QaGh
LgfcizgIHz9U5tRYNqKwHNkNtKQXh8f7vfQTL2TkRcEmZFjKQKSfIdJMs98S5sAAmWGf2KjZ1CGZ
GI+OCKdS5Ucb2xBwiyyFKV6yyIABDJu5R5eQX/8nJ/zlJQIRBrYVGdP5shL0CQIbEz0umM0WlO+t
EPL28lni1wbto3GJU2k9MGcoG32J/VJj8rq6xEtYHD3FW+vP+hwVW3/Qk+N8MBspygkzKOfna8jW
LqF0stIQon/SwkNcAknt00iIe0gNRcWZCSWNqEsBbK4sRlzMk2bNSqOyyB1Jf0U2QIktuY4Gw9iR
zZT/+VCc/zblR38IWitWwymMzHYEB/3qzDBWyQatB+m5Q0vmV6rCpUjhSvhWyyCywxUcAYTZ2Kzd
qQ5f63PduP0F4Os5o95TPij7YnhJBgZ9srtoGPt8AkORptM9/Yhnvptu3wqpuqe48ji1Re10jz5G
/iOUyx+AoneoyXqq9et37F6uSZ7kNC3IPX+3jvcytemC4o+UTstGfXFRkO49vQmZpxGdfmqndmj6
u2Z5vMHNeuXa1txGINX/lSnXJHarhTlAhV0nBbyxPPrMk5T+O7N+GI5K8hvqtEgYD2BgamqkdNYs
bjki7UJWsqE48yA2/lCImtynNkKa0NDzVNTkwlNg4s2pxPOXEsJ5aLlFmTEhy8/nSggB9WBCKbEL
pngLGguR9jusbWQU1sZRcrrccWUE/rwxLVSunlUZMEhDxaDjNDm6OcHg74whe/zSKoZOa6theoLv
rtUcayvt1YQM+ezOuU2X480+WREXfqvLvs6QjBuGG3FOXreNrPgZjgRxerhtcRoo5Mx/OMgb1pqp
oZZai32rj8RoP0mRdnNyzALmB41JDdIBzQG4m1GJPmmdxnS2/p7nj1Ih4rbYdtt18OJpwyR1zZJV
UizzObiE2ibTXgQL58N+yTs/ddylG3B0SIN0C6SHrayAaagjVcv8GZLS/EcfFqUX6hFHMoXFEvH7
OuYzIQU9SMLb77o6DZ/QA8fc8c6023I7MGgyKWmJ/zQH1yPCnd4JPUkVxCVWeSomSAQpYsa5QybZ
SgdA7mUjjkW9C0J+Ek7u6SF2MTIrggkoboB+/8oyz5AdoQPkt1fcKcg+XVtLCP+gYC1gdCu9Wfju
wHe1XWigQ5HJGYlL9/WgWiM47buZQZqV3sov6h1Vl2kIu3g5P3/ySLbWvbWYe1xERKE+N0AFUDnY
j2cKoasuOZgqO+quEcNazOfb9bbh4dBQqg9AwFWhsEIUfI3H6y3AvXMeti/AUTSq9rciLQfLlDRg
KQnXAdHPBkcIlrjQLqLvu4dGbzDZjHpG6e8raXAO+0SUw86igwSY7GXl+y0TJPZDp96qDBoQEFwz
9fpAxu9It/mDvfGJKkGxF9yCfaFQzt1CBlUuUdCXBVY5recGbUveNTNKpJQwhE2CPW0AUeAesk2U
fbEy2/AHMtq6qg1nVJkiNcZEBPb9oG1B0CGGVUSqsaucIBVZVYC+Us39VWv30cAz2IPzLnMbFqxB
G956DfvD4o/TQEzMO3BSJGTphEA6WsMRde5guI5hGAJdCaA7lnfroVvYvbWgQUmBZtR08qC4iqpm
PAe3ziNLGafsseZXDNBM1JJ2kacbx5tFHrakkrimozH1ewVmtgJDWK+w0MTfHF64kTnr7KwfbSSM
IMLEqDHtQUa1ePcj/bJ+JZQnFgrvud3N/PHI0Ro3N8zP7XDcGzAO5zKgmDWH74hcTyhRPJHTObx8
i7JyfNLzEExexd8s4ShL0Tv5U66Gkm1V/EBoNbO0KEsYUj0aFp8lytBtQx8Cn9IgvGozADCqxZxt
exNdj7vKOfzVrSaaJRP0uMoeUj5APkZ0jA0XimtlTIEFaaVqa7kCG5c4Mid4k4YEyDJpYzCjGWR/
mh0hTOVdK6nxh5iGF7RHZB5poosiJpISBlb+51695BvZMrPi/iSzzWiDZ+Vtwt/M+sYG6L5ztmpZ
4WQSCEOBomrwyUzRli1dCQSCdTvEiap6iwTOR2NsIP2YZqXSCKxe8xa8IUEBhTO+HIUpinJNEqxr
cCrPcW3lrYMbPZomXOff8D13uJgKU6soNRYTS2U/jYaVtcmnqpEYqGVIL9JYWUJdZhqo1MSR/QOr
QWBWi/f/gEPwVQwM/8wO9bJYSEPJRYh8O2U/i/o6IcRa9XfjS8if29f3bGyHFX8tUwS3v/s35CBx
Wy/HGF3pdz2wOf4dd6mYClZRa2nQW2FjyGyHj/9RsEHwY+c3bMQG/pEIiYzPkNK68Qzu2tMcZ/gX
h2T66lgSTFMsJzrg1LRbw71YTfNpRsJVgBKZUmysZOB61pxxn4DX8+1fvOG2duw1AqmxicjZ2z3u
x6Zw5yngClB/9fx2zOqoyH691O545Lo6ZougOtKt5+e3bT1PKG73/85lKocSeEFfX8xrfQ9m/YbS
2OhX6EpiaMrxmUZEWh+5qIy2uTzddi5+DIBSJ30ArddGhnr77hMH26Do2Ue6SgATYnCS3IOjwbsn
cLLg2pbyzLrbCDN3iWRHmg4UCKLw+HefaXf3AgC0C7MrGiInzp31Dgw7KFvhSXh8WxQhHnwFGyoG
AUkeWNwAlZRjYTbAG8c8kz+cP71B0WKmM1QAgv+oBQ7vFgzm0XKDMuKPOGRTexl891y8Hf4Ztx9M
GwoCSRy1dwXfMCVX33NL4qHB8/AcchG+8yhMGhFBHuiEukI1VnUrXRk6VsdNl0yVw9xbZsyCEmZ/
V5bsLE86z9rl2I1WEoJ3AQPqQjLRYV9UUHJTzPZ+e1Kx6HZbBJuFZ+9hpDnpmiOaW5PNPJsc2Vtj
vznL4xAcCPDYtlSgs+Xax0KTxq9D/D0RNQHxB2XmYAatybs5hLT2wwxpT8IbCOSz71QVLUSVRT7T
ehBXNz9QGQkYDipG94PRUgpAwfzplceXA8sZSwkx8v3fC0El45j0pJNbWovODyZQYZY5+JHifqsk
uvrbxIaiCwCHHdH6Tq3QBGS+Tz9+R4ZIladV7G9kxJzTw+Cl4iGeotWhO0+RYdfztFMBbE4NiI2w
0+KfT0rHxAC/z7DeSNQ4eKh138jLP4hqVc4zuXNh7VZQz3bmLE8TRTVyLJCUNNxKa8jhil5aZscN
/qjXCI3Ole/zh0YQaDPlKvcy/Heok9gcG/+Z0VdOKwZmfLoOwcw8yP7AgmWgUa3V8PjxqXXIn0rJ
s1pFdHWBBjvYZSh7yviFKygMZXj0MFFwS7ceU3NeVKyMkdEVKy5iQR+3IpHyx5CBsxCZdTYXwVp4
QjvSkxnviOmA4oTkQuSuEd4IjjN3RwNp41BS+ox4twPgkTay1nYpRbjDFWa26b9rYZYI6vDNWnVO
yDBTwe23ZyGXKKl7+fbwXbAOvQg2JAkVGRxw84XnHoWhTYnG2RTvokxU1y8IiNBH2VQoIb2RmrB6
prpcNMKpZnZnpBJ5pnHxRgMlw8p0XRNyeONIndPfpZCs5d3/BegIAkzBHd0Gl3+c3JRxrKBKeXWp
rmTGL3Q8rTrDupK+A+2fsHQBUXePsk43Uc8dJUYjkkPZU+89BlHJpEoMfLz3S/MlzvIIRzPM6hNd
ctGdPrPA8+Ro3Y5Q0HLKPqxO+snF1lENCzo+1yyhb4MLtTiEQtjrCoFFeR+K/igK2VsaJrJsLYZA
QXpZhikFnIpIeLzel1Ukw0Walfdam3TtNmYyjF/VqUwaGs4nuGeh/d1QJWdIUEU6U10LparNx9vl
1Si+5fWywV0YEF534oLaNRSGEgLSalGzE6xS16cU/nvTciftiC42yMmAmUxmWhWkInOB9NKaw6fC
2wA/Z0+eM7g9x26oDo1jP4msbvWyBF6/iMeRI4ViN07yepSHnObxe07YkSPCmSOg8wBwjkQtBFmt
8Ukp2JR1rSGisRB8O4EDVgRnIh2S0o7b6iODZHDCOAfmw5xKUoTH4EjbT+rnjVV0IicbJs/ycw6c
OxjZ3oNRQaVJppKTXoI/pLGWWsbOV40rhvqIEpld064RG545ywYSunNTY6RmciXukPwEmeZLgG+N
jsykuTD1+RA8Qpu5B5UwbjoLt4gg9S0ZRtRf28g8yVxtakf2qMM8Q6CHFsoMTwZBEy19zDWazBSe
VL5MX8+uVfjfA0oQ7MKxNrOeo7hoTj2zkCHY4urcvDxUzAGbJoCmJGQfHt91PgpRxJxZ+I5WlU4s
eS19/ZcQUkjmXStkybF4zGgqv5C3L06tuck+IThK3xm6vOBPL13bdWzwq31U1N23KK2M4kSUrzYx
6pzfQ2ed+7wINIiATtNGI0i5EzLPeQnxryVPtBca2l7zwOUfVvvf1dewOEZAv3/eRnaXSQkftgVo
BmhTk6Zk3hd8xSZRdaNZjWAnCZHSzvYyVLHqb4b5wYIovOxKplkslbR/8FmCWBkzQv5VMuE34QDM
RrbvhNTJlB6Zd4qA7ssu7nc0l+h+CzY5Ot8ZlkQmftpI6nj+sVJU3pXqK9H9tK3sM2G2RVTeM/66
WyR/kAcJMysNYnXK6taVr9sKbx3QEkhPY+LqFM7rPnAy0D9yuo8MHkheK30CftbjUkcN6nJ0uQ4L
7rKosmq8GJsWjFVhCh6P61+mQ8tvJ3IeNlK7LBvBFyouAI2AsfH+Bxqyl4L56JEcAXF7eaybxcpa
SYhVp2Mu3XxJE2UNyuLElBiPiKs2u0Ka2Y89v7tsULtHTZcIQ8yOhVxAKLu+twMAKAb8E+Kcu3q0
h99N+bNu3A9fPMCbQPcCz/jjg8hvcQ7HT8E/BfOMoYz6f6X1ntliogw7UD8z+yDZb+Fc76QlViut
r7G107g0+7S3Gt4ykzt7ByqnL1W+13cZBU2wxfQ/rXP06JWub+j1Xea4awZBo26lAzD87MfeNN2l
eMd1NOnymXQRjH8aAOOwsHr6QdX2CUb8Sj2AEkeQaxubEqdp2GVoQf5JjwMzUgOy+jkizaWsOSDD
knmkdCFJj1Oxexy3CURuCdhhjLWEQRfIXPylF+RbFwnRKB3CXtqzY6GBmwF4DK+HXSDgSDmy1jR9
DO1zrU2DANTTSGl5khfVuD0WImk8ckm1dxEs/iTRyKBSTRB5EQ7K0Vxc+yiiTIe0QPwpAzwmAHNe
vPQiv7ldGPfitvFvz0SUaiKOnKbsnkXAW5+MMk3Y7Kn9Jg/nR8ASCiDUHFjtuoXcXds2TiCL4xtv
6J8V8LxLg+n9vILN+4jTwFJcnW8ZPzhFy0K4LGuG0yStOxq4R92QeoneX3DGKoArwbmxIn4pnU5S
BZqouQ62N+7I3NChOUdOzCKT+bVYQjgN8LYnvVMt6Po286G2i4wWdvFxFtfyaztRHp+66c40swkE
/GcJkdzoq+yHq2NvUopOyh1rN8JKza6a9T1nFqi6/tFEepJiNUPxZidy0PVoWaeOwMnPEJyVrck4
h+1Xnxq1Svcj1ip0pjc0ghCXc40oEgA8e+utpK1rDhOHBVeDSbpggB4jko1VTvS9UD40Lq/JKac0
fxiY3SmkyOFi8pnb4S/i2pwzJc8VgEv6Ws8GXDHXTMgEx7YcPkwRozRXtfDxmvvwMjjx09nAMhA9
3IQvLu38tM50Tef2tlp01mMm37s+Qm/TxMLs3m++bu/gnwzoX9F/2NcIhGMSSbM/WsuW6aWMnLM3
oV57au/EUDiW2TitQ7TO/vOyRmHYlLvuz/O02PTfmpxSUQ6hkE85Hd5eFFNm8/+SZTGMvyyvDo5D
2cfwIetQdkp9IoldD0yZZjIrDcT/zpmJ0vQ1z2BNhE4s/nbsRg8uUKPXvdUmHdtPz+08fET7TXdo
AipjG+qzyFqOSje+WSv24z2tfJx3w1l8ADnBCyAwygLxa3lbn0qii9kKytbvWqgBSY0MuaHFHkZL
/H5LLW76PsrY5qL8ufvwOK9z2JraU6gYQ8q66cTPx8u/XfPHh7tH7KLHay53Yd5gZecPhj6CyOV3
/t3XWNmnTF7ErTXe4bHDThfOQOGJ6wc0oS+hGtDdQLD6I2dmPuNr9w2RPgnaqGszW01OEbzhHVbO
XCAm8GCuf/PT4Wmi6/nl45RM12Kr+0bz3wSSvW6IxqIUv1hf0Vrl7Xt9MiIZjReHQsOnxP81azCS
AGbqViNzAphO52lWfeHqiyMzS79/v9s8YUa0EnxXw9c1Vd8QDkZR/MeMg+XA0nemOYyIqHIG1Mrl
P1QUdVHYmUoKB10AE+dR9KT81FJ0Md3FhIcqM2H1oSckFgUSSqVJ8F+npsR0MQmPFYT6DIN0yAAL
617XKiwxHiGDa7z26Tjs1nUpjvAPhmGy4FJ8U0AchabPGqWEXNAHq7dktgYindVvwAWgr8vjY9pG
yh0bVrVuJCdx7GK66dpwY4RDwiOQkMYt0lEsZDOsL6N0L9MwyAhjYapk8vy34zr+i0xOBDO2nv6Y
mjK/+rrCEGSEPpFIEjGLzWMfDcoUsFPcmTSThk4A9GJFKx4wcB2jbHZo+71t+FftZfauBUNNQrxv
BhO9+V0Et6+GM5mCDSFNOrw/Hh7u5wMQGBNLJXzO8+W0NqDC226Zaqy6L/1wN1PM7hVQy9B1bf16
jeRIHaiE/T7z31Mku8tRmtblagXCFr3qPQJySBAxEPbCirsu2U4xb7t/Z5+rEGTKD4O0ARRwOBRv
gegtXf0jf6RAwX1jI8cFf7KEmD8te4YEuvZ4mvn7l2qFDLukcsrM9W3pB/e0IFCyymXRa/8iH99B
v0pVXk4pTs4JHvk6jHF8OkAfTb9Ve9Fmm+mGNpRAT+qzOnUf2Ju2kBWMdXdTsnwA3mXS1KdmDhHp
s7cI7rnWQq5xEeAJWRT+M19Gqea1vIpTxY6gCSKr2jXGw3HJ1kNZLdDVi8+OHTETBPWLdbsC6zP5
XN1QyGS+gIMOPHS2+JhDjTsic1ksc/Mc66qbKIl6QEhA4psitAawg1TYhkpRWFwczacdGBxlbF1f
KoLLVUuUMSaczpo0Ovy07/KtIImnqW/qom37qnLeq1ynBrdKSSsbYY5hxCVjek1p934Ptld6lBta
815Pd3D+cN+NcP95297Do7gThJ9hW/GtS1qDLBKTzaRxdWJw5/wkTeKxcHV2YNjS9Xvu0GX0+f/D
4nAcyDa6P54Y+jEFpmgJvSs6bnPNKrpOVlD22kX3OeBwpODuy/hGAjor+eVSu/PR7gVVtWvsBD8y
5HdVY2aCs8rMcZJY9AzQqvxJzpmgDcU7LO3gjcCP3tKW0kRX3fJYDIS/qsH8BwV9oDiNxiV84LUz
Fgjfqx5SsbwDUR2PEShVS02BUEj02t+UIPLn5XeCsRdU6Xu2MQItPfrE6smWSXKOc7ekRvByR53M
luIMkhKSWdwJ/xfhS5Kzwkg118N6VG+bgQ7lH2Z7LL5yn7VDqRWPBAHdOo/FeuyQPIjmFpnZWMpT
95I6mQU78s6KHF4X4ImHVudfL0km9ISuP0/AGGKnzQP0f63eujlKG4LHP2b6eveP2Kkpt24TuI2F
KH3hesOrM/DyTQmieRLEBZdm+GEZaPqxgsKUuLtcIVkFHBjjauXBoKAgXp6q6/LwDo3vysTuAI8c
IR7+6K8luSmgbIcEnDcQwvd/7m+QZhzulKnwTgdTVrdDgE9DF5m4yhgvZp87HJerojCRJqYyMDFh
uxuPIneWcIPbcyRYC7DDwDyLXX/KQnmzMKslrF477cwfKUQCWzIOzb4CX+h9f8UPc7kXEgR5Kdcj
sd6he2mExwiXvtc4+hJt5sl2tx9g6Lx6vx5f3+AfDAgIYSdvgbVnr/ps2Ej76e0GmYZM41BcRNxr
ri/yRhw3NAVaZ6RXsC6beFvMjph5+5tr98UoKkcui0J97/ewCVdIL22xVUBPKfgBVfzmGqlCOoFw
3LX2VE9Q2s2u2ENHHPYdspt3hSTttvFtye9W0ieKteRJWn0cuoj+I8bW5bankZ2CnX7ILoK9N/tF
4NVXnv+WF0reNjTkNwPYjVik9aijJP/pq+S5ECR3mfV8fyjck5Uxv5G+x796ddxQjT9P/6tPzj7y
5ggOM+MijtNDyAzllFlSCIDVc/nshcz6E2IsvnNAx+Px2FHWvsZMI8kmVti6CBw5RF81ieeb5X6k
L/JSLoTJDZJMMHyrDmTkbNnODecI8Xsjm2tur//ClzzWkaS0PyLXzJykbM1DU72+rO1dN4yn0q6v
un6eI6xGHpQmfsoKqStS7GNsMJl0n8nZS6vdw55u7oGdtVVeW1RAZNRX42Kf0tLakgHZNPzCjxiV
yZSp3huv/c6XWe0B14c5JaKIdoFBH4N+hk+8cmVfcZ1vmI3d3k8cIT7RcidZO9Tic8Qy11WjJroO
OZ4tAjgywkR6pPq36+TGWVd93SAliMcGLb7RjevPr8NlMMx/X5cEO1tNz1xTEIoMFd6phyk3NWCi
EEFvFiJK/QHgoyc6ZzvUYlIr0koBQn9WXD4xtaISoV3dxfplh7Oz6yYSPZguLIgqU6eekeD/MzPA
vD/MU0oMoCIHJP7aODFCjdrfEl+x/4hgZ4gf7jVqJNVNgvHLpIldzzlg2Yvu0vZmneCUVOc3MxSM
s+U/suPpiqR3oxB/FEOTvxpOU06K9OWBmrpOao6KAWhfOF25jynRXPPbG85Mx9FeIpyah6RDd5Jm
OVEWTGoGUov5dTE2N6FSdYrk/1lQ7pMHJzuEdmrovubYqHxDaFw8O1M9cmAUMp9u+C0DOHAlT69b
hlyC/sjoAiNnwYap5QeMqsgd3/ckp9kFOseINNMcea0U6WEBG4ZPAmRbBqEwuLM6ITqkZcaaB8Sq
0iRtSA2L5mnu8KSZ7QqH/lE/g0KVzE8DkFMwyHVOIVOVXVqyL0yG3YAo6uY7X3rIB3gu4P0G9Om7
nXYVvq9/FcixQGYthokqY/OY0wJNT1r+6jor3iwKSzg2onENGGw1O9H2zh8w85Z27J9eKOlBaUJx
1tlWnYyIgbmHLSMVwIJWSgEQyQAoAgQj0e6g8MWbxe1w6rLpPbhcVCOCTN3y3oPHBxRxDzedolTu
JBcsaBt+nPcG/D67CSe4fq0gN21Z9mkD+k0Qqw32Z8vw3Wn+I06k8S8Zy3fsMkLSKP7sSSoG+MzK
T1c1ZHLmlVOgatEAQhtsJZ3mQJfuYuZeJM9IYWaETvCFtZgcrj10qJ2mVpfgbfk4FuqWnlhaajlL
HkGughtep+v/ogHQaG4oShzXiqP798S+ZaoHajgtwvWeNeFkH2Fh0P+PU+8CbbdqqDitClmG93Zu
qaMrheyP17lgL5QuW4O4/ZLxP1xnbSERa8L5BhABaIIvWBhxEBQzBKsCz6nMAvtqQXT/gCsAu3DU
w2cCLNK0jT10jzepClU03baSnNjslzJf4SHdMbAplPr71Fz97/Ku7j51bmCItxvJuOFhQidYB+ep
qqjwwoTZmHJcY3pYYKUccvg/jtJlbPk10u5y+X7Qm4+z6vmKGqUGnHrRf71jFnPzezA1aLCX2Pf2
Kx1hrjoCW3wZ16IfxLPcCw0DwOqnlTL10RlxSj64OevrDTTVs0Rbb10TGl7znzeK3Y+1DT+luIcR
buCNjFSRUD9pm1vAPDYTxkNe3Epgod0awlj7tHd0D5WhI/7Dtmqbo+IMzG4mMELSX3eh6tHnU24Q
tjKqQbHGT2/mkYHvly5v+NJftpuQdbyBmzmgcjTYetilz6mSv21xr7uP/vM6aO2XlyL+aCUo5RKT
Q/ufVAS5EZG9zKAbv5Rp86ihYVZxEhDX2JPiGnV0jKpCeIp4keyAPu+lbc4N/dnUIdkzGEHV3PBF
dUSd+FTtrIemGoYKIFBd95ntIMGsnrU15OZnw/D3TtbZr/IqdK3hXGGuGlXv3Ahfs5bskNhtBFCR
Q0NznG1hihQ62h4gGOD8xiAkilbKi5dWXMKFtSVc2GJKBXL6G6r2c3p5ItSA8zncAVpsvHswW/kr
usQNEVdsai0gnq/jNwxxI6GoS6XKdqqSfW/+v2reXMpH+sYgV47Os/oYrUfmd3d0QBYBWmlpjRir
QxhXYj+tHpfupnQ7uHjBT0P/zGXHDx7gF+SOem0HATxngWNJLgE799Xq6N9jlNq1hcEOUJmATcyi
cl41xCjDQsIaSm8XagGQUI5nOhjopQIq9ycKNk4+kWUHjgQ76cXi2/V/02gDKam2qF6g1t8re0r1
cN751/dDXkO2NFKyxHxLQeWUbKgkBZchyF/Pm2m0Fzfr8v8gi4iOKXPYIcXfWXaVE+rlZrs+n3hv
qgb9PBLKpSxujoTXJ9KYF5LL5+z5JKkZqmAGpbOi8t10FehG66iqpqK1hSFI1574PzT8vZ+hUrf1
OfdVHnvoMSXnBLAfVJd7pH7pa0XDepghSoXQBfR319W4ZBl+d3/EYLA+FpzAvuc46Pt/CdMsRzKh
dXkpsjNX8iTkt4sIoX1/9bNQf3DlBjMghag6SZvzlFmF10JCuuagy4oBbnx/odJFhh9S09oHZCct
/gIJJPi7h5DgStkbB1kakM+bD4nZh1IxPwlMZ4hgCoO4RYw1ITmeHkxJFHjAasJjap17jZgD8tqH
2RQJ4MEdtqxT5vqdVSGqh6GPZhsfYMm2hTLo1sAkTCOYchOrXo13bZZjKVK6t6TYgWkDGZQhKnuK
4v3g8IkjpNqfO7fP6kZo+B9VM5KgzRdUp4RcehQWeCJrUzQy9nOdX4A9KPXUhTO1VcYnVXp29PYu
qOCzLRssvJQBPxyT0rtrYH/OEDWcLmE7D0rXGoNCeiRLxG+QPHDUQR7Be+DYH0+gnNiMjPRDaYDA
wLA5LpmHdhQBTM17jeAALYxo8JReRcOwoH/9GzKTYbvgeVCy1o2ovsklZNlf+/t4mRGpnT/WAKrS
Kc06i6pCzxgqlwz91Gf42qfiuY97JKRzlFUyc3vnkNp+J/VpCxm2OelX8dqbz/xyWGho9nh+N4bG
REA5pOpjmnb3dT8S1nuLILzrun7B6DZud18qHo3z0JqwKQ7fHFZxzgw1DuX5yn7jvxgmd8JKyqbV
1vr6auXRcH9mMmsFq86z0FHbX6hZHT5hQc36DBCgJm2qsjpuiwo69ep+T8XAprgByDwLB9AisUTp
OtoHWR6J8aGh/ioUNz8G62chszTsTEBSQCELaSKI1N2AujUvAKSpsVDReNKEg0sCqfp2V3uU2CXm
sDvfYSqEPRoChF1mV8nZXN0lEXJ/t1pew8Pizv0YBhEgnUxkIkgl4zcU6Kb+rXtO+GBTbUa5iO0I
zgRC0++byG7zs3XnVtVSh3EM5Egnu7u5Z3uW96aY5Qy/PecKxpUxjXVrHptbhQXO6k5YUNGX/2lD
WPWbFfKEiQ0BgSuEBV/aOTKMI8Tq1WrLB8p51rXGxzdpFYay6jkoHcF0WmI4huzzIjuM2y1TO6cX
KFDLGwAaKBLpN4ZFbtMQjA7DieuPduTXnsAr9Se4F1UwW9U16WJ23mEgmPZIX/YqBwA83iJAPjmb
lhO7FhkaWpBopcpFN7rIxqw3ahW+EY4VAIRqw8r8QoQH47tBmKZhV/QQoZiEDUY4Rw1iikLoHAmT
bQG0EO3OxiBnMvt7PZnDQf+qXZGhwqd3xNrwsTcO4MGsPCYffw8X/T0EBI+TlGqGEOUoYKDfDmWH
urZDwlWGdfxy2iSeKy2YM+4v79IeQc3xsZCbO3hE2AMqSm+3QTIbx1haHTR/I8UoruCyclxSTl3L
aF/Aechvyg60Kaz7SYRb4WO3G82E/NZmXh30pmyXZIFj042byR+gx3EImnQEAgECgDdX7pIE0xas
VLrFSkmw2vhLuLqKbK7+Hi8CNdx//KWmBCJKyQ7YvwQZundDodvRAsk32CJkMxQdjzMHKQ33QitI
WfhNwf3f0KoSEnX6UKrgC+8P6vhrM5Ol4eWOog2sZJwoeleh8Vp8YheVTIK0Xrm0+G0ImDguLe5z
yBll8jo8Cej40cg2dZMYb+hlA0tzCGgABYwcdsPQlugbGJmFaOZ/Rm9ASV5CAnKl/v2CeKzz75Zk
MYb6qpgZeeJAGdQl/pblAEHPgFV6hF+ZpM98oPN+kQU1Q5bsi7vQ0AlgXoqnkFWRMsdfMEWMSrQg
rXUY8zFhBZ/+obOcSjEc6eqbmycpO4X/NVIWdjhf9fkV0lUdoqoPH8OJIjGF/xvhnedvDaV9fj4t
watgWWBrP5lgd4fUN7c9IS/P71CGyQy+phlWCV3YFOKDHVDTrr1d8XBTy5Xez/0Z3R3CteQ/2/a0
d3BMP4L5w1wo6fRAOJdz67DGyAE6vcRNpRUtmiUFpadT4maRRK0Azr9nuhzgz9K1G6Vu8ucRnnpF
19Xb5vuD0r2WTb1EPgoWxDGiwvt/umDkFgeiekqLPLiUgIJ5eHrf1QEJA7+fS32h0JKL2t0MCNLa
Tsgrrq4PzqoNBwGdQU2NIlmDyPE8NKW3tV0GIazFJcS3eKSGjyWAW2E6/G9M2NFFh2chb90OxuVF
rPwTPomajoF4K59u4UGWNgM6CV/N0Hcp0sEPD6E9PYMU9YiBX+rX3ryNz2q6VgbGr+Mr6BGVNXce
oD4wF7tL0SgoK+WG02BWNA6Q37YVHy7Cu24hkbTg68IOMmZBMhstlNDmADcJZNuse6msvB+5AlMl
8AX9HKsj31H2dkC7jKJBD88Yd+xqTJfJI6+LbiNM+QNtCFU17vzHurqz0Un34o/F7PjJckzRpYPy
Oq/TG4FlpzAHW+JYIp88P7pAqBEgROWX3xay9bTcFX4i3F0w8XWXRwPo+7E7W5AaDbDbZl5B9nYm
jN7mGijQAYwVdQVHOeWQqosA/uoSl7sj3RzGv2X/aGhKWiP1SLrpmXGWpH2JLCPzPbiGucTVoIx5
HoxV23n9q55vCRa38ZeVGn94jPgnyf56xAfGHwMmLHO+ILgt9uIfRhwksk+zLrjjllvsDzn7aTAo
pumV/pdeHhLfqt/K3rjuO8kA7il7dWl28kd5gIGbCartPqDm4EHJNIznk/sZaHKdEiLLqIviXcqo
X7ZRxJ0qovD0Y9LzcZjvf6cByK1CgLFF7D3EBuWFkQhcIP1PSkfCtwMVf5SlOCIlGLXmakwcpSBj
IWxWniUphYpkGbvxBw91dkRfpXbd/MN5tRGSERKomE7iiDDGA53HeSLGm5lqtXXG86OVJmTGcxl4
Occk6h8nogMgsBs3J9G4FsZE1jMy83bwCe6aG45HMNgvAUMePuLkm4nAdhTBq6gM31MJWGkj/U7z
mM9SLvM824zzOajn06S2VVdRI/d4HYsJbGUWPlP8KkwEgIwq6m5SRdDIytN/m3dlmWIWJ+fnLJ5a
NIyru2jXRpgVW9YyVq1owTJvmmH34kC4PJCFPYi3yR0FO+HiHPz9hcGnwsCYfQjBGMyEVELZnCCj
7Eh6fJxD2AWsMZfQ6sZQXGM+hNykdALkNKNyYBXr+jP1Rszg1e8DpkBxdd/4cSlurONd02YtVP8v
nB5R5zo6oSHsAFogUsWRw8pfA53xkn+J5JvS5egoNqVBjUIxiI2J0kDblL4/QUfxNlpR8BRNOPBC
ez36128f+gmPGUeyb8frHqMGEgGaxafQ9TpT9IRtbk3MlSEw1yTAjTc6nyuB0iW/1mZ88d5uBJoC
+dye5uhNRgHhmAhHk17mr2HhrJOzqGDQvO65WHXXD3VSp746qk1jk39UwXWXB4NRJeF+pC6LlcsX
XddJ6lWqr3JsToJJriAKZuIqVtvFJ329FAo1vfwMePXQITK/HJROwRjeVN1RYKTOKRzil3l9pM8m
2FR5zC78NzbSxxQt42Q5lRzzw9VVIXYk2Yy8oXSCssJSJVcONujQbWCHh4DuWqsUCCuVewbnQIai
XJ5L5sEHwlmXDyiMN3R3zWahPJxAektr2J9UBQdI8TAFbQFSRQFf4TonLvo0bpPTH8z7Yxzv/v2s
uoVwjNTCz15lgi1Bp0bubxc0i3v3D2i921deGHUM4dYCDxCNbAf/L5uI0+s3CKfYKYGyrNWtZnya
5o1wa/44GEhk1ifj2HaN+83Erq/MU610f7oVpaIQH+rkxcPBTfAhKnpUHLbZMv2Cx/lK6ibcrad1
W/JZD7LwT/TYn3WJ4ybfCLTCgUwVDLmKOZnxdJC7eYvn9N+/+XeZYVWO2jx47/qTXLSL1YqskXpd
2J6o5bijoAtOc/7eCB3UGUzsSKqkQTv5eY1US+JtFGnhRZn27YbWTXPVc9hDg5V/afl+bu+cyRi5
SPxGNsITDMZwLHzdF69puPiuDcIPBqvU5zX2ludj/bWetx2b4GFJxf/3rUcqWl2pI7wdaXAigAOb
IUH8u1aqQ6GN5p26oJB4wtrDLho5zQSbO5DBs7Vu6QHuM6NA/QpvUayjrvgUhj4MBROYvHXjO9f8
hwCsGhmTr0a6OkrtfqpoXOnB8yk+9UgNJBT+XDUlgGUUcz6iIxm9fkq6MpHkZ2Eg1wIspJhAfC4J
/xdQZPdIh+KsPJecANXK6P3klVk+a9Gjs7ZzvmhpwpaivUEcYUr3644NL8ZRV+uvRo7XeHsTc33X
fy8phznUXFp2Qjm3JwtgG+37rI05sP/IoWr4VnZDAznnG5q6vnWilr8OcMqu0C2HSPxvUpWDf434
miArl8sFs31ce+umDazmfD0gOQrRNeELkKQO4vrnD4dMQIWKYqrMQjq8A1/Clx7L/hRA0D+uzt7c
U9XPCGI5dHIN+PwJm+oxRkX/ekq/dWHqD6L1gQKB4OBuLlj7FmWb1e1X7LROkXb6Y8cevMRoBqKI
Fac7t3SV2ysUZ0Uze229dsmkwQLvLGnPv8HJwpKG6+VMJK7tK6SZOyE7cWXGDdwZqw/74eNQ9kWP
sl0OfHm9H2sQdpDbviQTGidhiKUFC2PeD+LFMMykrcLFdHPfaeCepNEI4Nme/5Tx8uDXHbC0YIXT
mwAiQC7BkNIl13YUxWZOPnQyCTU2blNQ3rFgD6KdjXQMROUSDN7KrEH8b1TyuUvYR0RH3BRugB6i
K3g429cmebXR/yMk5FF+QVtxxoJGdqGBQWTXiJB3KEWjN5MggMLHWUlqGfa5MC5uIXVrhb2nms+H
WEDM/Jb06wwnsrw/J6A/Qvf7gKmfmpHMRpt6VPgtRytbnRoeVfBwssgJAVnIp0eaUjUymldAgOZq
FVaFWWwUGWIuEky509vFJw5Hv/TUsEYegNTbxPAp6W8a1mzse2Sf22PvNTUHQZ2/fo6fXXhZZshz
2FCIItk/b4iMWoWv4WQ8tIRL+N5mbBggtUlgdatNHxk0h/p2aD9YJDi+0d4lZuKH3rdeiv6mqOp7
NNdOV57dNw4L+iAzutmYEpUJnhkB2eSSJjKzdN1TCpH0mh/RqztEttWC4PD3VHbdxKv15q/MPPY0
lN0Tvbi9KKobeHqgrTJui/DFMyV/8m0rOuPzMl7d1Qq4szMCzTY7/Y1LDJoDt1VZbwmCEbQBk3+T
StglDI+xF0xoKAdhKKYufXZS84ihhqnczVz3glrai1k7Y3c2gWP7Lu7cOw1EXERQRPa86FEH635r
QfO+sJgeGupBsJzv+kwOAO/SwDF8jv48f9AbzKvqKqqJNFoyFb1t2JnoZZV7Q21rM39igmRa+4mq
1nzcn2bg3k0wOIJ+gGE6RkoI22SjPsD/nm1CMdupZcs5ZKpdBe+8MWgun5MLHKJ+kJQPy9JKCPOq
cHsWCClhW0eUrqyTSvTiEIh/1yQ82WWy4sIxfxHSpapE/ucWLovfFvUpdRvzka+fMMnkHVcDBkfg
ZyZeNdsGJqhfTbRV6Je0/lVvE+lklBzQuMz87/V9x3EIRvHHJvxuBesINtt37k75eBbEVijCZFFy
84MCfM7Rj+G2xahMVIbGwftFJcpptCInuft1hWeNZttxeptgUc1rtEQNgb0jRjDrydU4NTXEYzCH
6Kfg6jovjCZTDw1hVZRGGOso7RidEGwdl6/20P079zJ9ff6H313NOelgZEsXhEeVkwLSdqR+9fWl
aAtIuBNjJ9j1g8ND+lJrpxm3U9+qw1E6jndOXbbA9TH+ZWx4pqCdiFFLhwKjCciOhuLHWpBhFUaX
ZmL4ns9OoqPb0/aNnLW2iZXOmSHRADUt61+IA2P2GAoEK6IFPunGKlyXvNekBkC4OhVtI5xJkNq1
Uwo3mmTGxbmRD6XsGJF3t3AZpFn5qAMomTPgAPrQlYK6IMMLZU8SwgGyqWuJqBn2ZzJ+wbAwn0JY
JiVYaU4RQMm+RwYLsTd5oOsigwEBnCqkNmos7VDOKUcobBwtHFDBqAkvE4rR43fiZZ/cxagKkYqk
+KNY/FyBZwaS7B3AmbZnZZFDRQoT5dhVMIP3Dq7LsqTtk/fBJWUkudFiZEtSFknjDP2hkrLi6MJi
TgyTBE9YXHiWOvL/7fnmwM6deD/2pzpZ/k6K2wkq+Tdp3QfWwEJaQXG90IfnaPiy6/xCMv+9CK2M
wGt67NpZt+KQBqFTz4lk3jS2znFSle7gw2Uvm7tmrAFv/ETqTW6wETOiIgshxAmp1YR+hrb5H379
HQuVOk2fiOBnlZ7mcpvKpnyI4xLywsGNll7iAKJLv7b06aF0ZactgUcqmDbF1o8f7wdiLrORLia6
IzDI3c9RDlCluc+DuTF3rXOHKDa1ZyeeX+Sq8f89HBYstRwDetMJ3va4nK3rtNESuiE6qkaRwzM6
sIc7BTdVkY4Q7VqQMdVYYtB8dL/mlAV9pcIknIn3NMYO16HX/9gldlObRDVEU0Ex1hRSdAh2G6EW
ei5VMRZc9onVQi8FeqTODwppbEI9a4QuwBZiFFHYJpF3XJ8UtSJO6fjdboywDr2sQLVieEF8qvxu
ywEKzJjvhxSDMFjSjsXJIvB7nD6lrmLnlNYDEDUThMme0rgHGKLEtR0NFPRn7FJyIyg/mqKhF2Kw
B9nz/OjGZ37A8syIqEtuASMKUNEg8LIrRB6kIYAGwPEpKFH44U6kTpJEagehJA72TGCFKLWrpsHg
aLOHyshADijBqkU3PqjQlLoOLvHyXW2T89obDEaaLmeL6BvhDOH+B87YK1qq0ezSzfh9M3sNKjDU
7cXUJaC14/099SKvHBqj1poiNcVUyIiz9zBPqPUHZ5n33CI7oxBMFUiNWU16qThd/ldJjsDGHNNd
YWoA3mDsWvWC+4+PGn8qUHEBwlob7E/rpAdypTccTfTnRRctOiyJIDRFLgRILr3HHYdhiKtSc20L
krbxqUFpu8MWCJ2sIyOfETypGbU7C/mi0hweym5yUJJvezUlD52il/k6U5Gjc9RABSdA4aTY+Zoy
rc11JALfHoTsmaocZO+7arYn41W2Kj/iInCoUZP2ib8QegN3diK0dmg+A2ADjK2oRfML39h2wZ3k
flKRznmciRLf0UKc6AKFIvIA12TbGDAFvO6TIFLVdU+KEz2TqIIODzhuvlB57CERuqYiYJyLBdTQ
o/NqQRfk1DFLtB1YYgNcoH5rxkQhabbS9iOuXc/HjkllZ53GWOJj3YgV6KaQWECOMZGodClIJ/4N
vuA3zuAQe/ctenwV2x3+XnIhJyjQ/K/3DuNljb8dPBERrHz9BI4egkOZXlr6UitOIQ2QpYQ2LSsJ
WGsyLkL5LvMRoEdu6oDoCpKdQtmCqq/IHPqzIsWctog2jqwOtaTvXKYRTaX1rp3Z4z3B2Ioy2QBY
+NpLqoTDCKKWm72S87GamJt8qX7HR5iS0enZNXwtNzxh21Hy61a8cBfxjPwcxnjr8g2tSZ01lPvm
sdGb1ihs7y88sPaIflCvUAZZe9D5d6w3tWz79+NvR/QXVJeDk91r1qeJQz+BMT81AKrNLmpbJDvN
183iHTVAZapr4/Bn36M+Xv4JXA0LhTh/zGSTKj/8hPvIqCrH8R4XExcROdnx7Ug9Q9xZhTdOH1zy
iPGhFkfbQlGNryagzGk/Q6qmKC4yF29ePiG5yQcJHRr/gGE9uSMFilLm9RDHvYrmCYowIB8//8TF
WuKqSDg0ql6OohwJBfbkRbCADpmdaAU0cUhmhoXscHg93Yi5GK+xJA7oVXAixTZD0nhmuEJywePv
friSmStayZXL7CjCKLlLhawwClqRVSsK/ubdPWybBoaE3IoiqsX+lpxpAtUVjZ+CdGUFQJuqTiX1
tkJZBqmKeKDhGDhuzrSPrk3ZZatjcbyztIhzrIfz1Gon1g61O4gSwVdKKiIzRvSUZQAvJS3pvKWG
JLj7U8xW9zZsqXb8JIRlvdbNrtPfs4HvyAg94aco6Fgb2GIxW+jASnZWTVQ20YO60T0I7ppgItsN
8W5BL6Ns+LnSuTXCs/ntH4+vCYZ/3Q0+3N1pLVtqzsD7IJEWwpdDCRKRSf+4qHjUNt/BMZ6DW5My
nTvnjXymbX8m31irTLeqk8W4NZPEjn1XVG0+OtGs6KmHlaPmw7BtzGcwTkAf3YLktwhtMI+ePNzU
8XOohD+vslCSQIC4gF9ktBRn/Jj9cexs34tsQNXkxBHe4aEYT21DBvXDzWtGEdcWwI2Y9zjsLmyI
ex+ja/yyMmxwTt203OklQ9gewKHK2/vKFFANo7AItmrevh5VYuScdRnF2TMX6ZIUhHvBhi7APo1y
wSDWlQsTdtxuQRGeNPbWc4oBWAEfl9jIp59nojdFNoMhKzZy0PfCs10zvIyJVskoajqdkgcpvbOu
WHdooM6Z6bXlbPw6flDE5E9W9Ro8Ztw/o1ykweRja6/LsTCcAJigxTRLHWi+nEwIt6WWzYuku5yP
ZNbMmm4oOrykGSKe4aK7MFLqGoOpoxbZnEeSHe4PrJwESOy5gOelIgRHx04Db+9FAOjZVN8J6iLN
y6RC5cHuy7BJhUmDeF9z3wgwECenWlVPlrfUDxHPP6tCP4RVu1PLPIeouOQJAS23T+zkoPNDUTD5
uFX7fDOsJ5z+eixzHq1aw4FbhSaSSv+dV+5VAnibklC0ANCB4C5TeWZ112FhTF+CdtLofPTDsxKp
LIU13QzvjFghfTpoI0a3nxEwD5Cs0XN0rMj/6NsT38Dw2ee8L41L+lycbPPDr9qVIPrUll33MAHd
CyXs3vdseIqTT7TMNbVoH6nBqOLNszo3n9tGrjzhJRunFH2kNOL5lSdlqavH6hZ6RymBbo9o3qJv
W9FIq2m2BAnBZ88Zd9AL/YoxSMUGHHOC1MsdrmU9aDtbO1aulOU8hyKtJYMml/S10dY52fyHoCdI
pblQPw9YQLISoHVGCXjRdXXYBd6SiHFofSmZar93o8MV8/kEW0DYLCiazYhjjy3qb6XYm2tnX2OT
tuy0rFB0SUSLFsA3f3zHXpjKYU8UE9izkHusnOWVnAiLlv1b0N2nxH1cHUOiO3HbSrs61IDtOZp3
f0CNBNz97ebcD/2EKwVRXKSxSw3qd6Mac0z8hzy0xzmKbqp+8PEvwFnRiloOJ8AvDYi8/xPKEJxJ
Pe/rSd6bwHJ2NspZvNwKzC9zpTUxjp5cficNXCboRGRJjQ1Hm1IQ+N0pfH8Ad9iesmfKUIWzYt90
U5yDCwsFPPRl6hKtrijK39it/UD2k4ILUxi8fq2BEu+WeLQQHhXVQmLFKvsqJphbZrZMnrHH61f7
VA1unrf1buXEDr/I7YQcCkgIPej461IQrkwTxWtMWqQO2fdl9jYy+xi2R1BAmORmkUGozMVFL4TK
NZNvLBgk/AiL5YP6k1MzhOp0KdC/e6kg2CvkUfR/CaxgdUZbUswJxvX/NJSeJB0D3ir/t9aRzMH0
cGH8876gmIiOrqktR/wpl8YRUmeuf9cThtJG7cPFh2qs/UldZwfWTH1hjOcsgo4QcIeHUJbn3AvS
rbiBK4MtHqhgdE7oO3ArWU7iXxKW9YcziVWG8FivqxdZaG8kxvIXPkTrAJlPkjGCl0DUZrbLo8dZ
UXLNi6dTXO0T5O2lepHdVC0XxbzxBltKRGYLEVyeGYzxUeXhfAs3gMtGZ6mSLRyjauSaB81n+hxG
ZGitrn7Vi2Yzdg11Hpq/H7iIJca6MGANZ6lwJfRQpEF+rNb6fFs2OG6Vr6uJMLVchiZgAiefiloE
twE8n+Gy1edNH5USntxlAgR6VOafC/WitDWtt4bsM05c3U6464LkY3c6AhM4V2yN9vRCA6ovr6j4
+fL4Z3FCBw48wxgAyhrXKfe3lE7N3ziZReaoTMLQwo5BnTYwgWM0vqZsmAQ9gDOFjtWLCQWLN/WK
ziUSPE1ji6Qx2p7s4YV8KaMJ9P9h6IqJcXxjmIpF5DX93LOcPozopTDUt9/JSm1ERFE4rQe2TsYP
YxcMUNHwd07GY8aM2RvOR7mzZtEsM33nO/zE2kYWTD73pvIaVvKSlNbr9hpIa93ynv74VDZ6uWZb
NelpaiUtf7cqrZRx0gwj/YV81ZjpHMVGD7UxDKhbsbuLjzWJQwbdwxyZP/bBBF+yMIYjn4+WHUGB
LO/lNWlXo3cJFhLOElQEXwdVY00hYObdej9gO/FO//duyUfkqeZ8Pama0uGRR8SGRpoXe38dLR07
4xHBnZjWzym/r6b8g9ZkVnrQFYKkbprh7n+4ldmriTAgAD2hCue9loNsXNqHZh/ubcp2p0QrTkwE
Rd5OX+wOoqyOCk12sgyL50agkGYKtkKC4lHwHbaY5+X/p6kQt3e6eRVk0+y/mbrQZCFh3l4CV+Qe
tmfe9temhzXf1xiMjGSAa4KoeGqzs7/tJJZhHYtCYrkqi+afyr7LrUn9LZtkJ9eSJnUY85uAKL4z
p0bFKONwbkKgocFXBk4zzaOhufeNjXGTjS2TM5PbWExLqZ4BQbSv73H8bxcDc3DOb9o8jABbPGh/
OnZaMEjhNC9zlVjZ43kOqOHdS7lNQGwa9mLYe1Fgpg6wnJL0W8AqY1ylbggS6DYgH5Jp4dliVCaI
f/mdkkjNIfcrL/rd8xSjMgudS/aw8uuCNTCQCa2aoTrjHo376G6jqeDxCN+IBMOAzkANgnzh/dLd
T9M1YWJEZ8A9bLsUM3raBkrKwTI0EEPigSads/c9UWaPhDs5LyoOoyx1N201E7Ww7tb8+D2oodLU
fieRRXvIgVB3zB+bB+5cUDlb+MgZi/Q38V8sKrLF+cmS62Z/hr+dUDfkN/VD3pdiwVfEvGfNG5+O
qjsEosfaBp/ytiOxbjkiYmwGfe8VQ4v4sq/exenuhqojPzkLJk02ATOLcvJGsMK1t7PprQsuxx9O
lUPpqkdhz5ZIFVCXLu1b9eAXLT+R/VyHta9q389asZYCXi5lNT34cx9YUwAdNq3Yv5/tNiJrmop+
pidL0D6X1jKPA8JaEylQXsDUtvyMUmEw2IXlr1VkHqNxUfD4yG1v+JLqhspf5Jz0fld5or2zsJz/
VHbfUbyNPoBmegD5pYVqd7iszgHe1TPZQ4KOuiLJP3gQ27Q6wlpIZrJPJ7QKCMHqOlOXewbr4mBH
yPvpVtZO10p8wMrhxBjYnCWEypYx2zKZyjGX59pWUSVAcnn04QTey0jSIkXWAGi6Wg6QpMZD+Vyc
jjeyseGeuhsftdxSv50qKuL2uRNwrCP9CDkbqSXPP+ATioZPC/b6+WQHfohpo0Cez5217fmx92Bh
ti30yle8fy/EUbilN3A2meMJ4bMVHRZabpqa7e395TAjWUJpCELWhN+1+1z3pbPIwRSWEEBO6DeA
J9bzlSaFSDBoKv5YFnUGhAE+xdZ8aDC2QIn1vOHKE2x6YYiuY0WIvQqb2lN8+th63qB0RHiknQj/
BTnzMZPy5hB5AOfTI4vgj6Oh9ee6p06MB7DAtRz8ikYQXTAGz/EC3XOqTSwu9sDIE4xngyglXNR1
bh0H+D+9gwggK9brXUXe7vpGRPvvKW+91NondtxCbKHLPVvBxPB9RtuhYWBYR5ZXlVBcc1NIBOD/
02jU334I/jaysjwKb79mMVmYEHToAQJx6Qz6ITS4UsfWNV2VDIkvg8B0E8M8Za0ZWCYXvvwLhcHW
T2Gnywg0sLcnbvGYAxR2Z/wk1bgWtfrFF5DtR0FFTGcbnzlgGPRZEThn8LbKE/ClAuGMN5bnbB89
Rd45UnWJ3GZh+jlfAPjXytbuPwf1bHN4eP5UIhRcKMWOucXoP3vnLr/eZKlS2AFHxjUBLZYxKzea
GsmI1Zo5UYMXffAovUfjzwNYowqrbjtaVnZYK1NXVjqp30gI53IWYaWeKNRd6j0aWsQNiDVWPn4Z
cVAECdzZ4v/LKdD9re5yw/m5guGGyXxsCH+d5a9TtPOtrRyJUORdNBSV5PjQp11tWX/lYJSIBRJ8
6mHgAI4F9g7f9x+aVNEgZRqkMXTdPe+NYpPXS0emsai7MnsvfP0S2HTw/g1ZzoQglwBd1dj0VJQZ
HdXlaB5zNmEdwQTDvNkZ5AOkh1Pqu42QB1wt+BEM0EBPff6qVOKOGVcB++GTCe7I09zgLm15zFQ9
m3iUfQ7Lqo8MQbJ5woY8F0p5CpZNxCOQIAz48tdFAc0wZ9o87D53wQ/p19faPvKqK6eyy74FiV79
XsW1/R0RvyBd3ij0eaRpW9aBI/DjGWPxpJF3t9LVq6CZx5a0FvLNNL1WWeE2xHbBfLQ0kYkwy3r5
ancZF6MKVjWOYh5A4ii0XciNk4RqqIsfUdS2CnZIxkBGAYeHFSQdNDdHNFJ1SO/NdOzqUEtgAAWS
/MNcNEJ+Cj8cbmKGfyl7JevNMdKIBrATA/8pdbszv1lvC5o+H9Axkx80lf70YJdx3S75p9hMGOU1
VjdANSWBD9H3jTJF1V/W6ytWAr+9KaDfjQofpki0LsSbmfeFxCeUqq6Z7/NBXT9j84DkLpqHucJb
TFAt5ZYMo7isnqC21XbsjREWiRgajkKfrr8vPKvQdpmzrpWKyzW+cnpYBREvVoLSbRa3PG4CM9YZ
75Jy2WaSODMiF91DIGvzFtw315OrG0XjOrw1yOFT0gizE/YXgYrIjChYan+c6bQ/ZeL3mOJNEaUj
fHwpuDd7UiG04y1vXXpCwcjYBpMMscsCehNzeXawvtEXDoZSv3kiZiMic2WuxDLcbK+5ewm/Rhd3
buM0QHWINiN42M/0Hs28mFb8Hjq09ByhcBmKP81n/jVIePWRu5SdJL8lOmOP7XPhAwxx82//GEop
mXdgR7FT8sR32OBxKWaVMco/DCSXXydzuMQ5vQZqobtILWWvEA1/YHOab8hAaF3v5XMP7RhttksV
4TvETLo0M8jY2G1fnrrpvL54WFavtvnU1Gmt+xKNCXjFKmzyiS01GFtbAwGmEKDydMBFxCeVD1bD
DCulYa5xRrKwg3m4nLsv7qRkG16PrWZKxoimVCJdjAgzapNuYmmFCJCP4+03uRDeiwckfReM5sCL
Ec6ndcmRw8ad3l2h/JVF7BKjcxy/qAJr543+l4uXItSCVeOtVvcZvnXBkkcn30Lv0l992BHEE2T+
QjOKCxknoYqyFDyR3W6Ej06m1EwlQKkN2XXmiDHoUoeXW1Ij/g/vpyiFaccXo0Ykoe+xTrFYwVno
l/zGYZCqGxFxAgdyG+7hLAsjzYrW2EY2VLOXHmSwnNlg5Ue/4IDQiTAqJf+DgbTfAs29pjUac3yu
6mEbQeJB61YQnrdNa7TNAkXl2ettkF8DI13+dmSeqLKy04ZXYMyvsyJ2a0kE/aRXQz/Xw3c3mMHh
sRY+1NHxSw1hcy4DQaa9K4ALt5gmZReFwLpeS5XQbh6bmOFleKmzRbgx/yGStHvorWnEZ7itpZT5
d3iYrtj21mXaog6QHcRaTd2sqUY29dN4YhAe9QAHUbp4FS2OGEYYE0g1nRzWwHpEAWJa6b2QyHqy
xknLWwygVDDCfnX1XJAMFrIgg+3JHd71d//pYBL2JSyZzIOj0IYMeXzHRuaGLzJe+8hER4CeKlJX
nDDxz7Ux+ZZ44WUoo1CGyXg3lGJ8H/vsqogrVfDWFIve+ZWgyL5VXWeAB1IdLtY3SQtiewJq+xXw
vFhElaeNUCHPyhvlJXzxl1/fYH84GlO/Kjtaz7IuDuH9VMVIpwWf/BUtZSb7H1MjRNLbDUaD6kDz
4rM9xLCHMiddfMU9JHJN10rqc/F7wR+rVT6vcjyMLSJPdt8aA5oO+7ctW5FLrIUcK91pv0NgyVPr
wiw98cpzMtc2qvL8IuUk8y/w4fKHSDF/dkRgcgUthwxCL0MoKD/P+Gl/rgLEeo+BDY85tQd16klG
LnyhvhipsdJvPpKx1ji6SyP1JlO47p1Gs1UDRF/1TSud6u1IQMRYeOL3XYN9g/w6JDyoElcbitaL
XMpSC0FdEhkNsZfWB60N7/mxEjSt05MxSulyMsjj9pQ1Ecnl8o7sK7x2FUxLulFP6Apw2yv1NI8R
qPc2bE8CZsCtWY1Cs/Rfkwq212FSFbevYyTqTqw9XpYRFn8w+Fyi+/H/2KF8sIgwCE7HVUke5np+
tDQD11bOnwr48REjnQMaa8RQUlr7UR6ws8zcEB0BN3c042QyYMcYIabOgTlcjR8X1Fl5Fa6cBk5V
/ETbaFJ6kmIKdPdOaUykyj0L+XVM3di5p3sLqBzGSSZ+PxewQeSy2sU8/x8k5PBwdyMB49FLMxrD
e3dLcF4L8VdJCqW7B02v/tYx2jKfwPJKL/J5LL4AeOWdsjHcLYiQmasl3cm/KD9bGdHknEsmS3V4
5hpOZhi7LYAVe4AkyVOLF1bGpCVCR8zfuz6cetriY82a56HXSEENnMMy+UkpyZfp5wZj+xzTCszc
6dU6wDGPYKWSd8LVGIOl8ENmAWDp3uTUCvThRRq9Bmf83qB7KzhwnxJSkOGTlrBOmGYR5an4VSKM
2i4hXgJozyU+/8UvAW9kBDw2HvvDjAjt7rwamj0zmafl7pIth5DxRfg1J4yFFE+m4+aamdRoDuFm
DlFvBY+cwwheDI9XGhkLl3QoyKFLMDXF5FD4jUAYhJPrbvMJuGHHpmRwFksMy9IF3EogS2VNtC70
8iUhCoZ1ydWTcmbI+wxek3oReZ1yekA/SxoaLp0WdN+OHTZzasRaFWt4q+KgvA2XpHdTY1Sr78PL
1q9DIZJr4IlVJHylhSYv23PdfgK9s67pxZGhgNYZR2bnoB0ZXZbJ0K1gVRnv8PqLKGMMcdoTmWul
xFAxvB5hywJmZ8d959fkJup/2uK/Y/uXIEioYLBeRdzKHvOVsDxSS2aXbKe4w8OriMrzj3mAnrAp
hshArV7L1VK9UviCNwFKir0Lm7nnMC21ConITgjdHwo9534vtzc/t5+1roI/MVjKJMtXnyPcZzP9
Z/9Zp/iaPkfUnpDEx0wLbDHIWBCSgWd7iqk/CC516oNbCKta6QB2d6QESUkNC7hLhRrJVt9TRa3J
q3nQCTrqqzwYm4Q9C6GmlBDmBz1LyKGZbS1+SNcfJGB1qjvghbUw6jlUoB/36/UppEZmJLtPfB0/
QIzdZJBSB6jlM6NKgkv6yCDHghES3/dPb+GQAp67xswgZiQlvuzS4IhuAms7I5He8KeEbgBH14Zx
Kv1O0sJXQlYs4T4v1YOoxUDQpElH3crRtDOrU5LvtmjGBXgFMbEu2jJMdWUREJwHH8M8z33yYp20
gpVlg+rye7i/lNxg3riAmg6Y8OzcX5H+rx7PDECIfuSuT3uCQOLZk3h/qJ8WOCIdu1yuJcUR+NdR
JsV1zWwEID+4TYlNhE9E/XF9U/2uBWRFBMwxLHIdl5+rPJnb358kU1Q6bLPwcWGX1o5hAX3TWjW+
d/WKBs84MIIv/qO+mHR5R/2JxEpFlhcmQbjkRwYd9mTCGXYJs/2CDZmEZzvewgXEod3IM/OGaNLn
Pmvo2AEoO0T+sb9a0aAncUY2u5Z4W5EuzQjYCTV3eyyA+oOLLcstYepdVaX2M7ugookxQRFyLkIS
a/8jnv36gPDl4SDE6415JDASzvQ04GDIdI+qEFMnaIowHubsRDRkbfnXxeN0ee2lgFaZYS+T6evO
SPZCL9Jr4T5K5+iSIfJxTq/r+nD9IywYZLs1UDzb154FaeS/eE0VeOe/SRl3E/3kvMegBokgD0HF
DzFzIv2vafUVOSyd6d2KOkO1MzOWm9tpaaUsKQ07g2aTXrhQnnskFG8v7u2g39nVJ9pcRtNYX/nW
EG7G3KiCfpFma7OYQOgGtBvhRAVBoWfBj0pBlWgcBI/xT/8jc2d1CfCSDLxm5EnFUdrzGULbqsEj
1F4c8OeKy9iyItV37kBhsuKVioJknrunDM8fAb8wGaGCgQKHYxBJ/pE0W97nh8UVmnFh0gEBCkxY
MiQWHuqc25V2jwynyao5oYGn1IeI2T+ho09l8WfgkLIJlACRTrz/BFvd+Ksvz4qjg/K+kDLBOrmV
liIwar8XEGonLOwd4Qe/+5oSefgq5R8tQNwmG3Z8BagmSMuGNHUGKhHk3g7LtkCgl3fWietpqWAI
O3HSANuuViEqLnQADtzgAd+TweS21SJ/gQPrHk3KNl6u7H9asiXW2/PxmH+HmcUsT/YNhw3fEVar
Fwi6vRL6cB4svhwiCdeXcP8PUB53JSYeFMCI0jUWbK6QWcwAhIQkzwT03QWFUXD7C/Q+S2hMxfGd
AbeBEv7sBBZxqU5kX9aUm84BDd/VIF1RNMp6bLMTYncGJ7IGt8tpefPHxbXSOm/mjry1WOz1Gb30
zrauFbHFMtPieX8DyQj3V8XL3jPv6kONjbAvt4CtwQ1GmWCIdHs1T/SkZbVT9v+RjIJLfdsIV/Ir
DzfxVzqR7vLkH2e2auxE4xMhrjj6qJWyZ1IhnXcFJMzPmZgzJU3LpqBDtK4hAPRuQreQ1Nf5uzEX
Y8XTFAtz2gjDTdIf8zzpnAmjuLAs6DcIx7skdBaQYM9A40bAoCObwF5y1zxKqh1wzeHVKVFQx1ti
tlR4b/qNbgp8LBdfgYjYvHnwF5EGUTb1wxVbHgktRwrd3VUTNrZ7WcwozB0KTZVEiQgAiUGswLvl
qCxPHcBVI7pCaAM3INfnET/7IUJWtKCzoU3SoyFLCfKCY1c3IBQ+C2dfx4q9ibmjjy0XeO85R99c
D3wJIUbezlNp49t+/O1zU2vBPTXQUP/LZcYadZzJEMKdW1Qu9duf5btb4RR/M0TgFeOFqFYXqNiS
dAGmr8vjfRqDHjLpVRPvFJyc2KtaPpjhnll9QS63iNK90PreiOAMrmGm9OMJ7j9e7Fxld5WhPHzy
qC0eOCALtoMY78WB8M7TFAcnNEsQH3PBkiBoQjeeVVcfSyA3y7XveSAZ1lgJPr+AWbzC5k7y3hEl
5oIMH4yzj+onva2E7PiyCJ3FytRX+8mbfVPIN2wumD9nc0VBtt2nL/jcSqqhegzF3WWN9OZO5VRy
XFGgML//WufP/hWDRHkkN53N2Zv2KX7/0ZjQNz77aEHhEK334AfCILIP/mDU45WVaZjCkChGhjcP
MVzRvs92hmRyWjhgaB4+UJFsT+3FXPmhxprTvlKfcjRrz2lLk6vhH+f5AAw0CO0B39GNmRKzuV8M
ORpdlHnP0wh22udpnv21HgkKmwnKm51w3X1MVisEUfWf8eCzcJp8y8qtFJdrvukyvVvTroQETtUe
ifzHGeaw9XxNfhbRFo+a1EoQg01OUNrnh4sfaIgU099bnS2X1oKobmEfW4pOeV4sIzKx1i6tA/w8
HHBMkUa9b/4MsgkLzD3LmnWmV6fJ0snKrxR7RGe+OD90eoWfcmHSHoo2YXc6lWOAgyVz2zJi2NCF
7d3bYApY9622VTsAl/d7k5k+n/1RcpIHYcV49wJnrn5vDB8b0dltsJh9sng25reBL2RBymfk6kb9
LUGsjc2mZv/QcECL2e9PYP0fsGCRNbXBrNjTuJ2C704cF5imkKM4SfePd0nqBkFMR/1ko2DkIAhh
LLUTth3VUuORtg2Vp4jo61uFNizlOblJxbyB8eTlwR+6uSRzsFLWdk+gfrPchXsRNd6cEHloczEI
RJw/Xe/rxv8j4SVeS1dOKObyDVnyPvRaxcQuBeBtyG8U+hntKh2z5hv/2YLHoKqd6WRDv8oj8+NG
e7MlvbCIhjlI7aIBZclvt5qbyxtJFl4yX8uF5jleUQmAFwb44JaoO1Nmp09gRXWEUMo5vvBKjrcS
1qtiKaa5x5AJIH9pmpQP2d0XPHUwgvoKVs7QpwaBiykGaLC63G1jNZBEDRYE199/A95gedt143Ot
tCZkM2pNABTLAnpQ7hP+FIPwcUm7gqZurqLJoj9QLxxmRiH01t3kltT9lE7nG0zC4wKMXv6d/XRc
MvjlaX6NyJeMdsvWt/RcHigocCbjpQikeFR2xGtiDdhGEDrWNlizeFIsKSijEVHkvkpiz9TVxllT
ih3nUTVeRVzJll2BAp/u7bnrK5kFrF59JL8RQ/FmDWGY+OQRDn7WUuvbb3gjgl05M3lPRiZMRBhU
CizD0PrYbmTd6eVXQi28ZS+bGnR2PilbCFkjyugS8fjZdcopV7aTWe7v9XBm9kMhXONFaysiuwwO
zNxYyGYHjSufNx1+defX+FCM2u4v9/BK/J3uXP3QybOCoDR3EDwfS5k3swQForGg/lKKpusG2kF5
pPlvd0qyzNa69nrxaTO7eHy7OvzPZv+ru/qCfZgW7Ki53zKOzFG4wVAnkH+hEox6rjeXhqgXQHcL
UrMBCmNUu7SfIO7v+EMEVGhSaoY36lxRa0wElVfRriPMJ0ewOEo6LzhRFbfXwunILoScjbKvkmCm
RVmcRLBJqmVyuaXSxt1O3KUps7N9Vp45WL+hfR3bd6Q3ORKut630Dc2ECfU9VK8AqNB81ZzWAtax
KoVqMPnGomSa6fD0trtRtdH3YY8ZhxKiNeCXVpcmm2svRoVjLk7bUBadW4SNfCK65xrTnp0/MAb/
wDIXDuBIZa179E2sdVUCGhi/6Zme2szypEy9zFtiJrU+Yi5Rj03JNLfAyDuw3GzOimE1pYTD8XN3
GzErjOfCAU51wb0Hj3ZyxZ2qSEAQY69Nsp05Zgg09qPJKEN0I0QarObeWNUwzafh7lYWliWTtL3M
vkZ+o+uycvEfhMyzdf9voC/q0cbJ5Bg06FracoT+hIeG3Dvep2jx2FUiSnvcYNEIgbdo+3Sw/1ft
EI4eaWl0MXWf0JIFbdkGQCPFKnsoTm3Zx+dxqbjK0K6lXaioFFPP9INy1VkrG4WCfLbylnmqjefo
LK+3dOqr5qqJiWmM2ywRZgKKcpNxLISlKb4yoWUcRrCjezdcnqXQS44vUPH9gkImzuGrhHl5GI79
tDJEYN6i3LwxqYWl3KLOfJnkC8vCgK1QlmAQPmI4TR5jc2UloPIYOdJgxF/AQyStdXGXU16S2pdv
KwfvWNCk67p+YKwq7ToySXcyUprX1LU2XfYtgKalRQTMcjgzioamfoLCH2aXWc9/R1TmjicnpE1p
gqD/0YUA06WxhvEJf9+9XSrAjU8bZ60qovPhhTXwFVhpnyqQitnWlHksKs3t/bTHF/IKPkMhlbcO
z2BXsU2TiHO/GQnV8F8VbaXaG9JgefilP0BaFC1OXJpLskyhl39ols7bVN6N1zQUj8kNr++6O3KF
HFKeZXDIwG1aytgYZvyhugJPYi/6R/wY7O+x8PYFEGoJU6ciq1mhw9BMTLdxOgRDFrpF32l+9ySv
G8TQp/XC9YYBL8DG17SjKQT1zSJRyhbCp3y6YLVy8wI83ZnOs895iqYn9dCR4XYatz61K5gSBiqF
XomfDOoJtEkCRbgcidjrK3oNQe0f8xUb6Se2tdV/GE6/Ltm+8a/a8p4voZZGBaWK7ykZ8RAk7Hcl
J/R/ZBIr8MfVuncD4wRV235L0VVk6UYPAI1TTcBZJ4AfyrNbZoppeRtBR0VKaHC1E299NcRPgd5p
CBplRGA0/eM/upQe4Kl/Lz87E4aI5IuTH35l4rrx7YjAQ7VuTjsvakUlVkLGATMRnzbuuqkB4wST
suRGS7HOfsFI7MM4kc8jTAxrUGKN5Zb5rdBeX7m1d9Q9BVfYBCILJYjD3w7Musx+zdN/AWp0JQJk
n6ATG664aO9QmrCCh3t38Bb1N/Wfcjm4M8EJkm4mqMICd965dKpOgExO6DJZ7RS4gxdkDcdDcnoh
rGxTWIvrfzO3LIVz/kve95OHPc1Pb3uPtVESlqxS+HtFBCtsUiBHgY+Z2+3FAysJAo3pITNim1TQ
n5HclOcqlNPrZyEgk/7VTtqgPrPSaujmIWsiM9cFIjDOOwzZZVJzXXx5KxYzfhgJ6cIcgRLRRHQu
K/C7qOMGJMrjwz5Ogu93WqXdf/D4IYV/uUrR+Sk6GTnwAGluTzJqzDPSfhzDjA8hjiCJrgMGexVf
97NNKjqHrVhSirFsJZ6RSbTbE+ieZVMCFTHV081MTz7MFBKkIujQ5nBwj3JAQdota3DgiDpgfHJA
/KPTee/AgYRyHqAY0Bc+b9IyAo1rgtuKcCoDG3XCy/Heq9AWzw2DELxCCkI6OdxYgJq4x65v0iFW
wu8Ysdkyt97iaQLNT/tiBFxeZhkUEjYKMgB/kDB0BRpDYUpuYkIwwoUqcyFKGh8tEQy2yVKV0WbJ
pF8woKixCf7v4a8aQOxUQ1AJYVUQq/10ndMIMQ/sg4pdwVChNJVEbmZja/nhN9GB3xrDAoQ13HpG
y0S8sSdbWxivlkNrk/aSQQ3woy3B+MmPIy8AfHrEK5NNnmhzFr5NR9P8lVOVJ4AEsNInBLf7o6TH
90iFCLTUpV6nbCAYGzh59szbibYEGX1Lxa8JaFEU+I7srKs7gvT6P9m+6t/JMaq17hxGHhL+d71e
idsYeqUOCEomuSsyydub8hJCQawL9KYagSfJLdwXJCPBd549I42KMxNWwpGlsceV2EzEO/kVQ5c2
FPkOcILtN3EupJZwyQKYRBiGj2Q94qxCoGeifxCr1Pp+bp2jFZgSqB/yTTpmY9oi/+j0IuZ1uw3N
K3+ih+y42zgOisicuQ83FZjsWBlwDPx3N7voWspXIOQHcjid3s1YoW7Rp+m8TofSm4r6Zpi8sTeD
bw9pS0vCKxdV66vG1ql5mJ+bE0QZTPVw6+MgfStcucfK+j321ueYLk9lrSL+Z4C1VF56Ly/2XgNW
S/CCMS0yauSg2G1LirISyuhFncZe3v04gZDpIePcM+nE/x3ojvU6Zcc+/5A+iweA+Q0gCUBR/dJj
FYwQPptJWuPJRV6asGjK1cG4GdjfvubtYomT3T+29DtcJn85JLNBnlzBpGkQktnDWCL14GurYM94
AIwnW1xGUiFi/+9+fOOA7chjg2DUtgLDsDxXom7B3m9cIL3HZr7S48kohltPjVLpOdyW0BCcfKEM
hRmkFcioYU94pNlSuUpuQSfyBEt2TfX6mdI1b/pWQKy+0MyzWbX9YroaIAzAz/puZkNpILEnHXxK
TIoV+1O1IJJ4PVXbHdmqrBJ2mU/eHkGvnUV4XcL24uq9/gRXN+AjPDVqbDGzORhN+RFStomFZ/H+
XqghxbksO852Id60J26rHrh3FfcJg7rSW6gZ/JFjRx5QlpyjmTt6JW/Im2WhrKiThvC51rzbU5Ie
cU4iyV45pgl8OBGmsGD6JT+y353A4u1/noXsBQUW/JeNMLG0irjM55SW+TwzXlEurAtPgfGrdjPa
CKHeChRAyPZAD9S8X/rAtKKzvlXiYDpy4n+wv9hbrfZMOFrA/TDVT+1kIBketNZ/tdF03FEQUtDh
kATu1xsEHstLrd/k1E1BCPEJyn+lCaSrwLlNTTgBpb6knBPt0vun9eIXXU7WJObdkelNBxqeX5DB
9KiKHrrOHvrdIsnB1oKn/yLL5aE3XpKXyrtJXIRKQK976C6KKSnXwXmh4rJvSnV0T7e6yEWujqgu
w69Kh1KvxgoUoTaDt+fcgOlhyiD0doxshiMy0hqO6qZiMFnsuUMKQGDSjntE7aOJ++8+kktfWgZF
W87EW9W4L/MBMQ1YPUocmXDzUrIbSo3S1jfgmI3U35chcw8p2FWAn4OhGStLWyY+xDuwCBuy7QOn
od/gPSnz3OzGt18KQ/aoEu3PUW4OLS1N3J7k/OLeGz0E3c1a7nJMuwNr1Lzh91hJv5kEep8F/8RO
jERKEZT3kyZ6FvG/WZAqOK/yN3DsEb/D1bF5dGR8Vc9gTt9v4OtXZPxv6BQN+i4d88FuFGysBQt/
HxwDbn7IgtFinm50d3798eGJWjOf4AIYTOH9MLrMvh4/JRj0IZaCjGPtnXob8u5l4HHWJBpwL0y5
KvVBA1HWglC4Gpcn5BSFo3wuT4i9x8JfzmaRNLkB0t0eQoqhZD8oyTQfnertG8njCYKdCBFVmeXV
Vmj0Gv5/k4cm3BH0Ni9zzHgu/JaFL4QV8x4guNcfOlbGEAli1joFc4mFlLmTQhHpVrbPF5SPbpCl
fUvfls9iOZJFOQU2GQM+Q6RbPpnAVP4wbyroFEDsR83wnZfotdVecTwFEN/H6tQRFNW0ROQunnKm
D00e5E2POwlGZLiM/QG1EBTlrDfiYLdEZ5m7HVoAyhaUseDkYkoH7WOsSTQ4SOGnHEGzWkPqPJ9k
CRNXi7s5MoyUVQFUuSegxZCFs9JkyWQFmlxCn6loHQtKFh68aboUM6kvFNrw7Y5V3y/j3DB0/KTD
XGY5lfJlaQW1O6iuATE+IvJxIgi4+NXsWfqA2CTr17jYKgj6dJS4qQh/XsPJ7ulbQv+9//xA6MvZ
JVBJpa462M/MoWk+yI09cNxm/dnRWi4IvApNTtQs0/9aLqDRSh44D5QT34TIHfARnYxjSHXY++dT
f54NtQnFPsO8UxzIt1SPAA/uV6s7rRn8hK6dquRSj0SEgXLiXrdHgC4QAs0qDumOaJaaO6n/dpYS
kQs+rhCYekH21iuqM6ntMGUEiN23akBm1ZOFTQyl5e9S23FglsfUH8QfgkQ2dlApaZ/mkytpn/ms
F2R0vpLPAMX8b+D6xahwwSCpYkrq0UefKH9su+AeeXPV96JCmAFfSqnt3OF1PaRdLxLOiKTapaBa
7j+UXeu5VSQie/tFe0eXIdjKWwd8UenSEPbXCity7ktPH+8PRFA635rbN4AbfZ6E1QEsVtdxk/aZ
NCH/2S+qeuRsDGzPjsakH2gwHZ2tQwYB8ewRmO7BzknUG6kaV6jthokedZb2bJ1oE8rZoiPfwu1v
JivF4u0tWyCYOROBth+BXg9rry87ns2I6zOpLiDN8kR8IMwsRHwmW1DaPHMNK0sqRNnxDogX7Fle
x5873DM1jdcB/0Q3xrzFNvlKMEBAytLoPduDl1efs0gB5TH7Fh39D32MYUbmfIYBZXMJOe4dpDog
ogh0CRcCXVBfwMaasHk5JhDbZrbEAIzIVTAVCQmjUwDEfsHhvdmqO6Xj+5xrYimxbOEwbWxfBr52
Qsh+WdwtHRH+TMoQCnzdROwEuo3wd+l0SIvEcgiUv8G4ADmjELi3fYKqNJEQETYNk/j2u7SM26cy
/2X2OpfWGf5r8ThE3BiKOkFvdNO5TStp0SNxAPYfRHQ7xG9t/J2tt6PAuR85plKQ+lACr/MBJtxH
BWYOATkbAIep+ZChJWsPBqz/iygQM8uHedT0UbPfFOgYKydXGyllKq8x9lfOeufU2OiH/RFGj6+8
93M4RFc7JmjFouZpzO9y4rM3ZmS74RDlnSjR53ytStFl2NLGrZK/sAof3Q469w4BUjvCymrfJ23w
ZaQU0lUizfvgQ4YKGkRIZtBYdnoSaUW6TnqbyXkiJMeJhUo8YAJSrcVlEtpWjunCvkcf40UnJ/O4
TgXsOmSxcdS7v/mWXZCR9ykVAQvQPzywYSz1NF9Uq4OU/zOtYAzzsq+qGiNoEvXaKu4/iWcelpUW
eEuiGMZ78b0OM6XJLZRhIz0c610ycazdcVpI5tQcNYeD4XE+l+cpELg89zUhu+/BIoOnyWJkUv/G
wWu+nuLTfbo88PVFi2vRRkz2lPHeaBW+fsAs/tagSnCV1Nfa07+EeaOzr0qSuNJOPucMvkUc5am3
RvmIg2xzBpDstXu/OhixwCRyjE8hx3dtMWHbCEUJFBR+9HHnI60ik0t5zmRcYmoMZe3XTAQgdn6o
t6em64Jb5NoDSlUvTciaixRisfN5BXE3ZjnrDfMJe/CrpsfL+BnCR4QkP6ea37oIacF1z9NWuIsH
vvz3i71ervEJNaQFDwO5aVRRWAAjLFDrr9LCYa66CO0BJ2/IL/j2eQNYbjAfZ6glTaikdLLqqi0L
o8fMrm5KXKvOFhYVkKlv82KDI8+1Szh/70YaPK8rFpru57s3/HzWt3fRdNOT5OIUroUz/HytpR1f
g7Cr5gy7ocjca2g0OaAVKcj8h3+PqNl20eA80T7nwtbs6IQJlbGtAhUUQGqfUjcSmARPJE1cekts
agwYGC/YqIcQupoOCY4WGWqXTRdQ/++0cAre9nrex+x3xTW3CfdTgK6RiQAkWqYmZrK+4fpXpjb0
8GkqJjjEJ17zbRzGj5cAVt3wHIC8k7X7fP1IWEYuWAG8hEjh55n/pCi4fPrvnkaDWirfFm6DXexn
qXZaaKbuPLWkXBFi4fQShS81DCcObvruaM2/R6OyC3xmpeNcew3dEHRlJDhkdLN6c2hw9BsKhkYC
4F/Tk2tuJTLmO0VA1uPIvuGAup52zKENueAcZXPaPmeW3kWW17bydU+3tybMzf+8YwlMfeF5zleI
IoY9x4tCOL0eA8fjKub/E6p2DMcmXUmxscVsQbDNA255IkjJUfMstaSnetHdfG21gHXyYxPszQ7N
eHvoVVx8zMF5T8C9t4QkBdXVDrXiAusqdGPR7RTdkTrQY3haibuH9f4jVHgtB80ffav4K91y0bIA
VC/Y1Vejjm3gLCUCv7NexS8S538YnW/OS17Kikfv9/tkudSwOBv9lSaaYmqsUsNaV6WHgLr+0i2t
wqqCnTQTotIwJwYtEy4GKr7NoEB+pLROsJA7TS5+Qx2Q0gH84WQQS7flEdcUCD/bv/PJwlf50wX3
BI2bw/WyaH6DePOJf7EF49XEDuRKC/Nvyw07wjP42Hw4mkiAvYVr80/pOubsxTDz1K7ccDl7l1gm
xLB0arcroQhDjOEyXdtVjsL1wjO3kq7bszANpuKdrGpIWaTIYMg4B4rV/buwBGrVQo1GcKl/UQTz
N596srEzkiTDbbLtQBBJ0jSW6m0DF0AjJbTd6AkFVI9CQJ+WdrYBXDWngmqG6TajiJpICJ3NfcYf
MkgK1xE/NFK/p4EFGFYSnhSIjv6gfOzqEr7ks0LTJ5awtS89iVRuIHXT4rPET9Jn8pBirlGry5ZF
Nb/JL2E/a8mhWjLpjutLXwXnXEaaTYiVNJSgXy1g4wZbRiraJxSZXprrT0dFHfsjh+3i1maPVJgj
IDoMEc/RP6YCJvMl1eZn9/lrDTC7k+JFGy1sJOsanSKBvSc3Fxn+NUpsu2k9XNrpXaELRYXHO0Cu
Z/4/ZwqbL9lHY/VCTUKJNdbsUG1Ul+sF5IOZS2Jy7AZFCnobX9rm72/g5suGJvix1I/X3O3Rv+Sb
8k/UUF8UlinAASfI0CPgbv9D6pov/g6uwTM8cn6UZ2pzhRQeUpO1PaojnzEtFMicITv0ICsY/47t
0F8JY1uAUzqVP5q+umLBgM2EjmRT0EkzHWXJN5EQCmUvC+DlT59Nfv296joxkGwjDgyRHVApUirf
2bBdxdD+NqUdIX7BHmNzzArME5o+jL9yXdTPE3a0/ex4UkqQcrCHu8EQOxmeRFtAm0g1aNF9RWQT
2J6MwVWOI3u2LKjew7vUMbqZGn5zh4xuUYo+vq70aks4pntVmuWjH1VOTj/eRsDYJbu6rBDt4ROU
h8GEPwUIAlE9c4CthExmkrFSwS/qwleND/edMxy6gkNfbORJlxK/+NwqLQz+offlLxRlHlKYy4AD
GoGkO/DxmRlyJAHvkO/rQcuPPpNJAyV7I6iH30U2LBGNEr7HfVcQwR8KVBtg8ap2P0po+uJ/b26K
lBRQL+LbYhSqeWDgbg2pVAdU4Nq7SIndncZEJJaCb5LJSC4nrU77TPDJnefbQbhXu7yQ0/2Knkpm
MMIdzUJAne1w85hoeKTTimNtLm1nAh/Tf/dbFivPOhPbxycNWgo0+oQGBFJLZkp2z3Hu0w/Ntw7c
GepQSlS3LVJYkSTahtxf/EaJKK9KSKzKwNU+djx2XwJD9GuCyDS4B9uuy/fI9j4w86pCG0isDXzk
hIhfhxbQpeMbKvWmonQHLNYsyTJM3QVeo3R281KLz9ODmTrXdmAl5+BKugMzwf4DJc0DbhI5vUn1
4ijenVXTpidxAwJuqdVeAZzxJRAcgHbBbTT26+477d+bXHOLQlATRe+aur7FCFMj74ruwjfeWRCZ
g3yUd8BnB+E1JyH6Vi/fGWR5amBphPiLSQ1d922OlMCOduTozrZiT/GtbnoKetQ/5CuYFV7SyqKo
pGuyZ2jH1+cFipAYIo+AmCPZP+nEBylLz11Z+eg9oSSTkTjzmVi3Lm4bV+Zdh/On2jVIj9HB5+c7
jZ6UZY99RSsQWL8d+yWn4F25XQ0rgjrct4dQgwDtR2RNg17EpX9Hg5JFP3wWdMdIM01veov+ZBcR
AkQkfLOFDfeIS+VzWISF6MjpfzQ+fYv8J+fjkrTXWt7cS/OTGU0NVPC5rANCtWTH3G13H26L/SOz
sHivqjL/qUWMM/hOuv1jKEVUMiMNcztK5BASArzaNdpybFsmHHjOCMC07HwjM61fhaNWLF2ZjM4w
54gnv3+wmRIkqu5mAzSjOw0Ho+eEWoXAy6TiZZ9FUghc6KAkia2HxZLTIgZ9gDtNCT/Kh/gfDT0+
Ipg4J1c3RzNaIHjnoPzUsI//03FvPTYCFchqH6LiWOSara/TDVyPArpeA15SGNdc0J1IRTb3yeWg
32pTtGTxMwc46wM7UdmAu6ZWfj5Da/0gktqNsq9baW9SPEhauCHOvsGdwx9IGUl8LBUqtqr2Nz8S
4MbDUISvIoK/LOj+kA/crYqHInF1yisZTb1iEtPmgJk8t9ILlKMt5nRIsE37r9oNgFLjtw/cRUUK
alMeUjS7ugOBgRPXYpXYa3FUGTkKWczCcRJdVup0XRVLbPkY9Az54cxNsLX4e8AGLkDWHQQIKcJf
riuXUdMnx327ndiV3fO8g0mq6vUEeePZj2byjhTz2K4kLUZGdeMNDEcX66xv43oPKNu4bCfwHCDe
E7zwTyb8fWu6UUj5OhR8D5+IpcmpnTDhAOHuUk9XdJ0SqSL5OdNul86PhV2vgOmEE00d4exOFeZt
zthLBrtR2PTf6tVdHuj3O5GjlgHs0b1Hhfk/C4Nnul+cfPBeQh8biQWVkOgcPPkJXiRAWfIcSInl
QP6MnbHQMV4OJFGlaPcW3V8shet9haYbBKJU9DdLLQ9oQBIKXnbV9pexDa/jEJHow5XcclRE8D6l
QHTr+Dpqzm+qe6MjDmOV9GwsA6H62DoMwReiWiUo5s88r20vb6Pwkn8bmhynsSSKvMp/nkqSDhzo
uhjWsZtBsSGwvTPye9UPPNq2aTQ9Rn02f1kICRkTQWVRt7/naDf5ZwQaP105Pd6rOSKdCr1j1Mnn
kugqvbn0ssREXBa3HyfRwbuAZYU0X39ZtQYHIGFadwQvKYDaM78M4ZrvMOTH5zJ0R3MzNL1eZLQU
UwEGgbzVRw3Cwl0sFjBlWm4UUHgxlKHfAsmGGJpG5DDGMSUL0YX3ZwdCQpCyrQ2U0rr9JFVWreg6
iqfYOkJrWgesFuV+zeEVHHp6V/AEOXT8DJi2Xh/T8RKS0VF9siaYD5Dp9XVTUuVELlTsS8WZ1PVK
nZW1wokgI+rWLb2zQPEcBgMCiba4zr4lSbtFEsIA071oe6ObkodLdSuh1/EjGQO4aFxvBkNtFJvp
5yGK8iS89oYaewtXlDovnRbNWzcDBezkD+2J4y8mlqhzYkRkv7sJ2ja4Dm6miyV15ctsVbGfZpCt
ln1afqReMuYJnHbnp+6JqBHVWJWhfykQbbiYoYChRfSuQc0KggXhCHVwHwFVJPpIpHIds0iw1gy5
Ghrea5tDqDoaIQo/mqoDGZKoknHPVkBrq6t1nn2XK66s/v/yLCVdrwtGbxwPYjqf+Mn1EPyKoBG4
161PxX/dUKzoT/lScVhaLXTT5ovBRu0VRAwgg4+SZkVpWArKPOJ8wiWYyZvHEfaDAud5U01N/Stq
wy9lI8FEXyTPtjj2/LTBiSIPxJC5JIARIjJlnSwkjbmDa5RHPb1PqhZjEbYW+0qGvkV4V7DdJFbJ
DvTK09OXDzUIoSrON4n3sslNImGvGxCER7SAJi7M8zdu0Yg4BPGvsebWKBePfcJgKdsxKgPTCLXc
5RAUlx22F2RABRlArBGjkAytbQMpIcIf/DKjyVlMYQ6T6mGFnGiPAiMDUICcgQF15jt3FZFC8FT8
pige04KqI3f7JGrovKmHfG5kYrh1no/ZP23P3UjGyFnOBjk2uHXQ8N7vWx0Y3k9laBPxb5SOPKUV
AolOFCuUReM2zKuBm+OrrFPEqTGK7GNYeFrNTVCj6KQxiB7qXkDG+MFrxbKyhRRa4N/YgG5GIy2e
dmP0jKaGoYpVkyW1NYWtZY1rIhwm4tYvhPLC0bv7C9489ZmlOBWePAe3wq3RuxzTI6+qUlaBVCwH
efCoeRn9Av0/kZsZIK+1mT6DY9tt4/pFQSFhZGZydSa1gK8pz19CNttfJSlyRRFKl+oIpjJ3Cd4l
T8AKGSMqz5r5w2unTgrCMs11qq2PWy1OUQ0f8yOsEHtjXUirBFe3lXCqPxii3DOnBlHHab0ErhLM
Q3HAeJ/cYbrbhg8v2kItERwzn3vfIVvJymGSidSltEyG7Dr9ymVBOGHM96p2d8xXwIbhHjuLVc18
cjmIuVX4DkFvNYyFNlNjaDC5F+echFV87yZzXUOSHWrQtXCA5oGVMisPrn8CXWnalt2qx8h3uy/x
F8o4itDvt6/vhgnwH6pEaMsJlrzp/yuoEZJfKIIXDDlAqkOUi5wcQk3VvGAKcPw+G7LgqetXf6U7
JtLV4k4nKlE8dWR5rwjk85DRymAIpZm9kLpYO3xVpbWrn7SZ5YD6/ZdnT396SbFvJiAVhqo/dCj1
MgaEsMUdjgAu0wbqEGFES6AU+nz9T1Cj0j6zKVvGOOyEpUfoySfVoggbH/cHKMXhTT2uw4fCj+uC
XFt/SmyjGFluh20tCMs6HXO+GngTv1/BKRowGxbr78UKNNdsxvUPHCu3dNPfYOz/E3CuNMlb/erV
zw2f4+YwkFSVI6TbCbMV2qGkqjz2/SWXYUrYsW3vTKn4eSiCsLcofG/mSj4Qeun0T8prN9EcR9It
GsavEZDYclXRi0jKTiTrIehPRAMzFgTELisWiZlpTHx/jVyFdMf/Xzo/f9ul1v19PzA7C49wX1e0
VRi1MxWrVX0RRDV9KHROw4Ck7CVc6A7OJKJVFuZAWhIc75xG5fJzjzTPn/7qy9kwugklksaSnXfG
sKWoEp/SJ988kNQuPE5Ap2pfQmat1wKnVTVVyjUqZ6NBLrCrhwYBow6yg1OAcdoK0zIoeTvCM+D/
bL438WZs0etmHXdP8Nk+FfYqmZvSi7/74yuuBK86Bi2T5wh00F0IaGF1PIjkJbsLvr7W/qrijfsy
Ig06ufI8R3z8IfTQcvqEWMpg9J8I4Uvykr9eTxBXASqRKDUJBtGPkMLjF7qSET1jELHNR/4NExmZ
x76lO/MdkK138l3+GmABsnn7ACW5HlV0NlPinuNsDB0VbUVrCxGYobkyVRb+3Fxq5AcqQlgtONmx
m5e/7C+JyxVb9AflI2I1/ak9ZPMOFpQ3jmOrRVyjjJPLFhQ5vOixT9rF0PbZbnbCY05gYzUOmQyN
eW5nFmZuZ60cX+ChlIowWzo91EjiZ0LJek7EZKLtULJ0EN80RHcqIeTFkHGjNieXVRoDOL1zGNOA
ckrbkoxIjo+FkxMbLliVc9toDDYqAj2l8j5gP+FhPxVIzmjQ7H+5nztagNl3twU6ZW+D86G3ifjH
UQ2LmLwkuFNHPLPK28cJ/AP2gOCLa4/0zw9IuZitEaCwMF1lEwsLCyldgfS5FkmnWbTGBV3XeoiG
FeQlY2qJtGWbNRObT23szyWcljJG0CkSU/B+ex+MOfZn1tzz/Xs27sDkbB6E6rqdtR7UKW3Qa8ck
yNCVCMNE2eo2VsGjy30kaY1zKT3RHrRgCSq/8OK0WOrNNdnw7wTvoMU5+nHl4XppufKjO1m8ireS
RDwp/4K6GxXMcXURUip1ULn5BkMd0M7ycLkTrBu3/rcQIvQFd52TaHgr3sQS7UBDpAR83+jseWWr
J7SAhYse85puyW5J8cMgUQOlR6lUgyWFlBqTO/gijCNcJ7+16pHOCXgSv8du36+suhIM6oeAWIUg
x6Ak5/Wz59E7kXvQcsdYvHMPRoJK892h1BYT7kco83cRjwVqhj2iCxHhQiMCy/i5p18I0dzjS89h
dx2NSMNEzubCH7zEcmkULcU3YG14ZKjL5EC+Z9NCqNx/W6/tg76ThaHIR2gIz4Ir7QPbeDctW+Hn
Afl4saXiPHvpA64EY29WqgEMQdWFB6LA6+G/8UZGt5s+uwbbexj/ETxqAjrMuBH/LgA8FWUu3g6w
Lg6BnZ6f/BS966cML74/cVLSGaXou0FTn8Jvor/GwJsIW6M8D0pXYZ4kqJzc/e7oPw5OwrF+/ltI
+5z24uMy/xKa9rn9cSMxDGXB+Zet92TECBF7WFN8hll+WskjCnRg4Hzd57Q+uhDyICLpE0r/y/Wq
tftNowUxzG5nCawMSgNSqkV3boaOo8gKKiXPQ/mqq0wraRlke/w4H+hL2HmX4UijtJzOoUDyk4zK
iNcQ/BV+Q13LqjPU7zwhS6C7XopfRFTQi336DAiGF3QEPUbUdasXWTaRargOHNHQy7R/1yl6Z51F
YOs1OGD+9nQTpKzRdu8GRWDKySLs2M/6fY1elBfsmHTB1yRV6xfUQpQAGonEt+/TFOo+VzQmrxTG
1CcsjE5x6a1rkmQYhpquvfnyWTlfHDSvqMBx2Ig68sAtpTHVnbXiMHZmqtl9qG2i6VX2rGqB09II
sNblVpk2yIICd42x1ku8gudKTcsDcdUPWlI0+qczZafydrPko7tVMB/tLyB2QbM6YyfPLLZA8pK9
W+2Ntx2SoB3/G2KVwuH8zQDM+zK5IZWN9K1U3S4krZlwhiRH1wLIZplDIEp+yz+ygzZmW+D/pkOQ
gcp00koDduQrwXQu5kM+BWg9KH1oVqFG9qihGrCqm8SCUrhx3Yi2xfFAUzpSk24p/MFRyAdW03W0
oXIPAyZuT/9rFIH1HgxlgTkQ/D6Zw9bQQeDlYd9Q3XnRKAeNsWBgj8Hywws9EXxJ0c9nVWR0XVpL
iZP4vWBw4OkCU/lN6RfsWr9FB62EdMQFawsKaqZi9jpOAwXbwLx6nB+bMB6KIcHLUItyrHljszyu
rpD2Tp0Xt/LDJ6NNM2THfh2aRoWBUAXVPVt9KOPuCRUBpNwYNLhqes33bzMs0mBPUjglsq8jcLo3
jlh0xP1WCDkbUoMR2/enmAzCmzwgexArI/+hr3jkwT0h6ncEQBHQ5P+Dy8mZAT7gQL7PBh9IJR5z
rTBHnALG538wPVQxwW+B8xvBLlWddlHBWq8IseYWHsAvF/krbQY4+9VMd8Hw307MqQE9CZtaT6AP
Mr/4aJIlGK68W/Vrf4DXHLvxvOd1EDNAIJHytH9F2NLA9aU+BEfKVaCoVgFBa7z5WFAUhunowbcN
T8Q1bD5J1/kNgbb+cXI41RYt2GI2gskX1prfC2hEagrB80P7V5imeugaV+8f6ZmtKI6Vxgb7AZOa
XWm/IKheQ4vTmnzCwqh8pgJjgh1RY62LcZ/c/fo5PyY4pJMoMrI2itchLA9BQDs60u8xZnNkEJgK
7vIbF+wp3XTh5TE90peICxCU1LajXrokxeOAXjf3stqAIH7m8D6wrddAjcZ7jeuVDMTDw+q6G6ea
fiiwNUWX67n7jrW5lArIesVVhQnWChMfTm8c8BDtmlKsgNDWWvgUmHuJwC2Envqs8NnSXxFIUPyj
a0pF3OI5xcnJ5iwLdlrAMRCHlauUDNGG0Px0FspndrbOLKuIXiiTpxI5MKlKa5jy1nalic5xKZPL
Y6hIzQ0mwBgI7F+ocBz6N+br9sfogPCFDm+7oHydqx3C5IYaL7PYt7GuEit5u5dPFoxAzicvOjd0
nr1DY5Zi74wk5uiAAQMHFw6EpgX40t47WPvDcdo7Jl0+iMRfyCefPEmXbryoKMD0sQ3iKIpmLf+M
nm/UcMeQ54Gf/hJHVyuBFwGR0eVBDTkdEKv1TK7aVVjtL1ZzxcLwDnCitmjtfOOZsi0wvyK+MZxF
ZTas5nI6NRcd9Wes5bvMIqUkVLzZyMl9ZChNjbNShFSvpGb4RBT1wQInR85ZbJmEVE7HBJDEXq7L
xV1Dwa8FKxWGzsDeSaXPLXYMDzNOs3d+vo0vskrbQUdbqQC82a7/VXEoML1qxMdxhWl1QYv3/BA+
RojQfLOoYI9W1NugZ6nvNp6EOzUHfZ+/GCfQSi6cxxj0GOR3xYgGWvv9qxcGVS6MThJRGZjf/rJg
l6CYZbD/QF3CPwUzuH7UdVaK7Pn9a+cw8krnEnkZmdeUsYe1dA6mNXixBKvOapTXFj7WwiVYDVmy
Wv75bRiT4H5xjNGvZZRIGqs6GP/sCqpCWcFyCjL2JUZlsjRzTAuh/w9i/u6noDnMiKWwYgBDLReb
jUKqktrxzfdZ/HOjs6Q9f3feupR0mzmk7hVBm9Qk9Fvs/uZfajRX0ZuxAJy/prE0zJYD1JPk4z2s
cFTPeVRc0NSbnt6U9idUPxo9pLFKOwVS47xQcJ3fAX4aHi+WxJpSmi3SAwbjXWhqDUgfRj/xtNrZ
QDldz1skGWQmqSLIIeN8WrA/0JFE0K18ASUXhZmUJU07tvtcl8E3+xHWaoTdTgDngM8c6mm/3+TP
A//av9uZVjwXxai57ZtMuE8+anSg0jLY+BEEbayHFMn1pUW+c9hCIA2dv6k40APESrc/ZwIBq1Q2
CXt7kRDDgg8NgElcz1gisl6BGBPLyCnYYtTPADAoW8D2O5OOAJs+iLS9KcN9N91CXmMG/IdkDj5s
rH7TJLwOoI7Ve+Xb1/iasiiN2dhzC3aBhBbMQk/6cb0zOcxUp7zTcio17oTycaz/wDNpuWlF8mXR
MqI8V01B3JjR2L8HQAFu+ebykPgj5YRQ2bPQabn7dqOgvsj2g0X163ByCvPK1MRZStWe+2SEG4KV
Dy2+5nvzPXTg4Dq0qzEeWvGRWu/xxOfqZM2u2nsbgts4ApFO2Yr3RP3rfc9PuzxpnGKaGnG63/4f
LLajNEcA5MC/hTNxIi06YLrXdBxDK58d50Ll5szoKAKvtMYAMTgEIIQrceMKTnBtzhyOdsC3upUZ
XnSvWHWKrbca1BRo+TazpZwfe0osr4Eom4Dbwua7KHKeQ4YwIL5Y1EIO95K/QQhPcvdMjGkOMZCJ
C25nuxWPmX/n44YSIvEF6cK5Mntj0ekOyd+FR23Jt8A1bBP2/PXoUo9KPxveURZgBhqb0X0IMTUp
yh32MUlkXv5S6sC4pJ9aHMT7cLVz7ZfO3JyJ4iq6R5Oy9EqcKPVF1Xz0VMmO7TV4dizaCok7qglq
TitqjWs8KnjEmf2rHn8udXAKHI1eQnIgWQbZDMdrssSSqNJ3tIpXCnEoAYNev9Id5LCFVaIAUk3u
WoEhczB55/6XnkkVXxFxEAJwIxGX4E8Xe4Uk9pW6GJDEHu9gGE5/rEg2xhRag1NbkFGq3BLBpaOW
trw5yqQqruC42zpUno1RKp+5DE6NxWi+1bKqK3gTTChpEp9sGDU7I5Uec5uQnNDxzk944hoT4dv2
/pK88eqbI3IFmJb6+/YwW+S2NCAnKwwpXOzlA8ZZ9C4cegXZ1dKzv/2F7vCRb+t2lR5nwWFtvIbf
CBPw8E9F7gemO7768L6SVhyRrBUzIHBfQiKb8qvQSUH2Eqn3i4Jx1T2NLjrLz7QEYHCIk5crrLOS
cTu/+d1ejTqf8REJ7dqyNLIBvTzTclB8SC2+tMzuNkVPlbwsdmARXZEQDy52tnimsGOCdEjCscvq
sIh51GObpoa+6UiNGheR3CiTkyyVrumgYU9ZPKSC+CRniDcRNovaSsm0of1zOSo7SL6bw9xmIlR0
jXNa20rjPmi6uaYggexVMd+cguMjnaNMnv5w44O/Io0DnYMlTkJLgOPh8P9VeQE0pDREygN100Qo
m389Ck0GFFpoXJbV8SPVbYYhCnhWxh2VEbvg/qm3AGtSb4WR9ttcJHB1RKhBw+N596iy37FR0GgF
lceJsIwHRYTGgOW+1eGs3SGoFNT31VhuqW2efZgM3xyFmFG/kvMys67yMjHXEKG4ZjSIPJeiwCuY
iBiZ0RyG62yc/+LASw4wOaoz50HK24XY0XzkgZIWJv/s0cbEyD3VeCFRrbNrXMbUUWKqXSQsjxUg
Vz914j5VArjDG/8vWlUt7EwTJ2vg3DK/USrBGfHZgfKD7P8Og8vBC7szMD7rV+pHgY1O9Gza/+Gd
EBEbjG9HuGvHLqHUzJIeL9YlrDC82gLmrEdo26BgGaS4oBdkiyqNgFUy/spEmm5i5sZPTtZcJaIf
iWuGpl/7jomi1uUVNH8XT8lfoyV9etoBSyUoOtFBwuLHjgqicH72MYf6maf1MYujOafXkyZCy3Ug
XO/IP9j2STqChRAxirQRG104S0cAtPfzB+NxFCg0z8SzNmJVUlLIftFmJ8SA6/Ex+8EgkVQD/gZi
ccPfqLKswbAV8Ou6Cj8n+eDq6nI9KIaEelyikSS2Eu45vut6hyOqtGUenAqjSNfK1KPx08scdFdY
UTySsnECq68Ddbg9CIMf98iEFF6HCl3P/rKtlaofDEimBC/T104yi6aCb9Hd31Xem7I+5FtaX+Py
+khAEe1HTZgReQHUvd8EcVHO8CNfPGa8TaB8c5Yzy0VbYady8DqBxnzQ48/eNcWlpQPi+PypVCJ8
Tvntb7p9cXKUvsRG11bUtqxuJJqHSXn5gt51xKwHJNXTwCbwUUmy4SETfzva+2hZq6heTI50UEwc
0UL+SkDBFQu6zYo9jvh/oaD3fQAitg0woRsGPiS7G++J9jjlNJku3yuRxT2FwUuUPBl8vCoPfux/
MjrCHXuB9QuhVZdzCZGSddguBtJxy4VimJeyAnsuxgAQdqNvzCTBw7/op+RVOtObRFI3adoWTShU
uE/RHGiN5gmtfWBqd1IM4wteaxl31zpRYoW+CIfstD9dXrYTvYoKCd7d/YiJy98XqNOv8/pqn51f
I6G5w83HfIpmQhaqlc+i9DbrA0Ad49RUq1VM9oBlAimeudmv+4TSNYJTj1vg1rCfDItAKq7McieI
3ydCI9fd1GXzDMd/jQiFzNx0eHpfRgBll2e20P0i5T+y9bA9tx46iQ2XzzKXDX5yY7C+9IPClbW9
2L+AaPbChGAPT1DNyNuNiOGszbtLAWoybyEmtikTbI+TCM2CXxxgJMaH0ARF3EAliZtooXOG7aPJ
GcVFxiIn9DCbbpgytsk/uEhjtTOsCpLfISxD+ZDoU3HflHbLK5syj7WvP2uCASbpDkTyJ32Hppdn
oqcfAR/FX1jBZE5s3ROtmBBMuWqmjfQO6UbjUm/NSUKkIrxQJWkBSIDAL8WdhdbdR/a+0I1IdNn4
8i0i8XDUBl1GlhUxgfSDdB+ukvl4NscaPQ2QAbqnvUGHDpsAJULWe5/siCkcW7UQwuET/t6Xj5MR
3+f2ApreqIMnr5VFniUth227KTfYKdYxZDT55g1JoIb2zia68b/Xv93qRUodnAKJyICDXtVeq+rd
MIfWF8pd/gamaUJ1DdXwGb63hDLeHqOR2VtCrlcT28LSBj6rWqBCz0bKTwZuR51Qtrg2/Z0HY8Xz
GWcmWEmYQdHK6wnfVVATmgT1i+tC4P7Eah6UypF7HsJxgroeyUms2N7FyY+vRnGdZg1ACPoII4em
ohP+aqvo/6heQrP8gQyhibfKxLCoX30RspBwonqUH8rhdgSK8JWrkRnZ8SqWZ8j5740MGpmyHEHC
B/u1T/tZ59lhXpW0p4FybVZRqJXhhqpX9l36hk8ftjX426olgEBPdY9RxkiBMJ5oWlKn9LS0d+15
r9ta3pOsN5s2LQPtOVFD3OcosjIgxevqxKcA5sZi0ic1wsMWpxAuD/4EFks3L+pC5cpQ19ZtsL9j
bZtOYT1pbY5x/4NpLJYiQdFjLSw4lwaJgShiogKCnd+Dl6WYAGwGzKKkjfKxZfqcq1LIfIHErdqb
e0RQsZz26rvRJIQ6manWQpDhDj5I9qXC3cvwQahjgecUZqSk+izbreVtrjlqaiNS3FPrzkvtKnKC
XEc3QwyvNSgqN1P7TwT/a2pabQ+l6whPCr2e2orgpL9s7K3bmAmgXQXVoIF27D/gS5iaCdxqH3LA
j2A9oWqADYwQ+mCiTRpnAE/6RUFuXaJaN8qUm2qDgysPlL+AxAwJWB0qDYqIk79RkZczfsteN5JY
5sEkpsYSf5L4I1xqDdhYYKsmeGGPjB1uhA5Cowheiy43CblzrC9TaUmjMct0Bn43+kerMCQn+F5Y
yYTTPJZLUX2fe2BW2RsBxBEulCvnN7Xtsj9LVFODMwyzYprTyUQqmWi/yY6EdrE03Q+m2v5tz6r7
2F5eK4LO8kW/SJtByLXrvBRdQ5eke07tDYTzP7T5f2nLBffKqP7p4tWHkQEVXb/4fIt8FYXqhJxE
F22se2g+qjzk0EWV9BbXoEJLZsLU+NK5a+0DzuhvH0SzysDEeDh1o8Qi3Pu+WOtNv6MCEfaj+6IO
wGFJJhn81SSzqWBqg6i54NM4Wn5Sa6jrDFhGnpwnWMJbZMlKpVFSs7ll3pP4XckjoXrrr18jM1ND
1BQHnp7iyMjcJJYAXdqNqXg/kKtgDmSPgt/R9x7ERcLM6NRGGhkfFKUdUNTx/+k9H3aAkuAgugwb
WkjCW98gX+d9o7jMaH4q7DqiLAX0G0aZdxcMMMYSTbVZGCZpNEVE/jV0VgkmjvwlteZF2xJy8coI
alN1hIamm4MBkr3IZM2cGd0poylAK3ETL6kdKpgUDBxl8kt/oOEcFOe1isg4Ki0kRmF+mpzK5iTq
qOxGYjm7wvnSKZS/KA837HVfyn06dR2/vVYGFtl+FrkckuaX47MHzerMvwi7sWU2GiBYn+2w1y7x
T0+GtdxPOTKgQOOEJEFmruVMBS87qdz7PiPdL4CSKkKt38B1MR/RPmauqp+4lwR532zddowY1Tc1
q8CnDT5tma+qMm2EsNArpNrqYFAXLJaG5YwjU8xfHRS+ohCE7Ksl6fX3n1ahYv40niP5ru3GB3kE
lVdTLBVQ4TuJKQ7iMzceeQ0h45rbhWdv9DoKKAnKpZP2rWQYSRcQY0JlyLTs2G8YzP7nfGfiZW//
FJy4daR2XqF0EnYWtdtIs+ilCrey8NGF9w/GPHMhczCez/647hmknnDg/FEZ4hPQUKVHokgSFC/l
oy4A+2utyE2mTvX09+tDROMD9Y0apE+/RROzBwi51F+rusBPQy4Vumcl9eefxDs+StWZ4o7Te3Yp
migbX+ThhcTAvV5DMmKMF+ZzSb79s5IzJJvHqFo9ICT1DxInr9oGZsmNl1Ux31kP9Cv9aIdtps9H
ULXOC8qf9UzfDgoFb67zrmIb8oWekOq35uEA2ycmsEzP2rzvJOLuumPyfnMQwOrFEAyI9xQDo9yI
Po4to8qnz1GvSJ84lz+M+DS69RZfF2ALPx3s2Gpmg8KAQMYx9a7YhotCl0JGKsaFZXsbky/S7TbA
fCRZXnsnp8YNJdFCLNo3szsJpFJf/AIKaeIhy/vaQNkA1DLu6a4GKA4PP3rfkOmVnzGKOuxoCZp3
BSBEDpW83eyVIrTDqhWYqRrnE0tQhbPjSsM7foAzfJa7wPJChfCsg04xcGAu3f/SmQvQk/azocPO
hfJj6xBfQZFbDsCzOoZSVVyg1KqtRgtIXplT3+zRp7rxd7gvQzxBIwNCHlHu33rnzIUKr7BBVTaG
c/S9FBDBdSnBznK5huBSfNyaNZLEyi1gg0VuZ3BJpDc6ewSqq9LznB6Q8pIA3Xhu97YkEdrMkAxB
I8A4tmvB9MjYmUNfWfZ93vZMe823/ghQMz/IaIz9ulnJ2rPX//LqFB61/Mq6MTc8RM0bd5KKMe1/
Q0xHAnyzdSm50dZgLipTmZ617YHQtZqKgMo+SzmbpQuI6zs0WllMtTRtgY5l1Y66Lt2lSoF3lZic
IIii44EN1gMbsAzkdWUZjT4YHP4qHNrIZIbUhRYwztcJ+Rh8oMb3+n8tj+YrRpMJ/LDf7BlS/LQT
SkbVkPUIJUeH5xZx4B+WE2xKwO4choGPichDM0RCqoFvIHN9cnxKC+GYObbqQu5vOeq8N+b9VRKm
RkCLgA5z1nIoicS4VjHxmUq2b8M9ZwBTZnhBXO0hQZh1LmUFf3Y39kGNkpBdVS+XiFlqWPBpgjaA
w0y/N61XfTo7keNIuVueA2spWq6W7KunqQ9sC0SqhL9tWiewlI9wa9UXI8b72D8N72obhOLavlhv
/ow/lvw8O44FkCLk3AxWf1iXLSjvQbQ8zYDxK++O0SP4aNbd89Op3Wo4SU8icXJQ0ENdbDfgPEtj
dcP2NyOP0VIULZeJgqmvkBB5beVeABHMCkv34SDAb5qf6B87CA16m/AScsI9aVMHHbxB7n6tzGDC
y6vyla0jU9Q5soxYQ2tRezEDaj44CQV3ppydlMDtXsaSBZeDHX+QAUc1EuHBEctSp/vWEtJxnTuF
Wf5KjhuENmVChJzsWVKUX7IuexkvR2D44rm/iYc6ebc0LGccKEn8IWFq2uOE2Q0tpxEsLxnInpai
FEre+1BV6yYTKO8n9e0CT1Bwercz3h9fnTVaIGe+WF+7oQaJjY6G4mTe7BYcfXfhNvQTLEGHapHP
RIoaKH2/XkpyEh3TDiA6wEs3y7BHiALaU005QfuaXpFvvC3jVbfNn/dQFpUudsc+O8ueBs+dhYdv
Avv5vieOZem9OilP4rvjWIF4aO2gXK6MADoRYa6rPXidlKkXnCjabRsgOYehNyjZYG8PH12w/rw7
JoUvJlt/kQq6+c5RLgZTJkmNMl3plJX5cXnyY7mt6dLjwKP+surslpEJ82776aBWa2jyx2whDQ21
QtbFd4VigMIbwZ1JMYg4a5Hf8uQvWcVnTQ64K0wC2uAbO5LRY2j1pXrgqt5p6W0QwPEEya859W2L
UT4RJn5fHMGIa/kHvpAXYR1K9qxpy5imi/BU2mUiDCQf0BZu62pOTHYMwBSczHxWz6hl350m5K9B
VM4wCriC22li2k5SN5V0LMVGlo452B842IDQta73E3fCOf1CuOECVfZQTCieT1LZpBNPUPf7H7Q4
SzP2b7XMJzJo/HNDqH9YKQeIGsMIL5ZyXz/zRPnBsU9bL9c5uuBVaSaV2JX42T2VIFOlFD7ZlAv0
YJ9LwROCD39Jpynl+2QWItxBPmgjA7CdpDWXDEvf06sTliXZbP3z5Ap8ZGeSgcq3TDkWZ+f4HkLp
ldVwLRNXNdLN+Qe344Sombw/DPM7hwNbhv1awjiZT2iu8qJmmo9rt8xm1e77+S6rzeMrZG/Sxx8T
w/Qf0ayZ6DodTOCcl1s9/Aph76sR9I9OMtaRrTerTyN4cWUESl7gkGJgiHzRuKuOBPTX2qfJM6Aw
vDWjTeHpwdxIdPeMtelSDSuDDdFyEuEs1QB8cKyvl5afLdMO0I9owbMx/xTrSwknWjFjvJK/O6Rh
3W06rysqo9Jg4nwA2YN/RownSJSUC9KbB/1n+K+MlDoifiLam4L33IOjbB/w8e8hVybRHzpHddWa
662IEyz/194pdjNN+JJmAGwMC0Fn/f1B0lIlq2CxBsHueQ/ocgWcC6kptJ9RcZowyg322xdFTd5T
hXKSttVltZVudUkMH8WS8IRLHwBJClUDcLaNgD8brvVRISMipundukCw0P3GQE/sgfQSJs+ysJiK
L4PiRvZyef6PAumOLiE8HF9af+KYLu5lVT2AXHjr/7JMAn1Idx+N77MxyqoY9FvX+jhUf8xpidx/
+l1Oy/yz2wzNCx8JJBHCKrr6WQSO8mqaR4lmfwFkpJrME/t+615qWHlCDqMzXbm/4reaV7Y38KXf
fcVh3KQuZx08PuGgPelSn6ud41plBhedGuy8T4McFH2Dh1L0iDpIxKTTjK3DMMDJNu9p9es+J8uz
cD8r2fmitV9yYGRRhuSn/NFo62n3n5CXuyKAuL1ScaFMJUYsuzioGKRdpx+gm7LVu0WFzpRenp8+
DSzyNzmKcikWmyP4FC5uAEmr8gu8QX/I24A+q5cEFP7IhOryqamGuOw+T7HUu9ERZn70tFrBF74C
IQc7N/KpvJTpV/RsTdt0Lfg/IKUHNTZsSjaSIL+PDk+OUexsSF8/SiiC3sSHbORuV7FiyvbCdzeI
Czp1pecjuQF9Rmu9Jx5NfWUxlWoh11gHdWexiAywJbSGZARGcciwaThmSsEeYeAQbDu5Ip7Qn/va
b8Y6fxbDJ2U7PwTIB9JEcpKS26V5Tums+aSDF67x3W1DvwlujRSTaho0/Tvj32kXFUrknLNjJu0u
KUn3hSielwDSzqG2awoQxCu6b9rXPW6uKXJZQR7jL3t6i30r4X+Hq5KunFzvFrgdIhDk+JIUQxz8
651jSwNh9GBU3g14C8NKXNmG5SmLPZ3NwNnBM1+/R1qppqNJwqGtIxZBWi35puah+MhArxrOZLsl
ejwrYCUytBSVUY4YdNG48PR+hBNkdieVAm69THwwkzdRs9si0X0kc4TKJXZF24ZNKzvVRPvN+b+w
+NpCvZ84QaLEQZmoDbBZuVfzfbfoLUpF1JzZLeJLXl5S0BxgVaJefw0IWQ0jTDidptlwF+A2iwNP
G69JflyzqyWtIt1cJKt1POZ4SjAhpGmnulihRAf5zuJtoblfcvQkfJWGfxseT/wbVBEXvRiuQcvB
0FjuuFaqeFNHjzk8YKBx7xQ4MXHfBtfXKeqP+gXoDDEEh6e9NLOtmA+ngdJfbHnlbKRjXnN37ZtE
05wBWaz/sSYQIg1Yp3HAksonjDZ06mWAhC+3L3izSlKm1Lb69q5R1hKGX9wClpOybeweSiAQ17js
HRiWx0N4V71qApDi7pRtTxK8hi83rXQRwKQJ8mOnZh8Z7PYUzi8sV3N/SoYOebAI60+U93hbMLNn
Swd9AsygHrXOu9OW6s0lY3v9wzeQUQ/Vie1/v1ucZO/w6hwWW0px1k9mY4veQKnAN4ISpSCgU8MG
Ct5dE4tj/8I54qa7Gy5zb0Hw3U4mYwlBnbdULg0v/dwZgSxJv66XxZtwjMR08uP+Ns6F94q9Kqzy
ZzwmO0eWdcrNJVsa5tKwEE9pZx1Y22Bd/8lZYEIBj2Xow3sfMrabS6wH/JCIWLUc+aYxVynkENLk
nr/pTYmmbXKXcbMI0rpggOxpcaLyJr36lObsPJvyDLSaKYLEHkFN/jOvnFvP9AIAoW3hxGHUbNCJ
vxs0Wi8G4v9KtX7E1MbVIvioR8EzhrYac6WdZAgcnfw39CxBJLC3w9gVWbL+ngHexI9KzWywEYWi
kLC9xN/DD+NHD1RRCVTw2GdKcqUS+89Vcu0YaNKBvRjUKy9lAcqxVfExv+i6/e9xBXWEpDarSFn2
rMI2KS8n+iKYckijwhDk3tqq3oZ2GlWd0o88ubIl8nPXGrrbNpLPkVisINTkBkF7tH2T/eLofSIG
0LD4HWS382UtQUxJgz5AQ4c4CrQpvG3ohvp2axfcMB3G1plZ0RwbI5e/fk8vEJsa7rGRken1GwrZ
mQ5R0yDrrzuUwuruJXzx1znVer3obd+nzaEU2MqVWADbjoqCp9UrW49YeYRJ+78rpHwlpZykaZy2
Rr0FHMx0YMDf75afBFyc5OXKjwRS1jZKJtTtYaorA/AaQWZg2GZa+Bv+scS201wiZWZco8fmwEIG
Nk6ELO5WcaJEMeyQVIy+qsERSQciPs2IW7XrqbNrMIrifEx6ir5jHTVZlmcml053/2Vli0X6WvW3
i+cJ3JyGBYET54zbAKII/iWVFUlZ/kuHU3KQRkEfYF2kEsNyhXDYZkUnXHH7bUnfNSML4pm20+wy
SMgQT9y9MDuXTgaCLMqZ1750FhBDFaqumn+PGGDQLFIV0zE/0dy98XSyMwV6u6lqJvR5v18iqeag
HKJrKfS221wzhJrKXTI2+6H2HByWBZP1pv4oZG4uPbnKzZ2pA+vrbiBfFjFAmvsejD2wibxqodUz
37bcZMAtuSetK7+b3noS6xtxo4Yh/Oi2VbCLKRxIORg8QJcxpvJ0I4NLOglvqOw9DIX5/ypFMPFu
CD671gGpR3elDKhEGgRc1gVClXQi/UGVTyzRC1u7EyEBOS//m2NUrJOAgBdrLs5oJgu8DBYsIZkk
YQmqHR6Q3qb6wOrWAMOGi5pIWcYMVanTGiIL8HmGo6NurC8xoMSaaybT3IoFsOr860XM10boyvbI
AF1W6im74dY/+MKYp8uDwy141k7TtTI0jdUyKoN2/qUBeIFrfBb5S7EHwMpkeqBpMINKrjhzy5zN
GHe2xW6cP72HJsb210yLjAogciRio3QKUWZYoiq5HY6Ys1oMc8bbYyS3RIL6daLOdl6LaC/T3Gpv
exh08dtz2fgoLO8s0mtiv/erb/xuW7EOL50SrH0uBWOc0oSpGFavTojb9qljuIGcmOddu7JkLExN
oaPzgSDchrq6lqcOqJPBGgEI0EeNIEXDKlWaWfT6dbq+fAbhzpWMM8Y+mpkMk02GbF9zUsChp/BA
r8uT6NB6M3KK6S40bQTm8KFb4twel8ynqm+3p50XqRIal3pOnpX5awGtp8MuELK2b+YN/4a2yDay
TNZ/r3XHQ0VTVgsIUc447TMY9rxxZMVOCl5RoXDoDWe2ZuNUDRbBlRnC9mTYAGZsmcDTcg80OllV
+Qm9hlMZ7XJ5PqiaPOzpNpY/zlsW49yezqS6WEc2X6UyJQJW0uxXGVM1i40WIIl9sFd+KXG2oopj
eJTFE+R/5JoPRY6BXrHh0McFA9RVIWI5SeOXD79uvmL/Ccu0RhqJtzCcgqg0z89yDBHhHWlP6gLG
am5BRfeMNldAZqN/ChXSWnjtxJ+/jK1q4pc35vZQmEjo5a0qI/MwKfAh9Sao0xIzvLTLwW/KcuFW
br8li5stTsCQl/w7j8ci/8uLmw2GSgYBw0kxxhMrhHSROWKYdS9zjwm1MVBzm/mFOanRGiANH3++
TZntoFXlVTBA9igEMcRbOFcEvsFBnvfi0fO7Dkv5e01mi38iKSXBkOXjX8V4/1jbrWOm2l+Wu7F8
gtencvAuOBZaeWdqBC/dvXpZKrUxKjaX13iZYfyWFeDF1iIDWH1NsX453n4ybs+1sC2Sw8ON+TsV
GC7dV2D5mkhTcr8qRGm6LcCCz8RZR4Ai1Yt8istH8OyKJeOTbsEI/77BbFPrfCVowPgMLV3vXssy
bYDG9Q5BBEUvQbFoPogp4QQv7oM2XvAXPd3aaTI81Y5+Za1+i8Wl5SoK/j4470e2ONcESFEOK7oW
NUyghzvh/jmTsQ3sJ2H4YRartfi6iuoXGUh44F6tfE3yzhg256Uhp1W9UP+clxB6iEwCwv8QZ/fx
hmmHb/vtB+dUN/z+XGeX6KO6IfrgjJh0+m/i5mtXwm9v+nyR8JZonMRRkf8vqM89Alm91Gtkg/L6
NlbncomBezOsg9j0f4lftvYiMzYZmk64a4r3rL6j/cuf9KP0GQRXIw5Bk3e0AI33wrvlepZAa5Id
4FoNsVqf2IPK/4cBCiPkEMT65rTLxTpKrG0NbvBhisGc5jeZ8bw0ACRmT27dv4Q7J7e1adEmQ0gS
hNBVjOnk78jNwQC1MbSrV2hXBLawoRY3MywOW/tBJaZJ+zDBfwG1cVJLbOQDK+6KHdVtxK0ZnuK/
21VyY8/30DV8V9uK7eWRhWtOFKYA8Vb6YHmtBN1BTdWrv6BbzwtNUEUvp/K0mg4Uvcamfh1+reGb
xLZhPMR1TLcBh4IrUzcwWoXIjVhFjqjiOLY4bW4LTgqAupy0xtawPQmAznj1l5/HHzo/imPwec0H
RH4eHzuYm4toeH8Tip+JUQ6bTP+s+SlhZH4Btl60/AW1QLa7BkrmpmSRCtY74Y9K5p8o9ltaHPz7
VGrOZP/lNpHb8C1sOIRa/JB/Xn4MbK8V1eiY7v4pCh7zKRSgX/j21mXopqHGA5X+kVOgn2qNxsmE
EZjuuj6UEvLEdw2NQcUYwDqoQZL4qDmrSH4SFlcagCJT6O4eEYLadqAxMO8Ev6mdmLfNfAncPfra
5nMDS3a9zBJbfSBOKLqF2vrK5/zSOPtbP3myJQReJQFvm8cSrltjcoqkPzWzXhdmHhV5LfZCUVrP
azmCDyawJgsLPOBwCkir93zvwEICQqHsH/jfFtTbTq8CSSp/GrSXazhEqrr94AumIJczIsh9MzH9
vJuqii45Z2eqk1Z0o9LW2PfQ98d3rW/0GXC4ja1ywUw0K8VKdJYNcywBAl/RX32dMj5Ju7sanNi9
rvxVjkR5SD72Hpvx+XKROlQhUwLJqJWBeahkCEaKVj61CBM/vECEAMBAFUhVVw3GrI+/aMpluZk3
66ENtD9e7lgklE17bIbhnTX6T+ex+/Reh72FqSluqINLf5bx6nLDteSYggTmpGCb90fbvIqhiUpk
7Hc2/skD6+y6s6XqdXPcjmiSmXUiL76jiO7z10ap5we3is62F4RyNgExkN7ifxLx32eZdiqiutBc
sywnRtHI0RVRJj+wUzTOpo/ROTQkAv8l7g4sP6eZvFIfaJcEWIyVIp4R3EGvwwAD52hIJ1SfSvLu
JmtckpfIpyDZQBgbj3myJQPT6WaJZjr9Y62qjABhwU48sMMYEYFSyoAsvXjFsPuErqiH1U/lUYnL
v406+6APwNsxHn13zCaeFszJZmHxDyEsD0b7CxHUmgkWe0ESQO7CM5E/2ieybyvPaCGG+9v/0402
qNUc9ONX+HChm0pkZo4EpnCsiiJkSCDySdrIHCDWaKZwsA+OcvJ6BILODOFsIUaAMiYQeY5IMVqF
/MEp9zJdH0WY+8OVKUEj3EMJJNKViHenxoNZbQs0jgGfju5Z0vQofEj/HqXbKM3N4R2Etbal7dCF
GEB72Uc9oSkSK+NhzH904VlU4URHjiQhDUsGQL0vbBbgZgWPgvvy5lC91lhd4GpHN/CBt1kOpaML
LmAU3Oy/Zho1X2KMF/QkNxQPbZb9hZy15/rK+045P2zhED3OjosBwtnpxrzX7kfDHq/4gK5FLPFg
sI0Lm+mSxwUh1Z3FDwY5OZH1Ex2pqSKaajOnFnbzD3JlDri6TMHcqFGzI7lNVkdmDIyYPzlpt1Se
ZDQYvT/iXX3vDPKcCpvou6oofOcBNqoA9FsVL4432OJlVgluj61Sb6Pr/sZ3ngZltgs9/d/dCYZ+
I5UHm+T3WKT7YOPwdrjlqkx5XAiTzSbt1jDmahr5mKFLQFCmJM2Akylf4O2y7m/agYW6Mr56Bygj
IePVT0SZplWmFVJx9VRdcmcfhpApk2srvT2t0i99y8JtbR1J5SZB6cASwCYH68IHp/q0zrTSy11P
20+A2e2a+8eHT/bRhWZz7xJpgUhjnFmKuX2ukVO7+zADyDPBfxHQ6wLvShjfQrR+NNmNS/ngTnie
1QhtZLiHRrfqV2YQyZcKPvMAH58/pmJGajxqthjTp45ldkADpoJh19xJOxLHKcYEHzuDLvDw2WnV
zDAdwXqVdaZFGXEB4FdLVKwed1xVa72V1kRl+BqGacr8kRYWneYFJ899SfPRcarAFVA2giReyiAA
kjXGIb1H0OX1jL4ZpmKBxkQT6NT1DcUvU3wm9dRgxCQRt+0b+42RbXkAvyiu0cLLd8xO3Wgwx+jK
cVJVUBvLA61l/DXexbPLCJxYrSKFeHX9Y4p42DHrZllDB2UIFZ+r4SIUTyk2gAI8OvrJzJtigwpF
YKie6aZ3qE6Ib8XCSnc+Cnt60sh5lmUJRgTx8nJIknlSX0xbdhBGuiwmq25x+eDmbIjSGQReAaWH
E0wPETPB5j2mcHseBuG4c6zTlo4+HxrZ7J54fAtxK+0arq84Wt+z7DC9GhyR/tHeU8uPMBmRWAFT
OqEldOGaLSMfcZ8kRrf+xZM/QEq9OxsSMAIcUzk0Hc2ugVoLZv/VMTf2eBHuH9luTFWhT3b12Ilw
U6BSBlvwAwNNmpEjPOwjcnCK1BvaT3VK/QS6Fi9BG3cmOKieMM+GjnmNOHuQJCVIG+eslO1WBKCN
jzZTXBt7XRZ77bfXAG8QpEwJDXL2zGF3GN6Wq7s+FeZ/HmKUc94zvxrGgl0KoXSLymow1EL2RJ6n
iKeS7b6r9Lq7ihxb2GR7FLNVFXcfg1mJNgNH9VdZmcnBYyV/SlndJXlH8aTD79Ioqh4HAiG/3Fs1
MuvvmhsCy6d/qkeO3v0hOjNUxRr5WMITmjU+zn1++pSSmqIuWlyItvW2Jpts+5aAYn/Vxcv4YoYT
s3o0KGqbNVqOPh3FJgkxTEymZnPLhIFj1SXVPsAF96NeWaEf/8JHGnpPDh/Oo1YrDybBzjp7DGFQ
JstT/sfxM56mVcY5zBwBEY1bdLv+jVIBafJPtEJzJGWGVYml4crj0R2Xf1hVUMPJbOYZZBI6KCCp
aAn0hwzKy2KM7Bh460QLZSlk8PvEGhjIG1vn6lGGo4iHK8c30yJc+uf2t9ZvEZvk6RBJcv+9+l3J
J1P7rmhAao2bAC4v4bF1kvFTFHYHqCwvuBcy0JBIC9U3BPpwtgdiah4j4Eo1YxgHBEewtR82gxZm
uE1dU3QTU1boxOEDAZ/abfpXhyCIIcKOHRErfwYiIa/nGNu+HHYx3lSyokjSgBgrXsJFDg7pH/ti
y70XsNvRcRd2xmjT6NarPtORx36L0NSwGE7geyM7zXDxn9kRWB/gzzQRMeeuOWmTCP2bGkrfhPrB
pJLx09qjUOupphp0Ew4dkSHUwusgouWAaY8h0KKX8FUnFgSxINmBx4KctMq6mc5+Fz3ZXXsHg97N
8qmvo/xAWJ/O/tsvUDHDMEPgJjlgzYZOtF+3I8ktZQoQrPhIImhkpGveYNLLV+4Cur56wNqJ3SKJ
z3ThxWdt67lrytpkBB3UVOi3uc1sWEExGd937WMCdNFy8jMATDKu1xhdgc034qNN4F6sIl6zQYgk
AAQp4I0CbBcUPHMSJ7paD02b3n1iRS04ZS2ftGE3zSZNsH+gz1X8oub7LC2Fspppo57Z8OU70mWs
Hpmts3gjSF0DjsHVgK+8tbIwNvww/hDxYeNM8Ws2qhLQ9DuvpwyMxHTP5KK7d7O9StGWp8HoGJ+J
PnW/1LLze1zViCwK7yQh+EAKE2RUSME5el88s25jUsXujKnzrpfPQhXI+8TQijAHyKJLMU+TqKfc
ike7MOY1jBAVrW5uXZ6rl4CQGPaXe9vruY6r/xQwgkOr6qcjWnGlz+8+o6BLAfHW3FBcvEKs3/4G
7fp2B9+PGycIEwhLX0yPzzV6hE0tfVOHwIm8cwI3sa9mcjdMLorq0uqMPUjY6tJH8SbdVEj7ZYU0
qfJeLamD9cZkM7smvEeZ8lFpqenrbkz49DpT40ULxc8CJPE41hWifTjlKjPMyOAr/lvEfUDfu/xq
OJ1M9z8SQucE6xWTqbpMKzxDIhh9udhjvKzxR1ca8Bp0ZlOdws7tMfQv8eZY+IowPYHY0f1J++/X
mbK1lFo5nXu5+n3xHlZVDBsLfD81pkt3bsmlE7RVFPthhMAgb0roh098Ywa4HdQzH2edmsxReDxF
i4iSezg/5C7TyBgr8ueCDCBm4d5iR0FrqTzhQ/1CDFyEVIcaW6J5HL9I/gLgXeM+L+QdAhuLqrX4
ppMKpJ1aW8rK7HHYsGBgMkOdwVRwuVNepD8Q7yRmeQ8ZlZeCJL1RM3tU9C0z4uO9zH7u5bN+gxMS
8qrv0rNvAjstHwfuzZuP7YL4DAYb6adBAA7HHEPqG6n6wZMq6q+KnRLT8nJ9iLWPx+MNgztVAV1i
sab9+Qv3h8+OoQHo9fHiNT+n93/2KKTfTck9T9Pua1hKgmt7Wup/WXG52D1CElvCP0g4NoEIbZWm
LjzZ0qjtX8Y1t8ryIHl9Xrod4YXr2GatNblHkjV8oHIsZXKHVbNSNoVxIP5LfyXz9BS/DBHHX+KI
iy5ZE6YpkeTLrWNoRDFh49VrJHEnvF0dyQiAGEwgk0a4mCg8JXe2F0lWSM9g1pzWAMalIV0xtMmT
WvKTUP199iVYVxuoDddLns+cEPmtJU9Pwq8TY5ikJyZanRWZXAIDotKvyXs+950Ts5so9RwaCISv
Zdmw0oWByH55u7s76W2zGjJGl4lCnWFnR54WSc6gMQm6lNYE3qOiwZTSA6vT8DbDkHS5XF2lOFPp
WgwKr0BVAiIMnFZs23gHLUBPTgX/WQLLE4HxBbj33gIzdsSdqhlsZvsgDKru5G6VadLgCXrR6UEy
L/GeJBoG15uV5WWRPxF30qAoZvN7iOFdGbnIQj0am4hFkBtvpufdqNuJZoXc7Bi1oeAJGhA9sekH
1qtTxq2OzeDcuypWdIrSBFKawUU/vlxuIZt/3sEK4S8ergnooZCcUB1WqcbWOndAmjJ0OYx2C9N7
9Y6KaFV7EkAdou3Zqdw8j9zNuGrVqzvXQdYX4MAVjj3IhhfWKHp96wF5Ws3rl+S7wKTcRnSWdm4m
GgWf7wHGOARkH7zoQ3P3qR/sphTGpeWszxci/RxvbZG8YOu/pJVbie/MPMT6UVGpfCvMSJ7utF7J
NNA/2Cj2CEzsCD9TrjqoQ8770QelYGvnkMBebJv2uB/rxXcy67nzJ8UWzQ6KP4ditF2i/SF6aEPt
Yuv+6EihEVfjt0dv0W3862nbbRS13jUSuQ2V+Jrs0XSbtwflW6Zmz+2jmC4HyyuSQDI5h6JkobJF
ZUlaBkgUtP89tJ4GZ8mVTnQpJJRDft35u6/sLyGR/r9v5uSPQpxeGo3Ymi3rk8htX4LjrMEnc4Bp
u7zYfd+TrPweWlRptDZFmgq1SzlrI0Qr1BUatO1s7wInVbb34GhoxB4i4cmyfsk3hs5SlrbzSsZ/
ZfVFaQAprEzC0q6S7dShx2Ar/nhsvYtvLaIuzQ6H4+TzHOvoW40j4Ya8WgiTbgmI67046j29k/hf
+gXNS+3oMYGEb8Kcb8Ib1Qyk5PiLsBhLKfCswfovgtemerXBPPi6aQ2bcY15Ylt9H5ti7vzfq1Jz
nGPnWum3vpdXj/5ZywqOgPZc9DRSC4NXoNpjkXlWuOH0eEPZPmJpaVPlbzfmwRTCTrTo46y/XbY2
OJoRsY5vs7L561HNfMoAXGCma9VZfPefQrsEQIaUwUwXECOmPEyEiQgQwBPINgXMul8860Q86b6D
Q9ObR066yKMkXxF0xaz/YKAVVqddStGec6H3sr9A//PaTJOl6d0HwJPKP9+RhaImsXXd8vZFDgpa
5hE9mXWCAv4oc4ZTL0vit59gZWBT7IqBG1ObiuxNz6oC+/j1kJW8+3gFapqQE4LQrt7nzR9xrABJ
EFYNyvwhHoBYf1Igv4DNTd3c/aHuIh71sFsN1l3Z/B1WO/IrYmKrpJfxSzDDQ8ERFasEE0VXfsoJ
rJ90D49di1UPAZIu3tr08iSLUpnMWT7/pGGaNQ9FbQij0xCN2MCqZKajnwaNZbAEWw6bArvYlffh
AKI0+r2LRtFhLXha16eS7acTM8U53n7UvF1obAfKYO3340yP9D7502P3Ua8OKmNeL8Ljd+K54IS7
6wY78dK3CyUS3+k7b5GOV238t7or9P0vrM5Ojg1KG8Uwye/CD4XPsfTL/7Zfo3zgP85UU0lMQBKv
5XPrSjwtnHv60WhE3VcQIa0iHq062/aooT6ebPA6LKzNZ0rpTu4oLvs+juz8NI3ztBYayyl5DKjF
T4r/8LhnA7TVEi48LIzZIjD8pZZg+0Why9DB5KP+7JsEW3Y/ju2J3Ng8G+XzTnSSH/P9I+AeiPMt
4Qtj8x7Haw0QtpYxAk7ULMG4zI8SRSGzNg8Muu/wOK4WoQcHT5bYLn5xp5z4TYqhA9MQrgWGG+4W
XhYbHtDqjBZAwelt9LSqsGQZHlcpyDL2EMt0gM7+CVegmz+x+ZLE6rvMKPXZYj5hMWlvy8Xahonz
Jl1+zT290LBW/Irs+M/San6EC65p+1I+TrYlDAWNB3EriO+yDjF6gngtAQ40tvglu5z/mC07bxnm
lAs7oSZt48uaEiOfEhNMnEv5ai6LyFzZoBnAshfv+DCGlTo9qHEOC67SggoJZl6BHz7g7pfWgGev
t8ZVx+4og8Y5Qv7olkx6bsUY0Eb/xkMq8nlUW86bvsVVgAql3xQy4+Mdp6IOq5Y1yM84R/1edVI2
zUKWwkQKLLODZeBT9dCiXTLNn+xi7awjFh0HNaXXG4BtzWATPWvig2wrks6gjMz4QEh9FfwbHSZw
SfV0q9ZGw1qQBMpg2Zwkh0g9a3aIGPeb5Q3UBYMqz2raaCCVDSUfL4y15x94+WtrkTo3lgSIXMcF
C/0L66DlFPNt/YjOugXi0r3qE47aHVoQD0+X1OHTqTFBB+6dt/ahZFAROGBrQlJ0eiFs1Jgr89KX
IsGAoe5Kyl96aDCP84OUkOsoxtv+fR9WsO4Peb1EQvwM/yZCnUL00xu3R3tVpgJ/AL5Q7bx+PvcQ
A1p/QxBbHkhdlVx4GADgjhJVuAoD43kybVi8uBE5L0VDWUjku47fJ/XmT1bFfyTfDYlVgXlqJ0/U
wKzJ6HUGOsksrQ+CfseTXj7Gx0MaKwKloHVs0KSp29quJGsVxMIGmI3VdTArsQvxxF3xdheBQ+WU
jMMNgi0wunWgFQFp9YQctH15qw1/e1X0PoYNP+PGl/+RetnY8q3s+Nv7mRzNq8zCHuQ/rvZUnf2N
LhQDBEYiHJ9puuDCTiYPqbzocEp4JsVON9oi0ywq+zFfcRHrWpunDSWgzSQ6i3IzAWESrYm7iE/O
pkksm3pnq/74YedXqCfXSJXCiKgrNK0gOP8YQAKtdOVEFL9Xw0L0zT/oTI2xgIRWb3ijmpB4qmnc
dR0uQ8sPo1KMOEnV8uQTOqyTfurOykAHhnPnt7GLxQ+RCLKpgwKCGZ6viNavN2r0Vw5ZQXP/SeJQ
5b2KqOuLgJ3CTWmmRDx980jIPH6KY25bMj0vm0AF34jRGwi3t4GLmbYJb6BhHnSqqLThDyPUOvn1
Atrd9c/QabaWJOGfH0CzfeSUrZak/Pp99+lbDxMQUY3+0QAYp36qWl2xaf+FU6xtp8bCDmnqzPqo
HuXZovK86nYArYu4uYRSk/5M9klrcEfegVpw88P57J6/5e9HmUw+CGorgW7fJY5lvuf9FyRiDeDJ
jMIP1rdTzeSuaWolq07om/I0huIHyOn00hydOukaPHi8S2C668DvsAaGNX8iWL7rmToS8L9uzjY4
5tB9jCLoLg+0qQeeNAJx34CxwhJ/s9ttj5aO3FvWGgq5JvukdWkmFA7F8Par/pze4OQv4n8pQb08
6Pyq2bFO/xODkT8fogGSAQ/RYpacaRfjQ2HLgomL5GaGlGCngxxgIOhfPojMXUyE9C111GnZZng8
SanRcDPCIjv1CGHLndCTDzLgtn9TS6JkxQDxyiIUYni0QGcqDOhpC5Z7jY+j82IiF47BLrYOfKEl
4+XiVT2vYlW9/aWZm3vSJyCUQHzfYvC4IktVrJ1AluQ0nqAJclqTTj0iUN+tDrNAov0Ct6eQO470
jrfG0KfNIrqoZfc8Tst8Gz8p8LWJ8izw3ee5pC1COdZPnDXXneKels3rZIrmUOrKLC2J8Ip30tdf
5wgPSfJ+zXG6On6FyJxZmzF8x9Mbg4kR3Kg/yJYhuqrRW+zt0PSxPFqkbsuPpHEJj9Q9jSCkPUY2
6wpJhVMCtnTV1OYYJ0MPkunSj2z2vzsgFLttm9G3h6b9q+ItgP+L7MDpVLOVJAJsk9VRDuXvl6Mc
j1tbe6UioO2LkjJpEabfAq/V/u17ndWtG0N/x3tbqYH7YlQmes7tyiDtfrTlJQnNCveyvEVXHjL8
ziXlBkafEnBT6IoEG5nYsRS21l4+1sgpTXEMHO+Cjz+gJXe5BG/huQNgtduXlvpqq34hWR0rHPZT
jaVLi16wKidNU/2htGqspAiTSL7oZ7r7ED2GZZtqkLIcsiL0GGgMWtM7QuwAOQZrLIImWsX7aMbW
nuiGYY5KP6j+BQbUYC9TMI00EDSfZcY8DuqLMy+bjm8EDaAHJndI2TI6o6CaR/IeF7At14KnU/IO
4sQom5J87qJdMOaCbblNNiMU9q4f/PexG28CR1DuInt68XOqQvmlvxcsa1G1pk6/bTNdwzq5XWL9
1z8p2XaoRZUvIAKMV8VwCHZLCyZNLtBptcO/vKon+Af2qVqYO9yKi+6Q+10/XfMO/5YH9c0rpMCd
aHBvBr9ONckHCmXSo1rLv+3sRwdDMAhJB/89rH5SQF2N3jAjoRnTF5iyT+MdSNkwKeoVnYhEuxyO
WWTGbXko0ZXIeN3b57QDVCo76FvRFP07ds4vR6enRnAEj/v6912qkXSrtgPj3JjMOVai+TnLM0LE
0uz5KXXPTuA1cbyEkJ5rWy5PD9o83S0sPa9ZprITsjzyOvgzzB9uK/VGIpdjMFJhBaAKbOpTOIBT
nSa5dP4OCB3OE47VyfgKJCEEjkF4cbhtXm886XdmIA+IiU90Zh48b+iki2pT+/f69V9nQ3gtV0DW
WYIXWIPh/uykgATRV70nBK9MQKRXWoz04P1nrkb4oVceWhIQQV8nmcvsMfjOlXX6iUPUtD0p4fPP
izPBtgtxjUaReB05gOSHnzU9IsEopDUT51MhmUzOmZoU+0duPc5rzhgd1VCmZhw5e4ae02CQwiAy
x8dTOQmDtoTccqWd/LMjZKVmWmzGZlO9dgrpvPjEM2VoluPpKziDOWa9CFFjarcWUb5eQtsM6xY7
e9Hs8o7NPgiz8zcymKx3XwmNvKU6+y3m/AJn5r47HXWDvOy5lzdu4uDV9wzdgBbxXTBMHs63qORp
CktAPjsBRYNmF8oHwVkEfeLFRhBhhFUlE/OqeOqQOjCwP5oCQNkOet+1Zyn8vXEl4wa5XlyuNYm+
UXUOmHzGXYUcMVQoMJTv0hAs3BlYOXr2EeRnsWXJkfUTvpoWw4xxOoNjmr/SGYpg4Ac8Q6d9MuKl
qrgS9CacsnlhlTtFbaE14ad6WwIDfMmNlP/n3w3ZvQWrAwlTZOzOCFB/OLa2qgK0unQ9ymniyrIR
iHZVbES+dxjp6PZ3zUUaWWQ523nFWYLdF8YYB2slZ/UDLvxiEUztWXf186ikteOoDNUIodMKgQu+
jzW7X8pqd2hytCMjtMNxIPmXG1Kwsdf6efQZqnMXW0c3wCUmEc0sgo0YVMyrBG7cujz2N4wxjpSA
SWp0NRQNA0tKL+56avXnB/dnbcJ0Evo57ARJ9oBNyjvfXe4sOKSju0lk59PvJPu7WyCffhb4hGdt
mhc7mf0zsYbY1CrJNGSVt2of7Oe95cuJjzqqOre54dQGxloohhizakRy4UtP45Btmxx7ob00FNw5
7k3iClj2TaYnTC8DAph7rapS379AsPY/EfByjHJaqCbu/Oi6xdrU+c79se6tsOBryu4VumKV9CRj
cShFs4nj6phRUccLFa40JFSjaSQLoex/bw9YZ/0SiA5baI7DQwRW6rFDSulyrlygpvcIncGMkylj
MYCOS1mBUAE01t79DVtekYRN5cPyy0ShQePUaOJL55y4mwr/Z0fh9H1m14jI1TA3Cf+L9WbxwGet
EdDXzNCSKsWPx6Pod4hGwqBq178kOpm632xge0DXo4BGSerxyReOxzZ79dT1fBEDmFcYj+Q4ss8S
XZkE7lPrvJjeUZmPzlDSPAwiLdMwzWIxdEItKGatzUF8ogNelAt3d8nOgxfRGiaPb4fcGizkWoFZ
idxEZdOZkeq32tA1UlHphGYjWxn5WZY6lLxh6tcvnJff7biCWn5bNa0627GNWg9DBzLtn/BHfaPz
vJtSw03jQAVA33j598sFziyLtzPpci0pV2ptDTAHiUjiiPmhp2wJlEtDrYapoXK/Og6l7V5f6pFB
xEuP7nYGA/uzC2YzJ1rCp3M6cZaEnfxzbgoz8/CP8+nwOGzNCUJ1weXUtg/W7SQgWl1z13scE6IG
ZheLPJzTUkBwz5QtcIvKOtX5YXzL6mRjUNksQzRkbv71QRR611u58BxhR3G6GhqKMY/I1ifaU1Qh
5IkAbH9G0HkibP0yV8gkFe60trW6M/EkMiWyMBD4yOyRWJFuhPbJz9x/VchGrPiRmbOuJSJ+V88l
KN7W2zSZ14Pd6I+v9Lw8OWqrk7CxuzUiJHbkUvKZlWzFE/5Ps+xYW2c+enqMeEt8fqaAHAtBDUxd
7NRiMrHgUbOwJC68viOeZiEqYZoHmxoeC2XVGVkfQ0P7UrFyENhtxko79BkySXBnQQroNZ5FwCvL
BoqZF5W1mCwhiNK2EfffbVUOZClyrwNU1xoeiIihkEtpf2b0OU8pXNk39i3yQPW8gnazzRQ8sdVJ
wVoGCHP+G8jDLuS484TbUtICd7nHbPbq6x7O6ZZcBfXcwu4Fd/OrvNj8Si9CQRijsadI/JRIxUJQ
HECq0914gwgpxcyj5g/MB7URlCCxE48b8XghrPKSEt08Lx+KeKLv3OfhBNA5IVJpY4dswxFdA2Cp
RE+IE3NTq63jzn7Z5/Mcaj0hFIWXmXSMbdx6kOVBspzobQhl6HiZ5DU/E2llytQPUCid2URRGaIY
0XOVL5BqQ4qjBl84MdVGwvgKTrT54/M6lfq2a1svi9FJ77nv36qk9mY8XJ9tprpwed1GAXr9Mwv2
w+H6UFa9yJ/4dUlPUGcOKjFG+JgHdD4ffiMhXE6oKSIA7I9KzXLKvTqKcKdAIl8eUUhWenMf5dIH
/4k4qpoMGSMxYEJYtRM+VYYw8Bnb5E1W9CptRoNVKAGFDeSxk8HdywPXwZXaT9hU/17RfJf2uzty
FConABKyVEByQkFGUphVimXNO3qFKYQkesUedM3/sMjGgUUx4LQKmaf98MOloVhZXKl2qST+AxUe
NxKEMo/w5wmAiy6/Ur8dKQhMbLwO1AaDeFCtgNLph5lMdbyOhIs/As1LHJyMGXSrWeCMPHp6fZtB
vtdFUj0hN+IDiuInMGedDg4Vq+Q6dpbG9KJMf8ZRjG8+TJifk4f04DZWcUxp2aIE1Lscs07BfCzf
JsFbaEAzF4xt7UXLvG+BAMvAPzgFZW3ERmMW2ZvO2Bd6u23MdMqZ7fSXDCsDNcBX8rqDKKav6s17
fU1Itp4IjGVK5iBljRspUUrEIODo77lZfuwkUlr407Stf8iChgYTYmSanBQPP/DW082wH4IbvsgT
eIjdrxv1Rjwg1/Tpmm++h/XZztHpO/bqxo0F36aE7tvWzK/aUISOno3tzb3yntefN3MZI3Vdiw1V
mXR73V+Kihi+NHDgqQXOM0MvdkJyAZP5RDLhUr5GTQD8VneNjLuCDCQ07yBXEYrwfTOBNaM4EP5q
kfF4gLJGol9v+9B2TE3DRcOPHauWa6x2zi2WpW465eyrxsVnGwoWWwl2VDOy/OOUyidoF+CkFacI
Tmaq9z3BgGkWdE4AxWIHMoeH9aROUe2Wlh0Qvrhyq/AQ/xgObmrL8QYNm8HbbNEiCaSanNhVD2Oe
c1L+c1whDxZmM7WaztMvSP3vuD1t5Oj0oByMuV6wFjIp36c/jWhdOEr0PdPg1VVCy9eIgDIUlL1v
ogGiKwkcjpD2s74XZMhpsc7lLEfvPzHpx3GwFhHOI3EffbjLbD+KzwGzS8mPjxdaCgq5EDIkyiSw
glXVUVixvlCg5AVYsHCuCjTITv4WxN0L8nsz7fX29q6xFSAb+7Aenj5Re56b0EISwU1A5FtjPlpd
QrFW9y5VT6ziENdBQhNOkAlUgP9chTnnRqbtlBCVmezEq8iSK7O8vDb6lstZ7BfyM/5AvpD+4pOi
y3QHvTnuH1e690yoyrOn9IhpvD/VCi8lQ7ZnULk7K5wkDKlSanaDrpGKrUhAjXqqgqUUQAMdhqQw
VFaG6OW4i0Jn/j9y/jzzKrR0M07kiQRIhkrUIg19coRSE/k76FnSFnL3iYpVTRuZCw4dlAkDOcPr
+6sUB3RWHnSzdMXrmzPWaaI6xaQTfk2AZVPW7k4TLQHAyR9QPi3PmTi8kL/GrF74Vvn9pmpMHgPs
tPyPH1KRm0wIB9wumnKeK9wxE7hV/ij7ljpiBiXCjrcwYXU1dGIvh8Liqy8UpJiXCkcridUGwzQv
DjlCW2jKkEFT3/Yp4iELpNk1el66QvgTj6aaKXnEqmUvF/KQaaQI1wuSHvyF6E6tJWkGmnJbiLb/
ORuGm+k3rvQJJmSG/gbDBvlrE7uIs9GCCpMLmTpxnSUTkaZ0/2FFqAu0qJIYIbnb+ONdJyjwAtgW
7BL3SxEjWg/GVeRDRfeFHsKBghLoCXLGAUaDOdGJHflzghB48I5n1ruARCZg649e6wwzcvGGiIvR
QHKS2qoWK30QRg3N2jsz0psontCARodUQeav7DKKY2LLWQbuyfVW8NnjbEfe9+OFEPi3mrRRv3cJ
cJkAZ+qR9MDi8QR3GUsAON+wQipeg5rcUSPxZ0Tvhbctl0A7SO61mrlJWww2m6rdHU2jUvb7PzK+
Ow8AxNwBFQw8wTDYoeoxCii8ZUAiXIWTI7A/FQrIigcsuMv+Bpkckp2s68DDcphG3goUIB+zi6yG
Sx0kDkEkippLzetCkv4cptPygtRunS8aAFOTerOTatkxhTpymVLFQJXsg5B7USvyqu0WYE6TMlpG
U7XS2+0SB4u0N/guSOJpIGw/J7VMWNefC2wRapFQXW9o/Il+LBesnZoeFmLCxu8BiRvg8D/1vyUo
31RurOggZ3GnhA6R1X/I251vEEJCpyXQk1X22RX8LFlWvkMrMaX/eqahLDrkVrtp16lWdBKqtB+R
5bQ+B5HF8EltZQKt1mZpbehGWM1RzUWZ7IruExr8vJPfkaXUch+h6yh8ZhhhB5zVCB08cHcLWp5c
PYGJ9vfHY1SlFo48pkqnTKx5W5jXijPMSSD3m2FbOulPPhpgH0HgSceeDc06ti2Iu82SB44DVhSZ
W2IRHhk4vcm0no3hjV9g25K7W5+Z7xGc2IETE/2W/rAs5SnZC8eNt/wDqIUaNk4QbqbxJR+2mmYj
n1KxGmdRR8VhzwciTYB8waJSxbi2TV4a3w2AGTnFQcUb4+JXrKhKoTM/EKq8qhufyXYQzA98eCuI
SrXww9pthSpItUQMfB0ssTZqiXAwAc9AAasidpN3v2Nv91iQnUnOWzfzvDqXFK3gltwIV1aIOi12
rO1v1CdJeAJ938o27SZkMrTjUadLzf1oFIpfDFOmXuji42IZRhLG/8MNpgKVA1rBOxT9Hvn8qjka
myvq7xAzbXED1DVjreCBnjCH4Ls7MzVWP8itm9AFoL98tSrrOZ5T4YiwgSPOlQyZM4ra1Py6hZaQ
3+dMsAj/FoGV3uF3eznShM/tTSiZzQS8tNF0mJVqlran4YkvBCB3QdLFg93Mvn5GfwEboWhrN9hg
/AgqTuzb6SHuEoqXbBDU7EnIo18ivs54ErOsRwNDFcTXejXhCyH4sjFFDbQ6iWxNB4c1QYnknz9U
tfE51h8+QSzAgist59d2alc5smBoPC2d7CUzXf+yCd76PWBSQ407GlGBkY7sXwEuuiILeAbg7qxR
yuNRu4MKhS7ei5Vm88xKecFH+QJC+ctkIF0HVJ2QjGb8kM/xq9j813oJemcXu2c3YP0u2G6QJRsb
pguIpdK1i/TQhhE20VVbh6bAq4xZOY35SKvvE1MJAewZ6UqO7AaeGW9I8vDw6WgkRmMsWy82tNuN
WXdxwYteF1rPPxVtnToN8npylrxYf7vgDfiqKK+sVthZ2tzt568kAm0s4dcvTaJ7jv0Ozex8b9fe
xRd0y7wuOQ8/DyPZnWoTtZAxPHr0ZCLQIBm/xuUthL1m9lp8El5mIk4d9ihY8Gj+svKm4YJMdGng
jpGZuWEiSaXGycj6AlWkAWzjSm0+3VNtijUGpS3yV/X6PY+Y3K4dSCkbq1/t6FHH+UOlE7TsVN5z
drKenR3IAmukdWYTSaXx7v36gxpZOpts4XbgHjkA2YuSRCFx4O/ofJjWlJTfy8e0k6UTBkgbe6YK
WKBXjRzINjNfg5aYPMfZw2FV0tVqV+v/8Rj9hAzrLe2IDwd8u8cOczVkAbbgLkagdyceWn47szAM
oaCsyvLAy5ngywYeR8Y0AUeFGyOiz768rXklyQvvWlgSj6kvioLiCnCns2hWLux0hjI0x1l+Ju/X
oV1UVeOr47kgDqz79jRAiCVzOdP8Au9498ZxC0SpgsIGyzTyAKeyvcV1s3L+eWCzq14iNceI6wEy
8nhzW5RNNuSKv/0tCoBtO8Hzq/jTAaHf4ya+Bve55GHV4ELv7qqHzOTytT3mQcj081/ZJB6DCu1N
+658mE+ziLf72Ep9EevZbH9GGB4jgqOV/0uQZD0l8RqCur/0r1Jv4/dCpnwFOBemxde/5uMyEt1x
7+MhIQMBCDXdjRbYDdUnKkgO8W8/CNGbIHq0Dc6ovdSocdsy7/6MnwEDnqdQ+9wwCzRPOLpH93uS
mB4AwA9Vntd0BrQ+j63aJ6Nxu1gmOUXaoWjsDbZaJ26W+L1DuIddbuNwJ7/cc8QMOt8P4E90KNp/
MyKwPfb170AEkb9wQkNBf6wYzPmprXGK05RVbOpoav2XyBvwu3DBMHA0HoniL9OsmYocw0BN0/H3
OUDFNGKccqt27ECX59R+Puy0nqxvFU4DPT6lEcfvtm1RKzu955k+ZIG5t2D402DXxO5AFWNsuxsP
ieoYCXqlwFmRr8PoJK3GDCDQ8/rIrqwC4lKmINM+xBuPQYht4GrqtXQwxZuO4WJT8BNHwuIrA7tz
+eGG8r0ITRYoHe77UFJg9XtsKg6te0/ji1bDFfwdqfKS0d/yDOki8vmfo02d0009Vnl0xptcK4dH
8ipnTwp3hx9N6iaBu1ttoF1t+Zc/wj8XC7s5LpSQMxkmWi8htZ+FhzaepkNjbGxC1RVBWSnjJSEq
XEE50A2Y9r+FKVNL3aS50zmbzRfjiB7Dniml66fTjfbCUvMERDzvImyf+MsZ6Xe9Qoz65MLQHiFU
iT4GwOQp8ulmUTn57qp+maprp6WwQtizRaJ6UhNwPnpxlBB8RF74WmQncKefxbgZEZ5tfh6G0FId
AeiuMVKA92DamNxDGntVOTCzrpP9KzDimc5fyGqaQIm9ri8e0EL18xl/6sjAGHSW/skOaL6ROlT/
E+D/QnKHvTPQOb23aQ1fCzQUI7GNO2deb880HIQ2p+kX9nfcmV3Bifny62RrGdTCN6cGVhgRiLhz
S8zZ5IPi+960gPrqNqN/khy7Lw4F50ifQwR4DOCM4bsNKhrhFRSDzhl/lPEyfkmW5fsxdEYN22/D
3dc01xcvp/WQxL+yx6q6ut4A1kBMjLyM9GEMIvco3hhymYDf7akcP8J6F3lMH3gayxIeqqgwaBum
ZTpJQPNYJ/cBF+NsBIVEpvecf1y0Q88A8WYpcHHvMVrNTPUcJQXLYKQMYTWLKiMRg9wvr3D02/7b
dL/H5bSvnwmBhkdwSot8pt8e3qrCyerQ8+lmL6mvyl+4btjBrOSBFORBo08ZWdIXR/1Nu9R4aCnU
wOfpFXdKk2O5772xb06yas9cBlV5gQHlFMjHAXl0pKGptM7krbufOQ32Q4ymMNnOSVu8UJCNYg+i
JsvQLSHvf2d+faFAxnJ0J2UCY90nDxE2tKGdCGRt7kf96pM4MCWGut3PEC16RqAWccpoZTwz8ZnG
D+0MOMw17PYCA3z8em7MyI1P1MwOJ0ikPqygOhu6F80RMjdZUeWsXrkNLFv0Sq+purNBJDSiRcb4
8pEn/jrepEQIf8uEaLovpdYa00aVWT8S1I9ovn2JbQ1FofvDDRIbq7xyvP6dBkUCYZ6QTtorgcE4
aRZ9jIdK6RdCAfXPg3Mhhq2je5j1Rzr1z3aLw2S1s/pi8HAN6HeTiKXvkqc54yTOTuQYS8+NZccy
yoySaqAW28I8o1Eszk3W0jb/L3rq3JhdpuxmCR9ZXMvj+e1wHJhNZbmSCmOmwgcqdRdc5P7dAFPx
+nTKDwndE6gJb8bpUDBHKT9si4/C+nJ8hrTY9ut9hult/tFSCPurxn1gu+xC7gGB37I0mC0YG+oH
1V3ZM7Iz1OXULWRfLx5D8dqrGzNGZIOJ6birAy0VIfFoB1f1At58g8CwVhamH8blLISB9DOgmzer
EqTy2uiAzFAxRtgwG5e5KzGZ8cTc7Q+nMKVYOf73Vsk21InyFdkVoAjnCSqBaWWGN2ZSpjTpGlRz
sLiMDlwvCZcV4kaiirbghaxaf7v08QkO9oJ4uYdg28js5LJihfwbFTDw+rTbWD3hAVeMzmdCPP9S
jrXx8RpvGei3fEmSc7RfsbvLWbA14pqPaA66hGeSsV7/hvEZuHqmp1OmjX5Y7bN1lQXhjS7glk26
M+nEd3slZKgA9useEP62QaiH0djzl6xM9X99+dBKd5orOcWQpZ5+Nve/rWSAvLfoJudLAc4yFxJZ
eZHJrOCzcpvgUqWmU/lIUw4TevkoAjbtmDSukxoKy70MwJj8JJh488Voo77Uo85KqOcw5TY/BDBg
T5rhlxuRnxpnrbP1rPet6bMgY7gO6MUFeZokTc4GMGsleC9Zp0JWffHmzT+RVxV1RaP0psOXTo7/
HnFwlD4iV9skUahMHgTlfaPjoDuSAcjikNJo4WMJT5dWEy3u8rA1tuXO8i9ZGN17vhsjkVIK/5hT
eax6ioSCEyHm9wkIP7anRIN9vBiXcYmE2B1LtGPOx9+2Bp/ANoB/jZHpF1/iEfW3Jxl82BBH7t1x
th2iSlMj5AMY8g8FuPpY9TgKPi91nTKRwKI+RDWDUf4t8DAgmsfWDYNJYukr1EpUIeLgAqSkoLxp
wCnNWPfP/H59HIlCpPNPy5ej00ZJ1DfsyUmULOxN41JfsIBMNb32kuTvFB6V39JEiabiNjETTgKE
D2c0dvvLTB3hqjV3FZfyX8BP38YbOLX6nnGwLJ/cpB/QLBRcmzTAenSqz/h9Qm2nvmYnyu5G+W1D
Xlj5ocMzNe82PNrG/0E852rQx1UurHqa3T5E9lZJiyr4Ou7mWTSJfxL04mKz19JrYVU2lZQKspSz
S8FTVDz4/oUlBm9NkGT8Q3gqfGl6huVCiL3u7VeLMGeyTTWzpdGj3xuyDTuuindIDwj9fdRPcwUK
kTyYe76P549WU8E4Y7RyzttmKWa4e111tMBvjVUsi1vmaxKeUogsvgvJkEPgUtKzr3UjlpdagizZ
9U98obFACmkqfZYUUMBaqq8cdEWdxOf3IKyqRSI8LcqmPYn/tD5DsiTzbc1PgTwIOwRLQpWlUbwH
wE14o2FuAtG8L4BbsMWmSsEzCbjpOb0I22nXlHRYPr6hk3TMKO5OujzBoOHB0tQBQ0nzEcbHJ8bV
s1La92Xr3pNFxhTxYgHjgph2wWiBaQuxulaFP5dh9d7VE7JsqpTzHf4r/cDZMvcEyblsEfrsfaQ9
sGobG167MIgFeDd/fkRHt6OTQ5+uqZLk0TaFRxGJb7u1wKNEcZv4p4CIFtRttOZjNKWLi401Gnxz
A379wYilGTHRSg1xt3XWwaUSxmvWa+0GMwSKk4to582aE1L0D1hXGRi4ACIp3GBQnRFv2/Adj6VE
mNhLiKgqONyDJP63cIV4xtAIDM/b/zVpGm7KEFSeB8DHwiO5rLmt1cFPPSKwEPk4dnOHLiuQe75s
C3L98vyEL22/KKXRSoEQtXa0gp5JpYfRME5IwOkqPm00aRgQvB9y6E2HB3njSmiXPOquR6dTYUts
LO8vmV/zP/z0BEww0GBm6EXwEqvEv0gEValxfuYkhvS/yhVPvSvP6lfmSRIzllfAWGo/OEAKsOzO
wWEGSPdeBY9E1QftrywlPHCzAk2w5MHjR00Z7zO9Y9xDUAjvawdoH9sFGoTk8RSj6zEjs/3loIoq
FiyoKSCIXO2bzjtVg/CaCGSFjtGv3RB8aepdQbmOzZ0TkKj9kzcDGfP08OHe6KjfmYjyuk+/cDjh
ID9rAqmf9yfkGbw4K0lAiQqGgSyUbtaNl3T1NPxOU61tzIdBO76IwW422jFsW3YjBXu125DPDsnR
AQJjcA0fd53YqCe8NM/dsb5+U7PvhIuqvcjhsLWonNTUrOnOt5ZnPQ1qO7VrXAHsl4PVX2958UXv
9+RMVQA7W2T4eVJOTAVXR3WztPWVzGKcw4oH3/OgQu+KEiQKCW2uis42Y2e6KBkqtXCDiKqkq4Px
kyNIP0gTbNO14lUQICOxoTYWDyCWHVuIPEVYL7zfair4YuuEAEIxrVWLz9ozfZ39i0iBb8CGf8M1
+2eeRDLovdPNkAtb/mGNS5pF+feO0EihIMFLNkYkAXKiRLM1BkGQXqiQn1dFQ7WL/nlvVyzwDh2j
fvTJxQuO7ziIV0gCyWNJNiWm4bX+7Tsv1XsY/v08BSTXz/ur/qfYMHoxTn0sMAga8SHDMxEqf7mL
u4umWMnvgmQs9liYBpP1fCQllnwzbOH6seoR+iAGxaxPtpqBmGSNgbmzYTlS2yORwoD5Kv23BRoA
GUXRdf46IE+Lp2DdEOT4Qs39uC4cBybYQNpo36t0D+0gLHWXYP+tD9pxU/6HgXiky+FYe9CYXRsu
jRLvZm7k7Zqaem8/HbfTwpy6A4ojNzOgMXkB46rfSCgYvfLWJNOURoNBZm1yXthSJhn53SY3St2o
v1ed0crMuyFGvoE9HjSgPTAOWqsAsWxWWScZ+P8s601CpZ5OnVy4XXvtE4Xm6MZaTmWKZNXaHAGq
/y5JaJOx7557T9Km1q6Pq/cNZB4itusYgxXFEXjCadQQXV0+qHNyogkM5fR6KTDwYNuRvz6v/o50
rYBH6/EpIZ2bsNYmdj3GMw6dBwlz9kyFy+V5JCHhcwiTNLGEU+XhWGW3ch9bqKUtlDem+Td76D4b
JK5DrLwfogTZiD62jOrnptgXh4OPTJF9GWertZ1U672JHv+mZKh/cbqAfaBHx8cRelU1l9Twn4Rd
0bCbNaeteoDfI70S/YjPhsLeAQFU2U7mTEJjGhgiVTgVxJZ1ygUrpekM87+LArnVEuYf2GENpslT
4p2ofMLNsjETCEJ8MQJ4qCP/4E7wpVBqzBlcZ1EfwAaGcBGsLSVgKTdcGh0gVwcdFZ+e6iBtlEZK
p8D0jNnrZQwU1sw76QH00aufPtxGCsqkgUabc4cSee/3QA8pSIms5g6aEzyrJF16KIF+VE0CY1px
BJxT186VJcoc7DhM6SRRW9fgC1ATDsrfeOUwG77bPspW6w8dsLbopgrl2SXxH7ix3Yri5kRf8t9f
UqTObYtG2NYWIbupedw57K6fIVLPcM+8rJTVoZxWarSg12Bi3AR4YyB2Smsbj9FA+RTu/49HWm7D
ml9PNyp4hhDe3nJp9BinFAgMM5OcgBHpGrxvH6510DXK2kIR575zQLez6KjLTSunovMAlZFvAzCe
vjf0Q+2CmaqEeFkwxY8JYWaTOXCCovcxP9ailWVyBK7KSf/WHS1QCrgHPQ34BVLM+XK728tcxFJb
2BX4Ho1jIYrCQSfi0Wy2EeJCrPo4fJF79+kQRHmkdb+xVEDPtNKZfYFMqtliVhM6EgTOzg7DxBfR
sSYwEPuqygNytrGtjc3I+6KtmZ6Y4JtwNGQh4Duw81Peb/p8JSM/yQbFmp51wbfvdEGmq/c3UV3m
khiDDIvh0SSwKfrhdJOF+AdTycSMKmrGvxzy8MRNBrkVf0AXCbphexi7H3i6sCA1ERJJ3zXn2BsN
FLETab2p3ZCb1FKn+su0pY9nch61xR9uAeXYzHF8vDw5x0fFdm7IUMsgquoleprtspWrhh9mS4ln
XfKuwu0aSgd/pQrQda+bhKhguvZFxdFfHIR0qH7O68hKeMRxcH4vZVIJaWkSJH6BRS4ndojaXVgv
grHooJmWVmj3d3zklkE/NNVNQ6Q/OLdGTvHDIySgaX+7KEhFIrGxtCcyc1qExutrwSliuGCpsSQu
9K038bVQf/nybyOrmXSh67j+llnJn3KtUK34NBvTZ69atP6khvn4IIeWZDpmsGWpsx3QVjHm5e0t
2ZRUwK+6m4mJnYeLkZHH9yne6oz/T/d6K2uxAhkMlZoHGzLon3xuKff7XlCr+tR8X+WcETa0lH0M
n+R+HkUzLbzZ2ydTC4sdwUQDjL24Xxi0D0g5TZmy0Q8keqHncd/sUwxLqan7B9a9zWv+N2KCpzNb
TJWcHTsaRl57VcfGs+K9BO14FtV+KLCGQ6bNpcvoW473y/uocwX2wBQgJAtfsk/65qd05sneIpQf
XT4pANyax18JcVmzCYQLaf0Gi+A/pEdX8iC1k/yC4mBZTfVs7kG5TfuCgZgbHjF+z5JG2mRt/rri
4VLbCpPQWOVu0VAF+sAiC1YmIlBB+e+hwMKPyhdD5xo1IboK/kQVsd3iHkaBnnvCM7p7QoJpoCrG
fAqUY2KUPaOCWwu7gLdmLTH2RLaP8uDJmoqyghUrD+JcRlu9idZGpzzbp4T+suVNSnkZAZeF4jzD
snW/Wg4JAKj9oP8QXgdhkuW1ycVEmu51uFfA+0/uhpacQ4+2EV7aGMI7NunhCy0A5EWoYRPk9u4Z
NB7SjskWpu0FKZDloWDaLKBDaLh00CyFF4u010E9JpqfndxBIuAi1gnKjZb3IKyppY/HPjgvKZVA
bWyX9L78YNxeJvqJTTrDYJIjCZunLf/g0WrOQp4QGaXl+X6taZiUqATIrESFDU8n0NmlhQukOif0
0yP3KVRUZMzCiAdqLBlTrXpjwXjxJKr3hjuX2RMuWMSmI3BBKeXOWcBbmliUG2gTgs5vQ1FaQLA3
pNFEBl9wAXFoCjONq0eCcqzCE6RXJzsJoq7IX/WYi8/3X9MhJsGDxAwmmtaj5agdqj2ESGBW4c8I
ZqqJGJAiOPJFjUmEJoOjifklVlOxAX+ow8QBK8q45LT9vyK0YzXXSzgWQmq4pqSdHQzqsJkJqTHK
UA9vfFh91nGryJpqmRsTiUTF8J3586y7+MzvC53jCb6+W06m6opUqkVgle8xpeUfyIyJHPn8yhLG
e2w3bqVKxY7Qi/XsyI90MmbDtovXm9lEgrGS6HVaydfnwQO8jHQ+DJ6I0rOVvQij6/4vfymX1EtP
J+TYzMx6rAKdf4Uo479WahmjQDaLPVMVrhY+yXnrdEOSzYhyMOS8Oo7BboJKWkacISfrAax7ZbtD
gN7TjwU76TaVIhXrf9kWHGi3J169xWJhTYG5QRKiIFASUU1T0I5rxHza9W0tfE8q2hJN1K+/oTlR
XBz/37Uevgx/OKdfLGyNbAJwIlM3iohsn1/dUi1MzgsBJuhglZ7SQwdkaAe4/5mBodxwZV+Rzh/a
8oxMU8vw9khxDZOwrGdvtOSreiWTBiLNhf2o4tyMGNJ/BovDXOh3kMUAixNhPH9ISOo3kknOafLO
TmaxDY0hPHrGgNvxM9Q/QCZ5/7xNE/BiDFrSnWytMzJA/d96ztCvPwiXUGiS1rzRkTkn4twD9irm
BT0g2eXTj9yI67ftD3XQG7opMvzJzmMC7jatTVPKJmKAqr0UAs5sUWYvT9yno77sXgITnPNVY8dq
VfxigncUthp4DbMMzZYn5IAMNk0G0uV6jRdzVuWo09BCEJUcupBGCUQZvOSsK3+T/DKeOyurrURd
n9I/wkgcoKhL8yqyoLmduqG2BnzFOd5pevlteZkuZfoyOID8T4tskfZHza72z5UWIB/zMZJJeiaK
/Gs6lTtaddwDhsvbVVn+GdwKW9eiTozHj3YE1c1QCOj7pyI5wkN5oAyiuCTaJ74ja5LhFHyGLpL+
DKJaxcNCdoZAbYxkGMzgsIXdvtCt9ydLys8h7JQZlJAvcLg///SJqWfNbD3KygELQw8RAexyxr65
t5IjSztkg02Irtl+TH6w/iIO9SaVfVc4rD+2eGz5pxqyPtQdbgYHojP1rtnCZ0aiz9pHeJPCDREv
jeN8DMrc4AmvhXjuJbB/V41KxSCj6kKG7WcoqAJsLFU3f6H7mQNPWyx2jw9O5eIBMs/d+d7ZzV+m
6hyu20q6/Rcs3GuxL85GYncw+qW/urd/CiiquxrK0iA3m+2GndrP3pKk5688u5jAQRJUuN8gHfdc
LRvOTFEuviY7ZgXI7ruTXNQofEEzd5vWcygMPXLACbBboWb2adq+6X8rirwL1+5nQMhxTTsxMjUf
qWfWqP2CKzrlSMxaLDHzUC2AXA/hbLEiOdlOoDhZSfW8wwo1X0HO1FYMY9pCnp4X97H5q63k8w/+
8hr8EWazTTr2UKm0CWVcj33TIuos6JCbXUDZBglTTOXM4LvI9Q6quvtoJER1ngfOHfVGSKyvh8ID
ONp6PIkc6ZeLqJVfwcoBvXT/RFUVGKDg6rj+2o47YGYhx48CtSvm9Y0WNJB+8fw7L7mkQ72t2bJY
pwiukQgLbzdvS+HT02fkCu7aUOxxI2aniiRbAi2F8GqDU1DtFRBwKaMZnRZ0QW6W5sijC7YsP0ps
I3IbNjPeoNb5LrT0Z3QCqnlDqGRGJ4ezkCIjJzRVLwlFISVqVfBAaCw7LaksFHNKq4Vyy0MsGr5N
nM8Q5Fk6HVyO1r60snT+rQVH8SjaTwKlTtzYktc23988eY52Tc4hnFtq6nT+FD8QkL8XufMYu32R
4lBGT2GQJih0AcsznetSNObmPw9ftgPnhMvOOfb2sRmZt7QYQ+s7m1BVTXXSqY2v/07vz8SZFtao
Dtd3md76tNHWqNRwg75UMlI94ICFRW7RSGOOwhJeu7VjzDNLKOOjYChrzZQTWeR2cr66uDdWrn9s
b7uiwNvOFIcTMFrKGC/Evz3fGxBRir/5DvpgSCmWkeMXsll1jCZ8a4rSh8XtVkkaopoSRKDoy7eS
nRxkrSwYFaiQFS+F+PiBIvS9HfyUKUnTok8tKz7VUUeOjoW6OiofE/lnk5QzLezKqUT7GBjuUYCB
BePXjKflbjZvMCbgngFBrJa2+9b2b6KerOPfoewuoM2OlaR2Jw1NhLZ8+B6LYVSYfetOUQgKu5PE
Wul8VHiSNCSfEcyz2jyW2bzxG2mla6aVnGk4Ojhl1QJB7ldT4TB8fOeJr1IFu8HIwj45Kqi1Zi/a
vpuLz8EsNuVvjFcViQvralLjcQ7dhGbWNO4UOT20cJ2tfWuWbaatq4IUpr5q6dHgLmIioyx86v15
jkMIxxuZKUIvtF4fK0Zc3yLIOa4BmWjOGGYNbq1am70Z5svZPR9alSzvHKApozDXjaIJhhKAL3SC
G3W+IZzQSbmqlr3WALjoV8pK7G6+SUGsyOHZOsiZMAV4VOnR/UJ+PhWO/NGCUgO5VvC02ivVjp9f
6UvYquvLO/3d5L+U2EA80wA7ELcTokNtbFQIX3k9TzotqDI0wXy5Zb5lHiYu55M7XTCwriqa3mhV
N97akFgEDEZut2lVuQvI/9RlmwWLPgBnkDnbeh9QIAiN7i24kkjP6lSPiokmIkr/c2sft0kaNM6M
U39cY/CWVC15vgELT1+m1CaIwQ6Rdmvis8PXHIY5F25QO++bAOcFD4MWnzaK9UEX6soF/iMcbdqN
RLL/nS7RgNSDr4OO++oDR7yEdHjcmLZPneD9ddIMwZdevgYYjBTQj+HFsAyqV2v7BoKI2qe8YDJ8
hgB1YF76vH/yQU2L1scGTkRE4nLLkEj/BpDS/UN7oSIxfjjJg85xvx3LQKge8donSoyBtZ9Po1Ii
jznGo2c2p9IHGa7dMF7NztLQWQflvVO72NJ4OZvxP4j4jJMAu1aCTom+kw7lI/EHyS+tDGOE7Q91
cncrT/2hMOciF+a31iQBj0ZRuxpGczHgue3nF7CrFXbHgpiGJi8DJ3OLTmUKZOh/FFe0gdXHJ3GM
xJVSpfCBwnRSmSVBCAHKDOpbR406/tdwIIiX7nIhTZJMaKrr+lFDZOk0PrjjO5I15kTD9i6/8mPp
1Tq9BOmKl14qPbPSMrauK+2NKQhXKPcCDd+ZpYPmj920zq9BreF+2ZAVaG5h0OHOwXBRR3y9UuS5
v9vn6QRapOJTZX+LsxeMSA83dASEh6hPUZNHOA2TcbBOGd5/QqFkYeWYhCm2S837LIyYuZl55iSw
masxWoy8FlAt0YYdaGHpX4cAzBTjO3uyoA2a3ljzrcT7R2NUPPfBz0SwEqz4q4yyrgA5B8vGrAer
T2hhHBk+RF7/UbCUnkpo+P7Fan9UaaAr0ex7i0YsjKIcix51rMEXPltj3NxSju/r8UnAUJxvDTSr
oVZP6gDn8k8hVwPLJZpdGmpcXitRRb53dO81GtDWGjYDOmu7PNWwgIy9OIC4U8LIjv/0TECfKp3B
/Imw7OmUxcC3pP04tKXAboWGyt08B/3DIqFHpfTnVVqb9EXiNvzkLotiKa9YmuA/SLziPnBCnGdq
uHk+D/E9MzNbMNUUpPjiXbtYAN2TXXv9m2HgP+4gTW+nFGGDBmzt8S0nj0WvXlYoBDylDC5GS4n2
MzQRjplMwGv3uW0ahtJamg4gSu5qJ4CjXjqVFf23TiM74jrSbLJXZCAIvZcj/z6oOCDGfB0Q/HOm
HrQr642S3ptTS9GLmux/YstAi0tqJ0hqcCMzVNZbCTPUmDW9eF5WtRW+9lUa2kUxmFvFn274lngL
W8pg6Th95dFE4RjnUsOQo9jE+dtn3VFVekWAKXddZA9CL2T3Oqj6tDGUiTAPE28ldiYEz2v0FOaj
hIN8PVj/5uk3gIe8zO/2miDGWm5cuicPuDXF3kKgqKmgmemg7a7OH2dkyyMWdey9OOnNAKeQew9A
q2UC7X5zGjP7lnWOTwPha7zANlRB6wjrDOLHRZQ2DNnyZ6BRQsxmPBirlC+2N46cCWJ6EnxaOxA8
EIoVYwEPcIcYqNHEr9+gmMA8eLyU/wW5vqYF37pQOV/+1NFNSGC2vi99UnssQklXQes7rbc5Ad2H
T7YyYYJiXneTZcOA2WXDSsb7P+hSO9XPa2bgSaXorTG7FdS4JRXaFoQe/uYQi62TjkFJlD5LPdGJ
bYGzmNsPSjwXm2BxV/HJiGZxH3HGbNSH2lmt/UAV++nnlwXnIeI6DgwU/Ct8UoO0BBspY3rWz6SF
KNvosItd44+1ke4FkDHvs68SQ5HB9I+A0k+OX0288NA4qaX0c8RIDOC9hynfAj3qp7btWELSMC5d
kmmmtFS3XpYpTcx5QG3YNrEKYhYj/BKnPeAWUg+OFCGxPFDP0pJLlkn+Y6XPUvpFw8Lo2/KgckzK
60x+LDM6P0t110rYxxVQ0731i1SrTRrDwS7uwjx+INuBi87ovQISfJvrqiSF0dPyixxO+z0jyjkT
57ZTMreMKpznpkhq1pMGUtKnzlNzupJbXmTKImODgBwOqH3ibLDjwcfJdf5a0X4Uv13yiamfjO5K
OcKFQxYmhgVjyYuwKb8zuu8uiqs/XOaNxQDpaO1rorL5I5oMZQo92L/L5q9vPq78vU+euYiDnv0d
72MgH0c1RWQA4YXYDMRUzqzLu+gZmqEtxGb3aHNwcPt6YLyb16Fa1GI+EZVc7EPgOe15K1PeFI7g
ZhmM7/8rme3u9QtzxztmdNFpWcaj0SZezPqofBreqOAeQAJagTySqFpmWFGvVyEnUqXWMOUuVidR
TitGsYyJBwYqF517nnOMX2BPYfGJU90qcxbvpsJuKXeVkIS6M8cOfVALOWGb0WXSHEz8pzkVwTc9
GQCW4feg4AzFhdutwFcNTC3dTPJC22sr9CTUaOcCQRG1yoe/aLqtVromvW5hLVLXuU0k5y7cOJZ8
lQT2cqgA+V3U6BpbQevNen7nfDyTFoDISMgoIRrK5J4PQIm939phXvs7+mpUWnWkSoSuFV2KmYzf
TNC4W3GM6RUdXBQRA/w/PfN4Gp3BZLv7w/skfINAiCvavFxmTCjBzn4ejrmCvxGeoNyodC7KZk4J
W/kdTueNz1zWAPbZVCP6Srz67LK8sxqXULeA+gdYmbyqhByOgKvvnrDszIS3f3QV0hmIxE7yWHsu
VmoHvOk7luICxFXjjvm4V+6nrj6BmUN7H1pKDJ6mqxNCy9Vv8EsQyse/Hy6SuXOma0UHOkBgmCGb
RZx1UjeVheOjTl56geoRlHB5UFLqY2xcUpoMCrPQq40WNdnayRclDhHKdTdqW54F9m3aBo/vbech
wg8qb78M+GuK81cpq1taExmnS2z1J3KnRabcB9oG7fKxglQDe6d6g/ubYn/krXyBU55YyvD7EBt3
xO2s/8YmCTH9qWlqbyFnt6W0WdpkTyGgkqSkRVXvOBeWm9Mz7+GtrfyWdIY4Mqd9xxAiPZVRc/1K
FM293dFXvs29dbQrMMo4s6kFO8rb6heLeHJsdo9YUoNKRTNOFeL7aukmXzDeGhA5FsTT0OTuR29f
FyFp97FPWBi/r0aWet5MMU2nSbhmdF04gBhpPJChslygmDz0zGsHQFhbhPEqMXa3Z99mxZb8lDJ4
gASgbHvx3eDTNr6RLyFVpl2UqxAXiG3Cacn6E9xug2zuVPg4SdHGjPBXKjF/79a+TCGMbIodnsaT
aXFDiKWV0BXy/j5bN1ONG1QjCHRHvpG08B9M7b88pn0X/FZGaIDBCJiUCcguJqHXonW3xOeoQOT+
UWyEWUCtxYVPrXg8Y0Az0qfOlTnVcdFF2ai4U+jWhJpOURTHJXWrQchxxxnsp2BtKKIouBvXDLiL
aZ8oFLJ6xxGkieb9l0TwwfPr4fARMwrJhVriuYfl3Qi5LsQd4Xs3o5D+zeCqco37Xx2EbB9oN3/T
WgHgc6qSOn1a2eUqmDojGFSO23WDxfRPMa1EkMblMRuktzKObQdm8s4KwFQubMGDEETtVzyb0bVw
aq/Fc5s2obEzXP4a1qpswBvivYdWdkB5eX1csGHsmoYi8aKd9Udr582l7VNss6/JDrq9BSLNQGsa
7LKc6xuOcXCdFvASA9VeG/2EBIj/6yb0CJ3dP+pQc+az2j6WUis7JkUqXEVG/0vpgDsFd+CKj9pZ
9WhfAo4HPGxWPMsPzC0ayrq5chp54xdBbbzewCGvDCtPJzpQbOBp/Rw6fWWMrmBk7urE2Hteidnu
y0EcBtLPNyO6hsndGQuuggU5VTpWQkuXDh9njrZ8AsJKKRcKFOQsUr71zj4J7bAgbpzc8NwPeLSR
fbLXO6gke3GynsTgRY26yxYKNa9neY+fHTDcB5h9GDe+PEjLFNIp2yrf0sFbuP26CeQVbiyEuExl
yKuGS87ukF1Lfr6v0Kxx/G2XwXIckRbimAN7kLg0E87bpnAPLU8C7sH5nL6cUvafLI8OoI7X9sdw
GgDgkLbid8RRyiTToy+YOYQ/WpeYbUg0XZFksIZPV/WVW3oOJMFGUvRpDwgfCYJ2C7KZRQeIFPtv
APuBAM46qXEhadcTnCVKDOrIsVua5wQYlCdWuuVbYd54twfBiOQZZU+lutKZIj7qJzwlBaX2FrgK
LHmYkVNWHyIMAK66itL+P3rFRMClJSBb++pk9WwXlg2bEYFQZ7luzLJO8SFZECe7BPWQY/P7f/n8
8KaehFrkxbzoz/bY89zFOJJgr6TN8zvnQccnOeZfk9uRmsRExsLFYXc6Mgtt9YOuBsFSAQ7V6+mX
4LBQyMO0hP15n4w7ldo422uKjGPmgRZUwVUQyIV4sU6hzvtvsokWZqKrXck02ollZxv59SV/pjtz
J/AOczG1Ft2La+Ue+xsy2Bo8Cle4FFldRheWJrzXN3kDKA5kZu6gggNqNzaONUN4C/ILJBvdioYN
qZKzklvRkgLMJkllWVs4r1ajHa0R8ZqBSvovFxSQ/sYhgmzzAUMkMMpKK9gw7GQxYq2rQ2HR/OPp
gDITMhvgQM1/VvkXdP6U4/zakX+kEGDTkHNUmoemXu9fvLXhABr+m/kejuKu6SHeXREY3qtdMlmY
wiI5t+2HE8swQwUS4GXYFRgNAn/z3+Y2RFDQXs0QCRqpAmu47XrKvA+XuTeamDsVUKl21fXEfqD5
+2YfUggBMJZgb5o5QubEIhMTXgfA8kCvnO8WVM/LfmBjCh4pc5/6b6xyIS8ncY8gvfTiUhvFhIWQ
76W/BztvVEirEke9wrKPsGasu4U03+cVxS8ZzoLSwbECccjFtiHr3VlDgK1/FgVM6WZ2xTY15XwA
HNxLTDmIGNJiuws3MJviqypLj3mS3ddMCaoLksx7r1w2amsd+Ep2jaYze1vJqWqPl8BFMIO0OX53
Gq9esFLJmXTKJNkjjkAXxWz5d4JfKaKUcvp4KG3uZOHuB1/BR7khVt390JOK7dqZb3gFcdvfP4xF
MexJFiwSHKlVUrmYannF0sHTDAIZMmScjMpgPzHm7Px2bDr0aWU0HKIJ6T9KXoVqv9ppZW24nzY6
MXMmArCDRYbyCtD+PQTCzXNt/Xwoi9Ms0UmU+BlW7tplcCNro7DtE8/eaD62AwozRNCyWGbpRJA6
hXWs48Lw+/JzmtIU5By1OX3wkElJjiG0HZvgjs5ZsJmD2xAbc/e6SuuxT7mSfdCu+mDhsYbl5Qfg
N9XQbpVHxTVndNNKEPO1eZ8P91ODf6g3UJRXEORJ5FwGDw2E5iv6oUTg/ZBnbjcc81dJ0ZQ8fm/W
CilxLqvag/y5Ghwm5HztXIDRkKWlQ59SAc/zd5gWG1ODHbGGwkjyi6+icFchtGDMp8xmBmD9HyOt
BaIvftuU6FrqE/T8G/Zam3vNi5T+9M9aWP6F+hHNkVhmumAkun+LEQtYaZZzCdZVxtI9rNViZwe4
Nz4wOxUvIDPuc9qKvMCkqNzShErX0xLuH18bp7bkJsFuzYROjQokwmP5DvbWqnr+oQmoC+KW6lbM
g+ZzaxyZ71ufHpN0HEoSerZF08Fy2yNZET+ZhYUr9nK/R+/nNS9xD0WWLFf1x5IKKrYZoWGSQ1+R
Rdw6f/gjSWhxZH1QjDgVXMympipIgCsMNywU5u2vWPq+UtIpL380b6CifwiTjIXxiVWtcODUp149
ycMIcp30GhmHShB9xRboRgKV6C45munkk0UYHDcUlIWcMecfCXZsramVzBHwwNJQoLmNbK6t0K4K
zP8TLBwnnleEWfL5CVl0mmZGizd3p4RgPHUaJi7I1gJ73FJhiLpf3I75RjFznJsC5yntiXhFKliu
NE7hs+yQraK3+Rzv6SZkSPEwk/FMT4hMLFT9Y9YHzJJD9DZGMTlCyw2iSPNzwcHmyIqOUaukz48j
Bti0SZGuxDVNsG93Blv+kklMFPpJaDxl/AEZKn9tY0yDhCoNarUkOCE6vML8DoCCqAG2nBwSwTht
og48oAAAi1sxnAaY58pU1rBjzC94g9Vqc6u7TZ9qN4qhb4NVeRkkDrCf44ThRHJrHuUJV8d6EGfe
ScEhIX05G0WQHsd/eLo/4I4qElZoe8usHfQreZ5TkEN6r1vLLpdFDbJkmno8rdm/MRkh1GyMd8Cb
YSoV46Z39CEh3ma18HyWCrYFAxKNPqLGysXA2kYzg0DSOgA1wvfpEJJOxwX5aDt/Jr6YgltsBiRn
kM/x9BdRjxCmjC4B+bEwaQBpIXqC1Irp3q45rE7qBr0fCP37vd4Xo3NSNYNrIlXwkjP4Hyr5vGJn
PSPNgTqkcA6Su13ogPaV24g7oRJjiWLF6XMIfiRIo1ar38V+zfMYOLOrJ5ijkmhbnMmbyV10fArn
uPPD4wgw/hv0iwhQnU1+I6kYlMc4zhsrvBifHR4pZfCo4mbRytBlarMuIu6oJgM1obmmLf4xYKii
6iQONH86Q3Fe4JTonLpRMqMwEV95wGIpQKpYvrziCtBYM6T98AALeFV/z3w1Q45D4LbN4eYfIUCn
hQAZPh82Cm7/VURMIdNSb6sop7H2d6kkn0A31rv/pcQnIms3B2wwinUrojCqS1a+6NRmiZS9gKwq
pJjkHKyLw0qD/qPVSXVuKbLzm/49l/amtxwl5gMmmwTpGdOmzZAvqWRlueQXpMc95udJ+YsQsTPx
qIi1CW3BHICiS9fGrhfCUpMfrsAfmFM4iAtymQruUZ3YXYECs/nqnto6wh2eg14CLAApFijnDCr8
HDp1pHsjXLDkhReuA8jPWpEKfSSYJDvBui22eWKs0dpnNPYQUUBFjojDXlsMMjvMBVB79wdLqAlD
Ow7DzuvXVxsJ67OPPVNnmrkadZzuGlVmQsvnRTpEOQXGI0oTbu8E4x3suVXZJGnoFVSm1lDg/kb4
C4mk3vt2BlXNZOc8imLTnjc/D+elGk4cwGdVxfkmbOU4idg0okrcDfg9Hbtz4CRhAFXVgQbFhA5p
3K79FHuViHqc6a6wZjoMt8W8F/C9uwLvczohEgplQBHbGAw8EOjbl6BGZxodfwJtZR61Th8JEU0Y
GSL20Ovdhf9HUrS7JdYdnuUv5cbDyXC9elr63pmgjbl/RSUDVpPIF+xpdzzz3qzXcqmdKSoP+SsF
TsIZpWv94Jq26au+kYvW01jgyhTYPmQLml5/lrdeY/Ei5Rg8nUPQ6RwC6sFbPQYUfAbVjdcQ9VWN
WDM46XQuoTfNcZ8d6TREFaE5oeGnpPBCZp9pVOW2pdEMQRFpR8QXhSZoPvwZxrRgtrwYDgbFoo2s
Gc08WDCXu8FrciZxGwYAjG6UKSet9pPeBpqKW9GbtWaOia8I8mOfyxZaJ0BbX7L5qrU3rDnbvGA9
zjyWPW3S0ee0YuD8QI6iZuBZrJXwbAFz6VY83BlN4Ce+AN5j3rNi/M8Bml0ulGhlLOFTrEZ9QCLw
2iHoTUzKZKnvyMPaOPT3Js090VegxPkTy407MIJgylDtXoh/Mw5vL3ajsI5uwHMYBB8JxW4thh4c
qc6fxpmI7T+iBNNJ2IsFB/JT6OrVnOsFyM/oTvNUeGNDeBKilW/0jjAVuZN0P/ay1j758deBPwpT
suvXPXTe1Hozqtu6sv8Dt+z9zSKEwWmn5ElgYBjEjsl+cBp3yR5bRVNH6NGXSs1Myx72U7meADxS
T3dbe4oqWBQFjMFSCHoZvZQTV9zDFRyM0zDe71aAq83K//sfPo5Z5CuQEvLZn+LeD51Wwsso53O6
TfHi7MUHQ45jTcnoCwrNfn+P4R1/sx3AYbJmBXmhsC1WeZesFFJHwgVXKOPaYZ7+gkQUGBRKQIF9
vC/WmJrywcjKeepDXRz+C3WX9cD8VHVCH9c/84qdnghLzXNe0Lch+X70Pv+eUMpTiHJuGe7vozQo
fgSfRcODyE932fFjqSZl003D/5VQkofIP95CqNUvDcFTvtTD+QkC6tx/Oo46MXWKE87AuwhcgUY4
XXtcCGeqAvmIkSX7ewiQHQGzrflhPwvidwTRPsYcgYODgCU6loqtwXEsG+EKvTIrIhTq1jjBkU3P
jfXKRqzNUstGTWYZcB8IT3CKHK/yrhEsLgHczcljUnswDTTM55hTfW2GdRhQgcSkEhqT3H1A0r+v
dJQyVsbBw0JCpV6jn/67hr6JYhcCYzlB4OzLtzOVHB5gVT40t62pLdb585UxHmA64eERYaI4QexS
zHgtoJ8ZM5jOzaLgOJBevbPAv3DUB9x3LXdXYng2jRbJ1X4UDzmis3GC08nV9jM2vtsAxLcVpDa9
5K9zgB+qie47606r5TkokVyNIpQvjmtKgTwMUwp87FG5Ip4qfIDPUFhhZvWdjVIeWiGEuj1Nkb0P
U6xqseVmOUomPHRZRY7TfKHOsGKSlXF4jKI+VnKU5Y0Bvlvqwkk+mLEQXHHqo+RYTtFRmTdOyvHR
TdTMcE45OebEH/8p8F71tjZuEXHnKvTyrQL7800PjpX8Gqpz4wg4TGJjDVvWdkprLllWtBv+TqNh
QUxeJ6+3dmVR+M31dl8lxPDLZ7Z666UHa+cjYIdlEH/RS/hbxlZDlIbQF/KNvkBGxqTLUkBB7g3T
uf7npAQNhTBpCUtSNidwWnZokXHG7ORQcvu0nPPzK21zr2gpd/pmJ32VqsYKmYRlovdVhEBRXFz+
tuRpMgYXHB+Nm7m43Gr1ZaIEHzaQVORKg/wcYhGA/HM7CUmnQDTS/UvZBXiJPnnpcLlu0V6aMzIg
pAiu/Tix/mVQBfMmgxyn9ye75aOHdTDbUgrueYkMSeVJaMGXGGgYmCmn0fPYzApbbrbugFyrQLNZ
YnaV0X1mZEt7DJ5gjbCHKOHWgvOQ9QwTSe/1jW4z6XOQ6D74liZZY0FpSugnqwV/v6FTOPX6lW3I
WHfc+w1vFmSZzNo83sov7imJSry4UqNbhc94oGa7QzL5fkLHRaL6L7yEzXU9ty22ilM7fGc4Th2N
Zm+ApQxQfsXr88TUxHY+QCCMGk/gyomAPmuh6Sc2kdEwVaYqiIM3XRt/iq+4VOrIZWMW0Pk4MwDO
z+SlnfBiMpm0wETtdD14QU0NeT/+0HieMJiH/6rLrngawIhSEk3cOKaI/CTjDghJJ9zWtFcLal1/
NBlOLAAigAKCq1Cwy2FwTub91ljgnpyS8T++4rj0pDWHoNZ5y59UBzw7g3PhrCateKiwbJJ+tblS
j6jYU8r/3RFgbZjMOTZTZ2l2mgG8TyNsFD0pVwH/yBCszPXd3Ql1OCIO8zraC+2HhoGHTR/pp2bX
V++UaYP5x2WqeBD7y5H/oPpQyAfNOJYYJPWK9A8spD8ciPZNvojL3zUC/3lZd8KnTb0Q8RxAkMi/
EHvYXZkeJpyuWCxHK9k3XZ6DAD/02CEVZFHxXUIAus8Xa4p6l3mi16tpb5b/M9zmbLF8H+IC2y6U
P3Q6dkf0yD1F+RaYEGFj8MOhzUulsFk7zG960z+ao/EUi+LMASZbhXxDRpOXAnK3E/7nDhdAjBzK
Wg3vE6M4HjgQHCSQsWtw8IHFPIiK3Tc5ErKju0R3fbDrkwrB4iDkLvuF9tVDvOO3Lzd7AmiMWDTl
9RKVMocHoXGHBHmmeboMqHFGnCWqoLbyYtxxe+drNxBILQciwFiKjxeff3ihvK6w3qXjy5Smu3Qt
TYyQH9Q4F/jQyLVDS86HUCFL4ClnZj65kACxVisRvY7F7bJAz/hEPti+cGoIJHA4U7zZqBR0kNez
R4xFyNoo1eb9REp8oC7uEbQuJR1r1mkMpWQWnXQtvA8LsAjMwl4qo5ugFdzwN6S3ZnPaB0DJ2wQq
WxVnKfm0yt1WH1v8REsTchFe6eRPpdxpwEMf3B57CcKqCshrj3JE4jBh8ba7VCT2cAOUUO4tIG/Y
SwxaTB0b/4rMh4VTqS9A+qZD/bqA8VG2CcN0wPAuX0IleEcHRKZwXRiqIrZehlt51LQQdrCL54Ol
ErY2Ip35lQGRCKY5XYIjR9FOpzyx+GVAl6pU+MGWZFaE1mDk9ndkV8O1MjZVZr+DGNxUowvspT6e
DoUlAPnDN81hxlpdqdn+XhpIoKt+YmvntLzAtfdD5rNdTF921txWGWIayCyxiOy/yVmRdHCzZppw
PoWyuMRsyo2nmknOy625LI1j+YMEJjER0/19PRiiRJqBKcPJreFWUTjimVx46qkhycPcFjBT7pXl
SdIE8yHgnPpD657m6ft/A1g89fLE/n3ljx7t5tf54/K1eQsJmoNsALoDR49tWWaNL/nOo+setuSq
mw/UJEPNfLcHgTkgedjjp8qVlSiKsOm+E2QdFwjG3aA7vsru2Busz0sKpDTqopIzONvT5Bzg7uqQ
6j4Fq3irJjvXUi5RM0XWfBcaLY1BGDj5ryYbnusHiunBdFoG/mtA4jt0DW4isJnIs1BaASzneRk7
HjKJtfgzwOB0RZlHzgKcefA9/mKHAOQdjKfPqaE4FLY8P07YeR5sH5RPSiF5apB0BsO3EYioR3KG
wX8BRkGR/eAFNVg1FmaHohz6rCJQncBLkYZbHcWN9iR2euUbpt+QqfHrwmOfdvyL2ovP+4NrhclK
2YwGPiDEkMF2roNWtyG0dsdNhnTPB/BgdZSymIDXmz9YSSea0pF9/Ung2dDtXhfJ7CvPSrpNNRca
93jgnZeGdusYnKdoxq6Kp++eK0yD892d4Cz97cxndQeoXPQJGP+KN16xNwelJLLBuLPYZX/AENKL
jWKx34S6/6yYr6RIdBxx3/YDdRS5xrozQOmWGL/InK5pgDVVp+kJ4FDuBydgZhmMANaXAC5WO1Nt
uHQP6HaSNM0K7MZT0aMn3QB4KeWEC/gMNJTBHVqJrPl5EReFNCmpYfdR/T7DSAJb46H+cA8vNKPw
UxGbU8QR5QTuBHOqiWPV0fwnjg4eacxTsTQ5HOWPz5lXCD6A6O0FsS2X/fRzZ/mV/pKp0aGe73zt
MXDCPMo1lfapBqxvw64RLRX+xPwbn66bkVr3KoSPLEr/UNqFUiMjLX8Jlcyg8n7Qv9Kyuk8p8tVu
sicyhIcnE23xTtvgtwGvC5k1vRvTG5vVzCY63QSs0ygAgkYQ0pa1Ms1cTlWBT/27imGPaf345L+q
vwOy8zT1YPiWepkF7rxgakNFtjjeBh2AGCjxEJFi5YCXvUimNOpeAgeTYRJUo2EusduBn/tT/egj
EoLxGfRuh8TXUf9cGqVzX+HAtsW890nX6tRblctbUWNyJqzHmp92Hedc2RlRMW7rfOIBcSnfCjcq
l+gqJ5/y0O5n2FaHXojzEJFUyRPI+WRlOMLQUlTJqWMgfZC1Ymfhczs7ZfTIEECQOSEg969Ytkmr
BR7qSn5An/d7agU16a2gL26UeztjWEGoQTGexbVMEbac/uKVrD6qrpAWwFQx5tGFTSx+uumTMnK5
Shg4k1crnNrtX6CuIS7Za5SWPqIhPvrU/G4RgI/k6Q2OAjum1i24TbLPQqrbirmxOSM1RgPbJwL/
pfmFhWbtEulr0WyL+zWliC5mKDxw+oVocO0L1QYwZ3doe0kQWbL348etfE6wttGDoltTSnKorNNU
D8keyYqgaC1SMT+wLh2ws4wmN7Q+RyK277gbZA+lB0e//KVq4sA760GRhhQgVXVsEI/OQAAnYv/q
5ClpmDUVfYKcqtAqObBppDwh1rALPgohxOfiGVkQs4Rc5+ymmZjAr/Y0jP5qqz2rD98adQ10Zbv1
5xnfeZGj1Y+mGPaygDHoGPFib0mlHnE9+cvZ7b4a5TnaTBl8zOzu4R2CqAj7QvE7c+6t581iuz9y
9xfT0IRPtGeQxL+kt1gVSxNtWrrAwy+0zDqslL1v/oZXBpJy6KyKUIOBZ5NzSnGKHBoD9UaxRekn
3KOegkOLUuRVqwYlLkO4RFOYMXiP7oS2s8vLX+N00FroJBt7/uKQ1nvCSgJtMBH9N2CfYQ075pqt
iolduWKyrMISlvVooqJ8UjRwHnED7HtGTSi/mq1PeGmuWoRfvFd9B4wMnQ9caGo4cPkbF7e2BvjV
xHogUaD4UO0y4lpvWZLLJfppCzesWySCNEM6JhSQ22sN6Cu9KtctaqDNFpZS2pTNLve/mOtlziDa
MPPDw/gyMFu9D0Wh5RYaOXzXgqlBcpsascFjIan+6m97+Y4Sxs/G42deRP6kvahY4v4mkmInqbkk
qll59B6kPKzl4dC3v6DKSDHlUkZBP+G0CdHjjU2IYlHohHjbOYjJxJkCgUOpTQirR8leK9xMjMsK
5XnLs50AMY4Af7X+KMDK//eXNKwsIPkJrHgv7B/tzZkW6x2qobmVETHvXDju96BbUQeR/PRmBdzy
ChZ98T3vfaJl25ZDapygUdS8QpgrR6vkN78MF+8Qogft0B/H2WwxH2z69tIS1UBfjiX9LPQyizKK
8nEudJ7Q3YuEhIv1/nc/ugfKQq6hvIwyLzJVAxEIpGN6siez0UBCvm3e2MhoT1wZwjq+gkXnHyXz
jzufAXV5U+0tQljoz/1LZSWd508I7VLXMN+3Qd6vHiv5jTBCYH7V7IxzJ7gZljouXxQYT7meV65Y
lBk9uN1fxVTrQ+jjlElavQ9QTQ80hlPMKVv11EOJcB28t7/CZ5t32SGz0nFvAfJ7Oij9JRp9QRrQ
1JfgvZCoxNc+HidDgJqcdGQrDiSQZuDEBhcBIEDi16uc24Xry/6Ry1P6eAfTeJORE+Pql+TE3AgB
i3szS8mtnEYzyL0KxAtTYKyOsa4RvDdVY8Wan+jiPz3ZcDV7kJm49/DXt9lTgYEeMm8g7f+AwhFm
MLhElGjwzv7PijIEvAVFZIaTfT6QRCnrnvOU9kXc4PX8JJFcx8d53c1YyvB3R1KIBjicfGzbEE9S
PuhVvzBJntLzy1YZq1SmDnvIO5GInTkopASkV3pgUYuD2MHbeNhGCH5ET5VlWGMM6wYsybpszGfZ
LS2HTSs1d0znMp/RCEpZVpGrSEENPfjKHEokuwQtqa0Vad9tHNlziuHNyjAKucH5eA/8ddeyQzBe
c0FUsmEpM7uwzcq2k9lX6phin6Cjvt353yYKhzoK6oF7deVlTIW/qfIxvYEw7RWTRBVxO1VWlyK6
6CoLcwV+qcNXMwcx+WSxYE7DvZYURTeGnAgQxPlzBu1PRcMOwDLZwkIDJZZlzOiMjJ7YKzYq7CF0
K3RKE4uMI5pQA9dkwUk9Ljtn+s7VE+dgaSgtvtl5bTzHulWAtGvDbrRrceKX+QmUOrUMemzuxr5s
I6iwEUZ2BwZBJB9rYTVOJFgLNmVHw68DwgzDirPVu2QEDlJLRlgexqtwgR6zr1MbNz7emXP0TX6R
ThLoVFoHv5yWArX9x8oHky8btpp8mHj5LSdlBYsYCTkvlMyBNUipwzzL86UHI3LVn90NBTDF7tzQ
8EICHmuJLT1qpqWmOEot3R9SCHBxY1MpGUo97BnTvkX5Me8Nv3+IXG75NNB2ufLF/GknOZproWnv
/sN87Xp0iQptSFHy247SJx9cGc3GcSKKifIM0L5qzTckVtqKMivISkksupWi9X+4kwwuGyM84jhI
Qge0//o/0gPior/zjfmqtPbs6qfzgGXR144fFG7B+wEcslNjgpKwB1rRdGMzYr5rvofspFMtRUwf
uuw+vnvyB+4OlP6FDDd6LXxPmgZXLdYchHfR2HXtk6PolNyJT+qLJi+z6QcDRBN5rlcd7iIr3Z3G
NMJYYOeECWXAjd9DwUGeZOmDB1/kJtcbcAiDnL1oAwRs8UUX7HNL7x/GebY/EHFz8mW3gKq2VzDE
kFIO28kumxfs9fRFoG6qniF/d4kC9TKYF7HTJnU2pEhKgSXDV9PSMWfrt0SGfFdAXBr71bi+DxYY
jC1u+kOtCQsgEeKK2wwN7iX6jyikiV8TNLvVnCH3ymBw7VnZeiaYYP+ToGTAoMa5FMWNNemQzrRX
R6fja/s8xmf7iggNkK/luvIYl0Zv5l3F17P10wUKH4s+BT6vAcObWQKdoASZlnMsD+amr7V3tHeZ
4ByDloPoemNb00JPnRwwo23TwI/phVRgXpocOGKqxYR4gnLud+3YKYUfyAqmOpmHQ/v55AB4BPzb
3jZt03xEFJ8dzWwhceuDtuApZxmotoxsJv54KrJaAc6Fc2DCzL+USJCSonyLhKukuftfT1JLZ9kE
e96XYO9GI8fpiGvIB/dK5mdMV04Be1SCeeTZOPMQgnIdFlIE/UK8N5yFJOqb4/edgZ3amFse27s8
B7xQLHHTStDFIRBl2zAPZwnaBU0XNpFBjtf2it26Qb07rBJiqhkNRi/rSq0dYr8tBtUZlLZQ0L3n
n4oysGBA8vUUCsycDVDMKpTY4VdWr1+/hEGEFhV5XvY9X5aXBU0iP2CcTxW94/foDoB41c6T9Lsl
J4o3FxgN2iA77opbkMkBBbIF3dbMeZudqSVv1EMeUmixLERz/aRWNUtx9UWOf/RGB0I3JT28J/iR
m9LDr8taX9qOkwJt6z7U7Q6cCPhJE4hvRdBV5hcMv2whbkbrkQ7TfCxkG1MPv5zC/0Fg/1cy1wJO
iaF5TK5f0ghjcH2QwxR702XyUzGUp7VC/WyFyFashyNd8SPSFBESvcgylDOpnKV3WW8osjfxU5rW
JnRRwQ6z5gmlZx0p/Dx5+EfeOc4Qw1vKqj0owfb5YWqe/bArsqedD7pxxT8QJ9p2WZR4c25LwnEj
AxZghrItjaJKbyQjD5zJfdS/KE/BqNAosKeWsxjpBKJzbaoLLwdEShL32Sgr+Uy6pCukU85V5P0c
s1AYsAMnEdi54d6uZw4VNYWfyur0A5mkmvCw50px1vIiHE/glL6XasXexKXjbSL7mkM4mDJ23l/W
TS7Z80DX6rkMJfMvO6sg8A7u8d4j4YE5m8TFCu1njuGl5PzaAy5XDe5MxcFFBnryOnJnXXp8Wh5H
5SJs0kwTx3zRALhiFJO+drFrsbs4spw7SJ2SNWMjLSH2qbzDr+aBpp8TpRZG+v+cFAIqZ3XlNa08
pl+m03m0pN9xyM/2FnQ9JZZhF9uc7W+3HPQDKt4fRBBC1TLgngk+b9PYlkZI33jYu3NgWdcfcmeo
StjLqUCQDzL6476Lu1d18nsT/R9MAYckfNqRLgc0PKIYTHdxYVbYDX0+Se0iQHtr+w6E1/Bc8uWE
JvRv8iURyWpVBtGbvwpSLc0Y72JBnPDvilQVkbihKEBgWmNT5nr5hYXzcYK9LEOFEBo0SY1WCbWV
Gr3gWco7SpoC6VcLc87WbwxRGd0LnxF+fUY2/JOkVlaCS+PV4/sFaSkJ63j4pXHrJfs/1DQu+ZoN
TrgRXdGGn8gMtT10FpzxGWcoQR7h+oePveKMmKgxJbNtalwLWO45X9ubHcgk8gqrMIfyYk0gYb5H
rpH8UT6ntvazruD85oqCb/KMz28+wGiQjwDQlJZE6hTkdnQN98SyWOyVj7jB3QFuxsJYHIlH2PXS
ZogDGZtQPEHSmjqcipOoER0G37EW/bRGw1KOuX15nT1EKtIPwKWrU4UNyPWxGmUkak/TnPzKprj8
9SR2cRd8XaCDlTvUktOfWfIuPhIzGFSCoOCawIzc2PKuBTlf8hO0vuFQR9sEOlBS2ZrG0frXkmyR
/FlqrUXzqlqbwFss4/A/YjBFX/Ll5y/ofb3YqARNmov0MLKfFa6wuZqDZoWNky785ctxln0k9pol
OqUc7x7Aex4MPzD8EUyc8iVda7BgB7V4TaBlb3h6PmuASMl284QDT0MIqeeLxLMg2wDOH12kD+jV
uQOOm7/tM2iL8a38o/JA5x/RSIRSMyFjvxrQ7iOlreQzUbdP5VZm7GZ7T9yepis9n+lSu+nudO//
zshxUXldHu2UU8Juu65wgQ98Ih10WVDtXmIGdWGsghkvuJvzrBnYIF5eMamqVpPEQWVY3zvcELAd
Yx8ORx3+lKa/2v++qbdCgIAdJsvd79j7Q8bYyTLXuH/+IyfkQfdCKbTKeSB8ttfm2w5CMXCWugsF
UuUxLL/zUydFXMf+ft4eSlKo/tUhj1WqpfotqurwaDMnn3Xo5jHqzHBcS6OKwogXPh8xh8eahrAy
4B34QpvvsC/o4+tpUwb7W4wWALEGAxL9dmOjh4YQ008CVQsOXp/nly7ig+CxMH4S7rZKjcaIywd2
I/0T2oUbVeh2aypN6uJds8lr54i25MfiW2T9poXCmHlXVNjRlBx/KOwJ65q1LEAHxFkMtmAuVN7z
nTdeQQ+VozghXZ4hQcuxrLheumVAMvEM0BRT98RfnXM3pucqZ+O77MqMcMikePPKfuGots9IFybH
5zgal/T1ciozuhopg0XPDZkEVrp5I7Tf4NgMtDoPl7lfjlrz4WfZzn9gftdxKPgIoLUCmsOKJ8Dj
OJ7SVUwmmPtqPG0PdRHyaSHogPREjuoDIJPnX/UacEEyJJkVDzWf7Gg6sOTBFWYmeY6MKyjyIY5f
a32+U3dfwDRCNUNq1L3efgE2CTMZrC4/Ymv5tTILnhHg5bA+g/g1OkDgE2Q2WLY3vdzSg/ZOifn8
fwpQ7CGjnQOlY9q/8CdsadBPilepUXTHRnLDBGE18Z8fepLJgWSO+4434cFeqDy7z7j3xbWvVy8N
xr6HVju15smz1PLaQaSBv4Ui1qHYpVeNgYwe4mvX7GDuhiF4cOmELBEcisPC/qB44SX2dB6x9ysF
7VZxU6UlknE9qzk5uEUucPSrDOOZg4Ff6jxy3BZMOnkJtl7cK8+Ev4RdGKCYV6WjXMy4df+8CJt+
Z83+X+0p/yUnEiMtsi5W18jXMaa4MT/fxsNLs99NcnQNpL2lSqkpXwk+4Blel0uhBts3nHvYQoTP
9Iu0TEgIkWZ9w5DymZTp/gu80o0GMNnuEk5ikdwHnrJdH5eysUFcIcASsWxu4LevijP43JvAIyxL
rUSUkIgy0OSjcNaID1r/wzq5qxDrIGLHmERmFgRgL5ROgT+8YOw5kHALASFc7wvj2XCrmlnWBJ+3
PKwlQiKoNoXjLwieks4pqgQvKMpqe6vUZi5qE0hF5N+u2Ntmn1QIbfKYvN/mAEnJvf2oUta9NiyH
Lt4JFAba2+Uh9tSXWXJ15ChPKaiVtgfATXb6igJnuyxKLdiC8vMm4+P/q48IV7R1lk1gPc2whhF/
s1oogoukK2bMGIuo7q6lSLDK4+qFlErTmBKl3qiDO0oA3Cps15577g4mypEeQaDfU0ZsRjoDitZI
CwGqzNDmfHDRZCjGeq1Nv0Ln3rK01CG3nFug1smEAchErd4gtMIIKng8g/fPCleAd72MYdNHgCGJ
lr2Th7VwoEOw49WJKRsCY0bRln5AUroBXZPxWmqkPQlAMo7vUmchJl8ngO+xQggLaBDb4C69Wir2
PjqNggRjMtuH8bgV6HWEJf0ouNrry9u9D/BjW2lcWxgC5EhKyp6b9pHodbLqIyHnnvGB+CaOcKk2
2CYutb2/qEpHuLkGEmCr+eOYc0XnyMW4iHLD89VkPnRoOnRFBklFNBlROBga7/Hr/SN3wJ4l9nLE
2CwGMhV8icKnfCohX3XSo6xdnhhs/upV/XF6uL5wOtRzPZQwg7yu5s4qXODk0t35FaSvvyKM7KbI
VSofMYDo30YEXItLJdb11sT5+qcpcgaepWJm2qiR8oUI/qn/+PNC3XYFItLxf/LfaWwqJSj/nIKP
nfJPu4zl6E+8UdBTVGtUsgNDLjAOV9yXJCHwIMLaOD0nBdnCEiM+WNI/nmMRo2VQ2mqXGe5S5g8v
b0YayDMj5gm+9lyNsqAitSY1m7SEdU8ANuDWH82ObMTlFKoazDZiKm8PQguRgpVRJBbWUzlykwys
FQ6EzonVcoQU0TlnkTaXkgvhstudKhIeDE8VqXnbJbBye/ppGhu2Q5WsS6etklio6OpiliO24Ivz
bPtQ6i1boX8mEeR2cJGyhAUbCmX4bNYyG+exZumzMwsq1wgUTJKpxNdI85jFQlV8XQ90xd04yaaL
WdcyUNZnFX9b4U5Sio3MQ2/jSG4pXjI8Xa6s5TOsHMB2rWCvoGCptEWO/w5xQU7TAUekjKmkj2dX
XXXGIIEdU2VO4+94gIgjygmsg3d1O9AeWd39siuv1GCgoY0gRkBXtA3+6FX4sn79NwtDiaBx4bpO
eGmJcEeM79DlZ/apuC1TmlMBaRNoqmLdjJpty4+VivaDu71dea71figuIRX9vuF71etEBrOv9Cut
x/TTFFa98hgYkSHFYpxaJRn1/KGpn1eMffhUcwtNkFWJui7z5XLkqKZ+46uHVqEH2DGqB2ktZXaP
qXfu1cVMEPmAwwGfqTwAiUvnw0XF/wFNaDjYOiEg92PX8lwnVztvmxHphhpOBXXlCg+dyEc61uVQ
01gcj1S+o0Bi+CtuWjqwFO98gB58qQVhEWWJBwH6i4dfsaA3TYEGFYIH185Hr0UIvZclbyT5TVfS
eUifRWQTPVyorQZ2At9Oa+byvfFfcLLRWSTtyJ9CWsr1Ms3BnFvGq2okcGh4VQHzmgNgUZtVX40R
pkrYrWRzoMdbUbDKdxJGm+KfEp+8twqrrGRU68m/BmWtkzxSu0LKQ7BkSskNBLJgAB3fBto9Qamv
wtH0F3XInLekDT5a9WTsKQJ737ICQoLdHHL57QNruJLtesungyJ/HdMhvDWVQkGCXB54/qsQ0ez0
mNQ1X/i9MXARXmA+BkXZisdGkRpvRNUlghis1Ksg1O9QVjfzcNKs1hn8vYe7yzHL7FRgatJcGeCa
cquRM47Ky1pMZDG9v41JID6FPacxhra0gawI/yXUmMPzD663klhCauM0nlUXiQIhb47Ds3Hi3kgA
/USt5UPCUw5mNt+QuAGg22N5AuqoxXiToqhDA2fpzQW94/kVev782T5I0/WBCRskQ4affcw9ZqPX
gdSt5+5Qp3b5zuMKLftIABoE8GLxMJZ1VKBcVlrYmJX5bUGTw7W/P2pehjVF9bHNHK9vFQNqC1Ds
4j4O63pg1iC182+XCi5af+vx/LC1d9sw3Bm3uLt+B3CFz1fTaiEfQKGYxEaFVQK/7+jx4Gdk83ai
1AgT2w8xNvD0n7xqRZJLCkOnITl79yGN/DXzRbYaJl/mnAgVnR8HQ5haWgWG44qMu0q7QBV1BmXD
xh2L8r7d9VsTz9OXbuLJ4pY27ARZ+upATm6DdOSVlb8VRUFQNLJ4tTW3P0ldmWbxRPOoEW7Sg8AL
MM92sCwATb1nWFkTZ2PT/UiwYvEglbY79ndMGBIsG1jJ02JiO4Jr9GCb9t6sJx4JbuIuT5dAOATA
RUpf/ezbLvJYSrCwp/Lp++uk9Q8VgcJfbika0BC3gaAgQ/fJk1AiymyBaaIUl6VQOpiNGy6XbOrB
hcILrKBM2cjmUQL2pkA/TUqn2OQbFvs7M8vvTTq3wJ4W2Cg4FxvsBxQ3XpI6eKPaE1o30316N/2l
s04+Q0POvlk58E4PP52VwSbvv60fn597+DCOXgGijenee7yb9j6xH16TdA17DJufBhGkMVUaGoS3
woboRETeFMiAAe7k1CB0u6PXevjBFPT0xlUpLLIjXvF1P/IZnV4wMxbJ3yhHtvJlB9C6ujRLlTlQ
LNoCTK3dqB0r74m1YxOqzj5xAO9e6IG4UQEvLcRtdNzbl7laFhhinEseeaAQawaBRgNyRs6zmW6I
JNMdRNHW4pRXlAXCpgpoDfIj5Uo/89fAQlEzXZtL8JjWumWUQY3/8GKXt4BnRKvQ/zCcTdRp5wgX
N+7+cF2BWPWIxx+FToykllbjqTwZu2AtBqNLgk47aHwVPpG7zn3aK+Ilj/lHV1jvxG8nvUD+2xB/
Dwi6G/TlA0wCirJoOs8iFJubZBG2s+OCHRw//kZB0A4RK9xUTG95Lcf19ERYyBdieS/eivDB73Di
eAeQAgD7n3uOW6VgF/gOk/nOQZZNKypNZP3THXplYqQNRT/VQvfr0rfk0fRcy0BxJ6XGM9VkvS4h
p35LFshaL++zKHjvx+dxpfMUXsPeAsblIaoy1xvOrg+3mPcygU1eQhM3Pi0u+sWwN//OGjzeMjwl
UXBEE7e6Sl/G1A5mkmjjLM+GRPLTocQQidNXKDo9qtHYZE054g/xv+PkmhP+GkZ3Oq97HRHQHJ4L
9ULc6WuPhJcLFfDBOebcZPnF2irILKnuaZjX/FRtRXuGHRyFhSicfTkuirXUeVUQz8XGLB0QYw+r
mBgfuli1pKFFN/WUnwsyXa4q6lVzTcFPfAtrA3oBYqHJFoVf8dMRlNDjR1OEI3hCJv1FwKv2czi2
aqHs1ACktTmfLrI19XXMahqMBooilr187CKEpGf62KTvAM0qtRl7KxfrACbMSm7xXSmUvezNJwSd
Tt53SrS0UEH6+pkzfVvxftY+Qp716pcR6gRKYMomObqgGSwhWuqvO7ONv4dsp1EjtjEUAakQwkBs
fA3DmQe3M6166Tq/DoNCpE6kW7QQFAjhChuZG3o8ZZX6zEWNqfsO5uXAwOoBQzzU4b0ZXZXLnyIV
7dNiFKzR1pm/3gA8+KsROOlBSdDLcPAIRgZhh3LqDGQ6k0TpuXD06A/qqxw54ZyIk5KIzVQUnXIc
bfBI5yL00ifbxQGJQU2q9/IBXWCczAvOlpqPW5C5kwzwbke9/A8bx7QGMQl6rG8YnHieRgijXn4a
93JzeGWt9RpD/aF8E0ETa4Ev0eKTgaGKdWAdscap9u6DiMDtzji0z4mwARHj7UnQbMXk5g9c6GRD
eaOGWDmfBM8a85x+y9zXA81XXVFGFS5NkmsjDsWMqCnoJaE4D/C1Dv6jzUKJJLysMffBAVPcJUsf
6HTVHW9n9P7kHiQl93sDNFoP1K0Fj6fu2a2IblCFsN1TuDhYTbunu7mCPexjoabO7uo3KJzrvr/t
hrZmrPhXxFGquhItdrQGH/e3NTFRV42ivNtxdvi/ef87G+ePrgvvq+Jt0p8UHxB21LlJweyaLrh+
LESIeA412rYq3cN6HyzggEdkJjcKTN0r7beO71MdF0FeYvKqvcs7IAhASzOs2HHs/P9ohJpR32pD
ffJ5x+kY35dgNS+QdC8Wgu6hxiOXO9rya/NmnkT+tI39swNQgAA6SvO5m4g0zYkuCAsCitKSky+m
sarN2wblO8WNLY7q1AOzlRBGaCbwYt7NBTAS7u9b6DWLIRgNmcxV6yt3ftqLXLDZSlBgYovu5+wM
wL8lWwYy+oDTncOM77kMDCr5E7ohKaGlirqMAFqgdRoo7uc88Nxuv9kwwEUq4NF8gfWg4mbQKqAn
LVqKqbmxjLKfDzsOAQnD50f4YyAMttG9qPfFLjGRMb8/71lrUYOnCHyAUYmuqe5TOBQ1s9zGYfAg
p8SPejHzSWOT8jhcFyn/E2Za1tl+k4S6L+Of9pEE2IO4FaCUP6NnvY58Rz3sxxbq4Jxx/hDAm4U/
zqMsczbbBJzvyQcFDhEDwELW5oPzWapMh+6olHhIGIGPf9FkaF7c2QrjUFNRAD2TYef+GPD0USEW
9JQsELoJV908oTHJg4rIN7+aVHvShVhSKMUl9kZ7BQ1Ml8b/cqR5F+I3K38hubmNrE6WlKYjPC9D
5A4/2Vy8zeDKiheYpOKoRkJT2Y5evL/VXipvJqHRzV/PTSmfEwuArGZrxgDEwES1bJjZPdR3rnkI
3FRo/m5FdLKY+epxE1PXh6BJaUll/LwHA0mHqHybWzn4bWlfOmk4qkHccaxnXdXieB1sRoL1PPpJ
viULRuhFz21Ih2wXRtv+y165tpdMmgeUL58IuwjwQ6rSsfzPfEZkKrWMxkpReB1Axpy69DUqwMUu
xmHrMn9ez7/i8B11OxX6rBYBlbWYBtRlAO1mIXXm+buY3M69elA2m5QhKXrE4FTyEPDWxSno6ofp
4EDP26fyD4+ELEK86xxXV21EoLZ0A4ZswiIpHvlxrquXbsorGIcF6832JepjiwhECpvOgHKVSqzp
VdqHs5SyzH9eCJpEasn6LdI8Ml3Zyvp78SsgpRoDwxJkU/A67f6f2+QCAw+II+/Xh4XAkvekRvZc
AeR1eKe+LeDUk+q/CdNrQE38ndFHcxG+P/LCab66LI1tvU82ij49evnDSLMKsIF8TQoyn9cUQ60A
hJXnuMEDaxhJHkRxRbbleo0uyo8qrDVJAfatlkkIhoccep+6V65lxnZYZ5hPIbubx4f+IOqb48Ql
TN6s12MMUGEcikcS6QLFNiya3ami+oJJeaVh/VihkjhyGMv7/cRvP2a3iOnmAQGW/cee8HRGoM06
H9SuFDorOEeX5Y8qS62UWNYnsCoE+U57hxifZAlpA31bBd9ukC7PHOPR9bpAPUMUOIooG2b4R0XO
bWUAyAhD8VYlQyXPz+QYu54wZ57L//TLaoRfmJklbTG9DL8qAWlsa4waFfFUP2EqNUtiLJHb1yXS
c7zKGX7GZNnrHo/xjxGVpzZZfbJpLTyetXQlaIqKLb++51EnQ/Km949QMK2GZoaBYiBWobCcAeZl
HKoyJ+zrkGBYy+SgAhDCS8zHOIRJZtUW7QFXMqMhMElCJ/NZ+kiJLZ5MWIL3zTplcGHATOegjoBB
2syUnck3vkC6wBZ/9FX7RQofaYc+Pcr1p3cTb1b8nylgISNW7XTGF3C/8gtUUDSQu0kaGg3vwPBI
Fn+sne6Dv+7r44iq5aUr7SEZsCYFbt/Aiwv+uIRV8zYxJK4h+ucbh5qNvGiJjvRT6qTGAtz2srmw
+Ct6i+xVgIvZmF7tyvSwVfINMlidTseoU1rM2aPu14HLpxNwVVXtX0J5U1x+MSIbB9qv/KPoqiZF
tXsz1+gf47FwBVj/jERW3yD/t00aP/ZtQo1HLPblM8p68tpp9QWs8iKcyfVFiztohJOaTYem2yI9
0C9TUDWtFvWPm1QUIJhbtCt55YX267yFQFNkfg9fW7tRz0Y0fUFdDOoQknMOJ9U8wRvz8R2Iqbg6
ZfVYSAUp3FeKX24xn/W5KO+4UM4W5ZeVX8YW9xRjCZ8wambxGeTHl6Qmw4a82+AgYr1m/BlRJ78M
MJ3i2WpwFKbSP8JulErHzCTPhk/joaVh5sr61Qz7eHfynSfzegXF1NGlfGpGl29INjKMuG9qo5lb
rysaZw92vTg2JIE2LKvXPQHbZrllPjtNfWMyNZDckTiZSl/MOOqaN2/VPCZ0t8C5nmLtyytoYCHo
X0IPxel2fr5OSxJwqGRO8f7dIAHdyjiCDpXKrXfFqsNB2bnJWfhEfXLDcYZRwrwfbGm34Wp2AC47
f4BDCbP3TPZ3kDCIHgOVqZ+U7L23g7eOeWrQsyVImcsktygQCBlXA9oituaDOigeQzUs7Xinoedv
NvC6IRGX2G5+7aNeh8axIIaQ0cSFrdCROCnydh5ZK48FRH6I0GCd6vzNne/LX4luJc+aSNoquYOD
GdJRgGKZedF+zRujOAtWYRABBxKV+blZ1DGuklZJ9Tjgn1PgqskDTS0OAwRfg1J7IyPLs28A6zpX
YOzha9JZiX1xHdCYKRLhY9PV5Cbsd0AfdmZlaI/Pb+OHuarr32jHVDminv3hIPgHAthA9aa/sWc+
eku099S87l5TAdZUZdbCNbscl4CRL5a0VL1BPg/IH/EAhoCyG8ixfxO1xWfKKPLnBqSmCB7fRRTQ
GBk334yulYACzua+ngNR36AKLVr55cAKVUcRcaidcQ4TBYiGW5PKYdJBYYJXgmVJOZrUljL7qYXD
mDy44HaDOaxJ93or5RfiJ1MV/Ll4zolnck3z1nAgOXiRpBqWfqcYoh3gPkzcOYGETfPJkdt0+bWG
gkM1abgkj5uS403IVFWpMlA808s6/TOWSO+CSBkFE3CSQsrt8sYjv2vG2e+jhwN7pVNHRqrOh2in
VOqkDGAxMHIAvJDkBQauH/glNHqS/Y+ZFQo2jhDIiu+UhKmPwa8r9q8UfC3OdFGf7aGYj5ZBME0A
6Al6Lu/rzxLzwa52BvfEUy/JlpQfT9hOjqIZBB6NyUSI+SSqe8mrmIC0fr02ax6iAr/B0Od0iZGY
1j6sYYy19virwW8uguEgd2xC4RJCAlM0+sMBdX6+amIXG2diqA7sE+gwXuw3lliCuiiuTFI+bz0i
Wx87COrX7XuPbp9S/Wcpq3LCPeTbtmgktmMt5D3bwTJW8iHgBkWp5arYR5ZAqZakTu9F/nvNNvGD
mXRFDIM1an3NxLZER1UHPXNm/uRUVVWgp1u+hdDRnTWUHtBqMIw9Ccjj6RUhjASPeRmcGFqDXJVD
Gy936BmLxEkrnpNMwsOUgY2xd6IzmFPdMThjLOu+d2/aVhMhgD45y6VGRmngX0ZxV1BuQgLw01t4
bia8KOON7/IuSo4nHCLQZAX2lOB5dVWUjlvZtXBDIIzQiR9XgX9xu60qJqJZm4eYXQKRAwhSyQOt
QKyDpIzAsF4c8hsgoxTBBvkUAUSov6axV1NV7twiUdxXHYGBVEb81CkwdOg9ndFcXe2ofJ6FOWXl
PAueV/x4Fl91Q/LHlliRJb4WxNjG2E4HZC72qPFlItpfxQQsvBKrGU0M6Lb2ATXZsUbVZgU0C8/h
SLQEnCsWKtMlEyDUb896EemzhNT9OLPaLmYHVbjFPQva0GoaGXq3pUXHac+elKSKDEDaF5PnmtRh
D0vV7N8Qf1kJkhFCE4myafltEyzsB+shPNVW1wNEYXOrHqjwau6fktMxbh07hcRlFhTKPXLsT9Dw
/U9GySXkrVd2Q4QPpvJ8FKRAlPXuTx2T/VeETZDLp8v1ZtQgH4OFbDqHi0aK31OyGLyIBPgXhFwj
L2MokDHa2rBgGUG/Cb1Jv+rVrMGw5oZyVnpM+fVqKApoiUdsi/5PA9icO2XQDTmzQ/gN7nMCBztJ
QPbdLOgV1gyknAzJfZXmLzXrpTTSsdY1H5kmKoPbO2fLetFRE+xgZrhwP4UR4zowzN1Am2Ed3vUl
ONV8lcMxmGUOK4W7+r5RroaLwag5M2YeEpvNgBZh3XQw7xT8176wglSPUvhFOWDdc5eFazMWNeJU
MW1u1OzpThRBXZKDA/cjuZZGQAaQl7DJNhaU9PZgEgfOLtkdtqsVLh4pVCg/iOJkhxsA46rbK2xT
7ajFc+CBM9ZMOK0w1G5dx8ivsv0qh9/s8jwCkFulHdJFDQWGt0Jrs7vuK4M0kVAUsLQ962GLJd/w
W42HS5KCq0WxnIe8nW5qFvTRmYw3EoZXsAMOm/3HDO1umPQLnqND2bjMV8oUOn2Dmoilk7vlOw8k
zcnOoMVvJ8iNEl/PhzB6LBxtg5wpC9UE90l1U7XnBNqSfbJT3l3oTUuChGl9oDisFU64223En11v
pdMUAgd0Qn3yokgE0dSoUKkxG4S9SCnlLQdE74dUmmf8izAEcJ92ANzLvNEP5lxAA0CMnWFF0TUO
dQBXJbkMcxg3C6T/qSn7j2bl/sUDfyeV0VNpA1RmDmgKCilrZRBdGbahoUvZPbhZfruA8cRnmqfw
NBozgiFOH34tv+aXqd+AIlx1QnbyIKTEy+nK2YaUybcURsV4TmNamvkEs4PbIv7llqhIPoSbC3ry
kcJ1gvYof9FVQJ5k5PjC3mhNK1mbo9iP9PPTIWlhq58RHoP/uYJBrdWaPlJ0dki3X0rJ2MWDhxfr
IEE3a62GU0rOFOk27bAQIypNHcqQVlHHhRPwxNTzS4bBbInDltGA5uy9iF3uNtvX6OcsAL7oCqrk
MPtGnM2LkXsMgizCdAA5BjxDTr/NYYoY0akA6bFPatsrtC+qKA/x504aeKkC+TIFfZA0lVHklEdP
lopsnlybSjVOW0YhMZG1f//Yg2DP4/3Gl0HKiF+zAIdSX4SMYZu4/lkn9e4plPAvWzeeaGllzmFj
RJaKQPsgLoeq+bn+zSwv9QnSFZCYz+0oUwiE2/CgBct9uIRdyoa+fOkGuC1+HqEJ0AVyi7pV1UZI
MI6yDTtbcDfF1D8q+4ZJCpujbGAWKQ7v3yIQmdyMUWTCbnhWr5Gf3A/zx4RezVsYvonKLJYrt4dZ
x9pnm8n5vRdioa9YXYm/VASdQt8th3GWOR0/MNysIBB9pZsNg/ZRo/1QwlOvHKOZ0bLWxvY2HZ6m
crYsEqkrcJqPsnHqhtzKA5c1WnwrXmLAAG8V1ZgfbADRs+9PMu2eexJQmOn3zchcw5yf7/pMTh7A
0knCL94zLQONshsZWjbGlEo/ZFmtEpnyu5Xy9tjySteVkcUpBXWz1NCx214jHvgpFFGqxCTuqDrD
qrdNX7BpaflGKzGyFgTK5Tv1i7s5y1Sh/X+ebDG8Hl0i62a0KXcz8zDFCgn6zl++UshzbCAFYFhk
OPI5magNUg8yg4RTTgPLYTAAmhHxivOyRtDq4HCsQ/MZks6CMZqftCYGnC5GyEt0I0Qbe1CBCdV9
ZRvwkqETwGAHJzwDdjxDEA6iDXvcDbClRgVYY+SjkkVYVE6pJXvagNpRZICyfRCUJClzUN3p3WXY
VGAH8/fult3tfEG8heFHALIzK9EuZ58iT6tSEZOYShv7dhHHugkMnW34AsJxeWWddAdx3sX9LkfA
AVHyoZbI2IKVivT109a9qYjho6sW+TYrWuQsSeoetla4ml8+sZ0pdEe3agqtPUV2Biw/qic1SSGl
lz4pkBfrb7RZX80aD4geCRsl/lLKI4xaI2YR63MmJoczgWDqHVgink0Ky3kI1fjNyIuEXyiDnKTp
PrXau7dzW5znOI/BY0yx2idAnX5os6Xrq2MrkaPs4DZev69YO2LDqo75c8efndXXs4Huu5cRu73f
AaHNRNCloJCG27srRa41trtk/8G8kq88iwEOj2aK/NLjcCDtSb500OQq90YENiWibjTY8ig6vTWK
E158OfpcKBCvmNmaJKBTEA/9CHhc2e5xFMof8eLbXo+m0rE4k16wQ0QTfE8Ucf2aE9firKjzp5CF
5zf2Bj89bmjq1rJf0OjIZujeL9F933ujz6Gt4JdLOsYq5XjNqWca/bChph9MG6M3F3f8iHcn57J0
6VWvWfVzoYwrKJ4WBDeafPtP6BmpDlMn2bCzhFMCwbDrXPch2/8/Y32dBDa9aVH79Yi9OXWPnsBZ
aYNztvMRn/kwjsfQZ8CLFy0eyjFRbg5aP3pc4+DE7IEpjsLzl6uWKWGo9H9jjKqmehdAGidODpfL
L3Jcdb7ynvQDV3F1MCOgybjDVJgYYvQzmeR8KNISTk0ukMEmcGNeelIOD5VyVSSXmqmeQqXaE/MI
95PoCX5HKJj7zdXMbe33pYeSQwIlY1sgQXToA7vJZfJopRYlZtYK2mFYLoT2z02aYDKHvuddTcNq
uDQ1HgSUVdlB/KdFT5qkfu9dF9tvZHSgHSPgXIgaUW5Xe5pG1KLT4V8q7XzPDpT69heSFujFe7oF
LEJg6FsLxF67Ns9tw/sdLj4V5aLy2/ET0Or2UY8dBXjVsIlmNjPV1/8m02+9a9qQk3tEoB4rSw0Q
77h616bS0c00l7inmiO2CPb3Yn4Qg5h3r35+14/4SGWZ/3JrA2qGK14z0+YVsaAonbqC+HGdAzHe
7ggQkF1w8hKS0YMa9wx6iAshvPxbk65lto6rP+aeu5g3QXhyYiNah0uQz8XHSSSAwGEhe2qsUc7+
SNj994r4qcH8XskzUo82nOD3stg7MCJYPzJJZM8le40SPYYfFYjFPkeb5t93spOZoCDa0Vv8aQRB
VMUgiSYgW00tkDdLp0LoHC/sdHY7PvtP1bF6mnsA9VKFWYMFX87mOK6dFU2OJ/2YVIH7TVdUQb6+
OAkGu2D2HQ7t9WX2y9SgkOdNUrLdkUeo7shQu/cWUIjjyqe+IfSPhVnHJD4/pCGX5nQCUD3dR6OA
yN/9w9JB7NL+DXgSwOy22FncYftsA8jFIBp11TqhNNKLrRZDkeeTe4eIBdliwjqK78o0omULtt50
BVoQeoYqd2EN091d9B2jdkUoaUwgRtslNHVNHeR8mi3DkAqDWcSBX2xZvWBXf27pnD6ULqhS6tIZ
eu5Fwx95e42K0eZZVV3UkXqfuY/FupJ+z/fhXXLJvyCKHwIqDDUImjCPZZ5jl3/4pXPVRpx7TKj3
G4SBB60r/81HU+6W4XHPRTqXu3ZPMxxtO/HM2cHsVlRncqZ1IStQ1uSfdJzFyfTun3Tn88TJRI/z
DEBvwoNWbxv3fXfAWIXaZeNr5TcEqOD+MBMrZOBZO+8iF+URmjBRtFzXNocXXat6lWuyA9jJgwaF
odnTYMsVe1/yYvUPRsbgXR8khJhMk/JTs+pOw0gRjZpl5GP1UeHYhnGZ7UU0s6o++p2IVkTct6dr
xdzPeyMRD1ONrLwXM1nFy1eCYb1JZd75JsWJq7TLijjR/hK4IhrixRoBz4NG6YzkXa0cR8Fgh8Wv
aebAHkQiZwwqCBkzqN2FP4WYj85jVzQoMbUDjJQOAFeJ4yqXDcbITmb9KYqLbeCZqdBeAtXTmPG2
iiN+FonFDpma/a8B3euUZvIQaS9SEDV4CSdMFjUgZtAnyMHCLQ72LP1+lN+kzA0yFnva3RWZMi2E
CWRBmKy6gcrjXzQieQlfteV8NmoEosT1n5x5rIe+8B41SqnBtSxTvH92kO1KQsKbTk23ABeWNJgi
DoKHPEQ45VRzgVq+hJmZTglG4bGX9xPpCFYY45ZxTJoEOG8L+HXZDrZGq1VszWx8yhu4ivywq9fw
BhrT+dULnxxeESSmPQcHB6pcJtXK3HRwr2TJ9vZ8lxVEHt4EqRRmlL93nPLmsSeoIr8NDG4h9hBk
svLxFrxGFZx2ucg5YF16oM5rp0cU+yOEY+1JZt3IQjzUBDtpdX88gjF36eq46m9tzIKlIaYTGRCS
PT1fdm6l7qRsR6HU6y5+yD/O68PRfkNe1pzZQFAcCQMdM1WLpDtfoC9r5ag7faNz0/vFCEzb0vly
KdyHKDaqLSGF513I0pH9uxrp4Bq3I0f8NvuLf7ryLK6NeSAnxmuc4Mgva2qZEcD4LNuYwhkUvbc3
FDbuM9J8xQEq/3VSGepJq1ZcHL1PtJo88qedLodc3PpNQ4jytDSN/1DXsWWpGUzKwWdm4jc7sA/s
uXFgqxyKpQj/jb7IlRI9y+c90EB3xJbSkNODBJ0nKEqjqAoM62A9Aqe6ouSX9EW2WRLDHBKpQ8Wm
5l+4SMfaEMIiIwakgfU4BuS1XDi2l38dUAhJ/UxkA6QWehPzOT0RmLGSTeFzl79qqXd09stoZtCA
sk+YHPUji4BpjXcD5nj3z2hOnnUypp5w4CE70RmDilc2UIIOel82y9CKfEpQ3+8vaL8CMcdJ4Z6Y
4zghh31PMN7KsMzv8TBKdacnkGhKCBPFcmf8zydj2DQYzFxXoAlgxOKDKveoVIZmA6uGQ60ZhUcR
aNugHzZ1DW6aRfuv1IKE6BMxXFSF+4kCkgUy3oALEaSWqgQNpt1/tyhXlVx/s1woFek8V2VG4H+u
oyrLi8ZfOPxUf9PB4KhHgcGQy8ZmY0Q+lFA3xnz6qDB0V59UtUkL1F8RHqwHDI8dnva+t0juMmrK
jYCqz/286ZsxAtSxwMOJS1o1JhEMIiMkyCiOeY7AZ7Azz2noNjBTxc93oMuqYFUKSBM/JZ40t0Sd
JtlP+Nyous0orAb3GoFm8vjYaoq5TEJEyjRn+hSriVtnwrIls2H50NNOnLY+er5QgHwOaIxjH9yc
dH4TctcoSMYprKK1BvbWO/C/B0YLo5JwEzskQMiR6mtvWQLOvPFRM85tVUAJQ6ueOHl4yV5eyE0H
VBqPsKqwPtUDlYpcoaaSwJDbh5Wn2FFSt3e1CsRx2EcVQTff/dbQ43HiZ6qt8x6Od2bvkwzL7tqk
PnSXdLHhj9QK2ot/rdEoCPOEeCcTdqPba07ZadSRaBvhULEj3z7PI1QjMNgBearZB5bjib14+r+m
zY0uSZPo3rnZ8zJCVE7zRcpZr6yXPvQSqp82SzFk9KRvUc3niH5rYAn3CC7UJsLj4t0HDbDGLmyc
iM99XduFcvQgxZRZFKzfpG5gR9j1yFuGSJxZSYXXvNIlrGmunYe+6J5qDRBmSbkBtc3sH0YZemu9
jKdOnJAaEgLX3iyK+S9lIOb0vTrOX9/65wATVK4pNpcWP5QxTarT+KL4zjhgeRSdAdtYeJyLsNGx
1hiR4LWecfUdNoYvRcbNj007hdxrYA4UKNY56lPG/pnEfEqSaXwtri8djvOtM9x3PXjzZ7NCsPft
Y1iAsmbUUfjGXBouFTkk8J1Txc+0Ydsuy3OuucshsrXelXe6fcD9LvFL9Ttd6ChBoszBaT5s9alV
B+TJscq8yUtbKyLvrha4qgIEvT0BpdhQ2SP2UIjsu1etDhOKyb/KvfVOWi/QlmohbHTXtKWZupLN
aJ0FzaYxxszeH1IQXmPEmVjgDl0gJZO8BpK4ucf1UVC7fTVGkbFB5L8TzSkCHrVcKts5ect98Kue
zaA1x3z5VFxxacUeKg8DyKMQhLUGZSUZcfRi7rvBBDxEzmyMoDgrawqBhOGlBHCnGQeAUfArSLY2
8b9kG/hu156kM9N1H9jAQxHz2QTlP3ImiIGFLGcYk6EQMQFYlZc2TBPhChA721sZLzDD3rvbtMh0
VLZx+MLbMOYIhbHluvVotH7Jt+PycrSHeW+8VeI2Rcr7F3KwFJ5558Ke3DJ0KwaRnZFaWNSijuz/
XPi2jmPZeNhoRiRsVOncrYD8uYM1VU/3pn+WWhYtnQdt+Eaa+mD4cxlJdy8vO6b9X8qPWtrJrnVc
eoMIzzCMv7/yR4WwHONIb/lSBP5jZO3+hL/tXOnC0dPyOS/5QP4tqwj+EvY5MtpXr4EwcSOinRqe
S+iXBcb1Xt1jBA93aUKT3n8rgsAwYObmf0MaqR9K94iZzEqsSLTJ/FXe+Mjc/6PlMDQ0Ljn+Zp60
4jxcqGgoGy8i/NmAHhRNUdnT1DNAgoAcjgFYas5GGvUNrUeVsqflEGTAPwYQJTV7cr4aFYzxpG4h
fnoURyqFp+OVxsqz0/dj+9A0qQga0NceM81yLIY2TUmLtrWjvwYbBvo4No72o3J5c8JNlx1tj9n1
u1Ie4z056yy60V17iBScEwrec5hm6WKDlBlvBuQmUvkHPAscnOzdRsyv7NDOjmoSfHIvg2bMVQoh
8Wo9athQV4eABQEr0sX/wKtmRolsSiPewd8gchoFb4nEydAjUgU33sxbGyh/7pW+bbVqrs5ntP3e
tHy2jD22Ikxqm8xkzzeUupukx0KVbFl8j0L0sx8F9FtOnRoJJ8/rL+elbNCON+REHwlJ1wRNjoSN
azkFSTynIiKaXuAOvVmhl3ULLGZS0UZjpBfqD/hhPjOcm9AWTpyzgHyb8c5BMEdH3iqMOMg5/2w6
mcbL/lIqnqzUkLAz129wDW4ncA3eDsttHI17ea2jB4HzaTLGc20wJ5Pie4OtFsIKN9v/wZCawMF/
w08Vfm6xncEOn4yAaRKC1iQtmbZpZsUMIjQ8Zhvfpan2fsisfpoeamw1o0khL7FLgn5jFcp016+R
vv+Lpc5NXKC0pB+NpQm53x7PuUKlp9/Bg0Z+x4GnPgZfD1QJN2b1fsys0YVElJVGN5VV6gK284dT
83CHsgjnx5mA89R/ZjxfPcF/tqgcA1ktLFis2nsd+38+E8IofIyL8Mli2MjHKt2r7k9Fsfcf8g1g
dhTcl4TI1G/+5Lf84JKWqW/IVY+x7AQlzX+JiCiLsCeZxxlvMboQtjj3a3t8Rb4o+2jahKzjhend
imUBLttdn8SRFogxNcW+PEnVCZwKZx1eJoJ7tJh8XD0QgPaLi+jihXctjSN0s5U+h6Yy2+9pj3TL
ETvAeTF1Bqhcy/dVTFqBnIsJbehy1F2OI+LHhcWSe5kQAW4zLnCiYG2kbnpQ+n5nZ2RklgTQ/0bK
tnQEy0RslPeeDeOOZcOZbeW22RgcCXi/SChTWWFRncG5ni9/Ct+ruiIviuUEDdIRUQxiRlHvrxt+
X6jP21XsZuH8U8eEnA5lfecXqMIRyYFDt5ZxrG0PLBWrszTuABAOMc87afXUXEKM444MXmp3noJM
PNwmpEz5D7q8AkFSCSvzt2r/rqsjTe3d8GV6x8PA1jp4OL/ZOh+osBCoToo7jVnvEpetyOEsmY1g
55z8U2f8iYaCADd9Jo4six1aErh9hpztcF1sfRocqDCiAY0dJ5qR/BJFy7lDzdmUtuuO/UX7p2Bx
jd40d8oAvvYngtMB9dtbaZsk55vh62s1P5wPHXzn9efvEG+yh2Ykjkxkei+SOFzjSm1uQEwuW+SY
cu8fJOXt8mA+NzVKpFCUPKsngs/KibyIxhUREGxZ+0x915598hD36xuqFdrmRl3m0bGsm49PZuvG
R+VYA6qkrz46o6f3UdCiWN7nPgBQhFrg8oPkMMI1sPPVaFELtw3OzyRW+rWxgQRKCyJGMzok75lc
8oKWgmr41WY/sEy4xxcZT4d7c3Ks2tgLbQrIg1IsuYtsX6opB6dderTA6ESJ+pyhr3OcirE2HUIS
H04khJOT7Ng2OAwgjhxqNi6Nb3vPwBBVgvnej7hS+HNNeLr2Hy//foOlTHN0E5hfW8rYSmU1+qyZ
RXsrhNcFtEkixoUpyMr1sNOx31eI9RDH+dAfKfK71ej8a+yZ3dSn4bSJFiKtY3Uht+kpAyj+p1fv
1QpSSo7Ohtmn7FDOnWMvWHnpAoOPD9KmhknrA98S+pBdfWPMh8Mj4/ZDVjjUeCsrB6YQS0czrYbq
pjedkJRFiK1RMJhpUcl2ZTX/6/Z9cQw5Es9cKFB4tWSSY1+m/vz/OeN1z15tPnDB5RIfb05tdvbi
e5todbXJZ4R1Ui89i24hmlPG6U7i9AEvjou5iQJ8aH5uz3xIPLSxfKGXxyaSRLoP0qwAjgO+rsLc
gfHgsrNCvG+BONXGKRgYJNos+Lapu62GiVd7niFxkizVLDQnnH5rE+i4x9Hy4s55ukYx3DOQi9ym
Bd8B4LMNkG9ktUJGVC0+7wp9YtWD0F/uqbb2pGglqIZDLE00i23qv0CIdDgQPL2xO2ODEg24jf4k
j48SYshOiW3giOdVA1vgBROgSjU1ZYSo7t7y0rtsWmVBV6qVPhEeHG3XQz2YBqFXHMTD0bFIsWDP
heDMGRoWq3wN6O/j+WoGStp3gg93YLHN1kx3ZmL7Q1UAef8J9N06iCsYPYaoa72TV4E7KzHvyiZ2
1PZY4vihiy5XA/k3dIkHjpGqB1xK3thbgHoQzgKnEhlW5GwxUNpEB4L7UzxktvOTl04wxKMwavSP
/V5p8tqdFtay1r8Y5DThvx4uUuoFLSRc55d6RJnB2V7YAXjUMM0D5IM0LEDk74McEXYMTf2qnM7D
do1uG2kKusjN6NS1UuONvNtOPSVPK/GQtJnVbe3iPCn4Zo1TVMeQQMg8c5E2SwWNF8wBnqDINhQn
LLl/czi6jfJWp3hXMvd/4ku9lc6YTPuzXZdYUE3/GdUeQFkizrKfA28m4TCkl6FCz8H1riKT1viG
5m6EVstyk9OTArj+II1NHcuzp5lgbWuo621t96zRHS1uqqoQhGOpuVQhEYi0iDVm66181yEfiWlH
ueAKj7ub+uEnZ2UKeWeXI2kCABMq4GLo3WJidmwhLEFaHVhCgLDD5tWOzHtnC5gji/HQD43mlaWZ
Z2LkTqQKUTa4XDnPPPgIfG/6YVkzGWpZVzhooovi0Y93g3mW8yfV0u9cvB/UAywtdgj6mHDGv4sE
awD1uddznAgT52453b3xIl4gaI51DIOxmLI84Ywom3Eq30OjUk8tFqNC/KXag1k8hiQ/XS49dIFz
RHEsfLvi6CDkMRmWY6fXGC3/ybOfbBGvlpTZWrg6W3HD9R+Th0wytn3EsoIEHOQyr/WQD6z9QuiU
M9C9vXc8+5m3HJLNWNpqegRdJGwRE0QYX/96wRi2EDMf/ly0Yl0girpCfCAm52hsJD+9+74mleQg
UnhsVG3yCCnFBoRk374hh2inYP5cuoOJ8jTrrfKRS17msQrAsGUC2JSWtKsTwIrIv0q9+xTHF99/
PZuzCdF5r2/yzoGhL8u5Mv55DLY1TghZN4v3wlaitXYWDQSmiaclI7L3TCYrPu3U/IGUw4fTW3y7
FhV545T1kXsDzJCnFcuM+2DjDFZ7zGOPfqMAdPj6DjflZG+lt0XQ5wEug2rmaXCRZOGphlBlDMiD
ABQNd2GNhCmU+vX/zZPqAFNSmymrD9uNZvjjezwsphTDSxFRj4sP8or2tc52cQMjQqASyMAgi9LY
hBc5b2srqcYRx7NGTUNxKWl7Tm7R7uKwpfNPR5yZjKYZ7qm3p69oXoGefGGKstJoLIiyifq8tX5t
tvNhHUW8klgB9dWnHwRHd4P8hVJlnOEPZ6kSsZtBEY+FZA+nRzdgiH2AjxnjdpWM7B07Pigneiln
6/m44v/nKYNPT5Prnc3vk9Znmv6SdkEbL7rX2OVLX6hlZa28toGov7puf4OHbRC1rbBOQBzEPS4s
irCLQBQ4iDNj6rfqRWUFUbikMR07Y8dfZj38OIVAnGnqo9YehRkdLXHc638vWc2oapKzVW78573S
v6mz3YfJk3WiFNcivAp9gy3/EgrMo4v9fD8dqTC3itAGOjX+0nD6chf1zLRXt6MMjqm8WuBel32N
s69nyUXscPxyu9X0YCs3NLLA9GE8dP/0kSIxgK6/XZosAnTUOB+f9iOcBG2JwDqsb/cyyFgQb3al
LW/c72DaoKtCcPHeCBpzxM7Mjz97Q6qomz0TXD3C9bIdeEXo2m98FYVmHICYO7rR0R5Ap50T13yH
WRCyOcTUYWX0ARNNHmLMcHUGo+GClpmwyahLp8qeGLGyTN7lUBq3a3ExZhpqsiD9vWoRPxuienir
ALGkM+IZXbnNMwJUIzo/C87tTFsiRuRK3weKdZO9IxYDNRqqf+LNeuoAEn8+VXaHkOaSJbBlP5iE
ApB/BNW8fnsk29iuSK4UibUH5qik9B7FWQ4xbMJCnirxCDgKTB7zQiMmMkrhqjIUb5yDf0ByS4T+
SDNzXzmVml1AQLQ64SZRFI5706KIkYXxZPn9c9TysrbrV56LgkFFvG0jWc5K3/1LwL5VRTsVOq7+
9swFCihpN2sHLbXdrikqz/xuHmexI+UH+r/9SZknqal/AKLJQQbKIj4lzGRdnV8H1KziqqeI7WXE
mWqA9DfaSSs+gaO/0EQPo0en11zvwiK+lzcjeaN1WREovt2xWfe8oweSLre0WhhQrFP703CWwGt4
TUMmPKHrOgSmDePhCG9Ff95EG/2hv9xUKjSQ5z9issyDeS/N8AL0XwNfqP16WCc02CFwrvCqarVn
NX2ADENqJP3ldEwk3n1AvLJUOrktkWCTL70osKvYG5T7n0HAxgz6pIKL8fY+yrOAMuOhcf/eVLyv
wIO20Kg0ll7WkdMtoK74NWOR42WR3F81QwgK3o4NSR/2Tq86aDnTicis0/3tHBKA9JZjlkWdc+hJ
iN5xUV+pgKwP0aWmUP6SE1US0qjHwIo/5cGXnbWtVWPTJLDVWRwCHffsU9NzrTxsamb8RpZuvAYD
zmG7J3WBpbGhj06TMfKGSCyiGhfbBslC5qDLlxKS+7LmDe0DMyaaxLUzzrMpc6p7Q9A/3ui+5reD
VnGja5dYWS87h+qGo/ArXFJkW8AlkQQ4DCGKdY/biFy7g7ukvfWCAkjUkrwp9iyRDFi9N9SPvF80
SeqhO0DVDtALV3W748Sk2LWSmJjMS65XNDbIoypm3SQiHdBw1xNU2ozqo9k0OStlWnridXvk6H0G
ISGpK8OK2LD3mtdO9kpR//tpnk+oRtbQg+IK/vVf76t6ulqjtLlPJRFGP+yV8uvqWvQXTWZk20ej
R2skyToSb3K7FI3H24FHR5S7h/W7FmNn5vf7/k3SQT1Wq9KbkXnUiMPKZml+sfBxzRJRI+K94lo0
WLcG7xMp+La7PFT96kakIBELAVcmuluMtpjR5ljw3DHPh2TvSQ+vtZ5BLFquTqDiNv+Lmh5CATkf
F5CIuW4mnsdVpIw0bE2PJUqXfZ8IKpqc5Mqk64DfEZOzfz41Mus3lZLPfLD7S3bVp7cqUEgVt2Gn
GLLTaZVIlCke5PN6g+UTCnlPrRFV4VY6ajhFHqQZyLO95LzMM/ZBRY6QsGqtombRqyPNSveVPUUk
NFjWg79A+2mp3thEYBekvRgNtVqER18utLqtlRTVkQ4Yn2F2qpKniqeaiXS8/Q+3GLG2zRNy0P/y
NdtalMBMQWCWqAPPlCW0MoxlBPTZ3hqH3vezH9TjtbOOjCUfypbetjL09i2+A4Gm6DDX7quhMtEF
yaq0A4OhnGYOsx1Al8FbyiZtFXFUiBBuazyd737Z3DVSiOCM27LnP7QlGTf9F2u4zp/0CFFKbeqF
a3hr2N4GKT4XM3us7ICcJnTrWQ7VWdorU4qjI6p36wN7WiF7djAdEpGmBetbBIoXhQ9eDb2dOMHw
FX1tM861HUSioL0UfqLvS02eyPCqZQ7il6XLP9FFnvaa072/i7QnjSOH5ReyV6Fj9Jq1hbUqN5HT
ekdW0FyfF6luqeBbRYR9/VsgN5xI6iELe/UXRyb9qoj8l3tK4f1swEyTnQNg/dysO4i8izVBLZti
rQEFd7hgB16pJKAk61TZlV2fBQ33zBx2lHGyV1fJnv7NTfcY5DiAudGJ9V3zpu4Jk+K0Dpb1hL88
sTkRh3y4mC6Ek33hjCsKE+OUPxAWVzz/7IJm7p50ievNoCKp0R12ijMAvLykRT2B5vsy3w+cgeWl
oFVuO0RNImf9QQoMcHqILyXxFlkM2b3uJH2RwG+NBNQOCMRoDMam02ra2kigMKgsRqyYxql0fpFK
PKcUFO+UJSWrEU9jzKxAq4BB2mWBZU0MeffP9FZgvfFsFheZPiEHqjIPXn+FunOwqVg5D75U/lZf
dqp0s0eSzT484Ke2LmcE4de8r7hgp67ciPcmqmN0ygMJUkBSSawOxOti2rsGsYCbezIYig+99xbO
CrYJaWH52qfXV57CP35oCWh+EEk0z2DTV090UYc/AC0S9/uZRAcW7+P9XWvR5XbCvSivQiJ9QmXL
RbiMDxCcoOb14gGRNYWPsklo4+R8JtlwKoBVJJOGSA9z0ONPFU3F146iAJ7gnU4+cC6wpRR8aC9v
zNuLmJGV7KvVcvNiKWvrZnSR82FcfDEXDzdSwz8YfZU8ic8lDGm/ZeKtCJ+XChxh6nI8lnIZFs9k
Sdw2ZimdBNkD9e7vImIv3Di3d1DQmzIoYIadIdNrsd9QFbgdhQNcOAaCNFcUN5+fLY1KPema/oI4
e8N+ElwQaoEssunttu6QVEnv65VavBvB1SELZtyg1fyEEIiZNVav4zNxuqldsSpe2xVM245LOIVB
dXUiea3tfI/K7vSUiW4lgKZLdDwmxRfXU72VoZVHsVu6WYkoIRnAA3lUzUSipcrUYDr9e8kod0oH
hftY3jUF8h8Ao6i4MU1AChSKYxzjMhwCpOJkH5TT5XJmYxuEWPWLrj5hH3D3cYty5uCOmtRXTyt+
VzChUZYh1HNN5175pKO1YaCTYCvB0tZ45Mjnh1F8l1ZwCk/MM+sht0BheVULLtUdzZZt9rXgr8O5
iW0xQMwDqu8M5zyWoP42r/zhHwCwxLeAaN8ldJlY+jhIDykB40lUYhytkzl30xDN+2cIXHV/h7mP
CmE+NBTXjxzicKF000PEv1Jez56bkXr6o1CxDirvSJI+cSUcnv/wzaZKlkLDkqPwejTDSxjQJoOv
tRPorAn40stOVIZML+ck+lzaqG1IxR+gvM5AgGr9HDOrLfj7jsva2M2oKBshUWWJkz93hVjfZnbn
9aSKsnFQoPqqjzhsL5iiaakLKrnqSU6dPDnV2EpTfki/nrMCpIhe274RkrEKOn+50MvLni3D1i5L
nw+ttj/cphN3Da1UM7WT+5AJ24QDedmP9duZLP9E/ROeHjEvsO/zcpX6D29WQgw/dwPG1vs8UsyT
/ueEUsWyD4JttyQBW3cUhm12gPUW2BLdIX2KSEQbn7EMS96Y8sU4Lg4wc0CEFG4JsKQsPILSiRHE
w1TXD1VawByih0krfU3JC8ae4A0zHsaQnwehXbnz6eu4cDKxKm1M48p24cI2nGjIOQuJ/DSEwPF8
QMMQfmZnj7IVj+8qWb9StuYR5aeU6vaZ5YueNCD++ao7xDhUER4mP7CaIKLm+te8mR9oSOvCypi0
9EJsu4gALtbYy56xqQJX8wqgM26tygK0W72+mwKpz8GUwffNYnE4jCWgPicAZn73hEL7HwxIA/fe
+U+t319MpY6c7VBh0DBMLXez58+cg41ByFcpJXTAJy7Rk53Kg4ySQf14dqjMXBLHx8Jyh9qN+wvQ
CxTmk15KstPHiuwaA6a6t7VtQ167fsJCDSAYjKmdPHpk1R2cXSxoT6D9EKPmh8LB80mhzfRGQccb
GpYLbjaikwqfAHmNPqoTmGD4lUlyNjaWb9dgQcRmbj5oT9Og767kavK9ukc7Mzd3sGUGAaxCRa4x
ChvBaIGcoS8znPX7GV5TDUYNMCLCOCe6xsUKgQ72grPae0FFS5t1961kKcXLdFdvg85GzlkZi0Nx
YRpg/cRogQ+X+O15J/ckVGXyhSXEq4QRJLBnDurI8SyDSHyUe9JqLklTe0/QFSktUfwmmaDrjDF3
N3xVqq/UU3eBKTeb2feYLLvZXuAC3l30ciW8Nuk5Oat6y3zRqnmhl4z6+boPlz1uwM/hoZLp21d2
s6d5hrWqUib+IT3tdEIwPHgtSlbUkqgmkWBjhWpmx1Gffo3aDau2z7XGJb7Nx/ZYmY1qDlnUS1kH
hibHha1UzA6POVZ/iUrMVyOnW7txjRpX8ZOdgwfd0Mkl1aC26yNzB+aXOIUl5V/zI31SleLK64xG
GGvrFZNf9GgLi/IWJwLbo1ZTkfIknUJcNPwqWcCTr5Ir6/5EJw+v2THUvHlDOUQIUh/KVl9yBLrR
L+dIw1LMDHQc/KRlocISe5wcplHqNjWGpQRs5ew6Ea20sMNYzD+77dTsffklgYEou3vgdDTquKR/
2RgIgf1sgkn4ffFNBoEcVsLjRjlQQrAjhAfMC9uxhS2AfBsa4Mo2tGMsUT+dDDmTLA6Tj3+4CLGn
SFgBG/sdoMdqTzk1IV5AovNEbEUtooPkzcEir1Sb95DQgEjcaPKGxerB7pA2TanCNC9Sl8gHBI6e
bF1APtdejhqDH08InYp9WlP9rPCCQuUSnuY2t/ZxtVrmYfkrg9cQFXwRs/16WYTQ2ZdYKs5nlOI/
Q7pX734nPu8Jh5eejYSInudf45/Mdim9NrsXLQ/2d4yieFrD46S1/Sw4LvRfS0PE6+2MjAMSdy5s
qg3bXnc/oKenVYtuWULV0oMBc3GwCW38AQrwPCBxR2Uo+sx9ySNnRkIUr7chkIderXO1ZjIQxQEq
DQ0sgWXfL66oEVlb1ovtdCMYMIZ4sCIjNmamTBBEY7FIWLb2onDmkYhMZmS06duAx61pQ4rqlZRV
/IIprv4FhaRR62FQjQdGJDqbXRtUoXJhAbv4vSYL+o/y8O729WEJ+9BWk+2rAs3f1zmQOn7qCIF/
Pm1OjwCKioVKcmKXWr8Gc9ZADDYzmWNyGRkPDASPgu96uob4CBo3KIGY/+YjSQumQcULWamTZuLd
P+/N4b7yo6eFhiGEDv6/keros6exOMU5WtMlmZj7yNoush1KuYv4nIyEPBIpC5xv0NRvY59vr9s5
G2+08YcbNFKiRVHp2/T+pzXoLx0Xe63Myk2W3WuBAucUHFtQqluqdqOEhRvqScTTmp8tAuJHKR2R
MgTC/6mnb4HrdWTW2bSKuhkvTtoSXyvFUg6JpuAs5fEQGZ50gc3V3TLUjeUrI+Kg5kwj8fkMjsXl
8+x7gks4+Yr66FCSH9XDqGgmErEr3ysXRbf6oUll190v12TV2+OVYtInJxHQD3ou/nDZ7EgFSErB
YkvMKKiDixdPmSm9ckWaaPbZVcPg2rUuDpal9ceqm3XZJ3+WEoJWkJuggGQYVyEuetZbSpk8kdbW
CmgPm7LZgq1ynHFWPtJzrPAjZyIz1HDSNUAiubixDtvFrrxp3qLCktoREA2UzN+Z4sFrKKDipPE0
vD0V97GBAjXvh0rxdEvNbp8jKITI4CRf5OW7VFITQz2VCqjSDyArVanUIebaKP/+aQ1uFOJf1Efl
87am+WLq7PtCLgaOQUgelV42GqArXpnHguArE9by7h6PC2+zWsnoGXT1ORjxfXQgCcE8T1PUcJFB
eik84iNd5Q2tKbVHZx7tyNibvXknZ9gMYQmjg7HTnbB8KeajLNOfNUAl7cu4r3zbFodapcVVCdny
7RZIMG2T/x6xPUDjZn/qHLNZIus0Ef+brvua9abyWiJ7ztoXMljc1j+csQoT8HBVPNgpHM6edsNd
2KdCbYP/7nxia7pM27AyY8AwEAgX/gK5Llc41rOz8RONzksg05+MtvCcjbtWySxVU6AQWd+5oWtV
RFyrXjO/eTcfAGjQk/ZZ1fA151h1iW7mqGbpzolLfyD/ED9oHwAP2s3EJfNucwhZWB68Ym996bEX
42+l+AA2xeiLcJ7x+LfQ0v7cymnwfuKlpwCMo6z6BnYiFNXHCAL3TiTlJyCqNh4nMhEXLoYkG8p1
aDCEPZJNTc1IqbPYLScnGFU9CgZ27cgiNEomlkFlpl9ahDg6Jubk/bMF9Es8aplFuyZAsIAAEYqK
n/aRGDsMOZDWPraBwbH+BqU2cIf7SwI9U4brzDAOkABCUqTLNiWEEm2dmQqUqDf7vrA1Po0Y+GgP
QorhenAOmvmzTE6+oFdo5ObbJiN+5PYOt3NP+B0rsfh4VrOOTL05V1JghHeoIdNei39+cxp12VZg
lr+IRgVnRKDBUyTaDUnx6q/QpoJIgw4/M7XSwXmrXu8US1kEjvYHbY8kkZGNye6CSom+j6/W0FNx
qmWWqz2AQ/s1Xb1TSdICZbPmAMRbDai+F7UWtfrXc0ACuC/FFI6tBuafA22Ux7Vvcv83ryuSUyWP
DtISuWN7DNu6gjUpWga7EA2fAaUZBsjxFefEZwqTeZ2AucadVbgIlEHZ4brS4YGyLDaASidp3cQn
g75G9mCyT06WeZR4pcd+KKCXp5w+g8zj6JjriQ5dnOTiLptTdq5mVpYq+mm0ZIJMoS4mG7bacn2Q
sXNBKcUr6KFH1uhyypJFd0pf6lTKxKOMvJXqmswZTWrXm+qT81sSktgNdLYpVA+yJKVET0wWU9LI
a0CFw6SBc5L2NNOsyszlMfgL3yC/mkBDkqh4A2Py1ji4xnnrWTgofklhVnLORjvAKZ9WALHMcJ3U
Z5iJaQx4r1t/1q/TLBiSUMBbLHPvTAQv+OiyhvYBZJ4jVehfCRSydbXeCnXi4ThfQe0gkbjXgd/C
NR4ZcOBJJnjMkqVCh4+YyXO3WFzBh7mMaGZVAYKN4nmxT0z4ZC0rwjSSKa39HHVj+AJWryYm2jTB
a03G95Mv6QsiM9/nc5Z7qXiwyHMG0gQFkVrMVZ/aAzk2mspe0jOIIe3d6AxZw7l+9CjnI9Ylk7Qs
vBvVvAZgD+yWf6w9bt5GpCP0xjjQx6VKhYYjB7K1q8piPFLibuB+TVf01s/tCHMReFuinckwE2FN
XiwfQRyHnmfADlcde4vCq+BMdqZ9yWn0vrEFQTh4bF6ErTu54BF8Ff1xnBPdx/8CgPlR5x/Oj2Kx
TdsBzuBiuoSnU00urY3LKh6Cx22l2gVXQfscXQowEDBlwbbjhVMtuwpk8k4H2gTz/LyDZ1I8IYeN
WaH2XaRqaykNUqDvyxybE1fVk2IxWICz+akfAjOR0bJNVax0cjhBt71tsaCVXFTQlLqhZTL72FKc
zbZfDbNWTcz6rGeP+S6GHBO4cJ2ylg8f8m791QM6E6teJbtkC5vGFAqW7pALA5k/MTgOVZ6bt1or
mzC0QQbIQ352t5IaEemBvqK4AX0eOOMf2+SYqDBxlOJxfp9yrNsv1sWgBAMgVFlkrXoMBam0KQL9
TdtUJTDGG6+ym+/xZR3ExgbkROSBjtSHLcHyKx5VkzzTJU3ctZvtrWwzvIrmG9RIsjAONFcQy9Ya
VjTtBr7UfgQgTTx0FVB3QPHCoyjvEbiqTfT8lR9qlKu/QsLbj8USic3SdhOEb2xN4kjowmBR/Fa9
j9XDJnVMjwh0tDl1G24dvKgskXuHL0d+g/x8D5bYpWwmWnsFS5jNyOu8EPngtJTXV667HAMSy7iA
XKwBqODZSesR6IDr2cesv9ZW7Vn/F5O2iFwIDMVWbNgh6pQT+eYhX9dC9sE4ty2ZVRC3tUrLbTLg
guGGD1HdWvNt8aixtvc8FXv/clcpPF3yw/aPh3Q4+VOV+50+EWL/UzvRpRJVMhU+Df6fZl0YLvkU
0GeesxeQfxCDthKvJHk1cbvOm+81rLvJQecqHt7uv66WdCJ/03MyASRaWPQPM0AyOahk2m2uuljE
rhKsMV9e7nA9/MO+i08bfPWHwlxxvy1r7EjWitZIwJKbC4kJRtJt7uB2xPMNaxbYFz0JRfVozYt8
yQ/Aqt2rNkItJtPhSVza5XIeTUjPyFv6QtXKgkRiEBbSnbSJ0xkioo7lKzlmMfFDb+zOaVH1xpAS
HI75Q86rrRKtSVfutjpiUnYpT26mUoLgzDcPNXaPrEZKr3MUIgpp7205MiSpAB6+ldzB2nEfcGv8
KvFbMIxhj8230j6l3xepdVef3KjcDCGTgXT/NjTOuXYVwLS3UbndimxEQ5f1Z7E/DXljcCOkb+3m
aq440X24Hi7M8enPuxyxJlDgTWA8kNGd/RdtQPKyka9QIfsgaRjlSGuO1C9qbCI9xPAOAInw4qsx
dbs9KcbPAvO1c7/ArMLZCKI3mfrC6jwa5uPZP2ebUIqO74c2iYM9M77aB/A/61SjaxBlZ6dwcNVf
illam5KyWR8fgmYH+12lww3miKhApVd9qLk7qUYdsAgjKKJ6Vf8cFwtykhhOWs9cE5Yw1sjpCqeo
CLF2X1wlIPbiWszmtkma9WcIZkc6B3bZYo6Wac83F+TU8cLsufPsO2l2SvFr8Cs8mBzpPy9P0iGI
8Wh2vAydnlM0hlgTW7703yste0Wr4s4aKK0YLKA84cD9euy+wUmiIx5cMIuzQXi4oaAeJ78d1EJr
EhuZYZ6+xXlXQ0J1Bcq01+IjIrbBje5+EOhldqGapXnMzCuZ9/z5ZtR7wmolbgv/X4q34RCVyouz
NT/ZcsC1pzWo/iNSvH9sMky1EdwNBDACJ3x8exN9PugkgvqWX6g5xEyCQcgeyhwc/gkO/X6EEA2d
3zLO/nrngl7305FqUUf9ihXjmlVzY/ZOiFo8qz9EyNHCL0XssC8OVKKpideAz7hYg3V7vtWpV8Qo
2tO5u9n31g93spYG5DfYIctJAX0KGp454USonnpMWnmCTzvsqdsefd8wdD56Sz2we2itH8d/72n1
nc4IZWISFY4fxwaAcJWCn32/K906itNYSuoN8kk1GgBRj2cwdVpon4K3jSiR2FpzVHkwquPuGs7s
YJ5ZJzSWxr9h+4SUnjUXBJv4LXgYBK9ky8i1Gm0EJbWCTgx6IbHA6Csle8L8M/kNJw3sey1AaSWx
w2zQqU4L0mWXj7c3HtLGbeGB3MEcaP0o3UbfO33/1JKAx9duadDlEx9oC/YXwUWxfrsDWD2qCuqM
YsbJufyzjZhM5dX9qKZm66fJ8r41owqifAEbKSVQAqrZxQRz4dwvp8Z00YW+gVDB3MZPB+QPLbWH
N/3LCNuBkruBkLrNpuA7hi5+U1bvpJE2/IsETMV8nITPtwdTcwmlo83sWZo51OdAHwj/9x2GK5bL
ADQafigYqsfAefWdA0mbRiMkSleJlm1CwSPj0zbNp7mpeosXgiW8QE+hkd3SAkSkE2xKHhyj3LMC
oJdb3lhTCxGVuMYloGmOwE/ZLstsGIqmO4aAufO13YdCS0JOS3Z5k/tD+lC2/DHYxAQrjNqbX9I7
/3WB8uDSByU8YhdhGiHIIPOJ7k1v7dcvl1a7ER3qogXW7/6XwNxrq+u+CfHA3GVX2H8jcBc01793
5e0budi19+xhjr/OGqg8v09eQbqPjpyD9E4zSxzzKPz/rgdPn6bGmR9I8O94t0PffRFy0+bZDv5m
TQkN6TRpVXABQb8xsiTDXBS/0tmwzjUFxvFtNm8ASeGb8pMKJNRDS5/Gvz+eVLPc70H0JmeuPoKe
o/wURrPhCW4dClTUdP8a76IeTh+8Kvj8wFy4TtTED/NdMHj4Ne8sBadGkm7CcLh8nJQn7Q35iYqz
0MIB4My4WlTRNQJVhgM9b2oiX9kzkC4HTdwmZmWsp+rHnVFld7M4/tZczADbdP+wJP53bLFtMoMn
U8sATZqvIVhwy0hlL0DSUVIyaan1LdR0hlg9QwYMQfCu7n6LVbChd9pq0tOhH7KXtPqevC0jWkNl
tgSFMbpLLr39Wfj4OZTZqYw2Umb5hhUTFc6pyDl7byzAHv7dsnbZwvSEp/HiKLIJFvaEKCH52+59
Kv9gLnL45/xfLPCwQryV4T5XgFfdN99uWUalbGxP8KtQoCS6UNjyYNGiVYCtKjEkRxeP+OsTJF6S
zAq9pki/4jXO7nHAzeZyQKUtfBP6xt1+QY9TiyG4JXcDG0u2EwGJN9Dy/xIu0ffPkCLIBY8UK9bE
ZVXjpEgGpZqt9oJzICZ2zf8/h0ofvT1+edmTYKw/AqdbBdbpPS1z6BpBDpCHMl0cnU1udwLWO777
Ijp3cQELOhI4IjPTjAFdD4MArhpUdwBjxRg33jKbeJLtEVT5SiiZibcs+N0biYwl49Srl9Hh8JFN
gOCfR0pgeACMwjyXX9U8BpGWjK0ekptDqPQFyun27Du9HHnYD2doxFfSsvKfF4bjL7gAauCIfH9g
Jj3MisLEbxQf2ZWW4OqQHskpFbjIwOQxG2FU9Loq2CZI/8Iyx3Mprnk1537W5j59fWr8j3XAKzq5
DscjRwB61nBKDb4CitC1HYZBhxN7qv5RYBM8R6xhgniM/DbI70VGGBHAZ1nbc8tfeYilA4mV+iYm
46azDsGKJdklq388wKJ1f3FTD1uM/mU8FMaAO0Fu3qafj/zlVuZ/cdga2dHzQw4eZnXYQkdiBL8g
Lwp4/jOfvw9kJFX5vISZDGqJlzExTM/DK+rgEpYTC2yNceRIwrBp2M4gOvJAPvHdef63gJJf3Klv
v1h1eBmZgoOLLRu6T0KVdHWR4bF4DKrq2Snp2T24ymDDoAn2N45Ic8WSEgEPvJJr6/YF8yvcAl+e
3O+P+PJDTSix1P1O3Nhkn9CWzbFruZi+fjTuQwl1itGOOMzpuWxXfDj1muN6MKpf4+LHlXH2XOFY
G2p9dtWUpVLpiw+r9qI14PAJ3iCoAF9jsaemPOkfTtC/4n9FC/61QLt189Ze6bWcy+LNsCIV7BXP
aH2vAF/w/iTDWOlAwSc/sBvHG37nqVwaLBxsQHVsusw1FztHnra6GpcjZ0jKgFMeEyZXZdmEXBq+
zpLpE1ehAgUxQQZ2yvbo1OMzAI9MDbTnwGAlgP5psJDV0O/GOpwSICNxEL4xH+RkZ7Iq8yVtzw52
LCxlKJhS52cZdxDAldAuiCgdRcJ4ev7ffKDGvSk7mhq4aFO+yGJ4THsdbnTMU98lScsFmJX1WY/n
Pf1ZSyn/jjvRvmL1c1gDDeWX4u/J8SjBq6djIFcpfK9tPxmikm+rRTIyK5WvL4sfBc1S1xe7BdqW
ZrpE92exkWHRqeew2+KnDCthRZWtY4Sube63jEHTyRf8p4+utXajkpdqRNsssVvfNAIlLYH2+s+7
cpepDGbn7ps5XgPd4XNXSduuZ8uz8grePjnSE7Cs8WLPks89JZNakWdhMBi6ubzh6L18BVdRYRq6
/rDPn9BFxoBlO5QuqVXA4zrAvnByJpqX6Zic1bAF4VE1L5Thnp/mwvFi+44Pb+FNcxfVzdRRIqPy
dOYtsX8GmUX0pZ4dS/CrqlFDH2p6W4lPfObgL6CP8anIYMJHxKs6Dr0CvggsA/yIVuiSxNYj611R
at6TzpXpkuYYyltn79MRBqw7O87TrWjTxjJBNaq9P09Sw2b1ZQpDx04fddMrQhsaxF9EKDRvdfqS
lLw4jPtYN9+/NjXmK9C0DalVAcA8dNJId6RmSFv2G6kV5ak7ekcAceJ2ziGA0RZpQP2yZ+9siRk7
FxP6ctnCqxsMgBezyeBK/C9HYfJaBN+cy9qyraVfTy3q3C2iEPqmD5W3CKRIjOjnXHiWTzpjrZb/
kmLeEO/hODTllL1E/bizeUT/nmKNL0L2iujvYSqCD10aq2VYiRfu99rW8YrLAL5UtZwA2zDa8aeH
VwSIAZJ11S6jvn/gjx7/9WkA2At808wk8wtFhtMgBgFZcIN3EluHpsl4JX+ORb45uec4+Ws40mrA
maI2twcegRYWpV3u1UyiWLRPryn/aTZyzPHSQ7oilETWJ626fGzFmLO6hbeskQQTgzfceoWmNv3y
ogmuSJy3C8ct9fUwFQGh8sz/rcGifP5Orp4pSRbQAqYthGLW9xoG4RhhtUW97p203IBiVxg5mZcF
D97+xI9ZF08+Vg8NNxl0jRXsqbog64cNhyM6KGeLBouzF8OnsH+tB46m2wyGXM6qtUz8QdaGWTSx
vx0IIJKTSXY73p38UquAHdKEQpgF6Pkwrjme7df9wcuTl1c+IDcDWgbXIbcGD3BnlCAH6vkvcd7/
vHXbvCoGJP8zqhK2/bPkFxxVobKN3AADT4MI5qcu/sqYRkFMG/ZM+/nb/DPUKiJecimQzxMjM4mv
fgiGTvu5CdsHqSd0U/r1SooOkyQCTFMAv/H0vZNfl0rDm3nLqDXlNNkFm5TiwBXXPDncZOn8bDqZ
uZzpJLppSzww6WglA801UHP0FtFdV9yl8wUIZlro6ksiis907aXwQ6B7mGyJ6HiowxtPzlUamEdV
04FZe0MQlktdXuFP3JiR0aAHbl5Az5/IEuumWU2z4gWj/t3XMMd4Cj9qgADIryn0+4hgAVnVSQk5
1v3ykwe1EkGL8nFgAj7+G4ZImZhI2sY7RLA6R5U+y5aD3t77A6PvpBmwbV/LbKLuj1GbF3qF/Kyu
nOp5uaBnYVNVjvsiwr+cHTuWBBEEp3YrtRSwHZ+t2kP8fsKRPOY5XQR3sBrgsepxmjXbNa2Bonj+
XdwpBLk1m8Wv1YGWrFQwvgB59z1bClTOavqrwm1jc4T/rJnag2N1o9A6s1Wy2BoXCWKrYq6VbDCC
o33adU/23liRGb4vipCfuLqmHm2DW8e10nAj4SudE/JeKYHYoPXpcV5Ck2yIid2maoudIKylMRGz
PPCriYxAlJ51ZFEzYTQye7DF1cEJvLMaHG6s+fAt2zTht0wklpVnkRE67zMObmgHdun7UdabX1nu
9Z7HkpG5I2foHhzTX6PX+fXdv5+b3O5gfv64FYuB+L9nQotpZD+7vUpxK0Y3Z8wT7CakxCqstkTH
X0TNutVVebBmE9GCsBG+jj/AZtoR/4TajjzdmzPN2hBYZYADiyrIAXdr4kFRdTJVhcMnNx/Dtv5Y
hb7x5O/vuZVTHPqrJu840pxae6AyHI+RSV08rLVr+nBgDNnuxfSSgETI7acVZt675SLzXvuxGkz8
yC0B4nqPGPZzJoMamAzfs8GZnoSK485wI9JaZKGy+uuGksHJCybfLQYXu7G7mk4ABTDwa7p3LNyf
dHRiCENdno0uq2dbbwST25Dn7WIyoUt2F8WFCxYvzLjZ6V7PqZz+6Ovr8ABiDTJ+JIpHC7y3tOWw
DM9tMmmv/MDzSnNXeq988fKUTnqLdg5z1V2xnQNBwdaqrt0ai/KsRPcmtxSUmDfMVh5QE0mWAztl
brl+k6Hlu/vzHQvn6Bj9z12VSKATj7SuglP65y5RyDnPpC2qSzhG2OVJ8SJYr2oJeeSfu9KjYULA
juHhu84d+OXCZZdpCBLI/co2hAm999o+OVHwz2H8aMR+Pb2hL3+iXIN0CG5hF82xTfREJIJgnaNy
O/uOFIoSJJ4IgpynwvRVyKJ71uH7OA5wsLRd+K99wb89ixmB19jGV7FEac8p24a+z3GgjwUs3X/q
OQ/Xa9p45AV/Zh7hSrTcD4rPdAMdi0BnMU97ywBIVB2aFmZMQSUpJsxqqLw9S1NSZU2y8gq6f/Y9
Pls9GmXXHbUafJ7nkWKIlyFUc8lrk33IC/fLqeHnOQ1nrvxSlJ0MAmygLOfuNbxvdkGbu44R4srB
ooy+e9Vm94Pj3OdEYBxiJ76DD/5Srv2yrLBHaSJ1fTvU2LhMOOvzCoM1fFCwyHCUcDSATC8iKF7T
BTfGKWHirQVRLQenXHPLK4UCDhR9fTJq4DXu51YQYTry46FKFiafXnOODDArFv8SXt845RZyNaBK
JqJ9JBCVuAMQ/OPoGhz2LkXqm8buHugapTaex9VcUgT4NH8oAmnMmodfvG/MziP8jcvtYbNjIyxA
xzs1fiStVvEoMRVa7bw5UhVqKdE0Fv0GqcoJItu+8K3QTxTIQ1xnXfwuESgydDh7kAMwPcmhxcMX
/rV7p3VcHnOGYZee3+shkWS9uuYpJXdKxwS6LFiUVjd/auTzSd2diJV19JcPOwNCAFqW0V0EZOgx
VAfvg94pTEhkZnku/UKX+k+iQkMqFDMT/rTl3XiC5LGCL0rt50hMI4a01oG4BnaDxRAG2pZSyObH
Kx0seJPlbtf4kpfjB7vbQYG0/BezE4vpI1I6CTVIBs4orjxiAhsxouC/rO9cOP/SttboCTRUdcs4
TTHvN0qzQi3hwzgegdOC6kIqQ9RBUPjqH/+y0JMGr4XgAZw1YaHvzWfqXftM9QaNVKC7ULosje1X
ws8IQvVEKql7Ap1xeLumu5EefU8jlWvQy2Pm/dRVPq2S/pIeHPH6/rcn58JO50KinsnzkNOCQc9l
qbSEL0K0iDH3BjtczvFN+OtNCYnPMLmvp3slCR7TGKTs3HViuUmTr4B6Hoet6BKhyosxzSUE1owm
rQQ2oBItzvi9kEwSMOYQlm7nLW/LJAl17vPJ39IJ2iLVDg1bAsIU7iduv3HZe6gRGq4aO8tnGyz6
afS0BNYaRVjMiUDHr5vXq1DrlLDfdPrQmBmq3aSWUY6YaIGfl0mOpByxXK3RgTX66EkYD9TDDUjz
PBmAIxCNmZWF+t9d0PyokxUNxNS2qdaHjGj1ZKoXhLEmuEZ7QFMcAq597HoazdaHbm15Juql1S41
bnyElzeL0L5XpeRWsTVdaHF4nbyuiCSMMYGlDqKXIzLfH63rMkBd4F6bLLbKkhEvW0JEl40RGyNh
/+8OOZ2wV8+HiGVvwXil9d4ch3BSTqHZO74vLSNLqKxtLKOS3tcI6Dk3LBajDUsG7Tjogkod5131
ntiIAwcc86A/nMXquXS+ZBPhaCHU6NNxu+TVOHqaV6bDx6IS3VeSXMM28JBOmAiR8hTfbJ4+bnEZ
S4zHvBDrARSefzDDhSaaHaKEAluxE9unwNcWt4Nrd5soZbmR6CQGqYV1A9LPoO2c5QEBOtOMxsTx
af5vrMrxXPMS0h2ObAnx5687bZk0sILDVFxlxooiCl5EE/+iyqeQo1CqviettdH5aeLadpTv6XLY
o+3vvqsnU5bfND9amqb3QfQzM8O6ajEF8HgyV/ZWklsKkNHexFSWQ7FWX2XrcYeCwX+3KdZZlBav
ALILaIYE6BgV2s0UmI756ByIq5gTerek78LgWh5UDeYrBNAJCqOo621crEurx7uUDB5JBmMKDRO0
7XxA+foZ2v6cuYQdruFENIOGUHMF0y/dqeQLJMj/LZi5odWWx97FnYsxdxU1gKuQLx6ZZVyFYhNm
ejEK/KHdMpUvcDiQaCIfHYnwuNTWMsZwkeWR2c7J2k0EJJyQ9M9sNn9kcomxqqYymziW+qstJi8r
yPisKW2R86QHJONFXIQSnT1Ao6jgJIZUYMNaRhA35BI0i5q8tKmpccJW3UazwJEVZ77xpnXO7ssy
rWuAG2gz+L5uC7VIwMl56Mft2BmQvbKPrj55JmYJADKbd9Jy+rORvdGklrZoSzzeenf+yzmonGTb
0KzJ1pSRAEtGDLZkU3piLXThVc5VaRhUmazcByBpdtZrsLX5+VWo18qOkwnGkpyYxPXsPEdnhEAX
oZM6hAUhQ7Im1Ltj1h6d5MOJDj2iv9RzgdjGWwquCbU1wDM7zVWb/5xMgsvDP6PTwqqBfJhu6Y9c
bvABpyx+NQPCQWEh72BjTWrbAEc4iEyb8UFekFbqxuOpzhPpCFblz3nQR7mAJiyk7PKsNRQaQY2y
O9o1b/zL4WGBn5BcB5ZByC6qjdFKv16xOlguq2/pkZJ8KAkzJeeOfMXePWDvN6L2VdLozFo2E62a
zoXDQChUhmdmRU76NIIBww7eV7SnIERkuaaeeXiGYASoJE3IAzVGDgC4GwjlnmjvjWZ57EXIfgzd
Uq3hh6JJGds0rfEUNyWoWaqqy59HpCct4DjkjBa4wC/4gT+ZRXPDzg2PYjy0MIUv7X2zCYmvbngD
yBJgFqwZBoIh5RDwc2GtN13SPX6inBWgzP7Gjemz/Um1LYDhkoNV8nyQJVJq5Q6T86rbO8/7hpL3
kjGF+r/ieVbaKAB3TvigPlSEPKrFuhhRCCIhad+DK45asg1Hm5C4RDvNG4/TuNz31/JtW9iswcgJ
XaeQcqiRfZbY5bCjETKmzWMzYfikYYD/GDisAONOtvsLvEsRz3Fn7Kjet6uEq0k/JM4LfuWaHOY1
OzFBUzUUyw61DDZN24yu3Ce61QcQd8krJuf5s7Dd2/MGpkmC5g3AdnKirHv0eecfSCfc7k7vcm0a
aFPkefByfbjmHWgC9pbdkc1gQ0gNQj9CntCQAXCl5caCj0Ris/1aw7m9YE0XnrqlwD6II1LVaScg
9Vkp201PNSulNsOhengikdc05fWtw3Fvpvrv8ieB2Ya2Dx1wcxGvs0NB5vvRnEgDZGuoL1mpTJgW
3EouW0PkEJkH386Wh79Zlbnw3euz5uuVpnYvmpvTOaOGMCW/r51nLioSbDZaYV0fN7Y+cxmabZLy
meaPzLETDXpQqZnprUI7fRZlmIgvjnu++5BzF4/OgGIHu5+vjcmF2lZ7AB309MJsaHWyNWRACu1y
EpywlHCTS0AvYAZ4oDNwKiV6G4O6LXmQ6zTNtNiDYPv/RKz+s7qgMSxcq6RjqP+DwKe2SIULJz5k
o/yDnkbOTRBWcQ10pBvAtDvbeRYr8g2B+mS24RzxsU1gP0GMX9vNJF7dQbKzqbQXJU68uWIovv4k
cwcPjmIYOJA3+fluU+FUdqZW8Pv60YcZtGodArMsdyeRH9TU8UAX3J5U+DxZ01HLunfDi7SyGvVq
7e/QKQ0g9az9VspLHc42nkgZ4+YJ59dSSkjv4RVrKmLbs+1gBD0cYd5/M9l+sOklqO6ZhQdnGuLU
GlppOz2YKFG/ZZyKlTW/LH2krNwzbdXoxC9Jc8u+lfN3FLtJ58t0MOXwC9ikfh4+Uat4sXPuAYgJ
4n4/bdhlC/O42LQrYg66sZZZpYXzommZaE911WyCqEs+YZspD1axHSMuNnRvEGyHtnbR+3Zwdqom
R59aYw2P6rHqWirOzsVirHiT9GozkFHyt6X7O/BrJf1KzJZ3Kkl6mbgHc2JmBR5aFqtbNFGhXnMA
ZUqho8Pb4I3zplRqO4N/+ZuXsc8tVPfCQecSyC+rZFh22LFq7dbvOixQyFin1YZXdwZyrnzM6wEl
Yc4Sf0iEc1QuRb/R6JlnYGfW9WrwaXlK/JI2QJnBdG3qyaZjm/dHWj3EmgtjVc0Ps5tmFedEOjCN
XLueDkec4Hwzy+fIiydKDDY/II/u/F9q8v1Re/sYnUNE9lHFo00IHlo+gaipkcb3mWXMESjqOnr2
axJIsg4C/J1ix/VPM0Yr4uWA8kL93KZVghW9t8re4m1jZ2d66xoUi738RV0SPnYVSt2dKDQtj2Yp
whl9jx2lYMdIj9iFqBApK6q6/d6GR/6yG0Xv79Z22m/JXNAoC/2t5yhmVUk3ablJ3xfM74CVmU5N
YbNQIRRCsp8aKDtju/cxAt2C51tE2D9ZrLv/ZoqdCHnEzUWx8mV1UnJ1xe66nT1eTI5AuZbffp7v
nr4YWEUOQvec/1KZ8wj1pKsYNqhmP8c1rTBWKJjzPz4jAhw1uf2q/ZtkiH0/AvD9yTbCQOy5JBot
ONH+wjiBjdlxRU4DS0Igf2mqDxXXap/I0W1JvIlIoI87XK6Oo6imxSjdsk8X3EtTFNHyGuiLBocv
BEj6yUu/3tA37OO0VAqO27VA3LFGJ0HI9AW9X9aQfWvLvoxdpEzKH1u/yyCWnPOFrJr876uX307J
eNLDhXxQ5FITZyQpf6D1FJy3illtqrVyjp+ZVpYDrzPzfMDjlWR2h6kKizt0+I07FLWzFpuRg0o7
2gDsZhINKiOnpOnHOWTpCepS22/NO9Y4XoCJLgeJtTJyZhXPOw+lbIlFVVXU2Hen0/7o3tvdeqLk
1Pi09KAbRzVjH6cYVhnITlC9s6Ue2hAFGESr9/gYuk/OxBCjn0SxzePC79nZss3afio33LD53hVE
mPmZHkzgTZXkDG9N56NH+uNIqixRj3wVFQPD0RKVauLZb9wNgPSYSUHzga2YW91zygbLOaQ6SFKv
VMWy4TpqcrC47WkWGkbjb5tDnfmxLG747UIFTlVJzzkIsDvBoE6X/6B3ILT7npz2plwAVs2eiAAC
/6a7pg5Dhdplfo/7xDXTWMK2C3Ixzpy2tv0x8CnKmsKZQaPzrWKWVcrA9kVge7CDdzw5okt/Ybhc
4037uZSFsuXOZxp5vRD2/2vGT/KnfaCed0zE3y7zVhox7OSseXtgdPZWoC3uEj2lbpVcQqgNk+o5
qHmSfrvslOqsUBm2mFk5WgY3ce/l8SXn2zNWWk9JAxKnHhwK2JGZJ2qdb4/4aJypYmuYWHQVqIbF
rCv2jgrI+RdjzHfJJvVrDm49rWVTYAQd4nyFrzPid3lWGCMuBqbRIpZ1UjUO0ZTgBMU3P9yQPagw
rlR3xvnp9elee5i+KeQPZl4wYQG5JjOSpuQoyjX7hPjntQ5+oB/hW7O37QqtsgubYz5XFMT3eJas
hidsBPLuQftQ/rCWKNH4B4n1mZaVoMxvjvEerh0xRJPTviPqkjOO/NhrXv6aUhExxX+SyqUFM5yt
9tW2hENHXtzy7eVZ39u834pTaTVRg2O1dGgojtx8z/VNzs4mkObySwJaQSk7Cr44+ghuS8iAdMOr
a3Xpie0t56ui5a14HKap7hGcnrxS2/FJ3vDZNEfwDMurassPKrKwAeLvAmytGyK0Icl3/ap4lrt/
1SKPhgb0uFc40GBai+y9eOIhnMyEG0wMSzQucibzKSSfybUZb2HbdMURcqx8YWDYts4XG0wVSUVt
vfS2e6KL6PiVrH//epOYLyZQG0+QtNeBq8z9w4ZHxmjASIdWPF3uuNZGfAvx2j5QNMpM7fSOzIW9
VxWj4n97ig/dWcQ4JyaELDEO7NmuDgcofcGon026jkzF7Gf8lWJb+g2y4MXMa81OwD8PeWe4j8X3
p+p9M6EuB5C8Yf1OQkf6au0JzrI7tlr390kgrIuWd98VcJDfe7ZplC1tjvTp+wxYX5ah8Bd9MN9O
/2sO2JGSAw1ZkaAnfpOel/2fprs8jblU2W52eQb4RC3nTswPDPRnAMeCnZ/YmT21RCyMEbR0FN81
l5UzZbwaxGA3EeGqDiHQLHTDJytldm7W/eZ5t8zMoVOKXfwAI63FnNa5qmOWHhWGCd69Qqrms6ex
QaRKQdYg0lvqlOJaele54WFzP8P6RBmSOkVZGQOB6WlGhMofbzCPFxSh6TGI42JE9QLyY3Ng/dAg
HJVB1jj4pbSbDkddejc5zS0PSmaxwv3WiXBIw5Lm6ChZv6Lp2cc47BAj8a5p53UGdjhMssrEme7z
+Cwq7ZJ7tVqRW54JFEjcDheTlNLfCOzTZutDHoKeaRPWXggHEHQCrPkBPOonNx8fji9y2GN1mEZr
T7c9C84RxeuITlD7j4mtOOUrzCiB3ReqDW8/hhKHO3j26uWRS5A0ERfBapQkn57VpRysNUa5uU7b
cPqdVe/iHZ1RpyyuJYYfBYaMcv5IW29PnbiHxx9pJwehzgcEzjp0pfLcHrwir4XMM3Xq3gIseNqb
GW6ZS3ZVxUT8gJVsLgvfu41Gd4F7tb/ebiKGOLv5IjeCOc9XAFxrE/AKF1pTisoeCxku31MTcklb
sVYqmBjo9DwOsU/nMpANFE+ofD+/sd6k3pEJZGgpn4aSDJ2pY/nJMArRRDZQSS30Lo6JDDad3Dac
MxNf4c0JQXNKRtYM1GjEZRf0J5o8qysVfStdiug6fAW0ozdF1HGxsyrwP9U8blKpP6zRYpuAldz9
8gDLSvtLknnvPTQwrc7jiop4xpXwU/UDljCQRK3oZfhFTfYZU1zAT7oISvVpncT2VQw2raze6Dax
T5lr/vUQ5OxXMIRRwtOV6tSLWis6LdJEn+sfZYYwRLi+j7G2wG0ef0habZc66NfgWdNDzIWAqb/l
Pw9IngHkZs0vG9eX2LPCHjaYW6ct8ajUuKovEDXJzGfq6RR0FRYQWANim0lt3Zl+jBNll0pIJl6O
iE9NUPjgT+kMxyOwy2RiPG8lYznIJ1e3OSYI4XMBY7CNoTHQkpqwbCFsitKVOeaetzqWdw6I+s7p
uXNFSUBhdqwpmfLvRHyx2a7Ib3nOTXS6otxZgJH9YK/NfWO20MsBuXObK7PzHDJVTb+hb9jQ3U8T
pD8kfODp9AQptMWdjSk0JZ1xT7f6SgoF66DyRxRq74eEqAukEKaK/f4XpIKXOi90ZEYQyau8tca/
jJwiSkkEQ5GDKeMyIpmQz8m+T3WjfgUnS9AQzoBPpbI8N9jsi6GvDYu15c7PudPymJTQdjgx9f2J
Wfg5+ngWwedDOfv/EUYUosPYWu3hLPWWQFpVadTGQXV13oueH0qQh7YnafK6FiWaDEZnChwgukaY
dV7OSzHPpAVshomPFME7fAdhAz3CbEdmVuACdI0HVfaDCaAekO713PDH2eNm3qK7V0x/TdDsogfA
tF0napBI26a7+B3XoHTe1JURBvsSCmnfabrIlRN31U+vkEurKNSxi6WPE8KQM6FRer1xWEZF8kjH
Lrth5BcxOLWrtbUgKuWay9jAryGeWLaCPnkoQuF6TWVyOUZxKmzE3kWAYJwAtWdx/woGi/Y5mV9w
Tj4W6Oe7kwaHf9WeXZnwmf12AFdEFFE7yPDhR8C2YIZW6qKvAIFrTstB1JDDkjmnGWOdVgxe50Fi
WgLylz0wjxyquvn2/cSO2PLaO5GKEZ/YivuBxrtY0sR7er/ZG7uXxMD+0BtKcRZSZClaoJXUQCB2
QxzBW3Ss74RunoFkt6SUnKgtvw1P4wAukrGlD99genOljLaLdeytzYfEC1MUBUP3IRhgO4ITySwZ
gt7NpV8crUk1HX3AYQx0K7SXcjG01KFNHmYbrDNmyCIYFr8BcsUuc3EXFTj+WpI9HamAmteTTz1J
ng60tRXBeElSUO1efjKuUI7mYCQYJazfI8lxcieC2HH9zera2hAhf7j8IbKyc1df89JOaezUPOIY
+jbg7PKgrL+gHfDjfkoCnAgAHuqHb++Fy88Q2Vk8UxlPUOC14DEOQ9OVigOlQzHdnd7cOZr0bBZZ
MOyxXRjzC4XeFYY9cZ/SnM0+1OPbohzXpyY6j2WHnRGqIyroTbKqIu7zuIRxnM4W8Zij1DNamnd/
QCbqdODMJZZ05UD4E0ZGierG8Fgys6FIDnK7Q4yBInoLMOF8ZTKxpkf6PF6/3tVX1OuahehX15K1
BZvdDlLv9u+yTiBFHU3noOOm5yAzL16L1/zsYILLi6hgl473vYIu6II3iKh1vjX78oBvDp/0E92s
91FOgqG/FCDO0wFsQEL+TCykVCcUONia/e6fxMjUTG8bqiWw1g7Qu3R+OHHzyqJKGkt0p+6sFf1/
2UgczNtzxMctDx0S06wzL5pyRWsnYCpp03oHt9BM7Y1DHzyRq87quvVWpwCdjHlWh4JVz5vX03ch
axKIaWVv4IBUcYAaa1o/v5rxOIohlpe5Aa2s5ndNCm06n7euMH60aDrnCxQeBCIB5wtEpmQzFlsc
eGsgPA+Sb3x6Ufq2kJlRacii1UABLlZpZg9C7CMqND2WDfqrAJ6OKHiTkGLlWi89AB2gWD6o41iM
p8uUM+90VcCyA07wbTQ46s9FET2Bj2Y7f7vTNegS16fg1ZYqMb8txqABKldL6dzstGaD53LE9Exo
27abqIUU3vAaZT6Q3oFZyYVfvdpesapBEBSAxFY7y1f91JIk4SkRxa2WNd9E/5iRBvXNjY7oj58J
qF6P/08CbWY8Eae3gco7LMoSfuye7y/CniilOjqyhhNE8l9VA16IuUbor7kAiNdkDnqR7xZ9li9M
vs8k32pNnlT9MyUx/rc1PyJmiOU3ZCDbPAt0ShvHm1wNGLFoysJYQW9asN7P1HlbO9h7nW1oweC9
O+bR6doMwVxdHs5zNFIfc4Ek2Z9nWxdYa6xKq9O3Q1IAIPOH8jXXHynZi8NHHv2aq8dzTjBFV84H
9Gui7SJO6b0T4UQ1HdUqu+A/Rl/rVdIdobdTRTTbW3ETVUpM+7x3UXM/N42jEYApp6FZhJZTjOpM
K5B1yQRtjocCmalivtdtPbBvu8hv4n+2jqbl3S94GPzCe3txNSxte3GbYM6lknCkQiZH67xDx0VX
Hh2P6+qH0K8sq6nCaB2myxGbW1f1yF3wGFMVLL9SOr+3th1lY4k2i4jKBKe7z2GYbj2dhdNonKsg
CnhQmf2YbKjilInWMArmL3wHchkb8U8CRSGTiMFmv5LVyeKGbn8PoRPp+RZTTSE0/LbSgAsE1pah
ikb5tVH5IXdgkIoltH0/XIi8N/UtbHhRL+mg7jp7XSrqkordK3ozKtUBYEbfEiIWnBSHoIzh533c
bRdoqW4DdlbEnu57AvkblZebP6QZGXln830h0xm/TWm/Qbf7HYyplDYRDlrz5AJzIxlD4yCpTt0/
ne/lyDdXQ6Xq/9qrA3PtKCmt39TOEVq560PLIGsaJ1zTBITq5iFvUynvb50z6V2aZqFPFCqfuQel
k2g8uTkqBKQTx0F5iZdSXfczMnxUCRg27Qv4WHvzRdpM6EcstbgoK+YqyRxSto4ocbSwpNLIOX3L
Sdx+ciwybwUZjlcP+8P4T/AXztsSF9qVWphkGhpUAhTwtGcyDPg1ksdRLnHgbyPvW4prqdblNcye
kWG9UEt7CyOwX+xF54RMcrQzPNPqq7hBik6mqdFhKd/JMT5J4eUR/Tgv8zM+iW4bQTUGVHwggMH+
Wcy7b7sNC99fE7D81ngE8ydivo94LVz2ZMtzn2+x7RzhP1IZX7upi6uscst9sjLhdAXWtBiDjsBW
c833HxGYJIYTswFOEFu/47XMyek8/SHHzR8hmRFMf0j870e5i70hy50koFU0YJoK/eLX8VKkFEi3
3+zLAgOm9FDnVEXptG/cfPfw2mmstwnlc+A3BxxhlLeojdN888ix2HcumLzgwGJabJatueYrHdMo
V8zNX5IJWe/RgQioZwDkQBW2CyVA9hkccjvl9j6xrftDy5rrSzkBWm0bCxTqbrlzDXP5kUoZbPG+
qyZMGkxwIzRo9xb0JwdhbcjZx65y9KM1qG/EXznGCKFyt49WQmrTlmuAYEIBN4dsLRrSYEx4eWnl
exIgqwgAhI3QL1/NyveEYJ+pbuvnmwPdhG/P17w+cNH+IFO/dnAe9xCSQ4dRysTG/l5fblT8F0Pf
z1MRGU9jn0prf0hMaCs0INYysS2etnFlC+xa6EniQAQqkNLpCzhA2twif+HbXxagQ3mbdzL9fx23
TZ4XjmkA7dQ7JZLL+NjL6FX2OVODGTbWfVdX5usJuuLbpdQGEJ47c1mdc/ojZ/t0ZC6XGv0Rkngd
QXOVvKc/liquK/KnMBV9c0RGX1uSmnJ5xt51v2cewsws98N6o+rR8DL1SiBsFmksAy32qUPCTZhj
EMOYUo2bbUdySXA1vS+98bqLWyj28bzQ2oIi7qLgnUONsoCreddLQciriS9tYMtiIMWQZl/tiw/W
zjZ0KHul87oXcZboPqJvcHA4+e3+d6Q0qr6JCAx0sLd54+TrclkVllqstDswUc/1aaEv5gMZ1dEY
AcLuYI5RPPGcxjZ39SG3zGKu65LCt56Xd0Gqwk0NrL2bpnhZgdVRuUjVUjI+leIXSe68cYweEIG4
wrtYxLMipChFeW+0kpZrfpYVclJxBJ9gE3A6Aj+i4uYS45mHw1TIQvSAYRoMGPOX9eY7PW73W7gp
fDtEQfs93KIhqvgol82L/gFQKA6uakeOmYgm16FtFboZS4nVkZHTQigdJchwQ+UBIgYvyPbRNAbw
fh4a0xvLBGOD1Kx70EHkvOVTJaU7T4a7T2bBJqbkhB7IcbML6SdV8EyoANYNZypRehkOlfLZo46g
54lOTrcAd/gFjlNVDEY7rKI6xYdrkPVnJHypRD+sPL0Ki03jdnJLW8PnR3mlluRlWnESJn4b5jHf
VsacINRqyiC+vEIC5KVRYMwWG3x8wtcNtU4dQluDUeS4qGONa1HlyUCYBmU23A8KjvpZRsEy3Zgt
/OAGAbyL6SIBbiHIu27vFa6jyRwiHz8OOS6112YdmpMrLbwkOTd/2PNVOd/FUNR/GFHiZvIsgcK3
L+l5gFVPPti8Ov5STYa11zKa6s/5AWzP/jW2+5q4x6KGS5Q/gyXvhT3Vq5mb/To+mf4cxOJBpvCV
cRcTlGnxs4Laa0lIMLcdC00Ke2VW9l8lV2Pqu/pXSG82zCmg7kYaIAhwZGBDHq9NIXlF06p/TA3Z
Ky75NUXkv6+m+EGMVsmbm6v1PTeiYtHeDLv7fbPXpyKmamOkW7SKfoVlWQEdqrNm7hn9ofOpFRTb
G56MoZbP2LBLU+OGd5YQkxjaPPwMuN7u/zvGAhQOTsqsao5ZDN9Yo08qtOuM8pkgXCWUY/XWDAmr
6aQWA043l07W6LaC/lIFMxQLTvhyGPcjVot3+/J0vqR9YbJlJpOjvLrvQ5OJ72D23f71X7vSiQi0
jUIYnWgNo/eWHStk9SOyP8Mx2CJgK36XrnjA7GxDetu4lGXEFO63qA5fMFU80ODZ1VQph0aVdsNL
Ixx904+gce9OY8neTochnHNn78QePsrdcovhJUh3wuX7dNgXW5G9BX5Qz0WEI0I+PCwR1Qa2RnvB
qoRHbj1Rdhfyyg2OOuv9uG+OcW635a7jrqEj+i2gk4o2iPEEYNirX3WhGf5tDwJNR/LSlSwNiXXJ
uVw3bzZ97yRR5+bFG/f4f2lxB71Ipnnl6H2pNnQd+eohGiTVA7asx1QVHqctWIYyIknU9kNYwHze
N7dYZfqJce3831BqORfI5iiLNLIwK7+xBY0sEA7JNZUY3jihDs/1GZ+ZmNCVQ/wveKbM7iVIMebI
SDN+Of2Ukd2OP+Y+V4Z6rD9V4qk3n5jEuNH39NZnGW0FSwJQeBF67MxSRVu4HplpT9b+xF0Rn3Fz
ZYffbk+5Vcih3M8C7SOiH9fC8tCH7LfOyfY8Ubr4QS1lciq8r6p8K/nEiMLB1Euw4pCr25TIrn1Y
c3xyUj/qmNg1gnzwgwDiU/AX4uSPCukT3IkJvfL+v99zEsKGeULBcjuqAZYs0+HnJryWJ9JNHjjM
U7ftXgrkGYa8K0wdAMkxF4w2Pol4JtcrceuGoQOMLMVxL47IIxHTha2zinFZ6Nye96XOC2wfXfhT
alpxk/ihBDAFmG1I1pOZ7+/S2tDI/+ShtsXYQ6sfjBPhYcrNGM5Qhuhoh9zq4wc93i1tWxYNDsK1
jWQJLBmeBYhs0niwTpFYLgw2B7M4fL6XB2r/lQEgnzoyyUdaSAv2u+Rf6btv+VSznn7uqoHq6Yme
YWMbAtn3HN86O9CyUDGJqmIgTmOjs2t2kFwSiQxe/douzi8xYWHAMfQ0i+1SEoxHGd4qqFTOzLTQ
mmc7dmZe1HN8lQISgyd4Zm3JUi35kZ81Z79JdMSkGVtKQeHPk1N38PFFZ7OL63MVYf9cRNi6/z39
1tnWTs4GKKX3h/uM7GWn0hrg0xc7NPUoo1EC+sa+GWlaI45U+T0i9ypGjqoQr5L4ZVnxM6Rf7Xix
gNHrxtw2z32CqPQJxaHCLG0efV7cuchEq34o+VNbZpiHLTW+6YzKK/eGvr5vnlMpZBr8ufU8Yt2U
lPDKHkpRNGGQNYewsEI359WX+nR20IHn9XnNvrP9HHI8jLgFmYVqdjKXvDUPBl3ayeruay4f2DQC
fnqk/awAAWJI0jUkLlFZcb9EIJKpz7ub+CjvRIowuIZ4lRO2yL7aLlnLwV5RNFUG5JU3f+1YI+yo
xDSWw7gv8BOqzIxLZedFB166e5ikZ5R41WY9ZQ5iqG4OxnVBlrnfDLp3O2LMCHhFkC01z8Ucr+ZE
LQlpVuRm9jv9o4F6QxMpr4Nf8+mZlamY9e/kz89N7Xv2ERDgj27FS7Eqs5R7r7hvQgEa9WWzst6R
+O2ZAoO7t9Se6VyRWvgrginG6MZEwtCtdfDFl2o25N5MOIHpxt6O+yLGkq+558DJSKi4KuJzUdBF
2781uay3tLcyrFk2eN/hgPpkCBwve9x9GKwiIt8aTzbqjWbBev95VWvFq+ZOhkHLRixnA20FXU4P
lfHfHxhPXI57Ajpz+AWj5DGz85svtcLfd7D1C0XolbK8F0QFunbWfR+pEjwd4Bs8Xp4ERzQkIFtl
dwT9FxWxceYlyxvNO4sTLCgQ7f8JklyGzXnH0+NqTsDzICKY/ElfrQY9bYfnvUZDLglyeHKjv1NA
aJQKpe/U2EMBY/icsFm42YLIK5lFjIRyepOVbRLyrr25l/n/AE/32kIQbwUgTG1oLYg2TizRKb7T
N3q99VnY5nD6EGCbionHnS6xmxkfKjROClPE6zIP2j6vI6s4NHisbDo+hZVfE2bxHUig/mtgnGWY
upAEXSwz4oDZNzilO6sWo7/xodcvNDAiZDEU6QHrS4l6cjeFrNDQa2KFvtS6wpgP2bqBuu7Tzd52
+lWnFBwHSu0znex8eJ6fLZJ7Ml9KmJbjYQ6rMJc3Q4bm2N0PPDit+lAucgL/HRVrelo4gFjM7j6g
Cz02JYwoKfhodv2lMlPdQdy3sb/pTG8TNmjvedHGYwDjFzc8X8CW24gOERY0WWfcmDSbDS/Bmz6Z
PnAN7k2uYqnXUQrhWhUI5Q/UhxBfA6uIRfNqRyG73Bg0UcPnzjzc77/tG86kHgCn9P017FVo6QPN
dTz1IS692fisO8t2c5UAYtdDi+l0U9C4/YKC00JWxxyq2PcrRDSAJy5HW2SSuFgZ6oTo2oXLnWHw
xQ20kCSMBdgkqW3tkDCgFyfUyJJkBf6FnjGPKff/dRyk4jGHcvCaNiS9BmtzpJdiLi3IFiIDTJr/
wuaAw7ZTJRvUOTtz+OdLyEBdEXkzZDpZRavat8Z0LGOwzX3k95VQRsVsHAs266cVNQgTKgrcLnVp
H71JOmJPxJh8t6VQqThQ3p+VtMtStP0ktIx4tWXibivH0of/Co8TcFNtX0ypljeM5l5y801RIJKw
am3XOOzZr9fVwUDj6H1PGa/1C2cSaCuIkYyPXAox5hTGfeuv5Prgf7hK1Udm2PbUb6/lvuD+ejzX
HzvsBcvcTa+Pqm9qtAHNbJ52fG1/8Is+/06JwucKLwuVVUu6HkzV5ajKhSgpQJA/xNPwiT97zoen
vxKNvUsDMK3uGEN6agqjalrUE9yZfjpQxFNiCIaOcF8M5uywQ3R7k9jbjmS2HJ0wjtd4kpeyfQGX
DWus9/isZ/8Z0mvlGeb4RkVxCaoCATAnfF3EtKgMBn47o7kTNW9tj93hdTnZH2MgSuZV6PydD7Kd
c8tVZn7Iwl989GivpgCj/is8YUFk9UXpIo7LNfFvbvAhYgwze6iWW+orxOsVHUsZC1CSvWUEPkGD
pKwsy5eliXYvOOqVZbZVp49QIhWUBVLOgGMhoWAAnd71IL1VzyMMDrQz6RPSrIju4xINKtpkLC4P
tqUAKtQFq5WyB9mVjDCsixPAfYrlo6oDF+PpFrnxQFKrXmfjhEohzbK9KMcH5F73LUaQ/hmhsoiM
U+4ByYZTmLys4IJD8NFbyYgNgfcxQQ7HpZwBBa9NyguWpNYukTTCIzfIj8N1F7tirpHwNxa489Ta
7vCrfa9uC1eHhAByYPjQOnPXzZzKISBHPLMph8L1OUhOEYF8ZmEALmFIr4Pd5xEr/iWVb1hZ8YSv
nn94QcxdJCcNQTFmLU5487h3U/zQs+vf/9OlGdnXG+5kPpxLEFVSBJBTHLFrIP6vDU8Zc6jrtGQw
oqMouKBtR0GqZMOz+XblVoTr2iTF1Bqr7DvGnVw0DTGwZAVF51AW4B2yTewVDiFLrcewNZNj5S3R
KYwi/3Mm9ToBRCCzEyu2XDpTlbDCV0/xbAKBDpQWVpIAjvjnhFqlWiH1b7RpUbQ6eToKkMdsZ8SJ
Dsv1n4Ve+gFs9X5tTICktnBFudHZwY+e+H9zAtb0tRHD40DPnYb8Mszq3ym94WORE+j/6I9cbREL
6lhbC/46Zh7gVQ+12e3mbtUEVxRA9tEp6nHOOLOGEPn7gicn/LNVgUIlYtdOXCpMlfXAKjVmypVN
yhOkywXKt35m9t611drWgOJxezi/850LhUWEeMJrHz/jAmgqcUf/ChKyDwWbCSIo6k/iXH3nuRbk
bnO3tNszog59qQdX62J5Ng2e6togLJzjJ2Lk4BjLTb+3bWrXTwEymu61tan6ITKsP+EtfAxETU3q
sIzSdJwbEKUUvb/rZpmDwV9Gg0ptXSqQ1DKOqkZGmPFAbhJNykdbq3afpby3lRhLzqEypcV8ha9R
LqUdXVbwVFtB4nrijiDGrdcvGkVBNk1QPfi7EmK9Ftz0dnLZkPA2KrvP2EXCI0Lj1ysJnu6E73mW
KcBcxLlmvyPwbkH6OKKhbsFyb6NAFgKixres5nw4VYZgB0P8OF3N1DkTLQp2+mwuBAdbssuULlI8
wFWdN3qCCk4Kf6Hq9GT/j0hYVPou8rhOARVzWZZhQy85rUKwKE0qSpzXolzXmAirB1ZynQO5d8fy
WPSkEaAN2E5CwvC5QJYuq+dIuEDQ0bc00uG/9192I+Q1uhrYCJDd3bV6zNUYtw1PEL9S5eaAeE2p
pr/Px9FUsuDdsDw30hglfig4DMLS0bJluvrzCNjOu9Zuixcflttol8CFdc528ojQolGlv3Wi0FO8
yFZstsLB1h1ZDPZYkBF1d3yCNEpUIk4N+rWWckk8WmVpoV0+h7RAMajlfA4RpkoDcSoku/W0YreK
rn9048FPSMO4E+FFK8qgGHuaO1ZrFrz+zwSGhwTx6w7rF6i9A9GyRiVnMS2psevV9LISg/4vGgnR
0zTeQ0Dr5WEOSw2jJBMsk+vGkumXmFuHkWIhsS9uqzprwfTzXqXXmNqbeCtHf+TQtPZsR+5DpgRn
tXzqqCwEHW/p7g4/1viQ2Tk8SgF2a+qhwYEFiq1X8c73LXaNjruArg2ykLQSQ9tAzgdZ8BVnG7TF
FrWu665rOV+Yfqgb4EuscX2BdPdK78mhb8orDuQpVNzVvJtTRlNCKik66maBrFC0tujOA3oTg+5D
4wLKP7j+WQUhrPUSrgniWInhn1VQ3YCpr7pYGMjgd6V1eKjK3adP+Z6QUBoPNp8PZzUvgvz2UGN1
z/hD5K77mdJZ0g9TS+v3RLlKLMqeNch/QbL/ZDeSRG/V8MU+bdQDmK/9dt4Jf7c8rlJGKi/gb6zO
kq5o0kVZq9a5pTaJUfPT8XtuSxwPclBP/977fparQF/on0Ydi2EUd4O0+qcDi43ophTqKcBjP3zx
HJzqT9h3C6rdBCGtwKFmkJvQ4k5W+pcxQ1lcuSrAOkjUnmcQ3jYAsUDmbF5UDEeCrkT5o7Zz4/nB
BlnSDp6FdmcKt0063NjPBCZTZgqiswkAQiR2ePw41rPS37KVd6Sjuad0e7S+pgpi8sPWUkt06kLU
YTIITV4wpWp9bmnrgwi6J/l/l7n6pjCog1d7bRI33EqPDmb9HRhl1XEk/7jW2CxqGe4a4dN7SvPL
Xj6x5iy7p643fERToQD03woI9JTNTNXpz7ykQTUZwEWxFgUUw6nUMpxR8IWPxEmYt5oQ5gmS3ZQJ
AMviLniB24K1iUTPT8iVTCG4t0l7OPH3L3fZZ0bWrMsZgPFfKAECaHeuJIQQbxA8hCcrFrbkfqAb
bitBk45PD4LEW4CYPLJnhE/KJ9Q8tL2Rc+FlvWvYpG0ieHD7BYRSBdS6fvcHE0U5aS5j+Penjk8N
1JZVUBgSed7HMNMGbMilDG1fae83DVBtt++bDMq/Ln2SiBnkhmtfYG/3UwpgVqPxdtFMGxBohFOU
C5Hd7UGGgJXWzQSCMmdIU5hVFMp6Xc1SFWM9YF3jHjtsOHHTRp/9oXItxdcS24D7n761223NzeMX
7ICHLfbdlYOnFj/4p7t0K1E16LsND3kXHZoXA6cd8qnEsCygkJQ8K/v5lhkF2/rKsCKTI1WJBjpQ
06kMHFxchY0Et5sAgtz7Sgt6nrkL15SyuUd8BmqWUT/3d8DSi2WZD3knqKroYRfr36SAvJ7CtpUU
SU7qWfkIcCQEz4i42wYroNIUSTrMS5bzE0LuKk+/sLi4z8MTjVh81dH27SMkwEAgzHGXtLPi5af5
YFMdHNvxQ5szv/cvfOytv3lyazK/lCZVHjBl0xiiPtaHt79yQbHH79qVyBpg8VMZm7KvZGU5VMuV
mLKzodj8vwN1H4JiW68dbP3sbVeHzUIESC5u5T+YZM3qFj5HbmnWBY6CKOJmDsMf12yq53nMH+n8
4prnvMp7jZjRDnJQBnTuER2If3RUAmU2h7u1tjKE1tiZ0P8lt5/avWTtZpRIQXWpyfudUv58OBeU
CGNINzNyLDsLWI1ZzQdHzlXnRS7GmFQXKL0f52qpLGuV6cbBAVujAte6eRWVSd6nf320/P99A3L8
xML3HvASmgx94KQiTKSH3GZu3c6eXWslHrNi8jpbFSEc5SdUBPqH4Jfncjzi43Jh+NJo3Re77lvV
bwieQwt9Mrw9q2hD5Pkc6fyq/RgO/Uvuwx9ZVJ9wJOaBBplo00bP4eQ2LHLBD7KiLIycMv/TRUyt
4qNiSallX/JnwHZFUeonwvgS/DmEkqjKoX0VsAh1y/RvvuQ3Rp6E7E35XTUTvarkxOKVYYddooyg
H+PfZj4QPyz4Yzg0y/Pv7FERWzf1uYn1KvsNeJafyU6PGghJ6EJ8QP6bELu+RipCejsr7/6VYo9E
v4MQLY8KlKIYzoBX0w58iXV75bCTsnHNu6Xm1yLMPAGDQtqmetdrBwNWRx8bXlNCQtnyiOlm6VzM
iCs3DdXD6uvAKtZyMx1az8/gmaTCpbpUki8wygqfb3Vp9EBDW0doTguJxcKNcH5D/Q6xfvf/VQ1k
q18DEBh1xNF7dbjZNGpw8+4J9qYVjzkqPOkztHKrdVd0f1IJ2NeHnpaF9PdqzM/sfQKm53Ck+Lvt
S6UYDINxJX+/Se5Psi+iV0p5hVD8eUAqy8gotXANriRiM2GVgRlY5hQFv6MmMLqEFX6jFl304mIk
9iOIjvmcarpFcYegc2NzVL3kvH9cZqFuwW5EAA05nD0zItZUivzbTCijxP4RUJx5H25kKbl9n8cx
1Xwm4kwMM3HKZgI8IopqM6UaBjvYghJHQFCFGNhrKLCotONSsGcna6N0c4NCfE+hPfagiHl5TJIE
n5QI6RJ7s4b21M5tF3pkFofAwqOcLSzSNBYG1QnzN28hhZaiUO9z6TUkdDN0F+Pc/dzMFsP/ttr9
P2y0VmpoNShbGl/dH9bnXiVuIWELPef7e5vBYZ1F5IJ4+H7VTu1pUoLe77S5Y44SYssd2hU7Lmgq
w4kXdz/AKrOR4Z/fVxtnlDwJ1YQHDIDfuriIpbGAxGUwxSakLxjJvuH9EEY4yBjHCOCHORkm//Cz
3FM7q7MJE+aq2Ex14J2WWUC3oYs/VTahvecx/cnWu0tVfLvzML9xRLoNO2LcVUpm8IsNjT3omUgg
75rsm1rUVIYr7XjrqHI2ME+d30tZbYE4cgMBHlGbd1nmHcsVLTpovUt/2xqOZQNIob7kfUXUDmjZ
uVZ7hxQiR685nmBj9Rb7SszSGnsMP4naYIkCqB6ojEj1Kp0Hk9Iee2XOXFqZLpcETelh8rBWgJ9J
cpSqs3x1YhvVSU347tgoqMrM/ZeT22wte/nIWVE3xKnRIP1ay18H/7XMjARCkD8Rui7UWQ8sb3sp
0ee4ZuIO+5/dZfhD+y1FMKRd3kSi0ULj9cMVMeC7A5i3cUI+e1WCKjO0d3kTsE1224KHIZ4wwnXj
ZgKeHP+epcBUpUcrZ3QA4/Zgps+sw4hW2XB1F4Agj6GziqOCn4DXmwlgqqvkYMU+ZmWPaN57rOWO
3HqSM20zadSF8VxdcLBajvhs7P7kIeQUedx2SvoCdlz2fYtYTk3kNam9wVwibg8TQ9gscnCZfyWM
5HGnD9c43+FtNmMKLEYF8203ZLLOITN5Z2IYoeyU6/tN5HrYr1sgT/2w9GPaOlPHa//RG26NeNkA
D8eX9+ZN1pBBSdA03Ois1jAhM0hLLxB09iHnzDg5b5ecjMkeSU3U7+nJL6x21YLKnmFTMCpgQcmo
YUwfgL3FEmnXJ8jW8HzWb3bNpgPtEkMjuS6eyFhuCudEkvsKdCZ0jfbhp4pDb6pOyIwqzq9K0r9f
FAAggL9xfaZZO5dZv6MiaHH5kOiDwqM1YuifSB3YxMkQqfNZYqPFBd3FdN1RTvVaViceyvc4hf+6
yDg4pDZUCxlNttSeQZtVry3BdlZSz0RquTztkeX0SXC1+rL0lplga8LuFPmyMOtLhiP+O7QLH2WD
mWriMUKLNsAG2FRzXrC4ZdRNSeyNVuHh/virKCCVp1/+HdwiKyNnYFsmGt8QfAUA20DRq/ti4WRD
rWTyBXUioOqsUeRR0VW6lnlBVlsGleQ1s4Bj864SOIggfkgSDI5xPrNfIZ02VERCnGCW22HY1Dnb
uGUPtM+j2uPRgiXzskni2mt8BbhVzz3JJ374WEKIxF2x09TB6/rVX0DzllFn4OoIJCgz4SkauhJp
FSdP2ia4pGRxqWD9RMuNp3xG9vfcFHG2/j7QMtzhg+rNOy0AY9bGBPgRX5l/b+Gbn/Wnq4QAfkfB
5aH6JXIAotJoch/1NiXj+TSfrERklyVGBdAminw3RG30P8olWktUjEGGTkcbZ0DbDejVipA8EXc0
xzFxE2MF4Fb4BlUuQm5eKKATK9QcblEQ2fu8d3ShAjUwC3ZmJUnBiHnKhgPN6y4zCApHhk2ywCR/
Ez+FhAeZW6GOJt+oSHrHdxLanEcNKTkINkWyRx+IWHWE7djLQNyHE0M2oYiYxC8cMM03xdteARje
Jkxgcbk48G+ZDXCLmJ+iEchaqzj0/hL9L1+/utdb1QAHfRfeV/PHgf/1G+icNgcggx5GR96tq13g
qwX6jER2c/XzSDUpGVrrqSn/gOlgtjtepl1CY/4BsMnfD0Zq8ZrtUVbiMoiUwx39JRTsZ/xDIZzK
6t+MORZ1+i8hg7jHdZiRhiJgfMN5c598raigYxck1AHnkLO9H/VWWWESAfgZ/Nl1dxw4cBS/sxJM
SK0sD+xyiG74hTn1sCZ4598FRZ8J+s8Cr6Tq3lq6VhYeXpjpvFjpeUkMpvZh8E2dY6tTiYcZywro
eu0TwdnruaJSatfnj4pyA99f14myOFfO/rqPXKymj1HCHegChW5URlkHKvADXKkGTY23orOeeI6G
fRqmHSntmXHpmavM6xLTGzw18gV9DGlhh7Y2hAK4s7IE+Azqqk9y7PqS0GH5cookKqjK5rr/Q97G
X3ar33f56TnzxZP2O+e5q45srlEIegrsk+vDG1ftoz36x3jbRxR2uTbA5Uh6uUcZKu6vHa4NosX2
O9MibIRgyz6pVMN2r0ulfm7ig9oifSM9qrjS/cwRQBW4UKuVMj2PvzkwvqZllAdnSqB6tiMmn3Ux
NXuvbZHiCa3lruieJeg4G8AbVb1A48se4tkHxvgbEkMTuKm/14G6txMLmQK/DoRSjzadg7FTTAsI
EK53X9YRr2Jxw7jvOh9mjqBnYdkrhioEESJu7pMP6ZT0JIFOoazX1W/NE08+m6riovgFE6gFyk0q
DpJaU3SsHSDcwns8OC5y9+11nboEfQYth17nGFhCtvcrtdfwVPCTRwvNR+lPGWQe/PaiLtDeKY6t
F4Sj+NQBoJRXzOKeUtdkaUjwXq0+RvnPVKTeh55tjPMuYwQveo01oQzGukOob2p0lEk+PR8McD27
3LmeqKFLtLwA9Qr9DhqodntUB2qXmhGgjTFrf4J031vKzfnUOFx1t5z7BgIl+ETNJcB3/k2wAvPV
GaiEeu3YyAHQC2N759ZZaM+7jwdSHz9hOMvhovnnSp3uZ+51HTqZUilaCPEfEsqS4TivsBgzyZO1
0hWSeeerONQoHQMfx0l+rPT5nNrdTXMWFVRT8Gb4FSJnPrLlUVVZzVA3rzoO8Y8AwlY+2YffhgvU
bCF8WAElyDl2J5Q1ZKfIb1t9egA1s/CSyUVMxWgt8oASEYr/FSfI+Z8+XwO5G9OUL31Rtz5g0Eu2
/9XstnrB9RnWgAaqscwXzCehmGwupZ2YC0n0d2ohZavtfwG19ygeMs8OOnOor83tawOBsaQ6O4ji
9OTqbUurABJs+/BIdxS5Nkp16dIkcVM2t/wGOrjPfaVPJAgPtuwWWEXM7DlWDVdCdqCg0JGSJjlk
jVFpbhOYAA3utiI7MYFaW8V8fabQQsgNhJUfpz/fH9BBypH6SDPmW32PhtQ8+/J98pN4fXk9mjzV
3Kc+kVcxxTzdAtnMpNAskFsL6ulTNoLJtUpfUZ2G/rmt7ExgMW3dnYW1JZcD1bSGJ9TSQ894b/u4
Rk/NPhjw5DxND/KCOJy4+iGWhi/YsZnwvcncLu5VSNSSWwcsHtyq9U03zSX+3H02Jtq6Kp/DcMev
d0WSY6s9BgX4d1LkWh2Z0DHtbqFTlnqFLX75BNuwKuC4vjswuNlKntBbCnyddy1ujecZFU/ovymb
Wt+T/pdqaai0963knepV3a/qmUv/MQi2RZNXlbsDYjy1HlNUuVpX5nblYFfW5KrTrhGv++z5BO2d
FRJuo3LA2mH/1afsTNKztO59n+4tdE1zsb2gi8ZkTurASGV2kknfl7txALJPQFDzI4+NtvRNz+9g
R0K2qAidSiYaBR8ywfJNtm45UX8NiqjWG2mDGav7wYMkLbDCjqOR9yBS4Je0pwwkZ/L63zgRBeCo
FxT0kx7CyXnXrSP2fTUHqIrb3Z45QhZDxE/BClTig0xbxJHGEeBavpRV4nZEsNw6sPC2jHvsb/bd
rJUvdgMDS4wCgFGt5IyVcma4wNAMMI6wH9tGsky9efJFQG21e5ybhwVNmjInELg5HwS6EwrCZMNy
k7MKCK/2hz7zy0xUNfY0jGck/sPqdbqPmTe1fTP4fnqXTLPHIi8TIsTXF9SfTyX1vhSKOQTRuFil
Mt1b1Xy71ztBGWOtWnQWuFAh3hQp3Kp224qO7m0d+dKMhU/fxc2JaDXrflDPe9e9YKWuoI40Oigt
0dpEsUBqEX8iH80UYw3dDjmKsPO8Y1D+EmPOJRlDEUCgAUbtXRf9OX0q3ZNqmshv5u9EsMh9NbKr
hCS0IcZtE3UkES8CH5nHnPZj5XlFDEpAAIRHl8Zz/gteO6PqraqvD0Tnw6QNaCD3bjZ9cNRGeyI+
YYkGLh7NFET6xKa2cgv6t5uxnKz1fKx/H6IjmTzAyj6zzF+kA6bp58TRdvR2jUBIAuIqxZSq5p82
WPRuIXFPnOpDU4XmXRxa8TclAxIKBrw3h7+UceoUmw+oDIRn8Cu8/1+A4D0mr4NMyx7jPFgAQBXW
FUTc/UroqPIUtDxrbNKDWOgXIynB9gwC67Y4EACA1EfcWpTOSg9VcBMcEPGHXLDDc8+gmHv69amt
OrdZqJ9+oJOl/3oRZ4rArcs8Xo6I7OlsmMtzVttUJFpSha1Y+DABBVMtKmpKOR8dzGgOj4K9yreS
woShjrdN3qP7a3n8vsN5Aqj90jeKyq7jw0XXROa5hOR1fAs32g9lHDtaBUuc+x3Xmwx3gefHhhdN
kSZweUGvM0JhYYFtYogZdkZi/2aSiGX5Dsu1KY64Tctq1yrgaPZqbgCpTS+kU5rOXmM8kJINDISr
oGBWGmjdwDWyNqIMHmpsXipFh8vNIpvfiHQlNch3iXCMejQ79TE+Fmc/R9tPKpFZGhQ6JiZbNQZ1
ZAD6z47OqyYBHM9KbictoXhitjuTnELwV5ui1QPPoDgin7MSwYtAyUjNXLP9Jm/OoZY2YybcYOwq
OEEIciBp0ngL/uY+NlxiWSzmH6a3oHTeQwOzmKPf5PhmOMKJwiRzBCOsB+0vLYPAB7MhSaqYwYFL
Akk43KVPznElCNMdFsu08zbbocC+4U28sRYPUtvVAH/1nckLUAp+rEUfrlq7aANIYic3JXIPX6MH
sgNtR+pBsDFO+gRM6jtMRv9Yz8UFIUuy6UHgMktvcZ9pVxjpwF2+b/NPkM/c4gmNSeQ5mEnooIVL
5rvA1R3+/ySaUz/kgf/MSDmxNiWDb5q/5kUkn2O0Ug+Ov8TRgEHCgFT9ZKpYm6iSKOqyYN7amkod
o/zOFL8/FM7GXzpyVtaHe0C+w2r2VmUjC0q0VHiMC8afg6NvgoiOLDC3501H0SI0kptSyHUdzSlZ
YcwWJaJbCa1aVksiBD51QS0YA5NI2jT1jWiZaJNUJblssbXs8UARDP6SN8xTMz8p+UUwe2b4mxqW
X/m+fkLtkeqzkLXWlIZIpx+6CafiPtsXy2pkcOKGlvnZ75vRejdiffg/EAPsCEgaXmZDMDHKcOoI
4Ls+THOiqKl64nveLF2YbhJ8ksDCWoTQte6I9a5msXDLkpdcuDtJL7t7wKwRerveHx3/Io9uI3dB
Tw2tmMg+UPMunyer4oEOPX6Udsc8TLUIT8CnTUmNsuuL/BOJujpB5HUfKv7mkqMqRA+HkWulW2Ak
Op0jNBQ5d72PbbTq1hibQTQkulp/MfNr6iPRiSj9ejNoI4g6uyHjsiFJOWIveklYhfR4LpQV7c6y
wyIS7IK93GtZPx/yRujgFd4iEZWsllKmL2rzpLYFxvPMD/vXRejgWBfGOiQhzppRybvYYDdoNyjk
gz3B9jTf0odjELQ2lze6YVoqOjycTPEMWZo5Dt0I8fpgN5izBlVA+doKTAOnHEqh8M+UhJEycPH7
EVmE1+HLgIb+MQiksr1px3MJyUzqRI+YyRWjymF7fjtFdJoAbmeAz3/w4VUyzPDcBPpa6EzMZGb/
EuOkBMwNJubUhXbDMEWSGBt+EE836bN7URJgdj7NZ3jzqLukflUMmWdORtAARFcMaF8k8MwpZ4eq
UGaq94wQsdOGoTj1LtJl2hAmGDhI5yu+kB+2TCX0w0qKpHyiu63F/pxlzsVgNOpfTBh+BhtrjVOW
ZCKwOdSbKFA66jeKcJQG+241H54h7raY5IUEebDl1gulqlzg7uysEU3zwnQoL8MFRSzs0AXDjg0U
y/C+ezT4Ms8cNPGmfQ/r275QCuTjrAxplrsTZQrizKlxwPPGYGIqC/mWJuqIZnUpItI/iGVNDFoC
6FAedvIk27vlpXsfhJNnTWHe8myWKLyhHIKLcVHMUa5ONLBaKtNDpLOuYnbfvE/5PTVNIwk8vfmT
zHZbHnoak7TFtNr4GPSeNm1SSGG57WShtF5Xk3SRhHw8n0gHHXZBOHRayBaPsqpFfOx9jbBYG+3m
VoQj3tn77cyTLvQQxe0MUejIap12MI4L3Umut5+Yl6Oivgi+rra+rsLG4c8tb6mrPbgZRondQ2X6
J9AmCLg7X+u2MWR3mlJC7T/aofX5ZTw/Lp897E1f6YbcUrpKfedzth0pkIU1rDvaeaI5xpqzzZ4o
g2DFqChKaattivaQ8VDhwVuCoAT5VovlJT9R6B20+drzusQrRO2sAYMWCwfk2zkIl2p4KrT9QqU9
U5AKlAxg5c7qngnjAKxKdUXPa5+W+jnW5iySfStT4uDtkxZilDKjkwA4fyzc/jZoLODQbXYGwfi2
/JUdUV5eiF/yGc4RAZrXoJZpi0onZvD7J1XJE4gTFCEfjq046ny+M1hQsgFeWZpD6wZTUkvXvQC9
JVKVZGV/Z+vYlWHI3pfFI/WXa3pMQ9eb2eVXosUDJbcKHDNK/fjZUvo2vVs/VW4wE2dnLaWAO0dc
JldXIgVhYtHa2dhjn0an4Di/tmfA3aszlOSnglNGCyfUPtPrAz412n5w5jqchSItJjTVE0N5ODPf
bMDDPA4bORurZV6U/snbURXxRKpWVxHFHjazIJN2HHQVncn5lDjBWx5brO4qA1wTQTANTioy7u+I
ZLxefY2Z/HGCdOa6dlKVkmDZ7Vg5aA+W6xwoPqacYeENb8QgROco0zVErG6zUgKBtcN8cokBLz7J
SzR8Yk2vxEIdn0a465SQDHs/DwlX86n6LqO2SghBm+JBS8PFw8KgGtJ4RzUH/T0tzGtTForTMYEk
qtDdN5w7tCP8YDnOhVG7icMlFFDw9NejblgKwURR3hDcirhTewRqVwCnofjCslZjjFddJgN8DRNv
HFPVsg67k/VjyPtvw+vm/TJlpFCQm86E0c3ceWYipo7RuJG5WnINaH8kdHzEkCuWJNtU0WqNXiiQ
06wbybGIN9zjg3kdaRM58ooxofe2gnhk5O1pWZxeMwM5n9gUSdKbubPis5MszDj2zHxpIo45Zr8W
jDq7/L0aAk+Ja1Is0rgbgJxhfvL+WdSnJWopfuKcpvtkvV/54TczwrbvvxGhQ+M55zVnnMUJmaj3
jEyhnwIzH8zZgiUxu0fREVV7OvjKY3IMaF9LsYfm5ngI/ecAXTGyvLQm3MWYgV/HYqGXv2PW9gMg
w10hTrUS7u/5PozFyKV7/1Ok2tcPJ69Z4dzgNTi6OPsL1cKATOBNXyY34QTSXFdFA8qitNTm+sPm
CV/RbGr8cmk9eaE+pPzO9SNsid66GBIBnd4pL2KW25R6ocxhUV8WUYl9B1ND7t4N6ZxYAcGC630W
/ygC0m/KQSWP3vkCADLmwOEw4OGEIlU/i8agCo0u7uayFX6I9RJRDtcNP6ztJWmQ+uVwlJwgb2iC
F/GO/tN9me2PWDDKSEitYvlkTBoKQWRo+K1mLq2qfg4DkVWwMcPMN5HHycFGoViRffGCG8CQGtTp
zxk0z/QRCq4urT8BFbG54HtRpzObdlJy7l728KE5SdtJRrDjiURK8QgZdkzMVnEzcb+LHe9Bm4+o
7eSPqgDcWj00tZHQ/1Xi4igYSM1E/ppq9cAze8DTsB1XGb8WbG+XABgD/ZIJlOl9aqCoMoDLug4K
YEjRCpIWZBjry0OZAWz8g/XHSjE33WRA4QrFKK3M13FEvkp2ocxA7ZJfjfUekxeUh9rhQhkJ5wR7
OLiXpOBerhqDTxBwKpAuEN709dHZiV+vtlLGal65LSKp06w3Ul9GyJ+NdiRP8XfFPtVJf8thhfTr
vxuD/4K7FZ6Ak52ZfO4yXfX1dRrgyDfm37k2QS+7DzXb0TCnZY/kiHxHatJiWBu7BEu2UuHE0zUU
cXAbs7K1h48VNnYZdpj8xi+IIIbecQ93lXivr0mccJkori/cmbN5e8xKGGLM4Je1gBpEG1US5jyP
NRyg8HPZMEC0xQ/2sKv7AN4LaweGmZBPRcT8pt+cWFR0LYAUnolv6sQtmRzug7QG0Sl2bXyb3L3o
XyW5BoQbzX1hkVYv4YVOQqv+HymDKckOjtvHAacv2vVe4qHOEJzcWWyW8wekzK6ZdLfke/hgQPlM
dS9EB1+keqK+4I/dfCmpI5Jml8rEGPabu9ULCb1PQssQkT6I1a/pwUGeStCm5ETskpO7rvUIbzdw
cKlfpMkzUmwW2+CeEJrnGmRUeOXRin+bq30zkxXhb5OKr0c+dPMbhfo7SEaUC7E86vqGe6ROkFCe
mqPiPZtInhY63yAhNlQl7RpyYQquZ0lSJDd842Bnp097bot1DdWIBo3B98MsyHQlzT8HyL+jDjQ7
lOMLny7m+IPnaEmR8OOVzm8nG1i5MSxjHdxWe1OIGd8XU+TIJqD6eDPfhZMqnl7V4iSDGpMNJVUz
UwySCQI+VMhNGcNUM8rxCiT9gYIHqtPxGJpG6TbbRspbwfBPPqJoBOi8+meCNAWxrizVrKjEfImo
3JDI411oJhWk9WRvgcFeJ+RCYBpW2NPHBtIetZaYBGJjfGYIWW/CrgiKSErOpeVl6eOfdbD7qeNa
fh+KASFFP3kOr1rwLD63rY45DhntZxnMI7AMY4CXa5Iq0Q6oj58Ti/VSn97HGuhoOxKLvP9NeWzY
yn2U3Y2OIc9o2uDeWGyLKne2hw2Eg+ON4UTX48NjwpPRyXghvvXyE5oq/ZtsjarEtUppflV7q+Mh
K8RbKF4yjqE5V5ayY/vq16qCCyL+R54Exv8gMn7gYNyHKaoUOCAV75VvFEkw517xg/gy7vLebk84
4+DnPawSw98bMboThTsXhCi2JzXYMCcvWAhpL0yh20zGEOShwXaOAzyXGnnmNqBfb61PRtNwlEQc
aiwcUrc4o0S/onT+o4+qXf+KIP3U8yXnPFIB361OYSIB7Jh0j9BsQHpe/bM9CrvjtZyjkk+FjE+q
1cGU9e5GEAW63z3zfBNu3arDEUA8UoEdUkf7I4AyIIWBLJ4gih2q23hT+ipNRKvemQGfoFvwRRHO
kqgbnCjoJw04t5dUbX0TZVtFMh5E9wjiAAclKKbyd2yFsoZbzDR65uTjgXZlOi4fKZ51cNHe+aQ4
Z05xP8hCb5QR2gLJNOthvs4Rqxpua0mtT5i4xZLYeKuWbRik9KqPfQE9ag2f7ZISKA67S/EbY8QO
qtnfLj9/PFKPcqk117t3ilv5UK8J14skhHtKAk3cf+0KR+/VcFexj9sUtRjn+ZS5tu61E99C8ejD
LNTI4OMLbk6m9XuK+451AOfd/iZHIoDE3lD6NTFz1Xd1HL5iMuUiOyrP6iwNIocGB7DKH+m/QlEe
EqTXfpZcTEOW82pH0uFs/naHMtZ+GM/WL2Y4bl54HiudQWOxp0mKnyAn16LJZNAmc5G39JeL8hML
0i1T/WNQaRfPEtex++J93jbRwQUPu9HfzmHQQulmwlRZgF9ydWBkWBcj0xk6n9LOocaclVmZDn7T
Y/T27yQwGphB6kitkNBdEKc8jS3kVgZJHxEfpvGdB+ZrmzDUy45S26XBlmEG9R9rt/HSzcz88QXu
f/TTtN4JM28a5YsIGY313Qhkt/bSZLcvk5Cm9bdP0llDC3c/eb3P8qkeEn/ViQIJhTM3FZBxAG3R
WGoyJkwuvGBc7jB0p2+gANAxAiIr7R4O2SDOoUri5E2uOAJl7/uvkZZW02cC01XDWF63w603OU8l
ki8rKQML9DkV2Jn7mwvMGTwDGwAly5x9upavjhx+ZT9nej7RasQ30NVwLAe0hq7zMKj5tk6p5huH
rLYge7NzLiYfkNwiRsf9lQHAd0NlQvgYOWY4yhlwSDRYlqiKynC5L+No852+aQn6RQF1ZExUQCMM
Nre49rii2IZ4L/IowCkiOWHKQ6WnCEZiGZWWDdD53ytk/BoT9hjf0nyyd8E8sH1ts7SZYfUT3Dhl
vN6BVI8/M3EDEQzl8gRqSnByDUFCA4geEPNC9d6q99lNgkjC634/G6DHb6/ZEHd3vSE979yJZeMv
FfuZ/iO1cIk37ONWOUJnsxhjE1U50B15yKnggf7rfOslx37SV5ecBjXryzWFTCC00RVudNvrz17n
E1g018400JYKy6RGIyI777mMZe60vsNO7+1D3IrquxWAGvLUH61BQIY3Lz0kxkNJvYNaVJGD9BZF
s9WvY+c0aDOeG4cb1PMeVJc41usgt4xJSEK+STHhsMwEgp5E5N4Z9A9JbtfcE0Iwl8yagndLye+m
d6tj/ocgogb6E+W7kHgb83VXCsFjI4qSFsrZ2EiPnj7d4n1BGL2ZcxsjsUWGwK+xgXC0iRfA+4bI
2kYqdXVo1RxuvMAtBIBvUll1XwYw+LvDq0n32qZx6lMc4QgnmDg40jgUdAKhEkn0XnArO1RUqXks
z04EHB1lkZTL/1dSjZ0M9H6Zg1d+9xsTms2M6dLVmW5l+1/TkraI09sRPMvRE5PVVyXXa9nmAs2p
JD2g5d433j+j5WGJ6cVsnpbjUrdLk0eZ5UXNVSEqu2MlmEmyh+Ktba/8fS9k1cCQLaCofM8yLlDT
nPg/6UfCbKKWLqbPFiyyZs6mNL1ihBbfUJ1ZogDPKr6GU0mOO0kzbZ/0EsP0eOtZJVZPfH7ppQya
vk9GI0s33l/hgpj2/3nDHhtA019x/ObR0Iwvb5STVtCH6maiZxEZY9DNusdVbNmFnwxK+SizSuYx
UT9kHTxNJs4maGMMJQjNnhQCkj5BJXpPvvWeA3Zz655cG4x8Q29zeQp7eVfhEs5I6NMt1sYcK1Rf
d8cfZdSNeMp+uw2YfwKePxiaaQJVAPAvoF9SWJ498B2y6pSbMW3+puzGptHRIiCOBGia9SdtAO9d
Ge/HKYzfOi/zdzeWZ0vj3DMiHypkxridkkIEYKMJryNVA2tZRpAEhElbazXISQmTqMkLiwmDR/o2
9XqSZ/yfTcmssFXFhen9FiaftZN7X+FOXyxA5pTs8C/AaPT4T1kkdBLg1ELb1XX2PpyCaBf/ZP8U
WXuXMvCtzJFFMGnDhD6/y/pygdR2EHuro5hbRIal+FK0i0n18aYVo7n2L0UD9N3tLG+JMmo70pEi
brZo9yNAveqlXW68Znw8vDfNsgydsLI2s8A6bJKFpKtQpw+rm802xAUjzmQhHvt7UXxHIF/h/oGq
5HfRy7R06OPyAZWJqnCy87TtVgDpsAWeZCuEXD6ZVJRJt6+Mbih7Xi7yuTSPitrENG/7+b0WY/HF
i2akCPvbJrTFW7534ugml2dTqpJ87Hp/TBTrK6OXKvWnn64VUSWawf2qEFo4dAIrV8Nc2QeZT//a
dwJ2KcHJk92TPFSzecHsBHoeNS3+nNLkkBYmQ8uck4HqQ5kBr1ZK+kS4umrH5xQmRL+FL+mQyA10
keQJiG535A3CLlgN356HhufeDfv3IJgqnIDK7JuSxKaRcz1lY13IHC3OZdqcEmSRTtPkwR/yk8RL
k4Jw+ocy17GI+vlqASf+zLEVL+IZ8IG8p01OwRMX1gcutB50nQ/jU/Vo7MSpLg9RqqeIIHtBcZJf
7y5W2pa6yUUD9h4ucY7KS/7CmgmmzA9pYxV2d8zZ7RYBFGC05U4DDEZGVGnkQByxMtg4wFY4PrCk
5nxpBlRKZYYBCeH4Sn38palfFAGND5DwVh+caOevGgu3Td2KX2vJTWwQQwMBSiyfDFoydeuGuKPt
ljHHUTKWk9xRWr8GCRfetJTfg5kToONTQnr2aMoCn51JVRaHPrZ67ko5OdDbu41iNBg5+BV/9G9K
ZWNC4TxkfCcdWc+oQ7f5kJ1x4Cygtd//m0Xlr5rVdboTrNJb0DpclNGJrcEmq5/th4A5tswsBkX+
KDuA7P39Xw6aCQ6IbVLBqbBetE0GYnu3W1cSuuta5XjaI8zZAYKELb2z38y9aa0zCYP17gnhDUmD
Zg4f0OWVzPMWwKz8Xii6s8BJ9WClaFpQwDbO/r5MmgdowGr2CjtodBXJ4TLZ759lkn+ssYFAcft4
PZHyUValMjH+gMxr5DJ1Op02UI1ShDXGV+T/sQZ8rm+Evbe1k58wNpakg47uPkNgXyYKjbupRnqo
VxKH00RXMLdVWs6OTzOSFL22aez1mVyof7X6M5/t2Kpd7MpBwfwR+kpTlYlNEA1hd3fe0qAeFdlV
F6tf0n0VDY9Yq/RxKJCXWVs36uXJaPCsKByg7XiAgvTQfafBaZNSfxhYbHl3XgQ3ERwyGh7pO95R
eLSGJBPwmzY3V2D2M74r51kl/6KeiPxftIhpwyW1mV7leN+FTbOb7vfnQyerA/RQBLZ1deAoVjoT
oNZs2cB0t+t4z+QvD8FCnvrTGnSu4iouDGs+zr8Yj/B9zupTrxFor7NaKZPq+D4MCsi49EEeOq9e
Gx35pkSk/hlczK29g/oj781ePYWkCl85LPxRudbU6S0mUxC/+PP1ob+IYMKmVK6BD6E2uAQGJ67C
NriEZ9jVk34Mf4l9NN60JF2kRjXJ8xswO5XXIYsiEdujbP6dOrJJRUygMnLGbazdfCMIHQEjSGRI
rdOx/EmO+zwTDLwjVwriX0NncWjRf6B4X58LeAH6iTJrydX5FLty4AP5bM5NCqWlZmx/pYW56ZUz
F6MIXYnqSKQGLX8MzydVhXLSjh2rvjMr5RbpiM6oWTkxxO7hco4BPj6RJ9RwfWqIj+pVxl/A79sQ
dnsUmxHEiG/uFlsrvtEKksVvyQKMsWQzbYtgM5lkRPmWsFvTAhoMfN7cY56KqANM1dnYoWvwjFSZ
d7pWbT3Mv/TbqYHmxvxIt2cbHzY7wpu3UHmAmSqUy1YG+XQ5G1cKOKh8w7srC+r0RlmOp3iDV+Nu
v+4erhiRFBx4kxOsnr/FSxiB8The0iTg5pFbvRSpSJgnE7t2Jd6x+UANYWQm3Ay+rG9zNALL44h8
sgHB5FBAA5q4yKEeuSxCnhA3t7j5zdLcZO3WdzEJ/XvAQUZmhVy+1PZOpC9xMG9oen/miG1EYvP8
2gjpU1wS/8jNawWweQb8Mn1jGGjroaazqLOhY8JYu2Tat+gMrtyGp2CZJzr7EbAYS6LH8tWolwrE
ggDDCQ5gvoAHFeMLwH56F5XmEzP5bV5p8lFqTSB9n27Mc1CaRS0U9J9Z1eZz0xBdVm541yhrtIrK
ljIIWBmLjfrZY4kYqcmSrOCSogJaRTEee2YxA2utvD3nlX+sEXnqTFCiDCsXxJ5xpokT8C0NN9F3
4q+m437oY6kpgXlyBq7aFoHJIEa8A4ek+sf45RXcU9MoPJu0CvoBZkZPqVVVuxitYNSOOVdiKO/a
e9/TCL3dVwLeYvQ1d2Ct4dIGk8El5gkhe2F/CpqjQsKSAvpKcMr/xUg4CO4YvU3WhNR3MVBVg3j5
u4OFSoI+Bk7G+VOj8BWdfmCXpxIPlSD1L78H5Gx8Tn08/Zfd736iUz72UoZOXT5x4tT3d2MhD5U1
ac1rTnyUkXio1tecSPaEiIk6W55O0CzVAVPGcVg04OEAsBCryKkrVQniXkS2CLzdbA1JtSJG7uFj
VUnr2a6nWZIM43NZL/qw++qbGKFTvR8GHXt/5o3LP88op/g+3wPui8yXemCbmqKFJm88BQFKuCwM
FGDlYqtrS5jJ9RknOcgfmhcXMsovfgay4jyNfmXi280opvwj+tDFYkpSomNUYlLPfSZfbURKSklA
YQ9dYzyzUz8iUEHKu1pgwymW1CPngcyHUoczAiFTjcClsCQbgg1WLPfJ+rY4syW0W1rORJv0HcI8
FlagxUMkA87zyiopwFNBXc5nsY/pkF64Tc/2DxiQP8bQatw17hWXfFdJbM/RwI2gdHcEfi+B1qBx
ijNiON5kmj0kJYzjQW/nQDxgbxB7HqUooMSthV7GKxL2Y/+wQutFMnxAkYOPbKF6z5vVPBFzpdg0
FtEh5PpVwK9B2C1e/5l56166IKD+nmF63MUgrv23BYxAW4Gn8YshO6sWUqpRKs56JlOn/U4H9sQI
JwtYSBsx5IbBaXZuqdr5pgE2xQig7KXlw9qswDgpQQrCW31hOx++Y4Rq3qJNYCXzQcsm9scOv1Sw
6Tbz8tfwnI0pQevnBNRJWNMM5NMOl14ROnlnjXODiBQAvGd3imtASTDvPEn33ApcDV7MCVayVLm+
3oiFsbJhTmo/V0bYgf54NjP6awNp3+llzjVP8KIXXzN6bTWQVdH8lHv11jeOdK8mTJsTx+nYnrws
/UHT+x+dlqvcqed5ZAVoWs85agnro1xFGZiNvP8A21+b68r7TzWZZQS3inFaeC6L4ND2qwbEd0e9
Y40uSJmAxvu6J4w8GLnjgPp7M2ie03TfXuO/+rBQyOd9x/ycZHjUiql47UseQw1+HsY51/hFEp3R
YSAVvEc/38wTz4envA5djGkh0k8RhoDMazVwFkjboS+JqPowR/VwyUqg7GENOKLaRq2RyyjLUrck
+XxIByrUetFe0wl2KhkNADDb5yj6lHhwYnfMwsv8Gcy+d9h2vM6Lyk7sXGKzd40tpHzGSKtAJaXD
oGtW+pn+gLuXR1pOO+XHUQyNsyaLOZ1E2SUC0/EGtKuomJDimVw+pwb50DWqo5XL9g6jYz/R75aT
pjb0EpkijRY+wPcYbxWOkiTDVr0NtwVIigJaeW7QXAkNEFhjP16GOciJP16iwQi/GU0MkI4LOE74
5/doOsuR4qkq5Rb/aAfNDuCHU1NQhm8SMkF852D5NRa2+p3YNV32DO0Oltf6XU1GTR0oByXvxjNG
q0dgPmzXa3cLpbXmIqNqEOsOjDdIbNVJfrY+0jnNVOqEqoEp05kjROPftEKw1mYCq21MPwKIAFwx
i0B+hhBY2m14Kkh3KOdG75ilV4rH3RKz8EzMZRFhoTRV8Gv+JR3T1lzFKjG586RVK2Yau5bZfgLB
YG18gclqhetPED+OA8sPOhWi1OtL3N7lSal/j9Cq7h2wRxWT9G+OFgcG7BkpXmFiFkw5UySCwprU
EMqkcZkCBX7HYT8HXX17UkczYV6F/Co4k/L2RvS6OSmAr6IQ4cvV6yY5ztnWPdTOVxs4Bz1rXHxr
UHsq0EXYj/ZFkpo7B5P7yuJ5LxClMDyq9gTUKO8Dey/MI18fbFRY6PsCJWMdLn0NS3zk1Wf0hmz7
gP9HEYC9lhX8j5XMx9ZHqVxXjw844EltE53WJu5KQXBfKypg/T1ngIuZwLoRkFQcFG3B25gx63Up
YWrWQdEjyUMca2u+UK0fgwOahO9H5CDLXC9yBq/AGwxPjCsheQNS/7Ra+eOtjFIJI2CSvrnTUw8t
nrPVHjF2PK8JwDn5vUnAkWb3NYMRfGl6wUkuSMtfBqER8xTRWfbdv/bEYtHP1ibedFlt670iuCro
5M0Ji5dBxTmi8Us03FsGglYfvf0UVHEFCfFiWhS5+h01cZBcW0KUwowiDtV744fcgwUtPp94zs90
LEUdF6kMwhNLN27tAf8HkEMOwBvN5fYurodO3oSveA4Te2QoefevCfCfnip8rV9JCo+AVTJK1E9P
jxcVLHT8x2esFF01oeTsrTbSkb4Sv5TtDTDC0Tvz+kMLIs0CxFqSGmLBT8bfTRNYDu0hZ5Ct3xpz
pLBMystfXbHFbeRKmcSOaz+U30q+cy0FtFTyIWMtCGkdRg0+Rbz2eMgQgdR6zsqgJXoaASJ//ByS
DtzEyK+YJWjvGYnsfoVJMZtbYwKUJ1rEhk1mcUiVd4RlTQZkZTdW1w1dYxAcxbULi4EcC5yRKQZN
Azf8dhqwRyBG4nf05OMhHEj6w42kZmdSimucQ/J5FxWb/SiKYYSd6CI0K4JjZfgS6zylJ8IEFurg
0IsmR5e2PloKNrndUi+okZRcu78sbo3nFFQy21Cs6GF1Gt7ZkKOqfaS/ChrwGly57djk8Xn/Pg/e
naUlvfz/03O0B7Pto2spftHtwNnCsk3wm361u7UEekKwD2vwjToNUfy/tMc//Ra9v5OoM3TMEOHL
N1nkoZZl8+3p1wqE305AsxGmiUYJ6kuuspWCg3uJ3dTVsXhsSRD3N+xpWq/Jq8XzI+gQNhg53hBU
tJZ4cF96IblBPwJ8OoVZGhnnfise57WpnAg5TJ4AA3XF1TNJFSfSekW9Jdev+ustMOLlVRSIE5zu
KhREi5DybylZWb0bWZ6NmCwCHsmadwTIJxQ913H5LRS9mODh6OztCJuM6yJzFFa35nVPHFtnCGkm
YqthuKRgon2LHmxEsCq+i7bVHMV7kaszhkVFzHHySArD2VPc/Db1LPptij6zGUsuGjVoDCkpIzr9
Mi73mMfK5Wwyf6jLoPc6uuByzGBDA1YJz1iNtLAmy9t0PlqX5SIMbBnIbdQE338sm8HsZMJlxLI1
uC6Y+vGLahVx7JuAyTZfuKbIJBcTIULN6H/l3o1g4Hta+bQMr89eqniAGJxlx0UEM9kTPjLYXqwf
M94eeHQDZsRXGS45Tie7JhkVavgRSxzkBHwD0Sdai0lJ35HEn4LtS/Y4vhI1nkkUp8owhx+teuZe
g56HBEjeunL7yAyaP12vGt4MhjpKxzVOyN8JyuT40IlwIpF8Ywzp93A1s8apZN4JcPCaQIYkP3M8
ae01n/su3ODcPibdf5rnapZCnpohqglTxCtQqnZiAl6jW3V+iwes3TqB2kn3daaBdFgUrDS9Khuq
46Iw5n9Obm+DO38UdR09rU42Ux+6yfQzM4dWrZLz/mhUUGfCeavcc1yniO3XkKAnMwTTjlMX9nPo
4YcFz28XUObceLZWRqkWEKIw2LcF1E3M66XdLSKPvnPHABH+UoBPg+VYJN+h0jDbLfZ6D2GL9ttw
b79ypNyACeK4J/WQxY5TFhUZlxXn7/nboyQ/cCCsnDJ7aj+vhy5q/UcRQNSMfqtjwWui/PP6Sg/Y
AMbYXCM0Rr9F6myndL05Fl3MHpMAK86mgxnXV0/DfNDI51B2338DDYFw5slZQ71fJSd1hsSeXDhw
IRe+YlYqGxiZn11J8Xb7PUeWuM/x9Cs1qW6JKWposg8xr/jilshOxiWOm4lYEoEtWrbzNgSHXk2y
QNrYioSlcK7TwVOiLrJZctUvvi6Oxa22hZeu++x1wVKV3Up+rLPlsZA8Df30m5dZCU2rUIcHzUfL
8iXnoA9XnVGEMGySMioO4V6L6NonfB8aYUSAQCwbnKdhXP8N6Xz6KTpVSJFSnxojaZrlu3NHx5Ip
irBqAoM0NzyJFXgDVrW1yFrruHncHVXpjD+lQ/tyJubwys2d1z0YgP4R/FY1NhkPh83A5USOpVW5
FaCdRZns8pTuD9GzEPpy9QW2Gjcd1ijyni8FhNoUQVVZ0AimeDqRKKWvhapJrlAjLoYeUVnJZ/Yd
wB4hc6GClzJugUUEhvnx8/MW8O6DT120TGBoism0ugvSEAYGdUN/43TmfOI3FJL4wSktlnOYS5lG
Zr5WuDYqlOJCxdc1Qd/K6SKt+q7sq3/zTSN/YfXxuFC9Z4J6oYXTG1tMVYayypgtQnR9VYhehaEA
W24GvZQq3mLs9sFTukXBl3zsoEd8NErUJ3YA2u8j+PbBPErcJuJxrMJIO80g2apwxWOhOYo/v0yH
ThjT28K2SUZ/kEy87GzTYm+DAvD03kqBIrwtTcUWP2zZEZzVMsshqX0z9YZy083s8HtBmVdLKGMa
vN7ObGmMVQIdaXZ6fKFRHK3wnKjvq6Vco0MjiVUSK7eXPrmiwfCwoVmQ8MmfmsDf71ZS/7UIGnK2
lTqnomkGIRP6YI3PcAoK+xLJ/tKpn9eb9by29zOdNrTjWP0S/ltNPch++RPZNxjqpteMbVv6dq/V
YZVIxIg3hck3d5YAeRxxa/n1QzTBM6bbSYwxVx50u/ZYn16UyRsWU0hKNVG8E7OWnDsKDYaRGohg
xZ6FcIio0uJefEMLPo8F1Mt63AwrPeqZaSvJ5LjdiszHgQaHD+mfY1LcFrVLQVmnd8TmwdPeJPfZ
6w6/Nu8AWutd++d0SsVpcjO4bs0WxAYXdybqke23yiOJO/NyOLC2jjA5ub2mD2kf/2WevR9OziFK
GFD+53abBYOpXrzGjF6XAt/VwuDTITIkw0AH2uoUJ8M5ohpwjsJVpCaGpyMyFHln7ogwTw6CUSE7
PUF8GmKU6dNPqBpw/HG+Cp8fZuHIrM8F3ipnmmr8n0tu27oUsl9ugN2XdbZwc6KcZG4Em8Ql90dn
RfH9gpJqZPDZNoCsERmu9lUJT8+N4UvtnJilBepV60SVWzDTU0KgPJ4c+ebjw0YFKRgJ+VBox+Yt
SGrqOo6hfqyU8tkEqhDOvNEviRUFrxEHIWuk96Phs5apIa88oVV0wvqR40dMIhYN5L93PY6MOTyB
0hxR1LfwuCBq6OJQLS3Uld+o3bZo8g2flvBLR33FIwIdG4hUFFQRxBCgxNr8f57oIZ/MTQ+0GfKm
dYn3wS7XCkRWvxvH2+KsRva94T71Uhdg1VCgaoJvBRlB+HmtBVkKx+ied1L9p27yaAZuEc82zHgM
k/bvoeNj8k2nYfeK4n8+mdvuq5V7EBqBI8imBWbjrtMly3keTQ5ccvO0UETqrGvpTwz537o8XBxr
iQPxi9J2OwGmZI09Q1ys50k8F60ilAc/ZVqWIkcy6fR4aiDA8Zbja1kWLgZ+r+L/oUIvVL7sCgqi
WBr86NqFs4hAuKX5p9WYRf6ll2Nef/O4zmA2pFASL3yWFfk6jazzurDiDTFOz6zEAUNCUFrBG8x8
4eMguN5UBHHFi5slE5DNzbxeNpMMvlUME/W5ARfRrs9xQej+jRMh5Mz7JsPIkcqPPQti6l/lZsDZ
HprY9ghIe/erUK4LiBXliTA1dJJkmFO3wJa9Mm/j3DOjyoOg76hoCfHfVtoOmb6Occl/4WBdtGBy
808eRrpqY8zbQ7q/5FQlu495Iz1mCsM9MPjoA9DELM2K91aBr9pfnI1iYu8jNgMM6jr+8iKc55VK
2EvBpYtcbs3GUhwOUY1nS8UGMEc7C4fm85xhKW0vAXVC/IE/tsnmMCiIuVxyRwkN1cHyX8B3kw5t
ctDOynAfYJJVmHLMkKVzxqE32OU7GWS1fNNXSW30FNQWx03HgAUQq64ywtsuZ0kSmVxccIQ+Htqt
hHAzllY4JaCokNyOY3/R7/fNiq6kZvqbVRxbrhInoxBeVaj7Tx+cEmqpCQilcPtMMgXF5ckzB7wL
4Ix50gyL5zsylhZU8pC9qNwly8Malj91gLkR/cv0ttZsdSeJPLxC8DJaBKqnXiESFNvdWh667fu5
axkPm7Yiv8iDCaVFRPbJYpoOXJQVkd5IA/NX3DaYETPzOfb/5TJ0wq+4K785U0YnWY0wTrbwR1k0
EeO2DPvi1r5aF8N7voOk23oh3LCle73M9klaXkLmAUp5kX7zosX/MiU9MQBai3wE5NqkcUH+fy6B
pD1MovemUC7nqrtHl/RqJKVhBEj5Y5KN9XAAnAHYx7XsdjAeMtB5+Oqye1zZzEsI+4iJd/GLgDYR
nTUDfE/uVy1EDvx7IMY6qx2wiKb4rbj6A+eRwgF6XiTffIpDA6l5awDFs5R4o7L5p2NlKqEPThlP
6cSX+Zgft7r1KVXCSn5w5wHF4fZmkxYXogf1ISLu8r0dmvUq1CgDA+GDIH+cOwFT5l27poy+EtLs
tUH7JsN7Sb8yZJ7PPA+pWtcA7JY5psFyUmEWIDOhvjYxC58Jzg5HvFvNF8oGNrKO6c9Ljt89va3/
AeyZtXUjlzsz/UwWD3UOJUu6yB6Pnk6PZGs4ChLbb/ThmfA6ygg577KBQ+iHw0kG2Ru1K5fw1cg6
301IrsWlvTg4cxfG1T3G56TnonGkVP9DDaYheiRX+uivaEwdCX/JKe9J5eo+dDNGFiTY2Tj2BEzz
jINGpzb5rlaYca30biPOpU1H7yMva6EGWaBn7KOwgb3YcJNVqvOBvIKu7I2Er8Eq+yxjLueIsktm
2T/upOyG1Tii3S/cZ+Ljp96Ffj0fwL2ryIQ7CxAsdDBTWjGKhypJEAWwD0fAXUbDtkRZFN0Y6xkx
QpjzjZ+Ix0yZExlYh3GpZp8kXrOdPbKppfkY0BRQuBavR0Wo1ZeJOedKztTUt0pPYxAllTdNi0ll
p4YFcuny/6mOl/FYaHgrx+3Snulxu3K6eZVu2njjrigigzuA+nP1ZrJPS7iFhJWDRBTfR+SZ2T1o
hwSn2oSr07vxzgCg5ZH3tkJkjEav2kwhMrLTljzFrn3iiRqSDrN4MU/Hrz1n8hozxS8t3GB6JzEh
keulrxDlhAk8K8aaaQin5kj5eor7AL8TkybElm+riYCBjiZcg4h1vL32gWNas/qRlyNYhOderusA
ziqqZVZs2rBhUshg9hRW15dU+JX/O0lAE7E/8/d9UihoPzncTC5nWTtuYPLAPkPcS64k7bRbfVnN
vIza7QXdFy9Vj5sgn1M9lJidYZg2YMz+gCLYz+f/o5NQqbY3PAO+Wy7OYfdqFK18Jx8f8TUHDqvj
+006ENi+11JIHJ4QE4Gj6GGMKIcNDVpF+3V6hY17wKsZnnzbzONJuBk9XEfweSHpBPQMHHaEx1N4
hT9g5lCWSbP6Dr6Csf3/of/S0x9Zw0CRpmHsuXv4zzbGCqUe8iSwCBNipDFoS6DZPKiKISI9rbCL
ODo133ugcsE1MjJu3ryBNPX6phYk8FzgaPjX9n6fgHe7lfPpcmFxeoq7yAo72QsokebZMZ49yym8
Ev+4P48zwBM41rbZAtarcU1GXAflxHnuwovBBeowTYpy/35szMJasA6nuhwgspegAkEjNjG0uATu
zGparbVxNJFucu+2ss1Qd8fxd0gP0/hGzIJy5akuaoPu0eV6Mr9TP+mPlRJgK8nuKnI3/8i9TTqS
zlzFCWaaErxKyJ84KUoKDw4EqM3ITnbVP81QFYOv5SKzKSKjF4Gzg0xYqw8QaHCFWIEX2YIiVINw
1O9vWvXiiHl62FOtifb4SgiZFQtXvqExab35zY0WmUaUR1r4F35fezH6BAWHy2dkrYf0y5ACYx1F
+PcKSASWqOuvcs5TOZc3/hwp08BiKJwaGHJ22PohR+pPSJtgo3yDw43PtBnBgQeocAseuFeg7DMb
ceOe4L/sXCZYa11Rnl4EmgSkIZeKcdbzL0UQvy5XZXoUqQrdZjnUIxeYEGSH04RzEWelq9pXkOpJ
EpQNreEv0ivjnMkA8sb2JATb4IT/+ca77ooqzIIwTFI8BcmbpIUZGbj23UlWtmL41Mp69nkMO6uf
miTXCmy/OUbtnAEjakAv9D3FlodK71KdgHUheLYFscNodkAaJAsytQ46gjp33lFJbKcxawepxkzl
/Prvu0sDv1vR7xkgNMEE80FBIjjkdaLbuA0AMw9I6YbFJ+RRo8OUGYKIx70RUkGd9fF2Bz96FaK4
VkGsoZQ9qHPwHp/0GW6aMq+pOd5ngvsZw/9Rf2JyoSJLBpDMIkXNwQq6ZHJW1FnIkLzEWAPEqyMa
pVla1Gun/8IQBkk/2+CgUqE4n6Aw9V7BBwL9Bm+LRzK40HuBeBmqDeDUgiOtkUMxTsR63Sa/RMfZ
XLe0Y7SLMsyuLgn6zhb6QkhwOv91FiTdVbLqdJyUnchP/O2v+oksIn+SK2wriEoNQ5F0GvdPDhSi
/zCXRhTiokCLfYXqb7S1/N2h9Xv4J9oHvBqVP10oh5RtQRJ0MNaVcZHr4eEvS0mhtCNRLzXH+phs
4Sm/s//r1d1S+vkqTzlAkiWO6oWNYbkRLYVjAGA9nt2l5GxKbbQCax0fdP2Gj71cD82JKIkmUK5C
kHLQwPiMapHngufM5TVl9rBtgd+k3NuwZG7I7Z+q/jICUFv+9pNIbB9Jy7uQuA606b9IVOH92qi6
PrzKHOqZd2f3fHz9E18gBP9IrBgVEbBNQrC/0JKmdyh6Pk0Hty3kAyhyIQCBQ502UcqDx460Hoaw
QrWMVGyKf2lKyQMQwTQGw8R4T5DJ9/Sknl+Ygwu/QZkQFE+kwU+2qYXAjDfCDgm8iuz/mcdcmoJs
5TDROC0v6f3neuk/d+s748pz8QzP55v9ut7HRqWow42/GjiVILlxaUkSDOgvOvU9NDp1j9wrEtf+
5Ffd+s5HJw3Q0C7ZpWcKlW1+XaZrawAsBG+NNjcRtyYtNqAi7MQX6g5eNfEGZT7NskDvctCBECEK
K2AXko/Ixi2iM11659XG7PiH9jqcVIJqjMw2tfRQDNGD1Ma9YEB2Cv/SWB4cxE1olotdELFQn3Ql
yq18SK3WhtV27tf8IVzhzcdfpybmfhTH3gV3jTVYXYqHKTiwsDeIIW2KppCZh8CiU2yIHORFXP9A
f+MdwvgLhJUak2xHTK38YThILEXyZ+RQlQjdO9JLnMEuidQ/fg83J2556eP6vFVYED4asezuqQ4V
3HflyqUUMsVLmIALfj/yD3Xx5Mb4ir0uJBnOb7+L9bePHwvOxLtHquwPFyVflClPJGmGqfrwyLs6
LZojbwbBEaVejIFtsJvkQBgA4qm3qMsQQ+MLOURQtZXGQK5lFZ6fpim87BRfMTPRnju+00CtC6c6
fIvT/Uczbm+Iohbxn9Zm57OkXu5SF8McXTv8DRH3oUhdNK+6FBuVrrDkNfCz9SOq0w2GpIA5P59Z
dL+GI0h034xfjTf565Rx8FDu9zQlrp3citdYOuVqu20E3TCsyVK1y0If79f9hfJ4J7kX6taAEYQ+
HJ4GBMQULbWOgHndYCuo94NUDRfYyUuzMlp88myiLrrFMhA1VUrf23kMNJaUEcTxqIAFz+UEmuYc
e+wV6j636nGEfNnBZV7Q/dedBl0IPWtFlqtgU5TrVnDClq1TXuuBZvnTcpepKTOfStkgZjnXJ2Gn
P1LVjEnICZpHae+Ld9yMQga9tG5eq2yzMYrGZTR7qOHyrIJwtoK/LRbNoiaYyEhWQ+iqo3+73APv
qvD/Edy0c6K50Rs7W4Ks/J9tXjZ9xdvL+dbM9fRCXIjpk/RBxZoAord9DvHidj526VGXuKMaW/49
hnpUG+/tiKtUoRr2DvNwRxRYakHWC0+haYVEPBNQVOU0AUPc2Z51Ob/b5aVshxCsedmrIAsNChUV
FNlcxlLxr28vVQdQuBtfq1LCyHqfNsI8Qh4v2wKUEITwvwjytqvWuyXoD5uQHibse6KK9M5U3Cf1
BwY9Hwx56ZSrLjzmsbvzwxTCxSsXOqsHeJycXw4NOprbWo8Jkp1kirvxP1JE6hfBvtNE7TuDyDL8
uTbAn/17AapZ3jTyW7zx+WsZB9qKlkMb8v7CBFC2h0j60qti9dzA1sEFyaRocb2oH5EIstk9e9q5
yF6gruVt/GB4niBcd1t4wgJ135mG0LKYhJ3SMbM3X2Znp2q9VXElzcIDtcyhrtdAeunYPMp101FM
O0JPDouP2ZjbyYhgHzdpL3y0N5n0eEBKQdLWxvYPAlescZIKzlLoJxlDdpFW2ZTut0G38ln2c4pn
bysDhItQbj8EvQVidXCDpMYcnX0e4Ixd+6lAH5AjRczYmeR2syGEdqbyI82DR67kTJp8OSAD2Cgn
a8PEAcPI5MpIE1742vhkNPtIceh2ZVqAAvh/THs9gNWYp5ZuTbwyXk3WqTCeB7DxGL7xsXiyhjM/
N7S/lkFMXk2d7JzW9KBK4SIFENx93mMDKlawM3mhAWb3MWhdl+OX690Kj37wLjn8q4VLH+QvJmxO
b2GYaKtQXpaRiYK/pTa357h58K/C9Y2IsH1a1vXokazUiT42GWDMES9eVnhLyfrl23RdYdLdPBBG
XrdXNO0InW+SQRfcsWzcnLjJ/XrmssgZxPK2T35wMveLQZpc3XJc4alnJkVNtMQrR5s413gOaZIV
Mag6Z8hRWzN7ckb5iivn4VrY7qg4sKjr6L6MYfb670WJUJwI6oXmiBRKMlorWjc9CAzU3hzhYxsl
5TsY/RAC1nY7xS5Y5F7m/wfcwQURI1CxbvRKE860G3hVNfKaagMF6SdeGLfbzSXB+JMSROpSWMES
WzD22SsF/xPEqWCFIJgYXU9iCdWCkGDxN9FyDIdJ+cKqCiDcjgi3ZpJGjq6Wy4MjN0Y29utE1DoJ
eCJ9NHV7qPvBbo2IEvwejYF6OpnR6JaKG7pLzOI5W+xIw35gcy8CrlGHUa6O6AEpbVllIEPzxi7E
WPJUAaFMV4ATY92tBCYUSHyw8ZJKBTSd1JqZC2c2zGg4NI0sxfejHfiKTdBjiKQxDrcHMLenbzCh
nRwO0shkd8WIfx2hBHjQu929Jia3f8EwwaTCfbNMrrX8q7E8inVkrr0V2B2cafvJhuj/QDG6lQDI
po+a2+udOjR+RD4JfUzzbaLDmiVgjDInyJjdcMfatVr2h/Gtc3pbamHW+tH1jkdZkBTc1pQqY3lj
gT0TEKhJAgSa1PL7QgMN1jnVOgzzKw14Vb0lh5xR/KMb4syiNknlMwaPeuFyhLpcGC2UVC9hw9dA
Asb+9ybEFVytgUsOSRI0m43/ChgBJGt3SiBRzMkPPNqxhPLCq3kU0lm1jLI3R0FMZnbuGIilerLt
kHUnxfmTO6cShvlFMqArIHDOGGFS31YdAM3yzGvWAYePc3ead7kcZxGyKQWuGkgTd5sUlrt6I43l
ZhCRTBtX1jG2Pn3wWw4Befpnhu9nXSWDM6BE0j+Vvn5ilrjXBpMghjOp3ghmG8ZCbxEA93ksuhu0
/ep8bQX/cQBtzRED225Ym/jWDlk5o8D5rvsvokowtyEu4dWiMyXxUWHpknerTxLv+AV25/8ByLYK
mn3k01kZMni2nNyg1PbPmCZG2CoyOiQHBY+rcEkYDmWfkWvN2r1gu6N4LF8/0xbrDsJqsGVnI/Qv
SrkIgP/BSUhmXHrX7Qo/74vLv86ffWNsXzgKJ88y7GJU1aKn70UF8GT8pOpxmD4gPcP9ie4GP+dl
BMfg9xKQM4m4XHxQXCyZ6X2WBqwl1M/tS9iSdfxfkJHj1SCUa/REIQ1343LQ0LlMUcJv+zInc/3s
19wKVCO+eAwEK9Nyz1CB2OVnL4z8ABdrkcCg/9V8T6EVjCUXELjShl5FP3VeGR96oFGDuFnkA4cw
USGAKxOOihkMMaHXuiueSvf0D6/SNBOrOq3aXNHp9ybCWPYMyaXBrw5UbBCIqjD52sgeVnwY6wuE
NSFgxol6wy6YBWmM1gjtXyEWnwHhFqUICMhsOY0kJOaOLB1rapUip5aHMBK1pckBDPbEKN+C/Wa0
Emq/Oe8ogLvdDEVRo5AX5xO6DQzbt1S74R6iTxIplTQFb47lyFOkNj4VPwPkvjhv9k5Pt031fxFj
VLL4jk+jYExokZsHExdqPm8bdnMfOEV7QBBtoX6qxspjhRJYvc0Lh0TsbibOUxB0Qo2TuFGgUdF+
SLbI3/J+AvKsRZEttx1wQyHUjSa1TAr5PyOsmBxMukGruFBNFaQMhrbml8AcD9mF/9ryuw1Qms7B
yoNz1InnU5mUuF97cxHKGswBdEKKN/LY5w4w98dJ3opEI0bcCqWC/loBm2RA/n+cbiOOSuAtZLEm
TaHQl5Dmcr+Xs/SVrOioLeBY/F/l67u9Y6N9I4qkxPBnTBNXcJJW/as4ZuqeFgJvh5AAWsRc+Rbv
6ldxwiNKewDkrI7S7Jhw0T63c/FzILXFInaKMdSMsGRnTsj+JwZFdRiJAbgQcBqyo+k+KruyVWPm
r/LLcZt78nJH9AZvuGsWIFbwdBGyBHLj0hCdkX+6L7G2mklHhGk6zaTyvVkv9EzMsMMKKFegj2th
SdoUTHPf1B3ZvwVv/puDOPSeF5bKX7vzRNOCQ43F1y6x/X/24ifuaE1MmarzwvMEc1jOXmF5x7xM
MEsgc3HCP9UQjMy7rZ0cQ2eHdMmzgchPwxTf2NtQdZTxHhvzwgZj1egjDkL7b0HBBdLdFdfYZLuc
K5qJzduUOmRHvRkmrZp98vCatFZXuJShHi7Y2L1UeTRVQDXsFemhmW0FsYkOrExsY6EG3093Efg0
+mdeanEumTlSpykd/zuEEov/RAz+p06d/kBn1V7rebdE4ZUE/C3TUzuYT6psPTU7ZN92gNpNNuFS
8dMY9DeKFQ2pQ/0cfYXlymG1Q4pMy0+z2gEiLi+2++oXcQnyuWrCreWyFFNdLJr4ugPFkzPtjFVO
M6F5u7DUkBKhfcoeKDSvcuFZ+PIsolmmQO3ox/7hBhelRMPP1NUyf8O+7iaL9Gy5NXNgy1JX7MGW
ZfEthBGFV3jcB3vkzvgAs2ROHG17Jypftt4ukDTftpBvdWXizTCk5g5gb1SKMlpX75xZ36X2iOCi
6L4HDZnic6xttrubL/jbaGlMxPI1lV0z29IhgoHMcY9ZkslUSASJtM8sYy5S0BYiZnOMQsg++E0f
c01h0xI/Ie8Be+YMyjFVEupuvQH1jCAqF60FDyJe4hjySCh6/gtfJqda+RQ7XXVAKYq/dWlKAsjL
byVRKDzaVDHWR26Mv+KecCM9hcqbOmanZdgK/3A0h6pogfcQUerJ5waBV/927VNkBizaRcPCqtA8
uCya/6Q4Jw2kzheSzIreT+euVDH96MwnMnR9wTqm0J5YUafcw/DCDe7+jE6TVsMcRMnDfjmdO6R9
6DwhmPl5V6XtTz69yqfLvcQZ5h3kH6lzniSgAfM5Wc2pGEUG5TnrlcP1yXnJxdZZCMkiANdvvNNp
GNfOTITaEsFHpgtxjBilx5Yp1dCYI5IHSb1nfYviER062FEW47RCV25u8JUzhI9SlMK/nrZ3DidD
+7ffbyWkdu4cKJ8wVLOuTlG+EYxVngfb5fLaczyILVqCWepsn+DaDSuTm/Ba/eDZ1rDM+Gv+ycdE
2drGDz6SpfXiM2MGE6LUZ5vYmw6CgoTJjcMyY1G8gBbQrOL5KT/ZL9MGLztEyK9aEkmtXLr6nnCw
4hBeyiHNqr9fQF8SJ0yJovQWQEgeLxUAiExFwN9iEmp3nWtUUxgliNaeOyesW41tIT7Nkj8lwu2v
WQoSDutAbUR6sARHkk5G7zTIFPDXXWhFUp919Cg8koaxeGgZBQUqxek5XKR6A2HF8JN/R1FNYOYT
8SQLrpp+mEOMOoBdPrINAH9Qn0C+ngJjeljc63BUlA2OnmmEANd8A2BMZIuFWpsoReQIX0DMk3xz
UrsoUy/JZKsg4JJSLIqBUEJEYUv7Js7oNbYW3nCMPZhXTdwjVzDTgMXO7bfZ9+2Jeee1cOHVeKYx
NXlsiyskpmfG5vYHfbinuxYgecuifgPGwRouGB1cFroxGtg1muPGfAkpLdMlyYvt1UEJHZsyx9ZS
xlqmUIC/uYhJkkqZjSVqjy80Sax7wqww0VJmb5PzdfT0VDCforVRiKSI/T5xaYQJ12P+XJsjuc6d
4uvqF5p2g89QNBXxueabJUlUDGpvUPl0Jwn9ikDSrGSPvswIooaFzn0JjUk50WpEEopS4lQXcQaA
fgwrHYbkdQu4UzFci2GjoYSNOPMv7N0O7gyyYmiTQTUCoWbVaiIBCN4EXReulSqUoSbkHPCoLc0m
6b79BDsHKz1PJl164/uM2ADjZHa8pnlbZ8/Kj3I5nStVDhcU8CCF4ADgbSZXg24LVQAR2BsEJpHL
0VZlJgtGtSxb3pKR1jFLRSlwSyFZqzIPPgJF9M8MPKIESzA9pnIO909AOjUEeXsfBrfL4ToiKScP
aSw/hX2QBlUnfqp41T8yIxORg7/8pEd0599aCRE8VzkLDIZiZRHhjYCaTUQmPFJ6mRg39JyY+CSE
z0QD5o73GsrmaT3hOTuEdSW1tLdLyqe5qmOTjUcHuEeG1I4kxiurCBbzqNOqCByFRFMTfOtRMp39
h5f5FI0nf4PCWu93AzJDbF5nva+Y++da/Pyda4dnbdBwmZjt+feQudmcLAwW87HcXYQndvUsI4rT
2wO4xAZbYX6HHDA0+W8vinyXnHKgh62hnsT/e0PXE8Ox8vzRbSFWWwJMl1qgW9WWwyjsIBqwnnU1
qJEqtLwH3XXtbb/IspbDUlL/v4iY7iYEgWLYfTap8mmzg44kKcm+7pq46zS/czlDY2oBzG39muHM
B8e+BMbv92UUyTPLOXQyC1+r/kcZx8epyYT3kyXVvaAE8DBCWZ5urVnYtpgNb2fkiqRltVGi7eV4
nJpv9bCtlXFeUGWNcAqm2rAcLNfUlPlbWTQsaTzwD2NV5nuU0PmS4ZPOaPydkR9hjsePssdplXbE
tfwcXijz9V/XCVpXHySGklxhsVRnEVKCrtqcuw89Yr0VhK8Ct7g1kFYPr5fXqFzaEE85U7CZBxDq
BFy2USPOX83vBZmRHmGUpI5gRW+CYAKxzn2757OWfwVfuSIeqVjQXuWrk8TJGNV11x6RjOZdNKWy
4BlezYWS85YcM9SGHN8ekHdiwYXnIaOqrmbWzHiEbZ1+spRJbF+zCOS2+jyiGO6eDrB6Gd9RvjRJ
hVuQVYsW8H0SWe9WN3f2dZsuJ5S4HNn/NcoGjPNvdshCpWOtrTFJqkyMP/t03QBVGMgncN/E1Qwv
Dmz9QMq7yQKIzcxxTgZZvfn9TP/47ZCylRyPTgIe+UfTXIyhwaxbp6ncEydHu6RQtAsth2/6cx1w
/VBjis/a7JSBqqQxjJwosvnGoDf4sNPHEh072w2384EqDKcqPBe+HjliCDPoZwIJIV9C+pRrhjqt
C+aEH+s0C3LMLWG7VHqVD9wGV/T18TB1FoyDs5TaEkAolKQiwp2lqqFGeUe8LkfwnyELkNLRkq80
5I3tZJAkLo7KvXvXbUbZyJGsHuwbF/fPc2N8M7ZZS0YTE9X5GhZstJy8M7OyaTToNiaq/Hr0s2Xp
t3wAhEUlFD4yDb7H8KJXDsKFAi7p8+yAO5DAsNPw5nuTDE8UAIj7lGMQbDn6D4uHPQCLdqOXp+8E
FVd8jVA6Y+UjKOdnQ6APUYNXbybSGigVC4cCLPOhx7MP5QkE2sYqh9NiY1Riaon0sajShvhDs2dW
kpwv4bo05EcZhPj51fSPPI2eOZQDNBwdnxHKC9qxh6JtEcS0QKSlKcLAoUpDyB0z4bktj70xShRM
0b9aaMkZjMhKuuQNqBfW1qnIQUo0SL3YAwWTUiUdLF+UUpjzhyjDD6DvaAVNgf2GDk+08eoviGYq
9PXJ7mGF86ka4QL91DOzM1H8jnU8bJrdSP+YZpNjxjr+W8tM3SXvgHMqjRQyyJTxbwoHC8TpqiqW
RflR0F/zYXicjZs5Gc7sC2gE2mflFmdcsJmBEmd4REcB85grr4mUGOHHy9ZI8poSzCpZgpCUMhYC
PDByyZzqSPWfk4rcCebwkQa4bj3iXIb8dnA7f5G4is93aRsfAky4ewgAX0IBFXMyNuRovOptZJ14
14SDfIZusFJvh9VWU5rApNvUds7g1W2+9M2qBQOQ9RhAUwU9sz4NHxZFfqG4LnMfGqkqCD2UpQHb
ECQM5foDMVslGbp5ktE9YKK++tGEDCFExi6491/789sF+LRkW38Zyjp6TpbiBrd8bjORHIDTGfQO
h2p66nj4x4kaX23t1HyU8TWJEzTJo9gsF3eGswSjmXVJGlIx6AAqWwS8bzHBdVB2dvJFizc/ZMMz
goIA7nCViWyFQFg89z8Ht+yBBDM9oYDlS9LsrFAPh9ErnwRpmbztcOtAFdqcsVhcmcM+OFkgSps1
PTLgbxfj6hUt5Qmqna+G7ydn/WHfl9AesxCvdRwYlZBLB/veBIBnfakf8MkA9GkYjjOs/CdCO9uS
VV1MAbF4Z88+5x+Ndv6d3Kpaq8jrZr9jms6iGkURG5ljAPw1LFEmUrVYGoW5Pu3WXcEEvu7tBHpA
pkw5tbBX3K6V9B3cOEqa7O9bk1AQ0eLwsRihQxa/RtxqeuPgP5pGxifN4zGvfhC+xfLUDQ0Jsih2
q5YIeRvM9LquBt7DvbSOwLrGxP9iDGMlno69osYoqFYFuzTpRXB0PKMdTkkedJ2S2PDaE+77QTGa
0jOtxH4uVM+GE7r3otfNoj6u+Q1MXTDiWp5KA7Hg6cbD8PVKb99JEWKuldPdbaGrugSS6zYNImVY
ZIlTGViO+p4pCWVFE8OHCgdDF9SPSO/I+ygkq6uxpToglNPNPnO4e6HRTsNUscZdorsVBNLTAaBq
m1HDXGjDNSIdVFTQgVDs4AYD14EWUH612PCMe26G2dvMoA3UgFYvWDIsFaAlhJqu8NxA68gBE5/4
FY2ISHgKiAgB57nyWN6wb5yMow3LLd5S5RD3ChxKJsU6UlEem+Pbt/Ubg9jYTPDoUe4hDlCiUxoa
7e4lkmtK27KK15EeIYKkUGBVJzwd68n2I0HcnZ0KxIlhbxUxRxlKtGz3oMvnd4CL7UON8TcY8OWM
C02ei+wRFp4oxro5CzS+2Xc4GqDoV80rhVPcaU2jvRZNQ/vuxkeDeKlvIKR32rwhXZhHjrC7zgFf
1yPkUO3LsBW+pvlHEzx+x5qna8ObwAOSecx5n6z9avA2mWxKqLiriYymHZRJxpmfRmGHvvX/hJp1
hVrwzf3k9yyKe8trn4xCCjX/bLpUwu55ar3PC7l1KmAIldBIZ0CAhE7//mUJUjpu9jnyIn9jTh+4
kelkf3ktCXUhKxalhgmexcAcgGEPMxuWqfz76WjAnBRRyi9tO2g1R3tFntE+Df3w1ZwJZgselddD
QeyQ5Z4DCUmKAlzZxHtXidnegxiVSD/4WlEpktUojgWbM5rK1KWL0le3hfkEPECn1f4RNg4D5ivk
p528tDQjxKSjs8V5gUsK6P4fk9Pgf0237fMlA5jboeuwZg0ezPRRBQ4LWkMubW32hE1+SXnWjFWV
xLgCbXUvBOL69icOKRsvzwWN519Oy+6752aiSSwrf/pD2WOkGQO0thUaDgWc2hD54lsU7wmPht9G
hTxxuzugXTk4TM50WA8kc/3AuqEkPzGB5GfJ6zQaCLraw39HrUt7at9Wvxb79T2mBsTd+M+tXxKl
NOFPiy+L53pff7YUEi9MSK2gd6OlYbEDF6Q/yfkbEzr3rPlzBN9LBM1y1G2EM/XIUD5tvq5+zfxs
3hw5l1+cFbm6SzUY2/MH9KjoEqKiLfJhcjFbRROzRhDalg4FnEmLeVpJVJfWsSU/Frk9Ku/Zp5in
SJJKme2uPbZbm6RUbqj6HkMSSxCiFPZadjYbUyUtA+bxyqeNoQ57IQaHvJjZzJhMrIQ0sMhcX2nZ
zYkg7X4c98NDnfbpiw44uJImwOeI1SbMugChGy9aTuM7cPNPprSvUxQDdwmJrhw/msDsxI6UUuW1
i0N0XQvSaRNdWVA1oRaMG6k3b8WuCTPijZBt23Wr1hyCrDs8ia2Tg5FYyxdNppMMC8qNjE30hVP2
NoanxHCG2wHtQEgcCyeFAMm5lUPnaR/U6jWUSLa4zKVD8w25YDcxmkdU7OKSZkxnAjR/UPgS0dga
m1GvaoblDYaWJIOL3ffvAan6D5iKKQSUKxvALVl2QgEj4TtWI2PllMhtlbChuuIOHYKIektchTiO
z5X4EWPu1gY766g3iKnnEdDsUrw8ckwijhu9wOVD4D48LuaqhqiFxA+Z6oRPUJ6e7yC7rwv76Tip
/G3WlRPf6+R7EtQF4VO7hb4jnrAFmgLtKreMyJDNbufU/sDziQc69som9bsKFHfXbZGsPREynMVM
va6Dg9QbUteUkpFz6uTF7Omi3SaKtMywWcm7ocbTZDKWEKjuLM21BDicf+axFiSx87R+YSWJUIgq
zIQzXNHOb1//B0ErQnMll5T2kknyX5VWY1MHhNtwvPwmS8m0+Mvcpws8Mq6NwrQ1ZHCeNAPFv5ou
BHz3wVxQyimOaYXAOOcDa0GOZvcnUC0fRiSCPbQji+FXDpJmfSuVaiC1qEQsRKGCL/AFupQ/VUXc
YZpy5WJByjSpn1Qt8bPOAZ6yLzgdHULtG80Ybu4+cFH4l6AyljxcrxnTm5m7A5W0b/gLIe/pVEvM
awyh+R7U1Y/NUpZOaGjl7bXkWhoYruGw8n+SzXUf7SOD7iuOeSmwFvPCkPo8tYdjWq0PaQbnp+ol
wxYRJJlh6ck0e31HxGjimxKKk/Menxg9mxC1pb11soFnYLQIZBkwPkosowFULmM+4CgHwpMoFkRx
rwPiUqSaFnjbP/2e/CVcffgQ2klSjU4ps1xeZL652cVmdps9MTwrdI2H47tFs+jwYu5QSvNPAGW1
qSX3Bo4H5mwgJMDzbQiEeGyv3NwC8numYr1M9ELr1HurQq4ix8nTQIL8w/FwroOX1WTKdrbYC/JV
L8yKXUm+gbJXgGIgfaYGy0RG4dSVGqdvmEfHo0uzw8moJdD2thvM2t+ugLK+YXjeK/J0N+AZwus0
8raecBpw8Kb/UGgcLFXilbrbjYoh10JXFGSJaedcWKxdzn5hI5tgViaF8lho7iZuXXFuL0hCkKlE
khQuObLEuHIuAFynzMIfP+BLb1Ugxqz+KbyfVZCk/DRomm8KsNwqBmki7/X/92RG5T0rhSWCCkd7
h7ZRZ9WZT+XiG1MPDCSw76PkwAGHsDFZ7PDvpbtiPkeExQi9+4vUqac+xKFj1N2cWYNCTW79pLi6
/rpo3CGfhXipkLoH/Jg0vgstn/YBYxIcJkJU+LnczFJd71V1HMo7QBxpkmqFBcFbgko+rtGWt3Yu
RaiFjVAqLKgO/3s+DQveje33/HS6FLDuNzUk5t15eu/Ms+3PLmEHx0BFSzS2gXRIIWWea4YS6vQ0
XkRSMocSQH/SJXyMzDL+dfPh8/xH93cmxt4x9VBjWwntpLVhhHycaaCJzf2a1padfB1AVYqMPN3N
ryNTeFZ68o+2EkeXmZ4oM2wxhir66gboBB7nanmrGvfad/tuNIX5SZkNwDjImJAzuebI55/tsTTX
zY/aA6TqsRlP3SzmCIoQkOOmBZ9qkXsPIUTMHBjBti41RmBd7/ARkQTHO5hjmy4k6Y1IKG05Ew1b
FB6KviI3Nmb4WiFzt0jvj6Yo9lba/UDaY3b/MENm7gQW/1HmAMeFNR/eZ4psA9MWDfVYWY13Ryrs
wdrcoZWC2Ltoc58qR20dgN8wAyrr+b9EgkwikshB+4rr/Pqk9Ckuesd3dC0As+xrkZv32pmuOe6v
R4tiLtFC92iC0EREdxA0eju5dN2uT8hsRccS+1QB3Ee2wPWqVpdsVrnbQm7blPsxjM5MrLocJero
u2c4L6ICPhrEuKS7jOYS4+c+2tnAfPUvSWfUt23h7cpYl9oTORRYQKS0mnQuI5LrQQF7LaqPYwCB
/MQffI0Kr5JL3lIvzuIHQln+YF/qUvzY9xWcfSWYSc7hs4vIu4MDoxcDM/6S7Xc5vZX8+XrAw/S8
PchREKCAdtyt5mLlLkpuaixXNXW0wHEJ3E1FMkjHn6fBFbZ4RhS33l1Pq4hRuoygKhtJvrOX7R2v
vSxQcOftvnGuo6VUdp9UQUn76MvvTI42Srt7OyzTxYp2G0xLPlYnNE0DGjJdvGW06DYx0fn0QvIa
q/Y2X49fEfpMeGSnzMdw8/lULFl1HI9NJwityi7K/7PbZ9vJ2fVXrf1Xn2a2xXf2Ni485ruT7IxV
CalDSXxZTxFSrxeJNuKwGe3XXEsHOmeX/muyGKCzsss1O8Tyahg5OGJf51qoBzfP0gVT0Ophyuop
tj2OEscxhFP0KWtL4Sij6qJhOMnG3QPpvE/NspL8Qkt+WajDLhARsQV4MRJY3bjqWuyn5F0qHsfK
HdA7s38iqJn9ML2meiQgPgY2Hbswj3uncvxnPtVF43HnzfymZ77tdpoVivOTcOUL7E2orQADKYJd
KpfDPf4nu6cW3URs4Nif5H6NRVmiC3EfxkuVc13CWdfejDDPhlZTi4HHYm8uLq3CUp3Ua1lckwSH
n8e9O+2cpmt1D9/faSBTZqDMKO2RdTEJzgDQvQ3JYKv0oKoEzOybcXX6y7G0tAuXOsE8edrDWTE/
33KLSVok2R1Q7FD084oEjnhdCDxz1x5g21gfwHIBs89LH/j1y74ZV01hcOaPnUNggq8xlC43KkDv
jJ4YnYtOUL1OMst1VBnhwJJR2PGJbvEg+ZIkyzI0xxEk43xh3ldfKR/nI2pCcdLWrkd4rQf2Ts64
mMSXqVs91yDeEiVTDL0WPkkeAUPaCG2Yp0pZ70m7elFs/mH1KoOLormCompgH+abJKVfTNhZS7ub
e57MpRe/VsfCZ+YfB/vlDyXerG4DGFhT1FFPXGmMqFc3HIbU2GM6Ur81Eb4T298bVjfrvIlq7M9G
HaMHC+tRRHMPoEFyHv1WgGiYHU1IBcraL3wij9IDQctgNeKXLE7Dv61BSEjJZ6jnZvwuZ436sXRh
7iELeQWpD6uUcMuelk3TRH1tt4yIAvXoUXzc0nLn+QDDuT4QUwQ2e94WMz12XmU9v4gAvhpkwqR+
L1IQCjhAtrOUEtZj4+cVDrDvciiNfIZvyWfZOqRBYUO9lkTILdfMLOKrvy7JouYIgtxz1wZQl9iJ
TXecO/WBMopPWTvOPzqUuA4uQ8CR98xrkfRT0lBHCCzDu7pvZ5OfmRvqFJrXvmImhRaAyeHzPyyM
jer9M3UAcarSajTOe1Te2A9ue9TZ/2XyX0/k8pU0AhCaaHYuSG29ZNGNDqAj4rrj526MVx58DkA+
H/NSKbXksXaLgN9i+t8vW5G9VQ+ujK3xwD5sihX461WAFykXXgL0iOM9naahFvbsFvFc8ZMEI4wU
rUM35nrHgOtnJ+Fatfr67gZsManZyUFf6o+E/YCZ6yczloS312l9HoqteuGoGAD6kyTTG+gEXjpV
W5TiMJ1Bt43xFJKJbYUMQqAw2eQe31qofobmkOMcyWosFZmiP6TfEQ947hlppqPPeFuiyhETPWzL
ZHRp51ULTVp0xJ7g6hL0czNRTj5eg3iXWSWu1Ufc/QLy6TQZjOePlRQv40M3IE98y4FMJonmD1KN
D7fhULWPz//bVEGA3ZkACQvACyKMIGIjNMKvY56mvaHQVct3bDh1beMkdgp4k/UOiNH5lJwqiGHn
+KQg/pB3PT2QDTBw9PzoZEqUyQvomdt+msDBmd/Hu0OqGbBgI/1fiA1Hc6xrVyhaRieYQ9M0jIA6
QK3Pa827ogLNC6VVj8CQli3VP986UToldgdhbr7JR9eBGu9i1qkg4wgLGwtf+e5jyndYrRzbcL61
2RzojViFv3GbCHVae+v/ZcCMgjG9ZT8U+dtJKxYV+5hMreTCLVQ6CFCTLCEqQAIS2gQypU7ZJZyx
dFUNW1mUa6/tYUcwd5YXJH9fdG9WBCdBMW9U/qSCaRccVLQCukPGi+eW4JIH584u08Q3uKFoVW/v
HIqYkM5gNickWtLECZei0yDeIyoYpJXYvT2zzv12DmP0QnjTHtJKWgqn/zIX3LBbajyarl2EGqeC
THOtOEhzTOVB3BvAwEbLkTja0ag2EkIQony+bkQWNvWnX/Bo+q6aCrLO8yn7R19852HFapogVT5R
52A/cXOdG2BTgTaF1z0QtK8ArD2NUi6OxJXLe7X0e139Nin0njBRj/BG59My7AdsyVGRIXAucblq
Jglyh+sawuGldZx36XhOZ17dlzb+1UbK2blV4aP/mQ5j8qLIfnY5Fr48UG09Qk79UKtdAZ+r4qPQ
gHivvnxr8J1RTQLf2EWvVfERZKhgSlWeGcB2+g10uwasPckczgTA/Q0kot7w8QFz/8KaXm8G/5Nu
8uGrKCcIUzn3uqRrJFNphuc2+M0PLRrWUB9xF3XGpNU9PKhQcWvTZjKtiuNr4ekbKOUBniFaZxKz
fI6Zg78xj5XHmQKnZRSEYzsTON/VYYvjdghY2jct7XlIrzoF8U1D2HGwQXUvlwGNOFS50rbvGLNn
rZ72wi1kX6iHhbzD/62AG946vfXHC4gPrBI5Vb9VrlmIB7a12I6UmVOwIK2vpuhOnBdjSPWFLAxM
fyhw7lEP61tEoscXVXpuKP2acgqMc24qT6ANfFJgvpKDr1fTCER6FailgOnKTUx9d1BGtwmq1jeG
gVxRdT73Ct7Tai/i4kS0l0phl30ESjedxvhVG2Ef6RtomorbkhvV0DraT71STtNDg8RELzHxQWlA
dH75/G+xHiSYeT9ayEcmdyV8UmKD9F4FRohc8gDjrtt4okmnX1ftQNlsMTJLKgptKX7eWLMlldZd
Rk8JersXvASfs/sd9z6X+/GL8f1cJiIQ5tUEsRdAaObZzJ7krwSFQW6AVxrnN0QuTsInyOiJCAS/
0iKHEMjAYsXXIAWbSX0A6mVcMdD1lburCDVUhmLvQzJ4RsdTBh5q1zZmN05kdCo824vG8+dmkYxK
i2yzuTUvEg17dl0ulnJjIgoN5jyeJVOTdrxEfIcjOU6HUUahoet+qGA/eoCrM+FVRgeFqgZBwjcZ
AtNAPv+qzbYjw0v0h8KJEmw+k08FtUXZI0kbdIhaNJ7BFoPAI8KtA59eViZXmmR9fuw6jLTENm87
/m48gz2pFSfdxXUAIXlnhX3qtrpnm9npdyzDw/d9MEYt7X2yq3vCkRVRvQrcei8d0vpeUe9U0W60
hO916mx7/DHXtsPT8LckMCqt2GWBXiI8sGoAtL5g1VGZVcAA3xpXY7MlxLNu18KtxuTyHoTkhE5Q
RdftW+++EbHzke8q6gGFsXvrOvVDKgwME5R214UcgsevNKaA7LrdUDrdieCav/8Wb50qYGWbGFXz
A6j0+U+FtYUTuSD4a5Eb7b8K6tiB9j+NaZavjLx7V97pyeWWOb7qwj97fi1whIU4bjcKxEQ1dxrq
4l5dZRECjI0Xcg1qxdSGjDrxQerY7OE9LH6loL+RbraiLrVPQUhkZlywwnCZ4dg4Znm6GpDHtTxG
lGSu+YrEANGVSvjEZnIfwDbLWezByxyV35VLPRK4Fw1y4nKuBczE9dQDqmEV11dhZOofxO+bwEUa
G1ps0lPq18zTMHGTS8jo3zlIwYakAqWpQywhNN2jSxvlJbr3HOTv2elCDXdyaTu8av4sXsiYB3XM
a2jFnsVbYmde4wONxTQf5W99UjedX/7/f7vPFtcdU2nFsTvb47AamRcWOJAqOQyNVjW7L9n+tjC2
dRWol1AZkAR79R6NMSdrYZvvOLqcRLdt4bE9+cbML4XljLI6VOP9Hp0PcmhpR05vAHXpyqhaaiEH
FpYQG5aTupqQQN+Bf/1jklwunSpzWFR3dS2xLwCDiL/iPEq/SjltmuGbhsM1IbUVdzh0vzGz6Vp/
ub3SdxL+0Cb1u206zqvfg7kop1xarq97nv0XAkpuvW6iyWXPmjKzmNrjc6Ubr9OlxKramgkD7h5X
i/yv051aZ7C4MCAHimon/YL/HgMlbVEzmQyPNz0/1i95exElgEVJTWKnycJIjGVMRjBk5BtY9XMm
KBckmn93R2HnPP/C3QsXfJpjVqLPWvhCFe+d9l5Qq+CF2vwP0YNV9RzYu6qw6f3IVquxxJ1KGwVY
sL4gMh5w/9ID7iHVnkiToDBvIfXkLVQDIZFKMPO5p+FAXWhaRLfNS3V8rYG9v/zpU+GWtUDcDA9J
2XWacsE3mpyM5CwGDSFHROaAXzmRR/Xl+QdQ+J3u49xFopl31h3clcZUjNfgeJeFFhgRLB7vOAY9
Km/lXbRY8KXKPbe6jcAh+0KFcExU7GfyUAGMOt4lveu77cWuPHdr2ThzF/krfXOe7AI1rT6qTeKf
ema2Y5KGI3AS8oAic5kLfTvBCPO8Xzi0gvGk9Ox+qiukKXLa36da/AWR+GRZwTx2ZuqGTCyZHgbj
Lkv4u0QxoQkyLaiH91kHcXUm8zuHSdP6x9AhXPAKo9hw3U7u4ua/tMHspX/LdskviY42oVr8e8ga
LCryQfchNeXh2eWe6VaBRN26slrHg9KR7xfhwybf9m1i42Fh7DhSkr9rftGy+D9zmRm2oyzEfF2F
Nf8o7TtsDqUYUBrVh2lRqZiIPWsnFsDqD+Fk4Z59OreIj4TuTc8gJYUv1aNW+0LA/u7kR5yxZUQO
rHmDIaMkoX6w+qoH/eryE1bgxC4UMoNYYzm0+RAW07wKWYcnYgpZW9PbZGFiaAVG8koZUssnbW0D
FWx61k5h2x67fEbN0v+KKc3Dvm7l+ZaQUsbbNVR8r7agd9IOl6L0XgLvoLPOTGw91/dnVMgFScve
vbh0JoLwBmDe1Du15mcMXAGYVSDj1WuuaKDeH0509cqKkyqMjYz49YHsoCwwN2ceBHMEowngymYy
CsedMK9bYcobVcQqMjMTRnGwOG7zuhN5xPwMvs+L2kpTKnbmmqTiq+6lJJASsVmMAh655bZiraB1
2IZuCTV45OsnIvKS6duZG8SqdLiUmRqF13Fpb6aFl8zOxLiGbllqpC7VPTIT1aL7uPxIh6tdgKNN
dE3TWIJGpfcjwn1IMz7e56bgX86FW07OZhxb0XtvnnQXGEoP+07zkmLS4vqADoBz7qCpxhCEnIQI
tv69uNa2Zc00kE2HIoH0BShbjCfxFjxZjUOVA/5fmg1K+0s+dzLPMh6Wd8bC+c2kAaZt1uZGUz0q
oAWxdJdh+yrP0HI9DrARzcRC+8ln2XS7GblzmezCDxXhYme5nLFLbPCDAM/sP4VO+ChWMBwiNFj0
46J3AS58IMfOyxVfV0okTM8tjJg6sAZcLD2++OhQwqaY2197jH4/0caLjSfuWT3Z3F+ppIEaOBfk
NYin//uAVdla7bVTJqs6tPXIKTgHdyHo7iuaHwL8eOf6AtTCfTlha53YXdmt8NsMZyLI/Eyg846R
EEKHFS+ZZLOlBUDMc9DfKP+vNGc20+bLCrrRCCfWnmFVFvMQLg3f/MUO2hPJO14lUF6CWLATZXpt
bcn9/WlspbhS8IwtuRf9Dw5zihXzJ5WLRAAfo2lN9WVbjA7qR/OjtZ05CHhWCXFg+vV5KxI2jH0B
oubEzweC+6/TGJZ1dSKXfTz7A62bfhmvvByB6tr8QeXmHV54xEszEIawskdT8NuidnjDBq5c93Ae
9YzZGdtr4xKykfKC7uuij9J1jiMcbb8xglsm0sX7xJlNNShrisQjEIUXSqBYE4xzi1xGpSUxHIdl
sMDK6KH7Yk4h/1a3aWFa013p6bBgLbPwq0v02DH2MZ4WDM1V/dnRvknDRpJbsZJNvfe6sr/hbs1k
YArU1MtOWhPhQ5DBgPmmkc+yFkYwAugIWLLRkbOt129wVZPilQFnbsJsxTie7Z71blYr0Od7d0D3
buIAVi7A7BUrBHHfntQjUSdKxNMGhqfFRwWis1UBSlXWU/23B8bQEvx4C+0sce60LxRHcrWc++we
R7wllHURXQBu5tgc2ToZ3qQ5BdMzVzs2OOaVFrIipnEQ8lOVVIoOWDAHaJacWQiySXQZbQ3j0l0q
pNPstywm3RmvTrvJ6CJOdIamD5j6DeCibq3V68/Q91P+Bb/rSeIVI5D/B3GZalcaPXgafsNYJeAw
mlC4YJmB7NQFhOyLoLo4sNtQxlGPDWdf4Wfjn6rpqV6qN/5krX9BIo+IgGw5v3UiF/kauHqqh2+u
JkOL3Pv41We3ZwiV2peu8SwI/pkg2LlGyU5EDFTZFPX3/L1MObBEK8BxcHcSR8ZsZf44rEF8vkzd
suVjeygnaOPQFZyQIwfH6YFsDjlzeT5QYBrxHsFrf5BECpKaM4FItWVPdWyte5wrPupjiq8k6Xlm
0NeW2x1vwmDUv4Ss8wn9iWvtcAhQ36Lcgs7F+OJeqn70b9e5tKebQq8ozH6RLXCA9UC6OOgVKToY
1GgWk/MMz2PYuXF6lRnLdgOaBZcl4ybWMN1h/SjGp5C6WgtxIvex71sXo8SscY002Mze9YzGDejK
nrpOYHC/k8xLnni+Jatwj2OlSq37SuYya9BcV2dtOJZFcX/D4DoE/sutbJ1ucc632lyDsc2Q1br4
dEc3U6lUuIVg3aKyCInRRX6aWfft+mf4BNnwq+FylsMJ35hscoE1y8+X5iWFjEwEn0yFP4Xz1MDo
Vq5ETlkqZwG18oL5lfVPuOQqB7/v6ssPbif7Oe+5Lg/Ss8btotOivpR8BdrDVOK5T1SJoL3VnEPe
+cnVMDlrpL+AN9HnYvU75ZmVsa9mRqOUpG1g7WTwHcwANWadve6vGUqqO7MNtL8Omt4a5wVOQaq/
iovlBpGWEpeBUTU9f/348Qh09sUggBKrk/ZRQUTZyfSKWBeCwGZaGVCRX3qyexbybmySisvxUce9
mWok6+zBj5U8D/Kuyy7zI6ww6en/Z0yBg0U4j9e67fhTnTAEE9k8KZyX/dZiEiwL9+UIIsr5ge92
lRQjHp5MLZQMQ7PXxNeyE9zFhzyqU8PZ40ho7Q7iAZiUGvHCgHzdkodg5qefX1vPlJ+PpjR+/C96
Crh5P65oYICSwD+wuSDvlUGL81yM0yyFbjs2x17VpZMEgnAHjvaTPfQ25dfsxEvx5oLTq1cl5NxS
X0oIIbMczDps4dtTsuxuov8Si7CUpV31lpSaKZcU3ZE8Q9T7Pg8LYbQK9bnAYxyf/3dBbeqrqKbs
dPrZE/BALGgp9AdlTzCfuZR1QlDoVXvbts7PNPrHszcu9eJGyLhzt03A90Mx7Rns+DCyyx+OjHLp
P/JOizYOCzB3J7z9RgYbe19js4cIq04aWOhLGcO8vkjkVBJNUY3rHFUqTUsgcZzHq29ph9A+YT9U
P1/hCtz5jpPcfOLfzYv/6if627M71JBvcgr6zYhvpmlDBf9Rnm/ZxdrhF6icl2rggxL2SWiQuo/k
OrAjY69NsaL2aq0Q4Ff4wp0khwn9M0Z2uZtM0MRXp/pAwIv6WwGDtt9XzEhgAzYtEsDueR8Jj4Kc
fJaYdAlv1t4nwmbnGdu7wGdF7YX6I5nqO4OXNCAd8UmwMfbwZfYRE7O4ObfRRalNauxaXDXmniLT
rLGwpZfPi0SP+jB5psLLzt/XnPo7v/ju0uOmkvitgk7kYLdfr4prXOESEnCt/dJ64uvUkRBwhJK3
4/SK8I4nZK+U0nCsOJ/3dWGQ/qb2HvhVGqTtNJeV29EN/rd4bpcysO1Z9KCAc7MZ5pKECaf6suRs
M0QAHoWuNAvdEOPqlyvvVcksrgtFH95WFuT5Ota8tz/zysH2HwAACoXji6CW++y37goKYqmAWKw0
hp1lAQBPA1pLz7HcdSC2BoOJjRjMZn6sVztIf2CFrPU5LDu4dzBo1Ht/kOyefqVmkjMLIDmf8UuF
n/XXEVgRYpgxAgPX91zmFKOGtGsSzNNeGoBe6xf59FwU/XXbD8ZsR82EloWEHsLWveLJstahqXdY
it2H4k2KJrLjYy/+chHe9NVUMCvK2xOSBGc0K3t+CmDVk1MWH+9j9qb3R7QODUzPVXrdDmCkbYlV
gidyXlpGijYe38MUWGcLXQKQo2l2inTaCB0M7GXFd2Atv+d3KG/pzHA//8PJ7sk+7I0uPGxhBUEX
xxvSKJOS7PWnUWX3Tp5/GYihGkHm/UKs99yoj8d+J1zv5fkypDCb7hVHGEz0tVz0k3Bo+X7LzxAB
8wwZcjLU5Cgnx444HUsz4RV/JDPUabxlN+RuTcANM7Xfm5xJL/DfS4Q55gk4w6HEMkD+kqbSu4cl
F2AgIKANaft77pb0Jbo39RGmYvlFwuFTwRjH5bSB49zl9FBL1/nNJ0ehrckZeVpegzPQxRVJXfiv
JZCRgfOLB1/e5JM3wrt7yn+MbG/obFrPSUBffuwINPkQ+W4qQjVYs1NMBvadmHwQEpC6zu8nrhw/
IMdiG7j5UXcHI856xP/1uuKFzydbrDPHhuyW1YGt9LYtqk/fLxbghl/ssjGpmW67RcshpLh9IF/9
NhVxlTfwi51IPqg4zkoX4zin4wcqWmZxufAktJWFS8iSNy7d9TmBnrphQm11WHrRiBnJUdoiXbE+
5XjJStn4TfN/XijYi8Mlg/LLpSkgylsH0aDn1HMK+umq7GlLjheO4K9SBPafpq/JXkjqqyB36FGx
EEpOxVJCDGyiPl2mVshVLom95qnpGOoNJ/XJpLsl0wVF2oopCm1qjOIqeM/6kvVvAJfOSYRYx/Jp
QKWlreJjkezitdlCbe1FVDEAI5EX7joYmU7s8MYlM98Mszb2Cx8KL2unW07JJWRG56BJGFWGaVnQ
mxZx0Jcxv39E10g0RuL5Qk2NdG1b3ldKrtaAP80WiIHLN2i+xSEdhSXBClwfHlC7n9RcZDQsCdjm
t1ogUSw0ibWzCSmSTeZJaWtobnEEiHaT+UwRHn1RkGfBPQd20f4fPd522VVqFFW4ik3uHU9HjXjk
be5Oy4zD10fBQ0We/a/EadFAMe9OwwNCTCWFi+S5PhOwegSmjOg6bWQ2zxmT8jMMV1ckDCilXh3Z
YG6UrZMPDHxAjrWXs400n6DiZLpMfKP7hlSevDVuRhQe/xKc8lYERTj5VHQiFRRwjftW5IlrWdd5
2csdARDuWKnPghWKrOoJA/mSWVzMl1LxVIfVghUl+QXwPQeFuiNodZBfhRvPLA1pntfHCbXnEda6
Ey9zw21+FKfMUecGFYEBzm+6knQYGtG5O9Af9KuaNMzZu5VXyCEkPJP/eNDoJhMrx0wVGNuOgWOR
mRA+445pxmSVrwoOhTH9jgfYLsCAJuYA+tHt8WJ/VG0pJYGg8/WH1XN6qkoSA+Em03zZIbKCqfws
VJyhKN2W9Ahif2qSF6ea99XX3vsTL83/72TviK0uREFexNzYPGoujSsntD3QZNcpAnw4awC5ZAAM
unemzu+OUYXHSmS/+4JhMfoNNLGOf02KHNESx/x9HI0ZiB4sCygBHHJGDyFXGm4hYIN70Y+/66nE
M1vXzUaI8EXF6MMj0NUjiozhJNVYDsK1kFBkmR66T0bCi3QooxQRnDentVlHVLVYTjr8OtJSpphP
9XL/x7R4vVe+s0cDfT3rnZQrVNmeK6QTchySlB8tokbcsLTUX7TgithNrPlPm1nhgvHsmzq0G4/Y
DMHhcOdJQzRoBshgV04KQtEqVgclgXji7SRtSgnIRgd44U6puZMFhK6HTHo9CT+SUzH9co/EOZKY
LWJ5iJIpi3ZWDXJhYXskN6KlxVSeW07g8EMeipffsMGIEH488mfTY+gXZPnqbNAeFcTj49rbdKCd
gfgQ81M6VxH35DyXlbsyEdWrsbS58E2jzl4uGJcqIOPVS0HdAzfZ3+ZBmyhy3E03ZFgz3cG11PyV
vO86y5cDDLjkboSQXrYpNWI8d3fjKXrw0BPJRw3IObDBg93sPAxrwpVRdKNH8qLtBoX94bAdfbWf
u4xfTjxuH+vCGZXoK01plHRyupPDwRoS/tjbPtsX6F8E4OpKq7gMaVajeNl/5qHOrRtZe8qHIrHl
JfKovUA72se4rlAEliHtP44tw/OqLdAowNDT5BlMzPXDNaANSOTKQNl/0BoRRDst9Yo5PFe9pUkh
gkppXEp2UmGzc51xE3rINSiMZrA/bQP3TrfDf3v+4TvfK5TuD+0EE8VT6pWv7s51zVMxwZ9yRBT5
L7Geh5Ki6LoTBwfq7QXGnDgkmk9QPFVhBjg6XidG/+hJPuHD2zC/sWn0HKX5dDLaE4Tkflf3jkcm
YjQxdHJtTe8osdgKllNGr9/eR0P6034qBzUkpmhCqOgk1dsoSWSe7zyTYlTvhvFVQFnr+ztAueAp
nkOSmMK81jCz+Ekd0FeOUxNLi/GttKwf21Y5IfsE9mplpkzjJAVXI+iY43P1y1XR+HIE42bNQ7zx
ELOHPDcDi+gTGXuIIHlFQufsrHXFeTA+ukrmDQ7GIXblCPruJhaXd2qPM9UrjvPeWvU2H+ZtM4gJ
qiv7EOy/w2VIpfWHZUY4vKLYtmPWgolbE0qK+oiS64w+A5/KwdGshgmm9ER5j/XWY2vNcFAulZvi
7qc1YYGZQm7m7uu/YAgfedQMX8lNhJO0daSMQsSRQgRtTYZy1gwVctrXed+9Q/m/RI0Tnk5yYiDI
taH0eI+rFrW/UiZBTVaGNWxgCY/wYudu6FfLe7Xlla53Y+9dbuRfpF8MG+FT31cONEvJB6cRzVIf
HvWiy6xcN3pJECeiOmfbkRggywI1NPuRcbeRdVWh+FsRjUjE6oEeipsjNalbTHIsuzvIOMkQFOIZ
prTYZIeMYMX80sh9/MM3alYa49hw4zXtu5BSm9XuIe8xE2sb89kxKfE5VJSk5C/PLrv06Muf1AuM
hQfnXAaSkNkum9p2UzNoWa0DGUwmv4Szaw5JpLkzDE6VJhQhNXSTWTyNS1T67KYeyGT6e6wORFap
RIjxJzM59B82Ld6ex7WRb0+xaFnu45UjNlImrQ4B8EIetentw0HuQLQYZ1mkvAACgpJ+EZGO54sp
xng+KGYmDfHHjkAVuPw9tQqNu2+AUzNcZQ1gohm3mnYiCAiNd0ZCPrCb4K4RttWiQjDl9Sfxjxld
vsCgQzbAwVKwl3POkKlfTCHLDsftAMvLz1tgL9svYftuMuf9yD69XZP8Y9K4P6J7c2v0nbGkH8K3
wPbc27Yv9xVhN1nlYecebKYZjD0vIpgLMWd5VLMQImcvNWXc4Zqb8l9uBWziRUYFUVwAQzbIRkkj
0MnNd8zf03idgvD2M18gpewAVi7su2Or2LM7+LDvOmjIfCnKcI/5aZ15f8j8rj47hP4dE3gOg8ui
JqDslL/2uDZ4BxOzbkQ60aXbrdTdNiYU3eeQ59JFmNymr62CklM39HmoU5iTALGYeJQxULOLPbzm
CiMWqCDNTbWa7TD2Le6RwFFgYPaKGi2jZnRcC4zyrvod9ESnNFjIU9AEjocnGWI2iVw0yTrmqK9K
EErVSiWj3DElbPLxxo1Xa4fITovQ29GbQRukHZxZe2PZ9SU+oJ+pv+O1U2d0GDLyz4AjaT6W+BKQ
kEj4chUJn7khAvH2b7ewaERskjwCSuQ7XReUnSPqYLUsBBhbALkPWQtKNZErayjPEbc5FCEKB/Fa
hftCraL37df/4IHA/fkY3G+R5r8uNcPKFXxmzRG1buPGxsbbYLSsBRaRqclVe2qMl6ZQS0Dx4hi7
LD+TBeaZZnlyFXTx0zJ7TE+PS4Mf5IvacHRDBrGH0tyoEEixvyMIyA1B0cZoM2Cul461On6Xn6B+
yZpoczOAKb8CT2yQhicf/PzcFyAzO4KfKfK2hKPXOx84hVaTTlGeyTS/5J8bGx+WKW+nH0S/C6Vi
ItbnXenvCyaybqPK9A26/LfA5RoNgN1zzyWo5g98SPmVOaeoW8nwFq2PkL51k2nXNpUcEopyeIKx
rSMjO9DkD8TTsSMlgAw/sq3D1liDgO9hhDiuD2KiFheDN75BAPVIIO6oKvsgB/aFnmiSVAAF9Lc0
nRGjRnxkhPe+wGvY5zQYfsbUao/hKZ4tT7Du/Nt/MLy/HRGf5d3KFaNFFPDpNDlXSlJs6MBdoJC/
eWUrw2SpzJx4ZcfNG30RL633Lz8engoDl7yA23b0by2i7531GfXx6UdbBH5eMVtmNc5E5xEd2tCF
2d1Gk8CABrsYLt6bVBTpUpLdrpbGVVwury2s1u2BOdQ1+uqKL5BmyEBUH+Bbv17mkM2arpSqEK57
2w2GPFvVKLrInzWk5ji6z3x5YmcgqSQPeqK9z9dXpA8h8UguteUNpvUAlnVRgr/YiVZ5PRDLhFg2
Ls35dtL7eiPbBSfGT20qr5Erxa2srR/Ep9b8WEL14YTyYuAEodPfL4dLE9312WLwRVOCjrzZ0gUw
rtA2iCUHrhw+05UbBecyxTaBBSneF1EX/J7buwodc/xJdNuTdBZzQ0P3zjD2EXJYCQqRV4avL10E
o6s7ZFFtFlz0zkEf8jxxC6Aoofm0D0VJ1Ctmfbtk5L6e9wWVUrcfV+VdzlF9TBa32r4HCALWO0Wd
DURErIDqF4vaQ91SzChbBZ1d1rb/CQ606hWWHt9HgGyUUTwX16IUgf6K3Wjh/fPS2teG495KovAO
HljxYuJSe5rPRwaqkrMhMKIQqki43C/gddbjg3zQzcmPZuQmvfvg81sE+USVlgu43vmz4dkj5ccg
NUjAFMb21T2JMJDQlsivUDp8hhGeh17/yej6/kzRNf97s1Xzg8spjhZa+NsXgIU+Mq2Jxqg9/ZCi
/LA2ruXLeegI5EGWYE3iPSnrv84pK8FqyVUqkt047oZ2MXpAZQYfJD2Dr0nzD4SXF5pwgv3ctHiq
F43RGqSax5IvLPJ2WwoEHtJ5R0oW3VVelKbkG1DBSt6qNOwQfq8GAwU9xP37N5dxHjy9P4qPyho3
ejtNaseYdFxkgTZ98EBQkWBRa3wjqi49xL8hhPAhfznteOKcKDgT0rwPy4GoRc67R/ZaZ44Hpfz+
yoogCzsq6a2HyqEmND8b7xOilmCuHiNyGxkj/bkDdrjCDodW4ukNfy/Thv8HOsYTJfP/uh4cRmV7
p44ibgRTCGd30j9IysVDIksJkPSit4bEgktLOFCsnqEUZmrlZmImN6jga6s5m3/kmrC1Av0iYvAa
SXeQrzpOPRIiyVXyeUcucN7tSs20riWYbOPDObl3DlXp7+gv6+I3zZ1XZDLLVmqL+N+vKcSZCVjH
NTRiilQQM+lbj0exNM8wonZiR/Kuwlu3GZX/fiq0gfxC7nXvTkJpQQY4OW07IovBpcSPtuUBxjjt
Jmv6VpXA1tdU7tSqNj3olLr7EgjvGjxVIjkjgl8DMzysSY7YJCsG+Jwtzq8tJunsAa+HOSij4oNP
0fMkZsVo6sieSFhlafZ2rYSb+PDjoG1BCY8XqL/oE723Xs2XOLFQREXIl8Hn+pl6BerpPccu5rMN
abaw7/56JZamLzNsYCJl22MV9vczImQ7W1SNWbaWt+I4Dz6faZmJKcRXkdDkkiiw2gSTiM5fXJ3I
/2ZG3l0vzNpTn8z9uUcB5JEszs3m5iPoLQc0GmvvrVgxW7kECDuwz8avP7VMZwk+h+tt5SmGbg3f
I8tlQ9HMt5/knLJsib3NpDzkmcUeuArG2ITyc+oV+X5vzusNZ4ny5rvbrXmFuNSCix/OhntRHXRd
95qyqJ31dFXlAkNQtSwta/2h8UUAd/iYCf6CrACpRADk18025MxOnUw4JIfncGeGaKtGu3W2wy56
fzuHiY/KWX42RkIpRyCoruwpUrBj0eQrH5yenrMthAXdQpNSN+WSbckIlx36PgqrKziyTfVzkVE+
mfL3uKA5OVkzOBnBCT7MPm1AENGVt+beaIZ88IOD2cj1zSVeLBtbJ4UkZNQ+stUwpKm+Hmk+fnvp
bfDbjAwuINfyddbyeo0SmqlxwTbLrJCZ5KC3A8FIkgR3qg02gRb/i+Thx3bQy9jxQ0PxtbsvUXue
dSB8iJN+mU5CwBcdO7HM5OnzAl7TTwF0lWKxAODiVxwWIx60ITccUKmM7GOKRk+t41YiKEC03tfa
q0et+G6P360YeHldCPv9fA/KceapiH04MTo2iO3TTQU3Bsgjc31XThx7Jd2+inWOA8Ta6KGIMDHL
hd1HoA4gN/WdyvhCXiTKZJDNXR38eND7ltB2i9g/NmtW/EpYtlp9f1cqMDCGJDIVic4r3WyDJ0Fn
x8b4vmIQQjGKRXHvyXkoON4fFxOZWf8Wmn6QM3Yon5znacuth0rsMvtuf2yUZl8FwfXHXOD2BEKM
cR0vs72ruC5Egp031DSGSFN9nnMOfHvXkE/oTCQPFR+t+XR5dhhlq513I/pOs7cE3mlDeJssAhA3
S49HALDOYTZJWl6Kj9RQ3J3RZXVxXY0gPP2o47fqpEpigkS4ykJTYw/xVpqpYEu2j8ELxKlOXC60
+SS+6iJ59s68D2rXI2bXIDy2yPC++B70zHn+OETFaPpsf9mq/6lKMCwUrUIWqMEHCvo+pEPPKWoJ
tucS/NHhdlzu5zrDXLtLlN+U/HJFb+rWeQqVFetrvHqbMs1oEX2st3X5oK7LVK5lWdtbPTz9Ukwy
kBXK1Be4Obulf2QkBxGJtSE3F+5nEpLUu1trJYP2sr2W0caV3uDwV/hUgdp519sNoVhQiB4Ufv02
YMGXLKfXGHb6SbnuyVcbIiAsTSPwx7K7VgY56YOuRphGVGmA1dRh/YUJPKGInKhnQ1XzDUFNISp6
WOpoLpBOewBlgUwWEspM0e7oQJG2qyiN04HWH3BTEShJ/T0Ah/Eq60Dt1pjp3W7XkodVizbqzEII
PhZu1yxOXsLhYQ/McLV1HkvT9R0ZMNgRzqMnB5CL908CDpWVyHTTvXWgfG9TeMdYC2i6+/8EM5fU
nX9kWxxm3BKfqY3WPzR/Rl/0x/RUzyOMRHK3WZnbl5YEod0XiFanAxeQanVTwosa/ViTb76Mfmkw
kRUHsUf8nWGMxQiTAr0GCoxOGr27qJdWXhTh9qbKuyHcHERf22XGU9ImBPpLZFs0mWpigdCh60Ue
1q/ut9FrAbohWBqHkmCFCysl8rQR8FoPBjculqMSp9QBBx6offqDVSgnwVqJ5svgc0+wXyPyjQEm
Fth9tEA2jfBihNyzuv5RSkb0WWmbjt3iEw2rNCwW5vTBzO19KAX8InMwVo+oZ8a3bmL+ue/alN2j
P6iWt9hFebTTKWgAuD83MnlnE/4G61MnMSB6zP4+siSE56fR9EN7qfFwTyibDXQh9J0LjxJ5bj6m
+QdhPhdakF0ijBtruoE5Ccf4XZj99CnaLPPS7t0bit0PHEM9eVBuTxnf4e5T902yokjykukOrl1g
8HuVklgVNij7fX2aUOWFIu1fHmCN6DdZtzrMkzxWPHh8zvZMHCKo7rV+3BVGAm50mA9UWz1q8guT
PuiaXqTR8V9/QZUdg/vNNir2z0lsZrDqO1V6lnQQ+oUztp7J20hlYsLSkSEE6lC3ZqxLJ02JiCNF
2JOY0Sj/l6i54vKuBXdCTOCMdFPBNHJLLGce4Ib4KqeUKCPDMYereAaY63dsICMI3PrKzLMm1lbF
5X09SDm6Sb9AB2ISxV6PJ2gupHV46jFSNvI44xpXbZdnR/sO1PyKHO3rcxyly2O7naMKnV9T/FR7
QAoqzbjN6d2SNdo50fWCfK2t+DzPlH4hme0Nvf3dOVDupm19FFbjcAczZZapOaHKlaHq02qpEfxu
jC1w+jUNBRxLbxloCHDRD4R7TqUsBAy3C7VILWp4sn+PFuv/H7wfoMyOkT8lPUkhbH4cr4q+thw6
JvseCimgtjzKwZ5fsF3u700Og1hG+VjKs8BhAV+z8kwnXgugdPhbN7d984/q8y5RulM5Q5zyKNk2
YGVyRx+S1pkDqTv6Yk0MRyYwWBapaLhRd05y/lsRHyx08N9JjEyS0CtQRvLoY+N8Rf5aW+uPmx5x
UFMxSzNSXO2Qqe9NGCeHFv9nDLXK/zaNh50vsg8cF5Np3Z/IsUJvUA3z8FsQV7CNyqTYsROQZ32+
jT1KUG5UR9wNTYwvGfOGUpVh7HxY3vGg0PwwRTm10OP592JaJv1A5iBds9hE37wFMoeYKrzKqJ70
r2LAuDstKKxSknRPZSKatCFyZMG2UwjWRhO/nppqLcBBlKlcs5EVIh9DaOcEwKR5Zsd4QBl/2zRI
3UnHsoiPEsuMrcA3CwIQwwyfgyEwArr5HhQ4t6zDr2oC5xKgKgYyiQQYOKRrSXoGydtu/CoWgH4o
qcaoXFyXOFq5qIjtjlNMLeUAJDDeHffl2hK4ilg/wDEXTBeDvfzK/ElGcrtQJ061t/yezMGgkfnI
c5rKBKpJ9lRdUMQr/Kt5TJd+Rmh2OYeXffY8Iw5q8jfxYHXMALIx7HLoSN2ZpxjQ4dhfUKat2sn1
eidO4X7VlZzL2c406o2TsOPz3Zolg8Rdrz5r41vPtVtHZEsS31zPO9hy1ItXOLjsu+0BlkKPkP8S
fvEZfHuMVfd13deZDAz2qN/UGFPiRCHtDrhIcbPa5a+79L4pi7fKbsbBY/r8Uo0vm2XX6y6pJuHh
PmvX4sml6XNwa/q++0Hnyy6hPQO7qXX1qCBE9JmvU2/0QwlPNAebalhd5XbCBXNFQNhrPgwlIAop
JGD5UfFslV6dSYljoQR5utO7NphzJxfPz5IHj9s5qozOo3SYLmlG8IdY/3ZwNnIq+aJOjXoyxltD
fa/BTI2KS8EVO8OchiaofAWhNXIjh0aquQqNk1wG1osrIlIfGrYrjDK2tiVtENLPtM5HvkIxUEjI
Kqh+ORuvfi0MN5LTMkGSAcvqztV0SVSyys1UpKg1pyobPck70LqiXolWJjny13FFbGtmA79L7y2P
ljBktdz98nJgaHK2ZLdrGB/2VBgWkoT1R+uMb2ujxiP7A3bS8bepWlm5r5RvDTERchIQH41IOvbK
F9KcSdOEnAzOUmSVtdtSZaJjNf/ol8KrAHMn6eU5fudyBsEqrY2yMo0cD5QtVLyucRGWYIfi0hpH
tbybuDfZQl2Ar68CKs9sDKzFORqcv0QBPRnlRo4yOnSrKfqCMTW7y3dd3f0r4JguCrcO+gk8m0Jl
q1bcubWs4/Fxshj7PSgnB2Z7sYig9WhwZNfScsvQj2O+7jIV6JwWKvO138TolqevS6mEI/s3qSQj
8nNngXzClyo6kKBSOCX7ReOnYcOhygPDL7yQQAtoKyndNmGjwBWrZwa9PXjWAAuRytF8UkYAqp8V
+gURlWzgnqHE6IBpGBluGHWG+hSprjBg7CVeSHeqRAwHJiykKeA9dw2e/0vCgR2FUOppfZRD7kAS
l2DoX38qyY7zkTmcP94Y/OFDzr1KoVld26xqwefRUSR71kP45obF61aHDiwqiQsMyRtuW0Ca/7+8
WLFnKUKcn/Snr6oo9imGkleRA4kq2gqvoF6IIxLA7jNnVwzSWNW78My/0mT2ABB2K2a1cXx60s6G
SGl+2UohxaCSxvtn2QLSvZeQ/kzwK67sM4qa4yrXmMzDvzOaHwR6DItuPKxtk3TZnP1Yycrmut9f
TQdK9g0tP72KJ4+IAubO2erRpDSoRqA+S8Lh1fdpbnoNmK+39YsfowE6DS8c+wxdkYet8FMZWUXs
FrHzcf/DwZok0CINwXYvYedDQvZDeRQbzc4p93z8sbsQtzXWwE0CTE3Qlr89s68FRRzffwkswNOH
VwSH5RUK7e+OLiCJrGJc0x3vwwwGKwm5fxV5yZ4eVTeY5skP8Y6+Cv9bxqsR29hLtR3Aumvine77
8WwY8SKAekZr4uS8VKQ0YHU99a41xzK9n5KHQpLfjAlkoTUIhG3VRY9vo5vcpOPVZ4U+f59Xa6Zc
8xHyKRV+Q7PSvi4XZjtn6cgtgx8J3PSYJDnutfABN5oWuFWzJWkph3fKesp6yvbLJcI11jlNeB35
PxVN6Wi5z3VV+DfdYsJgFDaMOUMc+LsyrgMOFOx9o6Gs5I1OOPggf5BKoiNUYoOU47UD++Vd3q9j
rLNdL1YVOgI1QgytDk0Ga67ySGmoM43dSnnjfnbZnSH/S0AOHoINy1tipZcpLgD+gN4xBQMz62bw
yMITJC8zTaJ3AUiVgcnw7lHmMfUlDK1iwE7APPpPriEn6NSYpD83dKbTz+1vUrtQciU4U0RUS1F/
X6W0lv6QUODZx2w+QbF9T2LuNtfgVq3fHsYwBm9ZIkXFuJTfLEC3pV9E2Gb+kzaaTGq2PanIJ1Md
eK4r+qPSsDmTnVcWR9znJkxMvsIGmIkk9qqWoPhMkvUeL7ZD3/w7hpNyXsWKZIyzTLpBk5MzPaNK
Q+ZJxg5ZPrJ0ZVJEoN5M1cBlMSRaNJv7b1LvkJGwst3mAK0wy9IPyDGrn6ejuStlba06Z9yk+zSS
OvOjdLuxvpPJU+DRl4KBjzMsZm/ty6IzYj4Tc3LUpUYdiPiAmycrpq26bsw07XRcxRoZV/KiPyfk
0NtEmxhjv+9fpEeRgCtiiZmJpu26ACLRbFS3yNd9jTtnhwzV9n6qWgjhJISIsOqLzlg0ZigJz5yV
Urg7gCpPGHsrGW97E9FsRj5axyrd0RdaeGW8Iaa1AyhGwXFvPZ1HZxT6cae6eLsJ0w+RBdvH8kIA
mFtJfU0OSwujdsq10lEMHvWhKYJtZ3K4JbpoH7L4r7kTXFGtUH+Cn11CnzPWb1O8Yjjvcbchwz2M
E78v+JsC/NIfmEcJ8zLjdmW0bwo9YVpUwErLpnasI07ImBRKDIqKWmL5uLZfP6ETTtCd6LFYOafa
+QlZRcIpl6nNxnK9ys/nZQ+GxhNaTANHld/kf7m+mMEOjEF9Irbxbdv/J5A8yeU0l9IGWli9YGLf
1Oal+u4tSvNvFHK3PUIn2gAIoXLKJ6FLaZRuJEc1T4TEv2V4Q6okKRYVojSUFO1bRkdYhs0MrpmC
xaeDFpvhzbNVEIWm4KNulSu3JJcLKBrJEmAEyAgJXysElATCCxVgXFEvgM5LlOQ+cvr8tuuA2sAE
3PaanHr5L68Kuxeq2azB7v/LiF9iRQr5hNU/5br77H+H6xs/fkuDOqCXGlhA9/lft9Dv/DYZCPJ+
lo3Anme5cZND/0odBswTf/yQ78c6kE5hCdYrwDTQ8NbJDQux0cu/RzQeKa12UtaWOIy2jf9lrRiN
H0bHImh5O7vWkVWTfQxO7YguauosHlRB2QWEOwiMi521lu+4+dggAlKq4X7k7DL/8cbBvX4g18pK
qxepeSj1unG3NC9TsHZ7ILZeUn4Ew2VwsnhMCLMEXfRRMpXVanPw6lRmYVbPYTdvGnJB1vAdQhBb
uiHD8tsA5sbgDxPCYbryWE4gP3++qMmoQNm14kDXdzqe++ZRsrKugh3BU0wXUbhRX9PN9/U+UNRN
QFOtVjkCGgkNjtQQmPRpnUf6Zm/k4woX79kvVjmbunnMXkWxs+nrOSrpTvnPdRartPDYF2BZMigU
5Saox78Ed4H/sW1Ett387Y7zygjPWL+9GJo/AnDKlxpRqC6TdXeuCg7Ldi0qw0LKlx9Ow3dWfZw+
uGJbJupqaa2LzhNMPhQPyo0Hw0WT/1BkVmhOjdbfUNaAoMrNdCfbFZc/7b7kK65VZPjUeN5A2J9E
oASYp9FLW0fQ9udkNCraeo2W6o6R//m/NWbNvx8PQWnVPnyOq98FhE9n+2LrM5uAgUAkJPPT/DKj
8HmGz6VluYGH9TaQ61sBee10pROKMquxbLr3Dw8PGP8OFkY6X/PUXNf5VWRdPz0B7kvjWjxPMSHy
JG+Xf099Am7c8sCu5zmT6tMLqiUniijzOOuOSTscEpL97eLNtcpADr7dH6iXOVyYhPvT0Mb16UW6
bIyswu4kSpKVhqTjw06+FaJV5BnNujYd08d2hH3IiKHIHXGe2ZjXRw/LKObgFJIZvnrvvN009xqQ
0L5FYOIfDHoLkTJD8yOptn/FHljWFIybMbAx/vNC/Aw3lUc9X1xK0djS5rozFUWeLREaDYTLr6yl
S+NoX/5bp/46FSTohIe1FSK8ZMa2Am0Oa7VBq4vHnFIhQZ3BQg9emN5GoagE6q51eaCzEdUunS5N
6UF8kfupiQw2G1JQ1aVTXy5np2LyLXB23QrOQ87JcVcnoOznlE67lG7ZAd/0TzUOM67gYCMwg0DI
L2XnXume8LT0nxMwwXwuMCam1HCDfX+JAp71iXt3KRluKnoTqpp+FTpAcx0aJ02A4ywWiTJEojp1
r5NQ0pfwLXiZRuyHvbuibKYF/9knzDrMAJ+myYKF40gk36uyZol/9uaf6f/9OyfFL3d8hDMtp0IX
V6X4HOPRjfZqnaU1M3WjSF6T3NAVu0vbasY/a2MLSc/y9b5MHIV/lyYTS5svof8LMx/SuSw1y/3o
zL1QmcZRuU5lA/WjRqMwSwSP13LxmR+eqznyDlxv7/nGNqviokqiBPaTAE4Ov6Q6u2E84XrYFQaP
hspEro63WkCXPIrgdP4a3GT7Wvq6X5G47UsxmEwCOWua6X9oqCTDAp6RN3xt6iTBb03kZjl97ZJk
kTQsKruyt7Oh47a41NEpxQXt5amZxphJQF2Gju4XEFmkRcXBoE4XAfqhTaHGhF6/QZY/tB4vqVur
gRVaBxqaT/fqzB4nnv8UBLPAXcv0ZESvlmskqKvNBNzdslDclWYQoC2CwGgXfTR9t17x3odPU/bX
9wK2elY1XgBCEtvQnKwwIAeTu2qfCBegQH5muJZ30qsfjVbpq0IvwvfkzV5BiawiCrUAjKD7ag+l
K7480GqoMn6C5kDelGhpEmAsEYohumbnRpBGZXgEYzRqq4L7PFLwX6PxHDI4L6oVNQJRekHmbb3S
jsTCa6C/h9gLPPt+bijulHw57cocc/bF6EKT2E4FvDYTBHbFMgL5J+gvUTx5ca12Aock+cSjrKWd
4w0ApZMilTq9yXd4K6HyNmoUE31QPm8QTIADnRX4BReRVypNwRU65u/3lHHFxwJJ80iFznu+R0Qx
x6ypTCRdj0+XaT2wQ3Ux40fWfHuG0W4DqQaHBlkGd9jyiFE77HRZdzba4IC87r68JCfGr9ixCFMV
6wsLT2q9FhFnS7LQwDCKpxr+b5R7TN3ED5EJ9HH8hu4SYEp6I7sDVeIDX9uexjFVGe4hVz0qwvQL
ygUwAsSNFe7aR9SBOT2qBGDol+GTVU7eP4I9uJGRD0dEidS+PdQt/zEvzr68o/S0PzP+TTKBd3fr
jDdcNGZl2UvIcs18tPFtJBDVoq8eUCoqJTf8VzHj2cNoZCMM63LgTQK3mESY3cTDYgIAsely3h2C
CRh2KeVQ60a07BSYEla0HrTXEJ9kl8Tox+YOwUIAQyzgzexwYwH0kAVlYLNwbWmyaLbC6jji8r1m
rc0+FgolOHAHInohcOJcN7GLtubRC8WmNtQLRxkAB5okAXHwuLv+slPp3pKeNKcohZeeF8WhI5gt
vDu3/vVGeKHwT6B46iZnteE1uWGbMB9+LBBTFq3m4YRvFnfxhPfCVe28UALaXXkiQlQJdSQejKdz
mi1Fhg99R9itaonvOO9i7K6brA+WTkwCiD92iJOh+Arva8TBtkJfP99BXhw1925JyCxOw6cTLkmu
BwIItHMnRIDrUY/vi5ZPIovmPcC1o/OQZyX5/2UAJC5EEFqxavPeuMmypuUQ5XSDw2tw1nDi3oJg
XCnu3mJg9oV5UOazCYnyzYC+zDGvb/qhScYBd3cs33ovWBUxxfgvrtrJ/Ewzy4j6OVFlPBLLJlXw
+Q9NXuL9XkMjTqHOi3L5KfABNlxHgTchsF4oSaloj5k9gmo9sts3Jnwd0AYMrCqJuptBDS2fTNhL
A2tsfT3Qh6J5cDKKYKxcPU8lmTOtu4haB58IV4xd1AvtBS+YOXEwcqVP/TWfj38PBD2B8eMAoAmk
wjp2LtacLNiIfFIjHfJJ50+buFbkdMYntgDdw4z3Dy3x//XCtEFYJB5SwPe8d+3HQh6C4nncj3NS
YD7GdkoVddKltdJ7ScGQ1Sbi87IeusUkdFtOAuvhvqKkJrX8YTtNvSFY3yj2lAITWd/pF/Vbjwz/
wUW5xdN0Dye/s4TlaiVKWTi0Suk+u2EogrEAbNSibMzbzbt3MvIW3xji8WHd3HoEFivUIodXAZMQ
upQUOwXdfdmjvf3xdetC5WqNEaqlLYw6w04UBLP6dL4SeH+Td/eCM+UqKYZpjKbFwrD9KhvSK0aX
RwavlL/kufTk4mzrfnWLRayePYTAwg69scgbqY9x4n+kTw/xv0nzSKmDDeY4VBQvhZ5GSLhWNm3P
mUxHvaznI1YtG0vhfSU8/C2GODRASOVY2RxgUMzKQ/SGvDuAf7meyfq/5HLz7ZrzWmDH0Y4TdDlA
0FenPnGLxtlkYVSJ/SB9IgJJRNReUAjsJCzsTPpdkzjrOT4iw+L+pvmmoYqf9OnvUDM9i10qPtof
ro8/kFYZuGXvItP9lmurB3/h5X5p1K3z0skTBNUIsWqHMOZfzFnCsSZk1TPE/6mTtRz2IZ8EnqIy
6cLsMrDGRF92zu12rcAsOPnkO0ASB0399Xwfxw/gIXtb6ZHqMavGNDsTXgRykb4eAhyqaGhes68q
MxdmXBB+EH0tiEG+M2KDmgZB3yAbkGAQpAzimo033P3+8tP/ygP/jyoaf8ZK+5Ao18XD8eSExrQy
0GkFDH94U4Cg0FRq+4dWsiouyDWt9VR5pag354djCDeLVDg1i8ydIxkaMC0kMcynqyyfCAePeXLW
tlmNj6RIVLIfsQZGX7vu54SHnYfZSeJp0hgBu5GFd/BE377Uzp3WK8GCkIZ76OUC2OLdS9uKWOSd
eS3MInBwwY+Db6ttc3wz9X25bOnkPW1db996F2zgdM+MOAVApeqntnpBcJA2OueOFRnKU1zLGCn1
o2vXvjmeMtQKhgYCQuTafajsSOjwtKj5F9oyZXg8pAf2SoEV3MCdXTGqqVXgvEyam7jsxqPpMKi0
trQvPSzq9EIemk7rPGfZH+jOmq6VYSW8685F5rRQzVf352OfFOfXRY0Y7pEicZCR2yyDSDZ+kIU4
I5MvJRC4HMsCgDzx9ghS+/KRzeEskdz/AmqBSdgNIbLr/gddaSqOUbuCP4rqwV2uXUti9rbQb/b/
se/qqSYI/VKq0kA2CbqmHwbk2IfoiEuRhw9ifJw3J9vVyvkMiZlYFTCs4O3sjE3KakZ1Hg09RIZE
LYUrd8RjJjqyiTOyg9qN66Cl2ItUjjFNjSnjQDAF0MzI3KJ7ujBnYHSyLZNv4rOVkhAj2CCPxRY7
1syeyXHJ27eiPMxfqlAUnDJpGBmvURdqoo3lpVPj42TZtrI81/6g23BvS6Ay+ri3qqrxLeQDJjBk
UXlsLzGQmD+SvUNZ2qx/KYDgEsmkWXyHwVqI0OS3clWSWGSpzs+FhkaA1H1b5ZpHt6AUPV1rZKnf
puPAKf4WkXonTMRSSBNNrnWSSxJZHxLMA/APUXZAXFJtRvO6Q96vGBXOQ9K6p10f9pygJ0SxWIoq
NofGYCbmNKQZCLkH9pl902pfyTXrouHgaxDbkTT1zcCcXh4uxMpJC0wnUyUKvGQ89CGp+6UgqLpJ
fm5hNRMTejIH1AeTLqJftMIs3+xcjn/juhjqWVNNoLENwcgzDKTJAK2xAXVRwzV6lle/9dDjGd3p
3MV7Z+f3C7rbDo6qsT/LPDHSiCbtTfEI7/jaYGyx7ibcc68+uLRr3JRhnfG7Po/NCuuvDUR2YJY9
gA7kHDNOF9XMJyC94YJHWJVpq3kEWYKQxmNwAt+I0YSRs7G/8D92BWUetPAzQaOJeWa52C5ljvmn
meSx2jv+fBGTgur7Wjt6FLtliDz3aOn+za1CBjYOaGDI0xwkgT37Rn7AZQ99nipWr0IiA3YED63E
B+7JL6TezXQCMGIC0xOIR3ngW6cFPElwV+LN1VPrS+kqGZSyERM2qeSvpqqfijN1wayADLgvnuir
tfYwv1J9icFQcKXRSZgA8YJtT9o/3QIT0Us8y4Bjpd55e8y/k1PQ9pFXr7q0XvPGhd7jtp03vzJn
MXX79PUlkhFiIEad44RVhaU2dNeXA8K9tWCvJUHnbIQE34KStoVuREseJyWk5X13XaiAAvYdz1pD
dKERyKN164wXZh4LsZHvev0sEO02o4XRjYM1UlHVk9ya9zv1WykAqwUbNVUDSeHMNfM98Xe4NxY/
7RklLfDsJ06pqWg1ffuujspZiQyD5QlTpOIi7XIrwflhtpdhZP33kboC1VxQURccm4FC/O+yp9E3
6bw/6Venw7LI5WLXfjWadmoDKl1A+px444M8eW8rA82TJyyIY2/zHrnCw9LBsCmN4MGZ5edEGpXD
QSwBk/JKrgWAGCY5zpLdpgRqRT6vvbR0L2+QA0HnFCtue/YW85awoG2mStHWTYTPVRM3/x/qNbfF
UQd/T5ygAGADtheBPxuHvAO9QtOOw2L7E0zM08h4u/OmPfG+e7vZqpzlDmJBXboo30PRCOFrL3JV
IAOXe8G1iA2Qrvn2Z7iGoYGbT5YiK505aJ8pZkXNx/id+H+Z6gbtuKUVPYgW5OAjSdy+TVFhb8Sh
sBkgSxRBbuwpH2Nck7ozolB9E498K/j3PVx2TDqQN1+yQ61TUXJQty5oJlZAhE2To3gYGBMlNPtW
T3LuwC7cSDLiKxifr/uMyFzg6OOAiDsnlQgWJMJyli8EZSTYg6p2k07eeOAh0k3D7Ei3wYxb57Ic
SdKil9IYjWIBDrIyCY4NLyCvA31DFo4+VCq6RVlTEDaUXeLdWQ1Bpbys7Bqg4uiaubEHmBZXCBN2
hJ2yPvL0z+F7hhvWqEQhEBk9mf7KVLGFvf7ZMwosYZiggeMv2Cd1yAjoLtT28v1ZOjh5yTxcFPXa
GXE0QruC7+T5FZGdgYU5tSVoNdVeon89tpilZPI24WvudwtwWHQzdDUoCE0tsVaaAp5GCTD+cbMM
wOaYJnKSJMnAQsuRbn4pM7h9RJOpL5ckqXjklfUynb7m4XlRb3RMOCWalysE0Js2Ij4FILwMPIa2
ZyiTyE38jb2IOTFfLaGfshzTSpbpZVHrIsW9kmKUyiF4hdV80ZuMtfnkOgkg23rKddA7VYam5EK8
i+zjizWDVLHBjdz3zq09lmBYsTRggF/InX1xvL6+u55S8C9ADjyMmLvYgt/sZI/IIJKDG2oltTbG
M85GKBfUHquP/UPIj4HVVol3WVXyD5kE4sA3O6Z/iDIu1kdK2fRAezUyT+cA78d9FIjWyR2CZPhp
eKelXLGSZy3+DZ2kQRiwn5DkE4Y3O94C5n8OGZ0q7dqCc7U1Adp1J7FAAnoZaKAb9qwceoxVB1/7
Ay/dMeOP5DSp60qIZjsZylgW2vMhlu1KYQexoPSFcWHYvz6CHv0aGIP1h8WOoZBnYHqVReohgmmc
QL6HnffblSlQ+b+Eh7Gz1kvDBpTH3yiLLxXlM6WN+qOlIavgMtfnu2TK6QElqTH7zJoV03ZJxQj7
fAHuEIimPmT56vB5dDrXr1Hxeei1pt+irUfAba23tmDKJPXefPJ2rkcHqVl4YBuhL/y1jwj0DJXd
XKLJPpQNZBDLme2EdWq2etfwMjdjVR71u/96uS1NLuzMO/PwDcPWxX41dJHbEOfuHStv1Ld2fLFY
q1IOta5V1rd1DpkE0PadRCCgfOWTxiUzTQWxNIeSuadIhET4WUAUT4xPAtNdNmcLMkM33PlnRFHU
nOw22jpmAbaUJFgL7q6XSX00FbyExv0LMYMOb1QispxOD5wf/qYM6uRzT6f7w17Bj+Mn7uQNxcAY
hjHlpYht73A+hpnEJvB8w9SSR/evAgfD+ZJ1ahg5WlKgtbp/3Lpne03r+GtukMnI/ca4QzvTHbFV
Tx402rUxn7nSuoG/fnkHcMqPiBPnMhMpV4Xc+z2AaQ11HPsykb3rsz7Z5TdDl7W5c/WH3RB7GLze
UdU/OJzeWzN/Wmpd2T+zb1Wqzt89ni/byFS/4wUvis40htIYEH6SuwuH04XrWqTfeGHPSp+sKygF
dLzS81OVnVRzL6+VTC23UFYBy1rNuvCc/7KKN9kN4rAQ2+CjvFpF2DmFY0RT3VkUZ3aebPhvsgKr
sZPbXtE1g1ktLpaWgTafr5oo8hx7VgZWtTgBts/p103R8hdPr1cFPiK7xn0oCKIwG8QGa/kCm5qS
Enl3UwfyLvZRpbwohA3I3lWfjyXE5Exuv/R2MePKUixLuDjH1ke2BR36AGj1zd1t6LTi/hQaKfDP
jJKAKBTAIKE4cNdbs0HMGeNwi8Al3jQYL/vYQgC7K3crtLsuGfGhwJD+0sXYLGinly7TcBYSJ9bs
DfxDmIdfbD1KZiz1xjCOkKSYZ/oLR+HtuaQNJCMwBzs/C7p1HClh9e/E4Nu/BJKmEr5sJGw+X1jx
wIxr+mTKo7dePqm9Bsjjiz7zX/ILEj/u7GCpgMOsC+vravFv2tJ/wClSD/jMR4yAB58nwenHeDcM
bsuTDGBGX2dat8dhMXpQPh+4SL+LR4vYsp1xkY7P/69MnXYoeWV+l1eSrD7tPe6juLvgtZnH2r61
fIEa3f28Qd7NtZlD9zNDaRtgv7LA10naJ6MpGRQmEePElp8iRbnD9mljf+Wf2mGY8oie3TSrNXRz
SIYhB1hcgcCWQACJfvBzi4wopLjsiCr5R7uioN+QiDWAtw8ANFxYZp7og0WEGdWD8+J5rIudkg+S
MxZnFzjAt+xH35Hn3oZtFFA81vvMoaXY25YvCrNX33reaVs4TTfKffkLOU6EVvRIDfLlZvBu551z
RSh5sHS2eH01/fnPE8qIIYocCt8Flq66aEwg8kO7O0BCtCvQdETN7l9R2QWTa0x9EhgkyKOjL5KF
I/ykkR80O/Z5ty3/l8Mj2BfLAPiQSAdVt377EpnPfN3IFjMKU83SSWXCVRjtMwtzQ10UmXxOelrH
Y5NoX0Iom9C4LPTw3HeXjJFSgtUOr25XQbizuIu1GPtU4qU2vBao/mkzWq0y/LoRsXBUafN1NqpF
/GnFgz/rmi+EBc5R5NGr4N98htx0g2r+yfHQ8GihrP4eAZYK0KNP8V+ri1pA+ujssTfFgyYuaEyN
KbgFCrpZCj4Ti6R+VE4eDh4EDfC94mrPOQkBPH5qpkbWbp2aHhpecs+mDZsq1ZPVuulhIHeNI1zV
JyS9iGHoWlhgqAxFOuT4R5micW8fnOFQvHg5lLwjn2rIjxrj8cYPWegAp5A8uWMWyR3nZMff1I4M
kS8Rjrcx9XPdB+9BF9CGLVleWyn7KJ8JEoNuCSyUKe2dUeP4/1QnqP4sHdo+/HeA8OA1lWSox+Pi
PCny5Lbm2CyGp9NdAm9ufMYm77xdADM264EjK4k8wcF1wAhmDtC/jgubjTqQFuz/SHBoPssXFMDH
tduM/hrHZNZe4ptSvl1+YOhHBNeubStINa3W7Iqnwk5+r7X3Jzr9lJnPA3pMVKmRV+h/EVt6gZ1A
TTr0+ab4zb22ZVhdN25XPjtnmi0qa7rnIE8Z0OcN6iJm0q9S2sZkpalIlPL3iJUVPXOsiAz/L9aj
Q6L61vPANyueZ+x8F/hCNn6VEzO4Czqn074UfJmpSwKd+CQaHqzHkH5FDCV3ZSVCHluConEUAIZ+
zxSON/0F8YkkMyfwba569oQgoZ9I48Mn1pGi8KWp2cPi3whVgnKTS7m7Bh3HtA9Z920YJas0RgDB
WmHjO5F7EUhujw8SZlwNviFJrbGsOgwBo6y+KAJm723DTJlcXv0HVNagqFYifmv63F/tyi0vf989
Vj1c1hydbA3cfKeXJXlNDFEkCvzpOuiCjwZ2rUo+hY2784LF9jiQQpRYiVEnBY4U2sYtCmUgoBRH
MXZcP9hlLqjdYXShjLfnZhvZcOfYlElnlNmYuhVcE8PnFm0cyGeBSd3zlD/aaErSs4ohGJz1HOHV
pZTqAz4w0dtIM+CUItW/yitEtQOX3HMmklsxlHIZhb1hvoLsgqNwnGAU5GluX5j7SoVXsmHRBv3c
m7Wui5PqJ+t2BMluw972ANQTLPY361gZuR+xHDc+75rWjRUPpgMQ6d1GQfi0oPVYHNaiueO/vnnf
syFImiX8qgWVA6CFDmvVaG029Pi7P2VU4ZlYv6tD1LUQellSpzRY5pwOMp84Qpw/LJcuB91kAYar
lhHY6Sr1mCW5Ia/9KWDZz5rYp58JHDNaKaTSi1186AgBX+46AAVNojLiwQjKGUEt41uR/y4CTOv/
k8v/EabVBt9IowYXJ/M2x123f3vrJ5OM7MVAQ4e4/RlhAib5SpgjOO4kfBESgI6fJm/mKLMBNNgh
LIsz3+sBOYo1XjrJb/mdVDBHnQjBzxTOCyL0SHml0EFGuWr2wbDURoiXIY1zh3N2qJX+HlsRGv4k
A1F8cft5GjLi3H808BIjV62TSVidKzuvsYaBU4pGjhDxcifIOQYYLbNRtsN3C4D3WLKi5ec7x6bJ
Kaf3QJcOqLsgSzHkwp2fQApptYsTLuBbW6ABqUu1+R1k0qF89A5fkcTnufofRNEUW3b4m+gN25qQ
FBR1nlxVETKgGvCwhL69VFc7umpNhoFqdAYEdA6LBsH0yz/bKVjek06W3uVT744xalGxCpVR2ywx
IqiEdgioSlUAigRiUt5B3hp9MVvR/G3EWXFPaZI99ba8Tu7F5btBmV9JB3wV2d3OY2VqiL0ZTlFm
iUdPQAO3HKFl8wL8P2lyJXgVUUiROYTtKvA/AYtXlj0apMw2ZK+zzRTyVtbG5TgciTjEgnQl9rnL
ItXDNgaIiMTLuwYP2BqIhzA78JoI6PitrZtkIoYTRNDCOFuTl02sOmKnJlKPEMyPKjIXi7sz+yCC
eHu+UAX1aai3cgt9TJDnlAP8JRQHT6YBFL3RZD+ljqnXYwi+MtX/KjUJ4CpXq9swPOhQz+dirxRE
X9AUzWaEL9LlmkdnOmVJY4goDIMNC04P2jrcerE2VvI0mMHBY91ZZF8BiblMMRMapiWK9HHjWyKp
kDVxFhUsuQmUR33gn/o1/MKR9avjk3brwgklbNk51y/Y54XMQUP0vvhBtPi1te4uhZXOSmDhNX/x
6MncWLmhyhpnPIwOVFOM06hMADQx04Pr8MwIOo18qizxk2Ui5NgW5FtXdZp3Ok6hx7ez3M6MOzxb
zaTD6WNTcR0d3IECwGN+1Vldy7ALI1vdiHb3kRAzVvkWER8jzB3WrOMsLTMgYFjK3KRnWBlFe6bH
DE0eELN/pz3Ra7ciN4746HsQCGZMuEO+85pURfQoOcbXNR3+gE+VBiQlkxVTRCUOFRbjBaNC8Wl6
hx9/T1qpamhVnxw6xeC2v/bzj97RlAFmq9LBgwrpyiL3HKnIhc4QE0dTSeLnvyMbi3Q+aMGV6DTR
9Wz6ocYMOpw+2cl8jzb7Fcv7uWZ7VOQZi1TzmVR2z1cwYKREU0BAx0vnkFug43IRVdZBvHkha1ED
OkTqZqbIO+voFUsy+ot24kMC/oYZcB713G1/D6155W90NxjJ6GngNVxCz1cnVqoO5NzWr+nuoTPT
t3NL5iiwletHArtvh8wt18BGZM7fE6NDJy3AHjsbPIaaCCasJ58meY/IeXyFCLSgNTZIr5yXjBsJ
mnv1PKq6w7mvPYERfnKdyqCtxRQIgbtpw1y9gi3LTqwoOcBnjWtrVJvnN8ap74dt705Hrmg8/uOk
al8guSG63IB9febLKrzyVXAOxTBNO22blN27ZX07LHe3U9Mfmu3r8//8AXJ6okLp56DJfwzLOr4i
S70+YY1S9dsJuJ3d5GdJvQqiE9+eJj5C2Y/WTHkrrku0L8RZDyS+aKVcxEy/7nFVlpI42sMcPRua
9x/13bJi7LC6OJA++2KbTCNunBWnyihgQy3ReWhVmqe0UWZ55MuheBbNNqlYKae2Pe8X0hNPEb/e
I7gbNIb4bM7rp5ujetYNle4e9UHmiS7FKoRhzwpN1QeL+EC+cd6XUvvp3Y4hlzzJHr7ryxxEJ8uA
rv67T86/DBpcPaMC6kjvx29Y7Mar8JHYw43s+TP5ExN/Fxl25XzAKGCLxok/tTNLm8jEIp1BceCO
tnP+JcZ/TXh0gTfG/W546pVjwHPcwQR29VVWRo5MXxVeqHXi7l9GXl/1T1l9B0SNvQhTmhrZCQO0
EM6NJst8mLJvBvoUtCT5UxKoExRL0w1zUf46nLjuJwBCc5xB2hvoXr9oos7zGM7d2Ui2F4Zu8PSQ
+C9S+yhC5TT7noV6N5QCwsB/YB1VLiwawZHz9XdOTF+50Hzoy0U7LD8K7WAmKLPczqoMSxU2/KpG
sacklQxB9ZIDKySFEfbZ7NZ6pP9JmnWFbOY35pm54ZtolcpLk4PSioIzUw0aV7gHl+fPDlHnCszx
/faMu/pqxhhqCpPV+t/nl9UzYMlTqVnUwY43xr4tNG3mfPADbv1+z89ucc5vkNRz+AQHpJruQob3
P8INA7FHUy10x+HHls0zYvMb5bc8VfbquOMAFVl9eMZ3yXX/J3EJjSOuSugNJRJzeexs5yReAs5S
3WFClbVGVynHcKK5ptpD6oJC1J87a4ge9PyL4dViQolJXA+yiVatHTxgCXyY6vjXTBdyEfOmneZ+
5hnxo9gkYjTb+oILDaywt5zLh50dKJ1x3imDLlr72AII5LihYtU09am0uF3I0xaJAx4B/u+BH4Zy
mhWEYcjb0XW07jaUDbiyFFjhvCe0wmIi0R+C8x9ShH1twrWoVRUHRoTw3WxbY5WIaFO65Tom943O
K5oNxPIa0+Bksn4HEGVsXvUrHUMJJJikON86+Dp7fbOZlysnzPmNv8h/UA6QnI5m871Ic392rHsS
JXfeI+YeiJztZXk/bXOIMiaWY5VCm6ISQWEB1jvFOItilCT3AsOexIxhFLmdIdFWdSL6el60ad9E
F9EZuCNX2sl8JAAsdCnqYrdIW0IZrTR89bgehd9OzTzThA1PtSXU8CuWbcdCebHpcSkcaLvtbPEw
CrTPBGRFUdauawMwHHte5wGIgaujYMQtHqwfFcgIRFvW3KO4etdY3ZxAfY9wNfBKL5zO+MrP5Ot/
ugmguWftO3OKAeBpEI8OmgDmyZDd+utYFDejkHXyiyJWjHrX4CDxsKuOGzTxIvh3N9fU6Zuvv/zq
PwFrH86RoIEXXxlcwGQy+6fUbE1FCPuP2ZWs1xLkFXqsZwYf4E4dKqL7iJ+DKCnP9mHKMDPz1naz
Ua5Wo34OO23ynG+knEn944izQ6Vi1aM5+PwfiISs6sgSSw6ukT86QpyXe6hqo5UR+1EuJUybufnZ
JiLabvg5g7r/LT7obCjfFOEPB9PnHnKQ9Bdae8GL3Wuccj8O31vtTMuM/gv3uv3gsuKPkJ3PBkog
NK9Yzltml2oi5piRGOC9V4V/qn3J6QLm3qHG0cfKCRyDeXETYh0pLYQLtd37aVI1nn47INbL+dah
ocgTiRo/WfcHyyUNP+93TTQPMVWEKVX/+GtHQjSjaCF3xNr4JZZ4M2rEwqlJMh9OLB6oYGIRvFSb
xZO61nhZNhhiRlU9487+4yiUPUqxVS+Zh/ojArLPoBMw2VtZA7oEgkLOXWvFBfFN8hFlyXzzCAnO
4C8wv0Js0GyQSqjdIvS0g2PD0a2m1tzhtLWgMzSgqBzlxLLGs7rQUYlEfkaQdaO284psPrb/dOp9
+D1zZ1iNeDlpd5ggWXFXfUd7iIecwrzvFXpJ7PtC9o5+58OoPkT7BqI6qHj8jTSdtIdimxd9SyH6
KHmZTbvFNNjrv0V7ZvqCR7GrcrCo9IsCh0eo45YVcXIz3seJFgSOWyTqNXVYOEvuYJ6DNg5+RfN+
eabXObtlGzX6K/QLgp1tv70gjgiXnXxxAIKe7sgMVLpdx4CKTLcqzYhH0OOq4U0wLEMi+WslBDBs
AhVuDTC/lo4yJd6UYqZDH8q22ZcI5SqdjllxoPG3h5JJeEfRiFYOOsQ/+upWKKCPPgBZBgRsrsS+
a+AX5t9F1ip4yCK1VoCsVMHUAaQx9PIwafRhn/mBJreaVfnfOu43udJagNg4KpXonCi9/emzj286
n2ChkZwqupgKkNaWwMPMfAE4hzkwq2Hi88WD3+36Vycqd96Gnb4SWgjfVfKQGVYIDqy0Y7A5EEpJ
/0ecs2QWwICM53PrI1Sf5BwuR12HQpcR74Gl+0tbmOE5AyIC9DeeJwUdQ+q5IwS180lxkfWcJ+EK
R3gBM44aK5/rk2NK3icamOULQyy7gxYHmAQOK30fObZ8xu29xD3YTa/rOOxMMMHzpYBhvxh/zJfh
pOQ4urZnvat8fxXUlrFJ6Dtc5OpiJA9M3EcCD2m2zFWXxqAhzEUtF4e8FUZbcQWujTYct+HhBUiZ
NIZiSwpRBmcTpXq//AK6ldQ5IWxyQWlCKkY05+jLMFMOsjDDARPdO7G/dodTEtMpfWL9uFc+urcn
GkR3AXtv8ojACN830hc0ITUC7Etxr2HgKWzmWB08PO63AxShUykhG26G2Xay9IqKGztw02tQjb1n
QF0/EOMEbEKHNWqo+sr9l8jB2HaQUoVVlCAT2KkcbEkUbBNd4iUHYxl9zTj6UsQustSz1yUUn34f
FRWLkm2/CG81gth7BMALHGFhG3IIA89+mnAaPR6me2EPHEwOwsEFpt04/Lgrum6PjBdAKD4nWxm8
OcfWR6YV8ETP/Y+fotmoTnABXYGvQNbT88zLxFd6iT4q11nyBQuCKoiGGcsHATcyd1Q6J++O6vQa
FOqvOLjjzeyzvj5W+8cE6xFkROuJ9+hgyY/9wUNfmL3WnjfR6Teiz9AdN5kGSOq8YVVc+6m2Clxk
LrbFSTMAYD3Auez56T8liJENpkXxW8cyqyG+rNB60dcxNNr0qfI4mwfHVpbeZuDj0n2j2JE7MXvT
kk9JZadbVsQmtlUzv0lJaS7KRqnhcB9Mq8VQLy2dNXcKhzIArHoFPyFNdmD9SY+Yi9sSkPiIHQGm
EAgZdRAttkX9YWC6VzASmFJnd58StrEuLx2w6EwrNsRCvUfA5uHLK/837KCeMostm4nQPRmQB1wi
3S/pykGCLaYG5JhqqxFHcKUwOaL7cKHKITrAxOzwbjEF+TcokgXrvtbAMrWU/RniEXde99IHNGPi
zvGcYaRkCfGmuRfZBI6aSqL1mvp8/ADhn1DEHn/M0dDbvjQjTFFR/Aun/3/2w/z/ccr8CckYcsKU
V5fx7HnXCZuJZWbvMBo9VL+591eY2RfaVje3AVn+rGIre/q0Ew+UPTij04zjkcQQAseIgD00ev+k
PQVqU6lYw0sKBe1d+QVUkIG9bbmFy881blhbrr0vjM14K5u5zSdR3E3ej6owyQse+w9B6MKQvTBE
W3K9prdZwgBRbkwuurDy2mlAIrZBbdrNW3lyE5rQ/e6wBMebjCZH4XUuBK/WB2TK7xoSzw7H2R2e
IGw31R3IWIj6hDdi/o6t5/2tha+y7sOEZn3F80JBaYaJ+ZuBm/I+RVYlplkrdRciAWyJwuYaifXd
s6Tq1r+DsCGMPMFLp5/pls+gyTG02f6vXd1viWZXn+LflMq63FG/T3TkKDnRdR+hcypy+UubsIwp
GWsFxgrq0PldlbykpHPFgmvyTWEjq4WrEBxjLsa+sEcTMU4EwELjTt9j/0B/Jvyt/ENmH7RhFAg1
rZLz1iEvLodGGZMpY6iFrPMueCMzDGKwc1xO/3FY8yWfhEKhJxfrOgK0aMkBNKALHMWnAl+IyAGB
6BirYbkU7fpkNm5itLEoYleZgNhkWOO7AFxGTJBmdNf9MsSJn8WIoaOxbodUtzH0dmX1BWCXabHp
bC5dxgxeYtb0rcZYzQXPdjRCf4AGg8hLwjnVl+nDA5w++XB132Cnl3wBmjlEururkR/WkBEryJyi
dKXxWSkp1Phisb03Xtv3G5eU+JGZaAOUNO4qA6NjwDtvS+V5DrQFItP1oqLw4sSx+VFOiCjG/pdi
IhBXnsCOliKU6fibm2iQ9gEPViQ4SpxkhfL3SuP8w/oRrAx1uw0t4RE8w7ofF7bRijZ9kNyabOb8
N6goROATHG7sVJRa/v//DLjDGRBP8EBrbySrpxK4EcLiOpYcDcT8tRnYwQ1N23dbiAH1djbSP+9A
FOF1HzEA1IibjDUc312vaHehUJYG7QyqhTkIqx8g37LOBzLWuzNB0wpUagER6pKf0qy4T7P8fAlO
Juqxz8vbho2XeKEpfPKCETW2GnF1q2X6coQ0XEAqu2YGCQIGgC7xafXolRWsM244zLQe1i3DBh3e
loFS0H/r8L41a3/wkK2E1UmPrmuQNvyN9qORFf9crz7f88S/ljwlhfOnd8YUHJsrhDTQNi7RYenK
Sq3PtVQ5OtP7Ku5Okkb/DDY3ZHbbHcgnfFOFucpeGcUZLnmmZNQkgltLSZXIGllo+AjnfDIlCp7m
L3MPf2M4ubdTJP1HQHxjYnHRen6wo9YSXzJ/b/CGv6sZeLfaKB9g/B7FkPSSIorQtxxuBHukgSHA
XFwFIMTejKaq+CjyQyOP0YLwegxQaQ65jwfFu3Tz1rbtSWTpSuCYEAx0K/0E9UkdQvpoIbcZ2qFj
X7ubPl+Jq5XJJFDrktqjyMBW3iPv8ILNIg3ocpDlAeRUukhRap9TbqXzBJDkKGCjtfbcDzUWbWGr
VS+eS8vkPH/l9J7kIgEF1rICsJ9BnxmDveHIPr7+Em2IqoDj8UEJqU8hSAoHk+tANcAGE6H6JYnu
YokWQIDVaXtgjmhzGFN8zpbnq0Wg/hW9acimOEXQz64AIOhVOFA26wSRHq5OUEYcvIwX05CoNKAo
LTlVOG4TAcI9GYNEmXuBncePae5SVf0dVgcFeki6ya1vcsWZTlLmOK4pFqZ0Kf1ZBgzaVoytvS39
f5/zLApdCjBxXG+/UqyeoBK42ptnGCJD8VUdB7wb62i6NnkH7EmPe+p4adFQi2zEq18HS6h4//Sv
CsKBwOi60TJ+QMCUPhRxnllsM5KzHS6d4uWuhJCxDEf4gTVGFoOCrE60moyQoAJqq4uhHB1SxgFc
YiIvpULVI1OU0XGCuOH9AOpwq5iVdjsxZ9BxKzqM4DbdlBgtngSIMBXbRsHMqusH++Uvv4Cax5d+
Y48icQ5SvAB4PAGmvWo4Qil71TkDBRV/n0wZdSb2TqIJTzMPYCBC1GHQHaCoMN5f/tGSs/JkmyUm
bul0omMFky/wTcGN59UiUyp3DZ4XHZ+H2SZ4C9o51BHsRFvZP56fRCrDJr5bgN0jscI7tI3gsYNw
oG/PFTI2HddtWG87GkjE1bFBbKiv6vDnNuOsYIC9Nq5ChIDrc2LkEUNUjvXqxazvzFvEOd0YXUpQ
n0T65e3O+WDNxyRPD4nZFO3ZaYnUsjOO8fbDnw17SacjCu21FNgS/z0sEp6fH2o5X+e91QyT/4u6
KXbTUgGFFRrUHmCcdm+Ydnh6JAqrENm+0i+ZO+QZR3LVHMmAnalcH0ZoMQudBFphg1IgRcXD8poJ
cl261D8UPkUusANB+g9GyrEuHYb53GYC2s14AFDpjRTlXgxOWNoeELti5fD5gfcL5kdQIVY77RZf
4PdtH0Hal0mTDqCU1Z012irNMY93M2xruQTGbObegEKPlJrK6lzjX7d22B82zuHAJ6JzU3hS/GWF
vb+7/ypKC9UmO3RNbLUe9d/Hf6/lReAHWytTD/eIspk+Gbl97jYvo8H8E88Bw2wf9qjgSvnRQCj2
nbtJRD3Jvz+eVJdWqMYUYSnYqPkepTsX6MyRSAnw7viROUokmWYIusy2ar5u9yamd4My3PLwKMLf
/hWTgLuPVfrh6y6WVuz3N7zveCkJAIdWdpV+GHJBPMqd1LHc6+OCi7M4DaziwBRQOmF+rMOXKSw1
yE7pJTOlfwWB9dn/mByc8NQMnbMnBP7EJHjTbSRJLp2XbvDHpoLcL6FiVJNq7UreKpimWhpyB+2C
lm8KGt+ArpoNWyfjeUuNxID6fvZJr7QF+1KF6ulVRFhF4w0TDAzhIH0Q0AKMZPVNkJ9s6VM5cMHP
Rth76xCFyDwRw9qFYuiUG4+SZThhwW8mQD2HjI/H5/M6MU+A9UGm2nN2/6WrqvkG8PYD4JoRY2u7
tWfjwHVLsDklAiPSWGVRvlW04yTYJWxIFdHVZ/TzuL1/L9dzw4RhA+HMZJ1tPdd80YXDYiAUo/PP
0G9tdLloBKw17/8efiP9GElV84I4Jy/YS41CL/PUwBvdtPDzGDroz2vhrXeTeug37sRb5k38Lhxk
e1YYM/kjc/YiBXYg6t5UCZgu8YNyV1e7YZm4FpKLiT+uJf0MwztMy3gbaPmwuqY3Q8qm08Fbo8El
OFL+9yab41a3jOXn+/YCV+XV1fsvQ8UDGwQKxsogZnEjOPcZ62gt38G4EaATGqdR/5fqAVNEz+CT
qrF+Q/eBXr7JMdWFaYLh+TMWxQHVAc29fR5D8GuvbF7iJUA/GIVjulDOIohM8f4/DhNpp8fmKQw+
XGoPNkmxFgpfTtlWa/oAhEadzXcqVYDfGdPF7cFNrtQUAYHfHd8f+USSHFPGG4jCiLVoqsyH/90Z
EISXVvJZq/baGb2QbaSuWU8H2yyuMVwNaaqOhS3ys4Yb8tkN2NCk2/UmzbQY5LcJgcIwxpLQkViD
qaxplecy1LlvcC0h9Sg59dwsvSoUHTCdV3atyuxVBZZw6OA18Eu+rqIFM5mZ2d+NvHR438Ph0Bob
1unQPlz/+LZLeMO/20v9Vp4VMcLxXrFsHTwcbK/zi6nU8FNGIxINq+wTzt/4TAN2AvqyNucaqpts
Zm4xDxqD5Zbf8WcV+OXfCF0MsTWfn8R3alQrDubGd6kzphqGgC7fhyULfnrORb25buPrMHqestHo
zsUK+JV29sVRxhK4P8E8Hqe5vAgXvzfLpr1zWGxajFc4PjiIza29oNTeYQDV8DGzbTKBmnl5CnRQ
a/3oGx8Jegq84wxDRK/MRH6FIbmq4PyZ4yqkegNcX4EmV6Adc1PKlJEQJ3o4FoqYnL0/2L5jhoTx
yH3OGKQVADmHzNo6jzTSFfwIMkkB5UfHEWZSI7XCA2jDQk63Sx7kO9WnPLYLkI3nPTdtCCfWbF3f
uiL1bbvym6gme8ECP1Rf0fFP2O/vxjBRsizonmhfGrGUR7X6IeUhf7ip0/pELgREmXRYTxThWkce
c3XtRPbLmAAVvOxahcfSAviYxvWSxxj/wjHFKXpcsL37lzMJhE9DnAhPHu0GWpEcmVImM5rGhqAR
LLxGGWNcbd4QT0+CgBD4DYw5FLt6UtftgYUJCaLboLVbONJDCFTAPQSCD8Afbm5ln+AjXsgOmPbI
hZg3M74juY0MQOumg//aOStt16b+HfTOOrWuwCCakNTBOUPc5KGHYbFsRbMZcIEsT1kcZT4xEYA2
hifvwbpOyvebKLePBWLXWKKn2+ciiA5dcQuc2idSGK9Su8yVWEBI3VsqSAd/GtYe5IqHdRG90Lwu
ioWm3LItNLPQQcFFqvGx3+F4ApoRGr7OLd9QnQUsNjERBXhScMAD26RO7q5qh+JGvL+oM9G4laJR
J7kGyrt/OJ+kQ2HeldcnPkH0yfUPC+Wej9nr7hrKFXNRpN7rmPfLYsSOC0vlhN0VDTNlUcARjtkI
4uaO7cEEUTxAIGK+mBdIWbq3UZn3CiXCwIZ5OywC5fOj0TB4q4eI7Uop02fIlY6Ii9Ar1ElyBEiK
j+Pfl6EVA40RB5Cix+lU0+tfPTI5fK3QnCUYt7ZVMQURJhh6ZNWCCbxwHEyQNU8zsAUiWW+/nx8A
0nf2RK0yYlDsdX4TDwSbMqBOeMlNQqpl4x8ZbwntuWtJtwLVnRiCtb7sys0iL7PQ02zwZAeDKG93
U9EaaoLHSH4knTjabcMzapGgLof9J6l0SIL/r6N3RDZLAo+Ccdn2mIzh8xiLO5q+IpzA11s65tjY
if3EWmmtjpQfId7vljXCCqm5wkbsa7HRDVKIRbtLGz57C+7DcW3Mwi7p+c6d5Dknz1EobA+v5/Fj
Tmv3dOBs7h3brVKbRyQl3IKUHGrbVt851+zUIf4rUoSt/q2hGCXGxrn6AqUBVZwCQ4v4K1XvgPxW
AXhawUkfq7yy+IGG4cJgAkmhhmnGH+2Pr/nP89PcD5kYnDdeEY3p22D3EmVpULfQQD4WHXx6vRGL
5Kzi9EMsaIxfeXga1UrkJA/wcYew3aXlVG+q1C6ydw3D96a/+xOQoK6nF83mxJ95ECOokEJOTOij
b/wJ1eEnGfolTvYGWD49hLNALBvz/ahuT9zTyDIvLoy8Z653o8jNcnfU9h3lbPozFFt8UNlTSrD3
GD6Wj+qt+SWr9Vbs7OHdKaabwN2HNL4RC+2LmnRi9bT24fIiamC6HvXcIkntJ5zx4Tb0xgbEnlPo
3uDPv0LOI0f7mn0nvTVLjgXoXrT/vleO94crYfquiNPJj86hGwAXjQU+7+R9Sk08x46CvbEQppWx
uSkMfjoeJ7uUbQ/E21e5qVqYJNa2IHW9sx8+3IihxfVZid9dXWVHBglJxgX3PLe2HpfloWQsGd54
3tVi5lznJGx3qX84wa9C+FSaLTOesL15djE299jDvbD4KyhV8jHSqbkKeJxYCz9KsrTZymMsuDqd
9T+7jqk4lzeuEwDsjpn2sth2zNFXZOWmXa3yqi9hQMU8GjFvOY4QnmLWggQpG6WdjODKbBpHAu/S
Zc04P2oThQsFjn92BdpUT+6UNZkeGgU89kcRgR27/T/VV7uEKwv3G0CK3+AnMB0j3HtXpa4oIw/u
U5D7xHTp0rVRDiODdqSDIz2LuE9vIa7RG82KQTkPIoOKw638ss1k7fZvTCHX7/q1+jzuHDr8KE23
n2J658Yt2OwisCeB05mz5unhmMGez/sT/JR0aGytc/UzKWFyutV1bn+vHEy2Gt8AUl5Op8JuU2fM
YXBT7SSDzP+pShhPdLxk0kay/fyW+ZoE2d1hJERSJhgsO08rSREFxjQUwc5/58jDnEIH0Mm4S4nk
cKVE6jb15w7WccRbukInidGzRJwTYPbkI/ggUtOByq/IBT5DTSaZXbtYPsoM24gLQToM0ADJBefo
bqlWmzxBU+/6PPTcf08XIbqK49vIXjCvLb6WDM5EebVxDO2h4FG70CQZMdTkMtTlMabIZpskAr7/
vLy8oXzr60riWfX0wohiACSIn9DIcZRs1X+jxUBH3NeBFWSA7dvlr6dmXeQo1+t+bD/fvNPz1JYH
/6Kgz5/1qDWswJV7c0D9DuY1rlTrahkjzp1jEdUdxfczBSkIuv6ZwmSNtgwU3sKQMDeR1JMOYT81
BhAhOx7MYaMu3yYYhZ5838DN24lKxJRCrNRV4JV3wBa6fhCk/thNVK6XYoE3DySC38HFf9+gPpPe
UVzbvXOsyY0L+dYICVWHm+0X3OZeo/kTW0gH8neVKwdGzfKXvOL/tyX9uzpI7lbCStdDhRtMIXeF
mOOd+i+ARNSBVHU1aRIFT4hBCciXlJVuensZAQdSufUSB3EEsbcfe1JYXgVZHfs9gx5/AXoUPW3d
QZOmHPIfNcqYekNotsanag4fll2IMnAyJUwolYo+deYpDbkOzWsXqLTRTsesE8uhjc3kOTKasYAv
R5HcMB5mqpI/r/O6qoIJuFqj4GM6rQL8WdB3DzYDW2PgyNB9nxUfDu/hHLi6vUXQuWH8JjO9QCdU
mqU6WiqrwVQ28aWrF906fjemYSb/TpNZhITT18L9eUsLh3JqZ0e0VayW/sF7Cy41dc9dwUrskQbf
IITNv8COogfVT6CBXMPiKIRxBSaRvX8Orgr42EYQLKzFpz8dAB+D2/uNA9E7zZolmh6TnH31Rukr
t1CLNC9/vLlH7ZQ/vuvp0sRgFW7+W79af6SfwZNRRf0uOy4S6GiAZlmkDT1ecF7S4KyQ3aH1I35Z
fi91ZdnBdH3X77vdd1WWMLAz7jrKr6kB83ol8J7v8pqW/rz6QTve2OfkwlM2Rfpg8kmDdY1tH5Qw
V34e+W86QJZ3k84pkeAgl3jnnf7jSLSH7sPWcJBNhnCHklsNyPg23xvI4bCRBkLX49Ccz4w4B6CX
jCuR74IFNP0YlQqCvxLRAnqxsqXOsJTqt1f5fK2SMEC/NBn/QJ8mUOMqyJuiw0D7zPmr/JqSZOLY
7IhfuTvGqPklELZBc2HyMQo5aN6802QCTzmVWRyZJpG08ezKJWvKHIixjxJ1RIWu7WR3R4caNXtI
2MlR5aXlSbLlV7q+dQwcWaGKMry5I0gZXdllgq8YUcUKov2pV4PwPvGBXGBU88Da3BPNSqCa/FDH
C4vuKU+8q3QhlB09Sr8cd6YSRYO2IlXGyXTl7cSE7NIAr2LPyZUN60GkkXMdbcKt+qhn0VDG6Ppa
vlPsftff1CzV/8qOBSmI7AwelVzuSLE/NyhPAYC5jZP+Ktb+hdxXjzwoOTDJPbgHNMocqcuRpKKC
ACcusg83dHuPjg9W+/veIyPIYqDW8xtac7MREiDI40d/UwaRTQwq1VCE+NefSCTlLAUQdqxspOL6
ewjbf0n7gngGfgh9oFJ2muHuoUlujZBAsWntPevYBX8PDHef4L8Z11is6E5HfrCjZZC8kdG7uWZC
Towb5joGNzchSqpavofL20dU0ZFQfvWE5yZZRioXFWoFZQQud/lsQi6ALLIJuVdy+OQO5dGZLKNG
Fed2exNd4vzNgLDDs0RY0jVgd6dkHCBJvuh6fwVMdAFUGxA5JpHQ+dubOIrg0wLqEKu1i657uMx2
J0rUhnh8Bur+1H9JdZfp8eAWigNX26IS9yXQEM/Cz3vEd3Sbb+I9uTheKnySMFvHmNRLr43kVa/C
PF9yzVOyTXPPEf2hKHpnBMoVTHmEd08ZQOnAu8Wczl7JIksFoAH90xIc8bPsxqDbE4Ay31JYwRMG
73OIcxrnqwa7eutjEhpSGHBISbWymFS+k8QFYa/k4n6xdo4nKrnoRhsXajbzai63oUwWjX5xK+Oy
UL30sr4Y9z0gcVlg2Js1OKlPUO1jlWMksL7G0MSke4e1EzhTLlr2yaXuNiDFJv0Ao1urkkLLcXBZ
BqV3Q5WV+LoG164JOmFAryRyprfDXEu6B4VqWDF21t904iAsKo4yrwo15n10X8/TM3prCEh8L3DV
Wb9hoAKwiDOh+RTm0YLJOdI/qFM5PVNyzKOjrZOt4AzLP8jxw7nOd5AjPKGbMXkUznF5oe0DWpDl
Dx/UnklT+y1oOIkU1TH3LA3o7icW240Cc7LNOjLkqxMwIHNZDGTaKrNcYjHr5AvHK8RVsPY8jeHp
0jGNiAMmtBiMpiZA0vpjlueDhdNX4bgP/3kf2snxmSaAmn5AcVidqr1WB7u30fHm5LpwPU/s+zsr
PvIbGNh+UeLpCrBzwLME5ZpI2PeLkR4ZVAmLVOopExpZ7+Ut4NtxxMLAY41TQRZ972tEGEqRhzHs
cNtBC1vMz4MW0ZDme9xikkdeNJYyMKJrUvmYisvBhcmAec/dLdpTshfMqgMGmJyyKKxCnpyojEpR
+wBUPgRIoHB7drIUmu1IzPohc4C9qD2GnDhsjMng/CYS0mjggoZyc01YiGQXPKCtfTJbFF4HYgJs
ts16HswoX2uZdz2NU7LvZsejcUQViDDqYsphI4bzVAIK9IP/KPgI74rrnv8Q0a/4ju7oBlI++WQK
vH1Pbhf2RhS5Qnhawf6goPEsW6JsajsCu4elTsD+JPAyuXdoa1ZRrriOoS9+qXFuvsODwotUOYM/
8GpWnvF87+Y6dRiwI1NqFo7B3CdlLvCocZjAyjE2ZxHE9MCmZO7Ltkj2C+ZN4zpHT+3fwJiPCMMa
AbpM8jpgIASy7HGNlbQWY92/Us89SN5foaLZl58R+wOb/oDfE5nyLIBmf6SPFPb/L2Re/4cQGhII
rDOCBNCWPkxl26rXWE9nyD0OT2IiwPBVWLRSBjhPk4EPPHR7/J1DemkARfvzKLBSTqoaZBzby/Q6
pcIQD/Hplzo93uz9rCJUVd+0lAVRtmad+etjuHl66xoq0vJ4TmHsADdaE9QtHa/iGBZDKon4p9pP
5OViVodngQljXvkN111HdjHGKrUL67Dm4i14TyvI+vtkpKwcmUmymiJjNGSxftBSDN4H9Fn8scEU
CFLbgOU84pkT3/8IkpGEty2xpGOMZ02LKB1u/0esMikv0syDhuqGCunbIn6tNMttB1rlDDEJyNpU
PuK0RXgct9aomzolpEB/ZfxD6Vku7xbr3GyvA2WgFzTiZFwr34zeUMYuShbdHeuc8XJdmzMOkG0K
o5tT7nuv+BqsIDiSTvvtykQH/iRQ7JEMqWW+sv32K4IrI4mP9w/rzbpHI32PsFau0HBKWNol6bPM
wFlt9nGY8MFoL2xahupNhLgJbba2m3PPGArum87jBeo08wG4eGfPK17bpXbHTQV/2O9N4OYZ+M/H
pFe0fhkDLuq3Lds5t4uOSNpdNVHO5Orx9IyNORPVzkyJjjUqRtgJC0HIztXNgLN/wnWi5t6Eo2C0
0l42mu8MsOIxMiqrb+HTY97RwRWLDakFdjTBc3Fzy930d8GRPjzUaX2F2tqsg7G/I2f1mHqty8di
FROhsGVlA3u0++KZ9F+Q8vApdlRepMIBjMafXWTWeiVjUfWUiNvuC32tyoyCyBX4RTB6e/dcMKrT
N++3Q1LIIXenwuUBjxQj0sPQgBL05RT2iw+/I4Cmzb3ZNHHmAGVGtPJW5tdNd9bLLzGUO2FAHuUi
YR8J4buoFsfrxoz3+esOCWn2Qk6ePt1xb6MmED2qm57Yegz9pzbsi63JI7RakcNycewROCYiHVtB
QKyIxXIjtsIqMQiRYNASG2dJ8DPkdLwR4TS0fR5XCQqJ6likEiMMFiZpCmdctcPgkmH1y//XXSDo
977skqZR/qOEHXNGq+e0nzE6KUYdSRhgWna3ziulIFW02WuvVt59W0W5P6Spr7geAlck++4t953p
sSm5Ow/AL+N9IUK3bVs/0AcmEbtR7PbW8PNsXSdEetLtLvWDObkETRglqrttTguX5GMdv6wy6zi7
qeJtohzwIC4d1ZY2d8IuAraYtow0SErXdEbeQZIjp97gOXvndiu7JNfxmtQZKqzXAF2VysTigyZF
Vn5pGMuJ0hGdRUj9n5QEgqDBqVqoR/T5I0bb7Z9LmMrOk6+mbx44jjgTItciVZYJSt7xDl1JXsw/
jj4mzv7Sz2xbIdZBlz6xYBhTMapdwuSZs4Wpf/bITfkQW+AHczphskKyNLj12UVdlwyY4gQWVgGr
WP/uAqPGXDoFKnEGdIh1JVjwmzyucysxcJFg4xpwMb9oumxTzwUYaz4nHNZTFtr/I3Kbghol4G3s
Vs7WgxEKdUa9dOz1mhmgTjtTWhPT/kwQaku4ib5TQm2rx2ly3snhWnwe2VlIQjXruoktKgXHl7GU
pcO9r6CTZDAixdoMOYxgLXa+vTgI3V1uRjiBcY68GbU4JZ9oQYoqezzzLmXJR1IN5gkGTMOUGdKi
wiMGratbo631UlPub883otAgd0bgDee8gpwZE1vSZG3iay0NtuRgA2WUlwuBeifjNvvoiPMX7UkU
rCMgEXgLKI/CMDj0Fm6Z8X6Nn3MRTtOrc4y25zcyw27/s5fQgNPm5K1pFded6E/uxDamt5G/LVyc
FRBmEqK57pDrJZUIIe4tJNFD2aEhWzn1ogm1+rjP3S2cb5QP+DdCvgzVE0Y8MFOve4a/Z463Iwhx
XwCXXEhYHLm/HHQW9kdURqSSmTvCSErIpBtjX2lyRvQ+ywIhD2BfTQAn/FX8ezHmBvL4/d9F09aK
RslE1AxokWIAMcFtDOJ6Do39D+82SMTzOEUFnn8aidoPP75y8U68aqbry9bWNwXrNbbymWUw3Mmy
LqkRnBNaybNlwjh+zO898fG3FfgjppWo7gaZI3TOMvqQWlv5eNj8aPIE7XnQMl9vXTvVZYIf0biA
Z+r5Sn/yC5QLA3L6SkjfL/A+xM6fSrSTQT9QFne1VnH740qz/dCTU6NS0evCuj1d8k2Ep7bb9LDh
HBIQao02eX5qUxOYUtgV00V76eLGpsp5NxXd1bUsZrN2ty7a9ymrWdQf3vu3B5EWJBsNvWQYaXUb
B2d0mqcgOOfsBS40CJ6+h/crq11Dj9WXnJd596vLeIWDu5uAw40iJ2JMoWlh8wkf7vLSvLrwWUE+
ft5YxHbR0SNEXq9nV9/sG32RCbi8PpeVHWPmHunKWoodw/mxygH3yjItJFeL1mJAm2N81vOefmlG
F0jyutD1bz7vZ9r3ASADD5n2zIMBESGwBEBjssAPrj1kwKsj5PwEqbUoFxxRD8HqhjIa80AxjIJq
zRSjGkB5xRAQJJm67sfw+dkNPBmHZ8rg3evYTGheEO5i/5mCkZ5OkYNQKv4+tonJ2ai42j5D44ZD
aUhneXX15432mnwSGeBijiXT/MtcapqN+0vEM+UWWhrY1sfPyO1Yf42yDJZxzSfOguTropFsz1cT
b6Oz2ZFgOqYXLjSziWAFzkp8RPAqwUHlCrGdpnDrs7xGSyRf3sRfrmYtkFKjz3kN2J85eXCt6roQ
ISr/mP7k/W8FrUxEXrR2WAYfjHTNgq9VfV6GyX1h2/MwpSxTO8QzYWzylbcK/oe7QRB+qNbvkwVb
n2XExButElcl9P7HgaIiXe/iTbKqiRvF3C95NgAXkCgSTppG4cMu66ljFh8p8HNP47858nodCqz4
g5o8/MGPz62vvWKZsSlONHSJKWokh7h6hyKO3uNlQI7JcDhpEXDkMFcWzfgSa1eZSaKdiFgSlpv9
B2W+opk71OOgQpgRMOp3H9WMdExIVAiuNexpbLt4PkziTuRhMyUsVgjlvRXY6Ak/IP82sr/MyFX4
Wj1lXjkIPeTJRQEa9Ti9i/JQT0QVd33zq96/P4x9pHhcgUyDIDNraKzbfR6lyAWd9+bDF0mkE/IN
oZVXMQUBS5TruPL8jT4wADXZDClOqxMNucRDfKLYfOrKDOV/GAEgtS9rhSxTunmUgGvHpcB9BPqa
P4N5fTcqxuDgh/9ymEMddbDniHtw/Xeap9fGRSWhCNlammTgUn2udzkbusD2Kyr3duAxdsALJfn5
c6bVzKaD0kBBRRjwvlwDJBlCzWF85cqbI0xTqwIiP9QQKYYrI5gxPGJExaFT7nV6ir1kcIf2H3ar
hBNfV/3DxaHKVrAudIJs1gOqs619bdm75cZnHz57sq6uZFkB5l+NL/HmHd891oH29+8x8Ep3myDN
G/SjxSEjMnUbe96z8naDmF4U7+b143gs2eDkdCK6b66i1mxac0igzGPbzLqnUqfS2b6LHehYo3PB
V6SUN1pAPFG2TdDj4mzdGESATg+/mm5GOPimc6PFTSQWL7RL8qQe6P8CcV9q4HGF0v1uPQhcgoAk
KcR2S46AGGyymaThmqErBLe0SBIg/mWCEMjuZuDvbHqUcW92BZbc+1i8k+MA+HiwfuPVGWVpYVhl
10UqligovbYzIPVnxCBPtw2dfyfNAY1DRopjR3bO98+d1QkieoxL9HR8TZgTiA8xqi7TAwZooKs7
RJ5EKJlk+bSpkyc8bT9sApqJmSfJETdnjkskNuibAOWxC4s2sY9AzpGF44JMPR2+08bBSO5FgHqS
E6Z/exci1eYSf6J091fYNAcrHnU4XXkYGHY+QdNrnTAbJ+8WFQoFVZBESdbGiEoTiGeUItqVCXFR
w4hgJGgAGnw+QduABnDfmf4vAJy1X5Vx7B7R5LQYCWmwiWJ1C3QpyjExpOoD5AAJg/nR/nuga9Q9
vkn0K+3qAs049PN8pE1BOL25gVH+eOnB5iC+UZ+e9cX/Cb79bN2P75WmgzAO6eHt0MQuAOq7QdOx
YIZkpfHjLwlTxnxUmPB7SSWy9U+NusaB2wfuAFxBYRaQuazrMDHDo+xqGixLcGOyHtBU774oQ+id
fFEh69QtJUXGlIx90cQXzr3kixFtIGEtHg1P08zGZeCPfyinjAMkIHv0o41PJuBVBVlFVXqiHOhr
lwTlrBM1yRbjXeyb1vcDrIObldqSCNv2x/EoH+1CKpTsTjFMuvqzBstSy/8kA3Brid4O6CLXmV7P
w+4wvfScdj+HShl9AVOTcmBzrS8U/Gh47X/82MqYm/EUDKTBHTT8aXVzrFGjxeSUba8xSS58O974
gwDxzazEMtswjJL83tQ2s9H7L4LVQi6G3CoLG+EE0pdyqruvwQDlPp1qDLGmJhvnsXPP92p5Cs/5
R//qFhIBhqkTH2oSEX/hXEmUkKSmEh8ZgrXZSOgERpIGKzLuRz2PIR0djIE8B46Z4AQn92ca5yCG
CQMro8C6+pZJOmCgFt1wCL3T4K6lnJV4lvaYhCkD2nqBiC5YlMg5wvsHHgxMX33aU+NN4/p3rXr5
iGWRl9q6pDs0AmekSWQkszQ78iX/WZ99BLhlUg1vfi+j1XmxV/2DCYFt1dm0+w/MkX9OCQdQ8ywA
bqDpPGpQQPZFKUtuWtkmE9856dKht4ABSP3l8pBACkwU24Dsox1ExtjKXbPfA3wKgtJtWbeZoI+9
N5glIMy0qTxcSWzD2hVr00kRPlIlyqClqboLziGOYY02MJOkCvSJ3O1e35gN8ICrMyd81vhELl3f
CqXDaA8fKefPwpggtOD04utXzgxEAvZy9s2TnNSOX6i4fFc3nY1w0zZrIgMy4+PYvcg6JlzZr6xZ
gYivspOuN9elpRSvxZH8NdVuZPwylB75zZtaxsAl+hnwjI8KWBrZQFvBoPUt09jSD4+55v+9fL2K
MW5xcG4lHXmLzQJbdyMXlEJxZp5LZ1y8xKGdBJL+dntv34J2qD4zb4EgIWsaixs5yJ1pUPFPBtFC
P281HJg7oirn7/k1KaFBfhzl00kGhCckNIIl5CYCwAWC3PRLk7Sa7RD3b3cyX27LDFKA7T4cMcYN
O8g3U/hAiy+nAuVqIbWi9bxDIMc20I2MgD4quPbQUgseX4K1HGLrKMD7mIb5RwZRny2Prrx8OQRx
GWrfcZ/gpomBtlLKiVRxpqyR/rBOSPWy0I+jvZni4XbIcQx/X1V6Qq9UgTX9fxx6ahrzD/W9heKl
vzPB1d9CCq5N5F0ZjT0lVjvJwQJc8B9NGx1kO1JK5mHg5ylgOPtuH/ucy+0ZJJlt3x5yoZD3GOd7
Gg2Woj3pjCHC1ub7nNjBm5a129InNKC+SeBIliUO5tbbSV2RVIa+9Gy+h9umxVP3QjBQZcpZPR49
ZmHR6q3w/pZfVGMXzzTM5NkowTpkApdbAtrIuqj5c8g2gwvDYmwbKXdC+6kdeDmfy7P4OhI5MKUm
7Evp4fo//HA5FDv+p2wXQYDPbYCf+rZxfmavmNjOGYRCUjsvTOZZG7AnFqRPBv4auJQXx6pmF8Aj
5KE+tAJQcElhR04CfLS/7EoF09Mdu+zbR/98oMoeubgiA5ExyH0ekYAaUiSdMt1r0nxNIaT1yM5X
fSrYj7C9SbnoQd5/4B7YmHzbdhspfGiuHQVxQzgnZ0jiE89/u71iYDwdEWScM5umGQzMzNQ8raKy
6DVkAIxVitjIfijfv8nZXuoLXR3FHWBWGQe9AbyDOWC34RrGKzVxo2mfF4Te9U/sjoy2u41UfWaq
pCYJZENA4+HhAchzJAyALeb5zYKZcempWaFQgPbF0ldP92fH+zxxWQWFZAwkFDnkzCmEtv9vFg05
Foz5sQkriSwnT4z0g8DNsBIE3Szit715IOJSmonk6EVtRtwhZovUO5MBX4l8WITfb4x+PyqUzAFB
Nh5zMjf97MKQx6AfBBnCY1Qjh3CztGBRF2ouGvhPyv//T1pj7vv0MtcGs9CVtlyZ27Iit1T/RVqM
SQKwtlWd0KYMDf84EXzHDz+Cyzm65p5F8bnCALW5wI8pFb9c49941LzVdyXmR1FIUPw5fo46M0jU
CMnjUiG+LFln1h0i2EqGE4OjXpkH+5sFttFuhtIjnmVk8IAgGNJOQ9ZWUqPIaXdYjIqzegBRWFkd
xfC96NQALl3tH97smkUXK2bemCZ/IiksnaGRxQ+N4chN6Mg09llkbnzDqA/+n8Fzz6pSU8U0VDiq
0KswmcpK3HTITAzYScP0TTgthOhVoJwrOweMd/wvg/CJcdEmjigBeTpSF5fV4+KKAAPY/vzGpIsg
xYUyeHNZlinycmXEToB67YEG6ob5cZ++F47c0wMqe4QX3wVmcbjwBgQc2cEGiQU1GGBnboeyPBUf
vWSzzMLjkdS/hnJ4iitggf0CKg6Bl+6F7q5zp5xi+w/AKKIwlJ+s1UHNpZez1t1Xu9IgPGdRt2cv
Ku70NaUAWeJe5TgKGih0BO1ej5j1zJ/kqYXECXzbbt9l+MHRuRHy7jPO5D+yF0K7M1hE5NL9S8ar
wbYQKd05zr8Nh3d7WtGCDXcm+SQN6QQUF1lLl1mpAfS3MAWsok2EFZIJOhgy41cGURdAM+2ZRoIP
KYR9FslHyXacxVS200AjN/fz8iveW/0I3/C7pLjHfJpLG+Pm2YKH2HuxVANYaZacb91m6I3jNg5g
igCsxFup7TBTWI9ISooE3F0TgWNLXpZLQZhY0egZ6pyWXzIJ0XXLraQG8fEUF4hMWQUHx6TmBfVG
N+ORdoXbFCXTiQww+cUo+2wiUrLTGauu8KO8yblte4HFq6XDowTjdwK+DOixSZSwZ/gX2zRCJb93
P9OrqATXHpbrxqdXfd8zabSutYx2GiTa0LlS0U/UcnxHkcUQqhyzwhBsLMsdki3qEDQCLHR77iGE
bYabXAPplM0cfUDuL556lhRW214ZB0dJ5vnxjznMbCTojbD3yWmzpOrxiaK30y6HlYdXBxJ3ICoK
ht+WaVjXZil9I34iSpdIvPz0bf4mKxvEs4pUqlGC+0yjw29gXLYHgSa+5irHm1ODfl+okxJqV5/1
lnROCyinKKkQn6X1BkFIY9QbkdcfCC9yfktWvcoZTbBNrJj5KABmeqADHo/qeGZiBA36xeEZ1drR
bSONnwXlxWNjQM0ACm//gqbBmeFEeyESqyBoEg/pS1J+SLP3yYhtkmyHFvZ+vXYQ3IjrOzmtO2ET
bSU+DwE63Ohs0trPwJZ4thaHmxVCgMc/NXjEdj05TnKxce/sXHdmcsIORmZUX/VwIFNy4RsD5BOx
OqHpQqqJPCV7dYDB4p5rtNCqsJgo5Z/tD7Q19OTNZRbehxGWCyMFcQJQp1I0NFNVMjmegGqURMJb
BTtZXa8I1SSRl8ehv7H0OPIsso4eCS3BuH3u7XrtpDJwLG+sXoRe3Xyz6D0tYb8Uv/l0JWFuCgZ2
CtfLB9JQSmHj4NFcdDnv6Wu0zP7Wvw1AbqTws8EIrfhp5YR2s9ujrsjxIM/fkKHqr3KNz8Tm/32B
sALpoxs+eBHQnH0J+oJF+5vfbOmOw8tpAqN7sNusb6ENIvjSYJKl6RjF8YbqP7RL8n+T5U7+pa4L
7gAJkExQXgJxvv4wFNj4Cx90S8lIsQUdpzn6RJbydJgVMrXo93wdGe5JzLk/y/zhDB/OvAmzYAfC
dO2rOBzv9sDqJvsvsVhMTagNoA3nC/M6ywgQ+WUvLQOkA2rr0mrOGSmWMMs84/2IAJOtzcxGEJqy
iwPI5dstL2bsJJ3GnSpBfhJUdCg8ZULoYLvsCEEFGWhRKxIBhWdgeg+Rj7yYCz018jBQxh7cg5pl
hnMzlAymVdLXEsnAuPIZ3d9X/wAwdYVuP6fEL31IjiBaS3MM/er+3jCoqe0ndJBWNtaYcAj6xAq8
/UkgwQAmV/gR9dWCm1FZdY8Q1yBOq8WeCcGUh0dH42vN/jd1OVeBrlminDUvBDhcVG8hfR0amPbp
ZwN1K+NOpRO5nj34s9iwqqy1lbC7q27zvrMitpRqRYRY8RbzVLQCf2DFgitkMFRx2Kuhxd+nPDmb
EG7UmZPSAK289UtMMxq/bN8+EZeYRg5xnldHRMvUgdI7hzbp2VU39/wWcf0BfbrzscBoK5TR0oVd
yre17qF/DhLyXSmcQXb8S84Im8lcbdjLoIYaPV5BsBEXje0q6iM8UVfOvxnoCFDEv3eBFEfirkRP
frEqxqvMvWFsqT2n3ISoSeTutQezyFQn7+HudxEQpT4eC1GHzBuKEi4jZpqR10kx8s+mb7D8wvGw
OVZUUt8lVnfh+bMTuI1qhcfk+SqlDHzUk5UWanRcTtPa2xzwgle2pw2w5jjyqdrRHk6EDawGM2rn
Ce5SoyE8pNFXAJINYybUgVlRg+MH1Kv0yaRcMR9VNujavf8aeLgHoJ+7gIlguhPgaTlJSYb2DfCm
VE8yVY1z7GLzhee2zPGSTwoGnSXkW/bo+y+BTAzZQ4UDwR9ukX9Pk5la3kiuNZC9tgYadpnhM1wC
O+pBDxxBFwq6J/ku3zv/vy8uAN8f7vwRGmT8xX9AOvf8rpb0aay3JL7HdZCbNNbp6BqIToub5ZAi
5cCoYgK0KSF+E+ci9vXlW5de1NaQtKv0vgUkiYkh6fT9FpYAc/6q7zcY9A+MfdOEVAgOpGtv/Qqx
zi/Kc9zcS1j7nA+LJjlPh/VFiVZ9i3rh+VkmpoT9us1emtuQHfdwAksPw2wmnELgOLZCzstXpnpi
3q8tifcROGrg/JQmNh2JV3x0ll2IWH4DOCWH7Px0A9m3HBgnCYJfAMPpxRFkJggLFVhJBwAM6VRE
lxz2tC/DxK8xeVHAJpg6QUpF91y05XQW4tbIFWMUEWJ7Ij0uiaAxahhNHh3lV89UC1DgHeBzvTwT
EapqF4nP1IFFPYKoNHsDV2GK168ZQiOcTwmg3tqa+tOkD8dRh8EfP+QJIIV153ypIJhvASQOJqJz
jdPvsIa/Ok81wh7gbId6QMzcbstiRx61jcH4LiDCcstBYKK1IREb0wafMQKb/zNolT15NKV7MXN4
uduoGJgzO90tSS95TU9f8rapFp87WwASoF4mcdVSds4JHE6Cw3Mr+iqD8R8egkjQefTTFoTpBqp2
N5XhgniQ0QhnYDEEHUaE+xbIHO7anACqtZ9Ob3MoluMm8TWt493zMx/yCpNUaaklRxyEtQIwTxrV
B6r8uffTRXsoHfUISqVpYDrpQR+gBonGcjs5vodzcAhEAMR+0jbvTfNGmwfDWL07W5MlOCS1HlEh
gKHTv9CEbqxHPUbDOQ5soOcEGXB9P2rZ6c/5JJMI+BAq8Xlco6uJAELvFeZvn5PW4E14xo3rp8b4
Xp3GeW+C48Z0IMvl5nsFSPT2uLzoNCLeWxPCiJtwcrv1aaHT3myDm5XoiAsdLLhXy8xbhAvH/E66
cblqyDksgnrgOOn4kxADlHfJADZXu+dtFJoc5ki1rKtTte3RXJaIlWlYU0XMwg7JyUyRM0CTDV6x
QKNljXGT4EPUbIys7fKkQBMg4sD2n3vkZ2MhPbh70qZ0nSQfa2TakLsnM1HEA26M0D/Ra3QC0CUn
MO100mL/TRUDrLZXkC9sOtVQFYe2GUwkMcKS2zPJfX1tEQMPNGVcxNoD5P+oetD5NG8o0ufBzFhx
8bGwjiGmgzGa8jEn0luR5h6SNAV7ApZWlnKD9SRWmySlJM1L7vBv/0//31DqqD99KqAshoE5Nhww
oDXKH/HAW+MUqRogadxdON1rDThDiYZDcCzl5S+oLDU7l0kUlvu+U8h2JJuDTNmh8sabVq1PjJKx
Zw33J3ecSnCjLy5Tt81ezwdAi58JgbPYyIWw4VNO2NcISf9a/dcZqF5GM5h93Crg+TXC8VdBZv6H
ijmApUTTI4avrVMqVyW+tVOMiHzMGLaKGEO0+YL0Rl+ywop9Nq2uoamzNGCtD9GELtb0DK4LAjuX
WzC1F1GkNjtXXKXQlZAgwlPAd1XgT9dgr/74m+7+r2LvZPpa5l2ws2q405n9ufHCqZzExinBkcgM
O2Trq93/O0OSG+3MdtcBpYVicF4UcyYjknOPQ9ugwItkuKECe6RoBPIeEip2DfOxMlZmmJB/ntej
ey2EtlyY2W/k8iUeyMEDJyJ8fWlWctT1pRQqItqvIUZQitD7HZcfhS5EXGfJHZUG/+wi5ErtOClr
t+lYAdNGekIB0cK5irIXapfyeC8xb5NZx0Rpyp/0S55QFmWR2lOVA48EKeKxhnqQp3a1SddKfbNu
ISCzoz2leROkXjNZrGaauBRpFH/4ig7x3aJ6YDUyqrj79WRz9rV5TM/oTypyGyr5Dat7+R4rumMx
gQEy9rZlXtBmCc/VSK1mvzrhE1OI5jInwwEez/Jvyu4EZKMF7XfwtUTud6hhka7TJAf/4hlmfoyN
urceVllJSDzYPygVmrzVs1nKc53t9pc4kuU/Bm7HGX+GOxyHjZZy7TB1L5TvNhP1uwj6zSi1PAwa
69PKEP682UuxYQRQGKYx1RYnQ+cc+ERdiw1Nr/lppDMOINtBsO2dyGsmz7hI5mJr0bxPXefDpQcz
6fu7T4e0ArSd0q5aeEScHN/YY+4bYffkQ/3qOfbjVPXB2CzgkqlA6KQjc9MIijXoGkSGi0XDrufi
Tw2eaRx5tKYnaFh51Nyl+uHnx3PnE3XpmyVo1Xwt4d4pWN6SLRRgIfDkiYCVb7gJFqXFoaBYlbBF
ijaY5NB+VSFOHvakmGW8BsPHphn9bJ4HRp6285gKnsaQtpYlQ6ddHpHJFhrKryFj6wtV3SMSNNdF
a53uaUZX2SuuF9e6n7/sB1Ycjc/K22M1CMqNE1o7jPNCqQL/hX10EaNHZUgm6SoQhzvEgL7Ah67X
UHxqzZiPeHiGy6ZMf2xIDcTJEFQByLTwxBH9u67iaZIQBm3CQhuXruBqxRlaYaZfClpJ28vEgKIe
ZI8WQRlUSD1kFdink/g/2023kcVRX9GN+77f9Ja2in2KTkD3SbxOzhgBZHA3Xt/9Ja+9N3z7bFUl
L18/cOYX1xAkhT7XjFTqDp6oGFN8q9vywSXJar713swlzW3dVDwaYSIeomzsiXm2RfLU3TBPl4wT
0lRO2wzzSuUWADSV2PFIkjqgC2l0kOo6lrGOYL9qCiYcpObKK+WO7M8V6nqn2PxX5YL781kL4fFk
R6iqJF+Lnoj3WKKOlo1DNaekSRkeA/6XbnccYzLF9JBxOf5wub/bR7yDDKgeGGRZ6VyZIMV9yYao
utPdYVxY9+3EZDF+Wq0I9Mgbd9ncOJn5nzqBYm2P3+JXeURh/MoYRwelaDnZiyD/9v2QkubrOEmz
O0PrYJZJqI89XFFNI3EI4P6z1fETz+B0m2OiNg8bkJbs8pA2hewrrOlGV46FSMz+Kxv0KlGKEA90
BhHj4hWuICa8thnYznbpq+MxdyGq0clATAEmTxjcIzZLn/VYKPYiDPCXkuaTSckY0nN8o/MzPXXu
Es3jt3c2RJmGm9WA8UygDPB9nGfdFxO0reINexiNrzSPGOA964auCdWUhF3kicngsuN8zz8PDuvm
nmGhZ996u6C01xhQXCkeADUVX4+msulqTWLpPX5mLf6CVg6TM8LzYhD5LGgwzsgXHf8gSWJhZgtR
BdCCy7zRrv9MAYC7wY5IwNe4Mcnfu+mGfjlnt03QPFKfkfnWHKWrVIm1pB/tSQNgFvmovb8L8D7T
CPf/qmRG5g5AZXxm61PTtNKlbjOwEgjKL4arFE8SBM+byobt91N+CkcEgELaStV0fMYSt+U+1e+O
PVn1G/ZUPik77o1xsYhMMJjJtPmOZa+BcIQEPIZN7d5W2s0O7W9v74nwMfoIyYPl1nqB0zvirpcy
3QCcDwsCE6LxYPNsm4SVbHEbxdjn6sYmB1GTylKuFLMEZhrTNXrJBe7w+WMwaGswZsk64vVFuSAp
l5bdriD23ZTdqvtojSokZa57CGuQOD59VWXogq/rBwRUlyOY7OHuhR9tVuozyOzWsRRYp34UjqMv
LPCAu97EJ7KuiS4emX7LuJ32aLXMAeKne2o5N/wsaEZrZewZc7tab3eUgxGkFJYwMUeHlcbxE5dN
A+goXsh7553jkW/4IiKqd4m4ITLP67HIVTzE9VqEIvKQNg6r2o5NR/v51UpMjO3QHp2ZKBpXvwsX
zUbw0L369BDcMXw6VlYkMmuDyq9XSRPyLx3RXPkTScgqaDDf2JmHO+dRx4hJxH6HcTaGsVdV60sj
bK0YPpwoDrcwOUebJYQ1Uu3RKjncf7lMm77kJAiFaEHSxK4j9NjY2yPpxPj+uGscNhETdiaxhQEE
TvN1pjTZTXLuHzw6dc8MPntTGs0vUewCTHcSJnDb2P2MmEMJ5STXbqJitSjSDe2fGxIhq+eqtMGO
eZANG17PK+MBmgmETi0CBOx3V6B+ncXdtQn1RD60gaD/SEIEQx2W7aJd3eW67gCLGyF8JBzl2s/7
9mysy5gicRInUO1JU+63q/3VRH+1YE5VDaEo5R67BoDnX9rj/7JCCIT5DGPpRTIchICBeg1frPrH
4TJCyjoZZzWRGCrwKlcPdA2sCYreKXzHPFn1E5MHnJrjD5Xcc8QVRMw7EwByAiG5IXjP28JSKrxx
QNBnANd7/hKUTlzlJm5om4O9qUAwrDiBZbL1wvLWRtOB2W2yJr9aJerIPAjI2BhhBuAB/DvG8TX5
f3WThy81jIHy6e/2MPJ37+bUlwaaQxbuu3Xtt8pIlWLuCiGuPQ7ucxuNfWc7BVP703X3XfnaN5qn
brjubUAvf7rKhIjNqE1KHo7KHmV7lpID0BlcrDK0uY3z3aaI481tGaU6iUmqIxHQYAoMAZS9kkz3
S6PVQph64Oykfc6sBEcC+kVt4Q3aDOycHcmJFMboa97/AVbnbARMwyRAckSMfnBHNd2of0WAU/xa
QxOmJN3I9K29Jtf1CUl6e0Am4fZu0IdfQm1iIiIgJ/K+owsn3hRLfzbiEB3ejJiVN8gS3212E5VV
qmyjLzEShj5QPtY+sFodQSueQo6VrNJirA+7k+2Tp5oN4znK9aHaJEaNUf5L92Kk+7TbOIk7aebz
3bknYUyj+d0eMaWr6Xx7eRJNUngijlUWbEQL/pwQ6TzlBSqzln0W9j5Rrag/+HtHSfeQiiG71GOj
+TXJQc8nJ5MoIm4lQcn4Y76IR14ul+dUY5aUF9/yFPfg1VDEig6XY/EKKsYSNXswLEBhomsFinsW
g7LCWfW+s1/4bIWstwAhffmP6a6MReATj7Hyx8NRz5UhRp7+zCOte0zi2Luy2UpGckdSNoqxTKcY
vVQeyBJRAUJO7R4mZ4U6CJDYV02ASngx27vOPEUNMyGqZz8pKH6hzHNMgmQzPe1XMDHRuQFNhCZP
EkCt6XL/sDU9utD2X4OAw3aYekctfKeuIEbRJEx4dNzxJMp68CpSwlQDdq3DPXSnZRsJZkUGGHMK
jy3g4DfuYRCN5ghu+eucfq/43hA4oJwDfZuCwXnX+ry3QLtD7NIDk8WnW35MLaC62JpDyLOlRJ4U
D7s1PCJLIifa2g4LSGvKf8uLSOLtgK1e79Z4eXqvrR7g51qlipjJAlHrtGt+T7CSn4elzWGRMzLe
HtEqbROmdM5bdNPqsXZcNHpS1/QmZg8xTI4bW81G77TTI9Y52QvIJHmO8PcRKcUlskJ/xxPKu2il
1qfrBzZQIEww1nS1PYe8uWqBZgu6/xVGOiHwTW9/xQlJA59slPHVeb4xZu2dMNgU9ftN+tAmqnRi
7Uo1Jr3C+CufkTs+8JRFGQcMA0eIQWK/C83629KNrB8y8TzvBVcJmJDe5DeWvdiZZIqUDzop7/kM
ZhKdYJJAhlh2RMSIZRe1X2+NANyIVatCMj+j/qUWYk2NJZAcBqWM58HvXKAbslyKw59FVcGExZGd
0N0MscadU+BezQq9gBAuSMudUMDtc681kDSZhZocrF7m5RrRRS6VWVSjlaQ+/D0DbeNHZTsB/+Zp
SR/WD/R9t7LdsBML4ND8ZI6/Nsxbu14LbpPi3JMoy1QOOE2ct4cw8nMEA1FmCrZm9bWEDJv1Rm51
z/WxuqeJHjARoD+imaoPLnRx2SeZluIJgNi9dxsvEpNjKr+grGnJWUySmWoNeYagx7mrBZFpzmMc
kc6zwtdE5FiiaIBQs7zQv1d9XbaNabk6fWZzINDsLjfdu4F+UukxUb5+WEKhWMDWj59+8Ytl55J+
qO7Fez1wohWcUGCyR15uDv85TX9YlwHM5YP5zvXzpVLIkn/IjfZuibSB6nL5MSamAOjRuxyLFrhu
fX1RE1h2G02ke0FFfjjcboGF7xdb/BmF/XQSrR/1WL2/DtTKmlfZn/ydawTcY9ICD+WIxVjW06nK
8M7gdPSt8Oc6f+UeH76tT4g/QfoF7gLg2pNoeHEQ8dgIhxrSVdsDBWIwTieikVLhpssltcNsJhaf
Yp9ZHgcTaFB/A19lzySlzooKSuLDq9J1SSF/nkILbotGLT4EN7CGJQPRU9evXUakLQ9LDQA0El0T
SIJRLdyY51MyBYFOAwK1Lemq6uswUsb7KNZYzcXUAdxPYq++VBv3j4TCiWxnBH44FjEFcufZRMMJ
V2EfB5roBOy3k95QCgLYHWcgJr8tWEAVVfqZpd0zVWtyiW7OUNOVf5O9AXpbv69rURbo2+eafCvx
fj1VJtIotNSKv9Yl/SXawBh7DwDyTfQGvVQngyz8RfxF33Xky9u1IHAXo/F47euhA2WbErde1Wmv
zD3BtFLaFfhrSIBIyzWkMfbLUX556vyHUt+ogCARtQMWZ3Cz/uTSN2BeHeZOEKXoVIV0RPy99EM/
MADc3AGSOxq+B1cDowZpCaszqTHUGBHxRQVqhF7O99icEb6657GXocaFVMMHegx7FI6ZrlUAeGid
DV+dt0amRwc9d9r+nNnXtoMW4ZvqYb/M69Tzf5pxeyb7JV4unO4PjGVbLbtUo+2yGkwh5OpLiAsq
udx8Mz1E6GlYAH9EYaOgXhaAdHiCQMs7i0yh4qcM7wbKtms/VosbfKlO1aIAHkaEBrYTRiu8srOU
R900modZ0/Tu8+7pOd+9qZpxYM7ezbhDDuKMgkfVvUVtJfzQWvOLsfsXLUsK/Jt23i1SNfgVRX0v
4iNBVLgARhq319Botwg1t7D1sdDrwknD1Ve6gfZwjOZWiL9Lrcq82/hVOg72OvhNlMwriN96T3ae
Btb5SI8PWRweEzAUAUjux/RC31Q+fwVIYgXsgEZH3+g8d/Ts7HocKheioWwVQ8/nwCXn1ksS7i5G
9Ohlkp1u7ZFTFwlgHPbY3fKftQR1019LrjF7BF5tUJoYjBxID7L6qKb5wt6zKr9chgH3byMnCoRO
kjVtY1qC41etl0ZoxXAFj7yHwo0teqAKRje3ooxxR3gSlzMD8nhVcKok679RV70koXzcgf4qojI5
3m68u/iUB4396VMzZmmmD89aDGZbe2ErjU/1mylFxraY1lH3bEH9bCiCFQzo9A3oOdKU2mF110iM
DegWqK8BZuQG3YPXOdoTJupKrBomBkzqE+XfSi/KNowD2dtKQfnV+dbtABmyYcFY7ghOvZ66ujZq
RuKZ5Y1UkSkLEmOk4koxkHKxaQRtMCW73F1ZvqvhoZ0icUfYGc2elpHvhHVM8vTTQlayDPavdt25
Xrg6qC7obGPmuUsMly7dTf5KZeOkrtZYzoCYDVCLjs0jpzlyjuSOSKZeXsqwpTAwVZSAoRAogLbc
4l1G8yqKK/hXxCo+pZkJEu+2hBeREra1hNtaMhzI+PWd9SAmN/BOptt4nPWY9UyWY/xFejEvUQin
VQX/KvExrjDVYpe3h44WQwcPt9gH8vjYHSStdeoDM410dukQBJWdz5RU4akfZUqOr7PmW7M7Vols
1mi8xOxo12kypEyknO7bkTCUqzGZVVsKvsg1HIn/dE0eKI5XEuHyDu2sIsZDwo4dZPSr8F+08ytG
MsecH/avbXSF9MuOTJVO9BDtF6QcKVhnVmtAkNPtCmPwTYj/A9ZWdvyXP17gwqVSsQij7NKf0iSE
mZzebzIs/dsZ5TNBikbHQopvJRUOCgxJDZ99S/13kCjWVNut038iYTxZ+Rx2YeDTyLVRDR/c8VU9
LbwDOhiAO+4C6Rbxj5fhQWxrk6/jC1yzJ4/sytLpr5+ID9WyI059EYkvxMbNObdaa6f2Qye18pvl
dXDvPBQugRDCkqSnl6DOHA/M2iTl5O2hxZ4kL1LRqpCW0BW/qI3LieDrI8VhaQTYSX5RcSChsIN9
ilPTE10VwFD7aNUHHy+dxxH8rvGbMAP2MLNKSlRX9LxlvX//RS2eoHREcRj4E/0aFQRRDAOtMysT
Thtf6PD8x1PvpoEw5pmkqVduPVHQfBsupTw7uuPCoYPIzLLlpLPwCN4n+ANoFlf6v///TK0RoGTb
tZURU9RcKhC0EReeEPTiHXdK0EV+pe3hwYaorWMTHb1FhO/IN97L7Q7oqm5XohQcvIoCrJ5ZxrVB
RPLTi0ReV2hC72lk1xYcI1+fjNLnRHvFDTz0zlYmEIK4wjkm+65lMzrjT/rHxkgMYSzEdOY8CYkh
ZmbtFXbSaPZ7G5EY+1h81Ck52qN0nw2IgO3hCWzPsHWQR3NF+rv1E3FkMmGus1HxPFVrOc2602X1
QoHywypRJFUWg1N1ioIQ/IYP3nXddSGljKxAxTAd8MRx4uzEHG2Q09dRdlphJ4FDXtBP0KRuTd3s
X3Pirno8wr+1TgbThxQmS2YD+5tG5fGmixWOuNBiuXj1U5PMz8gXDZncClrqkCVEUFQ38ix2t8QR
Cm+9M72cNe7jh/oTAJ8bj8EseqOPxuOKji6a2dhbD5/CBNp3AU+NazU5GVZZikFcC8qOF1nFyaca
V/dyeSFKnMLgMaDxozzlUwQ4cKjz5UQBQ6Qi/jGHZZ2NJxkVQvEv6FhB0sBTTFhEKaTvGhdqsRXs
5Lsg5cSSdvokgKZ/CmKnTqmOBDuyztgw7AFFPfs/H/KrENUTIU0oEGbkCXZp0a41vtE7P8vl3cHp
OifVuKuEiSIOuH6jpdKBDVVsa9yGgGHhTJzt+4Lt9U9PJaJvPFrQU2EWCc01LcKoW78scc57miES
MMoVaxgDQ5neg15q57RYMchXdMhKaJ+t42+vaFC4cU1yPj53eeX8bv7mvJfiJpCESmQzydOOquiJ
1p9ZdE+E1MuxN0RpD7niLYvNQ6s0cwVyxc1Yd4w1KfIoIB18NSwlEk5q6PZKtKCfX5AZNh97/jpB
m5FNIKL2qfmId3ldDy0HA9fTR8EEq4pFIYZVbQJBZR5D+qQG5h3UGZtVm3po3edRLthNWaJlg16T
LsMqfGf5i3iev4WE4JXSpAIpu4xsFbvGXDuLOSpfirJPsfBTtJLk25emvUkfr79chnopUrPzKZZV
BeOY20BG1NHL7dsCddSPw8AvEHO3x2Fs5WcKyCu782OOfDb4mqekLGFfxCWp51TsuxhmPHrBaoCY
aooA78/UL9ozpnzlQvRsWMsQm5VZ1btdLD6LO8BYB0zIVbRkHnkEAUIOhdAO7/ok+tGVIM+xybn7
ULMhx2gVHLkTylekYYlvLDYEHSV91Kfas2dkGeTOP6okvqHfSz+br+g72MRRFewIhhaCym7LTyff
Y1UnMeicsDkSUwxw+z8cJr0VM0j7nYKluBBoX1EzcWBQ+jSXT5oejMJLqTUvfXpahh2j7BasC5yx
zPkc+kUkC+BuFLCKtJ5U4XsVG85inbsvNg2N6mL900e5CM7Ke6sHjJ952Ko8xSRoKs4MheZHAxAk
R/DYTq6WqPEaso3DWU9zCHCicggOnGY80yNCnordlImCpPBAonNveyMdTHupY6TEW2RlAMk9JwKm
cRNhWvfnOFIN6kxKrk3MnwPXbas95lcEmvvkoz0AkPTKybRY4zDnpotxxCk3h44ZQF/lERzYIROV
A1j5ZS6qNwKlstl94bVXaFOh6F9za6QuX5xrvg8KfIqNkaT5AQbcxH5umDfLnPHX1ZHNuhPIz4ax
QFmrAjxqnIOVOLyqiuhvahPd0Cp0FkzIKs1aNCFE9D7QTdGSgC3u3Yh2DqeLP+VDaWxbzy0q7oYO
WCmuOsUF4P1WNbmBdxkxQQmDmotlnBi83T/ivtX/jEQd04s/AxsSgLjJkxQGUDEDU2sIbmZ2Pj8X
6wSCmgCE5fx2fPXVETfv5nAybPqiTv1nmjXgFcGQiGvK/nbcrXm4DuHtaAC0JscNZIhLjYn1I8HU
tF4+LhDgn0Num1emmUHRu5n3Pgk/JpaEtocAUjx0INA2SdHk52/BPUSejXoKTVf5mCIt7b6XW1B3
X/zxQjJf8/Vx9Oyfw6otyPjtc2JTTwtErCUbemaXh0+iQr3kPD4zS0m9Un79m2bC8tHNLTDdx7K9
slujQcbARe6UtjtkiMKPq1+ijGe2Jq8qu4JktaASOQgCUIplKLa+7RMgHObXxre1+RHySTjkwBvL
Y1LyYsfdmPvTnWtCAaK33rQi8szhbQqNfOzu7+L/rkHb+1+CtRrGugMQZr8KGCCyX1Au5LptSn7b
mefcGQShtHt/FfB3SSCu3uCXYqj9fLAfLrympbnSwRxA4Sj7uv4RKBKJO81phDCt54fvl3P9BelQ
4HMlgxeenaWnAPPHOj6wu6a5bFp/gn5WUz2sJoZUMM3wO8lXqNThGeSvbgYE1hbmevwroS/2BP72
V4y++3SdN6qVVQqWTFs559YNiBBV6h+a+/ffwtwABX1EL0Bo8pu6JRCaipCrbAGgbhLPyqDjAUWk
att9Cq2I/+47z2fze/6hLGckGmmHoie6/WjLdHMwvTeb5Tf/xZm1+uApuZfqCecQI8OLDKFWt3IY
72z4oZyBDAwSyg9Vpah1k9PLcLudOxhJjRrhHnw5HfKL6WAVIk94zvW8LIhPuGRe1NLR4WwuUOGT
Xij09hZqfAsPJ1SWrnc2TyxTHF6NXaAE1NG//1LaiObCZ7wAw+m+vIuL3LyBJA0Ufc6RQO6d/RiS
7lJ62ER3e9wOrz+BK2U0lmW3gzfp2f0JEsLQ+72V1x3wfY+f/pImDINIdKzjl84DcfODbxO5lNkp
QlglKIvJSrkh2NBENpT2K8TA9F6EBCDU0OmH/5/sbztfwIY9fOoCoHFi/DzNeEObCxPKukc1xNv0
u9kvaN7nyFE+vRyHQJnodJd+27t7IOKBUipJMnUTKg9Xqz8v4DraoER8uc/jGlGkI6TnutUTM2fp
kHvp3ZmZCb+Es3j69EqVbh3PbphevmnC6ImTWzWxZ1QrlTiZIvevAIjHJ982mteUVsReuQYotX6/
MoamcQOFRTmwOOV30W9pPKboE307Fj6Tpj0v9tFCj6dfQSyFTjLETEjktJFyvtyQfs41+fXTWOl8
G2645RSQRwC3+/BZaILaKJHUEW4x2M945HaJ2atYxHt9QiJsSvyK/Wu3+CpfDr5oa8VNqXBos2qb
l/7UznxTin6GS/2CvwR87AiuCGY0b3D1qyjrckHIPVhmBFpWlASsDSvvChYp908C1d7AMkln23lI
f/9oPvediJEZPOqJH5O8FIX9YXprT+bWk9WYvsVAZGA4UKs4YuadaNXRc6/TFfYVIS+nqkH+eHbN
3vtYTKyAcByEjn0qglKqz9lJRrNOnWVGjAus1xkbeFtNrpqEZUSmE+dQT74hWFIMgmzvwxVJiv20
9qoIXxxeHIqAgBerAOThJZn7skiy6ChaxLj8TjyaYZnX8tZp9qIjlXUIY8VRiNeefvBERY2m3yYB
R6zY3uuoQk/FFUPO3Fo04NWESyCDL1UhzqXnu299P4Jc5/vo0FA3xFmiJ46VZtOmxP4ig4BVPgFQ
5VTolYcsW6Rwm/OIhUA3qaD8SSXT2bNYN0M5D1t5QX5WLkAiwVDDCRQszxXMHIE0nlnOe1CVLKgy
sAszHOdtk1ZQOdthn7Zo18EjlR+6JRRR818vAdjY1ihM7Mq1cVMbICDdtbozFzKHO9abNDKxW1MI
d1vGY8+L/X62IqVBsoGjlYUjMXpPTEIkv8JokxgKZfZ1uDKtzUyd67vjryPz1zSRRvk57c+EZbNy
18Qy5Ro6IKFxxc85KvqfOJd9UYLS9f0PzVvqR+ghqqph7cRJOAOFSyqj/U3fW7ufRe1evdEntTNx
kwywk+YaKb3OplpKQbUrAO1/UyEdnIGkjYxxk95RkzWYna30h08ekP03bZCZdNB2hMm58jkh/z0e
Ztln6eHZSkDlcJQD2t7bNDaYw2Jm8E9B32G1UpDQqehOBcAjj7kTq/6e5y2qshGL9CjVb+mlEXqH
ltBhyNP4y2FQZnjmK4DTNRb8KYZtPqCtE52s3rVqOndmXBilcONtfBsS5V4OKz1XDcdwzfXmtsnz
bJTgWzaPJO1Za5rCs2Xr1KD9LeBvdqloBPlCrp/fXBUedvxk0HijVrgkVy2ysf8wjDEknvOkkyVr
+be/i7JE3KjwRHRmIVqoo+5582zQUg+bp70+mKodIGxLPerJWJcNHfSMCntzyirSVkyqT939zOnG
B32+1CkzKGF1iUj7DV5ejEYTXunJRckyrvRcIwMlmAzBbATSLF9KPR+Ig4+126yQAMKAHEXFRpos
MFcQjVw4FstU2gNZnyGLW+pt6Y3cB74uPU205m8r+O51XHnTnZcU0i6Aw6RE2cPsU6OE8/baDxVk
DjRFb8J3SiQsjq/4YUP0V+oNsAGBe9rfGi2EOn/VXrHGgp5TlqDC7RPlFB418ZQSC5bSA8W4sKg1
ilsnFqpwCrOY/xxX7/MjyerJNre03ha8fLz4Kp8sA6L+l3RhinAwlNM2D+lRB1t6Lv2bugqTVnXe
70H1KxLKHlApj03X4TusLR17z6eqR9z2l3t6J/8+J2G+SsKZfzkxaGwcvNC+I6Zurd7Ni0JKp+ej
C270V6zNzxe4NIa/koyrXv+jFxSobqxkYfcJBCHijqipjEpKHUdh3edEZyKIyle6NoolzvgGC1F+
fZ4AmIpjRs0p9dND1i4570Kfllu0VnVKIgzYBfC2hrpEHSgL03IGQjuKk5GASPyFSMz2e7xbt0i9
qGQpw3aKwJcceKBjw060PIcitVhnWRw3VZxvV0djAMWk+qBeeA5gcBr6DNrz844xOrLFjIu0ZCs/
oLC/Nnjz5Wx1EqSdwAJJIiElgevRnKEjG0hB/5THMiglzoIDGZ0X8sC7fT8XTwwKWazgMiu+vfPb
d32Bfk6np5ksDtNMOznSHQQzu8u1c3qTIHp8yrrImE6t8ohom/2QOsWSEHflqwHlOezcEs6zO+R4
yyi5mSDT9BM4AYwB6mUitADiu5Z0T6yyaAx0QKEkkuYgsJ635D3AKJeXG1SPwDar75PM58QvgZV9
iddjPEwT1qw7hhuelx1spWgpAFAIHF8L2ejU9AEScDwE/qUIslxms1t3cheWz8BNQNf1LzlNdsTa
zKs5AaVldtr/q7k7NAE8BUcYrYa1KX5vGIja8EjbAJUz/KfY6TDPe9llxIfvM4HIo9XjDIN9p2L/
L9A8j4RzExRjOxkxmAYOhxs3P/8qWh02Pm+CRTxD0VKhEN0QSn4UKjYtILOZI26CcWMkM019PB2H
twqFesWsfkByRopSmFikdbEwJihY06UlartMoGq+HffG3NLaxcvxGHu1o8FJy40RWtJl+nG2/eNK
2IimDCsYRVW1DChx2f7HSYQj1p5FIhYzCifVFTHszbVlfQt+QcPywXVQV6sCq37QJNihjC27qjs0
K8TQVPHOj7nqis0ruFTs49qPfiOK9wutDEUkmAZwlfSYyt8bTaZ3SXkJcv9q7fyHl9l0k3sIIVAz
W8rcz3Gu3DoIMwl178+jv80TNTRTDWgkLTPsOQB8BiBy5SiIdm5ltcF2yE5jOMTsMmWfjJUFCCAE
iUT88XuTGKWDv+bj41i8a5hC+dhhqAo8MJdKZM50miQ2MORxDBcjdBKuZ2flTvMMXlcQRjnTLBcR
WZLOQhHVqcCMDqJmMo9iYtcOggkOwpXCeTzMLA8YNZ3CLct1i3eaZfxTQr7rDfaQOIw8TvcNW76Q
bDLocAY54e7/Sm7VNX5t6/IRnORAxv7wDPudDVUkj198R78K/4jeDZXrr0IFUlLdjkBdo7L5Ta9H
61moLJk9KBwwil0AP+8Qvew5BKX7uG09EC+VR+LpPjYdQjZiAE/hTe/KxNzIKO4xUFXwKPckplfv
vN/EVwLKSjlPbOibiPL5sU59Agkz7hUSbflJBBwUDQixoYQumv9TRldJjOe0o/RhXrZ7bCGUIud3
BXQfSdE6M1sI+4HdgXCsmdCt+U8eQIKyKoDKJOwRWAfPdzIm8zZ8PH7sVtmR++pmpXPmxnusMXvX
Y1jgIKTDuW1A/hzufK60Jd9Hza0ffcaDRQF9JoIgl9oqOemPJkYH7XLNe+LvQNTRgxEjV6fEkisb
bEBTS7xDrzkhcasdu+1mv6jMxz0AG62rNDNkiJFgwxAWZuQKwW3CKZuJO/XCbaO+2i2HpzUHaLBN
8ndjBsUubwkjbelc6tUVLgWmDmZ2yywjExBnb3H8Pc/6yy2BZwjLXZnW+gkmKyFTD1WzFgUBfh36
7Ioxawu2NrywsKB00ys27OOmDCMUw49W0brMY+ND1MH3yT9HizLkc2WdSvNrbBCajAGAwZuGcU57
ZVAGxjEn4MGfZfqBKKIlEJMP7nI5sITOHRnW0SrV4y0DZD2bV+52TQQX402oVwzbckLw1FpfSIId
WbfGIdyGJZXlKRbT+lY9t2AojbBizx+WH5jXfHyo+VQ70fSG7PxpByIekhzxogDWg9IZm0+7pFhU
ihVZrfVExa8YUTUsDuA3yLgvoQlczVpQ9ZzuzdFPfhRRaztzKJuengfJBOe6YHpjgAx7ua9CT39V
+9/tIcUySZ+kx9tNWhzmliavZg9qmBFXyBy0qDi4PDzrDbwQdg2um3faHYpUANJovCK94/gawvUw
yjNaHii0awdBDBOPCmtH+G+6/bsXTcx1Zg+erSWwmVY5s0x57G1d7VpiF+gIAIZygOI8oGV1PF63
vTzWcjbE0mzA7WRW0FmHtEbocrtnabFSP1EcrDYWVq0v5DpEa4/Opo/J6PhiEP0jGCN9kqaHzqsS
0Cr7M21BRMUAAexn0hBaDfYCWE0h3C8B/ccRxVRwBy9C/fBpvQD+9tofP59L2xjVeJDKC/5DIVan
qUADWktaBCBVgCq/hMOxbUN+TF8MRLbX5FipaBe6o46qQgTeqPlACts6V2P+BTxQ7pZuiVum//nc
tlwxubHtB63edCwPhIG9xt4HwXbJtYWHiPsLuvyG6cyrobahf8FF3HqVfPgUH4fA9q62nyd6a+x9
ThxAsTC6riCvsOuklahrX+dzDwuMGsuoYN7hfrTjh+JfOThL9t2kX8jlwq48sCuTZuTld+xrLGMk
RxvBMUw4twD0amCh3N1B6S3KnYLPwBGvipuJCDF6h05AjtvAS6FAdyG3W5CDfjE9d8mf38jHOKsW
UyzH82iYGDjRgSVvOSTzVCHLGp9FWPk5gvKcf6mTqF7s1olJW16gnpKCBYJ6j59V1vbF7VYjc1NC
NJvQDJvwDe2xj0N0k+fIAeoKimsCvNIoDfkMi/qUJvIXkNy5nXzYo+hnbNL6hPhL2PTv+NxCmAwa
LIWu6IoOuJ3+gMaY9Ob12yjPca1A4Byr5g6YomPa/R3pBLVurKVpVDewEGKmCL+VifZKf0dpSz70
mRJyE7m0BALJ0Dnxk0qRpZuWBZUP4NMegPKxYTtUbS56dzfA2aqllSWn9bkalHzwwLewGNcobmmx
K73vV585x+U7ORbPSOTDrmcnfAdh9o4t5GP9SLpm8C4P9cmhl5I6RtlHnJION15Z+2/+D4SYdFz4
uLI5Zw48Dq01fh5E0PZYIOuM148ZdvRtzxq+SjRWm+bmgKLLeaJ08sVuOH5JgcoXkO+drpiKd3iI
FCWfUajhP98Rn+NZZ0nnTZwBRPhdPWsYM8YOabsjt+/DsX7+rpjsYrOdQZ+m3NXGFIiXFWgIMboS
ZrFg7fnRfZIlDGjkPtt5gqVugdHVXAcGUr10fbh03cpbx4bjbYDEn+UkIQ8HeHkUAq5YXKcfyxrg
FDr0FADjM1ILX9P7v/Fi7dCu2ipMd4JUy6bdzT2a/LGlAeQnvog7I3CmfPTr4vL4YFy20qkfc3H1
OgR5Y/Uj+LqeYRMUl54ikEyG+IrrcXUlIVvqvQQ5+gpiLLQcXrhss9rW4thaCXOH11TPqQ9H9JyG
pK5X9zG4U0sGiddcEvGMes/3UEE5aX9gfZRLtuY6cyHdO9Fk298tmzSyspMax/uYFTvlbFG2PwBO
h3azZ/R2g8bZ0YIKQRE5BAtzoG6v0Y2/J2id9yx+w5wpvjGxNc7IHcqLymQ4dgq0rjdNpuYNPioT
PbloNITaUdrOL89OAOwwKwU/o2XO+UbxZirdf4JdVKGfuBP7CjOgGHu4rjPqhrVpOYwvUzGSUg8S
/tioUeyGWFQuluhkFy2EgDaDFt42aeNHALY7aWY1b5um9aIUjMjukq3IH1hbRbEaP3Tey3GTDrHl
wJjfqYyEA93kjVC4dxSRfDwqsD7ikEcpPENerpESnPsXZS18I6gdVGBXIFaxzKb01KyYSnmUaoON
K1W4sd/3nvVdzWZuwky054Jdlk0YCtPmxme8ItpE7xzHK6RzCrDxelVOC4bQa1SH/2D6V4DNAp+F
uL7f+Wnrv/Thc5Vr5PpVy5+4jZOAWRMX78i3YPzhtX4z+3X7Dv+3zJQg/ap8WQwEKbbdurVYxvY/
bI3z0Mky4SQKmnGyXHCxNafK85tZiawO/+5s1Itd59cdB+HQkssgm/audiom0P15/e9+UGlRa6DT
kEUFqYPkoW/DA7m+oUoQSMh6wHR9XBVnk2fOTtx+DmMYW3/d83IILufxk8quqfpiPceC9K7/XAwQ
IIOcIQJV2Ho3C+5uaHBXoOB0DvnTYFoqPMmVElUmOakVZTH1XQ+Xy4H4/yZ9moI1cQ8mzD4pa92m
m8bW+zENGORd5Trja8MJdDR2ZKcLCbT4s85YnTynfunSGoWrTJOo+Urgs02/vgebf47mJcHg2uMR
9jw/VcxALzSvAl/OqCr7kVj7EN7aZZXWRSMAMc6ollZms9zoHFV8BNSaIMlT7FBmSeqcPseXBIoH
pmjcEvkA19Ax0mHrPWRKy2RfLneq02JefXFzOczuyVFVksnwg7kVEkOZtGRJEydWtJ3d4L4kx27/
EEdCvsLKHYPWSA0Eva3m+8eTlc7JldkYSw1pDwwzjhK3hL4LTYbXRDqegkiM/Yr51zDBlPQU+AwE
CrPWqW0cLqPuJmRXI83ADF7QrPfaQhxSHB7aGUgF1rjsDrcKF+/sr2faaIKkjkGd5+t2Xd2Ms0cG
V+qPNbwnf5x2Q7du9y+q5mlxPTrJaherCEGKy30Oplmta+NgNB5PbFZeilhfledS6kOLgDn5BpqR
eKAuQMkyBzi3LHJcKwJWW3UjJxP2blH+NxfrjlXJDXprj1ZGSH6HsLulNW89hQ15+LAAdbPiufLw
hw+ycZMUyWOeF4DlTdNpG2DiPAvGKOdpXYwXcaA83Q94GS7aGvPZyVMajvGd8np69JWmuJGO/Fo4
YCARZZmXe4Pvg62VJgxOy76VQrXMAD47SlzRjpDtswxjwnX9MgmUuqJeaMdcNkQeLiOuVvKrFpaU
2AaU2tadNBTbOD1nI6sVfb/joSX3PxD0CgNb/sbOqXwmOB87Zndqu79Z7t8TW4RGk/n1EJmOQTvT
NimcF5W7PnNVLRiK0IcMyT8hcHCsEJx87bYd3/XISzYMErB9HFv6ntKmnPF/VnxDclAgm3c0EspO
7m6h4m9tqeP/nvDqrR2lmE2WC85Tle1ob4YUf/sYRTqmgiGK6vPKhw6bDlL2iOlR7dptHi7QVYsX
2oEEhKckt9WgluCOjSd9Ni2dC5M6NvkRPeLxcgHfvmMWq6HXLabzCwvEyKJSpFL4jgpWLCLpe6wj
X1R3PbLo7MX9/H4vr4XWm01gFRi8Rdo3/6URLz/tqUo26yzUBQNHsVOXk9ZNpMcOUrlYCTvkAMCU
QeqBVkij2tLqr2UyW2KHCzSfdHTUd9WIjdIXa4N1rhi+8wDr6oIFj8VsPBJa+/WxLrg+Oo1FQcmH
raUjoBm1vkbp+7eYyl4xqEjEL+VVMCwE69KS/Xd6bQD/954Yfgx412I6ovXBoXfpjB+hcq/kgV10
ghq285FGIYKyI5A/W14QIeYRmfeT3neIFIH8j0z9E06IFXVEQBkC42sPi1vi5mMS0pBqRHY8uKiN
msL02I/oB7CLglc6/mQCxUMMe7KNRa3H7G0yEPW8vv5IdKd1gxKO9LbQPosJGozvKihiF0NrbsnZ
0qTwC5aicT/uHHzSVNC4s50yrPFYaG3CXgtgWoZv9Gx4vJfvNNY6GhzP2yPS4Mru9CRRpIl8olog
6TxIHKeJsII0tyyFNU/Mbm8uFWiFA6qwwgsyu6p6rxXnLlHmJqOQeM3H6FPl0+XHwPv8p0lehilp
bH+4VjAOh+onAFIKk0quTOtmGTRGkFJct54ZzV4KOtv7HFSJyEoFHzIQ+9QvWbOgCpnJ3W+0W/zw
vssi1Fqg/v9/vnjq+z4WeUBAaJxsSdVco1cHuuWj/f+0drNQPC1HfBL3SWJU433+g77ayqozSicy
b+ExPRNVgGILcGmPSo5Wk1FeKumOENkCrW8/+2hBVVx4WVRMzDtT9KYqIdQboTpvhzehEbT/u0VA
Pr/wCygZXE+oEoEbWr/l3fUfI53M3EGYKGC0ayVj48P863nrx2h6i06oHyZf2oWaj40xSmKD9F6g
u+Yz19N1Kbtmoc507fwh/aD9plu6h72reWLdsZuTWq6IGd4bSSpKis4+BtT0IkepBtQ7GQ0Miaun
LqnKvfJL8Wla3xRNnay7KLfiTSfnRU0IfOGWv5uVhB2bAxw9wX0UVeEmUdqmcH6bwknn/WRB4io4
Iz29VSXsJ+Ge2+aXWa54vWLuzM8JNYvfvT5sv2JO46cQ6FHAFbSUqe3C8W4iNVjXa243a5TJSXPY
gNXeQoZAGBIBU6j6BhQp+gObwPls7s/J40Z7S4P3X4sEUacFxPj6ZSMm6zZY/Yipvo5FIMIbUCnl
+P4wELNPTM38ojcoKt9LUXC2tI+n60ZBc8kxRYtil6taqzxZU7PPWLDoGetkedn7jmfbvT6ujNMA
M1e26BUbtxVSg7MjCObGrvnz5NL8klp2HsGMAcD8BPh0xEiTKev90+82K1riaONf34bYfCpLd1qw
5E4ZD5xdnVjpB41X0udMSdsFqw/z/wcpb+12bN7o56svubCpd5lPiXkV795mYYZV2fJJ3UP8PN4h
j2My5z2U/GEVUmWPDHqFk3zG0COa5jHRMwieqkYvfJK0HbvehXkXITF9ut1x1y9DnF9HDixej6ZX
qYBsKhxuM9IuzpdEQ3nCsZIWhqiDYlIAjoHvzRBoua2j5PS1uZK9QmaZVFzP6JHNiS1ID19RcjkB
8AcCo8Y+9xoTjzu/d5p4xiQlzI7JbgOXnr7A5vvKVsov6FsY5SryFIxWY1QycJ/OjDDX8tCUuu2M
HPcWYQnaaupiOmO/4/kYn9hNif8+NuiOZuYaJGM1wzAVZxMNvai4kWRwwLPWFyM/NoGsIIzz/i1r
uj/rVY62V9p7vPBF150/opgrZNVCAyXOxBU4mx+vshopqTDf8WHu4KFabFvvoV4oJ52sb8YU+z3n
3v/ieNwxbmfh+gnpQthJOn3on0IWwJ8GIfqFdAO6LCr2FEL2V6SB2n+btJbtVVwdQo0iFAb1yT/T
w33x7Sqvu6m6FmHTeueptxDJt/nflODGDOtlSQ2NKdVXtkhQ+eKu7vZMEE7k3pVA/Vij5rrNZxzX
qozpOv9/KBs1nUVQi9E73Psdsj9609C4Led0Sdxim3XIjf5M9Ltr/C6aDe22CE++B6McmVYG2kTj
CakX0dNs+3zADdBpWVQxEVne6z5Dfk8vfsUa0skJYdBYaAtB4x7yVjYERMBJ/sWXxNass1xMHAmm
PqYs5zecGFURH/E4TrZfyftfPpNaIvFFxBDdwXuluQXPnuexiWuFw1LvkK4RLfNAh/lOJL/M1wmm
0a/mi5+c8yprsJdYUaHY/4biyIpKSsyZvHTd7TYP9iZY0xV7JbUxQNkL32c745WsCtYWEugwxibT
0e/YPN8sGkVrhz5WwdlxZOZ+8WNGi2xCTjO2R/XvAaDY8e8bL5iH7YAaHXJs5aOoAeN7MDN+Q7at
9R4bP1MqjPAaJTrIbTs/afe0yJza9fqQ/XNqigMw4aUWaWqDux+rUuS6rmK2jAZvsGoRTV30hK//
QLeFOgxpAKW7lgIPbVr09AY3av0g1wYMfmfGzdG+dMb2eQ7XuKiCsNw70OSrxwm36CHa/cAj8uoF
kaS/kpByUTV2ayxXEoRToemBaoZBR4TwGU8u+qj3mZh7VTFBnx6p5GaAPJhnMNQFt4824+0d1evv
4ygPuakyX6y6tmclJZSSRsiXtn7nHLQgsMGwjzqkXEI2dtYCgXrEapGlO6nEiGqa8L/cqK8ecV1b
vD1FDVAhbLJWPYJt+QWy9rvbcRQ2fzyRygBpRU7Y4p0fCwBu3C5pqZf0LVHec7blGwrq0ssB1Clp
3CblnTgH3ysGwSf+7RPJx+AiPNuwnEouX1D/W7AxXqX6a53qpQE4IfD3TM9aNKRj6pQ+YA961jLk
9iLWP4w6UDGYIQ/R/WICUDf0+9sKqdVaefUyJKI+I1kbolqS67ol9PsTDcmv9tMosR/wZ823kmdp
CFOXdYSmTLLY4jbVp8tiF41O7i9NZOgfyBNik6fXw2ICs9U/EvynlTUWNphzuOmIG1DftD2impe5
24zZxxLN+5hKHYGfZK8LJOlwJv5hbDWJx/nC70nHTjSgsGv7rgBjDHVHTJCtMypVhi0NPthICRaF
82sq5KN4UPUgV3Vcod4pGmVRkGZNc+GW9K+ce16kOc1asFA9s3MkGn4GlZJ+jQbELwWD39zoIS+h
7NbJmaXS8ELWqPYo4DuK3ZufvAeNwpRgUN6mEikFFTPspfxLVl/j6/WrThAgHB8ZJKLVt+p3UgpC
ODNBB42X2e4lBTKj7Ic55Rskj1tJieAYPcBCqVqpoQLSXrnMKcpuW4s+GFjLU2XHx5Kq61MbdFUT
k+NuYlyf1J9FgjCpcK1WQOZOo7yuZ3Zqd/YUutFBh+rvJ0z00Y6PV5wvencV3WkVdO3tAwvM8Yem
5hkFeleM37ygyvgvlrqLSkG3F6i9wypC9vCgghot3Mzp7AKflEO+R/mgdAJI5inw+T7i9MP9Ldt9
mJDmbWnvVDAlzkgv3/O7TC4+Bh7eekXUMHsAewByLjou0qlK/8GwvLxvWj8drX+NQQ88M3Aua8Oy
C76yTyMh25ts74g5wm+hXpO9hJrRKnAPWMxGbwjIPYjm3uMkKC+0fAFcCX8GvLVQ33irBKN1EYkF
7aRfG/gf0LcSWg3vYGDtiuKvnKH2fb9dXA8JsCvWO9esF5EqrFSqs5fGOAGoMY3nZHjfjXlqggMD
/W4TTAcrQHe3/UtCx1yZHWbKyQiz2Gp14Wgk776EL3FOr6b4qps4hsEdQ0xZgtcwyTIO2tj1HXd/
r/g9/KWX4T1IRolQOLdIvq/HIAeQECmJgTtqHkVmLc41KjofdTv2cr7xgFwtt2krpG4JErFR8jbM
DCLWnkfAKEYIkH03kivGQBIFmxaOkVSj+gsAaAYkGC8QEhG53abwFN4Bw0EsvJCXqwJlXnkpAC0u
vGW6BdzcZPlefRyS7mIP+hZFfNzH8/B+qA9hm4XnUOgt6qy/diE7d6oaKBMTpwK4TwZPA1OjLOon
lwotVkeP8aHsBJmxbphxFSNcH6WVoAxcKn7k9uWXzRWevqBM/DNG63s6dWQv24m51wGL5n2DEkhV
BKtr2Bs5zqW5rAoDkJSxOsrBDGojpaycOc9v+wRFzWtsLI5nCaYEf/64N1/oikDTnBnePxEVKmLm
eG/VlP+xJrd/zWBMNV67ziprN/Vl5qnSGgUvYWrPfeqyriGg4Wj7iXP3nikt9LXoCcDOZ9D5KC1T
R5LLsMLMKVgILuHMLXD62nmIQnXsAiKvImoF153t7GZK4qz40uSyV9Y32LHF7XGZrwqEqyjfAtyq
CGA79RYUSwTOR2W+aVep1OT36l2Az3IjtxDLoWgXHg+6E/bWnyvxJzWZdCMur8fZlPXT5aOklOo7
A64sWdgZJ+TX3xMZ9JQf2rEC05/S7hS+NmYE21KnEqwZBf0QLnMlO0UM7fAQgEZSi2Zpy2FBfBw2
zNPqPnvloiQcNlyyMxrIpSIVKjJ0QbRQnQNvel9v6jnE++sI8WvzJ7+bcg+/JdU9PzVqZI3DslhR
00wNaTr31dDo2VAGwat3BwRB/8Frc3T466FaemYXKlJMr8Za0d8m1CGTwnxv/RTb9znhUfZS0X8Z
mSEZvAZHQhWf5ySKiCjq+JNiewwaBgnAwr4JEE+Zqtz1pHjNki7fDLgxlVMhhRiNI12xKsPqjpZf
XqPyWqVl8hUwSWW6lNGLOPPZ++FJc/gTwZ+E+6wdNOQsJmqMAJedCC0f/sfuFCTUZ+GBevRBy2OE
81p9vaYRKbMNfaL7TOgP76lJf4JhpTKlV7ASUvGbc3LJfXSt6UD+dBFPKx3rr3d5BfKv4pw59l+N
gwMUmpJq0XvflEdJ7x5PTaKz2kh9qOUdRMe1TuRJPrXDPngOupytD7iDVGmNpWvuvAqexenkQBMN
Mn/5Qs5bpXhOu6qVtBxSpbWeRad86/ZaP8zl4pR60oJVit8bZK35p9Wn1xM1hjmI204A1w4+rRSu
o9chHYmvaX8xtSSlMBXDfezsYdNhPxDuVZtkuCC7ONN3amv1q7cLQc2897lsmHYRToVIa8Nqrkvj
vzJR0haAuZXVnAQMavtIg5ub9LXH+IFTcNzyLupRE2FMZa+UzGuzuIQRPNLQEan0bq7YwuwVN9iJ
AH5rbwf6PPBsG4g3yjh3EktPw0sUJU6XjurmuVTYj4rYT4t9G9+YNbrV7taiweheis7khbMUJzs7
R6ZHwLNhdmNhiT+gs948ByidRAbX4/sB2+HfysffxeQRQrNfjpnN8XOkWHNk3NKNIzyITq44ZIqY
8w9GkxbqilvZRgPRxydNehy+aYS7Oz/jP+0j9+JttPm1xTCnoqvnaf0kzrIZbQOm5eKEJ8LqImdC
f2Y/aAq6T5q7dURWN3t99vuIlzoFbAHtzrPFqO9ujufPV63zJypyrKvBD2S+4W8nFvtmQ2rm6Kdf
wUNgd40HueBFHoGlNkh0eHNpVDz9YvEwh4bHm8K/8GZ3T3sSMYFP9Dc/QukHyZruFtlDmW54GCS9
ffDb0ofyHO0G3hQHVZclrczddO+4gr8t01htz0QfRL7duU+PP+vQEM2lyazZROkRztBDMugp/mki
+GyA1t9MLhhjk8yHmGGMxGPgNQXK7DrpbbG/V8q2V2oifUyaevr0j5iGd5D831FswP4n1ZZGIoJL
pVs3JLjBd9+Ss++XUr/CZxwLgzleMoYXgOFr0dqT8ZCohH8ikpYnnDEBCZj47TFUg4OM3cHIRRh2
iZzpcsFYyju0I9hdboOgOO+ea/M/kdGfzfWlwDA3V0R1ZZQPVfvgrolRB6XNzUIhozWtlUEW4HGq
EnbAWd2Ya6uLCVDp1Ps7w8UZTS4VYHB1qxoZYRfdv4XcQ6l0QQ44OIAIXFHJOAMKhDyG1XqsgtiC
S45KwK0NLXNKG9wbmy+xh7hnd/gxsCOYG9M08UAnWR+B39Ss59HnGcuTgV2+62i61STQBwFjPx5H
xvMWN+j2OmELvSxgDMH6uxngczbm4DrBCXnla8OTaVMyIGRjYh72Nst39UwPG2K0o6YSFkwlnLIA
/LI4W2j3tiMjLw+naNjPovIfZ6rfdSA5nK2yvz33BTOkfRfvFcpMqb+3nG5VtkpjNu9u7wnaNl2E
iYAvQtlbUq4olPI8/uqIx48gV63An8WJ//Z3E84FpRMJ2zovYn6zHQBtBMIGcq4/SLlNKF2BHzyd
kgguetZ5lIN5MPWG+iyqP5wrZuDv+OUDtUPQ4enV0QGk2Pyhzzp/uHtyvJJ5ZgfhAJUhzV7tlj11
bKn8dqMzUsCStMZhw3isPRDX57J7APb750IRWzB6WY+q4kWPPXX9aa7gR+EU/RRqnC31YEiXRTvM
++D4rl3SC9kktRVZQfzf6pow0LjvkclxgpQoKqtwguRc8iuWII06uAqUW7E3IRTwFOZ6CJH+YM/P
8R+uJotltBY45oiPRjyooegjTYFvnaYhVcCp1XktRcNK0yQ48e6keX7wqv6rh6oUdlPCVw8UtlGj
TvhvMtSqDkTdRTk4nyEzWJVqlBSKqROUdav3htQthrYRdVt0wLkn1CItqYNa+MBUBmR5HdX4plxz
afUlrpsr+xM4GIFhg7QjfXjiMkHbRi4qngeXG/p1/Ipq2Qd+jMMBKJT9eO0VPyNakpFSq5RQk+ed
eQui4bOxpsh2wJGEntmmf/QfTblvoy9NEG/DewI3LzxEY4/yS9NL/+Gakt38P78JsDaIcBZauFiL
0S2fSElpKF8iY7+GzlZ+QnlnPiTxtU08JbXS+DMhrqtetsdCu8Cg3QNC3O388SbIMlLvAPrDOazZ
v9sjBXJjjbrEgOM4RSoL64g+bzRSZrvCpB2Wx6QucE7UIEtzFljlqKM1/+vNchA73VzlTM9Gr0wG
MvlB/YwE1Q7X94yEqurEiF3b6ha2Ng+kXprad2qa8rutyMv1FQpt68CWaC0aIiJWIYE2ddMrXb6e
BtmO7BXYiGubqnJemTrM9CFV9ctstD0Mthu2uo2X3ZCcsBEESBj1NvbKxtUqtRO4nFfEEzm4Er5H
VobBSd/sNLrDwp5kRtDXirp5tAuAI4sWKl7YVCSCuGq5Kq7iOndC5pzGrkbTKc2Cyi+KNdOM4yQJ
5VKibEFerWats9HXPmTCVslcawGxcyFqYsWKoflYUxOq8dc6w4WGNiqBP4Xu7UO08i/2T0FeU8XJ
YPkfG4cYbaQDvTtxJT0F1Y8NMDNa0cuuKvf5YpRfv8FzbaZayBiGMboAnIrUakCIwSZ1t7IAVLiy
4WNQpYZzXIMaGBl6J40288SocWpMnNXIjyFyP5HZTExKW99Vp3oWUxiQssN494mePpgvMDGKI2pY
yFhaa4ksocHrqaj33SkYeqOQAUdAM3flQf5w7+hp0viEJscX8HyVVJQ+ylU1E3aicIweHQXMyQiX
fO2ZlhTqVx+KsujHQ96QcRtM6j+Tl+aomXNI7cAewR8d6SJ4wBf0OnUdqAIQOk9hOzsvARWyt2+C
KscFV86y/VeUPem+sSHz2ijZkawytmDmyx7SNJX3ZsRaH4QtSexHdNqnlGT6jkyWyw7pDF7rJ1s/
5PA1d2TS/D1JbVDpMmFpK7wDMSFIX2fs7rOgWnWEzs57DIoUmnrJ1yLPE+MEkB+YfnvxZjfF9FWW
YHbWwi2EelPg8scDWBXAQ6HY5NvZJ34zwn7cvGZX0kbeHTRBaWas0N4XBy2KElo09sfK+Qekbqaf
QU4qCE1R23YdDiyiSJMke6Q4TksychNOu4TkJL7sakg3TUUZ7mGIM8OYXMIzX0OQCVfN6ohM6tf2
eUcMo4+kNHwm0sNMIEMGPecw5K/F6kf29bdMQpZFw4YkVGME2cJNEm4G7VSC237fRF5cZUGGPzMS
NlbKJ7m+9TWvc1xXHuMOO769M7veWWXXRv3mGBgBuimbM080NiLtEF0LevKdRwdDJkzMu2AQUOXE
xf7a4AgWEygc1oS76kaLjYWOkNPI/BmYlwDtltHRuW7s0k9IgLzFxmXttUhpQ7+zRHFe05A1SAvn
ipIlaGhyXLNOdvzSnDbwBNRNiKwtZs/rbxRRXkraEy2aLKWMLEnB6ci4bbmA2BNKj7dGz+/REdE7
9ODQH3toYNU8ZxWvdQUz/9BFslNh8U7WwxigIzRgpa/TMKoX2pInHTtaN+88YGMbqZzarBzf14sU
YcWjZaKYz5G/qzvjS0/X9Dj8k6o08FkbA49i+kBXCZIBeFDyWnhGJcEeHGsjWQYFGm2nX9m7kNWm
u9q70vQycibF9x/gkh7VMvfBePdR8y+/Fkkuvj8pkxWIJCrpCjtXfJHHZWCxvk/DO8zgfZdbJbGi
QNBNtwngtdDjLEXRivg6TEuzV5fH/ylhiCDGWnVFCre5y7zDdqvq8aSUfFUMvdIX0AIHX7cXuDML
KWCfMYeJN6AWDp0VdGwQGILNgX5H0wAtHLD2ztABf1sNPGA5bnWob1pg3njznjk6d2ujKc31mf2S
2iparoQeDpzTJl32j9XxcXszVscCk8txH7MhSX1jENFGVYVWvRSnSx4AkBpCky9RGduaV6yyiXw0
JMf4iLEAoAr4T9DxnyO5+6P5BqujtZMM73HMBJI2z/ZjIy1/6K7YY3mF0Ch6tuRSsCXrvcYnX1bk
6Bh8JmD9dyBtieZpIHD+TIoEFL/dYWYcuy3KWRI8X0KPvR4J1/lAbsM7HtJSkllepy9IceZPlSzJ
WrV525ayYsA8F6BMp2eZnLh5Ln96NSUGUJd+E4nyN954lD6wBptry4X7fGV+JgR57DF65wfubVcs
wmZGmTjlktlYgjvrkcoHiVC7qFYDICllcsqtpIjg+0TwMjm14t87sA7thIf7k0zCwu4Ob11thGvY
QdYwgtuWHLDyez6Nv3qz/O6g7XsDbnwy0Yj1CfIYpaFBqKYVu2F+s/YCSgF3Pyflshm6wwXvtnWb
XarZTXYuC7WKd/uqKYjt4mnoFm96z0k+z8/7ZeGeQ9hj06+ta8WIINQMqZk7JvSNye69k3mRISzT
wlUbsHF7J4FUf35D5gQ9yvxxqVWQMaGQs8HvQ3meAH6fLmfFbgTFpyK45gZ+VTCv9yzSFyOYNycA
swKnFGOfzBht0HxQSWnnHBJdCXKRGywL2goNEkIT4k/TtUGEc8MNDT3154Ob8tdLc9gnzRKFT1pE
7Nt9g0bGuwRY6htCsJWCHE/+xlUL/AkI69WDgebyKF915XUC4V4BzTjJf9T6Pqn74RTPZNBZflin
L1nPsJmAc57WIx82/TN4tsEW0n9g2jC3S1lExw7HVMCUIHWgRLFk7qswBtqlChjQfQXbpGQluARX
zEMPy0pMTx/3CDL/E6FyQMA+/MA1arDi9L3Kz7PseSk9+FFpHEZTrotD0Rbeq9r6MwmMn7B4zE70
4N9+n8f2e4mwwodPjbs5MUB4mqCDgWu7CcYFaXWN7lEGNQYRK3Lm0OZPDNK8GyNTaVz067wc2DfP
83/KrSyQGwZ5Ern2tQdSwoYBJXcl9n8gR1t1073CSEysQvubY0ak2dV6nYtj9fumQgVrqvX5ubOh
84MGquFbfmeMteKJMOvE81AQeOzyJ4sNK6aDBI7WNGOLjbZdsndoKxNdrb4c2WelsXdQAgX6NBt1
yTtL4fHxrYTkC7E9Tt3/gV7O8Mh2Zxu/WEsfSoYPPaqGPqA2mWQwSI0d09XCfh8NNWWtX51xkVEQ
m1UWesrI+MoQqW4n0cqJtm4+CaRCs91tjV4gLcZkbxf5nOZ4jrvzQ9bC5SXEJfbsmHoEEA/f/+NA
I990wLECvWSF+mUb9Izbt4FnUFS8Zbx/XX6zJLVYrFTTW53rlKTsj9gSTgiQvnwuVpdQpynA09JA
RHwyFWmxmgdnV2O7inKKiIyTIc6LTQrFeyufCN8TTgLDO/TknaBsayDmqgdmYJt23thm2LHm1FLA
Q0pf2/9stj5f2KMYixZgCVZ4nTDYLgXzEsp4TN2YqKE23gC7CLZyb02pvC1FejARh8D3uc+/JT5L
fxPhhIVe8zMWh+bDsPr0zHVGJuQCdNdBB7ePgG+52IDQxCaPXswEA/wo5fDlfwnsRZAta8YfAwgA
57d0tVB8Zf4YpITyL7B8KWDPwKDsiJwvKwHgM/6RaDo9Uchi6PPzSChBOW+bx3QZybz5dpCmiLEV
k6X2kUadotzthXnclZB9Efz0cNQxFGareHgSJzvGT5AA3/qe8R4Vc7cXFlSdcaIOJE2rI9MOQeri
1NMYMwON4Mtbclt+KHJrrubIh38FqQiS0Lsit7TbHhD/ohz5BMRDquGfCLJJv+hDsB78tR3QzgqP
vyHS6XLkpI7cjKgBCnyL18OwrcKoLSJ8Zsv4qrBztb96LProOkkP1NIM0WeQNEzDGqOCjJAoW+jj
Kd1uS3+qP60SMqWXIg9swIdT00l23LC+tIBM257uuhWN0FO6p4lep2LHSqXQMQZShn4ranQ1FzXV
toeStNZ4LEufIFPim0oDpS9bt2XDV8p6HeM4a+iK8G4ydhqP0jULEDLBKnzVHsTre+uvuicNH5Xt
CP7GVJeDYwmsIyIqDe55Wzu3onPW2p1dPTdZ9h0WxeqpYRbA+HIm9tjOb9nSXh3W7IjGFz2tQMDX
40yq6fcTZgk/uuCA6l+fN018Zdg1JScExoJF4tLAK3bAknk3zU2FKTZuybeTmneekWIuBwTai7rb
6yPYP7JI4a3ToXvfSPDxHUIyhOW9i8CuO+w60vKx9IEm6+gczyLx4xznYI+mFKbqvZ1nv/mBZ0xs
98ttmdPqE2hbkDIGovhtzkwpeN4llQNpO+4uzsdSdn1aakhlBpW46Z/5HZR9dPLfsokWL6MEszJv
J7wwPIAtiQDLJHkdM4Mh9SHMYTMblHd8UBU16wALW2dmjhVKR1d9dva6Fxm7lm+/9zf6nXSAcb1+
w2pX8RvF65YFSuX2IyMv8axftm2V2bxsfVWT8a1XtBct9hLRg2ConHqyNrHJmDINgtdbcqIzXtt8
GhS7WHhNFKOrovvyAHb0iIfi1wz6ZF57gqxgRoKQC0rUmjvpTc5u6LeKqWGNOmgcjmDJlvsxpxxJ
0lhiD+lyjANsy03A0LEzBkxRD7DDSI8eG43eDE+kyMb1FZT+XObPqT5+XYQZB3FbHRGBSatB+qR0
kMRYPtAzv55Hcq7/zlarjDy/4TZdn4QiW/0JQDiH8bKgf647shePiBQrm5cBJwTpRDoOtc+Aiw4D
+obkpoifM+bm72gVyR+jT/oiwsfKlamjSYwCJPXSTF0wx9+FCRHFMlja8FGR2NCjDgPG9mmjIhOI
G18Rg5BFVYVmHNplpA6wq/fTmKz4Bk4VfxrgQg2DWhKMtvFpliZHdsnapZDMMdVSxcPYG4Mb8ejN
KRbOy4CGUErtcXzVoX+zKaj+DBT/lACkr5Pf5cVqxcGhvk/x37gLeDXAkyS/AsUVjdhu/G9e89ZL
+T14dPaG4JmMwCtw1D7UBTttkn02Jn3XwcrraLdEdOtkaiHDtYr5mH+gV3rpJ3zxOCdXBPQJMo36
nAYZwuKj0D9zohy9+7/7ZgOIn4v+zj4YoHH9TI9fNkRRycRqypMfwokXLJcJIyVuufpPpblXWA21
X1lGHqED0RYfoqAlo/yfoqtwqGPo7wmam4iASZgk/nQbDPnya3dz2Hot6eZG3uuQdVr7PJKrpHUW
lq8/o7R86FzWJ58bM5HLdshGLU0nlbz85iUS3njy64faYsdxtvfIXqiH1m3mORHQfBJFsDmxvnfq
fWM+tK/D8y127jPi9Ngj+H3eOJ8B73tZ6YUXq/QoccsLHs+y7sRwnEZL91VyRIdVjCRUvYKSRH6w
1PTMnOzY/O9E4Dl/4K7GmQYT5T1q4CmE4523drrHnO21EGaQoA2qj9ZbRFJbGOW18hpRSHB2FbTW
HB2V9fZbWlf/TcTH0RyDePX0HFOGOTB0MQLK+VX0PGYjP59qgtLcJcQr87+OyQBT0H+HRQo8sEys
2U1Q8r0dX9AGF5bsS9BwvIgYbtQHdQQriZ8imxsQb7b8NlxLWQH1puiJyTS9JliXvGZ79pj38rQl
4PG3pG9BhOf7l8WRfh7CeyZja2Co8l8cwCrovAziTeu6ACjfzyiDwdovuqLisXkOfpu12Lf0F8pq
/4Af5+TgiopgrnkgbIfHJpOwBMs3SKr9J+Wof+pxV1iZcrIy+9axcrOUCKDFbo4jRfF2nIBpo0Fx
NFXCNNX6sf07HdN7wof827ES6OggfFy6C6MJBmoZRXU34auM2KcT9Gt/5Rzw56+dySs8r4Xm6Sx4
KgkdP9OwC3HZg8V3Et8CEOoYSs4DcGfzo8AtDRnsNZtKqNxFX+/D549znU6P1h0I/AcjI5IGCDnl
Fl5Y51508PE+0mHf4W7yFDjAnL1V2gUB1ph2qhkzkFXyqCvMv1AFI43jkKWM1sNru6ATbU6Pfndc
S8u0AcppqJhCRT0iBdI1pDw7o+J1YurjPhCzjT5p1nRyf25dgYGY/liUPywzMB6gpCTLBsOFRkt+
mabYUh6BFx9Irj+mayoqBJDRB4cj8xuwjP+WFUGGv9zQ/DlMAltpXptMuD1jLOhysd7VFcU+tECl
SFEKugblcIJGMnJG91DIn++sAz0cSj20kBwoRkyrbISygi/1VY7QG5SBo7iHeULglf1lQSOR1gLh
DVgHMmA8EdbaSvBHeUgmLB5yys5tcwh79HCvJ1Ia8cg6euJFOe3UYaSgugI55XAYNb+wmoGceOJG
Vp3YohVFWVz8yLY/63AenNCir5QOD/mR7AOr2u/8Yz7kKmLVxDibmMcBrv+zN6cnrl79VNiSu5A+
cjgJVS3L0wXwIbx5DoBRfAT93OfENgI5yqVRJYmcRlRZo3rsjAQk58SlopDAzJco/ezN/z1khCQR
un0VXdBeoWAQi1nH3cfSYudGAYhJAS/yeFesWByf7kPK4zfyr7OYYPjT0fjqLVL7aAfl6VxAF4Z9
iyX/OMIxgrN3n6ZyYMbO0jEDvEdvh5zuK1HI4PDXLoMSE7eZZ6BT+fVZRnnwzOoZBOpszyjbZoor
UwwvTxh06kHKXV9j4RpGNhQ1M5XeIDrOBpeIhtZFFhnjBlqWEoxe9Xz+Xa2Iw4FZXse2Oro7Z9Jp
ALs1A3NbPb/IfNDVy3dq5riwbkrgFhiHHPGUmoHWzbVSmalwWSmsUzqnTVJ6wR55Uyk6mdmo6r0K
9hm1ksnULk0MltIOh5Y/DViybCFCgUAISXAfEVgITzxKZt5bdajYuQNqDgtaWAhBG5FTBvl+6wCv
GIz018NL+4YFmSXpRyFhHDbRTO4qKtfK1RZ+YYrkCWD2KxGX6rg1JcsH4qDFougxw/Vkwm5+fM+9
/FV0V688nT6BJqJyRm96uogJn5b6bYFOkjEd9hubU06HimilS4rYw8fmJ6oQNAd3WUpxL6qNLLFi
0QRAeX+EG+Xiq52KLOuYCVYWQ7s3O+hFClfMSRyRX7+647miNWBBke8q6EzJEWsAtU5yiT4hO+YA
TJc4Hmi/FRtZJxNslgzDCKc/hgj4tWo6ByQLbs/TTs0cqQ7kYWzoEUD8QKIV4dVumM9agWlm1cOe
J2l9gAONteeTYvICHe4esWueNZwNF+Y2xPAdkImr3C+LckNInYJvUFXUHIiFLSoj9EHGpb1BxKpF
9yGLPB7Y0mXXlzKCuUv9O4QQq66NMFimIE8SxnMmPkkRcf2Q9l7UIvw3vI/EOb8l2c003rS50Ahe
vM3rnLSH+KkmEOQakd7aeyCn835RxoUlmlXNHPIVh6HfAbJMM2szyGgyCTVrYRHSt059jz89MbEf
Z4B26wf90Tp0fA2N6PC4MuVMrIsSV28EGyEuqShg/M185Hx+yige2sKFVBd1roXTlMjcRJYRWBSe
oxvN2p4ilwQPlPuMTM4TQrlpfJNPPUT4ooosLqQokAgp5slimqxmEEVW2J3GjD/KNiA08ctdVkIa
GawtfWmdNf/0c2l3n+ToV+fhPwfPvddGHYPJMFOB/V6Fuy/AyCm53DkUNnpObSjRR7IUOb0/jdsk
pA1f2BwZ18WNeNqeN+c5eKgo9el/haEvD7Sdldrecky75vX5U8IXf8+fnNbTC+7t7LHz/G7vuagh
vqjIuzxT4rq/sZMXQKSKKe6S1H5Qf0qMcBc/v/nOW3ENCzT2Rlo4nD9ReIwsf2u1EA/zfJlTIKB6
ea8acsHJaPs2t3OGEi3GYqcPh7cozXk6XvT0hpHkBgQJucLuEzf7u683AQuPr2xF/CZNJjxUvZdf
s154nI7V4U5ds/YwpoBXWGlgx/OwJAbMxHKH5cAfUmJH94wx2z1JbkTrZW/9C3K39Y+i7s9ejS55
efRSJFEL+uB4Meb1Bst12E+5YamYKRmQ1xOq48kRkFP77ugdBrueM138R1bCMnjztx6mnE4FjoqD
1y4LfYB1uajpIBN0Z6x/j5B8Yw5Tm1b8uaW5f+dXD7Ec9nZuJCbnTj6bHQNoJg1tuF/TsWf19xN3
Abs0U3NPSRcNU2mfix0NfJQ5/8LddibqobCUx6bXsjP6AZo9Z7bAGHhCJMN3P+C5LQs2c/CEoVlg
VuYYj+B0yoMo70cTzEufau2omd3kIKW4VIDG93vkEssEwUiG7UaamCJO5b2KJQ+5BLO5RYc+UYU/
nvxpbSUdbksHZoELDN6GIA5Kmjve7xG5NiXTqD5PAjuWt3Ntm3eHXEvF1lXZY1Xa6hGk3KE0pJaV
RoEzjxyAFllA4fMznVfJKDK14QDhgka8bC8aZzefaZO717yqC18zU1x6XCZeZKCTDFapKFXXuhyl
xGnpt3dXXDwzCOkgbBsBl+HnKC5gP5YKWAIT6GIvjXnn9LABfvn/CfSPo/NKso1CyjU4xNlVY/7u
rgVs/BY7dj4j2AUxpVsDseCHYnTcwqAL3TyetkGdxr6zujbRzKHs43gSbauDkQzj8IQINVFlYH1L
OwKN5nG2NUwxxAJVR89QBnBWeh67FcqGjN4mhh3qeApvvIgn1yBIE1KlewqBWmweanJlE6LFA/Zr
ahEoynPlCk6Ch6ltBGMaKxuzADEwJ3Nk0QGqMAFOIB3eFkUCI5iNi5/oBUlaYgLgXR58Osk9IVID
MhaShZylRVyMDHKgUtUYwDmk7SZfAMh6PU22+pbRhob+WVJwGP1Bv1bk0V8j+RpI5rwjKohVQGLi
9D5X5YwddlXTQEWRrdbebVjMgoFhsHurszA75b7G8j69tGp9cM/jUlUX3iC05x0eKbFIL9r4N2KE
WnTdRhzlIKspo4VBlUrVlaP2ghIbEBtR7ihK2dBCOiKGiHEzB4FtgklLri2eNdS+Et+AUqUO1DZC
ag36VVxnSTLw/OXMxs4H51hY1WSM6PGRTMG6sF0MNXj3VgGwqkDYrFUOA/4lhP11/6zQqWF+yBFg
fsbcMTiwTE1Uvq2gBfMAsEZm6hjZyKT2B9brtHLU7dc+jbmiSnua1g03NYIF6fFp/dtwswQdlCPf
6Y5Uu7H8Ud9+ha4tBR4+mLmYLOy56gWq0AP+ibav5BS11Z1joofKInsjALLhhPHszEWIT8R842J3
hJ4+IEoUQIH61oASUfH2WnDuiFehAWwRmkq1j16CWGofPf8BVlqhURG+sE82/82Y/v6bcf2HLnEa
AyvxLa9DD6Z3bYLvJRsUiMoJXyISBO5oO7ZUeBZci5DNHz2G2Qcs4wZHrKNA6JJzc99yYqqGAHhZ
VVDwK4+OyvPdN4E50xCIxDF+LGSIEHNpfQZQeo3xnkTMZ2kVOsjek0qtlJ5BawcKDLBXxBFZn+tN
Pc4ZOJqh6+Oir46qi8Nuc1Xjx7HRLKXSRRVU97yTdhrUr7geI0n4F71Ug0h3OYJGkWrUBV7Yj5Q4
nU0UacNFMgmy5pDWHoqy1LllZK/Nnj3sT4XugilcMEJic0oZSIa1wazzC8VptIeQYPd+j60YxRyW
VAv8YLiKaIiK9wtmoA4YEKbcgo6S0yFkfQ4A5mvuWSdiRvIy7ud6Yq5VyWGwYESaz8gcJqMudS0T
REBOkacGNwfswf3e8aMp6Es/bbeJaMxsyKx3OZ2bESjwbaI4SL+XVpi2vDNJe3mZ9OLelJGPRpbP
96/88HYBi8++kMrf/S0sMgzcZfQxaEdF+pDUSNO4UcDt5D/MF9yVnk/cmqC7itSnuDmL699LGLM/
ApgGJy8EoaFHT7iUEsq6uKQ6haNjdD3AmGsdTDeq/ElqaqgDeX4kNdAZd/HhgebKziXaaBIztsLn
1ACVQpBnDAc0bA1YczEPjHNxunbYq1PD6X7sG49AveoS9yUAWUi7MP8pms2Kr2zbEj/biX9f6msl
CkyqwpEg4Uh7d1KaxRsMIeE9obLmkeCGsiMelIHU2Kle/3H1rbF4BzD9ozQDBjuP5QwIXyhNQIZH
fWFfsyd3EUctoM06Ls1srEl7+0Dthn9H7/yj51//bgDPCV0BA6q+b5jUN7GSIrRTR+fZcL5qog3d
R7nBXGaqHzn8udv5jT0jmprAFNB3dr/xfYw9czWJrhxv93hLyNX3pQ+li+XQ5q7bZYgJcheettWT
zmfTltlgAH3vM8K/MwSPq13e2ny5bXIGDlvSzvg1T42ePNmDyrjfVo27VVPsJNOIdcFeqjaLYZJl
b7rbUV5ChOjF1G1/oHFIbTQ9K/misL/TMp1lHL3JM0yN/rHVNdGw9yP7AMSDjpz1QZCdbY/Ej15/
ljhDy7VqjExDkegF4TQf5idn7Kpbwx/CaxjxL4btFu5NoyUVhRakBiZU54aADYzoBt8e8JOE4eHE
nx+6mVqABHb78S05ktwteUBXM6DscJelGsIawuRIgMQkowPsqRQZottC8bO2v19TeHvRAN4vdfAw
ee5m//gDGhF2aVmGB4MHiFuK6nOj0mrQlP3hmUebFLV5t/VbByXyOKaYSFCf9C5BqyYWuPWYcyUb
o288NDQGCxpjpSBBUeVOhh7RTF/yvFrXocEYNbkQsmJg5FrceorRfOklgROavcYBVkEmNdi6Twnz
KvOZQhFaBTbioZxy43n6CPmef9pePobhSb27S05z2FNv6LBtsSPCQtfqE3p2mEa1sGnFqJr6uzH6
yRUvFe4YNzw8b5HhHBfEKsHxtNlOVV/1Ns+HqdWbYWcWjBZViTSxR2Jr0wY2E5iX8CUFrzAqkgs8
8tvjpNu0CB+JijrzNm2cIujkxYv4UkyXWHscFdT5IVzv7ePahACP15rXK6pNi/TYaIS0wX8DROp7
2o8+M+gwW4vDMCNPDmGF/dXgBqXC9p01RBx1FD+dXrI7IkKXIEyRssjoXbVjR4j8pQ0M9R5/IRKt
/UapIRskxOJol/nIW7lNZv8evjKBYQAINaYI/Amt+eAcbpztJWH4gl9URFXVdQqJUvLDxq2f4YsT
cNRcmjXne3yC2CHyGuufDsCz0WgU25lzHrnea6O98hkJTatrEAYqisKQ9MFkUhFzMz9oDRd1Hc1D
l0I4/8G+wpC4UDihU7PG10AwDe1GXFIIm2sq6n7CAExBDx9qEIeUckwBKQAsQEdvFUJZVRSkS/G7
1RhRTCBcEJc58CBp3w1Ex0D2qMbsgzVxD0fc3vQSYmMND7Qw+5RASO53hUM0ukN3uBPDThunkKE2
sGwrHkJFS31GM2gVMSsQN1lCVcqDZ9zn4Cjf2jI0GpYrgcC5rUiPi5Ht3v5t4GIDs+Qyv5aQI1wd
PImd/9tn45D0BMvrfabab35ImCrgPqx6SoiDf40q9lTlQgpzcvdB4e4+2LoaDQlHEvlJuDiqs6bJ
RuwwZOApp5WWAad0eg/bxvFrxgj7MHGy8ikGg5XDvn4VTEncGftczTEEay6CcPxISkmChYVXvBrK
lSNuzb4MsGTQhuH4lYS7PomvjRLN3euromi4YXVcLqkEkIAJxDNY9RyPDaOqyLrhgDcbRyYHlnPZ
7JiX3HqTRUyhlg6udVqF/2D/pY3Y5RV37ptFH2yVVuldVfnbf3v381MY9rCU5KvTRLz+LLYJ8qNL
Kg42OT1gT7SbCzGByx2+AHHh965QdSVddMj7bdwR2/zO/1JHjhoQ8BJYSauXBVBVG4kvord7qd8M
MO+fu+mVu6LHrgNQCoB3Zs6kGhnNUIzYLGN0YHHOlWJzSmIHgcG42ZHc4A167FhwxmwCaCmioV4F
MPem0shxfdbjEjE0g40vWzkuHOVd89unW3TrnZd62LnA+t3Xyj3RhNeGH79FjXWf6hbvLh9yk3so
8M5CwwWn3yZbC/ngpnrukWTK/9Fbc/rjatE+IGHDBaBFWrU+qOXCpto5Sikr5jgH994YYmE7bqNe
CBzzeeyIAPelBR8uql0GOFh+d6+fkKM7gOjrxtGHZzqm9CdtQXwgOdYNF2/AdNpRqF/7QNIPoDGP
FOCbvl3oitCk4P2l+fvVBhI0r2+0M51qFdRbRKtF1dhs2KLBOdkGYxpqeTuLR1zsdQ3e0qIyZ6BX
Onwt8EqCwiIrJyMw+ktMM9jIhJyr//HNB2+kL4xr/Aa3O0dFesuHawZglpaYv73C/f0zOfF5MzN1
sHUh6jam2b26deTFF4WMpeMJ8HvmbIo1DTM+4TqTJzI7GrKN2Meh1OlTzff34D1mCm/K1hJK5jug
Nht7i3EmUxmSCt62BxSWtA2a05EOnUnLex9jrUViz/5Z0ejVrHhoO9ce0KAbPmc+ltF6ZvxgCDWz
C+SUVtO2LHeNMoDrgl25mQIN0ttCkGNMnwJgRy0wsQTiifr2wK4sjXs9ojDagFnK6Af47marquyK
MwG4zcugRgxaUH0uInAxZs2Z4qERHZnXoDXGlusd2OBKf5gjwPvr/IUHa9deS4ssN5Rk4z3A6ppF
4EUyEJkKZkXOLPs8iJ8EQYhw4snI301iJmw+QowFPoPvNZ8Dd8WnLsedd1gWZE5POhTOorPbqw7S
88+j5TipkgLmrnKWwn6K8Mepp29KThpwfy4QZUQ1PIoFm1Jok7dnw2W50xELIaKVqHJr5s3wawt+
jI7YlUNBvKi6myv3TLaC1+NOOryhtGGVKNo6eZ3OcCzH3fpthbDODHgYrAvw8Wn0QJf1XuiqxFa8
amquYi42p+EkWaSK9DJnyTI35YFTpNAz9y89pzBAMJ8usL3ujgdckK/2HftXdI4gJCZL8SIRv3Sg
d+P9LnMLkjQ1U070V1tly0y47GdnMUfeuAkt4Omf3kUfslo7kkQbsqFSGOFj3pTMo/WEs4cXO3U3
4D6l46U4Wat6bcLppsMtbQjosAcXx8SY5MnDOoAWdeVL6f608oJoHp5ZQ2TKcDc42uRGTkTCtITl
GJk3manuNnO1t2J/Eat6LloldaU0yuAlUzjy6ebmAsh5hKJmJc+Ge2wn24eJLanEOOhShdxurW6m
RruweSsQZ1JK5x8z/4w6Dgh+LjM+q/VWeRXUtgXA+8CslP3ox/AHoD5c0fuVj5eW7JRS+ow5AsMW
uH+jgEx01CYUqjdnARM+1xmqyFqBEhfkL8Jvol4+MFsc2hj92sTCcJfzBQuG07nusYgJWueseuS4
oWy8Xo9qXqgNU0IpwK8Dh8kGkmFMZLLFw4uDfvWeyOKpC9JDLlhizSOdxMQENfi28WVqD/IimCNv
0KaBkNL959Ga7hgllSK6PpDSg6M/F2lywCF3q4Tdk7CaiJ3ESEhGqCRRrxnOZdU9MgNqRu+CHdz+
DXWX7gO+wCAgEkVZFWY/LLcLhavBIUNHJecCdyQyCYpsFduUF+PROEAvauiNelqGHrQqRJBYi80f
CHgeTa0zBNa0LPc0Gi9TF/dU4m003WOYMrS0mbUeo/vRJpr69wKUrF8uuzCBBHMhN8P0VKLbx5Nl
a7bf3HNPguo3ctQq12lhUksiGWvmRCZbLgraUk9yj9BgXrPRPwSUvl099Ob7IdLS0NJxEqeB+cAS
dTDwI3Tv+GkkE9ZNSLXYM92C8NMppPvmDyqxo7i2UUAllRMfGXuC6ZSKXbKpSC8HTV4INAGIIoox
Q5emiMLfKgZRBFJHWzUt+i4i2HaGbOFvk5RqUXwqJ0NQgbf/WsbMnQMdOtetw8Fbao1CwiDty6V1
nH7pjUcAb/LIG/HDSmqgWxIuQGQRyQmdbi2oyZK1KjfqsI3FHCEgni17a+6pT5KNKqMt7JWzxdGP
55iC7o2oukibiZhpAGLIgw7ZpaqfjwlMMGcYTMUK0YO/tR9pHF7kBm9noGV5CFhNjarWcXU/vQkK
NUGTnmhAo6ilnDYOPCFICLdo4jRSNTbBB3mbgUYiuwRi9OzhIGmQ0A5QIEXkWK1wvoEpj3TL0Hy2
Ekm4Dzz16V9AzpG2clO7nwS+dCL5hqsr7U5Pzs2+XAzCposo6wXdlmy5ZYhXa+aqSKEGDaaX+TvB
mJ2s8e7JsTVQ5xVlqZMzfuNbbybsrhAPyEO6iEKbX2ikUfeyBPpuSBsd7NMwpaT9rOhLqQ8uxw2f
AmKO5ENfwW9hB4e+teCSMvv2wFPt0pRI6ZHBNbbO2TxLjIzwF+Fq7Jye7klB1UWhCkElOHM7Ahnd
+paNklAFzcUEy4Au/mdRbVyQxBH6xOpKTRS3hJcwjC65ZQtQIUbcejROhvoFJRJEl9LZkPdaTEEu
nHvtCgal9N75SWvet2arstzs0jPY+ggG1llKaVd1DZvc1+W+ljqik2Nup8Nek71uWlXQO0ofUGKN
7TnrCs9FJ3Yfqdmku990Ht3At4HO8LBmLZMTFO1GlrtC3aDmqVSDiav36m6gLuGxrDlgK3cfm1Q/
6jkUfkS2fsfwKJ/gfmEm3rv/xJxT4d2pBLDFehPGewR3FCJPcsbmAXlX8FAAAzkqEd3Zf9+B9SbL
rh2lefCOXxbuIMK8sXLBWT3L/Q/WWmRb3nZMXh3pdL6SyOhCel5W7KG6tpe541nz6Y4KVKi9QVa8
VljSlGWkAY9qLhake2WREl0LugurC9iOuMpqI6Brtt6aI0HDUpBMj2ssZkRHi+IJhrQygJ4lyoUE
0z2YQuo2vQRvzgYS1K0bVV3WF1LrFwUXXcrxavCHZzW+ehmm5q3j75Ui2BTNkdWBp6TshRVUnZwS
unKtGzPaxarUOt3AQwvk0esenl1XsXOfa17PCk4rgLuDER817XI4nWgZZRVB4T14mToc3sY1e578
psAb+RCF4rZ+ktvE6f3y/6hBVp2eUKH69pEo6WGpDfeCJo4JXWs9JMHHgceD1LYIG8MlC046fXTa
IQTVhq3Ppy/u6apjj0+lABAUTNolnWpdZp7JAICA82jJHb4akFMA1TGxl+udGpMP/NS/20ll7GIf
IzwNpGBq37iyuf3ouwIwTZYA8sxL/5gwlS6jdQ6JBY2uzyx9TvzNgJbGIuvQJA7QrFy7shjAMbUN
6uRj4O2y2SkFOe/37wQQYd+RGxApvM5emjRFCkE4Y1Ho9M8Vmg4pERERhHx04H1DpVNSSy/cSAg7
fYsS2qvsDPkbIT1+bf2YMYd+KPZs1CAG0SsnnbiO9fALFfXpkV+hcCLiCUnqO43FYnBwIniPpJCr
sFYBp3qBU0m9Osavo/qPzNswtvhO2s1z7uS5W81k+lSoGSbJZv+gitF+ed96JOhxKbxL3F7qgc0f
lijTaMVaLTNUP1kbvqkc6sbdvA5B6QNWHApUeMmAyRd2MlEt39YRwtiDnoPsyyWjep2YsMG2Kh0S
zyGsKPJSsMF8QV5uD1ka3SLcRofAlGKIm5WeZt6cV05ZRom4TXGCgfZeeLqdSmWYbjJZ+EDqRYz9
v2BjF1cFM9xpUfBCpg/Eqb9IKcHmZU8y2+8sQUJZpRyfGHpFoPOmSILvhT2wxS5bBeubvvyOYw9L
ngaoSAYcaQLMDsbxDSd0FZBofK2abhxHqxRbD5Ve6QbZj8LTYEwCuNkpK8dJseoYlk6NPy08HmA6
zYY4zLheE/6DwS6B6iqLq4is/gEWwcJFyiX8I5ZrEmdFvfYUY8C/det4ObaiKC3cMtIfInKviPsd
zkvwzbov0G81toS1CSsqmDeeSWa9NEke0ZP3KN9sR5tfXbC4x1YLGVpVeUloR+HuqcpaYxYk4e+H
1Stw4TFTQDFfEBoxJY32U3WHwQ9npanom06F+WPckStgHzGRoaGamOIlkpCgMoWLfpUZppFxt2On
3X2MveIqV38EYR68YNszyAddtVDebYHkN91isWOePQ3sywBhe6tN8aEMyVIuUSYC7Ww3RUpWqj6x
mhditKCvoXNHUPfRg8NBdzrUT48+yJPjhb9/0Z35Izo624bvq1/MLG1tqw8LwUj4DQtoJCRkaY5t
7N0oiOW5a1hRilOZoEzcWzJaw09hCIXWEyZKZ7ervNhTf6ubWev2A2O32b5mq1VadmvvTo9hhhah
HmL/hqje+k5KV2mVs6WM6s2NYBTXtCD/Hs0VaTxnLaDiFzVy4kmekXf3J4fVDPDbFRB3nWz7DENJ
fo5p1cENPDmfgbRM5KaFMe83M9CY1KW1bRoG/wndh2de2lIWwcxmOZuSmJ6Tcx34m19n233pjYF0
yrvTVqoz/5z9fwsPPQhZYmD/z6LJFcaTeQvrO/z8wPf+j8QtA/fGYZbtLstWE3dsRVUHO+2WdgAV
xrTUHKoPNBEhVWBoYFh2a/SEe/yJ0qxTQhIZAxsiz+yxExfgyPyVDWLW1/sa5hgWIy0dSPmE0mMW
MOnaZmgIfLDkFj57qW7rPgfzdR95tmnn6QhklTtOKLaiMc/GASEh00mc/82A+nLZdb+VNcv1RqcG
4yjujhskAbH5mMq0jgEXooVM+Zz80T11Q8RlUeNJDRFDkPc7p87JlPXz2CTRH3gN4fZjqwbJahpU
GQIPhMegpXiaEo+plvTJEOaCWnbSGUAKliPdLjo95obgNDaWXIg1dnixVN6865FNeSAzDxZI7EHM
EUfT8gGWl5CVQGb+IUEbDpxCWfDOdnQGSmED0Kb9QzR4pKANydTmYKljLcmZIBCa/fvvH5qlmkQF
uoEfSq6nHta5HJ6ZuM+bbPQS5AGuTSEbWQsbzk8Dq7mRKqLBtecGohY447rJATZsDhWMc/ots4jY
Il84vlcb4/fa4Rk0/9Y2NyZzPx4ysXKJYbNZEeNWFXiD+iVIbO8MGvcmYvNsbKUta3q6ryoscI7P
cK2OG7t1/qAKnQx/qVSePqg/qlcuJOo4zpzD9Q0O9OyuetiXyAIByanHuyqX/vyiZhGkPR3Gh7rQ
U5ySUVr7obW7TnQ50W62bPzBMDjLyQLMB60uBVX9BdG2gGWnLEiMdDBPOjHJn1wt5pD+86e2zcpj
ew+aAvYRzPsHehxB+Wca+Nz1zx4zZhpLewoY39UBoY5am9soof1MX9BmlLjt1ClTzDyR3RY3ZYLF
5kdKlGExhME09MDokJyfrw9tSh8gxSMEzVEWImHuQHlJai+iDFpmcRPrlt2FA3I5ddXw/wa9AQjO
7F7QsE5ICGOYKFRvHUvCSjApyTXl6DPISZ7pjl7/GEbZFeCXm7EWLMPNI707aU7ZEa/9diaS1BbM
GQR7Ictq7Kndu64RiTwejSMXfbLpF1dEBvLzHEA0l6bmm6IM/+1f+k6pTOTPKLNX+h7yiKtp342k
Hq3VkLh1xf2WukMAKm1GHCXU/EHyrc6/LCVwqJ51dxFLaTNDRiDvD0haVwpehZqCpTUiCxi++mQx
kVCgoqCwM6wSM8vncbV0NO/7yc9/oU1pO1gvijn4LBNpo8brISgCuNg0nqcsZSQj77r8VzT0FwSO
XHitD2PXj1Y7aAWHSc9qgOIZhOarfV0f9OvU88GPqtVHIeHPwmZVaZ7wg8bVRkeTzYt1axKqdzuQ
u6arBznmWL3uBdywXBmH1x4qe8PkL8i1tXF7LKy3agIlIjMumP/3Gr/8YLzwsbs2w7N/9ho/jbEh
3V7+yKmK78IWqqJDHK7D7l8HUe+bQjru7kr3WlcdJPrvFjAbm/erkZB9KPnwWGpjLc/NSkY5H96R
/8J3frMDRi+fR2TCxG8rtZBaxYyJcdP3nqcyfocuiine4fj9gsDhUGXbtlqpb+WUYh8YIxkxsUdk
x6XS5ekH5PduyGJ4PJ5OiB0uBegz9gEIM/IjfXjvq20SFAdONarirYqKyp58S31FITPd6PPWu82O
quuG3hbZtT46Jb4DZ+9j7nyz7PaDehABKkkz+ImeM5nFXOGC2TPaDChqJSL51snNAu5gousFEAVj
MmsKR6pOBOglWf4wkmpzhrN2YTCcVhKsrnE9lLE9QjMdBiQtAakVqYvur/zSgSixs7bCu9HdrXA6
W5nVUOz4CBlErn96Uqu5tCOo8GFFDuHUf3O4WsKuKNo8g32oD68lMeYdHb5PXQaHqAG3MgrPnxRt
htfH+Y5Mw0LWREm3iHRyH9THcdfyjdxN3tE4x6bfoh46vjTwp5K5AoCHCWPQs+AlDKIMPczjVNxE
cLSbydMAROodvQoh/1l2W2OJ2Qd98asmuu1exKbTJg4LR5kPmYRZpi6m5kBl2Bm3vVB/QDy14A7d
eXC7Mm7uVZdvkA6e5HoxqEvR70fowySOPuzncegDFeTiLidJ0jK4G75xU4r012NX6VIgmg+OHV+Y
VQi+I5vLzY6Xb0+ggdkF61S0PCrgjPILIrQDeOlK1b5Poji36qtboHHVjnKfBVufl2fofJNTRhSh
8mI8o3R3B00jFnZ6o0nYluAd6u8yCsGtgV0jp7l4Jcvp5ErDrx7j5IQnDQE8OoOyt07WNclVNQyQ
4e2pvlGcJRhAAaMYDGAVtxxZJNQJ+aWLCZbqDPBdB52Lk26cQ8YJ07U3b3eEVNuJq5k1xw7x0uXh
A600h5e5afurxzTNCYpBxOICBhdsV3B3BLam7Z68EMSKp3x7DYoWBy3QmSY4qq71as5ZkA1v5ryO
ecRMuEU+HBXTSwuM3+bhXvZaOn0nGU+J3HcwC7x92wSyOukOIUd/SUFxtatN2/9g85VisfT2q0PQ
0RJJO/l17w99fqoBfz5L2L5xYP+gVBmvG5EhwumrErFhqYV8yJbhPbm4E4xUrdbJgu5LudaZjkwC
eWK92xFKPwKyJ3JR8UHZILy7TyyjMNlF50qIy3poTmrYzKp4fVub7zFKeVU2xQOeZzpZDic2+QhX
h804BupVhVz5jRMHnyyQBRe4RK3N3Mw4axvnfoNIqhdeu5afepZoQzQxbD/dxeNbUn82dWkV0xaF
T+qoWpIex4gDhj9DMaXF4kfdRwThrGW/paB0fAERQDdr7toT4q0DZrOqdfxVONeXjQNFJQaUfVNv
ZDLVzay5Giy4srEfLkgaGynLmzPbBawkon6TtNV8SE7pP2Nh6unQu0duqvyeoFaGS0YFR82deeY+
YWx/DOPQnpWdH8WCKOiAoClpRY6gQG1eoWFTbGjSjgNSHMqtvoFww4F0G0g1m3Tlbrtf2+wbzNPQ
Vt6N3Tji/VsNHCy4hFnBb0Qs2QCMgczh+FIIrqxDC1jxgIzTufPSqYbOViBiIiFJPYK/pIQAD88C
AfZJY//WFJv0MmPzRlClLtfr+l31s2Njg183O8+ed5F1SY8uxHM8nZs84Hv6jAPqEelCfC2JAcZK
jqwtu9/6/MuPIMgQoZ4hYeWER0BrQc4+e7KFzBlJg/5totk7+aycbQWJ69YTuZWV3yj/MVKDQoEI
znQvNGzXBJ4hgYd7YcWExUlo4y+Lqqja7XDG+lj5FeAtLfBGblYlXfA4qahnhz0rnXx5qpwTXP5c
pV15L+D3ZqNRFg6HQGOS0Z0hcS9Xkv3b8ujrK5qgzOUfcMWmW7FUHGXi1ifPEfmBuMaCwDWTpM9U
7B75zXB2LSSxlLbx7tyhT9G8zXwr+ky/PGDDzYocHt4KxGF1zvVWz+xsLMenx4xO2/fb8WOFRPAZ
i2l4LTz19BLhbhcjSYJ9UKthB8QZ3oLcz68fAWyjDM1/d0vV2h5K6vsz5zueOBPGraZqIWzxFjn7
oLF/HM4Ec4avN5zFTpQkmRnTkBJi24yykqmLd/7u41EYiiOPf+NXihUW2F89w3u8cDjqnYPVKRjg
vHwXDJ2nnaMFpHrHgCE1PbxR/Z9imRfw39ofyTGCK8JZvAvWXF/UNgJFbtFPtzKMq+YmVQ19uocd
VyoVsFGp6+b4RDDDg7PTbX9OmnjdD5nzS8AqmRv5kgwpg6J/pkEIbA03qzsRzzGXaUeQuiTSzHhr
xMVbX4o+OGCfg0Z5yJXkRC3TwLT5a+Oby5pfqsYydGIQxEqLQJysTBEYrJp/RYV21Tsc9xiipaiR
v2hQqGOOb3U59y9ra3BfPWsftY99lUTOezuOCoMg5XWRfr/6pWnnkW94f6zce+l9cV3VhIDGBhYb
DsTv1DrkVwOFdvoTcPqNYiIw9TTRfM/8bE0mW3aAfox1Xq99lzMp4ITUDRkh0LHO9nDXNiNrqS+/
uxeXTIUlz4BFXdihnzUeEyqBATIMfAd6RUC7VcLWlH1dHr3k990rwFJSjoMoCHNxgfx4/zyn+4Js
JlXAw8grl/NKJZkehgzi+unuz9/mD+kQG+Sf00qukyVCeey5OA6peMag3HcK7EUJOp7MWulMXnrY
dXQojbI/dQBiWiWeG9hHBEwl3YDLMyJKQ50/6yRD5BB80yFlInsuDTYOHFKx+Ybut52fL5rlo05X
FXZwdvsC8pM1vghuM9px2gldVEETyHu/B4ZzIXuMrOfFWH9Uo3322REInhrU03+GiimieQ0VPDLi
x9deIXU+evrxUTQL75+BPTq2kyci9AjHc5Nx8YtogpTReuiqOUu0Um6lsi4qiKvtplwmnLBjJDMc
FM1xN/AiHqv7609BT938wDWbq2cre933DtMADuczBHqq91ww6K1DezA2ldiUMn6RUmhKNvPpUqot
dXYjHsR+cA+roCP51ihHV+Ym3Ce09X8TIFDgfC8xtFtglmSKkZNSR1eDPoA65wM+QjauaueCj3Rj
aLudtsDXFY2wTHB/weD7fqMSj/hVBlg66TS9+pdLIC9REquAy8IFeDPVuwitaP0s/UPsf33G55S4
lJk2c8tJNlVZm0/uXJ9B7aMXCbZt0rB3RXuJq8lc8CSZAM4gN76hdo/5LyOhBUbMbaozJgQ8feF4
q1czMfBvusWZqT/ugxFSuY65PpPV4Cxz2f1H8/iYSTeq2VsEZPbvl6VvBB7AP/2G5C5GAz/wIfx1
cKDimzQPi6LX6i1P5Mb+iAid8V2Y90M24kdc26oVW1gdQWXBg2uLS6DVMbGmqd0+zUZl8WW3cTOb
GmVc5R6KASyBUl4EwZ/mzyTsUnJpV9TnHE7lW+HXpa5WNKy2TkuUI8YZ/yjixGXffBYZN+/aQu54
No0DzBuu2N2Digh1tC7a4nVdpCwyN65TV2u1QmSkk6Ki6vCJO/K3aplG/GBykVJDsoejG9UdgGTm
OSu1lshhUZclkcENz33qEBmElDHC15ar+3ggaB3VAGBOxCM1MsfkomP3zf7LR7+9fqZaxfITIUlp
P5q7wlPen/23rRDRmCf1IazWj67xQJuAZKH+LSAUOfCx4A8TL05nnF5In1Ooqz4ixUOXGvG6Nw76
nwTPHagMv8B8lJwgr+jCRCA3ZbTjhFnwwVYqr3zUKPwgATEMxe3YQ7pnvy+H+JDyGPlyA7DVNavD
2VK5SNsZF3YghNATLBPSfN7787scNH7lmOnZYrxh0uBjBPdkh7aiYtmncarGe/kNKugRSuWpFcs9
4BTIPkB85nphzN0/gByTh3xgx5Fe2vSMGkAbiWjXkK4Yri1IJ1xOzZmSfvKZcCTjoZ/GwQUddNwc
3LVHRII7nvFWhMTFaZhyXpeArZEXqVdjZLtow9c4gs8HFu3RPAO0LyaeX40uBnWByNnTK/jJtCzi
+z6kMJfIPDdQJUz6D1aTm+U04l0DgzVTbWulvoocOP52Umv06VgwzRYEiw9GtQGigqDWrYtkh0pX
I8tRItmrqqzOQy6tgP7Ni4QdINsqVHuiBT3QqplJhrRMp73A9emYTaghcItHwM/s5LLaA7U947nU
YVcL1/Kqwml492xlohh07Qf0fFYXwuEvJ55X6dwFTg9rqYsoA6CCLGqdFyFaK1XwBVKyCGkYL4nP
4pQvz3qBy8a/R4a29Hcn/Hhvq21RB4DgrPKDcrZNatMha7cRJTKBrU9LD8Ot7ee74UXA7vkjHRN3
z4JUyExSC+iKKOaJU3J55lcBS7SA0c+QsdKkXsI0TeBhicH/hClr6JSp8zrqgLAVBwE4g791t56P
GqtoSKmKM7x99aLDrtpdpYPC3O2V9psWU28BmdQyIshIfm+o6O2zPB/mDpweaMZRpcFbqrUkB1iF
fCFM9+fNg2b9byfBPd/7b0dd5NKIQTzaPaTGynuP9/vNvbKVhNpC4+StJG6JFeacHBi2VKujk+a1
HTz7J9EDi/4EIiJJouWgZWkNS0GX4Ekkm1iFUtR8OhXPZMyC4yYbCEBM04WwjpZO8XcGTD+1HE4E
LqdnlS0KT/3Ye81+QbmP0rI8aOdyepnbH14JPamZ7rkwlAeB9Gf+nB1s1l+QpphLTbRKEJHcgfVZ
bihVcyjVfQzNN5+E/ZZAQqDtRNRmLKGC8XaGrcAVRDhodiJIuEefcw8jBYOpSRfMi9sjmb+DUbsH
nHhL9T5wa8oFdBiKPSoAHKf/kTpdGpwh9XspKgqV47ekY/nYlvJiePieyd4IuSDB1P8QkzHqkg16
h1zcliSQU6F83b1D6lwtTsArCDxz5polm061Ds3AP9KexV+FxIyY1F+TiFho2NSLeqQC4K72Znz1
N+HFQ4ZV4thAs3HhzIpqFaBdvNsydbzODarJchX7WJH8hXVKxMQz0AN2XsN8RVu3f+isqwUkKPJE
VL9k9G79xuhbfAticJ7+bb2Jy6b3+UD5X367S8Mrw+4+XYfgV8hJebe7abWokb4Ny6NVXO4HD7S7
2NvPoZ6sZ7ubz3HAFw1BbzDr0Synrn7ruBM17bVJZUUEGyBZLo5yyO0Ix52Ft9qgdXWeoaw3CcqB
EqbL8eMMWLez57bqKxj6xN7JJSQ0vyy9kvnkHEm+rBFzv0eqMy2dxYLkfa+V03+h91DsWichZ14U
pMV1nwTneYNjR377uiC0zZ6K9Nee8XTL9AheL+fh37uuexHTlCQzgXSPn21oxy7kQ9sEFJl8NdJf
7ISYEsaBFeJH0ZWHf/uLcun5nYd6hQ7AxPp75bzjry86QoH/bIGrpmeVFnuj37W+OO2Fg5ZC0flT
ILEQRzGhmhm3uOfnu1HJfVEQRuyjj5cGxUTFIuzEUaDsd38v0cJrQ6GgDO7QmIDJabc2tOw3pn6v
fLurl4aKWMIMKFokBglkM9/3Y/mhN12UgAxHxWdE9zNIs4NJrkY/kcwdlxu+44z6tIY1aAilleY3
JhOKVNA+9a3avl68fnfekYeZbkYPQrgtCbr3W+CxPyiqqkI5+xUaZFksgKyoYZGX72Kx5WxMyL8O
Dk8ZSYgalz53o6b5NarEw24V3N7SmopU6OZVL1eUV655buvjFSHVyV8Nji+/Rjru7AqmXFDME3Wa
k6HhAbhzgdRhhKkudsvLx8bvq2IDqOR7WpD/fsNptBYIDCGoD6sDyFFKIjLBHyf2kqfhdW3MYwZj
Anx9VtLZsjDeLloGycFX8VjFBeQn5GKmg7aA0J/t5RoR4b6XHBkJSwH5wsOo0psnNqTfQd+KKQ3P
SU+yN4fXVXMepeZ7SiS59fHcyfUfgP1yFHbPYW7+n9ljXuwK+dKl3YXk9KyN0tX7/fG38VwFxwDs
66/eak1PJ+UaR6KCeNU35ighNnSWQOo+33a8HN62KWQPgjKGAbWHA8ANE2MxIQGPT5WPSY/DSelK
LOZigpL5E2yDmiAbZEddqeeIFUkPZ5qLv7f9V1sgzadaDdX1QM++8FNcOBIEeaSU0HTSJMbGyVQZ
UXLxg9GOrMMMRbXF6Gjt6DPLWa9J1LAyTHYnuVrVvcvS57Cc4ZPBuJQuHvfrRRPUE3r86pSGyYff
2heRRryLXsCUCZHU5CFM2Zr43Jm37Us+a2XGnl6+tvhdi8ysGL46Bl9D7oSGhFtpmfmP2CVeMqqH
dn7CSddLMtw/zNdsIu82DtuA0WY24jZks22uAkiLfPdzNofwYHrIGU1cncgrUvsIxWMwj2hMAlZv
xSfjfy4fpVk7zyLgQV6KXlQAZpxraHmSKGOpevWc1LFD6ImEqp9OGsJuHh+0J+1oIvxsmYqAm6Az
L0K1FFLxzI7vSKdhcULIN4RW11AR1XVak1cfU7yak0WmwEABz2iUB7u8vkUQkz8S3V1ZgVosUbRh
IlnfezPmMSDhQg+swY1og/58xi9GLLn0dzBaR/CAILghgc7r3UI2FCzqLO6WAGoNL6y7v3WtSCO5
OpSY9A/tTbUAkc/N04pAIFiwQW2MP01ERvkl41O3GVcJgpE5pOczwO6sD0CNdEXRMDGm8TShbkY4
ClFNGEN2yYamE6flMgWeo+yfSj1vvQ6onJ45Y7qqB5mzdkMYRaXHzNuXxIr2SkbRl3dPDA7MRkI1
SyZZZDl0nTgaMX/iNIjQ3FRVX9zhVPeLYJDIeSIVtUd1JfP3G15htanSIKEc/uAilt5VEVmVMovf
fjWsdoHQhE/LpG4qAgOeiVommtSTmP9cJ0iW8m/1BNxuYYsftr7lcGKwvGyibGb/tVwIIKlROnbh
jL1CvcceaVvir3n8XqS41KTz06But5haeln+xnKSz5LAud6xX+tFbAq4n8DYR81AX2DcuUrDjkHr
H8cOwv20HOABMQ4eqNDtNHObyZMC6H/wCpQ/Hjsso1GkwMC0XeD6VCPx8rcWgIesyPrUdg/hDbQl
h/aDeYxMmtMDc7pAxC8nBtvMEbiFrp7V/DiIVh+Mv2YGCzKg8K2OgGG0fepr0LmU0xdyAQ6u8k4F
4rR7zt80NMKxWE6F28VQmDzl/vDuIFPaLCXbdlLYJUX1QNSnoLf0n3/lZE9am0dgltT3N/a7CvGJ
fceErJ11+8fLQqGpIEvtzdRA/u9gL5EvkqkPv1JIgDbOsER38NkPMWVxawhKjQm4LOKSb8cIHG1P
5hnNHCOK6tfHyvPDCVIFmR9+UgELqJNYdAkP4/okbPmMRtkW2hJ686NLm+2gDpkKGrxw4BEQWcie
3fWpjrE7iPHIsr/TUSe5Qh8vQsBo6DYNnxCEZMoPN6DHKzc8qPflMd7+ZPNEDPylnROIZSkbuJ3H
LhlruJ2u3olDRaOpODkjGe76NEE8vhqLuZNebA/VkSr6U79BRLrgfG2nYhVrveBeD+uNobmmWmAA
R8u6RN680ZJ5GBFkZhaCjsdHumiwp+X7XOXP8UVXhgORrl0m1ey3e1vI/IMmFk4SQpI8GVCaVbey
vy3q84nlETmjkTAa32aDFrmvfOs7rHa2Xt5+CnadcABb7Wd1vwxAAfySOTmy3Mut36PvLB/lb6bZ
vcPJd8br6M/1wkDJfjjE9FQ70QweloqYiJ5YpH2SCvHX4iL+gBrHnT9x3Kzyxy+HIBNVYCxTGAa3
ZjNQCNSRdq6sRv/OPDvFCgYvEAW9hL8vZErhujV7Ah3FIUaB3jck+H8BcK6TknBdN29n/fmxRyz3
YkU9RjDbfwg0zx2l0aD4OHSJN3rRzEUy5xb1YtvnF8zUf+kmhtHeALfspYPEcfetDSfRI9fBJ58c
iq35PJwW7kDVhvBsal6uCbYKz6RzTb7TIlh6SYn5sscTycnhIQK/1+BqlQtVJW7fldY4L2+juUAC
v2M4yKH8v1IxyIujYTXZ8HLJUbjknKEOu3+MkVsjKXoOdzVD3metCOxcKJu7xncTt6JmMtrjf+YQ
4Ym+r6+QqTyRL61ptpil3PSwsbYUs65UoXHYurCSa7ZN487879K23jGtY8w6KwgrNoOHTp8zwOXr
aGoUwTCEOfismb1m95FJYHSZ76iNmL1mcs4rZaQPKmtgLIDQLKvx32Z6jjDR9kv/aVJir1UGABHS
SIarjtxw/zeeco2t2wrxDtnyWjB3+cxvATNIfBSnQABD1PnikBjOlU2EMIMrn00D0UleFxGjqwCn
EhRpRiDL5sWchThwnoArSmEIu6TcmrpTdyLmcTlrxI1FwUubTBlgYqRyt4G9uol4UPn/VQ34rVdJ
EncifXvsdg1mzDIVSwIdLVL7c0V69oi7Bs+tHStuhTJ7xtwE4Da1K6eTI1YFKaACA8s2lEtWXP65
/XNl7PD5yGev5/R4DstpeU+u0pj4l7Yd/KEzAmiWh9uc67meoPjqce1zvjuYosjvDEQsUo1T6eOs
Z/p9Or1HN8AcO8V9sQ+9/BT3mC9JvL4JzIxWP6Ra2KtWeD2ubgH4XXVDEtW8PL8F4fpqOgAdNkFj
Ck2h0GXYyustCSndntcbNEDH6zqcbckkJVE5t5aY/g56F93WLDodqdiLUfjhdF48mAPZMsWysrzR
gHhx2UQyp89erXCVT21g7rn5GydmKBCZfnya2Eh/4xcp1q+TaSuAAwOzL6xm1u+Ob3T0RltBDJlW
1cVft0Qkc7Nc7SQ3UGvRb8Cx87O3uyi4MRdaQzmWSKXsZdWWGJ3Jw7wQ2k2xoW4/4XmScCQUdmuX
mF6gycKvCFYuDftSb0nu5L2qejYPSgCyGyzNDYphljD9WtPZhG9gF3uBc8+d3Wb56x7y4l7Av0R7
gQHqSFdEpjLZRN31Z0Wmlp7FGo4AHBqkqobjXYSxuPru2G/Kz2D1AYERsUOzrbfWuxyGiqK6upGy
plSR+t5EUqM2i5O5KqlmKAMWBrMyCGJV2MD8BBTRWfRBv+v8DV5IbEs5IjY9l4tfMw7c4KsOhYvM
29Pfx4vAnk5TdVzVnY0CYqA0VfLcEi6shO+g6B4Cnj+5KJFBnxxF4cZ9/tXDDV0ZG1XsVIg0bm6m
0km9DKS0ZcrQVyYaBlZ1wT3cY312VBb5q7UuG007qo6blbJBC22IictSNid/qq8qO8yWoYPCgn05
kBOlMFQpGbRVg/ywsoHGfXpAWhzfJjOcJE0ikkaPlMKKpuRXPNEoxoQQcyIZmJUgqdWrMSrzSQy4
aOoRKfeAzFIVz4v7vssJFiUI/afF8UC9aHPzRHKJKG01SqOFOoxKx7Q2+7Jaa7MM9kZZ/KeQX5k7
HSqtawqH05td/O3w/T9tRWzAlDs77pcdD/Y9L0GedKMmCcxwG+4j/+wlXh0wH9uKEdRhbNJ1wkX9
EYz2S+OQNVj32m6LpO7AJXotd5U0Q2GsxX02ep2TklhzHcuqa+9mldRfIPb4J7qpvsavFF9nxk4m
cO33MdC9JBIBPudeKXlG50LrQqkUtZKND8v1P8+RMEAAcIsubF/buRLqWXOSLsxDY0DMSioJiY9J
n4P6i7voTqPf5kjlOTQj+9i+M5QGDpiUfaIE1OjMvEedD2Ott23UYY37csn8hIGvJRPspKOU3etn
gEukF6JJyzSZhV0jaGlISAo2+33AVjzXrug3wqvg1NgiOknn6Y03cCq/ildQ0URQKi5d5kfqosSZ
U/1yN6Za1/eXRvtdfBJzoQIEU6d28NSc5v7awWaiOMTGoSc2weLy0Bwy5wRgbdMQdijZ2JSVtW5S
Np8mNypqA5hWJEhbkerlWBhFdCe8X3CmfuEFmI08A3Z58goBjhss4uKbyBd9RGnHbnTw0EG3igRh
TSph2dMIESwoB9TrO5HSXxPyt5w7K7DSHhmPoow7JQZRjW3QlInzQ+hSTLsXrUQxA5I28d+M0IWG
z1ikdkcz/EJCQDCMDxUdcYfwYt3AeXpiDooHaaq5Hb679ucmRCrHb8tZK0mmepyZHldAIM7apefy
sbeEJfB0eoviXRSf6JiNUXA7V1qZXkUt2YYDpwM2euqAhLmcTqmBhWckwItWE9zsdbWs/fjuPXo0
kLb8x72czfB9B9SyyYiid9Fn9uyTmHLGzN37pVdu0xtXf/31hiTlsVDIdr6dOL27N65OEyDwCt0j
2CBZ3fhLuvdvS/eEhsLN18AavZHWh9OUsDF+wmIptF+6/0vOXyLzkOqCDnNrR1mm0o/fXXNc2NAp
DTC2PaVRKLsLWidm5RIeI/oFfHhc2EbrNhj2uMVn8SmPClkvxdLlzS+Ve5b4qVPh2f8K83CkyChY
7oa6CXQ0QAuN0LUkdE+iQfbOuDeKC+0JEDSnxXtMdtXZ23qBO7Lmwzg/QV38IWFFCL3rxFC/j6qA
jE6bIg/FggENHG0yKf40gulH+Eu/RJTQO8LqXoO89HIfKWi9A2RBO2AJK1G05jSGxWAkmX40d2R5
aKeNWw3G9OeB+SWbuEsvTV8tcuyNBCoMm29H0siQ1Y49UScYXjvYxu4pquG8j1IZICHPhP4AhGFi
DUxEapBoEMPwrYudTnJ1Y/o0tt9kvoZUuLUOV9SIJe2IYkwQUObL0jCOglkChFL7YBwE3tqH5HR7
Sqo3uCN5H1pFri+zbrbGSqxmBk22ozKzFbwFS08EJFnjYG0VhAXLpmBLWdoIo9VUMAUnkpUDAM0t
eA3ISqr/NRI8Uiv01JgYruF0R0ZdgHL1VnKMMp+x1G2ij198KJU0BDswgf/xZShvJa7Op8m0g9Xr
sr/wHmu6ywdffXBh+W6YjMyBpuGqudK/65/nyJTvgOM84fd6fd48SMcfOXKr6nyDHBESD5aqHN/4
GytU921+C2UKN+Cvb3BYmysNpYtRXK1tEnuqkEgrlYP4WZ/mKkwuUrhOYSP2+zcW6jRo6ZVKn7gS
GfoWOCvLCoT7Joo60xoQTqpyp/jFPgdXEDlWk3/NhnUtBhW9P1EiyTwB5Wgv6hwLGUb7bOAp9ZmX
TtSvcsW9xuPatIFeps6qnvBF1y+UXi+OD3q4AMqK7/u8ZxsLDB1VgAodqgFrlviKbkHTaZgm4j80
ukvvaZvMF3Qsj+18CjBytquVFPVLdq7AQ4x+3KFtJ+FPRucVj+8pD09bBekN5rLzZIIEVE6PDEZx
9dHaZ/zdmkV7bsljeQ7l/Mef1C+XgQPXgsRwZWDVvVfdtMpTyLmxaqiGUMoYa27u75/TuXcv+nT0
tZSaFxlh5KFVcco1f0NYyx3BPfyuy4PK2uVS/NaXYRGBD0rD7MCpkPBAdGUaC+1En4HZEMkOPpyY
Rfb5SEPUEjwVQMVQppV7Q4QAyLHagj/oL0VwuOa8DOhygJHD3HGVEXVJUBSmRMCBIv1y9cE0zLrb
uZFWZwfE9w0Xy7YXbGj7rA9lEO8ebUbhZn4wYSX127rUdJwvcytNXu6cgkw9nPWKQ5tkX30X2Jt8
qOon7rTbRJdFrfObq6f5gz3hQLPfcbLOZraveOuVdw/0aS3bmVO4P9ZNHwyjsQhcnG5Y7pJgwqkl
WiL1Y9DkGiZENrcijMt5+QDzoDRVmyGdUfSIhEZy8hzxcV/57mDg9oISQbtxtD63VWcN8UvGwVXl
5paMknA7MGsqtjoUH5Tc9HD7wV7tKLB/nyoP0xfd6veDCWHs08QzSI0dSSyOhAVD4dozXIGo5/fT
olKl1UfEJ337yktUYrp16P/Ig5oIqzouWiQv7VwlsZlARn9AOnUQVRpshwHfbRHom8U0S7kj36/b
XnDYen802ncdOjsjZJGUm/CzYYnr2wQ8+/EwSd7ToMRWN4sEZg9rvAw/yum6+503r/AbC3roAd/D
9vQrQ+6fVT1jFCzQZZA2MtHjpvF3BLtNkb4xnJfgJLfRD6J3tgaiv4FSz0LmyQ5YIpbJZQBUTUUj
O+8H59DAHwadia4Z127t9CulekuZAkkT+fYhadRcEQksqMcfN/3ysb7iA6ptlZzYF9+AOpAIltlT
CeGPvJCCu7y6Jm7NCj6ZRx85Mv4ilYtvPILBA00AmCmzWnN3TSUSh+nlhwcjxE815sJb+mGwA9B2
K3sGNMcnlebRruu/H3dyCyg3szzp+3x4fM87H7m6Y4CB3f4Qj8ifb5mbOqOVYI0vCLBZR2xAF/AY
ZZe6NpNNpG26rHYDHkD47rSDXZcW1sv4xRn5M3RRBVlAlvBJxV0QRAFp/DBUWTV4gRtmpq6tSKvl
4eAXBrs+CCO5Z4fp3KeUP7E65ZoI2e3f0Ac+uUmlPq8+SjnArcsokQDzNBF17JopYp5Zh/rYhz8h
oySIefeS1m64hqpw1/svMbKwrUilRQRrlB7iAG1rKI4R6ggRwsI1jzUpEehnRDPsEl+KWbxEF2lF
YnCYVhVeEQWimz6BK2Jx5GAwo/G+QeiDl5yzHCItzJraaQOL66n6lMOzCT+sT8M3AqlWn+jlbrcm
Oye/G8QOlWOn3YCmIoMxAd5ZdrVIz1j1TkvlGJJQ7HAin/jWX8XQDfPpa8kOqzqMTD+i6/2Gv/6i
YTY88vQ490PC861tGMJLx+Ck6l99XcZwUPSwl9vFKdkez3AwX2dPrFs/c7wqMq+cwqBFITsVYHm5
8rz9LGDmT9PW2mLMFRyoF006ItmpenRD8M99wKe77mHLGeA3VxsG4rPxe60GYqD703LXhj4E8/Ea
mjIFlSiPUr4btqOyalVedAid7NSHoAtYb1mTHShOSpsYibFCarBLNK3G+aGnfU6mvoyu6oiJEvuV
zeZ6P0E9gP9J7EYFgQAtQBLusyzNKYTLHd4dagJaaUcjMG7P9TzkMr7Z+68rctPfzFZyqrCMYaOB
TKcW/9QawOpuUgpYgs76ug6DQeOOP9o2eRWl8JV68aDfvNpc0eSJmvitWi/Nob5zTqvl9m+DeZi7
aGlaGcfDGp1VHzwVG0DddtS2ERehx3Mc6kPxE1c6OTjmos2hnXqvn81FqXabrrdwM+LkNRqLCqw1
hybTwjuyKrqgzJhiDghLWTbZY2TB3t38WpN+49Fe0P1hrn+BIlOacdkm3m8di3f4NwbUMyhyibF7
bysiJCvj14K0996Uu3hMeqonMzPDaTJal5Ww/5OnQaj3ZLnUZwD41wJo2YAbp1reVAwCdBvcEapl
5VsKjLEM1oz101GKzpoue45NuOgpaFt5sKRbmtn195ln+Nwc69o1ItDtGHXGoZyNUAecX14fSVmg
nlLjZty7EYmZW2Rqzr1J/B428dAju+GyK6q/hnNCo2m6d48Xy7y2At6fjI+cw+2qi6erRKUQiYoj
jzS1xOFk/jl1D0n+iqD4a1MTZH+w2rt3V7e/rN7YhQx35QDDAVyDV33VGUnGEPniwXbgebClTpDI
l2/T+11iCkgeDkbGIPPildt9CwwNYe+WkQXWMXDZKO2V0jQvaZ2cGgZGCjPVGajrQk/vtTdlJ12d
wdx9X3rWymZza6DHkU90rfEdHywm9WGbqqVWlPhDPZ7iOYuh4hx5quP8Pojz/RZ1S1ep7M0bH1Vc
PgNkmlCD20smv9hsEwDK0VmzN4xm9CdvSohOEZBblDm3INJDAN6hl7Rm8GR9lt+3QBZ4AxLO8MhD
EYNq5u8yJh+a1WiPhy1LnurmocBN40scWodYavzshIS1/htstrVVujUWUpiSiRc+xIQiEnccJNap
V8xuUXVS4Yy4+l9YqZWDz2FCfGRWbyUT+hj6GL9mWpbE5O9WajycMXWQesa41gGR1+ksXmYWRqYo
NNcyuejpk+WtO3POXiJU7SXfIBmztNXun6W3nBOq9e/zftRejd/Lm9bnAZ8kfrv6jPxZ2osCGbns
gw7y6gYAmkM+4es5nUbNHUoApDVQDvrjgf+J4Zdy4FWjhm1zncjrR4/rBOw6ukeZJTdlFII22/2M
jpDAbyyTuSuiuCGTT1dYmXHYIVwRk6zDUgoRO2y1BWJIwozfY6wJR3kIsyDgmr+SNz+XO9Ij27Fb
qUB6cGHHQnyWunwGS1ciHVy9/danKV7SDriAS7Z3bUBm7na2Hlg8ymZat+RyQ4XZnOTJZaA6SBzN
DU2qFnejJNu1dTxWovd+yyvPT1rRiDjGkt+ldxcisP5px0/PHUGBn4/HPnSBEuK9izvGwT3isUXT
qx+1REqrWlXalj2pXJ9uCxnr6FLgk/MsqQdgnd6u4R6DImodQ5nidbMNdMBgXjFoVfmQM2jMJ3Xl
b2yLLzrzLpYi6T/mkjTHLwpeUUIXY1qkSdHTE5efxZgobNlrYpLgPPRDqa04Y8tzxL8JpRH5STdz
btSKg6N/Be1tprpqYwUaBp/LgjL5FgygdenQjb77qCx+4wA4Lz1Wk0Sh9fRQ9LCQ7RGUX7zK0izP
9zaKPrJjGrJIprz9MHCsvidFlQYBjpetfDnVGGBhSOc/vpDke+hm7Ct8d7cv6EJ186GEQJbsCdWQ
pIflKVai23EV5F17DPG0QQu6KJJ1I36Qq6P5Oj08Ed3mUG1A4BhplzZ5lZyKtqc0hp4v1V3GMJy8
tmqcrRA4IlRaLC8RTsy+UDhl0ZZKYzQslP+ATa9vmCHMkEfgOAN5RYsNNT25vSTmFmg5DxgUBwcc
vdlhV+23kc3YwpWZd7ymWRPHG5QqQlTJ/yZ6++Mi1e6YHLe02gaEzbRJpjNjPHmAJL33RjFnH8k7
0nCPeri1+jRKms1TxAtC5WPrNZWOru06W+ImYaBcNlTvAL64AgVbqW3h3lklldZKcG9UHhBDF/rC
tQJZGi95dQqaMIUv1aHlT/a2l/7+K3nSupRcHno5Jl/0mhOKUQViYysKu39/Yyvf8kPs1Eez6pMu
0cz65SkaHbkAN8S4k8kTz3EENAC2QXylCLfJ+IimFpN0YiWrlnAh2CP3GJdQQBsJ41ffWvf3n99a
zWmxD/k/Wa5vTjWu2WLqJn2F29MduS/B7nB3ciAQQ0wAt3RPVFNTFC0U3NCmNf2Z8rEzdqL7csPd
BPF6TRKixrdziF8mwwFRvVWB6MoW6S1D7S9n7qZm1x6C4QCyl+nNRjJFBQarlnuCBSa9YJlBVJ+C
zm0G7VUrnObaD1vQcrKiYJfJF6T+3HeCsxpt5fG4Dx0tgL9Hub0tmW85EAmTIkJQloOqJY0cFdnL
bTva5p8rgOCnQGR1H0P9QqDfj7uXtZn+wXLuch0ReGJDKyZeWzgszXyJKwolj7CYdvD1EB+M11mw
FXfCDdJOXpOuzfHhDuw4oI9yqIgGYgSqnzYJHRzuEwvglwbWT/W6GTU2EezF+HVgb0Y4HjvWGY5L
ujs0s7VP/NgKpdn6z5OA0rJ2FEPqg4iYoWlQn2fjQxLUafjAbmAsqjQsYXF04QHPTxZOY6GS4xI0
tprTmS1uW7zTGoGs09VRd8WYs9jqqJXB1gHc6Xj8YAp8vK6xGE6w96FQC/DhjLvx8jzFF5Pr76Ua
5HK2M2oMS27NWdHzZ3P32Up214eSYRGHPdrJkc8ezVKMGRw4piaSRxkxCJW7JqSuQR/oRbHGiGU+
dSgscVUqTOSs5DHtdM6cWydPRjRRMPqc5qCQoDyTz2xRKwaZL9oTPWU7nxopQ6z7YWqgUVU9RXWC
10PmInAcMySuJIgfFR0oPa9gM60Rldoz2BJK3ZHMRAi+bje24wtDSKGYXvJqp8UyabyqThfgS5gP
4A1y22fnSBUOC0dWVKhUc0GKZGkVDk9iW9wbyQ7SEgYbejp3JYI8jKjpUwrPiCLD/xISxgPmffzc
Ky0epwCLV8NiTG4+mb3HW41/OZuvretYXnx/YDllKV1/Aa5Qi76GeHXWeaqdmIa9GuHo+X3aAREr
+J+IVIq9pd/9+0bQnRvkiHRXpcOb5UucN8oXLfI1w8YsnS+ApexhbzBvWL3kLnwbeRDemAl0a5Lz
jHpQpb1yRqGr6sv9OZRaOVYap/51MPM2iFXuOje1Xa+L005MaLbn3s9gStPmEMxSODdI5EeEB99V
gLQkguj7cGog+kcmqgLfAvPETZFvsDm4P/5m9hG4L1Ie2qmEz3hFxbBMqRSFuRDoTAejkErzdQiM
FWBC2KFsj6QR7UAXbDvPt8iLmkFFLF9fj9JqiG8VL2hi1v1fXsIwitcVrrJvA7lY90TpNd3vlxbO
7BbK1Nf900B2/1/FjVcSaXa59j0+15i3ELAES+kQPaGcmet0wq1kLh4EF6SedvRt3UCwA5IxblkG
dpzZq1CdNdByBWQrqJlaFu9iBwAE9nHG4YGPBX5TW8Ibkgm0KSdGh8MpsuqJUV02tuO3Sr0+EEzC
V9EctJIqwfCLziGh6PtLqDzzy7xb9C4GgeqBRgJER9MAdnM47OyFtMdCVt/HmR1zxJG1Hz6eqrun
HfGhwDo45RnVyiZT6QFI60JFR3WuHGG3qH8yZLLyHc872JYiaibNUGe5VBuhdesf2nVSjQmTbzY+
dee9/EOGnScFTiVcucLeKx1krJ1n0aZprzk+1qpeamaGPibAsUdJzmJVtsZBe/2x1ESNB3ufjTSk
LsRbLRzALapwyrwUo44hT9R9wbDkVAuNgf4VHYqkwgzVZjPvS2vzrB2fNYmEfd3LSejk0O2RaOkZ
s0FTDlddK54fo5qxDU8uKjYRhoMTCPOjE+cif9LoAsn0BDFFZpv4oTICx1pmL7r3Whn7KBnozQoT
v4y4MpGJcA48aD4LfDelzGfe2TrwLd5F63qiMN/M4xdxRMZyRdklo5QINbEk4Y/iVYh1+F8XoaMl
sVLnNI6Kci42HhpYpW+gRJYYUPE8SdWQmypISKDauykpHwO9btZY7DvidBmPhnPVT9dwRx9sOt0a
wc1U+tiEhOUwHf2nj2H9dwPpu4s06zUJT1U6vIQjtac1hmCNLOozGAAlsds9K2IFZJbwRC8WqdBn
ssiqryobIRPMhphyWpL6F4xuGZKIfTLJbtAv2EogqTuORzaZuhXJnVSKUY/+jci1GeF2Yep+QNL7
Z4QECGK140jzFfUDR1Y1dToIXdJGAFwPhc872BIjd09c+m4LHBqAHaybSw7tTnVILIb5jEtzcEZe
6Lc9Nre8pYnRXUJf7KUa5lpHmrrgh4coeE5MvhyoZgCHkAbBu7jks0m+18IzvV2oqJcHjPv2YNAJ
rmygd0oEDWby7LZfdzMBOiluAQGQJbVmC8N+D8C5kqlOpv5vWqrUMLuGWz+Ge+XVk0PpTIwRjtRd
ua69d2waMB4XKU8gzTLikLo7I1ffaMDyVZWJ8QHOunExx+q+kuITsNZ42Xp00N+btUjCCDLGd3Hr
l5zR9U9uAK6R6+9VFOhJZ/QImeqGtQIVMBu6RMwCsLo/jot2o49EDTDC8YP3a2jG9fBj6PDeGxzT
jgB7idum8HGcz24cv8yp28c/g4UEhgesZDxbbDNL64/MZtGIGiY+Rx33C+XLSh6pG2gaEfd3QCWr
GMnf5vOTTHaif/Uc3bx/8YqnHWmf8qc4fjnLuyXwJEI6efw3iy9ohBYt5EvQraW5VIbQ02WqKnea
4gjc17zkN3H6KKVk8qszMWOKujhbbkC6gQcXkweZ+ixfZSvUsKH/0CBEcNZwwUHJnv2kB+SkhS+F
LIlqxF9F7FxHSit5/BSSSkBzOnVpJO20CZYo74rwcSXBoS1pn0d1Fvc9oXYbGkoM14+wwlCE2wc+
p48OjXKuEce9wLolo2BOC7nv9Vt78kUBneDwL3M+kNTAH07qHOeQH6L5AMJDB4/g8d3i96QwvV5C
CdEG017HlXfngoGDNbopFh+ZCgi60wpfjFvM7v1rycifp5XBLb73a06C9iPshFRRf4nUOmr0tggj
9WExbi3dfJW5OhiQM0IB425zL8r6K3UrYUMywmt6+nSflvtwXE89JrjYnO3MQU+qYnBTuj66uZNv
KGPe8KzlRMXen5IEGD3RKwQrqxOGdGZ5nOynPdPYp7iaQmQEyDoEEsF1w69iDJwxCq3Eb+zO8/X6
bcTSPXwr4ubY4HPLkTLMU6TA3awwfvLYFPbpgLuc7jpS8SbKcSQL2Ih7CTL4mhq5Uj3AvRIicudY
yR6lmhgOXGCQ6iWfMDyYv+hZ928Lhr/KJA5BQJEmiFO4wVc0zm6khKyHfYQnPCpDJYJNiBQe4pWJ
ddbWSCEbI6FSCIv3LBct7HbfHILN4CBJ2fYVzIYsLd0NXpdMYQV566f5jtp92EGsFeUxEuSV6PBV
LKz7RQ0jW7881Z8uZuPbG24KVFgQvcQvRDYNKsd0K6y44FoPKz2dnUXn9pG5iLXBj71c2lRoU19G
pyJ/Md5rRJJS6nyWsKBRM77LK29V4Dp+tjs45GNanx6laZq/4Lo84DDTY4iDiqxIbFz/+B+xAB3r
I+jZ3DcFbedqhq19IdmN3zS2xX3F1hGYL4FYJl1JAoIWa/QrBRDc+nP/Qrt9CqUQS0NrMIW0YD+h
aqnrDScSzD65z6/0DgLRzqVEMoblyZHZgd1dzf8WOD6dDEOlOQSvaGbNCvhG4CmCKab9LIVeBUCL
0MtdBO8iCg05SMTV5tzTT7cMVKZ2AR7iw/ogxBAtgtcoHm/yXtIhtw4UTZTyx+O3k85NUCVGJ68m
h1heBkR6qZfsu5NOcWLhFioJeVXhfWS79MpV8gUZauyTW4gImCoL8/pl2jBm/dvmXyA+ARW/GChV
ykhXLPEfI8UmeO03BRpcXS3vojeFqnIkZqeZFJ6SYmPM+UAxxr9KbOfIHXmpv8F5fDTYDx+gF3hK
WaX0WYy1dzNbLdvZ+fSxrfG6k9lsHggrS2lWePFmBeAhOSbmU/A2zVPsayAYo3ZI/U39Hd7OvEZA
ULvJlsyVopGdtq424V02dLakAxLtignDPwGIXdBfoHsRm/lfuNuQ/xzSKHNlj32tVRnuPHPGB5LW
UnPrbDL9oJR1eSR0BkNxQYCS56XhxqbTKzcpkANCT9JpklqAHSMwSX04UxfK/WFqgKaK5ULoTWdL
RtjWVS6p0tvS6X2iRTVipY1qEI28MWtcIAIVI6ihmyCn6sO3aLvoeM9ILu1BIra0TedRqd9ESb6D
lT+4VcxHcdxoszTu5HO+fd7y5mK8qVWevWzzDnHanuCRvQNs9I1SAnSDC7BcHBnSpTLmhdMCBVTD
MDosKamTQyQT/IKgXbyqJfKSpACPl/DOcoAtTKLwPG5GCyQ4XSQ8P7KSaivahQ4Mb2n1YithzgKh
7NfPZV+VRY+rXE7cQ92NuP4h822DsKQXFTlhcsKqw0/DR0MaY6XmKk6lNtO4/65wl9ukgJNQZ/qk
y3pjNt8Iph+YHcvGn0z+lKtx/Qfi1iyL2bdYK3dvTM+ta3KmrQipN6KVSNM9cUjZKpSU9JkneW6A
c8QElSyQX9MuGesck8Mxpt3/hFH31hTvO1PdzoyIB7bcYJtX8lDqh+xtdLaYcd2drnNKbZdSludm
HQImR2q6J2BJ5B3vxTBg0jDIPX6phBx5iKY3HY2m298lr0am8B32hwG5VrHfdWZOu2LAXHtyqrm5
bFfVD21qujpAhYXejfttLOLysPtdxuyQDx8O5A1PAs68nRZQMmyvFMJeWGgi0qAjKQPxEjldQORB
vDpaICHwhSQhjX0LqpXhUwmHj10DtOSIHLWL9WTN5yqi9qQ0m0waovd49iEzA6vV4BRXxS4SCzMK
NfrTXxPyFi8Zm1aBNHtp+uOPSKBuYLaRYIHdcn9Vh7GVUyxGbxbO+AWdjCUlWJeqjN2dR12i1H2I
8H5JcqIlxdvEiPsPJYDwmNerRNQ6gHj6hAxsJcSYI6gwy3cfAAAcaGUbZw7QNsTl7XaD0snkX/KQ
BVXejOCMfEFUZeTnn8OpU82DY7qUwkMuO/bM+ajK6aoZfuzXnOcTGOpwXXoGNOsr97UH7JxTV4Hv
BlzGVsq+cMFc6rm4HFaKTPK/PLoj7jM4YNk7Uc0qGytmpbuIwUP9TLbney2XVV2MdR5JNL6n1j3X
PNRviskbPfJBKsYGr8rmq8Xopej5GJqQ3rWso5zuLZO6nIkmQm7dOnWfVZPzdUn0ZWsrs57mKQte
7LeHO3OQZzbfYQOMeYWOKWd27zg7943/2B8Ot6wSg91D11ZIERMgy8ltWWhIDq0MEqp0PjhgmuFB
po+LOLUYaU95vtJ5UG38dM646Ja1FJOgGonAArTPUQh4ULTjB2NEmdBEzMTKGwfh6nCZU81NSbFQ
GnnmkIbv/O+TnGoa9rhjcThwIPtkup59mOnk94ty2CSRiOG43N2Ycxqa8/jT7ykYky+2IH+8HiIR
cMnyl1B8WAO9mR4Yi4w66tucopYG0EoJz5kvnsM97Wl/i0iswmZbCS5+5wnBEYQC0UEbbYilbFwf
31zj+hGM80kw6CKlUbBx5BZ8LMa4M6q1i4JDBrscRYtowRJILYSlpm/Z+4STcbmoW5/4aonghTvT
c8dLpIFXC+otU8MNqdS5oYzFkN5q9M/9btQydMLj4goTQ/m/A+OxQ+A1upgem/uw8POUWj1YvA9A
CWoT9VgAOmP4S+OBYZsFQhGrUh6hqi4jiE64WKWaSipNNVAL07g7b730/6VTkWsUu5ELIRYjTmrN
q+hDsajjHuGwLDbSRldZO1GjXt3gGXmGO6ITEZ9D556aHnmADuvWF55tKeavtzJRj9LTH/w/k55e
4aDGJvexw+qYdi0UghBlOHm4cWqvLH+rEjDnb7QNlnXzoTTpTHs+7EcOSM/HaQg878qtrYbCJHpv
EKTtDLmkbM1QhmWBWvdPhM99ahsUsQyJmtfm+1RqdL0EuzUMFm/8dbF6xv1a59V0kZQLpLVMR1Lo
p1UKUCg2XCM4IWNydMlPJiknpG8ognD+C4A9/U+qReir1YM510Xa9NQ/HXF6HcxcUiMDddOy/inq
Yw3UbdoxU7wEKIj0xIzKSYEQZHDovlfOhsAv/CwKOBHj06Vbhnp41A0AGUF3rcz8rUuUAvKy5yST
LWQlme2uOTUcfjV3PybjcOrD1mJSXYof0aZdbpMM0VqacMjxhPNtk0iBRHFZDAEKmilUrkfMpFT8
69BO9F8bdEDsW8/6KkWbVatD4tPyMzJLCPvrwGYgvQsvzZJeo3dJ5kN6ef7b0CR0CJ2DS8OZVi8v
Q6w48sOczswiv0uB2WhB8P09jLYM5GQf5OgAHWFzNdYvuELi8r7/JXaYb/CORfw9So/Ck5qM22nE
YbBVIbOEJdqp5edSoXXhL8cSNoF5m4mmP/ogwAOSgIDvnvM4q2aQb1KrBYYI+6BGMb1OiJlM/aqU
N5wBD/28tEznOem72Lx8ZTdZXoFxb0nNjnfqstowgfQ0VLehsh0SeRUEJCL50C6Bxqk0hxkVcQwP
UH9qzIjDmV2RPkVr7vXeCQ3nITTQGxEfAYlUQ+XZ+bPaH1wHW2G49SkZZ8ydLPolgbNteXjiRxzw
OsFQsWxF13lNITnGIKxlvGUbQtFnRsEZDIvKmxWUCbfo1dcgcApT6wZeQbmOcWg4w0yY2Mu0UYQ6
kjLRXl8OXkH0sQHGT7fiPAveRUplY7Ufz9hOBjcWLI+p6+c3AQwtpOIzxAsRJfJavunJ9c09GH3i
JSb2ZP+Fb5Q1Q4tObKAHeRSToyAO5kE8J03UcP+owcsfwnxMl2bSDOU48e+nZw99apD4BtUmzQSA
8brxiq5DRruWblcmouNc8OKJXhbN+SQ8nPNWqk+26FmzcK/P6O0EjsdxAGMzryRnwKW0Th7M32VD
g6ifgf4lRq43ZyZ4jwjUJUgjMMs52QznumnJLOK9Y0J/kzTPuZpg1c4uobVSF+iPDYX7VA+Sgd3h
yO46jBuE7mmcheWCM47v26MF/6MDnqI5+pY4tRSDcOv1JNxmHg53rPlvQPSrzN5KJC7o4yy/znj2
TqKrF7FS+wJgm1l4w6pLB1Zws/UREK+TGvDLUAsA1jc9Ea0GHBvMlIMHpNo/Ob115dTFWTpo1kHP
DdHHcA7bl9WO87ROlKv+NI7UwDdnfZ42Azcni3Bcpp9S6dgpHXJ8vN/106dW4OTLgzwJ9WpbqWlb
4OKoOojF7RAL96RPG6zNUk0FYj71aXKzi8xWwCXPe5Yc7ynSXRHmyWVpU465j1zcMN2VJboEwPPv
aBvY5KZbuJoLWOM8A4JkCdFcPpz3ZNFNj2ChPEWK4P9I7cn/dkJxAcwEDXEDQxpKoeBNyRc2rlv2
RkswpGQpL25wbx2nwbHMwzyaEYpLZsmB7yeXams6GD093s7JcRuwVktjpkrKvfMx+x6nSMlCCf41
t3WAboz6KXNcfaIX3H+yuNuKGmMlhuboz4hzqV+EIHgmD6z0e1JsTRNzAOaO6mPPHYRuaGGfjrHx
y+Wf/kvxtbmmz6USzg8rx2et1wyNzy0kUzTDJIxVp4nWKQ6wqkWdCmnf1eyS9dY3wi71hHIsL4Og
eY3ouTucDtVdBpCio0N3UO4eN9cuesinoczwutJc4o8av58D5MI0fd/D2AmYNk0c+yveYBGKIUNv
iAnxfEcyp2wc3qdJ3Vhv4cmxV1pJNWngzla/zuk/6T6ndJGzrpAUpEvzQhoRKEsYzviD20J5nWSv
50h+FMlQKLLZu/ZqW+9UeO2LZKUsRHIg1QMzmHFITzT5ExUrLWeMVO/0gbel/3VCQ8lA8Lvs5CrO
MZaIo1iOTXOPvqGfpjAAcru9JjPvBOapZffImTX6055nHaYsGm7lPXQcGUxc0XSy7iJe06ywujsS
8Kb9HbfOU8+xCJSoymuENJcRHIjtrPyYCXItVPz7Sj7Lz0Jlw9/s1GpDpuoQovJ2uxTk3dQuZiCp
jqGrxUGpmUtiJTxWt22dp/YRZw8wVN2S18O8AsPfN/eX7ndxqpnnOznZ76uqif/rlbqlS624tvqJ
roB7n9+iR24tu8EgHV4Uo3XV0sQ88A80WHTNP4MMmN8zaqQmZB9u+bMNDk++jmFcAnd02jc4z0u7
nn20DtMtoLwrLCiypcVJ3DBjwHO71cALS3xZ38knVof/pqwlP8jWe/Ql/+6yka6RPdPYOiQLy7TW
owvsPizmQrFk8shuVyTu0lEhJrl7bePFyVzNw2ZT6v3N2CZKBvaTmD1SQq+pKMvNdNhqwQtiNeOS
6EvSayGkuD7mHHjtAYownvHPjIpNEkfWm6TYlMhyRfiRcNnmgLka8KNMSRghZ7AqXMPv+Ujb1ezI
qNfVFl+sf4prU2bhZp4hr330Wa2o1GerXh0UF6gAq/noAbT2jluXRwbC5SXf+cq3byoXZGyDvpTf
MDdl2kKIwwzSx2OLQWs9B2QpUt9hGUTtQynj/oDZTBNUC8CasPkoSlxe3aqdkM8LTixIDU9tmThC
q+Ju9s1Tjb3J9yFgDV4LDsUC8EQDP9o46a6RULfxc16wzbGu/P+txSMEogjOCzqDp7rc8LxXwXST
75e3jHmbPTuCsUDt28Spl9yuw3oAWgENPvNf2/6+CmcUgACPZxQk294sZH987mc5ZaIspfM3ugoh
eJNF+OYqi1DySMEbaZAnCsUOMB+AkTISm+D1IeH13byZfCpC9ubxZgN6JbKBriMtUJN6bUHcE1+B
GmAgKxDkJT40Dr//X0yrFNTb6tyaCpV6SGBPOTlTztM664xAdy5zBOumlZEON5moHc5wTO/2svw+
pZlt21cEBjczZDMwB5sgy6I1ugB5XWCKQGww6G3yBPWSFB6bM1ymcfbaH3ba0RlujulR0a+r1lqW
tJSY9CucVjDBt68lNYG6BnQGH0agf9kqkwCa8Y6VS6zgPfEXGAB7iBn5OzkaSYW5WwmEW1FxM/ox
XQOl+dY62cb5mbZZGT/STO1vfk/ypdZPEjKKjn97ucVEwiqlkmNdEug01HmOYWGr2+uwGrsCL4d9
84CbrV7O8YvtVgymmnPfOcl5q1G/kHnWH8LRSJvSqIAMnnwTPcr4SK7eaNLoqJRu6TKpCvdm+KY8
eMl7m1V4x4JqscHzNFWUnUcziZKfPBTCf6ML7jiXMsAHy5aQBl0H9t5WvOR8OQQ7ZI1c3kNxMPh3
wDhlEg4JFAZ4iv7+gPZqZv4rJaP5IOr4qa75ADbrQwUq1ZK3vGNNLxguzxPEKNRO8hotJq3duuKr
9EbqV/N6ZjDIzF1eV6N8umN6FZvs8UTs0LKhielDlMr5/B4GpLM5+siKkYhvDZSGrR7kpcBRpa2k
P/WYkKj/9lE2n8QlThjjkkb2aDcGJpxX0Wkggqzi8V9mTLJhjZ01uTPkp5N+UjPQoUZM91rVonml
yBgKsfoH2+z0024UbL1eovcyF86/zW9Ew3LN7ZJCzglCqsqS+7qwJeTeGA5wvednTXyz0DP/nNNC
tVSltivpheIxrZbWJ2/YxW2QsBMM2IV0o6iNgPAdB5OKCBazeCZvZkkDOpfRLG1IltTsZojnzwPp
617qjv9NDOJS/hI6KfonUoJ+126gEI0pa693mP5xmzdZ5B9TqCOU31FfM692D0HZ3PvJXqND1WNP
qFmDgfDEIxJ0dtJolOnn/hYmZtXQT6tQweyxCBrN8Ik0hwS72dctlaSLYL+vW/UjEsQZUlSRE5X2
nzG9gKCdkWocUClUBo9wW/u3PgLvqfAx4XZT893g8uDebfai1iZDxCceLyhfWHUQwhlFnuRrI2ES
5cOzD7Mk+SGHVprOUy6bAEiGXDB5P070Vt/GEuNm2DYAtUeUFh5JT4UqMofHk7HLZatAxRrKCOPB
8pbQHT5I/Fw+Kr8ZTQt7qe/gslZ4lgv37XL+bBJ21ngsnfWLfrWbMPxNi5f6evBJcf83EsXYhH78
C5tt3oHSq/d6J2CcN+wmFxymvRu1Qj9zgqkDhfQpk9bUsfVSpgCWIP7s7z8TI61yVWnt85xCCk6q
9s09lI6ZsXJ6mE0lB+OS+yOi++ccNk1mXMgTLoh/77Cme1TJVme25UlYDYVTMpJxlmdJ40gPy1H1
iRrgNMLDNJl14nuE30eNbo49YE2KSCNSOLwmsp8HL52MNvmaZmFLwdXwOxy1i7y7EBiKrJGLbwWc
JIpp7evI9LhXwwsl6gScH2zdwliGVS9dLTMikOrefdwD7AXRTqoEHv3gmmdXkAa3CJugccPNsF+0
/OauWgGMfoavSfVerlK82bqJN7zx5niRVR1t4WHE4ZwyRGA19WNkFlY/TWLlxHlQAdKwi0soLq8I
gLLVmsmJ8ak04QpDj6Qe0BlnKDTS0poywduLPAAbXSSfT4K3AjA49kMCTUg7BVieMAM6hISvbthe
44VQ5jZaHhJPCReC/MkMx94PKOljZZaz49ICUh3iqeLoWi5cisSBnxfSMOJkepHQHy2zmacTT2Fc
Zw6YJ4fUSCyuifo9k4QSbV9AwBl5Mv/h97jdE253zEvTWYg50Huu5aOAAo42r3lOQNLnbqg1SjYZ
zT/aTjX7TbGozeXkOG17i9+qGDEKmqkiBnNgnb7loOjoSXu3XuTF+XbQIYm2L9+n/xcLqz7j5QFZ
8Y58XNcSjUKE9jDjfEGQE0jkdGxgSZ0zKVwUJ0z0CLAn699tUTUS5fWk4oymdyZDaC/OUmWNGlPV
wlFTbT863BR5hRceptJAE2Zwq7m/YG8IMmozC6ras1rPOepJ+qYMnuD7ysVeH70ARyg7TisMkue9
UKwSewIC6JTsN3pVLzep5ZMyfrja5oDKBg6pWcSoX09i/2NbHaxqGXIDJMS6NkL78F8rnHAZCsar
2ViEHt82XvFOKxoDM7z9Y7Ctpf2JFVPRcmO4/x2rIPAGYWMnHu/IFKn49FqXaQ8KMmFzo1hTqHg/
KSXs4ObCL+p1xS5vpN83+GlBg7U8fXsa5KryTTYipUbGyFTRNWrfQeOjaKL5Y/d/7jPkRXAKk+Vq
aiUwbKp8v11iVxxQnn3Fp9Pj++deJOVRXDj+Jy59RWbhsrWW42lGCd/lAwwJVcJSL8OsxHYbcsQR
i9Mz0e6AKWGwr9PKqML6cb+HekJG83Omi3R4A9JLwr4Iu7R7+hrZy6+p1juoqCwcaLg6kqJLiNHr
vDPhpJ076FMgMi7XngjHFH7DSOffid9D/lvl6zsyAuP5+xt92DPubmLN7ijBt46f4ajv0vs+Eihj
wljdYizs2c5QJrkw5HqtOTCotVS+t34TUq+Tr4QdOyWNgJN94R6WdJipmbb5V1k3wEXyC8hPJqMi
/RGvMRDIX1gd3a2I+FHEenWmdihaPhGVtHhPVRisVll/0gdaKi6XUhPEF37XUTQZCJof8jXn5bR2
p1dzZTyAJUkQB5g+z2i+ncDVOxamF1rtNla8//Z/FAYO23/odvIUh85Dg28h/SYakHGvyHEYb+iC
c/cdzgyhsU+axig0A/btA6x7C18HJriG56X1V1JTK4/bcf4HYcEQWwHNEhqw8YJW2LdHv3opu8IP
yg9beT/vWchpfpr0q138nNuCKoc3YhyMTAF/IWHOBglMzduWRVJ9l+HeMQ9xQOjNULaLtte//LTX
8Yj0YswEriWCSbDEfIulyXNlzuAd674a0JNMkdO8ndSNxMZNDtz7LwW2KlDcTN7Y6ECl8TYxxNpd
+8YJ7TfeO3oCfGTMFC5L/EF+2wqx696TSEwTWvqCT0JunPEHnFyBW8SircMMDrQsb/rjKxZ4rrEV
nz55PeJ9NKXnTwDBlHpblhlQGmpsRv8OiNArNcWjaCPa25i49u8pvRq6lfYtTbF0XaCgTMAF51Xb
fud9UU8Yz6HmuPjeH8g2TE+w75srumHAHqV686I+YsPuKFhzqZq+NQ4V2qhOG34fjMN/KOD1C3zl
+JYMLQuTFl9W7N5hNBrmVR5IZtEP2TqhOlu1UHvKGgpsZiBrDrn4m4m+w9Gwrqwzfls2gp1XCjmf
6BMEYrAmRgn2QFzSy10mrm4fF+i4VqWlDc0ysWlVHcj8mdW2tQL1zjx1tAVHVde5OnMHkl+ewjXT
GitZ8PoGXeERzpLCuvGAbt5UDevQWQuDhl4AgRZU0HAd1RSY45opvdthJbKewA7HN27UjDOUWij0
QnwIOLMPIL1HhGacAoDtHhM8JvIxCOCvjKGqDGgAVj5aJ1shQz5+NmJKcDjpOpVV8fyzraT08u5o
odXgiEvIDywE5ULfaWYBM/GLd7lwvtlWHHCImHReBXlas88MY9tmlWrbYF6aiw5kRhIbINk7rfQY
Ricby0Z8GL+/QwdrhkvJITWUigk/CH3BQVdkCIurApHc2OUsEYtqLLHwLTYaN+ptwwTYqKtEilIw
XCy/g0HuLonUI6/7O5QFy66pnYdn5tw6k5o5AsGK8Ec/ni6nJ4qh0NW18Y9uOjMzfrADK51ypEKF
H6tiGINhbg146AIx7epYB30E7AkL1XRpC1ffTJzXmcP/lWKFjVctbHsvSzAMg6baU4StG84bpaum
d5enDaJ/jYjz1M/lvE/PZ7rKifiD1+2unjOkeTQgcsHKR4jP2rLuwLCzLNcDu89mDTDMWwCNeh7h
yDLnKagviXfQpdUanVRytzDQak2ETCelKb7eWYqNeXPr3cEwOaxRVTFPPuJ1S+iYLOF4Lv9E7Fv9
eZhIEBQiORJdlqAJZDO8jz/5JC+Vmz5pdDGSpGQABch5ga91CUELBEHhO7c0/HKQ5FJMrKQJjO+x
M1jgmzJRrJw92WMxLzRFSMMnSgu2R1Xto+pcM3KUhnbXuRkIXR8VjcaZIw6ktBCkMW/md+TcRexg
78galBWzrFYmQxwBQvRniy+gX+UF2/5acScdJ6na+ZnhV42ghPSyE/u4jsqQ+mfiqCn/eZbpqazq
MM0V6SN5hjCYIcj+HDxq/Ywb7G+PZ2xhSlE0q3eI4Zep1+h1+nN1mgkY/gSWbBVlTpaGtKDETwlR
M8S9RKEASMRrnOH6xLgfhMT5ZmnScSVGscIQaNibSTA8EtKc5FpYyiSFbxYjeAug1SsUOmqYgHwb
3+gHuaO7w/Huom0KzC3XfLyYTXEyN9wqA8+eb3qCKHeIUrUeNOtlfQhLOdO8smfw0749wL2VY/tl
DwzAzLpGocgrx7SyXC0bSN/0r72g3nVfWg8Kj1qex1NVgmIJ76nk+/jkZQObXmHho95TbbthODW4
fJrSwSdY6UQoeweHJVzzIO1BCtDzd+XJq23qAXvqKsSMEkpCjthOn+/N2OwNwMdxjlfhBctmqBC5
DQC9CDU5H/YbExLcmRPBGTV3A1zLtV3DCKctaUCnhMz3m9/78tuEe1QG1w3dciM+nrAM8TMEB5ir
/zFZtIQAs/pYCWmFr3v3Rlbv6F4eb3qMAUzcZMjQe9f/sTnSgCpVoCjjkPbdPei8HpbY+Pg/uyHD
m/tvcDKlHA9JA42Dai62uNI9LBoDCxwhh7vHEEGuYM++9fU9+Wx0eB67x3SmDom+KiSBsDHeVmp2
qssIfdtR2KExSw3Qjpea1yX6dStHUob94CS56wJUpcxm2T3jtdiL/Jz4APB5bzz6PvH60xXyP/eQ
F7/16QQRA+3tZPU3QIOV4VZkJhW62kp8jFCTsPbzeF+7ddbALm/E3iGLS1m625GFKNLJ3V/PjnQt
A5OZDWPLF5aW4JSKHMsjbyx9oErZTi3PId4g91CnWD/0WxkvTa0stm3lfvUeMoaRH43FDJKj2Jia
+OG3M6H16m/DtbInlLyWS4i9eIewnXLKGOBpqkQyHGfTElvnv4Cpk+JJ/RCYV5+PM31/Q+wzzH9P
dptAM/lQnp5C5J0kLGaB038puM6/EirD8/Ujm6qT7U1qRB7vbZFajQrmBJTtAFQEmBflO2FP+K1W
G7mb1QFfymJ/zgVA6mAM2aTjv6vA2eGbBNy0HwJxmT7mA+YpN1fDxmfTip/+voc3sLE+f2L2rgff
lvgihR4UBbNALZIZ1G4xtWU1FJKWP2NgSf4iHMAY4PxBYLPgvUk/geuDuNoJTDvw1PYflK9ZQO8S
tHYt2Oae4OV9O7ZPK1ueQGyFuUaBxMJz42EUk44CKCWr8xdP/p951xTjil3RobofmJxWP7l6gQru
ehxvrlfsPTfAuhjdaWjty9oJlvjHAh0gLlkkmx2qdNuUPfBJPCL041UJofPK4zCYjLI4rK/c0Eeb
YPTN5WWcwCub0OVlCa8Z7cEA8lyijC8mPwyqG1+64sVFYyqtrwxN22A+ZqYDrw3OAgCcD8eZcU/v
S4XelNm0Zr9U3+D+t5OrmsfAmHMA7fZQIjAcOfPiYbn1f2RIRH2YgwRCCVhvqWrPw9L6NzpfzaZB
2p97cD08Z8xjn9ufiT/9mauj5tRBIB2b3mxiwxIRaXEs6K70SgbRFuuhT4Hb7RbPpRHQs55fg+PJ
Jbo5gA4caYzuqAeCGHLHSJZgP8bq6EUrw52GCr12Msh22njPfVo3ejYL9HmsvpVLle8V0v8k+LTU
mcKinLQlterkamPOm12d/DCvIayIj5flLf1E80V8Kt6P1B4x5I3ZjUIxDFZ76M/6xaBYu+Qod0AG
2TFHS+pX03QiveOwcvcq4Bu9FrTXZB82xcSwnlbJGzydFtTRyVa+BGY+oJewULltXZRB0Y7PvP1w
ofOtOfka37elAPl6KrknRG+CxxlEHvSiK1TnsCLEtIb+U5XFoXzxj9NWnPTMCqvZbaiOCL7GFnzQ
wxXK+iZ51gylZb197nEXDLyH3pY7q4CVs4D4ERWZnMAy48IGwTvvY7sMJ5c3OfBVGAoCUWgaSNkR
sSZC5WOeZaGAlRadsjkD5JorTtDk1JAX3chnYpQAcITqa8+sZlBcz0/5U+GnA1SASR0QS8c5C7rv
xQ0IU1iDde5gcqGXWu0hbZDOqMYcqGRNVbefGO+cCs5Uv5o2sRO8898rnu3Q+kassZw5UoMrJ9bb
PGAXExzw+0A1M5B+nGNyFkGQD7GsOx6zkxtflMraOtHFgb+yZZMxrUAxQq/zlDR7HMlLyiCGaXG4
RhCugbk/EJSh5T5rWwGm2Xnw0UC0MmbnLhmvAKJgnTjwsW2oNq/keIUAy7yZwz5dj2p9anSkJhjh
+Qybqbl7/Txo7L8x0vx/fKXWvSDmcrjSaLh2TG6oJ0RIlRT3yvFPZqSV8nzQl3HO8TdxiGtEjnpM
yyFqFfUmKbW6X1wVDyLZV8qQWZLWA09ry2hJQE3siuTusnCt0jDxHwbGlhIz2Ah+4NX3PKZCH1VL
O71VKpi34feA/Z1r57eJy0zO2/ScO4MZ5FogCTXLbhb0ieOvfYt1fuQohB6AU+XRSFIhRyPiGdB1
O0A1vY9uDa/DTOMQka9tB1k2hEBswoTCzwAdbsRAIvgeY54+rfzU3xTZUgn5uH7D4G3yKxAwNASQ
SR7xYM8wXwh1C9qSemjWUqbbdpb9c6YcumbzZzv3AV3Q9qXMSP6ZfAz325dclycO/qHm7jSv8JG8
VbWDI5ezzMxZ9t3fYHlKzBcUWnrU/TzEd+zyE10xIYIkVXwzCH5Jtn4NDoe7X17WV7vvfRPzkXxa
5WQ1chjmcI9ScxnOPT/LZtzr20sEc3hSoYldUwzkqQSi9zsmacXl06B1C5EeERKlCaDdRgZr1mTb
dmn8hPJNFG0B7urAMPnqdDLiQpm5puFxJzh1quxRfkuwRGKzf7iCn+ApyLc5JHWhADHm417u28fY
CkBOzmF7pCyiHuWt5F3WRZcUZiDzd2iAp3CkxAiHSA/CyOJUb4Tncx1joPAcVKzH+nGxCQkr9Qog
S2ldAVLZusG7P1UjTJTIJekweE20kW9u1Jug3JtC8JZtvl3EEGFm2Xi8mt+0xWc2x03Uht8nOCz8
/PsVBC+G23vATBmCfq5A9af+vNipg3IK7Tc1DRJ57IgwBnKdElxJwgKvI6PDYgBdklfZdcakoG9z
hr6nEU9O4tD8MIYa9Xw07Fzs0gPeh0WtVvYZB+ZQkYx75qjin2hxJdXehVeljzKrBu80YzLK5Fhd
PI58Eqp74aL2snwLehooIFkBIAAvRmURlmJ0hSABnDkY8PUxl7AQMSJjqK6AAsIg5uwly3eeLspK
wHoATalSuOeHSF+EQ8rJXL0jQObYlD3sfu6YZnwH3dbiTBFurJpLto4vpjg6+A6w5iAe8kItIBaA
fc5i7ObH0jmBTebdLuXs9AmVPPYKY7sW4Ms9+3mM8wEOziXZ2vgbap/FgShQWFPDKKxEYwo55m4O
guayzds8QcA2l9VWrmct+lpSQllkeQpiG9TnpHPW2oxy5PbfoJHtuKyQb1jJDI/CrjstC/itAMBH
v3VF1uzgx9zd21Wj1cNO3wBopTmyUrzwb8Ge0h/giICX1uHD49hTqqiZVQ0Vy9gecjGeRHuOCmaL
7iYX/VhzwQfcoOdCty2imBQzh8yMidGsAl9k9Js1F7U2ylFhY0MEfFDQhmG0Pj7TR9fUTvAMBXcm
l/Ozl8vCYmkmXvcjj1QXvEQuc9yNRsbTvj9fZzZSjALUrK943/wRu0cyyEBxcoRbRilv1pJJVEsw
v4kPAS0MG9fMqrZIBGhgLGwCNr85DkbU5uyd8cgbL6PsRF0s6dm6rRWHpaUSciggi9dyFjgZcVYP
fzI2APfXsikeP6Ssq8Ftw2HaF65p3WrNSOHtNoqQ1xkfg2LgxU6HmhYyCqPXZuc0/0GIoq24j5Fx
edImlMrLJAHf2A1FPlLfSa3hndHXTRHuWn25+BMo2ghg7peZuc0ANtDW4kdtreyQ7IiBdXMlMoy6
rLlB66ZEdscGvfsu3ccv1VTCvzJOnIoFDD4jinUOIODeMosTUeQeICAKUirGySNhZiobdtaBIfqy
J23dTVa706CxKrP4W71syMSvfFCds6q+00EEtUoJAo8+knGzK/uMXN94OahxkvpjUSM13lOVBAfq
bKtLZclWTLrXhvHL4Nfab8JCLgbt2X5XKQXIq+Zb5fRRgGyHVA12MoveGU7dHsMUqfxsuIa4eQdz
1b4fF2RF2xxjSJqQ7i1S3FAMeIIdmc51SboPvf9ckkzRk9lmcDGU6u0kBwnVB2kLwQXlh82X9oQq
RZRBV2IRgPnaLcxQZKJ6SdUjpKkIHuRPv08rPvXQ9aUDKBsS5G6R1Yed4OiQVOHDmAaI2Rs5xSe1
4nyyBWqxIAlHVQUDLFzNegse6PQ5NCI42J9T//lCVKRVwYeXRUzu2YOB8useiksoBUV5VMrVDKPp
Yd2+j23KHMjDy1ueEq0Mp+/EkFXnHC/hSKQnTvHA+OdV1/OpFN+KgDDD1YH5C+4Al8w6LLhU2Ll6
dKCNqm6cD25K4tUPVRs/QC+3xvdfRZrY/U21WpxeqXNyahVOKDcnmKdBnOa+aleuh/GaeFW4wSIe
v5Y2EzI6LslbO3Yr/uDzpMIz9CePHk7rYoTHNQWeb5uj1gSKERq3H2b4RcdcxbGvZGUbuutpzMq4
uUv7ST5OCyn/aOQotiOO6JRrLzXx0jyfBVPIDslPmgcjxNqc9Fb7KMYnNqgm/sviV2gn/jdT5vEg
g4SBJ1xvpOykwrYWk1YpEUeN27K14/aMMG2lnNJ2FJjStm4mdpDDAi7h3YaQ6ylZ7zCtavi25MjZ
XhxNMhgElxOCMgHb5PWUpeUR3Fo9rrtPCO853h7a6LywAN/ZptZ9hqlu8uYA+FeCa0M2oJJ8isVw
yX5/VRqF2vt/a5v7AJzF/h569sbCEp53OfBEEgiwrSDL0Q0eoBdU5WwyzPpjoZOEPmXfCTXO6TEu
8s5zZJ6ygfGgulJTVHuAsHjR7cw+Rz5c0zaaijQ3D0kHfum+tlXBZ6HexGWSFQW8TbQ4TMi33BRG
2jhe2bALdFxVrgg7PIT4haqPPdJ3pgtX2LNdj0Fl9KMPNi6hKkrRpwtrZ2N3mnM8RIdoeU3z9Adq
1zb1fjR61g8hVHW+3LpzexuPTyPDJf8VujGqozFIpbRmRWuPQTfE7ElerUKQ1tc1fMmepK/fAEfm
yDuPQ1BwayEFdPlLZhbbpJ400vHS5aZct5DiYASm8VWkmRJzaPR+AhrlabPEXQ9+x4zaPRlstmaV
b0N+ax5fhN7eHf2qWBh/HU1m8xhFUIAZTfIosPXd4I3zyrfRwbcG8rtZVD8DTIsDLirpW4FsHedq
CcE77pj7DY6CLLJAAmV+eTMsFWv1ZGC79XhPxJUQxfblHFbHx/RN14mQD70c3PmjHiYYLuOpyxlN
nffPZIuc8AxbqP0iBsnNfs+UU4DCcV/o4R6GSL03KUyRI+ojoYxqP9oJISzNMAjupktH09wla1HQ
8hgem68M2AhAEoKsxePm1X7C+sG0AWA1FyiUR26XSdmO+01dxtcPgIOBLFZd18brlMSsxTVZfPPj
+Yub0Zt3vaI41Gboo7355yrmrBOPRmfOIrRIYHi5vQE1Kgo8zWvkDNsgiNOmTvg5QaMudZoFVk+P
wCe/DABu9CV54jZ4lzKmYcK6d90sRSgf9NkfmniVmYc2sXLbrU20YpnWPYalqx3UDZ4lhxqreI83
MKksRegrewYLGSZmolusmSYOL2vb11NyRUraxr/eE36y30cHTEh3AOnQT2kseZn92ajNowtjyRAS
zrsrnSqtvwN1CiMrRIMUmRvnJYXN8kLZ2874cpxLCv8yTGT2kgTPBK+PRcdoIdRkQBaNjZ7yYoql
SvjH8YSquTGdS8Y1FFLKS0vJedFTxHp2ypGqzio/Dcz8vYwK0QcabJYlRI+28bpG5VmnzODTYjAA
qYynq6ioG7oxeGJkTA431dyHHoORhg3VTbWTd5KTZiMtv5wCpd116owF2pmxQCoi+94PNlbjwflf
G/aHfPTgwd1LHWSbuzwUXkptzLSD6WZ9e2Z/BprIy+uraqghLdzdiSdKz3Y7JRvRYknobbMB+51s
aV64ohAXs3kBajWiz5QrZZphCAWOfj3j7F2VGb8DuajZDCCOpije+ppD/QKjDvgEYc2jl6eoH9tZ
iNiX9hxVMozGtiT/AlvIlT2RrD6bwLueYdBvHxogxdtiTldVhJ3bvGmlVzdoyOzkcPXcm8phRByv
iE67341M3hVnxgn+Pog4uRIh0OQECNi9Xr29yI7sPYSMMaind3HLVTdIoWQiC00bgUvPUjfMFsij
e0yQF9ngLwLNIu9JnH4vXTUlG8mO35cYbt86eEVbmRq5kmv/RocgcAwH04sZMoEYmOsFN/v1J1FN
xnN1bvfTDrJrK2xJEi+72U8HMfUeY8kVyxgJISNhjFpelrecwUiSzm5d3l2defC6B8Mc0Ypu69US
KXh48cFMDVeESJ8Oy6tiJ3RppWZva7vVbaB5ECfrCiRJ0yBJPGNWXGDB6ZWnIA+WWK3oF6prx8aM
f0rInfhMwqVrVXV+ZvOKlSpP0V6OJzo0usNJjrp5MH7CwFs4Fwdry27Uk2NnS1FdwQ0xx7e934RD
AYoWQuu8rONnWZ9R6aaFzN58JR30scdf5zzI2m/NoVXWVwkBq4xa2oFYcutVjYIV1XQXkF/DoYo2
/Kgksm7NcF7S1DKMBJyaRix9hu8tPncZAuxSdHdB5zC15k8isZINlOl+t9+nE/qQhjRHxMAUWt7W
5yLKHpqcPV6qDRKbgmEO2gzNDvaxZQACcZnw8tbUe6dRZoJPQ/4wlDl/ly2XOrIOlxviEKpweVPp
oEVzW5GQ14VZ24do+EBSir1KD85UEP2fDGgUX1xeDl79AZoGpApTJvp6mdktdt3NYyTmtCVlxjur
ByhBs4LrMuWnr2yN6jQppon0/jnzu3ax5oGCT+E5WhoKs0hcHS/peDZNgwTP5XeS7OXb+k/eD16J
OGo9etNzBqRPkUqAzEQMk34f9zHY/kBzGedyCqevV6ayrlOc4r0sGOC9kagAMoCOhxMPTjAJQPKO
cA8IiM/N3TxiuwTH5ugaP/j87fs/jMeOEwHGRm5KOcvlsyQyQ/p8GZH6+zh9VxRAqcJML0LPchga
iUKWB8nCFXiU3cNPhJF6fAfXM2bQ2vLvDI3TxNt3Kl2OMbJiCFOxU98k86T9tzKvmMztKNguDd7T
jA23f1sega/dDox16GWhyNF2KXVqN1O5JW7ZZD02zWIhqhkUBHmovW8qMn6pqpkt9oFLuBYZwLS4
PMjVBPJphV7Dvg8cFHItoeDklf0HmdiufRg0Byj+HDpGTnqIBgS4r6IGhgZIzt3Fm5CWD8b58xQA
dSOStDclCB0mM9jzEry9fixHwuvWHFZDILnQich3Sxe/B1zyM4fOZTFDZk96T0qGPgtpozIHSCBR
hKal6Sk2JeVSG8n5/66meVgThzSl1dzfNn01PJrNUbX0oTVNJcRSn8mlVJLzAAL8o5Xxi2tWzZPH
BbqY1QAh6WSSlAe+Vzbec7+hzija1CjbTv19FmT2Mv0SjQ8c7xokhzmDky+anQaagijlViZXqQwP
L8Ta+VGTbI5wHUbSYiwGfT0K965IzbNEg62khsOYR9wxa1K0dFhSTta10AUDOmv5VPuBjhahh4Af
aWH9HCNYIX3pPjkz9ZPLcoDWtUMceyadTGOndN1KdD1cuLBme9t5nQHGnYMAiQWWUWlprLgRam9h
IzcFcIwR3Xe9OAH9tDEs2aGxfo4DFDHtwD7KqzGUJ5rwH1QxI+2C/Z7pR3g91h5XyxIXbIyc4nXG
m6YdwanJYEDVmL2O3MMMTkSjRtDI2EJIGddfHenNOg1uden9KDxReDjXmAnqJnou+DGJnvSlMAPV
av/Jod/2fdAS4j+b/4bwfc8oG2nF4UHcibPcL3zTIkkzxaEkxcjD9ATFacQbbS9zB0BdXFdTpZiB
Y+tHVgqfdtxt8Po4hEkO9PAkbv/CGIGeYA2hliqN7eEYuoCraqv3mnto/+wZgD80x2AWscATHOF8
iiN2XdscsovSZC2tiszMzBALYUNsp1lrdDRvFintjjJMsuDjdgQdsWSfOBPSTypl3Xh/lacV9izd
qJ0EQIDWlSyz5zySMvu2IsLHgsQuUbeLMqhJ2LBn0My9K2mXSNd37Wx5GnirchpFLGxZMKfFBj4K
C4GBoz1A+JUMthXkZ4S376ypZwzCzHcbOrSpLN7LAZCgWGmK9/zaxzFNgJ6EplKe/E4PZBhgd3Q1
LRfWvpE8A6ADI8QFrIyGCMhKOmJUaRDWeYkcX273nCYOsRGHKgv+9KiG1gdTzSystiMRCkBsa8Ip
64fO/X3GILbNJRrNZudQIXV2RTHPjlSiXsOvlyxk/lyS1E6BwV5DTu7eSNB97oxCblzJ2jEeR8Zx
otA4/MReRFgl5CkKsCtR0m5vP6ZZdOgmyfvn90IL2C8VkElo9V3bbRkU5bIcstMR5Mt0YVPBxkop
diehEooXad1qZblJO6R8mkZqZPTq/+Ly3y0u5ypVXNaOmyJx+6GO1nqT0ylLgOU0EmUnFa4F5GUr
kqqJycfWb48zALwwbVZxUsekpVXWLIbV1GksXRnxs6ZwMvdp3TkEswq7MjQ+o9yHHuObv1L7OI/o
1qz35d8R69jrzOxwekS3fiONHKymz3Yj6hllsbjyzlKB/9ZKiQn7T+zFlIxFAJLlvEiSL7piWYfz
eynxYn24nMFFZ1uPUQfi0C4yd9DYVTMLSa2Du0gLkvmeIEwFkmR32VciY8k5Fn3RVHxe0Vz+F4Xt
/mHmKuSFQW07vHNhMVbvgAfna8D8CgN+K1psqO+B0A/MKZbGbaOjsXjDgUebEssoleE+zMmTxvrB
bbFaGkIMI3kg4u7DEcesjfmmoUGT77tbaia8sbyOGro2O6EBq36Lef0yCI8wHMHLoQqufPDqsI/q
ut+e9SUTGggktjepBMVWONg5gCNbmKeIfll97iXj+yUdKejOQb3rPRwznun8qAvrjIm99pImJgc+
Y19896pYFvKqhfrEBuRwr25m8bvIDqGukus5zM3CHurj9B8pvF+Lhh9/UDbheGrbeDm/2CR7FX3Y
Z+u+0r4ekoWRa2vtjeK43uw+BR5p76tXs8kXl/5XpDWYul5Aq95ufDIVMf42RvRZrMkR5negBBVn
oxvz8us9GV/eTLem+udU9DY0iPZkOleGPNmu5WwP9yqSJWnPQIMf1uIV7bNgTDRKyic5gpuw6Cr/
h9E2YSNYvdPdNsOy+/HQuYejo6alh7wwsfLYkUyZauFiDtFixNoWEz+YLWDdsKFoD9GLT24C8EDb
F2CszkBdrOAqP2CMSnAvk/LJcmhbYtsg8/6TJl1V/yL5ups8n/N4TfMyzkPB3gz7MGwp5eMY8R01
qgjeD9AQnQ5JTRG0M7oBPRdg9kVYaEhL76Ppd4FA/3bwc/m1VKp1f5y6Ijzldcol1dMHFurJ9VYt
2hSVS/G5ZZUCQrzFJ55QYVVtMmeBP064cGDGrCGokV9j9dqets/RuWev6YK6z76gCnFSHMeotR78
aNa5aqV8D/1WgaDY19pnCcbFICoWTM5OThOA/v/l9089I8fQYGSYItjMWTsUD6dp3OTtvb+TJFN8
as+6Xm4YphAl9elEhnGbouPO6uKhwOyiCoNLnGNRocB5ZhIRIW32IAFb3IWVjb2LW5jyGflS3DvB
a4IhuG99aFIwqXQN4iCKzss4wq51CcxLl0gjJ5stZfmXpy73mZY3MNpGAcIzBT+8aZiv4eBz1C1z
gEGbW+lYfMeSRUmbOcC0bo7UEvJOWyxnRS6+SGCxOReRFlshsJ7omjHq8LTF7LX7sN8RE5VC7zvG
xEQYZFQP6dwOZbs9Nfo3K5qc5zzViAgqj+tn+ux2z6m0UPea5ZS8cYby9A/9Nyd2h2yBEjGKCe9u
yJhJATzyoENpVdlL+nPvoFor6y0n6F0t784J6BKJGy9L6q0n26H+aRHUQWzPrrEgDVaMuOp9cz4n
bUdsDNV2gJh0vsggwrtfWHVsjgFdL233mE07JJqG8NXqzQxxBnPMIjlhlZTqno+LoHJUvWBkZOnW
dh8y3TIDjlWZD6AxGtthN/P6cOzBKfFTQof3W8dprw7CNeCpYWlx4ZA4oamVLzROs7cAWQ0vh4JY
ew8vyLkpvTc1995IkomAc+h9NwOJktZCfVr+SG14VLfjKwzxVENWjTVyaGwpfq6MeGrqEM/5tAxc
/pJFYeTJmQfHaqL2ecSMO9HfiTF9d4p7+yK1jRXbXpmijxQaA1tCeWKnaxMSsSBFMX34cc7Swv5t
Q/uFC0bVM3JUEcV2T1ySIzBT4We0qEyLAOcfd0vf1Ly+nzwnGWHd6l+wG4TGOS7P3AgbNIkQeroe
yRmLKKzFF9pPzOSYCIqZXRRf89zmSuUyVnr82kShMK1C8B9n3A8I/5KAoDJuGc7uM4U88ufoP6vs
uANnSvYp3XjyTp0VCuujybT2Mj4Az9L5kqhEIesRC+zYVqU9QKfsIHGB6wiKhD9sSn6GRDeDgWoL
H+t1dJzh+jqozEnFupPlTXf70vv7pD+WGDHXDbDSFT6Px70WQ4KrPiOFN8Wowg0bzN8Kj1/2UAi3
HXuYutR9sPhxYum5ta/NHHdy11yPXJLWSqf7b+iff6e5ZixLqTy4iS8yZfZt4gXxcoXeBVMknowJ
SIuNvkfns/grHg1DIib5oLyC3q02VT6MSEksE37FbrWuzcjqQdpt81EOzRl5nvTskPduv5T0wblv
4UmqRTG3NqzmT+J9+C6ca1FJZeTfhMqjxzo6hEOSM8wzv6OL+gTZ07WyJ6DmlOFD1ouOj89pTIiH
ynhl95fuYP4XB4CNrboeiN4RotiTNIhPkFpa56g/CUwEoZt806CpPdgc34ZgtvKT3cwAnYod15tN
T0EMw7R8+v7RhTl8QyoviosFXRHmXGkJE/gpRxk2di2U+tORbjCiH4nQB2ysHJgEkNTxmf59QpMW
akl+w/sZ+IQYkV0lI8UV4Tyc5o9+SymOSip5KZtRIiBB2oehYyasyIlIiT9o/Rn1SDT1koj7u0le
CxRkpkOGVNPQ/q9RfI/+ZIrYOi8f3ZroZrptAabqMQK8Mg2mEWGSU0Yj5s+F7aq9RwTH9HeCRbBB
Rxs67I9RkXlj/eiXYzN10Lb8Jrk3AlL3Hjn4igJxREt5E9yzZTCt3un8kKwIrCOTlbo9nU+imL2j
N3m7i+0gaWSrzfeZRSR8l73mFCNKgviYCxgrfnf5NE8eGha/76gkUMKohjEb2X9HlnrPT8eerxah
pU61Z3bz0LYjjmvvaMg2THEq+q6oJFwG+rWm2/lOfXQuBrJ2mN3j6i5NFfNXYL6ByhmFTTcydMIb
QJ0gTYuJOz8ZWExSisQ4XHgUcT5EqntEBKsobsb4gCs65tZEHbHqw6n/WPUShtx979EsRs53Gmsi
ZHTt++Vj6Ib+n530dTYd/I9v3Kvo7wte0zR8oknF9+C5SEVJcPWxnmPAtsA0Y/qc/MXCnHEIktfm
QemrRoILQhfjJyaDspkxyQya90BdH6aS1s0uyo6R+NLJy+ib7flyai09iAv4Dr+weNvbF5AQ5Mqp
cV2aJKhuQcT6yMvHevCPlLkJqI8URn0Naoy6KbcPBotCUtBr6QEPub5WL8GOevLLV0GbP87xyOFM
kkkPUfMZLBGBwr+NtJsjOyBR9HKhA1U9PrBhAaSdQkLh6SuOoVkJrBQrN3ZgmmYviITIslQ70X5n
Lpi2iXwKdjUjAycFpR4uAIywRi/z2cwuop94tFdJMSjW7d3y7++0ToVqgbiCjgJaKZ5P7V/A/bBN
eOqFdmt4xsVxsDHkmTWRfezi4Pqa7yefZ0sizcGmaLT8h9iDfqwubEb+n1YY15VX894aWXn4rXYe
McSugWFcLVbdMyQ/NbEfateSDJl7UVQWX6YVSqB69z839p7/oPNpbMcg1rFOR1yzNvLBnFJXP3qe
y955oUgccVFl86mTbJARPhyVzVhPLMuqEILriB2Tc36JkOAViOwh9mCWUOs3o8dCtZQtxgNI+cSO
Zr9ID+PrD4HIPKRBAc9ch/rR+WQ8gZVgimamKyGlNkRqBMzsmqza4q8vr2VA539C6FjvbLo6DUHT
k4YHJrR0y8qkQ4oVfe60eItdNb0PhmKy33tLv854egCwvyU45McEWo/uIyeUDOvs6anIjjfUc2br
+oSIbjm6LWOR6s3jMP2FpAj0l8NGALNwu/V/SSA/Z3SBnrielR6spmac4zNOofsQMrX+4mkEIOJc
2rHxIv+Zv+Q78Cb9yI84r83TTiWynD8jW/Gld61CCg1pBv0TK0S+bWjxo3/q3z/A6NTskyGIERsi
nlShwcQCrDq7x88iFVMGRt6CATW61OR/jYCvugq/FdWgTpOcMO7Cwd24Wrl53P0L6MBqKfij9NnG
3hFkgKbQf2a4T0tITgq22E8oQCx50rpmFEgrk4gu+jYFHUcL9JxJb60EYo1yHnIh2scM+pkJbjsq
BkKqxtuITYQc3NQNN6/e/1WgE9lU2gelhM3ntNsz+rs2kXT34uJTYbK1enjNmOjgUsrp/vBxk+Zp
iws81jd/dIFxouLIUU2wUO7H1jgoTEr8NWL5tJob2a5XF+0leDed7pqoVL359ah8pd6aSP2+vavh
lnmKssKL2MGMB4dzQ7IL3YQGNG2Tdhlkek9b8ckvNG1NqCzMnFaIDsxLIC1yQom4LckSGyHZgxS8
VuKDWCXDOyYDyERqQUoMXP2uhGjARvMEcJPrANmoSprWpyTvBD+vkkDiUOEriPobsXwWRSMxSea5
p4v3XOQ2SCLlkWE/dTuyxtw21iohB8/T0uICfpW42K2Ld4thbZR8sUNPDW/d9GkS6t/4z8nUCYCi
19GMES5jHIDLCEkNdzs0vDJAhMDJyoy7B0GIrqqxSrIuaSS1GH/8KX3RYOqehr7iCNy0Th4mPrE5
1cJWN8cBhd4OD11OAy6i0AiqibuxKttD6jXg0tvrPZGhBsIGr5vE4NHuaHyqHjY/WP26vg8cGJm1
vD555NJCY2X04dstvUx8HBMGKKdYouDTgc/XfnAPmMOzL+q8RCRzV9czL3uaU5qvhpbumGTmz3FO
SeA+wMM9+PBiumcPrLEfAAXkyAXsE6gFOe7xFmoVBcuYX8GNjuNT+iY3TOcGh9GTXD7UYvXd1mrQ
vGNiQ4H+6+bJyg8puBB7DnVOjKcIwOvH7WAsCLHv1od1vGM8sYDNK/AoeDtl8VPXANMJwjPGmVF+
WYbTTlf7GIf1OcKiyY9IgIe0QDhSbbF27rpxSoFvG9hGtWdwGiZBDDIXikDLeKi0hcjPUNAKEqZs
UJ8SAjrg0ygyK85s3R+uvrnfr5FJxQmG/flnaR5olqCDUByVOwWTjF5zpgr0Bq92TixkZXdqJk6P
I89p17X89BbblPwL48tfAktdw+WcUfAtbdwym5TgqeOVwrkUXVFqCvXMpjRdjIsF4bQYH16lgl8r
NB42yT5fH0MjN1oaAYYqI+9jH2n6jKyuZ3stpDKeClu8/hNbzBVyHH7BFzyfXgospgfUW75TC1Yr
WvRi/0MdAo7fruJ/xtvMX1rIg9NFXskRes9/e8dRIjCCUtuNWJ36T12og0KIlOYgPMrRqvjDArM9
6HNNKljw3qYo4nuplp55nFkrNSAtTSIkvZuyGMpWy/WY+oQZFHBbuh8vfxIMOCbZhCYhYtqOJPXJ
JF+KyqfiYWH6QGB0I4qcbNnZJdLKidlRQWb4d7IVcoV5PzUxHNlmvbJCGzLbslBVo9pHHgNCq26Y
We/dLKUpD4a0OrbFueIRMcOqwFeGy4OCZiUDzs23jz+Aj/BjCixXjVVaMPGVSZffEbTDv5SdyY5Y
cKzrXNasWe+B/fACa7covuJFh+qPJCksNM1XHrMxTIh68AYw0aZUIK9n3vmbYo1LWN4y6rZt2HBg
NZYXB2vjdUnWJG6iXkamNpxDUKel/gxjWJtqxnmDGyZmj4Cr5bnqzP7BR3YdzslRA9kfJMJ+NCn3
RezAHrn2TyxRdGaGPPPi5MjpJknAb6BNm2qSRqKfONYu48JeBrOssf3jPC2gIyM3p65UGGKh6ETN
+A0LwovRdTWAGXnTOUtZ/6SCcJEl/E8iVU17uclhyUkYSLl7ghM4ANJV22hiE2NW1UH7whDKvszF
aBpAILbbwEytZAjZcT3LE0byikFFn690PwwNM4k+dfifJgTBeTkYQ/5ZhniKj9EuP8g6SuLvcLNY
6LjzYpl/HlJZ16aLRat4QwEu5R9Uk8yFaCRMyf43qexyyfspAeqwRhVQeVfOQlIPwePtMiHnZINf
ZnKVGBledn8BfQ1Dyx0tdRPc20WnCJtNfXVVmswKVevtYpm/QomS4qHyDItdxayh6Wm+EAldXJ3n
4k4jhbUbuXkvbSI4nLt1e6d+lGuU2QsUMtjtyEQJHZaZgQg0cUvHhpbbjO841glF0GcwiVBGlQj/
YWNbD90GabpOqfWqC5YBCufguyHHq/DdoXZC5EVHbUFUEbISESXK2vj8cFp45XMfzTbQg8am00oA
MsJUDWPdelnWAQxRnBFWB/Gqc7usfUSmz9S8A5igV9hkdYodIibrqPl2Ee0kHdiU8bBTZmtuHouA
G1AnBm+L6UAs4t6yL/my88AJGGqMN+wm9prC4AuHTRWD1d/HuJsXWhrdPdyylU5TiY8VjThTXDj1
88yJkbxxfml7BXiHIMBWLmI08yhSQceV/iQYU1MJjSFI6j5FvIpRH2AoYm/ok8YL9sLTt6QJ34ZL
X5xLcfKRSEQ5CTPRGlI/MBv0HFt8WI74EqrkO+OSnEzB5UMBB84gvG4wG8CQo6kNfUaa6RES73HX
ygYFIbcaZ/spLk0SMpk97Ks/x2QnGehbWa7/sMdm4iybrDndYL9TDsJoyIgAnbkSdXG+V4wLoNwq
qR4GKk3tTRfv2DjnwpCNtvFNqQgEnfQC3PaDGw5LX+kF70Xsho3iwkwGHO9xAzx5UsM0/zP8Taxp
EGV8vixMIQVdXIA5GIfMDQPiDNe1obznM5atHsyRz1J3vQClhECuwzWNDG/ZGPqB4hFH7T13RdQx
FcrU1zarps9oK9GHJ+IuBG4kNSHwmMNTGH6KhiPeib5buwMOk8Iz/ERAukSm/TrdRRQ/lKDNZvtr
qQlctj0NcQLFpHpfQmVhyKQKl4tXiL8uvnld/l2sgK/oEZzTa0KhsiScVtCcV1ROQcMIgflrBOLT
ms0w1ZL5EqCKUEyroYR5PNof9iFWcGg8AABN6NzKQOaXHbPXt8cp2iV8tQAR3/KmYrcWxYkpPdhB
fDXhi4racAqIaQNCgH1vKXWIV0YROXrpM+38p2uJr7zfyPQjhhUbF1GGWqlSoIrUM/zNG03ZZXSc
LyYa5YVkAF3HMFht999S9Q9kU0+3QKwPVeIQ/01vRy4JALYvKoWMWttjyX0uKxW+fcMGSk5Gr/+i
AIizz9laWLPjFCF8PVxFEPTqPiGkyeDwmf0Zod3Y2eqHdxK1vPkqIQK8j5H1PN05l9nPyRNmp/71
311P84hHR9qVFPDiG3TSRPyUjprj37Z01MVZNA7WOezNqKdnHeff1DHWwqbLuam9PtK6RbjfwKTx
+kTJk+IVMPLnI8/o7VfT9/ui/wIOx9CUL7lRM6XsC3/Ta2efFHpSn3Fk5HIr+LOneH395SSN/WCN
F1CHemk9ZMf+vjZFpASXK/HzHcyp6ftrQWFpPs+ZGuHANQnxHEnxYZQPEiCZkcdI/QT5jM7sipp4
4sjwQ6vZfL36a1tGaOWh4oYJPt96d/coTgj2Kf0cGDDVYB7cQKZphxYvYyha0YLnpM137Vqt6EJj
ak3go7S5APdcVRae3hJpnaYX2m4UdtxGa7ESqh8ctiEPi4RqyO+xbngSDOPfKDCQtPCnW6ZlD8ks
Ztuw/LAFv5iTZF1WfLaxNhCmDyhaaZ2sjdq2VP8x7jL5q4aVLwWozpOXdKdp86O1XIgpj8MvUF1L
zwFW0jcgN18RH8hHBRqzdFiSE4Be6HAF9nHjD79FIdSKSQm55VToMlVU5j9xZVmNikTVo2Qv1zcr
mUuPpGZ6vA6nxgqzLVbV8z0kRL9aSUg9m1mQDtKoV7gtUTq7xox/8hp//HXISVMsP6zTs21808/Z
CV6l2OdlfZJYn7UczzRCBdNHhbCJGUf1n6BHhZk8uLP46Ad+teq6VRwmBM25F/fgB0rPkbrXL3vt
fJWsYIAZ7QBZdplZht1UJu/aHH9rUcZYdcvzlzGPgfWYMq40CSNcWdqFzV+mA47cs/84LD0DSWkX
E84LrXLblw0xDu7v3pwx/V/Q/HvwgpdqxsOZ6hiUiCoQb1KPwUOugen9rED+D6GcTA+hQGq0/a0G
ExjUoWZqURxK6cdqC1p539gkQea2FfwQMkpEd/+P9Fj3z2um4wgnPNnmRYceBS/FFLIT7s4lNrV3
7IqZLBwceshNpCVeitZodr44T03vT0u1AuCzw8AjDD4QSva3TPz3reNWm62lBDrVKG9TxQTfrjds
z2SPefyV3tYNCeX9mJZzyNDqU7+x0WLLeCDtBOhJ7+Yf2eW19sbyt02RJ+pMk9Du9rUuUKJbQdj2
jED6tYlLJ7AWhY2fs7uHgVVwbTg3hcLPEdCe3WQyCZEiRZmwZG1iS7jLmwDUQoQp67E/EPreENc1
9lh5oWOZhelnUCEgdRkqEHpl0Ycs39rUnPN72Rrx0qLbSNtHESzc/eUh0xXcFkp5izAfq+jmm4+a
C3Rq40si9CoOEB4vKMaPhdXTu6ltFW1Iv51+hcAoQvowpPQxe7UhDCVz3fmHp7hZ/ssUdcJzmtrx
8O8YGVqyH4ZVFtWOxOlX0PlAoPqC6npLzjokN12Ha+L0HXgiQOxUOwTd0NZa5i06qjHU1pUrmAAB
HzD8IeHbIJVLvBziOHrqITtcdAA/xCCDcBUkFP6uya6QTP8Mg+sp3fYd0yBeFrCglbFZ8G26bRRk
W9rbpbJXLvBLyQLLb0O+GDq3pgZiqjo/CKruPFJT5Z/TiuhyxlIrC8xz27jJMi6F6PWcBAx6oHVc
PjFYciLwNytsjwRclVJaVKSBj3HZyziwTzvXcZLz4oEGSSr+0gF29/88rMj+77vV2c8UmpmcuJwD
ced0EsizMDTRzev7nQ6s4EPN9uyEo/pdr+QdLnLVpYfnN+8yTAzfq8wdyihaxh0zGOc7sU5TA3K1
wNNPQjZnhUak93p0QFW57GkcbcisL9Ruc2pvXhjda9Nfm7BXnlLDNLzHozXtHuepSFCnIg6/seZF
RXuxm0QiWIR20eAKLecneGFlLTS0+o7ptc09xALlinXLBbkPQawZkVR9uZepQZj9avEOLr898fAh
z6BhqfC76F7HF9c5Sf6rfINUI7H8N6fhiQX8vNOP+iTwefUAF/JyJPS5HOQu4HX9Jf3mkaWcGBUt
7m7JZhWyWDORl8/YF6Q3yTFpnk3qvxJefpujG4AQP6UTW7SyNCIvV6uBTZQzJEcoFN8W84SDGKgL
nKCU008SkbTTuEtd4EzYr7nqhrUAySVUewx+EO3iMEwjBweaHv9C9ZtQ8+CYshBTN1A31KIGaf4d
ZwajV7xdVCiVrKgGH4Ez4ZxE1lC99NRKC4gN/PZWDKXxHDrqQZpJspSTJTX/KBrQRCjHUMfUehwB
XcuM/Qk+VJuI3GSjJ63HgoMBaHdXeLm4Wfd8a0NxhIUz/eUqnQ0+jDgy5Jey/rKH+TZhEVZgIqwy
som2/YTkh36qiLNcBADzBfwPG1c7OP9M8nqRClQHVMORp+GpU8bH7j8WHzsooD2WkXW8b5jP3gJK
rEtJ3iPyvlDMWtPrMomOi22Kl09e47sWWRIM7TxIP5MJj7L+FujZ+fp929133jLlcpvsvB9b9nPX
hx0qsa5ysJTpZtinm2M9hvQlHD79Jk7cmlW2mMYsImH3R3XDXWNBK9HyR12tBgooLSsXMguWSU6w
3OOq4UNRKUeMqofGYSKRNpcPXxyfKBvxHpTeejcSiy524pUMdwxjDutY0tUGL7X/gN7VSCAYWPWu
+vvMknPqj+L3PiPX1Nt8p/CywTUCVrDjlFpGcKTqhwXB2MyskRMkirBOXWIEFFMVxkU8uiwQWltD
19daeM04xEuK3/rDY4VXyaM3JqcZ42RdQE06bgIeyHOyrShbDI4+APH87C8oKynWffvKsBBmi3S0
vq2EeO/v0h5y4hTfrONVj7kLCiv59z19MstcxLBYjT6za5fGP+D5GR0S7wtpMb1QVmh7PtKo7iJy
hnHrAma3VzkuHaMrkxEUv+iXgeBs8P2YprVkBq1dYErDvrA/Dz+eqpDqV1RXXERBb28cbcfr/rZj
K7N9MOvYCajqSk7wIT8KY0XSw/B7l8TaON7PO8h8LOFvH4O3P9qFZOljqjf23CIF5oM6GQ0vPHSn
+M8bNVTR7z2W6hcswgahFHSegUWf1HFt4Ara1lBuDnyO46pBsPV9qRM6kYZC+36OGQj+6xnbpWzh
If6JQNNDLk07LqlsKecKP4riX1i7X+5+Iigdj5/CtVC/v2i4qeWtybAZl5YCaobF5n3rSjSwGssE
X50sS7Gy1Pf5ePb7IHcLmSZHGHgO1RHF0YA9DIs3+pIITAl+AhhTh2NqOFOdVDfg+wET9AlmoI7G
BcmfxjbtG2U50FTebTXv2kNUvust59NGGzCzEg/L3x1IwIc88aa45/ydmX1NIpU9ihpqXRSxm5/p
dqzWEOVhSRvj5cvDHam4Ov5RxzvCdU2OLU5YBzHLs6ctqpmQngaZHboNydsUMXj5WGusI2AsDrc+
jtEhWll8MNwyLPVU0j4mjbyTxl7qXGcp0Xokd20x1gsXqW8LYTxrM3c046bHvUi5UChZKV6rkFxb
G3Se5ifY/5A7BQKS8IX2GkJVTtrwam0vUPsZXUY2zx4W9fbGa4/Q/ejle598Xhrrh+kFRSdEtoLd
3C2hAvX79oBNJ9oIcnoHhohpN4VTAtP26w8vyv6OkjSgMjCBbN4eahC+LZ5o3J9L5956v3t7AJDH
slKSE0DIHW4/S+B1xVJw+K/dCqxQfA7Ov22deuDFxNOJ5wsYJQ36kB6vaDp01xya2+pUM2aLOOdD
WiRQBokdihwntrGbmbXBCSuVpgz+98ofrO0T+yTG7aFACfQxv7bE+naMQqfr2Whw7DQUs71nrdE9
bQsiHyvn07PeV7zyTzin+vxMIJePFfrXTJu5aRbkpzu+m2WnKycWLH3kG1mbLq2zj7zIj4+Wgb4p
jpC3QW3v1+vg7Bt1a9SvZ88n/gF7LFKnOW4QN1zx14lrG4RjFImawfWL5eCrszjyUOvQfQL7n631
m2dG5Vf5tG52KoZ0i+zYY5kvkUMSqzk8FQpkKCIFc9g/nAyqwDqQJGv3Rrg3FWK5rnIHOVD0LmsK
r88L8qfj3wO05Eq+c7keDmfx6epzdd+IdQcdvMoyDF8S9+u0/IbMvn4x9qXArJFXwTOzZxpb6cX+
cIvBoZab+45iMxZ+2EP5g+B9ph8RrKqrr+jLl8N2ZA3PT3iw3MEP2qh7GRZiiTFu2S4ukd02g47k
jvsJgW+C/je8ajIlI+z9gz+1itcrTl0iNFgp8cG9b1t4LgJOJjVFnh/OREOZKDPgirNayKbnpo7q
fVggWnk4r4orz4LNFGekH7GJD6qtAFDjiNOAc0EolPmbyoEkWaFnik2lZa8YDANXUmOEXrleO0+e
QAFM/0VspIe2q5Q4TPPEEZEYspFw5i9WyYvRpiWO9JYyjphvQZG2WVA5+1q59/uMdKgS36UeW5bQ
w4ohnwXGwszZahBFC8W9MIhVopLo77y45T7oYyJ/vD+0yvDzaSwgu494MkCOpvEYUhzZmGD2dPX6
q+Ve5mmlvEAK+Ki55MS+0XLrnJj8K8yVmN1aLh28Hfl7lSCut54tG4/yc2LXckORRYNMqQz28HBp
2f6IsOBAUS+x9FW+4oRDEJsLGytb8GSu0jE4qTr42zGyBwgeRTtdNYthbdTxoGb8cxNpBwC7rhyE
F8gZr7YcpJW9zv+tTUEe8+KVyuH6WYZgLN206rPlSM1WhjdcKCjA3RtdIl456QAaIeoVvn4xgIf2
/DPqR7hX2NaCM6aYaH/7AYTpst4CIl43hzmvRL2IsgiRZEDa37Qe8asbUxYoKmRy/AVkiFSFETrP
mzveJotyebYB64LFh7vOk0iYiK/00hBF4IZCEAxxsQaJnKRfvswZ70Cv98wNXDmKCdtIvSvZcbqa
LP/Wv5j4USmAX9ASan7P+/aBbt70WYTF/vVL1iO7jvAy6dduwfpXnVHNIir5ZQ+qrWiwIeuPqDpy
ETu8XJnHXq23wx6taBzVG/87JwHV0iwnPZFV9ErNp8/3RFSDcqZ/OGgJQEFnG1LhlcdD9+ObbeVA
1GoW7VvcUKBPbv58yYl0FhZaKwmd64b80neayFYUUJgjXcsckRxCWLAkfSzgLPGkMwtRgSWOYUcD
tXnfn2/Nm5vCcCszydIpo4iD0/9GSDxcp7E+pRDSQ02yvZkAJNx20YQ4JWxV+niTd2tpn2dkAvuu
eTxBqPFpD2VMg8UhMuazJSZYeSreXPJn6Eg2jHVmQgPh344cdx9ht64dF5+kMUREuOABEUzASkfg
TEyo0vAkPQzRSyibmcfN2r69xgPPNKkm7HhxDjogrDlvZf6IVpsig268pT3UO0kU5SRcad/LnJtx
jLf7m3NZTH87fO6nNZ49jiRAJu1MLTqmRfJKAq2MgTbHeGPI4vf3a3LbQGEiBjGHFgc7XszMaHGZ
jCyLInlL9wBwJqAd22nzQH8+mAfw/dU5SwkNihQKOjRORx57//xuma9Pcr8n59alR5se3R41xrwC
9Ix3Df7l42ges8XvfJW7yJONFSgvCSGWdaI5/OdWOkejPX6Lg1ErpiFmb2MhqtfI3q6BYTyHV50H
naQ6iq7lur7w2FaYveXeFrMidsdXdE0SI5ccZvINMynKbO5TkYVoXN3hAU/k7S/fLPzLj5ZNya1M
QCVm+FXqNNpRp+ZMghTWboAD0AyJXK15PU0j2G2pAZIQWwSK/8wseYBPhg8zVlKcIRvuQESQP12L
T9e06QsW866X2Sqi2vBfLxAQv8mO8kXnWomr8M666yBorUeyx2GKXfMiDYsX2FqFfUL1q+ebbIuo
hxhJlQB1hD+JPG1xIay6igPU23069QPrgkD0aw6Zj/Ev+kVVjk31FbHVmov3OPAeB4rkGUlNRB8l
qyPKaoubhDqizNShX76ilCT2+aqnXIwNiNq1ufJKsihGi4Zb/Kb8hlgFrmGfQ3xEGnvnkyzqv+z2
TjfzZr2iQYSC5gcjW4WH1dx4umxajQIBv5MNXLnZRJN23hvIACimHmptmZ6DIAZhjjlsEMqrlejB
VasQfY9UKfcYritK/3UTcHR98XiaaVirXX2fHVKwsZuAL4mwU2J0JAL5nozZOY6rqT1RdP4EInG1
+n6bb+ZDIwzo7vXnIasqhCDSvBylqEpPad2q6LK5ZSHbmMn+NCa/SLuytnj2fw7XS8luN2HQ5DE7
kwJI99TkU0R7B5IxjjOdA/t+QGd4vxNnqS5DxyzilHzAB4qpyuOgEUav+XGsFIBUeqbkOHHKg+oh
8ZbGzeHGUD0vDsZuHCGDthvW4m51kuDBssAF5HsLUZfBtBDduBTewhCal0f9pkjQnKUrKShc/wzg
D4LLuYzEO3J4RJZHMwSRr3n3PVKEmVpzsYmSqWkRxSPh7259KCLudQGkOMwU+Hwsr22D/tDcAtwH
guT63eqffHkCej1DCtjX8zOM13IfiBWzwQnvgzv7p30CySsaJvb/bZafKbOYB857K59d6Fu8hNSY
Sqy0dVCxzxk5WwcpqHNTIah9tVE1w4pkRY2z/UQsNVQ8dqu5QpbgheA0YaOFqekVkpJzVkWWUxHP
Qb1e3qdninlawnIpB9njiF7QUuCW3Rqmt+5RShxbxC10IJuzEz9LFK6PbaMCNyTJs5vlmwF7uDfw
C9CZ+W8Oy05sbjF4i0AvwvztCV1ffLq+Kcirl1hBafQpJEDSHcpeJ21JdO3rdwIoEd73dqAOcHDm
Cr9hyUWZcP+1W7fckBxF9TaC3c7/KkaIt0m7rsVZrrCZ8Ndf73slIWhqHp9blBIuHD8syuMTF3Wm
eeu6klT6RZ/U22sghm84aI1fFoVMLm7ei1pdMmUL4mZbky4eryv7pRnoBlXC6rj8YC95LVb7v2c8
gV2SifWE41xDRmcu7UKBXtsz/Cngk0I65FMzcZjJmQL3Ls7+ckl9gdwY9QvdoCu9Lxslch/q8lxa
4H+qXqVV5nQgyUNQBs/zRA2/SMA7XHy6yCUrrvf7S894jcm7llmnJh1WUFjpTcGqLMEnK4tzqO82
NOHGdmQmKnwlEjs+0qE630wQ9JgG9FMoUJdQYr4WovggkCXMhr5L+LolbrwF8n9Q2pB719KJP/HL
3GubRGLvLiJ6c6eyRherzTPX861H+ZwqTGJwzZPUe9xp2CnsnbaLjrUy/M/5B7n1Dx5yHhFXUp5V
N2G7KXBNdrWLrXV6f00ZvVN8U8VGy7bcuMyhQ48UGC6IECg0igaUQpdWa672OCWmcVj6UEjGKIYP
DrrponfaSXEAX0fp7T5O6CRs5fp8lSDpyVokVAc0PlzYyxE3HpQ8qr7jrwZajmN6mdreNL4S8KW2
oT9nY3i2zXahp7Ic4be4KYBCWNiMEgIn5A5GeJNu9E+4tKy0QpajiG3mEZNSFZghfkU3gP3rCsFm
lIwCnroIPD9bwsWh5tjhW//94ht1GrMRkhtGDLEj73tem8hRTCPBO+UIkKuHWZ2mSq1Fv3zMe8nv
4Ol++i2p5+D/7OkOsP66goQiQINpWvlXdyE2HHQmnVU96Z44uq6BID6DkocgblklyqG+FTTL+376
T87wTslBX4pKEWBmrxIPOeWbMz8269A0T0g698JuymyROS/CIGlNguPDo3HB5Fgbrq4CfKcbFwdk
G2vKNthz1Re7zG+KsQWz+BDO+MxbwdK619n/5IBbasYOZI9H5XVqGs4oMeYncgu+toydROCeL6YG
JH7SZdNiLmBzfw3yjE0Hoy+SEQ1ZqM+/ULx1YFs87z280ZuocYK3rx8v3wURmVuyjzfy+ZKMKZdF
cijf5+cjIUJKwZwOc5DDDokh8AZeKsNQMCQERy9G9a99kFYUPlZp/X2gGokeUD6Qac8VUA/HJ+TE
W236gjP2VDcQ/D++2UN6+CjO3sYeVXONzT3exDf3/rZzbPt8m9OZE+dt1kBQtLCuNiKw+7bPhPnl
bntQTEvNKVaqYcZFJk+acfb9d4vKkMT5GqKAwJXEh2HvLoTD9oPRwL4Qb8dj8HyffEdldxlfOVMm
HKqvp1dh4ZUJsmMGH6tB6ETSuDo6w17Irvn6WfRcCw0D1ocxAsD3udesSO7WOLSQcoV0exR+djDX
T/6ef1dCOWGYIHX02xMHffM4aEKHGv5GqKm8jFPetEXs+eKMs3MjEjpy4W0nJ2m9Mjr9rc3coAo5
e+BweyoKzLkCBocBRbUH1RKpNCT6OzWOpkevHIjtOVsAmZoOaRV8IheTCLInJpKbsu2/kJRKbwHb
fntgqiJONnzIUl5VAIbZoCecBM7qRZS1UIXLGFJfIe21UW3bdDk2orirTAJRZXuVYEm8/lAZ3Rrj
NlF3RFiZQGv86ly+Crw0EAm25Rny9ZlOkxuWfEMypQuQNrd92SVyywfdAUn3Zg7amndhMirAoNz6
Jp7M9ScY8rqyPGCx8JSB8VOTx58dHdkl24P5K3hImWD961gh/lWKrnfnpXhhIqJ78hhtjyXVEukt
39BNch2riAqwd9pxPxOc6D5iQNWZodKVT/xNTco/nkVJmB0GRE/twX/7yXafnGGwZBulYUeeULO0
aYP4cZsqwqlayNe0OQ/bJNzS+p1JO4NS52iXGZ7oGZn2njvVZG9YbHyyX27qgNTUNfuQtvdQegI9
NRLMeu+MZmqN/F/gloaVQbRewbPivU+/JAfwsNFoIhShalMP7NVWeMK32+R4G5XtSy1ddgArTGZd
/8OlMnjVCt0uL8P3ZBxxm9fuXsPjaPQozLCXEbQq1zz0cBcREqmZ6T0E0bVDjs8oCgjST+4of5Ij
Z0moWg1Q5cTcYCfGOrLhcuhiNaZmE/u/NDWPRpLuVl6ZXdB6Mtnak7iICwVYpznml2G7Y4jDJRE1
UAygflYYJP5LGp1pCZOLbseMx/sPhFZRmOiBwAf1OpzAQ0jWOT1jZV8CH0J8N7Fm2IKs1LABE7mX
TcddOa82q+S9QaHGEnS7v4AnfY118AwbrBF8Wd4ndDrl4PXQRk5pHdz3kbnCAzcsA91TQUYHscOe
kZKFLvPggDbapn6A3lnEpbSgsZAWba3T5KAWqtsiTg2WtzRsu0Nt/g/AglSWsgadWQn/a2DdlMup
HEPfpbNkIiSdJJO9sJC1Vhj3cHHM/q8yOeFKg0ngg6vUFO9RQhADKIbJBqKLAmnyDDatDn0Ynn0Q
5jCytUxx9cRUX03Hn8ZJSyo7BhjcmkJMfkYbLMWvXS1EZAP3Nc/U6rSRWItZarTlxvn8ML3DG+3/
l65aEMLjSOF6C/lId/CuFWXQ8VukrViZCZXTouCrHhv7qrfX/6DABhpRTVeKYAOQjpAyxHFKM9ws
cmz+FQc1VNuMv7N9bvcBrbraWzKi3AQJEgDs7vUH7IAME8W5Q2HP99voPfktVNlOhBgdTLj8KNBc
6bG9foRCGsZDOC/3xMoU6y/etFNkxhSYR18RBileZddjrZPpHN/vZWvIAQLee2mF8lLnGQl5Z/fk
RTPPit5Cstm2qmLOhAUMoSxvHN+FeN3OviHig0S16rT61FMYZaZ49ULWJkh4jKfVsfFgzwjMzou4
v42AldDD76PUKupjA9hQMOQ+LLWk5u+/4WCV9f2B/LlM35jmbHHu2RpXH4Iw4uZdudL0DE71YLc0
wUiTSzg5cA//SMHoSxDL7bbcAsbBURi9eu+ws72TrrsGJ3Mp6t+3jcEdiBPwtk2se2RD7G0IOHvz
1mil8xFHfVQVNFFBxYorShk/g1g1Ee71kEIqyIs4Ebb6+JvyglxP+vRDStolvcFv2S9O2XXbQTT4
kVDBHAyJzzIRHItwdzbx9ITdA0f93gcYlRW8r2uoD5EgYvyr71dRFZ68rem+f+6eLT1bi9VZ0/3m
lI+IaN/gDK7iV/T8FbrGMqQYUq/gqD8cjZwmkcQF1Au7anc9/8j+VyyxDWjwZK1guRljhIoswfMy
wjtCNhMbHRDQ5ljN80ix7dgrdb8+wdbob3gNqXE/SJ3QIqukqmEOIdGj2aU/xtYz6Oi59scH/n7y
X2wigsB2gftD/xC1S+gJg+aZWuLM+frDC2xG6i2dRyAHsyf6PPowQxtDSw5r1HsrwV843IBE49DP
m26fcxpQwOVUNzt4uW0P1IUOv2qGAT0BMqbB0WtkmLEHkaDsCPaQBUvfGeCQm91BK2PiuHFk28Lh
KYTzwsvvltEs40ZqXOBPXP55vjPuKV4ERZ4c3Bd673amp5m26+KjKMm1EpGcaNtWNlWZ0v1jIo+8
um54uRk/vlXlLEItpZo2bERp2DAwfr9ffbQfQBoo3i1h3ZQ5aizi7BT91+ariM8HAnnuPq9MzG/8
8+3meaBEIHnGbCzGgALCbincCWGYTb9al7NMHCn42uT7lo4wh1bwoMsBJ76nV+8Fl8kExoWGG/MX
BS4IBaDDXHHnvATAwm/breMcPJPXo9lOx3x18i2ThD3xwmpHH0KwIkFsYMQnah9H0soFwZr2H5Hz
KQNUgkph+B/2a0AZoR3rK6u2x3wQkZ3FDC4JTVulf3XB+dDJV+HrTfp9mc1MS6JjVsWXUPUwHru9
3DAHqp7R35kiIt7YGrd9FVJ4p7CGCzuyzhO6YuqrLLsOSKccHF/RrU41agQzE38rwdr4EKYQaGxc
xdCKjIqen2Wqo9MSNvAlG8/P6FiaGTKofiz8zBnBKkaFTZIkeQCTtzb5B6Dlv7KlBfSbaHIXI5K5
8nJUlMd4ZgGxJycEhVu68EJ+wVD51SD+GxsH89+jlGRJ6RzB3CNMPZJg7DMk0sibgerRUkWDuRwM
qv4GkXdY/3Y0DmoFBrWQWonPKooIb9NMvmva8yu0BTzM3GblIGKpOR0JvgFyOiTN6uuk+rGaLuz7
Vu9FxJse4bk7fOlnAucDUUYb6LgSoW7PlgiiovEaOaw/sV/hLFfFlW3hrdL8MEJJ5XdwDJb4QiT+
qYGMHtpA+7bc719nsIoFBA+GkXrQW3gO2Wtnzvg5vwr06pLB+I5uHz1Ti7PWWn7XuplDQsQsJSY0
sMomPk498QYQaqCYfGjl56lpIOpm2IPWGexUS6LdfflZ1TOtXPF2ZKzNwpDrryhJqqJLMtOQXg/p
oq3DJodk1teUe7OHVrE+Z20wlYslhrbl5/ayrpEk2fw8tJjiSwoU//tBAtWwv23yOldV3q8irPez
VrJdpwRcZ1W2EnTz734cbHOfgiavkyAKcuTK+en82QdCmhMETaomqwaBd1J7/eBwLvmP4ns+jp/i
1kjaxNbSunOmEYQ50sLcAzgwRQJo2bP202XZ2nACx1DobWtc+fcJf6NRsvriRuOwivCO4a+GGCTa
TgsJnpd4BXelMPS5o2FsH2mD87WxCKHu6uEIfn6ZoPDOvEDse4bNgNk7WnQHszVfoopp00N/19wQ
9ACT+kTvLe1FmJcP+Fv3uNJ+8aXOiSDYyyGg950aHP0COXuacZ5CxHLEbnm506pbWAxPgoxT5wVa
9CY9SPCT9hyXaCA7sZQEIa+T0UxFv1FJTD/a9aN67nTSsYW3AEMJgYmJMaaRpakuDnqBboBgtWwG
J4yZeRc/AsMfM71RSYbtqyqiOv7eRQKTq10p439GMGqBELjgdwbimcW/aQxDaTJNU/AszyAyj/sD
UW4EzE3HEKPGOOqoO3c4NevKp7B5rmU5aHSQS3PoMaJFdrtMicDiEM99irXVCjQH8iLxkd/h7xla
kEXOxN9ktAwsCITv+CzCk+P8Wp3USmBZ2RjWuJjAwRdpbVloyeC889dOD0n3tGQYmLDxoGswWIoJ
rOqiffnejPrCcW6fA1sqzMBDSaOqEglLn2fM0lDXUq7jWyEXIYvXV0ZW67US1SitP4KBb54c4aU0
x2DeRRyEQLKPXF3j4jz6aaztp3a8I9QYr7Ty1IVcYy7fw2MO3XSgrboF9GH0dyBqXlRtZfLSL7Rc
5f4qYMFar+ZwZJI5pR0D6Ib+PL7twK8YZOWJtn0MIaMviF5bH6rEGRk5JNvYI46xia1wR6uTiG2Q
a07uF5bHsD2l1iPybStLFgANjxEfhOBwWyeKV5rygaSMAETsh2rc4yVqrTXZqJUlbnHfUSxw6tV1
GkuW5eXqHOOFikUfT0ceEZK5LDNxbeK5DxTKbN/pNCbc8JgixYqrW0YjnEeHs0GnPzQzrkM7eO3s
VwrHkHh//WN2vOmxvtl468EKAsPO1XmWyaYupQd7P80d2aQqwj19pCX++vdlkxC1a57jF201oW1J
Do9XuRmdFz0j/D8OStBK++lQTTNDOxQBlRQCvWLeL+mCkPRKVYL+hpD6r+BQYMVWi69VhzN1Sqf3
/AUUa3fG/NunUV6TCkNsW1igpSKw9PKkY89eJtO2Wh92UqHREtCQEPmPVnjUe/UZTycD57G44xna
I1Y6W0DMjdy1RPehqUyq4co2Yp7dxf518lKy5YWllf04n2o28hLiYEKyH8xYBQt7Yo0Q7o3Jw5F+
pmx7++IoHGXteLzQsyY61I5RYqXnBpL0knmVUjkUfkWo80EwiWPct8T8yj5SDggnW5athE8Y4lYo
KdJjG2t9iUBjOe1o3DDKSZ8LdtYID+oi3Dck0HwN51CvTY/do/L8iL+QyTCABNOsP6GEl+BYE9ml
zE+H+8T175BxRdZwQx3UhGHQkpatIW/9SwGhpdFv4LK5A5SBfc9l/GQQkDP/3m0QJMR+3NLDhH1f
PMsGP9dcofei0K5dZDU5si2jUGoxwgDSI9iWvm80GClRiYikDWRDzXiZ+2S2mXbUIs5ubP0KKUZV
58lbOp/YThQtcPRBHauzIOWXj59xez+5GC3OTFECXI/uWqdVFjnWZqtmd95vnXQLhvWKdaeI4CAw
QVZ4uVG+7HV+AdZmJhjwBAZTsCUzBAsH+ROzFYzQOE7rfnkO5O7aC3f0rOCBC1/qR3YsbflfCD9W
w71Zoan1jYJ1Uf9xmPywwGji0NIFxeugOa2WFYywVmEfUS4pvSWY7mQ/m20JPbYilKQOnSb60t7U
RZhee6udva07NA6rPpOxtUn6Z893CRFUfuIWZoSK5ktqB1BAVTO3lSFyCPAcrmfN1wBsJm+D6MgX
hUfr/Rll5UiGZf8aA4CPMyopG6ZDprboSmEJpJ7UzshQdbKfKi8UKCzf36uE0qkXaaqvL3LTtffl
aeHOnJ2FWAdiWi4s7I8jopVpfQ4TyeDNgymzBWB2anX/THq6WujZuSoptzdES2ogx1UKbN+94AYU
tA+o8L9fVkncHSssVqnNz+2hFhb+NrOrzkuHqLhMr4SEbkFRqmtNgsohXRf7gFnM9j0bffklHI6l
xX1ZKjbKLPb0fcuWFSfRiH73BVSoXJOH9zr807x0hpDubR6EUyqXuTB60462p4ib+REMxrvkhf9z
YnSkOQHGXiUhfP+FScGOl94KxIcKmjL92SdWVWdr4TAv7Zlk6Ita9zzFt+eSjeq594gXN4rzgF/X
3gxy7ab1we8YpnH14/qNTfsaf6yt9RG3yinBPs/MIEf2HfDoSonvLLjhPx90jvjBjnIUQ8DUaje6
LDmA+GGCesHboP8IifjTme78Fzs/G7Spcv7aHMaJt5VjOitWpHNrHpVV64eOc0BCVDQSgF+FH5Uy
Ua01SCyJPW7oGVXO4MEri12nzn/fyDYVCZQd/exT5Kg0hfbR14A5721/iE7Z6uKIIO9cSGQOY5x4
sUjAMWUkIxjd9UdkQ3TTm15cT0HlS2BAvVzcx7gl2C/swMUgS8ht/zLfYj8+9aNwmmRvTGi7WuR1
ihuV6cnC7DIIzcGySckBZNNLZ4tnL6A6x10j6r8GEL6vz22TdXsVGv1uDD/TFlLQq+kpepSFoQ3Z
2lOkJSIt2rPq0IJjYxoWZpQca/naWRZGYk40WX6eeWa9FnU+Ry/Hfyfs2h2B5xgRBi6Vjzqg0XCm
waNYBHIEVL2t0HyO120L+gpOl6zVh4WW4Hz1I62xiPmFJC/R79gtKeUC0PwL0d9SBW61Db7ORluI
yCuUo8+DUEl9gHF1s+R7gcM0R9jUcayDQLzeS8BDqvGS1wExLx3M9M7EXGCMyFQydg75+dLixDzN
X6uS5tEhr39H+IAd6NQn9J+c62bBD+6+JtDyFxKzasSh3hJhaHodrxIFAw6dVSfjTxNDzGzKsAj5
LV2Jf5HedhXKbLv32PsMvsk0zu+4yKZkYwc0vxwVsc2SWqqxmojjKm7mMS/WgXd5LSsy7aXwD883
nt5fAsANeR1WFujVwdppalMjrTH9LJGBj+xEJLIPmtjBNgb5PUvv+VNjd4C6WEEbvz7JrHHr9bw7
ok0YCwIUHYIky2bU9xlMuXjdXNzIVeoKfk1SyR9TLgywoWG+CGBORf6UZICKo/gEQpMBUop+MZwE
faoweKyNkFkEmRp83PZdapW6MEsag7Bg1PfUzecF9k/weH1287FZ5YlCtWusInVNZj20/Y5nYpH8
HAS1/HIBBQieO2LWWtUUw2/Stah8DVFQxZ6eXuEqGEETidgg4HKTZNs3PhjEzX6Bv48kWhidfjjx
Z+fv5+cvwQ6lWh3RimOP+qU4NY4u0zaALt2wftDHiTD26/dOUCIsBNltKlnAROCNMsfuczOYqwlY
aGBqXKfKcLgTlG48wo2gfolDKMR2JFksh7QV+IFKHW1BC4BdHtbsa+1lGCvvanU4LvaMIqRdjxdA
K7RuI7NkEfqQl3n4N8v9ti/tm3H48Tbxw7SFtjqhkTBmlnb3BizwfJZ4ntNcr+CJ+J0z5Qz06ucx
CfoHCI72SaR2YBYU9L9tpTPvZ3I6WIreDWbm8AN6a44L0+5pC7YWixDrK422tvcyqABmAWEM/FtP
i/CWOx9rypdvDohWcg94qHmcbvnZjwlYBceXx+lfW5Yti0MAQzonOTnjlWmApYSP8YlcFPH6VSRO
dQ4/bYiyxf71vC0ZGb5oUjEqu/wae2Ei67gqhD+Yi+nSHMwBnEPNzEPXbgEsS3mSJvJNyiprMYKt
BHXCbLFvjK40preU/jHdMzhsF1bsdp2b4klO/Dnnlbz2lRKHfz4z2XZJ0eOlhTmjVA0c4yITkUrZ
ScZb3HRvJOHoAgezI1TV6JKBdK/asLb73jVL4NfrbKyPW4kisqS3+UQXvOBmnjJzrOCtWJ4gj5M1
C89uAlC//9JQ7G7TCIcw+FRkMTiUkx4xBfIK39nPp2gSsgKa4PbdmWYRyzN9khSJdcxCVXZfVHT2
IwXgewsWRrPGMRlM8al7hDVnUZynAeB1ZCydHXBG4eBYqG6Y+ExL6xvae51MtRJihRAI0dZoqRJc
Cm8KokSHaDbxvNWDQCR30xdHsH9PBe4/xaj02bPdAQPb2WF28kvYtiPFOGzwPfinAk+TAnLyvFIZ
UeAlD7fSthT4B6PHivJEWnFb3ACKvVLZkrYrmAvvzQtJ3rRlxNufBhnCHtNKQqdu6OIHT0G3t5zF
WbfAzbh7fkunkrygN9vAij+pZ1ZirWH1a/HrzJB3yRCALy373+g3XPouC/af666OtuxtRAuemalF
gq6oy4dzDxp4vxvEHfbR9GzYKCLHQsgSDte+98Ifpf1b6JQtUL6piGk0MaZKy1ZL/M8zCg+fGfhg
YXgA2KeP/jm2Q2ZOHbs7pTaqLnoKdn0r20dJQfDVLZDWychgZPn1Ol6vCpgaHNoiFzL8L0AdwaAT
mp6YJwimVtv2X/PvJreZaK8rcZR4aXMmjZ3/YepSDmDzuim0r7EwyLwgLLCIs+FfCHhZKToeYBRc
IpTJYzMIoE/IJtQk/nd/esOJ/piqszaLlmL3/XazW5jms1ky+jbsiKJpA+wfHg2LLVMEEC3jtU5T
FBjcYJpnUejW0gOFNYDMKvOm9/TDG3/9bkArX3p5pMg5PFWAi5Clr95Mdq34M3D5BQbyNLe0ptHD
F0RfUe8/RZTO1SUu16MTy+cTdKboebtsr4u6VdwAdSff6mW78MSwqm4XSFCZwcpEN1qpJZDnApIH
KHJJCML1KmdoalpTjNWYwtWJ8fG+7XryNm9BynMLETDG6kEEva1C2aCI8H0UaZDKAlFTI3xmMux8
7nZj8NistSHdxnnB7SdhGTwULBexaDSccB3A3Qj7lbRru/ypxtihCRSGUWaFQzaHZhp0/6/mr32E
pXXtZMNu+IpPRahGNpJ3lBpqo460LPwwFyV5qRCYwImEYV1g39wHWl0bsnRz6z8C7Q03e7Ig0npL
Wnb5OhbySN6eVv6WnAFlpaMo3W6Mw4BKztiPzxt5NnDVzznquPrJdxElfUKwtrew9+poJA+3Cuu6
jO67MMkrOsGB+S6ykBBJc0MydoUJHIdyy9/Q42mSZRFjBmV3mvt9SRrI9K/rY7jG59/7YGERw5T3
rgqcx+RbpC+6rthZSlF5RblEECk9FwCcIMw4HYwhLYISwsLESt2AjqqlPmnTuNolwrAVDgWYw2fo
vt8yzXmRL6FNbG2+Sem6F31m4xTNu8+5b14jvX82k8LHFlQpWAlue8aaN9bDKjC0w7mgveag3aDo
TC3l+hFlt8XpBWNfa3K20jZsExtoUvj15X7LuYd4UfchY444bT499N5wjZCjvp4nM0az7peEX1Ve
3zl9nb1ZUPD78nEw/VMVRRd19dOzkjIMtFeUWSyOVUAKvgt2BbxEgYiNfn/COJzooW7ls+EHthv+
xiFY7ndr0glK7ahMlIgeaE8jjOGA5TSr/piKsN1ucKFg+BJWjDPEWs026wduXA6xBO0dIJaSSOKr
G6xXYmY9jL8ID5W0ECZ5ma2fnSxEAcO0+C9kTtrsUhIjlQvwhMgK6I+H51KAGCrCXgZsSOTtMDCS
k6lgLB7jOc1xw5+Nds7e1cUMdWFfi/yMayrFc5JVLOSn1SkgoF6VEjJ9ZJ+IOxTOrIVDh3+eurEr
/WUys+5znEFTFT5USBwuZUYGbrcJxTDNM28dfdxoHpPqsNKu8cGbHQ0EA7X5m8Eo7FRukVE3ym4G
kNQeVod6TuMS0pa16lxgVr10zj94MgP7y/TlBgW9fJmNR9Ap4PFGomNn6Pqnr2Yqi4EjorMJrqkL
NdnLeu2GTv5qNIUk47HtLiVuGBsg5at0pNzFkPyExAg1/LBLUNa6L6y1V5JWSGwQjYcUO3A305LC
toZzA1q7qATnPA5O0QMVdq4nLrfx3uoquFPNyET5xjG9DZqW3tc9UG6fnuDug/9kiW2qVqGcHk0r
85oCw6PLYQYHOYbgLeo+BP5HV8cYxnis+U7Tpd+vDXmApag9JofLBEh/9g8ZXdlePB1Db/bS1ihe
aoCTAK8Q51DxjEvEAEj6wNLfDpQWxsI/b6shIOpsr0nJU9x9pM50wmEh1GP30OmIgK0ik7f4k9GZ
BV1rPDxJprDg8JFaLEIJjyR1aXw4QROmzbR2d3eiuPlxDvEyQMttlmKG/2LsLYRbCVvgFvXsNyiv
2ZdF/rUkkFawtq+Ca7VDXUChNlCs32rCPX9rsMR5heqoeDXqhjJ2ykqGVIzAZ4atv3+/BAPMwIhT
LOtnf8mY5uQ+N588P6T/rNiD8MTJxkCYAf+vSgM2d2MwmQyjF2pp52HghT3Pzk38HfWDeTSGZm0q
yCgaXHHcwjW2xEvazzQmYS0rnNt6PhhE/6vi5/uhRffHNGmfkkzwzBwUsNJQnIEGGsHH6V+azMfM
ZljySHihPVMpzUtdhrE68wcVHa7TVG4CGGvLjSX0LtZzTPHvMnN2UrYA7ZG3PgBbHo9dxFqSppUy
iCs4mTN7ilOzmObhpoys0lZXiTaa6m+zOJ7fBC0sm3BZmyjgbokBSY2uHTtp249hEnxoGK/mA7DZ
kP3DwJCMRPOhghfkDnd9y1vfLW5t4PmwExHofZlzz5spdoo35wEnrXuY31t5VEZJV+t12fZ7OL1M
erzyHXxyLj6UTHiqB792cxzUWjfYHh4iIaEVhRG3lTBEoeAM+nDreb1atrc0CYYesAkPZfs6ND1z
xYfuQbp1vr3Q2OMTNdm+FYiTnHv5F2j8Wv0AYSYXfnvRVisUh72w9cVQPVpdRFUdQtNWrqUYMZ/e
UZqzqPU9qwCvPu8bPKNwBrREnWfF2LQFaDSlH80iNuP3ItndUvkmDOqv8kICdi9l6YolvMBZ/wxx
+sywGkECZmFAmNk4D01omzV4hoHjyDq260+hC1K6zFgGZ3AXxTVVARM4zibcDKdZ9OvhqO4r+dJ/
RWQUq3RllMijdm0f02KDT9SpRv5H6Jw8/Vo5OoFCEd4lPqaiC+InLQ6BkwgyotUr+iJ1hUtHLxin
ELDOGtVB5j6viuzYTEch0lkXjdc0Pb9y2fiZkibTEbP0Dzw9e2yByCL0UwQgqLQbcrA62OnPWeD/
bGH2kMEaQlvMTuCHqSuBwk20ur7Ldm3nuRDLURzvuNA5gfgqVqV545bJ6e2QHkT341krxyOPkma1
EnLMtNCD8+3y5GkvFBq9I+qpoypN8uoApv6m3P/dR/A4V4zLK7EgpU6CTja7fp3kb/9JMIyrzGfA
xUJlfBYxtv+DYT69UZGzlDMo0ZEDORGF22RfAiWdpbyg+hHjTrGdeiIZJBEm4JHYu/uqOauGBo0z
4pvaBBlPku2nHvTuCZmoaHNMLV7WEZY2F+3APVIcbVggaC6EVad8nJUE2CCDhc+jTLNcSjbX1NgB
60FWosrLqXpcEECGzLQ+xxvpYhaHmoRGBnt6MG/bhDtie35Owz2ykfsDv7pYTjI/OhF8ihJFj/E8
stkS6d5gbMsDC2bRaxa7+n0A4O06CjiVBYxsuPX1tQTq1YMHVc5tb7xZ5HSmcLGHU4VcLRioSjia
XvHxqpxPR+fiKvoA73wv4+TWIkxR2JAmEYkZPjsIfRlEjJZ9TMa5e4Hcfdmo3zwU4biHKgtOOaJv
bOLQf/zvFANWhMsJO3Vz7Jy9hxaMm6xTejwYtXpccvFjnQe3h4BmYvCfqWcz3ZpKlFtbzo/mSk4K
p/GzPK148renMeeYwdpewhNqkNPd5KtCeY+uC2WB1X8VWwY9VnddS6byga1pJasvIJnF/6lQ5S/N
+faqIQncA4SRedZri6GbDvYJrGxZW2La5cDQSrk44OaA34sN8EJGqnkPFUVo9b2oNphJPnWfIcnO
a2Gn9tFsav0biJn0hEcfBckHq6qazsF3g3/gYQZEA6Hnu6VkORbPzJsFjVe6MRw1EGO3E5hgib8W
JtyfXA/1l+gNG0cBfjlBhn9doNhxcBBzq8nETO6/drvw2gVE3CqqQG7D1itRSRrqdqESKRCGrZBM
hxJ50zh4j8NQN9j75gL3GCC0JElbkumCKxvcv2IlrrTApBDw/VPnaFGKVUO9InH+8QNNHfaWLpRW
PIBCqp0fl9AUr1uOO4eG5unQEqhyl+4mj6OQQtnGYhBgFWlEX0MFNy5Uh2xtohGnsbgFQSqzgIJF
gGNMyKqOIxhwXlKODjt37ugFm+TIuMTyLnfRz5jq7lRUqQvXVrpz4imy/Tih+zI/NyF2cJvo++pR
kpRqOq5KpFuPxZsMJ5kgVt1Wy3++n93UlzNLSfcirgnYfmIJwSnJJERlOnnpU3+OqOU3TK/FyVE8
IvkYiWOx12KfDR5pRgKpFJgcyu3tgGEYPYJf7DaGhABjExzX1o7j1iUqtZJMBmnBYWdkEMwQsnWa
pkI6G6wy9AvuFH9ak3QZAn7cirRI2+9HnmU+OPIx2GpkPbnCzcfJZhmD7Ek4deeYry0EEutFQrg8
0FWmQwAcPfK62wRPMuM+RdLq6sGHYuRf7TZGVm1YMjBm7iPABtiuI6TpbJf7QvLTsJZ0be4Uigia
VaoR8tZvoATsxN5D/4IfKASmmBPmUscgM5Kj8guVIw0MILtPwP2c9TwSA6MlLlYr2ilSzb4BD5iJ
q3NAQlYWQfHVxSvnNwc+R5QGOa5g6nciCVdegisJWPFQPbsG3ghInpx/jHFg23DBg8L9lgpksbp4
hw1xJDQSzKKk5LfACRhEqwZTGxIYv3tLMSWpqcKet5R+bIMZIt7P3KnOfgqjHFB0rvYuBcRdr2uC
std0oZq1G1Dc6j9iFDSo7M16HBfQZkG10UkZFnHuIju06X/IkD3/IuAYssx0gvKfHNRA8D6EwiBW
Z0xjACpKVenFLicltNl8Gkf9RUqk6BR+pidAO0vJ2UgV0YsgfjrO8qJAnSnpgM18jHCz6y1jgBsy
M197XkSCbw4E0ZruI6m8ppTWfuLHaM3mnExFGLsqTMHJJRJpAxikbWduOJSZH6c1pK64j4rPicul
mrOVwzk73GxujC7ElmhZNMNhPS2w0zaZS8SFqzT3Eev9DtJljXpapDPQpSqiXnBOkAU+R7wTvctx
GJceJaU0U8crs0kj0YRsB3w65kqYZljBNk3E42rXd7E7FIP2QwYSn4jw5TKGtIRFIJTPdHC9PQ+Q
ZouekEH1nTRfzEk5P4ZK47FyYX77Siia7CHx4QhbIYPeKGd0Hb8Jasiy3SA0AWurWxfc9My3Nt0g
XgRtiOrCOjjX7tklfM/DQNEXbtvntUyzS37qwTzki9nkYtCJhJuPhsJiRlOGd6hsrJbwMeNNT/wg
r3UeEnIZnJ2tVmFeJZ219NfLW0sVGzqV//kwOW8C7aO5EL30c4zXoKUV8tBDJbu+dUm1GxYrCkX4
BdWap5bKAFAmh8nscMx00O/0EWWfDgnvxvxSFQ8evq0Irf0opEwk154hWgSGeDNnKc3V1xHT75UN
evxxSP/0jFI4B5+YKxM4GWexFHXoBhNaNvN7cNw1JKX/QYQJQbbiEN59+MRIDUEHtMpb+cb8HIKw
nkGpwmNP3BbLFTc+hzqeOrPVBPTUOgQOQo4cApr8Uvddh+IDGkhe2mNBIxchSBIyfvbcb2viD6bo
21jC8W3KDoMulylMRqWg7nrDw/VYUSrL+ylU9odtOWouBJMWA99AzmS7eEsW91S70mW0NOs1Tkum
Z8VV8gYANuF8UgKIsI6kr+NFYYYP9KXl8pEVO36QALKEdObxGjMIu7DeYECPJv2f4cimlIoHu8Wq
BAK0tcCIXGkLIe9AiU3Bcsr7Gf+AmHNRZGpdCNuiKa8mx3HWOzlQcOtgADyOClv64H9bWiPm+Hbm
DzFFFb1c6yF9vt0Z8TE8bF8H7+mf2Ikyrf3dRIw5015YcJH7aXQ4WirFqlmNOpGg0NaQwSUMnQIs
dbt6F3myCyEasYYiCnqdUovyU8sGuHIKzKFSJnM7kYJpF/D9qWHpkbYC5ssoN/OUaP2z7/TJZkIR
WuToK63FMj+vSV1DUHpe0qlA2ht98KqM1Jxp6f8MZxje6IVHtoWerpkC6ZqwnnAS2XaorUSrvS5U
IMUMI2TBfE2QSaEIjrKqJvfaXztdqH2UzCYmCShyrGzfKgEVloQV0VhQy1JJi4nLDXltcr52lKEn
INdLhuVkV1LvFAgCrMuWoyag3rG+dKv6jICgRg3jx+rYhnR3vXnjc8OfYfkMjNTSkSm/ZkmMtVMn
XqgwVLD298qWG6hvSeKO8L9RpESQAADyvGTbyq1q7Ql1xEaL5myvtAnTlNEkS91encM+tZ9OPze8
hhtodVAzyIt4Hq6rw25C3QkKRWSO8vUUHgx8kw926NS3ue10/izS4RH5508KO0bveu76w3qJ4MNS
n7Tdjxm0FLkbg6pL2nsHuEXVAgmPuSnXaC2S5zmDrMIuSq3YAbmXyFOC5K5wtkZl8EYPcmNfgwlD
PontQ5GnwopRtqj22ViwZwn3rl4VeDluWV8k+lzAABc+n+p+jfmMAKG4gj1SVh2qgsDUExjpjCwl
dc2/tsHMz07j/mRriFiaJiJ2TAIwTGewbFTiLey2mp9dtFZEZSeVyGw7PxT20WpbiyKR+xSWf0u5
R1X741bRQnYlLnJbif+L4ru/CfhG418ClnV4V0+Sep5WBz9+CeX5NzIc3Kfh7Y6eB2ZYRZTbDBWk
zWoXjhuBHeQT3zvNQ+B3NUCAFT80l2HIkXcyCyh+HyWSqpvSmFU7jac/8J/+QwpQDPqvbNgHiuNg
S2eJRCzvDi8aPKQOziDvYCa+os81fH2zbNOUWU4OhOc9WvSu2otxzeQ42nB3g0pHjzcTAtSdyzsB
xzGfUnyLQJuRNJt6BuYTIOfFyk+IL1ZwdRIqbwW6jiO7V+/MEorT/ou2jqhwfmHjPkzrzh7zTih3
M2jFTP2G91BXpXIU/h4wKYLEz40Pd2oTEnDkg9NiROe6qyv/tYpx7nTxV5wpXKwp2iTP90zwhaIM
U0v+lUlnwqZOFHQxWGMbk4NtbKxcBShzVG+NT0YC+Hbej9ROmVm9+yCYg8kBjbDDFDBfp/5nGbHQ
0/dcq45rUy0c9tezTl2gVTFo1stBXx+jjLUaLXumcMQYt1fLfc68DRJiPaHnSfozZI44IZFiO1fp
ycCnEzexv3MfJFd8cZSMVQeuwy9BdyzsTY9cIrFBzoO4WT4RojT5jFtJa0Ou4q4wyymJb91w4HXn
1ZUUisQiGlnZJAzFjr0WV6KCVhtiVNxnkMTpDB31e/msttdMiT4Nu58j4bHYYrvR8D1HFejUetzl
UuzCzeDznVp7s2/zA9Kj8J//yhC8UGKXu+/xQjR448M9Jc1g8gQhMqJT82f1eMchRdlBHesjHSxp
CE1qGISOaHYa/rdOx8/jS2HH3fiVsQLr+/ls1pmsUekPnCpC8SUsMJR+/yYKLV1C9cMG+WQzRKy7
uZj8nQsovDGa0mt/6rVSM7nuQcsOa7BPPjKSLoohuFR3s4JFey2DndHrn3oa5i7HQUs+o84uj3Fi
d05qBkIOFJf3r8tlVLER1Yh+blSvQrJc6Q4snjILUcfkzm4nbE8Yuw77Sw3nWZeKVtWEQOCXo/lg
JhTCrF06rmAyUJBPKcX8mn63dscEfsBt8f5R00Lo7TwFD36C4R0f0CEuva7b1h7YugJqNvgmzqih
/YG7Xp1dkXZwtdQnK0nkepx2DDBtzgdN13T0vEBjGxGozLdnyufzHzlRl3BY7tZrlkPprohHi8AA
fW5ZzhibnwlMcTIj5Qlhcw9OicFSx0+Jkh7rbwace5AtwCMUcNmcRfbNezfoFlzzD2TDO3VezZje
Ei3OC/lknt2cvTzYX6Fo5DG8QdFtwnzVYH118QWuQ0+nrCHOvzoHOfoBCmiv0JC4nq7n5UFB7rlq
C19h7OZj/BPDmfLkZuGz+J4OVUXPyT7AJvhjHXcWWEAXSenT/OBq2BfRYJUo6NcUl4TkTOoG242T
DG8ZnRyFy9+zfdk9RNRXUJm02YKs1t/0LfNLnmHL8odvVNu0e0h9+K978NH69zhd7cPCUmud5Rkh
5eO8P88g1aiF0KNHmc7uJbRI6ILoizTSvmxklszow2ONt//cQcqLitR7YKrEXFBb3WZOmdhsIqHK
qWMt/OZyOjSugy//HljQkTfsXct61x43Urd6ioQkd6lyYLKGCzTqZrBRbsazy4TQOCRCJFf4oMNu
OTt69cql5yLh0XH1M82+9gAFZKAAtnhj6PsKybbDlGon3ppvimRhxCkIz/e6t/zwQcZz2LpM7Y+g
iTHcCGYTFgmGiUwOS3ZFMbVQPOfeGg1VLHU6tHhSx9GEuvfzB05OkDlhF90A3bCYFcj5L04ppClt
rW1ZOQ2GW+1eZ/+Af383aFQzMVzSL9Orvl6d/R/mFu1rmhdvrc40UNCmYbB1YNDSUIVYh8zSrjxq
rlB1utTJa1iaywkh/SCIXc1pPXZfSleg20IcYAol1rdDwkNxpLERaLriqmH/bZsXioRecS7Dq7cM
E8djZeESXZot4CNLUuWN1R5ziNCRxXhJZhMMY0T4uAXSumvzvNbc/8SmIHkcN/1JlBog7wa1LzeU
Vy44xhJmae9QkubcwEL2QL23H16r/4gKfjzsXdo42VZudsXAHBmiog43PZUNW2xFEs2x1d9Tl2oo
TE8IzLTbUfiU4i/Juajw1cPDk60ww9oBsAvtXjaVtOoYgFzq0tOctFztYNBM6dWUmhAdHHNuzWh3
GC2/t5ubmCL0kbur9mheuab4NfiFbqwn2JZlrdM/9r7Gt73ax0kiAgycM4btAyOHfVugzF4hqWfi
0LnYhOUQwZDQxTThrvDRdh96LkHhJ8ifL0B1HiH45HcMYmP0NB9ZZ2mCbSCBdVfXPWZy/pzOl7Jh
nVt/kM97aQWkyi3aBwCY6UIQ1AyrKfbKy+cBTgs8mVwZC03LYHVgaQhMChS00qVsfoyW2CyT5AYj
W+Zu2IFA5y5g0h37AvAcC8jm1ZzJ2Eddz1Uw3NMe4dPNN+wpPMFJpE1Y6q6tPH0ty5tHZfEEPKXx
sQGChMrxRix2uzMW7dfOCAk7KCSe32JKrkrOAiaS1yOxXSUECHAy2tM+xaPzuke4z5QK+4LpwQR9
A6ue1pAgtAzxGj5qZIugPRBaD+NpW4+fCiIBll1iejXZNnMU9fLWBJbCuvWd5t0CdHIYDA/uZhWt
UPUITZUr+OSjI28WlQ9HkRJJymOVxReXUfvdFWo55nKXe0MmmEL/cmiFZE44/+A7Y+JfWS/SxZnt
8bFx3cjM0CafL3nvvlRxVLtpzuFxg0EUzASBkPYwiUIwB6RKe6x/oVKhWmd04a7R8yZtS7iVsrz3
/UtbpAdtpHNhtA4UjXklD5D+8GQgj+88VssYtiQNYa9/FJHqmuWOGO7vfNLwFUhm+ZzjCu+Ke/YH
FWKBxA+2FZu0umFywEXBEG3czw6RVklMPyc4Do1gpBQi7BQqy0Hg9VqYHNxOQl1cEeKK3mejYtkR
Momy2cPkFiZ9G4wU3ftVagEN4WZgbAJOf7SwiJIlP+oCKpxABQdxLGp0fjO88YzlHP261g82WDmn
LdAKsZxbmHz2FFXC0HRMYev9GNcoqEJGyFLWgAFr3SAODQtvKno91gJxoTky6EDu/QkO3K8SQZEX
CfNNV304slW5Ep8McvLWqxVRhASwxW0cE2D/mUVzRNVcjUM3TJaWjlNnfbXgTx8blRAHn77t1Aio
gkGa8NsLoJXgTQjbmV2U9s/uvdZa91P2ulEoIb+ZbB+dUQlZ2936Ph9n7S8vwGxI6yYg7Rwc7NOq
jSaOTbu6fe/qMJ69qhoZyVu5Tn+52Com0+t9CZxs54EI8t8rpR34FR2d8ObDKayh4i21URTdy+La
Dk98pVnQOnL4nRpT9Aifedzh0rIk4Rk73iPRgtl0aCAcNimYnkx/SRP6ohBJjDN2vVteeBg85Hsm
DM2KQVTv1vcQNSrFwT/3weqSdu9PdKhvR1/WIZ5AH3LDHbWiSLosWPi2HEOOUJQ0q1MJQxEj+kuE
4ejxcUNSZ3woKM5Xo46ff84j3jEKOhULtz5Ts6zvje+Lnwarizc3bbJAj0BFT2nH+VeM9vqbpG0C
9y0eyftVoEBUaBjFN0SK3s0Oncf+9TdPqNYP4gajQ5BjWfKlDiBCH81Bj8b0NiYw8cjGOFEIxRO+
Nf8UaBCi8/yavBqM2GX885vMH/mOGaGbAIJo1tIZeN+L+xKqyK528AORyTFZF0dey7bATuikOd+A
z1CwLqhOPTqEp+RaewPkYcNNxykwmkqZROyqaDOALlEFTVap2MRGLYe6kWlyL3rbtUlIR8vJZABN
OQ0Hhk77E+7vRcCEnPp5txBKPLE4zxnEC0Bj8V0g4k37CjKtGg0eEJHcS6geOcdfN8dgMgEfXSkR
90fI4ZQ4Z/CAVbRz8UIgQ/xlrymaozonqPp1WrOpfjW+OZBPdVkSBGQsxsvjlSpSBllmTMqLdxxa
Fv4NND3KUG8F+bnkLK0M+ubMxhKkhuNJHfCEBCLYvKsGD9bVX3F24mqCh91qkcBM0mabIgYG0YJv
LQYLXHRnpeMy3YwztxkILRfGmBjnd+JmrQ1XMQZJzyK7l0cxJXUJokRpaHdIiXmhlTkZF2OkYaRA
hWY24IyEIYbldPGKWXL29XwbVS2vNd1yPGscSbDHOPrsIUK2bOsmecTT5RqsqSG+GNIZ0uTwwCjq
O92UK+iljZaquGgzjVV48zFwUUCoQhWTE3z9URBWTSc9iPAE+hbzVjf1t6xT/veVWxWrMHYdRjZY
gW6nm6DsmapItIsczcIytw19JauEcpK+IBGRrf0VjMAUXY8dRl+o7C4rPJc6d6dxLWpJQwGE3NOO
prRsot6WhzxIPs0X5WL8bI7enBnJVdNvSXf5TeFi3veMyV4hVxYnuRU15N7wta8WU86NW5YokpeZ
n3DQJkJEBbYz7ejXUtDrDuYxCAlHnM+VTqbqSyP6BItxTHtt9sxjnd53Ps1Iyu6LISG1waQdut0v
6NBjLdgofferWGlx8DYM6wbPsvhJCKXNOad/vlwzA6yPdc+K+hFL5z2FXhUB7hTgDVsr0A8G4Jfw
XjP2K7j+L7Xc6UL5iUE3Hv3szxboIqKd7/t4/aizTL1b+OSzPymSnUd//Dx8XlYKhhKdgQ87T8/E
3KMYyUqWcDAyJRC5Zf/QJgoJ8WbG/MOQ5Wgijr69sls1mFFvnvE62TPnd4lzut3KS+dLoYnjDbRA
ii+/vzLeVljjbEzG9mUWWCWhC6MTVZ35wdaAPSg5baKSMzlj7mBxK0ysWzYoSa1WtKfGoxnMxXVV
Ryz0c7/xmRP+dK5jWe03ajt0Pl5bAhF5qdwQ81fp1ne8ynEVCChpHLgr7834oCobFUatJCB7FEbo
aCHfhe/Q4MikVME7Q/slOP42CCvOq3GxgIcm1thmg/fthAVh4jmP29UbHYr5bB/ND88BHp7Ec5eh
QwbK6y2Bj6UwJ+GYb1sJE7TAQ+PjCc8PUqo2lvLNbiVWljbBbjeQ5BbNaZ1nMn6Gws+Re7qUenrN
offQHiO6Dyp4eFmHimdYG+8Jyt6Spubmcil3ND6Nxz9OA7oFewUow7TX7khpVwVBy9o8ur43lmg+
9lJ7nT0oYN5POFH0KXEQZiu7EtMQJg+tfbds5ZAG9mBzyUO5uD5xmMiurJZi0ozDZ+bBbuSTLcjP
TJbUkw/K4r8V47vSBAODyBaxgEao4sdKqpigTiJhmja7Wj0GSICW74N47gVQbc57F3jsA9VNI2Ct
RUu3MDahdMM2LXcsZpen2QzImytY3LXenja9VmG6M4oirDSeVKq1cEZSKMpmPsSM9wSbez/DAa1c
NrcJDM87fAqa4L6KwvubUhwIqDFjESbmRuiuwz8WUcKKOnPaixI31TmFfRIi26k/vuCOUCOABp9T
kC5yzXGuqVIRoXHzkFn5pA9GI9YEQWOxV64yk2T2PeHcgg2KXSJyxYjpLHyMhVUQZ8pmOkW7OvzK
LxdIqfM5s0aDUuGplgLhZsPlp/Iva1muDNXh71pk7rLMtS5jBXND6QdUyfPvLQpzVUb0l56APUtc
Icoh4VRqHHxtCpk1yASf7N44mC4bYv4ffBL0vcu8IiE0WJFSFBGvEQcZKcNdkDOy2xLuGiX5SgcW
yEC2LTnxrI4X3iYdaV5rpmqEpN81EzyC0U4PQZz/i0b/bllFlkBsRS+t/kT9Vm2TYBuw3PqEtqSd
IPz8Pb9QO4PciuVjsgI41Ysza3tAngm0wxqFNyQ1+Mc7sf60CLei+4o8sbxbOQKzr7f0rssWeOrn
Q/+qyoUNr1o3uXqV6krbWNXx7xG7WEWzlcoIjp4FNtj1wHOTHj5sv5ijHBNaoklY9zMlSQKXcmsw
hv/CX04PzxN0kva+XeT9YiUaiMJX1wYTnLlb2aVHEz32X8TLSKWKwtzYjUTPMwhWdCnxzySw29BP
mf03WDDa21U3g4RC+jD/n/We2Swik9ur+hmVdAS7UCO5brUup6kuVg6ZRvzjhpeyynY6BXUPqXxX
0HF1s56V77iy2Uu1kFSkBmPAGryTAJ+jrJ8B0S165CfkitW31SEd+c1n08B/m/5tru2yv63sN2tA
fHQLDSWXnW/iF1q+UNdSxbldQ/8KRKISzW9ZLdXE5+8ZrNV6UQ5e+hen6xUKNbGhUy7Zeq9gf2HS
DAC3hkOwdLOdmrS3oZZ6NW51Z8U6hN3mIpMZOcC879629aD67r84JAU4ozvGajuIPMIKEM7CL27M
tCAN9cs87nvIMabcprQn7tQ3v1h8H30fXAN36Ibncbj8SZIaBS15cMnHizkutb1IjSm9H2da9j2Y
GG+icslLwVtJA4MJnCloG/1in07PORpK/bBCGVM81NhnLR6punETvNMr944aM9+Lp1CN8lq5sGZO
5POxJcDgE1/ryJ5YFl9/9mfhYGjS5P2MBk9ziHf4cX1deGys7/szWfM/ALUCn7tNkUs6Z7XSWW4c
uP8LZhpbigC5nU8WtReA6LIMpmkQ9CXBttt50iUrSK7oRzpQiRIwmhJlKL2z1xRh52WC21/o08q6
S7oGWnk4wwN+ZCZ+pvUP6TLJFCu6fXNDNP3wZNztb2wfUl333C6WvofKWGLs/+QvehcCNowuH0gU
/x6mu/DikbSRKeci3+DpfK8xwd9U/jUBjWjQO8zpEy7Q/SKz8mkyyRMdZmhFqZL57JRBsecE7fSV
2zApBPx380aTtJi613pe6l9Dsd5tjS8/92n37aptMIDQuWBq/cifsTvoiwkWj6dSxiQT3UhFZv6S
iu07palt8XVLdFauBES/nomyHLwefYjITh0KBR+Y412Ra0nBabuVQ2g506kPr38S33JmBBTkkQrb
WR3HoPzoG0Aaw7Mxrdu2fu18aug7JYCECb0mamMBElqrAr0SRd9LTYzan6sTMGpLk5DpgycrgAsn
izO/VgXzciEX12805D1V0mYmGMGqG6ctzYxzQvAOYIp8Wp3a5DpwowP8Wta2Q348PM9buKJx5ZzV
xN1Iz0Lj+/1CjcZJTqpHq7XqVDcMPvl8nzLEH/SOUtJMJHxd2OvGT2+4xqLVuoWmDCBlHwZffqp7
OumQq3RRpTtvBUjQHeDgdRqHyeE0/tecxQfFzoT5eTPEUKWj9m5YV+VVIrNL2GWBJv950Nq32qJH
xvuGwxJ0/wqBP8MB/PSsL/r0wecdF/SmwLEtFuDY2LLgVXgUiDuKWjRxGIuCQTAFhVvBpZRT1cV7
wh/vIKwjoD8B8Kk087wICsTUXBdeksbZID8Sbva5TUPafnvctewoCiedsci4S4iZAfFfvwgI1dJv
oDV8mz4KechadPWkWB1Guxau+KEcLwOPHc66plB7c/atPdaXmuWWmgzfUP1D1ZoOM5HhIi7mjE65
OIrZdt+e+TJXwirwrwjKGBSV1N1DhHpXXMl3YIkk62XiZr+i2nlsuQBVYPkQgJwLwxnvYCWypp+H
Z/0JGTb/UPl2whpBvL0M0fOYWKccVmIp1XGmnUE6GSGPjCHju+5ISBogu287IVHOK81Rv0LNJgqT
N09/asbRBtXLTrJUOufOEFQRnioGWRQ/UctpNQs1Uc9NEP7TA+j3Zzkq3upr4ZVeGBwa8a1be2C1
ichQh6a+QhdNyJ7GPlvn0nHj3iFbPdfdkzUroPDLxtTEjBSLUMRIXs8EndGIH9ToCaN4zzAYo/64
2UyfTG9RFzHtGmH9K0oz0o4qDDiaMNuayVXyRIfnhNp36rRQJu73OuCDCztR+u9C98iEqTzMB2XJ
G5lfDUnSKYQ6LDGEVWwvH2MYrGOhU7N377MRIke/JfwQOk/5LHDZxXYGTBWpMHCoW+F+UO2XehVj
LzzrFvWGoPEAFIb/PNLTpiqpby+JBb6j02IH5GSjwAEjYjCHvYroKtwka0INvw/MECxgptwdA+Fh
M3MlL8HfNjhr42hfdW4q5gnc8ewhT46oiYmCrVocaNufRx8q5uYN3k9lAFhoa2C1Hp1WAHmtqpTr
j+/QBerkS6w2NeNTFOeMCSFNERKXpILF14HhfTzoU9zNnvCgas7Oizpl0zI8Dwc0TLZZpuvqmZnd
gPpdWa6XadNKhlr9BzZMgZMk/1lOuU/d4CBbSFIsIkZk6PEfDvZgbJ7V5fnGwIaMNWGOel6JfCHh
uAH+VGoyjj6eJr+m/pnNp1FvOKa1zTJEdY6qFHdM3qHJJswZu1vxpyYYNFxXuY4R096xrCNvdHYH
DS3sHaGKOy2GdYdkkQTKmJ1O7B546qxJGD6C8hWqptOCC02ROrhudaIVuLtSPvK1JnqiAC98kr64
lzd5VjZ4iJn5zr2ufWL21y1oc5QYxGZGaKIjEdHfooFgYMHcpMYuU5IqUYsHxSqVYPyPOVdMoyI1
AyytX0oJm0HetQyJj9XuXNRxynRTlnUsgwE03dJfTFrVQLkZItz2UrIPtG9XVQh6K+33GSc5QUpi
B1acGBCFfu7X94fqcrhsAPD/ow6wjiN/WXh5HBiQI0jszsjsxiVQV6cRQTnvgfkmbsxE5q/PrvqA
Ktku6k2dfzX9ouAMYVhUWpzwhOsrd6JSjhpQ8Jb1NTuvcv7VqGdOCJdNrqt6zrWL3WJVFHbQYZP1
5Sr3UXORr2OFZt/LdwxzYgZhFQaflbDhI5IA3m3FNAld9/3mepNr5XOi6LuO6rQuYVn8/DbPe/iD
R+E3D961kvI3iOvhEWa8Y4UPt/Xi2TzH0giYaZs5VCgOvZ6IsXQ55+uSJyENFuMIBF1tYwJjbD6e
Ihanw1o0QB1GyJLq6merFgCeNoPzlSHm2TeNG+UshEGPTumfs4/juhRRBty35IUYytdjFTN04+qv
vCb3ufiaQ83yj89vkcW++4YyuXWCwCVJjQSghQlo0YpK5hNPsJjkbze5U7b3E2qLoDPQK4LSNxk9
TErb/WZNToKy34MdHl6jlk8L0HQtqLAla9LrHZ7+2M+2JsVo/J179mxUZvOIQk2SvC0m+3OILZOc
Sz2fvcJAJBuLfUigqxCY+e9Jz9I9HdsKpTpQStw4Yc/RKjy2YH8CD7++Cx4wo/gEco1sQupAvsNw
cno3AcJxN+5rikEkKPTfip2pr8Qi9Wzx+pkyHjlZ/bwoCjM155c8aKVdUvmUy/+TIRrLSGp4cRgX
cIB5mqvb3kiyTuUqPkzztyYhhNwXpdTzBXgx04L8ht4ed5nPHZ3dSuSHi7YKm7TC7ttLX1P4bwqv
8q4JYoJlw5No/DA6ZuKlkAIAeI0k9qLQC0q307AMc+6ZEziKKAzjcYikrI9GvMrc8ZC0gw8xlvDH
NAw9LAkynfZVUJKs5LxZEHx8wBurQR4IeFAuqeIXXQvffbWsINE2DXqWuWXv5QWKAghaEBaZcqwy
bk32gqGr6a5MxVRxG0bJiU71/IjPzowebQAKh8cmLysDVyhsagwGSsBMSnf/5if3fNDO0/ACVHBD
xcd9UArdCtibTklFBYf+G0/8mFpFsS8cl/ARKvokkC1vzCHHqiLY806ISFmE9tsG+NQ3qGifD0MV
mT60u9+089esQQ0CYt23JXhJdadv4hSIrONo35mKo1Sz5+GcYB/8Wt7rUsrZWaafIQI9efR1fwgE
Meqbs6KPwlHHVHyrwgQaZ1HIT1YQxye/ONDNoLpojDjdhTx7mn4ksymPkQxPCdInGSHFvAW1RnU3
W9g1R4QObd10nZvRAO9dqHdafPQHn5dzsdtT9wmwruX+eDtp94aNBVTPXwvOFzlTbeYmvzj6uAdR
RPC7BqN8gX0BlZjO4FT2Aom1D+/tQKuKaSoEcOOIXCoK0Nw3mH94CUYs59ygsX5JhSOEegS/j1QC
7CahrnNoHYGlcI+EuSJjBh9rJwiKWfF43jp6kRvxDA9zjMuyeuLj9xCvwbC0oLskRe6W5NmN6N6T
1ojdrTU9qYVaTc+LjKphYI8FlPWYkp8TxfTbwd/pn1YzZi1VTB/2EjYOwp5wizcTk6VD54BhEnVb
yOdUgCb1QYQHI4cRECtaXnyddCGBsXq3v9rJoqfTOke2R7lj1/1oBXSCDnH8bLGWzAsxXfhaG/v4
7od77zfag2kUtuqK/FmiLXD8cf5sAL89URsC3Ais35gzl0eMsOgXCM0gk2ycPX/TQeNN1tJCE58v
nW2WU/+KLpjwO3+oc/MAF/dtSVG7Do75GsLqcwuNLQDSizN0+71azxcQ4yG/gdfcIpMQoF8mDx/k
nI7FIcfszxZz1lgi39GtrZN6iFl+HtaNDNt1qA8DSPfzISQP+QCWLB43VfYidAK4aCWRheFWMV2x
RJ/tLxA+MW4Ajm9G7sDZWx7wcwhBBwkMaErP2+7rJw2StskVUKmmfe3tVyPWajT3OUJo95cqkHy3
yTsX9Bv/dXocoM6y65yHwFbbESlarsnH00kLvxqOu5l4RHAzNb/f3zQOhV/PLnoIxS8H9BWims4D
eoyBPbYzx27rMXMWZP2RdCCvs6U1ZK11+vZC9gaSlCAx5hvHodcjDB99b51N0gJ+wIR2zxKhV145
Cwt4UUN5B7UPr2xJoJlUMnI6yGtPsomACsmpBq5pxf1dCqXmCGCf2CAV1lOcCNtSeNhWLq6L2KP2
yn9jYUrIzLAeIpy4LD2ZiNaXo4WwhHWNjJh0yB9GmaU+9FCNzpFZEzs1rpKZeJEbO7P3m6g3BrTU
BZ4ZOO9i+pBb8uyDl1S978nBCadBWAPkxwyLvHKGq8A5hW0nQS9eK68zIr7e2J5DzYb/Quw5NoBP
TQXvD0vRuT6eJni6uAGH4g0S+Z/6oyg8PFFsFP4G7wEKvZYtpLCGiKF2tCzNlefmABdTFIr7IC3e
1/YEfvNPDocczcexEsuIGEgJ73Jt1IyqqeQUJBEfWsrasbAqoLB3ODCthAIhlpLphXmOUuFZGw08
Df9Cpz0NTjbJy4RWPohvZb9XtGuve48muTkZfxgFKZLXdrCBdk9YOYSTXwTxjPhpch6FXY3Hww9s
8z8yVL4dn4EJyAuYpxgeY4lpn0BWx3M4f4lG++5vCzHMM3Yn0OOoeuQrIlyKOAssKIiYZcweHvNE
R+EvvMYsftwwXq/T3xWdotOVI8479I18zOl/3U3OlqT9RImy1lW74ULFkqXXlpck0zJXWkfP9StK
6A1QAhsKSLs7ymCZlDQwtkg1gwboQoQRp+SbKEeTDzdAsyXqsYbTPXnScpXF17VSobAxyJw7BvlI
LbFiuf4E1hzOeUZKGoE1ZmKkC2B3EMALYAg/83n0qFNaU52xqn55AUT8RH/0sQo/HvDbB7g9ZRKE
jCLd5APjt09eO1IW83t1xEfrxH7BrPjcThtT8H8SYBE1cXe6wLGcFejDRH/1rj1RUzdERFOaHt7b
14oiP2Gd8h/BtqsNPdnPAQopP2uBFBFOwjNwOPfD9P5Fg4YxxjJFEHgLFVE+wmDVAMbSSJUZZVY5
b5wU/SU4qis4O/E1d6aVBA7epsC+RGmQCTS/29v33MHLXns4dhmg0e8VRaPgfJxjssB6hwDJmPHg
Yj0MXHOoZ/2zq9zHDvVnyaFneF5xzh60iwmQB+vRYUXzATt9ZR6IR6bjVSAQdSLnIYAAE4Z/XVMR
MFOmNLhnkuPsozWKPeuFhAJ3OXk6G/U/VJwpqBnLotvqBO/NTG46ekTDwrJ4CL0lIREbQJ69XK4Q
uAz3vs9orQm3mjPIdQdCCdhmcCK6m+CVsnSDgw/htE5Hpj7IPLWKP8f8YascXG0jLj2UhueLequB
Kl6y8fwqx9jnYORho7RwVidLMw2GmhzX8vo4zUSU1MoocOQy8eanhdguHThfLTiRZUZv75rOaLac
/VI5D2TBuaLiujwrmeBt1EQ5kVqypY15Y+OOP/CV/ukT6N9+4Mzt4g1hGafqf0n1lqmW4hxzN5hx
8Xsw1Upe/JYwIoB0IVi9wZjgNc61oBbpMD922FgASEs0r8geYzgPEk5Ctt2er6D9PR0nnnjQaHzT
rRZe+TNM+PXJrantWPmEgHAQIN/Tyy/tMwmy8RnF0DzngpFCvi/7d5kQVadpGuTg2vXVOkfX2ysA
cQAcfMxtN1rB3FvarfYQa9Gj1dp+xQ+UnjA+y8Ak7LnYxL9U9FsHgqsV8Ecsgh0WShJQrpyrSqXf
sMsYESXUmXN6bJnggZR8AC1kDxzBfTFbAu9dquZaUeOOJ9cwKrmwRNErPwTxKjupZx90CR/7Kp5e
YOuNfmzjWbbmoR5viPj1x4cG+fWhcY5UWB1LUkIMOS8b3+KrAhB1I+3pHad+x4sQkYdPuS8MTeY0
g6dH8iSzYWCUzsPByNRAKDWA01y/YsayqU//Pprdlx2iDj6MbJp+H5dLLEyjAtGCRLo9XPHstJBi
atg4oz0+PjpYTNWOlL3WTF4yC8BfGM9kejnXKpzjXX/b+kWgMfRqJ+AtYU9ED3JjvNYzDVffW4WF
UjegztPHnjpmEkWaX1cUJH8v0K3rUY+/FT9xCTVe5KSfyZvDTx9Ad0pUm0Eh6muVqCHi3WYC9m4V
aJPijVnXqIYz0LcdGU/ElaTbXZ0Nb38KXVmsk8cOpTSeQaY73Ks5aeL3LRrSPvcpL70OUMpzhjFG
tknwJR1+uDhY+dZBbjtXB0sLxPt1hlQC9FhqGwnyJkHubUQRh7ch0FF06sQDH5FbDSZCRKArw+vR
2oD6uwKWAJBWs8M+Hs3KQuXflsUofeiEbLSfRH/OeGZ//BrvCmYCk8i1swo1IXgrsloum9uS1gVM
mGG8CUcTYorMhTfObzed2bsgSPyBzuisuwcmzuJBTNY8Im9y7/StzBilntZ7haWKRrgNYgQSp0FK
wP1DPI8NUXcAfQQXe/7gKUKXQeJJEP/b/vMNz6bzsIQOHx6rWOp6qWu6MdsG5NpTOi99KTJ9RkcA
wjGHSCeRhh9jFufVd3ROsbX4pkOK+zi5iohv/X3b7Ya4+yxMvF+tJGLQ58OKXU4rW0MjpsfZuxX3
nKMMRxDdQpU+NqK7Bx+Ed5OZ6sIqQ4lvo2u72v9IFn6frblIxPuXRMwI+JEkgd92riT0ytvuWJVj
8MHdJ0Np78/Wl49jlQsj4rOkwMGPMBUxBR6KLaSj+ZzbuoSqTk7SNTD5S97R8A/z8pkYlvZcKN25
mWgxEbXDUxAS6y6BoeUogO2kly6EoNSvzsgD2HBa5q6TJM5DDWMSOMQOgMir+Fn8L9XagsmXSo8v
X6QiiU3dZRzFM1iJ+ktyec8m8B+W2tmNe7OJgGCG3gwDTISZIz06j8ZIRK6c/kDYiYDRhx794I1w
7xvnikVqzf7+hlFGnz0ra6nIt482EN8ejuJ/XS5tZE+w2kDdNdWL/fG/vRC+6meF0+i4wD+RqfIA
4+vsgfyLGPOtCLQSE5UH/3ItD/HOOgqZAVUdC5nXMfiIH+NbDePVHUbLuzKIhA80L6LFa/ofw/bE
uEQg/nDl2r7vTw2QtuZc/xxMH+vwVkXd3BqPUk5DL9LvIQWEl2drgbV0f+7aWa6Dt8FuckePIsdW
T8se+t7rrxwmOPzXIxEe1FSKyLj6JmxVXu9991K6uYAXffdQvbLAjd8vt2Z7PbeLYFgZTELtPgXt
iIh/3IBr1X5OPRrSwFdPNMOsz/alYBxu9nT3r++4/UbGYaVccTkXePfWouTf9oCeiU3okftLhMVj
XGj5x5uHXCGALgGG5peL+P39Ubp3Xo+MQZ/P2RdU7CVTMoxrXylh0iBkjcXaJlIv73dS/rlS9l6P
WLHS0Q1HefRDvYNarIPdN7aXbHXPo6Nil8dGYa+BR6dOaMsbZOaPj5n2+0WF1bSYnusMFPokRJme
n04EkSXAHnidrJQB2DPXyRm4awZvuzOp7fWE+GYjGu7xyFZO6Cjn901XGc6Z0JqA3PsqxcziDstP
XCMQFbzO8qZVOtCWzRMfClGzvJlxTMEK8QNACMLXgInrFdoL5pSMlEenCxwBniFhFaXu6llkCAO+
GLz0wkggm4flXt2k9Iur52fn5MxFhMJ41rNQqd4h+klh2tMaQoT/lEyWqyhNI+5coryzjv/mMDLP
fqo46w+qQAhspLN8CYQkHHiRdqr7CPbcI9PR8Q244ylWMII2ms/XNmZQEhgvUesKd9AIPV3WLLzC
KmpPwv/JEYv/5L0rLZsRL5wu7DvWE44KjVogTu9Igpt6r8Rcbs1xnOUWpbG7j3/t56JwI3aTw4Co
RqbitHaUsVHgXkD6nbfDjMoqsg3v4lFqOtl7rZ6tMf4Jd6M8MoUaDCQIBLoBqbDgoFNoGUSYejS5
0B24vTZGMKR4Lf7SERvN9+aht5gb1fKgaNMff3b5pDLjG2WFtjBCbdXqusFnU4Bm025J/ZQOdFLX
z4/PLlZP8/ADMc/dRWYhNYmXHdboFenWZQ4vC/R84ekkCepgbKO5qI7HLZ540hGVGYSMav2Jt0ZC
JyhgAptUw2gQIbPOhG8fIPt2ankTm4s5XNjEnVl+n0SLkgqpWjyaSAaXfKJ8FP8ELhRkhnhF9dlg
6isQ2lZwtUriSyMGLwmCOvmO0WP9jSsQpd0S9+sts9XwIZTJvyi4VmvWYhc+h0dXBNncgRj9EDn9
tVhO3i1ZF/AWastItXx/XwjQzn8FuSRDKrHlb8J+XQKNyTBWR2i0Qa7ZyudSm8RCz0kTPmu7z+7h
RAb+iQCnWITsnbPnFZEyEoqTl1BdAZbNbMyTLDIGdL2PqDKiXUk/kJv87rVsEmfC9QcBzZwHiqh5
IzlznJUfIRDmLWQRSjGSPaOuGXnCBUuPY17qKroUe5arAGO4f7N3E/L/xTDY6+BdL4Qe146rHRqv
HOdBytnNyHAiwrSSf0+y7+UGqOblXrLRvdHx5CfhBlDJlQNzFLqWeYW9dtE/zVBsctG8nn6yUyfg
KWnenB0ozj2fwCvnhIQt+/nfUq2kZwbKT+PMkldbFWJv3kWrHTgXfA/A58oKwB7Qmf8Hj2WfKZEl
KXJfpVFJxbsajSwuarBlAV6Fyxl59u9en5QWdp/qWt64KtI8dYRXrFKH0LmdVy8Fifpae0KK6FZw
ThetCokZV/ZDdkbb+cQe8HJr0YvlC7WpSlm0De+H9OiFqWyWT7TBUpv2GUIgDawPQq7Zp0OoDvpf
y1aYmD0ii8veBiFGMk/0HT3nwlzPYiNb0PIEuXFfaZnmyOQ6Gbv9tFMnnYzG2ujhr2MoSFnDITb0
Yl2is4pYl0zC3IKkspKdg1pxxWwFC7rMLyf2t5GEr4KYyRH1VL9fGNjxhQJoht5TN2a8Wa3UoNYw
WAIC/GvUv6GACxhj3cSgTQ8abOrdBKx5pAei5r2FW6HqFkcLJuCzjmrtUO4Mnz4PnTEwbfg429pz
/2Nr489JDmqtJpf0Ud9oDWV5NFQmUlCmRa+zVy0VpuTnPsNx1j6Y53oEUAGMtMxaqS889PMFofKt
DZoOViJiRe5umljTBf3kjIH804vF+lprmjMc4p5d7/cbUs+cXTJosfdZNGOQ+uPoDDk7HcqqbsYw
C1hSexqBjtJYqIBlOZJ/uiE5O70fAMM322K1WnnNlG16JRYYuXVifYaoxj/jzWomB/WZsuOxC0E2
oxAZEiWu5W7LlYSd6+dnZwkjz0ThxT7/X/J9aJBYJBaXM3BgLk5yVfXprlEM7v5Qu75mDWWx3Vqh
LX5FPfBFeVid/CYZDGoDJ0pdYwtP4p3fdHHx48GPOSmfu3WARu5LGdojLDSdCc0bYHk0jeO3GTLi
yPDTWDR4ykFqWVuKId47IIDZH1sCU+KX8bkXdbUi1ygd6hyd1xqtuKp3rMB4+uLZSQyz09+Gtyu9
KYxp3wjvwmwZ4XhVNQq66S+NiCwrDQyK1UiKWWR5OAyQJWlaNY0wePzHhTurgos7LtD+xZqRDt7I
7DULX/03inRZ+/oelTwoq6/AVs3LXm9Rj5xoccPNS9B+xaWeY13t5EGCGW1vhPX2RAvmFvyfzMRC
20dPb4TpNCT6EHQcNMetJVGXmPV6MyhjS92GuaMmhj6mPXAYtufwhlNSBSD471A2Kot4MGwCJtim
8ktznx5pt6z6est3Fpw8Dd2vjFpecipTyR++BzQTghLxVgE9+uxdAOkf3B0ACpyu2Htjy1siOCgf
g5N3GBOlezPkVn9pL6pOm0LeM5bOhMI63x8RlqAxPCpbBRZ4gHGFpIudDoQj/UfLoFfeU0fHcENK
PS3n0hNWXvVxsPtV5a0YfVsXxpu94TwB9PH2m2GJomWrOyUpq5i2rwLol2DIeUniiVzV5wdz3y3c
WQXkdFA9NYtW29g1PN21Nh/V7tRxj6+ZIt8xKATYqZFQLwhkluV51H091OkLtRjtBErzSh1Zk2v7
x6t9rhuHboW4zmcR5YAyuYkoBTnGs8IopMRA1yCctnKQJzs1zLGyyT0V0E0LduQnUGre766Ybyub
8F3kuNS4+WriQ0+cMpSqHDfF19AtAbGyqqP7bMkp+3StWVuJxhBfHw4wrxQva6nH4NavQsQClzFv
HNVrzUaHglvSYP+KjO1xFA9UQX0q+9FE5ckyrOjZAV+66jUcOxewtoLDzq5hXpHwe7wOAFOdg+QT
i6GL4VPGs//KiBBrk9ixMwNuT1/vyXTobgSSrNs7RrdsJOgeasMjLynVwIYYS5+gLttivo0mY1Uw
PvQPimmEANcBlJvRlyIqxqRJfvQ2d+cpxt1Ct+v19yE5dh2Gdqh4xhQMTVYg1NWJ8/IYmOq8eWEC
lWPI1G5kxXWlHPsBDKhcI7FfrXEXVebPHws6iOXtdJxu3neTPlQLSwIPaqyo9np/TL4dN+FCWaLE
LWRSXySG3UUXC1ZtoGjOovSYlTn3R1lo1HwK3Tm/oIoeu/x2rgUJlLlNBOKAXIp97bKMmnk84dYq
AHnAC56NK1phSTdG8JHP6UvalxEoZ3CHMtH1LaBRov3Xwhr//p33NH6mYDYnkhNuSsQv7HR1Kein
m8Ff00KJp1yz6BJbnI3Wr0iXdrbtjLdVcpPAvMoxFvWOP5nAgpbsWYs3UTedkYrgWJl1ZorHfouJ
gAsCHK1jvRzUh9OO+8FTvr+DJLZ3MdENd/rS5StPJAbynkPSeq9WeiDHm2p/eAiy00PanIb4YWHY
6T5IBVHPiL3ncOBX3mrq4KXKhnn1+NeEnDhUqlsxmvB/C/gBwjgRndnavz0De2hDMR0BGQyHxsu+
oYGIqHSX/aQOcEAOlYdSCTXj/J0Mk2/ugwNwtCGSOmgHGLSqh3z46g8IVprgS9eW/f6L9tPIT/tq
gnzKdbO4ZNeDuCjoAJ9uuXKY4tsKlWWQHRO1d3cXh9NrHribXU3aNe7MpIPnekdL9wsiH2W5V23J
lG1wh2rtWbZGXAxXmMpjLrafgWJ7SeqGyUCJNfDycJ0FesNNcizbilrLxHKnjSiCxbnjKwHQHwnX
TAYREuEYIce6lXQEsY5YO9UzlGLoLdRHWwiBgcfgjYOPSvzsd6J0f3twxhxvcUR0RejJvfEvi3wl
SlVy3RQTkOcnC+qCDFQQX8RyFdTO46wlckNPAJNvLq4Rz3oMgpVklGXiproiHhM7QQUUPOh8JS0w
NGHkiL2b+Qy43kyMne+kxtSNLxE/ouiAZhbCcArjut94WRoplYpVNjFnB8KKVsndYDQ1z8RkIiOL
nhXffaGbhU0TLjPLgVFdgM1PN4o1DuuuRLI6ue9Nh9Ku2LuFdCgGVPNOBWFHTyq0uel6VfiuD0yL
gOycL7jwSQ8cdssm/bq9UEgx19kwYmoUjjO2/c4oDlekGb2Hy/zj6tozoOvZQTBeu7VYTWuaU0EP
4Y0OzNSIyPMwQN+NImRoF4cmnDKT5OKCbQApnPkOSh/dur/HUyukx6H2INSguG/XFr2hiZ0nFOH/
YULauw81itoAqI5FPtsrYhoqMX/0X4o3vKft97Qx/IQAXBZ+uHOZBls8+PY+mGzFo/AWW803FxsT
shesrxeCtMNpss7wVW5K/ZeV2kLFNefgS6NGkOy6cSZwL4Ra1GDcZvPOyQS9oYce7OF4ANp0SFJX
xySQmSj+TuZZtD3TOf8/fmllvedqT388g01YEt3H9gEoG5Q1ZubKYN5i01e9JjQ0cOMUuLQIzgdZ
rZ74n3w35y8gAFOHWr3S2/q9P4PvZjAEcVZejtSrCJCMIFhhihH8jHXpMrYzW1RjQDkrH/Jv58Rl
0KlMocI+qySGD3bJeKXeoM3WcgNMt6OOe7aC/WcfaCzVqhPDixANFCnnkQOdHycwt7VkAJC2BtxU
RJjs7EWSnhHJgKP6CU8wRUEsPJfUoM4mbapwfyOeGpK9jK8J6lLuo/q2iraocD4VztbCgixes9x+
lkLUWAPRXGN3AfiEeavFF5c680hXZJMb28Qsq7+DaUseVmBHpFHPB1SwhZfmDz6OMBXk2Hwtww4C
7Z1pSxhshhD4OeBKDvaD0nCu87QHz68JY/AnSiYlzJ8pBmqSAmRvqo4qHP0sNIX4uKItN8sFUy4S
hhsk6p0ARFwvNDj8naaC7ePN2f0vgEjMJInm7fTFSFHM9M43o/orhPXmgQqmo2r2ZhgmZIZNtOZm
TMj6dwTVcXy8Asifq8kQGqT4IC6ETz3WuHo6wclZG5cnaLQKzyLy7rBc3U+2wMGY8QQyAQX71wex
cawvToIK8EBX7TA9S4Y9fUVsbYG3kd1U6RAj9rplFhzh28oLrRA2xdUMF0YpW/8iQ6do+6q6zNgr
9FMDmcl7ML3VO1Fr4zRvFQqZ3Djp+Pt2YYxJ3EaTqvj1iuMv59G9zdC2pJJ/I5wUJwWknfvlCZ5p
EZKps6GIyt8mtmQSSNVAb/bMV6U3Tvgn2o5V4qhlTKRJIbsrIC3C9j4HsD2S23RGF56n6Oxt1qxo
Ku2IVvo7J2WpzFAhcqQw34Lc/9wdk1BtlYaLXWM9oZHAnTzZvjLN8i47J/DIG+h7wFWKiMsYfrt1
OvHYM/6HS0X/q0p9Oop7pZ4+8rTBjw9ZIJ3Fv/IWM05a6isQJs/g7H8D4084oxstL6ZcgRW0Dafw
OJt8mXWen3nmhg2gOID6h8TZ4iLMZj3x8yqlLf5clu4SYUPL3L2Y9HefzG1Onk9HkQwScuvNeXQ+
CJGDfLq4v36TC2QqKMQc6iXSYCrVmBa6O1MzJjEn8OnfttFfg2UuR3XvjfdT7sX6Jy02I2gl21y/
zPFj+kY1RKg83Tad3Fr8M9M7fYcOt7AleNxvxHr5BE1hrUz1wc2/fje2dJr3gF8N+dCKfg9bmkm3
RfiG2ix+VmFwBK1UrFPmXVWYFFMq0lgCxv/wsXPteSJT4i0e7WSsiy3llucmf56hjFfg8/pjMFBn
1zM2N9le+Z9H9Df6fPDU+7MOHUHsNpF/Kqb7aMvhz0fKx8uhBgpw4nneFMOOytAIiiO/b5xStk2h
0zgtgfNvNkLmXzQtEkTP5tjUebHo5xUFfnpZwKlt9nxmrIu+3aQK8BUdSgWbVXVeFmNneoB9YMum
8Yz8hhc++0aoKPGGDYW84HjnmyfLA6k6vVaUbvIkYIFGOBxP5LwSMBII7qy3s2jXS+NRGhDMVgQV
QN5hneQrJL9oO0alyPOgOu1ejGy6ginupbe8n+1hruz8fJMly2Qi2h9YTR0kcFJrMrfiVyR36Yq8
tAg3QTLgV4ryWwfrlSP7YYscksfOrqGTY4wH82neafC2B1w61X6BXvx5AvCKI56ADh+Qv8/0bpuk
MHmBOwcTvV7e59wtszhyF/rQgmShWKLZxBrQ61FzTX06lJkdom5qMzd9BAn+VYlQE3heGZVi8+bN
jxEnuEvgd01YJjS6Pa9P3++YdcH27ciAPmrRdexQh/4Xh2moajTwgTehh2o6PGof81Y6rbwbtc75
YaWFB18DNYC55rlsmlo4bgkJzugZkBSwRePAYOF/2EykdyXaSqJxXbb6nesUwn1GugMPMfLktgAt
u2HvXvjfR5gvf4ualM05exsdbilLRXQ89DKVrANJcRUPnAMQ8HEUMQJ2aFIrpyq44Zg9T/rWCBWS
rYwLq9KoKBCIRP4GpvVKRMs6olBbytHHgBhEaNI+lMSvUHdm/wxARJUO28VcY/7dWSFjDLK0znEn
FxCEpq90Dm0fy33mneOyGbCRoDCXBLQ3yBVg8Oa09oTqnOObtxDyQ6HJSsQJbjP32lxTrzcnNN8I
TXYkzrNxGhnHWh3GNQ6A4bbErd5lHY2TzbYLuFTPoh9/AZbCkX1xeDIOdpyj/VwxwlkeiupPlIxR
uCLWm2diMr64uFXrHpYGCwvhkxXd9XtyYcs14phNv9b4zFJfhE/ZKez7FR40v5ONq5JRMZ0+rPCT
xz/plLHVG08X4BkLKa/OaMtR/oHb7h/gK4wtG0rmtGg1YzvwtFaSNBg0Fsv/mFodmPkARAiFiM4r
Q3nJWWjJP6Xg/1jdMAOn1DHozeTHBBSaDS15/IPmBDy3OGpJP6jkgu1GF3+mvB4b9NP8IqUxIIJ9
ig0QWIfrQxLFqsAT4MJOdGaSgS8Sbp3a4ckJwtTiPNiRC2vCoeMYY3wkh1E4JQGKobt162UHtNGT
UZv6oGXcuJrp2+OaqeZQB3pVLmnFNCNJnIhk+dKJJfgr7eeARynTNTv++stBCO5eSO/HmyMDCT/R
+UmtL/wHblnvYumS0dw+mwk86DcBivvcMAVR7IrnPFXxb53YV91kwWuy7tsJcKf+Cbrcan5iqy1X
JBYaRuPi5KJnzZeR0bq2Qp9bFu3157kS60fpDHvEq8wB12jSIMm3+vz09s8wWkf9z7Vx4tnIjvUt
9u2nZ5ZC33MttRLqApgmnsDNLNDZK5C32DzpZ5tiOhn/u3RR2//bIn4tDH15BAxSt7m73kvwr/9k
vuMSiX7VdDD3yRmoHC/HA+SH0CJjRrxEK/4kyyGIYJr1+mapXNOJ7N4fWdWqTxsAPTnoPH4b1+e0
T6eTj8GBg8ocwgcRB8+k8wxzH8yGtRUQpCG9UDwRSGA2g9+YJIrdcrLnAGx5LGAIdl0WB8d7g+cN
6reQPEXDd24FfN7gqF8lLicc3U8QsAjacOMNP+YyLqAiOrJ/x7G6p6LqfZ6Eg3hOxtXqb+s/2+gW
PTYj5SMTz99xymzAR8slugWHzO24qOt/B8wpsEVXuCH+yFYAebrPFnZrWQKbtO1N3QOtnIFG3pG8
dpUKPOgChXnDLCoOeA3yaJW1XH/ylHJCH49eR0H/vZxsBG5+gSuXUOD7EMmltJ2CcLqoMt680NhZ
P8bkZy6ZcDyzGlM+ouqBXAu9GCCD9cO5l8YM1MmySs/gEhfbHa2CM4GUTh+A3pTmNp0+6FDpVnv/
uj8tCnBgN5eDuUZGtcHcYvN1kPa31SlfdLxrzgdkZOc0DMed0pI9Z3ix1zLYKdag1pMG+FNZPChF
kHBjYQDkmkvP20nA5mI00hnkBjGwWBoy9NgCicDg6dOvLXOhXy/YEmWND7Nx3aRKKSSI9Ap7tVJc
Pk54UorNk4SApkYaV8ku6xfpvKzjWXvbrm8MueAYfO37KMyl+iStL9cgKuglDeBEimTtHptL9ig8
n6nKL71LE4wgHeVcjjmlN2VTlYSilB5B9Y6xR5Sik1qWxpqX/v9vv+mDnrvS4xCkevk2T2vhO2FI
8q1MObDlLtzcocmCxdpYPeJ0OXm2G/+9LjCb0rKe8S3V4KJEMTN6B2+i7iUQSpA1GrmiIEGYgSBf
GJnB484EZsOBJ1OxpwvOlZWeyW5uxvpqkcCb5JG8oPUxA60raJRJYs4/YRT8oH+zeTCjK4J7Se/l
i26mFSoQRYYd9zBntDQ6WmyU/FfqO0TW/2ZVMRO5dhixGAjY3i9eLtDbiIpT5c0nlyYJvpGXgy4H
gLEMCAFov80AHxP/V5SRdan14Tvu5hKfnTwOjYSKTvPdUltXg5NtFE2BUuwgGkgJ14P8YRCfRgva
uJRjTpXtFsdAc4D4gH9SHFiATv+gVLBtmQzt/D+A7uPXVFVmA6MWwEZX2ZHjQ9TdRBj2jNk8fzto
9ZAzDzOyaP9BibAUVvg+sgNC6oiQDlV/oJdSJoVA2vYjO+AnWZ8+W9kDid/i29Zf28AtqxQURNCl
hadmRQAQKNeG/Nc+asigWxEq2m/m/d3oQ3K58IUdz0YtVuecskRS5eYDi/aY3PQeAVZa6pG/vcux
Jc5yCyscM66+48nGqjw+BUfXlXrD5nMp0dhEJBmqsZyL7SpomNRTO6+7oex2qrBCyxihEugJajnU
LittoXM1M+BNvefdz5io4cFBqj+W+7c8xy4qWYXolXbJS2c1oBLa53rcTxnZVlt/BJxq702/Lufi
6mQoG6g9VGlBYLGdg69OvlotqZR3BvwzNasQTSzanafbexgVFcf4gj7zeYmNAyduBw9G2vHxK5Au
Vd9mLCCqNJOM0x19SUnnfXJSOy5ztnM9h+ugr/OBOEis0/W/9EYV65FQcRqZ2SKhilv3h/jmAIjU
uSVFaxq/pIXdwTGUI7InrOI28xP/i488flrJPOZHUY1/7SFZnn5JqWTIAHLhOwAE8BwWnZ2P7bA8
nFHSxoxEP/OQvr+RkoTvQ+4vQpss4pG9Dm3Sqrp8K9zZxomCdKyvG83c9s4A2bH1/XXuIWj4QHXT
b2qlmcnuy3RlhqMrNpnrJzfs/exstGzkPtp/i7Cu9lNsYeMBWUyuO0t/ncF5gW2NYwE614hyWEjG
mcVdDl0yiKwBWVwrSQxCxDwWWVksj3PQHjL7A3QJcE3NHq23SOrWgs22yR2gNeq80GoWjX/z6te9
9d1y2mZxZDV1KO8V/t9FjMb20aQeOFnTU9rdzDiChh9p952BPS+KirS23EbRBw/H44jewxgDVXYY
kwarOk3mRczVOIGByzNFyjxNjWNgVlI/XXf3jepo4oIstD1RO9PH7F9O5yfWLb83FA7z/jo3nB01
pEofP5jZ+Tnwr2n71tVEec9hUSEVLKxtYhmwBTRUyla2qQPnmc2J22AQGB7MSAkkY0Xvl92yN4Jz
gMm2HyiEqtzizNlvA39DD4prLa/EGeBjSpKR0Iaya6X0fQgsz9RRtzaLVDfZiXpBoPQVe9PBF/I7
24wCEx3QbW9mmojasi/y0kFCdpzNJuciBlErk/2fBCImcPZbFjmA6NEtJtwYNbU5zLenj0mdoP5k
M4J3ihDAynNWH86oQ14RIT/TtSTJkBrAxlt12qADoa8Ee37htrsQvR3nRjExb92FGuaz/86lai95
yUH32PHZ8JKaXWgKy2UUn0W+N/rRwt3PoikHYeLksgZ84IsFrQcg3RmQopgHtxrNbuMD8F9+pPO3
1E0QSbTp9mmHeuB9M3aGv/x+CD2SxatWq1/J01WRcm1E+MqzGaVWjjKpbm6XLrt0QtFbMbk1mgqJ
s5rx3jLyRC2fGxXtTGg6Ff2c8/SxsYxF5XpPVzPTh5KmFCucKyrakdOqb2urrKavzwOiU1BHZotd
wfeXss/8Y5a1K12oQ6MRMGbqMu8ETfqCaEClubbsNo4osrnYm/aHGqgLqFJiGvKBzK7K/QVehEuQ
nMdFC3v2G8EDfjD2uDWjlDJ//qol65zzgK8xplSBM6Y9VsfisT3avoKJ9o9y3BBcQG69jMZdUB43
LYzP4jvm47DsfJsklEWGog0X4CvNGb3HJDjDbzpDew7eJfQCopg9u1BLRT4S0rNVVIDXaWacEWRf
yo0B9cbe8nrtb7z2K1+OYmito6uzbxyP1ihrEMr37pReStqJHZZJ//hmqKjkHqn4uspV8reU3/d7
VIf5+eCeXDb16tjNQXuwg6jVNtXLNbxgLNg2ds8Zj8D1EgxuCTGM1IiuLgTdOYavaCd0IQTnFcR1
nKekVCLkhj2b6d6EU2px05ojwqxRJmmK3yUacE/iL+06Po2AfVwBoiTmR6xkYbEZEaiF4E8LDUjq
BybrRqnvhjTquAm7I9dyYZBDlB516xEaWIccopxOEuD6aHAuq4byLuDDYYf42Elat1uf+r0rpQLw
h/VW31n4jMN7eyrMR/cwTzxugGtQu5cPx+d9Ogx/DdEkDUReKHFf255bi9d8mPD1aGYuedA+jW6E
E5sboWdrJeLs+xjYQ6Kej0vAAu+W5rR5JDchRIc9HJMXCx0EO+wpjstVxO1RF8ij3Vawj/JgkW9U
lszYLbLxIU4XncoWS21ElFBBDF2B7Xaf26DI+Y3LW6v28LRXrx6jYeeCP/JEXBRfP3JgJOa6ktQL
PGxmGivtt6VE1W/ELjXiW8izA9nTZ/O7+TLZEeAiOq+VLuNo6DnvhTKUhmj//ZsrxzEKP55RtE80
N+V8ox2TlQKLdZR7kHGPve10vDeBAOmQicXEM6flnIFhm4AS0MFJnJR3WVmR3hJTdD93m+Iv2rUO
xAPcYN7PVsEHhXnkZvfqHXbKWMicCWFauo55HO8AoFJNGk7UwFuiP52W13me/7TSB1xaYP22wdy9
MUmPYgJ3G303R79jqlFEZoobwHccIQiF1HwaXGWcT1FTyc3aF+55vIRyFtQM4kKgOEjyOGMSUu3v
12kqOaxwPzmpm3SIqPtNaZ6ewCYlGF7Cypvzz0eeN4y3BI4s9DwcV2fdulScNUCzFClWlKW7uHAj
qXyq7UnygsAKB2Maf0lAg8W6Y8nCLwosoA57orl0WAcBjoNFT66863WKEFi3Y6mpAE48n/jz9dn4
2AkzlGaORe5IVvxcnPyWDw/4fowjv7g7sQHdmWrLc0XBFnqOAAQPDxDsHmw5oPZFxW0+C2x9y9pz
WHJP9rZZAlcNyVgFsPxUTUgpK2btnVGU+yz17o/IxTTD5nTQCRhjoU+v+pkGkt/4R4P2oempeAVJ
B/vSvvTkq+XqbcsSSphrEpLrJvZ2PvfgUCEyzF76zeYWtTK8SV3g0UefZCF4pC0DyApHq/zhr5Db
wwgkvjJeT+2DT4rmS4idEE6kjeEzNDtJAEMKrHeAUOfrRRM7zuuz/30VRSUQK6uoKogObZHOVcST
12h3SnHuGXqiemWoheFro4JsRyv1UomHgaDFSw/TtLaHYI4RQkPmfz036UmOmug6Dm011HUynbdk
ozCAJ3kl8puCXTKerQM06sYjhIed/3grs6bYtO8ly5GM/xjc9CEANgvrT7GZ7uXcTIy72juqmdp9
RlXaWpq82vySX7kAsjfNAWAzcp21HlLiDNrXRxY6JUo7S6ZXmh8b/iyTRqtO6kF2bHQ11kTuPERI
ve4CwPqZwu0BLFl8GB6nk1tUnlY5wDl+lcc5RZ9HOov64e5b5AMJEIRKjzL/+3YtydKbL56Lp1ji
7S4HWhcBwyKn5ITWmTMO98URjOysPdN8d5eyMbEqhL0DXqrwl2S0KZBQ/atTOmFknwrmuUT1D0ns
EoicxhmGYzpgaApzOjDwx6FhFLDCkEcq+IUP8imoPPrvGANw4EIm/5FWRYNYbT2d0YKjMCdWFmzZ
i3zL1RYKLQeJ/H8WhIWBfG4aYwVr78LQ1FEEPTp3IXzyB5Nvr/L7lNX0DCpWvaeuz32I7VFluXmJ
b04Is6ltLBMZOcmaNKOFR7svgcb19/Ep4lc83k2wCQgTL1Yb248Ml7hXvxbtxfddZASXHcU2npvs
s2zhlyiOuVNuj/SF3a+vhZitsazAuA8Ir0uwUnozvy9BntxzUHua22zjmvTpEwCopCLikQYi8Gv7
bKyZrvXKysHAeA3g79Bgtc954OhZC1e60dooOi/mU+9dsj80SuA1F5Jmv7Im5EG1HGvIIcOMsQxO
ezVdAz7q6jenzWaS2dunaK+NLK+AQ6tj8RbbC8x3F76Y4ufRdous1z4uWFHEGvs7ErCqf5AojMAe
lo0gHuhOc6sZTNlwbOb1G7B8G/aNPdES4uFvfFNqEPZZXfBRTcY1ejMDrivbdDLXZyxOU/fBfnij
P0JhJEYUeBTJ5PpIGgutpzoW1ckF06HjkFbLcz82ti3gD5X0D39OZIBDrjOi/qyF1oGL2IHxwGVY
P1S96B83jQDrFO0g2lNFg8c04PJDB1KnovdDMh5q6kXu8eL39cIwIcaL39Md1XOmY5JZNjTIT1Qc
PAJOJi4b1hMJJL5ED6weKOaQOmOqSlww8Rl3+OU9BrQF0X4dLzQTDvHZK7TR/qu6ax0ttrIqpW/L
pBokFiDQD3N2LlsUqYd0G9fBCfZNbLoNtYcFSeeUa8L05EFNgJ8lZO9FMJoA9Zz0Q58OpejVd++g
bwZT62PP9BCRySM7mm7/6x5FocbBk09g+VNDMSibm7MECatgVZFX8CwqWOjfp/G7MrxSPIFsvf26
8CMmE0FZv2EtDaIM4AkbiMLitTmee1fRvxUjHvJ0irO+X44oBukXuNiy1BKd2e9WH0ky2xttDNnN
KifA8hJh1gyHJmOMR/54bDCMMGVDWQ9YdUtoLOoWU/2cPbMfHblPYN2FI17qfezXPToj9Kr3l+e4
nk0nB9/RA2QVJDMU0poWTJ5gHQGlxjtMiTYR/f3rgOMBK6Fpo83aMsnAm0UbizRXChqQbJrSYkDg
eArtIEbVXs7OpcWgaxQjI8DTeI7jeUwCE55S7EXUw4Da4SfcWcB7ZrXrB9Xbz38zz+e7XpnIA4mo
GBCiykeR2P5zOHDty4RUjhk0mgHNN10QarDkJOa7G53QF4jWp365qng5ShMVVwMwxSFsYNHo8cf2
bMOcWDb7KEVZQiHbe+jdZOu4iFdZ+mPP1WIOU/v9uYtAxmk/9ivC53a+fYPncPabM1LKa9iRzsQD
/9WQm7P6GvkmqDKZmG5L1wqVJIiRi09lKqIquI3lLTGzuWk2/xCjVKJ7pP9sbU3IiAaK2zcGpEcB
q55iz1FnaItqPtgG7oFT+fBVM+P6IMdgjB1yDYjX0vFGJlo39JwlupJqdAVb9RlAUGB1pk9I/Afq
joXmG2oiw9hkbtwALODxXeAr0uLbS76xNgVX5SxgjTeJ9Z6fJqFJYbqYjfGw/kbebpQNA56I4x5y
PGF+7BF+q4kpkdsyRGoCQaegVwIb8pzA2P0dqJGAwLoaSRbRc/6bgMII8H5lD/Y3F2/RYvdHf+Ig
0qKA7d9j+JgRg7Bem3UlhV/vmYy+KTsoB2jQiEBF/ZutYhRImQShUm0Vam4nlT90AELVdlh9sC8h
7NrQckt1fPCaZjjiHuiLBMPpYMGzZAolEW7asZMVDXhEWiIHNQYEORy9hV6CKQmFW7uN1reG7Ct/
PDHdEDzV2jMie7ZpoS6bWiqUyyVkAzPD53LRePBY/b9V4kWtXE0JFVirstirZy7C9x18F8POvx99
KrGq57PP9dVuPZmJggCsOWYdrfqOhA2ca2LEoUaFHLh9spFftVagLkuPYJGYuourlb5In7kgp88I
zBjQoRUIBQEL13HaCs6vR/eVwqujxduG53NX5laG7floTUQ+t0BEhyqVq7f99QhAtSA5zCVt+Y+b
x0GvrArTQ01kZKkEUDOzTk5lOyNgQ/70GluGjIQvjUmCC1SXQjDKAlZZn5wQZw7W/h9Gv0Oz38QZ
Xp28IFcn/WxMWte3zz4zsU/sHJORI4nFFqUJieR2HoSzBn/PmsPw1edsSjovNG1DYpD8jiMEI2eR
0TBrVA7r44nXfQL3LUHz3kvz8HRU6Sh5my1pXmq+Bf7BvnD5+u3XbjozRmQynOhc6ifb0x607P45
tuH196nByTAhj6nP+Qijw8C+xBVpjzMc/AknI4hsYuXrMPTjRR0WcFE3j3lK1fIhOLstyrSuUnqw
18QiZgy/zX60OHajRHGsjZcdSSDAzNuWnMdjTnpdfjVnooybVsdRXYmO2suOo2FkyjE2OTy9FHkR
wo2nAhCu4ucLMf1C9yaHS37KVVCRQPnlG9ohl8Ts8sw+ME8S/5tK7P1aM0guuVOx4gtJzANnBtdZ
4fY2l/YeuwbyWE1+Ue1WhhP9AghM3h8U3nIy9+vxpHcM72OlwxetEfVTjIBMH7xUsjsSowxgvwU2
Et5lqjopjTTujolH4hU+MPo5Wul8cbR5ChmBl6m11kFPI0kHWibD4UYvHPr8i7hA8AzOLKlg8BUh
pCvp4IW6NwQLY9AoXrfCzXQhRgerIM8jMPlp2mwFH1i3AiMPq62HiiAtwYo25a0+uUCh/OLUxrvG
72DlUuJMkNw+KeMaC6jsV7raGA5t8HrEvE6JI1Kh3e4HNUDP5HKw0u6yo35LaKL5MlhKUSRlj1Vr
kQ/m8qpnGvFNWWGBUiohq17lgOQdRMMqsWX62cEtZzVAfbG1frj/zgZvH/EQCiJVjeFFO/axcQkT
lVwYRkyHYNmvmwuF3AVMc2NNessIy5jjR/lyNfjMeYhd/SVjwsNzAC6jMZIMXlbMUmQYLc3on4K6
4xa4sA3WGF66BODcFgT2kmk9RkDrrAoasraRzGwng2DU7B94vxVqmsl1bl6DiAXezZ6DZJLeCiGc
xLSpTRQ/INHlb94qybqx3W++jq8ZKt7GVrNulfA96QkdzDmtLemjysilY2xDfpa6Xz2uShy0OPCr
FQx8CkUwVlaTx2d2oiI1FNoPeaaJmND1a872lNckeHppOvHQHem0r7hfFBWLpWfrM8mSABTXCjag
/zah0a+rFaovcBjGBZ1oaUIcCWPZt2VOexWFCjt+HDbkafIX6VA/PpIZiN45fSwIntOnHaEDKT8x
BU8mZYrPjUVaw/dgcrMkyCH0Xbmxz/VQTDVd0LF3EJ8IPtlIkHGHr4rsyNOIXIerUUZV8Q5kRDfN
YkARUBXW4Ez/R+JSCsg31I73gp0GNPlTWnJKSETSjmi5L0+d+uZ2NFfsvx6U9bHBKJ1kL2QlFcmR
SA1SsFkUkzpx9lWpx6K+djawBvhqAS9WxXSo43LnvGno8ROKkfNaUHaznsozi5zJ3Jzy6vhRubJ0
Bdparev9Qk21DzCrT74ndNoDyMG/+74+i6290xOomoP5KU4WTTTjsylUFNz7YB/7YNuXuqvZBn6u
I3ioGRiQSWESl6Ule2T1F3vVFG5Ml4pMTUERhS2Dw/UjYBefSDTr5Vy9f46JlDYyw9tFJ6LlsImc
2z3LPknYhFQ41weynh6vJXR/VI02sI6YVOWFdmpEVvB0TFWV2a1/ldqzclpEx8YaT2v6igIffAfw
at99utvyHaYofbvK7T/XWDbh30XDvWpzeaSokgZn2gOgA/u/AIPjMx8zv4KoRZtEJ5NHkUVIazon
Ueii4by4qh9Ll5Yxk5bZg1g/nixnQ/lM1hnxd2cFK7Dc+iSiSL/XOYWo1a9hzQrMm86YhKmxVWmq
Z62b9YsVmAfqXaG0BAmOZn8KCWJTbmTdPS0CafKCmfhZCKj6j94UjYWSO3h/ospGbPbfUNISrjUB
GpYW0gnZY7jJLfx50i7N5OCGet/Z3SHiv62+qHG3MvzbZvBbEa8iLIavNCLZiFj2/kQNoVrMdMGv
LlBBFT5dYjuo1b4IFvluRQ55P/B7zEKd8tb7K/xo4hwScCBBirP7iNboDW9e9yP7tX/GlgN1wckK
zUbGksTVqeHt+vCGR8+YtTAVrJwluI6ycp1gujmcrjeZrWFXrtWHSpi8lss6moOwFn2czAiekgY2
fFQFA2/xCKQyS0S0xMOtCVNdCu9PSi4lEdlXp4l7E5JywMb/kzT1rkReWg+FCIipSybb2NrKNwbD
HPae81LBWzHwCo0CfValJtqgJZ/5GTtgkXxAoIk+9bcEcg48Ui+HZL1X4UXmDOWQpQBCO+Q40yNR
vFFKcR33xc2IQgj+yNjb5sy57D+ruQ7lsTUIJxZe3RYS7mMw31CJdGUFZlKxXcHmKmgWmTrclfhv
D+3bvV5JtiUE8ykL57OGycK45DPuER9VS7/qK/GZ0fLy2OaDTIAz8KBWh6EBKQ3JIHbJTVbrW2s1
45IG0RXGoWIA6umlFV8WG7rIJeRoHR4y/GABwJnAoqZBIk691hFNcdP0+7nLSI/txZrzeBuEzRRR
0M6N2Ug72+W51TqzCS2WeXIZN1xQ+iCNeglqBFtJd5nCh6vD3YTIixHcV9gdmg/w7kmMhz7wI5Rj
uWeuYqBHXpRVk0DUEFqX+iPhVh7sIodB/8kXgoBlbDscSohU9wT+AuLjjab4pVac0xtXVZTvU37r
F1oNgr57H17Ypj+A/E5VZ4T0nRNFpe9gqaNPAQVxHNDb162pPzUOz+9sgqAeKicbs9lvPrWK5jNu
NJJmTwnPPd5QQZxz3dn8q1/ow/FXN59VpjI5J91721T2D5fu0cx9tSVDwEZFhgWpCkBwcuZmf7qX
jgtgeKzGXfTNRUcZ1Fk76NeMp0T+LvE1FaQGX7hI5HIOzkr8RsEsLuKl6gxyq8G/XoFRGquLoEq/
7s9Mn3xJbfDtwvqRfPfvtHIA5HD2TffSnONErwfXkI0B/8S8XJRbWsQB5EkkjmuZsQaaLHpbFaip
C5XXXv4/7VGfGleM5nJwLvTz3dFpDHuuz9GAs6VAEBE056kKKjvaJ3N+C68caA4PZZjL0vAy/+R6
GCsUk1r2QyFBDInw7OJTHodDWBYqmeFLhsKEWovQrNjhgNvLgEd5hNfvw5VyZvUZgltsSHah3wxx
DaWMsOG05Vw0vbXwzwZ1KGusEypMMWQJmGSbLrqCPLO6IqIzY+53e9IlrIq4cGiUGo9AnqEhxn4N
Xd/UVyBomK7cZeEHEtsb9W0t3VaFbB0Jt85F5c7gt4GfIJgg04jBq/JxVIjIOBPYA5dKsJCHeyJd
t/1Dz0uWd1YdOweDI+y53Z52DDSKMQVTqGOXz3QquaDB54IT5kMcTjwQ8VwSGdo4UYgoyNkJC6lC
l1wZknJ00lbUC0ZhJ8nfBHK4gBz9Teerfr58oqqygrObTCBJkcimXThBC61X/DYbjJeNaPTV+RjW
Lag0Qa7t+7EuEvBvCkcyXC/LgH4P94rOxqD+tqstNM5c3UxS2s9GzFLhI2QnLCFBZyrE6ynqIV7b
jJyVgc0bkrMGRS5hO74h6nihMgNP2i7xNOLkBSHcm7POUqK6yMz62mX6LCbcdBA+g2bV//qwYdRt
fJv4Q9BlC2BY2DlRLfMYBE4/FyHUHLhsI2yQAOZZP1eHmjjbVF3mcCeQqJ1ImTuVPcx91O8GSeEA
A6MzNPEw1Mdb/vG97NSziHMo0HgBgL7KDZQ0pkbC1tq2vxDmdMUaqFzYDVJpSQSIvtUVLuw2ckQ4
REi3S/Y+XVlnDIJCYro9bMFjNx3IYCU/hhTIVIVReKVYWajxhN4nP/tz9hCpD8WC2LlIUvu1Q6bs
nxFYRJW7ScPhd57akPs9LswJF3nRUUG8971I4t6yp68CQib4juYJiLlNEd/+aWZpDmDH9nEgAQsV
4RlV4jDdppl2k3AyIoH6UNRzqao0NTPCs0QksxS7LITF3cAeT/U7DmX1Uic1VckB8j7Ni1OHMUD/
U6edlZcOxLlpTuqpqJ9ssqPHDII2VF6sPeyIy0t4QO9qAUh0T5vlFjk8g+1sGezI56F+9V1bXgt6
mGls1vsp0XzeNm/Qv+6HHqmFfjytSVDj/jow9EkGf8ICrO7tedQnhz6vfNFkXhoL/W5M2SnrtKDL
gQtdyXvd9bz2OLyRFG3nJ0E7PybIGq/O3korgS7Yv1XynlceD9f/4GYUT+otNeBaxUxRqu02scYd
XAUto/7NNj90SDsqFODvGYkujFq2Yhmwn+thH/Mx6amzjzbwl4goPFuISNRjhjYnNIKfCvnYLsxT
P9T2/z9U6/Ks4PjFY4fs2uyyEZU+henMBS9f2ZxFr/1rHLNwzLb0Sxp9uPYZUUUUVwH13HCbwW44
RXOa2sD42OF4XYTFx5H3Uyi8ogeOJygxCiO9YhQtMpRaavN135ngypzmuowQcbZZqgO+KTTrDBCj
u+KUoV1s8dCFpQ+yqH0hgK9rNW3VFHkF0hTXhcsbLoQlOhpEHWIU1gBeokAVDWzXJJGFYYLccCAT
Hu8edA3zAz6Zc5zEiAMctDPTrnObEKil6xnJeqBsyHpFEilo6+Ac3BgndMrVcoHg7EikWDDO4ypr
eCw2v+OMES1W2LrEYmpPS52lSkAX9e89ehoDB2okb1RbNyTfyKN1iwCFXpjUWBtvxuLsR0DJcEDC
KdPMpXN8W5f6lrVGhyKUPpGWGXUoldYYmtq7VSDwYWCVck8CB/OxJzQaHNbzwfHnN5f+v8jRMJyl
ARQ5MWg34ham7oigJMUVtddBHTJTGUC4pSI/bZwlK0LvDBgq9dr8MjF5rxW+VjMmVXzjbW7ujmAb
YfN6WfqOMsNFWpSY5xhjYWk9vi31/hcMCm1TXghmG6AF9f+cXP4iAQt5OGCYxad+6udckRgoepkg
LeQjUoCR5JXSk4NaFnmn48eaU7VYCR1Ytihs5SA95BaiofablswLLr4ABbR6XDfeSe/gnxPIYibC
3Gq4K3osO0xS8qF49FcCU6ULQVH1RL25PntvOxQCLslOscUP+RifcMktJYa78cziSCBpyhXnU4XZ
vWeBs3p2nL578rLFgBrbhSSLEpkXONVe26F35TQ5MVlPzSJXn3J3zIakkCNC+FT4jb88/9HrZc7w
dM+GI09ZZBS63kUeGTC7ZZ58xw1AKIJmL9TxHid2CwyZKcF6m5w6CtaABC1XFpTOUymCUfk/5T8Q
U+b2bxSbxvy8m3ga/FATy7uiCtKiNDU6GzCnIX27+o0nI2lb9fIWyz5r0G0/D4Dkk8A/hq1SEtA7
t6l/hPBri1sRsuYXiFeV8RC/ROTlGHY561Cg4iGzahdXdUjrowoxDMabYJhBqycOBgarODX0xVhz
/G3hfmjiUVbWg0mntzIt3g+NRsHgfFZTCTyKGkQ4gjXDHIaKVcs1zYof5rUsHVfW6toVIOkVSWn3
1EWg3rhmiiDQZ6wbDm1dSmpEYW/X1V0Qc0LI3g96VDggZim1kNSlQNwkzfC5btyKW0tINZIDr+aZ
OujE76O2h/9p11YdlLhT2PubvtCBmLZ/nUVDGNblnHKm2sKUDKZh5F1BQiy6LyjEnGr6D1la8Qg+
J1sDfBtu/1iAqJGPEKCvgBdwFvpzNSp+8wJX3GkIMKwviYcVQk+IYc+fbsQJGVUH+Wx1c+PhnSvG
3up09+99edn9pDHEeTYY6eMQ/Ko4CBKIjzFSqIGCi74TK5xgFtS21AY63r3GcpokKm8c9iUu82mj
7PvvEKNYFLy2uTw8CAhUlt9LLHMmrmUN7gwKacxMJeJj3QBlJHizLKkNHIKhQTsu4e/VphsAgnQf
yjB+m1IDkDNIM6WelaeYhhALGbl/aRslz9wKCbbZpIaI7lmdDiG3lG71R9zhu6FukZcTYcRKZ2Rb
2173A6j1kSZW7g7yC39dLbidBy+U0p5JSEaJTw6kfjJPboa0UuHAfY8aI+E0I6JWCh2dtkob58JF
sSsGfHEHLOGuqdDGfNW/f0VoriOOzAJ0ZNVDj+2DF8p5av9tLpDVembglVncndWGICTSCNvzAaKi
kPfRpRuelraY+u3EeH6e+ErDJXNDv5jgVFkskAtO+HYRFpyTl33P4xfjyE66aZQRzN9hFt/kpamx
pEiW3Sm5sZnSimHTj2cmb2S7AVySSXJCfyU51H2ZGbuZM5G14yy+OdrSUFp55I0TzKBLS5vSEr8I
EYSVTNt1rlF1ft60QNPrgTTuGX1tqVp+nhyS9S03Fdq5DMG2NLhX2GZye2txBmsRSFCgm03rxkr3
W/a5h/EyuB7r/CHwVnh84u+BsA29PnpIXMFqL95DcM98Duca7is7EqjpptqacbHWAGSmJaY51Gyk
099H6yYamYxtO+Uqnw15RWtybxUQ9YZVK9LwROEzwk3Auh7ayrNHe7c6o7TRdKw2iHu2GeGobkg9
jFiul3S956f1B7ECpWGpffQ9HZZryI3szdNOVmMcdBqISpLIvy2GihIGPqS1MlMKV9xnOhzTZ11F
2g1UyUF2jKrvyx+Sy0kyOpwzKRSjj+w1hNq7jUp2efFdD+Z5YMpmJEGlyqVTh4lp5DciXlr8ZJOl
HnPj4LRrDX0OM3ONE/BvyQJ0Tpoj3lYKJdnzQQL/d/dxLmeDWMuIQdt04qItBJm2nM2wIa1q3etP
vxfeRTvJoeXrVId+eecHDP7luP/fMV97qkB1RNtOt2e5x5u4JAblpUtCEu8kVxrrF0SfN9z6Lg44
bNR783+21PsVLKy/Nn6ivrPisaCtkiNaUIZ9zP2LnApkPUMgARybvjPHXrpnRBdUSpr9aPTzNxMF
Ylc5qZc7Xz16ZC4HeCdWO1/npx+kr4rskpR+HRC5uwlOA3h/FWAiS2ukTm8m2rqgN/zVyuYetc0u
lcpRDdXKQervZl8kuZpTdhHBD/fKaySKtuop8X+z1bpkA1QgeRO0cmUPmr3uCcEPNIjhh3q9FB3W
czDmVmRXZC8eZJxjJUkcTdTm80uKIRR/hPbdiuOtxfO7EMPXuoQ+jGKU7f1uNSMj7A7GH4tu16Kv
Y4N0Ua1FEGbq05GiuifXpttWlUAUzyNToY+Bphr5hnYC/uzUjlf5jrspm5S15R3AFZju6uuIA/c3
xZ97BmK6/2aGxw38LZ7g/gZAC1hfHfyhSQ5/HInbpnLGWUoEAYDbG5FtizrPukENrNg9XifmOWgx
JFLBG6T54eMIauLzLe59sD+Gi6X2R7b9PGt0SgF79z+R9y8GWYBg+6jc/a/uRjXANC7XJ19iaqex
agHF4nFAkoHZzZidzBqgONYezkyWUNJ4XqMxQpkFHQGbO9A2nH9Q1kSttTHnU2aEgGT1DW/lvDYB
rPx5Gj19LcW62JzQ83AiFT68MAJK1Jm/N/NlXarbCDayoYp83wKBzXSQgz2b8/Cz7Vqg1CWZT43L
9tNhHkKaU+w8HS+FuLNhF682AboXe5kJDE4A34BzXbWbdVu9ycBCSlyBiRIP6EtmLB7pn0vQ/sey
dH6wyC2jK2eNuAlq48unL8MYhb8sXcqeo5jrfKGoyhLaD4scrqXKkNemMNEjCdIQtDQgbB/YJMIv
ncMvJrAiW8x5qhcHvKgd/gV1gtv8lNRIlLxk4FhIZMKBFxeFVml1r+G1Tcy+T3xIufJKqgp/6SvA
M85acZXRy65/LR70zMaRduN6qo6+kczPY9jhMiA8dQ8ZCtHODHTtpLyfyyMPQULTKMliSUpeNaQE
ajPVQ1CCgbB+aNqo1BRG6Gc/YApo1ChinZ5F5cZzdvkpZHmtMc2P8iJKlhiXqS5J14FQwtX8ju5t
wnltwDZw6PKNMUK6Z+QPwBs/8085qLBJW5cO/RkR4NbKA4vqWSCaCk8UzAYIniltJFMpRJzGtNiW
O8fISZxrYOaEj8gis1+P65uOUvAxbpjGQuMbOglCFZNHs2kSnb+2VqBXFBUnRcgo2x4UX8yJxpYs
KnhIIr9/qzFAO82n+Pyixzs7csdVBTtGAxIdthhiwXY3vaiSZWop/iCllrCsOzVMS6FHTL711qsn
kcekcUJxHl89NiXbI8rPmE5dtqBgGu2MX8TcaM551Xff6lm6+eu0a08MVlt9n9zLwrr+soB4Ve4Y
r1LwkFEZMpf+mdgdX1/NYT3Dj3J4xU+ApPTibSR3/9U48gzL+7QN4X9dmetw0QyazK9ZNk1RfAJ8
fygHptnwNI+Nzj3vyg5wxeze//VTwofXyplbxrVn4+JH6sL4mq+W3K6m5eAX6kBOoeGuMEsUqNCs
UC9JCwBXBvyYU6qucgq0MoFCePXjyxIf72W/bRRigB0BOlkyVxsC+n7uL792XanVP7jH7b8Uzj/X
3EhhpRJ+j62eWG6D4o54jFMU7Qq4cOOSD0/Jk+rh5TtSCU9aZNiaJBRni43bbnzbaUknDuIquTht
qhOwXzOVZ4+KGYjHrBfzGbFv9dJCdV5EmEBfVMwPtiY9nMIS57lOwnaKmnfzKkkneSMPPFLfbLgE
epiGMlR8GyCMHGV1cl0GacYyGgTGtE6RRNXPx8CALNB9T7blHo0FahxWPjk9MNyzZhhhtomRT9Cg
Y67V7um+uRGjJ7gYxsLV+Nxjye81+kxUOpH21N6G6aogdZ8vudNieJGplrSbZRrjz+sqxL3ahTll
D8tf8am3JZ2cBp2PXjAQ4yL2Q07J0L2ocPNSPSjzmnVbBMYAv6x99tsH8bFxhNgSf7mcyvPySulG
TeUtR72r1ydDvW/D4TiCsC2QJkhhTaT59yO5NGOBuKdtkiGANnq50OE5aBApvwOMnepfB2sWOCbv
S+558mu8GvfKApyoJQ+cqi/6XC0BVVxDchhNKnDTy8jVGX8mjQhjNxzscQ2ybu8rFT3nYURDhBe6
uneetmd5vtyRVzeKH/WGLsc6zsu/KjopP5T/++IwHhhFSRx74i+/lYLjoCX6maKT2KTxzdlev2WZ
mSGIw0a0zz/9zb0n0vFolHo6/4EbbzB7PZ3llUDgU3gRQL18VqBjVWsAau4rIDbdr0FIgwUUQTF+
dvuBPFCLMAOzJQzemG+ruGbFHBeMfFEX29czgSPkTs9DAh1z/Ja+8tJdbQ/Z8CagCyurCzh85oGe
T2x6sfzyKtTGsuHfsG1hSJ4PpMkEig1GdJ+cyGWA1TuRWrErHPL22vFjogsYnFFxj6T3QKwxeSGl
r3ziv7YIP03GisiAhnpKT3XpGZI8dKr2Nnq1psA++uTuh0AWPaXjx3KxW8MjEV+78+6E+0CJXjSx
ZXSkeVr1qBgiVLMBf9P+jbAY7YMLDI0dJSObHRu0wTovQIMCdUbI1BjTDXuPtnFUpKgsyAIeEPB+
CcvRPuIbUiO8kymUpmz/2ohD60nMJgjEmWZcmMZ2kI9SI8rCMbgq7+RbgKYjXbca97mylJDn4nQc
1owCalGFi3lEpimk/6JhKrp2GnxhMyk70Hq/jmheIQ/hKxmMmL8XrmjtpgEXhrGgO1eQzxeqI2VY
nYfMnvS7RC9/EtOMEF9r7G2bgqU9xAA10LJaVJ3y7jbtFr4WsaioLGIq6jent3bJL14IeV1j57c2
0a/AlHoB5CUYSigPnP1cAzHbTzPkqE019thy++CwHVuLdZXkdsplF0RpeofrXuBSr2khR44nOeSp
67utquvYN+MLwX0sFgRAjlxw3xtSDd1j2+XY7sBqaUEyXXmoLp5WwFOEEWa7C1JsR02G/YTQHNZy
UuQeSz+hwwYrsB+JS3Ktze2FswzmaTe+gErEragpoot51PptFCGJoCZMB38JqaEgb0+x3KlSStyg
Pc1Qd6C+Kze32DobPHmfV/SQmz9PmoO2NAXe8Dff9GYJ76L2GICFVjHEG0F8K0NP0XFLFoub/52b
sMGu7SnPZolg8wNXEGV9mkttrmd6Nmpu9PcPp0tGS6XXZ+X4VdJOH/slwUHnRHrl1g+19fsHAgyj
yqNvmmAJcKPk058myprf97xxuBQntV6+R5di7ep7iJ4jeN/fjX0NfHNqw6MBZBufB7oZZG71O2CE
22wEkPMIuVEg45E83lEpvd8c+XHsKtaXIzSQA9wRbxtteKTmOMO/pbOmjkGy7jWAx4N00bTpDPFy
mgILa5YaTLwiIvOS3e3m82UHByJqi+tyqnx2p7PrWXPgKNjICpZq+7br0cyzAkVl0wnhQ375Z7dh
2LuUusk+9U/TGbwcnsEYZNp69udcgD3IbfCHWMqVBYxxhh+itD0NfSU5ImRS3XVx2Zp5SEOLVAp7
9awA0TfIQ59KkyYHWOvYX1rV7Mx4/PoNilN1/XuXmmGwHqJCxBZsksu+q61Q5YfBzcdRCv1IiZZ3
HfcH4W1CHTVBd8gh3dOfCV9SmJnKz+VeP0LvSkogJ6Ogmr6NZliOT51rqgkYo7s8kHLJVL0M7IfI
yOM44qNvbn4CdGc3KX/GMc6g/DzclfPgnTNki04PGydhc4NpXxz6ZI+Mp2du6kqgyH50d0BMUsKV
AxgiEnmDL/VYDEU8l+GdHZfWus690RlaftPHM7z6iWonkP8sCaRFvs9QAmGxTWvSoKZKJqLRDvho
3R7/XgZi22KKONPmrl8NBUckwdCiNa9VEf89YtX2kjPf/pkHwrWXc9eSj01mXhcPPqCZdqSOud2I
3jRl3ywLfm3O4cmWryFEQxjOXA4H/gCXv4t+h1FxD8t7KH/6eH8fxeRJPNlukYTVq7EvSAv7E79w
g9byKW2IhH9xZkkfay/udf+HVGd4n7rhchSZVQ3MBFA2fJJBdj+OUI4tmVPAXb48R+99aWA67Txm
f9haIk1p3G+cb0aPv9GPHkf2zaxhTx0yNCcYf0zy2n6XIRy74MBrUSiAR6rDFDBywIVCoWHSIA52
oWI8jAYglAJA/qb5PsqkhCAbDibzzPStcam/8pjfIVigrMxD/DAMUqq4s3KMSqgXg7RIwZJe2x2u
9NsGHo1YMJ8Fipg2SbggGCyz78nYZhM69MP2/58MK1+R47OMS7XUZ6ZpGlXPuIXlzPEI9+2a7sJX
ipmnE2EpH34nGlV2fGNbWq2fp7Hj7J8p94dfLd2X9zZrXU/OYqRZ2vmtLdHz880yeXqVf4U13hNq
pGuPiFYEXcnyZXPnbeuDMKEALK+iHbNLnK3f/fbkniocw+CbKGL7Mlg8i4K4C7rVGk8zJ3EhUfUl
+JKrdcqYZt3owAs0tO5i60a7CLTjusNykCTD7HdvRLM6TFm/fwACtQi3PSUx19Ehzv71KbnhNjbh
cB4qy/qqBvliV22OrxTETppKLWXy+cUvB+r0neWiD9SLzOQrM3yY/ZHjHkGrohfEvx2ommmI33Z8
jUNf+b0vEIwcEDt9uBJ95AYvhrMPkXHqZVWjSMdTDSJkNeYPEnv9Ei3FnXsPNnrdDPB+uoJ6+wAD
AvN/gFOmjwQkYOspsRtMHgWG7ICBpi8XAf+Qvvs+EEpnQ4sDMTRcT7LbO9+gYzkHkXgFhWrmMwZP
+XJIsIxj8H0ANjN82TgpnkAtkn144BYGF6jpUSLYcBMCfdSWoFXQinNMCgtCnPDvUlobBr2BqSqb
wMHg9HIiRdgjh7e1aKlsJ/0kbepcZQjaxitR835S7Rmamu+Vn7m2xdHXXPOz3VPtoU5XogIZ+6G6
8314iauUU+FsU3iREVE3zzUzHIj19KxHWCZ9CTgO7tSugme5yd6Ewu4ly2lutxLuJtGsfST515jL
tFkf8dVXW7GeEZPXqtfmYs3FiCkq+ZWJC6XqGFD9Q5Hhw0abPltlv8RBzvv/3b4XDvDrKJEX8pxd
/kNjFaCk1n1gKMnHmWwypznv7AmUw3hvXQ6/RNX6X8VRlXybgihow9r/XDcABMd5y5z+DgeX0klq
lT75VMv4ZTEKVxqSD2UPUa3K12srRMCvO9/4jzj3E3eSmBb8rMnzwLojEH0bP/hpwPWIdeCe35b3
NKusaF/bb1oSfw76jbyaI9BgNbnUbDH+lb+ClCJc8443zIJuyIerY2Rl7ueoaTYstf+lorGpVguU
nw4RdYr/kglnoltcZk8VWADGgs+Y8htfIBlcQTzE7A2N3ga+RXWV9xJaRg276ZWv/LgolT1UvvMT
zeg6G8Cq+W5Plfi4e6BYBdk/v7B9Q2am6MTX3gER2qYEk1c7aDBDM+nmRS0zwacXLyideNFGJsYI
jaSFhf+dfJN0Ne1G5xrxDBukgD8mjQNwbYsqa9uLeneDMvgKCMo+RPEUEJt2NZzHH7RhGeaT06yp
3D8GswTZkBsiNn7QOX4vkfToaN4mGFkArudPU/nShK/F3e5s4AXtoAWwch3QjDJNZ37/85K+Sz+B
KrwZjCorMsmQ4Tvo88UuoTMaaD56ILhaOGkt9YSZCnJjiegtpcl4fIzyqqPl+ufxjQM/GVBHtTBJ
dWojCdb50hz3j4r5dHL0X+aAMjWVcbAcQDmljBb/aqdOG2mFy4daC3YqNGsJvTwTBhLexqbZqxTV
/8dB06oPflt/j493LyaQk8HnzFaDzP4yWP6606Rdmvx7axjSpWboBuHJUbgT+TIUZx/reDvwEEf6
YeRmb2LK8G6RdhQ/KDrFcfkp1IzdM0i/ZlmnUgfX+6Rh26vMHySfnV9KP8QgCM4Q6HvEMIMiqXQu
acnCnAGwTuEJBS0Pub4Ile1ewJZMESZty5d/A7Ob+4xYdVL3OC+QbWtwEQ+5qWg3UInUH7l5kWJb
E6rvtSlfZwnWH3QWMDh+TbDV+2YWiDCed2Sbdmpc5REJNMGeHNabj8Z4hvkS3ZbOxbalfQ3biMct
loU27gKr7hNqnhuQ4lSDfW7lYLtI0GNlxWwONMtqjYwXqdAy7u4oE7EGnwDp2YFf4S/GkgR8rQYf
pC87xyH95b4PHwJPZmGb4x0da/hdrH6ormbUa3HVUQazn3DiyuV4TCBl5Oz+VZKsUTYduY9SPlR1
S6CI3qdlV78Zx5x7e2H35q8KrL84hnpqwU3SBLHmStlWFFKaLnRkFsPggA+beWA3GmoMfovxsKWk
QyCOGNlaH+RM5qWEWWl+jI45bRPKjdTP8cMLF792lrtJQ/vqdyU69JL0w+CHLftjo/55CisPL99x
g/UAM+uOf43AYwjVtDaDsgfpZV+pEiNm5nkyiOyaDH24x0w4Kl5C/QLQhmEwpb5Lo+a/Jg3rJNr/
Wx0rO+Z0MdwmJDJ51YmcnGiubzbGyVflL0//uQ3RQ4sZ46MczU0FhmIh2Nbf3pnmXrprieAEOYYx
r5lc8Rz6cJgsyODjoAn1L3fA0tq7ZP95J07FaDsL9NMvM9zdtVe18sHtLEB8gyfJFJxg8VKQ5vSz
2chpac080wKze/S7ojEzgoePga047FmLXZLEz+8+1ZoEfeT7Cimbsky8gLhgAVF6sy1ObR6nI09h
Vpa2mdgv+kij2r3dvI49QDtWu/IS+5RurKkzj8ph6q6bHM1z1Ci0+gJDXLoG/U8htNcJ0w5wY8ym
fBzkGVEnVVoL9r7SMOjp5sufmI/ITZWZgasjfGBoy6Rxo5jeR9LkKV/b916OyV5zAsx1ZUHZk9gX
vKFcNfhTHMRp+W0VLM0AYWSgBJeGOr7yslG7Q/ZyVeuk66O7VXJhbTXSClzxHu8zFMExOzvPoMUk
HT795iPCuIIXNkKesquCDz7WAQjNfyXgy1OYc0TOBTiZPjyG6xvB+NUnmxdzLKmnA3Vp6qRXTbfi
0BCKcM+iGozFDEDpxhhO4F62J/HBk+JnJ2y2UXhOZ50v0u27eLW9JkLUpbKEA3XXI4tv7jHWcFLo
xuJ420cECzqm1XbHT1bus+0ebJ+sKkOhkoH+tbxk9O5U1+gLRx6FQLtpEKee8jGXbL7RyTfZ04zx
POPNkNowKQA7HOahc79W1UIhg5itjbWtfNkxaNgWRhdgj9n2zbX8CZzo6JObkB4NO4tWZ3mzzgzZ
oCgw6qQYyAxoY6hyGDy/QxYHFUi4ltBmGkRSoIuJKsqlLJoIA/d48d5eeBFrut2AcMYxXWHTgmea
pIxc2AcUEj47kbNA3w3E7WmnohNYTu4J4uoDh1XKMCnsyD6/pAwsxLv0JNctJIEAxJCSbBKqUFJQ
Xgdm3dL6Cf3KY+4hTC3ZmVLMeZbgf51dQeo5G6RhMYtOWU8xnY2loodxBOYAbnYR7nElZt1/ztd7
i4eJ9UWvkuh92JfeOoHN66HeUqwiAfTQYJJSrwnBgjsKZCdRWjHY5fZuM4kl9VsqAD4vSkcKvSHU
MQKkpLmjtMoxxn1eJGFW7k0DdlnPwBFtyQsSmntKXuqpNcDqhUhvZvZH23LERmTUxhray7ZMxofF
EfdNPuw3CBlhdJuOzkBfv2XM6nnJXlsTggLmpmRzncsmPZ0WGWfuAmGQNrlDLXACkf9vkUVwHNkC
dKLLDxXGgUVD2rOXfbsc2cR2pmrmUY+y9I1lZNzi+MLeVFzIdiRxaWzhN9QJZxUKYgwdvqeRF9WP
8QGfrpWQz5B7lDVkoclxz6oYG3jw4QiHCsgnX+ADzQFkbTH7aoze4cfkQxrHoDOpRbJdD1j76KFk
5BmKFqrD+IphFws91Ms848vE+KZ3QGhdaBnrDEKqEKNSpaRR4xvkVLy4KWKm2hRZAXmMA1a8K4Nd
OgwF/DuIBun3/EWjOhkUJxdCguoDc0rAPXmCwKM2w3b2ci8zhKQGx4/gRvhSrwWetcQv/ipkoRJc
7sM8QyMT2bybOZjvM0+MKgPejE3dfV4ExJOBG88hqS3M0u0OXCQYrCpUV5EM1THS6Lc83soeMxrf
DtoYuCrS78ugYwE8Uk781r+9BiptpLj6QaN+Xnp+Hjum2Sh0zTrQIyly2+AVn2drI0j3ITB9r8GJ
Bl0K8vY5hVVgRld9FJcHH8bN5yKPfd4tCVz3w6wEvSyygoXM8e8GqFO8apbmY5tNYAzR7n+Z9z7t
drY5qUm7Av5f3QpaR9tIMYr3a3CHzyrPgry8lEh2tNBsOwSKsaM6cIJzRp9N2I0sqZvxpQsDiTVI
kkk+gqiiNTJ4rnn+DoT4/LbwblTGz/KasmZF+KWdAHmH55lCfKRqQ+vC5I8GttFOYK8Vr5uHz1WB
twyBijCm8z5kFv0rts6EEDh9PIqrj4NhnMEAIMFc7Ig7h+RRwQ2Azxrw3LPZlHGcjuL9pdctvx15
IjI7i28yzHax+H4nqXoijCe/eOC0HkPvPQV1Fpq/SJrsyu7IkzZK2/qsVnnRDuveWw7JQIYUxE18
JDu4D7GhWrErWv8f2zDsBGliBhJoQlpkpY+zWSxo5JbYz1ma5haa6x3f/OKkteymIXy1q0Hu/AU8
WHyxt09vlJrg5QnrsPZ0qyqjNsJnC4DyQnCoR+D+SfaZg9LKgJTXnpUwxvId7x5scC3pq39NKOOo
2wYk2Kn4n0F+Q0nR4KM6Wjfko2JvvHrPDReeVvhqlGiNwXslZr+tjgpFwj1TWUXlq7PrJz22dO3a
MvcujIaG6mY2BTvfGWv4cxf3Ke/y40icT94wfL/Pgd25B987rdj4vune0sqLDhz56D9HD7RciQ9d
kxovaVHoMlXoVk4gswi53/5ukW6G9KtZcdo6OQYWMkxUDTgy7+OARhPfXL4yMFeZhtvXiON3yaJI
ENTi5wMeVBkJp5q45MMYPwSGRmzGiRoIoJnv+M/NvKcA7CCDTx7rKW1VVjbcuv2DKap98R7E6Arm
WegbOQaPAFoWxqPD2TzzaMjPwMLECFJd5nQwlYdZDplz2tiE2AA+dw5s2Mr9Yitgwn4FyEE6foqK
cX/5rh7/1EYt67CpVlWoLUZL5BrmUH9NPVUndPp/ojnIeL7V49YeDHqHKmSWNQxoecac3dHsTe+m
2VuS8S9SKf0tms3VVZlwjbb11q9aMuzUrX+8BBxAfNhj2nMRsIwreF1sl6H2850kvsdzP2t/Wdng
wsqEol+UwkTWWbuBSgesHmc2XqLrf5FlvNJdGR38cPTFmOFSPQ9PAahPcgBG6T3lUK0QodVgkhGo
w3kdA6ihzW5Q8O0cOvmkkUV40kE7ImvUOq75jWncyyAhDPx8vLfNb+Jt8L03nTzdRN+rxK/T9rKt
jBrYpmhlG+agGZ9zMqkkZIxqbf64/biZF8VY7P9Pe1hQgF3cKKxSMZy4RlYzWbJZO8ujcgg3qeBc
dQoQ4w6VI6kTU00OJv/TecPvt811HY6jjIq7Mx/eMFyCmcZz5H0UsHq2XZAtOjIyAmRTVXvOYCyL
iWvsnqoijjttz3IgTAjKnpX3ZhSqf0tp67KVfNGSA2N2Dxx85xVmVwqBXh6xOcu6WgFy0QnVezIx
zjJeFUG8lSu5zhKu1CvMkBTK9NOAbtBIPQ5DSDWJOTXfxLPsDs0mN7RXwwhFuSnV3AWRbKYraNtI
/GJnnmFDAkesXkqyLJUlayeF5PGBwCKBXNy6IGDQUvnRIx0Z2mCIYPUImlvH0edzLqLgf2Qkku7I
H/mW5T1N7C5WXzZNePdod9G7pNwNByhd0AHii1nceJFBXBfh3CDayrtW5ioBZlzG/gBLtL3pVsTR
jOCxopVnmCwF1TyyYzGd0efQoDKnhgU8kGDSUpcQ8ZvxjjF7k0XWWd1BoZDJ52At0VeEyZRQiQ7K
qu4f7MB6oNGM0b2UIjMN2lBZ+eu/fHnhVYAV+7SufovbQkMU1EeRs2RLZn9T9FJjbCTl+x3IwCEU
C2AUIX247QlbBFSq78TBj++vYLZxM0JNfe2aJntwyDhM8KA8RyBuTsetQ9OacQ2/7fJNtS5dZP9i
PuM7txS1giQw9vS9W/9nMUDnOtp9NaU2FXoTBdUVeyCcG/SOioBZC3hE8pCOv0jET5ojo/071ngx
v+JCxs78/Trct+ukiOzk2PcWOs6SFrR2Z/3SjWaRz+N2K2QKejf5XFfmky7KvWUnBfJYNMxoU85W
jsSF4PHvv32mFof6TlieRXtSu3no5bJ8q5G9pybWBAXEwqeC0SkQk06U0fIMJmXl8NYSQjVFKAbr
xmXhQPS86hkagK5wFKGOQr6GuB9X5TT9IHxD9GVHSbCgZo1kSm0Lb+SctoFuWXxzusELdCJ3rOtK
KsPhblkuQkkWIrh95fqzYS6WyKk9/XwoHR0+HjwcaRoFrA7hx2s6Pwd/ptBy9vYqDkeEGpN7MhID
sXefnmMqYF60iwdrmhfC+Toh3B+qQ2UaR91yznYGDKvl00Y5Ed7aDAygSHnVBrKtPKpPm1Cs11RL
/xBg/zjz8WswEXu1+cP4ZEo/Bpr9TIwdLR2iylIeav9C72X65i8hVEub0azzM7zXUq4MLHboTgUx
16aZUxoO464U9o14q/u/8MH1PyA0ibKWV51dHAk6Ktid6+qZCcfF17hV9SIvmrqQv6IcIEXoCsER
TokiH+J1fy7E457+QNIm/i6lTnMQTSU/1FEetC7nmMFp8oRmQFrQwIhqV4r8vGsjlTyuQwQk9IV3
FRXl4/Zk5HGOHrjgkrNxZHHuZ4NvpPVDMYtYI7Nrsw/CkZFS0YH2d8y0qQKlRbtac9wVTG6HkD+h
FFGte7WOYrrhOE5jYuWKZAN6gBCizCM+PYFSu+4wwv2uWRN5MLxc9DNJ/rG8/92kugIhdLk2RNzm
DN8HyRKi9X3swJyMnNFvX8dSF0MHYKo0SRyl+AMA6vKUYS+qXQKTfdyFlK+cYTLTBXpzx881xxBZ
b/0hT7X5gJCEIE3rn4G33Gq1k7lYlBrc6ARsUBuOZr+uJkviXDdUmuJp7vEJ303n0OwW60P5XrCp
BroGE+PC453GXSddFVdU5QfJWKuyO7CIQ2r7FPBJvUwroxc+ey9MIyHR3+hoefn62YNQYsSTaepT
0J0Kw7O97iTksKFmDfSXySBtjSmwNVQ50tUH38rwtm/vivajIxPBl6zCcH5SV8bLqgUuFv7BiskG
Q2km78W52gXy0dYYBt4XAp00mAn0c3rYmCrT/wI4kLGAvfvi/5dR5f4lrcbUf92AMU2RhTfWleed
Stfj43kJ8YKufIwsJzRKkj4eESvU/PU7OTHE5K8TI7jS1yGELbWoFAApJW2n7IXoYv8a5e+5pdHN
hvuo5hQZkX0cDrikB/IVtTWCymX9TERSfRoeif0b4zwrTUnAHfkTGZAIyT0hqTWq/63gdduG2R69
wwVUCeYjVVGc4YbPeSgFY6nZ9EB9IMtzrhMQvEbXyTr4hc+2721MnFoqXU5cx69wqoBdqGVFkJMF
G8nmH+zSCGAb5B51lxkrSvY+HhgLSs1RA/fmX1pe4qHEgeLTw4rElF0r4MSKQwjaOV0jXFEkEJVC
7fQdvYf8ua8R4f3B5gAJsVjCG7zTUuUGG1xfYrGYcBCrPLHEHWTZk2vGtq/RTFOMzn7SSojSFomc
Q2McRIiDHt9DYWQnVSrqBF17oAlDzxUSAgL4ics2bX3VfXGMmNpTTE/CrMy1oA7bLqV+ALFO9dIm
bV03cmuNH8lvy9Wh4RSl/wc7IlDNghdRIELwtOriy2xDTOuelKyuVFi5+KTMxxhMcYdcPT+tEQdh
B3+EUY7mHeiPp4WcsfADT8QcSsDm01eYFkIl355DlViFqsBsuITY0bYhgZILAhA8/o2tyjrrDFDU
dk+2bsk/NahBV9T//15bjMXD2BQbBQuI9DXoYfbm5my2/3SYn6TpoW7Y4s0lZK3di+RBn60w1vjY
m41p+xiC9kmvWVI5z7SX2Hoq1SOB88zkAZNdL5Yyqs22aOH9+vziWTTpCiO1RsPmKd6xF6HqTmA0
Ny9iQkS1oz32PgOQNStE/nytEMxRgJkxh8Yqvf/UKKmfcerAnNfZTfj9UurJOPTaRUloLJvR4BxW
5C86tE6l2kg9M302MyBacBB72sdHGhkTTqMkectZDR/7dTLIMGk9VVfCcg2dZHhcli6KxDV8QSGo
Dw1ety3rrpsfzjjG761UYzUB498Vi1SCt+NzBYGGKlegzAG/+S5RrU17fe6e2rzg7+P7KOEx+0Ro
tqzQJirPXJMldiWWeCymSrx4bPvfB6yzkJGvTGBgsLRcG7j9gHlgF1K2cQFyoNvu0OVw+V85szkc
y+94seLyYl+jKYc+tyC31XyWKcaHU1hWpiGHhMQ/8/lkIjDQggRrEzyN0+XPV5hiXjfVfXWkUBTM
8Hzd9beeTFqcn4nop0iCSz1NRh0WO3TAacEZYYchDxcEnMqe8FlqLl+WRTFCHqK1giJUnZuEAnHQ
WLhWc7oHflpiHo2V4MaDFTeDrITMfmSX2t5AzepqcjP4/4Pm3uAjgp03emmq9x6MOfCFkyLbRBGT
lKnGnXPdICyIcpxvJM94rd6EXLNMCWcp6iizCQea9rsYPu4b01Rf+9kC8pUdKDFT5f5UDDIsouUu
PR4Q4CplIHD+biOaEDKiR5C+4yF6BLq87z7SYhY8iXeuoxsl7h0kgOLobvZLrUjONAlLROZqsDm2
G0HEyxhRkraT4Qzwap8jqRaVpmRUHiBtXjLTT9FqA8VPPMCu3NlTcyTWj00MNYtNRwBcCU70wBkw
prLmg2wAH31Lj54wZzxtz27qpShNRn9e2FUJ9qJE5PVHkEhMesf1Vso1Yqb6kmfS15Ev4dYmFBdU
wH/Hm8dWbRG2mQElECQBYI/rTp9Pbj1lzShLQa3BmM4yTj/1kqO7KnQfWIb5FUcUJTX/u7RwPhzh
p23zv97L8LyGyN+eQNGtcDvAEMTnkXzFHA0jtrDwCM0dm3Etu2vQtL0zvLpnY6dTncuTy6fsw82N
l89A0C66DzrZDonXJdRKJ1nOCjjf5pj3er4msvxvdlXbQSBKRmNVrTPWQBJeNXMfWPavcU7KC72p
4DwaCEaouHpkPZL7DV61h5UwlOvhQm5mfwo3NOHOr1DukBzUGQ83CaWIBbg5BLBEdBtFfRKBOuXJ
XNuI+WfWVCnzVFjp+cYZ+eO9w30UTm2tAkzKuzkhuSvbRiHN3p6gAFQfYUA5heeESWuGl6ZPCxHX
JguHye9t65up5c9UlonlIJEULN9GG3Km3rADj2XlG4fgl1Au9qKkp7ICvbQI+SKmQqxT7/droBMN
zA97XTmqK6cya5B11mGcwdVzzrw8uOYS5WV09bmshi004k+y2BzLjpmvoEsToiM70mwRAHiWzkHV
Jy1HVeoJVSlafyB2Uq8M6DKRL3m1xQQl81LbR0QhICTuK2jH0NU5As4sonkgpdCFSCWI8Cw8GwzC
F42FGEUpVRSl+6o6BLQMQQFzYBFiaQs/vdjaX9DOSxPnQTin19W31X+f78Q4feGwCqhdHjxUaNB0
5xZB8KEZlFd/PqoIU1kojV+zMZgbmeX6Kr3lB4SlGKrq0G+xE2jPbkLLFKhOMJZp/aioFhxkB7BA
7a1pY5G4YJFfekz/J3DOc1zRwYY0cMbphwezfCL/LWnzQ6GcjkaqC361OYYQzh8rIgywHzVKdQeH
NfmcsrpF0cO8n4c6zLmPuQfd0512+5NLouJDu37XbBAgja7+L9hqaQYlcsYB7sVO2MKy2Jxu+I+p
38dJg4U8uptkmkgt9jnS7ODd+TkHoQ8MD3QPctpiVOprNoiv5AKu2qP5slMZtAw7P0dt9TrrpiJI
TWJK7OgyyfugnM9//Jr/+BgXh12opq/R6JZmUV5MoHHsPbRiS/b2L4iXnpPbrvdhKYWVpus9f1mQ
2Yv1Vs4FSmIKygM9xNFWRxz404wrJqaBgtKTswA+nhr7agPILil1U5MReUn/MXe4dF3Iz0YXqp9u
D4ctSivTBXDkbhy0xRIqQdHf/hpOmtdWtm0wIP5u0qoKk1uC5Qzhl4EsN+w/ATIIAKwJl8CZNMrY
T212zlzQ8m6GxmMPo2cDUKbYqV/qlb1sH2CRcGt2ATQe8zY2DSwoNk4aAh9A2KzeeQTz76Z3B2Y+
RL+amVdbUUp5koEAaYHvqrd0RAAE07Kk4S4HWQO0bFVUQsw4Z6qCnRIKHLvzrgY/TEWhVhHIo2fc
blHTXroqDh07JKSSl6bPs4+eIcQcba/SygAFX63WrwbXyXUHUzcimGKf9GruIvFRXBpavaBbkfqA
NSkAB0RqokbonVDJWQYBeUtW+a9AE9uQ8Jdl85OPqo4X7egcIVsfUVt6ba6he/yE9ZxLBvJnDLMH
PeL9HkagRlo/E9Lqc5jntW5YNS0Xxa30Y4ya1IbP2C3oBdwWi3j8LoeQGb9Pe11lBMEqMSEeSNrY
Y/1JYNBooJCinaPgUSfEjHOllUuUM452sMO7xjPPiufiaAmE3+cnHiYU5+xt7waS1N2hEQz+Xhoj
gY2NCMlNdVr3TLMW5nhe6ufKCCa9G1tRAaDYWcVjeFyQqCtOx5NQSeksRJ5TyLuZrlCoyJlCl8Y4
mrqkc/tn8JqoCq8xtz3i4MDwVinlvf4HLTq2aGS2E9TgoQIt77I9/yUMr4FKoHloBtMbOiikU6tO
9pTclLLRA3XHyiCelNlWVM6hgNdkBgz4e3QHkAUvB1+CPT8zwz50l+T+rCiTVJ1pQr6vhXyNfKUS
yvZNjibd1hoOCkLhQzZHIa40GThrOyb4Turox22Ugsp8GJYBM5PnZMW7nj/dv+l/VqV4lQYyv0n6
ac5OPZJ7l45bbPLB0cDFj6d23WkfsLMyvMDqWc520bZeGzSrZjdiQFyBhrbplKX8NHcgxTg2sG9y
B1QlFduqjtTRds2OR2Xiydw51O9mr0JKUa2dIzyxWnvzR28kjuKaSPKem+2UAzoxSvsC4aoDIWyp
E/BTGTqrP4nPZer2cSi/xKidn8Cx3lcAQFj/77hMGdgPY5t1wVRFpPhZGv4iMp1yD2+sJ72V+83M
JBKVMTwcg3jgixr6zwSDIGjrfQX6pyJFR3FBTgO43MRBF1XlzlwK60USzZlnvQxUqc59TEK4oyr6
8D7kk743apXJGleSsjJjPFqiAPMhKhCKsp5mH5+BsgKAzaM4cA6B+2v4KG0DId1Nk497ImkFq2vJ
xBi2e791GhJat9qlXVk3Sf83gpgk5a1Na9G94D3s7jiSbyHSmQs7tfWaRjLVBfEbziKU66ssg8Or
zFxyi/TC0Dy+jJcLzSC9+cdG57J+frRi4kmxFD93rN0Fm0roQSVCiBrNPYSU0g8CHspnJS99Ytb6
fVFxwGH+bWFFvfsx2HhnxtHjqqI0alYMF9bjMTBHABCm5sxGpjKcXZUM3Dk89CM4hKNnH/hB15+D
qiPK2T+5Z1dbsP2bQGnomgYABPu7EeT7z/n+Eo1F9b3a0S6fXUO+EXD6KoYC0OmcCsYatVVezyw7
r4ey9oQdcMO55/wSRRARdFLiFF3tBBzq132+IYc5Lo1kgrUNPFZeVUCzFysztLvn59RDKh/7AcB+
ud2phO/TiVRblZ+me5LMWhGr1BDjRwVzOb3G8CuwZhicHCv4V4SICYnsoRPaW0nfCtXOD+O73ibb
0Px2Q2pGPOd7C50YpjURUlhmNswxPaJGwzjWcdnaLhGc4srsajKwgcd68RShWpU/V9s8kbJa7z6W
7YyqS9trG4axORKi6/EluCWT7fDCYLg8hxxFJW8aBKJoJHaKx2cLnuLDuz31gFK5pNF2/9Dry7A7
MuztIWmNdUcPcGHQpeaaCP5GvqRiuF4C2oyZwTyxeW9N3e4S6+YhDk+bc8j+thsP/DgwRg3igxSS
syL6N/rp1h0oYecRcShPPoLThYdtwhKIWM81mP34w2xqiGrxhWt04P439RfvbfF4WQ/rK3uPW1Sj
hd5KT6f5YUuEDkIaxpTy1CwGgGHvcikCNCa+6F2iGDvhn33XvwiZxpdcOtLmDr1rD+sVq0tQdNmC
2Tgz98jcM2QHctW6nz6h4vFw6PefyKblVK/1CTm72d7DI2QE1jk3qcCk7hAfp79e9JD4vatT0517
NCEBXZKCrjWlPNHvYXh/p3uKoTIBdV69BuDa3cdaHvXUzhpulL6hvLE/eqJOz1SmReaEK+U8fYV8
rgjf+gZdNEymuE9RZxJHxVbRPdKUTEzeL2moAVhdVxD78QqHngDzc+7YN0IStY9gzacloyd3DC23
NAROYKrLkAFpMV1QRDtUh8UxkRcMoMd2hFZnU9ZacedkN0P4ZycT5XGaR1wkM1n0sj4w4Hv7zvJU
adogAkPi5boqaPIVaUv+rmPUJ/iP5Z3PKL4070k+upagSOX8kNAEze/gDHrMA3lOfDZP28NpAMDA
h+MeZGMuucFXJ/SQKPvxOB2joxSwhtXmb83ldEWCLWt7CNxTOgmWJybdJ9xNO4N+Iv7hSggvfZKz
3PU6Wmt+ApH84uZfA8mK7tRfJECpees3yRm4r+sOHZlCH4tkNJmwmPcBINUjYJxMwuwn3171Tqik
gBFdqQirB2aD/3FelbfYeHVapYOxPttIyq5A76mxTRWQPIGrDb7saYHTYpGaqQPTaXDgu9EnjxSA
z4YoC15zgRZ8pG88E5MXeA7UsVsrPG4OggFz3GuRSUdDBhP6FneJOsWHwkO326RL17UM+1n5Nz4V
dVtSValC7/hxCfKWpwrcNgrxdZVxa2ofVz3pK2C2sMrdvLHjfOL7QOUMBCkGWk2JUvW2iHmDfSiT
CxRXtzOJQXksHDxQgGxTcvC/Y8v84U+UcThRwKNEtv97c/aiBHORN+WhP+E8LbaTFhMxQsK/nfmc
0gyreM1dRfEiXuh47Msy4Vs9Jygb8vuZ9lXi4MZPqhZJEdhm1NjeJXmMcTTivqrlGgccXM/b+WtE
P6I65GQ4MhZksTTbHupJ0prdFEZWZLt9u2oYFdLc592bHvPlmvtFWZEbgVU6T4mB9aIsXKmUJTYy
Ehdz6ZLTF8HmaROzW6SCNK79Ht/cqYi5GJ2mQcSdLG4u9/7OhLVITLHj/DZdx1e4YwJx4rCTZJez
gRUz21jXV950Kzsddl+p2sIWc8Wy8lmP+MKRDNGY8a6DhL/uud6RWNewRd1XLvT4v1SR53u0S4B0
sqZo7iAsmjD97ax9dRW6PFcOWIMuTj0aztXgAd8PEW/G6yBRf9J007gpBfMhS/Y1nqG+Uxtt0qVQ
Y/qw7t698QuikarPGMGivnubF47jqpUz0N83bKVbDoOiBGR2Qq8mb4E7QbSt8P0CPhDzksvu4Uj+
F/z8KBNE5xfMUWfEdcPuJFtPhOgMSX9fAGdhNINgks69MMnGfHcn0baeJ5tX+edHMM27CiIW1A9S
7vrQcS2wlUtHvdI7TPdOZS0XEDaUzzlTy6ALoObhP90R2osimMOcQBFFAJyXm2FqjxIUFXefIZAb
HzxFH/28Im08vSve+ma10lZZ0yAIx/AXXY+J0o2xrHPbyZ8AXxe86/S/7WJQ/gFQBRbmfA+PU+vM
mkVej2mBJKSAR8GT78u7DVY3ICXKjwQ3nqI8mFcDG3nQQrJgRpdLuseQW0tWzlsLpC50C0R5rJDl
aNt2eSyykVm/vbVfkMjG+rtkDdxQIp4jHmiUVfP5V/Y2NQMQHQ503zTHxQlhNck7+cgdI495QOYn
M+hEhN7mZL6NbprZnXgncJbC7UHElyjVtU9onGUGnUAJOHQXjT5yefMzPCtmPbWZpNYSZWhmWBhN
0mFINwJzl5sjYwz2FFAN/vyLeH7sMjjgZky46cG+WfjOFAJ4gG2CLpA19NvT9xvNlUmYBTgGPq7M
n7cAmO3fq3z4qDewuQ1R3bHZoxfwRmJD45ReHP/g/YGuhSi1I2y0HLgMUzlysJT3LRWD2u8IkBac
GHP8990+kIsBeHxsv5IcNRbPsh22nxbA2crCkY8fumgpUOHe7TR6JEfwyKijsO44wcjO+nR4THrd
J1C1i9JOvNwLj3e4EjlhrxJjD4+J8noGWyWbXV+ve8QgamQkedu24pu98jQkhiSmMGTYoHaRt2Zx
fWqC03k+rL7qWfDq/KoMqBGNo12WEzuXwXcle7BfuiL0e7Swu//w5pHlL5ZTEoj/tjYmdM+gLNby
JHz4LpEDFw5RnR9BOLjYSmwk4EY6VMBSvFWjPb51aR4++B43uwzrw2IqovJR1HO46KC5enwLpMxE
0TKP6gO6wJ1dM7J2jlVaTSAMlRAYlhSQUL3+K+pdNC75r/Hunaycyf9J1r1LmAB0XfsZ7p5wA1yL
CPSuut8yB0YkWlTHpVYcb04fhH+BWvDTJHt5gLz1ZaX/12OVyBM1f8X/pgXBRmTZ1J994ZOBx5wD
xal+h2K4QrLTiD1sKiDsuaUlGxgGnphBWuaMbKji4c+Woi2QpXiF0oImE9u9L9VTZPyaoNpORDy0
iXKO5HTWWuWAWr8odphtPbBc5kcF233NHv4tVXG3Gs248uIpJs67ZZiDe+TH7shtdRjsoF+S3QmI
aslyB6NvwqwMYh0Do3k+WOsy3+/+UsjuR7vDSqBCpzovJqfPg4Jujz0gGAYPBDhWCjFkVnRKS19z
D4ig/JmwM2XO3vdc2K43dQd3V82f1Rxh7pJaLiXzZI6ZY2pzSfE0W/P3uB8flQOkafbLDHLuzqW4
ODyMeraYRXN1aI597f26LM+IE6tufkYU/Nait9tSujW55Gr5g5Z/MbOuVNtWq1gOqXRzUd5Z9E1g
vOIkmz5BRRB8USXte+iOnfoy4U7ewfoXDFPip0ER5J2e70u3Lo+e6x//3N0UBd4w9X00LC9hQUUX
L7Bsx/38vpYUcBwyk4SCwVI8cCF3xK7tOSsCGgluCc4jX+tMGdueoYFgLzb/ScapxVmLBybVoqDE
+q3+UA1AG6DubV3Bp4eBb+bczuk82L86pdEnwdd4m5fpiCzLKnNYgU5Md77H2UWUfqYzSPHV3m/Q
nx2E5pAfkAZQS7Q8Etp/9RBmWqrtAOE6avdgNkhAAoYQcKKgzRqdytrgNM25ioM5QOUNx+MsdMYz
EIwNRUvkzHlp+ZKE69yncKkY83/Q2x6rhL0t12m+SFnpDNWBZ9R3fsZ8X5ozm5c7nB9W8a1pXQZD
7Sb+IzIIvC7i7Nn7CFb0ZI1gWf+/LgU/eszxlWujgFr1uzDRFwmVXOThAgn2QBoMz2+zPy0tR2pO
fYNwthsq5pEXrnbowKNvKoR4Hl3VWMgD/ySxuYn1Hrdo7LJ9gNeEZyYJwP0uVuyKLqRr1zMQ2hg3
k/T1YJlhyGy7CXwopc1MekpCSIK59u+P4WWSJyj7WQPy2rLopyYgHhLdGQqAJ1m8wjq5QPtwDkVa
xHz/2pBcQGP+ZrOeOSjr41gclLJiBsqIOLwllX+jL8VTIsi8BD/zkwbY2qZg64NoXqniT8WC3scP
rfL7NC8iwT9Yq2ljTdbuIxjK1n4SYSVK+516XZy5Q5q4ulL82emVVs4EAfaNuRCI15Vo/wGa/Cu4
FVNalBZJZ90BavJumONVpeDY384anIbV0eVT2LC5gtp4ZgvI0nuao0SEhd2GtcNdB+Qyp1m8b7K1
RNYxYpUes1BxLozUEB3L7e5ijC8f3qU7XqGhX7x59SqEnO9DkuK7qerL1+LuGpsAuDAbasqmlDeH
Homauw+jYFP1zTb8tWtXKHFIo1ULZy6o/5jWDJxPbLzZXfULrRir9QL8dzSKcv8gqQRRI9Pc1P80
jXhp+45LYClD9bkNXzxkAto3NS15HAY6y4e3fD1TflPKve3SBrIruK0IauTXdDWt9gpHDSAl2QJp
D5qWxPhOeFSFZSQzAnUgrqAhbdzNLrRWWs1vMtneTyuvMrU/OaQQlNLP9G0y/M0xyqU1WtpRU7jK
VF81GxsAkk9XmQK30IgW9XdGY+dIHWRt0ggsdYfAO9WO9SrkrMG7F1vmAr6W6b19kkfWWCRa7xHM
RimQeA9eXsVpRDeeozUEsXtEw4f6qPwO9Z5aussaBTNJGIDdG2l7JETawgJkHnnjfpVUIhlq4YGI
u2cJhHFsLrU0gwKU8nEtfTmdvit8ACK8UtOJDZda+7g/mYt/c+hBsgQ1EuxMLNqboOReSHfvR2QI
ADVbPimp9O+vMKDO10aoRWzVhCkrJ/8GGJgMfnKvSyuva2VtEcozFAnKz3gpesP4XBtq4M7Vpr1B
rrLu6aeIeaTwqcaqLAp+KMTdOfq47/NkEs5EjJXpHzK61yHXPw9D1J6M8OWlAcHrjLTFF3mVlGhr
F60CbUeK2iDv4J9L3cL37NoUoJ/xIuEkeV8dnu/bS0vnQPGWE/BTMojFNCSVm8b3hkhge5VG6Ze6
e4HfyVV0jXOzetJKShuoTchhOEppdZqDqjJA/oNG4A4ktnMS+ddDFXbzViurjCY8QlYGSVra5kNp
aGm0252o27K914ULNIgTmANK+UqTD7UT6eRN2fTz30yGehSFtApVIUNIRcntRqveuKey3HjDz0JB
tvbW4V6QLnpkNqCDkxRLT2+DJDWVsD8MImCyGWy+Ox054yfmCcJEd1d9fWLRTewPMBFxPXDJIyCd
2MUfzv30ot2Jr3eTKhHsL0hiYQ7bUy7s1ogda0ZxJ7ZGMask9e0a32zC92/zV9m3ylP3qP+rWjkm
xX2jUEVgtTL+xQFv/e5249dLsYvJz7GtK5mzaJM848XlQuJ9W4eGOmslr0JXugadPgg2roFLH+Ce
jWbrWwEi067sCnizQXES1DIug2QsQ3jtaMR9Wc9nda42Rc4mNOQu/Z0FIcGvEdmiMyks5xyeseAI
C17xTFp3ZkGiCi/1elKaE22bWf8Ybrs2SlDKaPf2fMxC/v8JofEQzSpbt/Y9X6cg8L2836v21QuE
Qw3xEKsUumHnuDHtO4L7UDMZGnd+3CMtrFwMD0zLwf2B30A0HhQ6mtfVbZpaifTUv8D8GiI5txZE
2urAO8We/snKBrw7ZHRCoQSIglY+oPdW7IFa5L1Y1h8U/0ZR8umxNrsGi4iO7js23c/FvATSENGL
Vgjp/kqQDVOatMchJ8iPDHuY5PdkTmwPW//9bIrEy49kuzcH74Rk2unwjj4QHZZ+TtLthyyQ0+OS
WxhgyH24XiP6Y2XPjMvQT5QNU8x5b5HFZWL22yeUyU7eCauv2y+3KN9qrQtaVsNPXBvvPm8AaLFJ
944wJEi529UycuQKcUpDcjFpNMQjbah98QFuopk6PuDA2f+eDY+dxwvxNtmBOWksRskVoqfvgQJ9
5WsT/ZykB5Fchs7rgGC07vjleGpRL04D94upX6XXF82tIL7vqIqRftmIh2UA/legxVuIRC1YAfhi
uPfVWYLxqLoVOACqgcNg1ey6A0yXY3kkApjl3lC9L/kat7tgM9xlhUtt4u/6GX187wR3jQ/5HarD
/fGyB5DH3/XhaLSszbsae/hnTvHETFciJ2turwiPsUk/wqlPfs4UBgY3wvXgjfsRP7TzC08ba3Cf
SCIbpUuMGlFJsbzHhmGTzfDvjckr403F3vuQpEDfY+PITtKYd0Bealaa1bBELvhUkPJuiafWGgS7
JOmfSz00L5XheDXqr+bTfcu7n19uHi2UTljCE1VKUw/Iv1QAZ+a/EqBfsK7Dzw28Wv9FB2IEQrzM
Sq5z+BVEu6Qpk63uMzxaybc6nPGBdyvDnUDHcCCfNRRKR7tc5OYzr65pLJ5KnNF/X7iCN0mA6MBf
mAoP4dFbIVg/dkag00ynVxAdtVyJYWGJNBEBV+KnEcbt7CBuuLw5z7w3cESLUt8OzlnZBIxRHJkX
YNxrfhU73Ctmfi9oE9B68ui9Kqrd/giNNcq7b/EEi8xGlPqmAtJebDjKoSgLXMBxy8KmllXu/npj
rSdvaFFdPfBrfGyuBtRNm2yd01ceW7RgrHXVSFjohq8T0RF2IBKCeUzFITbcrvXfkB1I5cPXHZAb
V3zZB6IH8OZTxhiXPC7sPbt7El/d3GFx2VK6YOeMYBelpPjBEd+GSuLEMHVgZs0NwajML5eiPj7f
S5bHVXy7Zpf4x24fawDwLDBYRsOdExBdudJcg5cMEH/MPRjzXEjtWgs4HFPTaxKMeCURgVQAH5AI
DJt3NXSoos2sE6zsldHQokZ5Nj3Gi8VZ3lR6hUyHp26Bn0N7QfTNbk8RgjHTJaCKCn9yi3+gePAu
xp8bZGI5r1kwFbAvTgviLhcIZtf69NIXpRu91li6K0bzAzT5jc0JCh4GVnXrat/HwUZUGNNOaMHq
97MJD7UkacnUCth1avzZwCuMeXsz3s6c4biDRBxt6yau5KMiX4pUnsVrdRW5iD5imsAR5IW8vH9j
tedH6qbjdZlDFpaZjalWTwz6GWWXR72udKyLK7PTpAys5rNQLnCaDcSsf9ML6I0Im4klHK2K4ODy
wBk1p0cgFkLYP+y48UjGwkWDQbvh2GHdjB332yMov40oQUb/KoJ+JkYuJuciMq7L8MMaYVBKffq+
aXgbO6F8TumQPOv6LotTXNteJQEuMXkwETAzjnWOZrvL2iS9tFrPP2Esi4JvQgTaS6g7nbjKy7te
h5MkJ1a5jOR9e18tr5lStgQfmbzpkl/VvoVQqbWvt7n+7KJad9RJnA+1iUtiwRS2ckyn477eBWfX
vAVDWXvPgc5zQr3628rAy9XHrDNs7C/1ylokeJHo4mYUchPtYHuDZTa7hnDDJ2hCZlDDZRoKcKLj
/4W6WMn93HLDtCwQtYatmqi1FNHrbUCBTgjDqQ1LFnDs/x3fxUJtMrHDpIrpH8lkLAPBYUjLPYM9
zYwpW67O2mSE6QWllNvgbfqsyigsGsJFiTUHEFkbWAJcCoIw//Vgls6wLiv7wBWt9btXrbXuHelB
kR4zTzo42Ya7zv+S2Wv9aeEPrajQq15rhngGlSRMPqRiok6izOeraZL2kFx06ML5PEQkWpG954JD
NI16j/JHrY9c+I+/RIIDNz6UlvueUyU2AvtHWnhTzPzAPuRC1XJQm9NQ0KBF3bLx15CbuxJfYKNI
N29UzfyR08lfUotRjV7gPq2qJ9l+VGa1b7TN6KGAwVyPmo2WLU5DPfw/tT8R4avtdA972LaBV1K9
Mh0plhDkKzosKxjSmCAOJxRgZ2GyGYYBTYz0UCtc9GJSFhSPIcXKm6TOLxrNvZ1zsXtVW9P/Fa0e
728tYD02XxHlKlqPGVgnFAWoAp5XoAVHDi6Sxp9cOQffl5N1x/xwmWf8dYvKHiNbAy2R7/nyJ3bm
EoM7NDZuLYtp3hxEyXQfNj/tnCzM4MkyPyDG/iLT60YN7j0WdE3ps6bjqZtOm+mKJUzV7/1EttM9
lbeIEB9mHxBriAuOwttHj/Epd457dgwrPcncDNV625J+bCYEJeADwlQjnMARNZJ2HyopdK/4VvSv
4msnBlYg8+1kyoLVrojWMnpn75h1U0dLuP6He3240E1f2JLfXl+piEXgJuqBeIcWQXX68AU8UwAo
ooOyrcGkhsbCTPcfVhXa2iJSLinGrTwUQWHNr0yJHp93Q4WLw6P+CK+luReZHJY0gkcKCZWBCCRS
RbVKsyvB5Ajwpnv5ZsrOxnxF8ZDiIdypbRiN0qjCnJloWAPZq5XQhTD1nxsUp6PZF6bH0Xuil2PO
kZBsXL56v33RpSbewaCUbXMt9+/SNHfSWZMm0cDo5rLOfMYGLfoO2aUVosVf8gX7XvVW8FnLqZuZ
jTQtmzRNx3zLS09g6k7+ZYHLBsT2g4kFEEfUIZECu4DOZiYrK7VdXk0T+Q+7J198iQJ2UrMfn+00
JElyGlxG5w63yJkzaoFdU0lyjlvnLEzXR4AbJSjFngfNDRFc69a0PFXpBPsfv1SC7h15HU+x9esw
Vqn06OkkxcEV9sLyNLnvH7G6Z4HuL5zMnE6JIoMAyerSqIUXM2LPxndzqI32Rk+geuFrMTiNhIUG
x9DHRT2KvV8kenxvAaSHAS39iaKVGuC+EW+aILV3rbcdQLFrgZ+00Py5ZZngzyJI418Ms+Uy26UX
gn+7Rq5K/Mewb+cZczx3JgknStFjfMZgJV5W+5VezCk/Wu3mn8q9B3oy3W9h2pJEAxcgVCixQjOd
XBvdJtQ3gh3Whc4SmV6wJOqfrYrCaV8WckgIKRLBT6FS6DifEgpcwBYukkRqaMJtkhtdLFzcXwR8
qmo1Ku2vl9//kQ1/6D49rLz9sNLcLltWaTmiE2BMWWKuAoYK1Ul2i2t+S7h+NgkrJfoC9JcgOr5b
EpmGVkqQtJrCHkPc1SR6nXhtHNZnq1Nn4bl9po8/fsXbXmph98dLDhP9PMg/Xu1G4iYatX8zfwNA
MKmKHUoWOikJkiTRYflv9QoOnjYSmD227FTkSuedp+X49lwEMyRSsBQMnjskufi5IWEwYXQUCiX/
HITvYP60ZFUpt6S/DA8wA2y9LKWCoQbJgJgmbvwSDpMHvPw+ovYhvu2RvEZpNXVBHfYzCT0jgsJ6
qEW7HyQOgBxjSJKbLhSAL4Vd12vXeUcqeSNAgzq3HBD+EaCQq7qBmJ4CMQ8Tu5rtzGzCGNOvFfAM
7v5h7ZVel7ELxR4NiKkPr4XGhFumGCZHfr0uElkt0sOR4XUNd5mma5lOwWUIAsqP0X19t10jnZQk
HsIigZ4a7pKELtroUwC5/l/lnassVsjASPc4ylUq8vyPjqPvQdAUA/dmrqcWsGJsTSACxWcobk6C
jQ2ZW7vF/RtXqQSvAKju1En6LX4vYvfyi3Q0ntOgdZvmOfle41UKA9o7d+3QpWWS5oaS/2jfstNb
nONG4Y1YxfJ+Xrh6RcIUE9mMJSO4aO4Pr1mIbtB9Pae3HCweXcclLaUlDHdmvkpirrEzrbe7Q0hw
WZ75hmUH/aPSIC/0Hwo6Dr78vWwNZ70NGJamu4GSwFLo8lrrh2gpFIeCWfSusBL6THMJVIV/Ci9z
XIbJVGghUztIR1HQfdGJvAPDAsMWRMDn4wGV/JHw6ug1weHEyQV7+/y9GHxR5hjZcX90943tDfzE
EZ/b3NzLXfTQJ7VSGfLxCKpiTz8y61IYmxKsb4qpf+qADXJyJSAi3Xvt040XcvG00b8KrYItIcKg
sCxemBznuJ0/cgTY2XgLrpXw6v5ldZnfN73NSaXYpIxzS2MfmdujwB64hDtxFYiJQmvtwgQPNQcG
UzoERgvaH0H4KM55qGduv9K66Mi/U9ipzwfhAKkTOiUt/7EkypcQZE0vgl5DIdQC+MZX41KWBjII
Bh3wYFUtBYR7ICf0sY8+FNtNXpl3wzV4RHC2eqt0Sb39b2yk1rAH0PRi5Uw/06NeOp4gG+EIjoin
WbyU/Dx+4Fxzja+/rF7GElP/ZukoshcSgornYA7+IopfXhMb2ExscHKLYiHdz+QgBCotZWWO+yFA
VtFYSLVKyE3Dler2WkYhEEqzjRzjp4/r98HlA8gafZRrHHEq/vrCutLO+BEc8Rf9Qt/xF6uKcJg6
wex9sopwb/GXsSjydH1bL/gdM8iz+gU97mv7vyH4Um2qngIAB1VBiUbvtzRDO0nIkMsER7Ent7Sk
aZcIzs8LaDXrZyHUXVaU2EhgMGUueMI5YWeDfHcYp08/emPBga63xRskjhgiv0rNJPY/tZ0W9VQv
nlNBhq4sifHEo54v1Yxb9qe2fiG7bpFgx87T/2Ee51HhT2hxgM2zkrSQyTsLiyYBc09xTwEQM5KM
dAOOD/QHVFchOeHDiVG06hDh1AKGhdKoPGUXK+Xi6wtzVqLLdUiLQuJ+jXeMfnJUjSAggjBzwmts
TprBCDnrKkb4pp1pqM3IiXYEKJ9lfWRucfz1O0qhZZETKELr64LPhd6EkloBoN/zAg9GBw6az5Zz
lGbR7uFlgbP9nvLvSYtXvFMIaYIknvDu0Bs5BOIcBuXZ2JYPPuZZpdYOw1QlMoSdIDtgcTxZ0lWs
DJsrS9KSFGSvzJUhSmqmdIZkiX5WMwol9nZhLpUS1MTaCJP25BkyANf26QjtB/0sR7boyaKOHR8+
MDV+WV0n1qZV0jheAWAloOveeAWpHdWOZ9EG2N/5d7Ocywb+yZH8PfZ97hscUzayNrEsyB5g1OKv
EeiC9HTEHtSqo/o4ud0K4IFEexoit4A2av1zZo9TiV0K7dn6aNeSGc7YDNoLm+Hc8F+lFzTtrQTI
324472kKFurQlUGdWY79GmPNRGD0n6AR9vZI347H390EoVLMbkoj1uoxcOhlaTJ9ALdl8bGJKgB2
6oQLG+jWmP5V7yVk7Iv5drIf3AD9nHDySwwIuT2y/fE3J+hZ/q6zCz09mhoZkuUweDMCZFVnp+L5
7owkkpf3+SPrTA4fmTzIqOhFD1c7tkRbIwLXbqXukgD8A4Cwom6bH3iL2YP40yb6fQGGKNZiwRKf
AutQTBOT1oG5fEFBNty4FRe9znyWP2WLI0M0rYhmRjXTc0L+P8z7Qzl07PP+SusXP17l4atkuEwg
0KOxf519fpy/BBUqa7l64vyo3/DLOVclYFPz3SK3ss/3Hi9sKS6CZtgBky2bJUkeDVLd93lGYfpf
2z+RkSZFJtTxXRUSTfO7tL5AW1oxtUYMOM2Z1yqI3VzQUj5UQlwnlLLGPJjQc9l0yqsBsnf1FIBk
LaQ7bXO37+LMY9N4kbJdaGYhLUl/Ky2hOktqM7QeC5QRyPcjV/CnhIkmuahE3Kbt47kcw2/x0Hvd
82wkACSLpG4Z2nhiGqdAPW5n1g7nFCKOtKAhfaZXxQhzyfA+9eQdWvg1zUnEUgaYulJp5L/VW8MC
rbTyBofnowNnE1FKKQn+Sq6kHy0XJL6B1k4wst5DMEv2cMyYedWuLVntdjq5/d4udr7NdljuPcZX
sxwpe0Pq0YwFEXAcfp1YDbavn23/EYavFrOSqg+mJFLy65fdOLkroaYq4WZtPjhI7LGqeOK9aTTO
dM6YNSPkFxt0XVOEuWyzJk8OK2JtdQVucmX4cph5L84P7glKZMr5zGmsYGZc++sbkQFe71+l2E0q
QjNXPZoD+6x8cMCJpibvT6L7AnCQuQHQ/BhopSWvu9t/xw32H/F3JwAFDRxUDE/xfBowD0pCj2D/
a/AHnjo5fVGudG5xUfB/Uieswci3l+mbbxoziv0ONBtcPpCo5BUBs64r7NWOoqYoHVTIDrlQ3gqe
JmJPfdMc4JNjCha88cQwE/b+IOEYADQ3abn2BlzLNiDwTjzmluavVGj5gKWoQ01spcplfVYcqC+L
FvCk+S3BOPOFdAvpXKTZapjGP4tvVE3VKSCDSLAvp2ygNLiaMyYO354Yl7koXRoem2S1pSiXhy5l
GA89OXTDMohEa3j567v+TP5dejzPkyUoNHDnVJ4GdrMHDczRlE1r1z/xGjSh1+DjR9zLVsSwF5th
F/GRSs+AVk0uCxmL7RvegdFDFVeO8v8sZrnGx+QoojiFV49X0oC4bqnruhhTQOoQaV9OGEk58C1t
C5I1sIPYQyyTdprW4HoqXsvyXygnWwyncLmXjmytegtjRkYiej00nKsNhfr5rldDu1KdKsRum1mX
G67pTMcLULQ7OMRzJSaRdFGhS/HhVX193GHEHnh2tZhU5ZgKasUkP862lTYH0qthlGuQGlO1tz0R
y290UKWl2xlbV1YUqgYowhUGJVkAN/G9b7Vgdlriq9MPB21mJgH9L9MwW4Pg3kqNjEJciF9WOwOp
gj4fM9ZvyERp16E8JjHmAJd5Teq/kRZuE7BkUADUDym894jOdCXM7nyvz7SSqiGCE5rmBbFVn6sv
JJbxpNi3Ic5GgwcvMAwBUDyIUO42Zb1P5HUc0yAfGFRW8WnRWyYzXrhbG1uKOwZkqpqAK3ciBMcz
7Wr93HHbKsCYlETFd7/NuySN++EIg23vcydsJnYsmH1tqC+qi+FzhmJLu8r1HnpRho8gPpX0T4ul
0W/55fY8hmvG1JSOrLvjpwtIBU5xDrh020PVUYw8h+ZSnu29jM2SHSELcZMEoNjCsGR9FLGumz6d
nwKNGc8+3iDMRD47aBysZmj/eaiCoEbmbhgzOd5tG/yXbx4HRDkDjQVwHLvo1+9Vs76NjPPxJRFY
1THVokA4ZQz6UBDgNGRd/7ImfqCOkelOYXogwK0F4DOj7QPncHd1gcW70GoCfYybGhmXie6JSZea
fuFFPJ7yVFpYUJA8pJsxxkGNT9RmZq+Wb5ew7N4WcDwWZxV9RdUMYOqjfnhwnrQ/8a8pnJqMgMUZ
hESRtBQK3RnXn+x+MnNaEn4viG7zJx4wGffeuzHjYv+NRN+Lm3zUeOFR4Qg0NiMUUh+EIWEyQylF
XT0w1a9CzhukXBaQymjqTHxm4hmi0Kr3gr9k+WNbBH7Qng3sS5bOuYMEv+euRYuj+35QePOMHHfq
H0+YrmFTDUFHP9jy6PHXAAtctmHhmAFfc6XU8x8KHw/GfTGicf6mMVHHgLv768BKG8CfRCEQC8et
GsWsKOMYkQBhp3ol0lNlAPXF4vr51FGXIc3NC3aKpjeieByr8s11uJmrW6Z0ZdOvzWXIqYP9kzOV
wDqvLlayNKEtAQftcD/5f0cprlbVFuw++FjmlzvC5DocX1UkjexTFxjL+j+YEIwuT426zB0Oi/mw
PslpFJKL/8P9wHKtsYXTo6NnV69DDgtuJ0V76djt9sYZvvxgB8VcKQyc78N2F5sup/nSPafcL4Sr
B++GU8QmbNg/yK37SaYVe2crV7PNUh+OYeKyzj2zel0ujsVKLtuIs/zEk86oZVo9CgKOUFBT5jC3
UF1qblqMyzj7Ks2i6Sj5dvkGyoj6MzfI43euGVhgW/5GAr56IxIAjsDaeB3KxzSU5Xy56mtPn60T
U8znHg5LwNoK87+n45gJsS818XbGA9/roeikP/n6EQBnesejLR4aFIim3fcnigVFHvKSTyFXwdBO
SrZYjOy0bEtlskafy5lFgJM6S94TWU251FWJgnAyDg8bgmcUPfwaLh0tNLNYnX5hS4xqACWcU/25
+4rkLg/AuD67zQKbtoi4dAeySj/woImrhv9+b7OcBzAqeC4BjT+FCMusGYWiFSh8LzTnH/08hfuV
uwoPnf0gPg+P2D0X8l3+L628rHhDeclkJi9W2ute9+pqKXNJqcE1M7mY2Mp2nWLR7+1fpDn3SOeN
VIrPnk0Z2DDEwzmtJwBgxRrwFQpZVOcFU+Qch9kOv5MbxWwg1AnyG2/SiHZ+N8BaBV7n9Ggx51r6
n9rR3F6z+kBkG/8B0ToTf/F0utmjrP/5uRtthYlvrdDBC7+miWmaAzO+AiwXp2I4dhlhsbWwpgyT
dENFU57bd/ot7zz7HFOmo0ICVs7Bc9zFkg4tlKlKgE577JRBYL3qJIA7jJ6P9oszT4kJc5shLrs3
/txFQQYDND6mKGAhVr99iyT5sjMoYnD2pbVtPARvKntqhiJXP9ad9Prj/OLT5TJcjIQAlFGa4jKl
NBnhwwryI2xkN9UNKiDaAvyXMSHOkjs3H+GrySba3l7jAM1RuBqXxvNUxkKsxjqT7PAVHAhiI0cA
A2y8n2HukMY/MBLID/lcdsjsJVdMWL/lg9SsvoBO0+AEDlrFoYUG0u7Vglii7ellSQ7lTj+vv+wC
o4jMB2JpSxeMCJrG244NcbHptwBaLtFzFeIuAA1yU8rjc/bKZcBv3OD1yGIwEN7Vkl1l4RSm0b7M
slAw4IYtzpbseHDvL/Gpb/nnf3SrKDo5UGiCCOOXv1cv6kNIiGsBjuDVQay10GB5l4qOyYNQUnUy
O1/Z1X+s1e9N9ko4bkP4MGpoIr87FvRj2HGobg8F5UE6pCBlLQ7S0zdZehtW4K36avBsaDxG12Yi
w36570hK3UwReSrBssNg2Ip0ykqaV5LqedIeF5qN/u0oCMEFVCiQOqFT158JOYligSrZ+3ETutpl
UK4s4lbJlzlPpLvlIZsJDsR6mCSFlwiD2zYSIxVbMbYHvhccBx69DfOLA2xrp9IM3H+T0MXYt/Ms
/b+Rv17v5tmRfdJLV72yC1FIth2WzdRTMtU/6ob8G93XRTCS0aAp9ISMzdAQYc4b4jVsfjB7nBWw
hw63RfNtYk3rBXoDss/rFIB7UT4P5EAp8EE/FpI0/mxkcYdfI4iEPK5FVCM1SHtvibcmAhMdiFPn
JO8X3x0iTGOmcER9IWgVcvmR2k/+V/cyAWsPgdf+ozG4aLHCursAde8VvsZLEe2Y1t+zJctLzGB8
PQfeF9rOrgnjh7EzSzWCblzBrVimdQtL+B9TUFy6J6hDAqQI+Sl6f87PGJvUcdfPbVubgA0FElrR
HW4WUNNOOZbJraQCinvS973ohLz4SGXOK0ZWEIKeR4owxYoCrux3dL+FIN4SStXhN3PnzRUPYwaE
uDXKXOVXcDoEj7PsLclfhwSgcrS/itEpXOKQ95ilIMvB9aJRIuagqro3CeMXQSnx5a2ccqsH7pSI
Pve6sfjflnaQFL2knKsjZQQv+s5ukCyNrs5aDu2xmWvn1IYCIWI1pa8LGnpF0hvbVZRi4G2DypE2
0ZhkhW3TizhWGKC12o2riH4usZWotfvSN0iLXBb5qNkmzdcl9qMU1D7xCBgH2kY8oR1dg8LqnPjW
pGTjF1Rd71vfdeWbFFiUAyJx4tCjq128sa0YZPkqtjDd6xJvryhpqCd/bPe63W6vt98sO87gbvIc
/QllaBT6DvPbM8Egzii+hhiwvoL9+4Vjah08Y2t0tAH47fOGdiyyfwugQLp1iYvr2S59+OOviBse
qxwiCugw6JXWGbUi9bsfFcUY04xvjHDNU/KxZFXe8Bii5/XIVRpgK31Ugou3HXJgcsBAVBvrX8pU
DelXHihpXQpZ40lt6hqKUubUMVvFUdTLhh0KOiCi3T0aRhU6EjYuxzU0oVowyKZBLPDG0/gGbPYd
e+UbVQH6j77BkiP3bhYxPsnmInS4cUTFDQdoH811mnxh42rn00pZHow61csVbK/N/ApNQALhr35w
5R7RY8JGQfMSC/kp+NWxLNhzvP9pCit+rf5h75Wm6l5UEqGDWMSu5EOn+fyhng9soFDF0ApXMZ8w
QRF0/w4cmPX1cMd0D1+ZiZJqc89FXodNM5B8qLb9+n0da3Jy+lJNYZkh6FXETT+gYsYoV8Fxp51+
QNTUMnk954jRblBYhOVCm9xbdxUlvmYOx+QWzOzzh86dK559cVdVm85wq4ax9LrwLnZyY7mlk9k6
sP+L+vJZZ9iA9iiXUUr0yO97GXeRqQ2hf4ScA13R/mJ/toSZylbHj03PYo+JehLVwhy136tb96FB
KWM0Bz3omnDWx/UMkHNN3PziGedEyziCHKcgbaYnOY5ummr7o4m2qm6OmKA8Au2FoffX5vuZR1dX
lIi6K04cayWhQeFcwYPPYPe4kqxcQLqtKq5cutaxN2d6IiGH0PATqOgauU4nR7XluEUJjw5RF9pb
3hDPYx377vZO/S9A4iAhjH21zECc9QNrzAdv2f++wz2O9VT/IV/SUv2zIuStX+EEWqltnOrR+v/l
kT27AhybLRolyRKVUeiuloe3NTu/iwMGMVbQ3jWJn72A3lD6N7OLAArYGGKoI2xPoq8JyXVVfrjb
YuZiZC9exi242HTgEh8YlKS814gBYB4YelnWQqvAK3MgNkMzXryMqy7EcuNjZAh9eMJOFZzkMVhd
HandeOdlWsWyCXfI9x0gUHLzastZ1MaHEYnSXOnC+Vxl613YXJ4OLdH1IW1U0hfzoDJkC9/+E8nB
pfx7N9yi6IVIfnCHo2Ke9QvZiqAVq1B7oo9GSzB3yQAeQp3GjF+66qGuUh6ZVDw9D4gvcaiYyr9R
3c68vrO/HwVbq3S4x0r6hT3NM/t8cY/6z5G+p+PXFL+GqpmnRDFkXffvLz/QSTWetOKj5ULiSGbB
go4GJDnMCau2d4B55ROozklbS0EDFJYpZsVMM3TBtO24f91Oe55qAVfoGQdM+wuA1WLKz5Yr9lqX
trPXH0IdOJ9lHbscORmnP3s+jKIMS6/689RJHZePB/4URg4hn1MNF9zsWEkcSyUpyyZU/i/4rNLB
ssshvkJ161VDcMAY3OPZQJ2I6lyJ926QC3uGP+MvFbQYQCgW/J8GPhQqDOlzmAEruzuDtDLxwWek
fGifPH84lbYz0fQ5SUxIazrWQ7QrGtusX80GBCpLFe/agTF5Dtyh8yfIllYApUz5tZAiLctUCHDZ
r0Eq/HXyqnUROpuWdl7LjOvIQPBanmhSv7WN1kfb7IYAkJP6dbwpL0GxWARQX0Jk39z/Qj3tQf6j
xxLwKmmhyZzV1EUBiRg9gooDP6H9xLgbD2JpCrIzM0yiCXVCA2mdFlIcnDACCj3+/dZI6WuQE0kA
5MBOMCcv+schZ8l2Soo/kqOHw7oYswbRoEdrVuELoID1ZG+eIus8V4eETqJSsAXbAQrUmTLMUoMj
A+K9TfO0oIYsFhnudy6sWnVUD6lw/Klq0eh4N6MqVcqtvfIZPVCSsbh9FsGwHX053bWqOpjt4TSM
sxRCCLO9AjXo3cAfhMElsJbOCoJ4D6RFSxtFMaQQK86Gk7MEiLRh2Wg/du1Wpu0b+Fx5H6QJfGWD
xULQu5LI1NmFfyXAiagCKhJmymR+FNHFRizUE3vX/SS4CfPmHlMDaXIPvOHGL0smfMsT3ctNyLTc
sM8aV9DMSjHyNUa6TGQPEmQ3pM+5xTw6+Qo6s6wEy2hfz7ZEJYbVf9j6jLOkYETjGgg4ngCiixkz
tlwobWuU4El5Sp67JWq6sEoHtRSP2/6a8h0AK2ERZLTLS81Pe7uH1oDefG+NdqFZWxGOFmGv5Vpr
NyYSXNgr5moAfdAm8nlhn2TfpoCcxyRs082V9HViPOGTXvywtNCTjxU2zqY8aPXnMKi8VCaFL1ui
DgL/B46nk7amsbkPVDE17gpcQ5vcmAC0hvIf0WVjd2ny1fkljsVYCcQWr71NKAJUY0frxhqy1acC
qLc+oxVzVVZgGJ5GcRb4h5hsuoZMllkEpmy+Max4TjxZkulaPuObwJmyGbgEhCuIjATNFVShct7J
32lS9iWeTmlO4uFOigNj4q/oP1eiRDLobkmYuxD6QFxs1vOGVGARBiGjRSjXbWlgtMAcQchZ3qYg
gF4tQexQE/y+5FT2fLNngO9eZLwcgT61Jhtlzhj7ViOzV9z7fSz+PelmrHcUJSwK71NX1EsVAEpG
hfkUMCBQBDGn9H9f6yqwmWW0/ClqBRYK1syEeFgkYLLcht/fP7u3WSq9wb6R7Ad+wBdHivUw5lEW
YUKusjSl87Qw3hLloCqaPd3UI1BoV1SU9T2u5e4+APW9PN/YWq2SsjqeKFWd51kcgeTkIqTGFo1p
XCsD8EGQfmaMdwKfbHIt63ADHx5iUFJbmP9bEMe//Ev2EOiZNzYot0rfEakpE019voKYwThXCmqa
UsIWMBSsoTw2GT1wxcXEZTDLVPhnfo6Y8Ythk4aDRIOJxoLf/FiraJ+KfovZ6DsP83aMshE4LJL6
CWOjGj0hneUbpE5sIij5z3nQq//HNLAUxtRz9kAJzmqliw3zYvY8A0mQ6QKpeJkFu3gOc8dACaJk
v/Ncm7mn6jgcZvpnxegNsfPrJh2ZJqiJ4mY68VP4sfqceCxjmyQllo1mmMupgP52PYUtEJmw3IEq
tG9yiCJOhKJCaVex/18+XFxhDTpLDydi1pRf1yJiw0EmrtM8XHdCqPHxRfa7cGKperf6eoZ7TFtO
Vy8l6NmS0alesbmwsluskpkZlF8DEu7vh0w5ZfK0hsPSI0Gj/XdrVY6FNkOT/xSXObc8RnNo75LG
aMV5WQE6lAxp/hc91xk49x3CyO+XQXzND1kF6RkBefEHO3MNsrog+svjEkrvUSYVvWnpDbNjvK93
5fMARqiXn4ktv/85/UBTlrT59WJCzCQeB1CtID0DMEF3LlBTCpIvY71DFNWY5X8dUdRYZp2dfo9E
W6Vng2InlfTB8JUw5ne8Ar9NIrYKt5iPAGFBgaLsKnDaU1ImnhLoAlyDDy21XteGB8wZ4lyBh3o2
QAV7wRRxr+IHvksCtWvlSRl+z4o4a6EwQoQULQR8vaDxre7mkYn+plski6D86cwpnnQiz2MkLtAX
QjdTUq+TGCYiqCPPLrP8FghbCEEkOv44KAY1ajlBb/ErefMJibsm3ox9dnAzQ7cJZj/Poo9LdQGX
5VfCobo512pOfw2E6WcSrcIxBzmu2kOdh3U9TzcSN6pLFS/S3Wkl1RyG6EN7i4whkhdA+hol/sL4
ePiKk4r6wFWbVJpru7D6SGwpmRMXcVDvECptXJHoR6xedYJPnAzgAOV9x7+L77ew7XKUv/92CTzE
4IBM1PZ4Mj9cK72ihMzo+FkKDM9SewCspdlnE3fAVlfK8twmUtDA56yqsH+POxi7rQp5i/Ni6PII
/pEuEQPWVUuzBD4KgCWi79uQKc2hp/N5HZ3b30XOY9Hl1zZyMg2wZgVjWUmhgkeeZqVLyu7ck4b6
WCFucUblpDt7NzBooy25QNG3ccx2pHnk1SDJWdqPhPRYnBf0pOPsEfpK5409kVkP/dMlT/qAxFnZ
h/QvLbxGcIUKS1CjL1nPwKZKJviScnXpw9Wi/1jLgKDZpy22tVSkFIUGradap2ZGhorfVSbVKZY8
2EzCuoK/kEnAUkuztJsMFp3Tw5Iane27MGwThmFFzHa6tSUv8yLQNhsvlaYnuHZsRD64LFz/tJJs
O43gQAlnvkcaoKt14UtF6kwR5s/WRV+NYhKBhtgrK2iDMrXTVwxHiB2iqv1frPFnRXm3xtRVKZeU
XLmNf/czX/owfiN7kGOXWv9M/xoj2A8XZm/AkshOfWGMwY6LLsx5dFeOynedkqlkjI/2Jb0tr5qE
hE5oWHYnLUTmmNG54vvEk+bFPbRDHe4m3L91fvo5cjk2AuDJfsVgnP3WfJwZsKMnlpM13vG/zGnu
v/qk+xQVgKttyNeXatm+ZSv+lA+1qx+Ofx46iBama8YQkH5Uan4la2ReVqB0Rn/CiyU8jpiBvdhT
n1Qc2Rn+ly7rSq9Hl2kg1kU69ITQCWMwppnW2irjlqx/wAyWJK5W1hPVQsON/eHvL+Xq7g0PIiF8
p9fXNtZeOojv2+vhCJ4HQeG+JqWoB3QMltZ1hcuVtKoJSAsdEj/LMXa/8jCo854nh3BeyYC199vI
a1XQYY7S+H3n/5jur/geY7tNOEuGCKTpqnlVqrWnB2lgGc9NZOlPl1Y1eUdD0oSU5JgmAjM8kCUl
sob2sr9vM6JxtxDtGPJZJqq2s9IfeU9H94ZrWt3OznJBeKOPqk651GZkbhLtV8QixDWUw0C7VgzL
OyfpdILcHJAKugWgqO3AGI/KdTH1NWeyrEFkJ/VkKqSrPSiibTnHU7IkkcuzLMV4SVMADtCmk6Zk
H/N6uE6wOS870RnXJyaRI3jI8l14j14e6PcN6HnjuWXLl4320nOvoMW6JWrRwkCZZTTpPnfHC1j6
iXG5C9neTA8HXI2BoLbjc7P/IO0o5WW2Tta3pqaCQhgucL+hEHAqSHunGnr4yHnPRqsR+1VpJ/Rd
zaeTCtdtRDzhO2R22nni8JHel2KqVBLcd8kSiMautzep1xZE1O/5ov2wNUrvaVQVKoCq1SaNp5JQ
V3rTflqcVUrpdfsT1M7uJWQRnRE9wUSVuSzT/E9mRA70yvWN3Zz0hS9vvpk4Ncqiwsb0yWtlaKQe
47mUpP+k+5xW71Bga/ywbaNp4VDdf/HxawDOHfuDLTqb1UpSb3Nq7falQHEYdWeH4m2niQNdTlJJ
+3Mxg694p0UEebOU3mydxeH0jbdKF0Ejc/rKvGim+HVzGT+5j9X2TxQTYFc++PvDNhokV12A8aUA
H2HwumlS2A6K0CdPivlNWAZ4r5RwdI6rNx2Re+/r5bsFtKTbul80JlYhQpQhMQYWxG5LUMMD/HAJ
I7+KadpO+K9Zyra5im0pyy613K43WD1QjJw8HBESak14Hm0UudVvJKpDrYucUogNgsF5GSDDU988
XISSSMNwCcJRz7XMonxSYk/jH0bMUApq39TC+pzA+60M0cFx+m7nHuYow1sOJVwbV2Qcfhsklo9J
wOpbpOsh8CW9/+hlnLDB11PrCzyaCqnK1oKO3UTb37JQ3neoEgyz52mTykoq1nj3z0E4i6CQo7ll
uMElqO7QbsNSCCeNjbUQHvcSot6alml6cJ+oOdlTw61RRJ7ep4SZBxukyShHh1YAdhb42ZOoQpLj
KfhtPva7Cw2ikQh4DWxFgGSblfrfZCYNEkVhRhZKxLMK4DUwrw7Ng2LiKyBBC0oELtEN1YsupZFD
UeTDZ1Iz1bNRlw1vZKaacrQEZnsSYPwPCDcXe9qEvgAWbkHeyDIzEN1l0uT1ZdGs+WTyqSFrXQNR
tE7p2/wl8eGelwfVyb/HQLWP9v6X4uLkfRnpFrvlVudiVMRMsNFIkRjwbhgDnfdUpMxINvMAEyhB
SuQC+r9d2xw9x7tPOSgMbSDxakg4+/8UsOlieSl82V65tFCqyZQexmoDPDXSUJRQbD9lxHgZaea4
R/U9+QhVTlozs7eYC6T5StmTqtKTvBZh7yi4FO4TaVL6dcEygbRunXliS16JoJOtGDuAjRvHqYV5
nXd7q40k7kKSixub5+vn6BeFWo9bveYIojyO/mlRUrS41mz/hmVNNqMv+I5y4Tn68hLYGJ2tHhYW
qngd7tX84ekvedgjON9bgXVfyiMh2cpkWinmYHkSx1UiDbtu09Lh2ygjUaixzQIPyRt4mC76oD0X
5YpnIzNy4Avm0TOwt3tukX1KZ75+YQquLzY1n5McbiOJ6gAzr7l4PknAaL/WzFw6jH9dfAbSb12K
UtDrJdn6uNr5LdtUdwe/ORMcMrOf8g1XOKEWwLV/eR4xCnD3nAGQ+Gs+v9xgFMNNZEd50MLLtpMJ
nrd/Pvz2jfj3F+NxOTiq2c8l82rHibqkBiDjcEL67HZMltQGQ83COUtURP6xTgpu7Ka3T0PrxJNS
UaIixOdfHbjcDWWCz9fNSBHn8bj/HRO5etXwf9g/Q4JPGwjfTmRtohnUYUa46fYKLvZ2u//lafQ8
yvCmHktzgMdtDPvN588mvT1Jc3jhSKt08NeQd8cn20n13EIR5w8SEf9eWFNmLKHXgK20JtGPr91f
blupDsXlDo/gWfWLOySg+IkNrtoS8iMQPGi6NsGVNgzv9Zhu/kCVg5yDveJqOwdGENAI4/gXpMTK
4Aztiqkii6POlu8nKeWDShiQCkIILNjYur0Fm79f1SJIp/rEp3+fSfq/Fhnj2g38SAc9fhP79ap2
BVDBz+MXBf5VZj8PZ5hAROdAFJioFn/F1EliCVQvKGF5kRLRSdgAtTA6vYQ244jBM0tfWjNUuWOS
N4IYEjmfmK8hEWcStYkBUP33U27Pl/gCDbDvgkI9S6eJT5mvym4RiNvIhudHbmEA2efnGxESs0W6
AyqGviTppX0nZZH39X/LCW/wp9lbN3Y/H4/xX1VwjeL2UC3ENIZb9lejMxOUM0eBoyLWgocy14QI
wSnTW+lSeZ1uUmJnTaakMLj3kmrnhMMVzH0RCpW5/O8tBH3ATTG2FLdySsLcwWuepiN8+N5mKTMB
lzEArV9HeJAmZfrQdn2HvQz2H2fminWOSvKR/KJ4tt7yjAqdvlkON9o1c2FITZf/xdyRNdlEk1qY
IKzHTMyyw5Fjin6RQGb8dodOQdiHDu8oyyx0wMsKMhjIX6wDjU2EkURPixb6U4YoQCmpBJZRxoD0
W95IZf0CyeXDUNH6R55O5WdCohtHmDZiH41jTp1zE7b7V4Amq4GzfBDuCgjP4l6rrlfxCJyD37/5
DPvR1IP3fReGtJ1GPZAz3Sx+K6La4OFQaPt9Ot5lGbYa0oxU2PzmjfDGBJbv0Zii7IJnSx7sTJDG
YqPi/RCcm3mGLpMaKlA2lTJz/kh/LUGfJYz11nGTS3LrkgMgHWjS2KGnypJLeIrreYskappYNOZX
Rg7gInFGiDOboWAkW2Wouc96garsOgMz9jrMfbTvgH+gpjdm2sAAbvHZeAmFe0aPyh5h5HqC7uYd
qeaEbHW9Lym2nN5adzrdYqRu+HHqglE3uQdqY2Ue7wEYu3aUunDCxDzOa5ptcQ0Cwzsib3Hik8+K
mx9RPWiIA2jba5Xj410tlo2SwYaaqVR3Uh5NeJ0BZ7hzi/EsMhZfeBko2omWAhNA5fPtzWzazXg2
GloWMs607fvVYe4QQjHjtMwYCEktFr9gAKr6nzWpAoLutnp1CoLOzfheZKEHy9Ol1JZFoJOWx8Ed
Y0w2D1HGOyoKee0Lymygwt3MTDr24l1r4wRI2R0ydI0W2IYqGLyU/Fof3UAXOapcAQKG3YvJPnqJ
3askekD+FOf5iEL8slTMGLf2RjA12syPZpYThGnh0d3Y0qU9b3UxGxueI9tS9gd0w/xGGLf3V5iS
YA7TSOXa/8+PhhiVlYb40tkCKUvj2By5Apy3RvfUFBEl/wlZs0/KAh0aP46CymOqhDCN/4i6AqLm
X3E2P88wjbHtlfy4B1J6vHZnSIHEe95RBmaFDO7tZw+DHrFC4q3Biwu+SES2YlYndVwI+jE7F7A2
0xHJPRZeiqse5XruI5AQc52dcXGsjvKVN+L+E62wHpUWSmWDDM6h3XIIcNUKT5JrZJWmDch3t7AZ
3bD5xMzA0fli7D9D8ULnN6Eu/SrqPoekKUB+VtGaAyVBEnXH7J0NodCG06gYfg1CBDX1I+c1IoA+
T2IOpFdcHS40SbtWxCKPyUHkpqo7jQqtoeGinLH71/EgbN+U4DYLlnubFxtjHKEfyN5wE5PoCLcy
2jpXhTkagNppp5ox/G+zwxet6+w8VcuyLAE118jA7xfohZQy4F0iHNQIHuEToC1GPVtSyln13EyN
7UkpDT/5bAhO1Pire75Dlb+WVEa7mLNtOlOXkt0vC6FNwP7D5MrLZqCdf/SANI2ydJ+wggAAKrVH
TWPLjUWIn67m3+j+OONKHTqWdlww/zjhcCIJr0oKU3HmD0EPedcsa1lHuxckWDNq74WmR0QppWYH
NszMuSqDK2Mn9ifVz9xO1CNAxTQarY9bFuwdLh99a/HNZIxZpQ4oQj9ZdQMRyZiJ+IVbS6+2OW16
Chy/QtYyLzWjoi95j4Zg7XCgOPLx8UT5FLYvocvx+j8oPmgZ9VxmfH8q88MGuC4Qt7c2kSfB4Bt4
IO8xBqxpu/f0PyI9yk3NEHkVjj3q274ejoH/+Fc6vBBZ56TRQTMPzaIeac9+e4RZ2srtSGX93rvw
yUGMZTY+tfXgVZljDbdzZX9d01S9nDY9JP1m65J0F3HV5H7Q91v3iCTbVyRP51qItO8o3VFYLNbz
ASn9FLtZ3K6DqzbnL9hn/LtMS+jPJdN2L8/meZu4C2PyKRZQyu2ybAYHWxQBrbqBwlqq1/ZXw3vE
UOVb9EAcKpDd92wk0Sbpo0DxSFJGSBjL8SHTOlF7sRPx0XuMZxvucSMUr7vXvpcAcVjd1WKX/VbU
qZkGBUTXNTXup31yKEuG8k4SnVYgjtJ2x3HA9+4Z6YIkWVDC01+PvPK5jh5cV2MbzZFdf7Mxi/Xt
L73TOIgHuW5IlyLWGwMmISb0qwdc1OGg2XKjz5wkTerR2o68u17z7eNJ75tAROMBDhOfjL43LyTK
C6YSnzBFSuVZ2Ccvw6OEVM97TTCYJYoMw5vwU3YBWFNt/KKW0PIGrCSqtnQO7c7E633i2BNmjSve
mKE9ZO35DFGKd7U6o/l5rDUkKUTL2KXpiVj4BOkp7czBwFnb7x7Y/CAcGUv/6VKaGh3BlhA8K8GG
jyqd5rjrWZk1AFhV1VgYmrzNRKudO0FLm064t0qe4Aa8BD3fFLz6PMs/Z2Za30+QOk3yR07EStKT
AvwI5shZA8olOGAL4EdS779eGmLRvJdt1Y1SBUik3TqvcT+aJHyFJ6/QYjeZFfaDzMnrlAwbrtkj
ec0PD2oLhgh4i1NJlf66EHZ6i3jtLTN1J+WATmAnTBTLg3xiH5wuMLIu2df9L524yrQLxBmi+nOe
Qa816AK4I6Uk2JqHOS9PADRYaRHZdvyo1Q85NQ/cfrDGJ9JNFGqvWpH5jr1S7GlaURqqa8hU2W1n
I7WhUNp2DiC7tL0qssiwVq3BWHDmE4wifJr9Ygk+aLkLEiwefnv3AfHPB8fyK4n3yjW9SGfUWkRu
s/lFpOp2Yp6asD07XLZ/YoCkWV/J7S5W1lJALMtY7nw12RicVlyrePfyqjto4x1iQccmrZL3/kju
6+c5iceBZexVPkN0VOQl6E8dra+RAhaO17u5+C+kONmoAKVZRD5202HUSuH3ma4kRnyGNi0BCzOl
hyBfKvTUSznfJIcW5PPEfMEcHr5ScSdwx0ivCxjaSqfMME5L8cJ86TL0CRUMMi81xT5eMxMd6869
/3t7Ki5rj0SvilTrIFTW6mtcmCYAgPFgadLo6rD3oH5LJNHa6TuoxRxQMm5VV6KwjCuUjNeBN4DV
cs7OtlwbOoWJyBoqes5jTjgk6ASXHPRagC0oFdYNQjJS5w6Bhll8cTuHn1KG1nlWEZ6OOJ44uDkb
W8tL5OlSPAsAhjj5h+dhnqNmlN4HA09Lyk7a/wpi87TaOKDmB+k0e/qelymYkVWQ+qJ72ScMajFn
wjfkTXqyfmSy3Ccxn61g3beKUFK19XXqrBIOW01/jQOZpxb6gbyHKnnJYdnl1cj06Tw4TL+f6mkr
awvlBkb0uXVtwejmZLqb6EISIEuv2WEbUdLP3PZtDwo78RwgK3v965HyAWu24eIR9bYlsjbLZS/C
+4ML89b1RLbTQPTecoH6IYonv27cPV7mgClZ/HVmL8PtddgWeuZQaOBRrWy8z8ajwgdEnsJ0V25k
f2Fsz9VmNWXyYnjT9ZKj0VQIMqs6xSaBmlgy3+77rOPPgOk+9mJWpBO+Q5kT3W7EtvJeLlkKhmsl
FCAkJ8anCVzyzumOJ0sCTLR1g+fA6yhdG1PnzCltT2dt1ZKcKb7FbQDvgt6LsIz7yxM6MFqgVBsS
LJlBUbja3nefmnsRWCt6WZ1xvVHiXLipmj42OfZxKHUy7LdVb5oz8mk0S7aXLO/kFC/oibwqZ5JL
WQ+tHJ6A8Vsj++JLtjJYUbk7HXGveUGQMiPk1euMu/DQRc/2NTyunt4a+sdL4r94iBgHG9QTA2+l
zWqLkM35BlwagAkNCIJljqoS5rVrbhd7MRX1K0HhkCoWcyUZftyvHxJvDl+xnLc1Z7v+DAfBhvyc
KzkBfXG/6/rbi8RCkgVygaU7bleUopJbi9WzFJHtdZzg8C/BHnS5amyxNN4akyRdQErPnrd6K8b8
4ijanUV/oFAMnxqWf81VjnEYo34bMiQUouxO8u6FKZ5Lb9Q36kc7MKXQaWoyW3xy/T2GskpdJXZc
qhi/psjziXrVdNxJBDSHtIPKxniqeQ8Re9VswI1/gCctPA57aXvkRpcpUbIm6QnaqUNiyYmvN9yc
8Ua41gaYBwym84Ybr2F8M+lJIGM0iszsxu7QuKJepSH9Dxcfc3lQFOeBitEEJeBp9gffMzknzx8k
V13gBvzFGSnVrcVlKSEM9u6cDHCHGJCk+KesYAuDgc5NdVphepBj+Rk4zE5SIo4Nm4TDprdygF5V
bGKKS9jcFo/JgAeSQMhP8GjyL6LiQMH3SY5dP+hgrsckcVZrlXvdpbzSFevCBoPQcmD/XQjhHMdh
W8HCzI+kaC7HSqFn7kT2Cjens/cFExUrdN0Fzm5sXUD5nZrmSELhuBJQWa+wQAYbgCZlHmggItJ4
sBNgAIpxvuBPVk9maQDY8fImfFEUuuQY2q7GH4mPiCen3jNDSbdhz83TiE4C9Dp3W22ED4JRPHYl
fD6YeOD3QtLPVctyv1+mZKN5g1KbSE0kFRvh9LDvlEfu9akTPe8pRB58pfPQASyJtzuBkbLPhko7
Gwk/EwpBsNgqY1lK9sowxl13FIR1pXWoyewro4T3O4uUjzcTPcKHyjD2xomSyBC5XkGtE8SfrkfO
i8dYK3xTmNV2sThSV5APm/weOjQHpPZKSL4+fqHY9AfEcC60ycYvswjOje/OCgVlZjBfffxC/g5w
Dialkt76789HQX9yOuQMMfPzckQ4G2MBl1OA83BI2JNye7Pf4K+LPcc0XHP9cuTxmQ2Z35K2FzCF
tlPgqA9Tn0m+DKhDg62tQabt7BAzsvrrFQ/kJeSc4C+7q/dDIwqU6BTaRtJQByhB4Y2WNX1RQQfr
4ddct/L5TCbDLE1BDuzwxT0N/2LDgT8vSTZMx8ckZCWe1mPGUqaMlv5xKOk8kXyv4vPR3hFRAOoA
o1k1VibQwtHyXXxnZALOJ5PZJkup3WnWmPDvzhtDn+8A0G45f+Tzb72qBCGumEXe6OgIEc6Tr36O
i1FItd4Qbw4vk08ftbtgUFvpmz5593ZvRsM/NZQWnQ2D/2hP3NpA389XzFv6mPx+C0kKBto+Pr/H
WgLUfYpkH+z+vDszR5VVtswlTOKtnLtPbcNVzW8OJGCBgwWaWfKlJkKJKu6vH8w1DICYIIPTJnLo
J08SZUVw97mLD96Qq6ri4CqEMVYQG4HYU8vAcB83VsCvu/B7lO7l3DGd88f6Pl46dZk0sxTJIp5v
Ekia0xMq4tsZpN2y0cYge552rL66OxXVpxpcFV5015ZB54MSeDOsFAJEuSZo6wnATVT4f0CodXH5
HB+Q7uXowjY008RzVbhoW7k1GTXzf8KFWmLUSrRcxLcFT0l/5HkWjY0Hu/PJrWyPvXmXZY9OSdN7
F2whKkOf8lmj+6NHthnOFm5grU8I3ROCWBxPgLqkjaKFuKb6Fn4XUfPx1oUxiM7m2SKVLdQyR0OU
kascPWKz/sn6LRYYd/7gRpfaT+feDi8vSX0rJA0Cmkw4ojVUfUatAPAmdPq/QDeaQE7Ei0mZaszp
6e6n56LPvuSLW5aMItOTaLrHh2wHNwfWSkJhux6QSFKc19F/xVhupB7Ld1elEvnm5RSN4lmG2vpf
mI29yW2sCvUX5S0IDoNGFUOGKZdyZ01YEzfXWgKYB/4id5i3TCoFhNIv9eSuxcc9hXnv4IRhaQi1
zmJx3eZBvCugr87DELF5TiSPGOKnGl7fjAJcSllkuPatcWs3P2pJwZBy3pjtC/z5qDWW3MPty2cb
Nt4aavx7489+A+c3gNUDrw223XGAwABgWgsC4JLaJOKLNk0asnBj7ITDYYfJQHXZJOhKTlW+Fguy
tnb72gGmLggUY66yiXcE9tjD09ivDuo6R8My2UQlwZ0MJGnnoie8dGgCm4m1imP5a5njZdqX+CUg
VE4gntCEcRNg6MmY/6X2Cpz0uu6N1RP5/0YsE6Zzb9hjfCeBCV+NOYsssISsaKVLZJvv/NFD3eyS
MY3+uCDC8XGl6arU+bovA1k2tgQtmVNsFnHMhvyHcE3RCLlrxJHf2snhncEIdtsPypc8s53oY3Y4
/7SfHuZ4UhKfjUNKfKy3Y6bWGXuVmSHr514MZ+1UYVF/P/7Jddw89W4BGkyZjw65y+6uqA0LaE9C
lxs4mJz/kFzq6k2vx+bsOzc+3pxxAyxtNxSaQV89RQWGoOdKGAwzuaHUvqe0EKpek/qnhq6AiCfQ
OZgLFLLx8e9X53Nstc+dZFF2SHwOio7U+EB/O0TC6mC9FxEDfNaAo4RKftvK3CA7JZ1UIhNcaDOj
G36Nk7A/zbSMkH38Bx+mr1L9NrRm8DHNqaoZXe9t/s33u0qKtB7faapWuUZiZtjmw24wLJfi8bHI
qkoDUi+9bWL2DTBVSj57NgCIvfKSU45TQ97Niau531ONSTedY2csYEv6/svCX9XFa4aFmRQpd6IV
qBe6hMNmGvjs+KLcvbj3f7Hcymnad4/EDgN/voJ2BFJV/1rv+S+lunSR9tLwIlW1KBH/5ps3rAGS
k3XcbAVkAGvkiQgrOfUdf4BhuuGhV7dL9ZC15WL1YVh7wuL35H9dHDpNdEO7McS0uj8+e9ER04Q2
/BbWW4qjvm5SsiafdJyReNGAqcYd3ca7795ZUrN16lc5arXqH+ed0iMu6d2SUUTo3bL1pjgoThC7
q0EsG4NJlpTSZr4PcWaCXj82SUKsaW7tb7EMy/BVqaonjlXtYNvg/OPtvp26mu1hS3Vds4x1rqD7
LpFONoAgm8dO7ggeQ2lMCWxmCnQQaNRIqq4HSTzmoRue1v64UXQNdp/nzr9CZLIKX9pdNnRigDZK
8vy+iBeF/FCu62tujwjPeFJ8w08J2lnNR3Y179+XNwIa0ItfRKfeYNJmNq4xG5Q4T+dOZUyVOGK+
SpanKACRzlxgxYBE1djsFZmxJM/PSGkhSmwM69J2VNQBb5Q4pxOYlO85byNkOVPqTZrgyOcUcvvF
Vuk7WhR4Wl0W/hU8ydiNeDvAgM8RTklSkjVfgHlWubmtZdrdMZHIC5gMZ1UQj5vALvAX5Yj/oCia
UKQWEHFJ7K5FhNARr5V+HMVIIY2wHqFq4qnVQRSZ1nHdBwCXOKVxjqpCuGFgzUGiSSjg3ZKd3+vl
ICLQe1JBZe6s7QFMv0hvpFp0zRN5g47OJwIAA5ZtktIo3TxcOL/UbWAIjCph9HNklapRU9lGnqeR
/i5/Tv5/cQrnzkM5m4cVoyzLbkFJt3yQZKvLDBN8EPrfUtVxuH2zAr5U8xsxYS2fNFXhVeURSSP8
8BZriQZgz5vhiRQ5xlBuTy3/kjBTq19mVR9gSRZad3RtVp5XDy+yJmACCW5dGuIOp5jDGWJLKby0
DtlU7CEA51AhUpequq5mAZGY8NiwYKsNJ0GJwihSUIEHXY5RigmcWcZzzjApiFwiTnnXtgwBEH7y
Qsay/5gQBMQjjurIhouw+1uDjNDKTz6OSG9ZwT397+mekVXsRrye7LzdxQ2HSZzc2WFF5xjG9ygQ
kWAqy+grR0eN6qynjxQal8zBBr8cy7vwWNuSgRZZUDw0VUjw5P4AwnHUd37SpH+WcoVm+WnzOXJZ
u2n4BwrWGaTD71X27afvnRCa6JbG6Wh8TEF9yseMC6d+z9zYBWE7o7Da/HNIE2eWYayGv0LoJqTz
/la/RLnX96naefWrDWPtVa4dAoA93iPpM5e+hulckGYa4VcKxz6RixbMzGoq5f257VX1M/ihJOA4
BBR9UhSN7vbz+x6ArVYygJmwkdhoJbfaulfCI4KyoZIg9PKxMj8qVUUquYfeoktOmnjeN5JbsIVW
hUuRjy62Cu1zwNAUIlDOUPP80p96CFrG1qTIIKM3FA0VSYwtZhiQTO79M0o59Bkw1yJO9vWBDXLJ
Dillhe9Mkji8zM9UWZUcB7l61qJlXxwSAxb6MuLIAlr66HJpEgT34eAFMsPABPV8WMFSQleMGryX
4MZhBM/8xNuS5tGs26ameYlyVLW+v1B7ppkV975DSuv9ltrb7eQC0Bwt4YnIHmDWi3ixyGB18Mye
Ewuhx5Lmj/KCDcWtGpbLKmNRTsM8gwhxDwM5AzhCfLlarSIggRWVUSFd0hHCVq9+WGZx2AslEFJb
BzD5+6wBw95ys81guQcSjUUyXTr+X8OwYlZXHJzgE5CiSQQJzHeQBCv3W1LapwpF3jL84zQdyLbn
AD3lvKIqFIpzHmIuDvIkiBtzsErS1ruwvL+zMNBIBxDLvIA2s1XwjjNPGhX40NqxNtkPk2hoywzY
FW1q942PUF8+5opLlxwNEd/hUXG9H8+6SxDQYGLed4jDISNRPkoL/Vl+4bBcYJUp0kMqUhPLAIpW
IJ2KXSswPcLn8D1vG5Yyt1Yddne8Chr7E6+nmJvdwvqqvEmx2OdWYYecFZhr49MnQgTNluE6D1wq
up/y6N2oCvBszOyHuY98Xjfz+/y6x4bo3U0NgSJ6c+YcuBVRu9rXtuKcrNLRRFL5Yy2N7B9kl+Hn
o73dXUK3tMeMqjvdWUK4aOZYdjhi0zDX5ZpDZ/OheRH6eXqQBARGOeMOK1PjZ9+BkEHGtx/MCBpz
4S5Q5KU/5iOskWM2UCXKzbaE5Hx8K/+fZ6zDUQDlsAyJndZE1QDy2WtlfQCnqbpvOkLBUSbLBGcS
hXRA6YJHua0tz9IlkBt7DpBFgJnw+UXFxU6GPJS5q0t2otVG/17YXteMgF5rYpKlU2RFuKohhh98
cmuKY4RXOA04jPBCUxEZTyaD17XpwLZ/anwcvWOYyyVZJli4ugG2zqvMrUmvvbzi3uT+iBy/UFc9
UMpt+MlcPTTU462g6yFd+Xg1z5lwtGY3AzPsa33LplMnj19/Ca79VJLb7a9nUpqbqroYl/MeTcvX
BlPCVV74T4hbdkXkA+Q/mceabNR2K/4dyONef7F4TMOl4wX29BN3JOTDP8hoW3e/WvIIz1Iayh70
lXvHUrkuCMaG7MzFavZ4l+qzdN0mDD8qJMmr2a96rOV98t6el4cyHORlrLVAu91PQeyAH85f68FF
rSZTsCIWRcoA2kKqokc/VOKlTwsZzYVBuPV4F3VcowjEOIWBpAmWgKayPaSf1hnk7lOTzy86RtyE
B9FbY0rCVx+PsSaT1HHA4wqmsSAPpkxnGLcW5kmjqjjbgTEnfHkJM7VmSZDOcKcHnyBf1wZOyTIE
WMrfkwkJmlpeYSEQeYa2d+2V3qReskIeTq4pomGN0SNECVV6jWRr8s/CGLjLcBz9FjPfwx6wyLr0
tFIs6E8uYKsMfhP4aooB22wV6E44bwfduZkQYAPNk62rmbOrvH8LZCAgom9aD/RxXPAyoFU5wDYp
bbtee5u14vAy+K2hCSg9VeTxQKBKNj4AQutRdYdwVmUHniv6jmRgzzEuTIpoYMXEkFPB9Y4m/EZc
tewBy/7AOEJY50ELVqej/MFfb3XbnBEGm3kgxFMITQcG+/UOzlXtsWkFjYKUsZZc7jbXxBM9ug+E
YtK6mnZttO3briN3f0VDUoaVYVU5wBwOy70QIz/E2zKhzQaijhEGbrQmaTM8Quh4PvZ3eyQ4kbB5
21EBD6JBaANbo+vg0E0OnW4qsvVZfMQpcI7YlGKvgGdRNjTu52x8iaS7uLiKA0Bwm6INGPa5aSjE
+g3rsinYNPABfwtAv7wSKbEuagb754v0/C8qD4pVelavpzeOuUDSbGRQClja46Q7C8SHJzwJGz6l
0367qhO/v/TcvThBn/WsMXUfCeg5wC6mu4I1W+Ct3RwL6dvP3VXLF6CWaepV8WHj1ONfubnjN+s6
FQ8GCLItpf03xySj9qxSn+Vul4LfZFLpej5JqHO3oIkDtFTLj65g3+5H2im8H0+W6id8YW6IGTir
kXE3GjO3sVm7SVsLVddrOlH52Sy4Q6x8eA6HtauXKKUkov+1Fat8/hhulJW1RrjmKwu6f5NkZfxi
t84ooqgU5uG3StbKIpQgSpWNZUNCqmPxcjw6nt05nx2v+Fqn+QttKMzMYu0QSVw6xn8Rbd68ikkB
JTLqm+3ROtpB3kN/FyJIHBV8DDXkHUEgE+o6RA/8uZx/lC8KPC7MDufBDZ7ThRQeUa6GonuFvWXq
cHw4gvj+Jlnwp7nxf8jom/PCSA/XFHrs/sHhW4uYmd3XiuoOifiUTi4Lrgq2x4DkkM3aChCgtbhJ
jRgfBNOLh2X39Z49984ow8OAbpf1woqnwCgqOaqjKglfGnzVsoJK0jTzQpfNvSgM9UYuCU1nUnD4
tFUXySXSuT9aSp7O7NhsHKL55MBpaVy7Pdf7Xo46XY6rszoXBYssF+/eqzttm9VUfdtmT72z8exX
RCAftCXeAzeLfg/BKm46mmTtplRog1yTHQXPgrxY+Qx+ZXLxPBUL4sCafIG8l7T7KSDBoIr9ByF/
IV3N8tf1lO8AKpBh7VRFpmyH2D+m8KMGu937TZ+tKAsRBfdq3eYD+OxYa0w1e8xiX6JC5L+B9vlA
g+OHHb/29zhKHA8IYscf+ssoKHAv6drPXmCnpdUX3QvsiSNoP8zRjruhAHpSb2ywNAgPq/BGoG/6
9Rbe4x8cuU2brDa/w1KmH4oyZrOoWSDTdojtJqmCeVPiA2WX1ed83QYV4a60So9Qre584C/6ew/4
GYz8HYXeQbJm4AoA+YEO7kv/sfbRlKfYQiW6rAA2rRzoJSqVRSFxwfHjrf2+mHJBzPJv/8qblchT
dWS+eK0q3O5mIG4RWIVBl4Aith1oDiy8+T4rhSe5lCO9HvvAofrIEak08w8kvH0FZZUbZnBEAZT8
+jRX2w6XLNmyDKG3PUHCg6aVIZmtNoZFEHgOlDnLskeo3+IETxH1X257aXXjOd1ulTbMoXb4br38
bgDqe2QTKL2cObrfD5xO6JWAoONoADqXZbpX/nopWSpddqwT1rgUCKGtNSknT9dC0O4UyWAl0O70
HXPjbxYLY5Ds3h4ntdrVxzhkfGQq12BQaYxwjFo2RBogqMYscKkPZIDXw8JZHX1K75PYpnsJ+hDv
uzpg9tY/Lgp9ujF0SkaYxyBp1yEJfxEr3236gzilW+nBCAI5HQP4tpriyhXY5++vWfnYdAL0hUuq
J63k8dftx+mPrZpIe657gAmQWGEHga6VWOkkKscJE7uFI/ZomxaLm0K00CshwRV1fOWjv0ZByRjt
CuvYAMM9AZjYrXCVeJ4f+Csm2P29sfJdNL06A6uYUrgAyoYUpuwy+vWFQw2Ur/tnX99Y0tR/D6JI
ItPf62uP4ORGLMzP24MGbOEMPl1uLFB6xdGi/E04hzGmRawdZWg7gPrtUR5v4L2AyxWsIUS3xitB
+6WY3150uGLd3g+hdU5HlSXGGJcVlPO9fL2jy1tkt5jxmbwIH9UXhYTmW9e4L6zoV1KpiV6loI3t
aD1Bw9V/E7+4I8gO7Ezf3FwrsV6v+aYWK/35jGS2dbEKxC9TBl3u7K4psMc4ykZ9UGrDYnnY3IpF
eV15iUpXRHEMqgZSVPZYrgnfQBhsNJ79olgHyhPNF4buVQ4ZPGAlNcCi5Evj92JVJEyWCjw1a3TS
Iv1qywFhiF8lQHTveRPsIsgTP6AAGHLnumvP5ndjKXJQxVy1VsGJQqYOdQyhx2IQQAeLUPbVXWeN
qBd2Ui2BLjXdh2afVFXhZ/dRb31x+S3fucG0iJ8NKv+6URkatezpehjjLMoAQNqX/8nQuQtbegai
nsO8dbQuHqIJloZGfT4hm2tG6QCEbhVAN/CIaTOskAdlHZ41iLNnNq4TxBLIUMp2m2oXlO2gFGmx
BlVwhZvER47UR9hUyK5QjnyOCxj1rs6DlTj2u9uJu3Zbu94xUMFv42EyPCcFqBd1Zf0i/e3G9GC+
WRtgQoRthXuGsNBuNr/Ddnkp3Lr5IxrtU7Jpi7du/LulcaCFKni/x1gmtZoej2eEPWtHlOYqYKfA
PSAKjt68N8KoryzkN6ilrb+anIhG5rRqeVN9TNYMKXQtN1RTBrzlN9DYij6NT9C4JfWWf+kFIqLU
/n+nMMSloD3kwLBLByKnz93r0n31z3ecngAfMGWr2HBFxJddthqhgz0x7yiFn102X4+i5KbcDSWa
6LhI1IELAinILldo3moncKCr8jk64gIOpYbjzKF4r1ldzZziePF1jByL58Me4lzH/WeegLds10nh
oXM6xx94ggGfdUZZ2ESZEd7QSzFbiujlSoJlRKf3lBzA9Itlel3WGVtTN7JaRCiyKueftp0xcPim
zPoyNRzaCVUCoKB9K//nWb/czO2lE0vbcj3NBFWDUM2WNeupg8xrO/GO++T6eNmvIKFlgmyRB6qB
k/847PxDJ60yVZ0c7ZkwDQt8ab4/S8Y17Tu569xCo+lxQwEmbuTdzdPTu2YdS7+EajNP62Vwe6d/
svaTIjnGIhhqTgj4K8YP6WWrG40PPmKCL5nhtviXh6i42Z7GMDCsqkcUhS2jKOTkg09aZVbm9xI0
fhfQEoMWM7u2UT0Uua5Iv2RkHN+7Pgq0pO1Nrc7qKNnOXr0Yweglx7I64eQvZcb+TpSeb5Mm8+SI
KOC2jaU8DhGgv4cOIdqKtQxEqFOqwii9FGl4u6O5iGuqBqmYAdP0T8KzrX5DJU3esOKgKj1Q/T21
Uf/sIUhYM1YUsMgdl3kMrpS37hMEQvtoi8au48Ugk7Ps6IbbjwW3fGeZXC6qHjORlDImQohPwMga
S/H77zGxLSsdBS8uFm07eJhcvBnOTJnLbiNSGao/f8ZklmB22LyA4VrBPKkyFtdHD/9kKLcTKxhT
pURLmrAY38WucoLR4sJ+HvnRDzTL7/xtDE4rNC6h+IRUGOhHWXcV5pF1aIUDzMqWLL0NqEMzU4uT
aKL1r0NNsz/5y4JPLJjKOXEyqWqc5aVW8G55T2n2Rj7ZL8BucgTcFWDiFK9yQPIdrM5HWk6cVysU
L2qA+GMZ2RuJizKnsV2L9mUNkM22d/mLZ8dCCfRFfdsynMTSoxsBuka9sTUVoolHt+/+WNAddfvb
zizHbo/EADaGi6g2pvTqVIMqbX7cqlFbmNShCKCSzO6heI8Dp6dsjXzZhKBeDnDcfMAzDhJ3NKSi
bVwMoJj3Gq3bJ5X3DVs6OHdSNWBfdoI8afvmLgF8x0DmjUfOcNhNLwVfGFhXoqAt6Uosn6jH/CsN
y1Id3wgFB6IB9RKwkvNdrShWDaO7MrGA32QpB4+rLJz0S0BrotzCmdP5TIFnXgh95GlzeXfY75ub
J/kH5ee5237cwoeGeTKLQcD+b3vy2a0FUOJaV7MI2JtSRCPB0nemk2jwCnOsnTGBCDUvrFOfJPoH
iyQZiKY404oED9J0Uq9/nFgkjLHLQ8DYR3LVygem+aAqptIEVQx09pio7G8SidupFyhrMRAcQdzm
/h0yYcUSMXJngJr5VJeKgfSylfm90TAF4sctezIXzqH05W6uq8g08DmBq9jmXloJzH+ihGnykAWZ
CHRqRNkjjx8Mp0KMr6wxdCGXVWmqtd8Tkio2MC+EQI3Xq5sL2MJnIxXImhHYrYlyq6TVf0MIBzIx
9n8jmCtv160NOMILfTKeljTIn8/XiqIVaHPZ7Yvjq3UBVLsh8NmlZp1rSI8q+5q8Kjw32PN8VSxV
IhRuPzf3wCG4x1tsqgYZQH7sywiZXQU533YpSMsIaa/K+WytEvWHaaX4PGHnQTQPguJ02zv0gAlJ
LQgqdZsfIcr1vHISn7VBPcozpIyOQ6rZohi7UhXjTY8qVoKgmvQRgMXanOdQr9mHVk7u886UaDcY
QsmrujFX3og+w5emWyG0Se+R/iWviCBYFKLSt9c7GF6KRFTRyHfqgYNW1Uq8Ui+1Rh8W5p101RG1
VoAjrhZdx5ck+pWGMDKrr/Vw4FiH+pRMSCNfwiGcfy+JDbAoupadZME7x/qXC1v5C20WdGL2/uOi
dIhH86PIep4wpgf1/NJ8lc+6I998D8H4ZF2ykhzqAYh43VukqZSwZPdr7qogtPsSKGkjWFErdo4z
QGQPll24LTB8T4o5bX/N10ftOx4y/Dt7yawUgAFV0UkMFL9U2MAH9+ZzPyufGemtIf3zYPo0wHR+
grKVP99xZd/86LmOoZSyQ4dUnZw7gQ45zL3VYYH9K+yFL7HLFu+cZZB6uV5ilKaxJFH36QCLenwB
TuASdLYdoPABECFWoF7qKNC86xpBBW/RNFhAewQlCsG5Eihx9qYs5gL648/mwnXF2vr77MhFLoY9
sK9mRvJvh9xe9jhLxJLC6ciLyU4lt7IFUPJHIomLt6wfyUc6kqxdRF/SeHDrJSQQRgUOK7DWLh2G
4jfiEDbMZGoHmOX2F6sQk99394FpGK3EkouszMH2oz7+De6RELIqX1XhR1CJLr99AAwM9Xl4PjUH
fwYqUg8kVj1MDIbKNsVRT0kkfmWbtEuI4ODMA501mt6mKeCBz52eJJv7dSDYCf6gnn+aWT0T/7Mo
2+L58/Jse/ZjaxZfsXKgBU3oXavzTR7TOP+vG/8STsPbfLMlGa0kuE8bB74cbBe0Yw4tjAzXH6Mv
KUWmVneg8i03fLCnQGT89izOjTwx4UeNPGFdEBe8t0wjI9b0jn651aC1brxvgf56bsvxKOEmN+Go
9rwMLRq684hZ3DZkrL+9cWZGtvwCfd76hFMWe76bbA7HxKn2P1NzrChVAbBS0x6RKMMzPHt77Ekn
JHfaB9/FEKzxwJRGCqejd0/HCLTEnUiYo5WT7AA8QUCrnW8Spb8u6JTTVV44ED/4VyASUtqneiE0
VRSCF2QR+UxrwIoZ2HzGxAzYv0DTf8pXhRGwVQwKfPnYxHKcC3xEETHxb0Ix9WEq+RAEO6hM9qOF
rwvlwdvmjh+1OFXNwb+9MItOFIhLbb1JvbNGUcDHnB0hqk1RvlP31tEcgoQr4lYIeE6xe9fyQy+6
BFeNhrMKlljWJuufegOyRrk5UBhqpmsJP6E/Xs6L/rd9VFyMA3C9MrS2KN5JMOSAg9hyZXb0u7iD
oBpiWdN7xzoB6a3sFQqsUathjddH/NWVuiDWd779PUhiu0SpK47RFvyALRUynE42k8UVZ+EMm6SJ
phm7wfnNDyBMplh5PJDrt4bW9j4Vs34cj/nZBTYMr6shOuwnjRlyE80Z0CWurB8QbWNwxYZm2rmD
awj+eSGtKjpLvGMvf4NnXrvdAuQeflvM+vxTJ5m+wl9udjMjAyswoqeeLU/XhGjrQnTtZlH01Nof
ozFc9v97aPWxyg8WgNwoBFZezyh8sdM7wzZeFwXVRdSUEXIrYxC5gOj8UmRxAa1m9EfFJLXW8+yU
rfmPCY3q9yUVuyoqk+cseUpbLQ+FFAIZJyypAXoN/FjtNSFE5Smp9DnLm0DfkyslpdPLX+vQYFgc
T+x5lr82CqhmJeUR1cRtJ1/Ia5KYW5k8isqMA4FVv0qJk8WeW+iko+TDox5OHwmSnho0pUAAgQc5
NTOsMQR+dEf9+TlUcHq8Em2j/ump2XXOm/PJWZ2XeFdZGUY2NdeJpWV1ydU7PM24YCX3/b+3/j+J
KbN7IqkfIe5coOD+adtzSue0SnpI9qydn+cUS2xXCI1HznMqNMS7lgJKtvfvTVzEJWRIMUesPMt+
OQ8qVbLP54Xopf+Aj/XziEfzWMnnxYFfAoJLX3z/4gHKSH+3lN6hkcKxB7uqq0WrVlzOd0GmIxl+
bDcVGkNDF0ZHHk55cF0HImdD7bHuql5SFKN48nF8/muvFLgdRmZ0i3G7d4qZQtKaRrCB80NDd5+x
sb7bUAjMfOhuSQdpvB5ZDQ8g6mTm/kivLaV4SWHzYOOUyz7STZSnXv1J3hMiVAkW5+3K2PN/a72u
9tbpxFqNUKf9yX+Z5GfV4IrkE7RXicaE3v65kPoTgqYEB/F1eMUn/JNtxqgmmPdYXo0xivWCdlxQ
hl2ROc7XrwGiHS9yiswZDwGTztDgdmEjfTWKwrOlWHtqlDvCw9DvAwz1yByPJPbOB9+WJdRZ8rfG
1Kt1AA/YeqcY+6uusqNrB9UMurD+jXRfoU6F6MBwzPrHiap6OFRWnB7ckB+gm8zZgSj7Pmpk36z2
6fO3wnscp+Z+f6jpL6ymdYfWnhECkBsbYySC+UF/CBGt2W+U9hsLqHhM8Cgy+5+kYjAJxTaMpqIh
lBFjsnl9fKjXQfmX6EuCPJye/3fBfhQc7896wQ0Yu0pUKXAC4/wojvta1owHPV6G+nUFwkjQD2h+
d2U7sZd/7t9W4axoxuwkNuA5m/ebWmqkqE7QWMBsP8EvkKUitgOvItk0Fki2Q55PqJY1AaB45SeQ
rdN/w8m76/MV8hLPXQZddXKJYSjQO/5XjyjkeZObsCz3I0mBDWDowI4FW5J6oov+Bmse8R1zTun3
mxK3ZXAGsm6iQXeToB3xDpIY77olEdfMbxxtoSXM6Zih4Ni+zFMisJruMaiCzSHr1sraxRwjFNMZ
cDx1vlRfKeXJ+7vpDtYbeXVMPfLerID8brQpbhvkphn3RBx/Mf/zrkqLbvtwIq3sipyOYa4/MIzz
efDr1OmyfXDnD/anOzgKhjBZpthmOgAZhZ2GA7EiaFV5o+1O0oStRFa+BRAciL+iX+lw5yHkesL+
NquFVOj0IIQTyCY3SFwCG+qNymANMf1ohlTTw0/rddbhg4umqCuyCwroR8mumw1sC0YQ2bIMjIdn
7xGuA6b/J/0yzOOV1DyTTAoWvcmJSqivuhm2k8q/IssmEv7v6/99zUVJiuw1F/I0GhQZmRyUVSY2
HTabAbfVGH+rpWTgo2EFe8DDTqqHy6ZtozamNe4P7Y/BNn0LAf5sxnjP3ikK1kmrkWNRiUezhpiV
Li9C0gGUlUj5YMOQwhXtpfF8AdF/m7vsUi8k2unBazc7EQwxjnArRwLJK8380fBA3ErpnJyguVoq
QUhhNKSCMoVbUJNu0g5/f7eZIy/z2jqhdL/InnNGGeEmqhdF0xafDk9CBqU7TMMQi20ZvuuqTHOP
Malf+46gIC/QP3IgGdzPF+u1d4pyQmcdA6HlGCY8VpVMMireXs+9E0mk3JCFws4Fsufd4h6pOM1c
K5ddhdjf5kwP54eEVuktbFw0y/xXOl1bwQyG5lZrjvmyb0m5J9yhDup+tXfdb6Rug8MlFvHOs1RW
1KMYdZ2Cf8ZJ9IkCi/+C81Gf3uJz9/aPuvCvIjhEwXzp1M4Rd3Eifdywgm7qoF81REkZ2aYtwF/5
xPXrwRbBg9otVD4yFoG/HlJ6AojFDFkxeY35PkWl46Dk4FLFhLwxgz8wC5nPqXJX+Zb9V9my2xyS
SJsTjEg0X/3aWykLRXWyUS4VfTuna15dSQTfsOSSVgLkE1UWOW4cfVib5kkQ4oYDB2sarBbEjegJ
m18FUqw39RNWMMqNAiEhzG5+tHyEJiuEnPwXUGAeccYVTSgbMAa26/SF1nsywsHzjLH3Y0H5ICDn
p8vQKnXK6nNpuPEZWg+4X9EPLKntQA6+CxKupw8gpcC/QBLwyVOIyO/MiUQCuQ6whpp2HjMeA/gj
DXEfgu+BfpNhiTZvNXLTuuU7SfUt+EDPYHDClQEmxl7u3IJyYez2GVr8KFFq+fkv9E/3l3Yetsv6
Imh2TXQfhl+d5NumcANqGCaTEO5a/BfJqsgVqHILbU3owX+zq6BYJvzG1xbM2XA6AEYVSEgIswvR
N/UNr6Is6BHzFopsWJ3DsxN8f5VtT6hAtQKf7XLfFQu6LZWZQ7oKCn6xT02sL0m2XKxFMO4t/CeN
/fXuuEfSmMnuJXLizdBTGz7bgaQusGnyK6PHnZKhX9xTaYYDfkgp3Jj+GPD6siyXMhO1SeIxOr5Z
CyK7LspeQCeaRHK7/97SD/tSnT8XDy+6eC2R/KxoGFTDnOIASGOaP9A3ALcBkCNfdnQSKF1uDesT
ubD3jxiITQ2Uw+X6J2esXEN6PgbNvCkWWroHSh9IQit7MeHi7Pnao+Zt64qLhHDbjIf4SkUAe4s+
4gvn9gnB2iVAPr8WiHIzv6okbB/A8tAcpFh2KwBX+1BC/R0rYcExMauC0XsKwsT2CKEHpLOjjQoC
4HGBbqs6NAbhiS8VQyxqYRg57GWUa2Pguca+ymx8urYhXqfgdX4FnI0AfAFyNB9RWSGFtvhwdG7L
wtjgpwTOHc9WG1qlU+HEP6pWZAhZuWNc6q8fmLH9Bbm6hB2hPkrYmeTVGE7GJHRT+bJG6N5ewrvJ
xNcqr256FZ6NtJVjQ6TV/fj6dXhnD1OtBP/ft2ZCHsPG+A23LoiUI5uxbHEib7PWbliToRvvuxWU
iuSJTpEj4sHi4Tgph49dPL0US+ecSx1bhGTmz+GYtPHweNJyCB8pljZsA/EskfoK+QCWfdHo7aW6
aDyzwiZGnynbheB1mEyj0xsA0gHdgR0/x3HWXQsahQmaawL7d3eGIU3xPXYKjFoDAgIcQ94hBmWC
bhBUh/OwU/fP9DRhih+ZK2ofbqp/m3+VNj7oPw8NlkwfQgidmHy+YcKbNcnkug58HWmQXzzYIJ94
sf3Z543DFJgaTymbolBWaxoj8MsbxbYFwkTRZRwfV0x7AqQC2ONwXUDUB70M4mkTOIy5M+MeddNk
7WHuxBQ4uXnhE2tHJ5Io1kin6XfCHksUD584BXaT/O6dm30N4KEQCtEwc+lLuv2oDEu8Y3vESaIC
vjek1bdrPJVB7YXkltJJStRSgvwOoZtkCtZjjD5bRUBVqYbdQgdv5nQbAuFKM5eyPDxuWak95DlJ
sZOMz4iUylJBSWfV0SqZeP4+UI4GoFoV8IjnXA5ZYeBSfclCaZ9PCCCC7CGmWhMuMLCxtywA+PRg
1Je/Q5E7myAi0AEf+KwGr3Lzx/rxQ/+Us7w3/dxKSw4xDsASUL3bsrwssnGnzwUNJI2EYItFiCMN
/cRv/dM7GNfrnU16agG+zSOSnssOaxZf//VuTHramuKTSoTo/MwUyXzLI86NZIRvPp0b7huQLWah
Se+s4DvmzNR87Ks6Jkqwz5p7U5wCZObsbfpBtmntE2gvKIoMRJ0cDjnPrDp+c3ZNGW2CF3JX/hQ6
8zvAOag3j6O2d9zslJkruHtJv8Dhx7nO7NeCYvaxsezCvW7VRVEJu29Hu7c6zYWOWXcTArIXiHP9
mX5NedfuTsAAvtLsgn1M9IPmvAsDRSaqGjZNZoE3m/HuAZzzamHbh6UV/Lj2R4ipI+B22tdsKZX0
NJ3L3Va7f7aukNLx8J1Yb3MF+slFalWXACHsRIFO7EtAHvuqO6Z2p1U7xNgU+AG//vGNSkNueARV
nl6MrbGTpJfgtRNLPi1Yve2sOxWmrttcopWjeteSHFUg6oY1+47c6FjvNxQ0Mg5g4zP/0W7U/aMT
FU9F7DB2VtTBN1u21cmrWisgwOFIhnB5lmb9FGX3wnnQPqBz4O20wK+FbcooN/l/6tBYKq0HHm7Y
6yyf3ayLkugNL+T+V5XcOnLycljA1vDsTNdv9VbG6MbOo9Lr6/25ZQlPT/y/UUAE4j+x5hIZsJ7V
TRV/6biSOcaDEwTadJHZDgUB0LECPjlAt0ALYfpgAiNnhokomQmZdlMoLVTJVCRL/v2wwfbFMFf5
PPurigDRy8opzOZy3jdlqP8kzQTzbW6OxQyD7pWG93VIKZh7It9Kll0eABslVqCOd7kiuaiykfnw
AMusrpGzbujxrrM1MMLs5IvrWcC9dpo74zePIsD7MxGe5mR89jwAeMTHHtTF546kPXoFbFIcTwi4
mAsXDVQDQp7tAMy56DCPLOVPU3sanH0eg6OQRRfeLWrKUlvw5JxiceytkjGxS0IgwyQuwLeHgXuV
7AcaexwAgKDTXqbC+IL+dPuWjQZL3rZzsa3JMJ/D4Xd9WJzAfE/OPF9n2tvELKmH7JWskt9nBDSH
wE57jmdggTvijxLHNy8IHrPiLzGHisbRBnaVqasPtGkKfVuVaB1Vxq2fytf7hUKLmJXJVs4zSQgq
s30u/FgMwr2ZoA35bIAQ2Ud8M4a8FleVNK9OC/OoEbGjlX5ny7+onYK5RxgYN/+gVn7DTweM9Ysq
mMJdXhxRR+Zv2YhX7XZ+7CuZY31J7DizLO2AeR+R3lWS93iCy/MKUmj1+cONlcm91PnCz0PfQTxR
ZHS/f/odtekjTvK3pID4hDs2i8++5lfg863B5OXhDJdy9UKdlP2/seF+aE1fkt5rRs7nDwjLhBvD
UiEp/CjC6J8uXmZuoQR+lq0uZNNJpwxGUIAgyQmVoOZvZWPEY5nY1SagKly7VJxwpTSLFFTvMpAz
2kU5O/jhCzbgrDq7DgnnbXYRCVEmN+0LN/eewORRfHISMdxxBcduYWH7yHpoNv6x0XpxyGTxWO2r
KOwaiUFUA5MhvfdGP72XfWD/pGDAldmXLf+W821LaOK4sjddbQlRH9KQ2lPUCKXESvnjXjW39lZc
rI7gnFIj0yK6Zro0+pNDZjZQYnF/NFsUWvYYH0cHQ8lqa6SYdYWISady88nJrPSCtVHoKJZ2T0Pp
59dTOhkwPofQwze5DQB6kbkwgOMKqv0pvLLxWNItwknSSailjYo+qysQqHeAMZvC4qeKsppVL+SR
BZKVXK5DYAQkQinANeREbpGpkqlHLlNAy5cbN7EG6njlKRdfkrD/SsAFANJmP2f+9FLqHf/0HHeE
YH7zM7awL6lufDXJP67VzMwIp5PNz+rUvqp+plfhLEotr62ghvmKiP7mEUCYacU1S9jIz2vNOhdF
dZoflH8x5QQs1s1BTal1nsLrb9bFdf5UESx2JZyuMT98bHK/xE9wbnonCG/pBnksQzdkL5YR3t6s
9Lltq3IvBoQNsBt/TN63OgY35rNKmjAQLHr7NBvdysOrZ1SAL1JtvwLHNc03zZj2GmGZUd8yow9h
dSvpOV2iLVasGMtXgDYe4nhakJr1vfCtv0T24vBpRsZgRIpF+RygOjMEDFgKS0W0ncHLfJwodsuk
1ql35ZQdhAXe33tHRZI1aCtEmrCCFtZ3k6XGH0MDYq4jdzsl1cmowtUNf9/KXplKNNhUnYpPv4KZ
fwt10860AlpR+UeQTBsquPILWrmxe5iRbmxFSXJgxetdtenYBMvgtUYHlgzaUwWHkJ9/WRZipcvO
hCGLQhDvQrdguTdIPoHdNatBLme4b67jiIp5iqS/1IwlZoAyHxDfH/tKiJzfMDnske/5XKdxqNnj
17mRB4wel7rNRBuiP4D/MlvHTXuxBDCQxfmxoa9WKf54QQYB3vjjYtoSC8uryVhgoS2O0QWmsgma
3LXnwEc7dmJFbk/xLcCM0sNRBxL2oTKzfXSr6IKsZ1vlT4XjXpieQT4E83sTGW1t5xNCtXdscuZw
aATzkjjs8Ru/pH6EcKfCXk4LcyPsiYxVTzGbp/x/DFFFgXu9CLEPiTewdf01cJmzpOKGvKAb7UuU
kKXAGt2MQ8VI1SGfvCUhAKvZS9qD90InLajvJqB/PLMU60ppvWed2mnBOM7wzkLYR7E2ej6+euJ0
FxsE+8o6lvFa/M75LwtegOJWNPOibR2QNRhX6YorT1N3RGBR3CmsBHK+8GdsdGLKLbDrcWzkzoBZ
kXLJLzhfP1yCXVZAgqOvEsSdyl8nmMLheGlDDd57P06JCOOpGsh4OclAZBlztKIKi4bfmJPR1QHD
pX3fxHjJ+yYpY0hKzwOXIkDXapP3iPl+nY+msbiTdYOJ5Glr9sOoez5jbaXX/WgOUo+8xbTJwOC9
dj3+PNgpw7T0+uLYN5v6jG5r53Ys2G9DErtfmtgYcJjlyUi3kLDM56ErN8EPsJXvkgBUIIsTEl7G
3E0CQY6/dAe8DdBxLIFPBflQmMiT09vjdDfoUB7PTo96n8aP9WezOZe5Mrlzs4eEsEVC+YuXcbEZ
YHxVT2lpedz/dyoTouywvTs4/wnhGjrixNV2csDPR551OL9QVN2+Qnf/SOl6waAHQJlA4u4Ikl6j
T510by4+KKmrLVg4Afo4bxASG1HQoHj9J64N20I83sjiputCnwZJnPhQc5+6HGP1I1PxkDNwfjHx
w2oyoIWV+LiLbugo5ukB9ldmLCyiZRgKy3k9TO6V/luJH95m8mY/tWw+Iy8wKM7ct60bPsTGrSHH
/7+gNqcu3bobfQnTnLtISoNfdLert5RVhPDfEAqliqPKCvRzNpMoYo98B64iQ3LbWehP0cHVIUWk
dlE4gHN+p/ZtlXlap39cWbnH4OEQ/eua9of5ozkuW7l57lkMgdIJ7IYbvrUKlMQEX1bdtCKwHRy0
NJ2+al1vVHF40xcy95hHOLiqfkZM+a8eY/otplDds+FzwrNqrw6gKKbnk4OOb7LCpz6h7qEg/aGN
xRqbCoLSAqocNm+gS+GbVttroOGXRkGbEM1rzorq4bTb9Q6TNvnSwBBbAwlDqDrtI/PjW7aPI2Yq
sj1a61+IhU8DKQ+xNvWME1fihm5swXvPf11WzRBY3PXvT6u4yGaFjQOnqylG2gg/8aMytZ/RN/VU
DuhVJ2k9NOqtko2UgsOYK1f+gHGR1k6d0TOqFsQ58d0Vib+R3M8vWfFX6grtK7wNelvuWN7v3fAm
Tl9kVZREaDwpvbFH3mswUTAuu/qSx3DvE/nqMnUK7c9E+CwU+bP4Vq87Uu71AjHU2Nwda8yex7rs
OzOzuidnRAGRd3j9UVMr+Nt10zCWTsFF2AsNIa6VU9SIfvNL0iN6ur8gARlMric7GrZn5gTDcXr0
Qyj/8ybxggjFms6jNlYrZZCF8H1DgqQtd4a2ugvnD+QFOpEWtFgLLwVfHG40Z6+fWocyZSDM2QKV
Bli22tXDaVpiNwf8DASJ1ZtrVglKIFitIIWxdpU0WzVXK/Zm5QcesuKsA7oFDzGywfFFvaUftrEP
f8ed9MwrX9MILDaDRJDIeGlSiJSfv8ELyzbzWUqYtFfBQhaV5XrcymWLCWMfUWF6ZnUusVbXljwR
W6+Ngnxwd9ywTgRyzPVJBDJn7iopq/K5DoFxHVDrvRVvELW0WB2ltT4ZCSGRF+AzUV1FFdoNBIJX
FILRQBX8vIX2WLlw89IK0ZF79isE7WiTn9V6bryfnIOkOIIrzzprUkLaZ2ZNDo8uxsIRVwUbh4nX
+v3xBFcDljPGEp7AdqNy7lVizCKCp+WWVyq1ag3DITPgmQNNejZGuS65SC7OHshT4SclNg1+AHqf
YnQu6NeC1QYRFzzmYE4LT36vUC/T9k8oZD08cvOXzwcgodjpBxr11T1ta4ubzn32tZfIPSwWq4n/
sOfOLt3JVns45oV9D/QMU6vDGXA0JYnWshj5vrMAvA21e19p1bxjfGmuiJpTArdCsdgCInGfD79+
AP+qhUTPjvU1xg6mIgdNURhoEIh1UYL0icoKn89XxiFM4OKmyex3ssdH59h0O4eyBZaN3G2iQxYp
WUvzSsDW/VAJsRCAUNOVL86x3RqUhmNDZuhgeYOUOR4xu+nJUxLKSv476H3Kv8lIvjM06yT7yZPo
keDSeULFEHEfw5FB4+XijpnT8+HgNuIMhQ3f3PhVer4Ba1aZ0qQiXYOhih6E6Cr4kWEmi97ibx6m
cDd3pSMxYg6Exg/38Y+nG9kfFQ5KuuZ72IK4lhxpqhbQm06NgAYHr4TgfvCIxHtFX0KX+BxaBKe2
o3ZCgmy1tB6U6z+zA3NXb+/E56pxAzVNNuE8zaBKuT7cLnVd3+uAm0GdnN8/Y0O/Xkef2U9J99vP
vZqxbbgUI8FcDYNboXvbnZ+r5w9n4+cq7IgstQApoLvSIYN8wSgSgwHLajol06yLAUWsCWrV1Q0W
lGswG/ZMAEbLK9ZG1s0S8q+lnWv9X4KvR5325m67wL27md88XbEt70aRNv7Pa2eSN5gSqf7ShGwz
PLryC7+/yzlvdL/Ne2c425/1yWNWAiG6nW4NwnACO5T2MyS2yuDC8Cyfa8jGEBZ+qXFXQ8QwMNhy
Q+Ue50dlby+xp2Nc2ZQfW8Jwvdq+kTKnPZ3tDnHE3L9UiIW3llDvoJidCYGewRczH/I+VEEQEo6w
nhk5I3ROZrKwHiMAGWQctIAXSmkzWZrbB7q4nvkVxBH6eJgMXIbAm94bYa/9hDfWPIYJuiqbhJ84
zKLxAZri206N89EvKMkC+wRqdTe0m7Jraonx8iZnDRhAiYl9ymwTRNsx0H6bBeIwbljR0nUgxou0
765ro6b6J/aQ4U/Y4FD7aQ8a2GfDoIXGF4seI6h+Hm7a5NeliSxfBb5R+FGhFFT/4oro7lqH3agk
lYiExOjTp6w3Th8NzjOwKOtFDOWt6vQYxy24i5VID4NUkVaMxikDRBFnKtcnDTUo1dedgCro17ce
USRtPAU7hBbARhkPz1JTjp/L0LSpXq4DwJyFjQ4wiGpGSLQ8SraM0Jwfh9Joy7dtu9b75PeGmfTy
S6O0Q5nBn/1E6pj9FxkVMhmnGWA44JuR62FYdv7tUlfJghNlZwC0Q/jCC1t1GvqQZ01ffSriJIvP
uLe6BQgPvdCu3vzi9PSnQr7MEbvrEj1hELnriAuRhKGsGC8IWyH5N79ZWHpLLavZuBUGUK4ZZDfm
xt2QF9abI68AaL7Edi3aze02k/OiXyxSPOzBpRKibJvxMmSRN9vtGMbs5LAKvRme7QBo/yJIk78w
I6Vqzry9Mftj6nuljrvsmwkwMUv7GYE4ZUUS/bo25NPk6XePjtSFNq+CuSYJVmfl6irSUU4/QNKd
Swa8B4JUesQwgR53ij1s2YHYV8mtp2ddDOkiubS/DVEYMn5iQsYux0/kEDJs5GJOe8su+X7FPewH
elxHDSIBj5jlOtGhkGM9FGQcKCwj/gnHaUUtpHpckAekaYHMSHxGC8oAgNiq8yC3CmPZGwh/P53G
B9LABayzFdwFDtKalv6dK6UlYqz3RlwFffgQlXSZlWaevntL/a+RXPNGj4LIHsxXX7sUY1++GHPy
ZU71Fjulk4FWEodl3J5cePlfUPNf0Hu5Yb2UYuVMMJoObTjmwikl8y/220U6bQFygIL8KCmIqtvr
gh2hte+Cp8jidPZTMZBHAP8nVeDe1xUgYC+1dkwGpVY4TOhbxbYquPAp7n6bOVGWaYdvwYd1Pb9w
5ZYqW1LdlsdhMepeNh2SJlpqcpfUev0QmMaaC11tF7O0s6/0GYjJQe4LLAO2l3nkSc9LGmRhMOOT
YlFIRHrXzahyNKbUrkjQxl9KtdAZ4hgSiCI3x7CWCtmlkCdmFrgTSbDAvoFSwH2v5ZmnuyXGcenr
cuewf/RRQiZ2kble2VB7IYhtCtRyU1dATFc62qp3tREwEmHxB+ujiWedKPZqcvquG/Sk2tK6aRXk
9u948q970H/gNVggGIjwNLseWaI/x6yx8rFGgs/1cHguwSsWb7URvPmRqb0ARDUc1Suc0zS0Dh5M
R/7ue0JCsV+lA2IkWthbtVHNoZG9aSTaxVZGKpfAVLzsidK1qLtmzKtd3n8u+GWpuZCS6TUvQkDh
3Smg7coHXyfxOprh8TjoK/Tn0mxIihsxhNvdh3ubXjKMdD9RZeZ8v1l1Z4pQR1xouaBeM3W9DT1r
ztcGXHv4njHrPlqvBcQXyI8iTtifAQozBLa5rv3eGUZY3gpnU34HCzx3ipZMfQJ2hZfUWfHdFyKV
VF695ZAJxRqlOJXEnWovER8zx8yxtSfGOFCaNLFjdqW2ru7ibd18OZIfynU2/xHVjgU/QO94knaM
ftI7PEelXHKE0wBIDqD3UDXx3X7M3nf00vYa2AOXgUui3IXhYfIX8Ix+OjmWeoHyXg4wb/nFfQJj
MI8wCWfoywQFTvSrdnnKIo7ftEhGVbldu7S/uaq884wkn1WwQ27KXpg/wyY6IyKBiC0wLkN1+4cC
urE6SCRCMjIz+djNEcM2IP9mztsHrYGWqpLfzUOBwZXv6+a/QuWtq/6tC/n3HrdTJtTcjH2oCm+9
H+nA5xSBD1s3mWclCXIvcZWocVyN21Famo1SwxA4WOFRfM496XFI5lknEgc8TUmLwEiegJq7P2Wb
SPvrPh8Dwjlzh2SErZfHntu02KB3AjAB0dHn8cK53tqZVD6SMg/vIEYnvxDZiWIPhfHrYrOjBBBK
niYBhe0B3LX6mjwz7EUf/TlRCLqzTajU4tUeQYpRK+ojm3l+w1mir0JBIn1Ekrc0NLgGsDmPnJ+A
LBYTaGf4j+JJuj6QdVA6sH8CzUot7Wk/w/uWOO6GXHEfkNjO7PlJCzj6Za3JmgqucpRFlcCEhUvf
WH0BH9WV+XCqR7x6vORMkAT7TljIBN4o52zqiUnQTpp6XU5gunVOM2hlp4t0/4xCWDARLz7O5Jde
1uDdBJ4ra+hMTIeS9qyN/oDk4wDY9BGTwL2+jtNulVovLTBrpKrTNOuso1tbwTYsquhSKUhEjmA9
A4nbK9sAp89E4SaDoQWYFVTBFj1ThHbHBoD3tESNtpHl5+NNtQbnjUVqYB/4Bbi9JHWIFMjnCKk3
3szor1Np9PLx4BVMisKfDAeWpGSakThCZLjBMFc4c64ikNNsD3Wec49EWrluj40wzHLpCmycwcxQ
tybifOBNYtHRyvg7sEML/a2aMe55NK8SswA1XWu86VyTKhlu92uepCmNcxy2Eygg6Cw8bIKLfUSj
XWh6/ZaWt2mpefOMtd7O/jpTXCzLyI47N788HeIlmtjx9pFYpogYHkA6cFuPTIpMXylN4XwdOJH5
wJSH0iWtX7PKSiskv1l5NGp2BkVG7LdxfIuQ313DzYUkMc1J/X0qA/fiZVwoukF0esJkSB+Xr/Yz
IxQKUzShALfpNyqHneB8VRaNTqgK8g0TkDr1iOnyM4PSBFR1upMv9PMLf1ciastXj6LxoIjRtE1p
yIBYGbYOuiz8ksaUy7ygoATWh2gjqWA7U738R+bKhlUffEjU6WmYtSmhiCMN2XPDNcbvK/9iNFlx
/fQGMfTzQ0PhQRzJqrgJKTgHNRh6RdbQEIsdBn5Vfo9oEoefm1O9cTFmuVUIiWmb8TArQLY5kt4a
KTKiFG8I6qh3w9D+yJI5hB6RVubHUvq7FGXs6ZfqJV5Yx77cdi2fLwzrG1QpmqzyzeAKJ01HndzS
o2Iphhi74zz0nhhphM6ShjHaS4Kmzb9Hb57NNATGwKDjww96ZSZ4VwcXNxEvtqVQ7p4UnF+NLkwg
3o8t8NN+arjC+rag0yc8MilLg8yZ6WeYiOTeoD+otqBu0pYD6HtDoldCSBD2fTHC/M6ZujUlJfXi
TNQHAZqzigI6escEOrOGPH+juny0Jtk3gUoryaKu7D9WZsYUl8mpQU3HGuTyjNbdcW4yIdlnBYvW
/b291WcFGRDsysyVQH115JaqSVeQF5zdK0bicGf9fZH8zE79aGojIh1Hd+6ASViqKz79ltTkXqUk
X/zejtXzJ8moelKJr4xflpcxQmGNP1gJpIP025Qa52/FEHDEpA44wud7HmhQv+SQGxwYMkLD2Rw3
n541Rb+Sj6Wmk8Oy0t4J+A/APbmedlSpKaw2V3ltxuTAHaR4GrD4D1Cvv5AffhixS9G8QVRFThhz
7MRYNz5dsNh7BjYCjnhHlfOJmnwVzIzrtNg/IAqGSMm2LTyY8W5Kndi16xSu/nXKzZfFu0yJbbpk
OJ8b3nSH77ekdac71uKB/2mGF458OBQlG5nXO92LmCycPYiTzKJS4V/DiHsLmmNChWviTVmeIE+v
hex68JYe1YLR1z6Nhf7K/47WMEOt578oRphikYcXPxsRQ+8TVl2GGR9yQhQorGZ7IyaP1S8jvzkV
jsjnAxq/fzhRImLl/uTOJ0BBmBznjfUmOoD0KtooY7gv8wcY0XWfNXNU4u45cePksLRMkmNNvKS1
nUzJMCpvsGTK2ySc9zhkDD+KxjC5nd2orIM9T8s93QThcGSeMfZWFixnzJPTkTrnvvuRopru39Qg
AW07G1F9egfh8o2DPmmwL1eM419PGzYESf6ZlTX9mziGywqKiDNv8jnP/Gnml/1k9EOSyTqihpUw
+yypk8MXrPIp6i4zHm08N/jUz2dE+MvMARSP/UE/rZsJyQtuq+hUxfyBozG+MsMaZxh3Eg/hbFwh
MWcl8VvhKLpUUc8X4/KJIWPYZlPV9LfeYTloCD4RRjLa1BsYeM68Fx01Htq72pM6CRk3GPOCip8p
P39l7Y34tbw4bwTyqkSortUlYAeFN5o7YF34HcVg8ZnR7sSf79wXtHkh+dLQo/AZLnBWwG6Snzyb
0cylPJjVZz7dvm/rb/T47YXsV0XRtvtXJ29eNbpGjCfSZJslO/JdLgT/I0dQE1v5vvxx0YPnhnWh
m2l8mfsM36PTsztcOAoExDFHq2lw+mBpZmMpfzGyMzMC3GY4PdbNtY0iBIafpf4JWXMNDrCj+MkI
bHwhm59g+AkR9upZgQ2RcC0afpYZSw+OJVA35Oimsg6bvNjc7d0bUq+OC05MXjqgh/BLu6PARXsb
pqaUjNiKM5UuDJ7EcDhwvYP7CekJziuGJRBspf4L0JXCYLzhqCnZa76lcmwyIwu/4cUulDkFy1+6
xW9KjdbZ3H+CbkYrgKcSU6Q+5dHvdt9ULfXRO59tB2RwBlWAOPPvR4gzC1EczXv7OthuDi2qEeh8
vJuV/zieLaYNteyT4QWdgslmOWpJwfMACoCjbTas7g5bcVZWi03nv7wajqMVT5TwLpB9+/DqS+56
RvgJlRMK6/hffWD0U4gVC4H+asQ3kDXXWV9R9lOjrHNdCFtUHmvXPIGqC/EHGUUNYHt068OYbOLQ
hCnQ4unWB/vg5iJOScDadX4aejIT7h152XTH5bwMUWmQmWiYzlAFKu7tLUj4hG6OyYv/NvnH63te
xbd7oH0DEGwYiuOO3eM2eF/t3OSIvSxLNKbDyEv2YhB2CIYj5os67xOuGyl4DJVFERIs4NdOOoZN
5jwN7c2xafZV/7MLBp+AlcQfAeEmrazcJntveQjVwX/PbLQzo0OY1qdQRD0nqpDqgBiNn02C21I/
KzbRECEfZJUalfqsURwkE393fgFeWaRsvVOuHA1C8o328CbZcLh3XJSSaFo357yS/+2JBDPgRrXF
2Nr0IfUXOgrjSiR9tCXRAfHiJ20j57mAevISFw68jQkRgpWMcY2dtnPDSpCXmB1GZTZC2Hl+bPRd
Lm0Es1YXGoTjF/LK/6ybpKGmpzp2coPyZU5lAVv2+h5hku/Dbvn2sixT7x4/WlT+MSIDoUZW5x6u
MUPKq5h1rRJViBmAzujhOJio6NZmB0tjLdlBdFm/4kRNMFfx9vRh7RXmgoaoDcz+ZZxlZ8eseFPb
qFcSOhELMjn6cHN0egL4IPMGPVJ7T30GeaKOpps+8/Du4D05bdyYcwTfZlLA6FvaINPvkntr6NHc
bqWGeXLLHlBohRmQr6uzDfg61wPaw00xuqErUvXcumsbPmRLKfZGSxgo8f8qAwJS1MFBukcqaUu0
T27HCfUVa1DsQWURcUHipqX33QblYFKK7243CWI51ITQLq7XUgY+hE8jXVYJw725lDa9VzWE2U/O
kizIQ4XZ7erOV5UlD+SehaICWNxmIAsMIBlG3phCgnCaXpvTsigTDeWg3gtTvv43heWbuYlNnD5c
0uWQprv4b8fnY1znhRohtyHJQ/IZHeOqZg9Auu8q/N5BwbjIRr18TXJkZ2I+w+EkV1rLw8ULbaj9
j5P3GQJtdxdJD4J0060OddmiD82NI6LP6dW6q5JwhkcF8OiOYfQoPG6FAGS5BPHZBj8vi68NDY5U
XvIGWhnaw+61/HAN+CJAKowVOpBrtV2rGkPOv5xWcFs6jyGfOPudq+o/hFp+XeQVy+MK7sWgSJmM
jfSsj0BnkhIwMuY7OksChDsygpOJHlhibcbkm7J/qIbqKZfDZJKT93NWGvLf7MdbK1PUtHztvamU
NtP48oLQIbh4L/KK9xgzTKumCBsHzGjnsZK57u9j29ntTE4czer41cW701uECpdY0f1UHrghbdkj
hs7tBf+jumGBgBZv2SiKod/7wXn0Wtgf52SntHhZ5sRni9jmoj7dmjg60CJKPSJYfPAHMGb91IWZ
1hOqoGuDSShWNmOw5ptjcCeo1DGtRhdDDudAcSpg/HbAxHuQoyMqY9lSv0neZM9+AHp4JwKeSI4E
oVJceTczAn6EvJ9KvdxVzTt/IWm3q2xKLPEOW49it/a+vCO6ZueHymMnS3c6MxdI8r1FntK4TLid
h6McHQTi0qv+N5qVPGvGChWxxzZ4IbwmC+eq99SqAW44685wfhMNZ0Al04YELVOPsnjstURntBQD
FGZw7qiEEVGLl9MsjVOViEUx7d7HqVxgYCHp2yxzp2jZpQ2EC/97BA1G/vhyrVIqr9A/fEmKuMv4
hG2/PpocsVXSI/RArEp2oHImvVAg/5v1b4ngi7JR2IL9XxRYtwua+gNz4SppMyxfzz8Q8oXoWAaY
rtTGIDNSeZRy7qBDiwyUkk54iibJErBcLFGoLW5BVfzLpLDbaJ5emXT2n8eFT/iklNdGttU87lGi
qiBmFaw9BaB3tSJmE+Gb6GzFFI/10v7qhLq58yDB0lzzeduubiwS5eODWzrUDgjOtHc6JiH+v+qR
AL2vzMAybaOaWDBoRO1vGD7LFoglnqYva8aGby9lar/gBnEto7ZGINL99FUbpvVVgXPkC1VatKLX
wu7na/a+hqHB8F2zpuufW43WOh2e147oecb7//PO1Dfw+7ZnGvebJvRoLzwM/ZlsGqs5Dyt+6ZmS
FdyQruahLHKARvcbfTlLvVyT10OzWPDwwO48hLcmnDufvwZYJUO2BPrntsj1f2FTC41tIbC+/R4p
xBVk4Zj/q/p1Dft/msDGf4Mg/jeuvw8dj3EQq8ztvz81HwDwovbDcczo4s6U/ayP7LBQKL2Vtjla
qIg0ldZXDxf9Zqs9dbjClpGzGN0Kv2+8WvHODw+sMnYpLMDcJv9u6h8P4o1kBMQXdUgh87zog7Zx
c45xr1q+mTbHF4gz1MJtIWQ4uqI0Cpo44zpGtHcUmARVZpiSj+JG0ry8IoK44hp+QpeWUVhhwXwg
G3Qqi6DNp54lvfGOpwvFIuV/sDN73cdBeeL+Un1l12+1yDprjxzJSrriJ/jRs05hfW0x6gFwFfvs
7sBMmSw9K2MXjnW/K0fZT+JMG89+4SNVpWrgAsXFKeXBQMKLxjl1o3Aby2dmn/sDzb+pvnXhAzkm
HIHS+XWCrUbcT+9XcUHhaAM3W9ZMUfb674A04HUTZl6pdSYe5pLLh1JnJkbVX/E2xs+TyF1TJDPi
AAgX+F2meW6XTcf2QFvU4uMQ45sJzom0VHPjHrsnL3i0k6WP+IjXDH5GhfdCkD8D123kSFysHN7m
UZWlPLqfPVoQJ4YHLuCaw14M3leGeh7zN1VFDGQMh02iMf3UnhfqUSHZshDUofbXpGzMtoQYuTLe
ldu82YFvWFtS3fHKc1AySzwY6wSDOr1QlhYU/KCa+zACcY2ifaOuTfng/QrcB8hEhOoauEYB3leN
WClKXoeeD11gTGuWGhLTPjzQUafyoB4bC2NxXugzrHjbGmU5JCxmprQGR00q7/IDVRL5ecdL0+LS
Xb6PjYl0REOlPwMndUubavKFxgSDQxMbf7vqYzCMicGEmIpzfoVq1wgr8IM/jB/PQa3gQ6rkQddr
dswwslD2qg+VDe8YZ3V2oRA9qpQf7dP/XCLeRADPWy6Ye16Wjue3TbZX0QMlgUph4/Fm4etfL5fe
d0xNwucdox1UhOvDXyxA4qhVx/t/4JWxGhRlEikyegv6E36EheBNgNPqza+5iX3WFUiuJAojHEPx
M30w61gqpPOGbjxyBksm5XxofzBLwBUB4K2tXJk1VtrFcci2J2ppAO+OQ18y9XQzkhU79Z4eI79Y
6M28rS5ZUWubrHKlia60MInnUvJv0G7FD7ZI7eru/GYlv42q1UuIm8Ka76HAlhE9MKWcbIKHavf/
lUqC2R9bzVdxqZT4o+I6Nq0xz7wh9ToW7YwaPSGoCrqQXZqYsZ1Ef0iIdsmOC6ltYzAMfUjWSDd4
Mn0KPVMGCQQbwTlmWNMrg00aUGxE1FXwWI8Zrmj6R6VMjbrqwpB1+slY+hmd4P210hZz/iKYPyIY
UwBc5fr6K9+xynnmGeL8eI+4qvQ5Os074mcWRuGZlY+QMjwRnw7aoBK3rszGRvBmTPPqKA1uupAT
tkGX8gZ2iKC4d5vuxoRFXq6O8h//mPpmH71nEsWfe1NMp89nTQjFgfxq2eg7Q4Vc6G5DSF6bIOHo
OV7hoA18o+niFWwfY3CprLIJaaWgG0/lLdBgNiOr4HTxTkFNPjzDmodfOeSgf7T60a1Y/Flm5H6Z
4WH2OTuZVzim98x2dZBlcaYno8UvwE4CHAHEDb7sYwkq2S6rUTpcDeuWCvH/DQ9Q50U7qcWK6eHf
izsuod9fQd9QdP3mlBAiTu+g4okXZJm4MO0DgExtPH98r/NYvIsy+mvAzlZdgz4HdrFWQPEq2igl
k7Ckkp23hJazjvgtUl6e7MqqwqOdlc0NA3Wnd1xxkFSHtbZfvwTDEG4muMQOdu6td6Ic+vcUR1LN
IMs0m2t5YSifRnjU82ofl8skhh2gMtNrcVqZSeMhdbuUoalFgDNeVe8CMQd2yg3ojhNPFd9uR/Qj
E1OWjV62bIzdglL/Kc6PjPSdFzX7wC6dApcOYb8Z1VtKy3CskBGQHtuHOhPVuQfgf2pj/IqymJJd
EijNm8pkIAPraLB6EyvGy/egGdnhM6Lqer7Z9g9jpFN/nB7Nr9ABad3cCiw92zuwYslIP/b3Lw//
QDwb+pDQX2WBgZl0pmk4jq0+hJuek+iGyupQMQdZWWCQDep7hWukGS51IMFkx3GbrF66qOZDDe+o
WfyLSRyaoNQL33x0s6hzDMx6aj+xJvnY6FDABdMAbktkZO+Yh7SYxxdCbKKaZNgdsqLQsMbDX5sV
+sy4Me8tnDlj5epvgG1hCpIlpPBcTDXHZYnXWK89ONNw5cnwI9Ip+R2ydix8Ne5j1CEdBBOktumj
uIloHXKQWlcF0ENxzAwuEfg+xb5oS1rfmoQyY28D9M8D7sOpWRZaNSU2Nc+BMtUuf0zgopneoo7J
9MytkfQlhEAFlrL1W1E0LrbzZNyMhJ6bVoqoHXSnI2LZzksfWaKHiuJv3wPflMyIesLz5W4LeTzG
vJIjlqryYj2nItpMt2P7fe40SBb0vHjHK543Tk/iTjhMx5uofwX/nUaNU14kNO2mottRsO5tTjLY
n8k2otsqA/KIHgaedkZiP91zG8jgZHMCoWgJUf3WLecjHCM6SIg/XZcBcQ1DgCI8vxCy0NY0LUJK
KrjEhtYpqMZ6iyhdpI8rsNvGtv9Ti78pb5l7+yn3XVvY470QRdEawNKHhF6QhLPod1ChGu1tltFX
hqdU0292tRxE2QA4Mf3+roq+dwlGscWM/A8xOvVpDBdDmXlqATmScRJwrJ3DXJae7aStCfE/2ZfY
Wx3nOSli7Hd8R31Rgsj2YU+yeknZFVUYT1DaGBJrCBan7Cvf7DXp4KfKrCJ0DneW90+HgVo9zOOb
LeYmjYAZGk0/aYoyxzxBqxZa4LqKzpvoc1aM1cV2NQBH8F3XT26LtDaKWnBS4zxTVgdqxpbmlNZl
4nu7VFrjSz5e3jFKPU552pWG/VEcOnqcI0XknPw7V1mX/3o0gg25v6Csj9a/9CjsLiqobXLCTrL6
S4Ec4M+pNOSo5dVlzerMWnhAP656kJHpbycZ8EE+VUwhRN9fYJpKjhQ2Uv8lG7/kEDM0r0uYt0Og
+B4e1kbYIzjb3jU9cKxtDwUjP+zpna+DaMcsqcHymNmW5kjK9C6jrLQGwb570w1tWaG661kjF0Qr
UKM3KsI1Gm3N3C81EK+HCUmFZXPZJX2seRWcNeftpHzDGHanC3TcQialakOLTVwaafm7UsCl+vK3
TBdz06nQa4Br7J1Nf3eKMAUkW828agW/BskvhSnyVpQbqS5hUcFT5Ght6u9xji3sV5edQvCf9dZz
ktQ9G+GMxQc7LICsGi0MzfJ57KC8g0PX3W96EekBV2PV47DYprVxIpTiJWplBuBOwhtzxP8zMtB2
+c/tjFydHyu4WepX87n+hXLVaEN1vDXd8CiE+zkgDhOHNc3aVumRQlstr9cII4BSnV/U6S3W++gc
I/Cz+bTE5S7OtptBdeBbXivx8TikrR724nzZUIqH9gJTAaUYo9HYr79bzbWp7jBoDd9xbWAgt69g
OM1SaDRz5U4FH8MJgwnecY3UeGqt7TRDiMaPSseRFIeFOEvgjPZgBDJ//Yn9bMIGatks42tY5qBu
ji0nNRNWjtfCe9aKftjMEhM7Br/HNtyymE4s5+RG2Buxc8ijNix+obiKr+cPNDojfEnjRIoziVGm
ESeGzr3Q8lzEyNVCX2AjNxwsbbkSi+j6cY6BtlGzAYnQuKHSsuUTqYh6FUmr+PEN/eFkO9u4U39k
jIQLIx5bb/V4jmnRHZ5G443U+2X/cHPIltHI7hOqg0Mfh5YQdoD0t38d+p6hG4IB5hunWxqMNRcX
KtwueSP6sPLwpJiStKwA8Lig30muzq8ly2m+3Umk7MgjpyvXOfOlRiM+V+zwCAXN+jBMsyxo+VH9
TvduTnPuOoBqcy4p8TCqJxUh+TRvNqv3QPcadqfSWTYMXFpWmeO7e7T1BaZJxzXYs6bspFmV+FZJ
TR1F0uD9Q4t6yFQaDtyEwHVL7ztHzH2RDQTe37Z7/b/s1SFqg3SvT9NPSJw78stvYcZkV/geZyOj
HQp8JGkVj+voBDYkQ69yYX4gsb1Gjp8jRPBLgGWs2kS4Nc82vhEche2D7iBUixpK+dDv4zBa7HQ8
x6K6KMT7Nea3WN5tUQOO+OcsCOcNTUA3qxS/XR/Nxg7VyiuR4TB8R+QfgmEpcp/mBhk6bo8hKXe/
t2P6aV354vqcqSZJd8BeQgMlg5awgYZoe6J2gv18mOuLnLMgmzc/sggRGVnDRWJA16V8FTXgCw35
8fuH5B4EvfxbGM0LQuLH6ta0DdVHLCXIBBFm/y6IaMPGDA02IHvRSlbh7siYbrTC5muH+bsNulUj
JlXbB9Lo3JsT6U7U96UzqwyhWU6uKfqPtCtkuoHPm6+AX0409hl0hTjg/sVWFFPLbLFwgUpMZ0D1
1waGcop/Ez5r6Rb375VQl63YHDByK+BUq+H+TKzAr9ad47s7nNPPz7iHbu/xY7t61MXHK2jq1lfR
nAGLagx43KXW22G159UvpMdIZjdoizgjy6T3K8rI/y5mPV/9Hl9XkueV8hRgbd+HdhA79F6U3XMc
nVoaftyQ1ofjkkCf8SYr0iB4yRLxYhYNfecLNlxfo0cibjxOvRXeUySfS41Xg0mXW2P+YC2sWlbS
OGaqk7NCbiJ0yEWOvjK2sGQc2RXkPoTmlJd4o+AYGkB+NsuIrWwZwvWWsSyGyqe9eDzNM/A4DRo5
7j7ap4ICIlKa58MLRW4wRTZ3n25J4O1Os4q/dorCupnaZ+opCuen+uJhNb42n9ue0+AhzJeBxGWX
/kStFE2PbfclKVCj/wascmWCGWM00Q3ZVWdnM84Qir87Q82bjO0IZYVjUB+tbpzAmx5Q/QUk69HW
78dVNHDbJCj2RfQxO+VYpMWaQDqiKXw7QT8oh7RgeJ1QwbI7DYNLy5p6iCMPUrI4dWRpip3P5TuV
b30jq9GJRskD+pInfhn8qs+q44erV1QwP0S0PUMyiea/OvqkINeEIEwbTizTeLrDZQZOcs6QGXz7
9ih8108GDww/IY3b3pef3FDTb6mnAfkQX4hOiZExXS7EO+MS/Cm6/Vs++gWaHLN9eCFoK4QitA3Z
sbb/kR7sdw1xP9KevfpPl6JCpv9xK2tvxyOYB+wQ0SbHNExCVDQTHmsQEvJ71AoQU76wcmzN978J
LQqyw7C1lMLjYfapskrj7MAOwxeB2yQBihKwi4cWszlwk4EGEVruRKZs79lUNf28RSPqD+UevYvs
babTSGxuQ5BiA4w3ynrdvsp1cNV7p3cN729PxVyj+aBd9J8fSZH6+EnAR2RebiBnu6umlij+Yi0i
/E8u9tC6xSDvjZp1N06QmIXhZ+vZ7JWwsej3xNI+JVmONOIxxFfrI7AXMbnNacWWsuIHlSTjgfdZ
K/eMJwVQdBSeG80bk90VK+eY7zbiEyPQl1Xo7H837RMe+xPDWomQuIDj7k8v5wJxyrutdrCKXW77
Fhl8eEPvWuNeomu+joRtZSd24bvjCkpiK4reOidVIdSpQ3+9/1ETpJ4O01wTo3OmqSa4GLb+v9W2
tEjVvkVOsS44HMZaVfFntjJWMtsETLr3c9OEvVXGtbMDWd2NmuC74+va+h53mDPY8ZNxFnjl4VxG
7FYvyPndWvo+YK3pCnxavKX28qe+9+ipJroRTwBQoS2+c3V/nz0eokDAuvBcZM+2uqAsNEopoArf
jG7R/tRzxAP7r4pwDq9/jBK2k87q39aQSWhKpOSNwbkswZhHVDyRVqSzXqvHuqldlPEHgsh2zsAC
uYF9hjAOzuD6zaejTZn+b62h8yRBehDAUThlivdWauSKL0/hpQfeb+r0RdlTScnx0VxnWdwDLX4z
l7GQ1nGpdqjx6MQMQuvQBZtEBjeXSU96HHMWtKdawCxRS/x0EKqWvOr+pRES5fpZdHaKJeu+tFXi
ODcjU1BbGAZXv1OBEpxZaZ75Dr/9wjrE1YnvXRWoNfCU2iYfwKrXmsW4bTmp0XTO7/DGZ5jazpam
l9hzewjQIxz0f7/Ryga1p/n1veh1erFt/nPUHqvTh/5IwVS4zuNn5wNIeDCszZ+0jdCw8icjID3o
Fdqbkmp7kXUHJnBVogrMu33chj+iAAM8tI9R3k8ERFcSc1Pgyca+kOE64hi43Zqyq1jL1ZKs1FYI
6CQU1Dajz/E0rQJzrXnlaep/0O2r6Qt4fvJD/GR0nHnEjLUoQqE4PwSSYskYW4Jn8icdk1AhvQ3N
WhXTifeMbMEMOOZaZeGmtjjNlsDodAhq+T29+FD2zmfrjXNYirS8fI69JhkdrNlftyFedRWQBksr
sLKuUMRsFPgtr5SV1yu5BdkC6eMXtZfmd5BZSBRx/2Q50c+DVOaeCDTS5r3ZIpGQ/mBzWMEJ9Tps
+3ES3xJ5CCVKg26sHoJZWpqjwzLQKqdIBy0dUNOywq3Hghr/s6qERAHg8u3bp7tA8MzGsVUEEeIc
0wOEUfdMr+AAxZDGZyP/E/LfTPL0tGIL03A0q6LTRTSQVygQ+1SOQ817TAycPyt9Odzt22y9mf+6
STvhoA6CI7JkKWUkyOqgSjTuT3ZIrCE8I7MIO2iuOKZcSgwkhH5HgSPsEaZqhmfRr6188bIoAnud
W35it1niwg51D18HrX+7SuGcB0K/vvQIgcpx/NYTxK69xvvM7rTVj7bv6wbaEJnT8JIgsPwyzjVd
eapzl2yStVCTdBVPWnQe1230g3Gs32AqkBsDJTsNqpJUuu0vNWqGPoNC2RHmO2/cKK/sW7IUE7PE
xeBlS/FdpPbK5NzP1fCHD5AeGvO4pbJEt4WYDL9DRMUvlwIJKywA5fosUauHcR1Nk3IlfqakPMam
VYgPX00yiqlMN5HGWhXYmq4f2xUi4MYkg8wmT+cqd/y4kq5+QWfADu3WkzEc191uen+Hna4pXAaU
eqCkH47xLRQuJnwPaLkrx/r3zhh9SCFDH2y5CGHpKbR4YriEJXP06XWtWW/yr/3ljZB0r/E5zdZo
tr01JuAWziW3cUpk1Mj7+0AJjqUsn3yhxO4IIIqdYuE/T8J7CVc6SPmbSnwZDki0ak2qUATpIJuZ
JzqFUQwador5tNVnfGbNN03Vj2r5XmYayLaUCemMXWI+jnd7B2i9ufViSOpvX0EerMhmgrG5GZEj
Y4e9il2kmtiDtchpP1jGJyNePm5Grahe1ouAPKo3pzbt0C6jAv0IVIM0nn3qgTgi03jHJwrFV4zZ
sLWe9xFwCuBNowwShOGlIMzafyGXi4ZQRnWQ+NPWnU2YS4G3Nn7iVzaItjkvHuqF+ePbpz2BW+uz
aQI8uaTYeQ02eP9pq6jBdB2BmZ4F/2TPVbLAdOAP/H+xY6/yHgtHP1imm7Hj6Wf+Wp8jQj/pvj0+
2YxGOdOk8NJN5SJRwFQDXkErcRWfSLn9XjGYC78PhTcoZXJnXik7nqqxSatJweAM6Q6Or6hHjLJq
3ddw35SYXHLM4vJPK0bzNURezcppFE+7Gc9G5CEN5IbzpCQOPKmmiaxRMktZB2pojb4JSvgJ08zt
5xxfhUo4rCIDrAUdorlr8q8mEDoghGDRwRyrKfveOCY9/FVqIomKw7q6r+1JwlDSkYRCpbwbkDWN
eDUOGlg/inq4pnOjAnE9iXDV7bO3M4GymDP/Sorf+YjCD4ymyH5H7F2FxGCUTWmeqhgyfy64mu4C
Wr2Ja2DmCdAIbw+Ea6yl2ZxC3lOm9bBwnpSoeLqAOgrat+S3ITDOHBgCC0j5Y7RUy1AoCL2hn/br
iW4qTUDCgHtNkTDfOt2QnWw5lZ8HUTV03nxdgS00rCUZXHNRRp9CJMsbL+QiYolnLUX0Y2Z7gCQm
prF3EnZfIo6whMlr84oF0wjUxvmcM+P2mBlh/BpSYMrx+1j4QrUn3HXo7ewB/gmZcZzXhdaCOhMA
SrA/xX03Jy9O+hZCvOlpZcpNxjij6ULmcxdOELAB37dXS8a1a91AdEuBN1CW5f6RGhxMOd8yFYH9
NO1Al+K5VDrSaGnr096KRQ2sBNBzwYgG/tYOQruFA1DJP14ZcnQyxle6PSEYmSQXIIU2tlbV+CrY
eiwlLm1jH6/FFZQJTm9J/0U0KvHqbBmmcCsxlBirbaOe6yFPEdwAfi5QBudQI1Qp4mJGT1Fk95TD
bXYk4Yf+gupIk6To4gMpYeCFghO0uEPgxjmrR7SEgj/w0jZjksz9vuU/Nla1Az/3i2JwLoFc9jQ5
cLjDI9flY52nuQv8olvrbLEf6ko2/kPD4ENZ8BgRiexL1va/CDN71ow9tAk7RN5q3zYKdJNVeQwV
CMiQfWIUTti2pMsyLbtrGKsZV1xpflW+RbkgoZku0wAHR2VJ86x1IMOQM7Eaaia+3f0jZz2zo+Hs
OmEuY6ET+120yesd1k1q42vdiuHPQka/1A5k/zz+51q9+r+O4FFkS0iwatt5IILQj0o7VJax6eKt
c9n0oT4uHVUWh301UjDeC7RR0UnPguOp4ImoMyAy2gxXvURhAs+DooryGAGXVlUyDBZYJE0ptDiw
d2Pp2ZCHJXktbqwTgW7oF+55Xwx1OyGKTZO4+qwSqqFLhyRcO4c89kbFCdgOM4FWt0Kg+66akd4G
/CnzSVcSsgOUTEfPMLCEcOJL468gAhQe6MyI0WWyOfHmmJUb0rvjgBHSzc77x7ALAFid1yOgH9Ib
kX41bvlJbYMGpIgwTncSu9fWW+jWzxWtt/6GdOx+jHk1OhFQYQ0HxJQuec0FeuhsyVEeICd0IeFb
EbK68s/RdUFcYkjiqEyytm9Qdcyq4oNZ0bwNzB98ZJGH5jcm1rPkqJ/Q9f54VsNruEyeWln20i2x
75qDfPXtsr2OrGKirMopAOCbwHC2ry/O4mDFQnnzI5mnlXkGTSgK7mcoOKxKLzIoflDoCUTF45/L
fCdTbxspafAUYtq9NcqRgqsR3sSdvhJv9XfZi6dBlljG4bFnMotNpTD3Y43UbhPcvZpKfCkMAxpI
l+NLQFQVVoJ24lYdhYWxgWSJCIQLlopdCb/goMSltbvRM2FUCRyfSbArZ1CRHrjjrMmEEqDFwoNW
OFMHZ2PEvmsHysgVAiApp4lN6T2ryuw1biJmj4aOUBytS8UtfmxlEIHiaBXfXeLhJJXCZe8HF3yu
PvbTxh5e2ga7BZcCTLGHhM3HgpVCw4IBmRyvmvR9WvZpXfS5DXahkjHjL2eZlzaPMLHJxJe9Y5D4
HKskyJSMGUBfGdayMcjrvm6Mir/nqrmCqF2DWGOMr6eHEnRItQDkqNFfBiZsVl+eCVwkH0Xx9aUZ
XGGOfl8K5Bw3UkNys5WURC6qbrN0TzPYZo766UtW2fvl+8XFNZv15JhstykC2v7SpZW8pd7J0uRH
4TbnOC7+DE4OjW+e7qPwXQJl8qucXwaUz7MawvWmm8uH+h1mj7dbuvsu2DnMQeV3CFwGpwiWvzRW
OwbhvcBVGQmxVymZ0HJi/RjJgBBgItm0wR9Oy76NEtvbPAwE3FrAyRtjGi+ra61MLwemnmG1slxM
67mwneIkPeXD0+i15stXJ1GlRgqXufWOfWDngGa/pTwaAR8CXU/7npDCniTWsOgTwG8VBhuHY+8j
TSH+6xPgTk67FcoLRWFer7K0ndvbO8aJftZeDfMFoGOADA5QcpnqocIiSWLLyI7hCwgmXi+MD0hc
ROpqfXGDwDwJ2peF3r7F1OtTYlwhClgcqIhGY/GoglT4iq3Na5xkJw+Bw/ZJG+IYYNvrG82juAVG
Sno2nOD24GE1FAqHfdmhQLx8oWDMoRT9dFjvg3lM0i2EBVWzm409702rSeZFnsaCJyh2nT2JNghB
AgzK4jqdHzGf8/+nwKkkxZNPe7A5zGtL1iVswxRpzjR46SYyByYgwXQyp3OmGgoxYfh6FMvawP/b
/ilAiDbwqhQo3KLLg6D0fJ/75yPfY035fGjwYYSQPZ5V5nXC3WJPccaNKjZUoVIgVI9SY7euNpRY
8HeHYehiSyx11aQ/cvi5oZIeoTK+yuitqoiqpkqovE8NI78ZMB1djjd4RuZALoCXU60kMgtO9oUC
z8n6DeEtVJe6OhF9p5BMB6weHf+1jBnKipw0w5DdQh3GBxq7uQnXP4iYAZg6E5CM7GzGcFJM8tgY
J8R2Zyc5qpBaUSBLJH2ENsLX/v4/rc60hmDy21tKrXhygBF6KI3oRG68W/WAW6J9mIdWomPa68Ro
1WH2aXeP+oz41OwoVcmqIhu7VPsISMM8Peag4yzUOkYtk39tjF1ZiVnrnwjSw8UYbvXKEbTwehBd
dbsPN5a257Ge7kjtuyQVRRbByLK8s6gO1mn5V/EIQVye39x/eqsc2HUnpNdMucaKti3MknqsgNPK
54LxzNyO/rLVm/ZU0Nf2v4fvw2m3lc+bNUgdPIuFkLzKAboLQlqq90DK2e27+G8M5wXTQ39puxGH
mvAL6fb8grmkfBqDOsNOxk0wGfxXmkt9Bc6gJcayDxTjIFyV1+Wj7tOGP2JE47uEaaebX/vJnTsL
Sx/2MFAEaPTsA6aPLif2Lh/0m62awFUJOB5MkdA9UAzqg2cRy0udFT5TN4zG1UQrIG9/Wuxsy7/Y
GLc4SY3aav7lQA1rDfJHJZ3vv1zcYcOto/e4+ClUSxEwLV9rHLYTw9uEbn1rFHCc175w7RunEAjV
od17Idu7OfMWVTIhrh/K6ysaQx9r1h+Z47DTcbuqUNfKTKi0XanT05TITVMZj9sGwSsJQH40pBtf
LiBV1+TUGoWlCuGTSHYy5H0U483w39HxJJI0Qn2988EQCjzsCesrXlTK8wa27G8RnYsDoQAYLfyB
t5cj0/zTlyeMQLvLe+0kjzBKeQVCS95jHJ743zkzr4K/kqCV+kEv8jAMODs84CzyW8OmIoh7vhe3
lIdglLkZKMFnLO/CyOikAU9o9voqTnnDlvmSlqu4gfwVvITWwW/55dQWwUEhd7qdPURh/lrongIp
Bx7aD0ts2MZeE42QZKYF2CWii5iz+rbTgnD8P6DTEKazMI+/cO9BxcVwllU/Ro8phOwHvSF96LVh
uglclboevssL/14uubPY/xEQaH7QKSFA1WPYDkrpmrEwS4OTtz37INVmrTlYgSSfMv6tm1euDLAC
WnKJj310Ev+GZMVktW5F/wLXIm0zoAoRRFGkkT0vaFDrqNX61SUyVAczuNBH6ZDrzG78Dg9/QL0r
OGr/Bl0nMrMaEXeIKJr3G0x0NID8eRDuXEq3YkPOulcgZjIgEeSxZdEJlDR63HDYp+w3Gj4jtRyC
Drer4Cf/POLyG851NzP11qhTROpq6y5qCZJPE5iMfqfmv8+Us+E+CClgpVKt3Rch9A3mUlkuAS4x
ypGqtxlOhv44aPXY0HP15n/Qa9zm2xtUbd5NnH0P1iydhNtjpZPsDgP7iwnexYntCjYl/lS3JiOI
E8MC78wQsa7+u4G5J821+rH+1uSJwhEkT4SRLGktjP/r/tT67Axa1f6mMy5MQ24FNHMNg99+Q9yy
DcqToMa972A1kvebXmbkgRZVmkFBPkfOZ1yTjY8ubru+6rDBWEUBwXbGFU1BdZjguJK9lyHze2jA
fvnDRFRAU6fJrNy/bh36saNWsmmSpnrHXBGUlz0/IQpeIZfpiVxLW/SngbH4XYRxSYYB0XcRwOn+
e3sq1hh2rFpzFPhVi2dKEmsRidOyZHGP5FeHNmdZyeW2XPsCpNiWQvLhp3PjzuRvXnwvVtgIvu0K
DhLAc1JRZWWvkRbCI4iRF2HSRi7pdCErAmEvSifisGoIgO9cWHu82ksr2NO5o4m2V8kLMzpMyeZb
BDhkGONTOjHvp4oHbx5rxqkYVvC9rx17ggwSDFi07Mb/r3x/jnsW2B7q2oBHYYQju6QRj+WM8ISR
A4iLf3FX4/P32FMHDn7HIAB1ijJ8EVVNRId4Uz3lN+DiuXMWnfLCiRZjhKSW1YJnK4KFZ25nkjJo
fkqTkKVg2gTpgR9kq5AL5C53/9nKnQCvO5ZQ7tt5OXtO/0jgTL+YYdakqLyJsusrZx8e5WHNdgGq
uMzdmow3S9sw+V1s61pOXCUcIxOwMuzHt5oOtoHLiMiFyeAcY5sBYd9EK7LQrI/1rRtmQWy5I2C8
02Ajrto3hKIoK1uDdljr8zpR+mTRVfpG+cyrq6eqQdZe7o8Ucuxy+ZuQhdIhlDVCk0Cv+TbJ8YlW
rJCO2oovCxJ9znJH4aagWi6Q8QeK9PYvozNutqGWVkiIZAcyzbkljFKBOytz7oshD9rN9Vg555xO
xD1FAm3evJgOBDsVI1qS25lvBgI/5K/LFoMph5ji5AnWzmtugKIR0n4IiBtCvui0FBITPvgSDLJm
UbwhZ/j+LJ5jGEpvinna9LN1cOVd1NEYfmduDhdVEsIMgSqaQCVGc/6UCeXEON7ANhYdV7Enbk03
IiWL1WhkIjX9cXjOKICT6KiWhz00B6vbEZzzJqPhp6RDDUEblQFTvLT7gsFz3C77gk3t16UZ4qa8
0PwmIf/qAKTFvXa7ihoWPUs6QwflPmv7lEaxty4pLtDXw5PKaVEHWsvOmv2svzDJkrN+m3vQZJDT
jHY66ADXwZaZISs5Hl0+UBk/YHk9UwW57hED4Kp2vA23PUx30BpAYoKWqBYJAxo2lcpmzTJh6eyU
LllXoM5GkUQDvKKtOyq5BeyT0YjlgsTJj7IHnFrdyYgV3EBg3ImWEAsL/xRHZlRBs3+Jaw9VZAqZ
CufiDOGc6IPrkK7zKnL0hOgxXWlno9HtW4UMNSeXEqMZBlUWFoY2CS+3ZyClcvv9lSZMt9c7ZM1G
KT9yw0ZF5NiWBdG9Ah7lRZgmuWXm4cdmgvWAk0mEfjCMQi/RwsfsNh8jRSVjOAAo87w15tdXnMcd
sp59FrQVS53BTpDZ1giir2hUGEZrQ8x2eRxSza1yPSFNVuokd5t1l1vgFvlVRa1QZHWVq7sikWK7
UfI/TRNxnkY4DgzOvFrnurBcDWDe+n0P5lVhFG7UqWoaqrgivXH5I/diqoDPc0bnktwHFXl2wdM4
vitkUurOHXATDQYFsMkwsGoh70QtVzlbM8mvQ0X6hHJn4Gznf/w3GKKmroOvFhe5eTZQfIoFbnRw
iJY1HwkUlpNRxJesbpqvw9RQrzphldGqag4/sFalstPiNRGnVYVS2mXnY4FPp0+baVk3GWpNIs0U
OMtairjd+BSmJh9nWVQH2LydKteR8rizJpEWA4j9amw6Y7T3ClqouKrIq75sLzXfbiHET2JoL+yb
VsPez0xUV0BFhRqQkSzmobym0MU7NXVOT191WQQeUY21fDtewLgLU0dLmtuFMItFxAHZxbyQr4hV
Q5nk4hdBp4LnpBIEhGy0KfCFdVWzzEQ/P1esF8AAfPpeGSCMI8RAaOfduFCr+96O3p8QQ1Mytt8S
hm83cOT0gsvrVxLqPFq84xwF2ctd/1iahuYGArCMs4jl1ruTMz+At4trehxl+NtM65fKveEaTTN0
6rRKdg7zrGZuiMvUeVI2MWfRgy8P/lLtnABa02thA8Yv+wsqs+9R7cPSVbsu8umCto7dLReD5KFY
mS1wfltjJgSEnK6N9f3uJ5vjPk9J/EIsdsidUB7vxwY6VWUjOaboTd/Gg/AtxJ4Sn+bX8Ek04Hcm
EYvuyfXURVEHFOLtFt60kF9ZeTXI/ZYWJNArJun907+LmY+1wJ2Z9WLOypi6TXJo+uQbs5kGy/Qi
sQz+3WaXxMIqO+BDUUmZu9B2LaAC8QQltWNj+yP9Se/xdCppiA2ir1o8DHFKxTHj0Gq+1Enkzssc
m0/j6jL0PERpbsXSBCs6t9VVUOlpy22iAi7e34eNGF+X15gdoJtwSyDs5VkS0EPJlyZutEPSzuK/
DFyI2OcGZO73nTxnDmZrYMgxdf44y+6s+ajd4RodWcbifZ/xu1Jm8jR1FNKA1k2muNVuqkeIrhHx
W49LkVE/uTveYxChQhVzMu7SrNkk5aWjuEJF88PrJYExX6bUPqvU4Q9YKzqEiT9XF71CDGlhVtpj
clmFy7OzEveauaxe+9KymuXBhPQs/n3EMMNLuKwFApFBzIt6TO8gsLOg6STDxBHBAipkKOCKuZWt
EfnMgyVjRUeOifDA6917gAVo70wHVx2VhT9cMZ25GN9p5X4lHTOS7acpmCbRg4Bkrek7XG6ELdqX
4z7knS/bBhit8eFT74CQGTQfVuuB9OYKJaerXhTr18SGOygBHVmwOb+EwB0XeNaIKMk5tHhiNyNS
64pgnb1mQKhwr7KBBwkDstRvhyZjmgUX8ZcwkcuNrXzJqm2C0nQV2+gQQu3kIKCWGWRQd3MS0u3u
qcpu0vxfH9jD5xlITeMMU0gDMubWhyF+lg9XA27ViTviMjB2Scrj11L0EXW9Sc0iQa2swHEu7qe9
ejouck9FM9u2Kw7xqDSooOt0sGORia+KOseW5eynVz+s5Rm/RbY6dfyTqp/oWrQ8ccLZO9Aw8j9D
AiIP+QXmTqGpamX/fWw84TMfvrjNbDI2+/D3zGs8MNcNKYDrFnInrMhaZn0mYztkxfju/YQVHOdD
hcWulE68AkMf2fnxS8ehJjs2NCKl1fLtGDAVgzyZMLbc4oyrDwwFrZCYAOUaElamBFfFojka5DWn
Nkvyj+iHKeS5JnbyYL/yf3TJ8Smj+JlNrTxtuGGITZruuYLGvsYZ9ue4mqqHSZbVH933CuhrJBBn
h363SViwoht3uwDxAQh3BDmuySD572vicOzYWtvA/NkTOaBBQZw1EbHrCiGqnWzBQGRgt1shgdX5
sPTNQIQkUiblGk2jIt1oX3Xv0VuLim4XxNtoCvoDqZlYCcpLsHF7CLr3KEWef7eQgdF0fplAeQCO
dffgbx9cKBaN2INfyG4CbNhzWBC0CN6z7WLClHoMHV5OG/McT8/o0OUqycKoTqyWDHrG+71HZhih
0iH9Y/4UHWnMapCETQxa1NM9e2S1pv3Te9E+2nB5zgOF1aojgJbCgCrKhSWM5K3gs2EIP+d4mRLU
I5zG4p8c6x5B+WHap8EMU+qW/fIcDqlUXktW7ox7I0+GsOGpAehnTe6JswUOYYKfTRvaxuKWA2gW
e4gF6hFzrSihVVFxLjbxR6BAtntGCscoerFlUrnsCt23pnJNTo1z1s5L4uIX4hPNhvM6gWD+0+Vj
ZjHUhbGLs8RBEfiFAFNFPkn7PKuxak6bwBqIKGIHkJEtxz1nNEiPmXQFqxTjYu9gl/eGJKe85t+F
mrq2h/M2Qqd8dr/a6ah/uaiQ5aYfchstWNVDUNECTl1yAgBI02XOJqw6OHYGN1Q1sSe7G38f5TIt
9dd69M3aM1hMHTaTz811Laudcxbm2mm1FFIlJRXrp9T4s0rFqd5tkjppE1jOZT84GPtGJOZj6Gzm
ObTvwd1bcp7yd79E7gGA9CMILGUKwunSCkJp1MPqsOi5dsDfac2d/d5in8vxGNWLHPtVb1mdPVrT
rMW5CHAZ3ghFTIxEjT8FGArAV7FsI2ZinFhhwwgeAMidswmAzTkDXnYf5Xx90peVP/s24rNrJlXG
kffiNp8GGgYv3gOkUBlhZ2kKWiAEB3aWgGzuVYFRqjbgxZe5dDzdayAtUfGfOl81VFnAwqcbsemu
M8xiE2nvrXquS51NQj3gjBJZOU5mCbNlr98NNELYMA0Z6t1G5CpsPp7kfcWOwAXSDx1EkNFskefT
+hlWYaWHcFH5extFJqxlOItijANr3S7uZiBpTfFnwG2CUvY4I6pEKgWdLDaj4dQKpi/CsrmepGtH
bX9rtCsA0rFlNg39b4iwJRQ/OD7snUfA/qcBjw7IE9o9MEOrDdquiMwo2AXuo5bKL92euQEHaE4x
IGel66yjJnxkkWN5k3sMv8OClYWCVY1q62O1T0pKNDYcf8jn2L9DIfFoeNpzzXrywMjaX9DkKXaQ
XTfaM2XEgY0t9Jy3B/wCitPP2trDVqOfEP/OMezjMmkWG29WBgbDD6l1J0oel7tb113Bz6fVX0RN
KjeVmLUSarELNp4wmhkeLlClYu+6w+N9cY43mdr1QGtir4E1v2lUhxCwJ1gd8ib3Xx68TgpPuxOc
vZjQ+cpjHvwXWsJID3VRLF8qaxU5pSP8WPpn6++3hH7DYxR+AfcChGpzgb+PwHWPX70RbG5mkLAT
l4IMmQE57BeUyVV1l3z4rbEmg1Hawi6tmv5oiICh8lOKIpRzfVZFONpmnnUsLz79Mh8jnHMvhH1Z
wkQ5jytYlJ9szGKTRS12+aywxqTeKRvL8YJO/dp9n+w/pi6YGPf+20k8TR+s843PqDMBereOJ4I3
Js52EPZz7XWJdL2FTr3b19DMoWRX5GxoFKwG4cnXbIOo41USlLnKDFExNjM4/PkEx/erVuo0jZcc
EJote50+HepJSqvslPu9h2rfuZY1/U/E8Lsmd4TNFhZgcyxHizj8Ev6iZ0SmKZwERrIz538fBBzd
57eftH6w7kVg8hsEec3N1BQWgcfG6059F5SJn5KcskVMwtcWYkCqfH9bjkugxURs7ePMzRSOrKKa
rqx/OFVnk/Pf0v7YsLMrZqNwONicJtU5MPY7TH/bs4ye87NMTo8XAVeGkATvMnq4kkHEIqtOkqWt
2HdurJSGeNz1l1fDn1m7SwfMrbAAKcE5eDB5097wlghN4xPBc+9rxy98hjSri0XbEbAVT/lwi2v6
7ZPOPkpvbCFdaTbEoVmzP8+hMgig7FgyECEAOPQd1MQNd41uKgz/iqB/rlZAJvBNZhunZeE7KRAy
eZYaLWKzY6xMUN5Yqficnd4de68JcR2+lFT169ksKQhbwW+Y1v5qNg0e9cYWAbqmFtWna/Pwmx5J
pFQM67KO9Ywp0xwN+KtoO8dLXltcwIZqPwDyj7Z01ff1DaI6467ZrQaxLiJTfjrFtyVXPeNdDtez
CjX91rzDoPKGpkP+88eEgftuK/Y0GzWYEAfi1xx7nHAl2mKW5ZhAL66CidYscUGLpky/3lWvoO6w
FfCG63mcAlMBfOpcXAiHf7iQ+fl36VKu1wFAWRUblXPUQYXCAGGE/MNlh0zROCGZwzmV+eHHlyVF
6dIQx2SSsZlKU+dDpRrlAx/7PlzS+9WDp8XZCI2dr/x3N/cuSkC1ufnPNOtxr05oiX2boaxaCYpo
hAryRGtp1NQxyj2yiL3eC49QKKQGn7YbGHUD6WrwqABMROmNZ/ZiPrCiYdq5X+rgMJ3EAQdbRZeV
FtfvKvxhXJ/2ZahuigB2t4wI6uc/VX52KnZRNE4L59gEoH1dn1h2mp2pA7Hv3id+XlN+I7upKjyT
AwitO9rM/Yza02+Ih2D9BHI9KdF5bA1kGZHXD2AT5eUN1q6HuhS+wWqRoz0mXslKKwJaBPDamAbF
+mcKZ1OP4nbEZYYALBNubfCaeYrRu8bfc819VxJalht1QNYTauZz58Si8sR3TuTnwlEno5bljLMY
IUpakyJw3ocYXEmzetZC20yj5SC5rrvMKVv0BR1KLMX355rarrrWbpZHYwOIvyoPsHtdoxVDWKKC
JWH8uqDADGSIFyfeL4yOtj/74r8nL7/LrY2+ql9yyng4oL3rIG02sQnPfgaqeLur+8cJ4e2GKhPO
qitatxeyXhjsxe4mVPtCjYCyjNv7cOS1POTliQh6+lI2eBv7n5aWcGiGEc+newwrlYciOGvTalX7
wf3KQ2rKRq5WKdTbXvcN+YGDYJnnBEH0mJfcmjY9mVWgZOUCgH+Ve37ecOCF7ddwaKucmBUv7S4M
Ow6Kny2gsMDb51w4x4K+Fdjfo/rIsBic6Kv4FaEPJv/l6Y2LcgQjt3bqt7Ke46dgUZ0/9aVI+Bqq
fAs9yYSOQ2AV8mBt/skHapmqryzh2Si32bA+1lOnR2XEZi7aGS3LsUMv/AFYolXlE7PNLxVT8NmV
F/P1KzayfHsX9G6uA8GeJEllejawAwgW6TkOxj6ocw0ksyHUt1O/T5RF4uS2tddrzslmCkRbBhuB
8SOu1LTiO15z+VMsfxD0UuR36ls+eI6G/mYotzijjrazMOEYEsKiVmBdZ6dIb96cyKPYfiw1gVxc
ZRfAsDqXk3uzYVgSa16e5A7u1FvmTfN92OdYJOCzI/mCaYtWDlqXETBOatWjs6/pvmEyFT3xWWUt
QnruxBeaITZXXaUlQKqTZpMJy/mBKGxF0w9KdG0GNukW6DMNAOTV2kKxT5Ww5bRNgIDAMaEmQia+
bAH9eXHyv0bJMoMCdSFMi0kKpHKzskUdl5QoSLvXvVcZueodjd4C7jZnNldHCXIaBP5oA1Lxbq8n
+mMY2k450cTzAzoCb6tdBZJ7hYj9dzZc4Xk+EJK88/qSFSKGadGlClxWQdFcxdqsnwMmj1y3y+jq
0Arkwb+xmtxk0qZQzCZqnh0faGJdvc601hJtqGH9MNEvEsV0cQhEy8wM5BK5ZdWhagHzT1yJoPyW
b9vhLUxDqAnzkDO4DTTI4/ja8LqdBifGqGQFGGRNMNhA2w1Mwfa9P4NmYXo2YZ30f0I55r/GSAOw
//olVExDm/J5Ol22TTsLLvINhmYA+0pfyWxcqCbq9vzTAN2S8Oej/LqiBzfbc6lKVhXEweHUnD81
fW8YIA3MJQvHnBlHV0+TXzczCRH6cWY+hy8pJ6qWQwe5wEms0I9b5Z/xedeXLlUeHJmDm8M3azTe
wRxQWvgET2svpJfKIKWEfaVn4K1hdPUlTq7+ZcQyo9cbqbFXiQDHskXA6+DC/IcvTJ3Q+TkB+QtZ
yAsAZlnjkf/gZvbry2kodbiASSfYNzcjl4zVD9rub4SCpRKCznU22s5+st5xL5WVyphu4VjJA9Jx
3L6rqWS93R6KuDP3778NeFJkZrcEyB3WMMsctFLNj/ehcGsoykkEIiZoVEOy+eFFAVvMuwG6XGea
7a9miPoZQT0ryRnV2yEsF+spbQg4gB4FGgh1ZfryFvncuIcIqpETiuAwqR+ahv+tNhX/1ikIZaEU
0hvipANQS7WoO2c+Pf/iMMNVYZEVN+yLBGPIDrP+gtb57ja54w6wOPukOehNmQpE808M1cjRILLb
Ptib5WFQAekoQ4ReopP1OqtJ7hAW80O+LJbNl0/V1UIV1fKwKUmFpOI/v8bduYX8PNTyHtYVRO9Y
1qv6NtMXLfBJapRtvmXHDzWii8+0StwaWhG0HeyTpsQtTqQjvj5aDtctElrwrUkltKV+eM9bWWHp
5daZ2w6aGvUW9FNqJPb51dKPtjrdICGE9HmgSY0hhvHl3UdwmG6S743ZtTh0JMB6UkFoV6SMIZD/
pf2L+YqsQzZqMiHhN3W0xuNv60t9FNrVHmqk0HkB0kUOaxHhImNPv+Ay7IPPxwoukXAPeqOlk7D+
v5uB/VsFQSH8YoiZYBmXxioi/nGPRPoQo+l/yERGenJtIx/lfkD+lkFKQsrgSOP6T82A/avxJsJB
H2SNV+qBeVGjonix5S5zHvbTFhcy1zi0vbFr7obUQddooR+glty/adsk0SVJIwzc46sue5op20sd
RrgziHOa+5w6zjZH5p0sys3+OVU2W+ITv0aiDTwR4D4tFuCO9sM8Qj0QgV3Ruauec1fu00J5tXRm
Ly14HgC32xj11vGXeaiB6UbF1BzRzuZmgtxgT05207+P3AxQ38Gsu+Rb1xc9lA77kAICStxod+wq
TOAYWw0WDBfZLbqiEOaJRpTal14BqvtY8FeQpASf/VqVqH7egHQfNhiThBOARObuMWhMgb+3kk40
p2PovxoRTSXS/NyiYbyzyFmb/EbiKa8dCCIjWC6CpyMK8o7l1k6g1nPRfIT3qxcrN3LFzAiKyL5W
3+6LqsHQbHfNd6jLYbJAjV86mH/97Ed6/Oh8pfrLW1O9gNCaiwyeU8ICHfKShd6rcGgLdPaiZvaQ
ct+YF6hObH0g2XKbN4dB3BhslayJlLEbQoj32vCM7ptJm0sVs/RMO/MS4s1zVNEEh5ozIMHYaCht
XGvM25i6X5r6nGDn1Gd5u8GT75+8hekS7mkjrWFfCS6rTzMgrWsbo7BapWPB5EEluMptYgLCVSXW
0YrTRXivS2uHIoHyHnd5haVOeKmJ98ZEYntMiVpej1iiyI6lyzO02wiSbVwxNjS8XCBLMudBoeRF
raTf3FgZeB+EWQXplYTexr99tZuaAL5aouNXuTa6W1qvxphvSqWKur4vJ4/fiH7bYDK6svrfQuxH
38Dzb9plT/7m7bfszdGdcASk2d0iTUwpdI1LvbMv5CePtes6t5X0Xm06uYZyPxi3FhEYcJwCe8vU
YPT5hBBd6xcuzVPqMq9Srsy7fmHLHdTFh2yMdmL5d8YofFJtgsre4kop/+gRNXiZRzfUh3qbaI2E
O9XKi9/n2TCTjB3HJOXgQ3Jf3h9rsHjI0ubdOWIj1z+dSDQAT9DmXpRzhwjB4qaRtEZ9JvAAim5x
k3NZVBw247HQnTkC6SZrYU1yW4gLsmFGrlFy6buH4AJxgdEpHWc7AiMJWE9sS/dxgT0H4fR8HltR
AmcLBKnJrYzBt6EdZ8NbeSf2BKZ7lWAelyqeIyzvk4bad0y++En0TPPc+dpI/xBX2iIl6ZRE8P1f
cO5Meo52mAjiUeE8PLrpNQhr/gPB+1lwahfSia7jFpqNeZEn6pYLTlEZA8M0UUdLUun1fYg5/Ubj
nUJZ0hzDA9LcdXOyovps6hDuMTTII49hS51BC4DCb58FQkK+6YYdgqAWV/uxdebAZhjqzETq37rR
VbKQGTJ7boDjT+5xF04uGVO7uC4oSWiRFY7tcjigGrYWAsaO6by9WfaP+ah3GAf5kgs/7mHleVny
yixfEJTSuTkTyu0RfbU4fOcdoSO44QJ/n8uJ8MzDc2EK7Kxyp1DoU8JzuGuXbyH+2nL2RUsOFG49
Tgb9Ve9bq9Ji3bu34E1MNVLeNmZaSKt/G7irZiEf4kI3lLfy5qeSFjgJSEwK6tQ9NbILJvaLrPOR
6zTwKSIhieUwTVBwYr8Dd10uImGY3o3ghghmIx0sziqkV5MpRnJdDR+p23anJC1Yd1mTL9uA+nJx
GX/hdB4iaj9ry3fi6OG/tDLih/iE+XDjVk6G9ZYcqQbE3BRZ47slT57HWdM5Hrj8sdjfXM3DPxEm
9TJTNG+dqteHVvLhozkwwqDLJv+IwYljjzJffsg2cHjik1fIILIv3f3g1ukr/GFA1DypLKRviAJ/
pE0HCzpQi0VRPn5JFyEC83dz3ETQJ1UMpiZYzaywCruh/NNMCglILoBtHmwFaWmAK5vf1Pmmvpdc
VhRu5ynt9U4u9MoER/MDJpJiPHtZgqKUPl97C0sqqFKKkeqsFk1PJvBZAimHgKa+yP4bALBo5IyD
Tdbaj2x/iYEGroNT+glktmbAAGTXReGLDRNZ5E/Y+dLjVH+xtM7pf714kDPxqg2Uaj2TNRXQcdtH
SWBosSQVpFfwnSbpRCLhBr+QQLXdpHVSA0LxvHYDfJI7WVoQYtHrbJTG6ZnTBenmOPvqM2eTjwFd
icZSBjGOMJL6LcFpfcAF/4mHHNiNeciH9BtBRQNlSZItpSkX5eJOeUgkYyqR0X8yejgCzcXqUNqw
EBF17HMoHVrSBUDazYNb0Ss3ITHJ8VnJWBYZA0ERAgwALyB7HB00YyFz5/XsPldwxLZO0M9lQxq9
wG7pB+4ndVSOOg5N0PSA8+eLfBymuNFshcawBOALXrTqghi1vS9djdEwynSiw60YziLwu4chWelL
LhFxmPcnkN756HekUgOD+FS1rwQDwTHnMrabKdlq6kprYxLJuDLg78IoOKGPvdCE4fMPElp46snx
dr0wJxYzyJO9IwBPaPlgs9lYh0GSb5kYQnkOlGh0TQBE1mPTZvlEWIqSibf/2YNH+yunQfZylUiH
zAV3h+qyUrf/380bE74Ok2QwExAj41VmXnym/goAFA96Ns8OfVG/lPvLxrNFvvOPV93803WeIpL4
yF/6BJYmxt9iZNSqq/rTlr6qnxu8Nh015Ar2AkIDTKFfOmT/P6Z/Bw2dMs0LYiJTFqH2baRt6waq
SPMcYgJg5fgFvaw0/UrtszZwj/n++k2zP+J8AMk07uIwe/pPNpbDU9gV1648whaol51TJjaeyxcA
FFa7VbIrmpX+tDH1VduKYZDO95wqTf/UdfvEXdalu+JebbI3C5Sc/Y7qseZL5DT3UhoKaLsLxfaT
wHMgsKG27cR2nsAnPkPTxAiZrkfkKD7o9nlTACKC05PctcguzuSMRPHiS9Y0xA67y/LJHajT+pTw
8cUKaBRPyFh8+PVHvvs+EyhzNmFM53bGXqcDagNnwUzNpaHp19+CiqPDu3SLxB3Q/tf9wEj85B+n
jI8HJYzyJzmKrIxS5XTOSLEylSVz/JzgilV6n4je6asG23W+/RL3CVvg4Eao4FDg/P/l1tdNT/Nk
RZEPHmK9MVLbKLS2qq4uVm3Fdc4Ifqq9g5929ozDC769FRz3L0Dpgilm/IJkz14fLUQ8ukhPbxeq
0hqwqqSaPyGhXpZ5GvISfLwr3maA+ipD7JXnIVHkwQu2gzNOz7QrAOYMBe+ywjwBqFdaiMjzdx5p
NfK/ozKdO8cbOU4vY3BG4wctJAPeoFpCvOCvLVStzX1MVC/PRXeEza0mXYB7MQSDl/Q9y9jhgf3Y
z+BUQXIHaWzV+w/ajD+aUv3Df7qiYiJPjafBMunlkM0SeJsoYIj5aDRYtYpBLKcg2rZS+WjQCOnQ
Im0Yv7/6f7wr/HuN+QRD9BeMqhzOcv574gpVrBnXVwrXSo7ZUqB2gstWYynsZ9fcz8xDv1spW2jp
GC8BeqHkUzagNuX8QGBIwCMHQj7lCWBpjrUYVfrjMBv4q3C0aRhk6uOntjNSMcsqQcdAuODnO4hG
t4ZNpISRDMRmpyWaA2nRIODuvXGRNwm9gUQ1sfTiEy5SiV5v47QE/sCjrHPYyF33cD+OGrB9m7Ab
EJ3FPFKfvEAY9bmdeH6/61w0APgV4/tYndW2n17jBvn2SDaL4OyWt/fT0BaWARGEvI/5C/QyTMUe
eFsznQnXf5NxB3BHz8dqFJJsaYS/MMjwNpoBxBv8je1T7JCjd8revQrqQassFQrR12hGe1KHdtDf
8eIBSuzDWRua/ngUS977WpBmav8NunGkWB8DIN6RlnVWfJrVP+sgEFWJN0A7KZD9wzAF0vK3Ny4Y
Zx1iOMKcW7wfAoPaAp9d6RWWFq9iNOXdT5FyJKiYIDKeHzNr3krrzFTRA3MvdRSvSpie78UNESAM
rnJ4Qp+xToAfQItyWgC0lkUppwR+nZwaijdInJho3hCBXOkEo8X0PbEUaMgvyy1wzP5j3XNdpxap
cxQwlwENS01tOk1JAZIisD4tTGGyq7ANJG19myh6NWJI7pMbGzKH7OdauFUeP992sK/MUV0ll4n7
IHNwjRb5oGdyv8AidMb2dTqApYkU5Lo3qKQiiCnKWltdWROOY+mKyfAc1jUyQlQwtSXehjV1MuZV
iDp973oOJzCHCiwPQ3AiwqdOwcu+A43HLC2OhhyzxFgThw/y7LPbxdI/OkKAeHbf6gy+HJ2ecLKZ
hXBhSfE7ICB60b4Ck9YTuBYOqIQEW+Elm8OXG9Whe8Xg5KIyE/gTDOkbdd0A8nHDCxX4r5GXlnc8
dqAcZmV5DvO2h+l1FfCy+YTzx9/AtIEdgr2yUgL3f+0z9k7HeDV0VwW1+rOf2GG2aJZmxy2ip8KU
ASQRf6szXsLrhb6FPlvQAhK1ViVMPFLK1f3gbPNPxvtfjbTsgSubMwD2yiZWErfsRD7HiXWwM2Ny
I8NL+EXtw2FIGheN9ZTqDNtohWJsKIB2+fTmFZ5cBuPq+DdpZCJ8X6NQgBv9hD1ALaqnDjPK/KGe
8X5pCEkM5ncFKUSZQ1n4w1LwpYvT1qS6lWkChHe5r82BPwaTqFDlAD6K3YY5/do/yLMZVRrByfFO
tUkaiiICAODgRT07V+gVuiqKXaDCXn3NDQovMXPuZPK65MHbUHH3jQvT+OKmDEfrduQ6mkJs7cgJ
ECHh9j0rU1SNwPUzERuurdJYtPU0XzxvR+UQeNxDuWbrMbl2XvSY1ZLauN91LAmrXy6vPuMNF+lB
E0wKPxLaxwapBGHHhFy8A3YQq3pqQrqq6uHAM28GUUvtEr1j9OC+Ns/9sUGQBd5KKmzGH4yE+JfM
ROGdIvFCJ/s65ErIQ9aSaJhSJPSOMXvHO0ehGltY6grU0RYNAblLZRxzsnC6JwAaON9KRmdQxgdV
oymewYgNMSw64kgZHpFXhmu9RwOswxI+LMapKOaUwNWwZXlMQw1GiAkIaixgsx9i8TwQGN1vp5Aj
fup8mfiQff7Kd27mdIUuxIrmbNGZBLNKT0kXHLPYW9LqjXGdUxhJ64nDSaNI5YU4b0Fi5RTi6DHm
opS84G2vn3SUlHV+e1ZaHGEMmvAKmlCjZvGygMRMjLfdro7y3TE093wFdk+ak3HLNBAHX27ObjA3
Tl//24iZ+DqHsuCt4tLYbKunk8Y9gbn4o+ECGWvCudUAv7vmX3JMa0cI1yeO6vkrEL7zm3mKQI43
PN0fKvWkJ5bZ7EM0SHa9Yt09fyqtWflqoQf/T67tDEMtRwcIx75In0EhxMgh3hyB9B/NEvAW9BY+
KmsB0CQf3x/d65W663kCMiAD2X19a+CgiKWBCHZ9re90BEmxyEvjdhIZhfXnOdkwhistSumumiQT
WXcm40hR+sYFdH0X2WE3Fm7OrjqAvvVvWObiiKaj94TthEsGx4jAxsLRrkZT30S08fgr+llLxWzl
rCFDcQiN3YJDu9Ot1nhhRvFk+liZcPEAUxHMUW4ZjGGttw1cfm0FHuX1aarX1abFZvEaN+ncTaPZ
4GMgvd0XWAQPljUnhWauTEkrSTTOx854ycWXfICNKXbYashIPReOjGJzm5njf4/Sc7td1+IMaaz0
sINRILI+ozCFWm8/owHr9g2ATiUk33GIXd/j6YlA25N/fwoO7b6D5vHfHsdAZ6MdQbayRMvRyuqm
8nmaspcHNo/5u9y1qZeJ/OKVTXDWdDZmwV/J0h6EKv6eZBe//Xqdk5AVQa02dSicm46FmI6PWbxU
2y8Vd8+Kx3Z2psGqdOteJJvLYVD4QC5iXogNox66w1klfHKo3OEOtmnq2n/wWZbs/BOZDsjjEq/8
B2dY8/scR1iTO1OvtQiP8MfNTIqbcCFUd2ZNrp3rB/tb2gfYBPvrEIl2WCqiO7MeSLy/svmHmGdo
xQEK65UOURJSjXSuFf9ol3twuz+IxgtNv5E2EKgEZgctu/hP23bzj56iP9CFYG4iCnMsrIN/eTWX
caS2iXaaCrIbscP5UHFgMCEyUORKjKrY0LeFuoezXbXipzBPyxMFeAfur1jU+VbXi6NQ19WV0QLd
C2NwBuDlqNA/hMI/Whlja3E8vdnlzQ1e2zUpU5FoCBr9W1wJ8TpI79ts/6FX+06mOh9w8egXJ/dM
eonuDOo7+aZgBJOBxIxwO/AgduUO1irAO6eshzxn1Z3mZN3RWqW+M/tzIcJpKM+PUyByvqs6pREB
oGhFNtv270JsakDsw/Qv6Q+Pr9RoIOGevya5my/sGTWAstYKHZbYkqB+xUYnSmsYZ1Ngl6vwhmgF
ZBxWiHeiGbte5AEHkGdHWH8vpKozgD0wOUMC4ezLURS4FV2fJQlpT2jvjy4IK0ZMJemKEx8zox+U
JkKPNK9Ogn9lxY73JD9q9Yb+KslFQJpJ8R+3CsIYPMAwUiPUiVll20h0l8+mzhbSqVgAT4yCk3og
woVMKQUkx6qsollv2pbLxcj9IVoVFU6IpJpRBfBeF6DtrL0UjaiQ2cukpUb5IikoSM+q00OOAyer
5f7fGQMmKevVUEZ6ppSewyi4xkRuJC/yY7FtWx+/79/Tbg62XBU78oaA8+b1s4lyZeTuD+C+jujj
xqQVfcnNmEAxFW/CXeM5rkWXsIXHmELDvhhlAoPltYu9S9U9fqAa85c/5ZVr8bUTvos8eIyBGDZr
L50ZIuOadAyBBssIIc9tclCQvP82nlkf27hDW398msGcglOcSbYd/XlrjWErIxQiNErwuqtGWwNb
fxeAgvfhdmoDPHiXhqKBmrzJASZ1vjpQLOCeiu56ei+7wOJ0t/fkboOb9A7XmjZhkyOJ0aujBUMi
PJN99KAYT7Mw3ZpKQZqUvsar61DeAYC0ljZ+gqZWsH6yVdvnaXemcD2/4D4b8nZaI0rbQ1dCYkKG
DNmcMHv4kQf0TG0Hiefpx8s/se6SbMGbljuzKKyMqnRsDI9IbnrpyvN6sk3+OXpOl5IihGj7pyNk
mgKshX0K/kNyShMjaz31wPxhhrOeKD5TLG5EwLx1tw+0D9AHR/jk6r2G2/leJ64I3YfoBm6H0ufO
amtgUeFb2sW6VwgprJdHFt6BA76hnHyptZxDGqJ8INiw78LaxAOZE3bAYRgOHdx3xedBZ1PIHdtZ
zKNbTNp1LnJKOMostGAiE3AEk7g/wS0qA3xsWHWFmgLFT9ZsNYjx5GHAY/KEf3HeU/IkJqnFbCBX
v7QC+JpkwouYCXPyNfU9pO/IBDOyaBF72/rgICoaZNND4TMBF+2wJwc1ZM37IVBktR7P1cM/BQxq
F41QbO2zWCSign2XhvfTV81lT7rwR2cvquOPfEzoME9DEqXBbEcIqPv6MCs9KWWfoJK9g6cqxM48
v8gvAZIGobv54yLhgyizcbgAc5R8b13HJVxraYCJkqW50GmS6H4QGJiyA3RZFLoFI6mzdaaQ6YQM
se0A1JrxAtzfN/X6ravlUEhwiOwj3QaM96KBITAJS8WnrhDjJqQbkpl7GJfxWDkku98UA0O4tS3i
SnEWgRaW6Y2QbO7fixyUHRH46PLqo8ex9/aS7+snEUtDKNUTW38r70RkiY0N5cwu9JJqKAI2eV5M
9S6Dr8op+6NXn17IeckdGClDWaak7xD63UQCa0lIsnkckvg1a1XKpCKcM+x1cZt+8X+xF21aNUi/
frklGFpj9cvCkeVrH8dfLe++rm3kfw5noqdF77+YyXsZNSg95rsZEu2nzj9ugbpjZfcsgjkJYrXI
f1tXAle+zzSwdD1a+3HdExr/djkKp/4ufXc21CB25aSFkBOCL/sRke4Egc8thvmpfznxUoTpqXzt
wfIWUDdDfrto1+tt9jwM+ExRIzmp/QBUjVqhc/JAUK2wkOSR5+mkDV5b5spT4WekG5ydDFZgw9zT
nG5pMX0C7DQU5Zfof1lcwxmxcEyee22Y8vgcHGwydGqZlhSIQp1niEQMCAh6WvgbvNF+NP6PUII+
C37Dtnxh/fbtqOrD1xDdqYPIf3sanguzp6+wX/bHsIW1qrMoJXMQmW4UPlJJ4RyXlzYs0ii4DF5y
9jD03VSACW99/nPznkhp2YgMv43k0767r8vWsPa8x8jADnUSH9fCJOQTBdgcNR5GpcDNhtpqe+bx
Bc1A3UCuSumYwC12BLc15zmlZ1OrE7vligRXEGDgRCf4pQ54xNtR0sSPvVllo2miLRDDtA5REUjP
uyfW28XwUpzQNbGjIZM2qEk5PWBKq/P2RAIM+D3cxRF0q3Oxh5Hhp/OuFTXjk2/2jt09lvU7glTO
qIMktKUunzakoAbqacAiDDb2muUHDnihcG1mE8E0APef0Uk3dg1G+cDVPa9qJkhJAtOrnRGvq7RG
nBkmDziVAfnQW1AOkByRIraQo+UrOcwXt33F5BWQRPtq/CbSPtQ00mEkJauP2vFnpm5RdJIWbuhP
AVkDDA6gxi5LpGYwVOF6ZFjmbzMVi2kEsMVE0zVRImu12J3F7keguMz71G14Mk8LyV52NqXPhlO9
Jg4YSPPJL/tZDOJxaW22t/5iu1cXXiblSAMCuDDl2ecTCGLTqfTRsZZSfgbZiqL40PQ6rwnPL3Jv
MqeVWs2jcs849nUvF/Hjsu/bSByh9ZnXi44F9ZcedsliOr2mEpZLzFI/OAm/t8x2mG8UBs6N+Y0E
7rbaRFQnNE1kxrq8/A8mDrRal3GeVOH1ZJvo8jDmm6yiMttAukqhIhaHB7y7NeKvVUuAbELu4Gv6
5O2iynC9rKUGY/SByLhM7wq40YxnX1DWohXZxU6RjIIE2QHhd76D6UP58IDPIr1D6algikzMB9K1
l7LrL9dl7cbB7uL4YOdPw6R0/RcutBYNOBGLzNtPSlzkkBwWJ0Z646YCOVPEj0syIaPAjQEyGOOb
65GBvFpucOancuTIFgptuwJbTPXBBA1Hzntl3dc2WNOmS5X8GD+UsLShFe36ls8rdoNxCeFkl3z/
JPC+KMVRQXJ6hgkrY3B3WV1humYzXl8b4bdGQuV+5R71rxBDx44xAAJtA0bkOVoy/1c0Q4SfPElE
BMC1iDHJOYTeizE3kCusvhl2yd6OMcjqw3yP2lmd4Lmrpj8wuKNEkaXTMtCRQSHvb4uARa9aBTSy
uuzA0UWIDdQhH8vhMgy+yN4CXbVQWm3raa95s1iS7hzhigXmFNT7Wa6VMxp9Sxr+tpD069Qc0DSl
Po9aTU6xW3osuUTGeKrbovPE2BonpQia4sekPSOsmxlTC6lFHRSRRgFGl1aIvyfv+8MZJjNCGixy
FMCypsD6UA7eEc9mFjgV3Cgkdaqvafqw30sAIglZLYfCDjFcsmliC4/LcoRy2it6ZIrngrOLISdV
HpabHNjONd4QZcaZrBnErgMytYV5jbvtZtNLEnM06vA5nnQ2KkBTd/9JtXE+FF1OXG3G8+j2gPFu
AFa4br+FoUV4/lAPxJmfHafdHqKYxFcuSy6pfiuP36JFPrfdhFZf5ZXuowSqcte7dp8OJEP8O/3b
Zv1TBerrprOG5G5UT3OFnIeV587R8IwmIQKvZVaskXyAqWa9wMLGbd0x7XS7O6cT8YBJ7eXFmP7I
brjK7A324SGryE3ANza2kgRQoeZHvlK6xhzd6ZfWDeOQMqdctUothp16gRGhc2dIddoa8TxZurC+
tXLiNkmMqt+59B/4T+wVWNUyv64LtuwhSuo94LmP2oYlo9AxEzebUmkeOgQsQX6W/G49gQEG92IU
rGSzIS37SzsqntIC6S5KQY0f9dZtFBn//kml+9sdwW0spt37vJe4c69awL8D44XeQk7ecxxGHSiw
c/1lzeOw/mYcxO0OJm42Xhl8U6TM8HY3Y4mw9bPXFBMQLyUejxJRYHyovg0igVAFEVG3P9DUxzGx
FGQfgV4mcUxuf2SYX9osRSgi/OKinNpmwlfjdJBa8Kei+dUcrLI3vUIbWit3N34yRN5Omn3ScKOA
G7ioJnWVBN0v79tpKqbBmCQPB9A+5T0Z5bpjc2DXPgJdYG0tGpTfPRGpmU+mFHXTVmYZVjxwa1K9
1OSovG1nKCkrGMMBVLoMOEiYEx2vL3Oto0Si2mZtMUXcL7jvty+VoH/wxkAYvzfrglxOvRHLaptF
m7RjvALZYYbZwy7zAXXu9tztxN2fYqe9kJZIvG1zv+ukuyX6LdlkLlxE1i1ewBtUxB1xY+4sQDNr
3Es/FDV/a42oCVMY2pzjzVss6719HDTwqsjHUE3carR8jrNcvCnzUqlkqm6KpRBplAHfw+3jUXuF
Y8Z9xdBsB1g+Sf1eTKqC2XO1Rmmf1PLrNNp07rO5HSzuZmSdqqW1MEaLEkNZzkJ8t1iUKG/IB6a8
SEPx05HV+W2ESI4Q5XYeDW4aGk6DOxJN7w0CKFt4l2RTaKhk1T6qi11S4IYcQtbQB9cr6aXvj7rg
nuScwbCm9OJ1YUH8JyFljpoXNigofCKrHWypd2C4C+B6XU5Lq1c7J9SgOyyYic92l2ahEoSIRGmb
r4OcjKfMVmneXdiormGYXKhPLuWcEx1QkPffB/5pQ35cyn35pROzZC39Si/VyMZKSGVGMSBXMVAI
PT7l4VsquVoltoGnFfEqc8nW7fC/iUUNPIaGmgWlytcV4Ksy5a8ja4OgbrmOl4sbweOKlVAnJmnk
XaDiSFNEK0AYAgs9PBOJ3FYC8ahr+61Q3n04YGECPK38llXtrD7GoPoqGqG7E8nsT11W7hUqsf/y
C7WSUQe/xvEKTpalV6JxxxnL7Nz/nqq/C5k/Pei2gL5wHo+7mqMr3vKqjRP2dW6i/n+ircr7OXjq
WvKdW8afCQZ4p+yFE86PX9Gkf+iiG6MbSv6303GluIpsqeXCJcTWDq0S9KcZVwpaE/XIs8a7K3b9
MJasIa4hXQuQnxT6yvlpP5axHb6ApYV+iYjmvsWDJSgk5HJp0UZFJnXbyXIb3mC2wpxqcmPriYSS
fQBF1tjuO2NhRc3aRMTbofH1MyR3w4YNRn0txNQE9wUhz8W1VDE/kLlMV+zRK9jKQLbMtmMmdIpy
AlDt1Y+u+sxRxJQJf/A2HEUKPx2eKwN6Y+ypR5HLLUc6vwJneWx4bGLrw0atWCjbiYExUdbp1Js8
q/rIVlg8gR9SOkINj2mSJMQ2TQIJXhI23qeA4JUPbSr6U76m5OwcseLDuI9rWFQJwicZTYSarZ/I
8JnRzDu82VT6mZLnZpxSOFjIbjlLjmo50UIG0aPGfjPsK1MTcaP66/qxlJzP2wkO3r7oiIaVaT4R
9MMrfXEujDDhPbvMwZaR10DDwhL2QlAD/bS6FotSiP77vYoMSel67qZGPb57VRB/V1mEF7ubpLcE
0TAZfiQD4QYKiMdzp8p5lfZif22Q1/3W+Bds0rbzZbVtVst+s9lPH2b7dNR4HtGekSCW3wVW4EHp
aMcSAVQ2/Hpeej0frhclZHITy/2B8WfG6vHzXvO58PhtEvWDVKkxyV/zSovyyc7Sj4Adnl7d+zPT
8wNymlv4m0Rk6ldxHzAsVCkNYLDkgehLgzOrbmwT6jGAnxGVw1krzCww8+rS93ZPS6aw5L6X5tr1
dbWObZRcOq+uO9CwZxVtCGdrThs3/ptcxqJpLtH1rOOcgxGQRAaz8hoUX7RSMGEj4T8vNqylv7c5
ByfSylfzNzcccT8DNV/5LxpqJXcgTVKQRX8GC2foYYg4oYZG03T7TabUIkg4OPgXsX86U3Hrmuld
gJdXCCgsIkswQ1zR4NgfpayVyu/WsMBiFiPBFJ7Xnjk60e493HzzaHKcpPbkLLV0nGvcc4t7//jX
n3P0Hucj783N6oZ8P5mhaPpFLMefBfkGqSkqnfed/eOMJ57vIO4mS9L/E+De+iZrX8dpq3OOLVfj
QTAPvvkwRPiYoBFCFmudtexqHVwmDxcWCrgi5TB+KciygwZZ3FdIWO9i8zOHyMMy/CZyCXcLF/Y9
ElsdYwdeo2E7sZ0/646KFQnAoLaio/erhyW0CNk6zdCQx89VyWMiiytWuzzxyqLjE0WmgmffACsz
a/U2rZf0TUwybtzvECmWGL/7GDDmaCYfvvsFOZf9CXC7edRW+USOReeu3u+huItBIHKUClStKrkz
b+SB173x/NksZ3Eg1rlVIHFBGYxPfHbVH+rKLlNJDfLICqFkR10K3Dmysyq8JPSfQIaVd4nP1FW5
WvEwSSrhrLyAfCEGjNmIUzlLS1XfJlwFHE6qAOu5PpBIwXstCUVsznJqFM416wORcMZg8TSxBVQh
ELGLVvb/SxdKeRKKE+XzsRqHf97NuE8PPYfvZoQOEP+bDMX1u2eJ7KG0rfBvBP/5428moCvCADSN
17S5U2bivvftIa/saVeOr4pWo4iFzBAuZl09sE/OaN82rq5EIb9rzmqAXeFeXGQNK4HlR7qjor9p
BxyXQUxrOq3Oci56schSNDa07UsI75rJpzMwC1uVbNwc7Uc6Y0XbNj56gFo2xxN06fHcJOHlXWe7
bIlSs+Jia5QSKCR0t0y8oE8PaOqx0HgfVJwaRXF6jP9neaMTY7T2pAv5yCVGQ+nxYZHDJju8w3Di
H1b+8yqJsTEtSXuZMy+cmF2Y+a1pkxWLsXx0TMSXKzozWuQ8kV0xAkVEzJZJc/DX7bRW5YR4YA64
9RVh6+ndvidU8ZsXugDgW3dUova3cFkeB9KAVt0UX8bNDg/fYoL330/XMfdzIzCQtBkIoCbC6Tdw
u9QirOZh3y6PKt3tCf1qUtUlbykd8edjq9V9pIPddgs6wnVIz9oe2G15oBBgnYrTu8B3iCqbKXbX
hSSitUd0zOzAuErlSOjgIYtF8kgIqCOnWXbJKqTBdA8NHLsATrVx05VkOrKTqtyCgV8dkUtB+nif
/ldm34SiwaO1uYIgIBmo2aOQDEinIjRMZPccKFoFwRzhKwXGce7P/addK9+4Petto/EQfnUo8Twg
xFhm6EA1orA2hKuw43GbtlnAQWVgcTc4Lu3I2VcuXWVvWEtj3c4jlGYV/MtBr7SHKPWj4ZEvGZ7p
zkICzsor24/WRC/eBoh92A26uza2us4EMW+FDMtUB0/zrRl2xtjMD60t7QRoEcZ56GbRSnP1ml8Z
Ov0wNzGnvKXP9k/ZUBjczJ5oYYtJRa9I5Q+BPvXSQTGZDiHXxOO+87GHySt8qcD4Av+mph2upzfo
FiYfwaUKdjzACtzzDH4922rnGNyIgZc3ie2WHhO2dpkvQzOaOpxv8gNJcD2FremPoD0sfVFhSUQc
lMKM/l+9gPptotW2URo4Y2ug4l2dD5TkXxmLkCA9+JevOZwCxbkbzOss3Gvwq2Tnr6fT7qFeKDbm
GVPn/gKQJ7PbEGLqdyo8XYo4zaJqp4S2o76av4cwTEzUzzwOQqtRIBFALRydjlquM6htdDkfgcSG
9P6/qWpIWpveqXltOcT9up0d+jOA7JI7YaR87HcGMQ10m72srkDzRC5XezBMEzqMHE/thDz59s3p
bQFUiDH225RFLewxhW8lsr4Dj5dS4ywRtmeExNn1bCzCOBYT6BjAUeB2l2CRzM60b2duKDeMIg5z
fGLyIVjN4Obt457uumX/2RLTaoSJcRXU3VP3uerkGX6Og+uOvba1e2mLPswtg8NwDNUMSmM6hrV6
hyqUzVKZNhvOcU+0Dj4ehKtbSHCGALlh2LxNz27GPgXD4cOk65RiQAPUVjLcO1M3czFB0gClRsIM
iy30H5AYhDtnUC8idQzgALSA3NwaAxXAEByyFUPcDG19zZtaui8BPRXYbjbdiliqRFgi4jAw79Gq
1IQypRMQpCuYMiTsdaJ0EVoPF2aT4pOpAkQG108c9WuW/wPGVxx0b3Dd/r7D/49B+nPtKCvG54Jo
MjMiRecRF1jzmtjJbSlfiotOyioT65iSpxsQo25GDtPtctKd2geiPJcb8ymrJOms342K+9/Vjlib
nOzO3Aw+1FsLmUxN28WiDq3hFevUMBRvbCmryqGdYlwgvd74ijYb4aYIv3ofGHbOMPR91GKJqDxn
JwtfUBflzKGzNaP1h8Af7Kn6m+UinORCU36Nn6PMngOeawOSjkZHEaGa456bzqx5rfVnBKf2mHnE
kH5QcwpZdAnrlYcJDHXHZrfQWi5cKALaiym9Vvg5u/TTLSQk+aD8HESgQjkGBjS9ojjAekDLfXX6
WM7WDR+mCzDX3yVYITklHCdl0cpif3Gl0QoOp3U20ZvlmG5fvoPByRPoWSIsyVGHmz01izMsuy88
v9R5lQMrElNpXShVur8cj77hzL7oyNLq92BJFise0Xx61ZrhiIDf9quCuANHYWR4boIWGBKsULlT
DP+1atZP4FAItEDFuhP7YHn0CbUP1BUSfpuJEWULOzS5ck6Gui6wyQsQWudGGdENJHBxCrY8ji1G
ri39nzbgHRLmPhYqb7leUIDb9svDVMpk4qL/sLYiRYzC69QOUm8dXmucp+NQmWXXtN2Ulbk1kbYw
+/V5HAout938JjHWsWKFRz2dqvwDQuin0g5pX3Kuxd31KRWIQS0nw6DJNb/Wn2LELCjxxTtafE/c
aQ7xU4O6qNvcqa54XWquikARZU+wpGAp+bUEoGGo5sewuiFfj9Qq4ChL1XEoObjhRpHltMpJ9nnF
uqnmQNkjm9L8FGe3R/WjVFxp3fmBMHWGNlty6AoqoZjg+VjExBDPNQ5uCe4sKRKg8UCWPM9+VuHX
vRopNbdy1mRRrmWRPbhJZPPDu4tqf+vU2FJJctPWs0nhJym18SoBHFtIzynkgp86z8MXfnJZ4Iga
Mwc7hZ8WV3s4Kpbm4D41Xl7wHqqdH98qBprW3YU7HJYhdkg9WS6hcOAxQC4IJ52qYbAKa0rQ30IP
Rp5m5Sy6cnXmREX209b24B4aio/lPJNupoO8ImA9jC3R2NzwwKsdqHFxP/nD4X8iy4jeB/h9ILyM
PAEDWhEAHoONiOalItwmL8YjHLDUtjHb/Syi7/geKfBkE88/OufnnZuMhLYqIYSrXVmDKOByTsZr
R/1ugCZ6TkLuGnywh1snVHu4v0VbjOUIJUdDBApEfppfYRSkNWJ63VEM+FfV3BrBIP+Dm+5tn2Hg
DZv1EY3WqGPEttJOjxbK6905vX8vzDCtJAOu9Gfwu6ynTlqktaJSKRP+e9c/DPD8Il+R0DmdVkdw
xjyuAW7xuA2XTwDEwakBqFrfRFQG3EAlQe0JvxyuR5q2ggV/bYJoQo/LSt1wDgde7rWA9V50MiEn
7de9ZnNY3ONOIKZSaO5T9FgpldduMP/MuMwIC6G3XPaogdsuT3dsx7xHtDOKzhCtNE1H4yL6oIls
v76wE300hdKKj+MA03zXLFLChIYJWBYxNsh47Sx+SmUv9JG0RNpKK0lMAPK0Fq2XIQASIhM9ovQ+
58jHyJsInOWLMcBNwk2Jp/f1nvXu62gSQuB+ZPAOSmwOIjwU566jldU64aQBER1POsEm/2MOmM60
d1ZrmPNOj/jcSUCD9Bjgm7WsuiWSUd3bWJ3D1SHWhyibSVEN5UJPJRJ6R1W552n4sRwpqFrcbQJF
Uj81lVbv3YSbcYu5jLHSTcSPzKujC4AWeCv7wdYC79nAdU1ZIV2z8IpR5SLltOduN7lYGb8w5AOL
ZFrgi5QxSFOnaRBYmMe4gqw5HuYLbhhiXlTfMtt9hJEFUm6ukj8Fh+dY22GjtSn4ZlTx3nJeJvzI
I07o4fXTp5Zgpt8CW5pp+b6zn/NIDM4fFD+efVaDKmEpZb2lQPbSKKzeqXWaE+k/8Y+33zH8BziZ
IzqYHFjwiMP5RiQ6S60d2LGcJu7+Ok6/vX9wsfuy5f8DS4jS/EPj1GqNGJqpQMEcM/S7v1Q97lC3
kw/jxL6HTuM2gfoVJ1iZ8wJMTSapi3zQTNTvUnUKV+e5WvCuFcQO2K6gECpVIfl5CKqeK6Wnfh9W
AgRbOB5Kwl/xTaxf8YQ3S75OPG+Y5Qj9w1y+0/BCtWn9XdWgBVr2Ea1lsMa3RJCta8oXOafn2656
EWoSME1Nfwm2A6kR2foG93Krt9tyOZMAFTLf+6qcHIjSBRqGcsTAQorQmIh3WndiSlVMYSbpzWe5
Rrhw2jLGgYeDJXw9skHW0Uw7pxRYlToGoSE5aaAho4xvzZOlc6vLv/BlGic/BnQIVPvTWTuMNI9m
UZI9f7EnNXoJUvwqRwhWfeZdjDSOwLcbECby1aCe6jsJYJ+N+gfb1Vft5crZf0iP0y+tCRP4QfUt
ho/tLFOhAoNKyB1gvJjBfWoQ0LoePZtAt5NndgzmbDXXlEFlwXpyHIUass+IV7GXsInCoO5Vzy7H
XgPyOa2z8fO40nhQExfHjADY8OsvyVb+skYHAwRdKKa/M9jitrm+OtaR0JtiuWouGRvi/m55vWDH
xFLgo+Ex2eEy6/94u3J3P5lVgmifW6g6wRnpgfTSE/OgE8bPcS1Ltsm7MGTj0vVdTLnkhUZKppyJ
iFr1V/MKmqMAmaMqut/Oxx2FQVRgNgqmaXNW4P1yeK538UWpWa6hgNSBExr7+R2Hj7qGiujMb2Ak
o9y1YUbjbqmly5g7pY/RDRSYYgZtbn8veI0h80q012iObNepzvcmeV5KSk++/N4hjeTHxzvSyM2g
nhNQRyXuC6EZKslxnojMgTasfCbWglqNJlW+69oNQUbMnK1szA6nPj02EY+8j4FFJBSWeA4CzY81
c4FC8/DsiIogx7UPM7L8KgC/j2RRUVLo7rFlZm7X9LQF1x+BiV3L9u5axYjKpEh3KuUQm7l0Q43w
+OT6XGfnQ0afMJ8ufofw0uEo2idr4tWokeCcM4c7yL6qmv786cU5QCUvVXa1/qn2o9any+FoU4T+
lgS8P+ikYfgcTlMIdocwJhIJfRsd7B7+FwIfUZ/rVDOsrpL4AtlD5ZWOoTAVWJOjaAiNoy5YMc/Z
X35N8c8JPAHOBYMdGMnsyCtiDVUDD9C67unKXkEHMewQ053HO0UeFulVG+fSiqwxwZfAppJGvVQn
WSuirvN0Ytl/tD+RiQx2QFhTx5rGn1I1efrIKXOJvQhyislrq1CTEvzQqyxivJWTTb6jebPRCrlK
ivTQcLdVb2SgGoCJQdz0E2niS89eJ/Ne8GknUnlxT+6XDNfqKtt5y+b4Zg1EBg+sKpxTaPAWLx9+
jimDR6qJJ5ECqvQhuiHmGjE6eLXRr5zHT/ZNe61sXXeXjrtcNXYRnGhyxZVMDcGn8lgHCosO1eD6
UPxMgrpTXaivo/+WJYumXi7Gh1vNITT90nF4zQn/umwb5Nqhn6YXZY1pKSCjKlNjJoUMjNkKdtXx
4S+NDrqIViFHLhV8HXtZoTTm+Ui3yfyewEaTt2PVa3ggyHkxrO7loNVmcsg449gC1Rovi1MzDnWl
EOPsabqCyxZ+Ntk4/YRC8FkNZqOvF4oGTTfGp3rpPuYY8TLJnFqSW2ez/k7yBkRIMOZ/rjN0jZiE
qL1ZkG/2cnSr0HupC5MoM3gKRuMQKDC110AdA6CLrMpYXk4LvUm0MPGnubAr9MW6Hshv/gynx/mJ
ZusqTndEdIS5LcHSPpOf6dacDXFWEEJmk57cfmPRi3Lkn8Ql8An70HpWUr/vubxKwHDr7wWaOLhv
tdtuncVZJaelyW/HU8F39s8dJ2DtioVFTBp+spMb0nLU3Xy4XIhXUIcz1wxeT+dcICE1xCb18PiD
GSRT4gXrfnZPpEK5XZ4nLe4NV7IqQV3YRfT4pgRriRh24u4H5MxbJGy9hEEUVACBemZOo3rw6sl9
3kXJ0hhF6kBPsYIx21S4QSDMn3uav9e/YZEonOZ3zwwmoct2hf/WM1lgM2NWAdAWcqTpAspNTiTt
lSUsWEa2MB5Rb+D3C4wwbQXKM/REP+95Gi9QVfrUc+SswMuDUXhSmzDeWHT8QMuKgpkjkzqXG1ZX
7H/ncF/N3PhlzThbrPhbHhHRm0jrcP5iGrLzQUzW9/xEfhNDLnfd+2JW0LDjuyioSh3pVpY1fMAV
JdH+PtlwW1+CiQJ74k1SiIU9PmkON0QzYc9Jn4ugm15LHj5n+TUU1s/CSAJITjg7odWzbeIjWKep
lfk0uuFDfY3Zbsg89xXEkeqY9zku64WRw6QFrQG0EpOWqA9LGedWpsNw3VSbBZ+hWTZXP/pFrtzd
iaVTwBOGAff8UyU3HUG/8R4vWF1mXyHXXH7eAet9LpNCb4rnsA6UpEL8m0br3giO7s/MA32aYFrT
E/asWrOH1hVyvk1eEUgJTZJboZpRPBaogFICcWYjr5stNpdoJcQkZycbiiodEgdX+PvSu63l9qVL
6hxpI6KpaV9MR3ypebU0Ti4LF1kxwq3P2guXwBg6wC9163uSNrDSrr1NtpAqmAM4Fpvs3M7qVOkK
MhRwaCtvOdVDbXWqUJd3X9SuXuz6cIgOBJ3Ybi1JvOnOFcy1iYMUFcLNxG8NOQaWhVVhCgGHm9lv
2cJwShqXI3dNzo6sgWwuGuO1wUflLkNpxTrVHQLNbTH6gax4XrfVupXY4RGaVkjD6jtM7x8Cfdt+
BqeOvAmdpWDhTqz5qIMS90xno8zvpEDDi2r0ZEMo669hbcVfkmzpmvTTdzxShg1M4yPlf8HzK35a
jwc3ixZrt1paxehKB4EF+vK1LBF1PY217f8ABzwE0rYWfyurj4KBU2DCz20iWwXf5WVSGY5uj5hL
Ziia8fmAwElnSbgtFdsUaWMd97Ch0RMJ6Z5VEpYh3SNA5JYKqOpF8qjZ5Pjz/ubYhUcOtZnTEASF
MBMZIgFXIfEcAPlfo+sBOf9IQFO6Z+0C1P5k8o9jA9zG/Hg0Sn8sRaTUkgBPB7bfEIjn7SlCs7k+
5Vr22RcZEdRed6X+GCOrLOwkNbm4OKyhpRx104rebRXuz2ZjRFSL/yHQW+lu5j5fYdU9prj388jK
AMbUKS+LwgImxKkgTDb5rqMp7v5A0rFpo+vLZh+wvOKwb8WuGYRLpEjxGwU/fGsAH6sgB9LOcR3Y
zLmINErsz7HMK+otsnQEXqBZR0qvek9xB6kJLq3vy67r/srgGgqsMgU35u7NL0YPOUj7I7ot7Boz
fdmrAt10/jg4DW9j5n0dxQ/91Qfj83bFdiyv2BWH9UeCJyddEJly/JvlhvH+aBEk4ST+lSqIgueM
K6u93+i5YPA53G4iFwlu+kVES+hO+LYOBJgh6pyRE91Z2n4QKKm/O79jRY/V4hQ0hsgJA7aW8J1O
0WxXUH79bP1MNQZLM4uPqtwecKDPLpArf3NUrUMAUWStUYFNXmDP7R2Zconh+r6XDXzi3JhKfNKh
ucyZRVMi0frB0KFS3NW2kHdyG0e9iIREAP6V1yceLU/wRpRSHqbfraIrIjMzPH5dGFhtfXGtWRnb
XyeyP57E55u9XXk8Pc1Ne4QfyNJLcr0Q6X9KWEpGI+Rzx0oDVr8q0aB8YKUt1KLgx0M/oZu25wVk
pgZkOO1ZDt+q/GKaUlE5xW208n6bCr+G5nEASwZEhJYNjo20ip053po7A79m64v+KNmmbj9+p5dD
ylDiGgkasOjBBkEqQ2cB9yU/XPeHNROt844M+segFDsHWxi+qo2Ok0IBrYNH2TXWLGKHPft+WHBR
G0NJ+Xlpsw0ZZve75uoa5MVJGppFhITjmZ8FnqORVs5uPZaaoNJ25OLUJRBlVIYmNZiKrt1Qr9UX
Na3nTmSgB+Zi4ZXf8Y9wtTVIbfWD+1kW7JkKRjIbnlvC1TVu3119RZ6ZTiepIGMA4wzNRIJhwshg
UFj1DE0wAwHj2xoulxIUF5ag7fM7TPr1qUWQYmWoWuxV1PXzjSUoVP3mSg3JSOzD0ufWNa0LJXoA
FQrN770WiZxOUkb4bsnZQk12g7sRuRhMGjvRHXXq53vdt0hgRtct9I01IRlkuQEN+rvYdprFXiJq
7KaxZgTpX9ZQYo7L+ir8H47Tgx0DluF/PU8yBVgSrhdU9pLCGNWqWhJKYMGdWmFfxp3SP+fK7BDw
KiodW1bF9fm/em1d9OTqorKPixhzGWQgRTA6otCV6QEporzoy5Ve6LluRmjMO/3CfO2ougXdiNhD
a0zAyWyLpDIhaqDVxezeZXX62TZm7YbGRY5LR3S/5/mBIToj8st5CggtbnaO8QtP9i54BTSOZjWj
+Y3J9AY0DHD6B+q/sn8GviU7uoD/fd64VrwrV31HP72/OgOLb0xY07bJafQiY+kYDsrl5K9MQXjl
ta4pldZpC/xbIKWZpB3YhFjevpU+JmxKK4WUIYujRLqVS4buCL+CtDOckPHvpggjCPqidZXst+he
2WOMPMAqQ8/7eIlk2wnh4EOEkcJvDRGAR4V2jyTtCwLAQzYojfDNW6MNpSva37nMFhg8QangYH2N
9MW3Tx1YdWM+hehoVbEuO8Q6S9KomUV5s7NKsQT+lK4ZgsZRs7u1tN6mMprBwAx4BEZvCg5dM1Q9
+/nfEXchEXAiU63+wlYZlyq1PzaKMdKrU684ySm1X2k/MXHdDGLXpRbaXL33R8xF+lbt6I0MJ0fq
74+6bIe1t4UK+ORcgEgA+qQmGPf+K6kLgywYaObjce+l8ioMS9DhX2E23fX1XTuL0zMeVbdxo2+Q
nUNpaTZCPaVCGOOyGMZc32l+ZOQ63oxK9k7JMcaogsv5D0xyZ6hitnVlGm82CwDL6cp4OTFkQtF6
h2ZnuMZPKeUjXq2v5RZ47r2ZpIJhkSnf9Q4PcptsehGIPwYU8gpgFDUc0+M8/JVW7gvhcMIb6935
4KBlGZLEYcDC21mvpJeZfY01CWgiuvZtyrl+NcYt7bGWfgPd2b+frwVskvTG3mTEtT7GkOA45tU4
eQuO9G/b45RbfF77HBpyfN5UvAuPhr+yLzC3AzARRjUjG9mMQ7OY17LyMraaFCNwkD9ym0HXUguB
z+DdW4FmewOdLTqVZc7mbYcwxYoxBI+iQhG8vZHvrgNrn5TsTNbKSkgFwn7XjH5n/J/4WzR0PpPd
6/KL2JmHto1TF4E9We1GCu9PS/JT9pK/58dlBvyEOAUR0bMUaIR9sZ8hpq1muUPyIPs3X0seOM7s
u7mfhXbzBlWycDd+4xXeMjvHnwd05Rpnhc3Yz4haPuKkES7ydYo4cg8wO0LmcpuY86LLB76GdU/H
jkQz8j8h/KYUUj6kc0RyarbvudLGIxCb26Z0UhN/jZAwELsQUky0exaPNP/VYYX3ZVZOzjWFi1OT
oULt68OK7QxFhbL2vdnIJ8wMsh4jEqUBNNWfgAaYSORie8FD99hTyeUKKLoytTLsnTMpfMo+UXSD
xp/PVJrNP2C/q6yM/2H0Wd1ceEVD0OxnsrJ+2/mGdrhpCKHZrh1k2o/VF7u1ZOr20zUSzyE/52gL
2OvJJGtWBSIfT60sftrlHJBtkUDQiFb8X0Tyn1QpGJJtRXrHz/avEI6frTlkMwnDEJ+6mzFpK8lG
izkYT2BXgTXIIe2wpJkiTIDH+pRWPUeNq75POmnaSRwuX6yKqQGDSUFQg7sBIlr66Yual3lX5fQC
CsfXGdNhWNyFbV/qIK56OTtbFc8VZEaxBlvM4uVk8OQB1qyXU1X1fMNcn+tqFAAK24aUGpCLU75a
sYFW1g002399rzvoYVSucCnFnYodHT++Q3lY3BjFndPrfydjBuikAAwXpUOJAXXc+aT3DmhcTEEY
9sf817fKAa02dR6yT5eh/QRuu60Mdc8kqzr8gjjCZUPMhXgqRJEXTgx3pXl7sSWMqjeS+PKXOmEc
hwKD/3CKadPK2SzcIuN8hdO2jIRO69+ewIAMpEmyrZ5aIt3QGMXC3Dfvbo0lLndiQV0SsdHsNSJy
7w3cP4i0lGc4zEHF1UdY3vRw+8Y7PegJCaVlAlt3zYV5RtfkQ/pWLRBordm/9uPVIJVTT/9hiMVf
ydtXRtXW6iGcyYgks6q1rctlqo+O8dIdWpMDOKBcyVBAHTIMVP+Ivr21Y/ZQh4etJib8u1fXvyqi
kk4walZaa8FhEYAtN7WmDXsIcUEuGIu1TZRtTMOn1e5BTx+3u3lEsYocOYsz9RMt7rjU322tK7im
67P6YhEBq+meOVmwhSHzAvG72sAmtf+x8FgQtTJcpyp4C8kZ/v52mTrfedmq/KRU564CX63Hj4pg
eMarX4cC4iOqnbrp/A8iY2JEy2Kf14ChyX/mo7wCanqahiTBtSR/bG/B8DdmCIzbBK0JFrfHzhDN
7JKvP9CbHk/p9+YI1qFlW2jzD+hdFuM6HXsIi2GUppcnXpVP/DKkY2bynNsprGgmICXauWKVG1zn
h3ubeuSUZUzAuymhzjLN9VPSK+vMBZcWQVWsCSpwTwenC+zf/je8RLljZNsFPNTomyH98P1dZ+fC
yGN/ddGnhDAr2yArpR2/WhxZBSGCdjhhwztoRpbEHG1Y5rMV6EOxpk6X4t1yMoIW1tIzZZtOVsIc
LN2jRZuPlHZIktqMDzM6xEAueCtysAiNMisQo+FfPBxnX/OiBXBGOKGi7XAScyqGMkRAIoiPMIl6
QFU+m4fceZnIhMqm3gOUxhwO4Hvf/BuYrEqaC9btqRoC4GYQowG/1yiJu/0/6D6h7D7rigtVlrwL
DkHIpgLLHLY22sYsS9BLSVbtqbUfbzwmDKDUmNTfPthBXMlB13MJSHveUx/V5g/SDp3aqadyRQCR
g4W4hoN+QJSCdt4PAoqKpGc239f7Re9EZFM1E68ly+15EZfTkFY5YAZep5UIjvdvx4xZj0GONc0s
AKvmVL7oiS7Km7dKcwSOvygkmqGFsOOswOSkdjl+22dXTdsjIeOsaarTMacBXafvR8NXZhibRhyU
SJqe1Q1Uh1N2LFlrMl56GLnCg7E7pELxoeYyjJCFycQhja8QTtcqi8LMIT9qwbVM+FBn3Z1uVEW1
BfUtZUEICrHm3uzReg+hjdDSwATGHI4KnUjPfHkpiTOpj31j8ElMp2rKagfRC6JqDEOWHr7H13u2
WtmHpOkGm+Lkk2RlR9VXKFBBlR3m63Mjm3kJ1IzE2B0JKeHEECQgtFRgEqikflJAwDUUPRPKdk8X
FHyfwKwyG17hhldNR5+IRDsha8NqViVQ4hdjAdBv3xvagCInahuOqWgNu0JAK5Rsnn+snjlKVHdm
m1buRg+RMffLnIEPWzsM+d5soptZfOZVIuXrST95dP0JUpKn1mIKkIwh425j3w2JQWoZZUSEBX7I
IlaKeJMbiwe/dG/b3Rdf/eJbJVm3pHf/ZucidG628rkwEhykzewgKoyUvvkoq8Q+VIYIp2D6SmhF
kyYo8L5FSZwpFlQxPiTyo6CPeH/pCRdeIHBg7ue4v3PQsctUVFTq5MgIBxbNXOROiRDxaJtdgo6t
tcxNQgmUaavbG4FF8R8Q1DqTxBFaUW6lbQkz19TDm4z63uBvlWbmen5fYBpuDC6VIvC4b4KJdYmB
zFza4fMbg7LilHc50wGZTjmnExniEqDNs83JfIzmcSMhPGLNVJeFZWYwhJFqkZn1zKt+pN+jfcT8
p30Ao+Bw1EoknpuB8S38onOyI3nwULw+DT8xbnu68pt1ooDXb5W0yzbA+UhZd74NMlp2WtEzDbD2
9u+BX7Wlow3paIcSISURJajLvXImhED/LDTZgr36Q3cVJwptDVPb6fL61T0aOto5E8r31MDKp1zR
bHFuyLIxWptOqJvwJ8QDDLVKHHvUv9xrpfojgeFEXpjm4G9b1MvByguiTSJHeQ/ML89KciN4jVp7
uLtU3qnXkn125Z7IbUL+SCQyqHZ+YGZvIVIxYeFKkvY5Cyxi87Ph33JJV1rrw+7vXOOvQ0isikrV
vD4YLqmL7RnZ8mS7sQav1LyfwP9Q4fFTzgqajQUb714DncvABo5pGXf2v+NyqgGJOLhhmq3B1wGw
RjrGcAL4AWMfPFAEatIIRHvXimFuPhLgtANtgzX42DFHhXqOeMTD8/mhZizcOitMrieFkFmsNrOS
0G61nwbZginz5bWxYiXif0mFrfcGOzT0xX6Z2vdnfshcainPqPff89Zhg3j2NmcJzQlYjucDPUXu
16Qor/nitWCo9KxqT8IcAX+lZZ3JrzkC9RnrDoig7a2T5FgHJcd6GcunMHAuAjf3LJAMBgnL5Qlv
Aj6uAMafwzG94gPDk1UrD7Qa3ZsiD4GOoTJl5+XkZU2CtMbDzLRan7+g+Qp0QOwFa6Yxe2gZsgKf
Dn178ZNcEfUmfwLC+4k3oSbTA86ozHYM9kqwjd7XU2L/S063BtvNMuuU9vK1Ryk8qVQeClxMiVlz
iJKxOhgT4uMPvHkvRX2qkGeduiK7uyVu50ciPEq8ykZdwT44hOTl+ho2hUxcLpROpu37eU8R7qWp
YG495wmi0qQC4liw7VpaYnobocfbg66QYqKvKBDfnTYI4j4ZeUP2u8kpd9JVRlTdhCbg/5SgXDXq
HaMLRJ9Rn2VD53zXA8MfOT7VrC2WrIvkLTQkpyjasA27uiRDKn256PxKqeKTjmUn+zFPTXtGvO94
JLqhepX93drGEsqXrwKKia32nmjc1/LkTqjuaHaFR9vU8hXZ0xf81vRKXGVOu4gIu29MfwezfSMR
0wBrAIgtKQ/EUEj8eYwk83mJKTYQktp4K4wQzpfwrSCqrJubyyJnurEbueQ5nqn0a8G5WzQ2tTv1
LAqsOqpMtWIjxLqMneueKsO7I0Z+IwsBD7/sVOsnlBOMMPC4+kVn3KZI8D6Br8qNV/xrWhKRnvwh
onIAhHI408l7SgMcbHOqE/ogjqg0XY4eqft6xcnTd03uutJiUe9c89/z81inC3XbSFb0Ck+eUjJC
uFAb9Ft2Srj6hSAxyn9v6sOyhNaLFwtn8OqQLmHLDQe+NwM3YCEeAJwZpE5C0frwdxH+cbyb+jMR
MSZbSynDE1iY7VvluPoWVovPoTZqaDcX5K/rHJ5IsXX1AbRNKPzWNWl1wQ43otiU8bAQrMzX551o
XQnW7CVyVFKIkjhARiYny2qgQMk7S0CwUr7b27w0VxZ9toPGFBXbmssTZOlIuhC2luzkqvTMfWGR
bfPN66tjPKpMTRecCfQ+ZfKeZSgE0NQQn46xTcnlolOdatRsLItYVBChImMWWMwUpjkqw+4t9DpT
2ZdcBBYmGgZrTAD556G5yb8KhjAZXx97/wq3wI2suHESUoh24d/oo/g4hHBuBBmZcHjyBySg8DM3
sYVmc2VSIlCQw4OV9tdeV5oBhUDgYMtBDjRcE6H6SVCtg2fj7VGuqy9TRBY0q/u5EhpIeGjF7bqi
57IAqd1QwZsu0hJ03oD0KpCVt4ftOreaTRkA5SnyX0dkfNVEuB3EaQDFwTKCghLuLOFQUwIrETvb
loAIuyCLgtRbujM6fcEtpOGm0y89hKpVoGRpQH/MwM29xbHrLQx90MKMKpWuGfxueVQVhWPgJ3SO
Pn5ZGWpwcRvkrgW18k4MQxa11iRIoEZHao6HGi4j5oZD+0XbvxApYlCtfwhMB/c17iq0DFLoC6Wl
KyXZUZm8F0bkm/LHZpeHYkdjXxJSow0JBTuJvL1gDlV09BK+d3ciH9OZ9E7laRAheskuDOdQmozj
4FSvviyndJIQDiXnwwufN/Sci1p5/hKP/R0rM9Edd6brxhm2d65lj9FK7ddEtc92MzRRHDiFrnZp
e6gOT31QtC4x9cm95m5ilhQlVYKA0klkYEwAEZnrXfeXFUxWRknWQyPQyyMDA/grSdKnXD7/w6OD
5K+wW/xQjh/nRfqIbH3mQQionQKZBH0OEpg0cf7BQSUp+Ga2T3dldMhSB9+K8+dtrKGIu3eW8xCk
RzXaeUDnz/0LaKaYKzLRdzUMseJBOZqqvREofxl4wY4bw7lJ0+vw4ybqFfXJcOxkaouRCc6G7aho
mv0uab6DdRtAzoxsMbWragGQ5LKjCxWNG6qretV2R8D5WJMtclDRny2mXFVYDxKMItggcbQGibQl
dvZaFJj85IkYApqAKpxCzLpfBKEgKQgbOYHx9qOe09Hgv+RD88AuTumS3lod+a1Ah2JsnGJ/9Nj5
Qf+oGGeknSXzKEbprIxFiZmmqusanDgrmXxxICYMeuKmIE/IKYiR7Vntxz42KFttA/TM1quX0eGw
2m9WAUzin96nS9Jk9f8tr1Gsp0ms/TZWnHZXI9W1sZO5EWbRl43ijYM93MDTTQn5osjHADx6DUYT
KnuBMVckphcTMzuO2owgAF+2GlsLBQ4flyyYcWQSd+sq+NuFMvRP/mIy2Jgl4Sq0+z6oGlHgT3Lj
yNefpf/ue1G4i9dtjvM8tN8QDQbtlzHrudeS7EWvInWJVs7pGGNxM4IVZ2eJgoRvagEgHVq6+Hzg
Sz5g3MehV7wHCG2Lp6evvQcZmnBZfSDpBsmL7+oqV8IjFxvQ6weuSYvHvYDcwjdsid13zMIhI4pY
7wFFCWYXCZmJIPva4DTBH0AiR1N8ZChGg/PXmEBtZAIAO8KdozBYHWjibwZnWtqTNUAggj7NaUlf
JRDPzBIrVV47b+Zw+rJ6OrqMFupZVsedypQ0n4KYIVnkLrTH8KelZwrQVyHcexxu+Fcr8DDdoWo+
KW635Tl3+vv+C5GevgBctbKLUO9iBBzlKbvR6bwWAjnKGjZsCLRvwPb9LDrTjAgSY1IZ9wzoO6JW
g2uSU0Mo07SDvM4KFc0qmcLnwCy72mNNf8EHvZ+1MGqO3W1XBTiwA6RLIjJwnskjcxksvPv4EOmM
uPLuSedFUtknn8Vs0/CP7evzzbv4lDJ0E2+Cy9P2NC3N1O84n/O8yNhaq49QC3iAVxeBmSEOHb/M
hJ7AmA5dzhN+lRAcJsutra67YYoRKxFlv4riobWdClGWPyohEmstCtYOK4p9YeUUNsyCp7xpAWN+
2ro1xiUE/XODqVnxT15rM7g5A7BMT/ItqJ30X++1DvriM7Jg4nKhv0AsmKzgyaYXTvOAItuo42B7
j6OJt11nhO5rkPe0wlVaj7eireTBU1Hg5Ux0KqLRG30hNuuD8kO/rsSI5mPI/fR8ZZ9JgcdgzYRe
0cQ5YZn2G/+x7G/EzbU1Ax1ZBTS5byXCjIr5NxoIrqMA8xBgX3HRNl8ejuv+fEPLvOhxtnkdvw9Q
t6zUHULTcNrcT4c6TP05DQ210bJ+GtqETHZcRUhRGGeKxKT4tjBvx0hrjcNXynL9LpZYWlFZFP4N
lyjkh5rgiOKZYXC0E4obTMuNJF3oHSr3tbMFW5md/v6eA/KZ0oFkQ+mEVn5DsGhbzoR5X5k+njE3
ochjdwY9PbMyDMLjFYMClQfaSS3CJcAZIx1u+VLgZlcDZHsQ7cwnmB2fyuSgSYyTrRIaIvVP9SQ5
KlkGvmNYMO2+i98FuHJgR03QElwll8wFsGPRt971OuJ9B3vszU5HPPhWiChLx76ZxpbwNvlAgOLt
jBBgWZr4t1+aGQyyjdnpjCRs9V9NCUA3ve1/SPce6jhHCpEL9HvQCGsmAfiYstksQFjWUP5tkt/B
w0MulWzLL9nomlMpluNjAelDcUM8TEu47/uK7DdSJvy16FxgekNFG311FYsP3HR/WbHNqpKNy8AY
rLdjHVVfQYtls7CmFzm9zqvjx3vbFSVuNe6NEBkYD5IE60eP0AV1QrO2hg/YJEMMT1ipV9h70pFS
ohZqaGtRHqVtaz8LUi1ulhdP1aV58TY/Dcl1SGvcMnXdYAahpDxp1uuAehrrYdwb33XVgW/nrb/q
MfV2J9YVmrlaWL5YCEpe90UJ5Q6HtCe+WapJD16b89w1FqxT8IlsYuYGTiWlXIL4YaoUSkJvrXV1
8nMds9l/2pAYtqTZMbztb8bV+soKpyHaE7A/OQFc8lR993AruE4qmDTJQqf6Bv7jLKHPRnq/XyCj
yW6sxNTq/FZHdGHXBhd3siyi6iAipSNIU0Bkxi8/5ZjaninreZI1EM0a9zXO1Ksc+YL/n89hf46O
ENUeAwcb36kYn+TsDhTG2ma7sL67zJGpt1o+2aHh8aUg14hSR0oeXXuosqftxU6tPB7qxHESV8hI
TRjayi+r41wDOfdnPMtuZdy39r2yft7odzjQCSAmxTIGA4M5UtgMJqe+HRI2hRaCExb3jO9HcCFe
HdoQKQGrIo6dbe/t3I8BzlyaJbf40wvL/vxg6qVL3mQK3PFpXcim+cn02DuWQPBIyyX5NjXj6paU
T7UfolGlGLMnhz+vIfBHUmhsXb1BGPeZMAjdGlS5jXwyPB8KS6fFhkCCP+Pq+M1P7h/zufVBtGo9
KXpl10e6J8IAHi9DMD9uMuyL7i16cs+dewfTlEiNxOPrtjVWCIC+upkn6bA6uoLo+rrviaEeq/rT
A4nyqfggvJnAzFusD8+Gjw44wayuQ8wHYKS59z8Ve2FbOWOdUdPqx50I9oJeRqRVbKkEk50NlgC2
LK6Jgx3udALtr9rzxTTZUhmDybwJORUnC2QGxUxOmmjFpdVQ5/uNcud+DdhPTBelc7NJUjL0ElL6
IVgGpopCkzBp4NMxYivcL2ZxtKpC4BaLt6sjjBHl5Yog226vNsmytpYafHg8BTzsJ8e/ve4pvZHa
K6yADbOQiJI/2e0l++pkH8su7OA6WGOTgUjXJfTrESefi8XlGAaIlnWyz9UMcwyuviJS5vEKgPsj
kxb+x4RPCC4JLyNJNz6EvyA7Pk6mcPaqClLlLYN4gDAymkn8VVFW7JpSKPIVklNYENKUu83C9tuZ
qyriXXPjNijrxJrhiokIkoX/SkDViWG8H3to2j9SRUHwrURX/DZ/AcVdJcM5oXKkQUP/kes25dFv
RTSMBsu/V2MEZEEFodhBYAvELdfeXim3ABCUN34Y+l4llqIPLYZmchbNvakSlvJmZL/snmltvw7S
As87TfsD4DaujjAnCwoQeELxe/kg3IzBE/SELHhq5Y3vxb3NEENAr0yU6FXUkIHQdsNQcFWUMENO
ORQzxnEZp7AR3Xe6qUWnf0bKT54HyCDIe/PgmDwCC7A+2gdOsGN5KEqEWhFf1er40q8kB+9Q8nn9
Y8eDsp6MqqPFoq/TJuRFsnTFyBT9oTC/SOrQNuhGvbTU7/ba4ugQ/mQP3u42pD5euKy0wXV7CdDp
+LVO43/ecchegOcjJyj61SLRTpEFUr0gKzrLZLoHeeqeaLXbh7fthk/6wC/cTBtOpNybyySPkRas
hFvBvbJyRws00V/oxAvYKmuEDFR0X/efd4ByB/CXSiPY696qC5YYZqdf7qmVyAniZJkxgyhaBgkh
0USV/UuPn2B9sSYevAExFb7G2ixUIQFHDJhyqPWuXZrUktI2YIp41hxSM6+dP563swpgnRUmBlYY
mcKYA45PxC4cNBQu1QWNxxPt7Yn/lqxWemgpz663fnFPmsFUznE0aTBofs8BxGzVr0Bqsaugz/d5
T2rqMcTsEmakhRpy4qG8Ovjphxt7HCBt2Z/TDDPWCusXAab0NYL1RPnyjj+1bmbIoXCY5+RfkAqK
P652rhhTc6iK7eRBTV8o8d5YepNhaKZCX7PGDJeYi/DFcJa+QQa5lzM40Io9JFco7GiVhinWGECp
TVF2Hoe3tb0QtkbwGDQqWnt9rUeraKeArqtTcqJnRNUeHtvpo/3vEDY56qew2V6wP9wiwcf0bkf1
HSAV17pDHpA4c5LMtgBH12k9eY5hUpfFRJjC0F2AuTG15bs1wj6vfPnnHG1sjMsopX/PIMO/zd+o
EzvO/vSB72sdxRmkbqtkpf9Ea3MGdMLG3VXWU+7QzgTHoK0pQ9mo2HbepwOb+61uQAmQoM2JbRp1
2/UxKSId//MSaQA0azg8YMGdUrVxjj6jXHk4dddv+OWtoK/FIX3OOHYnb7OnmpeV7nzdAv7JnMvv
zl+IhyA7qkhX5Yu8Ta2sY8JpHPmm8eLcjhHJHal7gi5HL8A/db4k701JAR3YgHLhOVgVKm7E7VJq
z8Wk2joRePmobEclwvJ90uTvKjqrBMRQOPWZHkP9wiOzsYvJul+hcZkHeX+0tbNZMukeqn9/uYZs
Ou5/R4zPZzFGSYkG6WVhf1saAMD6bKhs3zdXSkORZq7sXXW5jLEDj9HD2Mv46zT+urqMCx4DcCIx
bYr9EvjZci+QxCQJti1lgh25iOs8KLgk60WAWprRUK/CRCqWqFUyLbwe3YZyIrNXtnb7GdvRt5Wd
GUTVhM0pFdlwC17JWvlx4fNBwUINXJU9OQ1z2w53DWRRr0mZTwooR30LqwXM7awvRO7vVSHLfYbl
Xn6q9wndPbIdRG2LR3xdUcvJKSokl6ex5rJfasCGt6SD9BkrDRPg7KAGeHSDMjl6i7kxm0ZxunlA
odPDkZDpJmaBliZsAN4ehlh/PIVEd+ufre/037Y38jLGfzl+fyfjQHojOVpVR38kd0x6nfawZr/x
M0Q5fsebEmntr966jIdg3YvOQlzSvRFUA32ISGY/kmMVSRcb1phGe59Vb0gspBtgEakdGJg5d+Nz
kJMFfckspPRIHwwyymKdb0CD5cKKe5e/OB2F3rGANhTSPODqfR3u26jsyNS+SXkVsDdaS8N1tgkE
P2qIYweHouQzaowrqHQoix7V/JHHb3ZXGonoz3mDOQXeIfpIkznT5jg61nZSXhLgsmA1eWOHlD/f
cmnumdzRISWTG3TAO46e8K8cIAO8ZQKFuDlHvft2JaXFe6+3GA0dWdW5kVGKkwxoJ+BFatwpTEzp
J+twL+M4E+mEEgH9Ia+HDufWxDWnCKi9xz/boGaU5peJgCCoFFv12+2caAgWPFID49ytDoosalh0
nDFiKMx2BgjVMILIeJPpiU0swBWyBXlU8qGqoaoxC1fT4yLZqjpr7c3aJzn7RsMOQXlQHGoiuaRz
GhnIXLvZpq4YZgb5vuXQYCryKViDLoimv8mf7O+6kVkaWFZEzIJ+s4nnHtftHqbvRYdxr03RjQAg
IRPdzjSgNnjm+nh1SxC6OWUXjvOPUSOvHCxtq/gOysX4OEVxryT+D7PqqGzdkl1x8BAT0J2732In
0Vzm5qn+qlzPIVi/PJ8n3HIu9iwsCSCcNgTQE9aVWmPbSlPlu6SJEuNDFV4VsQ1kB+lQhhVIh4S3
ZXELSfAhhF0uhBxVUJKtO+ogUPC0XUGIejCq6MnGVtZ+nG4epqMovz9EimZbc6CTuEyl9DMX3c1Q
ynBWiXnbgU2i83iLDYfo/dJVTSHPchQ5v/1v9dUg8MSdqWdQRjzn0qVIDnF8186sd3VgR9Nr2GzB
6RszSLesYu0L13rgr/bZHd+V2MqGCaEY7DDbziRVVKLiki+EfmsUiN2/E82vOnBHIEvZGCr104kb
di4ZfMo9fuKMw8ZXUxmPgzRkNE8qwandr0OwsAkYKAU1gNBYApcu5m1JIbwlf/vW1Aih/M+mJko0
V0UzsCtmeXCV7pqyPBuAosN/CcA2LJWDC84LCyVNND02ffBMfdiMzsBo795+WK1gHWM1IMKFv9NG
rNVkN6DVx8/U6KsBj7lamNQHo4YXe/ab3Hi21ot6Wmg3DEnCEGM062J6V4m7p7p8umSIyEdl01d3
ryED9GNrbla+4byxbq/btZ+FeA8wF2d5iR+VReiMhKOujgQwubNsoRkaEUNXxEsRreoW6oDXm5ea
JWav+gSY4eOIUe1rgieALTX8p+SXG3G63t4+8xGwWUFje1VNscU4OgvZLriY9eIMq5P46WQRmg/8
CWl5l1qFQ5h1Qr8dEfDXJd4YRg2p2/HHbTzeovgi8FcbNZYW/qOieYW8IzRAhD+iFDwlXI5iukhd
/5BzHBcjQUGuZZsxwchOvadxIDBYlmwM9hNLwEN6sJaH7FwyCQWPagKIGWBN7s85FiUfRp8t/Uop
t/sxDmGZFErAGB8N3v1hns61v32WTBrbaKn5SAGCKjgOeV5+Kw6I3MV2uMRiOdWH8fHKV6vqhfOG
Spb8QAAkYh0mJ9xCpZ37leB5PJFhbkVNijeEeN8sIZrsT0ab5LNFiwifjI8Q1BpoLw8o+I8Jh3ww
j1muqotJwHfosmN2JsgGMrFhKBG4A6U71GbeEud3ACOrohGP2KdscKeu9/A9WuPmpvBeq5bTy82i
MZm6QbzIKZyZdKxWK+Jbp2jEkyZW+1s62lv6/Zs+W2Q4gVkLDT5oVleLALqvcYwQm/olyMXBKBXb
iU5V7HM1Z0TV1DUYgRTzB6FC6MQlIg7VrrBf6mS0VUPWSg8H0FqiIRHjWDkWsiA11mYuwvgMrLDS
YSagM/PKSbB6JQ70JGMgUZXAWu+4cpGYZs9Fo6LyeVEKw1F/d6AcT/5Uz0M36TsBQvvB3V5kL6W5
qbC1Kab+AsfIjQxsXZFuYcfac5lN+K1P2mdiXSLuapRwiMlNCukA6cvFTYK1CEiIn+yLkCuiMWbZ
Yc5I+mOrpn9UyoxOyqXP9Utsu+TPKM9u/Jw+5vK/HuA80lOg87tupBRmNZ68Odu1fY1X0kCBigaT
f1ZBVwznmadJk2Abp7XbAxN9SwbcDXL33Iyv0EBGXjOyaazbKAm6tI0/fipnW9676jWYBHpuhpWo
Rgl+I0+fIwi2cnt6GlqWB9onjq+vvpPptxqX1SkmR1+bH/uWTm1O4NuDycjlI4zsV2svSMakW1Ec
sS6mIAzomFtbILvrgvrJJX4BEiWnOmgzfSDD5BlLBoaOtzAlK+NUi3T1Iqb2WFbFmqipBbT6EgVF
MiY+yNIJYYKong6AUv8bnATa1hjyGg96zDOjfLig+xct125U+tucynOycpo0F3uZ5zk9Tr7WXQI7
cM6fTU1wuSOSM4FFir+HNbrWf7NBCv6GN+Qb6D9uYT1rlwAMqlhaiXVaGhlkpdJBumdm4M9qJF8W
oxkO6bWuaaj4rYeNhuIGBmBbEeTf5UW0vLWbRsKG/xhbDH+T3MgWvgtMSTMrY7/L/2bHdeTK3Zuz
peopgSioyT76uGVPyclGO3/GNLaJ9G94YVYONw3oou1q2DGT3O9kBh4T5/35hMt4CTggfNTIZHXK
h5OInMMcroe/RgmBHwt/WUp6ywOZWUa0gMU2/9fEdSk3dme1xMZSehEtw5MnZHfoJEuI74S58rI4
vddMAC4fN6KXJpwpnWQM7t+XQiYfQqiltt+mZK0HieckmWQeB0klm2usJW9Ll6eguBgbSMiqQqbs
GoUYABbeaATKQ9OSglQRUqHk6Km6N1TUPySNsR0+9+0aIUslyaaQkA486AJMksokIRJ5GZPUulwc
htJ1i001dQyGPLzRK+nbcLDw+5xygzNWjKKQHS3XeG1C7ZoANbPWA9NrvSwV0jyL7dUkXyexg28k
lhDBRpwVxqoSaG5sulFjHYLarMmJ/eI865Py3k0ios1UF1KLxtd9wuQiAQ11aePunYOp0LsRJAMN
kVKMJysk5dVrZQgrhisgGzPqLLPdNxnySyZyL99XJpfRQrbmP6xIlvAjA4DSns/m6WhZML8nZDsR
eSSxlC8cYAfhOWYCmN373MRrG8MoyTrC754d+fDXD3IjVFVpeyYol3lyj7TREjTm8oKLewm5NEpM
6Rhy+OfQRb6qRTtDBT22xx2APfYglNWaDgEUHQxNhowsd24UAvhZvDySss1rPG0F1EeT4k5tLgpW
Z1GiVi1f0f0V99htnZ8sjPaJO53CkVeKJA9Xvd+5/r+XY+W4B80a1+fOgo3Wp9SarLeahVLzAZS3
8WbN+ttnp1nDPVaLpFcCVpSrwVqNC+EiMb32dQspiZa3j65/++rRntxyiMdPdcWE48ZewaUOrted
iDPm13peUbhTzM/itzNALovPe5oABk1yUr7/A5OK0WUpkQkXCWFemB9LdRz8NdJbtHP2/5BHqsZ5
0opyq7eHqVtU6Nl9MQpnwXe8ooNi8Jak0i+n8Kl90hQXZWuEOxPripVTXdZnO0+c2c+/FRWTnmSa
3pjgP/t77w5zzV5DnUOpLp0tpwOYkaYVeK3TC6+8P51YFg84//PfyJnZvUxJfgJlm9BK43UrkAFY
p+lHUe3IPhi3Ihxf8iEyAHjWQ1WPdYRGIaqpRfxKzmypoFCk59am441qxLvDNfkzb2bvI81oH+5/
zUww8Mb2N6aBGB8XNN4H/j1Y6Dq9YbF60w3MQ23SqL3+/uZKF+oDDB2EGJq+DXHRGhRFOJP3qzcy
pIi6466+hLgxBWvsM0FlhDeTgkZamTacx2a43JnrqjmW4YJppf/iDeFpgi6iD9hSfasqRnIl6s63
dDN1eNBpCKkTZNLg4e7n3hK1Yce7PLUxVcypng0NK1ZUVXcTXYPqQWjKJcCEPuZd4eu3wyRJ0aYs
ZayVQw377M0hgyuRp0nw4lVXCXuLi6qvmKktSHEXgklhcT/rOXQQrCSczyULPN39FNtckYTnqfux
OqWF14RBUX8GlWEizsA4fW2Ywu81MQCcWUbDjMv3cFGH1x9GRNvMvxS2P2T2lhcyn2s6qAMF/TzO
ZdjDI48N146IOWkNjerMvfsX9akdW4+MWnU5tLN4UFX+prREuv5lENxKFnYzxHTsyRODWSI8xGYL
3XD2EFZAo9CqOYNb54LdrRgJ/QNAYGjOCoI8C9Ik/SMH/aXvEmQawUJpshsmk67F46QcOr1m+LRv
F0RUG2VUps+XwrjwwU+WiBJfx0ya7/hypgSTUoLnD5jpKO1FLDT0j7UQIBuJHVCqIFvk9OzbXNT3
ruUjyh3HnMIY6ZjaUdiTpUtf1/iXaZzkmo38+mWTcqa6yoLjN3sA/IsOgMWFdOF+bqeK3zgcNdcv
DiKs+rHaVC6PkZm/hA0LaWzcY7DJVwwsFN/7UZaj32Nx42nNOy7LSJTykIwd8JBbkSS+seV8/PDP
CjSNEKjksAj/oyiYPWf7Ut3cf0ZInldjbfYHkdihfSPIh7dddDRGF1TtVdcgvCGJDzMx0xbwgowA
ClnwbDK+OXzl72E5QKH3e+1QcmJPt8nspW+xsmOPlohQM79wp+LL1YJSsnMTA/BhuSeejmj0lvt3
LfFzHQYnjekEkG1nLx6maOj7PNPAcorMG2VSdD+dEyI5lI4uFyqlZymZjQjUGHwVu477UHEpui0D
GCMSnFju6TcbZaQk8vh3/ulwlZl/nEBGd4HnEy6BHoB8W9U0o+OBviLZ7d2UPHJJNJOHqxk75RHx
F0Dly3/EkGs0ip+9o0MY4Xw8gD4dexmoQMoj0BFMq5AfL471g/5rKaeTvQh7oL8emA5mJMyUrnHs
oDXQFy8G2qoMupjjF6rsrZ4ycbWbymxvu61WXjPjrnpyEO5DrajbbF2u81qkpTxWYZmOZHJefPqf
lN6RPaSXhp0TY2ySMUYPAoqi93CeuNd9msQGK2axqty1xFApmlowfrigmTfZJYuz/bNKBx9oxA7F
mRr5Hc81G0aC5pwv3/pZjxcN4czgZU63ShnmnSh0M37O9HusaaaJBwSOwGAav1qGEuAhzIaXHM8c
e8dmqU/P7biaThKmS6W14gUeZhNS3cy9SU3AXsXCca5pTdhEFs23NyhrpAuLLVLko8RyHhaejq2T
3u/zYVeLX9iXjjQGIFUP+Xq/8AX/4DiE20rw+ofFdMOfnZWXnjUwiXMb3HzHCl0PU0FpKiSmNMgo
RsX2l0mdXKdnr0xxMLuPzgz4tSC+2+T1PRf6p1Z1GeEq0bCNB1Oc+lKe0ZPFvcF0uK09m0AkXWKM
1A0fpOqkA/aRYk8qBdL33I+nBt9lZb2ZwCGQZKKNpS+8kLs1N3OZ+WDobca5LFTiTShUPy7jw/z+
u0BeeBdDYwyO9xX54U40+NM4wii11g8ZteTBcXlHUtgGX/T6mQSfKLlFpjY5oTeogp5H9eCLjwr7
nBJLEoa5XEn03ImbBmR+Va7xqGrm0OTX2nte6g/E0pon+WMSPX6ep3sgECSZ4L1qo4zIp2W1LGiC
8YXJBydE6Ol1Auu7UXcun6DGHCDMQbBeT+Jso9JyF5t09GAQv1nngo6bEg5s8hEaaNT7c4I0cxI1
Qi/kpEUn3oVFoTN3jNP7iEmWgfNxV+r36KJKwZvZPnr5dIy3+zIrul1ZPRVNQzNDYj24vOiHGFVr
K9kXAVR4scFXiJsSzI2mTdui9l2PjJj/fl0KBzrE1RAdHMPPjwHOcxhQgZJr0fy+DAbQxN10NgMI
jRw4pMWVz7pItcsfF5fKzjuqTPBA0Ko3RepECFJNVCJO5nD4TI0T9xgmto8U424CiYrqIiNQJccY
5+9x8TQd6jS5WL344kdmoJhYUamZSF6QLvioMYjRyxgB+KPmTMEGWXueAUrjrmqupVmGkiRTCXQb
8ujnxqgSaTFCQJUg2hc0fJ1AU9gtXsS/XoOjNKgCwCnFkq2d0MIGDupal4kxMLtmwB/Dj3CosZK+
aBVu6URTpZ3q6ewHC91mE8OJX5O5wHw+cIoJoa4ji+J94OnKf1I54VyMHqfeJPBWtul4kJKzX8mY
cJYprurW8l50dhwPBSERbxHAc5c5oMY0xnI4tWsB1ixAqT6jcgQgJmdTQxy0UguC27PyQq9zhPY5
NCJwYZCurQPcsEAjKlxTJUDXUwvt2o1Lhy+Qyp+4iGfSUap9enIgMlVJ59uj69PO2BfS1yfvKTUH
FTdxvT4XxIfHth++KS3+ROEffo59SwGsb/T6GOLrwHxeEy4J+aOkoOwh42Hk6QBPsBRFpSwGgF1X
Ra2VaFfnb4HaV3Ov/78d3qfbfAjuCk45IirAHyKwnsY7A3qPo2UnsXz9USJAykp3rnY17AVJQIUc
2FcHgOrfuMes3ku1NFmIoa+2+EAxJG4K8LpWzvtemI5MXKV/Eb33Dduv0Gc5wtonz5yF6kRqyRLW
iN0WghRkUG7K/3RSwqAmbOpwpJEdzhbgvY55V5zy7b4t1DLrng2U1ti3lKFbbCDa+O0g8ijbJi6i
At21THRj2kH/VITYaf2KdWa4s/mGnslLOkyEpAgMDDjQTvL3CitiYCw2kQgVtAr0CcbqHOirIgW6
FuFeeGDdMB4kR8q31Fuse2doyUchl2Nk8zId/KVV3OAGqyLB2zdZP4NFNBhxpHK+CzrmkoFepYRL
/OKx0c8TbTigLfG8I3PGragTvizuUraLZVoexwAS6y0oF94sulYVGyfumoR44brgrpPdBEnkEbhp
NVXj+0x4fx66v9L6FwDBZb/Jf4LA00cA9QDB3VyNV5Zc5qo+EWZojucOjf0+DEHVNmp5j3gwtI1v
hTo1U9Pb6B0BEbrJYpa0XPobb1Yw5MyqpyThX1VBXMleNKXxPUJTX52XqQ4TnNtW/0QL8uqryAPR
yUenbO/qnaHW8vEMTRRwiDol4hVq8eEG4sLujZD14d239yLvX0VeiiUHPw48l/tykwgUt++luaVt
mcCj6up4RcZkH2r2MGMM+AZ+CbxuYX9WRaLrwtf7YNiwiicEVZKdYMVHrJHu4S/P+vyldX+jYkBi
k8RdZnYvWaUdZOKPRQtzoSOXdvHlZGv+4pmgfjTXouztrnig7XBiwPB0jtncQvCUqpI9lEMJAnr1
PAuzzyaAY/G5fBjzi+S714VEX4Tp/ppHmIEuHbbVv+pNQkR6eEEoVxigIlJvrRgh3BjHM8J+iASE
R++qzqhql8cR1pnTjpuHND37B6Xm98PsooDB27XMfq9k2DkD5DzibrNIfaKFEo7L7xzIuyqH/oE8
Z2/9pWsPIv/AdmEu+E1Rr9ZAU0jZS0SIkkrwAwpk8fQC9y2WK5sNeRdK/vNYfBHCcdOKNlTsvb5G
aRQDRi6gyUGo9YKJ5xBabr2dF6uYfVQPDXQCSgFxNUquuNDktU3qDdoTdKtouk0YgnULGDglQyLN
50BpPjDrdJ14IoM7RzXkdNiuC0TGoEo2pMFJxLEsDLUIRhY27gnnPsNiRmFWycyZGQsI1bLgIDQV
3UOF02Sq46PHYhgGDZlgMutG51uOFCswOHZvOP/yd9UQY+Ot84Bcq29hXtBXMoMkUIpTEsMdAXPn
ROmACzvAbBVKP6FRF8Be/YwU51T3reXOF0SCtXVgbIYPyUkxEd7NcAXKO5UGdxhL1hz1ilOCdFGz
fEzAh0scmvxQMRaR8Y8cZEZ2peLjrZ3GC3nCY5Y1DomXSnGpIKCSvsYIIYupxb8WxKkVEjV7876k
XQK9oLKw2aVSevOUkQ/cRrsulKX15WCUvyOEo1Un8uqnMkeaoS37mIuRCSFyJql/vCN22dbdloLy
Q2MCUb9CNzfToxWUD8U2+funH64fx0apCvrVUnAlAOzg53WY4uUqnRL/BfAMjW9iODa24Irxssfk
mA4Oy6W2qibWPC5RpRoUuWD6DLwSWHgNOFcU5lpVnrTNmsO4Z8AtU77tgV3pQslEICIc1KQ+OYFJ
WDj1peRMjNFNpNIbby5HaWtv2kg/WklhDpStXADtFf41FDyGLKe2OWKImhJhM86s8Kju5SXAFRIZ
c74ZWdapSxrOlKoO8HY6DgW28vmtdsHYyHS4+c5/Q0G9Kbi5IJVgQzouXwLlC/LFJTC3LaTt0EvR
wygUqf+esM7EqRVenQ2jGdpkJshifPGXvljSRzM2F4jvDvOk+ChSecQvDbsxm31CoqwHTFjZ+uKm
8NbIv3kG6oKaR/prEk48oUmhXxt12NFwQ/a8glLT0aEdzFIeZhvXiUAqwYoKD2NqByAd6nphJlA9
fQ+A3VkWWu69fnDRNGuZS+bVQ+TXjvtNVAzTpdVvvd9CXzu4rgSBWiUVkiXkKBC/AAjfYi1fH++V
lvolIRR879JB/w8mq38WAe7ORHGWXTU4lRpaEQ9QHyKhHmQA2JelFny9/RuRmMd7uaQ+/gBSK7ft
ei70JCbOM+kpLl3QDe3zSb7qgq0MLy3Fx4vUQF6bAMtD1+93sgZZhXYWBxmB28GcqvlJZ3N437rV
PML+CjXixUxKFwZ/3dtUqDKa1MCOzCIPvpubSjrUSebv2m60dugouIGQmrTLTkANo11LC/VMXnE3
bFiMk4odw3F3f1Mnj7XHKbgjfd4qdPXBXZwW+bZRblum2TfsZMeTDsq0gTzHStL45OltnZxDqjmp
KpHygdLmtOc56Qh8MOEJW6wpN2NPw7z2NuGRPrJrE7SGk6QHfA1IXKnKQ0iNAlqM2AZk1b9oFBxk
HofgTqNWcCRDej5A4WcmEB4bcA7j0LB/oJoG2kIqQxmfJNDurV+ZI8o1csm4AeWxcougqYKrO+Nw
pWitjSaToVfoTtWjzrMiR+ZiFpNoBp9zce6bW73j/PyEJ0JhnczSTbb4E5IDi7fHVTDBx7/H+Cg5
KN55dpAGdVUpHSJzo2CS3O+dBLYd6oOGu3/UIx1EzZ7Ftga44iClfSgHv0rOc0S6eKVj7YYFxbW2
HqCysEb4rvex9/0NwMB64m10MIcTx3Ot/R/7IniYmCnMX2fCZk4KODXPcrESxFWQeotgAGIWmmCl
L+pHODmAISnRevix5XUfxQl1aqWTkjV/1JmSWKC2WIm+h+3NBfc/a9UHNK03GbxfZiCGtizcLfl4
JB+EPHmviBm85UILw/CfJ+nuYexPnrlJAe9e40tzqNw4z8pQIRxjEnBXNP6qSGhy6ajtFdXkql3i
8+Ywd3+Rnw5QrvwqcjjOC4WjHa3ybELz2T2VE0AeuXgDzGo8NmpyePct0hOaa1TzG8UE0ESzti5l
tR3vFwaBDAE0EqAguzqHWY7MG6gJMqUzcL4Ww7mUXsp/g+4zIZpRDLUatow/YGacMI+NBvsUEEI3
TwMH77oJQNBc4oZXhXgtYZhaokS+Fp5PR1jeEp1ofi5F1PwPQZTDhrkhXRGgO6cwbu8/0gM1+vIq
YixTgl3+9ZRc/3sssNAOTLzUZ63JkFQVQkQR1z+JW7o+QBZq3O6efZqsT6keT1nu/oGxtq8sBwOo
LRUUaKx5K28+eTt5Ikv0UrIcRUwOQWozE98UGsh1fIFQZ9vye8T+F0MdUX5H6wRGdkp3blymMrZf
5snqix9rLf5rRJsxujWz/ggg9ax/Zm+aptJMEg2svC9pj2HJszifE4XaxAhHrBGQth+cF+opi3AO
YwokgW1BXY4DgOE1kTqG0K337DwktKzOleEDddNnC0oGPrT3cp0+aXWTuXMG5exvRAJ152PUtkXj
mbnWgyRAvceDCY7f15udRv317302LXzdmlo0vJjaUc0nstXDPk6AWGJQOyY1uD9fOSfbS3eOh5UY
TKA2uc6W1SH/z38uPXqO5OcIvwxFmOt0W9xTmmmraWgh5F1NFN1eeQoCKiUtCFIYImvCxSqCsdTh
kZC3bozliikiHN8F/FTQ41TYm7lu0xc1nc+CIKYtsIhMSnYidYGbK0uIo8jzGBLdiwU2zoacXYf9
PscPW0WupxtK3C2qIECMWAIm1Oh3SuWyBjPkP8f8ZM1PslIzdEgmRG3bMIfRK9kzw3OWb+pwHqCr
WLOFiYh8SHx5njC8jvDa0vYtAWm7o9kbFPuMw9D5uF+xwAWmk4DKKO8hhrSnlVfDUfSHo3NB02oy
6KGaZ+gUmFyK2ZrEOopvXaSwgyuXtH6XFHUDeDnPhCars16Aj71TdVWbtJBdRr9yVebXqepxfHk9
Sv+9EFyDbSATv4Y41hmqZXiVnZRQ7F+5LCaqMHigpeNQSbxfMl+ihRWc16WzRVlGVPneqKPDqWkT
dCR37Hej/S2dRFsX7YlQ7Kqr4wG4OxirVXJdc4cFH/KtSesdw++YnEcpy8FspIDQDXO3a1Oxu3m7
158GZFC4O4ECZOIPT7EDZpHhWlBs0CXG7QrRgXZCONYXFv/oj1HUlljw/GkPntIsJZVv51yq7VjQ
R7Siql+MIICPeGkUfQrseKpSxRCp5lIAzroyYSqAsfmIBVK9tJmWgt5WFOk6jcsVQAxhD8EK5PDn
r/zPf+CndlJQs+V5KOL/jfCsGfnrtsGLhSjEzBvCwUCv0FoZdMW/5w7Ix3MMm81L7lDTswEmAgjC
2X60U0q0klVjHC+7wNg8WH2nC5NKzRxJ0M516T6HhkBqEI7maOiTsoIo1d5HEFQVae3WHwdCOYGY
698rpojn8pTYvNm8hDw1lE1nRTK4RV119gjE70fcypUAY44mBhIpY1dmZ164KGCt9ytsehBtZAhW
bPilBEVvC8nGEJeqDuzrh/ULcPHrPLMgbegUiW8YHOY9Tz//SGeMl1AFX56wsoZ8o+CGVyTYihTz
1/2GbIfNkz/F1cY/7o45zN3sW6KVC0daZ/S24X/EcfwsJeXVmY8kyMIxM/oLN+8HlqdtADu/ydXV
dsxNHT7dq6inkG+VBPI3hKYunapCDWmpb7iem/utf/UwDpUXFYXUkBAvXeFHP7SMLGjZp9SWajZ0
XFNgPU0bLJ40zFOsDnavQZlZrVVN1NiX6jjrno0EkrN02CTfp2MbuoB4eQ/YJp5NZuJ/+YgXvOTe
mJr+ooTNb9uV17OSlKVzVT54ncHOBEsMJluFeOBLemBzyV09JD7RCENx9cuc719tkEgRSZUEYRlw
OuXDZQPnSB4nGGlsWLQE21Dt3G5RmCBSHDfuLzTvI3TBI7p7Ymt0ISyw4BX4UhiJ8EvUktOIw013
MmJGIYC4Ng5Ls3wiqvu/b7yNC/tEQK+Xg6PjBjvp7aNhb2y8qhHquCbouYeqSnAqHQiij9Nrn1kV
jyKJdjKvpc8eT36h3lVkVnpv/aEPH/ZD5ALYlHHgq7RIlZh75FVe/6Sz2DSf8s7mwsjqtfMW8rXy
Zb/ULk6jcB/6qw1tjnU3onHGoZvyECrMsopZ8e8Trq+awhTlZFAl0Ukn47cTR4/XOHwLnpVrVirt
Odk554kVIEhAKrpV+u9+gZSG6GhhepQtnyTc6dfhadbpbUePPzauAZc2Oyoik8Uk9P1idV/c6ZKm
deJouwpRFg6j7lt40PCGhTf6rdA6zpJl/PxY9GnsJOUyb+eQnBw1OQameTOd5GURkyOuehGNDwNE
lbkrSA3usL/VKZ79T9T2Rm7YhKi9l8fEovVscw/RrTM9M44IC5RjeIpWITLeg/dWbPKcij+/ntIW
8EhuLiRh0RFwqyKdfNfnzyQ8yvB89vUW2ByunTa3qMjXr8A9+xBNzwonXdqri/ozvDqR7ik985zT
wAu9GSc4VCd1phrRIuiwBzvAxQHisFYA6F11JUIkY+I6HhYlonlEfVUqmRqxVHEAdaiuSA3z7crW
iBiIFJWQ5/cdaZRRosWcD70H81YryS/gznX3WBeWBvtGFh9b83RyxyNKaqsRNcKVXbSeAGfZjFJg
nXM0oJSX/SKL3c73+cy1T+cJn1hiOwLUHDYV3I+3AChnOQIskfJLLmqsJ0ADuSTpVO3egvrgyO7J
06lLHQ/JRdrQhsuAVqy6QeBgYlzTsP8s9PGWbM90eTcbRoYCIWvD5CS/nHfav7cxnykDMXXGhPeZ
mMEIqFUFqWiJV9TkA+8+qUZlTfQm2vad4o3qNXQSjoCCmgBb2X45UoKDvXRgeO/x8nOz7gQ9Hme/
pPRha+7WgSEzOtu3WJcafGlet8ZWVtNcl0NdWEcDO7u4f7ajzs2vN6z7Virf7VgqWI84mQgCFfAn
n4Vuu2hRj2WK7NFLhrmp6mu1Xm5o+fh2SMFiyKFe+RQLeAbcHpx0P0Yda5xX++QEhlo8mNMZFTdp
BeAPPrAr2JsIEaI5X9smPQzka5KMI7zIER7Z1bV1tFu2B4ag/NgxdhZXFqzl7liYAHw591lUuv7/
Ln8nze6zbCfDXf46Ra51WJAEfghaguVtCRQLUZcyp/n0YhW7vyZFlBw7byNnbDANrwl1x4cyxc0o
LA8yNTb/VJbEos0VDTOToNh1/iWl0+Yywx+btkSg3cwoh7D6K9BZRtTwYabRHK6KyKHUTpERAYGV
Zk7d7DQ2FrhT1LVX2Gb6Efy1jq8336wNeNwTA7/nyOVsa6ps0PvE+aILjoGXxIjfORHKSO9ZAMID
avJziX0WrYf7BkHxlaCcVK3PUVVvQugykgIyW6iWumZkLl4o8k7tz/BslmbU5CjMAR9NNTMw2C7R
3g/v6+fKX8JuCdoY1/yP1upKTvBZgmJx3WwK7/4AFqloXnWXC2ELcainzSRHZ0JqFf7xfpzQ7DbS
h6Kz40ottmiCgG+CFTLUZX95QB8a4jegcxm11RzSMBsNfRUohOyck1g4uT+O5vxyvdUyKU8OAc0O
Z239r7Qt9lyCXmkObCw7Aj/hwar+hSC5izzHa1vFiiuiVH8xEjlCqgBx1Lic7JUh86Nrg5dHKkY+
Wyhx8a5uEFUh45VDSNQOXknhOr6q7XX+p3tFM7UAQWIiJBlFYr/ypyea5SvBGnxW6ULtKn9aTHtZ
W4rQYvNmYPLgiSnRdMgKrBjefzvumpL8BxwZ+dSepC3eKxUr0kRebvivRJW8cReYLE+bhg+U2c7d
lHevLnOcEp9NVQUXi7M5zmpgHFAU+5u9N5lNmfVtz6u91vFeKRTbhl5aj7h4nIs3SnDdv1Xszzxp
V4BeqjHRkqW20jTe+CZUg4phibh1Bjmw7r7ciq+ZZfwsrOV7kwHhnx0K5/avYL5mYdnXneK3oWyn
OIU6zSEdq29vJG7RoMcH3sQ4KgBi74cNoJQE7e8QO9Ndl/mM8YpmXVDIs8qw/1JCunxoEYtZqEpY
Qr37tlyGrpao/SVvjzP+0R/dR9VrgarJh0dXb7eK2eLa3e735t3vFzvLMprDmjpgIqigkqYoPgSR
DWiTNu5XeEqNLU+8Grd3/khD1DYDSmaHcVaPWhKC4u0QsaSkHY5M9m1l6XzSSqAZtOP6Fe5qPiPD
aUAATnEepz8/DH5CCyA5KRXNiwsKDU6/mt1+Jy231cIaYv/SlNuY+hoJbiY4+iaFVH8gkbfOiQZp
ItBBbJanfuC/1/er3MpFCfPA57KmBCCyWzyxSxKP/vY3QuO6WqlqkwkLqCma+esK1jZmHVt8Et4x
n9tCs58lmwmeCVLZ8cGSihgIuN6zmlgjorOLQdULlp+4c8L0E6AZocFRDjbedTmT0kAkhCevPE14
dU3JmZUKymG5Swqzyvy+zoQOz9qcjzdWTQ7GWtpzocV+H0q5H7P++4QqJeohdzoTTF1ZOGbHcpzn
la7mSLlz2mcgewxFv/LAkaRbb2JyehykceEmLLdB87TlmWBc6vmRZ6K/Pv8TAR3N8UWKdFWMGjig
AnwBVDEPk+uBOdKuXaAX73+zkaQ7n3ELXMLlsvla5cremPKYFHjks/UYepz4mX7Hs41Z5clEx7eX
Ai/ilx2HgZGUCP7vkKSqoRdnP+TLOKWw1GruT3/TuVcaqKcVyQtrYu5IA0NVJx9fYXbIEjs2BCu8
GC075E5Iuk5rNxK+g518FFnF2zn+RyKh5eBeKHXXJwJfyk+KzQ9Orx7NPFd0+NB33BQrsFtImCAa
K9Jxfy4BDZZtAxj5VXIT4GCbgSvwwcey1IAM1kHsaxvFfkGYN1xhB25d7gr/H+pNFpc5UqaSnong
3st5+323LouncE5HGFdFNL9isBM3c/9cfgX27GDtu8dkm25Bt6y5XLEHQcbVTNa+DMWWmUXyEvZK
+cu9lQh9QL+21dIl+yiRSRv0Af9a3fOq8fpXCFI4+Op8nSXe047Zby0vmkglFFByHBBrI3z+kHcd
g3jBGrkE7LbtyxYPe8m7GVdxjlMxv7X34BJqg9AMa5yMFfqbByC/jYaG3DjhikwZJYD7UnUIkTx/
SJQS8oo4Kxusx35dKeYDP7WxNv0/m8mGKiV/Z4wgnU2U9GR0knMygW32yi3vm1Zl4sJqyAoPxAyM
tphXjLAwzexY8NG5ltey/oy90yuvWnHz3Lrbj8JB4I1+MtHDtPFJd+NzeipKRnPUG5LMTwic9A7s
zSSxFsHw1HUAg9x2v6pG2jN4aNDKU8V8uo8CYaQRvS//CI+AVnFYHNDX4RsP2f0E2/keyF7x98WM
EuFE8G2XOpFDMwt/TBZAtc4700QvWIaCrk5HnB7ht8AzOyGkjdmqfClwAAWpxya6oruuvElAxXHl
4zPYhH2TxsX6875dEt5r4MMoYLd7/wuGq2wzyz/Y6BbLSYnLHKe4uVqcvJjq5F/9USwQ6I/uJFfG
yeGFPZFWUu6xz9RVVqMLORpMCn0Bo2e+6z0yt5D/oPGF6RQogIiyzubD2BEMSop9yHZf9/4Zj/vF
ORpN8gl3O10H46bqiLrxmNkmJUHT07ASieMJPl/qz+sCHtyxLpanXmc4uDo0dPhegMafCaorkhDC
Od25kz11fqwkShVENmLpEMzhFqrE13vnFqdgaMYvI3leOee705Olq5z2C2gZOEhvhqXXo3j/DMLC
iCuqrHy8D+LGaoo7Y0Qn0bTj16DziNW2j+wuP0Z9clqE2WaD/5X6U7Bd4Ibje4yrl9J7M1vSnJqz
LE8RxIO2LRrF/fdh5ft8WU6OK7lnOHUCU593pdJM50o3RVVa4ylU6oYTG376PCDlUshwT2lPNOWx
NdLecwsUZ+vD0mRdNZRJAAi3Y2AOdb5glqm59gi0olCgoBqpjbtEDBVSrhr1OWbdFex+8bW3EjDr
aNWIAtEO6ZMkURAGmcUxk40xuTDS/GG30Sfwv25TRrefBikRSmJth7uBDLl9wktXYEHDng8lMtsZ
BO0gTqs5Yaw8L8edSgwZ/UxsZ2912xu2mOaIe4dv0/fQowxRX/+0mWL/3kYi/Zn0zikQr8lLQcJd
cT2+0JRITTpET+OYrE3nqOv78yvYB1r0KBEzBU8RoJOCTU1BMmUC+a6mI9bTGQIxmeSCeAKKTlO/
xY6n8y/IX2Wb0mV51BuFYXZ+w8wfR/rVajvvNcFehZNT6n1MzFIN4PlX3v6ItzRvIhNlqxy7vzpe
6YSbeGONrOSSjoFQVTP2mmuweZq/OTNr+kHQZHwCj8dDuTssc+xTzl0UXxdHij5YaCNeDwpj7q4v
yJ7LrDj9Jvz0CmQIjnWUFibUT8XuvhBuz6nWZM061Pu4u1jUA+XikeQjujG3QLWF4HpJnpeboe3s
2pWB/KSt8UxxIiwp+yEMT6TmBGuH6dt7gNRYvg7Fci7b4HOaxxMjmm0JBmrndAjuD+FBX3YdO5/W
STODS9hfIO2cisWQCav9FAWrusAvwJMwtK+nqWHox9vEM8Cy+TB9cOjbaM7rwiFMkbI7DSMy9aPF
uwUCq6hbehAfRdnWeAIFRZlSbaZhIo0ybNBPI3pjcFr434f0EKpfIeh5ng3WL53/xRc2DP3/Zv0W
mtcGC048+TG21eJdarAgDaZKc3/AJQk6rCI7eZubdIXDYZLTOggjI4sx9N0lyK52tIusRCMO4x1W
AbvWdAMWKEz1AskIsDp+ANM7q+webHGHZtmVMZnOCSzN76Fl+YQC8YH846uykM65FvJnBbN0DsNf
DcC5oZ+AQYKSaWgvkFlCJoY2Bu7mSxlaIAVDEBUyE0NAEDMFaYEGVrLLFgJGw8CQmMxjjIvNlZyR
IaZ7u1b+FWomVD6RKsgGlFh6c4cWX5c1QVnVkpxHN6/T4VnECiiEUAQl/+Wz8C2BsS25ie9eHbGq
ofKcGYziuPOwb9n/giHHvR/9ItEUZ3BzyjdyhlFl7x4nK+n3DhWKvKYTgDdAt70bMOuuGxCoiSQd
9QoyIZ2b28dGDL9qqfBfmXUi9yTY+9jOJa9PkWYcpsMvgz5U+OqxdU8pAZjDL3sqV2GO8NYTwrmg
fJUiTTTJozBRnwQSqL1VOaOfPeq74s5pJDC8Wlw8ubTf2geSdnjrdkcDy0+ccBCykE41sdKUkyqk
aMLCo3SPYqjWpoSRYKBiLZzMx8ypwJSBxw8bR7wC9YXkRQqqDoNUmMtJGtd4px5TtdXMn8nNuAxO
hDUw9jF9croTVBL+yMLRwP9LzonNHRQs+rsECP+rdFRvyYp4NOguMJ7djLmpUOrpW7dIULpbSg0q
yR7Dhdftn7L0G/EsDiEfSL4AwRsmubBV4F6S/FukOOnwdaKLAcAnLA0c9nIuhWN1q8KtgIIgdmBg
/SDTH6PBaI6isjSkKaFmwxWvXgdYdrUdSpTWMTv15ier2XhyzhdB2C2Ir2SmBBKGmmcQwg8jRO9P
0wKya3fTnceapk6HbeI8j6DPeKdUrnEQ4XhX108WtDkJuEglNZah4jy9e/34N5FxedlDN5iMWtRf
xZQRliw8Eo/9yA6jB3omwhbWjwfQ+rNOvbiuNoyT4KMghIBcOrZxV05K3u77hXRoDS8p51OiHalB
FZ5q3jTMrp9esQFd5XHKwvamXbLXABfJrNA9vkOOOMEUDRb+ASyMw4ZS/2U5o92UAnyQxTajbuV3
TOkmd4GdWwk9Vt65qF4IrydWN+pCWaczDmECm+2olaz1DfcGOeEfOUxnLjUfsMkuDuuLnohEyMZu
x5ZSAlYkWX5RYFaIJryUZ9Mv3aLtmkj1SbVEwxGGxeZFQO0B9HGG41gi23hYZ+kgKm50vg6h9Gva
he0YElgkqSqov6s0VkwbJgdBdQbLct+EPdeOXnTRZxQfc65vjs3qIu2a11mx1x3XTwfrKvgsaNRl
b+jKGzKdN73bUZvL/uF72ESR1LIZDYL1DiKJaocMyW9e8MRYSMoAPJ8NnsN0UolLFFdzJZdKfgOv
DL1LdZzMF7NX3yW5VzrX9c0sH0uCLjiYeGj0DxTwOed6dKPTtQtrnZrXbLJRDyG6NN/Arw7ELE44
Qwzm0Zfu0b89Y7q2nGgQQIF1uefT1w1W6qbOdDKVZ69Km3GZpPCEfucJ+X7aXrJgExX7paq5ItAt
GYyQFIozhsscewoIfspc2wXvJn0JJqC3rVghbFetKjVfWlyyTGJf/f9mfrLpHBgHenWqN+xdVJdG
2cN/0htXFRyXwB3jMDwKDA9B7sM0GMzCm33DqXF9hDmw3Gmj+o0n6XHQbFdguahuNQ8ixo/C6HBi
uTp/e2UGR5sf17teW/Nu/fg73p9NGUfzaM0koJTvDa2mSfbFQCIZULFyH5x6WM11KVbOsFrhChk8
TQCpHKITSk4ZiBZCRDmzTTollmOsqeHo2tSkES+SW8Kq0mGFzHsrkny9gafUhV2D2Gyv5b8/5Hn2
rOSkr7kKjwnCQlXVVP7q2hmG4xlyLfsFdAYb9z4ZfXNBijfi/qjb5lQUXcMCOf8zb5Eob38fi+bg
N7DrTOT3kgVHn4fRhmtwW5nJrZFWRQttjSbVGIo0spCuPjmyKoQIy2aboQGziXny6crcrNINz4Kk
kfTxKytmlRrSf+JMWu1z8+o6vMJE0ZWjOSr+XZMDqCqQtzdp3JjSFz2bsctUXpTv6QJMACt02WPo
wxgWPWF72/PfCtp1KvEcvd5rlHurSF3aW1M21JRcUuFWI3CZslynFVOJJDnhZomWYxIfqUJjkbT1
BnkBe4c0AeJD0g54T+gFDgWwbua5q9kyUfHI2j9FrMxSAZayyh9mmlEcfbloYWuCkUIGlQ+di3lx
qUw+FHmkww5jsY6t9oUQVEDwLK09C4fIwL+K0wUljIho02c1CMfIU+aMZ1u6KEinTt4vN8lNhCT2
yFT9jytvjiRX/larPkzA30IjNIg8HF2VmiDO9xSq7thBNr6ItgOhaTosApONwO6bH95wrdeHRjPE
sZqd+kMTGjmeMC5SXoJwlRxtBapLhJ3uIQbCmZkJlOrn0Ii97jH/ILG8oj6lmgUm4WLPm44GBfBs
78Mx/hSG2P7r2dxtGosalH21Z+pyfci0XR02bjPLH++YCjgqDAfTJHqJabzJ1qDJOFdWHWYIzel6
2uOoHDckWGXWhrlysuhszuAePOc6ljuLlQ8WDVhaqFHrRO25903AjS/1RBS+1XEhuVmGOpSMtr8Y
uy0bwOmGaL6uWvNpjq7YKBu7796JmR/F5ZMiSXGwdY1upiPXKPpDV1UawWzaiHzgw1FINi3Iql0w
YDh3n0VDqknYeDtna5rntzi9J4S7Cz2sFEoQGXzrpXeVdEL75KXymJrjd4C7MWwMS7nD+nGstyGa
U5+tMfcz6tKmwXHgWcdn+xRQERTvrOiS1uWaW6w8Gm7U4axw7LQ5RwAps03jvfO/qRxWZL2oTUgh
oUZiOVAZKecp0CyxAR1doGIHm69vYktSk2W9Hq8TLaBc7974U2nFwIloyqkBTXHEyG1y/GIj8I21
9hjuaVABhntR3ilBte+Lo1XGal6uhrRwUzGrTHJ7UJS8s8m/c8NIbOEqXsBWz8ybkl2yyjavPzWI
dyDmGZmWU+kslMbVUJ5QILLxe0I+VRduVhyCC5a01p3C7r9hqc+nK433PP7uRdwpdZ5m1UfiqNaP
ifLhBqjvTv2qb5DU6N9aFuZWGnYhyEODZtd357Cv39Hqp0KuQ0TtC3dy8Dnn9J6f5mlNSL3S4hxu
KR2vhVv7mPXGE4u2oZG5AfJjuxkr7HwvyaFVrM02rnxZhX9Ek2fyCecn+8TMorsqhsnb5Rl+H6W4
f4KiRFv12dgguTLFgZL//8ioCTFrZj6dZuPfVoP8XdNFCeSkv70mOkmmgn+tbNo7vGovroifkXdL
JB1uhYcgLa+F1Z9hSPOUnwT38L8PKCuKBqkFKv+3cO+smbFtnfuo9ds5brRv/mzkuDvKyt9dqvlU
p8/m3rcliKZ0dw4gONBypMo8VSGbbzx6uArFG1ARskb59YEjfdXsyT6q/En5FrWOdJQOalS/hmbD
W4UvmtQHEfXXIvUU3iFZhTHJu88wtf79Mm3OC6UqcslJQEOXvTaKV1EzwTtNlcjYzcH6zXybgnyq
MuUJZ15N+8yjnkIlpNAzqxcL9Kk+Cgy56Q2juKCPqVqC7/nhf9ziLzY9yvtDnNocKD5kzO5Js8wy
QFdKbd/u/Ap5VNPXURNMU6dA+5dE0IJ5p54ccOz+JLPGefoiEdkZFR4S3FdRNJtMXu9p+1Zrf8rV
pApZCX0IL1PQqLWbHfhUXq6itRZO/n48i5eedZC9G5xUDqM14RurVFCotlBzn3utJwqP+9QyMjYq
SkXUttxW1xgkna5cnoqCdreK2Tqwjxja/NDCexAICeccMiYEw2UJe8RE2FSY7QSuiqWKNv3qIA/w
HrwGCyxE3RZz2dVJpu85gXOUg2v4Gax9f0qobJONMJE8i/pVBBSivoQjYbRW6/frF27Q6+ftjX5f
ivkd4113MTyDHXzzlhYL0uovwZXvYpQwnB7XL/aQIOv09ovQIQ1ltLmeVsTeybBm/YG/Xs7Fg00f
wyLqJcid810D1dD8Zrr1QAWQq5coO2GXkq+RfGf78UOf4ZohYMfbtGhOAtogbw7c0Td7XoCTFXFC
1SGjQL/VSqjrKuETTtMbQTbAR8kyWZOAqno0ZeIIoZJ0YcMexUdZRjh+ITw3C+nrY/89tul8oshR
4l3obe+oW9sK/t5a2GzmPbblFRICYBcd4yJqAgr88134qOPRvUGMBzy9SjfjmgCpp0tK6CLlFfkk
Crdd9u9y+kCme7iACMUaAF0NwYUH1cSgtmkguH+Lh3z3zjrzgsffuFtaAHc0xE2wpD5O7nMQ8DQL
jU0WV9N/NAUNqSMnndhoZEXWkmmq8CXM/wnC76FUHKO3GUXe1ZG13GzxUx0jiHko64jh36TQcOSe
8hm48Sw6S++JlvtgEBD9vuMoAfG4N06mjdEqyBRbuN+MGquQW60fcbMdHRr3wewa8lgMtUZ15DJ1
PWSf0ZnWkADaXHa2O1GN+3ai39KUYPkz40xT6HCI8iOOcETx+InFSDoyu2lcThZvM3+V4iPhRuOe
LodGfCb+LAsNMcFc16aAdTe3478RayZ5DjQgBoJDY6xc2Q3kmzzJVwn2U89Mlo4v20TgFzdzjjco
gEbBYlx0Qyr9nblLH+LGR6Asqc+87waMmqi/dzYnHPsEL3DD31BEbX4Stl6UxleT6MeUQk88RNRV
eoPa3vc3LC8M/plHuoAzfRoyiSlJ7nM4DM4rbTezNJRqyYwg+ZCmdmD2BAjnt5/V7XoxIWiKXEIq
khwnPxq2ZQ3a9M3SUwFUxi6hGdl+TLHXv2mlwf7vKuj30XABqKApffZ/5mpRF76uJaDavBumeonw
xf66REgXa6dhujRg34pItlucb8idjQF2ZzZerzwJwE9A//4Grcvhz8TnbCS1KM2diOBbfONjtqMB
yff0TrMJP4ET+qsVJuUdAxe21+H2dZb/qtITXjEiSsSsQPBZNIz8y5VZa7Z+SsEH+vK3SNE8peJ2
9misKIZm4JGDhz9+rn/NuLdaFgY2Y9MyQvHRR4meFPmGOTlwlfgsCg3tJOfZaGcS9m01LZ11WtS4
0HFdpboHdqy30g7IwAYFL5x2OfCOVqCJanxoAHctxSZSWRRHdT1S/ax/gegSRAeZ+sWmQm5sM7y/
1Vk3fPkXwcH5RquwAEn/Zg8N+ZHnDGfo63ToEAbnSS3DZg0V0/siOlz9K5pGOtItFTxn1pi5LHFL
ez2O8bH6lxmT0RhBoORwhvdnmpVq+VNatnZIvvtXROGb/Iv+ZsN228bwRvNJCSeAc9ILTGbJxhc/
Kn0rysHn0LWtN/m8RN90oQhLejaUJvIZwSAAKLe5DILe+trpgm/sQxYjbKa90qYdOn4G98nX72iH
tr1rvQQ+cLwsFyldMwQKhoB0dKYBqp69VPY2ii+tYgu4okFNuN7E/JLoEtZ6SE9qhlopnEj92hmN
TEVxxAYvWMYYb4lt6UilCQCJq9CJwn973eaC2QvqR4ahVOjUD5GJE5Q3XnNLqKIF+rUHTcaa/c/0
SGiIWng5tSM8MvI8IVj6/o/tYDUKJFqtpCchzKOqCah8jy8hs4GrQsbbk8hGt/S0EMaUtWJYjBRB
aUXL23JbtZZfSWl9Z/+jKrz+XqLJTZTGh3osvnt+d5VDEFpvFMHIYRYm73Smw27nZX/pQjqqQIcI
9bUZ7DDIg2QxppVtOKA2faEYrMR3+SwCfEyLdNyg6ohypOtFjlXs7DZ9YrwDobK9fVbpubzyu61r
nnPC+XUqjA+aE9D0h3KzhSTKOjORv++K0DR5ULYqsx89Sqk+ZfPEUIXV1AkTOaQozk9bnsn6hOqw
JdzECMpeLqKlZ0rHg1JhNU0DcYi9FC2PlhLGxkk0V3SuYelsR/5teu2//UFJAigrjlN4hCD1SLRP
EdK7sI6IG/vyTNLqAUSV6L8o9e46aHnwYCHua3dEujUTTp0dPeN2sAwFEo/71h1RGunMut34wE3y
9glnuuKpI0S4HrUpIqFB0vywJFKsCpgbHdzTTVFzA0vWQX7LsADX4C5wIGUDC4uESz6jBKXrbMoD
SCgAs9wN7BHi+W2Q3rv8mRD9XoY0daSKctEEWDNFMxn6c38s+jyYJissq22oOLJx0svER9T0xsLA
sQf7BJzRS2Jb58cZ4qt3rETfnRusDK5Ifty/8phsKdIbgqZprWh6woYtSGM2sAn4Y3OCpCUpIuHY
0u/GkLh8vEEABsBV2Ajac2YFJS61VuW92RNSF0oQnkCg9FQISDk40IAaK2xMXy5SwNb94FBvVDMp
ey8ELyMiyjNizIbjI1c3dhofs8vUmZZOi7EQDVJd3yIS/7ECaJwAc596d/LHlE72UKA/FwL8Mp4b
9dCzGjbivWhLMh/MZWh/UrtZ3kAna23xn0BzymcrjxHx9xAYyXA9CNEf+FSqzJndQbCogMozpQqF
xkiCRUAShY+ytE3ak9G+lxDeICZueiaardc2vyvU6lwi4dRZC21ko0JM1P2LnouWg+fxM8hT1k66
09TlC0kUWyTQm7Lp6cwS/Q2qKF1ps9ySzVQ/F9G0OopanbmFdtRMqbc0Lqsp53nFK+z3s8RyOCfY
ncd3vpiAkF0iDyRuzLfmLEw6FPURbDLUJgKnyhiPXY099ujxdcmKnBqcpcgQaAsd5hEepx8rtCt4
qBkdKHtqIDfyTRkuac3e+KkODSpgCHHrGVa0P/NhQ7ZTTaxgpz6/MVIUTkzye9TrtoU7/7p0PCOo
p4+/uoPJMHlFO9thzkbxoP4LQJBg05Ya/l8jqwtRVfDLVPj5mpZ6kLRqbJFtdTk9PTx6E7s1gFg2
ZKSaUXlY+8ZYtpzzWjZNaGozY9jBMN4M64WjdiYWfVArBPjDoVcPgBonE3s3RiUpERjkaqbzji+P
8m18zMA6o89tmrVQbYb9LZHQdAIXZ54KLuMG3PJ+wUlnquDx38yytJtxmxPfCiEMNz1uANU8Hmth
P7S50k80DNDY230JlXeCkiPhsOWvA59EopuGn+81zRugT5OwuCCd6xxRgJtoeZwAIIUeguMnBrCi
loMXLPwDFlyAVYtQsFASOPdYCs0us9gg7bW3vYVmGq0QA1WMkMGTglVQk8HQoGc81B89oKA0DNXH
PdLM32Op+uzv5PmcvUiM++4D5tWkgMqtNcRZ8YbzQ6a23b60G2ZCrckwJcYTyAcU/KXNAHFF7Cj0
kIYU6KHY93xc+PZzR/xxdzZQlLwru4NWLemuYSyxSUT7lV2y8lx7BGID8lN4FMWB1dIRY4tImxKq
0oBNKOTcyXOYE0778dvx21qpV5lLrKMX9sC1XbQxl12lLL+oO7yZ8lg2JAuWlNzMHvCsvBTK6hnF
A2qFkuQfV390MP/7yyKF10ruZz+Z2uNaXzOgGQgXgDzzlbSknUAKVOMZ22zh5tUZX+Y4sk7Nm5gr
l3daddMJ5IreR7j/v/s6S5dw+kTJW/qamY+/fEg9BgcK34LspXYpNz1AYjLfe/5MaAlM7bUCYkC1
amk8SZ1XI4dKpKVpayDhcGGbpzhlkAUOUASha38lTjEySVeZPlpcHy+nXrPs30AaldaUL/I7S49X
YE8T4sUq+YychaZc1eymuU2YAInWCt28nQGb5YCRdHlxwInJLUaalmXUWjJrc9QdgLDYTummwV+G
kksUX6NqgfMMpPsHmEl3N+bJw7sPa2VNS0NBHEBhiQEtuVBUK+mXkyGIZGd15eUjNci+J3u45lpZ
Kw8yzLKBuDl/mRUuHKqoq6g3uvA/Zyucx7R8laSC+I/BeNNeNPX2Z2uuNXFb8ZXmPq6U+/xF3MhW
Y1sPjVrKAHWwSsTGZ+LO5ofAzOXVp2CL8uZutJN07509hY0Bw8286kkaLBfFwiXlLt2NUMx6bY1U
7l3UOtRsLPa/1k7EDRs2c4Io4eHN4C8ot6mWAPV6AU95NOX4RUneVk0gBRPwfAPrfsTMdMLLG1je
xOj9bDqjE/tPfyagBCid5Lt3nQ2nkGYB0no/ZOAbo3lBPdNVsqDRHBbJuhB5hEowMD6NJ7UivdzA
4BkyoeHUdPC00Dd/UPwbfFALqUtOWe4PtcgWh8z9QYJxaMWTT1BilZVxIv/L9i7qMlLi+AywJRKS
3jHD75Spy+T4Wc6cVTbBfJbMERd9ooYcNKpxn1tG4Vcn/LRhvo2acx9klJnh1foAGcXhRxgfCBUG
cPekVk0FPy5WhePAf7R91Z1Po+1i0WolQKKJZT7G5BWUM/BeK9OzbSyzqww6svHrvkTErgLPclJD
QB/BJ3dEmLgBGTrzoaPq2raSTdN76QPxN1LDogK+QG3v/vUmWp1dQTQ3LVKq+12ABeA1QO6jY9Se
yWFcknS16eILMIc8MTyIGO/9aurbnRYG/fBmgB38bJuvLkcqa3saA6BD2unW9B4EpGTiuz/8t2Gv
Rs95k9OK89LNh3KXmWYIabB+N9b+gLhxQoLfzxT0200jOhlasQcv99YEw10jKz0RAX3gLu38b5lA
PMDZpgGneOjzaGmptDf83z9IO2w4oXRAdYouFaFD+skSr9G2KPmE16bgtvX6vH5z9TGllQob7rew
G9CgiMxC0BSEmxT+xtxF2F1cj6IKs5IDb4IGT/3v9MytVa3wk3pm29DAY+GtZttGeqG2uI02SjXX
+waP7OHv52sfDOFjcR76kKnJ9POv98YZeAhz6WSwYF0ONk103yGm+X+l5n2dRa4G40SMhz9Cn+dH
a8qYXTqILPmQmApKboyl10zpCIpaGI2/E5knKJT0yy1qKxuv6UZNLDiIHkXYedHAPK87zUvVgJYO
DPLg1gUyB2d3MwjOQkaROSuYZoslW+crOtYR4S1zHqlu674Wrn9ek0DeruxoDHudngy1iSka2ojd
gTP9AiRSq6wMxf8HCRj46QCpm/Jp8suRLdCk5hZyQoGlbRe6Kq9OIYYVXYS/Jhm4juIe/nnBgBXO
qki/SP99JCMuiESgZ6d4jtu+af+UmurVjavbkVuwaaaV8DX4te3tA0ZHqJlf7XxjKLF6CnGTtx6P
9pmNHOkc/kcUZTgoOxCN4R1cmpvec/b8KmudYAcSszzTZ5SmCR3dDdTtgzd1SPolzNUMOUdDiNws
YV//92pQQtq2q0/+/KXkC3/bE6/4PGyZbOVWydLUzuZzbaw4fvb0WOwH2aVoMsZ6grELnIr3qeYB
zSDGP6bb39NgLcSGcIiuN8PGMzMUHs6sqxhijGCFmajwuLQ2LWmNaK+x8+HRO7+6hs7IiGo9J9lP
SswyjeJMKbzQqzNIdEe0JhYLQCowKsIMFtu2bIwiL6AhN3xNnhZMxnMCId2037vc1+fKk67kW/+A
Tv1nBxBkS2Y2msISiy0Npt+cOsj+TJcFMxfF9jIjY1zvPVEkgqYqMceI7Le9ar4cYV8r7tmiZ3s1
4SFqPHWhkUcK0HHuRYUnD+KQlvU8lKTYVrx1Vi6acMfDEGlFjUu7Dq59S53urhxbxv+LrGaMVTRe
Iy3QejrnAgUZDwPjX21nRH8IAjFaL4rHFhBNzBR/M6XX7AKPnidGB6pXwkvDSQIJCJ3b1/q4enpi
rm+drA2Zswjfdwr5mIGHZCT4a0y2rVsduXiu0Qxr2Vfal0MXKZ4QLrHghgY1NdyfUaQQwrZzriVR
NMNOYARyYLDnJJqnHlIy0alGfn9glT3DjzKNCJpdF81x5Z9bJjb0vDO23HzA9dQ3P+Bi17tbhfTf
SuhyJUcX6Z54YZqP1AwtAGwgsFc2cMeM1+dXlekaN9d/ErblBPTOiEgszDWjI7fCzqE6Y8B0Xxum
WMVeclDJylglaPu2+3MNXsiGT4rc0L/8ZnZ70ZPs0Ak7Wg4JQfEIAy1TrVsSRLFb2D2fxICqVG3G
7GC+MbgJdDgo0qtiM5lsHx2Q35PZv/kMDPfnTRlz9VVGBHNgfNIAcz2cc5at6w9JwR8lJmgdUMmj
/p0Vr9C0sc5K0YIqcwMFedkEfE7B55RpG4VmcWlAxsUWcGJMmGYJNI4y4Ew2Tz8Vq7snjcam1DvM
LN4Rx1kXwm7djEUEHCtCSMerO/8nxyDmJMdyTdQ1v/E3KZvDdCnjyz1aqnsbBPGMc5g2mBpJOGkZ
lJcrwbxygItdgLUz/7ifp+pu5JH53CyMzCi/Mc9QhipOX2GKMt9yp4H/1fm6wNgAEmZf8ulRNF0t
jHnUXsWVQS6nVtbbRE/hWrGRTAceCL3B9DqTaJOdJhZ/oN8poUZ3vos5oEUI2gLdfiHnGfVRLgwe
AJbLO3/jh7swaKU/vJIUqYJ329PG/7mlMr2oYkOV/UceffHwP8apPo5BH8mDIP6Ha2pqU+ZNUqGJ
mGHsAIK1Hvcq08fYG5sKpzZzum4qD0dBsUqL9cGoQJLvslPGoPKUz+BwED9Y5dVt3qQyW0rBKR0Z
QzBsN00pb8qFkGhEmWs5Qw1vkjuNJRx6eBrNPYjS6w261I6zRfTVGV/QwndBHX3bhCxHdcHTrqLP
07mI3JLfnEMUgprn518whmM3+PWntvarmciFXvfb3+XBzZP48fyFfnkdeXeaq9MrhZ9fKa34Z5oi
EHiT6/SoAzz9+8V6ugnK5sJPpN6M+bECQGjC+VR++qqnpDw2vTDQPa/3ITaRd8OtLq+wneBVLCNw
GnGSSQtwRJ4yPnrDdCrfFwUm9gWFD2qhcJ9znZu+7bTnuBow9MzxshtQIaTZVjwMVb4OerleCrDi
J4JsgTShAi/xJRDVUlM6+YOAKfxboilm5apHw/5kzEkoXfrvlr/LhqrBbRMr1PGGPFu9tBv25Rnu
V4voRGfb189Sr9lLmVhW3U3Sj3wwiU8g3/BYzMPeBn+4PVxc0+HSroz7L6ydGgcXw/9kLqxJQekB
HBcx1pwqPnILWG2LehDvAhW1B6WW3ccpQv3asADiUwHbLAfHDtYwDZyiJxaQxgeDLQpibUQJPQbS
nIir8KrfO/f+bA6tu8fGqRugsI3+hfJiP2pMstojf40C/k+duTWzIxq3yZBWJYZksTJYYHe57qvV
lvSDvKEIyQJVFXV7HyVrhsFsDwH7eqXu2YsSwpYLvHIeY/eOm7AwAwrHJuCJxnb28ciUnOE1AegQ
8OuHn+Uc3bicyzrUtjzz/Wj6jWroxBggnBWe4bwy0Obx2K31dhrE+g47bU1+Stx/Qfd9qPSdRvhS
8G9d3Smvy+Q5kkiQdbfWKHNo0ZgGt5S+VreneQR7ZlgJg60UhJOfyGmAmKpx3OL6NRUlz004vE/a
lMiNP5ZbRYNoIh7MgPTdlN4s6FHJFkJlZXYcAZhar2oNjoGjMd/j4ZV6BPgfBBdQ7Y2I21nP6tfW
y/qSgXrPudk317VJy//rhUKIQvLFShHXLR13malke4hsQKgNHfgePPtWTRGsEWITvpkMT8a1OrUK
bZh/yIq40FFNJUer3Ld6EJoMy0m6diS2Wk6zcpGtFwpLnLxeuQ1NmR4PhV8ZaHcsY0F2ZfdcxxFQ
A3HUk2rioOhpQDYgiS6FIXhHVqH6yLt9zIUD6zdIqt0qLh1uIdYmkgs1YvIpDMHUaKDeap27rcG9
h7uUS6MXV4Z2oQZakywkZIkWQhMXIdHMlqrF5StqLBPGoCIqKcxcjFSH8MBTSBmiKVr0bDwbRpTy
RwzO1g60S4j5Mi6WQyQmqorB7cYyyu3eJrVe6+ZmBenjJdDxYZKNqC8eFbOK1tkAu/sTeihAwNrJ
BYWSzwkQd5lJ89BlDIPa9mymmZIHfYV5mrUfZzmgQGcoLjzc0BLZa7trfFJEraeSYKbNSrejtdLd
9dhRAqrmnQBa8Jt64PNPW1ts0Q/huiw7INQgPnP0jGi7miWaRgCDsiqJj+G+sKq/iRYs6Yi1aYIj
L4Z0lQWfBa886BOVI5Pn8iPTOiXE08hx0WUeyejBAi8hf2P/AXM1DBlLUejkFmnrWtSBe8qFGgIq
/+2rt+PpaOmOeGZiJoOYuEopTY/RtAZWC3GojYds496uDfTI1o/m7VV4KohRFrICIk6vIR2rfJb5
MxJBuG/sTYJ/oHTMwZiXg7EK2p6rhFpeJO+0lvvDCbUWh79wUaRUc2/8AOx7dlHCruoFkbMA0PYG
/yRs1ZMlvXmu9fUNBHp2+j6fXjQGD2sAApJ+Cpc8PUUjzq8cHA9Vd0yOwIcCjshQD6d5ESDwmPVx
DvUdUb+qwNjUmGxR6ZiadahAGnqJgM+BPGDdibqojt8DNKLXLVbYyWja1X3uDIP59UXQ84oTPzxE
mi82jJ8k7USu8s4DgV7FpoZPUZX/WnvYwDZilYfz/1yvhTKE9QbZbPEuevxCi0PlHkLH9coJD52h
htIQbZwmFa19tlSBg5sOsh1H6HJs+dor+X2XSznVHtjI2S4yuYiWIETP1XTuxhRI3KvPLDoTrgbB
rOu6c8OtbZNg1iVOA3jefJrJZ9lc4amS17QV9ywnsgVxgp+eEs0nRQlZ1zQOze2OWvrsed59qPK4
wksf98/IJakoZI1Qxz6t3xnyUMJI9SQKUyzI+UwHcpaDlcbvlkmB9LBYUc1t1fSso8vHwSCqq/4o
yk2NkDuuPOJePGZ8nRTifFo5YEMg1csJM4Iry2QYn7zrWegciUyWq0t5WsjMu1HEgp/W4CuB00vH
YzvSze+JjyMY1NULrVNldzq2d4pxh07jbxMI9AnNJANIETosLTCNbZumq7LwNVNCRizSLa0UDvpZ
TxH5GnjhsBvoFdnO7X+oSuSQTbtxuRHMb99cZKg8K6jcT6UREo4XC7e3tH6UO3h+Pelnb4+DTuuM
8GpGoARxslC1Yadzn3+baZbmP+E45brzabKy2yW+C6/9hXnSqrZ6JyE70ylLiYu68l+kCU5tknAv
jtQPKQ3xdxvMG0To46M+QXEtuvShdRNKEgfbKM/fz8Xh14PCB+7kJ0CQRINf5z/+qxbfkXtihQiN
I9SdWuHiZ4Zqnf8p2RpWjnaO7WQSnJmxZYrtpy+2l1Y1Qa4sSp408Nkjzvs3yFWGK+qLOZ8+iJez
pIAulVF6FsrPUWL/2utK7x7upFj69c4ybJPQYPpIzamq+4PEviMAEcXRgT6o6DpT0hnD1eDZoUvO
0I0fYSM4xKKyN35HOxtOQSI5GCr0cb2CoS2ICFOuNFGZV2U/P1offj80Pq0xi2dj+L0A6o9MUMCL
Tubm/QQ08cY/51rA4RzAOSXw3qd+RlcV9kG7z51TU02O3WaI9tnFsIj+IA9z324fhbzY047GfjRq
FkScwMYwbUFhDknaNXKzbvNGXkUgVy7BEj1Qd1i83C3uB5MNeTGWqtY8EZVUCuzPLs8R2Sd4wh6x
1KTl2nYORJwNX+jbGbMZMVSN1FzWA1sGLgq79KuFnAOGO5lLnyeSFzZuCRv3apVBHVDHp/54VxNy
ERsA7vl7AsQeP3vkdBO+1nl+jP3WYlSC8Rxaz8oloNpvVT2D0CXPo/MFO/6cL9V3TD5vnvOsH2xq
IAzUeVMk96FnEpGLOiDxc+wwQQWyZBHH+fFcSn7Otuxx59rvdZIqoR5V7ob/QaFjOeLb4UDAi3Og
azqqkRCx/o+38QgHHdpwngCVbBR3RNa1G5sFLbCzvFPO9ciAkAhfazxhd2xq7a8E9ftu1fafNeXy
+3dturqmM24HTLz4AuCU7JbkZZJyKmgIO1jVrTR1RsRXAbb4oibC3y7Y5LYIIAuNsY4k5QelDgAc
UiZMceE1lnFsNlj5g0jcODz7xQb+qRJDL74n6vupJXKdICH2XEycxHzyjPydspK5s8n0cp1i9w99
qZXcSkdlmU7uyAA74t6C7bwxkDGl7ifGIX5a6grxuqrGLKIxhLGTSfI4vo5AnRUp8TWgzZRAfV94
m28UZTdxkfuH35behad/7ylWfLF/sZTLP6TZRZunLzFPE2oyMIEqt2Cv9IFp2g4ygsgmouRwFepZ
nzfJK+LXO5YNdW+yN3oh7SkuCveQa9Gs//LUcuBDwm0CWjdIyEhnRAwU8Ye5i94ACx38fhrU78qW
PuGDFarYU0Cyhg+uVrtsgVdMv4xTMK+dwZS9v70k/WFhF/KUIA3itJJRvivphSm3jmOMPGrkmiI+
kTvLaWoUCNj5M9XMKa7BkuCIyNMNxAVLC/SGnzreRvTZd2Pn91+Wwu/RbrGjnaEQ3uZv+dSID1M+
grNrDplYMXldDLtiEmTX12tWYqM0YS5e+8E/1jeS8wZJKYAsawYFG7Q/Jz+FpLlRRmZpdzkf4gdj
mRljuBqzpXWUkI8evuomINQTFnpduspNRHg1TgLDrfNKA/H5GFJL7RjGL7uQPwrBdGJE0s4xU7Jy
3IlKMB6iJhW7F1TU3q6rSVuSSgXCa6/94eZuI+eRWgVQgHSFlqQ7c3i9+IENsqaE7vIOOtHjp6VZ
T4FgS1CanoMs2zfQadbU4j/S8adQhWQ7hX0rucZdd19G4zEA/kfia52c544p3XnivOmy5xBtOHaU
xap3VxR1NEFuhWE0CLb1GMNQ/5/nEIKS9sTaQeh0PJQw1KJvLFdQawdink8QXhQ4+1Q/tmL5fgL6
DUKN4qlhnazrN6mwCcXxgMT4PWtxeFCZYXXLXO8yzRhbw6g8BAyB9qF51pa+Hw4IdokGwmz9Rk0r
Hlx2j70CKsqu9mUr95YEo7UFCe/eot2lRaFpiPguBDoSexhRija10DVcuBaruit84/1W4zaa9Bwt
vz+dc255VFbZ7JR52c2vR0leU8CUL/kmdaqFT/UWaMqOaHDSHSUXBfESNQHx0fmLBz4XwjZSBudk
axj65QmFM75iXWb3G0DVYEt6YavLL4fwvylBualATK3GB1BKrKZinKkbEX7NOYwBrRnjuVMvqHiB
hFlVyELMNj4Xnq3FshhGrJ1ctlAwxFxMu4QF3A4/CWElk+lWbfVnyE6orw6i0lzj5q8Pj2vGZR+s
cqpIkvk/4rTHTAP7iXSwlc1l7UtUN50oU3pqSxvFpGKQODLLLPL7KUSgKgUaQZoLAeQrvKbUzQzq
ODNoN4JeoZQPnx4XR+BwNOTcVgPI/wo8tHlfEwvqQScSxQKDR0bdjGIVXR+Zx1ttEUlUCzyL9mhP
IJxYrBhHsIqHtAjePbQtKtcyq8dhrnSzsYYZxLT0mTwabDXYxDMga12xRgcwaHMPVpnyv7DfC0+N
ElswnqJghcWVYdmni2gj+Z+1s8Eg25HIsKR3U9kgIDojozzFntETnBNVZ5kqkxOTdtFYcjYa0hXO
ukz6ukdzy2eJJvJrPtIHwMhIAVBAW0Q0WCGJmv7lpnb00S3orIuzs9Vbi0pk4KmCEQ55IVRhjyy1
x1XDmxW8t9/F/kSDJ+4LNCISscrSQPkWIvvFWQAoEtKnARDv/FkLYwqprXdIY0OH/9gvbxw7IW7v
8NSitA/c2DlQ5mJTpAxob+Bfji8E1lBBM/2A1yJLgY0Fp3nUNUJaoIn5b7NmtOCN5zkieuCz6Ot6
09xIxu7iRzehsPkkvjyzWyww64cy2aAcgPycvym/ffJRxXbp9ZSKGP+ui1+aZJCqhyWwi3TA+IfD
8cyvjk3wAEvXXGpwXVYIpxXp1EeCQIlWyKspyHnCd4fRtiXE9osBhbWaAwHsR4zQ7mx5ra4VUaek
qUUnhzdVYKhlZjwGZmu3LfP0tydj3BlfUfemJCuCVtXZDvRpDZnMnHwShGn6nDfTVs71uL1icra+
YHkytGPk+QvB6k/Yj6+aZ1HXN0qQBmxrbam4H9V3CD1DhsXVQXUXaswr5QU6WMoqbKhzn1ODoEGH
NW0hKsLLeEv5AJ3Feafn6osf0bfXxe8wemqB2IW8WCS6crZAlz+wTaZVwRr1UaTEqWT7aEzPAKh9
U64fcim3GvgSVzZFL4e3xKB/7juga2iiHcK2Hi/eddFsUjr3DryhjShYS5RjHM6UJ/lMXQUD3Vkj
ykWK0jn31HaFyvP7G8wmLTqjQvMQEYD70UIjSkNu2PGJZ4DKUW2xtKuEJHoFtL9nluCxsvlt4+pB
1admBb1pZXbLYJMHeqv4IAHW4Qa5JLWYv9K9tGhmy4NMqfVZSg0AnzSKqMW/UHLQNGJAUY8ULG5v
W1iWkiR0WPDxh1LxmZnzabDxyzDv1YSoAW26t8+KbsdCSKXjyWZSLZdaVhT6kXOGi5e8hlA7bGiH
j8ZXP/F6JwAIpB+tIuepCtpRIdDk39tCllpavxrom9h0crOXJw9sMP5lOH9atT3rjZYSHeg3PHSZ
/UKlkkHJABXSH8bAZ7DHlo4NiFKiUXE35HWITfepk8vjqhpfJx+tq3aW+umTemue39ZpqqvKg+r1
BtLYA3KbFhodTbkwy0bdMfyryNg+lHoiScZX2of+o4Ui/wHQcZSilWJ09kqQ+W5/CPH62ET841mm
4l6bLt+GrTrffIKLqwpCHHG1MS9ltdYGYi/QERStT/9NzEMquRyRUIM9V1B2fqVYtE462JoBfIRy
0L+7XcgOOTwpP/KOsJBXMMzOLdqu3Dl7Xume0mAgVfkXX1EuGSLRABR6Z1JN0VQ2OfWWf4/JrR6A
QE3IL6FQqmpT1xuMjYnjTVNmXI1HITc7YCok5ZC392a+p/iSq56XIjsVLERkPiNAaIHuMsl/T/bl
UORsIJ0Q9cAFpEwJT/Mj6BS6VYWM0HeVIWt15mc5WAsg76a91aiLSIZ8L3QKeWdK/+ohMEbPg7K7
ifznv7DXwa+faEIzD/WVTmZjR7NF+XAd3qTHok5bZZ1rvXsRPeEnzdUg12/TxUSswKMIpmnUECXO
Z3wWCPtm6uXwj3nUO8MLD7szfRAnEDB8AgAph0cfF5qQ+iqnKpN7YyXYB7uDppVjkoYKe2eAVeKV
x8uidTGGWqhvHTLZkayEIZxL9KDqfpGhHOvD6CS+xvoaocp2jT39lSFFaWzYhHcKPT/pjjTGFFdi
ayZe3N3uUd7yh9nHm2o0PfdmpwRm7T3ZKxhWuNEKH6lfqrABJE8PRTW1sSIvwTVKg434LdHU3N6J
KiY3VTRcdrbq1mVonTvssvWbMIh7H498ZWDZcMpcq2QWj/g8xds6V2zVN6W1k9NUC4ZmUX1607zn
sAjZWLnrcm8vcT1TqRBUP/ZbMHMChSwx/MEWc/Q2weHfmtMscKEEp+TUXPp4N2qTgWbm9knQhUpM
aYLaBW19C28KBFyHq6ku+jazbj9Dk8st+nwrPqCF842iSawF/yc030RP1ensOykAAATFdWEu46Sh
l3DM9vx7JvwzcOMEePnN61YJ8S8ImxWzOa7x1d2ypbX3jtnnQtzM0PhWuUtCs9RRGGXnrJO0BFCj
iwgjF7tiFXKSmxvTi54Y7Bm6nRq4SPuFqO3uL+zVoPLUs9ThpdvsEPRV8lfTdbc+GKG2D+4SxHs3
Nree+FSTzIpwaaMfDlXQE8SVk3HfJRw3pnImUbZolSSiMXegsgQ+X28YBn/3B1z7OjefpNUuT+sv
+dD1b7fAJ7PCzAAZc9DDEjlJgzC93pG7C28sCuEiNhE9TYG/rdbqD7UGSbAMYfdejb9aLDW9O9Mb
z67Jk7jF88i9+q5RldENKQsCrCE9GKMwMXK9OHXpfWpzpHVPdCXkkeCDYDG4JCZF5v/rPdA557Sa
iRJnvnrnyeoxrTSQNHKQj/oeiTEx2d7VhUCmMB7mb/TIhael+PhkRwK32b3/BCbzFktf2SwNCW6O
Ai/rf7hAOg8QnCdtFlvLZymCv4QkjvhTJko58jH9y4e9imXGKlea2nZjf/hELDR0pLlPoEiv5ZAq
CtVx9SeNYNoEHTxvje5oSSyto73r17uLCv3ySLBc90l2R3yznUCrJvDqM/wSc6x4l65SrNE4/y6e
2B0MTSKokNf0ugfFUOMO3jm1g36ty9rQatUnLIpdSYNZEXWikQIbhTVP3od+y1HHbY5zD81mZEH9
BXyzRPqyW38gTaM6MF8/mm6uIuT0UWbKr0u8xTzVfUamIWpY097txKulfenRkc8VKb3mwXvRwo23
mtcvJR1hIKS8kVG5gCINHo4jUh/J9O0JzI1D5/ljRP8wh1NI3JBqTTwRmJYnSrwovFVEFjO5Kuvk
V/14Cfb6Bp84BdsGDm2kXO83J7YeqxC7vXQdvEvszIOzNl3T20U5MYvq5+qPfkaM/ATFpES7NYSg
sWPV+u48ibNWdSTLUXSGMlcjODzVxh5a0blrnleDjNV4MJEugIMUlcQtl6YAvd//PCJTuJ07E0Lx
glSn64+6wHo8Sx1QpIqk4RxH4N6/Vqytv/YM761i2SdEOK+QanOxmV7J39BOe/FugIQ1LsTF6nPQ
0tP2tbNPgJZbce2M866DMkAbfzW4jyw2fbZEzPJnXNLmRuJTBdcwt6AMk9ALe63URdSNuzY+qf7w
mkHrq/Fv9f496Pg0HT9QNBbfSpV+XCjY+EUJmQVmZi7RX1UQPjtotZ2SPhmqPHHLHv4qUhVxlnc5
QaRblx4+mOj5acmoE3Z/FtLubKcBmvlV9EsUTxh5oDmLxGFXadoRSBgfoTcv7ZOmezvXw3kVabdL
PsBhVrZ2zIWND4FZA6nUatw25EC1FLMI77hN0aIi8bBWDLnQOfpqZdshRKsCNNYbH+wra9fh2or7
wTwyGeD1nAfvPYsJ5UoqvEmBOEcXxXoNPGB+AbqE5KaZT/JU5duqSzHpzyl/ML5crZX1MMjupqPe
QoqPX01utDI55mgQ/3bj45PisTaQ+EoBpluMdm1I/S4dBKu5Ozm8LMHiRWjdjpEPLGvH0Bx8MQXH
bRmooJxAtE6mNQ53gbFsPsiaP1jkyKaQCwdvajYvWlWzCA/TJ0YpT7UyHHt8DhwYr2RO6rmq/ERV
i3hkuhIE8kiR59MIMA51dan0BISRDwWkp4moQ81exO7ojSAP5IAAhok0CU6OJjSyl0IqeVl1+qRI
YoLedGZ5dl/ohNxKu1/wBT93115x4sVdz9ODot9Vlx2jUqxxuBxo2E3Fq+AVvs+YZKDBJU0m3+oz
mhCVoB+mcVG8deUQ8LIojmzU9AptYmFVpfi0quIBZ3Ly9hKFjObVyX/yW0TXn+jG7WBIk785fFqi
7eY1ucGD51WjbWE9p0Ay1iRFdRzI+6KsGWLdIDjZtmQiRiKbZEiXtBxD+gFNVhz74ZTnkImLd2BD
rOjLXUvn0MhR49tWa8f4yGX4eDRJgNghpGYTLT9wcENcCUXzrVJutG160YKza4UisGT03JOJngO8
QiMbeYE78QWThtlKkd3uEusOGQEiZmXjgWugEV5x2YyHlxraBPTES54+JSZlFBK6Yt2g6b6/q6Dp
0+om/sULDlVmTz/K9swHIHZRFbka/S+gqiXr69DUmk+wh2VsxQS9WyLoHK+cIv8NShhaIz+DAg1t
BTF42fmrkaK6zpxWAU4Bs6Uwpxf/tr8GJBzAzk6zpHI/Ir5+D2tBzFTkVPlDNSSNju4ObToNPj8A
VHgmya1s6Urffqv8y4OedyMDZhG/IockbxRfZP+eYRMA/PdGjdxW/zz43x4PkUHc+lvRD8ScbRes
rQoIC0tdf67+qkAhC7EKFVjfPLSEMjZ729bJyEELV0HqD30w4Fn+VYPs/tb5a4LaKCxccndg3QhE
u2kmeHIW60La0uS9Yk35GJzG30CjSTKKAKMGz2UOVPSut/5XB9+rNnxNIsFQQfLDW0mOHDirI/Z8
UJxs3P+9Y67BQFRCMAaC5XFJOIXo23LWFB+u2Lfq9x2IjAnsatSSSLf5X+lA6+bzKGnZme4YiHFK
c7ki//UTAaevHrnhSPXryNoVLRUbsU5J3qAwD9jYV3H7noANtumFm65YW6wC+oay/siSo2DR+680
H6nPEwthdIY4eg+St3Gk2URSLE4rrs3fVaZoLyEVxHOZi64sep2NBNq1u05mvnxHhkxS5MdipRk3
HVHW2LuQyafGYffvM6yVRts4S5lD+C1G47wWSZZGkcBdu0KFfplRn4rSe1+b0uYhRfRHTKTvvhU5
G8SwMbZvr6VvXoDKmM/1FoaR1dWczmjcIUrC/VJSy8EvID0ybSSn9KLLO9mxj2k6cN/uh4byu4GR
lyDPMG375y+Dt8H2dawWHAgIKWbBO8J5+pRpLRuoTB+RbKZb45Oppk/TarX+B0YHkL+wSSZkH02B
HG8oqKeQoMII1ZLVDMXancSf4eYUyHzLq08lvYAihf/5oAnqDqoWz86Jhxs3Z+pnIPfxhNha0i1H
vZGcNeRizr7rBHIv0uQJ+rCezI9uan1kZpRFoDMZvG6IIibhY8cGZUY65y3uBfF4PYb/+Vgp2Gko
mp9hkcxtq35R6JXmXc0T+Hw5yPGBgJUWoQTYlXV3of6JOnzA39mOAcdtlL7p7nz73qM+0tx0h+Tr
FdExktzgbMSALsXtYU0x+y8pxl1ruGDcelkzQpGHqh+aOp4VJBbtlnvm4UlO5DDi3kaGc2ygz0ut
aDksD6B6gr1Y9rKQDK+ycWggPFFgNmPVYBmo6wJKp6DKtzPaPzdruUwX/wuFmJCJPyqOnwU0aBMJ
1oVYYH4t7cYCJyJOKEVp22pkEfOa/FDN6z/JV9LeEHQrfMZcqWSYFh3Bfu8JYZ48SiNQfX1J2ZZe
YdwN9QcbB7/kMB6rhjhqYHfoFOrFGLCE/TyUkGsnbWFyMOxjGxj0zJet/dSlWVlmeRXLcCbEyvDl
150KVlz0HRf6awzxbOb8Rxlyj33nY9zfzRSVGgG8kHCcTQyv0vKKMioO5O3g65a6nBMfFMuWvVKW
S8uDXLoeFlVArVWLnwllLhoCN/6qYiiJRFOI5V7Iz8pmKNTMvQP2HjPiPzdw2ovtvRGKostxfCYz
hefQQpnoKTGNB9CMuLzx0MUktO4kJ5pdape91vtpBmuXDE36klKae7dPnQv1y33PPn/VaDfgSekD
KWvkMCte0JCuJ8k8Ni8trOZf7uYuBxnhyR5MmnagEUWx6PLZPd8iZXdJgqGQfNfOj1sncdgXO9mQ
pll8VXDZ4AalXMeyZ7+VCmfllelk/rOQztUJS5N/ggMT/RAihMuKowoDTnh9cIp97pSGU+Kuuw6k
0iJIuVuZ38pJLfWvqrl0M3SzIchsslxWmHKvbsxlp0Us5KOMAqLshDqBBDCzm467ANsvnvdZoSTu
AckjEzBTDptpPTIPKv2ujOnEY2OUwaDe6ArdeMA6bCEgc/3c8uP0eeaVhhg3lWPGplepmbNLY3n+
59SkQAy0Sl7lzutk7glrqLsgHBBtXnfhyBABCzFStITB5fbcEDI5XrGEwqoCiduTdMNIkRImNI+I
6YTDcN3OpYN9D4dHWkfP7tZth2/+La8p/iWCXCW7/C980BeWawfLU6eVuQ8unzKi5tok+DSQfYyx
bQmczW3uwByH12TqD2yFR+MJUt/nHCS5ZykYjQm14c1yVsxjq08/0dp01BeHHJJtMil9l5iKmI2c
KJSXS9tXaOd0nd54nD5olOK5qqBqDWi21/Quctk2obsIVQ+34xhVRHV6L16nMNsLMTJXvqV82TE7
BOyJYH3NlCQRHxa01zjZOO5tq/nFWYqSVtV8fBiz4pngM54z7YDK1RE5RlaijQcHjB4mGyRg6j8j
MRIkakY/UAw3iN94IjVWvgA8nyCBAcXoQN4+juE1hV2CZ3jmtjCDz2XkY6Eej8Ma9bQwO1ZjhWWz
4r3EVLedBahrWOSHT46zIF6Cd+6sqm7HiAXoOD27lhv0Ju/4Lw8uhqfq97ksjrXkHVFxfQ0InVXo
me+zUgG06pyjflQ/y8QLr8beHf9CSN+CEedCMmjcNdisfVQEADIRSdgxY6QKfHnoCRkJeFvywNPP
XeZGiw2vFngB6O/2EkiMrz6nqhgTXIfOr/1l2o2CMdetOF+Fy6WgkiBiZowPzghBXafw+eKwzwvR
5vOgQH2JB8DWUsUfquUD2lTJPHXFU9m5yYz5IGybZAHgHwyk2moVtzgKjF0CB5NW//5KaVcl8OnA
nP0s+XZvIGIxpO14/tuvIy8jYAMaEPlEeNDz7GwgPF1wFyDnGVSwx4QK2/WL6lRSHXniGz5S9cZu
30KjFmRTDwHzS/BxtEgRMlhCUmnCTupW2G43EZCNM7/cvDHXnTOjAYdy813F0JeQuU0S41K9qyDf
Fhl3NezSh0789Emqv9USegj4HgdI5DbPNfjE/jBhSkzvHf18X6jLxEYgzyQNm7I3lezB6fJ557XD
xG7jQRxPHoeG9kQI+9E3GIFKS0NsmZyHdCHFnkQexW3u9SVLpaKAmD/8noiBWE+I+zxM092gIBPj
mBKL6qYkftNfmpxnD/raR6zWJO8sIFksI9xcr4xYnK0KFeI8wdoziTOi1eosoKi7uWDSO1ZQp6Q9
rsUwazLXGUDFMLIyNopVWE7kkNfYPB8kK0oXTkvzvZlARW61tQ1u6GcyZFglNqkFkG4WsQ6I1xjE
EX3twBVWSrosTefwf+QSN/hV4Ss5TsSPbzdWX66WgCnq14YOyOuOS8zxfqMLLA0qJ7KxpVIO37yd
XI/3ddyIr0EW5Lq5KfIPGccXaq9M0CTc/8azmfx0XVlZSdAAfwu6UGoqrGm1or8MS4LKBBMRwu3X
VX8kZkzyH+rQc/SGgj3y/mXjODa87gGwTrUW82uXaz3mmETG4vLWSz863105yySsstQf/CzD9NEa
ZgfO+wke+DJLpPCkwlYaV70QTstFr6rRgu2l81xg0M+QszmnO/Wu0ZrCnuJMukmwD1Kle9HlLnn1
PYUECJCZ+LYZpp/5Oty+pgEbZLvCxCyZ3LXks1V4kCDfa6U4Edip6AhEkryX/ZsoGehUMZVLgNtI
sHP1EPgeyHIf/wIrUSV/ZIEMFzCFZOpX2TPcMvn4+HK/XoXrKDIPA4D6IbWbcuxQV7yFB2Ee1hd3
ovExaUw6KMw684iIepWchJAb+4AexiwVKyqNz4wxsjx+r/i+Hqc6WzhhpiAxz8l03Bdp0wHTOers
qJbF/XjZYJNntdVDRAufH1IdtXbZneLSrvt8tiOEMazuX/vHGRJpGxnOOIAhA0Hcc4gdSL4Pr9L5
AkxbeP/8bpOJYpNoVGJXh5RitJTPaSg++PTnAXKsPMuQpdlAV6ZeSdPBtJOlWvK+wflBTScjtRUb
7pcwn34b6iTbCF3on0UshW/564Go1Fy+4Z82a5ZckfuCLXE3jJcbiq3l151NMzuJKfy+IS8CL5qZ
G1rYyvXR9Hbvd5oHY1ry0hh+QHBxcjW1QBCuqjRf7cmirrFffOM7M7fiXWeeNkodh1REcCrdPK0D
S5zGkMTQ6kd2VNhXyvvQtOsGKkoqPU7B9iVcUevKBIdp6kZNJ4JhiX12hN9/mtt0cpCzls42Gv26
4Dlk5pTlV4s8XUiITDStw9ZYk1xzrRFicmmy0/ttqZEG4Adyee5QDvby+HC5s9audQ7YwddSQo5/
FUW/nlcvWSHwuVQb7uCjoxeQT+T8QeDCImAsDDqWCYWgyCuCwchj77lYSJwiE5JB1f7Yqr+iZ/Gg
KRudw1PSVudp1Lxvu1nuPPfVhWz6Hs45KpdNfdmWSMU9R3bYekLLKnzQi9+7kuw2dCIvXsoXoH6Y
P5HpgxHkV+LeHqCIvCYEpewK/BpDI82H+Ygw5Tc9cyaPPhsXu4N5om3myJLfUcs0O/kbNLTe/39E
KyawQa2a0Q/FBiXWrkeTm6ETM/VVg4zMi6DVBPaJor60YDF+EngQQnKr5/F1QjkgGCwckDqjU6R0
El8PBDPhAcHXwQhJovKQq1VnyWEFs7ryaKTaUesrjrk9AAXh5JuivHI96Ykk0vc5YzjWHaeczNrw
C/jcS4dwHRh5Uzuz8Nux1Yxl+MYCyjrrWlyAByYzvmCXRcRkcX8g2fw7UP2+j9yq0HYSUzvzdul7
/EhmugtiaIjEx+klTGe3JIFufG/A8Y+xbYtdT8OeDXyj3KEBxdvgykdu4Kg9jeOrXccW0pz+xKJX
VObwy0Zs8UkpF6bIKPi3G3R1GNuGBW/4HnDXLODAxrLRVMvT409DhoVhZLOUCjMdYHO5fV3xD4YS
QJ+djxFpvT2x6VS0Kh6dU4R1UMROXdZ5LAJPD9kgeZpRsYCW6pwB0gWvg0FLQn80K6J7W0PM5v4W
x+u5vO5f4oJn2RPJN1Ornqc8V9r/Ha8cyni5SU0Z92/srWxFm2C2g2wxuhpZD3PHSIoRbQVFnB1w
quKWJmbAFyZdv/nXYVp0mbb5yrqqT0nWGJFcA7KVfn9RdkofU0PfEB8+hcDcmS9q3hxBgNIKPfgF
4h3EpKBwyGVCG0m2wgS1sCr2jHd40N9ge9R4vkWjcgs3BJ7gpoLA+2gpYsU3P9C44KyY56j1TYGX
9XYUb05tPHHYxffOrKuS+Efy5URlHDwuucsKxkpcu78rDbGvf8nCDJRBpdbGlB2W/33O0Ve5hRsM
s2E7SjPNEcrAa3ekw3xEovmgvkODqaODUVTO0B9cu8ZwIUFDV55AWHMXQ2wlUXEb+npvPXbVy2Ft
D2IxOFoKSEtdGhbH99JelC1PrMnnxHuRdjpDPTSXmzo225lO8kMPh5YgcorsdZIw/XewW0J5TH0C
z7gwZ4l4hOL6s4O7nT46+P0w6dwi4y2GfF4dNHFive9Reu4RTyS5VzNsHhsJFywBhMxNZTQTbw5u
Daux+/F9PcgVl4bThIKN/KID8H76SBz2+fBWch81JN8nTY5Gi+jszolJtpDSI3/ozmiwcwKPOImj
NenGgpRmhl0zPLYZdp80KdF9Hn1dY7HEIzeTu+X/FuTZaXQbdh1phZ8us1URe17zDeNiFHwApEfO
f5NprD4cIxW3J2GuMgaXI/48RL/c0HtK/2SG+1VQWkc3XL9T0UdE1UzNHAeYUrPbKZkAAIhW+uOs
sbZkqVOyd8CaVpqMbgAa/TNAjseUbnlcrUmWDRWagtd/1Hgk/1whwvr4drxTQP0MMLbmvHA0tVvc
jP4uac5p3B4j5u+Po17AWofJmAY0YWg/IBHYlFnWFx+QJUopdRWDMHJ7UhdKqOzBio+CeQuYJvEr
eIYbC8AntpGPG96AGhPKBFgZzuJfRlZRK7XZAan87fd54n3JLqpkz1FV0xIkpJ7v7uYfto86JgJF
RIvEYD/F0z6EGemZxxDqxPOwCKKQTfee4U0T4m+2YH4ymhKwAQwY1pwFPXuAwvc4PD1tqkchTLb+
tsI+t1eQ/SYETUGqNBiDtmjsOEYYzpXeSqzI3YOqUTuto/2xfEkBT7fnkIzTvnYKv3V7Ulb4Z4fS
IwpAzrPtSzpUrhAlmgczCYWn3MPFnY8zTBR7TcQHvy+megIk9gYr/QG3LFf9l5FUHjyD272sQLp8
oERWXAjDkr01OL5yjDnHW/vGO7R9TDVCYn80WHI4p9sG8a6pectktJ6bef9olxJB4yt0IzwGrpCZ
ElgUzHHiIoFZ4FgrlmeF4LPrCCTEN4o8wyg+xo0XdOAmTD0YSARgVCUahB5WzU8I16xWQwM09ad7
iknrHtBS7EajIZaRXuCTj4hirYMhv12NFPOsKHxoBJ+D1yu5ykGKSx0FEJ4IHdwcBszW5O/ocolN
k94BCKypTvfOtkZ9fSvFNGK/bA/yEQlXCR9KKvjUaYv27z+zN2zSOyLDjHGqmhoiDMzeuJMpt6mm
rEFozEMdeOxvsVwejvN1kZ/160viQ7hHB0/qKF7hXhUGRGhu73spYZuwdTROI7TRnm925Y/e2+9C
AZbbvHd+GUNSkLaD37py9C9ux6FUsWXJueGQ307Lq26b9oaHWqvbCkxl5KPAy1zzCxUru91EFB9X
pR9zgW3jHv56aAYO7Couv/fjmYYP2Nu39PRew9/ccOlNoarGYZoUjOYVZGaI3qirqLDhuc/JaiZC
PUO5K8jiCJFurqXl+ZTJfmc7KbD1/2sUsuOg3kYC64xYZIkrc1rYxei1UmnOd4HTbPNm3GdHfWUH
ZFFkMEDMm0+K4cQjQdOQxq1ccpjyqk6Jyh7ZIZjI7wByQnP/7JB64QVzWs5wMHkMByaT29BqRFdu
S6HgLIlOdhZnzhOY5EUKz+jefUyuQOgSX19TTgPZXYSRSIYAVkFJY/yNPSZAbpYZK8cjOBNLEvSt
63fxP8Ml0SE5ubWDzDpYQzU6qJbwkDVhXGEhME4QPoV3ZaZ782ZlaBnW/YYQLNLaLU0uUNOUvJRV
R1IV7yKw8PyE89HMi4LZkmREVcVxS5pgb2fffrRU7Lm0+31L7IC4fsD98EXju2ev90OqVHJfnUFa
pcVeBIt5xvmhi39vIKoTxAmznWxtWS0ZzZ8atUgPTfIRI1O3D+TexJfXXou2BTCb6rUKhQPTellQ
7rUBDADC6qGqpNTjtDDlHh0czoyMNgGHpT1KJwf75RMcWMz7lcxzojam+CaRhXw/cTg5fpdgdQmr
81d4x9l475B+OH/pBwniJSR+/RGBSip9SCex+VtwnEijN4SVVQcLG28OT8szDHK4VcVwC3NJDGP6
gOhcACZeR1HfbDUD7cSDDyh2OqQ4EmaFwr0jYdWrr0aZrDcSrRkrhDFWfz9MODztCMuMyV/3ojDh
BMatPPxpwlWcst/gY4oilTt2WOlkSI7gxXLRMJyOdcaqHfrvPN1myQgd0QwkwcPtQx2Pdmwh3wdv
lMun6yN4l4hOHOZBB26G3eypRQB+2yNl2imiFz2lHQb/J8mnaWDEMhpFjok8AEdS/o6NnyzN3NCQ
ur/OnOwNhhTPaoObgBFBjzWV9oTISejtJ2VAPYYOS7n0cx8xtXq2L2WIbSrZHNykb96qh7MMG78c
3JJwC8SxmUTwhEnIVlJbz+FHNIEBzx2TCFjDiIgnP60Xw4g/bCyo05fO7v5wYAkWRy3MebQaYJ1W
ny/TwWrGROa2H614uSjvrf8rdglGqsmwZUkIkOuECKByhSD92sXtnhczPLXP5XFc+lO5VxRBgfy9
TWcYI9FbypVG7CSba1rfb1gPiDdmB0S7cjt0CUPKs1/H0t9IAGudC6e4OsL/5Fokp3wALAIIueDK
FfSx2n648aNGmizeQrjyYKqzaHJL6tuRvKU5QzEUcrxJ8rQpEJqL4oG4pD2MfbVyfHfEgl/fTiw5
gBtV286yntaAm5a13QItsB61Ei9agvs4QwuHFj063K6nSwIbXUjwONQW6a2KTbos1vje+uI5QJOt
GZpKy3ovq2Wn4ZYUNvkrmhjqjGiSDFUwUBX92OcdwpuOfP06ppiWLtyvQd1pz9EEwivk+2LbP8Jc
6eflTYc1B6TgKMwLjYX6SLmzcGxtMM5gj2SVRQ1ZbAdc9Y8PqKHdAMG3uA3j8d46MiwXb+D8w/pu
HqFHXNSmRQ5FOvt6QGGnsGHA+Rlk+7qQWX226lVTSyHMUtqwa75+CVy4dx/QpvCoTU+wo3SI0MWe
caSMHgnEkD6RZDCiH3bvQHFUkdy9mFbtaS5cMp6kMNnhCXXlGZsDvGbEK/U9hzwUAhuNwKR6nJZb
4dc+3Z+chDg5tiEbQXosKqhHVPp2RjQRdeIReVd3ohXtAReN9MDhfRSjlb5VWtoS9OKmNu6ylyRv
aE6gYKWjHZmgJYDEW5WS8qNo6+dogNf3zyjRy2hJOVHU/4EQst3YyDff2J6JpnmBHP8FcAirnWMK
Dcfml5sfGHAxPhZ2lUyzMPiXNQcAwpO89WktxpuVrrM+n1zDd+TeJ2uyRMoEwi/tw3Jv66vYtlGv
JSk9bnxgLi8q7HleENYSotj/Y0YnZU+JcIiFAMMuIzeXqcnJUcN//fQfLx3q1CYZiL/cHx3ILh93
2UsfKbhm6wGS/bmy79NsrEyKEeRWLAoxa9zaFCg5xRSaQUWBLLitDTEM6kxknEa2dwg2uOaUctzJ
PiFnocnZxMLfaAClppY/zTkrHuqnD0+yYm+/W35CP1Mq7zWkkkIxiR7WjolrDrqB2Rym5MvxA2G+
JAaaJEriRS88+heJhbJ8mluMkZXJf2ddaRX4Qli7YB60hvBISxNRSUk0k7jQ1QD+Cjg/fKB0u/9U
8ntM5SNyzwPSFwWKchgRcwVwLq1943d7op66Ps/FAY21rxMWJCaxWxSj9dgIuaFi4gcmjSkxA7s+
LVe/WGz68R+2MeTeIFVOoCdo1Hqkz791C9tkA7N05oiZ+wkClCNUQqvjyzvTOdAaTLyI/oYNH68+
2e5tQFsD2mVS9V/8Gp728wL8rg0dl+86NfkPRNHBIhT5s3Ho9FvK2ip7hpqB2LM5zKGwnvBfvFkR
NNvsgAFwOYX8Ij+THYepxD+oV1/hBEQHWdXi8lA7y9AyneeldKU594ku8/TLDblSknLSdWVe1Ist
yHo/+QKjn93Z7tdRxcFPAW57PA07vEjYzd4Bj1VhBzAbN1uREmGSakXBLev141GWk1vwp/RvotLB
PqgrwESVG9Poj51n8Odr+7w5K9+laqRAF2BqSqhGPoO0LAyibX4Wx4JCR4elBucAH2ZuWTHADahj
sKdmmMcZvua5SgQ2ywqMMqL31H3quA9f45Ygek/qTHk0runIDkQqvahv4oHtDs+BVx8mkHYz+Zo9
7SfeMMS4RQhFRNJtmCJLy/JIcfLYnptNUFaSkAenhuF0b0d5ZKdrBKJxpxyvAczGVcgDoQtGyfYx
P1CQ663U7F+T2RV620fLSskRI3JF4jvIQ//dezvPH8WG9TdQXldGS6vjccYmlgtQijZugsZ/FEGi
lNIEPYismxEC1Jp3v8rCqHM1ndssKh/DTr3dzVboOBgrooaexcX2F79SJndtspI5dvMX0yaUN4B4
dZ3y50zF5PEP+F6vOkrrjYsxgTJ9tVy9moxhBfOu7TUQ+XRkzVpN7/QvGqCZr36dsDAuIgqcr8dq
OiX85gvG8cZh0whclloetdPar3Y3UBDcNvLtv9uj744OgVYy1kqV58f2nxoL+BR0HASoIqcsFK5A
SNT0cKRmbwbUDRi2sQ6hT2tjnfZKPwxm2hKI7etvXFas3pH5MGLoSuH1y6CahrvAZYyk26YezAIl
YJMYLRFQ8yfZkXoxGuGJBHpIx0ZzE5846AnK4huozqJb9vf42mKfrwwK1HLVM5yMY7xRpbrOrXf6
uNztKt1LSxNizpkYMC2+tvG8v1socRMnI4YnNY0yG2Xbu54QcPlnSYy2Hz+GAq9FvsGLjfX8Fi+H
oilkoAK7wVkH02OjdvX5VXfWhO7pgpw0URcffe7zP56zwjG5hriu24ytjtTh0JHMQLNuOSO2L9yK
XsSXpt6eNrKrSrIXDQTHVu9rufaUubjlsYiABrzrladF7AE9Sh9S+RXBYjXcMJxqpQXz9dejxAAz
1n8wEmoDA2AM1T+4QFBQ08Ectm6bv+PUW+cp/SdUU4M6HZ6Ybf8Lriq0T0zSe3ZuD0SGLuCBiN78
tCq7/8UVXyCbZCKDknQQ36ipY3CjeMVJFSe1AjHqY3qm5FEaMtZKMGx4abMfpDGWgxT77csRZK9t
zqhYvhIGQWnp7H86FEDwsgJoVL8ajgtxaXXA/hMSxuP9vXTjXBKi6Nw+mHXovreVME249fFGzlvl
2xb4Ob2wACm2IshYcbv3gYNoU3glx2yxBUxtXmawdDx7kfdEP9x72lxGWLSs7TYWBRvYMoDDqeIB
FwsxBhDwIWYnED6ubRz8CD7ZaMvFfnRfS3ymKYq5GAjG+/mR5SigjVzjV/qF8p3hEssNznEj0HRy
NMiEoctlMhzGYMkjIZvqfx9bPlOjNzcjsxL4p1x+4+rabp+KaIjjw6fm86mKlAdP1jwPyxbec8kN
gjF5CPCLFZ27ax+ngSL6DEczCNDnICPVY3f/e52XLWFxdX2hwWZFo2BkK/QBezmWa9a9UGfks4Kl
jwPa42qLE7XbgdVbM6OR1pRuq3X4u8aKJxle5Br7IMBiGqqKn/T0XMzg5BgMh9x9lNdsWSzC+C+o
jqtcjH38skMULSUOeXD1krUqCgJWrdUf6cqLnsNZBrPPm9AchB6cxFgPGX/Ox94GLH+ewgG2qn1j
KK5gGKkL6r4ngC5rVA7aUHqGXEd78q793vD+mU8dvD49pfbcymasklwSKqSEVhspMn+YbYrDJMJ6
avj0XZGa/aZFWxX2k/ikhcGZZxcr+lvv/2P8t24N4vsa1iWqjvqGvKC9WJjqIzlxdvoWy3RzxUdt
lgOobtX5OAf3i3aq/qfWimTYoOJy6S+ronm8X/EtuZ/XRNCeOeX3UTDlimvztUT8U2kM2yiFNg09
GLIco6aEbz/DIftlL4+j/4dz+gJbNQtuQ3EAh9p5g28+ry6ECXq1PyJcsHitQjOUxJ+b0t4nkRY4
ysjNCs2aQfnfaa52TSX/KRCiupb+9qWi2cdL2b7zBOS7yAELiPfHvFiUEzxquptPJR3Q4aO4UoWU
l+9PlqNGXarxaWIrpB8Zk7B+LGJgedcUtVadKaxeg1i+3QqmLeJl1YqFjsW2L0Q22QQpnGMZLB+O
wAYXBl+L33oLrQOyD+HUyRiKKeAKWHyv/11AkahXj0sP0Y+8dmSym2wzp1p/xMwASRdZmx8heLc7
akAJnlD6wWrY2ovbYg5Eh04Mtf/qz1DRSd0X/pSaZLK/r9ZbUu4o9JitrJ+uYAbJq8R1z6Pv3sWk
Fg2UP/wjWtMv87a8yLoEc249qi0xzZzVCSh6NegB6kvCZCjV3Povx+MFn863N2VA2kWHF7wjdN6W
WXrZ+k9hFMZPEioxE9g8PtpawF1YUK/optAW+hshUejf0dEEQjtzNviCCvAVFDdqGpBvpAPtWhpx
hDfNFomfFOSgVm2EcKUWVpHoasj+GwS+FrqLGd0kqZF0ZuUxC7Oow9QOpop8cOo4gFG9Ooq87MOm
Xc4vJqw5asuWq9cT0A5O9/POsCmGOzZdgotpZ2rZbrfpW6CrRlkc2P5uttwtDzp7nBc6Byv+lbv6
j6MdSIlEXE1r6oxxym9fO0/GFRRjYuqJAtq/LP9N2B5BTVzA4vmreI5cE3jsz5I3G9BdSoJT2mge
DdC2EjexfdcdvW9PO1JuGZ1zczX25/F/FKABWfMrm0ZJ72GTA9lZLGd2LLHQHTG0J0OYWgMZwanl
j/X5QFO2eLIAFkrnTad78x7Qcvi0S83yzMM0whVM3xIarFw28guWQEkWqoT6VG73Ui6bYoCHe7R4
nJnZsXvfAP7L2Cdut5rhf9/y/WOXNe02LSDS+ygxS62k67i1dDLmkSiZkjXq3wfA8KBpezGvCLOm
Qy8fdEoIyeUNqmw62dOmPQZCBKThxLfYPv6IKi3rjn/KASVqlg5AQLXQjvNMxoj3e+bGpRirQygn
fXcuxsSaz/KeOVkbVAdaxkJlw+hA1jS63W1+8Tu4SrX/pJ4Ub+JRmmqpCuHO1Vwx2TDeP3BD3DQj
yf4gDbLSdd76ZknDBxlT4mFqVEbOfI5JIMXNVgezBb+jNEFw/vL7vM3wLyYqCBgotGLNoS6hBLl5
qMnAGMLuZ8rYPqqaaHJYbXUMgPLrZCZoG8i0DQV64IYHsHshmnQtE37YwtBM+0aOzpRe0OWxwdLQ
QydbeZi8TD0oxq4mMuXyIGlL6j1/iu2lHx4Mq5iyLw1KX6FjkKHBUK4aw4wCVygrGB4bAC3uSfo9
8rhsNlpZ+PuXsy64hFuNKV7eyXNNM6JaYU+NjUxgbPfQ4vuPE9x0LvhtiTkbdaw1prR9HDahOkXP
xO/MCL2DaTRj/MQKy4FDt+eiheXT/xKNJfaEM5d3acBS9BtVsVJzJdWztmtrE9aiCe5XUA/bxzuX
aJvG93I6NUDeyn54dyUMM2ad555TK9oNhcHuBweSJlq0pTCCLisKmh05nCAiRosS86ZtZcxLa+X8
25rbAAqJyE5i1q3wYKSS/3gXXAA8u14PkRzlaFpQ23ExQXYuHnpQkuUFogu41gI5+vkMP15yEk09
xv/B7W5l4KQxHomOw3XJCTd4s6re0d9/iajMpd4zKhgwspyVS7FfU83cAvVHJ6U6FBoTPsYAzx1x
mnUcDtFvfSeZTwxKNFxKZmn5kowWf/4w5T1SRZaulQzeX8MPfpKaTerzhryNWzv9SbNQnteGfXx/
eR9V5imISPtD6arJa5D7a56vjTyJd/XXQhoYFgAauS0mbir/VFx7IGsESHYPPWjRT/+9+PwM1YaF
LGtdRlTeoVhOdOAVM7hbqBD/lX4IriAQtEhpf21g0q3tWoEE7r+sEU+7KmdeCkcoit2CD0Btploi
O+pUc7iB8Z6JbL5OmK+YcbC11nPblLcE049YBrdHr7D8WAQ3rUMSSKJRwZji/OUta1nvWSvf5Xla
Jf6fWhAtUVua4NDYu4mYReT3DntDyAjcrkf+ylb4yHQJKQR9vEWj64MXk7m2ZoSjHdbJ9mmkYoAp
9SxAK9DmnXoQVP8sxZeLF/CQBSUfM13PpcmUoYQ0xD2vobmoPToN8VPCnR2gn9zHty/2QWahekUW
MKkRysSL++Tx8HnZNG6TCKjZAYlf0iDcus9JuTQgyPZfwy5Y7qXKUe/TPmy8ArcU4RFo24hDbBD7
z0Ek+RZCwgcV3EPyE/w5zv8540gmmQKl3XodkM5PHZxWJDaQmRhNkKU5gpspY/cTwbzy0lmZcwiq
RxE+UhTfNCMRJLC+dBjuTd/Onvt7Dp6spmXL02RWurVvLTz38ltDrCENj+wZ262QvRh7ADH+L22n
8LxtxhTDY3QRci2UP4om3AT5HKsEoFIXR7pstuKkbeyQWaLBYCKFReykicfj/pyFZ28+ZZtrpLi4
OBMmhvdzzIG4KgN0nKWSJZsl2mqOE6qq4artHcaE+bQwMZ/54H4dqavOzEjSX0NHp4Bnx9dbzTiM
g1HTEmfTFKbbpTITXlx3Uqk8ZoZ64kL6H5aEPBLV3Tw8lWncAgFrIgPlOOdyREDj01lPEj3dA5mk
PjXkhbVY8GcP1CJmf1e/u7RBYLMjHkTFXHb+BMp7BOl03unVxUwgECi6vy7XZr86Ckb3EwlRJppF
DKbS7HixsYBxODOMcQmQ7iiIiqAatrllVSxkYqrl0QAF5oNEysROcKunlWenpPKs62qlseaOqYTR
ZmkIkjhnBAioE3DxfOKB4SxBF8vH53Zlev752Ji/OH3bXbG43rdX3iuOulnJqlZ3cZYc7hLpvKyv
yPi/qHcKGX8PbTLTcCkLnjIqKWWMAxZ/mvF1D2pQbS6vhc5wOSp5j08esb1kNL9ieOxNTnILrSUz
xw0EPZz+N9Ifsf6zFXhVRPhsQOAWB+KN1TZ0Ubskfegqrd0pbl+fihiwjY2o+4FKNwcRTtvPY75c
WADPdDELadMsM3VR+R4ejrmeeVS2f4T9YPcU99wFBvAPD1phybJu9v7cA2mEHDm/j7qndCmjie+u
4dHRVOl40SK7xmCaBXYySOkuAaDfeA11KgBj2ZZBaB3IXmOiSx0uldrteRoowQHzfzOcNRBdaAan
ctuGI37zl5gKn2pB0DwYrSaoSU+GsvS5KNCDUyG+XbFFxH3JbR32uwPv8x+2KwQMsR+diWoPfuac
TvQLBvI/i1lx48uypeZ7AFHsxG0ty1Aniye5qxrWVHvNffAHAhC1dl1LG+Kgt92NdNzdci4Ptj5t
3hxtjwv1+PGOIqnKBwMYiTYhTT4MVkQnAuPpOvKQsH5gXGQAqUL5h+kYBICF6pMyQ+sSN6luV85g
TTu8Y4er4FgBTOvhzb036emCeF4Po+ykFRUpdPhXPAYhsH4FMD5/QH5Qr+CF+m/vUtI/jXDe44Rh
FRTryOEDHENovmX23+nrs2YLeAGIiKMecxRBrufGBR9uB0WBuIapvzgDTuCByPRSXquUtgyU81px
KrpcMAzsKoa+82HDcr4dxLzTCiLbwAtxr3y+f1rqUOX6Sug1s1vwYG2rJXrVn50STl14kvoQLoKv
nDBgNAO+zLL1Xyzu7NUh6vqda8z7CNt1hqboyzdE7nDN4r4nKDZgUPEzHs4HLsThaU7KK766nMZ/
1Oe/6fEid1eRNQ/Iw+xWPOfjFsGOvwlsKEoIOgjVVdtURJNxoMgtTLkJUAOFQdXTy8nCvxHg6C9M
63LmU4NGi05RRFie/Koc6yJVLqhFHiLz7WWD18VKMEUzAFwX723JI9f5gNyEZnVjr2jaHr5utqRc
T8Bq1+WuamGwkbihqzlFQiHgSDctos0Tdh3/D+vbIrlLkLgftSJVVoVM5QQL6jHqheLXLQ8eioq3
VJzv6KN7YObnADtS9VpeswsM4yrgb2Eitj7Vg49hxyBS6ISbpVjUaSsm2/ufzUytzgrRCdD3C4Ac
MeXxKa6HxY9eEhUtgJJuiXPNo2oxBucmQBVk5uCBNv4vQB6wgAWJaaFTcJT4YIDX9I68lzFtTVB+
heBtu52YT32deqzt97zlKFojUMT15XPmGQYSQ9bbP1hxfWoyCM8IF+txXvw7DgcF/1dVxaGRj2pO
h2RgAVB6qJejU/nS7INI8n65uN/YMhHgAeO89XyobY7mCbzsfrT6g3dVkD7Y2mHn4yUVlxUbzVSq
Buld/Rdm491u48uMj+lUl+KVDZRMnoI0alEHAxzG5pS6A/u9PFnk1n+d9+xaNz5T/vPmI3e5QL9E
ciee7OrleXqyvwNmcT2hWWO2Dk5yO+XYYdk7n7/qzpQsGK7/Dk97Mnr2qOKf4tDDTN6TS8W7EKac
CjQxq4SzyB85pPKRKwelau9u3zXTOVWkr6iaJ39e13lQtLB7L+5O3fdEbJ0Sv5nDSOyEyl9M6ifq
0ziTZRBXZAwgdSlMHquH065bmpMpPVo3YGePxS6bWDgNzW2eEeNtpSAcpSlsOauAD+E/wysG1/tQ
S2Na7L3aiCrVwQlJXjKB5jQ2Zc8kX2kLPPnrB/eAuCd6GHpm/UjP+RHrarbmKLXpsqGpNmskg6wj
MkVi0o2IGL5FHku1/4R5xKWkNxrloQVE5+YyBsu+gNKqF6NFFdTAvdI/aX36buW1T8ZjYCoANvbk
MKH8Oe+49tCARm5P1cFTXZe3rwP1/hs62sM0DV7+sMnk4HizrB90g9jqNntiF7KQ3JAbVlVgn4YE
ZOuupg9fBTjdTQRpGBMKw0AwKin8+kf9Xjz10bd4dEp8/nRwZvQHrNZxyTntnHiQVnMZl1dtj5eS
7Hzekf3gVroOcMtFK6/GHGsekKq9RAXtmDEIfEWWbt7EuT4cguJmcxWZLf7o+s7MSlblDYHOZ3Og
KV4UrBKdFz/PZuW8jxtPaXYd7RGAtHDC1L7WPReTy+SqsEpb67PgoOZJOQFrYe+eQwwVqh/RD2vc
w1/+oztrU9gK3eDRC6C5nKqpWo8zq2zFIjhV21549S2LPdf7A7fz5w/nZriwCHl4b+hZhxxCc5k3
USphF8Or1yOWPxntAKBL5Y/vNuXX0nwzb7a9ziHeXc0t2w/JEYSkevHk0rC1NLAFo0SOjoLpNS84
jGNOUmtNtE8eSsMXPRXQb8hjwkqd8L5Cx6if09H6k3TEvIIkfvnPCPgSmAxQP+YuyuCCCBpS8r4G
6CiaiJpvI8xKkQ1bmP+9O1/7SQBPDJoXPCm8H5RXvnd90dcMB5xzZO6YwN6V0HMqT9TfBUa+pFOn
LxD0qjklbk+5mEztWSCoL1MWqmWuWhO1zy45avGzO2xmz0y8uyObIcbi9rrkp2J7KExZWAXXQF8M
Es/VHMsp+k161yoZWsSeDcd5nnDZAhxu9O5lQO28t3wxOwhrFu9q1GRbTRfSzLun0piTOu7QEAh9
XKaL741cza5ZXIS0/39ivpNWjnBb+1PJP/gx4pm6/GdhaIqKqrvXcTXpIjT592N617AR7D6cpaPz
sIQjx4mMOKd89WUXTrb0n6DqFM8GLGXJ7+GE+u5s+Xo/P6tifGvTFJLcjZxdT5W5B3belHSVmAs+
oY5XT9CGMNJosuYx+MnWqZIJ1J9Wks8x5o0eGU06CRYWM44J3CKAyc0EIUNnDKiUZP9ZBVarOB7I
auHHMXJbv3ljfXPTLC/mqcA40mjqzttpjrDRD9dn72jpoQ4kyGoegV6HYEUEdktbf1hUMIjFA8Sq
lWokOAUegcrQZQmS++/e691EMW24DskswotsXmBAJWnqRqGhfDjutSNZkYxoqdLHjOve2G2twHIy
HNv+Kfh8mdntTuObkq/LSQDamMiZ6CSK7Zsup/jaG6kMNiuDs3Kytmx/kZ8byjvyRSGFnUDJkJr9
JJJSoUbACYSi/dXF8Dv/gj4DH45mUNse25WSeUI91Lcjyt1xJTuAgi7e+anHS8DgAkfaNcoovWJy
8P0I3G5fjOtLDC9lWLvWxouOhGig1WafJp3QR7b3lZYO4syCwv5VIcaZokJf/RChrNa9CYn0OWty
dGNjmVPycxZ5Vs0PRbWyLY7eW14rdUBbsR9KV5JZ8lYuXRVsIcc6rrHjzkOzG7adINPViBiOw+V8
bZGkRXwMrmsBXwBJNihQA8JPeKNCX8Fn+q0RKT/Rhh5krNEQZ7Mg/dEJqZ9KfiNQaoCMH+cM4pVF
pwh/PvJBPR205LOgUW8Wsw09XT+QbXW8A5C0N1G+gw2SIXktyWyw4rrIiVt2VhFa+nfZbYw0uLSU
xYW0WytBxec0O4618zFYUwnSyoL9FaVuFsArHTU6OrFTGEnpfaRzLWSbu0mJMMHxEPKdM+4+T0di
6kzitQNEnnnuwNIsswtITBh8uuzpQMMKt2MzrElo1sdw1wO+0Qcye4kBhSzDqKI8EVAunLPfZHPx
lOtk2CrKVpQFx+fwKWW3tPoRztytK9FRLVUQ2mfYPSHyxXauXoIC/54bihckURGnn0ESmEVsH97I
RCQvyX0ynlh4Sh3sulIRv8jGneQ1x3785oQ++2dUIAhb5u3gK1cZ+RQSv/ZiDd/3IUm72RMoUWf7
o6BMuDoBCfR7ZUowimOUe5mvB38AuiZ4HD/2R9bDpQdlgnH/Y5VINQeIsZTnv+QmYBSbstplEhwZ
iEOxSBOVfQaRGoZhdjdgwLrkLZBmO3JD7fLSS0GSMuPh6cwdu5eQgx5IwAKt1PtGJYWcCkwYqCDV
YDLa5bDLbm3Egv8HDBSck53p+CADaMuzOxrlZccKDnDqAeWcXWiz1BTjwT5FfND7vGDHvSbVv+8G
n2m6TkNGCWlK4Ise/+CHDPK8jAt6iUdnTcGcCdeeLw0vVdTLUOCCb+jw9tXSjWAm7KGsUWM3e/ma
5Crso1bi5wQIpizSmz73vulmQ5qhCR4xnbK9NIn6kUggmla5m24uftzREHw/waP7ufVdxFrwgTg+
blklBKqkS2cJxXzLADhb712CP59vEJ+GQXPV/I5HHLrzL+8pc3aFW0ywADoy6usLs/YbuKnmV5gY
jLV8ByWtuu8E1nHcIOHREZxYzY9nLJEofssMLPoCujHAoo74Ojt0MVEPJIg8Z6oo4uS9p+KTOBrm
ATuLnCWAZaSV0pqJx9TCb9piSr7pZq7SQ2INhM6DyQpZ3iwFEJvdCdRd3hhwgKSzy+Q6FlzqDGsC
EM1DZRC6nbtgXNUdg6InotkoQ/SIY5s4mWqB/sUIBb1A66LUJ9LuvABIKcJZABkDh4lUjRwKut0d
V0hejk4BDeARYiD9qrcc3NWUQ8dSWEITtUsQfzIwCE68oPll6RISFYk8O3DCuGoEImsChml+8xey
OkFxwjqIdSXeZJrIC7yDoz9A0OBoEHP4XJIAXnoxjL1PnNMh7ftttBgV9486pg34MjmObXoma4W3
SoFjbLYqRyh3gPUyS8tyJvp5ovBzcZn0ptzxG4RLdh/mS5Fy9cWHz905lUgh2YY3c8llu2hkrf9E
x3PHA7wOgxt8gfU+9TdFUmBDsb2KGol/CHErjvbJshc8M2z4B8bYfWcwp1+lF3b2hxb2xRtEeJ99
v61+YRKyq8siSuljbJF921zqMl+dxxcbEfYqy5IXmH5lU5Vk/n8ERJYN4/WT+njD+wYxwqJnermN
Mj6l3Iox3Apfi5enOwCfV02AL0QiwZbXrNPcpjyqsriGtVr88GqqJaYSWwZItyJkM+Jxiuu4hXGA
0a0HgzdLGOq8td/zrEZ1Qb276blNA4SrHq1xPqCq5hQHj+WecPD/F4ma+p/e8lEEfEeWxSHmhCDF
71EaKKXK1L26MSo7CsT9JmzWIjNT431mIXf2YMNyJ4INgmhcxkAsHb0odCP9qQjMkLSDLDMnqaaQ
6h6Yt//YjftLZoqI/iVRVCuKvPTuJ/OQ3Sd93QfEpsaNao6bFD2WVvq6L3D6MTfXE0AdEj3GMc41
7C/E2vhPf8CTWAsX/DKAhcG8kLfYJ0JQ483TKsbUFNGlxBoR+pxd6QX2IABsbc2J6dMpK+CGiGMg
++Ji/TtdTjthuNyDE2GO1AUoVWf/0okIM4d3wuSIajxhuWRSTtmuyoZAnswy17SJQ2SeyAcLxOIB
GWcY1oa5nJeZMJbhyqe87rO7vWbGqpuw4H9DDUUJlvB0pOldEpJlIeBI4sJsE1RykgOXXScTZt8d
NmkGPs4VjjaeFGyYvy+qHt1VqN4e3W2wMSzHT9K5xG0U8tSPj12EhyIeIlk4Uic8283kqckLkfL5
Rg0zUedsR8lQVvo6I85sUI2+CH34KPS0Ll9lIrBWbayCXwIlSYTQ1Wk0juX3Ukh6MonJmi1EghI1
EnTfNCSNYgruUi700sZPULN6ZVIUiyJ8DP98/UWPb89JNv442z7AYlIdTKdwlOtlJ/itGMKpwcj9
evkCJ+NeMjpTJ92bg8I3sj0wXeOoygc5nDS4gvHzQK6EAhPZFhFNhyXoKQ/pi8dhonalptDzl9if
fO6X9Bco7qF63D3c42PBL8+6w54w4momwyJN3ykn8thuWZuTkZpydDNe1rF3y7USYbundjdRTtgT
ma+RRRJpk518UEu1l37jRmClYOw+o/bJso9IUOPZn0GlwFTkBL/pqkB5XTV30FcmVwVkXJ/VnhXL
QadpJR35VcQAAkVr7vMOsWqSh9Ra+HfrohT4xvEt2K0rRleZeTwjx81Qcj1/nLCZfaGwRz3T0Bkm
z4ai7Fcdj4S4YpS1oF01kIDZwQIqfB/bcJJYmECuNuxGOJxtXWUWTuIsKtsMwDljOQL4BxMt36QA
d66phBFf5LiMknrnlf+dLrijw7fJ8v2V2Xc7dt9WTnQ2Mi2LcvQ6DZ0cAotAGBFZbYT1Ih0K43DM
iGpuL1VMEaGBzMZ6MiILJ/pggOPMA+kKzsO/Ti+RCtI3aLq6sMUjjpTnq8Nb+f7iAW/MSGriE5rf
mQLFrUATxGsIGHqW6V41j6hFxyIoR5oxwLYysRS3h1TnkAv+j+Ld1W/h/QgaMqXv7ymVJG7J/rGF
P/RaVQ5ufuiag7m6++KQYPLwIbg4djAyM65m8S1aSd8+/1CQIkCvxMqKkz1w1QvAycLuh4l3ebQj
7SagUAh3zBQCsj8Iidk1phTS+zjhdshYIGxqoLyVk+PIrNeyuKTXMZIfD2bq/c0VBbFEoIEKZg/u
CABpOJkkQcItfy3+BZ06wYjiE59G75b1GUOm9LtMOy4hpEipk7wf84PgVisCN4ky+EvtDg/0/WDb
6AqhjaFHRmDaRQLFjE6EfrvSmuB7FxwaSCp7eSbDvKVZZgvX4cKhT+TiJGbAKmO4ajdsVP8gfO82
EfpqCescjfjayjkGcaRemSKuNbT7bjeg8SdzLM4N2K8VdO3mc/Psfp9l8be8mWzs2VOj94G7cq/Z
dljmKsQSo1Y3SiMkqOzGR1+A1oRCqxOgGBREM0B3dEIbhfuk5f+xn12cXBmAL3g+VyrRQAATGQax
0xkcgmd2FaLc1vZA7QlmUXAGpd0NNa5YkDbBS24L+7fJubtxn0hpfiSbGF15qh9jSE7r/0SoT1zV
yd3oDbaTLuJVEuj0jCX1JDWUc4TRUyzKaKwQLFPo4QefGEaGPzH/RVRSq4Z/nJkLoStOS81/Y0dJ
k5fWJYFKrVFWdWMw2isT7DEsv50grq0EZDVgCCkN6E8tvL+yzZt07Z6mH+TWpOmkgL6K5GKdD2ya
5QQx0W/7sWkJ0v8vmlI+3rMNicyVTQCnSyvNTCXN91r1R8fLBGlraeIfn3Gm32saISl6btGX9/bi
DUBLeNu5yPfc8MN9pTZ8G/XpJQ5s75a+cqV53bOQstRpFo1Fho31lY9JaMN/ClcdHQZTVH/oFj8W
h79kE3C1dfJo4gFGmIYGAN9ThqTYVvsNqJ5aYbI5mpQ4lXmnVx8XqxVc8bg9uMdRza4DZ3wn7P6h
mbs0TjouWg4WT2Q101/eYp7rMsEx3qvlno+3xKflUF8Ssj9zpxSpX2ZJvxc9HvcrKdMx5b29r+Ma
D6tqxKMy/s89Pjzgtz2Cvtl7nOfQnVNelxPyg90jQOc+rulfuNiS6s7ArIR6+Cqn/2v8euBCiv9x
csfbekJwj/J7ZhiiuN+zpXUJLwLnK5zUDZgDHZ/PhpeHK7U2sW+NV912PswwMp25Sc1LXf8ae/4W
I1napqEdkRFEazkPOXIYOLDcA0Bugal+j/N4umyPRYsYd2iyyNt8DzzSIcOuDqdNj2VXQ+nnNqPS
yByNMyyI4ZB4S3mMJKI6ejk6iZoDvBCvLOcdYV6dRtktAbzBBJtsipxcDXTD4DvLCTKmJXk7q/Ue
C58erleOUziCRiyrxZT5k6LOLbeNB2YbQYFFouNVgVIRUnwUYit3OQcEWoNUFEP6BOBw3ivtzyqc
L2JpQxx6IlPgMujdpcVdJSYzeBvEWS5PHJj3aTLEGNbxEl7sv76OPAFWXm3L0zlmj909pL93BiGx
r0w6YZXenCUMiUwGKE6CtMdFpeh3+YRrYWbPcBBO5+iBWkW2poGE+BUt14RhUamStWP+F6rCAmQB
RwnVeolJGsTy1boUdmi6iYnATGEgp2K+KbUn4pagxsuAuH/0ZNK84TcL6X69zldgMfb2xm/breHP
4b7qI7wiu+xZBCM8DIyJYnjeDF1GfTn2oSF7PUO+NMq2vz4t5WXLsChsd+JetRP4pyGPBNrg/MIo
IEGZEw7alnkEcrtsnGapzV6PXCePWmCzha745OAHnoA+v09RDWvSxsrJODtKgKdJgsmOk9mGqMUe
ME2FR0eH9WNLsnRGZ6izyja99wUxqb0H7VHf3/LAx8SOTR234TO+V+rBVZ/r4itT6czljINLoSmf
2lpXp0+dCd0dXSkdyaE6h/O4aTt8v9CMQZt8Hw1fC3+k+52HbHqaIP2lnatW9DkIMDS6UEGPIYfb
MiNhZimjsugpyxV2wLDQ6vuBrXN0XwmItHkVO1vemsOrCUt3WjxpQbMNrl4Gnmt1n2HWlBrBVGp2
A1OGA6jeF9h4QEEKr7/fmn7ypiluReX4eCkXRb90aNT4hsJVwj4X2PKXf3D9ZPzaasYbY04n/IwT
P3d3Sa8bGGOygSC4m0KRGrAudCNgyDoJDYkJ9n+h4lJFN4PJgLe3KAGMdvvYsBTO9p6SVht8ZuST
/oa6N0M5ekqitEzO/oZs1YjGlUZ0cQWtH/CsdFDRGr3+IB+UEg4IytLqS4JnQQNv4Mz4pSdA3VXY
6I2+gd3f89EuIUdKkJR5c4psQZSDQuZDDqXhLOQzUUxKNsDNsloAMuxFf4w49qa1yEfFPR8CaOg/
lEk2RISCa4QfmFIURZJM5a0k1QYV1KHQZxnx27Hn0MJzEdSmlsrecO2LyNGegdnfcwED5CNtOhbV
aukFOgXJNF5lSGmKtWY9OXR0yH9zkvhMW9mP+E9CIIqR4x6zGx0Y6Dv8J1JLAZAdlICz/2RyjWKO
pBinDT4knJxzMIqxo908YrNAGDeQwho9YUb3Fgob+0CttcEJhAZ1FzVpA+jB/YARG01cRWTJj+C8
mEyCzfimPdcFVvH1AxInZiomNAnJbM9DyT/pTs6eJuUDlGQQT+AaGKF0gT6DTJG008fsblXvi0H7
ppLdtYXxtzfP+oN/ylQfQ/p50Jqvzucz5ChEz38qgtWHeqCd6XNVTBITNIBwkjHS7uJDI4nrSzJ6
YuHYwdKrP4KEUlNvaYEDKv/EbxYz7TuWWpeUzhLkcObjsGG9/tExe0G1O4Q82DLdxhiaMcy1i4zI
IT0wvbBQj/4As595Pr+1F0WsqRV16LozSffqmI2Vv6ayRmALAAYdcWG66Uueu24k1gQyBNlHfIJN
LxOrrPEGWKb8I3Vaf3c2uaIeTWBJy2H1sBncCK8ondDu1y9i+swcTm+CXPcpdmNUZwum0LdRhFfK
azJDPeKHo/0TUx57gm4NEgl2IKplkayr9dYu/757CjWZ4wPGffAWCaep4zd/yN1hZu3RwoqszHb1
LSBNQlKu/qhAIzrgXsQn4c2cf8haR1TMcMh/y0vrJ2D9qmoe2EtLXBxt9XUSAMxdgLsStXTuwpIx
DF6eZiD0Ql/gMGYHnhLmB92R3XDEisTvXPA93LcUAvj38OoPTAO3OK+ZiytPNPZ2KeKOEs6coIub
9zoCufIcb1nUjPWqqIDEyDMtSmJ9FzsEN8gL7FQbLOiTOJOURHp738AHWCQnyZT1KHjaev678wwC
S7q5MTVxSqd6JqQWYeyuOgxxkxJWa8O0SghSXih18WC2WDJvXB4srYl6+yFCm0jkCsYUeuHDhy9r
MgFvNN0iCEx9ndBDf007oxhlO6pRs1q24ZCk6YHxQNBRVNycKDH7DgJ/rMeGd0+hBQZ5i15M7znm
W7GDKV/8bTbVLXPhGgzyC2KFT3ScIgKyoO+ypJfl7me5xmsI2/XP1vg4cE2vmoArRaP6iWTYyBWY
LQuluzzbZmgpV5yl8//L6Dm35RL5tURUwZckFuJ/xUbCClR1lQTxPCILYtlNavn0TvHobMMGTQKy
tso8eWFLRWb47q7J1YSHyj5NF0p52buvB7J0Hykp98pWyXGjUaSl5buPDbkB3x6kB38lcLHG0N3v
acsIFpIU1kZu3bhgw2b+r0Cevi7+D+8PmT76nk2qfY46TWohsmCvnDaQGq6PYD0DkLqyhRHHCXU1
GifLeuibIjU1NHw/ipTrT7W7Mif4Api4vDevU2b4+CcaaFA2P5arzXnWMnfgfPOfwfFQTJWBpZmR
A4iy20DTCs3Nwy6/l2Gonvm5JnNQ5klnByhzh7Rm6R/DDGnmFFkDuQaht7Z+qYFMVi1dOYvuT+3t
94KSIpBIoupT8JMvIw70T8ChAT8pF3Zgj4JHq4GSjsKyS3G5taEZFj51oXXHnA8UeGhjEboi1qDf
ToxW7zKelYygHdPon88Shk3dgyKq/24DE/pZ8ejNtlvcEsnpI22nTQZHPImvHsPvgopn2TiCWdsl
ACQSt2AU+GmmlZUK+df5B/+RfgGQM0lECbS58O4j3/kMJIr8WZJSKPgb8xUP/V5hNS+lN2E5wj03
gugI35GM8yXa0NQpMgkCnT7rGIhDB13iVkkBEj0OdW8b1Wt2RXGHw3wQNLsJHu1EsTJxF2mwA3e7
aR4iaSyFc1ssXBP4pEfAZgc7Awp31FbC5xXa0TELtI/eqEWFNDx8b8ncQa4R+UcFZnes7QKmVH1Z
MYZQ1j7HmHD29gj55j0QztgW03+zSarehsSq6krYRz3HloSRvRUSr9IS46MD+eBF/ifxh26/efhu
kf2AmK3YAXP7dQRmFU9ubOZOX8pgZ4ak0C4lj4QIT/vZoq57qCsCRqkUGyp08S2rtJiM8PxjQjgy
gHm/I788fP6HroqmdmaRMmwofOT/CpPoC1z0l5nERDsjBgpIn9OSz2gPFbq1dQcg4xHFKJGai8Vm
fR20QH+oBayx7v2J91ANxciZTI+MMG8C7bzPDTZMXSauJIvb82WKQRVT3VMs4v/qz2gja/8K6ANa
6eZPV30Tab2mrr5Ze8/yJLN+wgGnA/JryNuYWh7QySkBciNJmV9QlbM/89XMomKLSZS20R7XnfA1
ygYubcXybaAJxU1KtJyvd2NqZoNzVnof66GjQ7mb+nxfb4+Du0QtgRZ3S0wFGXw1HDI05g0H6XiH
Pa8UvGL7ohByHWxz7aVxwzplPy24a2udyJ4kHTNf2ZJQUu9300KMyF9t+X3Rd9DBfFQaeZLFAkbn
L1SmDx500QGXkwDtiRsqX/cujJhMsONpFvDYQAJlsT7GRQ47lniy2wP7NXdjq3C/WDt8iSii+eJP
1b7Cw6n2uJOEA38uzOgj+eZUhGtK0XfT/LLOjFbfe8+dfvt1W2zyjn9kI6V0G2cgQvhAc0Bz/Je3
QHUZ5gWRS2ecSZSHmYG7XOoQXrzwI8ZGxOWBuAsnXfjxtOI9hDQYmXCaD2Y6kHFXZL8rv2pUihkw
ey0EDvL1W8m4wMFkOE6noKM166C5gkgVDgtMmS4lUAJJTHWGSckPW2ZdLlBpu9CbOMVxP3s18fvS
X6lcH2n3QufjKIBr0jo2Kl5leHvRCKM2Sgr6QzcoXbtUbHjFneeIh00lXqsl7xi9fmSOSdUggKFZ
nXJbhE36ITixL95g1Ed9hyQQ5ne5rWewEHv3HlHduYzbAoOIwajzVM5dLAxhOwC77KV3igrciOUn
mDsVuP6gBP50XyibSZ605RWX92tMdSiqKMM5VLEIixxJGGRYzEQjz1WZSOVW/l+z8Nsd/uVt3JMa
hrDrxJS9QrlFfqtPLAnLFS5NMyHh6eXNiaHAu0Hh70JflKFuIUw7KA6+SEdUXTrhbjT+jUzABIyL
R5PrsSdvGGkXhORTMOU51qsjteVARMSxqUgDtQejPDfThHWe1mEaAbOzGLSoxZ3EJK/nb0GTC9JL
ZK9Uxobd+qTzdlI5X56TP6cGYKanYMgLhiR8kKmjCXETUvOS7r+MxxNje3wzLWyR/abb4ymWdyE7
K5ZvveeTR3PyS6B6jZJq7rcOXxc1ZliyvydcfIpenSG14OnMzwduYkSGjVJQk42cSYm9rbQ6myYH
dcmoEjqzWMzSwBJnMMkGIDEFgDpxN++inTzyyv/db6f4/Wx/Rkk673zmlwCVTV2qHyAYWSTAA8h5
po5j6GliyzoakvPbQoKdTWMPfUxVNJl4wTXRARiGF2zJeotXETl9dllqgYHvKqsvn9I5ebJGU5oY
eSyJhPbgrzhX1hf1/hG3I+HxPT9V7TI/q9Sq272zuuJE5nv57QD8YfLnOShbipIwOmSnLkvNHVrY
MbJKLtpngEpwWowxz1U5R8GjEyhzvyQ3FgMhO0CLFMblhBhvAoMi5OjHoH8jyDCl6pLNuVvQ6Alh
zEkwdniajMwqVDkfwGqEfyidoHXplEcWfxC62XLTJwY1mlOwyU8XjAIN/nS6gf15CMYWWHQeAxHs
9fJta0a/hZ3s6ENVq7V8MApth54d7GvatLzmfOu2p9+ZkOwU6uERPs5cFU3wbN50aiX9SifjmHUb
3kB8qIsti24wikia/lH44JzOK6jVF/6zN8v3+YU+dGclgY7YtMUpY/ns6ximEqmg+FHyILs7Ww1w
6jNEuf5PMoA7aINAWVli7BG5EzFtCBnsEGYqKuoU+bjMtQJhgW67k/Ccf5jKltVmcTGo/XwnZQqF
01YV99hF/Tw4s4HQ1Yufw1TVvumC8DMOMYpVDhCT8ldISy7gSzA1ke9qLKPiAD78X3OM4E5wDrX5
dAU9mtKHd3dAXsjrrxn1xxEK+r2/fGgR9FMpHCggd9HnX19+1RkdN2Pt0mlzOrWo22RmSptilsDN
UUhHfJB9hTU+9ibaepYhrx0bEqCMvg8BnklhgOOrUC24R6DgiVAIvLcYqm6cIwW43rACAH+F+R1p
SsazTw+Zvx2pplldLxcYkbFhpwmY5jeQUyaKtv5ye1kRZqyZzJKo7RsepCY/Repwn7hqRgpqenIy
c2qrMFRZwo4rRO3j99N9wN4pe7rsKGqOC4agg1IDccjGTLcdRjfXmPTgmay2XMsfaBRWp35QVcpH
OziA3kxLHztJQpZ0PB52uuih/iV9Gh30IuE6N1ZwodiVwbagQdQwaHc7GVF1StrjlVVKDFmkB6NI
9lVt+JOytVJ680RzURxAEqf9cyQrsLLG+3X3Amr7vt65Te0VtB/q0fAAcWRrcf0rXae4RJxYtx+h
Hqmr1PWoT0vYNU5kvRibHijq0xJsRmGxBHHxqscq+gW1fj3Vw+aAZ2SXShmiUWQDP8kcYQB8KbBO
j42XlsqFAbVqD+F1lULjuhy/kHgF070bgDAHuXSpNVt9F+ueeJawZdt1efOOIhz2/Z+xtMGeJJ7q
C+y9c01vhPgK3eFpMdksgwmThPYgGvgwOXxi+Vi/oBAbpZBsjUKma7RSwpedKzvqeSdV4ncH0WqI
iPqSdCim2O3W/Dh0yflJ0QXm7bx5A0VFLn+y/4JA4j5nVdwISovT7Ho90noCBSEjknaJp5yFEXb3
QXcUjUqHU0RxKZo2LhCPtng0K33w6At3xJA2Dx3dcYh+3BgmmJ5CtZgbH1i46HRmIIVPb01SEPLa
BHnP3iWvD4uEtxpT8CQL8AE4SX9yy2Slhk2OpsY+sL3khGeEgpz32PNyDyVnp2g4wj1d43KH1twT
60hcFXc5Up1FFkPzh/egskCqYB1NuqczFbsy+d9m1vzUYDeyFtiWtGl5a3YEMBG/JuM6UYk4pLww
Gg8PniPeQJqkKn2grr+ScJ1LNbfYiy8Djr5skOfUTHcGeCkkHKwSn1Ylb+jptIHD5jdQFyxTa2FT
QGrkBKuVYWo+OcJSYJ7TLbQylI82M5lyO82WjRYxV/5Rw4zHxdQrRxxeUNKIn9jsUKnVlJzSeuIC
4wL930aaY10dTEFZkIi+GezLnmnwAXQPtWcD1e3jMpsekk6ExbWpyCL/ZhMmr97A+jS9AFXWaX+7
TZ7Jm+kGasSpyzE8exA34eg8iqU/kJq8yM2tHHEt0Uu5NVTmYziZQHiYgAtBGHzaSop8/9myio3h
dVp/EzbNhg6jaElxVItrTeWr1MyAEfVAmDdBT1xziI5xeexu5yCoV6wQChe9iixNPiR6teShAjAr
+FryXFJgYtQh0WxHuOODV2NgLP5CD47c/Ig5cxbqgZjNJdPZmsEn5qrZK/QYMSgRpLuo0QRVfnr7
8+2Zkbn7phwDLHJ+gUO2uM4JkYqMrVCUOhEibt3QZGCfKl8yTRpF3Ai7MoNzoVTtOMC6Mb2iq3ID
MfLDBmuzfxIibn8sXys7+lEr6Hs8YwONGbAOIKvVRk4sJvtzKXU+s1Z5gBV+uNQoRhzv74NNJgia
ngvqOY06UkIYUE6qF7hoSKQy0zJg5uz2noZuoxcbBQzUkOjsBmBM1KJ2v2EhL1Fzzr5uOiAEnzrz
YIg71SM8ncOgdP4XCvAetKKqtsGz00NT7Dzvx1PRRQpAf15ZrSJJIux1yi6e77zkMunjiejeilrP
PvR/dDkkCyRQD9+zddSt2j5LzMOoS1cejbiE2kgXQKh/H24+1eam29MZ270WDaMnrYkA9I7qM4gb
Jd8FE16KAUesy7iosUpPxO1IIqY41RDzikbTRY2saZ9+cu+x6yvzbFM80zDvocwnpVCLoWKwv3Ui
s9rY3fS4DugSZfVQl6N3jGZ0Y9s4OJGM3sbcTqQWsXD3D2Ljt/mcOvBSDEzMKE+SXUF1T0Zk4FzH
xRZq8UR8bD6zVBbPIT2MzpczCHhamY97uLP8NbKanPklZ1csk8EPNPHQaRGfxOq4H2ZxSNlDJfPG
qFyytypvLNOKHsqpPaJKZRUsPNsTAVaC4gma3nt/nKnwkTxPtV/EBCPJ1HswKTJW3zDBC3Ajn/xt
GP9kAe13MpZIeRYYGz9FXuukynmgr7URl0n+H0JweciaOnHJP2gpl7F07cFy3ZWPSTjixqqW1tOC
ALi2vFddqjAtz1VsTammaVqwSm8XdDv20nnYQuunSd64vqTSx/07y5Jp3ssCZuhytpfuZpkxkc94
AahoBol5a+2Hszh/d5CANSwKu/tj+mBYatBoyAsgCE+q03qgAlAUGTwz8Qy9A8Pz1LbJAiJ8kG5B
GYVNHwfhVY/G+80zGSpDCUMacNfRyu1L/KT4mrrVPAVFGY23oqkbdZ0bUAPVVwickaSk/SkpqOwP
CQv722IkA1GlrFDsPsgr8HvgGic5fqzfsPq4Q4GwI8ZWaKImliwQCw/0uch96Jx7vZs+JwrhA3CI
Qq/ZEYjk/sjrkr97+U+/kNzdm9K/HpAShUVzDSzOgIudyez3Aavhe9KhoeLYN749qSplUIzpIqr4
OkJlq/GycbmMwTqhkmMg4cVNYgIyM+4wDymor0syC23uOS98MdkxIDC3SFY9wGMftxgf720BZl+4
Mz2AZmKCrhevzuIeJCUXPqPoELvuTyyhsmua5uAbh5Nx8ul288ByBWZh4in8ToX49Ar+N3NeqVKd
p4H/5QqlLpbl6V5K1+XjexR2xbnJ10P1hHv1pFCAl3F0b++Dc9eXin69PUqF5EEDHRWQf85vO0i8
eiVo8ge/IlI1kWolCE9wO+BM7Jv5cMr7Osc+KlMpFTiTkXB1oQUwEbLIXgGjzJdztl+UzmpbYzq4
8/W93E+Xf9zwPH5th8Mrjh+M7pJZblLrHDmzvGPx+gJUagNFCk1I6fxhZAVqusGSRXqb5vZ0Mpqb
1tSqAJkF6PFws5RGGykdHgXpetHntNqPbHIXiTaYek8ydz+j3dw2ybpPhdDUeo7G5vb93crBDRRX
Av9ape1dgwOXOURnoUHRLzEjmktdTfTLw4Fm9+OKhmg/u2cIZpfUOvhRhvrz0+JRZEGuPH91KUxw
bNeHslJaQ/fOrKI7WEF3+pIKaJ0Q2tbaErsi2X8moEXAf7afczWVGiwGgEtIikHsyTPQJcP66wEg
hg+uPIR7l3kfrRkkpkWtNfNxKmOPLvMEBv6UkGTZnm7ceehh4Rdew9ISCZDohYsMDfaUeUAugTgH
gy/Zbu8F8yj0uhxYELvWLNoYksm562eoP9dP/aySBOkdv88G2KpQUMktOyBV2nIAEV+ZTSIYjx6l
ngk8alK/GM4TPaL55sdmC0uN0b8Ce+UIRXql/+nnAduklIEyTVqUByc00GBfyhMpyHLN3+pLgn1i
54X64Q5IB3YdGP6lC1QJ6twtI/CaV+DjOLERzZ4OAxBSH4LNOs4MzpPtqex5zt6ocvSfQAEh1716
nq3ImyXe3n2kXmrvzGVvVoIaMZxOwX8LLwgnT+dqrq5P38ObYL4fE1pfvg5IlwugwBlGh3dX4dIZ
Y4EMNofexfIonjSm6qL485OqxtMvAVM/8qUFO256eqTYzoX5pGZIk/6dBFO+ox0OyhXAuIiY7AaN
sQxjKpgEL4CaUb4x4sqS+wQrpjbWUqg55m1NG/Cirz6S4b3SXWhnp1imU5QjijVtBOBtFICmvgTv
KWgrQiegaPmFMLin3dkWFgzt9BP+cGlgsLsI6SAap2+ieN/wDVR/EsmQ9Zb7EDaRhIaP+bev8UPK
M7sWTRl+fgB0oNSKd5kp+hO6uxOdUfhHXM+XtSVG+9vFOeWss2CgBou9h8Ttg7niGkg/ZkgwNVFB
hSsD0Q17FIU4w7ecuJHVCQz/9JEUyQwadDLkcBbFKNZVtGPzlPgqjdhtVCxuxBjAJ/k2CCe261nO
qSvlwq3lgTgd4nVRWbdVneir0/jTIxEbGl/rwi+ah6YXRjdOWpBA9lUxWHWzHogLZripmDptMqtN
kuUGc+ps2r4uz52HC0Dv8wvaPadGxDN4yg2iWc4TC5GITUHk6Oq4xs9jX4yTIERr6BcVPKBYETI/
5I1ePXg3pa+Nqvd7Fq6WtEAM/1fuRfy5dfeqol4SIB8dsPnro7n9tSZHVUYJtTSVZocwn9esvo0p
oWF4oiPnAqRt2IWiBUBf3vUqUdahPabmyCEWx7s4Yw7JD92/iInu18eQtyX4lCB1uVAARDwdfiNj
N/e+jJgVrIqBLkv0aYVnTWFeDE+2RHie2m0ddpSTQD/aG2AL9jobvewT+u1Q9OJCXoCyMuZGhwp/
cyP+TukolUE2JH8yqVKWhOiXt40IheY4QMcfxEs6+oZb/mlPJ8FF8j68HbLfHfeAvXTXdcWT86LP
bWfDx5ScxOfaPmn0fWE3Ikdt3Tf2tsKA3WQvddwnUV6+M6aANybYf2YjGnXiG6/43nHcxdUTIVcQ
ydUbEzcQ0d6vxuaHZEG2GGyCgDzx/vquh0+5Uy3M7u5/tBwCWxdvwCUH5ix68hxVCq/qOlMwRS4h
PSV9QZFnDtgzdA9KOoBFGwhSx0qR8dUgZW7e1zp0cmrh6J8cSZTdfoOfPF3l97OL2tGF/IqUvKz2
1uplAw7kj5NYf/ABqUCJo4KfmZF83IxZvA+HF/2WleUpMi6brj37CJ1vVRIis29aiKiQTg0yYfNs
pfcpdPueAUWVsH29BH2+9ua0ybwkc+2DwRhg792RxkrVhep2eg59KZtGNf3WMgtF3e9D+eQ9Fqwf
uFcflIE12a3/i+Aagv6wsnRU0Pyi2+/tUuOrwZ5lq611XM1VsKrVvw64sD7heFw7lZlp41X/bLrJ
5NhiRqlydF/2mQ+OJC9rEm6ConS5cXe47Wa4KFAjI8NDr1/zBZUNMJLfGrgPj3XI+5lkUC3wI5AC
qGyygc1tJ9Rbt+N1HiRIHMLlfsrPondZ7gOUnqy0U5XEc3fFpGkT4UdzxgmkmMiY5Bgu0COwGUH3
JXn9T0ahshueK9nsToroKd8+Uwz8J0IW3ibNO2tGLgK3kyodKgDGrkehI8pf8aqCnmg4Rl7vhz+9
CcG2/aivpATpOGXyOnb7UK705WN5ont/tbL/IIL1jFpBAkaHlZXCdXd525SnI+mwlMe0zzdB6kLE
+2GH9qhOW14mnPym5v+jYbKZ6RMh77cV5QvrArhHQ03q/mceiHxONiDpkjkrWWoZHwsoRK3HhDDe
Q1HrcGQAwX6ToQN4T+TZDIj8xxJbuHjlK8eFCInCzvNrBl3eoonuBI/nnWTH/mtQ4wpXcCHsGA6D
//X+sZTfkcFlSTtb0kRwqeYkqbJpAKDeTzve4adM+A6WfcGygJ5AscT1rU2q7tD+aixnZcEfJ8mf
/+HqMw3OGjCSq/STZB0o/hgl0KiS1oWTEc/3FFY8r06Cstyoi6RPrSV+iaNh9BNNNX/XMYkpi4di
hE86erTpTeQf49UP4mbdmtK1hheez1B9xe60pw9r9bSgNAe+9Kjfw4QLIEReP3WmAwEXYSpgE70H
bZq2XxmNWe9iuexZtxBSFHAcONbaWAlv8s6uPp9iWspES+L/AkV+9wxnoWFyfE1pCPZ7ZviVoMf5
Aq1DE62fjJX31aTej0vBWLvmFeaLpJ/GhMnVmQ7v8OYl37N0wfUSVKx/IuhE7o3JtCx0Ly3JL3CH
oVA8fDrWRcJmmmduHvwrc+f0N3Gl0hoLjPyWEQnNOz+V5Bjy30z+127FBb/1HJP7+gVkDxyh+TTu
tokLO3KpOlAPOMWeKB8GFN9UJp+I6oNJMUeVamvSNNhmd7E8bQgR38drTFdLqCzLDRt5mzKKpnvq
XYvKtUibbuGk7nvAYy7bgOYk/JYqUPXjP4lXQqFUPpIKDbsIoCDw4nZrR4XCPZC8YnDnbxNHWIhJ
bU+ZHOmsC87jOYouOD18Y41B5PAMZLi2TkTADBW9adZFqHXFZqZDKDkNRuTdCelSVXXp4mEXtBMy
GmR2cDUmioS0x+IyTMNf3mTlIM8LQ+FxNllLPqWSrQB8LTOpcrTf6M2RuSm+xARWK8sQPWdXKs4C
AOnCIluPMm6TnVWmnMD5R7KyH932OMxcuEtDnHl5Y5cCdTpCMa8HiYgRepPXK7Rj6QVPnrAQD5oz
jxT6Vtlj7TOGgWKkY2S7RLb9LV6RN2rZYbGV/cRXYdK+2rt2JhPGABUHCKcB7a8PSQEwh6kVPP28
ckWC+h1ckqdzZqTTzzfw8QAXRR2qFqUMjtDsKv3IThI9d5p5LNbm27R4GE1lMKV0hSwbV/fWUB7Z
ZSSE4Ez725WNXPTKpMG/bIiSttjGpYCuXYqkOw5cQdw3KfHDHIbR2SSxez28IoE8X6pTKJ8iR40f
mDhEY0f3rbEkfTPw+i0A+7dDd9tX4liuIDB7Zu71SuudFLkwYNkQ1Mo8XGbS/zY6+StzF7c9ZZHT
jff3WM3hUH5UKsQnaO+Ehtle4XwwBYM/5c8uyP3uVXFzMIMTwH46hlNaxdQz35duezyr4pQf3b5R
bASY5jJeCKRpheLzKrmjeWU41r2dYdzBPfI+KKvNrf27otjM+SZfLlh3lmAzgQr3oCKsg/ZdlZNN
EpvG8vS3gxEZSiL6NO7QjHhN/ugwevaZQK3UXcMVo1a8jzqDs3zqLtFPDR0nMV3END/SiFSRkxRY
px7I2w51C0ynDjWuF2l8QGYAAK5TSaA43Y0x/vF6Xd4a8VwwQC3OlhzOULDosCm6S9fZX/xSrlcn
zKdxCHOTeFoE8RwiQ/NuPRZ060NCZcqTCvbNvZWz8hkTzkw6GoNut9PEZcsAxTsRAHXseU8BdyA0
iJ36BOd4rhdn0r/NG1DMwfVJ1UFPg7kA0OrzDWEZystmVlOMQ206HuUYs5iPnlk9Cteoloo6+qPr
TpNDW70hRyK6TFdVyicvcoQfzIYMck8+VyDNIQhH/kM+v52Xj8noISVBXDtUxC/G5FAfZjzgKFCF
hSuxZKgrDtQNUDE4RA1n0ZyomUWv9kuqpFIH2LemXfTsW9ZavMn8x3GCxfA0fzI8kBbkXCv23u2J
a1CQxF/RH+BnZggZRoLd0n1pNVUohcinMI/tKFH7vrD47Fv7JmY6PsYputN0jsGyCRr/HJU0IQn8
9aW87zNXInB68xGS/VkeORBEMcA7DmEMwuAhsuka96PDz551z0gv6mhCEjV+4mDxGVR2GkGEkttA
4LFnGqQcKI2+odWF3W77gbfeh9c5eCzYJuhhQD5M5QPHQUI4NDDBQcOVayQkCrSIPRgAi7KlX1U7
E0jXTLCLbRteMSynCaUJxPn+IWH6svz42i6UCdluwLcNsXMCzLRA1zoZvpqOKTFeuNDOQWugRQ2k
lW6IwFo0fOTV9TJ4TCmuAsbs/BOZTLw1QIg8dXs1seGStSD5vQ8qHPBkz3+xsinEN6BlCh8mV3In
eIxIE5g4cUYOXaq3eO4y1J/vfpmg2roWe9RXgUar0KNx41VMQnHKVC2lqSnoual7lMxvuEMWK0yH
1z4YVKhp0j4K1faGGRB3Sg6vmyZpsQYaRMPfOK1Y8m7Oms36bmcIRkLnu33vMIdrEi3m7ANZUsV2
kCuNgo/sYUHRoRVid5ZdCyNjlxYSCMZhdwrJu/F6EtIIlGHXVvTbztQBntQ+TlfWfntl5crr0s6M
EwlhLGuuqPCZMKYxKbavpTRwD6nQkYXDaDEtw/4Nrh9Pr+iJO55Wy1k6nWdI6qtx85bdmuLMAkwI
ifMXpRp4h5hmFNkrJHyP1Ts0YUhaSevXlWF0EDRA/V49N/EovbEKY6YeBJeQpQy/EWz5U9lL4UnL
WU5wLCULpp5K0A7B5n5WOyqe2UhFHibzGeC9WIm17WdvAWBDYX7WCn7bAuMmc706+AQw1jB7ESy1
AJI542dGLPUfzpCW13pCcgwH1BnSuLLfMDss2jOzQMLJe99JlIV78iBitxAiOO5FCoU16EHhTgsR
7i+ebDru0sUVejrgZFqgKdTwq2pLRfajecvVunzKARxCiuBKJTDgmIfyFiav3uxcvWzVt1P6Ln8I
Hz2dRoc/QkhTp/0U6QWAkpdmyP4fAdb3PWML1vkZRitRlYAmjbdr6tjlCt8ksbPjCmfPKJYUW+CM
Ap/g9sRlqqJhnAq/4uP3K09Bb4A/RbXINe/ou4eGnLZhWEKlj5XnlTgJFInyAbQvp8tZ59d6TZBu
K0RSzDJvi6o8FsxhSJxlGK8zAftV8hvZxHt03c1jzhIAqKfmqrTp7rMeN4jKH4CX5U1GwDRmGKP7
36aHYJyT45iKRbWuH0fvVvgKbTbu6Ec0xSEgRaus+sDYJzAK1aqajpfKa+8i25M6XAxrHUZ11WMH
VinKQqHx38UgmOcgg+6PUgAEhAy76h1CKVTbE2wF12nuI0yAgXb/GFouAACqmO0QP50XIqeAxhBB
WKk80yVHQR52XxVJ8Ei/4IQTOT0QPiXNHOJIZdbIZ0VYwBdMipdtRJFTAhkwkwE3e6DN8Pn2CYC2
HuN6UGns/veuxe+sOa+2kp2uOwb4AbwRwodDWH4P8CswJPpXA1YvVF63H+XD/ihnxOXF8XLn5/yA
e/OZd7kWUYbCAbx0ZuFIT7ZtTuMTT+TPKM6msYilOUKd8bM7w3FsYyaghGXXE3l70bWWu+9YOyGa
0qS62RyGSHei3jmIKv3zS03bJ5NjpahilD7LmUgr1R3OSOUehsZtfRVXc5UQx9pIUwLnfoUdW9su
bBywt3s6A3GsGFpQBx0aYuA6mea1soODg5eVsAdb78TJQN43Ti6aqYpd9nHmv/dnBJezk6JDpCyz
9Xr1ub7vplMnBzIdzjHG93tSPev4h0wx3hspzRgoTDHM6u/p4Xhv3uCfR86lYzTqrszdY2l8AyFE
1snlU6qFnuNaIMIp28GC/9tg0KzsFqU6TE1HxSLcW20lxo/Xu/dlyk3MTmOQkXX0Cgzxsa+i6n3f
7fN6BpmRBFW/hapB0cRGFtLQ0DPfSWO1Hc0lehnQcJvZ5ddpvkKaYn47s4PeHicF/xscsZknZSCw
8w2MBQzGwLDVEfPn2sU8bY3LjPWMiQhSjIrIM6qs3jomv00dKrv9G4RBNljofvRjbii6Ul/xeKq5
msD/WQo4MAeHQHiQf0ZxFgh11HRrhW1k/MeF6zt1lNbRpzGSX5/HVsuVvuLmzQDKcyQwUha3tG+K
fQBo3emauOufBWiB1TyzYdbgr0kx49nSWvXY88rg5OkO9EoZEkgIPUA8cEM4rWT4F83PXcPgA+n9
UK2TnVOs1NrxWhF9QP90uVndbsX/gqIcBjrpGKNQKWXSFISc18JU4LSFbwdZcgAlqtaD0myEewLr
0DofR/gH3mqwXm1ATnlCxVA9q19eF2J72j8J2x8ZcdywLqHPJvO4v8oypQFjavbj9DLr5QheNJUj
8/J4kj4w5LWmMfsrFvltDbUkFjdJoTeU8BA9jhGqEqAezNodGtlcpPwJ5j5pYEyTCAIVqO7i+xWJ
cIat+gG4Z2KkMZ22GpHX9OS0x9W5r7xLsXxpaMUZAmhoNHB6d2o+o65e7Ss9s7uaWcpao7JXbsEK
fytBQfytWUXTDqGkye9VlRj5/k/bRelhHO8oTeW1tWz+0yGBf6ryngCkiq40CwrBrebgqU20koOV
5Qbfx1jRYDdnGKt1Axrhs2of00JZmv4HNM5I1Dzg6mP2Gdi4urOTw8hE8Qr32LUJFtUpbiPsg6Wr
yjmZoEjw0Ms2vjykREtNHelrIPaDmfA3C6l0Mdtqk8vFE/41NvNW2rDibNfg9HYaPhnw8OCb6G/Z
IN3htNh5Z30Otlw78iUqcbbYp31G5mqWlGjBel+9O3YFA7/BQtv2Fh9oiS7kfPYGKT/4S8b6sbqn
1poGK8kFqhRDSq8h1MkvNeyKPsVxnLc6kbCAI4nfIxRy5uVgMxKHCk2crG5h7fhyLH/MzT6lq2SV
2ut9EoHfkzxjbRzY3O90jqPYS2V/Ll5ns8Gy3Gvc66zo7uGaNzvoLlKUA3pvlJ6GB6O5wCzpYq5y
8RIyQs8od8fDHfqO1KDp21mlwjqUdTwzIC3b+yecL8Mf0svkD5pZSaydEuPTKoCiOw0icS7Ka49Q
S6g7TzKRgLodkr2wkKhTXsn0IAo7CBZjMYVMMXigYIyYe5Px5C5DSjRut5QIgHdBStAptDSZzMS/
HUc5ELpu2gGvKAtA3xwOV/Yh2c9swagaAvMSkmlLgZjU9WRcI4RLxDEodjLFvSHzupTWWUw+16DT
VNY4vT0hHBNMcwOVh0SneINF1qi+c2fLKpr+/Pox1gddMlbofMX+zs8/XtlaVSGYnipg+H2zRa57
moNi2qbdlAzdx3uGi0S0+KcQUthZfFQnDt2Xo61rMaYS2ldEO5bAGrQeYRTBFE3r/DcFZYyKV+hp
ktWn9QUUUHz7QlOLWLZUBxFQUv2vBsDqL+4JLkxh4tbxVk1ycmjPnp1KoMZXIZAr9iX/zwt7lXVx
Ptks8l76isNwhirTpM1xtLEQqKY25LS7ZXV3cBpLwT7kTdiVO371CclEyGWYRd/F/O2VI/5xXngz
KneU4+7BTgVq1zT957BxU82jKvSs6g852XgFJ42qoKD3t9/Chx3XA0Yhfj2D3y6lOj5iuoqilaS+
ecSbKrfTVaHsqnftJlf6wJay6BnWWjuTsbBJRFgpSmCc4o0TGjXDm4sbedhtU3HlmHuOh4QBbRtN
9z36MP/n3j/f/ykebcuC88pi1AhDjUnTPaV0VRt/OnLGjIBZ0Ih9Ul1FDb43QoWsOTOAu927Xdz2
UbZaZ3yztRfDoBsDeZB+9bnzK28SB0Itsy0JNyRblosMMxsngtfkjLw5NR0ERGMu3RN5NHMh4OOQ
x/eDU5alL8vARpO/uB5v7HV5AzucxHhEuGMlgyS0rz3cKnwcJ782yRS4WDzdu6QfbKIfisHSMgAz
F7DsKplnkBab+YyyLnwBFCGYxMLjqRyZUYtYHXb5iENi8uBkdolCXipRzZbeFJoZ8vFSBKXtf7S9
JywGG1/n63g9uQ5m9UTC1hYKMn+lV8L/A/EfLoUbnCjEBTHxfXuzVAO0xZ/B1oNaaAG9pJgAR7Hm
BEgKPxM76jfkIfqdAdxcc2IGxLl6T15PDGylE1JxiahG1kWuBZc8OVgSfPcJqSpUnJq90AyOQLoQ
9/04HgBs+XAXIJxyxOIYZ2eIZwGUt4D98Jmjwx9AmJvijFdni4pTsB5ZP2XUE+J4m9O2QcnYn1c0
J/ek3L4Ds9Vtwe5Z1D+c3iQXDlaHL4vT4FLuJR3ovQPVL+vNdkOXUK0LzbR0G4u1EDNG9I1FN6bO
XikoFyMTU7RmM5DKmyloJC/6fDxMKGYxq7b9C2trQ51ki6cqLTuS9ReH4CWPa4T5tjlCB0oC/Hth
vQhCKkJH1WaV/YfC+mIZXiYlmzHDMvh1aAjbaGLzRVd638R3wCKrzPsVwWe/qCfPC9AvDQUq1E1O
gVYN3RWFN96om3BfsgMOszA5Wp6q4krlL+0OSL6F8bU5DrjH5eFfwAJrHUUV8kudFqp0HTzDpA7f
uNu9hxBRxwumDJzGy/nWalh5a7tRHDy9q4lZuIh2gNT1W67mFMNSRvSMW8fcP2iyjJkEaiSo1Ujl
pyIFeKeBO1MO6DgMhRqEIF7GW1Swebfhg+xacHXvJAeb+sYiQtBCuneII8WC7K73+fsZrII86quY
pY+E8TXMEyuK0Hy0b4Sw7CssHTHJFBfBJprzh58+tiTeSVj4JDerCD81bBEXezk/ZlLF4SALacu8
9jqJFTmuE7Bj0dTgXXvqElb/T5J/2APBvxW588odKALnFclGiHSwv4+M398JQ/4H2q37YKAJHY1c
hdhKzXWBEEyzCLpm/LHkmKBcQiBCxRF545RoAvO3bQGCRDtyqTnncq/J5aOy5OuwM4n4tcgIAU3I
cAlm33Q40JSnfjnPBXvZvLPuqku/B0OZdz5uw2Svxiu3LEU0wkyG9P+V+uSHyGnQUVRa0qUAgIPY
NsnA4kalsXtF2sgZ6H4iDHFUVqtpCxAcIaIbZ5LYov3pTXyxNgQyknl2rBfUe9GDfO0vrvVliw8Q
mIkoxezp9skYqrir8CIVUUtBGPAXAl2IhpF2VjpqGSO0UpumfZ/NREvBKQfm31QC28fuE3NixxOB
XrDhWR05EPQ5iR0Nw1DZ67mhVVNvqI4474z9sqUNcyEvTewBoTWGaYqLjXVnyH7aLdceK2u1c84P
IVeisQyRnCipcR6PONi394kPSk2yQnYTDwA3zTF7ppLPbxnhUbmZiXqw+smsR49Y2TtX/VjVCL9H
k4DHctceey0QDp3TSMwHBYdbXF5bm1Wt013PrHJ6sxbymWG54L7ZxUsFSArdSebBGTQGPspJfaVn
AqbVTtTQXvoWu5yxFsxGGnvsx+sDMyKZ+M7R0wxjazmKtG6HMDOq1zLtHGElxq6cBtUzEhQxbcP1
7C4lUD0fo0UBTZm3kzhYPq5ctQB4J5oy8/ryt04mTPI4FqUTKxsswDmf8Jo+U5dhwt+bmQWLWVk+
UBhr0SYDOMTMdrbyOL8g8NHEZPEXYbjDIhs2dLgn7qswvZ9k7zG/8p6v808Goh4Eqe8xYw7eUgwa
ALN/K1gkY3Ja74ylI0GTwcXwgtB5HX3X24qQ0ucZ0Wy67jeYESvG2kWbFa4BTjtTus+nzUvtksKG
eJivWqGxXxONw9Hz8xWVktNemEA3MiHi46rKOSNEqa9M8li2Yu4ByxJ/4uVCp7KUbgi69+hJtk/Z
/gBOfzcw8yHKdgxsYxvwh5kH67JXN1Ox2KCFD0LfEndrxuN8sWRALxmGiTEr7DYbYvQkNWTvH+g4
TtwTlJcA4gK+jG07gLQ1R65/qElkq6gWNSGtkUtdbKCflKKdpWb1u7/NpyQ5cK83d6ygX6YPfdlp
q2/WKX93C9rdWpnNszesMrNi76vTZJUR1mhrcwJyq8MJWa9DUyznarQe5JyNRgam+5ZxFnqIDKIt
xS1kkClXXuP8XmiVh62piKHutG0/VbdwYb3FZHb1S+Yi/8cyFCz0rmoAE66O/6tBjtwEnGupGIta
JtccyzPwnk1sPDGwXn5Z2uQHwadze6YbjsrF9DWaR/9NJJBpjZg02CZanD0NKyd56z3KBHD2HguS
2qhp8ejbA1o20mMbh9SAc30sCDYdz/mCan9DfP8+eW5VHEE5431JEjg4xOOebFGWjJ5PNeWT2CoY
7lfYdy5K67SxmBiDHvDUfjiYNUwi0iaq8aNK+9g0DJS302bvS/Cg/IgT06fQ6RVYYoaD+ts+PBvS
gdUDTu/gzUODd/h27ebH1xzqKoXx7Fe+TgndBgveGi70/ws6U2QVDKAYoeAdVzRYTK4mHK8NcS0w
iRQ/XrH+GeNaHTiCPOirxEBWYKGI8c/5mNvVqLYW30gRbLrNP7EAgtINOT08WraHmG1eiS/S+2j6
Mh9Payk5b8vwRrNmuFV2TB4m/8qeqsMaT+cpXD1HTpKEoKswnbpjA/DTmWPGcyyKVCrRElxG5kBr
x3amrXGDYKvqVEbWdNnnGDCX/W+j/YD7hf9i38uudPTl0ovQNjNC3B2MHydW6a4ikVnen3kIXkcB
opVWUl+BMkGdHkaCu+0uTpcWz28Xs9bxgGzDl1ByUHb5ZN1pKkZ77BzxJGG+1DMzUlzEcXSF4LDE
fAS7Fv0hJmSkBV2/vDU3qDrF8T3n7+qbcgOtMv8wTW4Q2uYg8YlxObft/7TJ/VvU/LfO4SjaSGHq
6cpyb7JYE97QQsM8TDw/6Na93W1A4/brIhleO000VErmY180aSDv5yfouEXPRmXdiYuRaBfvEBwp
t2AKyAB+bFBjv2fxuTZVmmI2FrroSALFnSmVjnwH67nMYYJ1GJSNqaXENFm5/2YRsEsZbhKAh5SZ
JcTFySZH87fhILYft/v5bHP2wLmSH9gmyJKYfOVlna+OnFwBx3i6uSYdzFKeyNSGjRI/MlqTsGdA
kTWopBpTrfTr2LeRRpyzp+zb12G4hTj4E5B88Hgd+EfYFJrmJSLJglsOo1ldvNmGKbv5AqLUF8Pg
pQeskxmWV6OK+QeVdFXgfr4F5ZnG+2bKk/eFACLtRiSSEN9BeQTJU6ew7OWtz1Dhrl0RON2hh522
np+JC929ldfM4z1w3oOSSgKlak89Bje3j4IOBPZF/slFJpnrEon19xlHc0a2OQHwzhGgokUMuPVs
xgeKIp89UnXLW+Jp9J3FlqgU6xdWcvmEQ2a9WBNbQ261opPGPmv4kt9mJvdZLwJXVVjcg/UeIoH7
GQqZq302iDtVXGsXD6vS6/0Hnw++UZwYFlxGzKWBBoST8SS2od9+A/xNAVnGxbC8LUdEiod0myL5
DsnLO7ybxwa0AQaQS9CHJc/FZH/I+7XPtaYYUnX0hI31Au+07WUjK2AlbOVa0C0sf5qfjETKe6Yj
CzD1z4UX9teXcOwpJjKdiEmjbwV3uprtrzFJ9eubCI+bXcT9IPcJsKK8ku8PhCL7Mf66UGmfoZHo
C+51ssnec1nV1TaewWxGXABxN3EsdU0vq/MJSNDa4cCiOPh4pOA99hYUIEhtG80y5XIH/KeVwMBy
hcMN5Qcj+7sEYtGloIZ/C52hYlPIZqnmoGDZ1aKDSSUAMN0S7Lcfq7hwSurqPs0bB8sij2J74qrO
eNbBtybDE3F5vuAQVaUNAZjTNwsmvQBNt/UwbpCgm2LV/HtcNlSVtDzNfjQinwL7/PDlFFEdYrqO
HJy3IWpWv3K7vlNnvHN9Y2GPs5DEZEwxrg3aobHhnv0kvHjLjXVrfMfm8Sc1ZG/k2UctQCJxu0SU
UYMQ2VYrLNOOkaN+wpdeGCfJG3oifsgYi/+OWaehk8hQ2yHsMCTjQE5aLU9N1r19e5AoSHGPUMt6
H3MrnO/15uX6qrbFbJ8UVlCpcm101GzPzFwgEowfXfhn1WznVqSohHJCJM7pB6S8Ku2QkdnVTTDT
AVbJSbmcy6uIn6hetZNssDer1n9zp0FzMZpvIgDzDU5HUp+vX3XbKSo3iNIfBHiMhRSBF4mGx8XV
IJIu3Ys4zTR39l0VoC4gQWXDrSxX10vSZIUAyHY3JIsJCIqJxmxYEaV5kbONY5eoGe6KXdzKu7m3
StkH9jz36tmYf48HdMj7/OqZaqvIirL+mYm8GRlLs/z2uafxFNXDF09w7w10OKGMYz3VrvW4pxiP
e5Y72eQ7A3OGPOpRxMXLHYzqMMcJzSNHKg4JVe9ucnHM+u4Eq9P+SAdsRXh9E2vkrlCgZjJyD2vN
dFWh1dU0bZvVzs/Y2LwhAaVncMvo61xKxO1ODJySIcK/sXoO6LfLefW3mx8l7aESA5d6Fg82SiRo
U8RgIsOtcM3qPSF48l74cu6BnIRnqPIBwZb47ClbpNTgSvJIa3GQlqKm1RPudlZoHpjRryc9mqeG
mdk2u3+7wPkdMcD/Uf4wzhSAWmTu0KNUwOoVhLVGO7yXfQWMipkQ1Rzbg2S1oKPfLLDmyC1QJqF9
vafMbmeAcDMoXLdtTEBWTMw20o2CWSvmIzvjNEhA40Otou7Ychmg9qd8i0Q8d0OtgIc0Qt6T6djm
GpsmqIFAoc9VYRZzXyJOXABZWfPdNyuTumGk7iyCEllgXa1rk7HF6O8i0DMpLb6njfv/voVgg5cu
QMPEZieqZU3Tc+AHsjVEY+NHflCSsBdEo1phqSepWraf/Obw9vCiUaHDUVzcNxqbRUSDrrx0UFt0
xFoOqZCw+wFoBvcdXyvpL6G+D76pq6HypTun6PFHCpo0l0o09PRjteiuc2d6cjUX6PTmpA6ZA3yh
0Xuhy0svjS3+YYFEZJ36revqveK7v4hfANQSWWhAfeRXgWSK6OLWz9aK+eroFQzkoqpVkXv1Vedh
XbthpzrgKhCxrxGCpib7Y7D1EInjCxk7Jb5LeBC04duAqtKnqgTvfyb4gqCOPGM70EIMIK1X0C4E
3uGDufhKWHzxJtQY+pedfZtTMC4Mj5wc8FQz1ejZvx4bmUrUoIAD9Hm5kC/UMNv8QRC/v0Cg7rCu
P2qHKpy2PBmxIN3GFsUy0U34BwrQkMwR8sP5/Nnynjb6sBWfhrkjytytrqehJ4r2XUG7vN1JD1Ig
vScJfiVfnlFlui636SvhkIeqazsYUyY6b3r/GxhCrHArQYoGhRyjh8uNxLgXoQ8wegqt9QU3Cdmx
kX+kxycJCgfxq8328nQkBrR+NklJJqi/oMhhjELHfwow4VQeKjJrcf7VCpTBs3qJvulfyirmL0Uh
JDF6KRNSaH5eADJuVSm4p+pRg/D81TWT0XQom0FWXLGpfcD3i6bSTTfcW7XsqmBTWqydAnSzGFD3
wLMkhcf55/O7cOCfYEcEBWchohf3adpMQm04oEGWlnfRhxH8k6OdlKLNzJB1WSsFFq8vYu8ZWler
700LK3dSMOe3IaSkpFr0t2MIi6GN1YCQk3CZxVMp3ideeEeahVV02XUJXmcqOkdMHuGUT+2S331L
SsGjfcymYHWCB/HzV2DSCppt0Tij+qXyxwNeJqI+zdf2KlesjSEeWON3+DFW+i6TQBmAboSkBOdf
HUVyEiqal8d9BsA9vp2zei0WuFjAuZ3AtBUMIEL5TQibNZhZhoPduU3QMofggpwjGX/HADoXrw8M
trXiYdNOVP33+imzOmRg75Ef8cztiJ1Pgu1E2zXYj1NNzLavTJSsQdhg2PlWjG3xLJKK+wC0PsQd
cmk5m7iA/1WrJrGCjMltqtGMUw97cvrdeVjCeGH7eHeYMemh7NA73sCXgjp4H+6XVDGDQH6jz5cy
VH+IoaKDemKuwn4MLfakj4u4DeSwvwlZS4rlkYkTjMiBxa5d4s27t/Csp4p9q5HdVZoB8bL3RJoX
p0oAvpqRu34Mxko4V5Dj+Wj87QtPatHn1B9wBtm5LSlQhOu1jMjt7wllDYehDRcYsSpwFy2TyzEq
Zr8l/O6WjgRTvzGY6YqSrzpH1HYIEvboz24SXHBSoC5gxqSzw4LJoFUA9OTHTrpIMaILUQXNim8H
NgEVXj0Na+5JW+adpRg4oceXH2NjOX575LrR6M2bqZOclDoe5rF6eR7TstD5kwgK8E868oM6kaat
RocbuaZyy9Y1YbdoZhyzDIgIf1AY/KwTP8wEULLPLwBCe+WwM3WJQmBjXFkd2bTnCqwXXmBZ99Zj
TKwx3hvdea8W4QhpZdklJuJeevZT8mAU0yVh9qP9B7y0Jzm9+4d0PvBO+8VG1irH2KSVPnGILt/T
Lu2CeaGEjd9xP3OvPJko2Sl6NCB1y7TeRwdq5VtETiqeZwRq6srUGC1e2qImY0aPYsEmF+QQf7Fs
0KD4gpHF1luy2eZpy8cCKJpSH3BRUp1f06Jvkfpd3OI7M/SS3OfTDR7WCTsHX64SXV6CeOTxFbdC
kYGrEXPM9ovv/+uubzGfORCgeEOPu3u9J0dE90pPi5NZpEmwjg9u39T/hFsQYcidchx+FIHdu8Yn
vtuxa0qzm7L1ZSM0YJ/SFkydcF2QUI+C5BL+Msob6rpK6nRK/3DV7ldO5/pN50ZvK74o/oXAAhoa
LZni/A14DChdFdyc4p2ZK9sr6xyQLnbOmxBYcuUDGTaGRqAmnmqWEeuUAyGWWGub8Ku0iFUzZLED
DA9sd6fPQ9PeCWnceGYOqh4SpWsVuzScbhRVEOp1rXzWewZHyS27yYBiYfqUT2We4XcWTFvqMIdo
qnxrzyxCROuUEu2pP2GriHevGb7RbL2u9ILnxc7tujnLikr+Qy/CXJJT3IclHlIzTogH7xHLN3TH
bAUbE4OUWD5SDVlljHja0LFD0k96xUm32oY2E1qmbUYh8pI/Xg/1kG+1vviuVfju88e2mhmt5hqX
cQEnkIsG6q/BRctTXYbeHp17GUq8fc9m46ncyP5d5RE/9xLgnK+IurkQEr3Hjwg29+xHhmw3duYq
7Ol3qFnhVvRnpI54uOc0hMl3bKCA6OniDGxhisC0sNpRcx3aiye1bF0qbWYkSg10OFaJcweIN+uX
frTLM0YZMisnUkgv+7Nj8i7z7e/qPSumq3O/XlMMnCT3rSkd8jLs8HHLBIy1C0iLH0vDg3lOILXZ
+dOGaZpnLAooC27iTwjkM+NIIbXJVzF29Ktkri64EqkX7GL4hfKFoRzvj21gLbruH9m7UPW9cT84
1m2Mb8SXTUZmz3G8g8HQzsW9yoNeIbmOeeCEdL0dJZHpnpkRh+zfnQ3avoK4p71pjhmZ+ggVpwzf
CnxE3cE8B47+CEeF4w9GmfBy2ZXm6k1TqQBvISkNsgK0Wj4Vd2156SUxPtcgCIIGo4gzKjcNNVKK
5XK6KNzldrJQ5wu6j8YEDi7RM0EvPA6Gv/RcyX0kE3EDcstlaNMs8ezpej/8hUuRHofOufGSwXpx
5M3k8JDv5MYMYQhmcWQG1bxrU05YkUeGIB6DN88WkPMIaUT3k9H/tC5TkYa5igUjbnm3yCyXLuoo
oNc4qpjVrpRQO9GVPt9oddDMuRTnB6nzHrH97NdYniIDxz2pb8pdYzA83PG1IcujKLEGdzz0Lt53
ayGx5/bVngG1QT/WuJ+c57c89hQ9VdW03XUPfHpksch+bdi+vTgLoWOfGcK4xVI4NqAqAx0pZp63
mMYKupyg0R/2CmzBBpobPtVSgufNCW18PfUW7Zer59wZeaH3jmIOgkx/XIOjOkmhtUeRBtjvvqIV
gMV5PJUcWoAzCdp0Ci9onUXbfL7AMeUs2cvDBBzXOFL/c819ohooLUsN0TNhx6UXSH7u9pu1W6iv
rLW1GwwOasXFHcJm9r34tZvJUvQTSh4tlvxlZpi7/YV+frPVFMWVmuyO4xNDghFXc+ne9ezIqMFV
HvW5VNB9XOuLxdbm2S0yKEKi/G14YpNB6TYoMHW/FPNSgBr3NyqQqMaTsiEMKk01//fmyAvObMEZ
C18+j1WG3DDMc8GQbr0c5/W65SNB7pBV9iqXmLD9Jc4HeaYbznCGJz687f7YVqAVKP13jENAWQRq
lE05akNrcKtW7URDKN3Eqp9lPtbS9+feLAAyOObqTb+7ThoN/kP3vG+IfQmshpAWRZXr/II9kZvB
Hmdg4YapplhaZThBAZHf/t994j897vx+SxUGZEypV2UMsBuhtpMhmT38hEdomOs8j+8608FpktHk
+0bGg6WOtFVBZN1Jr5DpMCjGkE5e8ksszhCMBSljvT2Ro5b0J+Yf1oRpaLgZGtllnOiZPmIkKFg2
EamladD6FcbpP5qKRBABAx9oOoJfOYHTeXz1T5btVWq2XgQlkJpoUD7O4sWLJf5XFBoj43FIYvP8
u8e2CmPpjn36wsaj3YC9+IxB5cu97hGINWmG/O3fLrt6mFN/IJjZdLp9X5oqFaSE4gFRMpxeoQKk
pGDRYY9JTh24UAoI5/pZ6uW7/tFE1PFF15pfkrwSOQjKNpqvq+ct3xJoeMZStt0PWp4DRydN5Odv
MvkSsZdW0woPkMwkooJHHhTwJ6hn/0JFEhc6ZxyyA2MeZYpBu2E24vcCt+G/SC03cD9QC1ZZrqZy
FS9W6zcRdXlMH3sIQcAbfergNZ08cWsBIM5DlyhalOMY4UJbK3xZ0FCRG/IHRSOwGGJy9HK2ooZ0
XtMxMQB1jBEm9QDQ9tz14vJuxrA8foggXKmotC304lsxw8pDIOATyEa9rsUfiI4hSls7A5uh8PAN
10CRvVt3QWM6cR/RDqdFZfxo6VaL6MqUHeB4E+0DpcFAWolR4G0PCruoZWpPcR2PINIGFByb62Dv
WVSJjH0HlYekKrs1QJQV2ro0s2Z6OkNHPVwXvCDrZhfKTXISdJZvvch+qzpAnAdrOaOdYc0w/10k
ZVA1qoY9Jqn+naJuaaFBIRTE73T0pcf9mRW2nQSxZU1OKW3cP3IrD4QzuN5T0ceTBDMXaU+4ZYnV
ROoFf+H6TVcC73Hj6LRshcDWv2nIM2Gdog4mT+mKPeBnVkFrjsBUjGTY04FjFeJBRWBhDcr4716C
2Dw8ViVSwBs2cTEbOBSUndW/JbC18onuB1VzqYOPXjPj4nBT7Td9+pnAabZwNSLDb+MJufDMvCYl
Lntfn3KMHNU9kUtPfwzqCoQuGw4u+kyQ1hMI0ehq0P44qvHZaSbNlDVfJ0EEzDhrcowE9o/SacrF
Noz6Y3Y/zqJJWS3kQx5TKyMsSekLpynqLY9le7iMywZH1rSCe2RKkilzsxCyYuj2yxRwUNsvEH/t
lkAZmctmI2FOwMs7GehUV7is8WmDDxSgM3iDNRZnEWzW+CIPwG8HmpkNsK/ZpI2/62WjcZAA9/0/
TyT7kjusKRoS7bnXDyjjeEi8sBA/ISHzgS0VMdmkpwntf2EpI0ZA48YM9PBp8XNNQdeh8OLFhw8C
2CUPktrkV91x68BTtCGbR3DsS1HXYbBVeQCiBsabREtOSpGBepWL8Nw9KVQNF31Y29vjbaV2vRAm
DiydsVx/EPRpLA8rqPqMfxuvKVJz63VO4Mf8WwvTFA99PpjzKY1aUc4/CvX4JoR993Ly9Wn2XQdH
cpudLP+31vWi2uQ+3rVb0LGlalm1E+g0mgAwuaJjsBuwY/h4riUDUxG+9XCaQr69mt5wBunhQGY2
AFX3akmgGXTyi8RXqW00srEuFU8n4U6F2Xl2VRC7AJA7pbuZBLEznE79R7hhGc1fl9OTYHGmM7NQ
LBTiipZXh31pWgeHIwf+tm9pHsN55T6RpA/cMXgl+VhSqz+uA/4buz0dwbURVQkR7zO1PQaQPIBZ
9WooSsWGNWiaTgO1rER6+EqcaQM6BHR+tvL/Y/KqrgP0/zK0ccqLFJ6N5LNPCwZ/+I26sZsZ2+s1
+FR9Q84FS3dvGT3EBxQsKmMr6BasjWF/XURJPkwjSJHIZ5vcP0gqDuye2VZe1iKu3GyTfMZmalsj
TNAdOkmxjL6kUaiKSDgXOcYAWhOYkfxct/W7pMEVr0rjQv5FsSfpbDN/m2VatGj05qG6ZdVqCfBj
0doKgpno2MDh7dxJHimg1c4R3GG3ofPn8KuY9Q7VE4nBnpS/fX1O0b6Ah+UFbnBouVnb4hOFXwBN
IfuOHP9LcQq6hQHzJZLdP3Qk2FRwdvCnJPOSqU3mdvInGmJRxcYuPIo+o7UKEM44Hcq9uc6AKwWx
jIbHl/dd1zDnXkdNW264+YWwxFcaMQKo9DIuaA1xkuUq2A84qecDhV3P11dgSD6O7wwgc5l+kqaq
gZzF3ER9O2P2OVmEUtML0qv4Gvl0gMaXhDy59ukG47MODTTJwNQz5BigZFiHY9c7S9emwxqkhakr
0RtZL8le62EMHrTGq55sLV0n17GCGQ3xCE4b7AtjFwCCsgjfxSsENPsiuAQ7FL6Z6Q155g3azDq/
0vvaFaUN6Khscbk2C9OgiMzl45xpO1LdZvIEhWndQZ70rwHxGgO6vYiwa1VJ4+evtGAWjbwMdK3m
GiUehFJikR1c9HnHG+IWibIbfru3FWi1aFf6qn7azoieHplehfIwlBKTBw9caNkfzD16HElbMN4z
2fo+cKkU+mU0p/J8DZmTU25N/tL76RdcdXdFdiDG3/7ANTFvwJgfL3P1jgyfQKPXFufMM1c85fqO
wq0ISwR/q53qePSqSJHti5nDzuiPsguP+E6XDeFTI6x+ArlmFZnhsp+7g4Cv73/BzScVRnEtrB3b
4UntuHojnGkzVGWiarwCfvnqUySGXwfzw07qjOTk8rrGX/bQP+ChU/S2IpSH+VPzLAJOAYhNNPtQ
yAT3MEabaRwNUULUifmSsxrBehJJyTc3tk17c4SbGtjSCX17bGEyGPI77oXe9sh1sZzLlrIahWqm
2qnAoVsDr6NNCRgvLB2LmJCnOO8zHGOLP4ukREhUdggowk5D2oGaNiL7F2bs8QQfIFHeFZJ2t42k
fJoujbi4FluU2vpvQ20v7tvZsG3IGg9Sk+Mc0Y3t9dgrbt+TCwbrkj3/i+9ysG3ogBETjxmIrB8Y
x5JlTVx9ZTpk/jn081KGlwb6/ECH/HXgWjjEqeigplH1KbsNCV2ulBKpYGC/fPtLDxJXAs93g2I/
XQWWRooOo+bkAO1nHRc0Ma6a/O+PywTHYH3uK/SJtEgKE2oHdl7QxtATgIbQtcmiiAxLmEj9Z3qe
BhpVWqu+quxmiPAGeHd5KW17Ap6KodJ7ecc2ID/TAHkLJQDHIsDrK21j/hWq+QwJER0uoDtv8LU6
qBTtgtyCkvdqRq90sZ4pBgh3laORicrtUMX0s53IvTsi06ageCwIMoKWFcgcDN4u/hQi6iGcWg74
KR7k3nvCuN3pyetmgxbQoJ6USOae4DMRneYfs4bOmMMNaqIaQu2eI6s2cYv+t/wqUyRVMLhpb8ss
wbC/MtwFMkMpwq24M4PznUPoMFMD+Wb97TwXIGv5WNQc/YOT6J8Fm2WljI+jJwm6bzcT/DIgMS+E
KgAT9SeZcZ2PdViEKa4eBs2a4d3VORVfg8HYnhg/90FrmwyTa+ZNFHFcgSL/WQmQtqpMmY8uN270
H5bqH8CScgnXbVFCkWrp5rqxRzWC7qDKlkR4cDgMr+moIKiNUc57krSekwfi3skMIap/rdozfem1
alNNwWiUtOGnjYptzN0l9l/5LsvKshdAJG9BiehMlmX/NmhcHnwldF8+7xpKVzjts59NLB9RkBaT
97fFEu8HNHeC4jGOTK9mwrrwBJDOhukdjk4Pa2rbmkG6kmH+fCJnnDwkkx4vnN9aj0poKkdGCblX
tlZnjrAsxtQadMCwTvBAtb8GjjvWAqGFkriMAUrrwxxrRVZphES9AZRud7Xl9AfmqDo3MKhttnkm
z+4cIMvbv2p6YsNPg9QLChPZhnDXEQKM8h/wo/7gAD22/vncZ5x9lWHOTfiTgK9z3OvsTpB0ldRq
yA6IdBeKW8viA/TaEVHACDYRLVp1uMtQF8nBHfd9NhC/C184Ge7N72JV/QgbpeV9iI5KVsqQy7yM
EBneI41cE9+/cCTG4+2UK0UZYcukj03b20pXcGIM9/ai+jNZl+QUNNesxM78qZzJQo+ZFGrLf2ir
Te00fqwUyYLiFKLMy/aYOj/TW9JeTMsU8D90MLYQUVHwU7LqjG7qK1h6lUJeUqV4d3DT+i0F0+zA
r3MJlN05QoQvHIp7PVZhDTXBKiJUudkSopEw592qfl0Wy3aAQPYWqjVxwPRH8tTpBqC1+chb7OtC
yewka83PRauN1UqAvQuG3w2eY4l8ZYh/gKT1GlQHR9Tr4E3LwfTtXW6JPRunJRtStRwBXIqzoBI8
b/v6AQk98/owAOPXqyaRaXLSThKdp8J79YIlmtwURi4r6hywwvFGa2vaJmCs9V6OYNc4VLcwja0h
hp+Fv9XRbGQZno9QNXK0e1m7CvMpLRPeNVaFiaXj46jm0wIo+1twfIevw88K+DKsTPlDL3QJkCHN
VGG+IJFvTp7NYU1Ir8BD1E5djsz1i0m3uA6iTUxoVp0NUUjWOvW0XmXlJ/5AsSDzSmO+bFq1aJV+
KwIKEf4fbrPNNVgB/xL5UQdg4M+SpPO+bwlmWfxIAJDKKWjAXsx2tQd2VdRLOljOioVSPREibl4P
QSMSvrPSfS0wQ9b0rUufuwTj0a1YtV1Aqgc/PvRmQAtYq3m+AWVVY+fyvxDKpna7/WupEfa4mv6o
nSuj9w1/Db4oW2Zu3/QaOyE2HZOTa3mpq82paQbCMcJHQ6QE9T1rts5NYr3jFs/wHQRzDnqXSmgp
S/JRW8+AjfbARsM+mJkZPC1gJ1VYBbYpaYRihS/owx0W4S43qkX7ZedebwA2AMRFiEEcpBn1NfCt
dyIUei8lxVLk2gJJmik4S39np4r5eMak9fZJ8lD5gTbWzNuF6CNYnNwQd5KB9/wpSvDzVuORpQXH
6sVrOBOy/++l5yDrCRrhm14Pub76C3s2S16tkl6IDseqF974jxsSzSHY6Zspe5sGrPRWyEDq/PZ7
dJxn7VWJq7ccINf26WADGv0gROze0tbY5VIgZpVhExYQEd2dlVtHByX32QEtWFcnFv/G3p1bFLxW
XOTtPVafmiGTieHOu2G25O1Z2vClqG1W9hS1WdvKYDkXadZiLJx9dKtFKBake+WNnREExPCBCdL0
iOOjElVz9nO0FbQq38bDU4taEkcgnAYO625W8yTCExR0yFLMSqyKhsfB9hIal+tGCsS2RkHHvSy/
1KwDtoC6E0xsgTCCD8V+yMfiWdKuTJWmRYJq+ATAlBPNhqS+AaszFnNNnoeDZNVjX/aAfO87DNmT
NcoPUovE9CshFGcwEE/capzizAHZU50LBgVj02/R3Cto+P/dWoJ5VQJzqeLXaV10YhhdZL38lWt5
F+QP0ieFhG/KWUVXiLFLTKnCCvzTyeVt7jSh6nZFn6Z/CZEABvSAI5KbB/Z4I1TPLYm+27jpyhwh
r6ydkn30Y462u5bmEYOsj6JrhFpZs3MDGfXL7fPT0dyos/R3K6xBR+APPFz8TxWtHaCa/Bo+4W0o
N4GFzbBFwERg7f9UiESjx3K2q04ocvCbs8rkgvlbvuyQ0jdKd91WCvNWjIdK2v+SrWreauORwmjR
tYd1FXvQGP3+z/RQsOslowMjZScAVGAyNoZVgXHxKb+bpU50L8GL72eT/2Gghn9KVMsxgueIpEL+
AM+Ib6F9XqwXGqpaGFbNDDfCYWXHojPtima9O60NjvQXNPDMvuH6jNYIwnSCnFnAvD9+yZN8Ddnq
mjKJ7etnHvybNhLGs+TurFGqC83zAW0vHSbme9xluwhIvrb+kZaUmjI2eqaa5xwmINSWxxakwbZX
ue2l+HXXmvZsmPU0EYg9TZO+tOhkUElZGgvt4iD7edsBOdEX+UJCDog516LtGA5h8FOvhb+trmQh
uijjEptNIK2XZaeHSGBMTkCn7r4FXtHho3AYvan8Ude2scvl0SIrn5Ba14eD6HfxXhRn7oyTfiTz
x66RwpbAoaDHrjeEzxd4eZorQF0OpxuCuB5+Yo3LLgNiai26yDNzuFwTgzedmJztvubrEo7mbAR2
tyYtUFa9/V12OupXfCrPFMdVDcs3ajL6dVYmD1HVUsUZMlxmxTasp7LnIh9/ApWntoBwFIKyil28
705Y5yfYTmO8SunAkkYgvV6Rx/I/vjVlhpfyJKOxny7OxwcP4kGOKC0+8LiqMNWqexYL2AfgtqCK
ZF3yWEI10Jtc0uB8VAbccGAdTWnz29FKywLrtg0rczCJR0IGtqX5oMOFby+7X8tZ87VaYFkJrWcw
zur/ypIKIm3/M5NB12qj3vjaULC2Gw9KzriU4ryVj9M7NCQZYkn93/CBkcd+WcQXp5isQtXn3uYb
w34LjnA/cV7W9ypH/tzb/LNmN0v9rII3DjgJon4Dgr5yMs/gfUglgWXm4OgkaHboV3/kVCx/PV6J
Rjw+K2zhib7BCIhwRKyXZtLVl+GLYLGis4V2KLYl6Vtv43sOnRsu+PADMb6JvEe8RTf0cMYq/3vo
bMU7P0xQi7ymMHsFbFvB6lYrmQtJmkwrcIx87mv/p6RZZKGPeykgZ3GAzI60Egk0+PG0AbQPaMX0
PvBZtMcE4wrggm7ZhI3O+A8To0Mx1zAKF5vmEd1/kM4lgNEXlR2FovrGU9PWuxdrqJlighZt4E5l
cpauRxU3Ltl3aL6G63tT5icrGtrOPq1+Lq/d2VKk316Ph1P2ZhJ09rGLCqTItsMPnXLqf4Hj5m5R
FB9+bZgf90yVOIFY0yQM/Qj8Fnm1vEpZCoiOS9TIny6gncHe5bIj3PJYR4AmuRmHcMQnVi2l9iCf
Vo7mXX1TLNVgVptHvZgA6MKmnCVTHE5StM2Z4+47yCG+g3rxvoteeqQlj3i7uCeH4g6SooyNmhyf
JDb+bCq6Xa31GNr9QKRB2734i0ge+CAn8U3j257pgcXnjseodNdCA3RTHJgwgFHte5sNONTKgDT+
TYL1VMNML0MWmT+BxrouKe5/hiOjFgUG62HfG7rS7h+u8VjyQDD2uetq/Al10sR6F+5FKFBKjqFu
TLPkJAjGgZbWirkieE7dbPLqcnsiTKwmOe2inKLuKdcxF9bWT0y4tt6Up/u7v8rbDDv+L9HvtFZf
b6pWWnoL3Na10MYXk8FMFDLp54no00eWo/wymqkTVt8iTU9dLzHhmGB2YAYqgV0tgBYfSdkVFDPb
VuWMVTTT/Jy2YkNscY/i9UDXhJkmjcuF6wInBiPtI+tkVQFNjnm8Gr6E+hOYCfHx7S3KEt0lf1l8
RGaEv0QPG5Ny7QpoWjmbraJqIvz8P3lWk8oUL+fBldXX8Q0JdtrN4wGtGQkxeporT69/EbhiF243
ebv9K5nfjJB2zqiRMaczs4CU3C8ESCOb3qbZGFVtGVaI26cwfKPK/15JEtScaPSgIs03Ovly/8Dg
Y2v6FgqrrjiBGOjCEZ8FYa3NpRZyaUot516zI6CkR08MnuC8N7tihi8TsZ3BywR2EaCBE0yJ3BMT
Fi962g03LoQj09fTawVCye9eSIO8CTGy7KoTLRpNgRfupmufDw9zDaJRxIKBIcQpSTS3Le/VBTtC
vkY06Bg42ijPSB1Fdt5FkKhOWjKY/teeP3Ww5/vtcGIo7mwx9KFRHDeIfKETjsCcfJbBN5if+Hl5
Wepv/ftzyippH+uUSCw3ODef4hiw7hukpsTWGNQsYB7GOygqXSo7TFMeA1kQb9CAs7fCm4LwQ5bw
rfLPeXq7SbtDGD9ewfdN3zGWbpmhAlQD93HJ8E2dae7cBj3F+R7AOZZnHF8Ir9d4hMyxMDAaqSEd
ToYBuSkFAPx4PtvNTEZuFjFT+IGw0XvKgbcWgfbSkzufO37Ya5S69tlm9b/rVYHrRkgLdVPQnOGZ
fdXmAg3arJH+nfRU/w4XF9Bt6Ss4anqwmS3F/IP0CKwFlCZelo+zuKed3WDGCn+wI/QbgdicxGh8
Q8dLgBEncH5HB+OepRb3UuiL8uKrsaXidnCfoLa2xP5dG1hOvLMf62PwMqef0tv5HVdMTJAaEgGA
0rGFqd+Cz88fM5XmcdhG2pkJt0FVrNqcbHmDhyqKIz4zZ034SVPJADVoguQMF0kCc4b4OkrqJoTj
1KjCu9kKSBx9btvWfP/uM/KjSLUG+IVbyxX2gjvPJYVi5LVpk6eIzEdrq5Ld1anER8UChU0PN4kE
PKTriHEr7cQiOVLJ5+9QYCZysFfqPepCgI5UzIKQuJdsIj6W/rVXnc049lJBUo6OQXovnI17JOu9
YWcYhjGDlFWuIuIqtC8OS1tvDKmHyjEemGIx7pfW+UWqbbhElNsjcVrgUo6wrBnQ29x3jT+efbTB
XLgau/LYDUrUl24eqnYN6W52m+2w9WbuVHf3VbF4FYu0Mk2GmPMHA+pkb1UTghVFSnq1x6rGyf6U
MEofrY9mYHCbFA3+uJOBi4aea0vUfjXArtutwxkNFonh1mmiQS3nqrkPTVvLR4fHBr5q96hxcGqJ
D2jalrZKpVc3IPPZCCQDavMA4vCUkIEDQ1583+KKRORg+3LhX+Z7TKrKYJirxLCUc0xt6xwsJB8d
0afptpAyJa6p5hrQ2nUO0VnArFdWtUvJ5o/8o34ZMjDIi+Yxbia0ablHIP/rzIzuHzpzM9/cy2E1
fGyTVsp7HT7jT9E/LV9sbTM/o+FJWmKa9NqSbmbKO2+bqImblz2Eng5qA0ChwmlWhgpasY2hcnXA
aN00npNQimD4s0PYHXPGU2zr1vXquwTlCrKQXUrRX8Xs7xktmwCoG82NfJazZJgYulxhYX/lbms9
QnaTQc+GGF5rNA+ib0VObbGtGr+JWZkK4dyP/NBxSGoxSULWg8n/vQmHrTMj9l0iK4YKNnC0ha6X
HSHzqJb5KaZ4BwUnj1nlAFIAABtgkbvMtt1ist//KfNVvB250RhW2yqxeVONyumWlDReeqlXfYXg
Mfaw5b6WiaaXLqL0xT0RCujGs50Ldf11nQC3TPwoVYycLpXa2avo+cG23UZE+fcho5W23U/yRGOR
H2WIEMPKO9COtQo7Fckpvn6Kz1+fYFggZNnKEhoxDkNQplLPxWunTa3BsxfZkFWC1AATMBRjbvV3
9OavKZ57Re7Ws9zlf2FEyM1ZzoPX1hg7BqGbIiM4bFZlzqdZ+yR5oBtAxadBeJqowAOcfTodq27/
zJ87L7fkYaGPEUTRJ3wTqDZ9SntWmmZ9MBPAAeuCkb6K6GgA0pz165eoNKCa6ZnwHCUETWfNtq0b
UmSuVEoBYCOnGk0QUGbtXuUcFVp8R2X0R7OpqSNW6ZcwlQCXceGiSOreu9NB/hCnHmKPOp35faUG
tTW41YR+YkQG3Zz5vADZJs+U2PBPV+aSEpoxmjGeGuagZzzsO6emsFtmvyUKYTQE/M5N6FqQtzUW
EZoLMX+bBQvDAaJLks0pmhqxPKOByXDFpqnAtdhSCcPiojtJjpMRtYtn4gs3GPueGml13nhNw4+0
Jc+ZWSmJD9y5HaHxiOvYGZA/+B2SS/7U3nfVP1R4ka/ZAGHKapcC9wR/BeIK+sjTVpfRexnoRYj5
fNAShRSPKeGlRW+UzshZc/L715tdu7Rt1IbqcqpcR54Y8LnrnNKNYclFKLxBP7xSS+/d5ei9J7ob
8F6KliWCDL70ZPw/a0MVx/TRT0LuYYjDbuFWFyht4gGT+u30ThCS7Z+qwCr9C/8t9INyZ436Q7JK
5sRVH880uBSRDDeVFCfBAyIkrMvr3WGeN/HKHjF6if/kp/L68iuYy/IwFI2ZzCHmmHhoaHqQ5v1z
QMNPT8M0hzNAX/csmSGn88k/MMmwEzmAG5uNfb8JUPA18kJuaX0O1p+90dvW5HUUFnTqjOfX6oY2
GPI/AspVzFqOARlt2oVJw4HYZe+lCUs482M+qbHsP7oeY/7mFbaImic20mIEoRLvNqcbRuryQcSt
r0rX0zKjiPCT6Z/KBhrdSOabPBadd6nQOMipH2Q/Pio9kVqGTRqY+h7RRpzpmxc21+ZOeucAPLc3
/vgT++1mnXw8oPDEjfx1eWY+WpFE2mZ61JeZ0y0XyenIq+qj0Yj0+prJ8lCxlY82v7f5Rv6dTxa0
GAUpq34s1OyDs4aTPj5csvAYJVJeee+K3973Ykv2zOe+MgT6Lid7hcfwxX7vUJxahUfIe8ClGYTR
8qxHOSYdpGBHZPN/5bdQRxP/Pw+2Asj2WFpnq3xksgFxMnnHsN2xKcSxeOGsTaq5Oa9NvQy5AhmS
CQ879pU1Vx1S35eeeqkyh0f79TLrUaeZZrAePH4pf9qhrKgTeLyd/Hzu8/FZmyzofVSy1SSdmmMJ
ptSCFBasb2Hh7/l2uPuOA1G4rDuvGQ/r3a5PaUARruDloKmqsX9JpCxeGzULpD8LYnqr6oWmJhox
D9KJ8jfPXQGjrYGIdnu4Pbnc4UYlhjm4aUWXIopyFuV8AGmz/UdPlAuVSHRllfxP4hKPoIcbULnH
y+VcWha5+enlZz3skh6GKN/M2DoIa48pEthxZUKgbC2jc9CU8rJUwW2aV//mIus4S/8nTEQ5eXdK
+PlTcg07xm7gIfbZrKyo6yNqyYONo378exzIch/726WHyMvzxGzGmyUvcajGyD41sJJSd2sCVgsT
kzDrF+5dQQe5yFUFHba0WwMmKUHGqk/6bPpypsB1H7d/SVOZtFvE+W3k4MZ7CTOdobLzcwR0kBtL
uam/BxTDFKbh6opk2iHESRaNK8dxIoQRjFqjBuuQOJ8xn2XY6jtdfbYYmNom4Tthb1TxczVUsoX+
VVAYAentbhho/gA+o4B0pYVassSEvK+Dx72SwgDYzPvA7KXHhFtKVnD4yEJmM25TFJZ8uXA1Ygkg
pXCvRO1BQDkjyWwRgy1cQj/eEvuU8DodlD45aiehYo8CoBQvm9XF6ZLw/UHZbSWQ+XAX6XK30QTy
HOYAX1Bd3k//UZtkTE+lHoqWuU16G99VpaY2OaSR+0Dzcg3bj/YjUNgIBAcBygpuHLk7ufHDWoRR
weOzVKtLFR99qPgknq3U73jcZ6A2u3xFB1r/Ale/6VJBmc+X8jmj41G0AsoKjFiVnNfOA5tJFfNI
I/TMzQgtUyTXcyhX6P1z5/y58kSfD5ljPnLjFkQMClz5rgtcJQIdqCFhXejhK+wyhDVQnbxCHFWU
pSjFvTmyneAIZf7qEU8spgKpdZH6M7FdEmFT+CRamzWky8vFYE3SDd81T5jCyAHo424tbvW2dEBm
lqhpqk5Z76WgInSCv5S0SfLjNou0XdP8ZgeAiquc2P0FY3qabCUfflRGDEmn/D1P6UfDg+vI70tT
LGkObwWshWXlLccCpDjEG6qG8qG1NAdXikRpiqUXDTpqx7mQuBf//mif/m7vh6GP4JksOPpdJLHc
WFwTsgDO4XClKjyLFyV5KPXAnPxAg5xN/qbo81KyhLxtxMAS2Vm5A4Py+9jf7kfM3Iz8QGFDxaLs
MA5CWIVpAiFmQnmC6aoPqz2u/8/TO92jXeWjEadOiuVvbxdKKXJoR4y+Q92RBgLbfpanVcXWEPG+
f7UXdXoiALgYV7JrSzCFga0hibc3f3sxquzeFUylzDnShXnNHIa4JPBetKZ6LHhMPiOv1IM933xv
jZ49VWOuMgO983H6wLvWBVWyc5Xl3PJOLvBcO95iEoLcrC9Br3mExC9QrywP8dtvtR8DI30UaSaO
aQMWw+lghy3s21bDyfgJJIbgXLqhWuRyCLzgiyUeSwIuRZZWCdmWN5TpZB559n4+tSBXVMyotu++
BwYHd5MQHg0GAnUlX6gbK7/OfgPK1iDFsATnUo+vFn9UkkGZvzjIoMqiMeAu3lvRlQJf4NnXqE45
FNRVbYulu6sy+poD+uxgwUFkcv4+m9dTtIfK3EEggifI4adC8CmTPre8z2ILKAlO9vFoFNygEUxR
Pqe0VoKlXatVO3MnFl6wjCZJvw3bLry+htg1K7Fb3GRJFPsSp/hy/5r/Gq52FfmfNVbvqsVLX45i
eDWrp0tIKf+1X33v1H4zCeTPPPQVXtHozbUeQl7lWJJ372g6ye0R7BHQXor6nbYdO/O89Cd6OMJx
hf7v8yBxh5rLdRIjUyhkspO040my5aS0Jl067XqBt/CCt429EReuc21NGCBIrp+VNtngTqWwkR1e
1Bc0C7HsJMni63Omb5fdT8+wVvwcVKx5z4xGf7vVa1i4/rpaynL9URF/iGSgOItb/WMcsivpTOZD
9czhd8UP0r4MGOHikXSzW0NMM5GEhN9A98XMKzNMlpEgQGz0FnykvahzGQq/7KAkjplJKe53zbKv
NaBHTsLp8tleftG2XMQB45hj2+buvdiTT0CnWxVklxE4VQdAwccxYwbW5GiDDxsefIqAfbnlimRz
RndX7QlQaog24o3QMdfSTpVOHJdrHXeiZ6v8ATAxeK3pSshYB0W3ciEmBPH594ubPrUoNWQ1oXjT
kEQV3DYoIezt/eOAzxu1ssCbfwkrSr3zUfgmok0tTJHsfNADJ2KFWMaYxxvIDDgFc0TqB+Y3qHN3
Yjp8r34MA34sL74iwpgeTi6wPX2PU0RcGhXSFhXsapTB3rOYc8jGYcDoYqntQfpgcW96L35JfmtH
CSkDJPbfjeXnsjLV7BkfTB4HNF7sdI71iXJTIxkS8tEg/GLX5+CMV6M0WCHeeWxc2wvevp5Xw7oG
9MYU4og0mv1M0Q26fouXTBw998TKHS+nh1H95Rt0+UoBdYHhQfR8Vjx8k/wOzm5929116XLwrj6j
lo+7KRn6Xy9WgFrSKYKAnXKkhU30+zf7Z0g1FsWNph8E711J5GswPkiuVQM4bSaHVTrLsv6E+oZ1
GQ7Xonv3Fh92AXrsnwvVhcMeRFNr3ON1yyJKb5Uy0QdYGjtXpEjfTTmoDrZl/Y6H2WXNw8cUbpkq
K9TbSQv4jbPhcm6DLO9D6Gp2VNF/i0yieMUSFHr6fV+htprmGekH127rceowRMVdpSLuhzS03qNW
zl+9hgSG03yrXw4qPWmvCm4rauW7rTiHDRU2P0Qi+kg21i29KuOffYmYgMw0OrzlL4ASb2shXbDv
yaGs+4ygGn/HoWDf5za6IpNQTlO6zqy7xwM+zIholOYEODuxu8YAYbsSMMohlpR86EExbADjDVAA
5yEZGFsh5XEBS6yz/jr+0URwpK04ZQCcrWzBFlM1rpEkwpafl9MwxgbH7mNvDiPdQWAy1tF5TYI5
asNEHORuIJ4GVv+XSIDt2Z0K0z2gjbva4W2Hp1x+WGTNDLUAWd4dak+IYckDHNj8IWIOVtYaSAog
9xJ0bD9TksN6qEuTYJaH6PbBPdxxmhm5x5cPg9iAVM2n+KXB5bmB/PxRqU9q6c9NVMSGr5dVvXYo
nwx8OKYKwY/dqRXbcH9DPPan5p8hM6ab3DubnA2qGcBXHVIBFVLD8P9ZHRE4mjBm6Mq4NmQ5mKMJ
QpC5SYRiAwbg0u79ZgyzvmZ1seDMwfNj6eNiFiUa/iCDpXt+hL128WJSZxqtQeEdM8gCXZYBr+W0
YbzlrVBHJr+iu2oFuoKgkGkea08J7Ec1ztY369VLD2jn11kbMZAN8+dLJfntnFviBk43UXyRZ6DG
XyNtHpiJu93mI3cKKjlAPJrXIdKaEUmVX9g+cx8p5h5rht8WP8GHgk+GKET+wjD/JaDo+VNRcqTI
axdEZVmGCUMxLZu2csINHEdAuKRmbckNVtEMJS/JuzQIGYEPmRKPwJJ8PB7mDBOoGF17hCxxVkHm
WiL3xzFoC1CLmoKs1pxeYuH+XvVTiuKUq7xizVk1O7M7HbjZ2PbVN0v9dxCiNurk8YOpjIqLL/Hh
mRyFfD8fUXxt5zFN2DRd5LEYbxTUngR6Iv7EDFHkd2/QdOptOk45tDS1FqxAIyl6wRRME8bb76UM
We8uZH854GX4WLmLnx53MnJGx+4lWL7PLLLU7stQusLQkcah8aQOp6a1uvDo/ndB+QvqhnxF+/Vz
DscIa5Vj5fROEpgsE+pVxxnT8loZ0n+/CHIwPz1gQYA0gksbsqtDdv/0lzBnoKM/qqQlUUEHd4GU
BR9VeIZooNBCZyGob/EVhUe4bZLzgI2R6FXBalVvuAf11nIQRmnoUgC84KIVeSFzz76zCqLT7FqF
7eY0Sekz9e0p3I26jtlHSoxwuskFxpYIMqJr1QVah7FpR8/2evZGRAaByPU4p3galfn/y+ZjCrOn
V0F4gG8UXSqHwWWujcml/OUROMxdvKsUS7lN+3tZkzirDHm0br7ddYFMmvGfNeBkJffjPTHECg9x
Z/C93e1xwemVa6e4FBJOntL5RHbnO4w76AQL/mWoS8KjqMCss7gwuog5Ut8upW+EsWdYrGcNHxtC
vrBBxo9Im03s1r5aptqV/pBFkSm++TKcknlcAYMZzVnrMF2pc+Z/i64l12WgonWPfjw2c/pW6yJh
6Z4ZvjZyJ/Z6SjGdajvA69vExdOlWle+R+DNgiYsBqJ8J/wEfSacXI/qY4froW++Qrp6icF700rH
Zt6BpjYfOOuqcn4Y3/vb+l9UXsf1940H/R0Vf07tLFGD6efpqwToLiOqk96+K+Jp6ga+ET416VjD
k8Jkbry9MDutFevFgx7vatDhOrygmSa/olyQR0wponlEAhdEGvYlJL/v2t/irhLisnLBlWW9Pu6Q
zUNuJpH+Wb+26CrpQDOkZzicttHC+qgD73SkyP+9EvTBTo4yARpoP6bo4R7B4BRqHBnGq6a6WXFA
ef+sGvoKJ4RVTiS2JtL4Ofw4F9RA7xU6rDsNGi18URj9FO5m8SL2xVzUclraxSjCb7/RbY/u+mvE
4VV+ZJyzEq3LF9lSVDf1E/ini7PH/AE4Y1XfvlVfFTMu4idtV3aJdN36wiEqn2iHa+BGzFhZeNSx
BvdBjgsUJtd688h7sDBk4Z6hfm25B+MX1e/my6OIJB2xikl6YA+T+4e+oJWlNgej4eG8d0pC9D/i
j/+Vaqn5x/1Sq+bJe9W6csRZMgxpS4tzPzvQUskqFaW5SmAJDiH6xkg5oJ9WHVuj4zz0PycfL4gj
1YsnEnySFghNnaKyQBtPLRM9Km3+X1rFkA5jVr2Nad0XU+PhnjjNgUds5F9s7a36NgrwHFqiYUJ8
ryPGFzVcfzZiAoK28wS+1rLqlXPwGH+Y5TK6g4pmNqHXPYhJZzVkln5nkIm8wVNHr0LrgCMgUFgm
Av2NRGXuS68vVqs31KD5zIZUYyuimToVANpR6dGavfcyHLXAm1Z2emFzvrOpjKh5Wi4/fy93DdUd
TLz9+Is/oaMtlIeYC18SxF/IQyj/lwuMdRXvkD0OyB6kSA2UP3rz5ZKhdpGzU+5eOXetYFGYXSZe
ig+6AsT2WVFelM/BhgcRsTUi7s3HzGxY+UiZebhBWhRey6CLlZBpcSrxLrdK0NlO+JCwEwsHABAw
INaeP+/E1cYwxmlLq/LBKco4kH6lZfTxkf5C9NlES8XtiZEFGl08j/eJTLXk705HRnxKjJYCQ8wn
Jt8Ou0sNipHdZ6oQpVpp+zcg07NY0zKnVgP522PKvxlniNT/XQBmtZBP4DA5sd3F4yBC8iegtDIN
yh8wOS+RHMYRwp3kFiCx1Tge2Ea5JO5hRwxk3UN3XTpKH0xFgemBlVxbtiaA55mRf7pryM9OSXE/
5fHEHOVv5bnO3qWA2V1k2Tmuv6mmHv373CefPOy73EMVfyqsK1yOmSf7ygFV0VMPfCUOmuIr7Swh
v5I4V7t2Wy4OCkQdC0rZcqacoznvyVDabT5//PzM6epqnbunQ/ILjE5ud3XmjY+uM7qVpiIDqu74
+7hmCCsnUjr4MdVYkPkA8q7suskQ6cj6freJYqGP9aFvJi+MPYNBnwzn00LNDuIsBpNUOg3WqDTS
mOFippWJykr72gaPQLiCMcVY+YaJK4VVwceKsPFB4+AqAxoEfU92iLJFQ+Pe4TDZtFA8Px41avPe
A2eGQsZM9cY0kjHMWgSK/XAuE1gOKkrSwzaO2oSCg5sA1d0aEwdw0/13YCemclKOPrHj9MsdNjXp
6yqo50T86Rm7wEp6fhK6HgEXY3jHIZodkm+tzzzdgi2F24D+PobrNHgjL+T02w0c13zpEkRw7Xm7
XahY4jYzxh7crJelCD8FekJV9kCmkamXCnd6JC656tu3bPWOibRmit+PDd2wU+RfqyPtYYZDLjcd
7fFRw847pAFE/fc/qDPLzOlF1ePOlwZ+28i13JJ3W+GshY9B1cT60QQpOJ1GPWgY6Ykl/3ARm7fs
ocRQrs/CcV1zqJu4s12Duh5PXQGmidV6/esKDKjU0vp7Bqp54U4SeIkiMi7HitrKs0RjXuQlXyvX
FReCboVDiAhLljp90OefH5ZYU8czUyT/1b7oZS9sKPpdlTQMQKE/jlJLS2y1CQG5V2l3PRZsmR39
RY/lOUfv9Ov/3vTAjyCY+hV3Fg8g2C/kL3mrbYPzfVD57SgCCv5a5GgUBPAkEGHdbkBVdg5xOonP
Fgn0kT8YwoE4HggRcDzMlky/Y96A+6h3YhuwY4s+FQLSw77tSfJJhO//tVC0y6c1FU09XpZ4D0FR
rJrUiN0WvES9NCUl+6erVLb/ZJ7fG7xVK/2DjGBOV1nlcJyu42CRuWJMSXf/9fyX8K+xqnOzn5Kj
fHWt44iQQgsM1lB9fufMgX9zNfC1KWBTRf3BZ+njr+u/0Y97nLqvKd4yXLvHzH+HenECASZB4XBS
hgw2jUXore9YLLCibC0S30cA9E621RCRq01rEzjpvsfalynMk4ZpFMi1wmtrODx66VpMhrD9pYPS
+AVVYfQF8hp2XHSS7Vdvnd2Oy0m1w8HSACPKdeIbbr1CQ9QLPKmfePa7xYLf9nkdW+ORO6y8cwe9
BCxHnjESCO/Q7QTr63qc1JZz98Plvk4pAdOWwUbEWdWI1Z/zU5DjbtV5iAj6bClR0f1b55BPbFPR
Gu1HcXOyQd6XPB+qM9LMU/VjSm8eapd8oRZ++DmmEmTZllKtCzDd6F54ZfrjrMhHTq/nwFEARnl0
GRzZD4xL04600U3q3I0+VxX5WlFmcUxwqA77KcIwvjZy+7WMH683bCyhjOL/lxGeLEFFw1ZNh9tr
ZXgg86+2pR3xLnuyaqyyT2g70t1Ax9wI6M1LwdDS5GfZWElHZB8FxR5UYNwbCH7pFFW+yaWECnUP
cIVXvzG+J8DZZZ1MltGpbShckvByXbCzxKJLT/P8RNSRTsthN1Mi18FTPhLbETmM/x0wQY2s6EnL
DicuYmqnATlhnqkbaNcFL1w5RqPZtolWcUV2N8Eq0fztPsszZLQR1Uzpy+im7yVOvIJM4u8/5zMI
RH+M4IDbfR32FfNhlB+M00v8BKmMFEVb1feeS1zXAQYxUcy2drgHmEsLJAhwaBltOmFhxLk01+hZ
ptYmfIMJpByX25L4jNN/85cKefJ3k8r4d11RWaNZnWUXFvHXmgOlidu7UUbm47bTahyX66JGbtnj
pq4FBX2Dc9xd12HL30NdfuGOIetxJjE76hI7t61kZK6hnV2/pjr1/8Dk31BB1WMGc4AdgqLIgxX4
ls15EnZJ2DEmqLo7QSPjU11Eq8SmraZt312kRB7uDin2Werw6+iuSapoj/fVXbnTVtIBmAZvh/Us
h7OgZDdItojWJM46Ul4hx1wsH4GGcWiL70VPe0u/Oxu5E+ERnJGeRFNCBKkWIcr5G/xo/nE6ylqO
6FiUmZP6lka0DQvvn7SGEAtLqUwl8cBBOsDaitmG6oxQgYi3g9ZHgejwhG4Q5R8UxifAeHCwNWzN
FS6qkzOjdZIwkbQndyDA5bC3qwf5jv/AOPZT0rwxTbP9oJzN/weDsQQfIJUElsMuj7OGHGyY301C
L/bBZeOLeghlRfwWbTxiawb9S3DyL1U3Ng/g5E5IQGSAkXwdFu6Jlob26X9RX0TjJxoxSCRdPic2
db3B9bxYhDhmoiOMXOFAbQhgDlBcCyUO+XFjHsvUZnKJypRbVQm5qOVEtkhYv1zxBaADy/MzoLc5
kjjiKorGXsa2pU85ZcnnaFIDyG+tpY9cK757KEZ4RlatGu1ZLY7b2m1jfZls0vcK7OuLFAwKqqT+
NFYFyeGzvvKFdbcBZ3i9/Ma/Ju/kJcEzKCvouuvt8z991NhHSDIB0uz/i6ZVit9RfAj+ZUh5KzqE
xaAikfOIdhGpF7Xg+GO4y58vo2Av2boWLbP8adWNN7Ol4ScmePmMwhgW2cM6mlv2boRBNUyz416C
6cF/JhXKvx3FCNY3RhjXEjVPQvAZTI7IGDjAljuFNYq3b73xaMQWBGVLT2YIeiVKtw32dWYuc0Jb
HfaNr+P0Y3HigYdv0xxtKxvB4gi0n+5ElpEROnzr9yuDMfwb4zae8PcxR79mNlrCOXEbKhMi7QYq
c8cTkmZAXOB7aA6qIq8W5fcB3zzz1QtwHMSvHw2nkwElthwfH34GRC/RM8NG3/6F0yJEqEE9DI8h
Oa2sZzu3sQ1e4LsGYqfI5UX3ICYc86mCu7T2JRvbvTjYCgGPft2NZKVMDANhtMR3o2Hmrh55/d/+
dWkgKJ4PK/6GL9X6ngMlPaGbe1AiGUJYjkyBJOjoVsdlyCFvjzK/yGgrfzg2omgUWzl8bEmsi1vz
vXpsJu+nLC8LCO7mCcC7unTMT/biJoACs0t6F1C/+4W1DUHStEuHCaNZLmF2EU8UhvBspRFu/FwE
giT+jQSxut78LS2g6vkkH41rXRSvakgJpPdlVOs1d5ZSL5DjrLHKUiw5VT1htgI8MLEpXwF4DmPC
xUtnDFZK/w0nJHntLSIIqzVGji03TA7WQwVqui6TYX8YvfkmiamxB70CoLUuZC6128LlmKJLgusS
ZhWUhAwJ2S36KzPT8zo6ftcuobyvG6Rf/hPg7/St83frcvYiLA4fgB05BUEgULZZnKkapgVwVvnG
d5JgiGPKu0EoyWii8chff5vRIzRkL78XeQiKPMZ9IMJ0FLltKbR5lPcRFqLstX9BCn6r5sT2uqo2
DSnjD3ongyFM0zEPdHC9TujnDVREp1G7l+m2Yx51aUOehf6LIQTGGIf1DZpHbYvmUJvNycx0nbBS
as62N/8n5oivf7s2m7WKkfNpmNL5iAVLFEfTeA33oK5mNyNIeQcme0M8Ux9Eq/JGdSMv9IfVjfEY
y9nUO59++uQOM8ok6Wv7X2NBLFwwaSmuwZMhFdA+/Q9XBHAdnl7S5XzWREQr1yueAO35f/H9qpz1
NXN5vsXmaK3XXmEBYEk5EN+H+QKdlLGlLHe8bc5l6tCfvhxYXUzUu9jsMn3ksk8EkjsjFvgFmQJr
DqmOeneXJi5mAsGglMTcH+KZAFjz6D693PaOgBWKAUK6wpLr2PiQX7QTQZ9SCaNApnNT5Gqia4JG
K9RmY2VGY6YevwlWSurhbhK+mUfwcT65UKFcmFOoSMDCvf9zlKNbanV+du+cl9LlOy6TnsUYRdWD
RyjD7qKhYGX3CDB+lhYPQnrdebLKO6+4aQvjJI4RmcO1moNTTi6c1w/0UhxtlsQNFjjKDo9/0AnT
KgLbOvZMj0gMLjJe9v/MXRrhajK1ZO62fP9RkI3qvh8JnVPnJncn51bOsnXCSczn21EJRGi073f8
jrZNdn+mmBFmGMbJqfEKsoxRyx2+/6+fSpcBMCBnCuuLl4iASwfElgy6EXZep5fqorSNpfL4f/s1
vWDb4KFLyN7duPhj19vIilBQogMa/83TkA0LZnnpK/V8hNAeuwXUBCAbFY38pjPY8mLEynn3p+VO
x8B2KvVrAGf7a7L0hvkMVVBTZctaN/1g+w/2DWBTmYWvZcpwCdAhkAufy6mq5uCtCddGlBsA/VCM
5UmDwKiY2815fIYYp+77pE+7MbvU4A5s2Dvxo13fqeTFwvkPB9znRb2io9MjuQc3VcO39KWJG4CZ
bO5oDC+gEOHel1kKGcoZFBAFmndeqMapnTLSukQl2QcZxuWXeMT67agr2KJ20JXr5iDed1PvHBJn
c5sKWqanytIiwkNAvd00oSnWwJmds4BgZcPsxtWfPnXYt+dYaxImMrwJvp4lQPUWaTDpcdLij9/a
mqNs3wzgUspdF3Oq3d2is9X3ygzUNFaAGxagFTfb6L/bNlZhfosH4E2r4K72Q0hUziM9218mtmuz
cXmWkvuNc/U396IHFu9IBCdtmtqPlAOIMQTj/ApfVbT8lkMLx13NxYxU/yeJzbKLYpMqc1wDW4hj
yZuiKHcK9VM661yIdvrTNInXrrHk58gUA1yui7i+nVII/TcDkZljLu1IR53q5ppPHNiOf1Of1Wac
F/3tX7Wmb/Gu78UNDT44mB2ryDvw+ZeezDsI4m6aGp/7w8IY2FTzIRYc0nJ3eUwumBiMDci7aFRC
vo+TJqtgSwDiAtVwCdW/timzv/MOowVXRK6OViQgmoI4JU/e1Zk7nvBaEiHx6fCe1jDmBv0ubyFB
Xnw1m5Iqt0zr06Zn9v63YxEIZ7aPUQ91XaH7+prt+8bxIqaWvqDlb3CvAF0D+1H2dcm9nCQlo/SH
I8DjQxqcUOyWtJ2QsyTiuHVefFwV7BHLFHUNp9e8+b5+1L9hvoCSeDaFkO8goeWVsdxnQol5BBij
NHrQUjFdWI04et5mcFpZARHxS/ZxdUCdze4vgE0sjnrmNGOHMcRJErAV8aZo9JXLg0/RMZGGHLBH
8dsWPf8jXuvguYxY9oltVcIJEKGV4QkLxg5CYSMM5Yt02UxmNgQCMHAQKwRNeYPxNOeYpVnYgxuQ
tMgHLh2FwHm0024R7TpL+tDBJbWrR6YTfb6mdnbw7cIpJRt9XuQqyWoZKveQO8VFEyGRUVcItmPM
oCCbj9Jl3JKL9so0pgAEbcwrAIqTPOD/3vY8MMkO+syY8uR8zb/AsZki0aezb9TLL9P381ul+IIG
mQA38podz2MmlZNHCW3xng0jXLxkPSd6ryXx3qGLlq0V/owR39yPxjdwpAspFFunBm743eoTL4Lu
8pRuLz60DH6vsyxsdQdrn8+KICqvQk9eAckO2c2jDE2ocDxRGqmn1Ay5PEJElo4O/J6dqqDoY9Gg
YEu+g1xHZYX2lXMRUJgyXCHarAuV9aVRFTy/YixPpQKROn/iWVPMpaoRH8Q7ggeDFFxQYhTd9zJD
i6trWa0ScWc+SFiziRoSkoHw3xtW11DdMpCt8+uPqzBl4Xcj62qi6Hw2d98MAGoPdjqoFCY3Upu2
VPM7BGK0FysI966JoyhJCNAt5UjRt6hjL6MxU8f4E3PbUzRz+kTJj7aUT88/n8yw0o17oso8k/Yr
KdH22Jw2NRiDAbuDP4WaXNgooq1MNLEUngwlLool+I4BCqDsv55BKXAKoIWr4N76tz5eSnbUWp0A
AziCaaA/d5+7Qm00wdx9QVrsoCw4PiSzWwfOoCT/xts4+El8Qv9ye3wzUWuIRMNtIW0V+qSSLkOQ
2EoGSN1paYRcI69sKK/9TtydsvAS42/Cur8oC9ElxbGma2e/u7JNwEncSUOIr1/7X+ZkMPhiQKj7
fWsABC6IpWTTkHU8UjGaf6gVmv8Ji0qiLMPJWSioMuOqW2S4076UltkzF8aiss6FAjg4PhIHBfJT
vhR7+sx3qS1Uzn5kSwNPxR12xz99DliFZI2k580l/iEV+OMBVrU4lxPEN8qCWzRyG+V0ID8OXoyB
hXVT6q0Hi8WpqlcFbAHzzaBH/eUAtyEzZuq60yhxYFXUXvpf7RdB+8mDyhKSUn0EaiEG2YxjHoI1
ugkOEazHZjwXQEJDEMEaLuwTGFxwM9rjYzxyu/i1n9kg7eDo5mJ4iqpyVxF1/xKnlSWaoYuLR03Q
aNI88Sbqymf2oYxkhmOUh59Ye7d/QS0a+XtPYueSe1RpubjaDoZcG6UFkmxbLEpDCzgAckHgmAnU
Zs5lwn4pNbiaiuKkVBvdGoaSf8avVq6Uma/nCDk7UoyT7AO3qFQH7fd6t+HvDe4uJJy4tWXbSHNg
6eadT3KsNg+y7H0DNzBGOMKV4XC2/t23apNNM0av9jmwLlRS79oCWL/OffCjr0Zi/NIBhjvttXBY
JPTvFwXH6JLcovFQpgXg3BzV3YOpDBfC3GN7llH70CEUkrdjIgHHktyKebCixM9294vQNpmyDs8s
y+WiszTnVmelJSlGzW+dbm0rzIwXpNIb0CKJTs6rh7osWYCUl2NjFCiYjB5d6HJjkZjodskxuQlZ
FrxXlWkgtM1I0iM1q2TlvC2X8+/NLZ6b+8HxWG2RBGBLwdBAqXws1XEpbYcQ4dwIA4pQd9PqZRH1
/A/9Qjryxr2z9gAV0TyDPomqSi+RxNUa6OX0Z4WrB7URyGigu5E7hx/lriq/BuEZZVk7T/wqEl2h
MtIlC8Nkn6LIHcEvmrX0N8SVWdzw4R7JE0XR6m9uBcqF90BfaQe76Yr/mbkX7zjj6vNQQIwxfxjO
cR4WzOKqNm2nLc26LNtxbuEqBtnprT0Qu9T+64pqWQrFPHoOygXidX5Dh6SJNF3waB+qMEWIa3le
D4nW04a5yq3O/M1Nh/NxZCJn2/9B66u5MFDS7qlh6qZ0H5xD2/CCl5REyNBE9bRH2MGOt4N19qya
NxygL0lGgwrTLwNY81etck+H++eakQjOg8J0HQdgNhGiwnC4v/bgjXvyHcCjhMb1+qdDJlzZGKU7
YLyGimy3duqjhQ9I3+1ecIl6C1wEUzHmaWS33/xJMOTx4eqemZIsQ4CrxbyvXSq14JdDhm6e0e6A
OQqUU95rCa4Fpw5WOAzwUgtoTTn5rjJBgm8W01m+3LD8lyyWIAaBkjoI8frLjtAMIK7P4zL2N6fq
GCpSpaEFmrDb6mBlcOJa6NOaAMpsSOsUzRvXuKYgtGTIjBgdMZY0yZ3yIhv4nHb+BJGqiScssGsm
1/aaezSJyw1vgDFU0hDoaYQ37b73llO/GE9zht4W7XhKdHVdJ8IHHgzDMJXJ8m4nJflL3hRwcTdB
40SGhOnc7a0dx/Yian2FfXuAyDAP2FOFAh382j+niPBIuW0k9kuFRXggEChpxXjXZuyAhAlFZ2Ay
9CVXfiF6kNRGFMV5OeeYMPTtYSixu8Y1zkyb24lerMggaNhG9RYeKcX510Go5WKcOtds3k2yzLaA
n4m5wjYYdxZUeW/CnjTs6W3L+ls2bnKZJp8KvRUzYjnH2syt+W4L5YlMQdAFdR8dT6rExiRTCzh6
HgsdA4YKhzFSXrZnSxWIy3uc+EP2wzkwfJpphAFvTdi9Y1uwvasmzvhJu9tg5DUlocDMkGaU9/tK
3IbfKLmoTuoGB3e9nBzdR5ez2Jld6UNI2rP0Gc/uEJPaXSjAwxPBRL8YRM9TB/P3LWALm02WN7P+
lFAYLBlmGMXhzZ+9UHMKZj4+I6N5MJCqq1Gvn0+2Ru0ZDlpUtVeTuj65YE7+15a269mBH+5DO+N0
qCOMhKwhSamI5v+rlFt/xOXu4eroSxJZ2UOojFhnwoFWbVKyNA4cg+UT65kx9WpniKd6mSJKoR+K
y5dVV+1fLfsY4a46JLhLWeJeZq1IE+SMAaDC8mc6/K6dx1mxqKKJ5YoEFtTWNINFgDD9y2etol0x
uUGNjsX4x7aQy2/nVujBUnn9BzR8hPdGjcOmJiS5kww4UFqFscP/h7ROflh3GJ512nZvo+1kD+L/
Boq8y1nicJ8l69uf+Gb5aTRzULge4/IP55GnPiHkaqt6mguttl3n5qhjoYO+1+UyImTLOcbois8n
DucPOCDnzE0892iod5RIzYNx0WBZpAyoW24t5d+cPCwVWYL7HaISYQe0p8h+XGMkLJkM0oCocoMC
dX9BGhDZ4poX8J+DqQpE9jkf8UMg2zo82VYzWJpfYZt5mL7gUq0m6sPRTx70BwW2kvsib1pNVJY5
7nHbpEpCXCnb3rezZRYYnIIhGh+xf+Her1lZsxrQKTZbEykybe9pnAC0p47xC5sTYltu8kXgMEnu
L7Hn1gXer2yXKJiIXmYWY1ezbeqCfuE8cJUyeChMMKzDE6L3x5IIHIXmFboFWl6nyA3HlO5Va07N
nsgDV2YUbYo2h1pyCBP0AKUWI/umfqnka6ruEggII77XIxfyqN4dop9L9ppvDtDQAOvmf24Xq9NI
bvwAbDBhDxcxRjfT6bDfAfpDKbtwXnqu5aDcst3QJX6wPs/GufubiPAbxZEY/AbMJ5tBwA5czU/V
W9KMFEriyPYEY+zy9DGcqAEVy3njXafn4P2uUU0d4rl60YA+1EqbPhtdcrryUaX2LpIDXOy5LG8O
XF0LJfLhUC+m1vcwR9HCE3qofnbWk+zqWFckHwCLQiALfUqlJw9LjaxjjG3QORauZ1PzhjWnKC49
TtLIhiYz4XYRbAXqv5RuVai8quBMZvIehnZrkIkptP1ErnnBmAj0cVuiyLRj8a0R5xHsc4fScdJt
ZvZ0ueHUnnwWUsvEY7BcV1CB1XfhRMbpoTqsePXu6QADGikycKptwEtZ+SMap/6MrWvE9qZTDety
HfC7N8Yz6xD9XcfrYsfK771jMmy2nMsiRbZ4w+jedk6/HT7QwDhpwZmY7ONs6qZg9UveGO54F9mq
6vMGp18JzTmP99q9gvcgQ1MRg/PPTTPa0+vSSZQFTjj/Ww72P1IGhRy8xbAaNo5kSrkcAdeS8ru+
nmbszjxys8/jIZbiqX81r7vemAOvFVbdqhSPl26ksjxqasWmxSFI7TxtR9WFeahV0475fldq5Ecd
8FeeENXn14SxD0/R7w35By+r0ots92pKSDnlQq9cRqdN3Aucv07xGq8GspAXt+i2AnrqypvdcBKf
L41Vr79ACJS2zMBivUb9IOzAalWVb6KYsWoRqtSSD/2xZF8V3rmekR8dgOvJxV8ye2OmV8nIAhEZ
YGZfScbCYvqVqjbCNLsWvshuvJHR0m5OSte1yFgrwnQYeEKz7XvlnXdSt3at+PUMdp30kpVfD0RN
Fg36Qu2msOuDzO6NQR4DLDK/HBFetztgBDzey9E1A8qWtnaehgvHWX1/aD2DIZCynIe9kUJ8zgUJ
JmOfiZmWYaDN14OfE841WjGiaIGs+DxCeOZVUx/7zV9IO3DdQBky4wEG1qY7wxXyHtLPtxe5qnZl
mm7UEQdICO6duFN04NUtcSW7o57I420Hpv93AyNIKRVAv27K8Yg2h8A6xXZzy9IFFcU8qQO987aZ
erLk5VC2N+2PnNWB1S3SyOjEWEIunmkTyjF7I2/OL619VC6xuZL177d6P2DkbMJFdZd5e4ts6fdc
TrwAtkWZv+hnpG5vfZ2UmJuHN5GQqEz9KmOQ8uOHO7CefPRO3103mVyhgn9C3C6/P/kQfm7MCr55
FBFidvDmulTeAdkGFp5WJfyyds5kygpLrLhxmtSzWGBtsp6K4BZ8ywJyAN5Mm+5PodK9g/8q84Rv
1erHzsTRtIAxbm/3ZrKseSP2MW/zk4FY18SpzbVqSuha8UTZNaUPKnKkMb3CNmdYnT6sMivp4fqa
LBo/UBabveaKL1ctgTqbezXRIeCvrZgVJBHTXFS1ZB0OVKYvzx8bkND8CmpQzDz0SSaBVkdalrwk
bXP7DBP8qrUcAlXDqyOQtdYIqxKqhQqP8/sJ5YNSPTrsOiQr1X78gsC+svU8kt+EFYxIzjIWhVS0
jadilqOfbofWDIKGRMATFEBs4VrjI7O/oO1aAJwqaUW5ib8K2xrgmgj4TOkAQtikiE1ZpXsm0w1c
Tq8PiHpw3P6g7f9QiAiYAAnFEN3mQV0Aob7niDJrwVg1nWfdYB1YRZ1vdQg8plG4EFsc+Lgv5/cv
pz3biH6U2XQfr7IpFD9YVVknDNc4iEPLTselI/bCQY3C7zdjGcYxypHFj6Ngg5huWiHWAXVs5ZuX
WY0rG2hc9i2sILrc6LkL4dxn5RYUH4/sOMCyRYtrpQjqfcbBQ4k2PZKrPnQ5HYhtRnhQfwuDzvWe
37tnN/JDhHtEruFrsX6nAPQXHNhGeK8M07uQjm/yMdipIAUOwLRqbOUThWsqF4M7RhgLnd5/1KuL
NlcC1WxOmGXFdTmJM64YbQfw8BMItvziCIspvkpIOQgmG8XXBiyl2VaHkc/7mhjdOxVRdax9mY4E
/OGy4rAkHIkmdvo1/Acwc5TarOanER6DAbyqG88Y1mtf+pcZCj9UuMLg9FQiud+P6olrMlKTsggh
2dyICsh5LGys3XAB7LXR414iw40T1g3c8idQnUF53n/BU2AUbN39Gfrq6XVyP1bJWVwsXTg9lhf8
2AOAvWrDEQSgF7HeAESxlR5CiPioAZnjO6BLZTV9pY+FnfHWOYRNAqiiVNtUZ+JkhYoHzkS+uUQw
JNkv9pBiBdvvhFmB31G/jh/Ig7kToojPBvjXOkx6cRzLq53MGexTaF2/1lx3ZayxQbTlethxE+vq
QbdE6+aCOhm15911+5X5hMuGHzVYN/EkqKYBsR7by6L+Atk5kldMgzs++g2n/yGrAM54tfnYyy2x
WzeufeP6vNgaQG/IxMA54eiHz4w5PY3wzdhu3fwGe6GdyZIX8EPUpOk+eQbbdBqtzwQDrwszGIyC
47MBB8LduMtgbOIOwi7BtUdYEX9rOdpJ+lXmp0w7zdaktboresJv9bos+togAyMIJdsg4aWy6rfx
2jFLqVadyOSh2bCgwSlBZ2aG9Lv/xQHjL4CWDfBlqUJnZs4qrOLfInm7w3OZ0xuG3yBm1VROBb1K
GPcDOI2GuRY9tdLCE3SjTyz3g8h1Gpl7SV6ak5w1vAghndxSZtpnyV7hgh9ejJmCBQ7reGuNgMTu
nip16BQYpEwsuNyEsIJ3J6vVbt9PYA0N1HMrN48PaamP2w86AIQ/Na40FoCc7pHjqu4B5WnNS5la
WmtyK1frbTVxZDMU6rs7ObflqpSciKiOk1wgGBrIX4yPkl0lwzdE3H/OC1Ozyr+2QYye/W/1Ypa3
ABUgX9HfwsFdjqeKZ4KDcL5OmIMDFRp1HNsH9ukBLLOjdHDPiGsLD7S191eO6WeQP8IGwMTrDBnZ
wuut9iiDn4SKgObz/tr6RoWkYizGsUb49cty18bUlc9OkVRRpw8t+q0L2dbdK0w+j4uY2ZHeciqM
BtE8RzSvQZeqvSUfBEuRnNtDaSJRSq/CFdGA7gU88EUiZUu9ydiSgx8D4IIC/kA0rGcd5pueb08A
uJTym9zmZ6OeTOoVIf6pk6CmAtIBMzfhf9tc4hQ8ES1AQk46NQqgHTEoRfgJe61YtDPqdCUtWemZ
iJCUDNAFKK8rlIbEkz8Ndg+GV+WOCfKx+rafp3oqacJTESn1sWdm1y8xGu3XM7jCnGhM1t5eFZ5x
/ik5Qpo2KCjQgPrwd/jLCiI+PizMbPAZOyA3wP3Cv7WchSbJZPLPXGKF4xzHdI5flaeNNXdqSvPI
4sYShVD2bkDBF4luBIbrjN0I3NvlSyebcLUu+tNk5jdXvOVFfXoDCd7KE2qIpeNAs29EYuOfULzP
z7XDyutmgj1Y9jHg9e4yoe/pNVwr2ixDc3ikqyyfi/2tKLWwyZYA0oOPUHEQSjTWIvRNF0Dqz7rg
cr3ViN+nM5rwRypx9KxpE+oWXGP1qhC/HS1anp9yrCGHIrkQaJWgKHX7dhzvsA/rIp3qLOdJSWFw
aXJk29JrnhYqsgJDV9YhD5W/n3z6tPPCwyIMGIJTpSl2TCv7gHVtEizubAUsb83EbqdEvGzHEwzq
WYC5ThdOWxMQGA0nhnamq7lQct5glA4ItNZZaG9adHSdI7mdJnK8OsDkr/rEHL6POoi6IvUl1+k7
S4miqHbw3AqPGJb+7VZiI7yxOjS6+2SQujOh4i41nR5OLff/K2Qa62isBgB0WyrGYBZ5AcfzO72N
CsTDuQZoNwni3AAxE/6UBQhrn2kYN3xJMM1kY6HGZXrGiY/YIVJhWHZv3DVj6HAW20W/kN2ivwUG
73kkLZYjgFa8K/vngkJtBvYjls7wr5DLYCqAGOyzuY/WOByoRt/oTDchEZBZUodurhBSNjQ3xlXM
hLVdw43KmTJ608OHRKbNtffv0UvlBW7ZGFOmxGgKhBI3iqYzznADI1U+jUgJDLanYabavb0zif/v
Q9+H4RrF8JsGHoZNr++t7igqFAHomGto+AzHjY1jigzyLJHu697vgZD2emHKm/SLc2Qv6ozn2nfi
mj0uEWEJ6FeJ6DEms/SkUF2ziTiZkoxooh0tiHHEDJ1r1K1YD0AdJcw5UVShheoh+HTC9S61g9g4
X9saXHJNClGNMFm8CFQc7hRbFXLun0kVZ1GXGlQTnkkH1WxipXxrQds+IFzbD9NTpUlmzvZM7yLQ
G1DOu9fQpRV0RJl4JG1zW+0UNFZbwNB3e6FIICEOAh8ckoRKizmNJHTsRIFGVVEbs0DoB42KYZuz
KC8QstQEmqeg273aW8IWCHzstWPsvTegmOLiS6kXg2lrQZ05bMKv3+xljy3U4CWwWjz4QonRK/Na
9+FdRRG1OeI7ZPsdzH0Ue8uv7nlH4nLmXss2k8ZZmjwFOplsIYeVO6QV/9aKwwoMR4VPCIU7l50I
dyIobggDUnN1K4ryaBk0Qb5nK5qjmyepo1in0eO9Tgjn6bSGxvAkZURmMQuglW2DbGX6SRps37JO
gAK0t4FPC3PzsMeEdd+h65P93jY9Dji3wT2zOgGEBaPXu5GVbIfVKQyidltICuD4zzFUFvsTgthA
yhc1hNDpYAvtFi7l0RI9qwEe50ZnlNejkj3mLYMr71M5seZgfLvFnxPfrj336ol2i4JoVGvQ7h4F
DbH20UphKHf5/aW5PBaAZaUTL20Nd+QOskHFxP3eznr6j9ENZocxmHiUFDgveIO6794sRiyZuH6P
Q8NiOIHUfYEtf0NMz/XLHtVzO9PGCf0fkBLKZvr7PBwiJiEs+u/oVxpuBd719c1YgN1pc8nPbxeP
8W1RW40fXOtgaTiCuFBi9HvTpLDnk7uT4y910vvH0ARWloLf4NCYIyl1LoeaqIJlf9gzFn/KF54a
l8OEEax1/m3NfIggI3hAhPkePFmYjdtaNbWdvjwcXR6QoQ748h7VTi/qoJAOlxknorG11Pu+NAPY
vNvoFvxVsAd+bmW9pDtDTD1EAeduCeQOf27+s5Amg4zz/FKqd1vXq6QronM4+eH8qmPU5/Q6J0Ah
0CVvjLKqgxzyUyDA3boQ09P91jaxzFOxhWXyEK9YWifLVvKqAIh2JsdX95i7nF0ZwhOUPNMVFGJ7
fCNgy7APtbjF4PWROSup1PQQNbQNA7o/ZW5lwSkssTPnB66wm/ZQS13BSjpgD5PTKKlohaOAIF/8
oR7dDv9WVCBLkvQZoyFWG0TyvccbkkDU9vA++hvecLgkAj8hVyWXsCwovggXFBiZeO6/LDo+9aJu
K6uE7FoFurmOGWe+KM2MoYQSrbI+Y51UwBt3St09xcFOeQmeEBUTnNXo/k4Jpqby/BA1ZJ6uFJwj
Y8kODUIgCe6//uOolrO6aP1Ll+fkRcvHWqk1RAOwz1Pv5UvzVE6mk3Y40yU7Xuvn7tvnSHsFG4KL
1zt6iJ/awvaSxogCfiJnUQ4kfnzP1c9qUs1HlZPCsPEH9AvW68iiPVl00W2D7ZOZ6jhgiWXVqDxV
s9+wCQee0KbtgqO94sa7JdTTLqtiw1qAdbSB5Mtu8e193iMu9kfziiwdE7OQ6qCwDznZkUEGq0be
tTXjMALvBjn1dG8lsPCPsjADBvbHjWlH3QEyUDhVUcJugXq09gFUG5rNBHAV/sfL8EFaSOK9/fHJ
RleVOrUcohrhggVb5J6BmIeuxGBEKVtvUyLl0kLgnu4UPF/Awrkt0cmzEUER8PHMXz/p9KdUjP+Y
Bz9a6f+wo63oVPe7r4Aojk7N2Vw8PuBI2kfNwCeW3j02zn5boMLUy73UO+8RtWQdSlhW6LqDZzsw
jxG8IsF+1g2afK2VGVIYeArI/S6WS2UjoVKFuoCKM/HsPYG+z63ny0JYKGz5CEW3WQUU2YHQO1rG
3sB+PYpc/PiAGaoDeCrxuoVq9XDfkS/LgNnuvGuDveWfcdIpDug5RVUsEYhHVrbCuXatXordPtGP
jsOjR2oho2pw+dE3/PfIF53PlmOoF+ryZWItCM3ei0YSvPpI/z8w/IcFjvTvXnb5azWsAD0i9bf2
BBvLA9l5hPlQUUnrR6PK4j0+3X0T+m98PFuxubE6O3QNy5hDhbEmWEznL3mkVp2bQ5THTWnHlqwr
phJsCDz2S5cZ4Tx6vAMbjCmPDkthO4y4+iJWYSc/BYfbnyFThmR4rS42hKlIViz4G/2sy/hDz6u7
g3ckKxap/azuffIMKdqIAhsW7WF5FopGNqZZE0ZZEUYdaZNQzOuUEKL9cOUp2xgCPtf92bCym8rX
xS/tX+DoTr2704lsLqU7OFtPb97IndpqVHd3Y99dU0fZP2OClTXvPAJGL52iD0wcWygax6tTDW4v
vNM3TWcp4CPQY+1mzouIb0N+g27D8ln5qWKsPfzDWlZa7dvKusl5R/hO+R2B1ULAUTpuAQNptQk4
+JW0fjzXKqFV0VGNBUCEU9uX3Lcf+YsSWM6sOKtil0LM/rax1ZYqi5lLEUcAcpQOpMfq3p11IugD
TcIExRFLHYIeRQiK6DgQDcOICjzLr5S6zKpSmmx9YJMN4PpGbxxK/ZZwJHwRIRGFipiJ6ua0zsIo
nGfVdjD94ymzi47uLwHugiR53JGDhvOjxmOaRu5FkNTOQV08aVZdjECzJAGzLk7FoJskU6kTi24h
OMOY7YSHpwMIkrJ4ayHx9PrWw0lfKn58WuYUWix9glczSRk07SBwaQvQaCZFl1r1yMK+n1DVWNNF
dIAPcHwQQ61OBOmehwWgIOW34p/r32MX4R5RJZAKwXEnWUTxPzKV6ZvMYKFUJI7xwttQY3lpDv3j
ZgomVxG7No3SRckD2cLN5n6osg5fLIFAgerJ3FHrgniSdy7D5h2eA9wEtpPth6cgVJiy0DJPEDN4
Q9Vn9ldN3AvcN4GOcWdEExmPNIN9fvLF/yO0Ct9tGw+e5osnW1MC2a3nZylJXoajrYkndWVXB4yy
ThokYj+Y6bHMT0px/Cbq7W/0habyojMoo4ernEP+94ReaRvpKK9veOvv1snaPShk8BawYH73exto
Y7kfpUDiew8SILUx//Modi63NX8IMWF/FmVAw+DGX8D9tBajduOaPsN0EAZ9DRpOXq27CzkiG9aR
xBZOoSZeaWsz2ALtSo8SORwzyCSeRflNShDDGHh90xXp3fuxwassS8MI2fm/b5t+lK6rf4vDIOX0
61bjzZWSPjJf3s51CVQ1npctaGnzevG+OE65a8UBBrXYEkY4Z0wQls8m72KCApa5EBzFdO8oZi3D
cZSAufP8J+MKuyzZeGMKpnWiAU1yaHrLjXrzZtFQkhrJnm8hybLXFrIUy8Z6+HTH4YVjkUgjy2do
trX5cerp+SVJAkdIOfPCaeU/RE24k0DTbCzHm5TOCbMPFfe608OH1cqkFJVp4F/d5Sw+u3mGj0lY
S5owsfx2NX7qPla1QjC75zNW7nl7PRz1hG/1CuhqgXWWybzBcAtXBsyyJMyMboyTgiBNXXir+5wx
GEWT/x3MyxY1n7imotKtKAsifxDJTgHMapy9qP+2nUo8E8fT02JppZ4APjIeeSzW744rRB5euISW
Ji0og0aZFHf20xAklADEpUd1fiuuiAzH2zQoStntyeTU89P3otfpykXi4SpkH86L6XsP/Ggvftyu
BhOD0V5Z2l8lNZ4ksDw24UtfTb+VgT0E+koZppAeSx2XKi4tPYQwYaQZVYKnJdYnzM0IbpqeZklI
JZZ4/H+fDEs3Ullv7RGxICbJUu7fGMtSV7VsF9Tud/McgE4bYd5aaiQtIkizc+U3c8MEEUmxWD4w
cE+Trs/ARSr/Wr/3WoIEewa7+a3Gi+rQbFC2bD/aJzJ7XMzhy9E202RkZh/LTAAsbjXQRyr9ANMp
Zv+ISgvv9CuZ606mws75CobiRNBBo0CaS+Ee+7mGEXR0dtjyqr4Oms8V1lJK7zov4BP7Vv5QZ4DN
U/oNDgD0cWI01+E2MjDjX41f03/xIjfqy8CxwWd7QkIjH80VAM2izPLFaF1ZN35nLFsKXf/4H0ka
74sHyj/i22siiPKpPfwfHzVjZvDzTfat4HurvyLg5byYBpdwMaJFf0cFuk4MVfuZL+FPfF/9s2Yh
/+ukbmurEZaPqlYv0dS73wo+80KbrtqhbeXeySfvffXEY0WcK3VMkM8HwWfVKTIB74NY/S0HkWHy
Zm/sD7ln9/PYWZc86aWctQaXcDNLAV1J1IZVb8TMsY6N8bgBQXsqLm/e/N5R+wZsCCUdy0xLuB0Z
vtelL3Pqw6PFTK/pfjY8hg5S1kP8HpGGzQDexjPKdWuVjrEE5griGuORNMjSHELnph+nhQIovjav
UQSLb3mJTEEb/zvpcQb1wzaxmHtjrRgoZE7YYvHUxuN01x4ZAYU2IOxUFjF0dKAU3ctphnGWvcjK
qYOeWltltfqhVCTC6NIVDR4MPduuUdQQYLV0lFKO/YNYwL4WCGjfwFfzdVCEIwp+Tvab/QQobg7N
XiJQLxCIQlLUaOpcbPrsYXZTtUX4khtea6sK3GG+6PgR0jHBvNManZSYilbmrLQLNIw73x7JSYu6
+Mps4LTnfsOgp9QFU6hcvHoO6SbRVYVMjOAewURR8moXosEd1vTSLB6dNH7qUK+J8UGiORMRR9AL
WH83bnpT1fUUmTfBDzeecYOteoN8QB/4nUPPlGvJEG660CnnfTsPbBGBXLvvobxf64EWLQ6tDNKL
cMnRnTk59cyEid1c1VZN1ANwdQU9gACu3HbhwUfiHRSCyoIGBTCTeV2BG0YMn95qBaHgnYgRjt1y
08hOi7yoDe4WoI1Gz0DslxrrGLHnuxSu+4XQ56eW9khzJNVeLXOcXMac4msM5WvRDrtdq6BC6lxO
g/DZTF93k+Z/sTbGaFCSJpWZUPJ48MJXX70qV9vZ5x6UPK8KvIPLAflpG/tLWTr4voiVjELPqNlk
sqCqkL7djTju29qD0lD54qiyMOvaqXiIpr0qyIlHzUiTBs3qaMqaFxQ+mv/iNrEyoXGRkM11u/KQ
wXF70+lRhiybjN7aCDm4Xi5kjtDxWfQTmgxcglvOhR5safaT9/cy/xNjDNpgtUNrvDS7epwx4Vm2
2wWPYrxeZDWygkoXrFTlMfzRULm7+D0l3Y1mlWnTGKWYKWyftZqG54uJMiYd0h11rkbvT1W5j8dK
htZfRhz7jhIbt0kkwdfKHk0pEn5zbt4jWNIbXJKxuDsweHIj3fMzVkRFxULx8RyZBhfLFgr3XKO5
fkUa+PufNSrNyc/hZXaJ8C8KRjHl5M03B4XW0nwVyL/BsKePf04enaBqy+LxbypgzeHgiNUYL5tl
B3qvCzOSVs/MmXZSLo3fzY6+VJi/HRUJdn6Nhywz8WK12AQzuo/Cb/qIr4KdLVJ7zuNOkQpenDtw
XRIrG5io1MS/w3klR9OSXJQdOg07vwT9caD87gFph1/Nl0HtoUoX1w4YjrQB6tFmMLG/fB/aUZiF
f0bIBZluQE212TiALUf4KJgXY8aViiHuKdQM656kQII/SsyG1J0x1PqUYTFQt3XFVea2n/ilcdXT
TZA8FYTO5j1w49I3fJBEr/6rVHpojujaHp4qMIFp2KjYC1J1TQz/5uVzVFDydMWPCpOwlAkx8YSl
ZFvIVf3KKrv2wMtTwAEVaJRyNE5FULVwkTKeKZAAE5F9M2sk/jVzjUSgbw6nIG0il9eTqnyI0plF
qlvEzu447kBxhLQeIuLWWkvIIjNEaZOqTSMlZCWdHQ5J/MfMZZKmW6/CSZ/ZZKzAQJZ3DbHWtZdB
C6PCcUu3nEivkcZ+UPpS9dPscFefMYqtaQx5Y56cUV+zUrA6KutgSvAgeOIjVxuuRZLVln+ZcefT
tOLXRY6ABts0lMS/y9V3zozIH6ldiFuh12hSTzz6PxWUo8xwKKSWGkFRZ3xHtaG9F+LErITTPBon
c9aGKOF7Ch2aCTxcGyNv9Cq0NN+eI3mqgF/CKL3JjADrjlRZMShq7r77WZ7SCMS1PhKc2QhVv642
LWmeVNxjA1jrGaggoECubwDtdGa5K1ytLPBHv1HDtKb2NEMq666+lQFr0FZ1UETKroxpK9erYxMB
NMo0ms0YORpFtSjOtNznh7LgADY7FYVqXH3N6cwFUReA67HVLWPuXYMrO5YxB3mbX39glKKumz3W
bnh3GVY0LFPETG6qEHoBAWhRUWby8sLXum6lMJiNrngmqy5/3HBTHze3prxky5+MtmTgav4Yz948
MQXSkHJQia2Dsv9G83EMtdo8qZkp2b6RNo9lAVK3Zbf/kAWaYEhrMjF+MTmiS+tYeK4NVXERYZTt
7lGEveiKDRUYcC0Rvmq9NCicJZIof2rz2JBRKMkFaJkddG4j4Iuxy6n9sebPynlAgqoRT5x+VZDT
d3QyrVFepWTNZzuw3K99RRIW1N6u//VFMk5yM3LPWnAXvxrr/jldBEguKPSwOEP4AZ1cLUxPyAuN
ECt4fKmuE3Q+i1mk0cSJNdWGoywSONxs44DkUdC1DIStNDje4xY4GeZc9QVOCIdnue88bupHQptn
+bbUW1ws9CkAnFGgjUm/BKK3VdItn1VP55DymWi85ActmoOz4OzWfN31u0DfYFCmyvCk3rUa50ZD
lWA3Yq2ZholY0ZMRfo6I3ExAjjvrfGxiILNTgvXYeIATPpo4SHjb40Kv2EmUw/FeqOd/SOr8S/GA
Y0Zx5Hwr2cADPzUYKuLnrbI9ctnIO9et1RIYP3qiMJhdReHpV/berT1vscQJ5pcD85yNpiau9h9R
db86nt/ANTbAOIv2R2rH0pqOmGc9Fh9bqW/vG1iSXaOw9b1JeY1rofAQGz2Zef9Y4jHX700rw98a
W93vc1SV7fS+8oL2MVBKNaFL4z1Zg7kUO85oPqGnyeJ2pyPKcAi0eTKDdT9XKGb6iUOWCB+wjJTY
ujO/DcJ0pBcZHkmVlLAEAHhc6Ue/Wwzx5oswBfxFlm8o2ue/DxhyH1BYLWQI+erWBwY6QH8IhWgp
rj0Da4RuqGL3rLAIjrgEsAw1m54YEg2zHh0KR+msHVkc1a/VLE1XFtFv8OGzhIXd7RizdVCLsBIr
7io/wDwFnmEtMUa0O79X4yR9ySeBffhKPAA0I17NK8K3wq7KJ/ic9sUv28z66yoBej53ZUekwWug
heC4WfUeU2PpGlKi+MaxfHAUatCnfxN6bibnnP1P/ohWh+IDtOxiWaUaFzyWEm605IAn7bo5DcjQ
0wenNbT7Se674bNZL/dK85KTcHqaimi2F9Jk3x1vMFIdyX52pHOYELrFwK3FpGd+i4Bkm6u6kSdR
FD3FZHHyZKBeZduBISx6SMUx3Z2+MxZazttZEAk2WeMJX/h6mniy4s3u8JyU7buurOa76dRDuMJJ
YAI0Q5YUO+EPK5yaGbp4dy+WF/w9VUL3SRv/SH46i1yMP9xjd3nC8HjBdnryv/zQzXtnpy8MXSjE
4uOJw8wjKzSkdG+ceXRVbTDnZYmyIcG8GK+0MAHfsVFLT6y7w8MCmYxSkqNG95iqoL1WSYs5FyCT
NOfNryQmmuoP/3ACMRoIij3F0jp+CAMmydU06LJZjSRsOl/Mfu0uYYBYGwM+TY96Cr8bXwOEQmlp
QqXEWKbwomgChCGdtqnmvs2s/egpTENTk4LV02D8yfuZwWfmzn1EaoGpd1qnVpAhB5BUCKriKLH/
Lpte+BpzdrFQSok8mJyh2zXLVdCo89rX0fDjNHP+IcgSyoUegPR8bDk0R4tACB7o+uRq+oNtsbhY
qzX8htNPO53TmwTqpl7+XEPNm7iGWKVt9GV90nWhxX1OjvNjO9jpMA9kItRNN/gSbRMWJY6tjsY6
BgWWKUDjwkttg8/KtqEUAyg03zWIO0CiGA9EGAx38zyd6wwPAPDDRiNJGKbhWEZQUfUJ/EvLsx+1
LvjXnCK8g9IDEArwSey+4cgCIDWHyQd/sVUa5MqpfFiXPOBbJgoTolkhbjobcIVvB8w3O/NjWzdS
FXGfxelZxT8N2XAh93hZKGn2k2WHTIO7T/HIV8G1jbGFg06JZpO31O+9+oyVBgA2gjsINz8wjbr/
6XHmVhOyeunwkeojy+VG9v9I07T3FLsKIkTRUuApKGLwkTpGoiBT2BK+3D2UE1bm1C/GIieakgHI
kVOhPqITKG6qU28li3YYf/UIgIRkji+7XOcOGitxwgi7AvEaSfZVpNVtcED+/BX66zHNthY3ch8b
THb97RofoqFnRYYjuh2+hncdTC7V5mGrIO1wwaUfj+QFbl3b8zgFpAX5YEnm2H6Xhi8k5brbDjU5
tDX4sqtzFPEgmRbFyXseUL5rJ9wja89ZDUXdWUwXmxKm8zqN33wfMjP2pbT29s9QGeJnLs8ZPmN/
kLNkdKNqw8xA+BLcjXVEJdaVMWn6r0ivu+xKardgqXqbTX1tCIMzG/CY5+xVyD38qS5jaaoGA3Vq
K9R1O+cWermzG8wrEs3GarYqRPBlml5tVcTNueQL5P0WghUqLn1oqRkRmnk4zRQKN9meVLSpuE7j
/og3PbGjJT8fJ5Oo3HeHbJW1OkGrZcJ+tMGVjLpFkCpgNwHUTTJBlhyaXBh23aS6oX99SUw6KiaX
Sc0VhctxdnroPeU60Jh+qnpT8J7QnpXhrbPGjk4Dd5++QLVufGqi2KjhT/JlmHp40wADFT6Lq791
aDyBVZ68K2d1fa9eE75rjIIYtnx1Ki9ASlfAWfjjaCwJmyNshxbz1Tl1Pc+xf8qd/RUbN/sbU30j
K6Hw89XZXa8e2f38ce24CKKlvglNc+afzDvjiZdXgxPZuwu5Q4RilvbE76S8xHXEbjLqWJzLLz24
rzD7+JVGpbTym4guuZuCl4c3Bt+iHd2GWlHOXR1olfoYY3KpOTuD+gp9ZXatue9UXPM05GJyIIuM
tD+tRvUd+qbh/oapI4m/d7dg8aA5ATtHuzt2pUyhHHWEsem3m/S0OlwJwA2VoOMWkM4C4tsiU2zQ
9OL96LSjFt5e40sksPYOTvH4DGofjwSCRTh4Mvn+bPEz2dwoBS9buXtzIdI1zdtjAY9dSA9R9OiU
+f5jQrIRIGmjyCdbDAV0hSqfV8FQV+hivS7k6Gu9+W0c816k8pGKM8ijjF9x0PCjdtt7F5nVshR2
9EzSQxLZqRn4CNo0wDSxguaox5KcBRiSmjmAKo0Qq3do350Vhj4UQId9AYB+X1ZHBCBJWEHheF/P
5Tbgj1Uhm1NnOPg0+tltgZ65B4B5NXZC5lq9H7LaIp4XAdijITMdsth7btBMNseUzkM2Czxlybsl
IgqRxsqqME5WyFsLHrxlOHUFjyeqmUgcm0Uwi/7SHkcnex6sU6FAk+ffkizKKjIB/2J5oOvCxsgV
/T8rNfTE6hwb7z8iG9TjBJLwIoxCZPku7wef2fiaHhWh5EaukeW9MvAtJy5FDijkOwIJxl4T35Xe
gGZpvGojuawFMGchxpLANzLU5+AgNUBcTB3SjjftUZYOwmW9RxemhV4CFYyqPK4CZzLBd50GlleJ
tqMAAGSfhDkQbttnS7JTRHCYx8dNkdSpBVw1G+lDk+YtvJMK6HzD1qryjmR1bl+7WaJEZZZedPrg
Fq3xCzJi6A8xLDja6fxN2vwtKfiT2+VnKHxcUSm0etUDPJZpOyORswCKHQErCeeAJ7S9G9YqOa66
zIM4RZGwDpy2LXIKImk4e+NQpitNVSRtI3VIRM+savj/nujJQ6zH6WnsFbO0ELTg6N4h5uN79708
HjfotPiNBCmQxuGBvQxT2EX+yi5YNo66kJa30TrtiN2mlT+hi6PsY6zJRqmEOhhKUWIZ06JNfrk8
8OXMQX0oUuwbzwvzCss6xzhlfAGx4DSCpG5eF5Ik9MbBcycoL3tePUyaI9tuCfBOpch1fQtgWmUW
a0vy0jEVBhZwN7afMaxN414V25d8UF46yGIJk00uI1cXxJ6UGWCnNFZi6cmzC76I+X/d5FsSgg/n
vPyhDNXcdc0FyrrtVZs3ht7m18UrUH0eYFHlMdo83sLWUn6jPeV6ZAjQPZkjNsOWPj50JRFEatFI
Gbftho9M8uLTHCIt+BuMPQXJk2tNBe70ap4+iYtMjPzFoOrIfZ+lrjrXtO032iU0sxohyBLmVNGJ
th+q2uANCssQBAfQSOXOEjPEx3shAalqxHvNTblAzE4pVkBtLV9B0cEyXE40US2h+NUd7UvmKHBu
IjmxyfDJINrmrlzv9VOJ0MHgwnq6VhqDbFEQVRM5vYlgJKElsrDiDqwW5D2sybrJ002eJKs4yfYq
YmACqZNMSRX/oI/IFSnXuwL+UNBwKzA92ODlEd6cHJWTPfxPJch/rjqzscfnX2WAD5ctMyYLJ+Vy
5xAqiNe1tkElrR2okgr43qzWwwXUBLes2+crN/H1HSH/Rdk7TKJ0FoA3PCbU7hLep0KUiP2oTi44
krbmCWQl3cGrTda2NlQlw4EfjcrlREycAz6cnUDzb20ijvywdFubj3a3QI5iMcFDHxLrU4HqEnMF
KqHMV5RLup9m07TEaVJPU9LB9oJ7pq1PsYsof3tw6HggW44kZbquO4rzfABpir9FGNL3vF+RoOcv
1FXcxVlDl0IZqirJbCrf//YJopx4C5FTzapfyOWQgD8dtb1ACS0SiocfBtD6dKYqmGtkdW1D45f5
e54PTddhr6ZDazkL93ygUOlh2IdMTHZSHafmEDcai1hNGawuLCxfIUJPEnUiggq4sRZ12kFUUMBS
E1y+Kirppb2N8z9icJBDAzWRzAOGQuHiq0O71m/hDqXi4q8Al56nUYVu/lNAPGYKyWqu6QTNbZMI
02pfoFaEyGjXg5gztl5dL+z0xRxxHwt+JNijBbWgeJlDZbERIVT+83UlYKaci+dGboTCDOR9TfuA
6KXBMz4tKucIYS1qJ4lDQ4E2F6B2XY7v5HcUfhYUQkgCPTlRKrKww0ElEVIlT6Q9/HLn/NtKvg2Y
OgJbIdlefm8fFO0qAK6iq0GhCymJuBKt7da1OhfMj8Ff/IrET6Gsms6W3kfs6eS+YrCi+wiNJx/2
oRPC4USoZ+/Xxfkw8lUTutrYCWaTjpNSmBmzTrVLfxoM0FWwi7UsctoKXsCGwrpXJPTuGFN9lZ7S
Q9YuZobICqGXiWWk4hyG46ggItsiLp7whPnC1w9Km5xRkOe/sAkabkW1+Hy0IVrL8LM85/6LXvfp
v0J7MFlZ2msNf7ycW4xOdo+LWkv86GT9JiOmtj8eBHPpQO1XQSRmtrItHuj5HI44wrpVT0fQEoRo
h7Mk9JMbd3rUDRckBxoydEyOhER3aqwV8i5hIjzUcbjuY14Nnw4WiQG/Q78vmjrMq9Z/uEW49Cqm
wd89aHXHMqtNx1HIserKLk8ZYToFMmHBv9MAGYcEtwOD8L8IS4lY5Dz/lVofpY86fiiEn/EL5/o9
zzEpRlLcRVWepp3j7/l/XsMjiAyE14gl4NPZ+CU8b7qssN2HgJJWLR2nrkN2iXowX3cZzQrqy77T
D+fI2xPCxK+oZPFXqGgbew74S8ZFwrsRFbM3qWIltMRh370H/pLBIkYID4JVB7ZFrnsW8bfByHBf
pwXG9O24LUKlFizksPHfulGkFt8TVT1F7VC3SOfzRO2LgDnaHFfls7cUw5HAD0e0u+xhBssRYBpM
XjgWIoE0PGe2yVZSEe3HMPoRKqK1aPkvacqyh9/5Z9Ox59GhKHaXqZ28hDwBWlcybE/075R/mMnL
p1/7h3J5855vogIzw+4u5VlHrSwZEuNHfia0oc/XJJtICMcpcXY5sy+upBPad+d0L8ZZ32izT6rf
FYJYYKvupRynbhpFV1eftSQa81WskYou8NKi9PpB8bfZkXKhrVb1LBww5tiudN8UdBb0TR/feBfA
/IU914shvl0ej3lQF66skSXq0q5qFe/D/k7r95mUHY7LFtSCWgKwkC3d0doSHLWBIwdhMU4WRmZB
9IZKyytvrzy45VdbENWTFR/XC59VjH4e44oqpBbkpxUbrYHWNCZsYqchYIrrqfEHbjopqs3teFgJ
5t0ZHTl/Nqul651Q8QftBxnLNXnE+5cdF+3/H0mP08HNHoIKpYp576LaOpFJQrztcZinxw0UjwyE
JGwBtfL1CP1+nhDNMUFgyP5jejQ8PcNp7XaWKnHwMh8BGBOFC+IVFElj9Z1YLYDZS/RIvsujOylz
7UqRjYZjqDd4lildTePgeO6baTQBRzE9QeDNAEsA1DeD03KUcEq8PHRFpUOE4CNanA+DCAg+Q2XC
uWFQg4IvWTUg7laB/wRe+VBhaD9MToQHg/7IJV0c7pbrPLUHmY0CjgJbkWuzjzZvNjo8rTxu/UIl
4qUA395day6VrSCpqN6HnDmAbfjwPuPc1fAcDpgoR2hqN40ZRBuTq8A3+T+1qVUKe6leJHLMBoAT
+pVH8xOkQzWCMg5MAPY7aSqdxFO1XWUGoDpgO6kzEGanbTRdX6xfbWydYxm8+XbD2InZZ3bodpsz
cie1bmqUbQvhfh61xP/Co15bu04TRUG/FAZnB4KsTpuNdZMbFQh018hrPQIbAzH/iAabsUnyCfOE
NdLYXsWkUYaSbWruGAyzLfRt/c75kk6ITXl+O6kq0f3uwNavu5odSR5VJ8W2wY27tf6l8ekUcAjO
t6n4uAbo+HWHC/hVa3u9vw5dofHLpMnH7IypLiTTD6F63x1sPbztFMMI9H2r83rd5epcl6m+yB1T
yOSose0T3gI3cFuaIVJcuQPNWQ85EEO8wwLo0ZPi0c5ByLVb2RQSNS2e9uUMVbzzUsSd+EO0NBxF
TnQ+joVwRgbW31EGKwc2VToOphk61n+olxxEf8cnGtMI02OxjF94ogul7T0qWBE1vXfV09jVkc63
Am3RMIyLhENmeyEEAFNuRvI7/jCqwJokEcaRsvaZXrXgiRs2i+qtuVTbsnJihW3o+ysi6+hlcNVn
2yma+FlMmxYcmp2mQQE3r28L2i5jb1kkBE5L1VXdw3+xIBhqUFCUDaHSmlYR+GnpaNQuJ4Mbm92n
X99srshbzN3aDby6XVc24OSX2A2QZ4OBOneyaF/brmyQS00BkjHpb58CCEidAJSZJl/uMme/crf2
5zrjCYXo5ORg7C9efYovoGy6TJeSuCxxvEQ4YPYiiH4tbNM5hbjQftuR0vyDrtWpPgBeQFEn4n9b
vnOCv7NbJLGWl4WxqnHXXWv74D4NeBAD4vB6WTubrU22GpsUD9DkFzIzpXJIKcU1YKpPbfyuv1/q
T5Dq5tlMvEM/iW/xANXugOM/iSzH13Tcm4nxWrd1GzBmXtVS54pd4EwfR6W21lm9B3dKWKVynkOB
2XVPvfz+Jqm/VyIR3jrcxlmEoFolLxwgGw5AOAOsg1rsPvJ4uzCI07Mbimvu91mBqPOb0LH3poyk
wQaYVFJP4aK3jKTs63XYDjw21bD/kO+OcXEhhAFq1tvnE/Z4pIEuVJNFKIxG2bWx+O2hr4FvVKgg
D8yzK3inBmWj99LPC30HgcSlIb6nU9ctYNtzOLcVpyA/mM7eubh3zqZMO+ir02fXeODIZcYAMaOv
OMI8me6Cvokb1Hoxvwy45ERmhfp8hYRiQHPPyr4TGCzIVZ8aCzt8FIYdpmN4MgvmnUgyxoC9Zanf
5ah12mCy8g1jvKVpY7AOcIOgcGMAc+ru0a8esxtbQ/K36bRo8LxgkmPSKNG2bFk8Mf44s4IG0MFf
BejpRfsAQVC8OtA8vY/h0U478FjzJrb+CVpXbjGlgLMJyxZ9eTyIjdZpuaoHn1i+P3ehomz18e8/
MMjRFdaL6GgW9sudkxHE/9KYSGW+rYAqTv7bXH1MfS9ja0LWR94j4AegKTRM1esL7Sn5EKgG3AsU
uQzJlmPlILqiNvSQzKZd53wlnnFhV2Dk2Y3C/3HjtQ9qsSHDn/JfnAyyRkxIXGNkVYANQYJ+WAGq
UaANMndKDk3OZ+fViPE43zNASDutCpv5N5N34zRfIJe0VJaAdUZ8uNCyG60GtGhR35lLIzoJDmZD
qmJi4LpcN4i+QpPsvz1idt9Roxdi89XRdYcfyugH8w6HLoNjOI0P32jsh6ELnK9B4Y9aLr7PB/ox
sZxJqJy9JtKWn4akSkjBQmh+l2nt+tpltJNaEYFJCiKnhbxfmfBJ1hZ1BUYu+Ts8JCmcP7u1EQC8
K/xvFTDdgacd+5olEqqVJCi4iywOde6SxanfXpMOzETGmidmdznrcRYtQ69YL64hAsMuDmE0bYCL
v2pqkghJOFN7WXj157C9K8c1sLbs6f6YhPKGj0KFopoeMOHcYsasbUfypAszt1Xw/OByhEKUNSxH
TcG6JfWDoGltQoion9atjESVK9Hu4fGZ2kDNZKFQ4c3nK95V0p+/qJnShCosiFW4OlMn1/lvnVEX
lfGL1jhmzByJxtgCruKey5Fq/H3ViaI5B1GsjBxZQS51AihfgA1/7ht/xyC9PGR5WMFZ2p7WtnzI
v8EbZAI8uZ21aDloYF0Em53Qpma2/yT+rNo1u3+7jNn/YCP1fKshFk0CKFsaio1pm9NYvR4ic0qx
sMFyXjmjfPFC5c6qyuVIsQ439HKCgNyUjvkYWgMhDLFBubMCMrRpZz/XGwP6KsL0Tz/6waUah+ce
/XWT9+lSf271ua80ac/kAakgx328rN8goqJWF1gQPVIAPDA0Qzxus43Zl7vJurHC/Bv+OeVri5Pq
OhxjZBYXAj09dmWxTUKdDJyaYgykoDdh3NfLl9oZm5GXheuu5sd9V65mq84qrE9MS0L37G9n5zZI
hSgty0hyotmRU3QAKkjGrcHVe8auZGsa5AnNs94+twSPZ5x4zhxclbpEoaGOixmC6btNRH5nM2bd
tZ4Mn+D0JoeyqtixT4Z+YG6iumhOd8Vl/nt+AwSwK/sqrhbeZEUiObId+PGwnQ9AcQz5F63uM9fl
9oBOyIh2ceAkLrK6F4L6WQs4lmOZP4Nj5ciNSp9mvC4pG6mQBCHuh5CzLArgOzHrgYR7GTPBwIz4
6LQJCbLKTW++Sj6+mMzXq5Bh4/JE+J/I1DtC7Je30oqAOIY/8wYEeQJCuO22y9Fcx4hCuSFkD0aH
MqB9y/+blsAABCIbXpxgehVlUhP49Rleuj0roCbBr/ZGBZ0lL7LlAsVEjV+1qnhAN5rkIqvbuM8C
6eT/fQWMjpc5xTByC8nLHI4GLQ6WtB22PFLN/ir9B5LVVaosmqXIxTXmAR7vuS2cnxjJw7iPvgnp
oFdqqsB1jLHrEci5upVnltnp81FC88vTiqVbEyEf5ziLC7zfI214n1gsuwa5aLaf1W9w65S7z1IX
Yw+aF5LJKvAJ2gDB83v809Vja2RaF+M41lzzmhsB+MNJzxJ7OrjEASOL8Y61jl2xQsRSnQiA+YxW
auNOWoG3K/7j9g41u5gprGeFUOMA5/1MRFLToe0x7fOmKlco1KW5Juts1tmtgNiOmshVMlQClygM
smeM0UORKFh48GFAvkkQEMV/XFkP2B5/B0cwGTwZcjXZ4BP9ypzNedyfXBJJCYiK2vtj4kj29OjC
9HI25YC2N8TED+6tTIGlJW15Pk6VbTZ+biSAwZzoaO6NQUUpPSA04/XFWAi9GwNSZI5iQ/toNkSw
aVWrd27iprH9G5BhrZneaRGdVm8DfeeL8sFlhgV9gSZLjFGNHUiT+igNQuYXi3htNQAWf3awRCDH
JUKw+XKNZxjsyWNGAgIWkJZwLAMp14yna5Jrg/JBUEYqwM8t6Hf7f+6HmE0zMyLdaokz78WW1ItD
ZAWBdsT9V1+d7sQHbLnVTBTUbCBCEFN8fvjLaGDBPr7InlJpriUBR2TESgmNUzWeVTMW18Vefn3+
cM8UfyABR9e1RNa33Vs13L9IlWzWKXzXs6z41ZiOY+z2sNC7mWgW2F4KD/w8Uglmbf1clEqoQrvh
FT7/AF9ShOnsKBz//t8+hXnlqI5ITqcot+U1+FzDQsnvwO2TAXXubZW2+QcobBFF72mRDMXw5iHi
QQCVWHLdqVTH991+i2lQJ0iTVCf4iZy/O7sYriYredyP5+0/TExHatKhEPuTvpJ9i0bnTuHjL2KX
lX5IFNJ4m2oMZSuiEzv4n5WoUDAZkbUI6mqUwQVYydHPF0yX405CdeyBWPs7LRGui0ot/J1BOQ5A
OeWvgSb58ctDKQviOeiHE8BnCLWaKNmkvOVxb83HE5ipRfh/BaeIDDkl+mxjfB4Ql+RY7eOBsAto
NxHei3exBz6C8xCSD3Q98YpGF6GkpT2wL1xWLHt9LyTJaBnDZjDpZJEtzgLE10KGn3bWRtAvYSsl
no55hWuuvjMpddRE+1XrfEMKe5iNtdsX6guDZ9GnBu71u9CbQZDuc3CQ6JUh5A2d8+9qeGyL7sRv
t3AhtId0LZgENzVvCuPf2mvtSX+hpYiBqDaDqP1VGU+6G1ZDKBdepebZp1Qt8XBxZlD9TFzAdJCB
BqbUBV+U24sKKhte7BfoK3gxwgMhyewMewLrjGLFB1N8VFUTxSUhDXB9VgNbPAn+EZUA+Hv42pyk
lIYOkjIcPa9qWdr7TedWa7AYIILq1PboVgNe5qAaAU3hckl6mbX3Pc9Yx8LZDkFfomIvLzXgrxoR
ssrwX4MS5VZ9K8Cb8peCNDagsu0kG8GRD/zK9teokEirSp4SmdhgsAp9lwzeVbfJkR446Lf0XFqo
YMcLdqi1Bbe4kLr+4ypFS575kc6o7tDCVefxEXfJDiWmLZY2YZbS79SzrGoVIT4N4CbgrHU8wUNB
fBO80dYiH0vQ7M6RiPIM3liu96ElApIvcssectixpYovOb97T3W8F4MqfzDPQyxHKqrqZMzABBUy
rmmCjdCna013/w68LQCyj+gkGt1PIZlZQ/l60EZvfhsQDvIQhClhiA/rxmXl5Yn52msPK2BuPKN0
/A39HfYIEBp7WGWZJHEvw31zMA0uNJaSmlb1b0khujWneXsBfZS/B/wa+ucwzYTcaPk8BhiWU+Cb
sinPToxvH83h33zgyT3qDMySD/e1Qucfuw9R9v67BO2wF7E9NmJxdCrnXyhz3xeQGtfBh9CpNPXb
9Il/OjurTuZhKqeyivCLLnVB6Zct7kqdiIaq5WijtRdHh9TPZ0IMaFRELudChlnkw2+8jKiEDdMc
LJqxHc+JWCPKn3Fn4i9ue/oll7O/lMldUVaByxQ7hPyjCEcf403o4sbZjuGnhDkrt9jx1jb5aUUw
N7Z2NnJy4QdjnY0goPLth42Oou+moKAGM+rLUlXvriMinIabrZV8q53ftVfOJ/DPPdiQqiPRA8C2
ujABZuSSKP71c8EQPa2fG2TLUq43SdxrcxvKEvmBWJ5uZUNQCPG/J/2nZndKCAhdkFkJfjRWGkJv
6Drw05lYqbSwqXB8K2ITyMOkwPFcFvDT/ieEIkkTK8UGJ3JBMl64YnzQNEJwn0d/a9gNnSF73BcK
41TZ7K40I1EouwYQUu2Gvap+kZr43Aw3nnIvXF/sJNcUMLjhpayuxsOyaoAnTc2XUnXa1xZ+kocq
B2RznKB665DVOCbMr2ptzXY1DPsBKayi6MVHiERgWOBwkVquS/nOVR5k2aJbKwC1mkF5V/1ZdTOz
V84KPkhRoR6a8eBr+ql9GIE5LZegAwucbBGI963+eORHbgPVznjTVt5yJpluhmwRUBoCWjjaSopJ
BpjRQFcS0gQiJc6xfbWihMJygeLQWdaUVTJIYtMl772M65VYdNdGQhJ7/sW9jmlhs7aAgwS6Jqid
MHpXyj3IOFq0AghT/+fgCWTh/bFiYSwh6Lo2efpPaY9VveeWFYgJuEcfeU9I3XncV/AcKlBrZWuW
7uSJxztM9rdqKQ3ppv17/utsbYF0oHv0zsH7JidGCNUO2ESUHBx0ahQ19AbQg3MkOFddTGcaicJP
QtuX7HtkY9l0NJ3wJJ1Uo6nOsR0J5I43sIfh0tlIx3rniS/hLj0xJjGZNYy+kBRnrPvm6x4lPaO7
i3250zh7VtpjpIkR58f95XxvWPCTl/7DBkA9+M+9DTnY8kqSEq8mW5TD1sUvqdJwHKrEKzUdIhg3
FLMwfLg/cw++LHHBFolWLbCSHDX4RwFfdscVP7qlQdZB+3u7AyMsqJreNSkSyRZNYHT4VWsv9dem
Yt87Tbpxic+BQniuc8UIEzSHW5yM76PD3rGi8xorNR5ZByWKHc3xQx1s3o8sbzbSZC34RGBOndAj
hfZ6xpYv7UMBJuu2kSUq7fqTlWmB6FO8YOxW9asrS13gz99KN2yTonOihy0nHoQ7pN9qDPm7VKnO
24QvGRt1KTae7i0leVwEvNQrRblaTQgChkI1+c8++6jGKnsUpY61J5eb+oD8inOQuw7Dpnv1Ah9F
SEsgFr8HLUfBLx4q9NDfZbwGviNqL1sAXZosi1gN/YkoXE98YARBS/F82y2Nwn2kIl8wQZSy7m4P
2PUaAq483f7kYTo1hrRuQT7tUirORy6osjSHWlvUMcTspm9vmb4sgwFI0OxUTj8ku9h3l1V7tVEJ
ur6Tfe+45HZ50Se0WXBUXr24fwgu+VFXir2tPuSvLEghrSJb9WbRn6sdp3xFf1h0TNWTkZ1VlUwy
dXXyxqVlm/WSEFlTiZfc4yt4thGJuIAvW6b1swNyftpdWxA5x4M3+/Q5/Vas2ziHoVLuv174zbpn
9krItuk2UGUZ0XWg/gSQuIwyjrSboqFPi8BquztmnYeYI4EFgl5yMA6yP08toINtwDEsIcergQyE
1tY+CHir0eNuJaICaY618h5sPW1knVDPkG4BzOPMVjyZQ0SXYU2Q5INioiuY0DpWAuQP2ImtgqkD
cC6tvN3TM1mfZhq6Gnv1g14/bAqUy0oO1fNZ98cpJQpd0GNMSLLpOIbHDhnws7vYsamhLuqQbKwD
nd2eD+Sm2eB7et7Wmq7fKIUonexmRBaHvaGov607Y3sM1WFHPEqSGGCFQ1eX/zv6B3Q27sdf083p
8L8RkedYegFZbM2R0Z78xJEnqG5WACJ/KRzGb/NTqQyFLXjWc+ZqQde8x2KTiRsAX/EieqUNfCwD
2AlqyIaYKeN3gRHn0owFhAhbsfpYQjTzUY2TpRa5GOOPcAs/lF++oT2685c5ipbS4fArTGvM4idV
LlyiV4VyJgcdgQLTjbAEysx4ryZsz1O3KPsIQapfkdPTWwvaztpd0MA+/xVLKJ6aRCOX4a4Ncfvx
meNSfpnKXz2oB+2AxliJ2Jzc8/jD6sbD7713sgTwDElytdcAvzfkMsNnYZ0dTOPwEvtun14P9oHB
Lvzda8Cc+T6aifSCA9F3ppmhu/gNbpu2cXMS5ToaWohnPxMBrSLNFmGtJLjdguFpWYxUsc3xCRVl
nmiLir8GdHSmnfq7TELqODMUKDgYFTxH4qwALydh/T9xzCrTXgTVnD/CBFKlhTcXNbZDZxpXc/qW
dpWK6G3RVLbcWToQgr208cEAyhChUXYaY7GqQexyjGYa3psMH4GrVYjDTodJkUDjlMPRagj4lMVB
lwGXIR6UdyEEg5j8ZmCySUJTLfPLkdaXMemu3wMTXHpz7ZhXweEyUdRzr6osY1241xIrdRYcuOQn
MYnqPAsG3CT6wTMLvxlHDTBioNg3KbIKmQ82kctGFH0bCvl42sbTrmLKoGxw+drnmzkjVIc/NiC3
uJxWHjk01OrYNu1p4m6HQI+cGvFmOsNU/ViF5b8JKQm7Cktwh+qBAAtXGA9toM9gq0gNY8m1RrKO
vrGFdVWTNhTOq5N7/G9NqVd7pqTCIAfSSG7699j/ivIqJ0xlilPf4fpFOYZQQP1crrHDVGI9HZck
vUe5P+3wiRs1YOYdzrdx/ZywENq2jEafnY7mVET4iGCQj/r5V16KPjBdPPyUBPUQEJzkzbVNQn9l
F3rnClW2xj7dbObgcbhDmjFrui2RngOhZ58SaPHJiYTg7mqiKm9DVJv1OkbPYH14n0IWMAdgtjIK
CPV+eQ8WJVSB2za6n9MBUa9ZXkKqbe7ZOLHbxKbILEY1FvbGkJu4N4cyYY9daUZHEU2LMYzydHaG
grVNyfjd8/wsLS+lbZigv5K4ZVPyV9kNlwRUMG2jb0tB2w5DX5HWJvzDNCWl/S28sC2n4KUpMZzS
JkyNxlNvOurPUqgQglkjYuhDlyc7v/yp4KA5VuithqZTy9CGzGYOPOgDMBF1Zsju3pqfl7H79tf5
4Fz3BQCCmWftVjoD2TMJu9UHHlezUnp7KYVGsaw271Z9HPHRtKnBzAbom57gFys1+mJsEVm42NbG
ZiBfbrS2CCOpZfWGWBC8MMX+WhUpdpbx7I6bzMf7cokrhBDM4XkyyXFVPvrGeJStLI/COruOmtgT
/RhNSPnc4GsHsB4M4nE0PO83lgfSPDjf8nBDidraWOpMIW5NiW8Hre4Wc1PjDIO8T9NzQZGRb67D
7X0+NinvVyxjyLbzKQP2TXopSO9mUsbi5KMFonFU0rupwZVhEm1AfFaGwDW9n29s88raeyfNsstz
vJFSQrRwYl3F7VqsZ739fhR/0BrtNQqsoyvEmokj97iGXL8zDKBgIuZiPCjoy1wTXlYzlqTR7iMj
IZ4KqiLMN3GcRnBdmqYOdLDwkdSJIbw00q9fPEgqCad0lDs4SD4dg0XR2vbD0B3k/jiKPnQEjs7g
VyvjLCqv5fzgWJxRon2JaVVGWbKqa3bUf/4+yU34cyohM5JuAIrkcu26ZhjPyEI3/o4Tjwxc0hmy
I+hXR/yva5+uSdv5gj7f9WpfTAifRkKUD1IO0ADRsccE50k1MTWCuLaiDJdQuiODF4LutXNvPuaU
BFPvelNpDThaQjHrd4o4qKqLYeAf3nIMk4c3fyHMMg651V3CnicwhBlmWFftf19SvrTddVQMWHCP
HEBRi+Rhzl9tWzwsX3CDy3aHBxxnqXMMI1JOFVTlGWMtd9HG7jXOTy5u09wrdr331s0GRs/4kAhC
A516xBxdYtj4YEDCnCsW5c8PwqSXr6d2l77J8CscFk7RND3qdqfSWtGjhQ8CwIcvrecQhWxGht38
dmVUMOWjG7f1wCnknM/jaCoVOuqps42J5R83BE3ye2HTCbEI0uypAF7IwL95GkFPOgKB3g6YACO1
2Mo5Gtf38tFh+zyQfQFOVfiBMLucYCdzUGB9LdUlD8cN4+pm0I0FHr3kioubOjYPXRuPo5v6bl7Q
/ad6vjtDuHTSE/PO/q69QFzIaUvCNUmh5KGQuvuUJxjnPQspzBlPOou+gSn64DTqThuz87elyyU2
bkUibW/0Cm8aLJSZ943IZlWRiTrBGcv42Foo6ktWdEzZ1SLHCZkVpXiTShNbui7FLR9wfQAAiF2H
6XVzAI3bwJ3ik5hMxbcbdVr4F38pAPkQeENfTho1Klz75zu0IXLR1o4amZ19P71xiz3rOVTnZDHH
EAhzXseMrVBPN359StGzkHKYGpE2FEnUD02pGGDj3QHbA/M8O0qbTI/trhsHE3IKIyE72sKTENXt
R8nkK7zR26Vq3LfCEiUnfXgM770MW9tGNwT/i9YyoOHuOn0x8SUex/aQ9s1GvNx51cDEeQpNWCPJ
qbQ4rhxyuCAMhlidxQ4UfA/xfd3F/4CJI5Ox1QBFhhPLmVTYj1Uwve7LVnUG7gciTiQdLFs3Thtw
/s+yes6RmrVTuGPJULMojLVz2Mrc3X1ORYD1u4W0fm6MTaDw+eKpJMZ1CigoydP0i89axp3IW2Wh
KYtnyugHMAU7Rfd3ckj/u+8pnr2+FtwGVyG95FuIik/xgSQ5iShOREFP0LQKddj1OEyoMtn58gjj
iw9F1bIh+/tMbD/bd9CFGJk+vk5aV0ZgydHJrWqMkGGEp+UANx+i14azs4idS4SSvyd85wC0x+Lw
FAw/VUSsenCp54BDEGvBYTysk9bfDZ9rh0wfc7khDGlwFjiRGdGmBmKVqdN6TG3u94qioYQXcmuq
yahvzJztcc1RbZChztZgk4B2eSNgmTt14bIuUpF3AQH063N7dS/XWvjFbaecHQrVfFzFApw0TpDc
20SJmv7Yd2YTQ66EtGjgdl1fOKYX4DvIKytuqIUiepKxxksU8OjAYpMjOkZmifEnbtRg0UyaEbHU
ENT3ir8HXBg7zn67Ksej3pbS7r+VmTzVOklsAwFanr1OVkeMcBwveROEHQvv9n1qOX9ggDId2Ooh
PeYKbjczhWEj7t7Ij9R3PnDXZBVDRCIoucwD+2+9gPlOXcyXjrW9fJTy3JxZ8LVXtrCPC6RHfPar
XBMKfF0fy22tJALjEdgWSO5klaMsXq7pW5kh8bTK/wzVmNFpjSrKWQqMFUfrLI8qcO7xqcia2+9W
DuHjQwEGoO0d/td/HmJZv3f0FDZcVCRXhSX0uQkLsVO04PRkU1M6sW31AXC5+m51QnKYQkgCjVKT
UlJx8QoDhraiJL7YmEncfywTcQ2SNpPrG7VMaF3hkAjKKfRxi28+v/Eyn+wwwJPyl7+07eJ0CEP8
0WhACbt+3Qrg+eP3tSe+a53dJH4TUuOeMwJvGp9d04p2wJESLK4gjQklXDEdLjk7EnKJ5Aw5P0BQ
6+nywVy8uKuuNvk8UUl13RSwFJsKakGLofVMGyWF5Bju5h2/6jO5go+gYyGv1+MhrgpVx7Nu1A9a
lQNy0igcBSTO7XnxEuLfcmToGCfAyvEXP7i4EZ6EhX4p1Z5+820cLauBQOm1YirhTLZnxE6DunEO
fSSUJsuJbh1hOuN+ADER2RVZgHOEfb2LgcCNNAgEW3PmjLsDq2xftcBmFL/H+2xrjI7kDkrsOQXb
J7eKREq+02I+VRT17rKA7TBTrDwWh+peF/qMaFyah2opf0RkvBx9RllT/joQe2KuH2Q5zrQeGN8P
0NeSzVBWMiBO44LZdZSRGZ1mH2EsyzwPwAobPEettznODB5b8Ifpup0clOhxxBF4dkhi+SWPXe+U
qSGRBMZJFhgMr7oPiJUfXITVxTKkHB4HXgXaTVjvJB6kHtoVvZxrYkVs/82DdfNpOsQVpfSxUGQg
R4DFzpKJBHulTgLSnFcEH1RW4gkc+ZzRQ8nqYLG4H/aFBSRDkqPTs0/Kx27CygHAE3qdjsC7UuXn
mblQvUVuGVz/N9rHpLoGV/Q99ekz/FSlbCjbGWAYXT/+SXYzVAWfym9VpI3cyM+QE7LKTk+BJ5oh
5IG5mj73SsJ4IZksa8XMrkJwTpbIfMeuqPUeyZZ4TbyoKuaUdsSpT0p59oJl+tujjt6eh4iG14IB
LSmHkKIGEGByu1Da+GsZX1zfluD1EMh2421UqoMmHT0vogfeA6NygXsozYTTOe0vThPyhEC5lWZH
M/WjAKT2hpKA4Sq/4dislwgE5AKRxDO1aG7n+2ywnyymoSsiJBFFBttyXphy6hyL4oCTkpmQgH8c
HI8TP1/ZFQ7TrYxDwOl1AAsAHejIyBzVoMY+73DtYqGaKobadzQh6J77lodFXqrkx/wl4+A/r/2W
uIfSlsXL4j/onfb3Vnflu3zbRfj4eyu/osKtFb4LiO8L6lxZPNPi/F+4uCZsHNNzuehKv/S/eB1b
eMnOmdzyRzBRKoF5f1owGoV6RGPtfHzZMbq/KpEYdOciuFNWpbqPt5JL+UlIp/Xv+nJjO+rOIPH0
/mkuTmGNDsTrenzt41Awrq0xC0MPSQiD/gVB3koaYKBGhJUYNwWSd96LDRYvLDgfR1hKa57LHIXB
dx47bEIfRYDGb/+3knayDsuPoTI/TpZ+oz2k4UfG+xVZ36LUhyhpQ1/HksDgsLMUKPMKoMlCYzV1
z65lADpXAbU+H2lXKgaindDXUpNp4pLLy6AXlpwQU2bObqhADnXy0C5r+sI1tgLP1uRkrkz2TZ4z
QqrjrFGaFGgN6d9EGxHt9NFnPje5DbvBkgvO2wzd2/9qrzt+fTlP8wDGBOZldkeWZgJHNojCCYDD
fmI9TdtnWj/oJApmpxt+jXgtukhDa46WApJsRHLVoUphxWur0fWkAeeUNrFZgaFvOBzkQ+B4zUXN
XBUNU9AYK3ySZicdLCp0k85I3aMGpxD9Zp/0BCJ6bnhDCimL5JYmywVidFjoUs2b5Cyy5htY4dWf
iC067zdsBdeZTTWHDyYzbc91UITSn+/QRpPzJtGL7mw09te3KMu1YgMEuMXqG6EiXZsLvB4hARA6
ukTcyfAHjA6NYUSMLE133ZQhXfI4lUBdPO5WasXbFOOA+nEX8zydIx3qVxsXdquhSk4NaOMhWKCI
Wd8QHcby9XLYRk4M2W2DILyK3Tbc/VGu+b38q7H6WYDhbIpdO0rmS1F9qRIP92r7GbuPmssftrqR
hwKazz2N/LF2T2Qbg32YfXRULXzAWITpin6v5QjaT9UQBvo1P+q9RdlQYFNq1anPQjfWHKTihM57
Ji/wxso/bxDeXo7diBTwbvS0mNoK8H0tWuMaQdqXSUx0D1JOXwgXNbRT16aQBrqKNTI7yNaG3+aK
/eLlizGu5JpcdUhbZhd6lLMYuiIC2nVGOZWPgaAoteUwD+us9uDaXwaj/wbgHHM+3Og0W6wijGgC
qD4su76r3AEC6z++PJnTmFppwWnRG2RLmRHdpD8Vrs75VN+2pbTuVy8UkC92usPCEFOD1uGjjNp8
AyJgj9i595LXQUrJKghp5BsK9ktu53aqGSLj6rsmzQfvOG8kfH9Q1z+r0GZgH1+wTTOYShpxjodT
jLhVaSRZUxt3AaVKy7oP3JSiX25Gu5PeYehJY2yZiAZX9recRZD7f1PXVEKRaIgG/rm/Kx194xhp
kOO48nt9SGT30lDswDx9eeYKponSZ8Bqnw8+CbBd1s9D1pE9e0X4Ipg2oK07lFaj9d7afDFyPY+K
/0H8y4TpBHBZS2uJUUG8FKEUQu7nkXirch9U/s0G/x30FCzcCcXesj+Tmg5T3iYeG22bY0cE9l1M
c1NWekwlMoen6BlgA4jYUZQgF8OQvos7pX+E1Kh0A4pac+ibaEX6x/fcwu3pZHtZ5xlRiEWabbMx
896VWVUHqLHSRIww4nEPuqXnJ6V7K1bzZzKAdHz3eZA4CGmchEjc+3aX5qRRHZn83SBiGvB8chDC
YUvyGX9GbsuQVB+89AWgfwsInucHn2o/zzNCQkKqPluqbPm0mfvr/sDTw7/g1w16OBaG1ZkurQvo
zzo7YXWr37mwaRvi1XAwIfn2nc61PEPTuqwtEz9O+8/b1hKbIFb7DhbB+3mTykIYsUIx4B2xX1LF
PJbK1T6+ADEAQcuA/dkOhOfFKV8XhFVuA6KxaFnb5WbeutMb9pmrBIIZ3+N42uA3O+oR1BN9/Esq
incz+HfoJ3/sCeOA3SJLsUC6BkPZqdnaVf7580Rpa7mxMkaNZzO9sncu01L7Xmjwu/LGoIW6r4zY
AIviWhHtyPBt1gX8k9wsE/UH/0ssKWLUmW6Ddi84HYcFIADv1YAq7+bRCYyZPQvoqRdlpkIPl/X3
C9zJLC9K+jK+w0sEZj6zmGKtbwuB2zqrDDR60LW2bVXNaosePlUfutLkkFEgb8VNKnACteHjizS3
vMQXNqBf41DQ5XhlXvlX3l4Sclp/HH6IDICyftINO/qoQG5UTuZvBvX5sce5zvL12V4QWCw4nELC
q5/mvvOFZNP0V63kgwAcGf4osi6gBA3XMgZbMb/zOMD7uHzqi88Jb4CCmmNEfgvmAbPXEv51/Q8G
RGRQiNE3wQOa0q7Lt/cWx/pesFcoSUYt2nvNAm56BFmDPmVQnzE8kvspdLYpmfjmH8ZNMITU3V6h
PHnq4j6s99CrRyiJlokO9wbac+RjVWYODp1w+5PM+LmoKrLFaM3Dc70H39wPYmIiteSPtbcaxvgZ
r7gC6My/KxdwWzLaRR+6aN8z/aNUmbqZ2PvACuzyY0pJWl0ts7TG5BZtzDPsX5oC4kVil8ObVIjs
Qk60F/6OUcIZYcwKNs8z7P06dt1J3CvBf1u9MjrtD6f582d/16opOMvnbvEXEnh4OUWgbNSG7kJv
Trl9EDpz1yjlW/5RX7Xh9NQWIo7s5ws8JwrPi6Hx9pBAHB4ZwkxC0EUpuGs0pLP3k7WwDaThwbsN
MRsoa2mMaGeJLuPsUUDDE4pbEul9QuMO1PMzuGtn8iT4gl4Maxix66jLqDpDiuFGCnhJzxlzRy7u
oK0O/SyY5NaRD2cnkMio0DtJD338fvKgdvEp8Sxxco/2jq6ZAdvbWFnQ5qvxOaYHsPwnSFzSrgZU
8+P+ILq96xKTOEKy4f6DSUWNnII79pa4f7laGCZ+Y2j8P7LUVEBs2R1PKn8Wi7qpHQreYgP/Vnll
mdestluM0wsoeihNyO+x9/60mj4eESyAr6OW9+qVfDKBZr87ZM9WSOBXfkVZcQwc3ou562gW9Twq
xTYRBn9FG8gyFVe0DnyUZeD/8qInsF94OWO8lt9XpNpxtdASBk1UDUzaz9jQyYcUQ2CQbFv+Hu5z
rEhF6WWaY0aRxZg5c8/DunDzM/vOlCKC7g6bpx0F0nwUKe1VM6/WbSg/nCJOrpuUEZztyV5edK78
UYbvV3hqhCL5Zn6ZsQdHkKltJOTJmGJvhU1F1O6dpsnW1+OSOeBtqbsLHQ5C++Fb5tnyJdVslHGF
N/bQlhiEBwlVC9G3peKhrphXhUlUSRWxmtfkvNHYgx5pVd3bEY+JAp4Ban+sVBvopwE7/KJ/3hUI
X8EYEPGXF+Yc5Ah9ppYuCvvajzXLfOFYP5YgpF+ZOEfifUGmXgvxWgpQgFrbyks82oSbhqs613o5
yMzRHpyHb2kwkCcRhHqCBo/zgdsieD1xV82WO+m3Rlya0+Xu4v7S/Ra0yc5s5WHottUc7WPo6KIU
vO1wAmHJja9qetIOY6fZyQOFzc5QKgT0oUllZUG26sE0/QYzxr5mi3VAikzSlKeTYRm/o6c0Iot1
yA8CziRbjZAU0A+5/CU5HBuEslvCbuxDafeuVLR5xL6jDWXRXaM7Kh+p8jWrwatGP/6P+cTYWY/C
YVlao/xAhizzQJZhRMjn8XqnPSDK1Lf8Oubt+pymJNroliNOeUifIiAU1W6UimNF9RR5e35RBv0c
fD1nW4C48vvX8xf0TZt/wAx/W/Myz75KVVam1ji+fR8DXmnZl6+7TTOCqICnd0BOCgpdk/C4uz56
IrkrZsgCX0qtH57GtYu1aZG+Z9Xp0gWEzqZFQIQgZD6057D2B9UVPmkNdDEd6yUngLKpCQgiNerr
PlRAwHdxWMHZ+XKP4xla6Eqp62VC+1tpnNiBAU1c98dTK/4KacJYMPT5aOIAYauuwXJhOsebzApp
Ohbu56AwVJ9t1fK0x/qppUawzIHxHUAl8vhMs1MPy9gw9NDVtKamdz7dClCN8J29jexmrxmy2Ckt
9NP9oh4ytN6lgAR+CJkCr8w0Aa6zDDN7z7NA8PFII9AtH1DZO8QqMQSXv/WDut3r26TBmmT6rcwr
z3hjZn/7u9TUp81j2dGxQDMegYTKyJ7ZhStVv8CnV812On3mN8LEWxsp4qBLZFszPNv0o9RLuJOd
KXW0BD6BUVvYlcYKioI26x+X0TG0F38+i+8qJL0QJSx5UiXNUH74RuWmSoGiWksrJCAcw7u0GN4G
QJRc2Mmrvu6aNf1T6mYzl82VS3HtUUwhNLZvE2K4FYkaUcLXsIc53RRfAkF7UvOoAY8gPeYk7MXE
+yeC6mAN7qvMgQJ3UwB0T1VwMeMyoSppEsboN+FFHIjkCZ3RYa/fMbNW7cchHgagHnVa5lZegy71
ETvk4yIheYofrjxUPoP/zYMU/U34nC/CslyPGVpDChQopFW8kUlaoGLqNLJKfFa7O7Ahh2zzwwZP
rauN2pNZ+XoXAOeM7x4ABkxzvlQ8T3xpM50oDKMteed7Ejd7gMOqw2/dzL4jqMxViKnoLkAtTDZs
jHFmtjBhqAWtXbSyVmbg2nMoq0PyHpuyf5b2FSAKME4nbMRZt1XADFsQpjST69y7oZ4wwFNtV7dj
OsPkdxDU7ykuiMp95E33OXndY1iwi5PNQcocn4GXDQ3Sst6K5Jy1Rk6PBPwxj9xCf04ateaCtCGM
zn5Lg9RLRK/pwVZRd6p5yaQsY3xh3GmCIE+gkmc9zgefbGlEleVHPNcaklEzu5r95n0sZf/NArjy
oNDqYr4XB9kcYwSXSuOJr8A/wnG+uq3Gqiejh7tnU69giWHl198fcWbtYNwZzTj12I6XLOdQAFxi
YtWVwbKU/Ek/7Jj9pToNM8gZ3/Vrzz4rcR340ocAPx8437m03kuq+SfoQm/+s1d/glc5R99NgGHk
EmIWr5L2jS+A/+T3SimO8Jj1cOXeB9h7Xbrn2dxbP/JckkC9niwIbaIrs7uJQRiX/lvbywP9Z+re
5CGQvnXwDYtR5LO5ouT6KZX6r1IKhb94mxHfoULD5J15GPE/vYRU5nwlnB3J1iO/bjdEOTOPVg2M
diqfMq1z/RUpFs/nLHRN4C0ETisVvTHay/f6NUJ/txrwi5PL+QJOxD9kujPUJC+CC22H/6NbR/Zr
FEukUaaEk7zk+HauL4enPnpszsKkaDIqU8nqnbxG7SwrCk+kZOnplmmfTDU1b1fFV8dVTxeLPLbS
jCXwftKiaM9/4PcnR+lXv9PP5SOefca21CkLL6Q9/rZCkcL5r9gObXU8zVKtoMwAl66ycMrH1tdu
xIBECwtAkeUeaMSMqbnD5j82qeGShzbgSlCUyOoTvzZmafc3YlNM026ruK9379B+ptPQrGuq6WNm
l/t7QjJxH50psVFfl+xQ1Oyj3won9MbAznIQRu3aZ7r1oR/GWd92m9MAmDIsClnQa1nB4mquc+xl
uiWlMS6zp2UJl4Ayml8DLA2brzmhbSWKu9FNjBqJA1abycahRiwKqaHyolvJB1/6RVBrtmmRMCJg
07ccWUp6bN1x9ZLi6TgXTu1pPsnW6+LCd9mTnm69/U/4T6cFfQRHmI4L7BSrOSBY1ah3Md40jE2o
DVmW55+wSkYB4wdVCqKUhfIBL6nuIfGW9DMAAyUh8J7iKHvJPwDbQ4XEqFYw9KNyy1TCdJzIIc3d
VNdLkxrJqhfm9iF5c2ZKi2XGFigNfxG0eBIFWZXSoUUw0N/dS+L+iAshI57bcmjpmRKViJVk88SF
rbY0KwOi3Mik75NWFDGzQJa479NXI5H1dD+uKvSLjCSht4mKzY2mWwxXaPP1h99oFlzsGbQllDmX
FnaoHBWp+tuQpLy9gYDRVia/CSXaY7VDp2a8eh5jsTcWWFR8hH2Ee8VuyQ8GUIg0w6V1o+Oi/0Pe
wfsDYnc/iWsRKOSj/3ldxKR2WC8EeRa28VEGnu+VC2l7LGEXmCmwJdqtx97xPJRVDLDpTqxJfwvn
/SFIfSarhWacru7VT0HvpbdUrnEM2JGfKMPVxy8NsQQ3MZqTyhrNtAbjaHl4GV/PqSRgiG4xCD2b
vSAwOKzv1EWa6Qp3SKWNt+GxnjcO540czCS4ry5Ge8kR6kUE6uPAWDGY6LHC19ypLaWPG/r7F+NT
+hllTnUu+aXWtk4DrzcZskdC6igl9/ANAQKurtFLHF4Ft0pD1zlKA2uFMvljzYPLAMkSgga16EKL
0V9Ey4zBEOsLspru3DkapaRsPU/iybqbhkwo3jMm8sieK15XlPJqt2VLUKeJOojNdqIAtItZoRJh
f44+nTcUXjPpOBagLg1JJOe8H1RAdvLd8WuU6wcqn3uHiH+4iRcXu9mmKHuWCNoO89Q1YRDTtFV7
ME+crs2h2PcsK71LHijPzfeyaPiHQffObkUWjN1rQlzSd4d+9HfHp/9UMI7eaHXUiPkJopn8oLUy
hH2V5cg72q5XKgeHeOGn4LfnwZi5ke+2PXsFWkm+MGQdhbLr/GXZ0CwBLqgf0u+Ox5ni/mDDLvEV
+bwEX/0H9WoiO1RTC0SSNE+9FFtsq2bgwlfk/Yp42PwQTH/gJoZNEM+jZF/J6fEpMGXrqXFYJrgk
5nLjHoAdtvsFXrNUbYI2yB86bSfXrxnTmNewBaZce0bAtij7zGKKML8ewc+ZigMy1Hpwlp9PUXL7
zlKlEJZS4xiC9AnposYHCXUpL8Xi69j5JwyH7mPGZCaVK1gagUR8z1f9lOeQQrgJZ17WGnMZr0nX
k5U5UUIwf6YIj94igsErITWqudpYyLcqjaOUxiRSOLktQip+czv6hDUd2np3GjqRrYdJx4X0APtD
LXwIBwCo4/7lFGSoPgJPJCjm4nMJEWPf7hvTOFgoiqRMJ2GH7t92vg7IghKiElfVTqZt9lbSoEjG
phitteXB9MQvQt6uB0bQOj7Pdcx4PaqasqzcmuiaGiyxy8QAUMiBP1wF/hjrYXYaf06/gYEjuWdQ
ajkWEzSF9mspzb7f62iWZ9aunFgJFScRmxxS+DISsn3uwU+2zWSAUU8pRQd94e00E24ts16Q67ss
8r2z3f+KjPdN7Vd+qWkHbEopWV/A/xAfDY4Xw3KBiAw8++2czlygbGaj5nZ1e/PB4hw5FO1x0n4Y
inUzWDcsQHa2zChGdt+474BXQidp3IKpZPPj3qk+PThinOmFWp8LLfCeHwOOsvw7jt/qVKXJyCfy
oUYgBHyc4WZDyqleJnKvTmH1IO/hVDCZs09ST59MIg+EJ5fvNj8a2eHhAueWM1uEeJ8+DyVXn+Ax
PWP7jrO//RSL380XWDt4Lxfn7oyO2kyEenZLDg49Nik3MrKnOkCQft9Pwg1zMNJck5n7+5+GcQrK
56OWBL2O2wJFrM2dG8Y+TtchmVFGdDAFJTPWVApZLP8WDLZXgu9JMOmT10zgyEKXalNmgReZgXbG
QcJH59CKWxi6anieJtM8zmotVQs8RXHZ3Q+hG9egpZzEqHVYkQaWBwIq73AdktHZY7JK/NQ0FZo0
jLp7CxaymRcpjJtpD2Hn7Z8eSkkmkQx4lIlKefHSexs9CZmxi1pQeECTs8c0I/PdvATRDR3iWZe3
HLj8nD5S3f8hPXHP65p/Wtk+RWmxMzhZa1xz8tt5sxB5Y3A6wqSSnOVqsG8c42rZGB+3E8a8GY7U
4LJSw2QianCrRWrnaGJRQJkiPEx8CAp2CzizsOLmbx0SjHXhDUPXt/K4acdrd08zkuFBn/JVRwQ5
dwdKymJzpu/iKapQPNzNvd8iyyzKTy+0UJyrgcQwBDVs+CpCdZM0jb7KaCa4XbPaIn7N+LqhxECx
b6dMCpuKg1GqAzPNFODUjGblYuB3tEheyCTUPea68tPk0HkE+VNpwfoPdzr6km2IIWCX5qRAcOxd
TKu+g0dzl3vHNa5Xb1VL3hYC200N9r5zKiYzm/YeRj77zbsYadkjMCcyNds6Z8fO0lmaP/RdKdKJ
hCfKTXPTOw+NZV9uJPHFj5uKh+UTruK9+WKaNYVl2A/gNSnCoZpSQCr2cVM54mFZeIxGfrGosruY
0OYrcv2TQ5SmFoQjRa06ci4wzsdSXK46JvgO49F3tvsvgnE60zKot7Cjc/oNtTKp8CiZOn9yanXb
Hcf5dPQQzLB6AGtS0sVd7n2yGjBZJY3Ioe18Dlc5SdoDVuTnRtQ7tqTvVOgBWy+DhzsKuTzWB0v6
7pegO+c5LmAg3EH6bMu/jyAbE9mYUrDnjzAw7E1DveyZ9jQ5iAiv8lNmWsH6h346rYV+3yy+dGv2
WU4dSEuNeEWANn5US7y1CTdO2WAGVcSMMe7dKtnDGDVnIV4VJ6ewtDjJuoRToYsj2pTDOgM9vvCS
AfTyJWK9M8ZuQSgGY8Hs4bW3zIwJRY22cens+I3AFe1/keuFoc08ioBHIYULSh6FEGxYSiAw6Grn
t3P5vjXTt7A5W9Qk8cpUKvMolSd2Nxo/eK1n+dplMPl6JVbLfIk7kAjxtz3Q1mtlVIXM0z7/Tj3C
Btg8aaDDzZS0WSTPqd4hm03WAhZFF03DVUB6dbTG+KuqWShCBJhlVuVvIZcsZ3cAKSp57lozeZ6Y
JfLIGZuOf+gELcSS4NpCEXDcEjZF0i4Fvivq3/wxWBqOl7Nk5GwaJGTKWQ11fhjxHzGgvAQYrAk0
Pu63y9Y6ImPfbp1SOdJxpTt9LnzgdNTn/DeX4qLyJdNhHxVYArB9Lf2VjQmeupijeii9Vjhu13NL
5/xTG3lAvBw0mZH2hu1NKJIhqjOnVn3yH+jLRRNFiWbz2TSt/WWeLMrED358R3YY8zbauer5SCRl
YSvc+5XlrPThUxLZpxMz5x28wvPCGf5oNyt8t8J2xob9d+gDhyg1DCp0vJhFZKg8q5It/oxVnzSD
Hut6aKFThHJsom/h1Xwk5A2f9aXDQOU9WOU00gWlH766tnzbf9xdP8Z0h8M6xBuvO0/ky8ON6RD5
Div9mvLSvdXMl5Zs7UtKBoVJLinNd4JLoxgrZQOaIz2fmCuqAh3CfpGwUSAkmOIalxOYGZbeVLOb
3THM4/Kr34XaJszMlc0UfkNWvv/AE+ipTbn75DjIwM6lIw6VNA1DRHK8QWcks3PpP/uB1v2lyqcQ
XwwFYEshfXwgGkJKvIeolrUuzQuMkZD1jAAuUHy3l8DwcqzvrNtwBUYmFtGCR8CjCxJRCFFeI0hK
Q6ScEQQtePp0IZDkHq6t/hye4kQ4UwYtIaYZ+5JwF+ZiaqTi/Zsy9QCXgpOlnEodHTIOHwnlMt3g
XkLq/3FyE8Y3/eQOt5X/lUAzYTfHEVjjKFBx7WPwyLeJ2oLOGLUDQ/gt2sllwCOY28b8fqCT1Idj
SiXaY5Az64gXXtkzv4xlGako7M69voMrojWTyqk3iGxUXus5RjK+s4eWJrnotsiWgOAZiPYG9i+4
2znV5Ov79PxsLIBFRfXLm4XTx01mtheMk288Pj4AG7SdpmgNRQ0TZBXWgG/006HVl/9W4VnravUI
NpMiyf8SyAlDQA8KQYbEuJH+XzSk1L3pVpdHVA2/1ytHZiIdH9h9SRdM/JWNToG74Lmk45j4fkdT
rPDwFUyRcQV85DOQ/0vxb+j+Mjcpkoi9CW7rZ0YABPI+2M0dC6NTTD+Imca9qjG8U+Q1IEe+DES5
TEcLTfIHWj75/71kKXsgpLSL2pXG0CJDTr/J6yq+wP0k/w4Hea6WwmgKH+3/poH3+8gwv55pIPRy
r+RZ7CktDUAR5q7kIH7rGRcoXO3C48UsSXhQ+PcBiWSCoCr17CvMirzQG4EhLKWH3RMWu4rRH7ZZ
FjPwlfNCFLdXQYqDOGlJZf4cLwQpE8wZcWys49I6xbjGkRJGCxG9lDrUjkr2LMsxfYXPM2C2lV2B
mNbbI/p9a9QUiaCTiLHKuwNK+tWs+ZEcMAgJVbZ2DHN6Vsej4ldILnYfEyMBZLek/ejpdezJvkTz
x+tKFC17L0ha5vzE6wVmdNoh5ayyCx5kY8HTs1cs7oFsvhOcQimfdzLLYA/VrLCLPi8a71oen037
rKvCpVQZrFdRu2oRRv0T1JL9zIxEKQPx9MKN7WwPD7HD2kjIdFHC2eLvHDtw1qfTQ9xM8o/ftQAW
qxN6i71drBWV541T1xaDEgUyFYyo3CR2PXFxs6Js1khAQJOk7AKhxjX4RVKDscqcUekCUWPS6eEN
5yM/t/dz+tU57t1IwsiT4uHbXJzzw2ccoVyPyk/FhunHgVUjIdwuwS8I7NflBhnfIzYXQWse5iYT
fvQ+4cp4zoNclJEIPiLlfmYtpYvBfYLtKBgsmKDB8huS5FO6cK0+PdSV0KpB5pNBvWliPB1LT52y
yOwz/5qWOuBmkra0eCXY4pTGJyLJIpD4LqMiXzczU2FIgZizXuRVjO2vQGB9tnh8npu0OGxCtfwj
x6UzHFFn9T+NXzCZ6Fghf+p5No04kyKJ3zA001bsAhFG6k/yjjlX7xEU8njOMkiD4stYWDObaKYH
NbhYLjhGQ2g/VVf/IMDoMmSnKGPg97nqCyaASADt5lM+ezNa7P7tTBIgoQ8LdWUBupO/VrSQiBng
bWzlka1jXS8b1o0koshJWY0ghqHjc84wMRpC6h8dCFT9FWN0BxCbxHRFOWnQUaSO/dPSJVBYJ5+/
NpkNRGqYsxbBqOQMKHYlv8S1w7jNpxDKPFE7VvKoQjEftxkorKikKlBd9y04UYJRiBv+NsVPNZWT
/Jyr2se+3VjZTyAEafrDaAqMeevycfoFCtrHCQXoggu1Qdj793EOYbfwSXJb+EDrgngxSplP67As
ySg+r+P2i5+blWbqxzQ+LkgXRFlqRLGwE8JbiSLphtWo/iGi0lXylSqj3qg20oMiD7HfXnLXZDnz
cYKneGyDMGCH+byL7dpO8QxaLi6ZNRMKFn6KiUGMr8SJfm3y12Scebv2JkGSGILNREiJGCzqnVyq
7ebYg8UucT7V3PIaV5yoA73ooPkvfCIYoTXNCZIKJ7W/nrYqSsQmUa+pUQ8p+w0LL6aBue3KWM2m
gQJ5R1eg2qTNJ6csmw4qFVeOrFouI1M4v5xygCRdXuXyc4iVun9ZwfHh68NYQ5AEciv9+SHfWE//
Q8yzwtG9A1YmabUxmjVvb50Ab+eFB0J+mRhuk4thJk5l3TaKYmpF6ZM3vpoX2mrSUfnsXz7Tcst1
aKJ2BGIq09P6GTI2vGHstgJleresKN+BP5/8u3x1DnLrCzo7Tf0yAOSDSOOVGQalJC7Yo9zRyy/b
jgLjXBRqrrnCNS4PKJZYGUhwRWFLao3xG62g0YLkfw1FLcNI2wjNxkSdHsYS2Ua7BnMxCmosMNrw
65M/3BTTKkWCwKVgbINPJKBnnLynj1hXcTHBUDH+A94jaWynOD4xCpEZLF/XmXEoWmFhhXObmVyS
3DUMPvJiUGnvtYrUWlI15JXNAuoaBYn2GiZmE9v90UqVEt+ay+gHVrV4jc+UVw/TdpSU3YXrxoWL
GQw4rM81aDJuFtQtsrzHb6Gq6UYczYrkQmMRD0UFCwbUrKVxBsAjqNbexEavybKVN/wLX3VfOpb2
bYOmTVsSzvErLeyXx+kxs4ECXElJQGuCofMc/czfZf1Gsytpld/NaHUl/pRDHrXM6mhCn1CS+0gZ
FYDkyyNwAqboaKwgSsunFOSpZAotX0uO82u6z3/IpIXXTWEh+zqPxeAGyiSS9dmUuJACv1IIhnBt
U8MlsTm+meOYREQuOjTY1gv4ko3f0wLKDuV+z2MvBjxBRjHvoSHgEcoaW82PgEk/HdKjVVbbSP0K
RGU0rMHo82hr7UQNdwtMlBkCFqeCI5cWekYKdj9As8KZ8Crxj80Bdq7elaMU4/dIi342+Yb5doQY
5wam59rFImgafAETHBL4GdHv4aq//2P3UwKjmXcSIx89+KWia5hMavjfxpVOy40baynKtPJmtIVa
s5EoTk0VaMaysFdUYMhe3BM3OcrpIAhhETDpJAaJJMCZ0vHjQsSXBTcFfIQshxC7otzAZ1q19V4x
R28ao+kchzFN0tvYn7s+Q1BGtkCjZp7BXN6li7lHC+ikR6xOpmJxIHeJr6mAHBnFckGGw2dK25Cp
EBmFxLLlDDiTOCC1BE6vNgeoRmORMXcat5asNOlZF4FcKpcjTc3uPqAkxy5/IWMf5YUlAWeh/yJX
IshRQbg6KvCAHoZSx8dTgBOljo/GkQm7WMPLCY5bqqat1bqxpEg6dTsetXiq2PEqMLvKF4fWyMFe
YW/pTKyBOjrkJ6+PNqJFF3eKoHYepeqZDjgjNNY3hAax8gOZwsNf/Wa7X45Y0z3CLhL+1H2C/5jQ
pg9IMYnrcSzFkAuGhQF1lT0DvrpW1nn5Y+JroUAC7FIREaMukw0rcnPwkvMFdX2siCL1HOCVRLJb
RUx99U2m/UBCKp4vYJTJq3Z+TsbJPS1vcafkFzuxjk9e9c4PFhnWMRi7nBJkeGcQUOvt3nDhEu7G
n54yrtRudyxuXqRegPqzXXmxhX7effJUE7rNesaI39EqT6xD0/vc+z/3sk47ZudJ21Ghc2KNvs+S
UTT05P4eVrFNodUXBITtPUEwsuxlonAe/U0a0Rq6UPXGuoCYswk2madVEx/nRS+b+qEu20k3vvEh
S5+cnze8+Uf5W9AY6r1atDh+YFxwo49GRAdKg5vuW/4fL/7UVZ3Hy6wzq5dQ/T6xXbnSy5Wy+Hu9
DiZ/+un5Yn+Pr35akQYy1pEuKfXJixEPzj3e7yejmoIYIzLn5H0xWlL/NrKrU07SJiRM/eyxYu9D
YnrXCP6L1ZY8jllpRjCx304RxJeCorS+PYCFIdP9Xm+WxxWoXXAQcMiaAsfqu4cdqs0toiKh33b2
5AO816p4/4RC/9BTqD3tr5dWM830bQQsOwqTH0I7lccz+qb6ZX9CyXXXrbUcCC6nYgcm3qS0JAdH
lxm9YmjlwXlKgUWaM7I4BfNVxZiYO0jQarbXfPgMd1VYts2SnOz/occoD7fJN/HHccbpoJHzgB+E
YW3WnaWTvrmzfUdw7G/SPLc/9LLpJONfgE4NwMNvypLyaJZeKs4ofeVMq6dW/KgZ2n/wxlsR/sme
6iGTrnlR+2zLTZfN7DgYjLaE4N3zKvqP3kKFbZcnojMB9v66X2D2zw0smFCHGCeR6ETLdSmGGOF0
39GkSS6qp3YrR5U+S9ByklPnVJ1Xsq780r9a1kjFuKAmApRh3BA3icTGQalAAV/szz7I5NKIcU6x
VVr2cc9bVvUihwgnWD0O1Rqd1sHoQ8cEzAytS2ymXckv667EVFhPCwmUUXsNZnYxFr3OJBhA8DU7
gSE8f5Q2XLLV4+WzYsQcIAUlEnBQpprj58pth9k6Kl4K7K2YbcvJoIC7k118/vZLRKqZbpFUBayX
fq7iFbVXnw4Aeu1m8wlYUvJj9aGvKsuCtsJGkZSZiW8ganU44E3AzvKi/weBoUmXak411zITbXZa
Qf1mju2DzCaklcCO4KYXPk1nWgge0aK7lpGUiQ2dedw7DydRaZF2qRyGK3YQKHvMCog6EyrGaTUj
Nc9Ats/Co33qBrDy9Q9GY94xT0Q1zqc6XiDMU81m/asXFnZJ01tOdRN4Cc7upvutd1EHKUVbTz6R
AY/ORCTLVdIbR+E95bLNgwspogY6o5ojLoj52Npa23+lWvQNAxQQUGOiNjEEdyAyBbz5fZy9Cq5L
Z9sOBeUFM/UcyrX1TfDCb2rYou7b8mt7wr5YhuuUZ9E6MqwlZZXIgMtC88tj3mI8SU530t6Bs1sn
RQpj8U6krcMjEK3dnY38S6FZW0t6FZkY/vyXm0GGs7QeJfnugRtYGzq0lhp5pLWcFq/q89/2LCp+
8gaNJluHBWbGf5rp777hOZbap55kXtk9lcz80+nEChYMibULniXBjH1gNsYHW0ODsPzi/y7yqW+V
mFEskC9Fdnv2n3q5+++3Ue27qPf3zQf3AiHyq6yQHo/t1MuG+h1eWJdsn7HKnX0NIMEQa2ubcM28
EB0Im+nynhXI1sLNSfweEGQ1t9o8BkRlKJIAGRiWdUdMc/lR/9e0pjo6e9lg/rYHMwesXcN4mGSF
QI8LcutEJFIxTEdoNdACOwJ95tNS7qMGG1XOmfj7fA5Swp2lxGEHX03+zs7NWXrdB6uo/Rod0sFk
Y84/gxhfI4UOFkDwDKi9tQerU1Y8/S6KodxYIcgBdSzN7kP4/8VXxf+j61pzi1+H2VXhMNWlTaaH
LTambYDnWTac7NYPFVU6kKaUT3HZaABB+JNcZiYWc4AObBFCKDxerYUoXQEZGpwy9m1LaGf0Q0yN
XTVsNRvvOmPwKCcnsqEIFPpSkiYgJraEYp13Jvh2OgABu+Y2redKw6XUcuXwpz1IkgGJsFXkGpQg
XzgGMwnMDIL8eN9qliqOEHzS4OfO/Svj2aiWyhkOI6twqyUjOmQ8sT+KQGkDNyD+d4iY5DJw14eh
1dphHE003k+NSu4LV6JLFBfLZP4FzIJPUoZeQdSXGuZFJ5iiAHDSlZMUAPWMR0aFla+kiDUj5QWk
1cBtthehqzxKwPpdb4U0ut4kbQ8rOliMmV91J2Z+zt8Ku68nOMUGhLSdwUOuFBUQlR0ju/Hl6IkC
FKzhPesAXT/4OM6GVL+S+FUtkT4mgygDRrXkYIiQPuz38P8QyJuRNAABY8DsBelwSa3t3IWLVi/7
u0TVfSWSdI8oHDFn8nouIZDOztvfHpC0T1El7yqxPnZQjoN/R+r2joKHS4pqgkMnOoGaOomLFAno
VDqDhx2PSGqoeqrvhRKUDq8ld4vaOpbOxKMdsVzE2ocvAqZH3vWbZM40QIZzqL6Ry0sHD3RX/Y1Q
Bx3JZmu0UfI+5c3qbMXOwDj0eB1AgsphtFqAjc+eWL25p6khom+V6RrtGJFlTBBnUBewWcr1LnJI
u6fgpkwa9H1os4zj4uIFs3V2ukI6mmb4CK0dOqUUqjTNdUChFFcv6Ir5t6HafSgTjuAjAAt2FMe/
KM/tOWeItrGiGmWLnnj5dXmLUz8dBX516tGBMV1FYfS9++CVsIZIYINfZAzBYA8L2jInhHuht4+1
wLOtmCDNpyfDlWWyyvqS/NMjVxBSN+XQLsF166Kbnqu8xXMxGOnfNmx8Vk69nQm3TGX0t1TvcHW3
gcAHkvgsU5/26SJM9RPpsYizHH9Krvy5F/tlZbOD1JrgUftHYLkQHLAHAiWgaCSnGSZH1VTXlMkO
qI1yEMP4+MBcOJFaM3FEsN58eApHL0Mtar89togcCeUDgPNAxnhOgVFCpFSUqJQKYbokYYBqu5Hc
tG+PPoAxgit1f65dDkfpmDNiJwUHmdCAWe8SVwviwS0J6QowVeUqpMZv0g8u5M6UVMYkvD0aROwz
N+LROCXQC9I56VHc6mbRjLmWmwxz/t+E8eXRK9L5wdGz+ptOrC8zV57+2bAvIF8O120340UjNXm5
3ddu62czsq43kfp/e1lMm28C/G5ptbzzAiUU23fBV4W82JBd+kCJBYa0c/QE7dDu3czz/vU+XKua
wtDU91mD3OJIWmmAVkakE1BgIXzVKwXw6XZZDpHeaw+j3m1f5BDRC7/ro5i0uwayMD407AmUT9aE
M24qjALjljU1TxiIWfVs50bhAv86Xeqz3SuS15vI8YW2irN6eacKp5JLhTXBFymu39cuFS0ilu4P
ftK8eNUkKz0qtgjAc/9mYcuH6gzF6N3TbxbYM9z3q3eKEsoIyuD6mllFBCUc8a5x0E3wzgJfcZSG
+5bhJIR7y52xrCUTpr1oUpF/pLbk/gUFiBtBZ/xDSHQb5nJZLo3oRBksT5I0N+AHgAF3YGhKj3jD
Mj6i1JHe0d+GvXcvGdf1PeNEFvBkqkeFmrSDN4ZrZS6iNZ+DHlAsUHDCNb7cPVaaFZORcWJ0/nA2
EJ8EprgFdvKmCjfTjW93hsW2lUDjMERHCg0np7ijNdsYs+Jxb9jdguzBXp8jCFbzynjZvE3BEhOF
akV9Y2IT6Fd7qEZoSLzsAhgvXLIJ73comcK8Zi3yCob4hOaTfRqe0tnVRA5XznEGKecWVTCutiY2
QA56Qp3jYa9zY6F7F/aA18e0iG9/dQtQ5dTUpzL2yb4u8nhWNOFnrhq2Ad88vvlKPnm8QHkYW5uK
a453fcDTZ6ww8Nnr7XNTruIJG+GbG5uNlknUckg90urWVasq3+lTdcCeD6Up+Np0ysG4GMWpoGwE
XdQ61NXrWMZXWvMhnzzLNCIlQ6l/1dXSdqcSZ6t+7GR1y1EnOsgHZPfop/N2KAVCREjBuZmmkyue
NsdNUmScVdFMMLI/SjrBs3MH+fPxDvgHdbgJoiZLbH+5EafQHfm4m7esKT+atsXl1V+Gc87RaH+E
MSqss7WhTfWEAS+PhR9ZOcAnnolVyBFfweHrxlHnLBlFJkYz4GFHt7G2kXuIDW4DpvnUUR0ZC//u
qDF7K9vYMXBXbDD0NR0vcz/gG6e3Jf9A/gWfAhBYTDsy/1ReoUmvC3X20KVj72lZ5CsztNeu7cdF
Edc9wcnEZSVrV4nqI1Ae94/I97DWhZNBddm6NEhB3/0XeQdMRQi7GLkZAeG5raWTLttbrTor1JDJ
DYAIm6s9SB1F5Sg1WELk2eAwTpLFV0g3EVWQXI8hG0k88hCUFefu8+fdU+9Ycq3eGqr6OkA5334L
GGSjfOS1iI6wB2QD/mOnh26fyxJAO0cCbtlMr6Wf0a0hXma5MzIiD8sjalqN14+UMy+45iQ6eZ99
kE5Wc/o7TuLWA/u9mxp3WUbkBIqNtPbBLzEsi4faIFefl6xbo22FYVGLsAKww8EPcNCQ3rgizZN6
eW2PsFP+WatIQ9UklgGxoyMVqd09R+6UnZ6pBV1BGzEcGGJg7CKYSOQVfU3+2YHOzHtzM+5TDtDl
lrTOT/Y+5zQZas6OAcYg0VhOs1Ca7dkUasDcKydEnyMLOmdqFd7m5C7XriAhWpeTaSg7LCcYBljv
l7MTP+7GNpQykP6xU2YqmZN/4IrWWuV0EZFElsy3KKjmL/V+5Pb03zxm9YO5XCWNbo9fKs+7SVZd
1CtsQfs/XbJaRVMDCD2FWeK9SuSpVjyFxf9mddtaaOPaTBLiyGimSu/Fkk6NxEtHkIEi7wSRBR23
DNfjgR2hLNe5NYcCSAedoPieu4Iuz9p7foESTmHI7ffvAG4yJy55msDihzlCbP+ywwbSHnYmmfD0
Jke5gA4M7V4jEBgnT8zei6Jgp7R/2hXsvk8n3za84BtFp7eB1c8CESM+qs2COlmbNIyiRViFnoic
uGLYcy/4M/Ur8k6qz8EWzW6uI2gl9XTCKVQRihU+AiplBLd45/+Cw6muRgOF2pdKtdXe6muha4Zn
UGJfMjQMXETWTVx9d7ROD/Nmbsnb1g6yVGddHV613Jy6TYgIMOrbHDUCdR4e6wCvK/uKHqfY7Qxn
snhfP85otpCCQAIRirBK3Ryivio/eRh5uEzS7k5cQrwhleYBrHI/9nw74WIKhhUwQF5Gg+DMsXyv
o4ulWEMRgl6NdOeWvL76T6reIp2/snF84HtTPOXCYhnTj9sSTkAlQ1TRKmE194fMElDL88XVXsTL
g7qGvMnRpc6Y+awUpwAstILecHdpyr8v39Z/VyF3UpGi65IqsyRoEzU1Y16xpoQ+lCgS/Caht7Fy
BXcKc2PtLwvK0UWh36/yI/M2L5pU8fafYnjbpJY5kdgAyXlV7FURLshtjvsR7DsLFpLmzQlH7XsD
uFF82TYopxdkNAfeCaDDhpFg4x/R8C6yrPx6wLL6z4DvzKJcpBbKJm0+y3eRv1lukAd0etznuiNN
w2idzGROWCLW3ggyAYERW17DEtN8/ppJ18nii7D4MVFYrMyuKA3D9/eIyZO4lC3emYxp3HAZYVZV
6Zo1rARMw1yADgzBprxlHMyTYw59HFUWj3d83x8+mgxCRXWIF56k7pzDsrHfK48KRWy5QjOo9FxM
SGwLkar7SmrWZBwsCB/z6FglMAbx3WvSEKwfyaa5Vvw/HG5/9E/rbh2RVzjZed7Ub+yA108qHxSt
K/v9ZYEf3lgzyjNOXVZd0ZPdt5blehnamf65kp1bD7dXyn0jpVdIZok4zGy1SOT0LnAcY0efOp5r
CpNJ+ezpy8tJJeLGqw0SpIThd9IzHOhXfg+llbbmyWpnlM15IPRGOveiyn+jRKITOUxVo45bVn/s
N2qq1SPISm5eMADwOV4hHzoII3ngcGjSe658x7A0ZvVDpvDOBNSq7XJup9uZHt+vem84gaSkl/Ze
8bpsxgp2XdNTCsuChxTB6AXf0a327uZHJJPPUV9jbl54Pwlj3z5R2r2cbrZuP3Dne5zPoxiyte/R
K6h5X7lMefUAta5ooDqYcqO1zudwWqV0vZQ4xiu3Rjsji7KniAoafTMX9FTSuJm23WIu9o8aiY53
ryXQbFKYI1vdoS/RtpIbk0AV7LlfnKanuLvK2Uf+A4kRzpA5DyCFrp5Ax6zMf78MSvvvu8ctVjX1
lSMriaodRz79Sgy+ejHiuwLHuiPK7pPNBPyN9XpKmn4GODeUX4oQy8556XGoMOZ3JS7F+6xKK4kV
AwHihGCZtGx7B40a+z2Xpw8sR9CNVcWX9hBJ7VpGdOpwcj3Eb2jpeJliYbkqlnY77z+6XW9GUHkn
dE1k92y9r/J4Ikjwca2HdOgwy56NAJykko4vRgOQyaSou5WG1fq3KvCbQsFHFX4Bz94qYBqD3ev8
tCI/80MuKZJct+RhY7jAGAMovyEVI9NQv60hcpTRcNMWyuHdIF8nwX3t+kfMkPbevVdxPEOpmFFz
6y8wallXNkgrGGxcvguXx76z+9zLyhVZ0sVXKdVTL1wa6ClKnlskRkjoyGyV0MzeUs9J/Ad9iJnx
XJdv8AFDaJXuS12mhPYRBrACOcV8NzYH4DS719kLTcMZq4l05mz8b6pSVUd82gk4ZFq1h+KllNZ+
3KamFjKJMOvYAMrhAP9UzJbpW2d3cowhn/eViYyAYQ8osxGzkMk0SiNnRel4pMtkQfnz0Lov3WE0
eyngw27iAKm/mC628Z73WJoaAOUEkajkSOBAhW+tddgoelLS5l22sVtt/pwq1RSBa7N16nKQIMq4
G17kAlFAWBQGyKvGKHfWLI81H77dgLak56mB4WMFhdBrQ/ZXNQDMMacwsnpx9AXbjNqPHNL0FxLq
/Nml32eyjZkiZ1y8q5me6pLe9JIdTMPWvtoCnNC7edhOMCv4HC3Yjika3ZEg04TIZBlw54qs+4Ef
yc42v/6J8MAmnvi84E6lq0Y/a7tIbR6+jN4Sy1OzPbCT5YPCwfJ9AS/wkM3HyQX9P3pYeYYsk0zm
qftpmup2SJ21oym3MFjGwiUqR2W7sb48bQwUocT99ez6mv0pEBp4ANndIgj9BcRYTFCQE7XXneCo
guRzKLt28XGGzLvVxoP/LvQrxPZYj1zL3vKu6X+36A74bWTy+d6eQFCQ8FMIFhNT+Du4pSjhdCFq
8MhpuZdMYMPIkzFze3dNzWHn4+5dQvz6NwQ6nVUWS3ie7PUyLYfCX+RvHMfpK8Kt3u53kuge32AN
/UrkEpKoaXfszYfy/5u7JeUKjOjnHieQmSxdQBDXyjihHKtlN+43XiK+c1b7xQ45FcUBXXZo9Sea
6vDl3wIqbvef/1AZFTF6i0rA1WP33DXGKRottfk38e0zWc0VrKCRAU6ZlhIPx4uSwsdbGjV2Hq3x
j+SXW1CKFM1+jgyoyPSzQHTsb79hcvIAKch4jjiGUKfsDIz6byoJQ3PDszNl8BFVQM0ALIbCHALm
3nU43bPDG6WWjd9R+wXMOumfwZ54az/AbFIGoGlqx/d823D2IapY39gym/9SPXuIjbEA0YmDLCwz
QNWK38xajPRx6ik5GrqXRZJCzdxQocE6eNQua4TCN3plx07DJTunzEzkdx5na4Q6+ifCxKGhPf6B
+G2gY9wcbQbMSlcVvmyaKF29RNxqgr3amvP7Rf2l/2BEzcmf0b5lp1W/DpZ1vmApZh7nC1HaOHho
qLXpOIFCSgS0fPfwb70vwBG1vN/l55LGx9+2/EW7pWuQf8sSynPmaN47vWCJGcq5811SO3kjooSC
MXb61DTBaPl3d8r310MgCsCmgJ7F/13ycG2CtZofO/S1gDdKqHqTiP59R1Y97kfr5ThjE3/6isPG
rfuiuv4RzuAxKrxZvBSvALsufvr4JlQ2BwWfdLDekg8jLzBWouzwnIuWSPHoXbSlzJ+31edQbBeb
SUssXJ8222pXNrwwR8BtNehPE8yz8OmJe+1ZcWdXuk0jzIGmhvQt957BDfZni98IexH5+mYKIQ3I
Z/l4zNI7G0SiGH/pNwRwJ1FULUgEv/GSDrP3TRh+JIWAuWv3KspFe9FXFzYT2nQEVNRNAOUsfDPG
g1NuD9fm+PcrvQXP+FlHUk7gUXGj0gFYQDkb5QPzSDDb9Rvihu+4MU3gz4WhMe5t0rmEl8ZzEQI1
kvVRpm1nGbX1T6WjiRYkp9zvAFntX44WdNjBYdZ2eVS3T/vUuHEhkeB+iVhaYuSscNhUxG7RrkGQ
ffE5knvrHRuPyFLUvjlKmpd2OSsDb9OTXLaz9ldKROR79gqhWDXydmqhAdD85SDzNl4sfwnFCWhA
6WGEzDszomOz5Z7d7eVLqu1s5HnE+5RLRqEa68hg0W2P8u1Up9xl90jwOfDgDE0rxOvHJizva1W3
GBjlSpApKelbpKeA+YWLhRF5tRIupk79ieA/clEM9w49y5/qRF5CrXhrG/kleYYtRKNyWrbi2eur
eEY3ItaSeYWM+5eIyC+ZjQfB3rocvf0lUV054WIJDRwYla1ltwy/JgpgxwcX/FX7lzqov2yOmsmg
XuMGATUp5yUFqFCnC/uNH8fsa17DS9YZCIUreyU482S6AMeqpl06UPmF/quZe4dx3+5XWQQVsSKu
MbMR/xQUj3/MPIr6LCxAB2Hq9VjUODJ8By2BP2Kpn1KQ5PfCIVghEtX/0hR5abKZJJVnKjcGj+7H
cXeXgP8AvvKOSX9ZQcXpe13I0q0o+GmS3knNA4x+sJVdqiP0B8cVEZQJHBHMZ2uPFhYGvGcIwPMH
wh5iR5lR7cjsn7ge+pQbNb8U2iyWBFbLVxuCHoGULHKmETQPMrIKc3dEVabz8dwxtXjhYDwyBQEO
oN2p86C31hZAUunk3fOaADyF3Wqdy/MtZG6cQbF5XfBmopyRuLXdcYO3kMbe4HleZCAVPu2OUQH1
C1LNB223PCBYl9qH0r1125nWr1VecQCGIOUYhxq/NmUHxdLokp1QpgbZemudEeSHgWwkooeHuBfN
CJABp6/1wCFOm+cDGmrTCZtGNtQPHYCAQAPoUR9Z/RBiMSx8C/+wKoDS5q0Idj+oHlEjv0z9r2J+
K7hBGgMpQgCkRe40VcII/WfYCAitGIjAdrTfXS1qtrHOvlH0qXTy+FJHI8oXRH+O5NSKsQ3mfgQp
xwmm/iUYlmfBcPsXrOXVw9tlEXIAL4wTbu7pRbCF0D1Vqfz5y7QWsXwbleWNd3l3rmH4Qkb1DOv+
kYO9zf+bg5bJD09m+69ZMJ2sPOMbz8q4R3VsmCDM2C6cBrHByIeBtCx7/riP/G/6/Et8V6bdsTkD
XUk6TbJfeOfvJYu8DOh3qZO2D+kh9DdDv8iS5Rl2WYd9KoGaggkaArbM7ZSJlEbHF9oolbABKZ8h
GGanKxYxlnF4dFcU422GnUCwMVKEpT+WXhwcyFvDkeIbxaXp9usM+utZqqr0XFkg6SfUfMVP8fit
9lMnK9y6U+UsZg/R9eazguD9nL6nLNd11D6s+rj68JewWaG3Zk5G+Nwh8UfZ5eWfxqpIb1cXjxG/
5Ytcn7BYCKcSLNzlN20oia6K4VpAe5/DeDK+btGckG+qLyikYOobS5thHbJbA1EdEAjUhTfZToRw
YaozaJ4b4uztvC7yHDe3Ps6Y5/W2Q6HbO5eok6O5ReraTHNN+sDAARx4oRcq7a+d4DekB+id/NqH
CMw6nY701i24QjK0TxXHXuYVBl7b18Y2kTKhfUi3kQ33KdZPxuv1pA7VZLcedcGo4Kj3lz/eJMjl
okPOrOmymjqOVrYUdDT9e/xeQ/2hvuBLSTIMyGJAasVJKjnFAkrtvWYNIhk5mdaIChSFUQ4ZDVY0
hfP5WqEPIsRSbT8UzbJ3khFtpeWa/SvdzC+xFzydPhckprP9uZ2NQcMpUb9Edm9rkjW5hlA7uejH
bFwJMildOBdWAxX/9qm5cJ+3hARMrzeIWGZ9P/TPtc8d1GCLmdFTsfgDXtiYztCHrDubZXMtd8at
tKggQMVMr/rPZtcbxfwqS4v78Ek3PcoX3B8QuRE1xRxrvT+ADidVsKcUGM4p7eLWoM4cZuqVCvHa
H6+oTswfsd1/Ble59jMMu/Z4sJhxJQcLTsNpfnigKImn7NbiOP4HNpq4QgXGEtA0m2eyQq5RBK+V
j9Ewzf6CGfvtG3kmCi/TTC5rY1QgZ3u02hiWtYZhWD48czEc1ytyeT46iwI5g+dYB9N5cn3WmfJN
7lh+V0hGNGfndFuDNDtV/bER8oY+x5TzOQUczhUi/bUATKgEG597w3Hi1MhLiw4CDWC2edXmsmtG
fzaS5Hnf1x6imsCqapeCMb9K2BQOuhszbxHxkCp+wsR4e2KQJhfNuUCiWXh5ORd5zeH3wpJnFlW4
hS5eXCZyv6cM6zapbtPga6fNs9GIGB8CaMfvi4gv+xC3ybi+ggau0Jwem/FSQ4LJHcfOeYOehUyq
Rs5mHa/kSBnoUS905N7G5ExdfVU2bVD73oveRe5j1xNHgFxnn84naoWQCoToSfrIQ2WDv18uy2xQ
1kbLCAlKEx7QyI1Wt4uJCQKqGhKU0sDAPBPm1+ng8rGou63yqZzAPr5iCuUwZLXU0k3fxtHOXqYd
Yd89jNncNU7n3SZEFo7+J+0XsaUtptKCrd8Tzs0CVh9/P5p1u5jv9D8oX25QmI1iDb5bWIngXhjG
sK0q6GKr34M3qsrna2NTH5LnYK7omPciLMdEDOpZ1jZa2gCVc3+yPeAAkabMbfg+Yytx94zEtbIr
5We3c2MTzveJk7yEyzYCB7OlaFFcI+MyYIpr8yLM9zLV7O9QxuQzuWf+AR/RTf9KfT099F8S/bnD
u9iOM46uyr2HYwm785VkSxiwceBq8tIaNFu9IEvvDo3X8+zS9ypreW8kWPVJG4OP9TaHsZTEAsNp
wCXB6U+f0gTUur5eGLf4QmDKAb0Qv2dCRhElUp/m89KwWprlhsg9S2o0h7ts6MPEdqG/aLkSEJYA
a0tBUQxJSUfITx9qJ6GVgyCTJOdN60cK/kYrJv0t9/eO4F25e88JmyERQO4CF0wcCTjKm9XMX71Y
XUr1PxgaaOFkF/peo1mNBJ/qs6MVx73bx8ukQF0c2jYGoHdEx9VpZuhCdObhXVb3oDKW2z59zj5U
JOOjhz8O0TRtPdtlHSRszzVs+Nl2Ssdjj3sK6ala89G62O9sCCLgpI9HTwE0fnOFuRp92ALDZnQ/
SErzflMP+P6Z67DyPQ7S9KwaxtrLdbbO5twY2izYlPiSpXC7t/qHruNX7OWp3IOqQJ8Cp9Nekny1
P/9n9RF0yGt1HOnP5NhHyaqtmtu+njJydHqh9OCF+ZvjmQ+f0xLFflSHCREyy8i75QjBco+6BeWm
CAD7xh9rHqhpa/BDZpOnHxnqxy1ZbghZm+zDjRAAoHK044VkFSVFc/lN62hvh8ffTxclcqlmpNm5
pIPnh0I9JG/uF1PhClBEi1PViyd7EEjehKwo+rW+W3kZ2eOdDjQVT69STTqnuGqcshJA+kGKDS6W
GwMt0KwqzfdlQZaYtwe/2CDlI431hLltdEaTJDMz6Tx7YNZotYzLlMVi/OJPHqfc8PuH8Zjl5Pll
W9UJcyuOaKRk795QhFCaC3sM2Ad7G46whdaGeZQXlyLv5fvOfA/gKR+eqXQdRhtJ6bhhtQrlolBr
B9cZXiDmv17acGKItGHP8TyQgXXsNFNaTmbaqv0RakFwSlVZSJETzBIC1YeB+qqs2Db6uoJJ6+y5
tFQXK2hYpkqN+/dA8O9X0Bb9RFoRZTtYpi6oZn6lBV872in97ATjuyhkYsMwrbAuUTpF5EJr7O5Y
ErtRyuQe/I57igv/YRQW0/QiJwlyQjUs1LYxbnAZreNiB0thqzG7zPYwyHOUpPFGVea+HtYvdzag
JdZF0+tHmXISm9Vq/0+6hiLaU8BQeG3khcczz/bV/d2HGJLxxvnER7RTJwIfp7lU5+s4/DkGQ6S/
sZcOVDYPTPcDEgn4HNIUxsvMMTo8HpF/u7wfTqDiAgg2vKHGuj08bC/gKNAb0LVPApnJUNk0434I
SfQHZ4sbkebl37xyeG1Zf4KbSPXP5FxytlnPlwiipeqzop7eVTWBN7zvVtiSMPuo0mMS92VYqWTS
lRky6XtOkOntqT0U3kwgUrllVR8TmQtHJQ/Sh2VYDnlDbpUY/HDY2pppjMXiSxlGC33nI9bFaBsp
Fi4xh2N/PvHlqEAmjhmd5S/CvikUwgFIYXAMzRpsPrlJxmR2ew6dYk4yaryqwOVtBg68pw3Z2W4o
MBostV5GwGX2NsMtuPWU7PfS8xerb7pH3pVAj0iS9t5gD1vIdDlMIAsbV6eYBK05075XtHsTt8UU
zihVhg9vhELvR5OGHK+YzPbU/6GYrollFbfLTtHwpi90brFC5SvQmSVsjnI0LhF2YBVBdjOusFk2
jQX5Rt0TtpCt5f6p+1p5RItUGSunv0lesRv2QHt8Drn1Quurm+Wm5tPE3dm8HrQnm/vh8y5CqmZ4
+HP4NwYTe5x0P2pDc55I341HgAUtBfzzI2NO8ZZBxQnMsKMKwUmd1Jfijtwkj/FeOUXq1o3sdX0v
dI0wjpqVQPx+k9WgLPYQCm/fsUnEb6KKjpYoYSsDo5EOweBr3MTWawIsCmv+Ct1BpVXtL3GDsrcc
61ZR+UoLci8YAUhmftzLGAccMjQsXerbZvpduzPfN/Bsx5Dl42swVJgV/gUysXnMUuL+FuqNFJRZ
rDIi6jkQ/ACRk7BfU7arO8rDPKfpBrzGoMLsZswmyrSKnlL4cYJhsvZwhsxtwrsfAE9u6oOuYbGH
gEdvoCbI/jAufVvhQRlBU1nnkh+/qng/LmHXwodI+JfFgOzO/qnVC1j6k8veTFUQHLfE1DpU/j/y
LIcIhMAtShtIP6SLyctU6PR9QJg8vIJm7a1iI8U08kMXidQyOnm1meb/D/UACXi85TxppiUn7+XJ
NwU+wLnXD423IaVCFqms4hpBu+RaQKh8rLbJGIri894IGeqoX1xHdecTRQ9Sxm7cyRarUozg/JO5
X5SdDQ0TVVS+QP/Dn0KhwKZxXl136frFJ/N/HWRLUmar51VKxLjj+fpl3WrUb+CDAYkqvzOym6Wk
FevfKjzITNh0zjDXiAQhYZEI2lLS1j8O76RvUGCnUf+hdtr700oFenxleK2am3SVgRzjfSw1MAy4
3c/d915rkTPWThJj1mv7p95R4zS/l2OezNwdm1PaItYe61OgVErNAuiATs2zXR7oPUO81dVlTT+P
KAu6fwP7eAEKB6jYVdcusIv5HTKLz8UwqpZxBytwdwo2ND3zVpFyDs0dayaZ0RUC0cjkXx8pFT8H
xTqelH9nJC3pJhAMumTD1zmqxo+4OteNCIH74uT7KSY7BKKiecFExLKDY5rspHXCT55xXfclIwfx
uurwAuqyyDuloBiR71xulvbw1ZARJuibEZNGlOqmxppBUFhEarZs08kY2hgGcLFvkCyRtvnlJjYo
rB5f/H6y2G8xykICRFMkxPcPMUlmzwuXgHZtf0qYh4/rdBCbCqgm6WRYcyb31AQhj+YTN9H1sPJl
i46XxvOEXXl5BfSEdUz6JZ+NS0CEG2wwDB1XcGCc4YrzroxuCxaqxbKo8roctPxrsX56vv0/SLty
RPehU07RM6kevpJQzELmEmBYKZ76lvdxfF2IvVUYKJHZBw/HgIOJlCPJTPiVs+RIBBWJdElcOVgg
ontE0F70f4AYTwXLmoG4DPp2DaCm59wQjgD4eL1BOToi17Z6uFK8bWEC0V1AExCxFy6xxMOZQqcI
e846+5dvtqwQrUJG3EVYVDvyTzQJx+hvAbD8m2KlKaLhHs1tPelkZbf2/8WW4bg1moSacNav64RA
vM8qp4LRenL7akp3auHvf8KAnmkKkJLo72sEjeTmmivpGAAdceH+ap6yQZtQ8Hb7VGz3PeXvbcc6
+/EF5ztK8WDl6gJVuFscsOV8dpem59akk8F5IAhUy4jxO8JPUcV83KN4ukPJ0sOKkZEZvtYPp3J7
z+WDLi0FCu5FxjZFmM6AYZB0MWcJSLtPX5GBDr+Smxd9aMCRG0vYCLyD6tNxCyVmpyGDuCfr2HXs
2WlEL5KWJJeZr4Gg0vLcjTfXX6MPOZM0id0bxyjSog/EppPrMSXhfCH7+FAg49ewWlyy51h/bVHA
Nfhx7yyhwL1VWxQQwECGNE6/MUMh0HNRtFRTBqYswP5iwgUBVua0iA+z1Y3pahXltmvXe+pzv1Qx
Lf6Y5Wch6H4ZACkCBMH7Bg8xIJulc5V6NSyqbVkyngtHa1I9QNaNTHXemAZYgiTiWx7yix1BeIUO
NCc/O5G0lD2jqTsbAYb6AngHLaYtYFkcSUIia3x121s2b+rr6T0eF3DCHMRdiwV3Bsenx1wUPJUZ
/zl9TnHCiN6nMQ8fVcQvS0PSbiZkjPlaWSS1v/lbuV7GhgBlZ5/CeMO1FQdpQRoLPivVTF/VjGWw
Je+LDdgRAWTX7xLDDpN9or34PY0sXahiGwxci77Xl/d+qMhYliL9dULgMHcDXmCz9xwcL6zBQRvH
3EYwFlWjMbBuugMpjGlQQWICqZ00OceFVaPNMZjZSp5G3Tr0lJLWg0mPYa0xZRsn5VaBbFBEFHWZ
sZn7lIbOLp8LeYTI3GVWbVyJVaJzzRFvuZBfWNCbVpnbZ0QC8RUZHOputIPZpJOuPUwBWDoGdSyC
zVt1+5nwNj2Ynx4d9XHlY2Zn8NF5Q4P8H5juBUcVCrr3hDRCdB9jznOEFwLDRK8fMiKPsp/PCuVI
BbAwEsjKW/OlR4Ese1hWxfX6JLM1cALn34y6eZNJs7FIPMjj4ha0kIm//wKqWZ2El3hTEHxv0kgS
6Yz60Ar173Q3gOl3alIyHq7w7v1c48TEa2c1/CUoNFSkOrClOybXzPmvCy3/YaQ4Qs/iS4Ce01ez
oUf3wJIYLuqIvEMylfB5jGm8pAhCnlPRFTmQjoQaZf03qoy43o9xmlGKu4czQaJoB97aS5sbepaV
+pPlfd4RyXmnNOW7ZN0fSKKvRHCfh2LBTJCPCigfJqYHm+xahDbrfLePcL8DSniMkzKFaiNShEn8
PXGP3fEdZcuS1RxWeiRvPCeBEJhBVdsUHg9zpAKc/snw92YX4sRENAa8BydNMfoziHmxnabKMPsv
b9aYyqzcm0ZJjkc8opAYGSAocBg9OOYRQqlzaoD2d6rvt3yDFGxb9QzbcE9aZiOgGlY7DBlBebPQ
jcy+EgHCbpBlqbcA3M/pkRLTKr0qr3KwvoXkoplsmN2BX8/LivAi9NIhmJVB5bM1++MhthaXWHjt
GJ0ZmMaJptzcRP2TRXq00pQ3iJcL29oUXbVO+Wx9cC3EIv8GM1H9X67yBO7w/c+TxS9xWMPLGXNP
nzpw+fXoolsRJtBP/PXIbpi24az+Nxhijoekmq0Zb1EzisgRy2zJfG8U4W/KuhXe+ARVi6QjQ5cU
2/25Pf+pvVoGQ3n9fbk4XdkvZRB+E6zaQLedWnolYbOj97TSnUqCoqTdfn1gdiXGsO1Z8s/PbL3t
C60Q3Di9Qw9aPedJPnPYatLSvxr1vgXVSToWU/6js8w2D+my4gPemxS1c+xzoSNCFJ8jFs8/cBKP
sALGuScMxen7n58tWGb1bl2KW8arNJPvPBfXBLkdyULhekPGx6DPHhIAPdGy/rWopI/IJinqPLt9
dZj43Dk/oUW4aBKG0ee08OGwmWUGtOJpd3DlvM4TJXYETodQKZUN5WZY6joCXkVqQ1NnA12pMCA2
3H4Hg3t9YRjpQAXl7YStX3WYnl1QloiQ35PmFCYT98PWr61R6SF2zdn6WM8q6MoBsfTzvPs37giW
t8sjXAgiE8lOnhAmHMA7IstPNoMX2EaHOvHJiBP7M8lXqRvFSEQiACMGZxb9ccrzgFl8GZaZSDJw
HNw0YqI9JGd7yz1JsB63DA1wJIzsLQhIhI+jF44POb8gSJiW3j8C7uIUak8fNrUSbPobdk9eYrCi
HeJtbDhDMtTr2tqRdYMfsY8iOcgvwKccW/hqKvICXHCKTPNk87osWZWCKNUimnU8Qsmws6RkQtDa
jZJvD8sVl01CyQchteuFmmK9mFFVF2WBqVAMpNWfzZ7c7olmJuLq2L+3Z6mDqZLYU8us7WPHkjJ8
z7ZEAcNIqm6Jjt0Z1DvhPAPiPOSexDQNCC31SoK1bHRCIysbOAHlr5rrnDMngiSBYHgBEj1XXg4p
QgiRs2DPEgzJy4JFmnRIkwK3MYRfvmPvvgRjQMtAw5dH0Cdu5BLqcOGSSHArMIB9eFx+bc2J4CMq
3QuX0v6ewa+oNzHijd8SMWLWrDp44MZygi8DZezAvNGHf3FsUOpBlmgLEw16BjjmT7gnA3uDvr3E
28caXBO3UHg4CNhb+tEWvsrhfKAFzCIjbv3syO1vHaH3DK6tLjrukS2dvTtrlez3nAdFG1h3icRu
nqLVLkMEdQ08JMHgQAwzTQqlV6uZDPoLCH9OTA0GpS2geQtZWFZZQ361dM0rvR9INydb2bnSG7Sd
R9K5JwJZvSZtPN1Dboxoa7pG2NYvheS+GnmdncPQICLblOgF5EwcehamImQY4GEflSHcvyfpyKnY
5vLDeqGCt7qOZXvEJT1nbXHdiwbmAjac+8OgzpAEpmyjHtw7dKZi1pPuVUzvRKm1xYVmo4h7jsud
ryvdaeW2xp+20D7ddAaJqiOthVzeGJdfaUNlcFAbcnhV3gCrm0D11LdGiTa+n4kpOYm9hy66ca0Y
uza3OYDDSWoXYpp9969qONgFOMLgR806twSfBuNzQS7I5O3rWk943uL1HA8KLtkePikuUIhL5kAN
56s8sr0sH2aWc3L9xb5f4UTkIaKts+lwMHjh8v/gujWoadhhTwtdCP4JFMT3Gt4L+uMs/6G9JLa3
vyzXUNa/1x7T7bQJX8MMVFfkkuYjvHdmmjnqmFMZrdh7+FHxGXvHuoYAAE0HXTIrzpZ1+7b+oVtO
m1kM2FHV2JQiWGOkTRvBZov8xb0olqwv+8aPOjBNXSnSbeGKSkj9SDvZi1wRW7LJYu9GD3IxGgg7
ajUqfJuo7aDcLc9gY1YCbqFvwaulP78HdpPVRSEuW8iw1raTwWi2Dl0o1vgnYmW2jNGAgLfxZyvY
TsSp1LwXkSW2baDQxCaLa9Al6OfxPo9IZHyNs0hX0BdvWjK4K2dyxe2neAbdRBk5cJSYyEXBClmz
4+AvrbOPALd3uDFIFlJ2YwQGHwcqTMfp+z7Ipn9jMjF/3LoHmp1cISACL1UrK5U5GfCd+Fs5ofAv
h7dTJRbl4G1hpU0loEbRT4Rp6qSYPi3PYOTg5AlAd+vSOR10GQRFVP2BVhRTZPSSXecywq+W7TmX
BzeN2qS8mO/91sE04/yEXJYV9uvE9cO/Ffc+gdr2E5B0ps6tnDs6mdXx4P9b4JlVT21FVJ8UGWHp
elh83E3I4YpXMl2GDl0cxNAOJBJJIH24n1HlqFgFtNva4XqIusOCTGEGFv2EmBz/UKOA1qmS+vWe
WCwaxzG9PNq4D+fGKHqleDksy8XvQ6DVVzoTyfVSQLGX4GGAruI1SwrRSbbX/ZcWHM1AM9+I3oIt
V7WtCJ8DYF24QQXy9k6C1ym1Yrr240Anj9aRkWBLAlCeZUiZeaN8r9jIcTD+ievUvr3/2efcjNds
KFo5PRoxx9IF3vXVl+M7tJG10jfpIeqZCtHJa/7cUqMa8yTSfJlw7Y9bKL4CfNGz4UesewPfaLEx
Tv4y4nkvMZGrENnI5nvjgbHUJU6OPgDaAshQKsMmcbJT2ja0xVkUDffsiaz5zE1tSAvlQWzHUR0e
zwseT8lnnLMonEJ2z4kFXOcHsWdGPjhYKxsDh/FicrklqaS+u5DIwGkM64wN2VwOIS1n4I1MG16p
oIvdp0lh3qJsGfNjUNoqoFmXrCwvOrv8pHCF4gNQTcVu5YAaite964FQIkNf9ya1Wj84uAvzVkGj
cGDNYTwzjhurv2FVjocNOFRH4e5TgzHjY1DOCR3ivTtSwgZRbnjOn7sK96AWpSReZknYOuaOFCs4
n7uOyrdqREplwtlhqaTAwFQWzDNle3UONDoE5+pcoiFUeV4dEbZm90Iig9AcXaLO570265juoFnz
eDy5vuChU0+gS3BjMs7KIjk13XlyLYMDEARZdRhdU5R5L5NjDqRc3lTLQ2VfahgIaTPIxfFt4JvO
sdv3zCE8jvjn8mXMVHo4n2jDjeIG5nPw+1tLw3JnWy+B/DpnwMBuHuZiOGlAn8wCeeKXzTUiifsO
5R2Z+CmWa6uF6AeVDzksYWa2xrFQ0basmbl56zkGP1SSeZYky92YC3Vqt7Jq+N5zF1WSINsVs55d
mwI6Z8zeWvk/5sBQiLJWvpxtgXniDtUgdQScNsSV7gSQ0WT4f4vnbanlO/9pCbWM7qwO0z01LXkW
IQX6IEQOv3JaC4kxpdk+MpE0TLiQcq9kNWygPqr65QqlNrvrNi52p37gz5Z37npLjyFasHLDB8XE
x5Jpf8l+1YZ/LuuZeVnoxTR8LHht0xgPTX/u5I5m5bUnR8Hb8vagaCc1Z0fDk+KaDFEi3Z+aaoUV
wA95t7/6N4fLRguvKup9z0oYD+yjXvoCUqXMd61ID5Bjltuj7ZFUx9NN7CURI924MOvbvO3fNuBu
O+l8NQgFqTLXr5V6ML6P2TROskYUen8lmG0MR+h+jRpjqPF/Stn5gt6IKtsRjG9ytlIzOXj516z/
zsoc4KkBh/kjROXChAu50EGsgbBP8dnKBh9Gp9/5f/PDx2Bg2J4QnobAbKZXzh7bG9M9c06+IzHM
jjC9/JRGqhOT4JMEgRIERXT+2op1M7Kasl2Z6N6qWEH47t5BQJpceDtl26FuPv8RkV1A7Gb+CCJk
8NSFw8GRJcGtfGM4mrDAGIjaFblbkA3GEDjYolb6epNNsF/EQkDEyrcXWleP0Nfdp2VOIkgvlU9u
k1qysN0DOhp8bi9bbl9Or2ODPvuSESIbqcRSc1JR2IdpPRR/QFId2hiX1bHlPj377zdfxI1XUTcA
mkRI69R3Dj88kTb0vLA+b71/RIz/r0SL/ibGbnfUs9CjAb39nM47vJYnA+NoBhrXw9m4ivVJdjvS
QYrAqcipWaLGbAXNOdc9Sm40zJKe5TCjFS8fQu09JMOYq9mBZuEH79qjz59an4x2ZsHo39/K5b5q
MNCWyTWqQJH27z0JS5AazrZiDPLlD6T5l0KlihwH9NJX0CiLVEXchtFdWZBmVxF1BpFv4GLXq9Tw
tRlcr3X8CQ+9Gb8j9iFCC3zFOXGHKYwZkUDPZ4YOVvqsmjhUoeNl0hxSgR9tNELgbE9YnzdqxuzQ
NLnHNIc9lU4gNQCu9vfUGAOt7APeQulGllSoDL+O/38cJ+qvZsE/V7QCKRRQveWw+TygINPmH2UK
gCsdBYn0ggXjZr2aoaGOdsUNycPL/Pc5cVfUn/zkatJ6V43vH7Q3tOoRo2LqYSustkQqS/vwmm7m
PS9OdtR/srfqjTFqymPTGi3Ru/Sot3z23CbBsywSKxO857phSGJo660Mw6Xjlqar5PBXFhcZ3FjV
ssva0rp0UpFLk3Nf5J4Qkwu72Tqr0Yg6CICFcHcQuO64k9zO5yL99lkpj9YHYpGNyeypMUPUnKMl
jDUJl2pYOWI13Qe0y7TjTvslDVcXs3r8z6qe28RxNUaHF2+EsD/6PRIK5o/dksgkm2lESJwOph8l
XVGcU9xa+myGB4iof2wypacX/HKWscB8N7wza/o8pS62L2I9KYsa6dSLKSs05wnUMZnXSK0FqZaq
bprlee93Q4lhU1SX96pqFcz3xyprCu/zfxayCrz+MCKNKpSLafwbqfUKlc/k5bWj2Ye0BMTBMVTw
4TE3UlBNAM+hMwRRoClgPAhOky8fJRGQ8h1UvBFfdgsac66uIg0LbnjCKEswqcZ0tkMqcTKTOWCn
PM+WpXPu3e2rOp0WataCVBOtKZK2fz7znuZMeW6N0z6L2S3X6GN/U1RusaPoLpBmvmPgn8GQbxSq
9sotrrJi13Q3NZT5TBeGdBzI4aUW/cBDkkQnK8a6O3yOwfV5ubLrOwwTooiQvcopn1LDoqGwK43X
TjHBHbzZLHA1W38aJ0UHnImcj/lWwamzY62GjjXly+yBY+yThUgF0BjJj3ha4WvYKOJmh9nymskj
bH4M8eqERyZfV1pWns0MncawJAlwdTRpQHjasYVQgtbYShsIhcOmZl4OSCNksY6OSpLl2rDJSVt2
zgkPPTfz0Wh2S56vBOwlgqtZIyHcyz+Cyy1hi/K74OExzJzzn0mSizWSlr54M1FgzNmVoOHFVzkB
iAKzAll1Hq59SIhRERrj4kO3aun8C8mK5Lk9jSIZXvdIH0MeNxW3G31dcWjtVKhD0nGxWSBlmBKM
EFdIWA0jo6/pXguys4UX2Tfk30cwLZUGsg9pXWAsLEXSBvip7Nd9BNb9L7K2Q6iCfKTzSlNDHv4Z
OKfA2dWFya4wYbMNqyde/rPiIVNeo8kaOruTp/husZrwgTjtuw/pzUjtiCFI1SEqsmkeGUrPfUgg
PwPLPyUeg1kMOSgSK5b4swuu547zdw5XHLIPom5Wx+D7yam2ov3yzW14fhLBjDlMedPLzQkicdGC
BzVivGfZQN+SaoVadk0+97/S5KgjH/ZUDHzGels2ZUVwCeqTXPRjAcIgx1taNTZEw9U4LN1NKExQ
3ojD01EQCyUpyT98m9pZZ/ASd2VCVwDCUHWbNHZLI8tAwBDF3dNgx90qFXqn/YUaM2hUexNEeUi4
NIOFO9x1j7Kp533VDnvxeEpuC5OUENz3zbBkUJpLkQ6xehISS3hEHAxpQVgYg5llj/czrF0j1uJd
chBmDYCWlUv7wVT2FeewvdUjZVNbQMvrGVJXHkFerEJRtuTDXO5RgQoOPaVMRkm14WxGjA8vhWRQ
unkT3ZBRHGj6jCW9JYP7jXh6HVwRMvAKwwLHExmx6NkY86DeLwCVr0ITQ0xo9ViBj8ZwNCV70quF
q6vy1d/IeOz/iRCUbZVuN4v7MZc3MNkqnavm7fEv/7Z02dm/Fe9BUhcv1vpYxtNUZ7V6oRUCCv5n
vcv2HrwoNtjNkWnS2pH+cgsQj5j7gqW8jLcuGteAZi7+zXV3b6ngohTBQR+cNyw/yW1bKflrJ3ws
K7HZjZeQO8pppM/n5gQNl+FRRzOE+zIJQ0ekFGDhLWZzgXtPoa0OEnk2f1FIvq4/XdPjhuAqCAF8
K52E6epLOhL7uFvS1sfdSyk2nRcq8YoFXtv50/BidBu49L3KSbrVDHGq1qSO5sa0la6UEnzHBLh9
k28Ip95mLk60C2WsHyF90zWqjw6+eOOwUE1rlHG4GQqemoS4WEffpysns44xBQHm4cQlUtiTMMzr
E0p4u68dbQ7E13jmxA1PUwOBEWa2EJvgNTLx56/Pjmr6coIIuJqNOE0MhYeA6HegboSKqKjAWhxj
duzpSultx88AXKGgZsGu7cA46HRPS1DLFhERNq2vuSB0i2yJuXQrqntdOWFHuSnDf8VEWA1I8zNr
97jhqSswm/jGIcooCIa4lva8WSQ+RtaraNKti5NpmK3oJDKt4A+gGFZGX9IBpqfQSbIoz6Oj686g
4YNmpnAlJ5RHlb7dkbtBpZbkO7GLBZEttViEYPctqrD9zm1jukmTC7TGNPDMQut5jV/DJGfTLV8y
lzWNnLj8yangiMTxtUc7ljKqzE3UCIb3rmeVkSSqNfUf6Yxrf2hYwLbuNcRtbJMyNIHmu7Tn5zg7
xEpUkhPHwf5QRrvnTv2d0KPriUTZQnW2XiAnPrjZQIWx6GcsMZgBpW+H2bvug5znOURfANxxtJzl
BOYevxME21XYEvirTdKCr7tunH82z1dlzhNnjiLHiyvcaRbiMlYba1nKTeWaw3XIT4Y+lsDAKzmX
JX3xu9AQdGRSXlHYlSNz3ys6tdyFtu6NuYpdkdWevLfR78MhUOWZQk5ISe+j7RS5d4viibA7On+C
FggsNGf+UE3ECa4BLTU5Cj19m2+LXxXmiIQM+kFzp/xlxkbCgr7k4IMuZAmHV2zwOYe1wrgUBaGh
n9OzMyv26mjAq3m1OO8MVE4FkPRmCM8A3nabYAPYqDa2Hzt+bZ1xJYSUchXGkoAHU0UjbnIemmpx
lO5BimJEPNovk+ENqgj3lunZ07r+bJtPAJtH5LjmzfYBuWSb7LBH9LqlY9Brw0hcNQDW7SAcYGfJ
5/1Ps+xAv1OB9NlOfXrX6K43WuPBDewbI3Tmwn7cwG6VWZ6+qJb6NWTvka7DEZTKplmgfu7VDVgf
LWqce4b7q6y7B/Phsw8PnHUUzp13hXfLfzaVnF1vrc5Nm6zEpxZ/Wgm8Q+IhXf8pP4E8g8KkV9cO
J8j9ZeV5F3gXsxfyot5Sq3y2FaK595XTu9MZvW0MQxzu9noA1zAtLOA3yP0cSO4IXX3JUYAwt6WC
aiqAhQ3sANvgDekShNVLpYUY9Vx1KCll9T4SX5iLt920irz+/EQJWHpI0048BX05i+CN+haNqtJC
l7b9vAXWBw+y1gbVn/vhZ8Rf1F8hlZV1rw2xmQwG0a7GUdUTuI8e/5VmK6ykXME/GP6w/7802hY5
GFOEh6xFkDcTlb3GOkIjAJHH0eQE6yBWKwVt3F0lx/MgSQKANpz/DrRshreJTGua84K6p7nQ/rrV
b1cEE8lFMrDy9g9FK5T6bgsRjJDsvtM9sCrSCd3+JFMGxBY5K5DcfKHw0PzzG+EaVCjYTC9V/0Bc
5aACd4vorm6CbEJ0yWAQTTvZcPGmiFurlNz92JtuysB4Ot7cmcA7t50bCBedCL1uVJhKpA/rFbuY
k3cY2S9oVU96oEti/lEqg5ltjlQCpGwQYQxGtLpqnMvZqJExPiVVNHJjxarFuSa2qAOTXDe/WfuF
o2YFHIZqEPJVCgB4BH7fC8vUu7KCZF/vLrUuyuuvKF2cXBSIAjMLdt2j4FOk608XZsJH6TtD7IXq
6NZmVz67OPYz1x2eJ2vTEUTPW6Xufy9g+57g76SwnY+xwVDwMEO1l5tXHkOXV546jIzbcbFzwCpt
FqOc6vvmn2H0wdHVxXzKU7vWSEFtymhC+Uiaxvb1Xf0aTwL4sfVYVDETIGQbNxnHxHFN0J6YTch3
F6nXamanKnam7/YT3mlgIWCAeg4VrEEQLnKzam2GkA2Q4k5HIB8/AKE/dvQCHjI5Spw3+rJdh9qb
pNA+D4fJNzvcHfAERDG5g0NKQJHerzzgavXb6No0gnx43ud03uWu6CsGQaUTjfokEzUcWuJsMz0v
49WPIKcmzCGzwEvWZ0AaMowmD90kMfx1STlIr+NHJttdkkGq+wG08ND/hJM+c46ngTUu0F9jlmw2
fgHN72Yh9zVqPj4KNc63ADf2wGhouL7GZ3hKeAc7uDWLLa0Kbag4GjXYmfeCNWEWBPVCQ9TuY8vX
lXtze8U6TKx+OVBzp5g2Hob5LqMSoazMovNQ+E3IlKyok+2eE0vtuZSOUeEcil2Ps0ZBZXJFuMdc
C39+ugFeNK/GkwIfntIi9T5PelFYYQq8q0XwyPZAZukd6aQhVokuxRJzA1QCHynH/+54iTQYZ911
OQRzAP5ooiCAuajmrR5CBbkVDEbuJyUQVw6XlSNAqjQiQS1ASRzxglOA8wzLiP+HlRSvXzxUkOIZ
UqbmP2ke3ZZjFlP3GupfXRihzObw0VjEMUyN8bKfyvUXZWFFxZeJ8NCoEnKPgcSKpV877YNyKmdi
QuYDXtCYYytvRnzItVrjh+lV0kN7uvZpa3H6pRC28sDJHXmX9uM/mGVxT60tCx8DWcDg+nPXDYBu
pkUNWFFSUPbiAycRR1ivyWLVHMK/DRgL6VxwEg+fkHulEy8uXN3OA0jNb39kS6+iNc9aaOdyYWbI
PzhBXOqgf9z+AhQC2E/Ru9K+9UMNlFUERYo7i7Mr1lsqv3okHMnuO1my1WiB9+i5/FghurOkwJXN
9AXner+3aQspo9x9kebyOi/o9mm2O25/vXSXPpk+vTmwxC4q/A65uSsTGnFS13gzAA87SAMQVuwe
wJelUsvXyVtb9ywy0JyM/v4RbDy78HbkcPVnqEIsOumLNu5UuJM26bg4QlQi910ihW9kiBAyHapW
kyjesIlw6GjenErcrOTy+pJ+u10vyUdJvnE0XFJP5b7q5JjueBDFbug8V/5PfizAIkhOlMjclc67
j2/rAvzk9EjV1f1Qt/8Q/g1hIgrk1dPIly22sfXC8YKqgwPUwqkUSebvSfUC6RFLg3Kl3NrkrqWF
txx/UnC6kbyctAMWXW4m2cia2F30UDeMTp7WxjdU+xmN3uy7+tGi26mo/iarPX7Xx+egxPeLuwcc
hqrMfv3PFHbAj8lplgjAtTYMfbXJSk+XjUq568/KaYNhL0bK1U/xQfowu+vHDZWGw+J8D3p9fyrq
b8WdCnpfxrqW+804XFvmHRUzlBjcMi19O3uvcPYvyPGIYV0+MxhWrZu13jMkhirHoVb1zVWcZBiV
zuwr9pXKemccJQZdt/S1VXuzXHpqVogiw4ScVl8CtNhg6+n0RwmmBNf8xaNRCh2f/bKOnbhekZ/t
cvUAQc2vKMZxgY5zh2SdrO/UhKt8WNvWNcNRHIbTug2waLcXBYFuJgl9k1KTG6hHajU1TdQyCHXd
UCkvy1iWAI13+QqV8ZaRYpSzIuesoVQxhFPZXCb7NkgMDCGanbae/8zOPv1T8pDUINnONy1VTd62
kPwNTlewRAfGVptvjKz3+AUef6MsklN+QujjrwesaS/xpuFBW+tsVtLIJpD07Qpe/KYaUKrHgfBi
6lelOosesa1/H9T8pDlTQLU1Bp+AOm+Ch5mUob9XLaLUKTKj2amJJs4YJrVW5rawbdVXtwm2uyNA
v8S0prPISiMjByTohiN7ZZIPRgA5tHO4UHb8uPbatf649Wl7QyDmg8QEFWUttZ9NNgwhysIJLWni
OyyxgxMlqHem6RXp8HRhHPYON2O4hLNDQo4UajactNms/Phf8zxH9d8GPCCULgX+j02cn97asZce
ZcUekrRKVF6mKDEz5Iic3ljqQCL7mKAPFZfREkzqFJ5qk0Sj9JOjDujLz89NbwCgm2MYaHpCBZNi
BbCurV6gDL7HEXWdvZZQ8+aTK5eb2NZs/YqqBz5flG1RNN+DqN2kE/bkKJhzBC6/fI/DCfDBjBuY
9uMI+87qg8vh1/4gKRh6OGZpQCL31wE1DSk0yz3AlYj46h3rvy6u+KSo6lq9rnwPc5MRrJCnc5HA
tyuqmKc97Qx1Fi5bFnWnH/q6HPpuS8kR3XdXa6emfpGRuiPR6dnlyTv41p0mFhW7F16tBEZonzZM
WpN66m4Y19zL5frvVij9+/6CwJfIKHxEpQYrBpNzhfDXuZG1d6zwLXYX6iFOm8F73I1tHWg826TT
NSvahQji7lpXyURePH5oEs8sEGQB3Gk8FFuY8tgbPEXCXfOHcc0QlcG79UFKOJzlxPix+qVCDN9y
C3xz9CBzjPzp/6xrEORAbPlhgpumIegxeqcaueHUAp2sGizzbvibwP3yPRYb4urtv0jk/gteZJWS
EQlRiyS5ks37OI51XY1PI1HcYf7czbfo97ehHBg9CyFsi7LQYJQxMz0UIrpVp7a3uy1c/OQUPoVb
Tgfl+qQ6e1Y2IfT+ZTTFH0ygXDBcRLyBqu1ezayu8Y6YEKBcB6/PPROia2Iq53NM45SL9hfE6Dl6
BioZMoUGumAgkYaCqvdg0ngYbqyQVUoIOn8jkBGYV47I0wpo0XoQUcfsQpmj/zEDcKu1AsbthCTm
rD2aWfKeZrAlr3zbbhIke4b0GsyIrowGTr4NE9rviL/efIMuzQVYwUKN+A1+ggytI+c+VpoKayBa
VCL2/n/8IzGXQB/5fSHYmvF8eOxIB6N1yIHSbyzdCsJPH/aNQ7BfM4Rzx3gDnfp0muCLkRicTIAG
p2u5Novukzf5+YDRHWOpNYGhhg1AgUMmrZiRDFrD5/s6QAbrE4bb4hV3Z+4FtozItrLRjzuvHi9k
RvRzm8+kOv5BPpFSbH7+m474+MWEk3dOb6XjgbPZija/YhaATV374+HaxGyiFaM1PFxENJfFxAkE
DozPqnOqPAHZhjLhSCn3NrmyQOZ+tnnNb1Zp9fisEN2bdIGKA6w0af8UcwBn3qUa9p4qS+oiG/qJ
3oc4/4fy5Zi8Bda/oXk8g8oZWkey07Y8Q4J5ghTd1EyBgL/EhKHcMco5gQyBoKR4eQ11Wy0LRJtw
Slgs9TAlEsFzhekS4iyONfLByCGrjjC2zkqUWdaXJg5w/19O8ki6XNGr7m24JFUj5YyWd9TkrscX
FdTsMOpxsVOZVZrPVSBB9UYcdBGI6oF8Rubo0Vlh/ptMfF2vymVlZg/tqIpAYMTu00KxAwJIlDof
dw6xHeZtXY2stF8G+6LwrRVUAqnbPJdPXrGUH99BroyxuAEF1MgW4+1AgQTYdQ+znWLWQgEEbo32
CbuC2KY6Xcq02ON19FkiChABhG68tJDhOX79ex8qKBJOJ3USSr5+3WkCFlUG2CaaSuJpARdD9pL5
tIDPbxHV38fIuLANQKROIL3cggTkf1zHLewWroTzcjvj4k2eF2eblC9Hc/PFioOs/lLWU/u0Pls7
R4V4dgrg59rY48zrw0a48gQRuYHhu3NHNSYIJxvMKRFzIYYknlhoYDLrWgaJOk2l9dReRBKFuXls
ZsH8XbYJxhqWEJyw/4ATe9G1FhIvZiTrnU7feIG74ZHkF2IjvpDYfMmOoM8KLOlahkIYwwyl9Xpb
9xD3FP3qWugYQ9bxE05xkj8NJowwL2SdHcL9ZbxpRb2RTylsm1hhkV18kCDePB9JaZDgpgXxRTvk
8nHxdCtUh1W5vl+kQ9wNwNWmPZvByxl5Jf2ZH2OUgHhNanVjXA9TT4Q4rlRbCyZ+6uRl93HBC1gV
45hjOCnhgurxBtnwD/pqugNUz08NtHOyO8eStbNgTwW0ahvF2vbx8DCX6ArLaqZRX0v7rQDQo/q+
nZpeoT3A18OeOudYP9X49YYXXovutnTEvxK4AIdsmFKupMAgBLddOzjNOPMhKyN6HMSU0CeJNTaK
2kEVHpCjumNfHRmN2byGif4ZBYS3pFrais9GikBEQmLD1+7kIUOb99xkiDL7U+FlUUJj3N+4B66R
btoryQz4+uJYf0CkVNR/KhqEx7NQae8k+1tJ/9jns5svXcBn1R1k6blM0OP57Gk+2Av6h4LfKZ+P
7sIhwty5TakIYyJtKQEDS8FiYDcTZasbBxjmwuL+kDu1VkUFUDf8h3saVWQBnN/00eQ+HH0Ca3MN
LiFVuu0/zfXkclVVWNuJtqWLP1K9J/z9Vnaa3ZsbAP6REahP3FzULGRuFa3OokkR8Wblq2lbgQRn
JKXMhqx/0ft856htxBxepRIIolCAwSm4e8Ph8ZCzjG8AOD++gA+wcySwBXsKen9gEEsuZyhqGlmq
Z+L+z7+DypHOK1Icvfk5nmKDD3qGbb1CyKDsPmBC7cjkWInueXvlcyIpLmDB76CbIrWFnpCt5OTA
JSN/pKcifHaSCi3PM2H/8tuiXf/biqP8eQzkm/bEdjpgwZJ48qgBNQ0FIkmJWqzaiYsuNrGweNgp
o7snBaFtAuA8qI19QXz+4qnOBR9pLBXoMidHRe+unbw6U6TYtyIM8ZAgjoDX8jbKKRtFSlFjtkzn
xHuXxMpVDub5kI7d1QYTXU/zt681y8rndxDiyQZXs95Mp07ODeTWEXJv/hjIUT3zi9M3rD4O87wU
olwW642dBmD0yPvjQqwZBGBaXCioi9tLDyNv73X6lEhKtmHnAXnu34hKcR7sUTlpOR9knDY9Ilqg
e2C0Fx7OoY3g18D4oof3nJtuoVjMOJhZTXcRrAzFOh7zp9X35il8nNhCpXhlTebxugqxIyShe6Vy
LPP3JRf32yGgruM/VZrrGGzl7V0zNbRcucRjSAreHfG3SmYoYh96Fqp3U5GdY8KrqGbGzUFb2aVt
Y1Ct9CDZ6uFHyqj3WdOQ+eLP9Bv8YACkuwLDV+Fg1NnczWnW9wpTY8bbdZHqWGXy19/rnWGJSZUo
ay3BM3f9T8j/mvRVyLs/O5S1DTyQzCZrdgpH6baJK9aUMPJnut4hCl25cxd8Afrr6Y3r2QlTyp8W
3hVxWoHm7gSnTCxEeVwd5g/VY3d3ODKaajrFy2lNXrA6kPTyeQxuxwriVsOFN1f1J78eOCgIroXo
CJgSfb2FnPiMlR1zD/3igO3lZ0tYjERgouGRQS4IWTA/uQzC+qjbj2B3W7yGD0GFjTdTk/I9C+ft
a0XYDoQRFzjZXmLNAs33R7VtetrVsoGUg4K3MqZMzVJhbOv8ANoUDTpp529+vGdFa8jo5FxkzREF
Pni8n8e3bRYvd0Wv1u0qsVW971I/QjnBan1FOtrL+yYORIFcJgQ5nP3c/DpXPs6PmpBKN4u3tj1g
mN/V4sRGKOVQ0A2PRMr7Kpd0zJ3Cq0+yiiMc1uHHDd5PBGPxKCq02Hxh8eP/Eet6CIZDhidECabT
R6V7BBPaSg8PTh0ihxbwP4Wqdy7VOV6Zc5uloHwfNnZnPWHQMO+VwbAnYYd1jJt+m56//lYIRXGq
+QkbS0jOrMyqmj2VJn9mUVvzPrmGEr+Qr3uGEQw9R2I4rG4r1hbB4loOrm556/0mvPHPeHk8gArc
NxzUF4bZw37ZhA3sieEV8jMwe3D9EnyF5qvp9nMN2eBWstfbUIOrZChFixNWeZjdhimzh1lnyQ0r
80s4PNZMnWwtHNgDTOhKnECKpiNqKAzMuLPbAoFZKBSBlOj8EMZ5Ozhzmi/QDR3GGM+nSo9HJkJm
M8JNWWS4/RJAgNuuC2L8UWRA+YzeZ6YcvsBGoHNhCLPWU3pZL9mogBoCkaRJAuAH2wGVYLC+ol2x
GLIiEHm4d8GGMdpIIEF9r1HtaYC+Tfp4zLgXKnDkeoudlAU4puSKYs/IJXydfXCU+JkkHSPVyaPD
+K3vayGXLw3C1VrCyg1SzXmcKJWn0gKiOX5nsJgq6n9x6xHYmu4ZYGAXZtb8EeeDfCqz0ynEydF3
WFsnyeDNd+qGkw2sEKRkfaJ4QRyGO/uFKgxkkmp9U6Rz5hUbpsdGoIxleKekrZAVe3e45f0hFM5c
gyGiXKmLRzM5+t2HcUppAYEeFTFXEnocD2WDvz/iyfuXpRysYR/pyp9iAn5NWnuKHZHruYn15TSQ
/Uobg+Me8KcaoPWkj4gHY+NieNmmiO4mFiAI0pcQyH3vnYgIzlzGpAt9WPawjvieQUiVWnpMlG8d
6LQs+zaua6cuNtt0bXxX5+aWgq/pcs/zKTtDPASUVcs8i8PuCSBfAUXiLTEY0gY09a6QSDFHB4kS
/PXBcPhsVnhAlgBeBI8xYxrnJ5dSGuKsT1ZpjN8A08Vqk63oiLaBGMggSVWtw0yL2c71JF6bgtkf
LInYEuuKVRoaDGgZ2uKEr9YAVCZHHM+dol+FYYkQBU+/8TJwt97baySA6k9qwZBfDn05Vhis+Oiy
ESwzv2XbblBWKyPvO0DIcJlomgrLrpZsL1MHSvwj5Owu5fGZTmnUd+pADPfpYxh5TPzIuVBsk0R8
ZUk5kdc8JWUBCk/qiW34YZ6Y91LN1BHveeFZUCGlisEdv0KIXx5AswmO11eowu7KULnbPeiSkfOj
79F0+4t0fLdogEB6DnixJvhE5Pj46bNuMWpjUaLZrk4vfMOUMK+/tYQLxjtbVbW5nH0q7esZxjrN
67C1I8uyWAMAIOhvNkmL79hKIPoVbB3vT11nBPF8QDEep6AadcDajG2zbKaIKkcA1qzd1sQnNBt6
Bk8XMN3YEKEBgDm9Wx7FeewnsXn2wJqwbWTBLQ/Ae4set9Z38YFZM4E5zCbATypci7R3ZSnomcTC
PBn9N4BUSNToh9Mea0GDPGaj6ETwgIwGq1/G8O2Y/3sQNGCDixcjERl+iNrFzXCz4YzmoBeqKzaN
4PaUd5CoOJV9nBdAK7+CCMQFtsxGX3LLnfR/1/mCRto/4uh+HdB5SDWlC3T5zk0tw1MFApb39lJL
8AnyU0g09FEe18WXc4PCKvQthPiCjTtTZiFdNkCJD9q5gOC41JZIu666HI1cpE9INSyfA2NjdWId
fpuug4zqAdgSdryyv2cNsLBeOCKkmwr7kW+VUg79KDFvGrUcfdJSBnDrlujUxzA+B4Km8v/8X4IG
16mgQG6Xq0CWPP0nFv2+M0c9c7mYkWEbZFAuHEkM8mgiYVbNETKpTXnW18WE58hX4wAmXGxU+8bS
LoVejnIR6ccR60p45KljUktIUXbH2qxMgFYj3Go1zb04nFBo6cTKhYsR9IwujkhJW9Xmtdrh5oB3
UrmQF0GgPALJ2d6vLIzaV7ssvDHQc9e4jvx7g3TP8kthzjbJoFHAxl/9G313Gw3G+28BSUwQeMDc
rEeR0qZCUeoFhSJJpei2C9gNrwuKJTCe7ev/tddcoiii9eV15Zj491MP/taUPa3SLWN7xQqFNdKB
qeXs1T6w3O2vwqdpPJBB1/CG1i7piSqElsmKRikqZjJmDMN7smY8fYg2Ub7VnqHCSJPOYkWBAhtA
4eoqYeJWNzjVgqhTRvhAkPV4mVXWmsAcRIR9hWMasL5N6Bo/nkfiQICwU2XLcl1ShQwsf+1ptQEO
+TwlzX31kCZ5PPVxdErnlLkbDuMJTf6PpuoxzJeCyKI3qGoJzQ4BnJUpa7eyLJ7NBYeXgFMXxOP0
ZboTroBFulsxx/Jv9S4fxs4d71d+ThSwqExhSwGVPIyLpjgWpj3kz3lWgPWDlAaj7qgvxgn2sVVq
Qls4zB+HwHIITIsnwiDNdPktKSChgT/r+HVGtX6ylpzK8kZkYNkhANfRdv9ia04LHTYZYarTkPAc
iOag00bFsL8JbnsuyCDnzw1SK1N8TG4uujoqjlz+U7Q8Zu2eSaNIEx17VdVvNREcalMLRHAIlc4e
ooooreRPWnTLe3LQWOiZnOeSP6wtuVosfPDGqhqrRYo25mMardyUY2jmLlaLrKcyk1rbXEdB/BJO
JfZ+/RfqyGkzvpuqnaMghFqlFNufTJxvfDOaqPeCLUlquBMBAOgCU+WzsTYpuFxM0cdCm0/mUf9I
0yesktUq07pmqhFeWC/Dd/30g6PNnAeHcNseMktva/3Xj6IvmnNYkcSeRFrb7IeAqJvqD6aKuvR2
jhkFAUr3euj2P9tpdFcSLlMrGjKGavGO9peir1jcj1MCJ/rSU+r8BsLfWwa6G6jF8W2k1FGcPrFn
tCUJp9qmBunaIqUUldaV4gxc5LbkcddfkGR5W7B3vcFJ6CrpZ4urVbnfs9IvsIOAL6+i5bTaR/Jy
nJTEJjLkURjCiOWcpdENdnR/SeFJYJKKZniqdixe3te9sZfId5Mbu8f7tdy1R7Ooc4RUOAoU0Fl+
UkJBOWGEVHofAjkXEfpnUd1UKMpsEEfF1uNzF5NN2HEowq10XCGcji7mMvk4d8sI8qqz1k+fzCCh
DVhlm0lMpNA3LuK6zIVZb9SWvWYZLpPiP2R5eIPVzPsFnvLEsx018ILS++crlCFzuhUvFMUNEO6X
/notcWtnCGQe6ZOQgL8mm36fmbcfx/494ugbk2Rpar0mPd2W1LrgWKG5Z7zaQUR4cOqupmJoA63B
/Ix+4jYAIzaMs/OvrSdMNOTDS29DdrOm9UfKUckvW8w2/QD+7+kaNBv6ML+Rix9A++7roUhPMvfJ
535EyVveDNqgYJCDhPtj0jC7sn9ldCslQiBgzDpFgMd7uTf5ElKYewKTe8kNPKkjMciOi2or56y2
S1i1OmyK342vkpKIHNHQvATu8/YDHBKz9aHbVT64od9IoA+Zr51i6PEw9bvtylEvbixzENLc+E5U
ePosKXLtbngCtBX/N7REtfXtKELfPSZD6yjjYFsZTv5C9yGrV2vD+/XPQxzK1hNr6K/FimyDArUt
CuiO5txpccSKI6lM26NL1zpIwVxgli5mmECbacSoWu1JMy4HuWfMYkBa+zteqry7/hK9qxb+Du7P
VQWL9wzOTAH40ygEQRwqrTIQkOFYqybJitErLIYM+Z54B+KuKY6h25+LbQO9ptl2Q+oEZVOBtkLF
th9eXbOkALB8mw81ZGTF2x7vokJBxwdAn9YBkkvlWotwNSNOqnI3sXSerxFMkYSlKOVQiGH8likF
umU9j3iEW72SJAj1ZwQ8wPbVnzPfKvBRnKNRCHkwBCT+3FOSVrFMcg9UrzaH3RH+32zyjRyJ8bRE
jpTkNDdJwcJKIqru52Sbres8sCJqXN+BH0b1zE4wEENVpOLGUTp91vmlaiTOZVwF1CLESDq/MOV1
KgDTCpemGmJv4kRhrD3sr21ICbk5TenAxSUMRI1hY0Ye4Z3PbT0UNyN5rwr0RiIEv0+5Aih2+4v6
i5VK3hO67OLVFpZn3NeVubJ5dsHpL7UjFICY3ZbnD2dS2YVtRHOxkDjGFtK5JRpDYtClOWY4S5tB
2T0HbTDUZhDDBSPobBQ1SOSYecsjGMyYXI1C6fmIvxXEba5I6E3t654rynDiEROH9XIU41OYyyoc
xoenQJ30ZpJPTnDwut43Ml0KrCxkJ5oA4Rkg3Qbl20C4BN5+p3qY9Ab4TPJ6pBgyRKzZZmC001c4
7K5TV0yDtLKqjtEodQTiNLgCIBlBXV7bRISasjQZrbfXkp7erQ7bkrODhWSzbJCJitZIOLh5aF/Y
U8f/p/dM6hI0H/83lUeKc4yff5Ruhbx4wUkNCS+k8e2gJW1dBmuY9OPob6pwkq25qjWvQ51JHohf
FvbCXwdH8JsN2uns3s3DUnDMRnsvVjb0vSfucs9/GfecpF2fxBravtnhBtXoDekFiVGm5j1r6cY0
BZKXWPjIX5glpxqajGgjJyDN63C6004YWtVaobCXJzACNx1j8bsdBUv6axsB1yegIFiXCbaAbDe5
lTujfAg601pGLKsMUV6b2DVHnKHO38jWVomBKb4T36VV7EAG85I071gYYZ3a46U9S5ol5xqiADrA
l0t468/CB/oHIGSmjcmBF8q5ak6C4eclGk6Ej/n3UVFgMFfDPeNvgPkqZ/kq7I+ZPpiyOXe/CGYS
VXiMUXrAKLwFmU9CadXDMuVpZ/CsWxIOmYD8fqX4+i3mOYQgtmF5bO6cKe8v0QRc/9GDQhLkDWXs
fk3TcX8iZDE2bNJmgTHUdOyvWYmOLjIp8gSXWtqUxke4FUG9Q8nBPzfg0jJIgAk9zLZd6l3WJ70c
ic4PTBwkI3y5m7ADO3Dhro4ghx3jYUHoIwB+k/0i+6mcZuo7mOwhdgdNxseq6BViAZMWjBx/+vC9
hN+74Xuuq/YQkDjojO/xQ2Oeai79M7ixw+yEh4YIAuxLvaMtZ7/7vZ8qIOba1FwI6a9U9kTIuetG
d9FJpqd8igLcXayN2hOpfWIw7Jnk+wePw1ZVxOEkKM+xSbryLBG+2wWLFvJR53HPMnE2R/Wcu3dx
9C/53lM1ob4Qw2yBeV3QBWYno8vEa+iQmxK7eCsZI347qfTueTstqMI/O/aTYya5Y3dnD3AZNxri
RfwrWg15vA5XjuIcWmqvrkum8bypQUxvFRGuhwKcXNgJg1UmWkRzfev77KacR73aCxWy3EjLc9pE
yLs/nTwN9+3FJ15BhhTHDtEHL2cvrmng/EJcewirbYyJF5718APG83d7u/K8/BaGgBArzFWp9FR5
C9A5NXc9WWM1kFWO0Mpng0PxtYwwhBnFRcmVWymmZJbGcVHiw9EtEI3B1WHiPqphorK6mEtaia1y
xcV7/SHBGiVX+vZuD9M7briCL+DmAvmjJk+COU8XCDQQiUPVdE6qsfkkEttitXb2/59i9O3A0WL5
PPR19Y13WlYFawKNYs5aoneItPjxWZcsQEjtdDZ3kxX6xXvBvS1PB24CXdYnGdY6ABsOt7yetTPw
yQu0PPBrtM0VZnNwiEoRC+IdsQRW6KaUFgMKlYm2M/Up1o5PuN1jhGbQTBpURljU9QM9o2WA2ljG
f3OQHJhLg1eL6vTN0rL4d+INBp6O1iOO72eINSd7MbkWnO8EOKNwvo5EVIUnXt3iv3HzPvDfCbHj
/pNAeRPtBqYKZYX+CRmOoCBgk//X+x8r7XGUU0iEmNIPxDmH+/Q+h4EgzL1bzkwhYMmapviRMHcx
xYms84JRBjDE0cF/mg3c08YL8nzgFvK4k49QToHkj0B+BGx/l5APbK0oO5k5aNl28B+1OjGzVjG7
eo99rhXT713lIw/bfg3P4H6eHIPSqo2Ty0AOIFHiC35mdlDp052MLVVW5pVmDWtnZScuX2f5Hu08
7J81efNsGGjcGntif1XhCD1DZ6iu+yPTHjf9Ku8IRqlL4uYTG8KD3eao+h2wxMZ8a7x52b+K3qfA
8ww5wU08VvSNP+nMmMNsay81iGMpCpunRNh1+gnCt2akBJWSfSR/EaoSqL9HX6iaUBZ8PjAEFZkM
5tN9OB0nX6iHXBqFx8/YlWcG9CIoaHpqIZFXa0ffBoh85BBWvrXFwZYSH5fsbtTfPB5Q99YTJ4rv
z/uQBl78YBj7k+DZBdhA/9BfSD6Usr3xfbZpSiLsBej4XS4/u5LL5+t2ruHAEGydtI4/Gdzw8t/A
B8aFgWg2RnIV0lbttk7vBUC8VZN4Bfc2UdCDXN1zpi+gGF4fJoXVH0bGLraK3qmD8DMe3pBMvbt3
g/x3RNw/1jyKFG8KV3gdiDsFoI2id7M6vN9rdQdhusNjgHlchnGZkRwPNfA95gHOexNpPADMM6i5
bIoL0yLiJn9u/89dHwd3WuMTAqJdjS1ohfsVTKIpg0eCwjeSizoJSzoGxwslIx3IN8mUkDGvZg5n
kqs5DzDRK5RKzocu03cL9Hfzhu7qvoSrxDR8+dIo5gkaJy5EN0yhp6db4ar9/2fMKjHoviuA0I+t
oHBzmcFS1XNRDoJuCg0S27Qq2QwJK+xzmM0ILJbvvKrXMA+MxzxDNxRwlRg7ajsgMCbOndtQmSW8
mwW5ZCNN13F43N5VVjPxWhyNs5DkeryrZ/DRyNLMUp22Ub+t/WzVzdpER6KbAR8paGeOqru6RLNW
rSHvXWkn0QyYjjZMu00lcBZlV3EadWGPdQvo0oBobEr23yIK917n9VK1fcc6rK/KNZRtpDLNkrv0
tutwutK48fMiU7m3Hd03AF5N7k9/5OsGKFMm0z1li2ke2bj1GYonV9p6yPTWTmVrUMfhtsugdFse
UMVlkUqluCBLuhLOBQDxgqFydshESXJLI8Wamt/IPBfLZnIhfjKjHvcvu7rSgQNgjxvCfSjnJBco
RzUGRTsno1JYfQr/t46PbIglxXt+B47bki42dbrchyrjzEnNSy9BotQ2STsumRVVJrRtmKgYRuzj
saVkGjS9f+5M+R3ffS+nSx77tngbEY1wyEkNq/rhTnXEhvfzRAd1I+nH4exP5KhqtbPNZhpPyTs8
Q5B3sSUdh2lNg075y7oV45mgu+Qf5yVPzHLfAUuMAlMXiqJPEZIQ0ftNFSDGGxPK7RK2nDO6WyMB
HU4Ji5ms7clR5xk2kZcnW/LTIsdbcC24fBCcmpqwEtlav9QSHSRS29JjtZttAnDomPUt+Lc2R0Jf
lf3epWHMa4ltSFqBdj/WXm8C9Fej9gNFgTZJtbWZLtS7LNO4kZxZWHuXGKBCFmGkeLPuPKJ1Mu1o
ZG8H7YCjrudjjX/qoV09ili763hbukm0l31cA6hcI/qMRShDaoQm+hzWAuFh7OWxCzKcJ5PY4LtV
g5Z7qie2BSfq3qYpmqIB2tZpedXPQxHZAAWHl4gkLaOj3tQ74DgLlQWO+1E33f9xNOz6xxYZd5wT
ZHPoKsXkpr9LD6fjEE0GXLC4HBpv256QNl4Ou/QWhGObSavA4UR/iF6HMVBmZq+8K6gqLLs5is47
9xycAL3jIyqcF61ZCi7Ha6JLFWt92QmFCz2MU025kxbmA/pSmMGcUOTBa4WeqJ6aVLZnGLjIKf/L
gSDJx530Jfsjp1dCAGRuMNHu40rZmdrKZNkP7aUvMDV1VKNaaj+MYKvRnITJNn3Dcpy1st9CUnai
wsXZcx+fonnRPuz+QS0BgJxzyHZhkVBrD3Qo0Qcro7kFdg6Ok3D5ZcnhZSWZd9Ps+tdmu2duE02s
1kgbgoD2jTuDggAt0oKpHiHsyCUpFRwDqLU/0fgA3HIfb5aqdXp/Rkz9Kc6O5WRJioH/66aE46Ji
xJVz86hgD2S9/wSSk1rhNBswZTCBN9pxPY0nH5D0FF23PS3jMVw6S64Jl0ppAINo1KmccSA8i3qq
bCu6i07HmAeuBEFEcU4wAE5KSD0qS6vC35STT6oqBbnY/J9Jb3JIm4JwmSYW6RQJuG7JrCDnUvi2
EdHblX8XjrUO17wCPBGb972pB7eRHKn/9m+zgyP/MdLTOOpz8EV27fRmem6AS+sGGSdxU5CXXmU5
WDPGYrGYXZTpwyCmtpiqYBKIUKm6PkEQjzlWYnaTz1XijqmpisKEPXV7h5jWJ1SmTaP5ciHh9PKF
QsmTBGUjB9+W745wXz0XazfZ3a1DsUINIQlArK+kx7Q2545kroVXHnwq2vpAdn0QuHByRZRbqMme
oBRDw6VXtoK+V1VXjnB2xsaYQ8q+SKk0pGlvsD5tGvLsbqg4dsuZrq1JirKBTJf9SX1QnvoC2mqE
Zmp9/ORouz9RA0Jz2gMLN8GT3qRwFdJXFZAC4cYnCtMl+ZgxfYTiZEKvOTiglNohMTUFFrDrfsNI
4SfcMs1kJYArojyWu3Asfj/ljMV5V4d0GXbQ7p7wfvZfq5XNDmem1vSMxSpAFacvDHhaAqkTcFyi
DOXoqtTem5xS6JUW0dIZCUPx9BhRUR0ZsZThFajFHeTd0bSo8emrJxfcxWKTMjlvk93sG2ywvKDL
uD3Om2tZ3RaS5qxHDGYi+RXz5Q6MldezUCmAvqu/APfybffBNz1cqXtjXf2l9SGsG5DP4kBXFoq8
HdLY7RXOK98D/pZrV12Q14bq6Gc4Hq/6OmXvU428DvAhfKiB9Er9IUQbCRPCnrzctSogSdnBKsHC
msR7PZj0YvnbTG1pMW1UQfJXnLqrcWZU2OyvPAn7jDv6k42Yh1RSDo60tt9XAXbVneWQb7MFOTEY
y+T8NhdhPwjhVIc/mDZPMW2I6vunxqltJiWsdmlHK0RFlrqjEdU2pTEoj/fs6GZBKWoIYhFeIegJ
Jz5Wsd6CHqWlzr1Fe5uErGrY/6LKAhFIIUiOnZOAx9mV4LQEO1p7Yf8/Fh3zoE018hWHDwwdy5WS
OV7GJPxu+JIlgBt03pwj9kQkPW7rIeO2aAjtTbQ8hOBPSgjK6RpQQd9CjCShsvz8xI6mrBSzbs5t
gdeAMuFkuCzg3jeCjEDiEksGNWl/z8XfnQhsi4rk2GJSsLWv+ewPbAjHJ4UMo5CEAdrhAxsjhTqi
MAg3WH70TS70MLbq0gFsT7t7V7AP2CJH4Hjo1yZ3tPAu04caTcicskpXe+mkXgdZJmCMN9aqkmBb
wfh+Kgd43Ix+lP6J7ixuQ8hnKrZUnTi+QQ6QtgFYQ6pshU9zAyJh70zpXwIFk8w2uwHjhm7uVS47
0yiY3vLeBcemcPsixTP0jUdi6GscbwQMQMBkMcgyMI5tAPN9GI0HINpbj1DIKjmIL5X5BhosJD2+
8+dDjnfisHvZYsNf1FmcWl3MP/q6MqnJDs4VYOSEvifXMUQWIsR9GYvCgqgq2sYD+HkEKu2/b7MC
1y8r5y807/H70nJcLNEJaYKJsIMgeu9H4cUmq1IusU55i6Jk/v1ePoa9LTqVuYfdihQP0LhHTejE
disyXOtz6sG0PGETkwXZu5g6PAr6xmRGd6wjMXp/E7H144r2h96/ZHYSllQc9OdqA4JipzK2l5aI
mzQIYJ8C2QHJfhbyc9pSMQD787E+ea8yRnPS+x/JvworyTRVMA4jXhRykCRPIyrrwZtBw2byZu9V
CvaYIPWQ4IHmTjRox4faW1QDnc8f1KOjT6U0kyYttMpCdQJAdKyeqhf6tge0bH2U63B55mYoyN0X
bE9tmllgFJ1szb3EoB0IiZ1TuxXILIpzDg+6RL60Th2nDjechtNryDqpIPlpBkkj+xQioVjQbO4m
khS6b7kpW45nxYN4SsulNoUxUUUuyMufaXOKs1got3W5Ujm1gLaJkjFSVaiVrxKyq6VHEf9H8c+X
DfINzTbEU8Ah5f4ZaRGI09wWnsNps7zrUJM/vdsOEaDgN0JHhHZwNcD6uCFPc/gtexHJu8VCJXHS
86s+zEk7qCnPyp1cigaHzocmt55Av0pobEk+zI36pYje1rgG8RZZqKe6S3B5v84lZ5Q4RKwrwSMc
0Yt7BwokyxOAVEVOViAA5Ccp4mXLS11WcvSIO9xYB2DjOxQMoqi9tIGLCpur+hSeyh5aYywqwIpJ
R0PX6bfycRuARNf/7AA86/BWXJ34awKIFDrHE4JxxF1q5hlpSzBr1dbpq1aDE2mbACVolUrgkyCy
ndcRqVnyvFd637lhhZKjGObGEOW8E9/XIk+kj2TG53T67THb5scyTG0/i4S6ENFm/TA92rj1wf6Q
bfVcx2dh0Q3XqnaKc23uDJWNhbVgNgCnQTLXPABc9jikGSjzwucwh0WJdfhg5iRAXM5ggZyq4xol
4bECuzTSp0fS6GAWVorF7r/JH6E2/X2x9tFOzTg1rMZ2Gxdlnc1dWTPjUH4tKe/A+vCKbtYh2Fc0
ju70Z4z0Kyx4EV5l/XEBYnCJW+H8ChS+r+XCbYU4uw2GFheo+5xIkZQ3eGTCX5BO3PFkyDv1J2V+
HHrivG8RwKOk6O11hu+GqEBw9mcAeU43r450CVY7wHnTYrmRDpCj/0TZkEOkpUUOgZ02lTIifJoU
E/8Aktuiq/e5L4+b9wjaYZTAbrwvbZ40jNOAyiWmDH12L/2znNdWMQ2qAoGPrZdSLBauyzYaAAAP
t8Jqenzpzd0RSACga+TuWrJCcf4JTKQbI+fuLSWCAIIC/ep2PkZ6+14E4pZcgp/J6HVa8dNr9gFi
T/pDAgA/dXuscN1gsEydZocNnCCbps+YhpGVShBDgTfEslLjZlGQUtyy+WggOdSEJyIDurZGGlhW
N96X566Sc4WFmdQtrrju7aDHHShDRjJCSWHDXT6iuL+rIgJe1QikHdHQ9sYqBmweOzyRQINPKhYl
wQfwLL1qcIfO0erHrjldHiFrNDoJyjI/jZaFpOEvpB8sXtAZOsg+3DNhij+POGYHaQNkN2UDwJoV
GfdukiWmUZqvD0U4rMiW7WC8qFBOdpEWBYt0WIZB7N+dCZ2N6I43lvSs9qrzo4BrykYGiCrOEnwF
LjHm2MedNQt8YseLNSLgaGBeFX/ceC3VVFcX3ls9WN4XnVpXBp+hii7BgFG92CXhOjPBLbYSyRCz
DnIIN/2mUWo3JyEy3Q0i+D8wIegH9w6oQVOmjCgyPetKnqIoVYqBzB0SFO+w8GDiZa4tSL16zD48
xVfw/EBex2DpAdLd9yQBTFrj2qOYsf7tk2F2QSy4Ad7klhgemts906PUIS3KMoWNtcdfSWVW/PRq
SZ62oIpSfd5iekDX1QTnGUuoohq6lWLTEyoIFajOuMiawdZJ1OdK77E+RteTQ/BhNe1jB5uoAAxl
vWSVTV2bWejCZw3iXjf++pSGjW5WSz9LDaf+A9Uf6Ef8fACM/rVz61WFs0I1UXQqbf2IsLmCTdhi
1p/9Ss25GjvjjjDNkOM5WsAhFfN5GFe262ybPH/ceJGn1tjAweUjLIhQF2qtIOGIdlL10RoS8rK/
8ZIGcV23squopGE9jqCq6f+eyt0ytStHrERns0kU7IGd93g/jkaZbKBocHuBhITSRrPXECQEGQwq
W/EwRNXeGCu5nnemGrTBZTLSkgmiS7qZjQcwLtIf9DcYQoCvsxbvMDnjDffzhK/zt5FD0tikuR50
c/OJTFtib+yoY4xHm5UWiGIZDiAFik3aXY8PocHG2HIx+5j/SF1RlY+X0JaqXOZirM5UOlTgmGs0
VBZwEA6xViTNNvvRF8LQdptHorxzcJj7DrRnC1WxzqsE6a33VTOLNYty75c4gBAEOzgpVtCNOocM
9pkmaPJwy6A6hpgosG+htMVRgWgAi6OK/1AtBm+1lihfJd1I3ciyog2kniPKrsilq/4Tzd8UXFmk
KFNy+NprwqzzgmQFv3CQ2Gv0w9+uGuvCRk+Y63lQ+RPidoU/crXzYiWvzqAaUwbJbOdjWTbo20GX
gDYCC4Zlyya0aCorKI71V+7tV8b3Kmmu4/V6Z+qS2U8ShsPB3HW+DhC7TcXll98kGvIMpz18rHzk
wnRuzDQpwwFnPXISrtPhj+PwcbhFAnJ/J0/h/oE8VP/xaxky0vhW4m+IP5rwHgrQPpdKRlJAv49D
v07LuhPq/LVYj2lpxi63re2NZ2hTKtGLrtTimpKoc0NIESfozUMTQCL5UHIQT9N0mEt8Mx4y5oSo
FZxotJs8+eiZ8TgVBO5QrOp9FyHuawjQSjDA1q53+aQIOVc9Wm2R0e6oQnj+ElgPC4YMS1IUxlWf
6N4BzytkeYl/AgDLr7r9LkNWsNkisimVTbl7NiqGy6GaoUbkHzuN4wK1P4YsTlfopW/6FNG3zoBE
OCTdruP6OXyzZXk68RZqNRtfZ9cUco+gztB3Azg5Zy/mvGurOSJuFRulLP3AELNkokQbxs/zn/Ug
JULs/eoGxOaSlaeZarlXBpi9MXraUrge3cdsqRqxU2FlwDUC4gD8VVklZ2ro2yEoQpP4pQ0dgm5V
/H0oYqYPayF8z1DbbS0S/xo15+BuQDb/V60J8pYaVow0b3kDFs6r4XDBT8ArtVLHFxgGQMc7WugW
V1gg7InRnMk2Vx+7cuccTzuZ4sp/GY8jX+VBQ95sjLHIduHm0VqwmKdhBpEmIzrBmWjgHU5k6Sp+
dh9joPVqpFLeA7SeHZl/4H1f3BmA2h1tO2m4Yr1AZdtsYVqBSHaWyCUyRrtFBwvdDxkeEnIRxFnD
gEETkWz6jqcC9X8JiwomueUVdy75bQDjWHh+EV0/gomqzeyEze71CGijMHc6uNmsS0j5nbND3Gvs
ZkLhFnW0b/wI5LsSAUYqMJJivXq1J3G6hXqUyjYMYXhJgZ5Y79z7WTEMGiMQQhOb9yy1XJP/jPvk
G1Rpd39VVURI5w1X+AkJEmrE4/veCtCZt4kPgihY7SbyAOxe3v+lkxwVgvhdiOZ080liEgHcYCOB
3/uBYT1+PbUVx4EO03My/3dJ3NdY1kBq5+he//yAgXUp61J7fVy+RQy+sJWbaNrJiaSSeTeoWVFj
hwKGVA2du9TQzJiCyNkOWbvyAmmO2bqxbP3Y6q1E2Z/nJyCg+35qLo3P0+YPnKrAtk5y97Q4gpSf
slFuu1kOJpeB+dkW9RETVpbJ6EtO1iGh79p/F4GskajXESocX6xYMZC//bXdL80l4loUxdoh/hqa
9YNIzmAi5f+RStPwthiWDVgzH3P/EzocWxYvMuu4kXKF3f1WgvDHYUSINBfnHlpK7XyRfMPwwQ0L
k+GoDXxhXoXVRFoIE9myRV01gwQLpTv9CMIJYI711Yks/Y7dQ/nlCaZ7LikKGACsqaYe7Q0CFt1F
1BQ2xAadUqVItu+KFdgajO66agrefKO2Twb2jcOGnMa9/OMHH4E9yVH4/xqeztFXyultlAxeDLgR
Tt+l2p6hK8/HFgxLlovdz5JV8Okxcm9bE8r20T5dI0Tu6YYC6kb58nHniKvwhKbdSN8v012ekkHu
XtcqMt3dmGRpHji3plrmsvrIgHfF2XWtBhWQUYbHuQNP+EnYbWJIaJyqbYaCcODUQfv+FfuJ1ubM
9Ua395pJdWjXTo/5V1qaUv6eE2ZBcqu3XySUBF6sKgMGv0V1O8p44U5bIEXjboKUYwyc3xkGcBDO
EdgwQiFXsktMfr+BXUlWKEH0P1yvzdZmRQ63/PQjoPSyGRhNBcemSd4+jJA5KoVOataEshdsHtWJ
jC3J6HC3bZFT0WiMPZeiih6dzHyaAYhpGUO0Dvc8IIlm2Yfzna/tHbdaKx/C1cuyKxpajVGt9LKl
YamlGm0Xqi0m547Ype260X5iM3zDxaKoAvEMiZeQ7i6dlKp9gV4ApLC1u/3n5m3ovtSQdKgM+CLG
U7d/KtIWZc+xJ/K9Ves0//ON5iffVwdbs3x0iMsHgd2P08EGLCakxD3f/9ZGggNf+/QQ8VZ3qdct
XnOQXxaCGNV/Ig4LxOA2SHQ2X0qpwDOvKmVLfFyE0Et+aBSSx1OzbuZOOakJoJgqRzkBq39CAAxy
izq4XPNb97t6wnKXeDKJdn6BmvmmrfcfVy/EiR/rQItPWFYKUoep9FXu3QxwzYUkcQtHyv2euSQ6
HVkl8OTheS/EMswiipwKevN4Ub8ooF0mFtbehH0heSBr/V5ZhpkvnR+P01Y9HrlOiWBirCLTgw9g
UsSKmy+oaL2NkyQz1wHQQzxY4ZDOWcCc27qGq/RyckwcQRzSFnlArL4+12O6fwxqoznkMHMZ2KxW
e3Wj0h8HNmiyOnq8S8CJbd5LKlP2WuUPtwmV0FZqaniUz16qnqHNzs+ClffogS+xcBaWbA8MzaUn
xDDK1wZCjO1gQiZYcPfN9Rvo7HKLlPs4wcQdjLyJLC7LIV7j9I8dK4LSteR4bZdhw1cLOXaGjzXR
yOMY0rJXCmBXeQm3d+95wBtCPlQd1RbJN8jdqpZ+7/a10bZYgprJEG9UuRyNxNLup8MGzhZIKNvl
h+Y6XuV7lsdEwj+R28y3wP1tfTO1IPcgzDlKwrl1XVvHuZkZZpnenL1Jw0pZW8AB7x+lZQE0iTR+
dp3Fte5TcAiSQtHJKAEgSMz2CNns2m1XKRGzN0Bt0CT2kbvQLqNboORXWnGTFE5J+/O6MQFyD/Uf
4O3P13IWjcbSgr+TB2xhcypNj3VJqP6BwIRm9lyAYmAK0LFHFLaBBcSZ+yZd6+3Z63nPXwMeFzX2
sQcnC7bXWu1kJ2dc7BwSqTkl0uQEtq8qmn8EtLe8dCi2jogXkdDx2kKLIzGuuA2OndtpLmpDBJRJ
ucDMu1vHKVdu7bILTbsIjDMavDP8ifd9kOZUEHjxBTT1HTE7NbJBkNItrVPlnKsGDWVLPy3I3mB7
16xTDRNGJYJryF1RSHOpGCCBOvDjohAlVswOHLBybXZc01BUW0gk1bcBIi6qXHWsSYLfO32Lgbus
YO6P0puZleYoXwFMgXKKqj1+fcaZD9tHRwtNksAlUNQMTDISncJLlYK7SV1Q/En2DlWRSzmmSqgx
DXj+zTW9VOyGLYq+DX/pBbDlZmulAn5rM7PO1jXz28jAQAdywa01P8RFEyvxwLw15hfxrc4MpYxQ
n5tvD2SOpNrVyFztU+w0zisjDDzes+ufwJxjHITLv39uo+2QrkshWnnImSGeArHhW7KPeYbm2D7N
h1Xi01c9BUVSG2hnS1rFFBgb6q3O/zkoHJoe8/l5A/IUUgZW5E6hbqGhCEmgGg1knXsx+8bSJhRZ
yoe6ezn/l9D7+ueF2GQbzsHsAMffXY27NAITxP8GFyRw6ZJb2b3BGRw9FLz8Y3/eotj3vgFay/5L
Yv3WjQ6LXgGjT1/xHuO2p0+ka0nbDNuh8AVFsp9KiR5hpAFherKVGVdC+g6/9i5HhM6B8LIA8WLO
P6sGOzaLJW0J2tffz+a75uXXwQ4edwHIPhmzI8LBs7YUPOag9Jr5kJBo6ZMN83QhnjqZgvxWO4kg
V8bKo6H1OtRkMsdXffa8O4YFt5PdAm3KbQBRq4KGmpZ5OOw4yf4gtMR1ef+hJfjPQgIWcktYmknF
tUDhivPMEsNlAxN2scbtivMZQJy9OH9UijZaYJv0f7LW0HGAfX70hny7uVU3v3PIU0SiYGhVLMpo
IKf2va2oo4VMJjOcN3+YrrHqqw1apQs3j8DALVbqmSYJfawjGjAoy/SU2AG9+shCo3hP7eVCJq2S
AiE+vOeuXuG0aQpZqLCPt121SvPoGc+893hz3bnol/K9nM+94GF9vtc3UiGDIaZ2HhPVzf7jP//u
5HL03+2SuZQ2zDp0t0LsLOS/Z4oAa/BlVx5IAB9MdojZ+fJG/nwDoqdjGfRFoFnXTM61iG1rWdmr
Ba8WgecVLJkFMVS6EtXbLo99zovv/UpTNHdnh1vMcLLHFyyYgz90kC990biBYk4a2bjr4gsaga4E
VSSkYXquvEmcFe+HSa40KRQAvO/5F41LwIKDIusyK5I60sAOvNuk7VR12XHO55EIDyTz7M2ujrPg
FwYDCWXl0w2PBKfqN2Wm1BzsimPppLm5qQ2nnscU0rQR5UENvYYrb3GOxR0FMh21i0Ut0gp4R0ID
tyIxo0egjg1TTeGGGL3Fm30+oPnWQd58ydBIg5p0OD2iXxrEE/0m/fBIv9knrhyttl02JqTps0eA
19kaRC/oTT65zn+kVy+f7kbnFvDThZjilvh4PK3+AAIvxy9jIH8HZFvGvzoJYd9WkCFmSIjdZ7wr
2Qj3YuQJyixFR7VLBf1+IPDAb0cT/R6pVwbN3V+EhiAZzRv3NXfywfr1gmC5ymSw9reHvbb8oJHy
V/kIRQSA1kGEgqVBwKK/9d9sIEC3z+jfuVUjoMH7tMqPpMUBHwL9ftnKuPj0JJl4eytbpIdDrMJR
qPRimFHzD0jixSNcQa8Ruqm3u/qYyvU/4GkK8lbSMckfBVNwcOGfjDFdTesdIr6cCI8J0hLYfhKe
hSyXM70T/dGsJwSg292oBSxG5H565BFSlGHeQ5ahYCtX7nC9c0NhxV0ZtllrPkbIp0fI2fc9LgH8
UJspjjuikUE+ZdKGIcFKmZcZKIuItKp9BwxhlukUL3Sfzz2AUAgMK0MQYwmQYUjdPs7eliGopCmY
Ztc1Uxzf6kT+9sAJIzPgFAppjOA5cOsz17cZ+PCg+NWMRoQFAIVU1oEq/tbm+3OZdPh87X6/W5Go
MouxObTQSIST+SUudX1qAO2K0NiBQJC3Jzw4Fsm/z6cIVXdq8RCDCq3sBiIvwawDKBDGlLzzpbNd
4UCkAczrok3yrEoVoBlYU/XrD86JowR+eJK9WQFZnMlzW2FcK0vD3mjVsRsmQ8cLTfG/6Qhbx0Wl
6/bM/4I171ml88YfpzHSKRW9SfxaRd9sjBTqFVaAYV333i2+1Zd96s7UR/Rvy/L2RE1QwIQku2mJ
WdbkxL6p3J0DqPamwnHQQgvFlyzoqg8Uq78risd5v9inVMuFraAY8wHunaDg1xlW+CcpAygZ5g+n
vVfi6ci7t62tZwWk6Ea2Ure9Nb+Q6h0srmsLutL6NYPfOhH6KH/l9ue+fz++hkyzF6MhQAsGPcwH
RiK4RDSjeEEHj7APZnQxEPUZzwvViLEVOkiCHGjxtH7ii1op1vSXPefDu8zHnqwzqU4+A9SsCP47
SrncBCBrlZQgM458ZuSwpZLrLyLpO+DLI+m/rsnCWmz3/WEB49LN5oEZNF6UC9eKCNhAvIMG+Uzn
P9/II4JwUS7smIrjhM9K3nDALPh7H6SSuMPPw4fGruYHa8/FzhuQKUrMf41DCL6s63bOBIZ6bPVs
uJ0agtS0UG5jv891NLVksWAWtaml6nZwhyTIjRQW/Dh7QeYWCku81yGADpgbZYZw0ctOtqSyAdCu
3uh86qM6YLKomj01uPonKAQSmY6TpNIb+S7NcHTZwM4bpbSRHsgi+rTzLt5ZANMrAWWdaxSlOXOb
CORmgXB+6m9OjNhlV8ndnPLQnM8JDRyxWkb/Bx7Vw5JnZBiotrtNAM2jImKOZeM0AxOhe4iDcZ/P
ThSUoI3vzxDF7PhNWHIL4BTF3pMNzOaSil9om2A8dHO84yWRPlFKen/cnMXSn+wwcGeHLKnDrljS
QQ403lQyrNpFGU49u1axJvqv/q5FQbHRk76xD5G8LLufmHYMBlNsrG1tVyO4KePyua0KYgaxZk6X
f9kWRXoqTa/TbAr2a1u+gDoVlc84ZrB5fgJtoTgY3kZulXVV8N28niex/HzqrBAiROCsqwtIXawv
CbhuX3H3V+Ie89kA2PhNs81qagSgY0w1KwUrp6+iVW97TT2uc4y8AXUwO7idZhZln2HbY0SlWNx2
Ku9BHfq7DY4C1UMzsweLi8BxPTQ40JnZVyy0aTv7N6I0+7MiEx0qRf/boc4nXMuX2sVbnHVYdxgc
AUJhYbrXVZHbjve/06zUaPlDAUcX+IjG8+tX5HH9+oKy9dbwmr6TgufZ1ExmWoSWERmU39tsDjdq
Gwue3U2ySsYjMJSeYxzmIErxWEBLQ3ngBAXGjGlLWE5xwxWGP8eyesWv9+Zmf8Ku+S/6zE3xhxPv
xNMyfj2vfVHB1lRUxbblPKAjDWxF4SH20AIf0Dtvk4eQlwgR+D1W0j1QkYTqQ1ynh47brJTzSQr1
J5OaQBJXEKsZageuce2RUQYezK2YzuHlfLEeFOTIvREjPuj3e2u2XCQ8/titBKn4SqxOE4+Tx7Ts
ZyIpXoqcRsuXNmB0x5QD//9u4FYGYpt368lSv3sfh2U+86FQrpibuIjAi4vZtZzZLjP09fzPdmr0
gXySE6FG4jp2uPP/cvJz642kVJ0xDAWmivpfNfW2XWqRi68fX6mtqQxlkLwcNPl828XGjKon/SIP
0hkAaTyIPXxcj5fOYWCvb0mwzuYDWUW7NYDW7YdG/vDdyE/yOCexrRlp1gDn6TvJihPJF+bk033C
csbOt4k87eUZizyJONdWkv9MMtLwZgl9f0uRJ9JLwOaAxkOtl1zIjalbfxwyl1TYJQNtV688M9je
YjUKaRP5BrPMtP2Ou6lNmSmc0l49nCQkI1oxWidrIGLdk2YWAWQk9SagUAwwh/P8QEL5n5Askir9
CefSGbcDgEH2kk89xtyO4xHLC0Hw2W2yVXhO4oLvMroZl74LT063W0P1gXzTSrlj3o9Q/DNY2//M
Y16KZDWgDXw1O0gafFhNIrsrTlO58WZlcOrJWGwsOPJFwL6EPEN0t4IiAG6RsvsYHyjQbz8p23IJ
LhSqPTIvnQ37cq2alnVWAK8gRQoe7x5QUmu5chz4xTfGQo9JOka/laotx5F4alRPT6ekh8SKIaIh
p8llequZUu7zZkEOqxuht6gyscVs1Vq2bDK2nzlDhuNws0+0cuA1oWa81BAFS0LSNNrKFUWNZgxi
EwL+M41Kqp41Ib7JNbRZDMw/KEU5QzfAHomRZgVIKe3SJc8fdjiIC+meymK6MyjYxDFTTcGXPQ6h
tZn2r4RJKQKgbPBXySb/TRCAzDY98IYrTIJr81wgzU/xKCFHVrpQr+dfK9llj/9MCNSJixMk0F23
Q2bUCJ8C5OISC3Qjs+PlgR8duxJhmxTca3/WXH8bzaKPu+arJsemVQ9dSCDBnPk1t5VjMwFo+U6K
OkF5MHr3qb/kLoBexovw3W3RQxC8iB1ZdEwrf5dHmkzubBLsWs6WzlGNmYybjSUTKe6OK3ylKDNZ
YxC5ywA9aGnvOG1o5aMo1FhmU5AFkQ0JERnGA4VmPzw8yhYDO6OxP5BQpgYSUG0t3P2JHEPOj82n
w7tNz3l/zf4Kpd2OxE2yUG+k5TL3rr+5BakW0kzfORq4qvAXVrygOhZN3U1QDlnGmpPM8aJ2c2Yr
xWSEY1/LaPfj/x2mMhR6RXG7Ks4YcvyJxJTvSdj1auluTFkkb6ns5aEd4WHZW2e6ZEVL0AcPBmZU
uvxuK7DkapTG/dUwjDys/Lht3pnJmFMvXOigUoRTQSjlEfVby9kE7g4TtFDvp3Q1qqsqnriiW92X
9MiKoloM4fExhoT4MIIMM9Pz2iul6xj8A9cW9vNe6kK3Up1gHItEx6gRcBnEGJFiZBnUzA9RY6to
Xd67+remifG/tOqSRwYBuUeG3ajIhsFhPwgQ8TXTOv9YY2jnoh6kVOIMdzO9dw8L78dIjfNmMMP9
TuJC/fy/+pGOFvATnmW8NlbcAldr+Wu7C3qQ3aDRH1/r/CCK5IRf+ErDAtPzyjSRMoHAeG3avMtL
5F4xHSacoHYaB24553grIsNq+1SHU6OJgEvbWgbIamPw7YSEF/4COFYFyZv3FY7itOTBAfI8hnvj
o7DkmbYu3gi7ms8WMFX87U50Ban0V1Hp6Ay9gbL3XwZ1jb001nGQKS15BR0RIgP6HQq0acgXZC2O
JDUoMTMIKHoJWCZ98B5+Ea9/58gSO9A+d1ibabK8G4Mj4onuK95lcSbMsfAr9G2ENuTe5QyZ3hmb
+Igd1KHOS3+U9wxs8cjQd1BhFg5VLKgtzCnMIBYQ+TY6viTkVp1mfiKP2/cRb/6TaIGBsRCsvJM8
Prynouq5ph6nUoGrA+xtsIxFukRJYOVmjOHeVdsTBwXPBShvXEb/AC8P43NPfZZFoWG08Vi1fONl
R8ynp+b665tXYgTRF25owrOeUjTg3SRX4HQSBf2MRe0sPck/gppBOKBqAp4Iu+OCQSZrew4ZnTBH
ipDwY9lPS4rbpxEsBiWD8De6yB8xXHVWDChuEmmUMpckORBHfKNn0tPKTsD2QH/53kmMsvm8CqV5
h5c5H+pLrR2NLFY0eaBo5nrVK4h+379sPR1NK66HNc3lZz8OtQhlIU+92GUauL44VXP8ljkz0dqr
WJt4BBPB55/43+HdADMxbcirErIJ0pDJILYg1SrK+FF4L6ky88KOIpuq3n6BZNzpVMfvYqymH5ej
fIq/jKtNgChcjQVR72QZeGdzJeB/7MCMaIK+FNLgE8ydvCGqkqbv3b+2gvg0hU986xzGlxzm63zu
DvwODZpr8m4kpniO/pkrfd2/xssL3vMCJjXELJtAKd9+sNznoj7LYGT0C+4/uzURm+wSv2hSiOTQ
hZ08L2ynXsUnDsqsruSK0Tq6DwJ9r8EnaTq1P3xBEd+CwWsBfxOhZB6FRCkmVgKRACMG8W3Ye3+4
7tFXcfhRn/jzehRJ/0DmUflsXpfaj4JbYLR3dp0aeRR1YTFqQ2l37Ykvvf/hXCMvLfpvlwCuv6PT
50+q9xI1CdcQmoLgyiixeUfVFpwNoCIFA4lmQeh5lgt35/OPbSsK0LWu7sIvbyQlYv4fbjZGP7dW
F2R3b75oQj35Trm+z73gAWiqdGPzkAfQYo9xuJwokluzt4N/8M9vCQpSXpg7IKC9fIlyckrkT8Tm
Edk+JsOGDqbD7qI6wVSUSH8OGDYAM4CN1wSCgLxhtyge3BtbZk5H2zWmsPi9XZFwfs6994KwfCDs
MuxjfIXJWdx0CA7HWPhcuGfZsCNAwDEtDi6yfGjKcwWeFUYYTt6/cOvbzY/Lu6EkjzVIkiXeY0TE
8SkcSZyDQUxSStMqVfVzTcOY6SUfoo44Zb2Yv6O8qRA3VmjFrFjybhy10cxthd1iJzdHB2obwO7d
A3Fdz3bE51iuhR2MwSJHvJIvRqvw62VyqDActyoOdPLrwWmtf6d76/mEd5E/9q6XaZq3oQzS/gXN
PU+KCZp15NguPnhJMUBPkxjYmMrgtETH5Sti7rfvOxakT7sDslJzh4IRJQlxi/w4WDGroB6DO9kM
QgwpgJES4bLdxhfm4X9ZWXu6s+hN/R7RyxfjC/6VKz9dqUv4OXQhBiXFrOf2N2ija6Y2DGt6Na1P
DJ1QDr3mT3dA/HJATlIfS+QbYJHSTmR+UI/BEiaX+aWlyAcJMOyRElQvBfBUCQIrcpZX+03kZvnx
WR7edN5oUpkTLHYT4omr5OH/QWFxw6ueP3oFqv4Tq4Ba6pTSg51HPOsPTGZZfHdqxW+MaUFcWo8y
xVJLPYCnZmJLfMNNQRnYXSppFY7K5d9gHB9c+NTB5vunk6Bi8G5N7io8eEsVgQqZpVZD54hYYkG+
DXtL9nKRFmg4rXHLyrRx3Pn6Yaj4Tb1LNuwP50qPPJnMeyheA7etexwasIqIgvMQ3bC0AShKa8f6
sahsLNVzud52OZV/hCFnMhe7KbyoeW+pyZYrdm1giVXJM8X2XIpGULqFtjuvtqfUwBL9UXY9idmf
cDEj5uxhTq6uLdWscRXqb5xT0L/da+CatWrlR9AfIlKtm8KmsAPV7b/mHc2HhOQ8A2FLtgz4Dc2k
OuNlk1No69IfzHmZgUeStA4EBgPjyOWtxhR0wyr+nUhZADuP0/D/1AfrOJNimF5ZAQw6jFneBvU3
ZXQHYt6OVkbnPHgKduT3kX6rmaNoYVDui1WYKKgMiVntdwprNOZTIwZoCOkDKENs/zVXEzIc0Bl4
fKZbVq/nK0yrVl6++g+2jmK2vuA8b6QVYbzVY0dd1PXvUwKgiDMpq3SWXt+RBhDtS9igNZ/xxS7Y
wLKDtjuHBrMEtBOkHo4xQxbWW94EJuDiFWZqjEYn0kDqPHp+0ErXUSiRAU37kcXBNs7YH7QQn71f
d6T5OGJLQg96CocfqzgINx9nizCJo70a/NnZrl+1z8+gAXHP5IxpXNhBoqWeBfEK7hJUZEsr48gt
mEBZg+6dzuNhhVoEuBkw29DXVFxxSdwOfcoh/SGKicBcXJrZgfd88N3UiOeB+YlKhDEjw7rP4Eip
QHuLpR1zzJWTyivznxocZrc6lcZ8FJVfUZFBArX6ol6xZ73LKU5nkWpOjZbmi9DMVTt3aheFvQFj
Ccq4/OfgTHvMY0aS0JNEWbnJMehZzeIEIxeQ1HrLc/u0ekUDX/1NmRkUZtoTG7rLLvmn3XUCXR9H
otrUo8SuR5EnPC028f6ZlapBIH1OsX65zwIZ4I8H3EgXt2cE+1BeY4LA4UfB9VdXHvnflpCSfgw9
RpBKrE8em7xEsFZqBmSe6J/ya9S7OJF7tEocB2tUysqYVdLkoBkjIzbzWTQsunn5inoBZCVTSZbs
HaQbocEs6JRVcJHNsC6XLzAjQcERmuZru3pbfF2Mn+4ArKtHYVH8R/HJBjiRIKnf+o22o3z+2NVs
fDqQvkIgIsmIhzNyIELPg7CzTQ1WkVVicpOEoAUd5dPgJSZM/593nYa+noXXDSRtWi5BNgneY4Jy
qld7PUo7z05VfVGbc6TouoTtv9qBAmRAGBpX+BqADwL1D+f+wdQaYdrlt9Fo73TGkS8KHVagDQ9H
RCCU82znhkmnouPvce6MlxeDdpbTvW0vy0PewUV7aLMYw+1waRF7OvFcFUQIv4m8xKj25f47rJxC
tZuD5FSE+bEipZd7z75aT8bvLL7Md6FJRjH0QxUFZTg0NvOafuvndIHWkWpawn6UkNkT9QWVv02m
UbZYI5lhx56S6kGJEHNi+VcX+mxn0JL7m9pGzr4Y/3zJZ39j8NN5dAtSc5hsk5Ts5opoFkvdtUuF
mAqW/qrsZzGQhHgy8ODIiYqNikGlimqgdO7SN3VEI4fet0W2g14ZNtzg3vIkhbQ4cZQaDJQ4JuDF
6PL2x7dKLqYdFlZAQLtrDDkAfj8G+i1Lfb01fLjtb3QVAhknn/vhRPUuB7DAbZfrLq+b5zLAXu4Z
PMBiorf8X4KY/Sl4ISTnSy0cG8Tbc9N2yrjPAtOhdcFEY7mlcJdgki9PsIZQRYMpjQlzRotniiwj
jJX0xjoi8TMlSmf3K3Vk/KuAqjfeSNg/QGm3C0PoYAjm2/LgSpmtQBGYD1S8PhqsihKRoWjoNa4u
uR25SeCMwgL5d+aZjNFGIOU3zV+ptM8qAVAAvoW7A/JQ5CeZonQBGYirDQEiI1WCitCLe3DHcQq5
JG+2iNaWXJvUjf00QQYmZVJjABv6+y8VTb37NybuAFjc0MBOAy1Wdo/66UFcxEkhJKtWYMXlVnBh
GBSCTOiNdbM6AxMYulWMgn5cOnurg6Yf3+4tMkwO8bYgJ//aRKnwtkKmU+Wqjg0XgXexUbacODDd
zWE53IWxLqyOx3kTvHypvAAyM1nQJbm2/h5DqXVutRr8wbFsAx7PSuE0PnK4+zw6Z2ZBITr11KbI
IlAhqmlyDBfdvYtgnMMegCi0WU65wSkV/pPU8jI6Lh2J1Hw1iAZkWnQ1y0zBgfzpKHNFlwi5aBwa
cug8BQ04dOlmEZyzSV+HRwfwmYQbozDOrXzrYx5UC1AfU3HlbozdPgHljLMW8fXU+pjyG5v/2MCL
EYocRmhxT3EchRqq+mZ3/Fca1Vs/INMSGSScQSBJm7aMKHUNHR/oekAdvFWcYJ/2O+1NU6YlCSkw
4QWtAyz6+HAetdaBXIIwDRv0cVSr4bXPws4EylHmR5ZwUcbCEcVI04de8/QBPavqqZURF+UNGu/d
iv/yl9fIzjAT176CYACmsRNSSC/vvNPf+2wgM6qDqdXKIJtwUF9dP2/17h4lx53Tn6mM1el+JFx6
WBsPAKZJH0qoIzLGXaTkwGJ6dgjikHBKpQ17cbzhef8h1M9T6CruTFUmLWhMAA+X5eSE+QzfGfwR
1DKTVH3DhKpLvLMpnKUPP5MMP3hbdiJKAzpAWBUD4mPwuQOj82So0Ql9Dl5K/UaCbQKbkmPPtAuL
0H6fMv8U4eLN1XhS1i1wlRQ75rTWmbDJi7epTVSo3bGxksPakzxWrFeEYau02ORKO5sdNY1qGEz/
Z1uv6JVPntap7lumLBkuKOfDx6cK2qNsLySPbbWgdA507CByftG/lSFEJdmBOlNyN7dAoGZhf3Tv
or8F1pv0/WESyPwA+HtDOzVFEjeiaeed/3GA0Bng3LHt6+H1v6SzhMPtRdWl8siDl/R++ER5DtDF
hnc9ks85dfAeDvfhVtMDwsUV76Ve+TeoViDxBbaCmBxe2pjVmU3Wcf050Tu6HU8U2DVGsweiGhaX
hQ9SOfwhLG/Ozzza0t40Yo6IJETADksI/wKSsCICXWCr3N+YZgMtVTb7A1gVYMiMmVgDicoNXgSF
K/lCQ2fIYwvZvrfGdoSHzxpYt5ej15WinNCdVgt3eZYKbyFVo2aM+NPYlWpnmg9MD4zGM/jLyu08
tdnermt3fUYeBAfhBY6yPmYJZ2YmVnzVYTkcfXCnG4ThJpIBLn+jQFXPrrkoG6fGcOIo5VBj3qyF
RfHN0LO/FENpDcZcQTOs3qVHHsSxTp9f69W7dcHCjcfVuWVDwgTFwj7gtiOW9xuyCQV3l9YhafjP
UD7/6mQVVGeeNXeMY9rWoQjxDYEamQ82/lqRxQclot9YnyVvfgRSWo5fu/xABfRx0/NtFKBnT7VP
3n3xKtK0ED6lgQi01Nvetm1qfTJF2jFEp33UOT8aYwWOUkg3+8TAEdQAjuAMfqfRG+Jbjzcbp42t
KXiQ2y127kkQZWKJpWjhin55Bdqb3qyBJL7Z44/7i4/BmlFAM8Eua+RHAICnu2qKI7ABk4KS4fRy
Y2dMDRmeobKoy4xWAGoeWQPZiArj+zSrYt9I1FGDBrKIeGTVtouTU39V/9SFBC1iEm87GHmgKnQa
PW+DPdZmIuda5byKnS+eF0BJF5C9EVYYH+MlDHJSeY6PXGEwz8b2/N8K/OTGf8q85OyCZdIxSHsg
uWoLtoPNdWof0FO/LCfAtsPoi2/cFe5AdvU5OMxUQe6p2jdmpXyZY3TwianUCawS7hpWWRS83p9B
vkjkqeH/wDnOa643EhX1qAgHDtSkvDB+PNF0c9aS+FGYcL55Qjgo7Vtlix9opxLwvKTg+dYF/BGG
zHkzpwRwBQ2Ucddq6wYRG6vMJNFrag+EAzz6u5Tly4zd0x23nj7oJMtYSr9B8dp/k4UnMIjlXGIQ
HVraBno5zG7gptI3T3aOZCPfe73idSapNwCUzpb6k2eJV67VZlgzKy6FiV3BeJ8RddIS9uP2R7mt
cRT6bTurpZBnRRHw0xlOzz4Au8KR3x0yhNV4yNiIoDNnZfhoGClhu6V/oNR664VVZ75CO6OsnngA
jOuuKAiuWremvaAqL4mJnKU0dR+yoPPynZFHa25D7wiDGvpsf0iQAZoKK8w4RGH+l5sXNEsVSXs8
XHGi+QaIMqqgIXuBtoMMr23b/F1933Dgm7yCa12sRHqrcelDHIsC3J2rzcr2mknSZKoNUvysWcuP
CbTgG/B26dyZq4zWVDEaiAokWiAHNSmKCXpKMo7HJ6T5ue72X5OlHL+A6BNg5ExBd+tYCvtmgjPj
DJB1ki3iKv9CeuC08cYNcsd1/OuyhsCiwZ2NkE96zz+eYxwsJdibU0mw9UOOH5aECd4zyOM4g6Br
evt9KfDss7GyWcG4KmDvJYI09+H0JMK4vE4AmjXOXuwt34D5UyYsG8DaFylg0qxDjdZmoE7fFomm
UjRCSlgZnJFeq1C40G+gcTdIi6zQQMBjeHyong4ouvC8ag3xZamArz/1T2Gs7LpMVBnYvrWomdbZ
PnrBEiUnOQZJc1AdGrKsrL/NC5lGMAqIySgkWqaPeii2VxXoHc6wvBcJq0LhiPcGTnVuuejD4eBI
ELU7l3u9IzoF8x1diDNUa/zROy9KZofq36h+bqCMA0nlz4ihzssUDXs2yoxF4FZmgHLORFPTOESq
ZBSO/hDz81MsE4A4ICHOYnrmP4lcMTkNMCim0vMDXFsvZ+Du64z1i/dTxD0RLMZI400gHX9zXq0z
gAyKi9/8/h04Im5Arfifk/4FTicLXEbiMs6QJRSjxpkvcY4KvYRAp7FZK51j88JTF+kW29g/G5T4
qxBTHDw4l3VrZWAfrOOud5lBS0jZ79+8qKvPi5ZaJkM/gvraYq7VTSOwwEcMd/WmZ6c1nFz2LMm3
9+Z6PMV2BP1Yv2eMkcC3ybtBzGgcflRmnBEzhMvYXdGg5jZIfnbRej3KcsI1jSo+Dn+G06A40vu7
J4E0N4lAp3YzWmV+BOaUDt8qe3K79y+9GpCA7pQVULutl5S677wXxW6KPAl/nV6uA+a4NP7Qj1EI
/O80T9DLY0vi8CDzaTfnf3xxF07hKyuRAX/xXe1d+wYyNPxqAnIbXzdPNld2B07gv8YcCgFq6cB5
BnhXEC1R6szXfI3qulTwYupgdDmBx7vfTdJzfsBrzF7lcbDoFwoIVoM/sHnQcugsFkivUL+jX3uW
wF/WGpdWFZ1dLfdWDa9qg0S+4tQ9GGzmNy5xZ1ZviuLswVb3HprAQDB7YuzNsct1ho9FDayKvM75
i+U63WAVVeSbLWX5v/zobTmnrU90lWPkvF+cLrpssyfaxkxey6V9Q54dU1PqqKSV/Lq+EygXb2Xy
QlF9dw+64fFvcFkC1lCXxfZoasJdeNbwF6AomNvfKifQQ6A6FA2+HAeRGeTutXkJLSo5fdKVLNsO
26leb0RLnRqTqNlE0+b5vGGZoa/0MWAenF3sMSDBkAsbkFT3yre+jbPNXwfDKEUHlnQ6Kp6k6L7s
OY791J/eQuIITybGyvj0yQXhIhSTDHezjo1G3+WJwiehdcsTPAqTUdT+YjM1KOnT+rZYSZjsjgi0
gtHS3swPC6vczyCBpPFWb8wkhWm10Hw78SfI92i2PNnBl3bU5w/tH3UOhJS9deATkS8eg6rGUCqv
qlD/RlzAsuQnuIfMexvLXWPqGJasq0fZWtSXRLuNvMmPDxeqIw8e+9cPtB51dPe8uaNRBUr3p6hs
ebkuCFOdrLUi9JORy4nFwpJWCeQyGJ/kkhM9mCCxP2GWKrQuaowzUacBP/GAQbbH5xnIy7Cnad9i
4IEH2iSa+LChxc9r1/xx3ajbqeZ8/oTjiYsMD84HtN1pWNGTxa9d8DKZHnwxD6pXXP/kszdrV7pP
/yBwvhXVEEZQbgw+d/Zh3zRomOxITXdXPMAC41S5FkRhZuXCaCT+wQpP45Lu3HWbK6x0xI2huUoY
GJ4ED2543kqEoHC8ug7JmZ/KHGYaTRd/6jBZfLVF4Xh7hnBdSFShUbDUQE1XW7b8g8j9EPh+5H/f
KnpsRVQiu2+4rhxs+fBgJbKchvii/g/fJa/joyfUu3rE3+eLrdlkZe6ihStgsHprNAiG9/xO7a0o
oYXRe7d2UPPso34GfT7e5vm54HY9FuJr7gZJKocGSOOQGcrDZ0NanF8v9O3nPWtV/ONJtplGByqm
x3y6qe0r07g0sl85UjAKwTsFhOMqKmpFlNiGBsHPyiq5F9Du966qw2sSBkQMzNyAWCkAYP3K/1k5
+Sbk3rPTmxqm8feQ0/BT7gnvf6X1t2/R0mnD8glbfkzsLC0dqrApMlMQ1YjLH/7sCtmpiUjCKBBJ
9tg4fo1sOY2NBAJBi+Y1hspq2ZV/HVChVE+Y9cIbpczOejSiB0NjrZwDLNI7hkmGZIuCee5AnCLw
9lovu3PCu/3SBFfZORLhx7TpRzWAB1uokfTi9unwVrcwzXvZ99sNE85x5tBxEKWVZsIZx/gskSpC
d0o9vUE/XJWVAVVkGx5PUvT1+81JKAtEc0/2C9czmvY2lSRGT1NKL2JXgQvkF4/mA+gTZE+CdcLb
fOOF69DiFPrHEJasFpMe+PubnlE1260znp/S4KNLKGP9O/UnA1Fuhwe2ZSdmKdoY2f9rHQJxiWyR
3OXRiANeNcN+c8qyD/XB63hO03eNZVe7VzzAl2pfm7FpOUKofse7lNxikeRwRKYaVGhmCC7oqFb+
T6CzfLcHTNanb1RgjmOlMOPzCUl74Q23RsXaGuZ9mfMLtQ/4x+N6ZhncNNaAQnixc+OlgOZod9q/
1ad7v+AnwpB3L0RFgVOk8nbo0EuzLKWH5necn8GQPa6p750HteVsRS4nznYI/A/bBy7MJcRJn+qp
nm/Gx/QPK8rfmtjNo5uaTOt8zM+qrMi9oSibh/pN/U7FURKr0I+LVo721RHtLojC52rJlbrx1Cjj
qGUluWhU6qjpS3184/98CgpvnshWkdNVh+WeKrCr67WVOZSo54JylwNz3fgLiZ73Wak9X2aPKUuW
ymTuGEa1QkCDdQnCvsjGxr/3ZAx8cAz9BIM0qi7dWTHExE42iG5+UEGEDxtflmT9HXqBjjXDmaRh
vbwIVJuJI+85X8f2qRdtCXr32/yKR7/EAjItkQeA1lpT0AQj/SYDkb2zhK/bFbQOvMEs3KMvBfNx
/RpVBWEXWJHzdjmMnsHRQQ6ojq9Fvr2BWQOiyvsqmYPSFojnnd2kn9raB9p+wNFiXB7B4CwhJwbU
o1/yxcGpflxXaOXQrIrEtEOGeQxLz4YxtWirPIDnvasmPn+CEnfmgcDzyub/acpNjqupj0mJ1U18
g1iXIdQx8/margHjXCdPzRLLT35LzEDRS5Tg54qPXL8hjlkaNpXiEA2N01Zff+kWeFNwpVKS+Llc
pZHDXAuaoyF9eYFyBbENYxTDQfiJ8GxTpspp/F2mA19s33n9MyLbrDwwg79dq4HanmtuzFlZZjJk
H7sOZZpfq/Xl2EGT2uGZHuniCXmtZHGBnMVWKIkFIHwoZss5PJHtAIf1WD5aspj3Mspl/T32mrUT
JpQgPI9mlbcOh3bWUghwKZBKvkiKxiTFFzpRjLV13YtKyC2ePqzYJYzgCc+MbwXTfY+fxjHV/MHK
1GL23uc8NpNTfsUyCEHqoYey6RVDqhPl0X4R1RB8gddV1dhUiHlLYJ7LKZIa2bYAqDKNmF5tkzTb
l38ecZ304u9y4vsv83GP9Dyl0Kj1VFCLf/GlEU3De8PQO1z1+2EBwHyi13HL61VOoZw8uPMH9JpQ
A6vjQXvVfs0rMW/PANvNflIITCBUhzTvetQb4b0QX1hOe0FVOIVC2sNBWN+Pj8cSx1dKrWoJ2mbN
vMqjXgs6m/ACmzNxbmuvrZLKv6tG/dFX4nb61BJCh10fiWczirX1WA/Oed/JxvPC2UersZrShcxY
YPH2lM6lVfP2MKW7YwsxdQVlHsK27zBbP7tzP9cUZgd6K+ky6HAcKRnPuWxnr6XuD3JvCtZIH+O9
lk12faxG2hVV5nSyFO2uzg92+MuTooJv/Si31/18caRIrfwbbfLfzrDPVxb/q3x3VTkc2EoT08UQ
uE34v8WUtWyuDDW074jiZ2BvWpUi0nt/ipd5333p2EPUqzv0EGY/C7qkUVRA55Oi+g0482fNYpbL
0yQ2awstg+saZlq7AK0bk7h/Dv6xOwGy29eAEjQfN/qM7q/0hS/UDqF1mG+hxUTcnwYlAGNRKujz
NsEb9RIziLPpPOMceu1uUfkLqOG+zZDWKaQa/zbsbmOnhHzg2iKOFn+4zrPQKLyYzvFgq+waoAyF
qjPtrJ2j+8g/leWbjksWCOEhq82xE4GFJw/OrDlvr7DLL6zRN1ayubKsYWTicoHAUQDc6Jl1i61u
JJt7YYFGjMz390kiylGpLsKwo5eYnRUWfJWGsR7cOJMgHR2Qumvjw7zyOQAErw9do2osUBjUIY5i
yCINp/9tVUmcRvUUAAd1MTwU5aclbqsOAq/41bRXSarFUeH5SxiM8eejj7045JxRO6szw1AoIZUX
xvTDzRB4vCbiuXRoXBONusCGZXJ45raQOf08UZ3wcNr3ir0QsxZFBP6J16OegdtecyO2l1MUZXZL
nuzE5sEnpDI5dQMIEjQ0iN+tA3IWSAM9oPF6GkuRaMEGwPkreYb0CzJGa0mjxTHQ8d+iaM2nh/BL
Ls8RAw5YrsjHP+jhNBVD9k/ruQiazxsMTbI2ptz+xI+JHmxKHuDyjl0mBnS3rayIlKCCJ1n+wcTX
XAnBHNmEifAd15THEIHMkdMAXfLZJcXdH8TfRfJwYW9HxwowvYn9iUQhARJv6M8VzHNAT+8t3T/3
+uS8FNNG735OM66p36FSM1b0J79SBobrTaP6Kjy4S95kKTL/qZG23VSZE2ve4RI1vWtbTmQdUVHP
6stjTTb0SM94Fi0WX8vGby+nl+ZIN4F0CfrkBry9PACqOQcYq+KzE+kOQYCtMwgtAYKpd5794mf0
2WIZoyAqlbxHmnc/w1n/SFRdEbN6eTFq+DtZJw09PwZ+afxIJVAjRSDv6Zt8s6u0YOmr+xUhvd7h
dWXML6uJJYkc+Lj7UtymbGvo9txjB6or2k0OozE6opsXsMcO9HEkMLne4yDPI959JoJUmxCpjlx5
90O6IHmz0HknEJAkGkojamD4oODbVa0Kkq73qExca+HSJkbsabXFey6QaHrcHCvf3kbC0Sv5ayaD
pauIuc4KOkXFz68F6Rly/cxy9LFD3VfcMVXvnOzsUGhSmVTPo6yRj94dN+YLdZ5rD103lhPWdQAw
ey5j+YRTvJ6SrT6ZJZDVSZ8S+K3pIvNu0qNr/M93Ua+UnguU/1eveFKIsVkEhrMF1a3+KUXELNHW
B6/U9p+dSZ10oJr+Yva566XyuV8fBvw//afM0yzAVSMDetabRcPYlrQeuqWlgXawNH+ZsCwckz9j
XhnbwjAnRul7vGsExMBJaPgaW0aaOyS8X+Oy4lfPh3XkZKG7asZWh2upqjbDSUNSRLfWf3PXU19N
Y37C83EAgNiy0+njnVoNjr07uCAVOY66DHzYniApcqrT9YV01kW0W6okNASnexT7+EiGUAfg4+yu
6VEyHlYXf532NFKWxHhKkOzoT9Vt9JgQCYIxqDbWyjhrxRU+WTAIkt7AuhxFgFkxB9BW1wHhMDrQ
fKspGb+f8cQfUgq5Tn4gVAIUxnikZPrb+WkNNvj5Z/dV+6tzRDMW7n93Rm8AXaGhmTINHlftQp0h
cq22LuiWqUFU0Lw/q+Cx0E03DjjJWgsxbTwr7kOCtcYEcZkgidck2AnrgbC6NAJb3RD+dOCQmSU5
mt4l078jpx2IQ7ux+Uqyh3bGSPJEYcmvwgcg6CJ0Ca8jZphtQyO3FmKjPRMPWFKBx4KkdskvFgNT
NdrGtiykRzp41Edp3of5Y8lHfZpgt/+1GgqbdmBdxRMsNWbV1iAazP05vzl2Ro7WOVVHAUwa1449
0Dcs0YqB/hqAXFBvSUZHKmjPexY83W3ARBAj0eVoo8IBh+KGjAMBJrBcpFUZrJTH0c8Rgp545aaJ
BLDdMlFbB1TLvqTfGzj48ZlCh/Gy0Lo5JMKcYdKjOQ/DGQBnOyXAJz5dw2rAwezHWF05n+tnRuof
SYqDRKZNQmFXq8QaQwLMYPj/63N9qtD1SCOl1XE6KNBkMPrJj1xSp+7H6kWQiJ4zLcQ/OR/ldpZV
kHt1jkHnFmGU9xqn8ncZtIiTJyvN6ssB7DHfU2QaHo/2fh4TvqtYDRGsENekfkt8SYqO+PaCIvz5
aBgNMPXPIesdLb2vKGppBrpJoZVSObQzfK2XuzF8QdDT2cxZysUkCx01mbfdnVou7oMe6Sz5TCPd
iPnqVKTkaTOg5lrDY895bJxLRbFdI1jj16fNGuzJLt10rDh1DgeGd2zbwYm6dxpHkBRey8p1Rg9h
VyYh2HPB6KirMKwhWUcnQG3FBntG/wHbH5aFMHnCHTQNk9oG1adA6dChEprG3CKMHaLDQyFXXDw2
McAx3aXLWpv9vDs0q2t7kFWsJbR0A/jsWBjJKCstNwCvloMBAa5yYCUJ8xQUKZ/OjFQeii+6xoSI
XAL4566oxKY8NbK4OUy09A2GcpvMC2GHvxBi3+OOhfhzPo2Vng0lhEUwWlGE4UfWxL19Y8iOPWMI
UPunY2YMtR9bHuotsB2I/75kabg2vgsMBpreYLCsg+nQVotxXEusyjJPCrp9x1NLBVzKpeEC2yAT
x6Jmv88S0rbJbb3VR3/cn8L/fQ46bgqOUe6/a3PXKCoNCJfO/KKiG8AWMPZA15UQaIREyNLpft8x
Zjo3X9KrwannN4SRvzHzILC8VU1YdtV/oGM07p9sZVsmxqHIOQva8k8qJcYdjtmWiDDJPdFC467P
+ls+uqSbvbo1RvBkF8A+AN9n9hJKPiD/MeMD4NO6o6VC/4FMxLpBPK3fn8QmSTV7TwSRroZYYLhu
rmQuul59OZ2S3bqULI7uVr5qm/LcMpsitMfGvE83sr0FpAMHIHTpbZOdtAyDEGluNoBOTPfpqx/Z
TykybAbnW3jIIidm9VlLmMMmhMR/tZyE7mfJcsdmcBQuThibhIwYZ36JDkPzRILYCVj2sJimw6U0
IPz1P3KLMpB5B0W7BQLIa3dlOvQfO5smFpmyBXtKnf60nvDzKa5u72D210uNG1Wn97/F3HEywNlD
BjFKTwBN6IhtlTDrtEd72Q158xFqEfMqk6VJinbG5fJMG9YBWG125nDR56k4Mmz8LPyz56HAi9fu
qfEPzWO7Un9xE9GnI1fbtMI5y2atuhK1bOO4whGTsQ5j3tC/evRGfYHyeTyZ5hp5VA7TZPZXJsfn
iNAGl8dvkJQ5hBjM/DBvj95ofuScEDTpj6JIU9/9LCdYm4Lr2KtCcJvjjcnMqnZdeO6aQD27pBGK
cFQfC/mts3/FgEV7Xbh6v0wXR8W+VCB60X2Q+C5Oaf74x0z1/RhFym8jNd2KajcqgiqVkxSecD66
osmxOAJjZW4ukUCCHTVg52DTU8cOrV9+cQHO/zjBG3kKUPs+/UY5pyraF6OmhgMEhKuh7cNU65Qn
A5H3zAB2HfHMDOU4nNnVgK2N1E6+Ih6SDoY8QW+CQZfSpFy9IV+1rCMtdqdIMuNqdfgutF6B2rKL
Pqjh2zzSn87GB0O8e1sADyArgBBAbb1Ghaexkhzri5dgF0uLh4wQ71hJ5u+QQ/A/cMnxfMGM9h+4
3qdQxaokTWUqemnBGZhC7Da/vJmED/0nBKxX6rGdQyGh8bpmXIUIZ4y9nXSarISx+Hszjpx/5Rff
eK0ao0UyjUJbBgqUkonwInMgshldiBe/nQKk+HVWngMxxiN3vscNdCNGsi2SblsUUDDaRAU0yDOg
wMPwykWLVcrBPDhHJmlahAH8LZ19UQ1+VV4e9LXghz9PK26XNaU+LnVAo06NJqD3EjxrdmliKphS
9YGZpsN80J7RSIwC6IXLRmnl2gF321Z07SpjYbPwac28VMsDHrWEtfCASqsdZzeTi84IuDy0Tvem
i2I2+5lhcx5xD2q2QkD+sdDhyrp7f5CfVdZ+WIV3FrUUgCdcgskaidrU8rgKFj2uwaSQIeQ+WeWx
8OCPiEjBw4rhprKOr2qTvrxRzlTogFQC8+fIhrbJ47B+rz3zcZG2ZIqx4XjTxHMYU/iegr+biUa2
OC+2wc2MY3rfcDm3K043AFcGIkyxuAuuWZsvJ1Z2vslb423W+8tOA9v0LCd5BKxN5N7y0j7Mz4Wo
Hw9wW9z7VNT84jLBZOPX4Lg4K9F8ZoueuGEhUUowL9bk9qFn/4QvHvA0DQtWpdvx3+n1XpWhS4OY
gAllVz/29gBDwOI3k9yNoNFd/fg5PYmEIzaQIKrpJ973NRITGny7xqvVrvpjzKHT5mCPfUhdmK4R
ODior2aLQQXMUTlGe/Y1dcI2Qf0CF8xUPgUIv6S1a2oKzFLUMMfH28YN1vOKl/hrZE+h5RbRYcJL
pTkBm9y3O+L2Bh6CWoPAkUQjevlHuHRwL86mZ+DGAo4RhK2iR0SMLEXCyucppn4FsIT3VZyCXVGy
8oJAW0jpfufiH77e6cIPBkxHzfF2dIDn8OJcIFWKEmNU4lirgFn507d04lPZMImhK7eZ5SOQfuXp
9HWgGZBl8uJYopBBGfvZDs2dPodeYsDDk+W2Ohu105Fx3L9/pkwyYjERteyKqeqVBMau3iJi9/LO
bfXNPEAlDjT3fDL3Wk8rvnqr/EzoECNE4f743+QzKIa8zxskj3Z9OnVQBSjeBoINUyzztWVBkKYv
M/m7rmZhJdPf8qj6dVVW69GIXnJ2l9sXd7M3RJeePlT117UySOdjb0UW+nQk8EZo9hsgQEOpETtf
rwkLb6295PllNQNJhW1H2tDTXd0QN8xLG1UkQXo2olKTLKjdrny9TpbK3V/NosrHHc2U1esGI1oc
YC4SfIVkS68YY+sNKr/+r9VBi/QVBZVjZmwP/ffbxWFSsoEC0ToZra7SelPHhAtQWVn5/kW4VQU4
Kpi8cfhdsizcouY+RvCTCNJKWEk/U8X06ZBba5C9EEgEASQwB9/pfL3C8F3qvdsvFB+QZW2RRA7W
D9I2kzzBx0HUcgBcDFpZMwxB2NNZOw7F+z0BklfhphNLZU3gexD16TWlh0kDufhHVsO0fNHodYR1
BiNME84phrpF5YX3ticL8J34mpTxDlrdV7prxFSOcSz8vXQ+98xkukw3sDuJEv7LVaGoGMdZ/a6+
IPkc5vgrZErVeGo4DbqYIjanhwGmbNTYs4oLjLlZBhw9kZryqnyhk6iimEsAwDX7rmzuH5eRAuI4
aoMu2onHEAueoNN7DE+mUct/nWTYffui5k3k79BeNvA4CbsWGyNEv36Kk1VrhXmdBxVlL1snbxd6
bIg6m6MXlcUTfIIrCWdGGsTQYruB1yOZzeJSoIX6R1JJai4UgDfl7Y8daPCBTqLz6hBOznRly8xl
shtshJBLdGlGS5aanNin8TxdiQf8hWtdr+vSHNbMarowtvEsjRi3CQpliYgzcg2AT14BHt7qAjXf
VZ8mQ76HptT9ucSW6O9Hd9Is86GwJdODTSPFEZAJrZvOyQy7CvboD0hasQY7ZS2trEG/98MFCFUK
oufYOxp/sUyt834zVrvBPPYRF46IU+K+y8YKP2g4S6eSdSbs1tXLt7CPQK2i8g4IICEcBEqb3dmU
YFmRKegrimf+OC2H16fAD21Lg3dFWBDL91bjqYye7ov/ZS2EpesOFh8P9nYua2STx+EHkkzqH4xj
YfbeNtomfuVcLi5MoLHyrXxaouOvbRUWjROq9v4Nbjnbd8TZ/5PiG1qBOp0vj7wUu+lm62feRYmD
9a8+upYEuprrEPDJN05Ucnkr/pdXRLR7q9+vBo6cw1XZBsYNIGIWltv4oJ1kb15/YT3LmbZB2H44
xyf7lEbqA1Ijdidr7DpWPfq+rdDgzALYtJ8x0PjKFpnm8YrUSjiNZ4R/efr3NPmlelskst8cAJHb
Ogd0iQGzZe6M7wDh8VH3grLMcQt240XqwdeAt/9VxEl4tK3XFcEDZ4h8T734lle32q6vKrrXazd4
2fuPrrTjiq0+AO+IRbu7uep4VIvceXDvRIor29vgFBZaI6MotnjvJPmhbu1ubCmb83O//74Vfp3s
NNPfTg6e0KlIUtZSgC3ECvTPpqwYlOlFYDJkJCVnQWRmb94Z3aHOzId0bSZQATNBCoxFCo+dWvUv
TM/jKI6Zw8vUvgQQdZjwcNxb/vhRs4zGv0B65z64DBoOkR9SoFUR9ve5jdoONI+WRgl6u1AdAkPw
fcVupgTBN/UtXHnAMj5dw3+f4vJz7WSZ906pXdzR0LKxE6gt0N6BvNBY3pUE5BjEqvH1YOd5YXb1
W3z2OyCUSxSKkFtpHunkybjjLT0koErBIdnxdlMHL+rNqz0VsYtAqy9+A6XJhRlqzypNI2UPgQgt
6n3epzKKs3Cv0fknYk5tptyJnDmPGjIF4gKKMr31+yNBwlcVJOXD3aMLSBlehOnFQKrxb2DariHf
PEN0oobLvU+Qs3C/6+Hp7vyqm43gJSpCx3VjzGuww/Bj5xBe7BqUcCDtjz0agbLImD5+5p/Bdz7O
Cb2aj+qCctQr0XxSnR6Ufd7WfZ1L2iQaXTVQsJL5QnQNo0YHYdB8jqxYktHrEpjAsbeLQxplfvXI
vTL4edNwdf/2MBYAFkm99LhQOfL3MpaGUJbh5i65J7kGoTx/Wl0cgxHyzphKyuVWdbIopOt2dB9F
WuhFJZi4QSSjkuQEWOoLfSNIJnRFpzUtaMQQy6Urt/aLnWz5vIOlAYChahvUQjfd3o918E5OJGWK
P4w0L0udAFdxulUGnbThCLChaUl4BqqMRxLXUagcx53Ii/OqWo8KzOjlJjE1ol6lT7nqIvqxF9+R
22c+n5bVwIsM02ZdqHLv1AI5g14WNXGPpTP+D5SebKVWH8REQbY5fdtEW7JmBTxBWQa2OT5gOMdU
F6fPCBngreM/5diJvsGINeGUj4UFdwaJCZWoBRwo4WCRmKfSLPDZCUva4eDUn6xLO2SZICaGZiqk
W9fcUMlQezvXKLoOvZXalu/seHiaQXdGSpt+qvmZcFXbqSNZm6lBB3+dea4k62NqyZPMGLl3vNQh
Bgtv7yHpujaZhZwHSHkJdQCsnyLak6gnP1+tEdrXrJQcyFUDuXw+Adf67vR4k5bKkwpbUGI0I4HF
Vd6B55BxzBRO+8W8V/D5zn8gwZJsr+gwB9uFVTRRBBnwpLeFl9K/JAvklbLYk7PH6MheUU1mlFmR
0mYKpnQPAQhStAT16OCGTt4qUDipO4fgHWID7s5ToZC0HSVN/eGzgHJOrAI7AZpRxGvvDbBP6T/G
S4PLZ1s/W7DM/ofDw4+AlM3vUKHCrFEmEeUvCDGUjgONo/Q7dtxp6YgK2CMQVuzc2FTjLtlItDYi
MEdHEaBpvdFg820diGKmYOo5T86g5skFsWVasAkHuLa0vlOEfDB19RC1JKFUqEguR5N9GsVk3c6p
FoWGagj79P4Y9rXYdpPSgzmpZ5j4Gyk1vMslUU2SRzOCGiTSpqSlLMIygAjuN7rLYIa2fhVBR8I8
SgQp8Zfoh6Oxkm0Qp7hXuvOZI1IPxixssPAr6kO/C1PCV3358GeWJ9W3XgWbgyGt0mYZ9yBNq0D9
ajJZ7xGWQtBPWgl05KC2NTNEsO7nEl1nVPFgjAonqGCdweP13l/HPlKn7cz6pW0hX1WhEHJPBAZA
TEdd888yOeXZeS5HJJAweSpKBG3rzaCGnMt7RmscM7qfhhuvy226I60roa8M4JLDgqVDEi1ZvN2r
o3FLASkdgjPqYtj/YD2Tz8s/4SJFOCC/zZtlm6ilvUY8jesYx86MeAqPsIHjiV31trY2jOO6hHMX
VcN1j5GECcW9rCg3uMiVfvwIvyzn+u7QB+2Ph2710gUmGqjKJj0A5LDHsWjcqoURcxZ9afaZIB7K
F5h6nJXZ3wKmjc9WL3K5gVdEG1aVG7hj498bgSA+MbVaeQhB9IxXl64XtV2Vt1DVQJzdsc4tHXsW
aqwcvgzL2ZsWvwDa7xsh0agod2Pbb61NeUU5Ir11ng21dXnXi3WpIGHwguVBaAW8QKMMrEyVTXpd
nNiuQFBKkX/PqqXRus4LbhTBM8Sv7xAK+GOsPrZYCj6FbOyvO1v2nXKxGRmw1dpfakCIZf4VSetN
iHpvEHtYNIg8kaAIzsqZYDCWuapOS6kdL0EnAxSlX3sLVTfvaTn14Y4qjVc4B4cHPz2OhhdKCq4W
0j1KZreJw4S8KPrfIccXtfizoMSqReFL88m6U4LuHyDF2qyy/NZprevq7/xHD3KYU+pzDYEouiMm
9HFX+XkxxGeUxlrQZazkLF6xWj/WVPbF3kxwDa62OlyoXt98aDlnQCip9SUpww06aCxGZK57Lb7G
BagZ34s7tIBqmRMZKmPrYjh+eTO9hKjZqks4fEjSqDy4pNcrput019j7nO6nHtxUtgSK+NFaA8N8
6xYkwidxIrd2CdsSL/oPgERF/Sigqd8Fg7vuJ0VWJSaH1x6xNl0DLaSvH6NqPqjVi8ZUgd7JcwB9
v8CNfMF4g9Msb3oENPYZu1OetybFtYTSUfc/k/Zdyh7kWb/lSZn0KBOlUPWZ23DrwpEoEDA6dz6I
Ru1ojUquwz3qj02Fgn/feJuNTivoM63lorwnXLB1Sa8+ji8AZcFvdw02p8UjE/bbEu6AgQN1GOap
a2IEPDbIVjPnFrrvMfDrSh8nux0Kvhx0J1RuAoRDCXUc5NtsSFSW7Uh+Cy+plzcjk8t2A77zkx2t
vRQ9FRXKR1MHBNlsNsl4czYg3arXNFIyZXxJZpWZWhWe1A0/1CgNupK9yXxZZxL9FLJ3VnNjyAZm
yLbSHTDFYk9J7XpsyUqKY3NWvOOQZ2HlsbfjXovpDlQ/IOeyBb+TkOxGUTIN+nlzxqUN5Req28KG
jTV6qSnI/WMADgelIhtp9giFtNdNe4Hs9J4JlZvk30WswG2q9/RQb/T+H6omiiIf7qzY4BNSNz5Z
mQpWXb0OH/jZM7Y2exiI+V3JIhvqadI8U5xAVqgqOP0t6V1IJVSpi7j61G6HyU2q6HqrgEwFK2lH
NbAGBetaFpD5QW/6ALE/MscYeSVFKiIRtTvYCk5M9MmKvT5IO8dtoLSwO6jX4H0x2erIRvy/UQAg
EWNS4+FlAuGkkdmDv7dsM0eJq6nEe4lwkod1479v3vmQOCnnriAofQdE0U2ni1d5gCMyOIGeALXn
lLKi7F+NnzmJda35C75O3dEHG3twD82MO8i1YgWZDA5kMhIEYntrn0Pvn9ay7ZatYDEFbftz86Ue
W1QoADIheWFhpntiJa/wtDo9J7d9lI5+btKWjblZ+F4WGdr5KicXRRuKWyCAyUqt6e84iOOMACCl
5YTtwTaIzvFpDKSQrz/KzO7tipY0Es6a/Ra0oG8HOk4JV/2mHj5PCgv95QAhOxI82u7ZxLQCWN5Z
x/yA0PHYWM8Rj8GDiWXzmIbdio34moW3i5SfxFIpSmWQ+FsDVzUCHF6vfLatUTM6JWiTPpTsyuf6
10Ku7OBDc6TJgQ976gx6JY9zpQMoJN6Dg1fdrESAHrbSzLuwRjzXZHk84+7OQsD6TPlLcR1Bhc0l
y191RWWKkiwet+3rrrzPFeS+Xsur37Oa7TzuLRNZPN4342G2O0uLBh/leZrBcokjc+N43m43J5JY
BcecZ0YxZnqM+NNM8FlqApHH0y39De41Yspu7BI/Xtek8W8zQ/2i3RmBZh+rggAAj2TTbFFeNgMU
/GMM2yMo8YzaAlnw9ykbS7OevF9qZpd9lOgpPlxYEbvnbjWkbIW/60f4YSkxqfKXZ7FGD+qC6xxk
I+gnVO4YzqKxG5pUdRdlRgUqnqI6CRATw/GUlnH5J/ghGctoNxvhI7NNYJqQSVSq6KwSgMFF5ha4
EtTr8loicYcItHNkf13zkD5D1ZfQz3I/Ef3InMz9cKv50LrmN6c+psB2zPFpdHuEOAvsgx6z37bQ
5hV1JgIsOfnj6AxaE6cNyAHbyuOSRHHZsqaPfJssAje3Rv+HCeFTwplIaWcmR8X8FxbYE8YHRlIy
GMJSqGwGXXyZ37UQ6A3JxGV6Ncic/PFb4rIiSlIqMGdK7dHpb2zy2LPRL7tOV+OA/kXVAOQabvvd
3Gj4yJxkc/EVJD0emxWe81LT0cxKBb4jeiuqgV/0dpYaF5sdZdSZ0phw2+gtbIJPMtaN4kf5NCpm
ELXqsh0SUtL6rp/NpxR5FZPbNVbFLhPT/loDEoyeJm/hzCpmr3jsYr2d3m1aDlKy3NMvHe+WIQ0Q
gleEZ3DWyLBfhMij3cPKflwT0lh0oiCDkf5DOnnuBg4sr3l1Y0TEdFChBXzW3Iow7qzDxCaHxtA7
YuDPZIaqGfORz1EBza+aQ3FLqxTGfhXmi85HJan11/FfmFULUHU43xubmJhxV/3eflp9s8+ECAS4
COqn8mWxSJYa7dt7VxFo9u8uiVbPQdv3+o5RSuZIUfvNdD34VRH1YrccljhDVo6alGwlruB0w+Y+
u/18Y5rCLsWFKEjWl+tU1qQ53kS5bglinergUPHRJApvS+E7XjPr7fw2Q4H6tvd8IT1fgfWGyaRq
8Aj3Hd3WrR1wkNz3QdrSV/09RitdPk4Z2ZZicEJKr93aM7NpVzLUr0+TiP9vuJGn8PoTfCn/btgc
nhF1fcc7mg5uhVltJ63ZNqmYirUsxq8vMaUAyqFIVJBnYpAz3g7n9QElisyiW3rNStN04OsUCrQ4
V+VC4V6mhQ7PYgTn5a0+XZb55NJFQ4P50alXc+LCqD35Yl5bALPRqisIuHc2R1P9pmb/aC1E4oPc
si4X361SXybn+tuhnSQXf8JGClqplBXkSOeEaNbliL0tun0061uAjd8d1YW7mnWo24JtKR8yxstp
8vStQEhY1ZglMpo4SGb223Uf1ugbJH3vYv7s2vQgzBe5JvD1hBylE125c+qFOCxQ0+X7CdVKppVX
dv1t/v6FVDtX0/onWBLFayhehFRmfzBVyuQQMVp6gT1Jqrc1blRFk2c4kjgQ8LnT0wiQHoogysK7
rCin/cYQjQD/U4XmSTcMBvdBlgkOHYauVZQ2NH1tSpBj04V0Fcj5CepJ77VrOOgbgJs2WFeIo1/y
Sp6d9Se23CtUJSt56Rd9hEITqHf9tJMyQ/EzLWdTTxHGlFRFIzcU4VEAx9CYNXPccjYsXeT26XWA
Ctstd3rxuJTGupQefnv9udVtzrqf2vWRFTE3swIFsgClyBzP65JRzk7mEjH8FTZvldvr0z1ZzfhH
lFP3+QlOURUQ1X8Z+0R2gquMa88otlSbsUFXt8M4Zoa9nNsCVfHh7ASZ60hG4gSovHD3xMNDVNr1
/ZN79vWHI1voL0cG+zetCPdJWm+5AccNK0s6JiglnB9ZjViSW1Zd+ToW4oSC+vjEse0Z0Deo/SV9
7f9jaUNKrTJw6rshrCgpoBjDaxxahctdTNsbzhRUy9LVUUFh/phDb7lCrITcQz2XvMRZ3W0d4SiB
TrwykEhIDLzGtGRwauZmk2ikI/cF8B0nSAr6UVnHly4YpElWB19xCqhP674Tt+iEQpEMJpWGO56/
q4VJS2l5T9vsZ6rrNqiCCBU72EiWzJTD7F4wENgM/tiTnUuE4jKr8dhdQxnujeJ8wS0Dlmu1ooMy
n9bzpgZgJxuFvG03d8lM7emsxzcXBDknpsEmEL2VGH3OWmde/bOKvTi14yM1CLSEmK1a/JG4T+Ms
T+L7lcvbl3wFDbCyErjubNx33KRJaMWHHzQJNq7qPjo07zrf3iWWkNRJsHIFkoz2SzwKMPKSDb4H
FpsjgsrbPKFKMPq4pmRi5O41TaQec7cq6oRsw/MlXP+OBRl4t+4qhwnsa/p6TrIsWWySdrws1hs2
IGDXIjyo/CxUfo4cCuO6WACggnQxYwZSr2MRUH70ztSYDtXiqtz+wglG467CEr3yp4guoaoh2qg1
ykboRN+SzWQG3Kqxjw0cMiabonMglLhBsGMdQ9QtDpz+YT+riMfWBuaUJ9fdojNSBFWg1zLp+eca
XNXN5THVV3fgIh532riOAi4A8JpABxqK7Elb61+RMfK9DCVYBCbBj8gwdssH6of3hyqrhqn3EHEp
vVXtGaB1byTVHgGTHg+EPO5HrD68dfSp/ew4AQLQA5QjjpQLjvJq4ZKa6SKKo6rTLzcWj86GBQI4
H1qSrEWDapBZhJZEZbfJpqmLmU/OsNIlQi6uZMob2L8UMTLNEOlFUPlTwx6/EIQHFeEjR7RebKpt
lt3vvOllbkhJ2IUK0FkiZZ1pJ/2sUVNs/MvSkmpPINEjelh0QOIjj+z4tw3WMtIRqjjDS29x5g9l
Cn1EoEl/wfJ9RbnLchMxNSabm7hAtJxdB3aQRb0R/sbqzOChCeBvvC6JdiqtsIX4eC+/GmK/MLzA
JR9b1u/BftFluiPTWVIERXXTw8N8T0AL2ds2rI8UNV+PpTnQGElWCkg3I8AlnwRvPzolFrEFrIMW
frnOGbUHBRnT4qidNyHxlEqmW3Ejx965G7WG2D/a6XLuwMgQrqN9I9qBkMreHlPvo+cBUMneKXVP
srRqOHlpF0D6E8lG1zvE4xc6z96XJT5xLYmo08ulZ4gmkPuTGT6e4qpKC1Ij+OQwstt9yKZSUnN1
nfn/W8uB2KDk3uuKUS6SFjaFyWPSoEiDy7cDXl3da6tVvOS7uXNHkbRSSHOJ2HE0tS0Te490BoG4
RzBEzo6XoFA2bsBB9LiJoZCIAJhoyrMpOYMe0ERXkXXpdy0wMqZnNQ1bFXmFIsQNlU/qmsIep5wy
vWCSWo+EGWA/dkOf4zl2BKmByxknrq3jIovBdf0UIzNfl+EIRDSs26FC9cQzxyMYeic0d1pZFnX9
ANKfzJ2H+JoTt4+lQAQnbQnsbd1AV5CqZPyI9AYkfKgvvTWH2TeY+TaRsZUJBV8w1QMajlHQO/U+
aZkf84zQ/5xShbGjnXHGgZ466erzrRWwwJBrnXrAPkCYF5b1CPK/UkwScbDqq0YmuJHJ6ynzHtu7
CkeAUKvYym+uloW8iVMWj0vrAh8e/3827Y1UF2XaKQ3E91JwGYMW2uOHAWKxqKmQawJLu5fB91ua
sJXf+EWGUrMcu73/kW6SvrmgpmOpkjc3Myw4dG3XXd1M9vHtkwo7eSgcD1MtKQPrg8EjaMsz2wkG
d6ohoXeqZLm85o5v3vsRXzeUUEOZc8IAzYjd57orzUsIGIteZrDe4gIFvsmhdg+k9SIxpdxTD9zx
ZFOZ/u1u22eF4WEwFKExxDW6vnay4WXUolyyQBqMD1GpR9L3ApmOaNf7X8/VSyl63ruO/AmtISVA
V59/ccjGIk7wA171ZDzGPqY+Y6FGHcQdAp9oNc2pa7kMFSWC0ovqHdFe+f7D3ow2vaxznce0V3XS
PjZIJPvzV30tAh+ZEyJ6oOQCbcpEfUEK9ZdzZdDPjQACRQEtC3fYJ6qoL4JzD1MvOYivYIPpqrma
UM7C/lVvu7gsF11sA7MqGb9r0dO/xvvHg9xFjaPSoIcfFOs1/jHDhN5iIkk1p+cpeWleD4YHvwlw
YDUx/pZQgVWzay6gX/vqleEUIPeNGwNE/E9GQrp4q5LROueXSuVhhR0Q7iWqsePx8kmJEUnJwgKi
7o3WZ+B1thWiyFZ/CSSiWZLuvr2YgEQkOM6+si9mHuwPrQnf/NCVDBb+IpPYGm/pIVfhqHpMP1oU
0UE9aPe1v+EP5/9s1tVPkuh/CQkfZXPGGy4Te08B7S0OG776Ilz9LjQCIxx0bO6jE+KUVKWsp3qd
CGcClPfuXmYBpRzYGXsWqYLr8dVOkQfS/n5KZU3udJJGyMJ9NkgvuOtwIo7xRYbJAVYrFCZi5bJA
nYwBlcLcs4jwv4HH7nUimP+zV4cSp4Qx8TROTahK1E2N9Rzn5EORWVAgPfusLct12YnB99s/OFbA
00jFLyb6hPUYELfw+RS+FRzeCQO7LYne6Io8xIMKM4Z6HyTCqksbRCcbc+W1ngD1l3WFZtBhI3EJ
9YEICfU/dEAWoEu6CBxVYyGnADziYK4AY2wwtdcYZ1s7ZHX8xy3W99tr5ggWNvxJOId+E2+N3VVX
xOaDk0YEo1DIRzoXLpO6NjTpo7QDQMXmyc9z5vEH8yN8aPFsGKPWG+j+gioKtVC8pGLh9Ug0WxIA
NGOdW6jNKsqlA/W5XLMV4mPVj/TUl9SL+sXjSsjSp+2EwoNoGY9N1ZJdkD6gK0Ch4nMUhlOnLNk5
OZgnivNAAFXLK6GWxsboovNQIcNgf010Rpzen9Fkfh4sU+fiC5Meg2TubemPtQgo9dfA/cZ0n+I6
9oslcPUeaS3d583BMHbTZJkH0/E79wrPLPcYxSSBWX5cBETdF+m6RkYVpTeHBF3X9mK3INPM2jJV
31bjkV3BNsR8E8HJZOdgsiFaRPwloezY5OOh0bS3q4N22fPGnY/PdlcZm3rDK9YZO7HhuvAMm5E7
LtM4Te98Xl++iy6MNFs6smVEN3RFqYAuoPWi+XnisN1bunMUCiSEcc5pAC1mPDAirNs26zb6IRWN
KJRynJIvgsSi4m3kI4iA2GXVaMnBMwFImnwLVkABNMmTqtrIC4xZShX3lpAf+LCFGn1lkVlFk35r
SMQ8cDTBxEl+iaT5UAgkvz2g1x2oV0jDSJjLeJrUglkmg8cWyWyY0hL1GGafRypzgX1PdUsVbIWx
wYsetZH0FlXkI7LHj0CSqCf9DGe8aAn2zMQhFAQHd+uAP9MkMFa/xccQeeKUdpdQcwLsIWvWdYyF
7kffCqhFAGWSLaRjM0wRYo/QlC1vtBVPY9DhEO4H48pH+milqfPI4p/qcq4Tjb0t5jZ6yVxQVa++
IhWDycu+i58oHJhF1qylnTSxJNe8bBb1RUCltfoibxVR56xPqWvWEbiU7HqOYEhSOMB0xC3y1shk
CMhNYPWY9FkyYK57HVSt+P5UdDrwfkKONAf3a7FPKxID76dV54l5zeqKJe8vBIVJgllUUgd9PQDP
SqQ/8YWARH3cNpqlUcDPeEUuOlYdzOrUWAiKG+ZzW4VeeNdzfE6dDN9iRIOINm7PLojYCf0wxpqK
1XW3E8RlzCw67k2Tfrr0YoCsrBn7mT7j4MP1jgJP8j3QOphugPLQPamEc5O0cOzs0whZkMUn+FP0
RJ68mIR0yOhFE7K/pALKMTI4Ti+eaIy8/MvPf4lWuNwZDMNjtgafRNfmZwbH9x3OxjodwepZCYqd
Ou+USSTzuOvVPc7v4Mxm1WOboHhgSbmThF9UHQNNDSHJvkZmmlWTmpjJKrE9+n0o3gSkq3M6PXMG
jFcnZbOdjSzRF/G1JsnP3N83EYktmX3ywYtSK+0BFZWaEZX3zXrq08m4Oil8d10/ypiuX4RI2y9v
1+bJx+k8BJPqGrVkH6zj4asX34ZALGVTQ3jPa6zRQBvYCq2S0Xa2rE6hhdn4FQcLmQGo/jAraP6X
sMnHmlHMgHYOoTWdlAWepuI/NtJLBtv2sny+5ecqkoapdqtNfGCewWIDJ3R/YqBH8tlpjfH0vYAK
TeXWGNIWUeOBHfcEAM7otFEghn/pG/hNYLq023VTfjIFmdcSx7NLGRzyoXq0OkRlfVHYB1w1QtKf
DeQtt7LqZ5MjDQ/oYmsxY1OAqGbrOlvPkyKJW/tFvzmoenx3QPfhMZP2BMTkOh8UOg8gpF4e3Ow4
SJj7CuzTctH8V9V2V80mtLiVc0d4T5iApMyk1miE+IIKkQ9x98Ve0keTX1wuFI2E0BIe4dCtFZWu
74iN5wcpRpDoiF7QCizFreHcAQGsX4H4outHQozZbaahG/hWM1aumJfmM1R/MFJDv/kQWGuFHssX
UEsBx0LbV9XOA/JgGqTK0QOouANkrTDvQVQDJoRpf5Pz75cSSUPMGTOV7BRzVGaCumsvq504bszh
X7w1cbs188cJ+WCEtDjR/UuoBRf36eftoc8Z0GmZ6fT/1FVMy5YQJdnaVm2oQ4hahowII3jl/ZOt
xgD3wewaQdjX8g56hWH7K1BEVzkuzgOdtb+aR8cjfYfHAhG8eX/tn1oa+99QBk/oF+gmqUTfA1oI
R56QtPtskLwd0f/UkkJWH8Un5LFDFqC0EmdslV0410x53LtXSzesO8mpQgYpejH2wetz3hbR9M/N
w3jxIMa+seUOSrCyv1IsIhewC896WQ7zCObSE0Nt4FCCXjlLQ/Bv3s14peDMU2h2BSdIVgHVZCbQ
NtJe8Vstq8L/18opA3FNu5e5l2GFQMFnxfJ8ChwE8LG5ic732qP8NQPwDSI4EhNW22xULtwt8+VD
CMmg1m1P/XfBXoblnStqXE5h1qNWEoWZhu0CWo4hyAZRKbsY/CcKibYbQHH2hP30qDAjaeqby9Vl
9evQScDrVT+gZPCDof19xBhJk8VWdijiSpVjolIo/y0UtyCvDPwLxlK/xFzvr/0oLCKASnYIatEs
BAAV9Wy8gRl9blDemcdGfa2g7vHa3Do3OfL2odph9MJ+Yz8ioGOwc151/wXhASw/9z/ai0IUH81Y
/7E/y1Xb+4xfAPTUFtXAhkNiMscrb/k+JMcoyRabppb/tzw7d4Q1RrIQx7fc4gdZvSdgNlv9RDlL
oeF8VIGaxm2ubML+vBwtNpeenI8uRDXA3nR9ioKbt15MX4K74E5vpEf5QNTCya3KEiK7S1uDV8ML
yfn64OtmfxqNO/FkuuMY83cA007WiHuRA2BBrRmeschFdrndx3j4qAdQxtl3Y9UDSEGaUieN7mOW
KD/Knhm8Agfokha9e4ovUC13cImD9SCTTe3LonG0peDxI9HOxvp+Rcwx/LVdHjuI9asSgUj2RPk8
9gyC5MkFi31iu12iDQ5nSoFc7UaQOKFMdZigwMwfXOjG49pz87yvWaXsH4KfcCBEmfobqx2S8Bpo
y9Wf+AP1ep82cK+O4bGWPfLBlLcqSqQi4lFzIO2g9HjgEtgpWKKaFwf/UG85dhrqst3Y7wk24+cq
sW4T4VKTGchHmOWF0iW9YcaoaYdwtSJfZgFbVanW8dzXznPfJa9XynOmR5MAMllYZ+2/WknmtRzi
mpwkSb5G/rko6Umogj6+9d6FR4fxQ/rN2UlF0+9Ajjzzh8HOX6r+Rxp5SGrc6xMEPzc+EdpKbaRr
Pht1ztn2Tc1iZ7lvg/OXd4Fcbeje0KZM3QZFLES6f8xlroYB7ZFll5yD6BM1jyBYiHmrfhw2l9+A
M1XtoagWDgIF90PvpBn248XP0Mz6hiKiP5RLkM1VxNIVmQm9j3YfJcO7f/SCLo8t8lyjG5AHMo/K
LMgHNt4Vu1swHE7em/1Y3b9kWSCUzSq2tB/qzqCalXDmmc8mPj9+IkLrLC8QEL8Xd7bCYO1THB9U
dp2k0W9YqurnL+r2EyiwnLKtEWgAQVWdhFcS0fq2YTY9Q04LyXIxQs3SMghFn/gwRVzORxSUVxr3
QupOK45wHij+IIVA9khJAbzBA8FSyz9RUvesnTNvHPTC1QPq9TmavyKfWJb7sR639iOe/gKr3G9L
7i2wE9VdmrRrgkstQu7i5mvJf9VOyeXN/Q5+0O0SVlqFda8h+GEXEeBYIzZo6BOl1waGbZmDyBSu
rC5X9CreCm2bnrTboeuuh9vKNbCT8v8gyTurA8am2FMkgxbEt+yC304Hf/W7P42V/r7vFqrxptc0
ExEWqPN9EyCl0i9ZekBMv4i3cp0MuFQuIGqZKseloGUYthovMBrpta2PK84cAH3ehP/0MeIehxbH
6SYTZ29MX50xR7YBkG8EwjtSCL6DQgna6QYrOsI4rUcDauyTwQqLVxERdb/jDMmpvAISReTGwukw
Sc5xhb8qOpOU6KDQxnjq6tEAxPnxc61nj91m24I4OrB8oS0kfIiAXDdsDO3WzHWgwUcBf6zqGEmb
b+sERQUvGyox9IdFwjDSJFDKM866u93F5O3fNUQUeo5D3VviiRtS1aXFzMh4Pn6iX6RM5gOvTB0k
PWJIP+u3C6D+K6MSoh6oPjZG0HGk4GnFM1CXm8Cs6INihzZrBzO2gx92DbztsqAKXnYiP69VKcs5
1oL44gMudQVYa0r26nxuvhD6TZFtYWPKK+wnjkfl4JW2IsXfQpmPOXyj3NjUltuQ0SoNWOXcgGBE
RGDDAfXmCcT/xowXsT+cb5NmtSHwWkXxJBKw36mlJRFA2rppKYkLEzlzHL24Mk3/R1qPArEvkc/Q
PIkyjqXwa7+DyQj9Kyjoi6rFlAEU4twT/D3YQFwrU9W1MAmDZ5Kh2VX+Nr56jj0szUkfRUxIVpMX
jd23T2x3UB5j19MzVMWH5f8bQZMtjnUOd+7k2h5aAhnbRkAjn6XV03Dsw27vubPy8COp1ZpMDu+W
ZcY0jfQmAkBqfCrYAneH0Wy448sMOL8jY3h/hAAiRkeJ4hdFHchRl5GPteeYmnMt2wHLfga6oN5e
26+X71uqmYL0024rLMdi6S1uHn8oFKRmuuf5JEpK5sYf95McGQFs0itbisNPTTkOB1yd8lumIcph
l2SueiD9n3EorRN237OuUG00zKmPtuCJ7p9h+lsdECQR+s4nZTmU7FRjwF7RoNKdWbb0YVn5PoXL
nDiM1tLKM5k9uKnW2W2kfDFLk+crkSILU8/97lglKhJF+C4aWvcFs34gTGBk1LmKVXDYzqvCvl4q
pOztVAJ3n39P8PlRCJCELmJIWzgFTBQA6BDedNoe16lOCYjtcSEirrLh0sLg7Wrua9FzbK7Vdwww
AO0up8oLLFTpU99Tr0jEl7qNHqE5cvHpcuqw1i8MW0sbZSPANvg75UVqwAcMAkzkjQ9wrMrxbeDv
4O19Z7NiAaXPUdgYjwwkKxX0EnyiIgEtO4PKDEVtOs8dMob4oYy1bz0AZBOLMEFimzC+caAaT8WI
3R5uxWmAFEqjSYU9UJL5TNFOBJPsQZeQDVrzmXv9bdVWdd8YQOWN4jJysx8EBT/loj3L32RUftcH
VIu1KK+2AAEpkblfKwPzld2o8m3IDCV6YUpE092T3eI2PufHYLiXApyP+mujRZenJcclH0ugoWWN
ek8cowZosHsOtZzTno7SrQop7VVtf1NS/8qrQYYyzthNrgBBFgvT2ky31hm99HV1LPWjKN+H7xBe
EN/E/tVDIFDDsSHNG1i12LmGnlVSnTCprlZgo3w9M0Aa6zj7vIQblDc/26l0qnhTBmjodZy+SiUj
GWtKi4r/alEkhlyVGqbpmyhfoieqnfe+drVmNTRZSPnEdPu8IWqd0oBc4OLS35UGkXjw3mbF6pME
jCSpotMZw0rQK2v8LGp33Pr+xLyDvxvStLz9VRqJQ5ywdzBYc2wCtxG6QXWErJX5aG11/x2rjHvD
wfIqO8mI93jdsoJFjl34sd9CJSAv1FCh6dSe58RFQsZw0ob7iAOtlBj/dKjaK5ZE7ELyAVtS15Xq
/2tX+mJUc1vhQlvT+aPiANFsya9SY4n8cHu1EVTyK2pGJkW8F0Xa0oRnP4il0q7izFDL7jLTMFDf
/eH+h1ZFRkOkvzf780HJ7CimwIqUTpUqWhd7haLynw4ZY0oOkwTkDM8FpPbzfd5lEh8KeFborxcC
fDRDORzbY1ic4EiCH9t0p0dd5NnO2GXWc3iz624ipgPt+tcDYzm+IUF8HJ55rja9wf0EM4mpliND
+Yd1+YZDPXyJHf32TmQVzkio0oU4fFaBjVhgXEvxmuLc4eCiEIYBA+WMF9hLqo2u+D5OY/o8lami
2m5oHXexUzp0p78243Z+8NEaKxUSAQv36K4vTVbv62bpUWp8O4TnzRKfZT0zz5Hs2OSvjbELC/lY
j1HiW4di6LxgXUZpjJw9w/UC0gaq83zd2PkO9nVMARld+ZuOVyr2x/lLndxY2D+VMaTfefbsoGrI
NqYTGs/9Of8pws9EMQa+b1LV3axjDK+n8kTofwCpzlKF0zBkd4nnFokTZgMO7DCEfxxiaJelHsnP
CEi0RCqgVcq1lQ3zGOmne4Ajivs9YDr4FORDqVcf4tNzr/3tj45jbA44D7A15QMrWtrrI0PEfNqN
kwrzbyJvwcNc8V+11Wz19VnqkiyVuuv/ZXSXqStfxk7KQjxs4VRZdiaMAMyFf1ulTg64J4m/RDXp
GzULGeHJiy3WZDWGZ0e4rhtkUN8wVjajXPSMKZW2BmdgBYuzWaAl2VLYFLPeOfPcTlr8HPDH5JXw
le9va5oTWnv++Ua0h3jEeAGIZRndiFE/ACN3NvlWX8i2/zq6f3fL/n04CNNctSNPbboqZhqjFayw
UHUx3OP3MwGU5FgLz41TIv0eqG6Svi19CSQ9zKqyAtDrKrMLVrUHjEAnOuciZJVwudrn3bBKl/Mc
qXtZHI0bMerbdWVtc5WyVbB+arXKbYJXVrpa67uXQZa+AHCY8Isd0Tg8l8hbmoqkSFuTbAcJfNZB
KjtVQAwuYQPl2d9ecgg5vxelHH9fIJQhXz96SyBosywuWGFi7081lqxYPsYFcjVke/Yyb0jLvcD3
pY17F3SaNWAHv1fGO1W12TC5tAfXfaMUtGCZXn5YpBLKY1HRGDfQs2X3ZpP/bfYJbnJ/AyuW/X2B
QhiBFyklyhtLF0OCK54tW8SGghB0knHL1KuDCpsbC4+Clq9sQuIKV64MgMtuOsTNbWaIIXP8MO2Z
LM1Sy2OFhqO3feBviP7Cv9wGe3JR1l6CX6Gjtoj0LOD4byrX2oUnQq8rJif0i3lkmWZ7RPvSQhYR
yVjtZvwn+O7Bk+3pP0u/QLdHzC+BLT4ZfF5VkRN85PBf4a+qLNfVcxb21OTfFLoTkyiZouUqfj0t
Wnw+T3r3snAOYVjIJdlpKUXg2L/boy4Zy8imk+rD9Shn9iOQWH0qg57+ZHOib0H4a2lMvwem4jrN
/C3GJH3Pnq3voJQ8d4EeDVVob3U7wgGBf3rWFosqgAqcaepQT1i3DgHxFhjFFq6JoqJk8ZQBTwXK
HtN/A9PD6Ixce9f1ItxXo9y0IBkm9mV2zkwU+eqME/iRpVNs6EXKK/XgRrIAHJQMGwF0g/T6y6AX
HBBQmWWMY4V1nBpnHTQwZFWUmeIFvP69aknCmyD0uRsnhLop6o8UHX5S5EGIMFNbtv6hBCcyaj8e
2UyJ6y9vxiF5F0n74mh6ik5mGI97IOwD/1CdSnwaAsf09VbY8P38QAP43w2vE1Cr6gbPYA96qP17
nNb/idSdZjLuhrUfIzy6bM0WgjqCajz9hgf/2PHDrsbewCkXUtGVQ6vT482QMXdoG8Jm9d17orlZ
53P/EeKBbIW1yDYMVTLKXx+m+DUhMhVxIUg8QSNv2+Lt7jYqKNXCw20akGccycc/IIPT597NTWI/
c8G3UbL/6r0LuZ2AsStwVhygascHWbRCe6ZLPFIi1l8fpvzI/fO+joPav0/pzrI+2yiYvqUCJ923
T3OaJ//ZCv6aYi4JSiSnvAqlf4V7/Tc6Ovb+10sTR8RvARZK92tGXBmYsWC0fPW1hdMY/rCuC70f
dGqaeXe5X8PCfSSTXWDc3ISIycpv0QVcOK89uUExSu5reDFGdwduZtXYo4H9DlDSgTUP4HB2cTqA
/jz/YTCcptHU5K2qvwSCIh8/VLVeXVPvTGK0Qv20DMFoApI5UeAKntyUFc2TkwPYlnxed9NEwuJx
ZrPLQXCUbnVfXR9Qa5c6Th2DVIk6fD8qGt3FcYz7f5sMekMrz35eIrUh8xD+G1XGOYz16roC8qtI
zT7A5visZBG6m0dn91jARnXnLpCLEJZA5tvZCP9iZWZ9VKJw95UewXNPHasunwHRQpl6MzeCzB15
Ll8i52W/uzIipVUKV68+2bIPRU5ckl5cL+MfVzxq1eqbGioFLalt4soXAlZjnd8LiO4/8omD/GZz
1AXNHg2Zb3qUL0HCnodcI/kKtYf9DoY+W5WfBNUhRgaUuOsEvG6kgbfC9jrWbzXJrvvslBlw13vE
mpsjf9zjg7f4ETDSYq7QbXRuIqa88JSAnaEWuc/Qkr2dnHFFsE4WH4GzKgrQpQTmyudWi3ZJWJsg
BiuObrOjbzGlkgCxfmxxVGYWe1RaU2atE1B0dmPIXqUmA/JQ06uJz3WzlxXwBJBpQTq39n4rOkMu
NSmawT3mNVhrwjmNxxKyd8Y7FHtSKn6gnrqrsdilDBwMIM6MbDLhxQJatsrKtcj66c0lcThO5JWR
QbYofF9C2je0dOOz15IqB49PKn5BqDrV5z3gypDiNKkyCBgsx6iOzBz3IppEZi2XvVam5Q+3TJtp
ko6x8u5Hd2QikfP5kfDz0Z4O3MBkgr26++/JpfqIQjyEXdHIuW+aQXDpuPrupXvK1YQKY/b1syT+
xmTUlwuOTTVohE2EyTWqokZw9tFrfBZcOJHHaIRkaYhvIdDW/4URiWOhd2KE8EW84jXoGukfpTGc
S2oyzBkcgay1QhNSUZzckDOEDGOBv7tyufUf49ICuRnQ5wTg8JQaf5ICDgjtHkQn0gokW4ZXkyv+
WpzOOJa//WC25xWbeow+Uz+MB14LFOw9v5GKupl0l48thHzQuFfm11yaIiv70DefA87ht64y0YMM
bzjvkQ95MP5aLLt94u9C7bhlNnbPow+iYz47lNXo34xUh6plWpVBGTDuRDIA4TlQgAHoD7ZkDJ+8
Y+f+6XsP1zyvNg5bXKLHgaMgpgHurjZSzfbNTqzlqu8zPevLBQDYIk1QWSoW1ZcN9lRmFxzSNCbE
q0jMaxz4bM3szNbEB4qB0+3hNmgUEJQd7kp2b9jG1/+Q5F0mxiP21fVdQS0HPwo+uRA5MUPzT6V7
RUFCI1SpZD0dpG9Z0BOZOqj8Tzf9SEnlhPj9aGOOfN2E3t278w5Lm06hxjwgRc/RH0YTFxLfjz6T
/aO67kSKfT7eaHlvUAUZpB0VEbcRFWNeE/1wYkgL4JJNJu5rcJmJ35T+LVxZzOEZdXlTDF0chfLf
I5YMO7WKv2YeJoBf6jS48hRc7NNfjfM8PXzJ6x3izAvo7tXYrkBeHBQs4eGlF0+Dhqw+byzwFAL3
hIJXHqFn48ugLerCNO6C0447/+G5fFVxRxmvIr5lvccTy6UidYRct6dvA1ZJ62dttNCJVSaBQj1c
gcVW614BVsW9hJTS/YVt0669+nGvCeLeHMAeyIbWa3oPdvqExkL3Mtl7I8fxx7RGRjR3aMGOgTEJ
TBV3H/3IKTAjStXnVgFs9Zw8YsP+LCpV7tXgTs0HTH28nV1PZWniSKdcznFa+Dgwab4rddZ5vJ46
rw9DrV551KdwgnZk2Ucdw8TA8+NTGPy8Hmq8aEbSCaUoaaraNp6zv5RF7JruLHAWkcpT1RpOpY5Q
5om51Bnia0GbaQHXr05/lDbkLSgFK5VjWMEBaElZXx4Ibg9kFkKzG1wGekMnd06jo/rdcpxtJzgK
+RG6j21f0qdx5qxI4yHHOp3tZHQD2L79LodNFIK/xJlMdk/10izQIzvUV6g5dig6lS7M+GoReQar
haVbapEzROM8ERE3IbXUp7NEaCz9bWTva1g10jN/9xZLsCQmQCqFuDIc975DUZcpplTI/4JBIhLB
5osNzpwtNVKT7AG1j2saBPVkiqhh0CgvuBK6/L8UMbFWVhoyfD8AW0GdzoAQTpgDEQY9/7xi44+D
f6hgNyKl1Q8BL4AFwmBLWNM5HvFXhvPcTxP05xVYYbyFJO5VlYlhoZ6+hV1YLtYSfU6sjQnej2aK
znUPQipsFUV9k1Dv8E57oO+ex2Gp7xGRTT391hGGinqkO8tNJT+erQ4mS4zYiKxaShW6+9L6Rrx0
m6qhE4M/+yLjQxyvnalLT7L3HAyjqtYDsODXdTunHLJ17xrRPLbLUSynG3HB6zJhusg5DroeP5wB
uDBbTsJDVBFviAxuUb84rAejD0q032aywOgYk4/X5GHJnkOsUc6D1/YWYD1BAajbi1QUUE1B856H
E2ejsLbqmZpDw/3t2y8ttnTdnlw4XjBEdj4I6eoC5uakVWP9BMkcGba976VgjdTQ4sAJRbF1C29B
zpQxPLSPqheBqlBCzLUz/BOX+lv+cmk0HiYMSQCJk0VxfRvivIKIxB0f7TwKJ7Qg8BvHlX3fUGtI
lCvnQwroS3NktmCM7jBVwS0LiS7+37CgxyBE+fiOWj5z241AUkM9fngirrQ+c1UAF0I4GrrCD4VP
/MVGlCbiRUa9c1sB6vK4+oi6qmkRjhjQLfe2u+9loIrnNzcHFC/FPCJQJYAtdxjD90uri/wUx31L
B4xHW2XeDYQI49beLK3pbm3OlslgHO1ar4Ei02TQJdxzIUFKrx8G23rnQK05lYOGI7cs1dOJaLWE
Dc+jivHzV42cLhTaiwrWJqun2J2mmhLz1OlKk1QP3oxojf9VZuCMFo8wJS/ajoFkwgUha4+tJbGc
kSuGCDuF+tCQuwEQKqzo5fEi1EUmRAC+w4nnYHFOzwLDdxEThCKjOZLgH+P5R3BFbCguw/1w3Med
rqeTD7ieeybNumCSKU9fkwA0ccaxU1PgnYm6QlEw2RmwvnVANKDDoaGl5bg4jAMdPziC/hS/F5cW
zcgNISXbZ9+a6UPKqDNdtCAMiMAx4jgTaVvwfnFjoBB74kXYn2WBdOfBnpDkgYmRXM3lP+tXQbCP
lXFht0/EqdGEgaqvMDF0TOBr6eNM7fO0eXOz+tsdlmFxn+tmKmI3vf2dvbXJ6thu8pWLJxkfmvFC
cFYWgkG71T+VeblG8rGt3Qhj88h1jI+gLUo7Gqb/zAriTRo0WBtQ/Ttn7jx+86m2F0DeheQvSXpA
/S3lnoUp0JLS1HiQydujPJAjJESI/RK2hzMKIJm1fWNX58afgzWDjidY4vwnvGVajXRgPrhGLeRl
Zl9SQk03/+AbkWeSoss1UTJ9+uwmFlvA0edg0qBW2MygoJUvfm7/NmxlAIkH7ZpNkW80W/wtFdrG
mjrJN0BALJKLIhzXGKKlnQK9dUk6M3yQYfmiMQyacSlH+05eBhzE/S5BlDN5d6Ws524uxQYzKTVS
bl8Kih141tmxVqIXyT6rbMG8dIRdgjUcRcQ757OnW74lS+3825tbsXiRGfddC4+L461syQQFgLYs
SFeItr1+TaLYag/uzuYPDr7jcENUmi6BeAv+A6aTmOCtjEkbbIZCnsWKnJBhP/I95ODkXnAgtd4z
u38ndJJxL7GnZjrpDEQE5qroyoKBtIxEQc70B+NSRmGNN4u0CBHcV7aB0hddEIeyHSOtft2QILys
bJISDAXVN8NcNhv1k9TWx988n/9Q42P35iUSzOMXbG9sn/WrboT5JrnkFwvwFHdbQtZMJ8QkZtWq
T4X9ajvCaRQwhx942zm3xf3NpnKTOJnRELCCCN0tNgQI3/BX/3GKiW7D8IUP8IUi5E3Zs1H/dPh/
B82dnqkCE5Zd7V7wslNN1q9CDJWmyrUmZ4O5ycPZLfotoJfY2x2AqkWBk937rD9A1YgA+i13LkYA
mjVnidtAJTw03H65+Yg/wUfe6SH2OkshahrZQSAwJtqqo6LGaARRBiKTbJRqt9s6k2QH4zifJjxp
EjmTrnASUezWnWn28ou6h/HJhPzLYVLzburo5NpUvbuLaNqOeQTlHznqAG4CYjCpunDx237Imoqk
3KqKKZuzDtcjw/Qw7gQ8KNTSq2UWyLSlUuy0G6LEExSZe2iviubAdmx5LJQLA2qm+t3PKsC2z7oH
d3fC5NWYS8IOYCj45wQeGJig936DJAtgM2dcSf0sCTIOAB3MSaZzgLE8AJ0jR/NObZMVtFnWfdmR
eei+YmysUgsmsz0/30Q+SbJ/gEdMnM5hFsxtCbpS/mlnG+Ocz+VfUroRIiWTBNIuLbj3EPLB2fKS
3dkCxtvMa2f7uNx+8/o4Gj50KM8iLiTCnxKgsz0SskZD3BvAe60qwEeS4CJNoidtiDe61aVJW13S
Km4X3fPWeCC8SuUmDXQ3Z9DmnauCGRMq9qb1dnOGp+T1AlyWuSsvvsLaujEFNP1G/xJE9TveYScD
KKYFSJ3kHw6ecwO8tAX7RUjqYMhbdVmTR51WviUxMACtY8lB8IbSH6trLerkMk+vTJpw1HSotPEF
mpYOzN5829r6Nsu2dMuaK64xladIXHFU5nsgFpsj3bWUwRMb1Wzv+FwkRBqIFGKz+bzkOq3Ngjbv
bEjNdOuHg4gMqJxnQFfR0KQYd8igbUhecxVJHpJm3VVorHQEwWLapVdTiZjsM19Riex0O3lVm6ku
gFIigax4BNAHpFy7J+ap+ERMwCL7I2LRZB/bG5VEOF0FWFQ7JJBsOLzk3Krd9IviKtnbf6fiKUda
koVYZiB5kR8obwlCrPmkjSc5yg5lnlKy2CKGo6+ZPVPgEkYrTCbNhCGf1OOP+iqG9iHVdabZE4lj
s2p1xFP1+2QcDBF1ERT8NyPImsbW832B8dX////Ed2JqaEdiqlDsznE/euAmUOH9id8pjMuHeidv
lLg/dq5y48l4FM4IkmRxxNX0a2ddmKg2T9OszNV9531p6hvr/w7060binfWCsoO/dmhJFeemV2Ct
rBG1iRqOW1q8fuek/y/IqueYIAH4dibvy8UyXtlgHWJ7MA7O4o94J1DIdt2OBg6i2CMK6pHOH0bE
6QQPfLimGJojdYxZC8FfkL+U+H5WMtx9tWV6THR+B6JR2+Wrhkb3F9t48RsozZBUynYQSPLx8Es/
cS9kLXpoVeo9+G1S137Vwksiq6WsVqUxDSN/8PgFjbDrpgFqsNpYjiv6HfGDYwsYzXe2fs66HHtB
0elkH8SMgpuSSvaNLsUKWFMWA/D/SIgXTZjXdv2TqFK+d+TCwIVlbW/heXmbHr/VXUIELf4Bu5BO
5f4tZeIm/Bx1ZDHlylGQF8d1EYq3GMhEqI8ZJmDhpm7OAlv4vMjdCEAqJz3filox/AM+s0u5QYh3
4f8AP6tUKRFodLRCcBHSp4ghl1RpaRPyga/Xiwzs5TQydszfkgMIppFqLLXcfxhv23IRzvdwJAtR
/Oc6+6SEnZdUBySMeauh3VuYKreTOiLnRthTTXyPkKZ/wTnbwiF4NqXioZTAmt9cBUW/DEB0tnWM
yyM7Nywe3ralZtxT9I/K/+E3ptX2chPuWeTLdUSONXDVLGNOCT7z6tYX8s0JrNU/TTJdDtx2fOnA
U252bea93lc8aybpoWvBgYKYBWTzMYAfF+X+UPYIo3uXMzP4UQ8yRAf3ZzH2mYX8YfHI7CTUAYKj
rvDzjg/KQrwM7/6ViSdEAEJ+rZ89k5SfqvKTsxQX60ccoIG36qFmNZPzOF949eaY22sLT2IyK72c
2IOj1zu9QtVSdjJJxS2YT8m1+z+OqhO9DR6l517v9T85YjOQhi2iQ1hTcXGFRXJHMnZaJ1vCYYAV
pdD9ij8SlBX7AWc6GmstgZhiz9lf27hbAjitgHMsKHTFh2vmO9W0tjWmIDk3GktdtPFzfv6octKL
k19IZfIJx1jYwu54+PHicL9FeaSm/vi1mhau5WkeiC4295TewpVktSbAj97Afp4dx6EF/mx1KEuL
/VtaDUQxZpVjdf8TwJ2SrhkDBxam48sjxpCi5ipYyiCvn4DUfucZcTI5GAKSSiSwAWYHEnuRY+54
UHsNwj5P4z5uRcNkjv9GqaVworOiY0E5BMbeYY302Y7oBxJccZbpqWwpghzeRSsldvPU+ncSvpox
XUCEqV6EXfK2eynHvIN4s1bglNrqWS/mOwt5grVR9NIMCVRFhucxD1b4SbgofxD5uy0s2CunDjCK
Pae+F2uSG9UAJPoOpy8wfF21qkBQLWLrPxF3Ib/GmJLNatLTy6w05G6eVweo/IhfcadrcB2D1k7I
jfwlNY8T7D5rSz6bOepes7cmPwi8MRiG9jBqNYF3iB+XLZJ2nuU17skfTGtTmyxeYJwHiTjbNZTU
NgqKxlzx8qYd2oDzrzihLzSNW+bfk8EBZECh35eDtwDUtL3882tEhxdtoe/W4UzZrGkxns5H1yON
yz6l5qK4++K73hzpHQfLHXT8DzevZtSdfLvJ88qjTE4DesjPyz+AYeeAoXUaf1QnwrUIYRBoABBI
iYWOFvzFoUhy64icx6l52UOxsL8Kqz+ZWVHO/NNm9U0oVtua37lepoJm0FxfVy0Idn/4yhUWoEGW
QlV1gN+RwbfMMOwy1RfKoFx/P8sAbc9OhylpomeQJKkdXreYL+ijXbeMh/R4qNmYmuJNmHZXbbek
3Lcvd8iKCfI6BnmgRF5WynwA8on7swLca3V7Zhq4j6Lo+qo0FEHQeafMYvsGUJMHssUcqtnSnzLs
mu7XWMt+dE01FHBK5hJVgZ+rjoc/rc2kufBmQ5aahqkIBREFvrSDDDa0XGd82MXLoPlyssw7z+py
3kKFwq8cy9BE4HWbGXv1bO6eDecLKRvgRg9QYBcB0XTNrDedktzyd19wjVWw/mORupmPYWQWUCU4
YWpDNiUhtbJlrN2ifpcmERGRADa8Ps97OeFM9AfpDpMfP1Y4QmuufWoTYrRFRmLvhMZjqFHLuKv3
a8olYfA78no1oQOSpBG7vMkEgT/osNidM7dYDLkzTTOZEKXlnceXD879c7RktKMdEQQY0b2uXnf3
iHke/RWmFr4NegKYt7N2v+8BNdnMeWNcA+6qN2RQRoczonxE2V0bebOMkZkf9Ay67M8XSwhDE+6j
+GrqMSNEOF6eQGuhEkueOW/S2I/AhUzyNi8bd22wMmB0bhzzYJHbDIY8Qjzl/uinLaqDrigWSFEY
0WcrmTtKgqwnmVm5MaRF4A84lJsXbKKuV1WbFbDYxj0MyiNOhAsZL3oF73SN7qcvjpApAhpW/57S
pB6VmOArpdbjUbSEx+dhn2IHt+QszJ24g7PBjbarcb80EU0O/ZzEjX6XgxnewQgxX1mjeLV4RB/d
v+tLVlDry3dix7Euw3y78cXkuP4MaFd+kYbmsWwJ9ObRxRKjjyOEGbdEepkVnNQD6K3jER2nWlHs
bW00ig1RMHaGkY4Y5Dv8HXeVfW1CWD/EZtH/e9FnZXQ7vRdElfshtDH28VqPtQ5LoASSyqfYzbRP
FFMt0RRAPBAmBfVI53ImItVKAClR+PIiIvOOb3oBYBR3Ylye/RoY9Ykku19dEX6jDPQ1UEg51Ajg
cZk57JpiT5MDni2hL2YNdN4Wb+M/sLn5ZdSgCAbXNIQ+vQYEwVOHWXHhYwrWKBnPzF2cNZ38kkfX
MEPpK83AWDy7NIJBrC6Vw4ianPgvH2nZYOlxvnUy064CQwKcsdjLtExqpdV4AbsPXNNJ1SxnJ0Fy
yrnW8shVQLljHbstagVEWLA2zu7m/NUq5k+QCLrKFoN+QtBqv1jKWOiVfXcnG7BknR7fhU9Ei46v
6lL1RCOW5yzEiosR5eUK51eph5s6iAi7HkaM6j1v4cIQ1lNYc2gvTR8Y0Ft7hUM8fA2ZnsJjkqwm
qsChU1PGliOGBb/GZhRnoya7xwuYRcJ6rY3lyQ0dmvj1V2V3DtJNPYUHFFUMJ28dsTQ9EYyEJeE9
p6VXAFlB2HFhDobUXDL7WnESDPUJHYpj7bVzOyn9tpzmT0OrExPHEqFFd9UQnOQTOnp6/cDZnuJK
EO5s0H8FxcXLE+OIjtTbt92+z2fgDgdMkCqy/7xWSYnnF45QXBoxPB6eim8GHvNW0iZoIuP9Mllj
kv8Cl1kyq0IaYIf+RJNpfwqf7/qqXIW8GPcZ7rz3UpSKN0EyTbXoQ93Kers20Qw3ZHPJqXAtvQEM
Q+pSRO2C7ugzG+tsPwuWESb3dPcdeak3mrUCOixFrpzCZ2lJU0oNEWOdIEDJ9RF9Ohc0RQmqCDe9
66gc1gbgDGijMQegAQrp0bd7M6dgleIohAULjN36wgIsWcURD1/0rgiZsQcSEp5PUn0Fl1N/hzVo
nnyeEot6o4pc3NLBrrijGpAwHr40fR3hAxt2maPZ+to6frmyueEL1sr72TLe5S2GU6Eb0j/rLjVQ
5G4I1dLXiGpi1SxYfybFX/6/ag2ucGtnKRcMp4VSlvibHXrF8uAqWW1K4GB4CIkMnKOVBndy+PRl
/xoKX0HtEMHKjMVYB2M8+nqVfOV22D8jALUOpZYy835rhs7YIwMlYn54wYR0qT1RSjgcQ/1+iuS9
rtTZnCWfFF2+/nVXFnlMGZYvuuJV5ddFsK+bK8uLOaSMepPTlOX3z/EF6CkTZmqk2RWmDLPEgenj
PD+CpAo0IIrWm/h+fESzN4zQDQlfYglZhLi85gMFkly5Mp3daWkAiqaC2RwtPIofZ5hIcOCvDNUl
YTitqWx4v1iwFqcZkWsmy9DcApwAJ+2rfUOEZpoyMtUSTeWCTnk05pRqYHaRG77slneWrCpTkQqg
85Pwn9DXrAhVVPnPxG+cn+kNa72EVhJs9ZgQUAK9S0d+wezSt6ZiQya3tCnljdZEn+U/8fVJwIYF
q5YzXXiX4ioCe8lUKm/p2byyZ/vF5tta/h2Ka788tbl25imQNa9vcVNyrIuGSkbrrC4iDRp+cL+d
Wdkd9whMcgRzB0xHfM7mQLQ46IL44dMRVRKN7/ksX1WUBM3LX3o4dZJeJe1XJmC1B8991TxqyqxN
ehveFXlaAfUm00HkFIGdlInVMpyvDCggG9SZ/M1pGCMPC9HFqcCvMq0vlBU0H/Wd78pmV8pz6ogC
k8ck00xCfi6RksDjN20ib+PSo6+RDU0o97d8qGYcy7aIEnIM0QklDMW4zvTV1lGrr223L/bf4kQP
nRbDUotREczxIzpEKysmdJDNzAnsh8XkR9Bxu3Fb0xIB27XAr0s8L7B/gn0E3lMq9L+b9NRiJe9w
y8YH5sba9jvhHwmnv76JkJUjW+fO0Z27+sKZNBmwN89r+f4aaM49WmCN9/GUxmhDnS4H0oAHtDgW
ugSzGyURyEouIXEkcZTOd6wJuYCAz/97c7o/sweD/uXHskXCJ4YkknW2xZh7VRGk3dHng0EqhJLT
2MiqdVDtgQ6TMGwWV1cq38wb/4zDsGs/wSY1JQQOMhqWjc91qSMfppEK0B6Jgff1Ycioi0MCHBCk
TGWvassPeo4gHH7vTiJWJ0HXSDJZin0n47yoKUdvbqydRNR+lKrmWhIZADHSchX4as2cR5LG0GX2
MWVQBDEBvlsyNzmzFNPBAsh8ExTCxZ3oip1eJOIyVY39Ix8Qo8aUA4HA/HdAkZbMP57Sh+esLPwn
zAQ4zhDD9jj0IHyv2rfa51m64L9dvrMJc9yforKWfK5BFAe7VJQefztxmO6MJdH0HQQZxgeZ5yFO
oBCy5Vm36ILfuGZnlH22j4nWdqj5oBKrnZ70PMLj31wfDhjMctMbNrAAJ018SKI682s5Baem5K+y
rpW3zuzwTN1brMSEM3eBt2EYd16enMT4tYXtgo30acr5b0CGvDuaAVTt0NYyy7LVR6wYiFfuc/vR
WG4138yTpqLMyOrwEhx7BvX/sbFp+6iVRYH7/gM/ZxY2UvihDWCqNCvs9S9AN8AN+1C1xhEJJFaa
6O/4iI5h0COtPkTyZQpzPLT7Q46EK9xricZF7rsTMrJgBnTfLBDQ1jAtlxsIzs/D24xdxhlThXi5
ZxrTvEyX8MNJcCfOvboNOaUHj7xLQgk13Aydkl8L3a7d/MJap/IsqDHveoIzAfbUWXvB6ZVddl3V
d1xHiUwtEV4+nzNMPoz3EendJzHubXmKvv88ED1Kd3OEWLXb4LjUrCIIUfFfMkJNmbHeWbq0/LXs
6PVFNmyhsh+ImtPZzkVh95tciwpBOCC45Gk/wSCvZK2Aq9B1m1J9krzL8ElMugWOi28NpihxsfwI
F2BXFagh/z31HANG95pYabL2P5+MK7NJ0vahEgIpkKEyRLadH9IMmDpnHjoiy5vBCDj7l+F8AfuJ
dgExk+yWIxygXXmVYjyUU6wyz11Xkfbo0NtaAimd/v9uypC25b/1b82ftVjLY3JsDCR1abjsU7rV
c2195E6r4FuxTGRaxqQjFdu/Kn39znxFu/qkw7PXtA8Cjx9OCZ/MiqUn2QF27axGovtKh1FGqCnW
fzdqA0Gskx2Q/Jin98a+3S4RT7fWb0/4MiKxatXHQBXi9GSTrA0zi2nY2+aZ807oxUesYf4dTQQP
YU4kAHKf/UgOg2BZCLUAo3/fu4zHVcqLpPgdv/R6q2b2rV54SLCb6gnxBaAUOflUAMnFJcPplQ1f
iqJH/J52JYMOeSLZ3HSd2PE3SXSyB4KkHH5+hDTgVvEyvweSXKYVuBaH98puC9BVM0AmpW8AAbfk
In3SQmixzpP/CCbodAuSneib9A8K9R0JwXkQm2ctl3XlyUL760tIkA3cjB4SB8AXz96MYwuqx6DZ
HwmnV6JMNQEDzbtDrAAHBR2Gl2t3TU4F3rJEmzW50H5yeJ8UudSydaLhN5X3QMIo0jhNjqh/x4yG
i8i1pqIXhnV/vevVWsj14ERN83pcO9ZKN84CSUJzpSDc0buv61P0/8QjG/dtOpniz7nWmr1RVwQ0
ftBwRFq8KjsK7IoON+5llbSoC6dY6x1lV+Neu9a9C/MWyRO9Smv9A02uQNc+osX046BotHfrUaAY
/iLtgGMZP0SUIbSZxlIsa0MgGn3nzwILYCUXDRDKPTdO0b3kUj/boyba0ll6Rtc7DXgfNU+FGGGF
xx7Tpi2va1TntiziBQvBXpkRukWZSePVbvQWhvJgcXtj5uhKxHr7wp9qhl8XJnKx+y/8YJkoqW55
xyaNpcunbGJEoIuYLyN097HnRwd4Iqyae6u0s8q7vermPTnH04IOy3E2nJBJUyiXoOOhvpy3Hs+I
gOgnoGbl7ywDlhP4z7F3BMuX8yR7+2XZACS794Pn4D6cDSmLmg4RE1ZjSKcguEio0yPvMV1kOfN0
gHUv7uwzAV52u1gp6OWEHbj6VE8A5ZoAhZlP+U+ZeBHo7s4QfsLeqxLgDLIe8ulfB59wezw2mkbN
kLKLYYkHTTxAqjFYj6xh73XIoc/oAGp4s9e9CyliB6ZOuz5ClvFQbIpYE5cYJ+zgaG6H3v6nyaXn
hMqfUITQiYxcuCBBXeacg7ZIY/ORhxkwhMfKgMCfx9fmlVbVfVocWXKh+uMDwP30AsPszHk6MhQd
+eTevzen/Y7CgaQg6ProbUbAs9kUgElWSRzZAiWqGa3cI6XROu0pD09OObdH+Xi1TudOGzpU9Pi7
wag2w7ONn2J6lvjiR8mAOIGHLfa8DYZCzbI1ddaXFddCEilm5fjkU8W4MFLXmJZRibmviQa/+1Pi
SiznYDwF8qyUI5SrfZZO/i6Gtq2seX8/x7wBux32TpBS0nhs+XpjbLVwzZE9+kumEamn/1t5o26n
Qfy36zqsUwR3kZ8hwjtRpk/8VvRpKdEt09LMOuwncN4X0peQlYWWjw0ksrcuXqJorcgxWBh4kem8
Rr8YLCZ7iK1KjmvnUIXJoygdYjoDWmfUOVapGqLMXTFYfMAKZ1KeL0BT6g51D6XtCcl9sChAzQb6
XLNYMSEButbF1fgDL1KQwHBJgOLkXZsCNeln7qzwJEzhdlifHpf607fYPPiMLI59xBnti67nJO95
22F3+bUEdbCo4p5X+nQtiQVfVYdIzzA1wSyGwOHWVyXn2BZJKqb/8Hw4C9JO3djxMzZS783DmFWq
RHQVH5X47shku4chglleOJW1Aw9JukupB3nJpM4/oWrVwcZm+zPy4Pb3ycHbopYTHXP2sob0yQB/
M+gzFpKc4kmJBpJKt5E63HD+nY9zf+BnrX40yar6AJ0tPZVky5e3IxY/e/x/PJVo7k6JM45TvmcR
tkQvnNjvmm+trcdDGco33tfzbxTrq7vTHVDpb+P5hvOaGfCizgxWcOn/lmwptPEgfMUG83E6ZYGP
WCgn6YDYGXY+SoHHcBHnhKKaQimXceMi/CVQfJDfcLQQkLfJbkieT2OdmlW3Yowkpfa+SzbX1n4d
Hli82J23roRCQupe1jXrDUOLRUqFWmn0NMvL0+QbAyu4SMv5eKW7TzmkVzBtgYCyVY9+9O8GNS00
s+Kn5IpHEjUgFVomj61R9nW2N38EJ5cmCzm5aBm/5h4eiUArGecmXR70th4D7dVqNcVD9alvKKgq
KFiDa31mbj5NX45/uYafez8iCPrcDymmME2qPYFj6Gx0IRVhM5crcdBa8+1Dej5UXFbdVz0egLJ7
4+6iXhnr7rF5fjfSQ/i/K3ifNKn4nLo4reHd3DPcw92PaoSS+HU9RTH0gihEExQIGLn0voaMT9iU
u4BF5ttBlazC/adaYztdTKKUw9M2kWwoxBUpiA9ttceD1UzrtwzWeqpa5qkxEV2ivwXrBo5aji38
4uunFADkUtVjwqGdDitcTGBbRs/YYO5Tuf8/7cl2XHE1tJhPRmtQanl4WCDxCngOQv0yEVYwFra9
kX8V7vfm0yp1fSUD8VtAsgI36kxWjHmJhxshNx0ktIfkj0hRpKcnm9TAaJoEcch8x7ddysuUSm18
dPEyNES5WkZYzFUkEkCdNhES8aNM/EhXnhzX50bq9ENiq4qUmC3MKVGMoObzjHwVK4dXGgxQ/fgG
/Y0Wc1RYqUnJ+w6vdhA5nwWib6dDZTGaIRwDpuh6vFukpAZrifJgCufx7orlWgZ7xnttWCl1bu8y
IdfxDvI0ZQ5ZksHi3Fzi9Vtq1LwS6eyXlXGIV2Fxsnasv8LEaiw7EmWNOmk3aHxjaAIXBZuAKsLE
4fHMDMuH5+ayN68qSZYZ/cGZlKDp3tsT+4xGRxlONHN7DflUtvLbV7xDep7vsEL1d9REr1IuaxgE
c5Xpw+wEVXVtNhn8DS6vVh+KVHQmVQ8lLS5v0ubnCJq3aT++hMEnBBxWjJp0ZlTvNxATZJPDppyp
LCyeBNIGvBqepJ280GIk0zqzH6dWK4FW3azFlWTpHn2vXSTeZKyKLIGsVTppJEiAquQplblh93gZ
Tn2dJo5adfLOJFB2vyLI+fsckys7sz1k7yhMc5CebIz2MobOtH87jv1WvIIrvPLPQZuzm/hgqKBr
YzcyuhPwO6w+qogNxgbYbqCvT3rYjlLxxT54tJWkTl2GwPRyGSDbEiCDjxbvVEQz53DFtnlL3RHq
ku1EcaaoAEG0muIFOaVAa38rZLoZLWwvzQxTidl9Ldmmr7AzbsmuNoRqnpawsuxk1nGUmLNnaCJ0
7nrpEEWMUx0T8mvF/rQ2+o0fD1zYBJL6k4i9QKOuPlmlhakJ1J30uQSyQffcdXgkrPym0uvMeSUU
wG9B2/uIm16DguIY6Euf5q5w4pdDyw2DPXjbya4z4UHdB7d/7jakXo0QGismJlqwvm3jwYM2Tbtz
5PgJf+hrF5yfCWch1fpJLyYnRuRwsgryRnYMNOUnTinYPmXtXn1ct+WklNhtXGax466Kc+8F5WAe
CKvSVVyJQEK6lgcBmbpiDKWZjmKTRonjSYU28An5ac7ru03JqdGJmSzZk6AQ0zz8BFZURk03X5Zh
idaWoNDBqjrWjDREJepWqQ7K83KgWCxecN/ScGGPPdRF5U/x22fbAkKMMNr66vcaKuoPN1JiWRdn
hj5hd0Hks6+ZOzx0zY5JpSB/2g/PrMZ8yid8oJb3IjLbn5zQXpTbInE+ImacmOKLUtEHPtGzSfu+
N9YGLRzPsyiueo7N7NajiODCnqib6ubw8m+vNaCRZ3BIao6sfz4cTm51vvFuqS1mCE+M0N24PmgP
7elpK5N1HApEadKrpp3piAh/u05vY5G+4IevPdKz+qNTxAM4Y0gkINEdAErejfTZqcAHTIy68siX
FZ6cBz1uAgp7BDJ5aQXUU2p5uNIaowJd6LY4hNn9uSeS5x6AxhliLpDzesYVWueEbQmKM43Epl81
F2Xv8vKk4W6ujiYVWmvt3MGYK1YEiDxGLwGqwqcXLe4gR1aMSvw5jQteq7/20uYr9Bc8ef+OHfWV
3zgAfFVkxHNNS+8RLfKmDSSFIVahUOQde3cE9Wfq3emPV6SzG/nRG1HasjuO7DxxBQzlccvG1aiY
w4lrVRDuA4CKwyGPJnNxNqrKb+1jLfN65AkqUnKOjxgetenYjn07HA50RoIIZ0rNgAezH/5uabM7
jyaP8llRXs9jiiNEAi+rljYcwkZR3wE/r1YpqwF3ZNBRZId/6eFtoPEDq9zGOfgFgz8ZcUu6rPUz
N5Nk06xdkD/PV3ROYuZbt8cKVo7lR48AWdQf0e0CDM+Baehwkoow77KJdqrjRbu8GF1qskQXP+ko
CY2J5FG8YgZmWe9RgG2Wsw5rCPzpuSCp5EH8JD1Q1uUCEOBwb19hs8yFSvPDADcIQLrAhMTtOwsp
08mj9kwk9FDp4F/80Szz2jsa1HVMJjeD4O74foYf68U1xTrXe9ZJrTZsT562Dd19iGOplsPTUW2I
xAWxrbCXMFQmHPhyuwE4lcCrRCNGTDpGKpV86aifqFwXpsyffcOdsIw2e8TFgshlHPZmPBD5c6Oc
knySmCnnboUTOlql/u88/+nbnucav9H/CMnEaDZxXRkiksuZ8SmKv91FrmEq8FpAlSgyMN3t/ba/
bqlPe2icdXmMq6/z3XjVqfY05fKeXY4EhytI4vIEFDManOuFWFvVyV/VKiB8ztJA9QW8SbOyM/4P
fcC9ri4gaZBhjwa4xVW+WGcZcZ4BFYwEDVyZdOoOXPRrut01/A3mskTFGCSxnU0rfcIJ1rWQo2vQ
Lqu4oI4siZdA3Clh9wlnCEcwoTyKkYaIPAzMmpVU7paqyURkAykL96of4ZeJBei9ogVST8UV+J8x
/k7myVwavD5U8c7tmE/UTlkXkI38H2wpL/cozIYU3SlTfyzgQPOfox7QnKodU9nWAfcHINBNFiWQ
zsix8pAEBLj+PeD27RofuCnKOi4hyViFpiDGiVKIo/xSEmnwcvPgtWHia6FAu5cbRv2VBCJMbXJo
IosNNez5tifupqYh9L6KSZ+1GuduFYLG6qYLA/j/V9pXKPh5Tg4xLUn0s+YVlSVFk5I/y5B2G51k
1Nk+IuKKSJKnnlPmAdLCp4b7Oa31OI7n25my68AD8O69GTpzeOsPxI2ZVcKZfFP5ebn/1BG1Q6zQ
bvLdkPd8K0XMutol7z8JiG2bBQiYeXR8+kmNxtG1pqR0D9x6etf1Tp15ZKkUB4WrLJ8RqfjUr7tS
kwskSAUaprqTZe2CoakOuUA2AYTkhMoz0Ljh+EKOnR0aAibiZwWYS2htkLhjIJ1Y3geJL5iSzcEU
T2HWNjgrHXrs8ttd/+5fiYIZ8WPRFB0KeM0/aPt1Fx2G9HCz2Mbc3003Fc8kd3NiD1E1qGQnsUvW
LddSsHjUqktjf5EgKfy7VSSSHFA7Gz3kL6laYpUETbohh2lERb5369R3QvRbNQkQObbcNBcLmsFc
qT+P/06RQfvCX2ef/C8WQrId8Nf+Kby45PBr/koS2Ni5UV0x1TYoWhw5yEwlH9m6HUL7iD4mbdGF
CB147E5GZi6kPUMsdU/LjPwQfLqgS9P90YwHU6omBECKsS6wKPh9xV1fFr1z3kwlANWL9YZmB8ld
vBhY6ZAu0m2F/gRqwzu8DnUu2ox5T+2DsXABQaEfKknOQm1ppsWF964LsnAAVrQsaKFctUrmmD7d
vMdX+QUePlA6PYc/ne7x+NQhq3Yz8U8lSEPcmy+Z5xOby1v5FgZHclxAB7k12hb9nUg4JCtRX7vF
lld+eGD0vHWwchosD+i0dDcGT+a1+yS/JzKUMl5UET70m4d0WcDwMmC9ngoAvetNjFBv8xk5I8ut
HDS8IrKMj+bUkhDcH5MCYJe+iFG4i4S68+XxOWpO5CmPjcfe3JBAc1WBP06OevOSTD+6hQNjkYSz
50fNZGc5V1fRTN2Nv26cCkJAXu1L5kxFBbbFUvdvcAQF5zzGqW5vh20dFp1iiIQDcgSuBt+iiAK4
p4/GV8HYJaxd/248p5tq675QML5HQZMhh3x9BFMEaUJbZxNVf/E3zaR7z5x21H4oOY8utu9fJtBB
uOyepqXSLY87djRPpp/N1SRCHI9sOjgQhLOn7b7pqhsxRpOQ0a/PPNh7zMRarT0SX3/mK6wY9fE5
CKJYp8WmS9/poBiD0fGYbCC6zIxGY5SrOqheW9kaSHORkmYjTML2eqZmKyas/a9G/Ucfh+hRrDpz
g+BI7rFhG55FWMRgp7AQk/FC6+dVD49sG0PLoJuxHgIPStPpmPPDrauTGtPdgCicT0NPUrD69GQu
u5jEfaxsHcMkbRmsL/bcXpiSUmZyp8KSIq8966Q60ebOiviD+1TnLaQ64yioUVIkOSps0N5ibPZI
cL6Ia8V0feTAS+uZyPzFCOd83mMpZWidOYatRV7Lao2bEumnA1ghkPKZVWibiTi6ygUdfw7aUhiY
DjGGLXuk/nf99bYjXJ/oLCNiMQW+fSxHmRbwdkR4rjcxriRgXsjz+b9nTLzqDrkh0ollLnhHwWp7
ycfiqDAVABd148RNfkPQXo+h9qPXP5/228FF9MqhJMhk38tEOqXuut+hbPyTRhrw8T6wGV3SfBin
mbg3dMXViSloZWXP0vRrWlZYpaX/f3+yUIQQh6SqWjJ03Np+HfMjZlSRIXut+zfV7h7Wiea3+o8b
Y0qS/Syyz8tYtzHVTtG9wDoilEOiyfVJLSFhr71g1Rhe4ZBMhWpUP8kG050yUrcnwF4GO6i2B8aV
kUqRZ2CZc3PJYTqWKhOjHI3izx74/8QpfgoVe782j6FtRNCRmgB7veGbWLOXIGJGX+gWzqk7I3mM
pPMrN9O2boffBdj078JuJh9imytg7TcL65B9Cvw+XiJc/cF0NjiBoQhu4wEglo4j9Irss2PvBUFj
6Sq3+Y39+fCwnYvhxKyYvozRpOaoKa6Q5Bc9aU7wRU0Q5NQU6AzMOdSMEf8ZBDquMA2cjR3veOqO
HasLIPGMHYDDYjt5cKA5h/9SgyR7yLfLSeT/KpKIjSEJo00mrBZ0FfruvEjleEcBFy80e4tseN+V
PRTucpZdeENypXaN/ABFU+FoyWX27Qzpj8zJVYlo8ZbcuvYllaGZt/iVNARhWrpf/evHCpW70yGt
qA7wdh7J7iAFNB4z3oGf/naIwCXnoSbtqW94tFV5I8WCqOzRftzHIeWm7euOoRcU3MPxY3eqiHMd
vPWhI8VWVcy8iLDETKdGnGVO+pIf17HKThGywzqoiw7pEES5QAwKTo3Ls0OhrIvWu3waKIEGPM5d
92gPTDgMeUDFuRbbCPLslC2ghNQ0FM+NvfTywh9P6fLVS3lrLNwMd3erMCNPJQPYo+ZGWPHeNzBU
HV3qzkfqDc00GcRfBBLmVlpZ7TYPr5JtBWErAMTL8MEmcX0w4cEakNxaAJ3J469HrO5i6qP5G3qA
w9ugJVZMiG1CmukUiicqqEzI4niQq2Z2pxSYrvU/Adch8TNkAD7JliGPaynxUMYAzTG9FScNdzc4
3QuamUSFinfQ85rMprQ3CWGYaBdp3uwgJE+u3b1vbUk62H/vP36053kB4x9TCHK7/CkRIKbFSvt4
IoNo95CK80oTQOQHcalwawmx+MKupWxYvQkWs5SZQPvwMsTJxVU1vvQs8lnTfMcQzL2aDLZtMU2W
C96IQuZqNDnpNjVunE23IYynooTWKp6x4XSv4Tbh2mHDeIFYDpXNbYdNM1fw2KvoUmzaOZSzs4Sw
/c+TYwRFIMYcW29Dx36B+usBjxcdSEMlujfbg53gs7+1NPZqoirUupQlUpKy8KP9KyZHIHn463rH
1MdRIRHn/ArX2Csiyy+rk4s0QBXXIiMiqKqvFpY6YfXfEeZqiWx2C6Smr8rncX6UUCLIWCWVNYwj
8S7BMgRsOW36yJlX6tJNkrC3bh/O2U4+6HRbFDn3gKZWsTC2F3YJ7Vq5res0BpK73cNJhzhfYn4R
pita44nHFcagYutV/0/NB4RjBxGjOuEYHYTrbyQVoVcMc4vvXwRHRhjXWIfS6JTQEacPhNF6vC21
LlvorBHYqykbATnHAVAOaqE5kzVgiXUzUwWrsza9vmMbSKrq/etuIl4JXWR22n4iD23e/SDEB4ic
Lj6Vb0NvlZQMctCix4WhXQvXcZ5XQfsWF8o11rrsmrfiZqmE0ik/oYJ68NJsQc9+OoNiuatgIUq3
Y4X9JLmxboQuermFwq2Qfa9sAQ+YkL5XVW0mLYabk64CzaSwvDCmdqUjuoyD8IPDvzCL4RFEhkyB
UBJxOi2gE40agKZAp6TaXXENNmQKMPVNY53xDvMBgYPssugxAscJyVixdvp+pF7cZyhaNOPb2FOZ
DwjK4zFGWAaRb3P0Dbtyyiu+FfUM0g1ozCw0rAXeghUKNPpSgLlc36coryTqtasQacWw6CWZhjad
0nNhAcdpL9Xm80vf81Q12AAq8GmW2Z2sjlpVQSxwIK6wr3nxaR1/2cAp2Yk8AOwlJ+wdJUB4HjnU
SrBHID2fwbIytvpuwheU/fZhDTamilfcXOwMzAlIg9dOa/1UKOtq4WJVIESEMcUw4w9jQjV5Bl77
1xyK1G58uwQNKmLruzGaUoJvab92ZHzEn3U//S1/TU5iyYqxs3wXSsS67KWEI2bl3vOhQS3mkeBV
1XV+Ic9SMM7xQYHXgqlMjEzhYRvBE002UwlfnPx6gx9Q+cTQbuUOnNZwkEUaFKcu8a+ovpLLedce
P018UvNLkyN0jYskgB/7Vfh16gtuUDa62AX/jxvkEYdc+cZei7zoUDfrkzlq46qtwGfUkkUCBlkd
m60ubtfw/qwA0s77AUYL0GCv/kU8PuHLUdbZonkuXu1voKnKxIM5nuXO3jJpxbiF+WdtxLX3q4ic
/j1zKGIB3rlkNO3EUYKnzJAZJHYGylVtIsuSQuDfn38E+gGd2SZ/w5y3/E19nvOJKxI4O7i8eyIT
/jxxJXFBIunYulHMmBtxRPz12jvxjwefEYkQDHpCCf+rVvC0VKi51LMC0W7a0LtLu55ywfRuZvtB
lV3Lcw/WXCvTWAx9lK9b4/St9W4fJH8+ukjVyjdTJLCkrPNLT4u/oUIyv8NFS8L9LxMC04Djpiiz
HJiLzL4ZGTXfKS7QDH/y+Cc2MnkQ+faawvc3fOgVffdyWtUd/LbBpRrx4woz4KxO4MO3qiCD03MN
WnfKdijN5p/t2uvgtH/gO5hc691AoGt71gJcoQ7RYXQZhcc8P9m8z4TO+JJ2nU1MvCXGn2/gbhwj
z7jVW9K+VVFsAarjGhNkhI9CFZbK1NIR9YgbbDayecx345M8aOYsd+Nu9656ku7BN0YfKAxnLPaL
MM9R9em7oiXL59M41P6LzfU5KBynsE6g0T/nbaX37JD0fzywJhdzqsuvIYDmn4fkF6GkhL/Wa/eV
h+YBssNV3e6cIpPgUzj1HidLrBPxwrVL5XfXABIoAGKN4c9b/B7I8RkvJuDa1F1IcJHitR/8mxcu
JjQyZcTeyMWqh0AvdL4dUb0qi/k2vMVoAzQx6XiEEHz8OnZ1kIvfMJgh3VF93sErm8AJ2kCzsyZb
oz6gDm2tPeEeWS8otCn2eNKY8UCiGenBxs+l3EuJg41yauJ1SJZGITZW69NwQwCnCuyUqHnnV6QT
XKoEc5au0aZYdaL8YXAuYUxdQGDNX4GmM6IFrrw65IBtByunIZ6T+fg0GqMTYPSdeB80zMKAOnsd
Cchb1KaYKnm9hc5DNivBnX+AyIQGnzpKBDJIgF/v9iSwRM6CXm1d5zvm4VDzkKWQD/WrhmHzXC79
tJKwXuENvQYmMwjnDFNmQL2Iy+b0EfaWEDvHoAIMuL349fATmB/Yz2IKOxQnPletuF4RrQmasPah
c4UvtX1aj3tIjUvwfeZMnptgp8XKbEsMMT2gHKRRRi5lzacz91/4WkTRS5kzjSdPSPy/jK1vbRwT
B+uO52yf2w8WrR3cw+APEWU4L+CoodoAf38ezyQVX7BcMAXDN0NZgu089VWMirvEOnbhEjXVdPPn
AOaeQFA4Ud52zXu88LCLXLg9Eggei26ibvXRHy5ztW6jH7sDZQ/jcm9ukmwP/tyEzLNyQye4Iqo+
PeIZUBGNHDCj9oJjLFg6cwdfAxWnoEICPIjeURYQ/5H/clW/pYO9na02v8NMUd+2S+23XZ7pzTEM
6TI/zr6CfL1RFndoQrF+AQe1qAuYVrw8TiYHRrrVxPjzzCgvMHbQFHvmSPh/5G9CKrz5j5SqSk6f
t3n+dGsMliAx/FP2k+tUANGSLX5tGLGRV6OU9j8nIrq9oMabu4EbloRahMNva6iaUA7tYCzD15jY
u9qB06XSsu5HSdM+5lpoO6jgIvVaYKQcpA/oso5Z4U2CqSH6Wsq0aJgMYt+cIYt4rkYVbtKiMzo2
DKkxH3b2jEViWWViUIfGmO1bWGpafDNQ+PAwaGpevnUsac4ImJmi1IONvXuRr5yLncIE3BGMMaRR
p5aT19aieT6EuLA8zeD73VVwnVN8bh9Xpc2IgtiYyWHADYtGQU3Yo2SbqSxsgLObSAHXWGSUmakF
XOK3s5T7JgSJ9fPnS0jAA4fHfgMiymMS3e66Dy0bcyDNwHFxmleafiwwht8RTtzF4cF+ceL5TbvD
KYl4Xn55g8VC2j/rqsJW5pCKUbMH7rzdG7RrmWOq9YGTof+FvDXo/fpCXGM9ohqKXF/gCPKGh6uP
eyDePIcVN6DwwMqkSieVMwEoknKUrpPZmxslj1dsT654CAv9zC8Zai5mGhtH0SIwdGljMQkEcfan
slp0lo6kNQt9msT6D6HRXudRnIdrodQtQ28x4vDxnqRmtQoBKOhpC+jk87SwmTb2UjPJNQd/CtpC
K29fX4Aqr81Ubx98+EyLixE6kNcB6ekSaHmefbRTCiWOjhFL1fODghKoUt2M7tpQSKbDank4MuDg
MJa+NwajhygQwELf1l0+/Kry3v9DMoD4TaAdCBMVfh4EK8jVFNLfVOzCLgjZlsX2wgZuDlshAtkd
/axnSn0VKdf3i7YhIFjewiz7B+u+KLC3uW3qu0o7e4tzUT39nvC9yvnt9+eBE+/6fiUeSsOBA6jo
klpEqjQV+3ci/kGJ4hqVoLN52IpzaNzUMDOM3/MCf2bnGqrPyoykUPQy3vWX0aYL7S1kl4PPHqud
hNsRp2b/XhpXHxyTPkTTqjeakWUfqNQLGS+ZxzSGEo9pYt6GBS1HNKq0QujWDOHsSM1DhYDS/khk
NJ14PY3e+imEnTZbD1d8aFlVxzzECvaMDLIWHUpzMixUIcl1jV2xaUk3QcXt2+dUCZ/mJBIMkx3M
HvFet37yJAjW8otKj+LGqt2KppUJjibunsprJOzy7SQofAL6O0yw2THbMREt4rk3UPlL2Z3cfi4n
5HRZo/H/k+AvnrRS5p1Kn3IjF47Bof2dhZwr2sAD1Wugmc3vGLOMO+4bVOtjoFNyEwQ6vG6OQCdD
yIY9Sh0UoHsf8K7ghY1uLb47/p0aBnioIzUT4aFGSL+8XGJ2Vnz4OAhSEJ3m/nnfHJqTajfSwE7R
FgPdabZZoumfL5c88Txsc0D0PWnCSi9oTc0D0MUvENLMdfAfT4t+bs5EbaEk0VNTI/6WIcWOa80l
4UgBO5XUOgY2LQcsXHBK1/Im9KeOMfbJRAfb8rjqeeKJe1+sUrnjzqzZsj/q6n1KLIewbFCzScMo
ZOhygVYqZNrZnyQJHgqazFnGsNS6+ggit5kW+IExPpahnMCjKRiWXsvCglqtvRFlwLZmGt09GMys
m2GFsXejDYCVi71FXp+iTh/oePVLzBmoclHvia9VNNxfFxzgjmCo+mwQvjeaBYTvnLo08Q4VvWKm
bE/8gs9OnEfek2Cyp17fA+/ZfsMJehXI15GYGwa6yzLkedVtXgko118wuhnCjwV1aoIia3ATi4rt
K3QRfdQy2ZqbT/5BLZ/vtQ6dCtCKT6Aq1ifXt7pF7nIeCQNd0vW0SpCwQjlLsN/9r3/n+iWv9m+u
WaRms21MdctKY/jOrhiSFU2fsJr/jSjFDAo419EjhcH+FeQN/JY/Sf25oonc419U+SExv6hf5yNn
2eEiYv8XsyUMWwXGfPAgMeFkyTzcfGkeHMbQct0kPfDsLOvNrgRlWfTlbm60oVkpaq0vgbecbMxI
41M+UcYWxwDLBfV2l3E4KopFCjh4Y9+xp4DvcAGo3ckeKZWKspLo+cMsfIBvALcYbgN4lJg+CkxK
eY3ZY3uTiwHJGuZOAbfMabvKq9n/t6GcwSrWgF2Bf2l+7olAOYa4X3tSZ4iefdWnouAfRcYV4xIu
y3UV7wQp6MB2Uq6cQ69dXEev0R2FYRzUjC4YiPCEQHMN2XV0f4vxbizOAHl2I7M7m+hCtRAwt0eb
nnRKpxVAM38IU2KBs6zRhV09Phj6J317x8gdvRacQRKTLfW4ed3kPCOlbVSzcFERsheh8CoKPYn5
OUhtbRW9cjVXU140/8vhJY3ZkIwvZLKFhIi+prZ3RVZfDb+L8CxOWNLWlhkOmpZ5iP0cVPB9wOtV
BUUmTSv2r0Qcb2KEtg3rnUrgXoQA4BfosSynBSQKhcLJDwKOa/9DwDTWMWmHHcS32haaoxkhqQaU
RNLEgH/Z6niuayzp+7BGCz2A19X0fpzjnPsII7N997cgr/MMSOQZ1u1rMmtWXMBOScsKFDT+v8rj
mbsPvog1GoJ8TsOeIjVxGw+x33gZV8T5V6YH0o1ocV/hopjpvfzVDaALAt9XnrgzPQ+BSBCUdJZL
hiMo9S9eMshh4LUBHjtbS3sLR4ng4vFn+HfQcOryDOxfJRs6c0gYW9OFWPTSncYf6l7cHRYEAJHh
si2cwvS31dvCqcjBV3YwLO6bovYKxY0iFKOyVHZnkhry6RsDo8xDTlXKZELnBCmRFHBpymnLCDLW
hnLKprWg67fFx4Ph1k0q09rC0ZntrRsCsf/0GD7icahcyTm/IYc+EBhmdh6kEKCFXHuQCawVtvVP
+2/h4OEMw/3ZTOhmxWdyJHg32w/OYQ/63i87R9y4tcRzHZzIvJE2SzGT/9irq6GKM3GXQZWVB5oX
H8AVHAg+SJ+Nj6uPkgqWBFbMhvN7x3w9B+9WZzPSAyIxx4hd99dMQw1cppEPwzdH1rzHNp3mZo3V
OTW+ZaliFiUomuSCqGgqNZ6Z9A5M8ItPGjP2CDe8oI2BMbWTtIYRCxWfG2tggRNGZ2GFKcLRCieA
o/xOBOiYUffQYYej9j97cBnK4yMV1MBFh2AHnOeGCIuypIo3Odx71U9GzFj2NwLJ6O+VFfEK2gVh
SCpYUACjnSyRF6xsFHrQs08brQYv2hNZkGOcDnH0DqwEOt+s8nDDKysMnT5fhciFEwmVzzZo7sqk
6vEMu25I5l8t7mKgp+GZDpaMonsqaMqfDYpmNo2cM+rnmMgPV9nkjdhGXgfNVzzq0OSt72OZjiq7
hG0hFmOJ97WULBBAeNZRnPr8BINarrledfnTRjSjs9AS7TsSzd/AQ6+PsviMmlhfdFxxUGpxe24n
GrBSsMaxcQDcJBkH994MIsvqvucY/k7GXjTyQzLgotKPZE9hBadVOd7teKbpVfNZNrp5GGsaeEcr
4hGu7JIJzsiiU5ivWTFe4BqKB66mlRBf/bV/uyymA6Swx6K7GDMh8++TA8ozY/Y69OhzUnAZy+ls
W8o1ve16p27dz8je3HABFFYQaUfyh8WNlwEJY53pOX8QSq1zNcpyRDdCm2AgGAd/mqPgc2nGx/R0
QvFlwGr3TAryUKQMtsN4+NzLvQXtkPLvYcr3dhFmgE7+GBodlackABPGRK1DD3N1Kc4CmP2+nLux
PaWK3972vuAo+sw6bltIWjlMuFPmpJLUM758v1kOFTqB7JP3jb0mmKuW7n0KNPXVB29cv+kmbNYp
/JEqB5pnd4R+nVd1E/qSCnSLluYPy3Z0JbLbpAeN/jUbBzp8V3N+kKv3ltYOAHsJS7TWcl7e6Ypa
4pOiHmo/GeXtj8yY5QSABBQJD0IPq6hyMiQvvdDV+5jURsVvB6/dEblBQHFtHCVszODLudfEH3FR
ckJlTzszeRgvV8xOf1ylhxFi4XLKgUHWAQdskPQA9Td0csKaNAxp5Ti2xNKAA4DWyKfIV4yJpz2X
bI8tS/puksPhGUchahKxXDhxws0hNBqowSrhOxI2uAe6cVztEt97fqAmG3OBs0yHWDgp+Ot4EDRJ
cCjR4W06PmhFerLdXlocf3P6SJF7x4WiLUDjMQl6wDo6mcsYRmsatuS0jTRAg7aFBXQcxqJh/0tv
ygDwL2dKhWYPje0+j7fyObVkewScT1FRQks3VL+n0PRXLpIOtVumqBX4pM2GZTc42nR+rPGtkjTd
B3VySbMCJch3E8DO78RzF29FP6t9zu7oRzCBG7RVt9tEKuG/xUKPmTfKtGSrIh/FSgexSau+mFUp
zN7LPGQD8Jv8s9xsl+X65luSxJiEkq1iG9rUJB4YIGseN7u4OzZbfuLO/yFF4XiU3npk9FI/BG+D
mVzwnFqRLVcfvZoWXRckMXMCy+68U2AvIpTZHECz2itAqoTDgNI1RK2uwSw5PC4bVHVcWMptczmu
ZQGlNJ8cK+QNWpw2UfQgC55jSjY4aBqcjjSdbZOHZ4toeeoeiW9txMFB7Eht5ylD3364ofqgv1yQ
k/O2nxG1c7eSG9R43xGlfB2ZJVKx+rAh13mGmvjfHtjHFuxCruvU+bQpX5iyWZ2HnndL2amPvfjo
A7JExFSjxpDAnVKHFLD3G3gi6453LIC67k34CQ+ZVhnx6/YexvLATNtUHxYzk/qNqNuHBPifD25I
zdfAQx/P9uqfXsGIHnU3J6ctgWp1tWL9ihFQgGlH4WbhPvtLc1TVTfuJFLJ/FU0/WfFOavvk6bWU
XYcuuoprc1J1kjxm/g8LwdRT/xRbhIIG0h/pYtAWoxevaOIqo+OPVqz5mBXLbKOCgbjlvvhcUts1
lMQt/dp8YUmn6tbspQvc1rmiO54EsMjEb+jaKczBItLnrAQAzb7jUrMttOykQ8oIhg0El7Gc9AzO
tQEOr7X6SOQM27VZeqpvkzPAZxZx4BAJTMpNjknXc+OR+6iTTH8Z89OfaI9UO/7enhsc3ag58K6+
gZjmHtozwEaHzWASI64eyuADRMX19L1nyQUmr6ouqr2raUwjnGro303vbjPAjP5zmJ2/iq48mdXU
Kb5SyZ/C0FBMHpQVYMNIYgHL8oBri7c3DYh69uiOBhKEoS9QkppCF3m1syRPzX3BFaVAlo26SvQi
OoWtIieUwYQDnK1+v2nNDS4t15NoDvQpE3eYfSqDQQLq4g1fMNpsUAfwaTZQ8RCwT4TLxVO8Do7H
O6J5LXc+nDnqWtjJVw4HdUXYr7TaIcMDAWeaWQ7UWUPAqatb2XoUPIAx/xEsG7yIH4pMHgGR5rLG
cP53J3C/t/uGb3ota3gF7LhNzMI6JHDIaxij1LrW9TDyUCYB93uwxeZCVOcMXgaQorWhg09ppbB5
Vbyp9tRp1+9xv3XUqqvmjQa2cGPyIfhWoMhNUtjIKvxCx/81rlwh1Z8u1OTCsrOp7o9YtknamIpO
rAXWPd9/BIhPTEUKSJ27e7IpKyfWC+V6PehScDy5nOYmTlmp6Ps8Z6fA5P6/tPgieXBuSSXv3i47
yzgdsaIDUoU1i4C0DV7FtckOjP2B4oQkbvNOXqXB27VZf3xOmXEhnG899fDSi1J7TsaTY2ubHg7i
nXI/rT4K6UEQ5Ss91Q4xa8oWncgSoRtCJUcfQyUqJwQClDey4080ciyq0rIBzQ4k/Pws3+XKgSB+
76i+GGvkgP1qfshhsTyw+0iAHKlRS6JYKqmQhOJ2T15CAfkovowDwO2G2KpUCyvmEmIpRJHeg6+/
IHS5cZ3iD5itsmVXlCeI9wC4gUfieafn2Oz1//XW5/xoVf1ApHTdc9eFwYqX4OX3L2V7vTu82mGp
2PnViC5geaWrY84HIPh1Ppbz7mFWC8SDli5625Qd4WdgOHHSCFY+Sez3AwmWbI6A5mk3Xya2ZSwt
wDr6WIq10EYE+psooOoXkP94CtRwL5SdkgPC/rrJv6IOi535peAvzGJlB4C4zDripdgDyQFEDNdS
wMoEAGWEksTuLel36zrtAdAFajRX+6V+WudK7/j8qDiZTeCSof5Ji+II0ob6KxtWawwbalvpfzfC
VgKrf3UUeYhU3uhh2XHUQC3AFHjPgo3yGyktkwVRhyfWDwgO+yFnPcNek9llh9a98yq5rEBRiKXU
hhc1Jq8WM60ESnI40N4p9K++mqiWlDCMMcJZ/U0l8zuPMYkd21ERTbds11AkT6J89zbqyLIiGXvF
1pTIhlHAQnwkTZJk6sXKym+zSQBfHLQ4i2XIcPn5s/+2kb0WpOwB2ahBUpjlwGkU5mhhmSIlUst3
Fa/VMJu1+4wEZqTYj7COFsBtc4Eud66JzI+B7xgZdb/xULMrqH1gmCBPHBpWz2sKQ2PHulpqaHrj
l1E7s6sh6AykKB6gmAmkLUHKpAWmXldXf5NAjAZFdn9Q9vVfE5qr7784vR763tD2ldP4m34nLOtl
vABsUAOqCs3Q7CX/lOKJJ4DSxbzwWy8m3JENdx+7MnmjK4SUhzAD3XD5krDynsQdJVLvK7cpvHon
+8W4Ms3B1AcUwlcOZ+80MZ4WgP2Jkz7rXkYIelRSRc01BzQkVSeYS5HU1mJKQNVCD9Enoe2P9CAD
fj1wPsenA05L/s4QCCTgd492ikbdkN9Gj8+ghF+9IQvivIQIAXIRWxx6xHkf36zBQKX+HCp+EpyB
65rFNKx4pRXk1WJMHagYTot8yVl5a6eiveYTURZsurrJU1aHURvmoOLMSHafnmJbg57vwBNrcy6X
Xww7YEb0ZLGaQW/2cL89J+/WdPQxMwjhP2DqcHjzRPpi4iK3rllvxhm6pHStFBLsB18ARvoDV0QT
o5dCPg2WlhsiRmKtAPDyCw9rntTivS7UKnHqJex5yBwhAelua8S28S3eTmjKYLZ76jaHRAz2AlqF
RUkjz4xQn0lnYrSD6SF9IVtVAyOQwTrH5/4NuE2tnnOAtAxpYg46ACoiWIVPtf0T9OPX2W71AK37
A8dnObtXH30aVgoA44KJRVv4QPtdLqlKmbdeHqvK8rzUZEjtYW5c8Yi7rHOeax/TqcCY1UIJclvs
c2kS89K5i3As9t8jooJOhze9rAiwPq0yEz7udnMqyiIDS8nXtL0ccolysFMhRgvVIJT7TJegDRGu
P7rd5kNW4hagEEBiFpXBHVuwaZ1WbPZnuIJrohMDSkLgHfNYdwt7hpjrHtMF2bYtx8al+CH0qBGj
1JRRlmnXZlivV4OpKcIaWBn8J8u8KH6EzleROPxHj1DUaYq9yzmbEgAbwgFCz6I20QgoFiUwI7TZ
PG3NBZkSEe/k/Z79Hx/bjBfeSk2HGfmohSqqO+tRoQhStPOPaDg/UzE7iBCEmiR337n6ksOwwx7D
5JjujdfNO7jPhk4Q6DRyMVZIHWvzXCI+Iynj1/Y6lksqzgCkpMqvrQVozTXl5jlKiM/zYlAn+R2y
W25p9VG5PBCg1oUbSTsrJHob24EF6vmRZw6uHe4Vm/xgxEtttvPrJ2rmUBqOspt77WkBY7y1PgoL
LZspGLxWkDYSv2UJcImmDuH3UDUSB+CskDGFzHqgVZGclEy6v+R5HrbZD4hHyWntnnbNHiB8VLmR
rAABOvwWG4n5jtQwgnsKVxxatdcFrotVyhP0C3b29ifo0d1OQUTXZYWRjeMkwDRyB7RCiALBy0N8
cqYZtoiJqV8sAphh+32DQAP1VZQ3izQKXWvH5DjEXhhUCFxryUDKeVomhcJlTcxjhsv5AeIgsAhT
Q1KpkG1ErhSNdQ6oY+Ki9j0TvVuxUyW0EtzGBNb0cqSU+V35oEvOR2dLscjfKtj6tYlRf0N0/amU
yAHcWackeMmpvP3e+Uxy9q2DscuHbJoumT6rWbRQY3Xb+LNeqtkkftED0AXzbQNlgoptTCHLvdS1
6pp8t04mkfdmy5YUpVR36SZddLpWT/8lveHOUX372p0/3uckYQx5NtE9DY8dHdDb/RON38deTBLp
YeJUfdEx/uSKm4weA3HB8mRguJjly/fLCr0/+1r+shkr88BcnLZ4BhQkXEg47JAzIsP7JCROkQqS
Mpy50L0ABV+2UReO8QsMgFVaOj4ue4OjaQfhCli5+ybIxL5m3lo9GMnpaQn8wLel4l/Unwowz/fQ
pgB37wUBl578+IOApZxbOVG05RaqnZj0mFoC7Zrtm6oOjiFR4/5ND34k5LU3KOJON+iY1qqOcAaW
ktFK7D08DP26Mz62VS5HBhMlL4BApPL3KnIl+PtTsm3TXATl2JEmhpyrEdsX6+B8aMBovtIVH0NP
qbS3GGzKpO4StHeOghUOTAHWkVzE0YlWfDRYCuT0uoy/TbQLXXfZFUpITiHDVY15wT04QUf+U/Ev
hH73Zchvb+3auyXfYWy/N15mMJi4Lk/RFNW+MjmVRHzPZdsfeJkyf8emY7gduuuBK0MxGutGSm/j
UaEvHaxKdW0hpSD7pF/4Ce71Jbry4FOAXtiMwcZOBaQTJy6OfcKkDMuGrnF+i5g7Kn3kz6m6q7TU
HyavTDqe2rMxoYnm30zXnMPosRRucjJlQlxZ3USrYufbvG64qciWXnYJJDp7Qh0VFaNfn6TEAWo0
+VC5UNuV7Xg98T70Xhm+YjLhkTZksY18uLyHdYtxK8tmAz/GxJXX+jh76ndZywiYh/inbun0f1Up
NOGCnJ9OpiTpqph7QJ/hkCP5FmT1e3koclWU2510N+JYnIXwcs82kcJxXbR4Mt/aMGXZ84WNuc1y
zOcNQNRikPFLqNx3yEfNL0rtHJsAemTL+Jjrvq20rWKK2VZkM1FlBMTHpvKzO1NO6PioPtBQ9/nE
rc0sWFPiI48hl9E0BX3Oc4fDjunSvfarZ8okwSYUsopsbsCeq9UbxqJ2Wkx0u5KBB0w4t9DM1Ecq
fsW3TuyXkFcWCru3Se1Bb9QbextgdzHn6kRmzg7s9WwCwOvms1FyWRuZjI8xDSaYI5SuAC5SfxBd
lfFIuxLQ9SY1MyvB2FsC4krS5OlKDvmpLSVmD61KMpGlHGKXuKoGcHDzNkU0cZngMPfsycA4P5wh
e4G1eKolt7mEF3G8v5WpkCW5nEirXvFYEjg0jPm2hTttqf9iFb3wwNzkEMwpAwJkrCR9m0wOYjgn
YJXfBdnUjiwa9jfgJgfqaURyRrxwySQrao0Kpu4L9ShdG4y1gB4Dt9DYNGOCSYotlUu0zJo5P2a5
5CijV6MLRcokkt2Htf4g2Rom4Ecs1T0IlI0bmH3lHTnfbNMORYP+b+m4NCISNpByklHU8Kgadq4B
1ZwMXMki6drI1lpU9A7L5pCCgSQOgYsnSs3kUJC4HLvj3afdw2V5p8dDpEEBr2Cgwof7LBT/7TxW
vzvSidt+lDGwu3HpbLtR90nRdhzL5wqLEhHe8XnZivrFW3DwcDdVMgU49TNExCX884NbowXLSb3O
YfWN3TGAguXUU0e4ncRoBrSP2RZGdfTZ+LUNBLJ6W6c4GGdqJEiE90cKXs+DWKIMBURnAD3wsGOs
eYV17SBqwpBnMdVVVMci/9eLpFkMcjVGBZvnzUeOhRO2l8clipEnRz+BnASzFDHoew2K8hvEETrX
dJFvliKyfKR4uPa7f+aSjWzddPuPVhglSNXyPtfQSsCOk/5JPBGlAKU+LDzdoFCg4eTaEdItCKHj
uWScAQXrHK0i7KDgn/3Qm6m6CMJM4wdU8zhGu9Bi2CKfiLpQgBbO4bSbgbilDSU8WSBosoVSgGyK
gyAQ/RlsBtSCtIIN3I2po++C6GVqHnJEv0if4GbH/zWlAtcyzRZgK1OwFxJZC1O39FCszR7OZo71
UjIs1txttzawxBQogYki5+7wtQXx3tZ8P0qIvNOg/j2cCVsOoJPyfEjUZHMOzYFXUZ1gmUvHRgo9
xtCgCfWmvowG3Dp1mNuiVeaCtXEK5hMi/VN56uuihL58otRMRCJhICdj/2eUTscO9nHURwXi5Wgp
clTH6lSu8u2LavTmF/PaEG1xHOyabsfsdVlAczqzqHBFDHKlff7feBYxTMTYeDRYTI2Fmfj2whOV
FzjA/w/xael0sOC+zxKKWpdOdzTYOi/UZg5UmT2zNz1n5cuAgkCJU5LPW0ksx+/9OL6JSITtdgL/
keNkRYejcClNPoXO5BTthfvrN5QvQlADaqq8ewyW/KFnNCeHIoFyRmQIX2VYf2HJIGZldMt4O0T1
k2Kme5m6KqNTRmoLKfMn/e/68Nj6IYEyItLXGAZM+F089RElzKNWSvVezlzIMITRHgt5pQxkrM+c
tQiPtPcBSOPPkcovK7nhjnM0CCv8qX3L2BOnhJSbQaxYcJTfS2iL6eqQihnQn/atjXsUvV/MC24o
vxq4qyoSU3guaZXdoOpi2qYthemXxxSkpgPIBTTj0WR4ru2h6J8iT4pQQuvlyoLtBIDX79WC7QX6
3AI6ceEezArRqmItzZIewW5octvd/omNVLyVpDr4UnMxNgl67QEXdsOTVNKcCfMWn2BknZkzbEtg
QTxPcrgrK7jCn+5e0osMZIINCl+KKg/vZ4solb5eT/ss6KOojrfSXQ/z74g5Tfn18jCyxQ4xSr6z
mGPj2C6sI71FKLCZhHI/kDRwmIc2oN+4c8PvjlAo6IdyjE2d8+VP6cpC8CJAojyJIxQsFRzBZS/0
C9n04baI628KMeoLQxjd+VMjSGuwUphKD1leXUOq5cuDrQ9ROA2zJkoQR1YewtHvKJSMh6aWV+FB
LMg0W1BBKW2HhahIgX+7jLtScDEhqVHWCTRiQL1DQBmqRYC96uJt7bxHVJn8cEj9BwbeIbUUO3yl
iRfNkYhJxTwdlWuc8OaZBvylPZbXs/rRcrSAQu8zNRQuJ+88Zt8XRo+jbuz4MOid+hlYMcsmBX6o
ZV0j1zdga4q3QbUREs+4i4xn9WAdX5TbhMTyLvhZdu/ouVBfDoACYShxJAasOId2EiyxxdJirKmL
D1+ClRF7bH/OijD2T6nmyZ9S5f7lEZGEsaFbrXOqbnCL5lL01xF8kRZE4fzyMt/4z4M11FaMA1lr
pLqhWCG7jl0aN/r2wbhtY+7qLzOHks9jNo3ED3421oBQadoWyCoGO+rKePa9YlV3FTeZBslVF7CZ
UNyZJSYANK0CnJhAaMD1Ux+pyVSkhowawuxJKyT9bUIMJkg7tncBoUnHURUHwp4d/HKtd/ICl8yd
qCYX0S/6P7SNVUYppQ773dfcRpOxGAE2N2A/fgnWkORMIRlIlEQlXRvNa484OotosmxhOrarQO5g
LTMn9dzJ+0OLLtjsDgTCIppHeDWU+wMOMEXBfKCZG9WHBspb3RLdZX1C3vktfHOzMMhBNyC+4Ix0
FymcFQdn1gdr2FBhaxSV0MB7sQWTRJkB74CCo1I6TXHl4vYM3MD7Qj8Dnqx1sdEoVXp8cNRmhZoF
3GCKutkg0BosV6SMQbDdVCmUmE62fwnXl0/GItKmFp/XSW20ILShscjD9ocvXyO0ORyJDOrkuVs/
tjKHNh9Rp/LJQnBO+Aj6xuXYhaHR7uAxZxEbh8g4CKRFIzcjy02SyASwOfE+dun/Uqv/keGiLSzW
VpqAmr79UHGXPhVwwb1IHXY8ye+3nopQEjww5FvLctwKVFmxlY8VvkHbbPT/iZP6TRgD8Vs4NcUU
ibJNy1tCRG3TnyH+BZXErf+XbIWGXhtNwJdjBZpe3cow78yyFtFNctORXFtRM3MGOIqHaHOfnoj4
UkV2+ej7ZuJQLhZmky5gjntc/UXvrpUMbARBHk1CfmprVOtXfA4kAzSMYCv7a5Az3StQqnCflGuq
TYbZptJKjplcxTDoUX46Me9mwDL4ZEUqtOWKmkv9IxP/YrjJAIZ7g03dK97f2D9d56pxKruAWGtQ
gOswm7lbWNrt0O2E+CEugmO5yk+D9ae4Fkh1AHzLI+S1Aqs05/UcZw7q3PosKiOtRwvySqsoBBEQ
zUzS1pnZQT5ndlCMaiemhKwZh0+ls9c8vuWeWZ6SZUpv5tHW5p3S5JB3bqNAULUbOldWeuCh+yH+
sL56OwfQKQ9vnkiNp/J+XOU3T/ryAK6/A0jLh/UgNczi6TKZB5QHclyi4/wcVqkKSUX8mX/OCSn4
xcwC08fKG/iJcUTGrFi+k3rg/613kD3bmso1QLp62pD/e2H0KZcQFaR2E+NXkLbCyaesXcEUZTPz
cLtWYzgidIck+NXIvS0vE3PUGUPDiEzFxqAZXqCKRD0wi2x0ZdBkKQAm5xXu3CIBWJd7iIyhl/B/
mmbUhJ2VNMCckK91E4v1H5QkLMg/hm6hlyOXdsFpx6HT4rdSp3Kvp21RXPiEn8UI6sTmt55F3N/I
a/mowoG6jCwgP0DtwKMHfjLyjnsOFBdDx11iMzy3LkOPGQqtc241UCc2fmot73oI6n5ITa25sVtI
FTPu7DKnWKw7mq0iJa9T178d/sutXCkNb9LgOzCAQxGIEiGainvDL8nW7coGWHi+kVp16wTmBD4A
1BPUQMzNRD8P4Rvr8zX+RBEuiXNNoGvPUVJg1M9O6ULWOY+bSwzjCc4T9m7stiSZ3Rn2LA8/GRFu
Qoc7dZVTq2024mNFZWXaysIJBa0M+yKbejiub52d8mmpwZj+Qki7yNKY50dt2Fp/nUuQKF/oaJBv
mwWm4h3iKpukqKA1Jk3lzrTB/jmQzKYjt4K9QQ8B/5tIXlF7MiSwc7ml6Fq6eeywccyoOp6K7AOI
PrZgLdM5ndGLNUvzm3Simi0u6kUp7LOAzs/FzaC+L92xHB7Xk3XTJE1/+LqF5ecPCOqnbMFGXRMn
8I3+FJCn5EHGI4cEWqzsvsEE3qK4RlDTDEzFP19R1/h5LF11BL2/RofSbiy3S5E9DvQM9RhiwQx/
TlSrZsOez2CJ6Nd+P2erUc8L/1x/8iRh17mVG5JMq81rDWjJSouZj9S7P2a90lq6JgzuW17l1BqS
FpzhhBVy/SzqbiskfZtcwrBZrYlFZ5yohxPypY3k3MyMmKs0GHkiyKMN9GDovL3kmHM17iuoBV8H
l31tNxyLOL1TK9LlTzjKpLvZ8WxAGxUZGJ9yerdBWInfd5cTboCzqpga8x2VPbjFHeIypwXeb9Kw
ekjq8IrkBxoH/2xKDqfJM0YKjUggCf0PU/rweRPjL5SAA8w4L5tjGsRSTbjpYdXOr/hTKRvbHeZ1
JnLeswqhUk3P1t+ZBHw6vQyWd7+DhjPCaAFFBoDCzW2Wu/QdhlI90DklOW7rd++6afaTZzkkj3PN
KB6844qj+lbG5S1HFX1KmC5MVer2KXPdNGOltsa1BDPrcwuL6HYO+hHv+2dBx9+NwB+Wgm32YBcc
mxS3pTa27LCqETxMc8cB+fp8iaWUDIy8YT10nmxl3cCtXUWSX59TFnPd58580ZKHj9eoRYFEkPE7
ZFm8lldQq3Ru+v8cEhk9DYq1TYc0DXka24mj1KWQ/sFYhaF02WB6D4qSG9coaJaMs2Bi/ILsXjQz
asHAhghO2WH3FbivgG29GEjQRio2OQb/Ddp/p/NTs/0bV+J29JITWJHdlhONbFOi5Th8b5fhhCwX
oQ1nSxQor3HJdJQV/Frrrbm8a5oT4dfIUVe/2FRHZIa5+dmZVPitHhiGFfnuT/BdAlcUQcxz9oOf
bYBzENJLfjEK4JGcoPWK69YWkvR7StCuiRhtCjXk3Qn1nQs7gBKLdXu6qjziTC0X+RY4mLLJAH47
oG1hL76W/Qp+W01fqcyqHMSMqv+P+eYO/bNSC3sdLrE9R8YANMUYm5oUYidlcRj0wBa1om0YeJ6d
kfJ08+8abs6/+Mc7Dz0uXhTBwLzYxy5OMk319n7NXPtscIjXQyfU1x1LAYZaNwh3srl+wFCzI05t
gKxySesXonUwj6yLgeWzn4nEMiilIco/w6R7sL9oo2cEoeBGERXpYz6OzeIYZYikiO3SxP6EnZi/
C/5hhblFyJo2RLcvGJ/HEqxy8jTx9xcjBhXFTg//WCmru4zlqHwoVxsXhagdkD5AZpf18SoNZKZR
Lwd6/7SNKxgoVmA964jEi1bMH5r+xfCJVGaPEFeHmFmSQt/roZTf/KgZ6KcvfxZbTQkZbkXnJETW
LmSti1bWq1mwsTlsBe0k1p0nYfVSNv93bgk8wptIGdaCg7dDEtkMgzXWDL3s7/T4wNNOp4KAOmjI
FyG5N2sTOiOO7PeCBqkKN//uYzHFbaSs6reQsKIectCtPw/sA8sBS8jgBmxiq6o907Nsl91vG9gT
TYaEvrP+N11HunasChFDUbhaWaAkCHO+sATWU4ZlheyOWLrvyosjAmoTwSy6QJwVoQif/fdwrI8a
DX5rZnTzbfQFs7qOdTa/L1XkISX+MaD9vL3pAMA8EH5bjqiQlfYKgqr5ejd4b/inDxya9pOBc4HE
QIWKXmc6SfUXwwyeWdi5/b6/APpNdrbIUSS187FVKa03oXwUfpErdGHY+CM3KoCf5B9sNsdBoOHu
6ep06O6zFoVT4K47D34ehIzPePK9cW8p36VKTkeJI5YYUFPPZwht627N8D7JJ+eYPBJ7OvEOX+6C
jHtZV2VBszDSpKH1arvhEClZs5+m05QlR7yhLBC9Kucf5cwW0t2AXKKEp8y4EdcGCO8sjehgD4fl
93AGNnCj61wPb1ZaeX+ZRfEr3ecKbcFkuEOdmM1moEX0qVYky1nzitMK37RIQktjaj2HVVoNu3w9
1Zdv7pNylhfIwTo7I6fC/7oAcvaVhjuACzH6r/CDtYfuRW+R2dFz+McuGlhMTBYqdgBfMFQQq7nh
iLVcIEAsfkF+q+7IA0AfrpqHTNx+lXW1NQRwwOn5QoZYjV5R5lyjiHVuiknhrXZOkfcXpMhAUFMR
9xgdQrNC/QgpmdjnGtLHtKN0EyLJB6pwmF0N2+4wr/6uM6lQB0vI9NaIX1xSlYz8TFGJtY5Xt7XV
ZkhBewMSG+/RfGUA0rhxBkgGjs6T613XSCEynH4sLwBu0ojjAhHMJjGy2HvLYgBzXdDpjTsKWl0h
wCHjkF4Wq492iVuOba/YYDaSAh9wSar1BIOx3N+V2NVJO+esx5yrayaVVWKtG0LVe+BgXLff5GT5
0fM+OOlfRP3zFYS6tniKmjE18UeC0JrCVDdgu65PQP7P6kRmx7Jja5d320OxTeYBJ9wQgCXIuqMd
oZs7bFCGWwuctH4Mp9kXdvw/ISscjngjTzPcB+ITRiu1ZeaB1aPzLzvh0CVEmCN77zFrjGFCAU5U
RIHRBBaiBwm0YfviS94aGG7exP2UXo1nes526/qFYpp0XNTVyBpk6hr560IHsYCzk7Ldyl11KvGw
3mEYGCU1lHCHQXKxgnhzDz4IDpm9WjO76JxrX6srE/eRvIGP8Q8RutlUzS0U+ZWvJc/8w+PKxZFC
RF62RsWSqgYUtngemRhIlk6oQSWW9a1YBnOxKdzUZmoqWg2PVMRtJI4nyCGAYgaXfehmWE27BCOH
tLbIcjxX9n6cm1DIecAyPSPhHJXDm/yhEYwyHR2QDQeOs65bJHpiGHCRoBkMN08MBGOeXC1QqL8Y
lA3Ny4dGCt8KKo2Oz/CGFHICzZ3PrYBbzCxwL5MracAwSXqqh/la3xxPa1E1tE0aS4X0UieGR1hD
lU6fA6uJLyPeg2QgA6iWgFskrfi34+kpYR+A06l65LOtfD/TY0B/qTUh0PtNM6+B9wVa2BO4riC4
JPNt2sgRPOL1xsRjMWcRz93biv9tXsC4V6aiifkpmfQe6Qra9II6E1EN9i4Tt43YwXFEqzXYe60Y
yqCYMEbCi7atnStivH33A5JBKGe8/O1OwqnHJNMEJ87Sz8keInFhvebwFryUOqtj/YnqRyZXf+qu
BXhfbe0t0Ys/KqyHQJ2KXkZUARxQMd+Sbxj1vbzFFhrPSiLd8jKZeeyLIyOXp0ESY28iMS2A0EI8
46ro8jzonNDS+y7g7wLbzvLXpqJZnqHICto7f5ri8ZPciq3iQ0D+l7XuhCWe01YEHVP2LXt/Srhe
KbTWNeByJGifHmq/cw+/h9m5efNKFIWztw9qJp+hKZSMIFSJ7WlsJz1cPyDhLpUCyTW4CIFqueEB
kxYNujU+oOT7EvbBq3ivHMBxt7Jev+BoMUoNGQibJ3t3wAtIVOsGsaCH8nr5V1MwuGrwqwj0GRSW
OlBNXMQ/X9+5ocr9wzUt5yMjN/yx6tUAMreFkautc1zKVtK5VmfD3ebDllbQODPBRXfsAFIeOyxh
i1qDhbcwO3rq56N86LEtPAmikyBkJtr86KYQF0Kf+Ga1pdeO2ZisaUX6/GyjaYzy2ItSRECrerx1
LhYeTBZ11ml01OS4260C3Ow5R9r4ygWywQX/ArE9tmHagCRg7X0K1aQnkpYX6OaAg0UoTg8FHOoI
75L0WlY2amev5aETPreOdL2jWk+hzQPxOu0UZ1MJLZ78DD935Q/bWua2nNCGQDPdJPLg3Js0jGS2
dOZ0dd0Yoy+s0BWwvCGkoVDHMUcVtOlzcfhglIMdTLtWpijosFrMZ9JLgq5lGJIHr9mpvVSzoUzB
DMgLyc333niJUeouBVeHm438vPi8QU9lGoCZRzhCmDYIhiIevxDbdUhZo7GqMwyko/qXQrrz25im
SjY45/74SxvyyG8/YvqHWRzpBCzRUG3ALLciJnPSJQUYf3JxX4LXlc+CuSnwoK5IXuA3UjcHOJON
xrH+L2wVF1sGXp3UIzlNeE/r+IK/j3twhdL7KpGwsnpo9xe3S5uKec/93vGH6O5gWiWPC5VmL+M9
EVQAkZPHtQVrdV14mdlO2fm7mErCOev9BXD91gGaNTN8tx1W7X24zHD7LHgfp1umva2rf+tUPwfl
WQiSl/1RyFqOjKi+H4YJCGRG8u65ijmirr3QZnA9Ro9TDu7jXgyhvGvtD6ZQeF72iFqH3XWawP6D
qYz58hAZP2ZMSdOvG15DI2UWwDj0///HcYXDLFWFYNPZi1ORqHiqhMrBZjPNWTLXI/Gd64M0PfW9
lL7Xp2T465YFAGK9ns0hBcf1fnz0cl57EHoM/I6JcH/bFYvEx455UzbpupIMdKHfly3jZUAh9q7C
cWT3E+y7Dz1mvIeL0Q/9Sz71eWTfdWsuKP92WJztJU1pEr9eE+OWc4kTlltGc3C2buoiFSyxj2RA
sKADbEVBjtY9o16IPkpZTYtv+Hoy9ww+IpovzG2o2SJME5dfyjYZ9TcMhG5ty6jFnn/gHaaHsuHC
j09YFefU0wkhkEmi7DRdNi6EtWiQ7AoR8RuQXvnN2Zoy9iFViAu8fPBo8QOIsFaCb5o8CpJmnEYM
zWN3TCOTA9Q0+k95TcH5lNj8xtCYWIj7GOkwNmiiudLGrCUKnTDI5qmvvcPqf72FytS3FRrtLj8j
E0Io3+gRccDd6dPp/VS8F+N6hx68ADeiNWXGAtZXvV2pf3cn5EI+yWmqWvYpD25q1PTLlJHJWY+w
q/Q+Vd15uNxoquSwMAp5vCR3FLj2CgESJZX+7oprbApfYDEwKcW6yYX5gWgdUj6spvhv2ZCDRF4d
ns3pJI6rgKgphOy2hBs+y4vNq6Sv6xUNcbmbslA/lLFiuVU5X7VzTZNwAjzIrn2TR8ZLXy7ElGtz
viLwHbfRfNk6EIpfktWDIGTvzKU+vEO61vC0EGnZwPzD7kjFE1h9yqJRp12FfW/Le+vC8DgaKbAQ
hcosMWE2d9fMl9/vyzDqJxaMSdoOEVwNjQwF4j/uCZDRwbIJVwmUA1YMJ/L6iZKaVl+6MUIhJOS/
rXsWaYOBHvaxGuLeBwofUe1vb+YZnLYvA1pdBtUFKeEgKvagHABNa2PcZsnso/lxnZOYrV/IfjA9
82oeymj6K3vLSVOrpsroJSQ1thzmUnWzdAKlve8uRKckqTv8luprvSc9m0MiO3PeS0A/BdfYE8ni
TaMlWxkdq9e/IG/ekkUXQpu6HZdFXz+oTe2FtTgF7d+2na7MWd0FnhLs9hfSDBB06TFdBwNSVQfQ
YRucL2oCTx149K/wYrepA6DorfLL3A8A1YV411rnd8Z55urZ8BB5jIBsujjP5dq2ZxssoTTAuKo5
ZspXxUiNcZ84+J/4TYq1qmlcRwEZVsDVfJbDhPLS81eHSGPSBmHnLxKLZuVh589IWaDEJWLJhI/v
Y6saDktrltQ8niiPoHab5aphsuNlSSZefDEt0Y6JprBCUuVIriN8kFnNEBntJc9gED0tYFgjwKKR
pkD+M8qeHIIqomKi4pnMOTeIkorCz+eQJLeZ96tbyQynALxGVJ/jts5361bkOKtiPRnQNRpP7Zyl
OXPlgumxv7J1+oaFNt8PR+N8N6f/GG7xi5az/LRabNhEbnnlCVXf9ujfCzfbB5jUmcavBoapipPR
I4fD/yC3gxCqPClfkbmXyaclFyYIu8cMGE2yjOHrsLujXxtQKjKVbYc9otL77G29hepvd4waJWsj
U0gTmmjo/I4N1tGILBMnzcJBs6GBzl3m28TO8k7ye1ypEM7DCFqz+AGHqbCUh4tY4mYaHMAKXLz/
etkusiI+CI8Bo+X/39eqjgtxbh+aby+L9mU1GuI6BKG7X5OPmAcWyZQQchbLw/VLxQdnS/I1/tXk
6YPSB2IB7bZL1ohCvav0hnG11EiCgWV4uyRclm/vD2ZIfbMd9CuDYIoLTsdNgvyTANh3SQcLStxs
6jb7vNZjAWhaYEfJSNG+cMCSwxNqrU6/wkDRRzsZwBrXPTJ4l5AU3aQ9/ViFrehPpb12EkeEvu13
AOkBf5lNGc1c6IAcuZsd8fuPymMPJs2uStMf9cpMH48m4v3k+FXNKhraE1xyqI5fZAgUjWcY6HIa
+yEvJ7/zOVr/z8w+2k/wsshq1cd4H/C5YEi3HabEECxAG/+YqkThuxSzAu5Hecrk8D5STHbHyIqU
+RyguZSiYqaAqp+1iu4rqKC0rKDcWLdIWhENoexZFhmQbJlKBjgsojLWw9MRPE4Nz/1Vq5mpmwzB
anGGHCfbueiuCw4xTzPKtQmb/R/MWAe5ijFexCbHftJxLYhogGpwj+t/PCkjCNBgTNzMcMJQrlWm
oShxcevzrqy65LymRdWFBXvV/aupJ7elknyLdJecGQppC/minLkIuDSrJW6Glzuk5cFmS1jANAtC
9fvNTiPY1n9jF25xt2KwhvdmFbpU2tqSD4jyTRu4pyxhYRY+jFFTmcJgJx7Zdxf3aCa1oNnPKbLf
Cxb0hRHWzFyr0l0W1L+KmO2A8d80XWPmfbLMnDJKS/KJJ2CV3/vJlrdFl2MU00zbxrVSLaWnxBHG
VvQ0yLZKOxcNzqv3w69CqWWik9IPx1e39QeoXUjNTuwMKgWv4b4/Qd1VkGGpr4A/6u2Tj8+rptJd
jF09+lDSRpcjknQViQf7DmlBBhdP6LvZa2HdqazZYpHYl6aawnXdEC++/LXIRQZU5iMhOND/0c/4
UtWUHAFDyEelu5x6xY/RZrjsRuVLEZuE6PlHKapG2DZJ5tOoiWv3B707EnieMSD6hxzfvWXADQFr
uN4PNaFJXhRbrgdU8Cl13Dad1N8dS+//LaWGaT0Nbt19LRkXJQAnj0H4NoRzovCaFI2d5j2mQQqU
ak9pLNOpmUE71AqPQtBNTZbnUn++phi4Kd42UlH1dvLnIKRCSBlCCk8cGiCf+zTH4LegYZ6L3BWC
zmUNaiZKaje4YNqBFtIOLoAYJIeGi6rd+oZ+VC024L3PfOd81bJ9AOthXP+dSWhoySrtxZATyvg9
70DglIWMtKNppeyfZcGoQ7rfjN89GpGsWQySULNQl07MnC5g+/IWF6Y97VxpQK2bS8K1UeJlWGDv
kTP+Qtx+8dH8QfoS107TpIzxEX2QxSv7yVM/2JAaNFHpVpMo0mx/NQxqCt4zaqhDx4/NvMELBGs3
VwMhSvQWNpMY2LZA4XNSCacDNAv6ist3rxJrsFablBPDueM33vnVM6bUf29iBJwysvDCZCt0UUZj
y0s9YQn1W4s4tnmVUoQKRD54fkLKzPtNEnsBpzO88l0TTlnX/W/Ezkt7fUmw5MDrTMwr43lv5gPG
1bI2ZVlsuSEDCcl6kGouPQiEiD/Jp4b60GLchHOkVLddOgl+yJt1QrMrxMuF4O009m/nFcF49lHK
wzm9ybyXdrANrbL+4R9z95Hd5TuElk8WpbLCRqvq3KomkQJdIE6i5C5ZNO1EwZC71Mjhm8XlrPZ6
H7ESjEyjn4gURXTU9MVi5TFyzUyko2ps9yOOo6pQDKp51I6Qb6p20r9hQch17ukudToZeKZHX6g1
wGZZ8f15++MmTf1Hrqc2RLOb1SBO5xr9tdXj62FdYY9cHTCHZaeuKTG/4ei8oFILbwxB/N/ZF8mg
BJqLEatubCmLJthbt5vFGQ71n6tnKc713WjmPtu6dBZxkooMXANVpHpbl5JIlDzKCIjY5dmrkRLb
Cb89wN7oI1/cFtwlgFtUj0XzHuE6zfe0Cz9xSdcj002Iv7cFG8Ck4C4L/mPto/OhL0+YUWrMzNXs
Ix76I1aZ2Y2vVhHAAuCktryNy4oMirrASgyPBhcG4MhwkNiTEz2juqgvAtnyvI6cfQ4FKUFG2xlT
akFR+Hgek/FSXo8DdeHU499h/d9Of06GrkxqZLhotCNulaT8geU/tTHf8lkMDT8Xxwxh991fNErd
UlZZM/Z3eAB3qW0K4rkpbJGVmKUxRJqclV9fBmOFlwNENF+KeOt8IDOZC8MoOuZfnkTL1/29sGGL
0esliLR00Tq+fSxcww7QMPyqD38JewxS3n+6IwkLcVX62I2gZJUIHOFF4RrIRSv7uC9bON8AXRhf
x1xBcL4ALlBtYltnYnS+OMa/6y/Wo9behkkwd19J2iKlesu3B53GRA9BJXNeK/faZDHkkIuTX1lR
JdboRus6tAHVAfT32m3VZwxIEXxpOOi3kjZG8pSV/rbl/LCXIRFhItwNrlrQL99frhup2Uz0BaZI
J8w/tUUBE9XuD9iWigJhEcCPji4HvVu9l98mXMCydW/S/Ve1uVrocJg44ooC1lRjzLIXcFhYzOK7
UsuABSfcjJaOcm3wx1Kv5WQ1OJrU+/PgqmdSLJJMZ7KgizG1PGw97Kd5GsKgLTaJmzhh2nAQ1/9N
4zzxSFgj94st2rE7rRPVE0xuuHHu22El+2h9Jy5KUenvqIiBIz+CT/hwH8KFSojZEovEvn/v6Wsw
zwwUOB9g/pZ34rAu4CHlouWAe2Qu6l/AQX7b/g/8bQMIjZlw2+WicV6l8s6SHQ6hXdKUL8b6T9lf
PJF9TwFag7mR/KrM9bOpEucDrHJdPzIOJMWbdZ57HViL3EI+s6ng2DOkCrwjTXL0i5LI9LxJLtPJ
nv8ScFILpbMXYAsb3dw6gaF7RYqb/Rdec7YlPo6PP+QNXlZwt0J8blB60cnr7dQomnk6bHV7x9H0
Zr7I5jQJs0Pvv3dz5ztFZZctVg67K2gnqBssW04Sx2NYBv83MRlmcNfVeFEWy9hGZfw/btT57lgx
Zp+oMWg5cBTnIZMHAB4jY6C9tw6Z/wFjgJCN/0NktLwWFQb2z8apPzXNajoLhJLNaivSTJrfWvSk
QYDVMlLQ5Mfp4HMBelCJODJKJD4phb/WEG7xjIQ9kiMWW40iTKQHfYQjpDagSsQt0LBIloBxpfPI
Egglk59vFlOd5Rxyabg4N1fw1sLBFspSi3U6vRPzNzjC3X+4mH9bX7rJ743sWmytM6r3xFwi3xFx
JwIoiOiRKHCSfMqQxU1Ea4MhTb4yOkI7ihVlyxEuA70IEVe1I/TlBggUvcFzCX+0YHdYhgSxp1CE
KLJPkNLJoN1tm4RqXSYyIHgPnIYidue1O3RrQtOP1mSucXoIDB1JYH5phXU/E53pVVygSDeZvXQl
+LwE/Lf1jznknc6QPWJD6YT/6sQ7TThuWYPzolq1uuJivQGYursRKQg5xgDkVazafHcfqeTWekp8
2y3M3EdOSEfdv4lzvIWyUdEL/kkyshBpK1cmXgTHDdtme1XCyglUs10kH7FY7RsUf138cHQhVML0
vxKZ8jHJ4/UPNy0aWgpKfKzkiLAqh3NcgqtOclp6beiiXAdAn9MMEm495dpPG80SJQ1UD04x66kH
QQ8sIe7zDPKPQfwbdg2aj3IjFqU1pwg9NVsnrp1keOgz9+3Gr/+Zie691z5ZYIvyfjK67HbAQXbU
Fsn7ktBYYFcb7MMoky+UZr+dGwm06V3JBZ9MCb/9i2ysCQR3fy9SLVjCM+JUZMzZKWdkvI1x7ihs
v+jj9yHlyDjMZEIxLSmzkkcJb8K6KV++CYm0A+ENTbn8T455sdoTmj7QBJWwFjjahxZKg5jEoFGe
u8lwrMjzuBcFfNK+nU7HJv2t7jGl+APkmdkg2Rt+WVb9jM2azpirOeN+NPL7n/MK4lYJ2Isk3nYZ
rPKbg79W+7kNG07000gk+8uMv+K4vkbYGugkb1lW06F58jldUYV/iOLGdJhcbZ1huZfzz/p88l5i
eThiExVHnJ5RQPRtmSAY3uzGtX66ulzih+B/AnzQMY2kjcpxJSE0l79TfEFc5M0JaeY34iSKqtDq
rOPU/OOFrCSjnvRU9OWSGDNyIwv+1rZeuCmR0SK2+ZHcgG+K3oYQcnK9Mb63/J3zbgAKqqnaalcR
ZEYxQYh6eNIgqaJbzeuIsUaOMfKQJlbC5TWwt/kW8r2i+hJ67uwTL90skrjpgMGJTQiq7PPgOzCk
VQ2pQQ7rOCTCEeH+KMeEhvTAjSAfNg/OcdTHNhQhrsgeWGMWOpReZC/nYycA3F59gAiHGR/zoI1Y
tUiDJZVYQKAQA8fuKl7Msqo37eF7oZMjTdGW7AXTRtHNBKA9/6XNZ3IKwETYHnl3zuJDRoZu7vAj
6yg8u8ZmtsTo1ksaHLJAOX6OVI2dmLx3RQB88F8QZQrPwNwGfkk0gUi6+k3WtBfbBBRmCJaU8wry
lVic73DBPw1M4qyGAgO6kDV9gkb6e8Q61es7OLkoEYacp/5wsJsiQJ1dKsK6pEX3SUrLCiZK65fv
wzuVzuC0w629GTUk9vVcjAJRhfT25AMLfnCQsL8wcb/xsugG+x/WvaN9+xqWQp+0eO/PaqfkskF4
dNFAxU28PkW27WpaBrzqnoBpG6DyGqrw48Y0em3EM1VxHuAIYs8FI6/e4cZQWmajtJ8b1GnV8a8g
x+KfamvKqvaWfGQZoCCS22nxahtWZOUUVLc9YfxN8y1F+eiDsJ8j5u//DOPnq3EqYiNSR7Lu9xgj
yFhfc9Yv4zN5tKEY2S0SZeSNKzXUD6n+u9Lby+54aOk0qs93LbBOFmuVD12QWgUsvKEvqvHC20uI
HOJFc0FDI3wUKOemc4XcFa4IqzXarv7D0pO2I/Qv63LI7cwMw401kuH3fQ5iNZotFvhPym+oFXDY
eeIyzPAyOL2nw0y80Ql7mvF2pcVR30nufgv29UuXEdUSjo3Egj+XoZIMI9jILF/CH8L/0l0yjjRP
r4OcGbMd/w8sqBgGNukWpbdkrD0r2ZIGuqyvhGNnz7IvOAC94Gfmev8A+BG5BuIVFuj2xg96IbcX
H6onvFmvqJKhtr9hPky7a9Yt9rYJAGcui8AGwqixy83T1k3b0Ha04oqOWi9utorn5ZMAfshtFRgg
lMXpwk8MgwOXf+yfhheyJjToVPHc9ZURumIwC87z4cFhmxX4vHIL4xnTwaMr3Fws+lZQk+b8ldt4
05vNyL7hqvvk1Ym0AdysnTJec1yLiMPXaLX28CkflRSieC/oItoc8CcN2JxJhVoIARYyW+Uu6/qO
ftYrTECwxri1YOxyBYcN8bG4K4eagdu+ljoDS2++VF1h8jpvmyXGdvKtlqy/UP3H0LEVRXWWV15k
TTbyzLROuMIDAU00x9jYOd3H7MZEYOs/46PqP1K94GrByfwDbUJu/jMTWfrGCJnYWu2gNre5IfW3
vtJm+OrcAmEdfyxB8e7J1WJLTISslzzFsrtsVxJAxLd96H/zrh6fgF4tAxDu1boFWawF9MQ0dKvH
bLpcOF7x/pwTorgKbUkgvIQQYlO/Kn070xi5VS3nVXtP039VmtYFvCiTRhnfgvQ4KP/NlWf7oQ69
J02IX8XiIiPNKkM2EiH0nD/njl1CVLkvUmY7oiQaQojqFocNhLJA04usupwrYVthdq7SFnvROueT
kxyIkgBriExe+8Hx+O2u7OOM87HqLVAC+qbMWaZxPYukr8NVGddnFbLWjYzXOFv9HBS+rFklHt6j
VvJ7UAKdX4rkWnI1YgTnfz4/p4jfEnpDY6935fBb9NNG2mep/N+44mGM82tgCxRN50aOc5RGQfXu
RxH2azpC5VznHInCO85wWlK7XIBd2blF/U3HGXZtaWQUORB1lPrJji0wwY9hdRJvlcPkxgODFwl5
/sdFN8MxA330rIfx7/vI7lk9DwOz4E/INvT2rVS+6xdQS5fKPUge/P+XicSE0mk45/EZCP7Op2I4
l7WIrJd1tOE40m+FiEdPcf+novVHUJdphE3/VTDzXTzmfV8XTxISrw1TBeY+Md/GNX7a/+z9SVbf
P6lvIu0gb2X7Sq7DA46svdLFxrXnJ+8y3/1a0XBieYo/JRZXTtp7Hmz0XQVtta+GbxZtcI+tGH5S
XwEOD5d0ShD+HArN/bE0XFGO5EesIkByCySZGGeNDnTV7gDqrCvEhVNKR+lr0VvdQdi25/45T/Y4
oCQKDaa6ndl+7xAubAViXpShB8qWZnRPDZw3ymAuA6eIsFPrVWECL+kE/XaWmo7WjxqeLRanx8WN
nP16dY2C/IjRPow5LcsuYNQG/Pt1rGdT1E6bQWCLGv9XJT46vAsNyGJKvMlOlCsnoka0+dNpJmYg
SB8LCXMXZ2vRLlLvlQkDIis8UFT9ZazVc0DYp8MtceWXjsyUd9eqNGuIEJCSF0i8gP1OlOMVjDGI
LRK3tT+U1uV2extyLFet5/GpNTB66cp0e397/f6hvqIJFOWSB5oX9OiOQLitxrwtX9zGkzdh1JVB
2gSVgs2KUM2Vn8Qt6vHOeNOFVv0OWXMNPa3Zb4fHT2Ny7q1Wd+XtFftizOCsFMNlOauBzeVfxytG
WthA1oNQcfknRcny9sniUZYLG/pPoL2/9zYuNruQguclDH3XNHtIAqyzVOUgSNVuqziiaPkv52oV
P+n+bOpifp02QT36MN7qnqxQNN9XUzKhbKJ7YtvAQSc6RSdsBz+XmS4ENjLCP/xuNQKyaiDqCaOY
3vqQM9HfgiCPUtdHLFs8PGK46UviGCmRBX4BOt8gD314ObYYyjIkWWiFOkMdHrOXnjLwiwU++tmp
YruxyJUK4kSC7yLoP5CoT68wQQH17FoNnYk7pPpSsaw5zOy9iXzOneAw6L7NhGBTVGsv0qxwshKI
ZUDoqu/GOaemAHp1oTw6Q5IjeM7rhmt9Bur7pTBtMwLRhRkB73Tjogf/KOA12TKKHOxxxxYcyTiv
925w1ZowK7NB5mtqDKuNyakpEc6IkGgrNY7dMEK0SOlE16LsnAhDjyrNwsTKC8rVcPJFKI8B0yYy
iqLTCbhRtUzJiTnlJq6ZSFu4jgHvIocQwQj1bE5YnZJeoOYfoNe6Dzr1guNn2S0DPuXxhkADYOb0
BYF33at7Z7vxR/h3AoDurZ27TMqzoY3o8dLQhO33BKqyjyqcZMVgoTfg4y5Ot2XuHxEkXKtARhOL
EqINkC70pydaNZsFuTTulV7hgRHe2xlzzZRmmUELMe4Ugmw/AW9faIqAageWsKPBQF0bUv3Lpq7/
e/lIiuJd+Ik/zN/LOvKK7zYZytJ8VcqJd7akIBgKVhY9JEk0PWEvnToHTbrOxlXh53PLQxazhXnt
Yq26wkIMYhKY5r/JkPFmSYka/1xSybaYslIO5jv+QPUyS8brjRnm1DMlMr2pMpPdiJ6uFSIG1sis
CmgVznLr0+UlV/4SgAQ+uS++D5DJTKMiq+E9s84s99noE8UDnE6jyVX+kbJJuJ8JnXVPmeDAOxsa
JS8iXj3g4TTWABUHn7m9NpQ6P/4ba+LfBVHV/axSbfOSHrjme8WUbqS5CJQHPxqkfx6KsWIiY9XJ
GX11uN0zaTa1xW2r9FjrYZVzosEp7MHrQFb8nhlWnnnwPHgEIognjNZLobM967U/3dD+mxCJXX+D
/Sk7BR9PzM6+99L7UDtBB2qiP85TrSTCEzKNA0UGpgGcOZGgcW0QuCozFf5DJ6qrDlj7ePAngLas
twWwo4oh44m3n6HdAkulHzVifLSzje0gjT8lqooFfkZXMOtNu8r3RU/Kun7uckKRtDPu5Fn8Vteq
HS5siDNoc+QbdsNmIYdf02jZrOPH7xqB0KI2dMt2DujemU55qPpbZeNMTa8faRMZgtpJM/BprpXI
M4zh5wV/cbR9aMqNZb9e5QuLkFtnFiD98Ag7e4RS6fvuZBgI/NGEWD9vag2zg5oXU0YuW7IxLiy6
02/Vm0/LAt3zZgPVjxdKJdqrWrPt/j7oj0BMSvDinoTVGvUerMiserT7lyNE9c/s4K3buzfhOdhI
WGVNLvX5goXR2UbXm2WroD/ck9axMVrBxCLJ6toCwDUBQHQ7bMWsXpPS8lptbpzvLS/hovRyP5vz
un3TT1d0tr6Y9P0zQ1uhSENgiWLfAecTrBo9ChZzk5+xbdkC7rzCCdTNgOPHLLP7ASdH59De23BK
/lNnAB5Bm2MlxJ63PeAm3gp3ngZWLUCkuji0Iad/a7+VCWKuL5JgmZ537s1WQQXBPw5/a2YngMs0
cE5DwjmiEADnmJiqC96pPAo2LGZsFfy1q7R/V+OkJWumWSNhin/u08tl/GOHe1yHNHQQaBZRXcDo
PJcA6DWR2QgND7AqvcNsJ/yJWrjQa/Ou0+73yeap++e7vW2UPcWzL1OKB+vSDAmxAhIBx+j/UJqG
JyZcvT106lwC1+dN9DRkQHjnqF2HcD1Yl7Q5PZjjcsnm8SJQBsPCYiLb2iNUn7bp5pxonFoghCVB
NjlVSrev0/B+GqEyLTyKkCREh2KRPR/e35XBwhvEMg62qbwsvhq2WWwkv9ucHzJJ/2DJqABlzNJY
ro4TXspG6T5DGzVFgui2NtKbdZakpFPekCnzL9TkobgdeSOWGOaMv1bs8qb13WOOA1f0YNDHyIDN
PzCrhzGRcOHh2EVvi6mZVHxLGxb7qm8omSjXlbgXIbALRx60OgHS3EGyzjcv79ZkdCmqAbIiLSNa
66pSpgHNkOXlzSZR/a3enHyjGMhZwTLWbYYQwugiAVo+qkLkCxj9vdAE+pxohPL7PV9jinmrTrW+
pqjrFHjBrOaXnnrlFX5o9Cc8BE4gYcgQoPJryqk2Nk9DZQhqgPz+ZC5alQ9i3B8ccCkJbD363AUb
X6J6ess/NmYjSzLFZJWUwON8M1wopW7LsM5/qyZ3JB557Mz7oVfLAWK3NC51L1lefo9ttDxw2bji
DGfIFqVYlb6lxdZI5v01y3nTONVebdWTIJL7JGXYUOyqmQk0mE9oVT2PJFlTcFnaKXes13pbUx2j
1t4DpK+W6cIfGDV39og95ebywmjIZMn1pAT5d0JwrwkGWI6sa9CZCBgU/tT3+hDLqgmBZ0mjZ+5I
bl3QWQA0wtTbam/LMZacTptPP+JSEVQzK6juY5aQqrXgQarE+/WyX8NsCYy0jOUZcU/v5aTo/o8O
Xj3Muj/y77lgpnBFlAjigNLAa8fWXoq+LCCM8CnMAHTzE9cNeC+BcTCl5Ujhl19+H8G8x0d8VSqg
zQYH/YPkCjRwlGIBnhngWfT7sbUikSap8z7s87WtUmkOLFyuUd4Qq9FJJzef3OokmIhYyUut7IV+
9Vmu82oKNVk7zvzWmUE7ayQj9pj3M+ZkXb3ojOWeFAlJSLDFYifLa1YsXmO0JWTF3bmTe3meieyB
jPLAA15FX+cva9Seu/NtilU0sAmCOQPYFJbQWwQHhNwrUNyCYHzr3pZZnX2mWAEp2qjGbSo4q47s
3rjnWYUbEi5OAamKzLMzXcNbG5e0J2cYg/OHre1LGy2vQq6JM2xFmbhwTyCbzEI0GVHptQZazIZW
zzdEy3UBe780xqlF7xZ5apADWofIGKogEK0N9BF8kYZVwTYmIkQRwwkbpCZsX+nbkILt3bZNHk7J
kyUiEB/v+rw05NoyVNH8gmtHHPVcb+QCZAIa2oEBfLT5Bzm91mXZyfhh8k0DkMZujehnreTKQB/7
NXBtm7WqbFz5ntAvpWnuWv+DV7tlHxZhnrtkYwUdV6mlRZdYVQHAPkSaqfcK/KR2tFCN68z9cl6l
4ZWjxEUiiJcbZP6I9B/EaAoXMgwxKgs9iwud0eN2whHozcphP87bq9necGidF/Po4CnkYd8VQVVK
FhG/6/prvTOwK1jb8o06YiZy4+zFlQiFXi6ywnczU3UIWhm7nKhqjJC7Yz98z2W07HQUCIDZk02k
o4GQ1BPiX6nYUC5j/0QFcu8941S9uhvbAait3WPBykXMVYUXFKfJAV9joXwwISoSCstqvBKU35Y1
VExlRHcZbMYKe/MRnj4YzK/w+EHqd3q/qmUJCd2pfPmilJg49mDTvpSnBv3c1jtnv+HefuJLnKXI
KNNXD1aP/HbVJX9zCGcVRnhhbx81Go6T4Jn/j2tX6XUnNYYyhD0xfDcLE8+HAP9ra0TGLLRdyvd3
2Lo/bvgOGf8juG5CaqNHPC2XTEyi8OZKi67jIZb/MfL4zzQn8jdV7Gwhmp6EpKsveaJMwZyhbjsd
RtMsBOBhrV76VmJKLyB3yVwdKzONxnZjUAA2Fva8ri7UwGMlGcSoiWlLXbvI2yZGLKjoRJAduTv8
M3B9tpYCNW8AdZ3mt89bw3/nuvS3UWW+cKKtx4TsUQrA5aBU70yFz4usG0+AJeEdauJASSp5HGjv
MigUzjVLJNLc8IJK2GH9evxsAJIYmoApncwuDkVPlxJZTnFBpEpdY0/glRTcIgdbcViOg3tDkpsf
odne/3IJNqfyJHfsXdN1XxPSW9ENasYETKd7ux3/tCoKoydIdOga6iyI7r1t5bFofRryVVkH7pv4
RwwtycO/+F5g5NndgT4hdva4PH3HXCK5prxBnfFqE8MhRo3TxxRtFnTgEBfhV+NR6on9SpS4gyIm
B7Y/G+rs0xvqOzf0TbvL4++iehxLcLv9sJacXKjbAcAskWytAf1hQIUF7gYp+Sf71WtQew9C4/89
2CFr14p4tvPBm9H6MyVRbGhn7aECay6m2+m2ujvHGQNgYfzd+/82ZnZH7hzl2t+gnafeG83clssi
RB+AhPfIG3pCDXZIxK13A28tQKOYpIvt0VrRWkbdLldLkkKsbmepJJ0ufUiyZsVjqYdpV2pPtdLb
8XOrTpU5aC2PTgOaBBUdyrKkUTfSNe154PxI5wKFq2KIWQzwEIMOmapdHIRpWVN2VYQHlgYc5kKq
vqLuP1IXUl0eivOQRWAhwCr6vDEH3/V4kdF5ojHJdBiZqZij+xDpONIRvOgLLOxTgHKJVGL4ySMx
NVsS48uNjLj69q4U7N7rRvw8/BdTY0BL08mvUz4hvuz4BEN8aL5cuJGt/+BooikbBH+zExN5Q7zc
qd7NvBHCaZsUtSxmuGI4KAy/WpIq4Itiv59yYq1ttwUowUkTiy7QNXn9NML8e1q8E1u5xtxmE5bR
DhY6mB78CchGsHmi/E32V6DSS6hFkzsM9BunUqYd+dfgqkm7afHotBrSrHGyondutxEEfihOz2Sc
4RkpBYGfytX+L06JC+F1K0wHrsw6VkkWPGpsNNeRViUHJU5Iny/aXBe92aC67LdyLNM4Jo/CTi15
QVt/vTrM9nb//orEMouWhCiphwKUhVVSDCzsoOOP1zJ88C8L2lBXX6p4gur52WKuDFHJziBtiqki
hl7KrDZtL8NWRtKcok9xi772fwQT5Nktuwx6OdYQfRLzHV/jfuZSB+oyMTCdhsAO8p4+DNN9Pvvj
pKfjjn3Xd/LRAVXKFEYIcj/iCqsEsLqBAEEMnHnB/0foHjRXu4F+Bu0KJmKdGb2ZlDEnOVhEg0Dh
8C+mzqr5BNKyAMbc/lpYcqICyAy7FQ2n+Zj4LfAF2/4Z1sTpA+ada3bct1DhqGkVQIqC81TPwm+v
sFPOzVEbrRWenwp2CohLRlOhthQTS+2nHfam//FvKdd582MFOmdnQsF+NKhaZEwbHEZeuadyFDqP
4eluH/IrNrVlQwQ7eIsHO6ICFLIIoqEAZZ7+zmJpe51hoQc0mzt7mY/zxL07RsE5Wboz/d0bBpGX
U4edfgoi1MuhlBJNNmpu6JcPT23SGj1QfBiw4WfNGozVML/yxB5KggRj0Vtvu3DKxCIIHwg8Qwpe
2zS52aXepfSa3sL7P/1PUGJppQqw1TrhTncbHCc2+utyQqRBij+PrldMQQvMAmFXAVXJHpGXDh5P
F+QVYJdZVmWZWJLjn/yVKgAJGRZpb1AyT0yeIEN7kI6PgiDMfIP3xqd4eWR5SF4/8+VLvGKOo9PZ
V70p00FBDwobUGkv+6yNTcixRtTt/35qyw8QOzM9omGhlRPHlALlnFc0HP1OKreHWZ9orBfky/jb
c3k+GH0ixPy5qDg8dM3ZyhJm/Wt0TZSgXTYJ5TB+n1G1WuKNc4RPHLiKvmvT5e84DHpt5ZYFM8tD
bN1audaBeoSvKJ5t8lZQCiHC5AoO0/Tb9LplewczWJAHQA3aP1bjVkd/geit/7UCriHjjyJMKGWi
7BGhHg9dk+5r5gjYOZ5WXDjGe9h3xRYwgrj7h+aZdCzm68NQwq5onRoHLCSHkweRTOzVKZmHhZeY
BzNkpOHjbJo14/4aNXDB3QyWUVm4PUKWD3DbHAaoCpksVbL64MZU7tmm8XEjNQGKv2eQzvdkm2NY
vK8Ip8vL5nhGU9bLc+KKjsG0YKRf9uY04z5V1383XoT3Z6TQ+xX65NQ7I0vGD7jB2XmXcLyGOdor
lCHsVvoZs6BzHwcjhUkS9mhkl5512lTcUT0OgusQ78HWkAFguTy/3/qyNUI4l6iEZE7f7imrm5Af
lTa1Uz5ZVDw5BPrb4vt1LYdlvEoMc9Eqv8wEneArAC9uVg++HAKsrrukY95I3NuLP/baooXKdxaF
XQ1Y1rO2NSTL/vgw9Z9kpuL89zSlpzd2cJBmOa+U5NNTyWGLfG2LE5oInW2/vGRIKpEofMiRHuPW
hpOzxopfC6LiivgBY9AP6QDEeuPZt4w9n6Bm/dObRU2RCtR0Yrdz0nXL8MecTlCEZ+AVmAyEQamF
Jj9sbydKCbKECqjN3Xg8x3txq5Ym+igubJM3YQFFO+qBaTD/dJnM+eabPLCVe5zE5og2gzZY0gGY
lRxLji+wwrE9kz1WIYFG4mMuirxuZyW5KEHEsFhpX7GcWn7+qSo2Wf1oU175KuNbn6UpKSvavRMc
3wVWO9kwzaW4gOPQXtLfqkVJ10nBuu4E3x5HaWW/vfFBaIueRrVkD4iT9rOkPb9zqHUYU02bSqtR
c7jIae/buvncUxSYwTGxeU1jm/dlaEN94+4R99gIEKPshHbKegcAcYiF297MKumNkGDzbqgaRyGE
5tym4IbZueGX+5mR5ZAgHvbfFShosblNAO7342iZJ6GGHyQEBGR2xWZlEpetv3/dd0DK3zgweZ0A
XnwtYkFgnzPROt026hLZPN0yZIAP3vqd4bXqgIojLD9e4BOgaETGUelK/1jO8PPNohuaEyw7TigK
58J15/OPzQKYpxZVYOtOjkoNxRnTndYMUzuEjVpOihfOG5PmyRjYiO7X27x66VOXmU/X2Sl/QvF/
8fysGaawaeWx1/SqgdSg4H0zyG+plRErVyx7tPL+MfeEYFHnJdmXhSDBAU2X8e4Y/o7AR27w/aEd
VpJhn0P8ccmwGB1vVE/rsIPSoREjJmn6MhQ4eVlLAQ1cx07U5WYjEqYEI6vBmZbHTY9j+wY6yHGa
VrQLA/9pzrQYCSz9vmTY6KefuTbSVuhhpSoGeQX0woN241UKjKmwel5YD05Rz2sIu3pi+aYNkYvj
h3eyOE/x6aIo/0vXGOLEYM88zam2mxG5g3zix2yduW3eb358Gry/juM1uH0pGJCmBkOQ9IvB0MqE
ZMSftWEJ6s/gTxOjmrIfTnfQEPV2AqIgYiRcd3NZMvzb+DgEBXASyC2SmYO+to5ODMrL8kcvkhDV
lLseWP68eMD03m4UNDT7bw7nveKSITzoh/J2EXsz9W3pmTgrmcdBar7PenQ4JLlkFAW7eDINNgR6
k8nP5AnBiioXRJvwEMvaX7WjvgYIwrFDlLANPYNwYrf9cjda2FjZVGvnqajjo2yl0R15xpIrzA2G
ov+jjaxO2K5GBgsEO5WDoTUfShc2tvYaSq2qbYFw/DcACzfOB87jIBkYBROkVQYP+WUAkWH0hvtA
InVcw2KhL8I85bDm/NqG/GdU55vcweBmcPtR3dLBi24gkcOs4fIEoCOlAMp2ZFhzdN14cal8xKDK
y9tLMR9eA8Bh/FBTbyu1edaSZaq2OSkAUVWraZfsJeNer/Z874Bl8adioHobtqNJq5BTFvlboSns
jFmb6/wkl/bmIji+UnCswDHs/16KM0IKUHELmrvLn/s9kv/6LQswJpX4akMapx2o9//J0i0p/i45
R1KUJhlprUB0SS9djshqgpYn/0kI3BDEVLZA35SWnD07Sk486uu9qI7Fl8Z2BS6cGbLiaR38p3RO
xfn3n+GBHQMW5aOaJMz7yyhrQQ+WNMtoMs5xd8jrH1NyO/k/0V2z36xgPfWipP6wxmjpjxvsl2FH
wuRpI+i8F9os5PA87phd1kkfbXfQNw+t6O59adiV5+B1xcky6F3geN1hOtZMcQBMvya21qZcOszv
lpJ8Ftdw4PMEjXc9EExV4XVIvOmNgLFaEsMI1U2rPBGlv63ed20MkOsUyXvQml4dFS/yLUt2zRUh
l/RlbShcBe4dvXUeSpzlkG2pWDJ8u/nT278WuEHw9YSqVmu7pypDKY8pQ6cLR35vvLxU+3R9Mte3
JqpoBDFHURRO84EduSkSjztif1uoxWxC59JGv4x7LrnXyZg6NVfGWOZrs9x/E+3AsX+Hux+56gwO
fbjq0XupMQBgzPapI7VIoL/xa7rmpl8sKVJ3gbEElTxFMIOi0ZI/cV9YuJprQO+DM5ANrGOSnjG3
19gQWOzgdYPIueMQ95mRM3iJW9AWxRG0GPvTOnWL+N+tjxHDPespbxYDaEeKI4D2MU9Gx5mJy0vH
MVbGvCIGwUzibJHlUz2+yy7HyyaWVC0h46kN7X3/OVPfr9MxqF0sJjl6Lhl5gYnY3KQiojxDGwuJ
596jzReJ81g0XW2VJEfxTqbd6y4QtHrsiGEC1yn6AcDUDJOhs5/I4HxOil5/cLZDrREg5un37/Mh
a11oWLPfU61GSWDVbxkpDLxNtjNr8TZ8X7rvNONSA22go4OjUlgUt//vnKU8OlBTVzdEixzb3Xes
avulJ7ImGhjYkG3uIDhSqF5/CuMEYFxGa1NNAEen899Ltu1ypqDLrEyx1/XcLl5oLKkOJomGlc9f
XNqYl8RgMHGPPJHHf+svhO+OyA/amidr5m7ENylBFa2wjLr/TiekB36tAMdDCMnZ4Cvjc2pflsen
1pnGIodL36AP5ooY3FXbpN71zTVT4pso9FATDD9n25Iv89/OEiNEEjRaJ++YMSb8pLyv5PnM4Hg3
O6/z6zgoj+EVKd0XatEH/YDwhbD/ZfzmvlW93Csq8nmX8jtWNSzU6QwqWQHqtT6qMpIPwyWcd0a7
pSFN0ZIyerROoEsfhmg8xwyP9g9kKoxHxHA8kKQnKzV9dHxEvEPo2I6XKW7cKtH7Z6qoNlarC44Z
kbMtGjxaufmfrUvkBDJcYimoRvQddMWRgs9x5vhcUrG/NkFKXK8BPfmO0eCZyNETXP/pnwW0MImg
o8M4nfY8B38VeUfs7u9aMVLqlwN34PNmXu1sIr/9fKtguPTjDwifrco+etH0YJSk2pAWoWFvQMb0
p91+h8YPsf7yucIZr9klse+irE1psZW2dYPCaUjcIdqbYut3pXcndgE5KhXpHD++ZUb2RxwANzP6
jVdV+1yYGaKJPHrSbmaVA3AbJGv4MD0hGMSxdnRvrZhej1jPeF8H4i/BVNSKmudIvJmxroq+XeLO
SZLwHu/QZMlFHMCIv6wIuuTFBRPS/MmAFQJTFIFUx3wZxCBWoYf9dajNtQDct7s4OCognEN100av
re5tJM39lW08jtHCJYG3uCff4gor+Nnlb+4GHPJWF9nIkGZfKrAVaNI3KCGir+SDgD/JC/pXJK2b
GYleVaQEK8K4f8Ir1C/aaAnJjJzFgbQWm8i5mTkfWfDW0+YpEzHNbnr6A1F3ZGvVDHkhJZBz1mz6
27yGS1NwDc3MxtCecjnMAm1TxjHoA63l7keG7y4+M2AVHf2LAFtH/UPaCuM/aPPh8XlTbNOvMQuQ
oLvo7PVvl/cxKnQk9qwL514H1D3OXMsNKs2LgPyp0z+ZT/nAfkNFEenRbxm8bwVZudOLNU7YCoY9
jPy5Uaou0EO2Ht3NBuU4v/SAdDKapmv4WyksSTjRxwRPhyIFQA3ikZjT4teeWwTjYsn4AGX3yYsK
CPff5R7coo00wvdz52QqQlWtKUKwzjuS4RmlMpMom9LAocnd2jGSGcqKCdLwgyC8PFSNr0KYJBcM
stltw8+UWVmu1JK4pCkQYTR109xlOseQHEV0QnlZF43YRBLmWCpbjaUEq+4qPp3r9R9tHNNV71Xn
Xf7SEY70W80qB2zPAXExyhxTqgwrzyklxwSdGC6thdKoV13uaF9tBWwCXaASEV68u98GbLwO/Xdh
+cDEEhnjlehOhujEupUIusdeH90V05NCaGggrz4T5xfSc9oxJHOo+9ycb0KBXADt+RV+B7grobRb
Zdjg98gbi8iJ2SSeBy4+9cji7E0pLjxF9oAV6INZ6MFp1ntTOxNnUUlc6LiNxeODBoF6doykroxG
YccdXvjvXqpBTGXEKqXsmrPavCIzLzMB2+tym/LTqjdsaAPT9WMjDCD46ZNrVee+dQ2jOVxTtJrb
KtLT1oinzwPMfCOx8XGmWJ5xERCzUyBLvndKWHfNkE+oMT6ZawSPihzNAejOCWowy+1+BiSz54ke
i73WkWNd2dotX5+BUwD+qOzuV+I5WcI8Vas448WNKBW6fJZoqU7an4JeKFDMBq1gWzQvsbooTpxO
2sQA5FT0wlO3OfVKHjsQULHs4b1An7MmHDg0ydtNZsv6SGapAhhVmuZDJQdgJmp69v7Wk3pvQpN5
vj5mgiKdX4j6sehEEY3MslCxyrmMSxPk7Q0GHELiRI77RP2NBQo97M3woGf6FFk1dqM6VUjmKhg5
0anALRGIC20cRmsKo6NOEYMjgowyI9S7Phlp0+gftpS3gpQMDt3IMtsp5833mZMgyPjYlX+3RX6l
9fh4CEJmeLG0qh0672GV8MOhftz9eQ+ytYCmvWn3CznP2AMhobke6QVJUAPldEF4yIcMdYIbQuUo
+xeUPb2x9fMmUbpOvU8SI41k7+jmymDcVxWCUlKWT0nQw5gIAwSYbVBt4CurDlzYnOyg4mvlQeMi
UhvQlT+1pGDRDpI6K8M+Pm4zNPb8InYq43K8Hm/rF6nWTxFdaFdsvH6Ry+y6HpXlK83LxykVUqw+
pLcaFx0aC9mkUeNt2TgQtJ4OEhO3t1yh/tzA7WISCYUgFIX3+itqMWOxj+3WnW0HrgSNN758tviV
PuEA+vHM1KH0WJLIXNAj3UWK/mh93O9B91xaN0gT7BgQb6rFBxMAw2TPy/mjCjWmVBJR2QeiGE6M
P6UWHcsy3bIkeTaL7IQMcBcDhLr7FxTZ3FH5sitr2jOHyoTSlwCWvowEai1S4M3WhyVPoRtT7nDC
GciOiCy6zSaAFpUB+hvvHL1x3gtKXurD63iZVb7BCxgUM0a00kGVXOi1gnCl6zOOxZ+kxeFkoTuH
4rnwE0GpO5Y78J5z/Vt1Nb7yuPQnpWIVqMCLgWu+axuQn6Ty2RfWb9L9391oevLjGURAx8ng4pJk
o+ua/aOQOJ2aCaDiEVr74bazXWNMr8iHbLI2aVO181+Jb7/oe5Jn0PP6X0AHx519z6SCT7NzHHje
04FnhZJOOt8pgl4wtYIZb5iwII3axaGm0/QCup72t2xVBQiuXrj8YNWwMkkWzqLzXBddlRC4PPed
zJkTt8lVKl2uycdugjMijTD1Npb4WNnw1QmV66xGHEspfB3JeFeN9Ylw6gFhUTc28yGGWd7jVoei
K2yeMFFRLKgbH+MarcmbKubHBxVG2TtvdT2X8I+vBH4HZmMHpMXYpEtiopeoqdZwvr2rFtjx4iHE
8cHzNGZWEHO850O8E4fC/LpZgIG+MwSvg35ck2SXsasapY9V1UnyYM4wTEYUM55AooGyPCHCsuLW
HHp82uZDNnoDXcjgOutRj5a9QwVu8/HF6Rn6hrkrS5Rl6LodU/6FswrIk32Pk3pMxwXNQGhz3rdA
RA6CbjghZ+RCfmT6be7yMT65biy7rdunQSFfEBxx3pIhibsR29vdirLMIVWo9iqCkfNWK66QV/8f
G1X5YXv65lLGoiEKVB97vQHZQ7HY+maZTaiKTe/gJ/SGdOV2F43YLpA8VYZ2dUHtWISIJlTxC4AM
j9Ux3FTYmGvtGzAuy+vISMgjurP5pHPGeoW1WjPJMpCjrTksrMjBi+/1EGoGW9c09DM4zhh7QoYm
xgj5LLhnzHsNGkJzwEy0kfe+sIK3wJAQon9bqw2E73veHNt5nvOsP70pODy0Geq4cQSeLvmTzNaw
xcpypwMs7FPqRcFH6LJT9GcvUaj+lEdPi6PyEO09v84eBgCQSH3jZGoMnLIYYXmxh/OUl3FH9aZZ
oJL8p3v4YFkyn6qTG/a+pw5FGJ+BSzh/rwkJC6YI2X8yV8GhpJ+2Wxub6GkOCwtqev/wtO0Y0OBS
IGmdCc9fZXIsRjxcWTX0viTEi2HaF6bi3NdMb1EMkZvozcZOo1FdfHzDRtGA19QfkaVTUl4eeIeT
2JyT9FJH4erPMaJmtItMgJe0lJyHs4F0fthp5mri8pw0FHYIXgocb3jURx01qSICtfk33JCQqDz7
x1A55h79ZtGZXHDJR8nIenHyytrzeX8XfkvlTIlXUPHGHhUNuKiR4J8SAWMfda6MfE8bGJbRTq0Q
r2zYoMzg/fO2IvyFsRFieZebQfqIHxkIjFkLKJ9OvmsgvNW3zZ2FJf0jsbANcmMOKC1CNtTz1y99
aVKm8BME4utJVN+2P8k/Ys/n7Oavi4Fgn+LQZyXXLgF8cQ1UMWTxKq31gsAzGQK0dZOqmoF6KmWR
Cy2W7KOBG9J+Amv0sStXb/myczYtxJGcCIkUp2uxkTuOeynIAnISmbI3ComkWkZ0P1yKHWXtR15h
UX3JYYy4wrIVTAAe2x1Lg8kWJdKicYXcKftn+QI43ysEfj6QJbpbPn/ZSCObVh+eQAIa+nv7rhaW
kvrxNySQiyVLN71myXreGNq7cUTkNHEtPNIX9cQKXzs8NDKFlr9uhBp1dtlhUmO1G7veJtO9Pt0c
9AtRBWfGQ94VJ8o8R+/ZuSd9EUQ7aIjxmKgAWpLu3YhQbuRTak/wcqBNErElBy8T8zoJ4cAZE54N
o+O4NZRvCQnC2BlXa2+AnEIvVwVbHVybS4wZmTucPrRhsTcJTtbvmgRiu8KdFgIKKAG0BG7LMCAa
3m/ZHm+2mN7/c+BciI8HyS7mxWyfgjkKsgZ6JBAWjZRO6QSKjtlf5bPh+4w4o48yTGZtzB6TDnIP
9osIszFIXH7THy3Py3DE4Kq7AuVrTDOPe/E7YApxeUB/YOmohED07vI0U+RHufEO5i3jyGTg7YOm
QRFO2odP0DLXecT+4QB86+yq1zCdX2LUTtl9Z7Dmyb12Oxf2At++NFmDNynyJ3Tj4DGR9bw0Jsn/
M6Wg4Q9JHFAjsZgMT4qbyLMSy5lgqQFE7xdRN13WaqVXZh4a3hhGF2w8LKGj6mm0I5nKx+x0Nxkz
Uh/9Su1bjSYjHg6dEqpRdKGhzVR8Gtmk2uZEjw0nOwrnrGjE2FwlnMQdkEYj4Tli8l3UCDOpFdXv
/sNVan2eyMQ5yTgBzdWgsVqEfhOp/dyfqiyRIpK6O9YGQPEno2HvXhUzOCBzjGDWM/Wb+ZazWffN
eKs5VGO5NFSFGu3gg73gNk62Fe0ENzhFnWzpaGDGtuzzL/k1WpvgV3RArVf2L0isPknYBx1MNPTo
MvGtmpgFN434gDDsRV8IfCH0GjK5ParwmW+p38ageqwp3vgLvTVHzRQTqSs4d3Ai09tXq3j1ghBj
TTMWKRven3knlMAJhW5QX6gRNt7xAGtHphBZljMwkBD7v1sP1mc0YBDNSU7wvKHfChhFKwAn5mpf
Z5DwO6epNPimgpZJ5U/XLM9BFgZIe7QLJRvFVqz2tBN8RiUgC8v4fR3D2ujy7SP+fu1al97OS3W2
xbheTS36LOXYZWdmE8gVmIzk2QyXxi2kHPED8qP2F0XgRE+HLxwnCY5CfqcTWcq0Fkv74BH86kZ6
bGA6kPSnXIlGpJAVihjJew5VzcapzTkzIEqEVCUE2yCPlOM0WRqn2gzKaacLnnLga6wex8wg+2i0
sJEytTx29kxMqVtbgQzSwQMtRS5Kx3lSUmEZGKlXps6yuR+o12F0G8WM/w2TAkhNjOz6acMEhQif
19wBSJwv5Fj6Fn2gUpvvuz310CpwlHDtfWOCn6dCtSUt6UN37adOqYDpftsbuEbz2GSSwERTANKX
iZhksX3MFUxffWeBZA0aX80vFWL7PquxI6wGNMAPwLrhfDHddHOM68E/ziyzWCWqzVgZ3zi3/Lo/
QzDtlUSCNeSV/Wj1twxIk19pFbO7beu4/Njdh54i1HmyrbjkC9mtgrt1A43CflT6dy/XGhOBoZue
JfJQ6T9EGAc4q6Rg3Ij/5PxJRgAmOlOML0LJthWQ7L+B52UoWOFq1KXmj4oH9escpZwmoZNob5Y3
KzboqIJfpotoGxUrcz0GQ+bwk/NqGs2QgVSfPX0DO6V4Dyh9nWHBQSsqsYcYiqB8CcGCHMUiRCbD
BRnw88MOKybfwneTKlnv09w9Zh33VAT1p6R6bef6seyjzJt5huE/wqRo1QovJQ0V0moFiIG/51nr
/fkPdBGZH+YHpsZ4DPQXx/VW0M8g2mNANLakwfFLjDpSojQ1xUp0lZ+iiPzG/hltatlTyes4qmzv
ikFnssLN089GXOz0+0AYVoaNh48A0W4N1zl3JlE2qEjMhAcxgy+gNrROGSTBC6txtHiyUFgGnXCa
eZuxzTBLomnLGXjPVywqtGGcgH5tk6sPOHUAwUDyCvyipJFhH9rYlL1V3GOCG7bRf50/n1f+pkRl
XSmGkWYP8r8Vwf8bEzfW4mrNiXmwIYfDtddPP5twM/LjdAho1Ok7oLlUWOGVYzgxsCslKoaKN+34
YuLSEAtWeDYInJ2dhG2e2VeNff+juYbkSh5gdxD+H0CwfmeWjw4odPBlYI+WtLmTJUXl8qoqTgy8
/StxKvmRTvBTsioL3cP+QXd2YlePyqYIhB08wDGObvfWdgH9Gep+hUqnCyQXndjdH+zFwBpaqO+p
1gb/k/rRLd80UytkBBNpVs9yDquJblkCywbQhq0BbacptoVYVT8c8exm+DInOw81bK/9Cpco1kXp
p7NcC/iKFopjkXOQ+9/y8gSYNMz8WPtnxavo1nhFKWkhv4Yz/p2d85J+r/yrpStG9g4LTfOiEC2q
2QIaE9+sRNITpZjqX499A+kcLmkHmb9ccRecTOoKF1+G5U/Vo24p+05Rh15/GRaaOrdPaA6kHp5u
AafebbUYXHoIDu3W5agXGpLhqhC2MRtYW3IWUeJGrRaQhVcmW+vidyCbhke1Fno3KoaBgCI/0N09
J35yHvtNmrcgRXV1NalNktQTeBPLf6RFa+ZeyzSqIQWi1mNaoIGC7G04Ke94k/AVmOvjyb29EF1h
peB4icKlcX2jUylicWhmgWS0V5SL5XkA9neIRiLpWXhImmup12qjyWBZZ2KS4aKXxGI9XkVM5VqZ
HnOOv23jFC0EPvc1A1v8de0nanuG/oAOcemF04wbWnCLXoAd7y0BGTg02VTz2sA4JcmyviJPIQ4s
MfSPYLLywgamD/UjrjRyQ7VzybZ6wD1ki2a1TUEIC4rfV7oAiHe5UKIgo5OmHfj47ed8X465XHXG
5CcJ0c11hJy84qEcANPmcaW/a4C8G8Grsqxstw842Laq0tSVEfATCmx7g7Di7NIZuShNfBIWmDSv
LsWkFiE7A7Yj9a2FDGrwcfujeWPbyz00ngEXTxvgA2Cw/XBRz7avdcq8i5pB28izuyR479tfF2y+
3rmbLU4DLXGcanrCyV15v5/u54d+HNnb1bCZjJc3IC+1xUMxycUuDDRQpamkFNy2p7kYNcvKBt5s
hi80GVhXQTmXeAh06NsmTFRSGSirCDAZm2y8f0+4j+Vsa8IhOKnLCOXzeCPNvb2GDzhLZlVlCGT2
yjzRTOA1qEgFKrqpk8SYEbbIQXOFCA1LD8OTHvwsn21oSIDDuonzgoANAe/98oAq3YDzjJZS52fr
Bg/TFni29vSZkqWIOgFXJOD7Toq6LtDltfMK/gLrxRP8Vc4r78Qo8JN3fU7+dp2MDagDeV4/4zjj
A3ZSY6Wth75HwJlp0A9q8NpvfNjicDiGKJTqFenSrH3/3AUIv1/yUdiBHfTuBEwCc828JKnW8RBE
qS0rJK4SpV5/ZkjnlML5GnjPw9YSVat95EX4ug3ECNihBNdesVxCSTMxahVNI+qdB3CjnsFfFr3U
D489qIj/cZKgzNuwQyqUH1sx2QoCMYc0mYKg66aPhjnnJ6rNhyQrvHd+54+yA13S8uCW0e7m5JD4
fk5Ix2hXFhVxt9eprP2KS8+F7DKQcjRwLdl5+6ITfmvFToAGwSZS5B8EwcCx8yFlcGaCbB6nuI6p
voBvapatQP2GqrjH8lUajqeQI+tuml2hgQoE5DKQRfLMYtGo3btvu10/qjGnLY/lBCsmyayzjbS1
0neiImnn1jJ/Go6rD5IdXcFvl6tXOCFpFvoqFx7yySOwbdV7Cj60u1BshczjqifFZeFEK6b3AUoq
uRmvnKZegcnQkj9WoKbNfMotUMdQDSugnu2xzFBkOASoWEQHN/87Fagf4bqGh9aKQ7OxeOVn72L1
athvFuQVW9uDin8SZO8wn0HwKfyp/i4TnmLQK40Lm5GLMT30B8ZL97DmQ+tCYRCD/eRAcipNK+Nk
QRX1nUJsX5Frofijl5roP1quwGnXRpoull+kzxNYyNJjSYcO4I766ZIHK6thrO71FbL6ShYaUX0B
tZ8i5qidzwKoJqdbjxfK4kGKW9qq5OQQ8Dz8Zbo3i4vJftuuvuyX5XaJmFRSCoI/hZPxtoxIY4+d
q8+EiqkSHSYn06BL2ET0R39J2F4uOBNoAEujI3p3eXGi+TjlQ6zPs1WmuEpok+PN8O4hp4AB8fa7
IyZH2aN9L7KNsDJ2/ROtwp71WgdC+Vq7UWLMhftqf6yVj6b3umI/PhhbXYX1vpjRRw8M44OBCXbT
lpEZ9xOwyqD74283pVdTW75oYQUxiv/m8COCbFGNWoCPe4cFSMwb14PF0Tg9v48PXwl6zxWJ+csY
rim2Ao4qmHF3jR3vqa8dDmboqjHrrasxbnkoG+LOG8DNjt9w32XRrCQxveMVj4lL9E4/bD0G56OV
SKrUg21HOmPIuXrYSSacob5vLWyMTwQ83mAsTHx3/gkYbr5qM/m4wp1LijvPE+8Uk6PqYCmnJ2qN
Y/+OhzKOYo5JHpGWfYY6RQg0RQGxS4KlNiWA9E9stFO+pLuPG+81rPHSyfojc4ggP4pOFgV+U1rT
FJSiJRGVnQi1c0I0RqZauWGWNssVyPYOIIh7mkL2byI9AnsrmwgOTZPHPxMvytI4LaE55quXL9C3
3aeEx08RYdmUoCfB0Z8+mqecaQ7k7Du8vZ4kvdEjXmOVVmpwSYqolUbDZp2ej4Mi3/2Tf/VTZRzp
oJY6MpMwVLyAnI35YFZ4x4QFDmpVMNTc7ZOmObr2JpND/wPXTeOfvXpb5vidrPlRdsM1XkXwBAJM
qGeLEX2jfGUqxuNKm30Ww5qMc4K0iJztuBKfqTg8TQGkbe30qWDtUfgkiznVYmWB6pIauftYI5N5
l+affHx1V7dJAl8qlUWhIxTVUG08mke6NWMcEPcJp3sScgE4ZJSSG5fZrq1ZSZ1DG/Msj6SBSbw7
sp2529IOZxCF+i+w1p4/GNX+GhkTNXV1gq3fHRjeaQtr84LF7xMzVbzgTHzDAsV3C/2V0r26Fn+T
B80wsUHjQTkjAeze9s4c5KQW8oJ31jyxuMHaXEHPyCEbLU+a6YskwqXL/WUAIV9WKBAzSi0ojiO0
su5TgG7r+cZOrllb3i2E7bZmGyzI40lwgY09xU3ri2UjlvimZKP1C8wfU9GgdJ0198o4kSbAXZsc
ipPE3jHG8vrwQ2G37f27iqJQrXpJeqB/85ogH1M0zhjbiJyMZIaTRQiVRNCGlb1o89XfNL+zcYY0
geSu+HlI/DMbypJsJuyCiItqmUBGx7EDsFig5daMkzBsokN8l3/h6pFL2xqKXT9pkxvo9o3ymFJA
77poZjYFSi2QO9cCtEyYh3rN9ca/Ycz5hvuYi/7sEtgpHsFd9JqdS3v5VpgZJJy0dWOAFgTyPRR5
j885LlXK0r1n3aJ2mQzHcSViDmGeD87tQczHY2M/c+g9vvnj7quFaWvFnlGH6GguKAAi/vGx3E2H
D6i6Osl9obEOPHH3OBUkSL/1qmlgzFbn00IUMaO6SXdD3YdkKPQY40DG3FkBBAKoMK9bgVE/tlkD
tKtPTW5ShUDpljmy+Z6rdiQz20Nr47WV8yoDjlm/BpHgZ05MyuDlQ5ZU3paIlvoChn443fkWrFpu
BgB1ZEx6NIMCMTHPoIjmm95enJnxNMpxb2Oe5FerjObmZWxiLmMvpBgFcNIs8z37B1x2MP/ji//9
TA9MG062i1QLjPWEpy1Rd/aJgIsEBfyer3rnk9Vay1hKYFjewrRlkBO0z+l2lSqzcjKSAK6muMkE
IuM6Dg+E7BQrQ3DsD5+c7BqGUT7WiElI7JGxQVYdNGQpXa/b6BDfNsLhTB/PTozAaplwOE9eAMxV
8bgVU07uYo88WagO37ISxhO4I+PrMT1yLVYn3MFQE44gOntUMj91/BGueIqfPTRc0L93tFqWhFV6
UzMHFUmPJ6d9diz+CqGXcwVWb9ZENMSmONfebrCBFvqBOSLgR3zXlaofm3QxvupfvgNlNgDHQx8X
7cpAzWRRAqZvL6UeoRFKBKKz4xOfvVjiqC6+MGHArYsxjRTQ48bUA7C/fJgTPoV6PIOkL9AdbbfJ
ummW3fkiZcAyGrF385wYYDWTj8ouUEuAFHCLdstee5qJfPekv3IEbIblTeeX28ZC+uNjVIQz5FbU
ZUwA7rnqEkLUIGuuItD0Nu47pbA5WGs7eRZ78MdabTcYV6bt6H9a4HajHuZ7keUiJy6Isq7acqA2
M7WIzUzVlOTMubNI2hksaYO9eDhuwXXykTm/UbsNdi/WBkoeRc8UnCwNw4uuaAQgLLGRDazgOfdV
00TNuT/nkp2gxp0sJMoqe2UpP+A1ufNpWOOhtI8HW6ACty6GmAoEfs+nxGtFMrSQWTEgbpVHNbv7
vr8WN8nJSK1ugKJg6J3Np4fi9wcI+O1fQjy1mhtFmBp0Lo3SHP4XpozXoRYGNWtXCplsSnSaEY7T
kg+aPQe8LKsGWQ0UiO1TLvnK25BgTGG699mXEmlK5Sko71oHCBtcWwWLfTGxiluKl9faEomMvjf5
hBxOTHlhx5Vl+t6a5PSUD2IL77m+1my9OKq7WFVJLsMy0uoPvKawq12yq16nknMfvxpkYI6yYBpZ
mvLh82dVxfpcHKUoO2YlJlS+KsDdxAVgzx2O/rDqvKXKLxbNX5KQgS6J9SwyIkDTz9L2WMRYC1Xg
a6GzVoby7bGSNrTbvZTAObHJqgFbCwi07rB2052TheJri3yVoiLoSk9e2+M1jWGz7Vk2hgcKlsJn
KAsMj3l7WNqyWzeB3eDBr6K1d+zpZb/Xxuo99tJ0OgKYP1ISwhgZdPuOEcMJOUiya74jxiqss26Q
cG4T+33YjMJoZAFKjW4B2ckc9ETgys/Qn52smnoPMxYu9XX7ZFVQ3Am23jhare1M0LSrDQEV0f/Y
W+CT7grEO9ZiIFQxfK3PgDxVxSTW/nCsVQd1dM9Swvl94zalNR4mPzF/aYe+iB7sd2TSYeV3sBhh
WRtBnL2111aOjBhtrqHQIXzshvFfOlvQdxRflBSLm8HZ1I5vyhxgb2KMCw5P8oKhbsL77r2hV9eC
CAn6K+M/a8coI0I/4xOyjvjv8bU2nx14D8UPtqCzHOTPuqZdlm/uoq9EFWBnPYdTac7QCbLOlzKA
HZmovY21yDktNA9T/1OKKiwhcue0ARgd7JhGNyGCKocPbfDRWxbTLAz/P0JTZThQwsKLKTzQK+td
WVE5uzxyUv7j/gb3v9byCDY8qnquQqaoyqRX0nVOKpFqJJBBceDtbYr1+eaZBE5tuvQv2+u2V+BS
YwVNke2arNDj+9UwrqSQCyqXxQGmbrGUY8rwZtAWeoZ7kiRMTqVsvXTMda32xVPpPAQwACnWYfY1
ToOR9rPIQb/QpM88WB8nfDBecbOm2hao5PDUckSjbf24/1MYPJoNJyTxZQd9rv/9Odv+Wu1xF5oq
hg28hTelKwvOA1uQTTnRWSjO9qoOX4vBdAEnxNEyQxhw7kBtPzOb3Sq010HNpVMpQGLlqVRvnJOw
VB0BFRovbC6GYlFCc9kd/RnAjV8VBfUnFARayj5amDBb4aziF3JuLtyYrgrtPOAda/+T4vRPmF3C
twdx5vRw7gTlZPix+IboLrqDC/Tc8MkuPCIa1Dr1EjLlSucrbWvEWxjNaG+5OsyArzzBG51yBPXi
zIxInU0MR0Z45B2ah4eUDehO36bfHxbd7LkWy+Dmj9UcjOFaUiErhrW6s9M/OYaSIHFSlmlTIOSM
OUQ4a/6tRiTCEEgapJlkSrGlIPlNp1N8+LYemPK8ICPMw8cNNwvs4kT04gGy3UFKDngPnZe8xel+
ENqPtg2i7Aedtet8r8WPAY0DkbvQBsYlibDFiv7EmaldWdgt/w+oh4bPEExZmY+un3ykldn5wAEI
I6dZG9W5lJ4xwNJ29cjFurxgOrKQT4HLNfmDDfMPUZbgnfI8Y/a4gMX2uZquF1tfExydkdWd1AAS
qyBz2YPKE8TASiEXSQWOpjDiDDT3yn/aJg8xrS6nsiOPs1b+6bgqEdzQ3TVhocursN1wo1LPpUgf
T2pNoTVSYDKNmRpetwj8EPGZ9vkE/w7ia/8icg8ABWMfPDCbXZ1v4m9hSnXrz24h3j07SkgcqCJZ
6aBSwCs8gVwfzmCSxU2VmRbyv2bcARr/smGX4yFhvN528XvhXRoiUfKgUmnY640uYncbsrJA6HwN
QLIxJKKtdjcFu0luzUhObslqNY5IvoS+1jAoifpFGoYL6WEjbgq4pfVrHmkjBhflkp1WgLNq8Hjf
jvpJWhLfw+uL4GRATGcSWz/q/ZQhMr/Rwk+vI1PxU9kW+Qv+4XLnbWPMtx3B1PI46XYMLLcAwrB9
pHo2ZyQbnR+58IPeJ0b6PMhBwtewp0p+rEfwGznxcQVi5seb/qgCpY2yDRlYcr73KQ5b3dTSTtZA
m0KWWcFL91b0qgLvpZQeGlluOwJfmIZrn9eyClhjRhrY/bkGiRMuZk+diyCCdQ9Np+k5iniNGclO
Bl302eDw0Hhcp/oyVyzWhN8XX8/E0JGaQEKznY26VfKF2MOBL+D1FXssYmYDUi1iU+Lo4MYmjg9F
AKtVhDctj3wltfasf9NG1mfe3Jkd6FxWRueDomrXy/y/x1tNxkR7RSaiL91HM1PiH5K4cHCyOmHG
FyC5119iVvymFxMkc7rNQgrblk0JNd3TKfsHjrDrPee/Fe5sWNlzamIFUsIeegekNF4sfTH22Zce
0pAxQiEDBU+tH4uyDSdmsA98TztqjP7EUC551KlgCnL5w1OV6QQ0JB481mHG/3tZ3nakqMLsJtf4
xeP9e8gZuo/b9tRA22kEeHQT3mW+bN4IB4A0BXAgbJ+YcC53IPuS3sutI3YfCPPkluzlRCxym4w5
S/0D938fl+tNBTnbXqVCCw19Lzx/s2iqSJdtko0hegFQTjJdvJqmalA5ubBLjYA2y/8q60tIfb/w
txxYB/sNVs9ASQ2bKIwhkz6cKqZx7FqLPdGItcYneoR04Rg2+vj0HAo+ks1G8k9a9ZAUua9OC9Fy
8GKEJbEsNr4a6FeInL50XeyHlBF/pDgeE2DUIc7P78s1klCQHrOzo19E4cgAllmjUG4OzblDxkY+
H6skEAbJLlmAiRg1/zo1dU8ItUtoVUR8HTWNpbxAYO5SJmurSLQ466YzGwsG1dghWkrS8FhpkxJw
eGANVI5meBjc+DD1hoLN5H5uFR4z7iRFp4AI/Itg9KFh4ouQ4Jgq0nGJsoHX07eYExt+Ns1MG9Ni
5ahF+WEeMf8TgdkastLrv5gHIliUqXYHt6StNaabnQPjYiDdqqDGpmPFekRAYl09OvH/EhvGGtbU
ZQBQtXwtnODJ7fVeOOC0woXrlrOZJV+Tl4gBAek1hb7zR9vn6cUBBrEig9nEZlT9Oeg9i6QghpnH
fTMPQzWqaOlrnzFp5dmLgkeWDlcxCM1MXSwsCshkGCP7ZIE4rahU87X1o2L0ypOqPVJJcRLgCmT2
UOMZqLFvsE6yyfAMifIHxzouTf1+gUbC9v36TUop7wdHN/mm2pQ8pgdXZqByCfsl25SrQV6XXOMq
8q9974jRbcWveGoR8uE0IXOGtn/mfYvgD793uYTbyFW4BKUMvUZvsSy9OObPCVpVRdjH3z7ggS9F
lIs3/FPsihjH3H2za6o4auVxzAr64tfWrFki5mL9NlTVeUhaduT+NdW3y4L/LpUV/Ha8+jGSRgDc
YDhbgfWE18PguRH7TTuCUGAbshzLKTuMS/qjiZemcQe6+zM84XXZeVtv1RGJNE5j8a2CJuWmXICZ
eUMLLlCZoBgFa73mf/MOnNNsx/o6aTTOkGsjqH2U0mOLizTEgjhw9nQYRICLftcIoplK597007ZE
SN4aj7kXv6GMj/ZYi3qSeRMraA3aZHWmh+zmRe4ULWrJKXiHkjAu+Nh7EBgpX/OqiXJecoh8Izru
oe5weqbXwkVFBZ2Lp4hHRCRHR3rSL6H209qAw9ykJvm25MmvKswXvlqZe1kIMUHy9GJBoneMcV4V
gnrs5+J5tQmcy+IGPHAnm2M5TJF7Th7A383h91rPDtNN/h+7AbSc+DO+4NPPgVKNzNQ1G0WaXXu5
ReWLeL94tGQs5MQkq78JEp1WnklWUKNmuqESI/3i2j1ndVuUnNHtVJUrh17fyG07P/3SwVrX6mR/
/epNx5y6rQ4kgfoDnhYHSrSKS1t7VkkqzoP7KfiSrOpGvkG68WCgWUzZI6Yk606z6ekatAZ2AzJy
Ns3EoyuU3yFnLPLojnGzbxNKPT/vuDbLicfMVAvtEWDeKkCX7pjfVmnCk9Dz1AldqRZWYjnRbCwY
EwjNoboEqN2XhKQwa7QXhIPLk54dQ50ceuZy1noimBe472P3+wcoP8zgMMNuMBrPtnO5sC7E8WJZ
FJBWj4Fdfbk4awfQuOuP/05dc4GoIrFfxKY5zOzo+fSX25K4tSVgvDo3EocjZf7fggk6MiSRJ3z6
HbIJk4CC43/dtpnj+mVPYZndtr3wtRRpybZ1AZGIj7NZHwHNtZA7c7NaXqyUUysRKLzHB1RM+L7Q
d6OYBNDXiA2Ddly+EqzhgCKdiQPguOnAOQQXAZAGtUm6DXkCttWeGi+vdPNXk+1aH59ODH3niUiW
lPyozC5HfjBYnrxQ40SlZMhlWe/EdlNv2cci7lKv3SSBBfMhkUkVwKYtTq+pnwUeLWzaCj8I27Na
Lu6rIDW54eTgkqxVfJfwgY3EXSyZ9JYZzNmE0ymjN1vXPd8920ZtZ60uVzMnv1rJWtzUZmBEp8U5
ku6i3sn/BncaXSz/ONG7FgmGCr/r2dJjR5maXxULHuA617tgXSTwBSVYzC4feijbn3fUoVYtVc7G
Q4R6Dk7lYX4Oi2+n26X4IN4bcXv4waKvswd2x7XBszWUFz42k7XAYR0Kk6MAKeahpRwf3EkXfsLA
sNElEQ60bKGt30o/sY9jAgTXabMASPJgEHSULSfDcSMSeN7yjlzmMjBz2ykHhVvvDCVGmy+bkVO0
6xYLpEOt/F0TSqA+uh37mO+2CVCdyxe/kGoKlqNFpL8dh5i14QK1jZHJvcH90HSBxSQ+tsANInbq
FeGH1nvLhTactnzuWC9HPdzg7oq6PcX6228+cVEDrWKQF8b7AF+cegOO/PG3uqvOAahnpZsOROeR
JekkjxISMGBZLjAMnB0NBHCTJMGNrz/qRxVnNSnLv+xZpb8kXeG3OQQiD93IdGdiT9nYua+Uvg0c
/JsBkNJ1koW8Jz2JyJ2apYO0MssEayVXwsRojSZoCPCtuDf0CtorcUIpXMYKEgER/IICkMYD8HqY
Go9sFBBKa8mdiZsMCZ06a58p7tPbqJ65fTEt1twjNbLpy8/I1J829qyN/3xVxDjwPbR9Sa6w6+TG
O5hsLJUOmes8nqeeVI80GyGa/leTchZwoRKbG9z+gz2BTffMyO//GbL/5ER7woTdz3nreg706gtx
IfboCxpjHMuuN+l6rnyRlRnjh578sgePFqfPQfvgmGaYLGiKTRJ+BRm5VjrU6yBWYUUuKqRMJLMk
PsQT16L0qzrv0v4NKPBbO05Lc/Tke2XC0g6c5DXQQoGGQYW1+IMdXjf2A3S2IsBTqBwE5rNwzKrn
Tro7bH5EWP1mnigCUurs1rvy17LcTdn++cuLbU4yqtAcHliocgmjg62M91XLmdpGZz388OMyy5yy
UIooElpcuinakVCV4oKsQZJidhJR+9jk6A82kGmnKFy1AS1bZ7p7P4AyxMpMjBouTHcoPQuJr5aI
+knfcibAYKIzzkqcdFQIecx+6tvOuO65rU56HsdzkH7GqC1z8JDwGLHcEBGE30GbVsdemfh+kfAK
Az6EuyOwqDsZTDPcv2RqTfci9h5sTcnw6ThVNxMycneMLGE2l7rRA9v7MW0+9URt/k/To2AeVkDK
UpH71/Pp0YBBjtRqURhZ8BRTp5We19HFF7ouTZlM5mILRkE+PZAKmXmUG81Gg3evyfVnSpyRMxaz
GX5FDKwF4aM4KLK5clzrRAsQeTNuLmRJ9Le7AOg2DErQZ18x+W7omHOXWEsWgiNAJMqPtHS1nHZY
5KSATNdqJ/nBkU3NjJiPgqIeX+ogZ90U9ntrDGXr1GPIT28F/na37QSPlgyVY/W0tiwmaypRcBGt
B8TRaQEFmSIsE7sazdM9zQh/jBAqaNcwTGWJtWhiik7yDpwdAdLyS/AQYCEdSvI0o8zbjokkaw3d
6P6pjJ0DR9NhRNiw2Wvfm73vdoRWz0Hl6PLpCPW4dP9u+qzjjnnZzjyYoeLLbTXvrenG9IKhgyDx
FGEeRz5DKSFwRgWRdzbl98EEbxu6xeNfARX4Sh9/D5bca35KLF3NdiGZsR6UcJwYHZRQqkMSuP8E
Sy+cZyRBQWEsDvcS13FRA/NcFCH69N6EWQIDWXYMZM8ZDJwunZRnLiaovQ7Cqbq7i4up7BGLb7Hf
6FyiRKRTUxdMEXja3nKrKQ46Eq4TzhG8QIH5Cqgqyo64bRFO6aCVm1P76PzuSjMlHwFRPnkqjd+5
pUUN0JQbam+ToiJZtf9F/VajUN7xpkouvdOxbYuwTi1EVZMFoISPqU7PP93zgtRG+bY098FdBR+d
b7tik/YNDqypnEz9k6hLjxo2E50qYaPparNcmsuSSlKdY0wC37Rp+Ftv3H92JvHgWUpk50BVrAAC
RNUycBpn3hVe0bYqH8OzAZhzXNdvICuDsLH3PZEOl+jn6Mt+msBR5xzkAmuAw/2C9Jp6qMz7M1cp
kd+a1/RCyBVR2NMgQWYkTFoULoRP1qi6fX05pb57IzXzjc7W2Th9EiIRbl/+3rSyxlW6hOUXzJDs
QLIF/8qHNHsc1u6rPqQfM5cq3Pc+DGJEerqi3Gz6qGLaID2vbUgMrk4WWMFMDRCjkqu2rnDzXZQ8
nAJTYB8m/5YRBcD25p5jWbXp+kjhNytXFWiOFnT3AxGw356BuHmsdMPsV6JUkMAazF5OxIz8V5gm
Ax9K1E4TbOcf52KKVs1L2om5HlOs3NwWMNCrfLbCQ5YGOYmCgsC58uaM92ehiDkFv5lEyld2b8Y/
yYCdNs65qQdepfIRrTas8nw9IJN5tsyoqKJvqwU9jG9Q+Q5/Nqo8OI9snNdzP2jSZsyNlPXJ6p+l
bLsBtdeCCMFaCkq4WE7baOPsl9f+ewwxtn032ecQv5ntsJSyUz/9LYburQj1JZnD4TOpwTTzFDZH
m8IH8TJTmhUW8nJOKBR1oG6/Nd7qzFKfgjX03MgPvlZwbwwVHKOQUc3SdUfRB1kBHsPMHYYYnBd1
3xG/dlTr8jQ4i/XTm+3WgWMERoKfln6FxYg4JxIock291plXVSZA9b+9R+RkGoWklSHufLxqPFKP
LOFHeG0+2clQ5XMQ3MRC99Oj1lHwnL0qq9RgmGkp6xuGc0VeJT0sdxgyK2StSmhZ8dY1BQQ//fQZ
4mvb55nORw+9BZbxOYP/lKsp9iFdFgqPUFSprMROWnonEhMD2eLovfPilhDFCTmBjlqw2hbMIoZQ
gfzAMpXcARHrdZpSi6zOBB5Z+9twFtWPzjW85xZ95sgG62L4mKmEIqJg2R9CQ+WE2G716xdG+z6+
ZRrWwN1LmRvnNcWku3WxdStZdm4TJVq4uYplMsrITFcXatPgJPZObMO8Hc0chdYvSZgVvABa0ops
VVqtgJm52ExAZlL06a2xuaceAsE6BZSxVsTIlbUsU/af3YRMhJuC16vIZuY484ggC+ASTTaf7IMY
d4r9tp4+p8+N3iqZOuIGwOv2TLRUW7GA55tfxGiIgNT2+dvf1cvVp535xQIo+kANVWP0MrjrbKdw
Ajrli2PLO6cq6+3JTum5HZ80j/kJepHlS52QHpXHLLe8Jq90XTRH7OqkPgkI8bgd24G3fwCNcNYq
NoLaglX7gTGXti6x0sgP6c5LGmBjSNz3ywp4h07UVp3eDvFC4ru53Pzomz1gPAQ7d5g2gt1OTlY/
gpEpUtRG6yOu9PYXrzkD7XGI/y64jR4/pZ/67XYUZgYM7DVp3wL7YCl9y0dQUndS0jL85vuF8vFT
LcSa8Ivw6xSIpkq0Vnq3me38qBQ3tVlSPc88Y0xmyi5qv3hd9csnh7F74L2MXPxSe4iRb1IqJRrf
09GahG99/PKhnPNYcxHEQuAeZOFGNBdG3vfLXmKvBtczYVVwRbStNim3ADb3sJHgDPwLS+18ZwIy
rdGs0Y6kG3BWPB99p7YwvtCsebFo84NjHopyxxBWaIiCk3+rr7MpAGFJ767tCXs6Vs5sGB5ZoyDQ
OeOTXsDWf2ZL2bWnrFFCgYNCuyYFQLFo10fONUu1c8zdgFd0ipA8TpTGIwfp3KlsNKnCDdEYw93E
zsyKWc+VTSb5R5O2ZyoKbsi/iohFqeXzeTq3b/7aFo7Czute0xUHAZCTK2FCXn2xs1X+m9LADoZm
ehRsxQQBtcol46bWysVt+omFr8xI6X5kG6NgATaWDJ+Jd2l49cvBkXnYIAclC1ZTm2wVjenVc/Yc
hH7IZwLWuRnUifHyWOGEgx1DKDL+sqPC8RIjwiLMD6Ln/edVTAeDoKkBtLj7xsrpFmjKIPFUZbf7
lo60Zz24VTg4Z0jl3GIzudQ6/6z4MB9ovvkWLGWcIZP1sqCS5RZCVEZU0p36pj+ZzkY4ShR6RZUL
pOtaFVydykhndmpLtT/sgHQlhxMw2lbD4JgI7RK0wmFYSROuUCRg9b29576bonPJMqK17tqRy6pM
fCPR8tgviu9lKa3qJ3tUx2qT87k/NAsA7A6C0+AQYuI9K0SyCiS4fxoqNwOe09SyVh7JW1FelXsr
Jt8hjRDVkH1Fg7aZI32zH52CMmGYpqy2bH8io6rGKU9Tu3P4HTziebn2uENPyCTDsLGXBicG/TP3
HYJ/IwJ1h9jbXjku3nsMrIUM6PvdVLhspx4QQQkl0AN3auud3Hq7cTebe6H+uVK77g4sH1VcpKeH
lrnGI3xK83p7O5U5Z4f0xPNHckgYPz7AO8Ou6+Vk7P6ZwUs7tb88ZOlgoZRJb6wBzvmv7v50sSup
KqiIsLmPRy9AZrv/6OPSSKf65FNYV5UcCzXc7FaYiouDcu1o7mzkYBKFuZ9lDP1Hwz/nOWkgqfcc
srqKPez23JB3J5vHAS+ecOpkkQEF3bRq2KY7K7xVwAF7E5b0hYOtMzCZjLYogntsdgj2a+wBr/OX
wloNEA3cU7gb1qQ8EI2yCiGOwHGLlAtTI/AXo1cP4vaL1EZDYT3Xof2hAchryFlXV5sK9jmi85NI
WQyN3eOeXsi0jJo1Atv2biEcMwSAnUHp9XEajNV/efZtzl/IKypSEjFt/DYEPSnKfi8bAS9hVsfN
CRS6ow9zjiyv6p+4LefD2KQQRdylje76eNpgxKtuLA7m3Vrh2QGXzVWuxg/0MRuKoN2Pf5yoH9Fs
vfF86bpsO2Jgqg6WpGDrZM5ugVRY+jP/vGHOijPGTRpIEVxcsiUcxVmNoQnkvFUYhmnMbJHFClLf
3ySf6bz3q+u0+eoLRPrdxr5G1kcoepDD2ZorDYNl6bDJ/S+fzuWnL3/Qq+KoW41TZd9pGhwbmLDy
R+X+sCQaE7XVZ+OiL7mFo2Srze1B9Alw6WEsInfy9/ofqGHbJACujwx808mHjnrQJVWL/PKf2Gsp
XyrML+MGDPHfXwHJdrPj1qYT2HurgYwgYDGnVmMzg8XMUWcKKzdo6YMUFPP6pthFS2Uj++SKUK7f
HKDYtVjZGhal0ixZc3RLUPQjdNlUp5b5qq99P4wUfheGSnfRpOfFhAhh0d/l1ryZY1E/kuiT/AoB
rSKKQaFSsl5M6SVjkTAcydu18FYdgCYAvTLpZZV9yWHHbGge0UxuGV0Mp9zHJxnJCecvQXeiSVAT
5nsVydl31L7GovFSnpVLnea7X/yhL5ZmOdDnvYzeA0fIMyrJrWSbIvOiM+Jsq48c+liJ1aSd0JXL
nCCglPb/PwalxDHxxt/OKpEjjTQvnithvHDGRFr4fDn9/1zZxixSRtskhfxr2/A68yftKgwDbFLe
Tr+j5IGCxWpg4daTcxjKla6gZ9BNJZYrAoaNRsSF2LPMP/k+wux5Q++rPkIt0XI3mkfef4GQQs84
UR8RZ/n/uIzXN8E/9Z1wNUBZWVXNh8TvyX9lDG3ipfA9BVoMUae9H1q/6Ga/TKNVqmPmRR4UxkHd
UOZeR1O8WoRGn5faGvzkLR54kUJB5UDt8R7+SJ+T1fzFDvlWDlIEb2fV6hxVB6iS/61yt77tij03
dbzxZvYvqjB+DSQm/KbSnOAQ9RuLKLcCP27ye/hN4ncY8PrIFlTjtSQnCTO7kXNEGqYmqL0aJLxX
kdV6CzMZcKKTHIq7gbAPMgG5/IRQXGfg63UHBnzTbuVHoxGYH8Mlrev1zoqv18teS9s+QGStIBCS
HoUVCjiChjmDvAA+8QNZlHtJfb1nL8X5NpyslkAR79KZgMBET6FHJJsC3A5hm9dwbKBvTk5BOPTL
6QnL3eOu0WaI97fPeJrBg0SFa1C2xWvy/n/VyKnDS7YM+MYmUyzZ+tBwekDJXH2qv+5MBlpEwojn
uafguVyWQ75iSryFmeKCwB1klgi1yQo/MW7uszUNGUMljiTaEZUT4Kl832bezVs8AHk8dfGx8c29
s/ySSYdL1MA6qyJRM8dYSMgcFcOqxrbUdMkKcRIhFSOeq0YWZhcz8aUKA3WJSZ1cB3bSP1/gNDGs
LKI3dAYKNuh/7eLIAAkdyFuSRU8IIrpom4YskX0wKdvYwB8tnvR1HQQrJyGRqxC8LJaX3Um2in7G
1aSf8zSActsiQHDqb1o5+UU8VBPPHT1JZbO9pHLG98xOZ9VcXwxvc3QLZFetYF35KekZI9vJqzxY
QDZH8hIP1W7LJGW58BReMO7r7if278bRg7XYnk9C6PfP7FrvnJLZkwjakbWoaWO54v/uN4DSH8C7
jq95VjjSPBVb09xBTkH+m4aiNwp6YgWX2SLilqbjWfSwxNPa1ufDjP9RonukxQYvZLJu1IxgZR7K
ZgWyOq1s09eA2J9aJn0+7Z969Yq5hxy57QclVB1C8wbqXpcWFFbJMaRzwPYORr0g63UUsG3nw4mr
oUuThDXyzbOoY2Z1STzX5AGIe7Gbcy3nX4KONBK7RNV7vco6OhFI2owQR3lh1TiVAcdfYCHRiVO4
fEQVwc/61YSvU54VkyZ9xEqYbDKNNPcpYCukAy+Xng9O0szxMene/EtezqAvcmBDtBri69AO7CXc
DG+VXvcKerRGoidTbQsT2KhqDFa/RcMUHzM5VOTLnqZP2uOBl1C3YhFn7AoDAIcE1JqaKG6ELy3I
VM6gNbIQ9+3fk48Ii0NyDu4As9MYiJemAQ3n5ZL5FhOltw7Cg3GAOW0jolCCYXzsXd+XLk2mrqfs
PBVhKC7TF1HGaLCbBTUT6rss6p6mVEFrXmE50Rtppx5vZ07Cx9ZX/qpS6OyQOwcUm2DcanV3Yc2A
aYIckVG5wOPFs/5Qj0OVNdJfeJaTHlC143CVsRhIVpLap7md5AQZnyjrwo1F/7GcsPGmC0W+iNui
/WGpeUxXN64tR94HdU5liEmu7j6LDYpKJHzhqaekKmZvmrkaE71OBo/MIjcVsXw8FIJdhVOM9ScR
2WPlxpMFvd9q+20E61oStMLqORsv1Ls5y9b0VNbIAcLdkmq/Hr2ALV4oflobRfK9ewWOjayucGeS
RglAHQnki4lh0ZyARI6XBJEICvuAVfvaBieWBgwjoDVff2SH25in3u0FhK34g1Uqzdnm2evcFIpj
UkWgvfd2UISxthbQZfhGvgmyroCQxsagJV9IeMJEL9nmBjZhwf1j9GMZtlOa90Dt5Oci2Xk5D0f9
GTbnMYskudmoREWZ/15mgLWNFSVIX/yYdwDqOUPNnFoU0cNPvD81HhlFqJhyNsdQUCzZi4vD7ZcO
3wIYv2lnsSjdTjwAhh7UEf7NDZZIBgTiV4P7w8i76byD5SHlTyqH+0opAHQ0XRFGKGwdDIwC2nKO
g62spbtGQclB8kS4gHg/LNsbwAhOd/6AqdcwP23Y6AZH7APxUtUgEBSQc/4kl2qE9N2FSEqp7Vgm
WKWEeE4C6ebcDSgAGWalxjbeM6hja0lGdV46XUvKow1f+nVPw9Ov3paMYbazeIZD4KJOPxUOJr3V
1CPiWAXyKT+4aulFxATm9kcsKwdYIDcE0aQEJih9gOB1kMEMiv1sM5OLlOFfzPDy0r0GIXLZxqXe
SHabVmQzww2W373W7L2VVrLIsSZ1EjSsTuLnRNZI8wOua2+nfp5oGKsZtWIuuVn4nca+HDSrVqwR
QMF7sUVJVr1tGRYN1ial8bu3SLE7LDOwDwu71b6bI16p3ghN68x82iPCLerX18sFM/lDZs2raTEC
CDuq0wM4mdkpVrLOgFe0c3MzPRKiYG5bzwo6ScnuAnQola9J6qJSkBWlAXlYtyliqkkdKTpkNUE9
4MVSFZY/6YCt2Uui4ilfom6WUNIEbYc5IrRmBROouS+JUvM1rtwqU+nsZz0t5Ielj43iexp0dTHV
mkcngmEOOc8acs4h2YBC7BSud9pBeLL0656rb197aMJvq/nSES8pcSgvKzViZzBhcU5cu+jKZSSY
O/1KuJKfnGd6hW6/c7INX9M9I/dtPlGwNLi4z2BTzoRmXdRQWGeJopXnfrRV4lRQz6gv7YS6gZC5
zdHUEuATm59YgEloP2uYID10rQA0PDutys8js9u9EjKWColSiEjsyKJ5HGqhmUSQgYWXOq+Ye9wG
qy8r/h7UV3Oj+wRY93xXvG+ZRlVySyh8stqF4BgE7lpk8pUBrxdw2ooRBaM0Ldya5EUK44m0pUoK
aB3Wv4bTZ3Cazsa2ilPI8c5pTF7TGmR+3pBAZuHWLxemq9QVyVA2KvgK+qlHTZIhjT/eUMlO/eMF
aJZNKyjDTEMD4ZOJv3LixNgyt3KPb94ciT/IeKyNO8br45W19e+Apqqeu7WkQvQD1+8QRDao7fUG
TcTiytrJN3BTH+uJ6rfDPG+DNJ/4mpwnc5nKEzvx35KRruDYwFWsBC2T/kSBGZ4eM8km9Gf4t+3s
pFnWmytcm3f4m5Rqz9VlXxkXkkmelX2P0KYiwswFyJn3umUaDUSTQda/tp0RuqXGpr1jFG3k70Z+
DaeBsZYPbKv7oUIULHEGOwg6FKRU8KZTi8lNU/yNZ2T53amIBzXTjJMBpE6LIIc4NEUt9K7zW/Uz
pFVicQ6rIR9ejdIFD7PEP8Nk47n1zJXusSwPk71YpEvo+l/WfSAuOWNjZ+oE1iTdQtgioXM5L458
7dvtB2epNLKhsb2jBxaIb7djbn5qVjdSE1PIY+5aTsC5TKq2rpYTuydjtAMsP9/vuovKQFPIwsi1
MowRNFM5xsiE+TtWXq/SLVdpfqKa6Rdf0MI/1euq97ZEI8sbKKyHpBpWuVKMU8nhNqIpn8yPbHIP
0OZKzNE6PHb/K/tF/jFPwDS2YVMs7Il+eXhF4OC5Lu6hmpWsrvAqKxbyPeFkcTQrUuvGIbM5hH5T
h769etKynPWs7K3wvJ6bg90cNIQMteoPhl8h+vg66ti6ZijC3sumAzhjKbg47otSe/ZHjgijULgg
TRkcxl/SktS4FJp3BBlspFpaA1BaVFgCcf/mXRsf+Sv6UBqrPGl2W5jROwAuvi9F/uJpXDBvE1/c
+hoFkIXz8OIJVb8JEEOKARx0kNeuK1i/UsKBZmhLNWPzX8MCqUgU6aOH0/QNQuQierDfyRkaac3y
67SNPIzfWemz6W6aXaYCzx1vJMBxGruQ5wkzNuVfNllrLFJjgtKf+1hJttakh6dDCbHMOA077vvJ
PfC0VU/gr5xmUqvu6hB21Qqt6XuXA1es9AD9Po3db+4CS6+ZvWKYtb4cFyoDkkBYq9OKjNKQu7QI
UVRAABA+vyogvDZCEOIVypM0mi7S9r0kNAdUMToaedKyzakb607NH07itv8Ga+2MUWhJhc0nMpRm
e/6BpiPMo8LZldFeBi0Of4zHmsleyWh2eLVVjiahBBhhXErN5sJaQ+AbBgi/GJe3PWHJ8syE5aP9
XwD59tDxrLHGr6aRwznq3vMO9sg9TaeOOkvvfyhL3s8oibYGo63N1HRqnqg1KQH62pvkirumWaFJ
D0bRvAQ7b5tCq5csL7bCBe6IzTLYMI/Gw6wWvwrNfcJ2dxcGJ+tDWhuJdNZJJpG90NdtQPfSy2zj
RWTN9AADkmkZVwkV4/mUhyDNDEbENukWpZJfdDJv05wbQmgyZaMWpDtJWN5ts+jogTgYfnlftcq2
LefVSZRIwCuzH/LUprfRcEHUjYTQEwt8nGHmXPPIP6kMkpV8nBiaEBzgC91TH6EvLzDtERiPw3+h
VjMpgk7Vnh9yo2uHUV6esBYmW9qjEVpxw1HSTYGF7WbxKxEsy2q3oMoM9beV4qmF8SyiXoPnmHvB
rh/SqYhFb+/gZYSGDlLU1BD8y4P7GDXvNrwISfRXjib/kY5dIDhfdUvMm0BjvAU6FPcOG7Wzt3or
cDzqkqoNdyiF/Lgxr+ileMab0tVotaymYhMMfAV4pNNgmW5Dhz0qYlscmvMsXs1HjOyXq4xg9rbO
tGYz+MutBE8aMbwuMQ4V5A11CUexv0Tu8qrR0rJNpZGCgiGGvgn4jtqAmt5Xy+xGOWhhvS8IROuy
obyVNRtkHiORf6yq77EfzsrfnpEFgj4cDAKWgvqFzTJbofc1+3+b/sAvh7aHviY/nbjtvNAUh6e8
HoBME+xP/lfYlwmYqvL5ihtCnsn7dFldKTFu+W1Wj72CN8UdPAVJU4aimsmIe/Ts1IqRLiKTZd2k
E8O2cVYkX+WkAB2lz+A5uEkclwc8Foo+gl25whN8v4fqYPTbLMbIJkbPq7AIOVehlEfy9TaNEi+M
/SbLQQ+U2lbOw0OFWwOveF4rPssS4A/63BFdkztNE+adk8GCrLYd0hm816MLhG2sD2N3QVBSECzk
rNubURw97VoSNPMk0ZkHi2W1kOjlzFBxQmpXaw0H5AkYwVBtplqaEJJle3lDKm+qY19juoUURqWw
/q95T8xC9A9mwCxUocUS4C0cm9osGBAkltpg68aunG1LqS17W7y709unfIyh+S50KzeMxOhaTLPu
foT9QGjQXFMNja+ZaYl8cN0QqY5fCFrbtNzdehRpgqxrI8E8Mcf5bcNH4GRo0AWcWycfV3GftQMb
ovS5VTTSORiCeXjZ8euYCd58kBdOuoF0EsZAHzcwnSOP+qBZFZt1qFt0Dyne2x5s0H8blBB2naBU
ulTlbqYPmMK3Nbrjf12k9kpTAF7VX46sK9GIGwdchu2saTlwxsGRTqpZOcA/hCbwkBY7wEaWByMs
+mX+vEWfE1ehWYlb6m2MhJD+nDgN1V5ZY3G3dq86kBguy6LqbY3IbTRxnqVOkxgZIXHiezdpbomf
a11xG3jo/CuLdiQATmO7I5QgMGJFt2xKmVSzAHzUkW2ReOZCRQkGDy4VSIGdxxAVEDC2Nwj67sSO
6zg1oB34DKt0tezGzcGD/x6hQc6dzGyQUj2Gmk4rge2x8yQu5L/yL8LtxOrkQRO8bKn7dvcjF0FE
mDK7slELhiwsWSxTrCQ100vN22yjS9zOIaCyx57d5CouwfiTJVKQGFJQ0t3Xulz0jgpTNp3KIFit
x7i8YGJyIwyHnsoBPTIt+Zx9uP866MNpy1Dudh2N7XOXk4lG5e6E6+XoOj96wulkfzhe/GPybBQs
YIjlAIJPMcAhZP6v13Ck/D2EQqHRBCDK/TtqN7q4+YRcSIvfbYuzGbLBWbdf4o2hgYDXrzfvH1zV
gdvMnF0ZXqU6RIt1n0ohhqVdwWfHhLhJofipCVTvWnipjkcUzXJ/lZS0SFvGzrf0YoCv/GO3QUgF
BvxDwA2DB9EKuzpbdziL28UDZGRAWFb+piCeE2PFPQLavdk/y1MU17JGgdC/zlkDmciTIXvZFNv6
JsV5DLYptI942WtghAWB9D5I0xkszZWrNpqRpPJaPtWch3iQvKHZlBBmwKSXVZGod98Rr/ZBMXMA
WRuUQYL6NEIIpg/GyCbKr5XBm8DrWptPirn0dq/68/Cg/tsxyxfNwgU+bD+YfNayESk8P9DtuJ9y
rAdR7rEy2kz2Ig8UOFSZkPhJOslOXfMMoNN2jrXDjyC/wOdbAs5DdnTrTRoeX4oy3EwKMG22lBp4
z3vy6GwjZkiwjEoyPRSqy4Ej+4iAqUD/6xJrbKtV9rs0zauF2S4wIOaFf7yZfLfemMbPuXTLNdhx
33Xub2vkXGj1s7M7i1JPdW527+NH47P9/S93fEpmHqwxF069rkiTHjyf791GtW8BNIY3d38GbLdS
81wf9FXtL5UIgMZKpNyy+8Q+ZcZUm7WGH1PI+mh6jU/sPkwSf53Tkq5+cahuJRxRokufGvnJ8SIH
TvH54LC53OmTGrUbu5CFv7leRo3jPRQkzLVmHUuWiler/Dv68AAx8MBB4wWZ3DRREn6Bb6WLiR5a
1I46TUlvzImPRhT6I/rqAWzfDOnKbB6Go61Q+Iwkwo3RAgTBpMK5KPxO1FbO5LSoHGb0Llobg01T
26AkOCz9GjSITtoZcoy9btvzgfHkxDO+YfNlx4R+aYmHO74eKdEkjdTSNfQ99yMO0xKHzU+wV2w9
hhB5iyz2OpOIDl/8S1/jVdXRvP5DySefZ5ppisD/Ki9h92jYNwzYyfBXOtg0tkSAZbyknaWAd4hD
q11FbH1x0IFySq/zsocuiPW8J4ZkGj9s9BCDm70Jjs45kW46hlRDlz70bM0wLzAZSkGxdX4mQB9p
NHOqMjyNObmytKola+FYl5B9AO56kaSE/j6LnJh+4LqEC2+KuC456RpWh8k/FbBc6RSRS0r1MjPz
Nz+v0MhhG0ojQfis1hdNdcKzgW53PYneddo5ZNb9rDD/HUqzn6Omi+LZHzNOHUQBwHUbHWtIzGsY
ah5YXU5bNIHk8IQUK6IVzUp6n9c8wlho2MzMixE4Rf4BTrJluK3pv0BeXxCMy2grZRLJcGOefVH0
UfL4PHDZ7Xc1QWnMi8njOphOJEFfujnB9QxzKBBG7ZJStGO9aIc5by0jezbSt2NgHwr5ScgIslhY
1Fgs48WNzkHjAOVo9CEp5bKvQJ6sN0vqvfp1QGMYpAPPuDvxS8SIUa2N7mxcBFLfreY6rtvwyAWs
GNaP9blsSnqbjd2HHBY8tfhgBOVtLHFauwIN57ISI2l8NEVczp79sZuaMLNHPh9tN+l3qSOJAKdB
D9d9GEnFRl7Ci4Y1o4fHR/srjx0dth/wP+dP+S+4ChfNpn2BaWw0Ox2bvVstgq1PVs66Squk8edZ
uT7xjv6JYf6Q2s2hsXdVc4PSavTR1OJpIpcsuJ5XzkDBLyE+sr406mmAuJf6Hjz1Pcqhfkzm+bL5
cG1nagGUgOVdeNblULdNx04V7fzV8e5x1UBVwJWd2dj/XVUm6Wvg+eU1owy+HYf7Y7KGvBGzO8EU
qsOgd0EbAp8YyJQdb3OylOldVfC0olAmISdK0289440mTJVji3Qz4tNRtgeR05XmrLOuOKVy3Wkn
y1zvV6/bCHefBMLNyWv9TCWokyfF4C4TsPy8EXWtc08liY+qk02F+8Fqxb0joRZf4PjhJFmureOJ
vc6h5tA4Dzc1dnakRA1gLvct03wrdpxWsHXskiH6xrTVxbWOIABDl2OkU2bSXi2QblokRijREubL
4XG8puR2zg2T8QG3I2C3/UefW1N03jiZHtNgoECdy7IUJ20GAv1SQLiLAy3MzglSGOw0omWouuY6
fAkUIhkg2UsB+smVzW3M2PdHkDTOEeOLfiyG1SS/qOpKUVCUmin46l3mkAXFHgiD0rWe1uiIYJqs
kBOlBf6pcZw1ZK17YiR+DXJ4jYBPgBnCOItnDuCMr2xgqs0ItQBjMVHn+F1DuUpcZKwDOG3RPmZ+
PDdNvrRRluwraX9bF6Er+KR6URwTzHhGJOQzkWv41Mjjwc4U3I1f6kdfNMuQ3gMjC7kDTOSmZh6n
9+V7yWKAAjb9VgDm6MAclklBAHVu79GVlxrctPKRVSsPkqI0VG1j2ag34noLHULjY0Fn2TUI9uap
cLR3ilg2zX248XHC3LrRQk0GQnM7jsUrq+o2LJrHM2Zf89O/qLJrIxfWo9ADlTo9wzpHnmgttk7x
Ns8Wd/t7isAWIx1TI3hJlFA0hThfbBUCRuozkdXYOO9C8Xs57tUdU7fKil+jdrXOviaABDjIzP4f
aAvT4OIO5ahc1oxNoxgPeR1rCdfi9Db5VFsTKSXoYIGJeFVAKtUNjQmRfk733F/7FvJo4n3zpgjF
2CB9jGRl8bPKDe47ffOCgDSRRSV5l3VEvc6hk0W+bbrzDHoP+UWvZVp4ismWxJyuu2wkzJZA8550
0IRMAA3p3e7xSXSdR/8iWNn4V7HcA8eFdJNRr2n614adgBhhDspmaH/bmbkVPDbJDNKmq8Kb7Be9
M/RGuAYCXCaKD2rmqv8hZkKKqQ6B7wgylmNPoh/mSrViJLCXLTkaEd9/RmLvprlqJUU1LgzpVR9m
Z814SvKX8eC226gA2h47lrTz30zHE8+7MIq2jrgJfuZDQerX5fr2U17RSr5RZ+ZNY82JVLzcTY6Z
u0MX7hYzI+qEWS1+rdcu4RJ4ag6e2To7be+WlbTpQVJJ3Ihy0/ZdJHxJ24nAp9N2eqc6uEWKNv1u
WamyFfLQSqDnCrvU3nYPjrrbPagb6c75K4WCsDUHsxyxBjIrqAIeuq4FjmPPLELMhtdu/9cZcRwm
78+6vwtP2qvtSNjotNphrc28v+SHQx9pFFG9oVxhbw80TZiCzH6fyEA8r9LisrxIT+w7SiYDH+7k
VTnzsfenyCFqpmIL+eNomiK1ZADR8Tc4QSaIkIe/v6ZVKDjVMjk3z2hY8LMPjwUSCeX3LH4bKI98
25ItNJdHhfObbhVtNG+lmN8W8y4TcZs0DnYd3guojD9wuYDUoInVUivj8CKVhi9DO9bbCDDh22Ad
ixr0KgmoProU6z6Y2k3PhxV6VtnC0W/MF/kbfQS5CFK0awnRMdtWuOxm9TjrkZVBUEgPw8IZH9a5
H0sPF2G1TKjAVT3FZpn/HuG5GwfMTXtonMwiDaU8QYsDDNDPyXfQ8rAQ1n6w15fpX9fDD0lhSKtb
yzYnsjSk+pqdKks1jRpSdQ2cyzHBKSlroBN2cz6kHWSYkPBZxkYE1aEIzNbvn7TUd21byC4zljzs
BeYryEmKI/YMZKaAhlB/3jvOjFDqRNUgS7i4x/8N4k6gaiO5QaPEgH3ZFyTaDocA5a3fmer3VZex
LCpXQsJcmSNxsDUHNwX85zheC4U9dpXYMtKssfhALYrtQI4xSTcg85uAkPcUncmJe0Y2uLyJPPkz
NZnQSAgDa/drxY5Bwne3wI+/YLE3vo5h34VZA3zQAzt10xtWYyKyIdb/NEajbi8Bqcv/93ymffga
65auWnAyVeJlAZ9K0QLibpCldhlwM6vIqD8h/znwW61Zt0Z5WTp8La6R0D726weeiE2kOrrnQhM3
YnbK7H06jBI1E9lVMyKlLhHC3PqHQK9/HV2YP4UvfZkzYYfNaksdMPm3nQ0/pk+Mk6kZE3PR9Xc3
WPKzffreHPggIzmp/gAvp1rxLLBJYHGJKFB/XcBRvlQkxC0SYHbKPLgNoMmPrssfe1aTgVgziK57
k4tY5xaUBESLlIwOPHJ6PRkLJSXu31DadicKeC6VQo+Omn+zdmF0881E6fgN60Ni77rn0Iuqlb1h
tikr8BtUj/qvr9zuejy18pls7JMFXwUItS+AIxEL2+p1YTU53wUf35SOi7wfiwvs4E1D/hz44Nz5
9c00fAhxvRSZGEMV0Qv3Y5PgEF9dD06jOLpVPlvKzjQv5+q4pxZAZYnUopuPjGnjaEIp2gMVGCCb
ZKcvGtcSGgW+yNc47NWWfNFRHQXe93ZEExEJEL43dAj/AV49q7wYU1796xGJkP+U080zPjM2qLSo
YXFVsGLCvwFPVbln4JxuJBlYChqzPOnIcJCL7u8kRFTalAAdVm5IpUSz+VjarK9o/FE9L9lEfnKA
A0Euyj3bC/mH7Z0UBb8+lB7JQ/qrLVdPbZTYVXxSzxT6MLIEq8sY6ebqo51NHlzadkNii7oqq7pQ
KA7do0O+EjVlD5sKR9s2T1SDzmmtQdC/VOmgxUxeWsHT0jJbHYfEjJedlCBt8Frr4dvwhjKSexNA
FqjRLH3gXdxcgouCPpSVrOX4RnbOwro9RSR1goM1b3MzPdYxL481pDd17HUOx30pVLJx3/FCrXfo
S97FGe8L4jBVfvohXfz/+6pnLwJ0WQBRsgrzuFXiv0teWrAy0C6XbOwjvrvv3VmqEKOWqFKBBSv8
kJBv7M6Coi7vMaRdRKvwYPp57zeG6rBVyKVgKEtpdyHT3iEpM4HEqSn0XbIS6a0UfF41qDNHFA5v
J7zXW+luBcElxUxRR+ZkNZXNhoxyAIUoibsQSDWy2W3HWy0Aom2SIXZYedW3oK43dMblKT1oX1K7
/yjF8Xr+94Own9hAsfkFXkTkgYPdP31dAOVvvTVQ6IK+4gNJG0oQFyiw/oyc0TXGOSohS5FGJ8dp
lPd5TgKZ081+P5c/gl2ca9vHQn/+rViI5WvEXRzDAPpTHvNdG0en7YIHv7IFcWL+svRaluT+Zg6s
wVLPStJqjUbKUFKgGHxj6JbVn4iUBaryAV+UBTStIIjSoX7EkMAbXZ5IdQ5H/YexZdVhLhfdLSpr
Mxod37qpzsfmci0kYJuqP7B0f9C/RwZEYUanxxalyKHPD8ZvOHLSB240iuiGHQv3W7/3AZnpf3S1
fSRLSKdQB6NEUnKvK0Mo3YaY7FXJ7FL9MQnX/7lCiaTbX0C+0AZmpi16n5JqAWpddiq4CPeBvb3m
0B8o9609ReZFy9Cdoktv3dbu45ZS+DiH/fciIV4FgKvMQ+yQWBj0uJbw/HaavH7y3gergWLuxPsZ
F64/TSdv6QGHQlEAoxLWL+QWPhhXjz7+LIH+qN3XIS0H7JN+JWtCdb7K9N0+t2vmjq7fT9Hhdgoz
w544/68Y10XcZZUFPCjQojKVVMMDbNDHyFOGUKf/8dTf/642G78WeuVDvv4B65qDXSfa+SxDk7I4
G0ECjuZcYuJsx6NOkE3NKL6qm501y7VY3l74xNh+Gc2blXmBEXPzedA6RHVWadK/FmxFDv74ueI6
5IjMkQZJF68t8a25NPHUHXCdyGNKZgwLWPHAuC/dn0kfViWUiDB71OI5bOvVsYzDl2SaLD32g/Fi
8W8xNDhIBLStYOY8fmN6vvLIzHnT+RXfUh+tz0KGAsdl4GB3KqcfW5m4YQjVXtp8+i6sxEPEDPN8
D/pe0kCUCmUPaaTOvl01457lxB1Vul5/vebkFweujhIY93vx8tCh9lHfxSWQklasMCrKHPAn03lt
7GpuHlINHB6sBb24m8alGbNKMtxLTClHbYCXIIMhJfz7miP6MiOjPvXV22IQJO+PjUTEwX168xsk
2sLvFKXCghCs4svaajO9EUNlMXNoCLDy5Tdi/2wkAtGJHw56g2VRUBnLwLFwVU7YEJgbODVbrfDy
pDs2YPIDFzk7+2V1cd3T/flEUphtgjKfUDit+PlINBb1aWPKt1Wq2Pcb3s9Z4/Ln8Yjq1y9JCwcn
E/TRc//+cp96Cfz4v2KKZ0b5MIoDTqeecmP64mSnJA9nJjjGk3dMcbM/dkC/CcxXOa5unD8jmrEi
hBnsxK6Bg8mDM/V8yVI5B3owcuWcJflW1A7NaBTnXbXesZ0+JeIrGoh+jB7wsJWMM/YJNzMl5f6w
1IxbcynFgluRjhuLYTvKmRIM6mJ+zWg8V4d3h72p/S6dWJR3rrM5pEvUjy+bSpt3ZtKOJk0zZtKz
qPH5LHWnLso171r+nP0kUytRSSQnZJ9KGFQGsPQHk5fwmCPbGLWATZ9CNXtCwMUqiIhdIVcxPlVX
WosDm2FWVG8FciIBI7NmDC28iYYFurkbeUS0eT0oZDfELrCfG8YRvrPFFc6Gj5KafDSO/jwtKCXv
0VMcEDctmonOzwZs4S2WAAJrxnjw8VnD+/CBQFeUMd/9YBKOV2PW6vQijVTii8Rwenmy/kEuYBJv
yJHRbDT4D+rW6xu58nDfHWVCUNWzqfOprAZQVvnST2/ZZ96o2BurD4azOrvFs4oZ8aChV9vnFdmC
qqPki/CPmElvrgeMQIFR2pDUntg86iz7fXmxZEtm8irSRXH5rgCkLldN9lhP9MSd8ZkkcKL7+az0
ZVRl0dr/lNM3g5umxU76M3cZV7OW/sPwv8Nc71Z10gs3JI4IaXv9udXNmi5BKj1+CEkwvcMftI1G
i64HqtLwfkDeGarWvhF00sZStF2VN5AlrvJsPyknAGkz3wAvAzS/+pjATFvvrDM4b+SKbZDi0ya5
YHcVV1NFLmUEXnsEM8Rab28mUJckTCdBYoy5XgCzkW98gzMq+lBG6E2p22JAt+apCmrX1WcBzQXE
52SVtXC5VUBQnt8qcDegPWcs0pBRanwv7VqDrbxKG0JEnby+T6Dy8MVf9fNT0zZCEM2tQcXfbzDe
QSX0z5q1XaK2/E2GNxH6WuLMxklQ5SSoNZnr8PBEKJPsWMNbJ6W1+ZfAeoDJEeCxdvPPf1br2hM/
bvrnodSIPROabjwA+oAc0vsX0IPU//LxIfwp101/uUvBkjnr+wa/vMWQWxZIJes8FhW96pFOpLHb
Lt6+ooCkX+gMz/ORRAA6/CIxYAzHFxdxnS+ml0m6kctdMQNNub+281XYioIRjIR4Ue/e0Dgo+VO1
aZiRMn65FE321ePgL77W28aoR343SZSXnapTo3u3iPq8BnWe3sfLrajZWZBorEKolKGB/lE+Ki+E
WVSLycdpPlmLZ1Jv4VBcwjUjvW3K3vLTATi3s3dluTppvrNrKYy1awyWCNiJXUBqHHR9k/1PzW/5
lEkAUs3JKa1bTbWAo/iKvYHjwVyZbnH1jEqtik+oyTH2xCtG7c1TSYSRXcUci9r+xz/4vzOHvtl2
KKIVwfKdCR1uZDr84ptVVDp75M0is4xkZLCtw4Y7yC4xzSXJLsLbX/7SZAYOhKh4sfUmDZ8H0EfE
ZSuFWVJzCABHbnW41l084YLnXF1ro9K6ulDjUTkEiQhHpJuynt8Ua2+5/G3fOoZmfCFhUSjL6pC8
hmE1M/zR8hTIlYOEZYjeF/trWhEG4DImrfswTkhDaw2EZQijm0LaNsBJPitDZ0Zze7CMCQVTDeos
uMyJGx4A5XNjADt104qViqMGeFd9Y5DZTCLZwyzj+cE8mC6TObb4DSIl8zzJTOtGcAPeOzbV3tdD
f4wn140SkbH44X3XhGTTAncvsZAMR2+qCG2ipHMZ9Y7pTqCM/c0F8k/JXpFFjOY5+YdexLJ065D7
cfjl4ml4ajRSBspN1kAKBb529NNRshnPoykc+rZPEKVy/Zx1+vKdzcUobBpyVq0mk/G8taktlzID
1Zbhr5lQ6FBGgRA6ATg+iORpUVXjfK8tomCuiF5VvqgiLegzgX4gaGVnW4iuiNbk51AodpGG/T/z
fUWk6tJffrrt/PnmcUgJGCzX2yjaSt4E406NrWubw8idMeGgiKCXV0NBMf8we5qCjCs7q1p8KXHX
9ZpZBkU6lV1Ui9SlQuCZjksU6+A0HWjQpNMJuzPd5ndstHfr8RpTnJzQzjRw+/IyTp+nfpOu81xf
im1J1Wn6NRwMk+W3jeKelsokEzG7lVhqEdso4XwaSfitJjfb3eSxRRVn1vI+KQgKefzoThy23wel
G5FbcPuwTFHSS6rZdKPeokSD3fGRiegxfKctA4hmjCvOUgR784U4p9aBZClv8CN8TApgc9bBVA+H
PVrSxU7lz8Nhde3evjVkgaed7qqJfBP+mFHWYcLJiB/JHlx2xYsTvXhts6dIlqdbxg8SJDku9Paz
TYTDJS2rY+NLMhCXHff4cPKkUgmmY7v68RMj569GyjvemzNatrWtloUcyMwSQmNkB3i5EFN2xDSB
SHvHSiu8VvcRtm768KelDbyPR+PclrpSx672b4V+ePsfSw+eqSXYzyZdoUHQnrTL/JloyQSamsMB
E2CsO1ARlBSXbqSQaDJ8x+fD5M4TPsKk/YbUQL01vFoYDZYRmj9hBmm3HAnQ6QsTTmW5cwZ0poA5
wkeZwTKibDCrKpe/69kieZSl0BqfwQOnUZgXwwI5w11eXXMnNun+GQcwCt7AGJgzKbT9ToEIjGlZ
fX0GY/m83w5hh02HqwcJ+3SlmOJfz2txss0dDuLH41VaAmahX1fZNhEYzB+UbC9lXU0QhPxC1/S0
+4QfqFr7yTYuYqz7bj7iq5dEmCQlv5Pl/axVNOG3rkQ9Bfy0Gpkr4kFoCq5EZM5FXXrx1UmvaHjf
08YlAIEUcGkn8yRrHnHr/YLt96b8H5Gbb8aTCYjLNJ8ZPC6Wg18AuVIyqCuM7mQ8kPJUPQbCu3bf
ZuWFbqWup6ZT1OKhmO7/XUQrIUvXe+R72S7AlyN0FRyZIYB9rME6IajKTlstOTzOwZTEEf94/MI9
RrvBR7BfeNRQsVlDWOfYJJ/f+Guun91zbBmqqYarXOqwrCjMNw2XqIpoddwr8ItZtiP1dCNWP+n5
o6uMHuBL4jcDSPR/L66oISBjdBFngCsdtFAmgnEpTch1l1pqe5ErC+pk/EykEUbkY63bDyp0P6nW
P0etsv6uUUUCjKwNhx7uOBf2dymnxJkSKdWHom8AtR/QH+eAWxy2FbeJ+mbffSjJ3JiQQ1Frkysu
53bJ2SWlFqgl5N6/jUa432JtxbN27HXnVgg8FHHUQC9zbmQzYTW8IKszb5uAkNFeQjR5Lvi3qHci
E8WhidmvAKytY7eHEQHzC0ZZB72raQJelCLVoDwfPU664/qD3dxd0glhPjNMlKBFw5HB158OnhvY
sWMxgEK3ejPBOetw0Dn7Edh+mhiwdJvvdIT2K7NJJ5lmp0o8XpjN9VNcoxkLE9LySS4K3y2RHkYV
aaW3oNd/dACf31Mm7KI/AUgPog3ZTXqU8Z+8hC3xnn6hVSleSmOJZbhmDJu2RvlrUiONIaXWLewh
4V7ML5QohePOvhRr71JVsT0Xy6gBSRuuvETsUOkBWII3cXC3VrHNXOt9mFADO7X/3ZGRJOBznN+T
hdG/zs0JcG9QnusqC241SdmecrMURVkXYYAjOe83ckTQFgFF/heUKYrUzdZNeV21Z0PmHF1+4Ii8
iCWJh9IqAFDIPGR5h+v6HxFMY9bKQp/sFdxypxULomRIaCj97fVVxf06uKhIbwfzFz2S4h9UJC5g
cSHomDCwe8oOFBPBRc1cyGFcUg5O1bS5QqOEK9WcnYXb7ZOL7oYkfr6VQIqT19gy5qhTgMjAzBK3
RyjmVO4sBq301DdlBAp2Bu1g0ACwvkCXSHumXQ/igeezvhYcC8K4gkdunCprKoNTbsIH57YAZkGa
B4aeZtyrgSwyi4w/+Rd/FLpReIwQoQojebiUOSTWrE0LbM4O2MXxGLroN28qB6Z4SFCiHIMDyPvk
RZyIB2keOMN1kUEVH609iumP1j9V3lqLWuhhQTTssSpD38Ism8DJ0Ps6wDvSrUeleF7WrjSk/Lwo
G/cD7t8IWALwLwURs7k8UJpR2jovV7NJl3KDgexoToa8TAR1InJ3A10qmsfsjJCtKb8hNdV0NGXc
ybtemO890ukRaIPV4tLbx8Rj90wThym5FYCaLzSU/QC4sYfjmXdRg8u7kxwz3USGTfPZb8jYm13F
gyRI5md32Hi+VBs6ZBCcF7OWoQG8/e8MD4qzwCLxCQBPfQ4WR32eHjiUgEFAJX/Gy1kRD5BngYLa
7Jh5R3AyGCYDFQAc2NlErDCQ5u5E7XHHzObHeY/Sy6TatKtYNHF1mSZHSkw2AH0Rp9Q6PTIdkKJi
R8t389jwvPIgG4NUSVdtYOvI4N8R1TwGZIkOFNjH1Y2Tdu2vNsW0g8MklK5Ll6Lqx+guW7Snp6xT
/SEEjzirhENhBS5JuGfHVau85BjgitHgPwDrHukeJ3Ewj5bagxkSJEKjZ+3iXM36cbsZkNs/tEou
LNd1s6r+Vuei1Sa3JcNaM+HkWKZmb6r8YNL5rfaKK9KnIRzjV7LnH6Qt38fKWhXi0XuaDFFMd+mT
89pxDeKb802V2p0OsuutSuzQjQeP1Ry2dJXeljWqAxu6x/6vRLgeK5/p1LNiEOuH4lKbfcUzhITY
aOvDff25Z309jXbjD1UTV7gkMaEviGVMr1/4Pn+7VRxrakmo8udTvr3Ub31O2Tn/CWVj4hVLAoWa
Z8atdIcSYlrWlESeqaynmfRIpXqa1zEq5UlBPsyYMTPPWBBC0h8WC9ZslWQJT69NX0c7YezwrChk
QuumS4TaAo9J466cWSmEHoRQ31zJKUsIr0y/t3TIQWaOI29nMl2apfD5ODQNu3pAchJrYf2uwIKr
5GNZTZCZHxRpI5qTu3SvP0I4sGm1bg6bkYVuFvCv3kT8uclH4e6u8Q6A7GT8QKg1RfWswCX90YcV
ltiFvfD8W7hhEtnahXFt7S6Itr3za5I0MNFdXaoqqXz+KBiMWpGoQSv6jAklKLaMBCio0PoiK0dv
HmmsHSz+V4XnV1dsU2MxDOoB0jkNT7xDF5vz+fcRBAMVE+ZlszAkAlDTBtN+Um2yhuVbf9MVkrCj
DIyCjS+wDyUkGoBUGvWAkTYQ1fJTGaOnUcC7wdZLqyPBA0FpY6amzucxvhK4Smrv3BM4cgi1nF20
5M3PGAUgi8wzlzZlsDghU6kLOkTdsdyr2ghWqMp7IXtosEEcoJIWqyscW9WiKwDOCac/R6cu8j/J
ko0equq7jTqOq7NAJbiAUN6+FMsdT5Owc329ApLQ1RPuEEZIrnoZ8PMpBnsolsFaugdK3Gq/6t9q
MbBg8AnWzfndxTv/M0VJ3vTaTRRcJDm0znZwIqbmJPaBHq7Ed7OjHiG1a8kyW+MLZzvmzpjZpH0f
fugqMKl6YxcppscM+bwShKK7KL4aNM8V/q8FtE8GYhsOM6J1KmlDkQqBnElRRsKbU+Lc813ChIWA
wNyM3Y59jL63misd34y8+SuJlzGEmnY6NvwyLU/J7vNZiwQR8zw5dHywarnz/xHGLSGoaqxNZnXj
7GAHze7rWFak1ChHguPu0tGaqszYSAUZ6JMctxWmNq7qs3q8UNQGetqf9OZILNilQNy4LQTlyoCR
xrPtiGJyde/XsNg3fzEdRmizzmhyWVO23TRHeEldUmwHwfRebgISpr0rjjwJY26jMO5HkXeEwzCH
uXZ4h7w5fEIfDl2t53WumLvLk4tMdEFQdoZKGmO76NiMJaQgEJC6AFsfVzFZuMiXXYX8cgqQFHM/
3UcAe4iTiasd+YgjHB/jJ7WRLTiv3UppG/prCt4XaUUHoess5xu7UtVZylQ9bQRv7fxaKNk0yS8v
YLL6EWEy0WNgxBnfMjlwuh8FOXEtzY7x1b0gNGW71N4Do/fPTeaezjbX/230x1l6ZW00tniReC8Z
ACaimPUBiEkUiU5t9c+j2THzzvAkdMXYEmnD6ttbJJkUaqKf0O7GhVGwVZETwENGaSHuMCVsBntG
0mhxFIEE49WDB1tE8GooqYO8Lg/4TB1vpULBPd6N11Cl4c81VmTkS8azlbz+t12AuP9tiB99K5RU
0FEDLRea5s/o51W5v3c/nHh6pKF2Wmuumw1w9goyP68nb46FlTESJBDiv2zvYtMfZvIlASdaKMdM
A7N0xWS8gGy6lIv3zYqOMfMG59tgvkG9iz2pOKiYcjbqf9gn8zjqTZ+mGwEyGtS8L+Jybg6gPxg6
cbCYDUcETGX08RTVfbsc6/tZBnYVe3RnZgxeHBwnKRgjFI+0fY4/3BXtuwmjxe0RzxJQDmOUAAKh
JuodxjjOqTJcbwDe+68j4Zd5wJJqIqVZS8N9bCg3QFECx0kgDUx/YsaGCo3TTt8C3J5vtW3gCf2S
HMY4cKuR9yESlCybF3IzufZwWx3EsgzJJTsIyB7k+mLSWKEzXVysC535dOllGiyXPgzYP5baM/2S
cAVOLtWVljoPlPRzkk1Fib8IqHRwJLya4LOeVQr8GxP2JH19oUxrZlk1joGNbjZw55SINk/5NabZ
QeWjcIZdi1vHvEi2sZEVk1YlMNiMUCEBaOwEvlsS0ByAbERH29i6e+Oc6ykMupfwBOgZKCVxSA/K
tbGDCc5DWCks3Q97BurJhuiVnOXsfZ2SahsA0LREwE6QQ1J3W+nzUyfg+E1brIg3Lvzzt9BkcxYS
KrHRHQst9ISN5DroJ7XZlqeVq0I74+OKomZqgIyN5iNeWipTZuVQ4B5e9NPWBG5rtFNKcKA44AKo
0UwG4RgIidjs/LiWmKcmYOmFS5gd+Q6L4qyleueoDkCU3JkvWQxx8Ea/6U+33FtmJx2KgEtuAfky
RaKcA6BYEOBuOQOVTCOSSdmAjYujNQD+puKeX7p55LMfDTYsvpUWZ8lS0tPrpoudwk5S4kY//DN/
YS24QHzSHFUS2T9OQ8kHTEE20ozlOs/O4enYQHJ5sX87nEXLdO9D7LT2TtPl+Znh5mA6nG5aQ3g9
oTJb3+6YqZo1hbXrhLoArO4F2le25jeFYR5I2/ALZOw2DHNLia1Gb+gWgZNFNoMqKENqc438qslC
Lsaz2Vscy72+WCjgKraN22ocpqBJiBZteon6fVl3ydsfFPwQOYtehWAqBNAqHdDO1+bk+6oeIa/G
kbBR7RvgAPVU5zw9H0tXDBHtF1+Ab2K4jgxjDgkTh0rHoa/pNMUkwBba6tPlmtn0yEYIinbYS0Dw
/lGeI2QfhheLvXZG1BMeNDO/kahYO9gftnUHy3FPTewphcdIwBjOJOaah2cLhFcfQobtTFiqWuQC
TMgeI75h/xOPfGnNc2EqVZ1WuqPV4My0d4IAoDC5Fgnez4Hnys3y3G8lgCQwZlqvQnqFvSpHsVEs
WAEpqmCl7uJXvMlWae8cmM3LO3FZqa0WiB4Eb5gOFPfo7XKRcKxpI9XCkWEggInU5gY80WVZsBpC
Wv3tasdd6hH/dNhFBxaI63fqprMB5V3oov1LliJF7vTdiOyG/ARSeSSbGkIETUk1Mr4+RFK0FJ3Z
8TyTKSpSPUVpnqT716W3UShRp9GdOa74GgZOjFIB8eOrucZPhYKMktKUYK4/CWNFCC++t2Uvywm9
CIEPe1Qv9jDsCYAeLOXhoz7B8D6DQ7gDisbQ26h7frBYdZiVn7VaZfsK1BPk+TXizR5reMxyQbwP
a8FKjAmwbjFY/nFJd85aKsVZhAJRK3mEWA+80XQLJ2hEAvvXPs7Lj16AXhS8Q6PAFVabiYG8kDza
UIbwfN28sNoFzE/m1aPBxvEqxeu+5vdm4IKMiVBv3euTBulFVF5Q+A/BVPIHrn6NvRN0AVltuKoh
RHUDj/669VzYO+uKbSBOvcRiV85/PFQPnhgVAMn6eoaYMuIecyIWBT3Zg6H7JLY5sH2vqB3QSptD
v8TtqwJ947aTx3lphwW0wVO6lIy6g8pXRpuIYDw2Bbiq4mIG2xpffAuhe15MFEVq817ketUNGnAi
viJyxM9bbKi5eG1tBd2OY2eXP7+9uk2N/YT5cJRpbQHWxT2AQPgNa1+rJXYdIv+fh/3xj+tSmZtq
++XzvnYyaTTM6Z+7UOOMCv/x14wUuAK9YARt8gQ2qT1FbBGWgZeGqiQnVrlBRQ19j6q6YcxFjUc5
pOxK5PGJsSiv4AA9pgobSdjuRpRW4fK1pe+oycSy2sFN9abogu1rlz59Y5ACg+/QbbBNPBWwzZKc
N+pBXU8IRrRRkgnzXu3DWgfBdcwGBOUkqd2XYkxUedFR3wJ6/QRQCfah0LzTdWNQccYJZCV7ZNhd
PUOLfESWqJxDvsPAZX2jmfSYQs0XcNdd7H4XFDgHkZXDrhb1g5/aJbN/6NhyfVDwvkG94wAHl1ZB
MqUjXjQK7C4XuREjFdGaa6/Uk0UWL1TLMWYK2pqm7Lo5WtW8LcbpBzeTBmjqPyT030nogZbVotY+
jLW6106OQTjt5QwWvZP8nMCNMpDUqpFA9//2dt01Z5MxX1R58AymrkYF73jnWiRPUTJxSlg/FYWq
NmCcluPTM6YmkvatYCxlv6d6JKsNSXH9cSsF7QIoLCO5A+sb+QQUVbELOb/FAc+/yxcyCx+64q1/
8DglVwY7YEuLLTq2AzSrEbeRsCz/POSqrf6WRQHEJ69f986jfzbkMOrLCqk+d/0VWrMFrlKTmZNG
I780jsWcawLXwXC7BKZJf6XwML2IZBU8p7qFWv+T69IeKzJO62QH8lXYx3F4a2Zr/t17Vk+N1eX3
6jWEmBRAcNlAymVM/vWQ6kD5V8TvWXe3TsKFNl4vBH5mirEuEb5Hom1S53SlpPHZDoWE1jjgsbGc
EYOGbIu83rkv0c8yrO4hHR5zhKi8xewxZ3O0BHFQnYaYvBaRWICzvH1Wm0FwX6gO6ko2DmnZXFLV
pMJCD+AFx6otis32jr+HvVsxBbq4xfn5v3tt7zUIgk2lUGB3IWuscqlODPQ8Htr0RR7/CaImG1m2
AkoYCn6h3SpvgFPPuqA+CKYy9mfA+UYHLlQlQ89EfOoVvvGZtMEK39zEiifA2EW/UPbqSQFzsbbe
oHm0UweC2snnxvH3VRlZHwsbvEWGmsha1mlv1frqCs8CrvHB3xOiApwVWp587ocKMnTy5PNbK89Q
wRYaurrY7hh/XpJWR7HmKUeqnvh4YimDw2lKgPIUiI6uTnXfGo8ufMKfVxmO1x87uX7FXsC1Ir7s
DKH7RVRMRMevXfE18RWDldBAuZ4PbdBjGNlobFiKItBejYR8EK+9d4NuloYhgnp/lrvmDghIZPD4
VJnqnzB9YbD6rm8yJg16tkJnqOLr/Ef2Zfb9XAN8u4cILN0fPlpnB6/ziQko9BYqrpK5+3dQVbqY
+CFgDwQTAM36w0Y3eO71dyi89qayc123YBawBeeHCHeDay0fODUI0bmiGyUeU4XH4Yacq6Zr3KX1
2zgJh3LOgFltzBMv7EyvWL/hT3EW+WKW9RZ6cdSij37aGGKWnQhWI0cHk209hgEan65L2kx6fDkg
bcliv8Ldj2BQHjycoA8TJyby3hD2XysU91HfnF1IrUUJAlJd4aFuTEOInZQOdcnuDxV0xSN8FcD5
WPJROS7jIwudPRusWaTSDPr9D3GfiQ5SWzAtiV+T7/1fAPzMVBcepoX8bHKJQjOD5GC1EvLQXDLb
h4qfEgeeAetyGU2oltaOn0oB45UkeawKMZ8zfukDwEdrPhYzO0ZtrL6hNpHD3h8fJ0Mv1Unuigd8
JfLhB95qBH8THtS9J7WO/WWrVgrkL9Zta646Cd1Pa9baVCvDT90JVMR0n9Fp0UsXUEAjSKjaC9H8
VF93wAd0xedEhxt5Oq7XJ20SmOrP5zgQ7CfdWiz2YSOiDejrxFPSg+wDLuw45qW3c5xMlMRtLVtz
WxjAimReqlt7KwdDjnR0n01xUqPJdwr3vJkhVvDZHWA/b+B2NPd6ImFjH4JtM9oCDh0Wd7x2aU1O
ANi11f9WavHhy+WZ/BnXPlU0Yg5d7Wcn8NnrXfryql24QrbJTCD4oBH/rFRQPnxBoWU27tJ3nDwR
9uvnEc7VMg6TSnXJrpVGP/JPx2mcll/rxZmC6LiD6+Ht69O/Agx/IyB0CxoolRjX+8S9SGl3WiDW
SdIQSfJdiHoROGwTG/Wpm0YWH2KH3cjYZfsGVkTLp9Ywy8IQfiVOu6X89glnyxWiEZ1qnEjqpaZp
TKlgYQY15oxbb+wEUr/sDLwZxfgX1HsFsfw3592RD7hzUozVWsiVgmoUvvGD/9D3afzEbpslQE55
WGzXnU7XkSrgsk1vq5OyZYg9YHy/TztRF3Fw7h24xx9EfU5Fh7hBL22GfGqWo+BZh6nBPvszu+Yz
ajfWkNvAXO4HZL0i4LBnwVIVWxgNYlM6eCDFEbKj0/jQxs7z7039XsY5oky/kN7PTkH3EU01Gpyp
/QcSMbkOek0YFLIVF7sqdcBcjgoXMv91eYf+3gvD334Vty/BjawrEwu5wpxwGsxH4Jkg91Z44HWJ
2e8FnG/s1rq+vuUg4nUWsbmPC/ne9z4wlkD3mVnQzd0molztd3AL30PGdYUoUoGoaOE3D3RbKDn/
7Rni6hykil/zjbkTVgjgcsWm5ED7HMMa7IbBnwbpcs19dJoXXPI3Mf8pelpVnEy3TgAjPyMip7im
IEpWdP03Iguh0pswBcQ8R1cAl7zYx7K0cr0AkIGCeuCYY2NYq7bKyFXUDRlwNo7mmII0QK3HTOJC
XCWw8ocI7ke8zsKiN4sXYMC0XUBS8/tbqdlD+vyS4lxaWxd3X1xyaZZ8tznnhIQ+StM+JDk16PWc
XfG0ri6DPKJ5ilEAAH/VAUC8aBo6gaVeRDWp8bz19ZeISOfDyAcJ7bKH9wrXQDbSKbztJKnXhxOo
ggUHXc+r1e/QaunXdokdX5qxbbI/92PSdsL4jhlSCVXPGUWNIdG8fqq2Pm75Y7GUxPVl/Jskk98Z
RTuB4Nw9Q3z7kDfmKgo3d5tEY1xdwwaHKZD1qUBX4W1hFCigcQBtQdzrmEHYPQ7Gne//W37MJ6M8
LhsNKbIl20c2JdKe+KTA/cyNAk8n7Yo3j77aH05WU4lw1n0YWu4+xT54T726MKrtwQ+co+CeM4PG
8SqD5GnD6s+YqyqfTTQfFMN9geFx0ArzOYDah/a5HZ0dowu/ZCZBW1a8/6+csHVS799YquBBE/cd
9chJt3wP8M1ANB+z0mlPbm6N8K1dxn3QPBN+WRl+JPr0mGT07NdJGjNjYnnjev32+FNzgFSzVb4y
r4Y5WVM9NIEGSGg8NcFuZplw+oTJXJdmXHCorjpXK3+wjnAQwM/xu25V9Ix6qSDp52nOIXgriHX6
sy6K1zjPxDiTVx679pw3UCjfZVGvykeCEbf7j2E5nRtzrFwTMNrFDlZGk/9NJIrIXM4BjHM2sfZL
KoL3oiu2YG2DS6N+8b7RUE2ZSv0TR1JVTt/Iw4APb1w2L/TvX2gNkaDr9WKu8/YeofXBdzbS/ImG
rLGWFD0zUWm/HteiL9kyOfvV1ZwoC2IvO/gWpB2IVa7sR0WfTR/ttHHJP4zjec+rKuEIQdigVHTf
Y8l2A3bBS+XSoaQb0KkeR5IHfYAylcdXUFiTngB8b9snDpwKW+WKel7WWYKw+eKbE+FJpzE19Bok
0gN5NGxho+3c7gNlJf13QJN22wJMT9qHzrrrkwjWJ6cBzD6nAhaQG2VRK6hqhAehufMFjsCpdY3A
iDVtiiWJlQI8GFuvkj2KZYlvJGx+KPFm/dFss8WK3zf24URNWqzuTqo0Eawa5aJKzZTt+u2aLsIg
m7zamNUJPHHx2KeH1EaObB6jXu+9OJFh9/jid0l9sULl+H56QsTEbT3yqpw5366mKEUbRBafzvci
lrTWSjUnoNkiDBHJimwvsS8kMdoBdGQ4l3EMP57mCcJwR/qR18Nbybw6MW2ceelLFviak0j3S7Zz
a9YZvYpPKGCKT+CPw40M8XZmeYPrXboAGFyj/LcSfwW5VXzWsoqILZk9ZajQL/aSQxZePJzRYpvB
gNPX2BPW8vdOJfLfpXxym+8Hsow7EhJU19P5P4bPe2fbTL2bDcau26k9qyhCbXWyBLy1bFy5pbeY
C8TLY6QmtHVZx27Y4jG10d/5c5DKQOo257Jc48GBISnr3yFCGZ/EunD151mTFXj+Qt39pz5F7Smi
0UridcyeItm4V7nlwZbsJy7vqQXzQROCkRjiNFsYsF4TpFgodj/c1HdyHMo/V25q+89OUr/W8TGs
UBFBUIdLoXGwcrHya555a77bkmg+JSUgU6+rC52iKltglf4I6Mf/Z5lGieO/kW6k5dkTyTBNMuyT
QzZoT2n03iLjl455f7IIjfDZnDSSkhYXrKG+xtdiuqtCP4hcpjxAg8vVJ+0MdYH0O5fZnDX3lgrp
r53nTSReyM8ikvqJotOTPc4DpD/p7vl7/oJblcLN0jwcyRbG2Gdi8SvDZ0NWJlTlk8GwkfoEdrrf
DHM/tE76jAtWLlgX5wX7Dpiy5BVTQ4TPvZgqlATAlAj5LUEM19uJ+mWpDx2NBgqcE63/25/LqwHZ
XuSv+0QvjwbhCXNgibMgNhgScadxXSaCIo9lzAJfQYmmooOcYrH4JYau8OrJsYVxLqKA1244k/iQ
4EF3vWxnapgq8iajmWcFwNsGH92rYNMy7Sr12GFzTfvJ0DyGfcbHIEiV8gHSMoMZe4o7//t6z+Qi
uH7Mav90MebEregRxlndCO9SWwlFmfuYqB3T7ISVJ6AdnQBtyU/Q1AnwdIWZpJwh57p2NjGAqtt7
bWd8I4WIvMjmbKi2cP/92kWPRib8X8feCn0YuBu5hJRuBXvBzX14KasUc91TnSv2vYaojvADksjS
0/2UzSmlOtSw10pxmO1H7GP6rPpbTyc2IGLDgEL9TGA4KbMeFfOHluyi5txULdZiyhCkLX1ruTdq
1CZl/aY609yzQyw3IPpIOyTA6VcCjrPelDqrnhGPkZvSL1Cj+a/DlSjlleoYWhZvXhEgJ/kJo7LI
Q9dLK0jFqKGtJebQRgnCO8FhdRV0moqhYQCl+ZLLAPnHh9DbLK4VZqeI4EJABrkj3mou8ERqsHOP
HQcWtQIyVGxFdkNZM8A0WX5WafrcyJEm32Qe6pQ2jjno7+kRzESGwt9HbDl9D0cZFo0yxiJ8RfdA
UHZS71auCl6XjVvlKZlW+0xjxPlHKsC5/PBAt1RfddKLAWVxKcKy2hjxrbnCCbb3WdYKVSznFnAZ
HAhIP4CqfzSJ49QVCDeNETEkpZ8LJJn2sxqMT5bWHp1sGuq0s+oa6ddDk+G1zkLXDzacSeBv7ImE
bqAxzhsGkrg2uRFt86Z1B3OxaLg4366XtYvKzEwYlqJmR2uSb1XFz0ma1Y/FXiQwk47GLrA6VIRb
MrFX1GGxhVBZNgMsQ4Al2BM77F90kT+umavzTsxRsJiYkHpK0TX11Gaiu7P8w+ljnDNUibU5fG2Z
f/JZ7rY7qj073a9QJ98/VQTMe8/Dr3Yl1qgX2eaSDDN1VBtBMjtfXm9xSZVu4fn5cXPPj8xeBNyw
X3VF129bG6HrQM8DP0xt/ceptA/xF5tDWyNnzu/CcwY0MXODKCMUBoHdggVDmZLCoCD7a9HAixWi
awtRKe0/bAasBgNmHU2rAIgYXCN0NWyWkUjbN9dPt+kpAQV9kGCl28daO1f525VWkgRaw3xBBDgz
XiwEVJOZz7ZQsEbEmCaqP+nOYFN95cCQIgq6SzgPuCqMgzki6KFKLSi0YFNXmsFo/Df8k/nNNqac
NESPdNS1rnb/72nkXftf2fOConagkGewITOZkHuqXhgYSmainBFV3huUuLsxpzQL+XSzVT/MRFd8
uKJcbD9bA5fghBx01ff2lMzrAesWWpxlRniziU4Ek61tUhx5HD7GogzVvzNcceLoXdHyCvUn61mV
nowqy/F34qzVJZe1raCdddPyh3L35b6+V6CklUx8a6lLyozZzsjWS7cPFT/hl1Q+pRRsrZdATbIr
6GGyA5/5Fas2bkaXNcsoHo7NSTNLbZWrH1Lw+Xq6Y6hRUJBJSCUEzV9NTWclzUSZ5v7iirx0Miyc
9O7XYoRkLqrHCMymS7MdZmuw6q5zPrb6doCcYrmrhbR6WgW8BUi0OJMXMmftrmZTvL5GolcLJp2V
ROPrDz4Ca/UCp8oW621nCowojO9fDYonYDUrdNNb0FWE0AOc4bHJeuFexIONwJIliYbueeY6Gf7E
mYTtuzl1vJjU+vD+Zu72uNK4hKtc8dLBaA/usE1wLe2TVPpfbYqMIjSsAjkUoUCnS7SfiVumonhy
ypSk8S8F4xjBie764J4V4kORdI09M9CI/c/Ko1xydehaI3lh7MZ0mMZcum/M7nBvv2o2Q30WoeBg
HM+hglyY/UlVjym7ml5uNipfi7Cj3fRTD5srtNYguIjUYTUMStCVM78B7X497+rEkvcGsabPo/7p
Pn8SC+5cURfz1G1GBmGYtfszp3gWFS6tdS7oqnqYfMa+lOdfchso883y2Mdf3s6H2oQM6HLNmUQ9
CPhcYmu8/IC54PVh6CbRQWVQ0DySvjffebsLZ5thO1bKn8IJbtIKt/99yaS9o0q1kG14H+Z7GpcS
A7zik/Tm4qBWGE4rvL1p8Fnch3njPKYQz96MTAiOteoLBglO7xKDSVIVn0FO4TT+LdGAQlyGMLYl
R3x2hWZz5TcXtrFOhgbUZ1O2IELQcA0bN5Xnystgz3QuOkTWvcCk+7OBvYwEzBNwOfpIulN7UEMG
KrwwvQKEohs6xwx8/tZH3fJOG8+MqKml1ZZN00Sua6GpIhSMcLqN1LDEikzRhr46aGX3MAhT6hFQ
hTjG5c7XNDP0iuNiZSNu7e9+joBVXGNoUVQ8dg5oVx+lirGAoESXeM5+4rNAcmv3DsEh+/v+9/DE
TuXWJn/UxtyoAHk7o6JPgLOhCaf/p/q4kUkPur5GJE4dFV12tXGqkjid2ACsm3Z35IbUv7AuJ6dV
HtlQxIt4Q0FhUy6miJYrRyO28ZqCJuralt3BXkCnH++lMtdWHrT+c2mS7VRWPTPxpGu/QLllIz2K
+XfCT17npuH3zFjZkVXIl46OLKn1iW8wKgs/pOjg8o+z5H6XVbnamFxsFVAZUc2n3mUpIbLuutIi
EBzdUDdMa/yTymExsErlg2CmpbGWV8dfTUWmHKjzfxw68TD8qLbOUvfqO/vKsaEGCm2D/wQjW9/o
pqykSD7J4xOBza+G8Khiv/BwX6T8wKa7fzPLg1QlS0FxQHLXAIRESariqr0m6HSmlj7PyTPWiOHH
p2Xyep8cJlmcrg6P+jX+i+Djg19WepPLewqrj6x2ObevyJcgLBWgik2tY8xBvywc9l5mbc3NfKm1
1ExstEy1p7o1wo5tSgs90aQc+FrK2LrnedX9nrsl1hHvEyKHBkTQ7UncOIjCFA2YDKtnmhCsyrUy
ukxXSiptfyMgmT2hRKGGRrHA2zmjfnCpdvw80U4O5K2t4gh6Zh6Kkr1GitP831q937MjJw0ZvPXV
WVlZU2w8y5UNuUdl57BUXrwD2Vl8hks/En6SVzCfVImCWqH/VBnVgDIiHD0NcgRPyeehy/hWH71d
lWnnUrMW2UzHH4f0qvS8o2w257YDCU/R9m+i8eVHrf5IfqK1l70K9r6fLb3l06jORzKZxd5Lbd/u
MMkr0O7/sFxYP4V4iHv1g7EfZE+/EhOPi4/RPz77ICSLIN+xbOZJ2FcXBtDzsrwHbst+iZmhlQfy
1odMIa1ggGrltFTyDWPNgdcneMKURMyPORtA16kLHYQEkIwnS5vxb1OioK5qCXmPRv1FineVfxQM
q0InLbBNWHY7FAKROmZS91gyJk/cFj7zcKIQq5vjgStw79EAj8IM+h7hGic3Hysx8kRv6b6pB8Be
jikkKCmM0qFA37Z5JFAjlu18rvkGJ84m+8qZ5uIu8yZkuni7xO2lrdto6L+CC+ZQniXpy3KdhXw/
iOlUqWdg5WVUqHOSn1yxh6x6uo9QKLPdkzPK7p56odGAHFCWORKbjvU+4iyLW2UHXjHq6eR1bEj+
8Mdr3ZOTiCBIfo8JugLwgNbBBcFR+lyM17ZAXdsYmwHt3SvKBaP70udgWAzU0JIUloouFvKPoA5o
Dj/8AbnND4/Znnc3tcc7e/4cRZuws1/N0ffr18MdD2yRJTWIovfFdRP8fsnj1J7HOS0DPbSob0UB
ceKY3H6AmcamZBfAw4eVRFFOBVP6wZYoZihBkyiErvI2XuMq4Pczqa6CEoSekUC+Nif5vwr//nO1
D+tP6spxtOPRULSNz+IrcUlBU6FlUKiILZLvWAKL9gnB7C7cWQBzNl+YgYXLrxi+u0zCPerLUbLG
JdSe7vTeFCVIqTHD06+Zv1GWmT4bwBvvue0dmz8ArU+wa1Hd7d/O+iKzndT8qPJJ2JbQ1MklPp79
tyRF5OyniPocXm/7yxaFvTNk+jOsdYynWyZ0ndorSVFQ7STtecYSJkh8ujAQ2cHHywT2rtxw+qwg
+cUeGxuml9FGiq20kjQ9etvNVJMpjN+UMKjjmQBznJ7viGJS+hbAFQ2xMs1p2/mPzeIFiS6TkaMl
pcpIuUM5GjBxvoPYDjd39nWvsmHj/t9mJHpBQ9CTZoAvxgO5Fj2QtZ1LHuYkaPBU1XjO84/4u5NZ
ADzeUcA7OsUgiKOYQszpOBtTMFQ6Bdob7WCU4uZbnesRmVIRNp/bu4emBhWPLR36WwvQ1mh0Aedc
lU4gqRW6KhQr2HSAn7ijkgSwtncSJi7CXUlGxCPTW/mLn1znpJzlLZSX21cBOUIiNO9pfrsvsSdH
umWLVQa8/goEgan0MmRbLyJ2wvSocvPKi5MyBMEsSXrFbqJ0Z2+HzjTUbmJ+mgeVRJSiEbr8H/OT
P/Y3FuXVB+4++FTFMvH7JPy81LVsy7UmO6+oe0ypzlAY6p8JMzY7LmTxXEyBCkA1vKV5Lkw08gDN
5GR4/C8FKIrfYhMdqZgYXbjhTm3EK15qSLgGE6LjJn8ejVueZD2aG6uiTZh15hp149hfAtFDm3iA
GPk/aDnmU1EtRFCb15pXzH8YsFqeVWRu02MImBe3EW+hq/91BAob+UG9y/B8nu5TN8h9CWjgSX23
UEoGFORIQQ2ENJsrmkgkIDcTD4yaro5AH7o/qZkh3/IEJxSwTkg9nZuMMp0QcUzDcOR6Ngas+bfM
cxvuDPUB1MsYTNJ4Ebm21/JHUGQmrrSisxQVzkLbRYR7pY095I63ZXmW/BL/GYoywzFX4tpNKLwy
CjWfXIRquUTe7fURqsRcGOultFLiH0/DiqqpvVdpdX4qZCUCqr+sslj6qNoFFAOmbJ0ZIWv2dSZk
/HyTnxp3PbTHoUzrtK00hqeaX7uM4QmFn/KXaHjw7gvk+FvVldO5QvkfSzgV2ZyQRnsVihp1b5NE
lem7czQUmLCZr0OluwBXl03OV+E1IOVHD876v/tbF6wAY7iH00zr4PIXdebtkSQn0tf/RhVUeF8o
+xBwsqdN77yDwcyK5PhXy5Fihqnw4hagKSphVEsSYh2RyYkafRcT+XOzx5o9VKUvTxgB35PP0oXP
TqsS6SabSDs3nBwm8GEOFy9LuN4V1m9DdsfdkfOJqpbcYb9DdNNB90/zMiTR5R+6ZIg5JSQ/yodg
9VWPgBU21CekhvW590J/L0dO1PXbP1WOOsuc13aYQuxuIGlswpQ8tZqRIiBfUlY99yxX5e6abl8/
I2Sps65zun7EOnBmef6Qr+mj5oFiv5RoqzxzENBynZzhOUSHeZTA0eEB/RxQttzFoO4dKq+/MaUc
UplN5l8E07TZ5tozeNTSUSbtfJM8R9NAXhdVDHmdbr7k6Z5U1Wxy5W3rqOzJ4yhtiAp7jlCPJLS9
gGnTEnStTx7nCJJjlwBAA86CIFUQ5ANK/OXa+ownaEWqdZdIjWBfuac3d+cKCS3bfCV8Dc2GnwSW
OzjuiJn3RHHWxCmTAjUNt34GXSDkTXSjH4QxLZu5UvrRwk91YBbDUBGtN5sAcH+tHoggIEK6k3Zp
sViBMBKvdrN4S7+1DJzZeJHwD+0H527I4HfOYUyKUWyerReDoT+Dw3dN3KsP90i0PPWmcOUK+d4Z
SzsQzKw35mK3GL8enYnrQ2KRaxlpWH0ryQw94nZl3/pGkA8CknvR6uF5yxEt3iS976rn6DIAekwx
NkemEfjEHlTomDOoRzUWhTdw0xHwy6kcBGUhHdg9owWCB+tbV6W/RnbjTJ6dBO0N2J7B7amRmYns
vA1UmGzpw0CumNpJxOfAYZ6v8g3Fe9+uRPycH3Uii9dP1ULM2tcrdk+iryfhwFiZYCoceEcmpxaL
pEq9FIQf6RvELfsCb5NNz9Iff0MiwJHEhSlB58WXQVw/ZeSxXoVn43TH6cXMZNA+brwer6TTKGw5
VHCMxKTkcoaNrSbpKL2K7VmIHJKruhWTBMqcUMJo8u2h45MxlNDuh2thxIqBwWOGZqQSItCBhfq1
9Q8aAHrBWzu4DYjYKINccV3thGmJRsF/X1Z/WK6cc/rS95/Ii92zMhZT5eyB0IMgC8XpM9640+E/
vF7CrOkDopPl8WhCT0wDbiEHCrAiQfQ2o0rJu/hIXutZ0LN3N2TpVDGUlGw08ZqGHeWbaKiIfZ4F
USsc+48vpzxBZO+F4DSD120QKrWhtR5YpHnc3lhJONV7u0GVi71XO4l27RV+NjRXjX6F3N+NvTeb
otXDdmh2KWEMKj2ZFy+1ZAcRUGTuK+v2TDrkXf56N251mFxxrjpF2H+fL5tu4ZnmDA7W95aeqHSD
i0x8S9w9xIs816pGHN+Cw6Pz9nrIXLaNL/1zdp2zW7P76kkgjyNdvMGnOqtbdWhoeHfuw/cEQ97A
LeYSD6NqqElAGz+TYsL8WGADC25NhOBXMYAQZQaOcUsDzXmtCAibnoBk+i4gmzrbbjt3aho1o6JH
ka2Gi67ukCSZsKmMSkU4/v8ty7wiHc6XNLjTf+jNU9Nys3bvmLRbiQ94sGv8NQg4TCHitKT3IRMt
0by4+OxdqLBkrq4NfWQwlTVhDnBbY4w1YVpD5NmhOJ39nAXxaESOVqOWVZGBzSprL3J47QAXAVA3
VK2DmPUBSRLjeQ4KbFQ8zLY3j/p8nW24A6UcnJBt1LnPp0GjRilHtbEhTXSwZCLn77GVxfCS0QpJ
JOva02dijRttna0wBYwtBCdGNJBuRqa3S0Xwsv/CMZsncwLXPpDIu9wdjeKiPx7FwjQaWi1b69H9
wqL7FCs78NcaGyGtmNp43O6ejA0RRyodBmFEPDhGgq/BemD7gx4fH46mR29vgo2QQXzdA5RN+/mR
0BYLI4fPw3naD3zFmgtjIjX8QD/ycWxcE6H9BQdbL5IJXQ9R5xu2Iu9Hsg2xHNxNVqqr95PZ5RqF
oRGuAQIkfJLVREydEDO3BuFBIhgoldi2Tk2yWpDRsJLUe1G/m2wBS3o/nRIbbWPVTs7mitSZuZzE
doLDTOgI43ZQvgSrNolCvFkgPOvgiaRGeCKeXFeLGC9ryvj1aA7Cpet7EOr59jdD6XFldjj66zpL
9+ck0SfK9oaFTrNNXBbs/i5HOVp/zs9tWfusMps9ZapV89h0nNNrH6bJc2Bu5OnvgMVwCVsysLHB
ye/K0Zh4hXWnoHiDpJaO/vBIEO75lLMWZDGBGT53VCErOHne/PjkwwhimpHlYSS5WSoUe1LLMetq
GFfK0BbS3OcEMVuiTfS5fsDHuhNxqccWkp7q77NnNoQIQ1sKzYLHPYn9Hd91QEeQopwO4SsWybVJ
Qpa146Pb28giwfIzb9YKn7hsKtMu4jPglByanLQRAw8IEmEcth0kPhqXQUaDawOCnqBiBjY6UcyJ
K+eEqhK88XFEMeuaCeYvIWxi/BuD1BhsCh6WpPY+weDb2hckbIZDQhUXXmSV7uP+xWMZVX/xS7g1
r3WghfnVGUypYKC4yzDnb8vcN/7pQVRL1+7ju2/jyaYa2od4bWN9oZH0uivec7dqGnZaPWEfiyX1
WUxrq659GvWZkI5rCcGnd3tb1dMsA/CnEvxUiCrlnbrXvyF2UTSC6VRzl+PiT09FUmJ0mgyuBFOc
CDe4wpgHqcHOK8UfpOPy9E3aoQV9fTDt+KnoD22t7iuf4Bcg1UxShF40Yhhl0jgRkXYLKrlS12S/
Y2pO494jw9Ew7rEke+PgyvPgIDncWvja5GkIipMCjOdh65wpXWp/kYQ9X/A9Fle6tb+2mnU3DNgV
R6GEZLd8VhSG9hmmNUGtCzyQr+sv1yrRSc9rESorFuj2vUBSr18CVUbpeki1VJBbcpzvAeVRj/ZK
EN9S/Iv/M2MqI0iErCskOLJf1KOwVS9omgEN6w9RsV+dh5M0/T0IxhVt0arVtY31Rzg1jCaUvlFv
VELXvuHbnyYz1ueluJtAZaQHjOoLgwpw8IeEBOo9l4kOA6A2G16D+pLvQ7mjD4go2s2MvlFR/llS
McAm2SE1/gO6ZgVNK9YK+UAR6AmaEVk7loczILEvuG1l1zzIr8fSHDgtvLV5R8s04mHzXoCT0fzX
/oDUaObJ9WGhKSHyiCwGOJYcs6VT/8mGPgQUSuVcPzj1Yh7qL2k6arST2pQH/YcFZ1mN8ZugC5tV
coWfHCE4g8EF7UxQRDfMn1MIprn0m9aq3iBnSyw9Jg/vmRmYVgQF2zrw9AqjtI/f1jf3uxqSyU5B
byILiDHKUTiv4gg49zuA/FFy4XquoTGLdiZW5DXdOIq75nhwQ5ul+kW07cSoLxu2CG4d773dLdob
hlR/nc+cVJ7bv9lT1gRA21CH6kdbxkxGtix7xC+7EjdlIU2rfMRY2q3vy/UzsHpcGwcfb/IUiUCV
Yx/oAlv/tS0KN3KdpI4XxQWxzEiKXI2nj+QFhoXW8PlNereJhO9OJVMGUd1XA+MC0ngniz3WN5yy
941457F2hHNMDTgyB0CMOOGnOcq4k4O4eCbJxhxGckdNSnbiNhSMXg62/fAoYaFz4Y7l/C162OGv
Nvkq8qMoCY5n1z1AY0zqWzzgp+ftcFDaga+43ZuMYZ8K6xeeB6s4hrZjpzVp+0USK2it/5CZKDT2
QBggLKPSCL1h8vg0cNFWi7y5YGCeC+djzP8Ls4Tj0D6/ePI6LcPSBy737H7MApurroTF82HVdU9m
t+ZHrXUauT54/QQYFaw3uz/e1iLyvvxfEZbz0zE7Srj474iP22lKy6XIDjwRZoXR6toI1ICaxmM8
4+RFrND/t51uR54+Mxe221ItZxMukOLgtk9kMiSZqRyOoeoFwxL+jHnMdBpocAUrXcREVtf6BQHR
UslbNfHxxb0X/oEdW52JmVNY5+gyXRDxGGjG4pQsAZHcVnXOkz90YYb4ijUXX1w/LsALNDaJtOnf
CEF5AaB2/1rHSrE4kB48Uk1Y+AQe07tfxGFSHkikS0jbPhKT9rbktMVY5bvkqdkRZEguqDEY00pT
yh/FUUGwGnWJjAO6Jx/DO6yXwK6dqUpOgqdHJG9gCWDop24wHcGe/sXLirHYOM1HIbYV6aiLUfHw
c9CmJ3me9/UwFgwQPkvS24ZtZa4e3eDrYtVTwQuHoGChKaAMb/qsV0yxJl+gsyQGwlDpSoDsg8r8
/zBKZvtNpmOm4hqz9v9AuJP2YFkVt879ssQRWdCuewwnGUApQ2Qu6kP1Er8i5lFsxv/5tutW8cV0
o4MkP+AeMbT6/jCxRaQVWPznWSUpZqVPzklBmRkDHBdCtQBQc9WHv0e++e2IwXG1uFLJLtRmUddx
E4GGKlieFPCFNCDdDpkmwdd1wAVe+arP7HlIR6m3VPDvwlEEYpn01rHByG7vCvZAqQRd8yYXNWcG
4ami5rN4dXygltrN0UFMIXDqusqL18vyKIddSPQcKprH5SrrIoy7f1DHx3am2rieBXjt6VVAvP/E
DqtHWMOGasImz2mTGD9HClE2AkHdCUfJ0L21pVTF/WX5kBtddNFHZ+dd3ACYa6EQVUT61JnPY/29
ppa2cAfqwahtPZfT8sQZzKDqp8pAs9ubVxkwyWaASL7AAVBcTAneYx7iD2VC8d0kGbD6lYOyv6k2
X13c799zPXjOp76cb7tGRlIDrIkTxZDw/RIr+lVntFEsSISN6tib3kUTZh54yVwOEKja6PyY+1zh
Saesoo5nSQUzvleWkmLHiP71KQjLxWk+fKt936vFdRhL9MEIuFe5DDor8kc4HzgC3g91nxzrLe7E
PCq3jp6p/+XvY8Y1V9L72DxZCE2y39O/ZBAzx2qe8n8kU8R20UqfKaltLe1+nGp34Dbi2dxFZdQO
BEGeOW1dW3U2q3wHwQceif8fCf8fYcARjyTzFnpH5OJvv1uRmUtP7dfMdgwxRK5iOUm5Q/aNAuTK
+AEh+mC8cTo8JlwKBIa0Ug3LKJXIKRmUz1FnqsC1inBP36izm9222+hWH4kFiE1icS4Klq10CwU+
YQfphKzwmNuCH/3O1kleSF1s04x2DlcqiAhRrQpfY820psQtUXYTHEZAV1b7iMkIVFXsRZzGtYiM
1xycdt5uLZHpQJ6TdfhMA/8/55eChDX8+5thFEi15cmVOOM+ZTFQwPuJbey1R0xExqXiWpFnGZhG
9mN1FJEnG0XAf4xcY53xZCyjrhxKpFt8rPD72N0ikGLzF1MzGzunONCogCbRxNcqyTshmhzcE2vI
p6ug9jlIVIRjEXLNG0iLc1lJOf6H7F1E+XbQHPz91buwnUAooMzGf13yPmKrVYE87q6EVDl/26e6
2w1Fs4M5D2MBiHSTYu7RSm1zPT4aD9d+Hpvd3BO5zB7VOdk68P92FhcvRrhTA6WlTTk2zReZtP1N
XmxZ76UkDE4Jr02S8pGnlmbFE4wEW0gRwdNV9YQ/9P+GuAmwLtL9ZoyzrXfk+KcG7Q7+IVR+JMkw
mFJuidp5pkbfyNZ/bvS+mhhYB2JERlE6zWkE47xm+2yvjd8Mwwf5YeFzRQ8auyxb1EEVpfWbe49V
3XuKq8mLal3lWrPt5HM0EsaC5qPYxbEJgA4z/teUzgD47yzKMWWp1cK7yO7PtPai7aGjNik4wxaI
z8GiGD+osXjPBCTmgAKhkF0nrl1CHEFI4RFJamu2G0E715SnFB0DiWfUvcblwRoZ39+PY7Ig/AwY
7xT/3FbAVnV4nzc3AVZ04LC3GCgsMYO/mH+M6xljJOkImH+8lDQYeB6vJdJiRmWRWS7eczt1Dbao
rR+gUTBeQUqV86nVzddGECaU70bN64l9k1SloI9dPLbFtqpiaWblaCbVCDAKKlGpWPZ3a/BYZaqK
D/AJ57oWcVKcaKR6YnKIMZ81mDf5kzdJgHKUSClAraCSdGHS0kyG+5Vg0gpUmfL7gROEhIq0RHnA
aP3GZKRuT7mHuHVhLbAKhUxiRD2NUBmDXmvPkzo7TLr3xvdUqsyfG53hnjsj1cR+iXo1t9ubGP1d
eKEz4MIY232FcS6/vNueSevKZgh29ScihRFrLt6G9MamgXxlDXezYwjTKeFxsS7OMVJ3w6+rCqaw
ZmQLkp8jY7++G5t7p10gbfLq7I+1zEMj2J30oDQsveroiX0AlBr412oCiNAKvMGko0L+TeBsOUy2
ibbivbuR84IQgpFbfYUFizQsxm5Za2yW3XAkaLs8hlMyM1/a4kDqWNbuVLb8IX8gn9BvU9WNG09k
wZVusSOFdRDtx+qkUUjQPSCW+e9LK22ZvwD8xgkE/1HAP/yPK9DP16m66OFgSTRsPdvQh6gWt44W
3nzormyScpPpwfr+OYws1aFLREtCJiW+ZOHjwEp/2yuV4NG8wno7SMUqwmx3jPflyF8Xh9HkkGxW
LIzHvMhq8xlMBatdIuV+lfBl7s6Pomv5ro0GfyNBbHLVPsSk2mK47Z3ovZ6gciCIx8zuMqoCC9YZ
uXLLetS+RwgpCWWbonncxliZfJXjr6eWJC91sGSMSqhLl958/kgN3fw3i7cHy5OYiDeyfRU3rZhd
wdQ+W7rOK8xxL2NHPSe1JZG1AwL1HR4O9W8hxE6nJ2F0rlAj+6Ic3bBTmiygVuhWnNbFRE4ycyDP
onVBabGH8N3+PJJ/o0kolhn3HYcMZfG7toCEkmokysPcc3cMk8FCnr35henhxCgKgf8FSbA6oJZL
RpkijeGwvyhApTsgZxX1SCGPWhXTrawtxGyL3oRrptbGTVbFDAc+YjSdPLuhsBzL7ByZGsYv0l+g
m+uUdZx0cNR+0W7V5ngepXk+ERruG60hkLJUwZHNyRtTO7tjCShzeIi0q8fXQg75TVf9OeQa3bAc
qLgl4pUTC0LzbY9JpuKIjprit1DjmwKDbBO7uWfU5yCwnzyWpG8QLH/yYU55vSQ9G2hi35Uhbns9
FsNgna5DQ2An/buUmIJ6GyYoLh8qend+vO1BLOCb1OThpWjb0u07gFI1jvxymTpnFYM+/D07TGyC
7X83ORIoK/GzGQUsMoDgfWWm9kE3LhHQ3SRb7/9QffLEzpTd31XpYXh43EZ0Fk9PUfaXD/J5L+dV
nb7F5FjEXr4n12IQJg8rofmOyecPjq+nbceKaImD9zOw00LGAJsQpQpl7hZeshldmqYuuH6cBEZB
Iqel2bNWethsBkWjcXriouREOC+l6LHjZd/9iVGeGZnukCW/+6vdSHkhGnM0BPQBRxFAKuIQco8m
zb4tgYRPQNLL8OxKoTTMAufGNGDAFvaMZf/uVWXDRHlO5t1xEkKnBjOXrfC3vPMpNmryKOUpHCXS
Qv1PNTb6/NZQx4/u8sc6appi+NtkO/ZHeJJygDjEx1JlXH2QyUS/Hj7OXxvFOkjxGt9B39aIiMto
EDqi9hZ4GIt/z0vNJzbqdZBp3CBd5RCMHb7VvKl2AwpeJFm1cqpCyDc0o8TDaM+WhLpsCiIrENLc
SFL4x95hKHoXFz2TH9gcOxz7rsBB7eh6ezLZFJjRrkbIkCI42NC3rnJdJHkM6pFvn5u2AIKblCmT
mZOHn0cDd+ikhBOkDRV4Kgk3OD0rY6uHrAMcTTrVi1atW4mqT5jn/wxQrjuzcuwZ+enjWuboCdLM
M5IdRA1+Gms7D7XeomqzyGLVHIty3Mj/PiY4MmvfwLdextwfppP3YWBaxIC8koK544zN3Vrbh0kH
QxRRsbQ5Y8NzJ7OfGpJrOSRzyxMMknuE+uYAeOZDslhTB0kI9ItRIIGvwkUecOvrQbt+EwDehAqP
44uJp/gB67sqsxurF84R8vaAwJapKdvsgLekItnt2jlfSSzKU6H+A9Qch/FucxZeZ6ZyhXjYNQ43
+RwGR8OO7rJN/gbMWVahrqMSIp7WfhBp4pkWD7B66X4qj/UAx0hiDB0/mVNi4cpwg6Gh+pO04nDl
gAhgAoORjDOoWTTuR7Hfc5s8O43JGrWd4rwMhLE1F4mTyVYZjOOI5/x4Jwdd5zMm+O8Bpu2EPjHN
/nJQsDSe47xMQs0GYCkL2GzaPEpn0Qk+uN1wph0vrYo4322o48zGL9y8NAuWhQJ82MBRs+gj79RS
I6OSZmnvM3jslF+YUX/VvMQNPg1P7PEgc2R86pQka+4WSff1ibcLhBKDWduNar2DaA7D+rwqWHPs
8sbf7ZYOyGxgylGIBnZTim9YTneFHV35bTCDh/mvjnCO2NTVlo3K5WydJk6xXINshSvGzvpd+76u
DswNLtUm4fNYDz+dAdQV110I94/bb9Cs77CQ6GA/hEM9kMjNLXzRmrC+Weby50y+1YdcU7lkO0Y7
ybMbSNTbbIyvxhAKIAuLCKCzfLxJTlDFa8r6wMZHzehFRhN7gMcdxNQBAIL6i4ssg8XFrvUVHJBc
SmhhR7WUE5O1axf/hL8BjR2Z6iUZ2efPCw4jFEdeNNvF8ZqhgihDrWK2p84VoOGJHAQCBUGC4BF2
K+cG6yz0llFlDGWlmjwY1/eqDvxcr9zapXMtkGurxyWS8kxQJmSOp+lOPLIQclRjIwqgxLv5gqtC
MkgdD8nsuxaXofeEAA/CHWN7fEY+byRO6e1aWkSTBnC/xt1+L2lv4DcPEfUnr+vb8rsj3zbWGuW6
Ww45/rLW0sDIQqk1d7kxzUpfbH98WdRePNQXkTKQG3lwJ088285zUZ0kNJRJ6nWFXJDRaySBKVkt
xlF7d0RQrEPR32GgvkFuUB41Gw9sPWFCnluMXOEG5mxYHRhSbClcQ7O8fHdrt2Imo79iFJPSfBgh
r3UFFdKy/vjg/8fsAB1J70VrMpHUd7I0S27NBe2cb/+3W7HpGcZ6Duvjdoa4UA0OL+RP/0HhdR6g
crOL5lNeu1+n5LmpDxkMK5ZvAjhr9piEkohmLBfigwMoQgPmf/vDOEZdDhKRe8ZNjNFAYrz64ydi
PYrwvUFzlRH2WStimeppbMD+MEQ79Jd+RtqCi7KmGZRwvz+LLei3gORAmZNY16FN0yVMgjCoHT5H
7z7e/7iEAgvDLg6BgU/jRyy4VkQsq4PZx5QMrcOd55hAYyAUZuyQVo3806Uscbl58VLHYePgEVNA
1KMmqXfpIdNCQll3N8DSyIwNYhm/6Ld8WOZaA8Og0Y2V4jl0mb4kkNacm9kmPMEfh0dCF4iSe6aj
0biXeRjyHJf7X6kXpWwJ+R7espThuONblus/PDl59NhYMqBVvvVnSXZw1vqvwksiwQ8yRZ66XQab
TGYgjUdRyCru2Aj61DecOMZC9aZnBf/kUKJLMWFluYzH9eZzfXsx5OTMaZzh2rvK5Fp7NkLY/RkT
plPfiw+69GkSVe0PXujDaQv+ttTwFX0wh9Wy1Yn/4O6NoTWz/IGqqIzsZ01A9PVtEAiGt73ncYlo
AdFyynk8Tbjoks0ayu5CYOkouywwH8+1ufZka5O3vzosZLcmpAMD3fH41YbIujyEfN7KyjpK0TcS
xBWnlF9ERLl1iUF1VBAx3h7OQlGrQ6/lDppNszvXya9Ou2G0dL8ohdDBl3c+N498zB3NCxdlCqEj
bhe7CiA9rUi/+AmQpwY7WqEGdWSA1iZSHxAkEFifTsbgISdsCh3WT+cEfgrtkNljd5+COCqUlzLV
v3W3cUneN/nqF3YGpoxoFhyK3lzLysQuqvaExSbDjHWmm+GX1+q6dNBq1ke9mYM4Rs7AELz4awRG
Lve/IU5hc28gIolq6TXTDD1AqaqWlzepYXbiwfVwvrF2FI7wIPPvldTRsFrnj1gbKdEho/fiaTwP
H6QNWN6dfJZkNhFIIN5s1I6noL9XHgZwmdovy9Wb+EUwOlfCMsBXft6GPtrlug9gihie6CP5X73m
ILC7v1JvnOBh0g0ITldXXC8eL5hg5beQ252MyQGSBSKDZmGumM+bs7NIRh5LDQR+GH49yBnp+hit
fomndeusHz+PWNuUqloXnMdUKGnMOFc+udG5+0HLXXuaYe0QuYkdRYKTNnMuAHUAegZiVlGpuE+9
fG2JopWrojiAnSp9OFo05D1YpLWnfbsduqkM0T7urhoxDVvnAsXMZ7BEcZcQvJ/LW1xpi8Mgikut
BRplB2ECZZXdb4BWcIviuNALdUt2YzqH/AtUEoiMYH539bgYzYhmkB1HIUE3bG+mpHAf7aG4Dkb0
mZ3N6pmuI7BJLXnNNSbJ3/uEQUWxMQLsrf3sidEhdgae7fCq9Apf+ym4g122dFh1dYVanowZHdNv
zEJs+OWNL3lXP1EoMLvi6l0IYAOHuIf0x9q5xpcxuuWv3KpGfi+u3hm+6O9yhuaPU2SA8y1Jit42
T/5LmkZOxenwUK9uoVDwH0aqcojfYtpZgCnxERxFe0WG6gMakjKyhRJAeIoTRFY3Jy8Yu/Kblimi
3kqKli0fpaiiafD2pd+Jo5TAq2ViRWR31GyZnCx2QAcTwgSpUPbwZoXQK9Vw3DBltlZ/fin1Ztdc
pe1SAz4rdH7VY9T8Ra74OTLMlcu3tpQMao+/th6g8GRf8cCMkQYCHL8E3SbJAnwFo0ECfU6LM7fS
TeS3pCDlADp5ocY1gIfDBxpwGpK1qm8vFbpOlZOK1taYyClyPwW1SxNIT6mO6G5dAzRofCi2d31F
LrieaefnZSxPWgte/a35gso8RPH+6V1eAFCScTreUY+kPql8r8X4yNtsUhO8KMtQflG7JKliIkFt
s1WKir2DwLE7iaFDRzrP1VVAYllxBc+dCf53OB2Tzgy06Uv6UM5aApbIdOJ5rPp8hCTborWIJeii
t1RBFY4cCjDa5zE5fAE/FjLamR7uhGylU9RZlPqyLohD7rwFwiuCEkwniSW6oKZtA520JZNGsbJk
OS3e8OwEk7SunW93Spx0lEr9TKg38gRVF8FI3ygC3nSBuk2Lf79UlT1li14PxLhZm6HYhy1TAj06
bxl1es3O46tDUNN6eR/o8eNuRbAZubZQHlOOX/AbO1kLQPnD7VBNXdLvOn0rHTvewobeipSroD7L
ymI/h2PvPiQpDiwaaa9qkDTx0Lt8/BaBWQFAPuAzr74cq8eSj5NTWRZapJlgPkO5n9EPbtpz0sWs
ZK8g+hdJbiuesOa5rAucQFkblEcVqQdSCMgqwuOPFXVKUKW+uJvElmQp5vcOwdSh8McaT3vP8adX
ectNMqq78cckOVumDf8XGDejpRVgUXTOGYUOlZ0t8kwdW1zwUewBISL8uSDOh+doj/zLs7n7ZbYA
f9ZO3JnSr+sGgAU36mxyRLd2Q3te3Xh7wz4bDopCG38e95haK7xk8KHGHO+DOqpq5EZSqpifQP1Z
2ziEebMnb8r756OpCl4BDI4aOJYi43Kqchz0XJHoc4GMse62D1bjuA/5f61dZtmWMXcxgNhBmg1o
M4Kf/8q3JEA9I2IVOAXLHEslGHAgZavOXpuRK07QMLnPYL2EuI3xUtJQliyiCUXu7v7rcvWJXgqN
/vnv1OgV3tTf86/3TGTLMJbFYjbj1GMLqS59wPE66UquW13TL2GFC+UCbZyId+p+4+SIKc7OC7I5
fIHhdRlzy7OI1kFlTAXlt35oQYx8RYvrMpF5ZVEv5K0j5iNB4PEDNocWmCvpvCA5msqTUvF6hDiL
am/478OSwi0LOUIfgWMLYtJ4Gl2vlDw6o7GXNL01HNu/UEctS11bhaKLLYyxSbkR/xolDNx51hnw
4q7fX4A7UFmQCjUJAIiqmPvzdxUCIHmWBmZ6pYMqzwTzHuiClK8DvOXjaovDznnbyz5ssOmbhzFl
7KWjYrGaYFseViKe5GpmykKbJHSgXKUugGGiaxCWkVVcKb8fdhBs94RjP7s0FGM8IXhhaQcxdVzs
oRg29UPleYpS13wEDRcUngy18cj+0T5H3fv2DNWTUkLq1XcIJ+nZyZ+OjO3dTs5Uv0ZWK82qus/c
FuqQ9r8k9zKjLOgrYekvTP18efaDgpghJT/jMQehC/14UHgxPic0tWh/v0/xMbl0zr386N471z6x
zgUQhI60Ry0tIh31GTPAb0fvBu17y0A36UurdnIealWwYk+U/SjhT1C5n69h6zxaF7mo2rRI2PEP
pcYNYHXz/UdahqcJG0vsMbZ9ZqEZBJBGot7kPD9gqZU1jChkvHm4r3TnnrYejx+YBZMTbmyMd7Hx
n/NWhzekoIbpE8jbjnAGLM8OvhKnlJ32XeK6WofzakixfSL79Wfpz6rWfb5nPUVWKougvl6GUPP+
gOOizt6xALBVPR1dF+/sZ0jcr6AgO/vAL/iOQJWfP9zwi5cxT4IlYKB/3WQukdMJB3Z3IIui3D1V
BLZC9LavD14Kdk59tmSxsJ/DO0pwKH2f23KKGc4nLrQs1/C2JSULCIZUu1LQxehT7L9JTLNqW1wq
9c65pojgmc2AKpMI8a61MmEgKkKFmhd/DFUZ0GiUOk6ZckqwItOFnEJmh0okJiZmcPLYbgbj1/4s
V/8V0/uMu5v7hSo73jxAsvMuMXDHLBcJp0m07J9yRyjVLHIyxHAo/UyHrxenSxMkZrpD0FUckdMH
V0Yc0CqqR9jxOZu/pG48jO8GRT14eFNivtsrMoidNVrRtMzgO+o9Z8BlkVkaZTm8ksE35S8O6yi0
o/qq1XA/nENw2dwB5AN2A0hKrmn/2Sv/4WK3AfuBZC8PIiPy+5hm5U23/QH97jXpDsogNSaFchYL
ExulABHSNjmlb8ftvrLuxAH7U63ezuZeALr3KLoVdEfElV9a/KZarQNetROVuHENtPXq+fKEzkOE
EAPoen8+4av1+xGsp4GH8BZ4zUZplBP0QBC31kdou1WasVVcnIhS4F/217pShf6bCsVGOYtBh+Q1
jvmQspebeqtmPUUHZfFSAcPj3ygXhtow7Rw7c1V76JnRZ9TQ3oWpFKmCI5+1R0uE7a21vrmzy1M/
E7N+4Qx76dUCC1nQLYDiVP8PjHRhgGGCUwDvMEUMqwqffMZ45g2t0Vcod9IduUD0BQn4zRtMGyWN
LNcv86+M0MY2DGmUTux1ED2IoN2ykVL5Y3TlqiNgNY8AvjeY1NG1C+HtGBYbYQKS5QtCOFs1W2Ro
HKBcE2mEiBhhnfUmr/CHq4wtdLOsb3+OEvdAfOLE3sClTyu9vPNgUOpcEe6yeX2yhR8RPt2JGm14
Y7wxzlTTfWMjoMbdWUPboTNVfsLB70vRDVixFOoiXUFxcl/VdHhxLvzchpvbPlonsVdu8cxKtoLs
rxotpUWNMqaistrUTkqXfK4ea+2/lb6OeO3JBgSLlrhdkewn5b7LJxyY1yQ/dcZ3+RbxoMLy7pgo
EX0A5Nt19xRBmWU+y6OJ/OSrncxG6KuBUx9em9tJP8FpT9Yap7zcbmFIyehAjRMmKTO8RYqj2iIl
GrQCpQgQ3d++qWKG3b4KvjU1enP2KShXoMudqznXGTQHMoTm4nfVIlfl2fTK9QdwQR7iwML2YUiw
E+8MZdPQVPZGOClPn3md/Y9h0RKfju+qDWLNtJyxleFW6Xi4/aDs1MhXZttwu9caP4g4LFEriZ8M
xdHXKWR0VkQRhXPInQ2+YoQ3HVmqCsJg6T4pDSx1KJ5EtoEUjsN4aKlaRN4yV/sRi23qOWn1pOGS
qaje7J25DOMLYemmOH7qMET/amR1slKWuFBX2E9L45u+/IA5qSRuxcEIaQ+DvRIIGtMnEpcw6I9j
RExjPVoC7bESQfbVXpLeVwHD8QElj40qI02fJRfxLzWjA05Q792sPS4V0jN5lQYgdiMtrLrSgx5Y
WKKXE/1riBhyR2lDkebQR/nHf/KtAOs/5cmecbjxu1XC3BqyAITe2delRqshgMW12KNV8QokHiz8
V0VYzuCYWDzOF8nLTyDHOjagXvfk9PbvZf5eQgRDiBM6iTfXNQ1sA675FXK8TPTTcGu1118gR/Eg
eg+pu/MYCIq4kh5nlW0ajNWwrDv1y9lt8VbGnlh1THYLDzCK1hH5X7G8qGamMEENOsTUAmsHJsMp
Y0hQD56Hq/6/dpvgLiDn9eCmIYGqKrP5GTXpqtNPFYkTQ95qP3ArLH9+NdqOo+H0y7U/xvB1l76l
zKyXLnSIQiibeDNYYs51yYBtT0aEfxo9I2HzjfSeJDCo4brUHHZNT7EQm83FMEIe4WgdIWIL35wG
V41K4nt3Vm9QgfWA2GmswzajByRGJwAOzScsibVxJ7JWTyfQub5bkmdH0EUZIYoFfO/DRcdeexEH
6AVzHuCzhrbNz5tUipHMv4cbYs2jhqUUE6xjPtvhtJ1W+sILIZxs1Rz9s7Wf31Rg27TdskxSbRyp
PxL9FhnpfRBx3FbMc2t42DPA7NaEMpmJs+wHX8wFGcKdgJqexoqtFyhvA4MPZh321575rAWnjFwj
Jzuouli+XxWwHrfvQUROnMJn2yOzolrynKz+PQ3KLfQJM+8/ZnDksgdjczP3gfkA86lqAr8qlZK/
I+Hv7hnOjp8mxTimuNgoUEvl9zlrmZkwxet1mtcEzbZPFvwo3fyDzWGc7g/8BY6eHfOCh+Bv0RPv
nX9HuKTdqL5RTAPOduzD6fZnhJ7gCSoTfOcbjOtLjlJJBVirCsSHHsUhkcrb/JyhJnRhTAEryRZw
yjYevpDXbuN4v4n60pjJq2kjBFrJvfGFfDZt+khnSjUVeWpKyF6jnbf3YNcxUqMexJ+easyIT6Tn
cUhNUDcc45wejgdof14N4/xwFsXgTdu8aW4UShggUiNH0t3RTpBxiWYr/I1U+FVP+BMJHUdQ0uG/
6sMtGrk4wJDxRl12HWICpRb27vC6x1NEzqP40pfozNHUJYf2EZkvxmle9tSSVW5VjfVSCYj7FvuT
3zlkOg+ohzVvc0z/nZBJQ35YE3bq8pN1cRNOgIZt5UGe7R4mZ2EiOI64svhSX9Ko/x6Kjf1ftBkt
cc6l0fyBFswkPAj2ALHsi7WbHQjHvd3OYw6M0z/91USPzdse7/fo75OTMZbRQkRzpX2H2umhwb+p
4jQCxCp132co5uUwEWhbzrZW6ZIvnHvyyUPCym138VZGBFMkNAPqfrQnn/9BtsmvY6mPV5DdF5+a
0+knSuA0BWkK8O3rCJB44i5VgRJEcWkovipH3PLJoc2eAccGoh6aWyXER71KLzwYjmBofnnz8pM0
GmIjjlUJtgX0PiuXrQatPzeNjrcsRD+L9D+xv2UTS6CAPcQAL7LPWaNrtFWYJjQf2VVBN2lulRX4
tlvYw29vJL4tak0fydIBzD9fJ5ur0kdb830dRZssvCNIBtEiIY1WDsBQblhqmyv1X6dYfBSI8C4S
HS9PzuCBxIty3TiQWvTUXnheDYMPca5BR+tlBBuHxMXcxegJHuhNQkmWrpIMt7lHL4ioje/yZ18t
Ruu4ywJwWmF0qlqHOvX6E7hw92CHZsg2jEXKg6E67I3369nZpaBkIfKwnJ1otjGI6qMPGCA2icse
I6QtiOLohu3QDYU3ALMlEakV/SpgrDikukjjgEWjmDErky4Xb3PQTj8p0BJkEWZ+f4me/6OSh0a3
tdX2AIp+6xH5CTTdDdfpftYYWmj08IUYAiUUCgfGj3wTMbknvPaaIXwOQm3QKyb0ppiVrrFLxfad
v/Acj41RsY4T5+E/Qjkietpn7UA0OAEZQ3kdoEGGhDFg5yoehWN4HSvH6o5Y4fAjvUBfOmMcnLxw
rClIMXdC/C6FC2vL4vlBytqzVfNrANmPlqX1lBuS77SQFWSfFQRz7XP+oE+nWLgpNojEIiHxKAI2
AIZzolqf62Uh/8Tgbl+18nmxXNfRWCR32NcQ27aTosLhohmc/kL3XgMuwqjpXcMNl2IA+pwIk1Su
KvlxN0nx09jGIftcC7xOsuzaONvoJUdZpHXJNW+nXeORS8xjBemzimE0wZY5UYydGQA1cEjLg/xI
fchZMX6b39FuKuTcKLfH9+T0H0wpa8dtpNxLKcW4JYbehGxpwJ9BOkOV7oG9zp/3L5D0pgvKR6Hd
l2/Q4bog5j7HCywfHglyBgTfroBYm4AH39xv/Fn7fHavCS4D6ySbnk9yoG3KfxNCcpv3Y+GpmS+s
0gUW72X36mUKBsaYxw4diTPjU8giZTXzEUjhJkfayum/SPrMDh88/+RUdcA4yj0OIYr6Qmjb3lh1
rTwZkh4NbyRyzdBcbNc9Lt0u5Vc7xxeDz25oQtmPxoWklWyegYFkYyCdCObTH9udRPRxmzhuuDst
DLoHh+ObujHXKmnv2Fk8AJp/86r2wxfO5m7VTsIjOsi4vHiEMb0xsVNDNzmhdUzlQx3LaQTDXybn
S22h4RlFlnIH9i4sQ5jDdwGtiyce6s1TmJjkqQ1+AaapMlqhmiSx1j2kou1jMV+L/WRQdw5b0166
0qeUZuyyGMjZYOEaoXgP/VrdFhFHfFhFAg7xDPMAYgy3gXnTecWkI8rmxr7zosS53bbg4ohwCTf8
WV6wc4xWCAwdPQyyLEuXL9Fxxgs3mXmk00pPXSPV+3/y7N07ocSxk99kDnySEJJfkA7OKZxDGxwu
Qpwm9b2bkOsCrb9ts8cLB5wGCEX8s5GulplcQ5owX6EdRWXxx0SoJ8CaOnK3saxrBOnObARBKZfs
RwrEFyfFP+jPjDuVPGUbAnGGEymzEyDh2EW7+t5X/fXF3YBIfgjPpz+tiCzi65k+UjitkSG2j7/d
p/N/r9BAAJKPD/M/fukw/78sozhPduRPo2Af/LwgNMypD6sJ1Czf2PL/l73TT5dHHU+xvUWMRWy0
DFUKMQ5w2vD4K4qVtc8uE3N3MBZxO+9J+yJ9t2dkoAq7Z0FIiR+zSIfdhgSxozLi78ITjkXG+rvY
sgjFz0Es6EBasLI3NGGYp9XpitwA4vTH4uWcZAeKAQksR5g3sa6wtLc7PoljGznfqencz/sp3iYu
jOcNQPVvCjhwwfeXy+e8UOd/5yW5Coh790ornss8aK9xkOOLI6S16T/58GsocjMSMqbkOEUyPtyz
o9LZf6Ot1uSr//8sttuGKqOyzbCTG4mrGLGJQcOeLrOSIH3xL4wCN8a/lBsHaYuWwr7zLO7sq3C6
QsUcQiylbkYEepIUMF/kJt6Kp2PpQVxw+stjqPJ4FASD8WFLHRm8CSZRp6y8Dmky1LGr7mNrGWrZ
sznbUa7urQG1aRwikuledxolzdXfEgsoTB2IciycUKYuxKhl8vyc63ZTUrA/sAKbizIu81PU2BTw
7JsNgopu0atemwSe0+kPxXJxJLpzC3g407LFljhCNP+EyYOBcLWqDV3YvPchDF00Dv1Tmi1W3eBD
e2Ff1rxmqSoQ07g1sFrx9K7PqHwMlpDYL1bnels0qbiK6xLxvAAp9rukEickYJ5tPDYJ+d8QAHv8
gmVKLKU2kZjM+G0oxf5SXIDvT381Jdn4pXxzbcUiia61F0Yfhv+Yacck3v/1U99EAUiFSV6VMjPs
5ii2gEYglrDRN6TzAbkxYhEvSKU/HP7Xo90MUjXzTuyaNI6ZESls/Cct97vd87S5BZEYMSJ4YJFM
SDnwT3+YvQCewvOZL4p6JYWMECk9CT/iU3OT8x6S6Z3ov89EN6xB0Z0kfodwqLPN84rnkZH7QO+P
yTG3Rq+VOAhzAWStjSsgxqAyaKaS8QB03L6HJqtMwNf37B15GC+s5iyYOxuzV5cLKqAT5dJLL7JI
PK0E4FbT5qy1YqnryH+/Zf0Ffs6/prNxQDDSPRbXWF/DjMLy1iWdPx53kzIURbvGqJg2raD+X1Jl
AZcnLzlDdcGBJWd7OU0cC8rGim2UfdMiZ5xI+RFexNXMum/3NmAgEETuiRnLkVAJJZOefZW1fUjC
lZDzqZqPT1XG8RvU3UEmlS/Da6mGva+ukcEzNH0Woujkk6jfY70YfsFSNxjLZAuujULlxA3pdPMY
2LMc/LqpkBgzs1SXs+t9bmvr92yAtoGpDtg/DdCAroKa8V2P81Dk/1SKX2SxbVemHlUb1mlZaOoE
cIXsSO99AfCPuvEX/cCEksjRJXIz0zLw64nak3ITeGtqrFfe3DbdceO5KnBVKECP2TpQ6+b/g/N7
9g4dHI0lgCEkyg8VwB3NcRa3JH42CKezneROjkAsA42rvslgOOWHPycC0pN0L3E9ODfa7zoImkwq
BnIBYh6+G1+vx831zIisAeBqWEPWCWduB8W7wwOFuyzlQgFzsgwWKeBzwNHt6f+EMtccMhQl3RpO
YQTq8YSvu7SAORrlSseE5kj5vON1uZTlc31SBgzLlBnC0Mj4CYpyk+/Lfz9XYPP29CF1JSV7FVtl
SE6m9UkV2iM96HJRuJbTtwoZDFZ1o+3dhOCK6FxsmNOEVYaWZS5dUC3VcYhulUPcK+5t5zGWS/0h
eIEIB1haA5yZWYo3LfIjj4iTPHcnW5YDfifDbWG91UaYICL8A2G403OKnvJyyFOgyowBfspRJJHT
lZn7Sg1G/RtawP6JT9ODgbAnp+/AQM6o8RPNKM3ajv8TbznXXVPipaB/hycseysiy3fBip1i0555
JVifbrTlV++vyPPNmdIzN/yNKdZ52bR8mfZ+K6UVSqQ0c/KjivxJ8yJfsXA86ygxb22Cm4Mcysq0
iDOUOKOL5CuGjTcEHL9DiUG86uE97OplyrueJaYMR7p0miJR7P9K1mJKN/Qym7lfVP2Y8UVndLg4
hDx8/vlfHHsKNuMT98M5T8wvKp0CA3MezmJQLCuLKsdsXst3BEyH5zGwNyZCmaxmRSh20S6WwrnE
1cZlfwMS0UT4Gu2Wy/TPBtpqJB39CdL7Q0Ycu06PEQMg2ABV+T9mSSap2xz/MAREhg5oyX+Hg3wY
Z36nKK+4MRS1F5Nt4gu6e59srTzZoDWe6/T3Nu/hVlV+U8qhGD3Ss5YzuVZvk2m4Lb7OKu9OMBd6
+Iw8zMswFk8p/ROzKH4WcTnxQYVC5nibPTEKh/1Hkc9vmsImvofr86zM1nPcAKBWQI6Tu/cRWLtC
KG+fRwuUHrZniBgFN/ZPX8PdQqOo6gotaC7OdPaMbkdi1RuX3oMJsZoGE+fWMjzKG5cHJjfjeStk
I13HWrEbjLaF5wqcjc/nl+rLumIF4Av98MtCRQIMoIaj44at3BOhDFYgK+E9JGqxobx5f+D0LlhJ
mbaP1ZlRxMeWYkEgNDRwmqLFVWPsx3Vu3BnC3dbwhYsbqJip+pi040x3BKUG/cWOE0tO/zuoO36B
+GIjK9o590GmElw1bRkRvGgjLKQkJbEeMvBcbeOZaeGYyE8yvywb7vCuFFvV/oM+Fv97CIkxIqby
VEPJ1olHbuFNwBCtGa/eXqw/ADa95dIAreTWlIW8fQpjs+lcOI+AmOE8zLawrwpUKrzam/o0RLD9
FHs5fscLBkvh0mAA09fM79/68DWtpFef2clr5dOxWxQCQpVjOM8cr6MnjFp1xxo6ckveY0HKfSmm
th9YB8I4LaWSz1mKoq8k6DKe3NxOU9KB43W0p1S4fxh2hjkfgeNMf/wzXj+Xy/Wt77lnaXbTAHUa
mfA0e6qPQc9An0aJaEEX80cy3TBM1brf3oGn49eME2rpDGqxj4EvuTC6TlihpQop2SR6UH4xiPIY
QAzvNKPU71wx3BoEovGbsDf9yEt/Ox78r6h2azGNXN0/pUrBfu7AUlk5fsnWh04lEy1Nl0U4YLQt
RzTsYNFzcPB1/mxUseee+D9dYxJGCeIt3nxSwwndglaKoFdp+UvNBZbOSiF+qNAY0HbrRCegXris
dYsns9I55mXGj+eiG1nfCMmc53twQSDGhIsBo/o6i4f4TiQvMlfqTT4cPohnPY+2XZkgoWTd0+eH
WXJzaZ220lOg0v+FyrASFQqzTe5VCJK8MyJSQq8LVn9FSGjFDUe8EVCyq/1Vy68VwAtt+1jz/+sL
nePFkDqhX7ccPqagSxGpVAPnU+weaIdioVkMrA7zkHIqNIm90hR6ywsdmaJ8VlZbxDENUeRXhR3g
VXD1iO7s3ko/I9U81/NaTsDp3gXzhBePQTweaJat4nUaN0aojpNEHjsKbV1zoigXooVOwmIInc66
7yHrea2+GLTg7iWnrFJtrmONcH1N8XNCvyDIHqqLNStvdPNNWhBMKXP01SLnGo2Z61Jf6BVwhzx3
T7TSg3cxqM0n5zINnx7ZFdQa2imaf5eEC7RWkOaT6krQnAaRIEwnxGRbtSTfau/Ts6btueG7hR09
KD4svQ3y3y7FOUmpCbUdmcCXtHG65jqSc5QLwF1mRtLaBZmHiNQG/m54hSXR8jO1FthZqv7+Khlo
k4y1d2fiY7eRXVW8/dkO7Nnd6UoK+DYILOUAhq6rSeRdmpobR4SHNsmVxtf9KsDwO10sqNuDTXPi
3uM4BtUZBkd5EDIYYw4tNhU3WLtfQBXuIJAjFuIR0GtQ/fu3lk/db7I+p5gg52wtsM62Y7M7cNe7
nu2hLggQ76AIJvDjs9VySKpP/MH8bls4IkkS9gwx99xIIthsL3KAfdwObh3jCBg+NOsKcWuSrmUf
0SsP3Egh2qRJx1GD7r5s9hw/GNWJrj25/88EmqDePBYdeJAcAY+bpX11fgynaIzEKQT4a6fMf0UV
LrysfHw0Zbq6ilii2Eg4Sxt7bEv3h0wZN/s/JJR107z3LWqjJx3i9R1HjhtEayaRGo2bIryLzCRq
s7QZgNFnEDCBmw3ccqbQwi/hTfVHKs6yIobHHmiE+wYmBcfjnxGWlA4g5K5CUGyqwpVx9a8Mebo6
dduYGmbZqQDdgr4pT7SgnSnfyZDo7MsEeI9dKjzy1NS6O9tX8MoYM9T/gfYzvLpYCWWtz+COOhVy
x9QA+WeA9B3Z5FWGG9RZZMlcIue6GBm1gmUWjxrLQ0sdYcd+A96PlUg7cuFC0+i+20PUijU1FXLL
V71wWWgUNKYAIVaSPC7+R2AArJlbEwMZFLH/rPABjqoNJh+8LeIylcbqfXRhH4jcovWXl+UsNZ9T
2PIAIq2rT+cjCzmfQKLHlCiNPjje9VtDLJRdCn+9bWc5szaGMtaXnzQ9alpZbl3BAmrm46XrDv+/
b7DXtSj5ZYQpc6/arF6SrQBi9dnKxo4w3I+EZaG4yRSAfrrBaB/HKKRbCmKmJJtiKNlbhtQKjqfb
hJv5U9ZRZwm1O5ge21JfW0SOqSYoHyQcVoFhIXtS0eVeoZpLd/HAjlJqMaQcKEm0Zp3rTq6ZdylR
yLKrLEeXXh5A0lcbT6G7f36rHw8aEeb7CdxWFCJQQ8hRzElo0CxceP1EjA9bAyk8qv5Fme5wQvvI
bpAgbS5Ab3Pt24fW+M00Z9muykCviSyhY4ZrtH/m4KtGZGAavlIV3JfCt1Neq/60MHqfHWyrZ4Zu
TDmXIaIQn/oguw3qneL/IEU0Kk2n6rjIZBbZmd4ICkTsElukQyx0NMasuHJkkYSDJvwreh/tybKj
ZRlnOuUizo/lNn3lOCDFg7EaxowNsnf/DdYnD1qGbdrGrcZQzxQ+mhdA5nFpyK68zAJdD17JjV7U
OvAj0pwcYcTLPVZtnnSy6pcsjR9VCmvxXI/vXfQLzDZCPQXmWDfNjs4e9AI6gm2Q2DLe92O0qWvN
NZZ+6TcF+DuDlSnK/Agma0sICQwge1nma7t9drA70ovUbYZxHNsKOXZ7RnmdrQExBRObxc9f0fNq
DbF0WmfydTF30wW+pIwiRSbxnlIDpevWWZXmk4EcoGWySm/jrtrM9G1miKRnjWsE26HrPkcU+7od
/H3LTS1q1vEciswcDgZ3e72ZaT7JnH8uesyKjW94fHBvWaz+/ZwhRkJEfYPu3huoLW437ZSgVrLC
qnUU/wggTYMBSPA/0i2Fs7ubph8Gf57WDQJyM16PFxiaDU4t5LhKrsaPCAxWjQuyO8GO60cSkIw9
/QlnArd5AG5f5vbvAvoHLWXOGMN0y/a8kPyRAPwDYuwev8ifJiG9IujXpVKvErad6+rM921lHidF
quaZcdjJ9QqHbj2Vd4CbFlbfSgJWytSCExUJpPbtGCAGekvYDQT5NhNOVmlSvPmMNPxlYFf/MUsq
362HthD3ULazxTQE0rHFqBQAwfpf0yiYjhev7bblWIp8om5X68+iYvK0qomiGnINdJSxOJ7ShM0V
gjdGPazb36HhEWVCtCUzgByGothUGKopcJ9nflts576MSkmhxGeg5lcV0Iwe8RlA8FHydOKzmAoE
1WQpFElaZ87SiS1yokmoTpp2+2hvmDbVM6x9FzS3szsoNKDJ01O1nQL7Wi2pRhxpN1PVmPhKuJd/
zhgNgDEJQbmLpkqKxY7Xe2PPiYl7dFyPNap2m7oAmy0bJCD4LvK6Lj731+V1GVnvuYO3toC1Rbh6
8iedR2cl1H3Pp52cOVfoTKsJhY/6ZGbp0Uov7rQXRcRIju++l59EciaBf9GpgnwbHr4cJKCKldEe
pv1MpM9bZ4M5G0L5zc8m/ED7Pk2pjR7J8RlsIEFRoHce2yo7806v+8kV2stvb0ou1UsyeGu31KvT
Nsnif1u9HTlYNNa7qxL/g5CRMHuWtc+1op3wlDx2GFrscBXTVHkILPaynAZNAAVqiHKBqaZwrmZQ
NpMRP22VIYI+KJKyN2wzCLV3bYeb2MATGC/cT0q4eMhvagWwdezUfSuHheP1vgHRvkjjUcfOUAfl
iS+G0clI5MK+fSoBqJ9bu6OPWi0GxyILdAyO1dxh66008yhscmyxgVXc2czl2Ibe23yCU7uXezdf
ob2gRy2rhFAXC6e7H6FiL7gpu+FYCpvOTsEMQ4qINh3N3fxkZfB+jRlYnVo5juiG0lDHPuKTHJOP
llmTvXifSwsgCJa63cDypNas8frzsFfNmqde/FhjhintkYlsqbX2W5zP5RmTAOM3AoDX/jRaEz/3
yb+oAOjZG8nATs2xqJD986B7bt7yNxhmDXl4vMrQOVeJtlUGQjFMd4/8myH6flqODqnSUPSdMVAE
4YZINwU44gFl39AubD1kKNCYbDAuyCmbTKjXHQmFSO1qYEbT+p44a7tg/b7lQeaw/RbF+eCuKwmS
wpnZSWm/c/9PnhrZeqGNpVbuufO4hwkwUzccgckMQsK7qh7INMK2/qLXSWLdagQua0IpA0rpyCn/
U2NY9vGnvmHZSLjA+PSiSEqjqKJCtgZlK1uL3cNBEsCuwoMS6PM9wApQ9dp4qanfWKarmS1srZLK
K1lD4H7a1I47KJfg3XBdUiyo3Fej9XdXPpkS0pBv8YrNN8FMAwCt2edF2NDpr7+Crgff//SydMMX
5SEHawlIVZDvDv5gLgcxvoIg2cxRn+GSRFcJNlfQd+qYTNOSskxH0zdfWVFFCC/p6GwMEuAkQKaC
ZlNxLhvp2/6BF+g/YmGtP/NfJsfbg8B821zIfVktsJiznKafcspHoeb5BtawKzr66d0p7J7LEtnE
pzdkC+T/CbbbXZSW6NjSBWqsCnmtoAemQETDuSdpynDc0nEpN7gMqR83wNqh1CR0HKDans+jjPVU
GYp6goTzrQrEXw6gaWxQiVZw4/y60B+hKeJgXdygnaHBroB5B2L4tiswtf0SdkjfGKgHOO4v39cP
OY4A1QJ9EvUgKp6k8t6Lia7VVji0TGWp+YIYGXMPewK+vqDz9W/RlJqDX8s/saMp/ndn0MydZMZ4
yLYjvV4KHvlUoB0YXVMM4YWE5rvzzuAZDNT92usnU9WFJQY2xHY0TTSwGIE/YLr1Ty2JbKqcQ18m
aM/12H0qYR9mHlujy6O5IazjAJ4fO/UupCbWw5Gvbqz28+MIUieThiGFHG7+BDig4dcnYbzJXwMS
GYWeh7aPAmRxJ/CuJQNGDZ4LBJgybOcV9IzY3/XKnT62fhxjOI+jzTKOX7l5urz8cz6eNx8k69M7
TosvWruKhHtbUGNtLLz71h58RuDz+hE8KzgNa6KZ/+bim+X831KECLCw4TFlQZLggv6vpaU7anow
rt/2ZIrsz/wqVKaLRt6/QGQ5iEJL2qmULIRK2LwiAXgQUlhOMCdQIen//iFQamRlet5ECi4ARg13
r7FxK3h+UpMH9qKxxcoweINPTx2UoL3TNQl9YqxExCd8WJ5/zGz8oD24c/wEwAom6PpzdUgCavoI
t9t5HxaSg6R2cmm1CHB5v1lD9GYP+ZG+F519zq82gsbeJq/CK1ilC0J73GS0LRcAeutUrHDMeh+K
iDM3+ehx3FUHScN9Fy000GYWQ4XrZzTCer5aiBkC81CI4dXCp87Xb0jatif7Pj6m4qmZkHyYoRIO
/+TrVr8X97R/oO4e4vHNumQtA4ofWPYW35DWJHzJO2f8qV6W/4qKkf1arrzGp2vyzZQw7KY2jeNe
4txPCwXunXE3F2LwGeOW8iTLTXMMgmFMQSDZzw4qylscazrQ3Si1y9sbxWhrTGy+n0q5AgECyq+V
MoDg1SjqhptK1IcuQ1cIkKSvQb2g8yIbn+SEhmC/4ExjTICAdUGW2inrCm2jGGR1KsnDGFQRqD5z
ond7w3M96+QFhsFUg6rda9JSMnb8HeubY+r5fgIoffic8IFdSWgt085SgCPK49PR+Is1q/h1+UVS
KBJyqikJGaHVsmueCKxnxzQHhvdkeiaPaBTbPEmSe0HmIC5pqvxqbsh72VmM7DyWcrRSOxYEGfUB
Z9qS+ZV8I7NzFDMjMhUxszlZGt3eYSjgctm2lA6EKoqX6XdxB/JECagilopng4FLZOTW56xJLaro
pJIo7Imzd8TMQjnIV+YC2KcbGa3qPU6wXI84Vs4KC2xvnctwLwkFuNrvS2awKTTevv0z8+0fQOCq
yLNxb4ocpyreAmhaU+cmJDvc/o0m/FDXfSdoWQs0QTw6mg13INCPEA/s+hZMkQtf3Z9xfqIas6TN
9DdV5bLoba2+bzFLn214xseCWZ34G04wgtQuIHgSJE/YA0gKQXaqpKyeLlPtdmaD57VLZNFYrILw
HkYczHq1iFnHyI0H7YCh2cvbPAf89HT7PzeEJfjEmSohJW4QRyGxL+RUjtGNKqLG4SwzdcLs4SER
trCFpZs0SAaFg1Jk7Tmf9RLnO3uIOC3o69ukXoh0SaoKysdpC9NFyp8pBf+1+ItcZ5xCGVl5C+H1
NvyNw6VM9VguyyO0RCP1es9Qmc+PD8uA2IzbfUd5bw7iJB3gyVctINmvzdOvQCCvDaqFhjwc6HdD
KeTSO8zXXve9vy3dNi9X+ACKenpT5Xsyc8ttl8n6kD75acKKVGnsEKRnMHDOW0lmeyEKZ4RQOXRq
EHY5rbACIr4lXrElP8e71l2GsmZse7YT2iVixaE3JMtBpoJwyGU7PwtgERnwcTqstiOFI3CSOjMl
Cj9uKEKOCPAdb2YjRuUD/3npO5n+gGABWpPXOpdndk9mMj0zyG9Db+2Wr1xrtwBUjYHnNxuiR3xC
zlZ3ORFk6XhaWw9tPEI+VqbzZOTd45AaEXEoYGXH6B5tHbc9twvDHOpPOvFsKPAiU4x96HJ1g7FC
7CcPaUfIlJOPlvjgmvYWOtOpWlGWJAOtA2LCeS7Cb50WUlOlgHzPikhhbna4eqP+LZSlvIaoRwLm
8dPyXkBDmcXX4NEFSbCXG+WgdyT53izYzmlJz5KJACb/rKU3UMCnDfbc2Pf088khFka3DBFaOK3M
QF7qriWj72TaFtgod6T8f1TVhvoarbvOmFVCKLOo2ON6+dodScviB5KdrYC7/1sHn48EHI1G4qsv
v9n5qVHcQApDnFnoS0TSTGeZ1ecsrMXmstVENDayTmXmn4L9QHrhIny9YSimSYGWdnKWG4PxuUKX
HbfmXwehnutOQdoJuzQ/7u/mkwyjGQ+yLw9ueiBc9Cw0mU0KWEORB6aDy65YzqLI3y+ytorIo2kQ
6eoK7dh/z40z4HEtS6JQBXw0vQ/ermc43jIz9fxt03hKkvpFZMhZGmC7F2boknuext1ZpU7G3j/7
1vv0pZStSRNqio898SMwQOmmHir85qt+3KiT9r+TvW/M0a3JdFAyOTaTA3QWIg5nA/rvoFPVFfz5
fu3TEvj77LU31u6d/O+NR6Sx3ffA6vwfpw0Pv4iOeNbkJz3yyPizidR15qPcyFzQ2KGOdtHePJyd
vy/sPIua8qEIvc68TWt8o3irec7Aquvb/YQRJxVs/vgrIeZihX24qFHreOXAHP2XsyCe8y3CF/gD
vrpnMZTkpic5HJ+ArhCyn1O7LTtueDR7EYDIodcuQBb97DAi3BFy9aWHav+6v7XoylnEERhdqs4v
CMks66m6iNfkFivhSypG5pOn4tnMSzMW8B1+aJ9V+v7RR9a2Q4y+0mLp83Hd4HhUHsvaoH+J5Eub
y/+EWGS3/eejhewU0l2/kRRGkpiJ2VFFVVDqKTfpraBruX/A9TCz4ZKBz2V176fYwKHaMYnCCgaJ
evw4J41H0mkGV0MVGJFAeMdBqCqi7hXXP7CIjQ9jkCpZJZplByWJPoJlUWGxPi5YHZW1VUH7lvxR
Hk9PlQ4db+rHM8b4I+Sd0tOsRx+fPDqS+If2XZTC0cGfEWyj5XPHDVd1a44KjhKM2nMEp+it4Rad
BdV7noI+DJDwB2izCcwNPZorzJ0W/H1bTskDq6yeC8bjNN7LEE5uBP6jvUpc7FCv/EbIE5WN1wg4
fd+A8KLxbg1EY8ty8WMAnEQSLV0WzGqGp5yW8nIpOVDL7vYLJlgcaZugNK8XB9yOxVu2+mUn8H09
jeIqo30GsjPi7DWyMHop2nTuKuBVOxUmD/DxtrBvKf+R0IrMM0hYb/HC+SXVlcS/y+iIWiWlUEB4
UcYRi7ruQ/ZCszfy+/TO3bohvKnD2/uaXPuvCRwbuCrDVFf+1MWsH9ylGf9O12Gb7hCNVChTkTS4
hlGTJ1oMIGfkniPnrT3/zr+rMI+6igI3WybUH9kBOjVYu9poyqgpVunv0MGPjF156G0/0R3CrNEo
VgXXxO4tvgkjNcz7o1mXpMAKXOkfJ5zejU6XNnaTpguwi+emIx3MLkYmN+LucnvCXlhxY9NUKmDo
lFzT8B3KCJTkZjIG0DnJHeZFlORJg9R9ayA2ckVvSSlZXn8KAJ11C+s2sqDRLsvaxf0Swx7t/XNx
a3CGQvbqBUjFCNGuyEHuUaf5wxJCNq7PnMxLdakvOpuVn1ea7RanOFyWqPoWF44QLX+8V1TKjPT6
NRpCYsEMJjNkeCjP26yJzBYGwgK+sycy9xKscc4aGMdqUPi/ptxsfe4Pcb4igx9ffn7WSgNQPU39
L/++/Wlz/QgVoWHrnWL5drJljUva15TI4qTwIOGv3/Awx6X0sHEtUMh+DpF3510uG2fbQ80n2D38
JPQiYCsFz5wg4YRjKb4KGo5oOzptJ441XLSrOI+YU7YesgSjZNItGBeNRWsTJSe2l0CvKaip9OEC
CeVrDySaCnmC/Oqvznv8ymvP3TL4QPEbioNFdrtnO/sF2BhzuWFpDSsuA3Zke4rSHOw+KeY77kN9
a1neu/cTE9kJYPaooUBDgaVexooOKJnppivv9Qj4oDPBKuTOb+mZ7G4Y//Ks5xon86Fc+Tvifbch
M/R7ZPsApuT82WqEmP07vtmAppj0554iBogBTVCUnAqpGbRH8qacj8Dj/LlVJ+S1OOtZwYc+kpAy
hRy83TI8FzSkvBP0jzTFLT4q395qYLRoyHzTFAGdsh5uxiKBnndI+AYBIgv6WoV6ck3QKxvycii7
jS5uYjyDgkTWuKk/4v09XMC9PPbKR/2odHGydnOcFcR2NxAjPwfCciR7KsQQ7hnGXxYsVuR/ndlh
8HExjApA7nFUk9BEbFINlBGI4ec+iCmkAYmvuuepvetDjT0GiReUBWlN/8B+PBtJppaVazZKb/me
sJSdelIPnMrzvl3JtQ4TQy4oxH/30OUb8zf/vB/OjbZA+BM7BXI18kCRKuqYQgjqhR+7dIC41kIg
UHmv3hPqbXHGheY5Qk/D0Ing22PjP4HSnkr7UL+Ms0VYD2TFfAYvapd88O1Ns8pC5LYE7jaLR63q
8GCtS8OZqHbheBHc8Yf9SF5ERhmTAJBtj0YsB7KoUaYdXfToE6/eBE79LKCgncU9RevVeC61vCsy
9tvESf2FkQ7JhVcdOiuMgaKSvsrP1wEFXHRTnI+HlL09BEemhgmQMVBSTTHQTlBTv/MD6A/0cikZ
GnviOgPVDkTgUF1b8om61X0gsLDvRbe2tniPoxxM1v9YY7AJ+2j4OCIWclwapSuCdc9wkcxun++f
r0KgCpmrpVbuBHeU2akqoMplaBOnzlmBLsmvtsVVmM35bWERlkTPn29WvDI/z1hPRULiD7pTu4HV
z0Ef15a/SD6Euy/Ct23PYPaPXsfSOpoumxyx2b9THPql034ya+m4lFmEOS1mjgI6MwSeE4mkFYiT
fpcWFl7MCHWiITZjFKTQKf7INGeelcCbCtAEFz9EWNfSxX6kBK+OLvjTlBIlVt0DQ3mx5MchNWzK
NK9AzD3Pb2AqwZkdos0YDQqI9uD5IFbKI4Sv6Y6eJtLmxCLsfG9m0IWGgO59YSw42aXy28IUPQxw
neBT0p5wmdNItZPosrl5B58RtADTFQC7qP2Ulna8l2NnK4u0SrAYXIXkgK2JvXqUivMsxIMsdj6U
Rc2J5iArOya10tM4riCepPPAInYzxpzRznRbO62wVkMj8cANCrkTJlUbEhxYG+Yqsgh0393ceTeu
FyzP5EtMcad0oFFiUuJLUy1oWkFDQNma74eP4jfQkU9LPwiy28fIqrkRN63D56p020w144KWBOST
sZDX7uSRWVrUCA4BoNiqeAZpqzpcZ/9YsrImkSOdOiT7i3YWimDSeVMRBRtUijkzIX546od0WQ4J
sc1agaKwS0H+oelfYdNiXo7FZvuuTd1ud7RkooC50zdBwsCS9XYh+JqsJ2wM6OLdFbO9ZXNZ04P5
CecWqMDa7aLkNbaMdEHGdUA6yebuxRMp7uMkaA+bt7hlOTWAKBZx1kT2heH3GrAxatMXjnJQqF6o
KENHxIVYeE5IfalWaPBhq/X9V3kPt1/17H0NiiQBOLkWNBGf283mWBw9K+u2IEWLQrsv+s3J9qRc
/hte3qrATEGB8HMKdwwiDoeITUdqwJvAacZXc29nSsvohIHTgJu6T53cJcZHHSGvrgC/8ZcVh5Gv
BMQKauUxjU8g6s8YehD+uEnMuNdxVtzZ98HySgU0Dgc+lmoO6zJI3mkx0iPCk6yw+MPHCcZm0rRg
R9LBOEJzEXOtJCjwBRLtURGgBv6jSU6TTMi3NqCOvx1hXBX7OQMIvumFAF7zBh6fdf5V2yn7VLkA
pHmB2R1Jt07MijH0fuT6Ypm6jkODky4htm0ODuFxBms7k+gegCK/giihnbwpZcHVOyCWX7TjkVC0
yxByjU94c29+qVtEXr1MDipKyzstjKEOBVA+2X7RChso/ZiL36EcjMPhxli3k0/T6q84YsUBHKKB
84U56kLNik1ntC4R9mYpKfUp/aANqqCrTXnhknqrBOn7v4/qyV4hYXPMyF4tk8hCjGkrGsaRRroc
FalYhKWhwQB27vFr4AldSmGxKBYSgwMta5RUPr4QrZDQlEciWPOTbiXcnJ1wvdVGXlTdyVscfrKn
S5zVo+b6/APmgdVmdF7LKLVG3LUe1H7EH1I3m4BzXRoDhc+3vsiRD3JC/HyM3NDXn566XxVZ5iDl
yEGWpT4r1ORTiwWf20cq1awwLeJwFTlu6DCQgh/UgWaBe+OpFVOLmeLg2rk2a3TWe4QwceNVouVI
xWXWzBfo6Lw3DSnIFtr6KjyWfN65/2MFDYFJ4eC9XeM8sxW0blhwABEtu+QK1SWUxs/bKi3LQ5hL
0/NZCZHo0j20pai2FbuFmkSyUZz/Qe5WCawPCudIsiKGizGAdZ0Hh0Lz9BJc2Z6LDzWKGyCegws1
ZAZWu/y8vMEyO6ME7jcVLU/yiS4vQYQagn6kvVk1tFBFLd7TTKPxluiKR8D+0f+u7O3TfOlRBdbw
6JV8hjCmTZynYlA5c2a4jm2u9lmcgcQlZrSGiYqBMJeLEx0GhZ30ZYj/eHpKFQK+qZdXwO2SEBNX
MbZRBdvsaKCoCXECM5K2SYduYyswdt5VynOzKdUQXn2lUgqj3hJgHNX6XmOuFYqn6dqkXIJR3tXW
J8D2sFIrnTJsPWCBSNJxwS20t/twAUxtoYDzE0BkFOSxJvoiZj2soDdvbfzWyFKsTGYAqStATYqB
RGzcNS8gratrFpukZ9YZHvzoE4UH/qXmAVRqPwPyxLvaPDxeUI3ho0rJMHxFU5CH8cANmj8ND+L0
f2ElrM4RCpESd/+AVnrRX30K0eij0EXB2ovjqlLCvz3+eDOm1SD0L857/nI0NHtYmrKeLWPZuTXY
myATcW/vf1lmTox+COHwMSP77wUdc0wmE/IaAvoSMfb/dyzGxND80H/ZJEb0tK/7GrVVND+i4YHF
/LHaSisR+smDtuHyBVzpTVbGXbIMPfGb5dT7vIEXqEwElwty2fqlt3NhuynyY1FvueM/4JPpCcZv
6rEHGizXJfI+SGR7+1g5Dw7MmtKZmg8uiUfO5kXNObHuY9vzt8StRKhLsnI6JlsMC4PL0Rh7lrrT
/wUQvknRHVazTZAdNskBiX6de7QxdTTVOBOovCG5jAUzSpQv360euoYPzpZzrraAAN5TqktnSTSe
pBA2eb+3H7e90jDsYED5fS8vks+enJVd9oFQhx9Ia1gy2n6x+hebIa20ggI4A2KryGsCjpgOSifj
peri0NDtN69EBp/2cbgeFtNJaVdhWopQT130tMej1WpJwSPC6SYZW/s9cDgrS6u9C8Ln+gi4Lnwv
WE29MxLkQ1OZf4gTQUJ1KaoS7D9L98wJQrco51rwY50b6sXjpn2wf4myslHjbgEDOeeX2hYQ+zfM
tXjPs3cbCGmd0VPXvxGSM7Ef6j56IxBDDTYm/My02qRSihSWt0YxS8pYo6fMK3PVynGQENP8TXQX
AVeqxTG2yqxLzqMKiYcjCK+hVnvQ59f1NqSd4gyvRsrTWzSxrfSGjjwLQnhu/JWiE/8RUKEreqj1
7fD3oLsFFkzlQDz1ghynrGXfSuMAnAsvFU3g5LICF0c2qdFTgHgGrZa/mJKvdYsHWLszbSrsr9ew
Co/i6Mh/L/j76qvOizaCzc7RTvbjNJnqc1F9oGp+c8g2kauqY85Uf+v9vqwUell+CF+tJlW2nC7y
MLqz5Y7SZr/53L6KtbQ6B0EF8vR9zOtK2NIhXxEY3ag34T/6JMJ5cIPtyxcQ1HybHbxxf+zLEDqt
qUdQzOVpmLzahZm0mUnFRFjXiZ+5VYLLuCwgYlC3EKqfhTv8PcGQXWe5hIiOqbWypPhKWIzvZPGF
UaDRrIjynW1UazMiR5y08Y8OYTna0kmPd2E59529u11cP3nKHvpRLcn7IXRDj2wbomq5SMLD+ihk
W1ys4BfU4sO0PILJMVtwiqFxUkzWI04c5ZaAr9Jrrv1w4HaS7xTWSkxL5q9HwednwKtXi6b/N5k6
MfTpRdCUx+2GPZ8oVA7571jggaIv/Nlmpczi/IOrmLWerx640+fj4lCOwVqv30+hYXvaKzwOzj20
ClvmmcbdW71X5FcJ1kq7lQswQ/XeumKEACXT+fRkwu7/kFFZd9P+16eaH3dOeL5xlHe2s93hO5Qk
kMNk5C/W2mLDarWFit5G0/xkigfIqrjy2U2HhPBvUMLobkRHddVvKPuNSJW93WLJXZqwwOMDafgP
oDcmIZ97aa3pHwr8HVVHrLUul/G+sD85Mppz2nlK9sbshwa1xgRfoBHIBWE61mkgyE8Vl9tS5zAp
lERIM9I9UF+dqBzCJPT8t2n60bGtB3mdYPZTsXzl01Xa6CI4SEFtR+nLFlq+f9J1obMkfaBdv1m0
etf8COJi/kp3t2eKfIfGlj6Qmjy9DZzJOfD8ceXbObWnq4BdJjjQXoqbKOZj0MRCi5ijtUmoxD6K
nSZ1bcnYRcoDw/hHcmW3qVDt81FqKsxvC//QRnC6j5gySL82VJfASniF4AbtrHEcFNkz733f7sK8
mlvag6fmXEKpOxNNlWmrAO96PiEVTaHLV/XVEIo5Jv3SCbPt9t/coqVKUNlFo2RtHolI8oE5jurT
oAKFei/99oJCJ3oT5vGBP5AWU1kyETakahlp5GeenALi+hKyOsfIvJqIeRDrkZisFn1yH8v2tX32
2Df+G8RY2idvl9pIjweRl8UknGq1cvTmdSj/7LBJHXJ4tU1O/9qjTgS2RlhFcDfhSbLXIsOqCobE
8aLmvKBHcdgdk4ThH7w7XuVRvJDUKZMAJA13o22N+UlDny5zKzuSmn3YruL61EapZZlCSCzIVs2d
hGvDQsK/0QXKIk4tPejMVr3a+ApxKMMrF9s5EOtzcaDoHZdV9/SAVft/mfkmwSbQ0x7+NIhcCM1a
DK+hFswQBJl290cQNx41Uqd/pJwVwy93jC5YU2/GZlsq83z0kWWXAGjb+mEL066Jpx6bVMK8/EI7
UIs+SXvLR3sBf4CpgHdxzhcYs1fZoOtZ/ZUMfvd6Y6UIkFG02iNez5zKqJtS9oU0WZZCQpd0yfAQ
rzn+nCDVMcs7QXfpA1aQo9sdxF4zjtlVs1IQXEOWm5oLOJVLXlSErm/Zc7I7kdPhY4SyqPTacv0E
ZNIPLWVUX1pwwEkfvTdsoJ+gKyhqb4idkN9hgKxhr0ustQ6mxYeWBZPvwF5OSUGZNlpQ88oXKQKt
0Dfl3VTwQVo+TNE/2klYZWDpqLAvLniI6muoXf8f1yKFLoDOBQW69787pXzdZoxDrY8SEzk6zQmr
eQuXVLEUQHWUO55+kutmpVb96Y8hxyV3mQkhbSQw68PgHnpz+SMTEEhO71M0+PAOuaqHRaulpK91
18Z/vX0HmcQISv3iZrnbfEmv1tH+4KICEs2DT3tScoPc3SDx0H7XLDmmX3ToG82qtkX0sUgnDB4W
mTFdy/4z9wqUi9RscZDvN36U7Mrg0Ro8yvsACBBkezxfyvmpYm8HX4e4IiUoZxudot4/jdo34ITt
yIou3F8QtJho98MPOCDC8D6JKjo8TDAS3FqOqHrLFyEHVZojv93AYGkBlpxHIGs1gFo5grbIGtD2
wjnME+ptsM0zfyZAfPcPJjPtCTlSFtdfIEsU7vTyvFaIOMicXxtSqPsXnyXXv4bZ1WB/D1vbi6B4
MccAL/6J3Rd4u9/HvB6X1ogSmVvFQqmbwRBKx/WPGC4Xzw+3386i/3BgUj1chpvShRv4HRnyFxzQ
Jj5z5STnLjisxj2q46/4d1TzXCYWj2JOZmy2ljphwBu3w81jDak8xXBRA+p4Xd024s4ln1AqNyOt
rf52ESipH9MyI1d7vCSWn/BqcwyDq9lDKXQVnj8MHgzN7wPp928aSix6rMDIVsAq+iqN9/Ij/Pv5
XT4Y4lV+9fZSokVAyWQrqZZipm5H1qAYW74ofZgRjrVfT0DhOK9PY1Gp9a2MlVKmLO92DMJ95L7Q
PyCTTv0oyRAjGBxCI9km8sc7WqamXUVuZy6yb+ZhBtmAtgfDulRTpmr66ZSQwk4DYO618zYB5tVB
dNOY2Pc3LBu6ayn+rgyDUxUNPN3rgdCaRoHcvoRs+g+TKL5e2ehPgFxzgkY3QtlXuwxTQxrlj7AA
yRzVjpkTqQIIeizx24b3r6qPIgulE6YqI2oKw9DMRVIwRbMITol7916WPJ/1Q0QiLd9WE3q60JPE
rJlkbqRnb4E2ZR7SWHrnXjkk1COmopdfyF34I4k7h5pg8WkK2jaaMKGi9jOP4Iq4BG/S8efSUuvO
ClKPN0GMoMqrG8ejwFEfTC3vV8I26+TbayxjqZfgfBSLg+DHz+cjAnFnY3lN8NyubdZ5ArYQOLhz
cXDe5A645DFZgohhlN9yBuOVJq3JqwpokM1sdvZtsLE0GawMxaJfulABs2uqcMHL0ejuJLNbgrgs
rs44uTDNVYW/vcxsIgZgyOgLQITA618ojUIbB4dYiVzsJNrMde1A7EDuCs+N+RS+ah+SL9hQhtVT
dEvaNwINOO821PRFQECW0oQJhxFYpRtLmbtI9GCiJj3M3T+xT7KWpAJ8R1nmusglDUP/MrPWTaRm
Wq8tRscYHryuXHkvk5koIVdfnRAl5OB1CgfdMauyy4q2uB4Lz/CGQg690qybjxSwescW/E2DeNu4
P7WgJAbtmYCROJP2zai2N9HorR99p+oLY2Y0a38r+V4HGZmN0L58FGA/rbChpluKFGB8YOguON+V
BP9YIPiDjgsD0VgQKLCqmakWkDvqxYQRMrIB16l+4zANSmPw7IoEG39ZolMLnoazj1G5io5NY1Em
7/eAW3OQ9jHG7H1/awQ7kbs5Sh76yBgbLoeknjNJ4D3xtc8067q1YH+BYA98iBnCmsKulutqXEEZ
Jgr+A1DYyT9TJt69lqu1U7T8vtqTzszSSNtWM5Eet39kaZJPB8I3XkIlDuyelJZsCPTL6DPq5+tr
52jfKGM1c0Yil+CDOIK1hgobxDDg+1r7r1aq/dAmbJ2xp+zinYoBxOYzKjQImT459ghejSsry1RL
rDyAwJK48fBXzYqR/gZjO5IMf9Lfb97SZr6KWCTV3bIO8pDkQbrKmZ8bJVXRqhzDf5BqkjGDhN/O
QAFUFEN6KVT+Vg9tRCYhpykxE7cNf0KpYPiUFTSagNpCm85uoxNSeTYA1MLCMMyfLOqMkyLwiniq
+wfPMIjW3y75GIiYenyZi5VFfZeJMYgltqq+CUcZOTfngA70KXFAbeiD58xp9+cIu94VMfflTa27
B8jqiQeLl/R/xaRML1+M/NtRLyx7C7l0RTHEU9DdOTYVdpFWg5uPDRFIsibbIb8ZJKPlvQjbR32Y
pl7QyqLiLAEVz3YeK/l0YV26FssqRMs0KAY8AEvL0xSWFU+AcKdfek0VWY49GRzf629JpVwH+MvN
DRRoIUJf6FGviehDUUE8PhlYSc7lyZ8rF03Hd2pboOnjvNwEJAuHwDeVwv+URm5CpA7zWT4ej3Iw
COyDQfD+yVntb0LJGgk2yQN/Xy+/5RxA/S7xamirhz/AaByyUr+nbKrxEay9jFDsysznmPwHXFEk
/z7KI8UyTO6GPPUijCyexXaoIc/gu/VU12Z1Hj6D0gRPJUABNpRDqDQFjqzWSWR8QFmQTcqzQhYy
EtkKcId+RuGIm0vU+BBBUvNQ3XbT4dVdt4HasySOy3gOYQkrydWK1sU47q9eu3Va63I8q/ch+TDX
XwpAqIQuBgE/Xfx30pMaQ/h9F9azGastyYeJx9khBrRGSTPx/i/+jywngNuSXEvLD5x7rrGk+kqq
/GBFbmPbZz4AkJkcc97wqBPoOOGj8QjfGmS6zf2MfFZ8j9nXOH74TWpT3i3ygxVf6mvNxO3BY+ur
XfgrY4+sZRz/ukDb/uhUlE/0Bk+2jvU7K7RrtVDdCya/Lj3vapfl6SFuEnQWnDhdUh0vumDRJRRd
dr+l0DEiGYVFe+7xVwoebhTXf1j4M7OhV/u8dCy+/dPfKWoHqW25o7oAqzfM+/2tS39DGgzKfhWB
22qfZGBpJjXKwANKywdKGIYw0cHfjugEU80JEYzwypLTlLmzLDNgwUmSTxdCBPvmAytGpnZWVydf
FnK4w9gwgXFUDRtJLXk73XNdPb/Mq08dmIOd+1UR+anSOETO3nLP081iWeObSph31OcZJjWuHebM
oZmr8P+o5k7ydQVxtXd3Qo6OrR6ACZuxoY1qWqzNLPfwstyDQ/YoacwCg7ytGs6/Jbqev6Ngbdea
rckHlS5UJmZsjAxSpDiavNh0L9hmtPYLTWgztORBzrGm8wNf1e6YIJaYyG/Rw+AANkep3IfyuYwV
raFslPxvWeoUuvdhhTBkv7JRxBEOGrXs8UeQq4LMT1Qun51rTtzBt64NcgR0jvfl9Dh6r1M/9zsp
7Aul1JfqcA+Ms8NDoNoeimz3euvDXg0uFfpfWpyuU7TB3hmeXWuGoYeMsOzqkXoMyHV3phDE5L8n
+KooyDcxGircPLVA9zJSW41gsp1r5sZNkWQSK7qUydLt9+Ry9h4E+zrIj0zkEqF0DctTZRu3yyml
HaxJqv6py2qpB5TJyU1kze4LzIvYu853cBjuLkVht+il9UfWKYcTzxEZ/35EX7RHRYmRVYJc4Dpx
Z0LFqOsyNncsS4UTdQ8vrrnxwazzrilPZ7QX1YmGyjQS5GMqLL7jXEB2FJadQo+M+SZr689kX9bd
oGYciGtl6AkGkF0qhkiHuaiB8H9xdUN1djhmL3qfIoPmrvEV+O7h0PY2rgub+uWvpG6PMPcEhnAS
a89sfutHCzC/jM+gQFCrDY+Ku5JfedVXwTY3PXH5XhgRqbbDZoiac31sgILhPFmSKmiI4TrognjH
fqS5/UUZpp/uyG6RuXHdo8n46pVgIvqViaidFGK5eWtwoMoJbMJiLOVWONRCh4LKTWNEx2+MCq0P
XPsuh6c2gxalOQjNu2+9tBUwVTJQG2gtF1b4gQdNzpP8+i8noLMo3cSwXniWW64lt6yiPDBUChYj
vVJozN9eew4zqsXa8Rq3do/yO04ZUpU1irzCbKeTj7bhpCh64sz7UO2cyulpvH96/plWjN0pdEIH
IV917D7FSCdgnAFFf0nCTyeoJ/l3OmyfCg3jD/Agpb8P8wXQ924nTCMLqmTlyo/5gW7+fYaTiFFH
wX7n2F/rVWTrcF/Xx+fszzF2DlFkPYYznfqZQm4RTW/sbXv4Nal76dFAR7PvKT3lHfKCEB05XnXl
yokqWmatSeI4V3bp6yoAn8FnpDKSDkBvUR7UO09bWYXTZ+xnSxUyLw0k0+w4L+ppXbvcb4hyFvbk
zXXdc1Y7NcEZYiIdiKJKRkvWV7ObMiHd9EAW/kYSEpZNU3lgVPvTjp1XDFs/1EbUHJ6acV4baxV2
O1iGuTmP+dGC1fzm8Qwz00Jy8LIQpiXaUIqPOWPuLZcyq/IdnmYcVPVP+tPanMWggSSztE7xhWa5
EMoE7nuIplYvHl9Ym7hHi36HCbAueX98aUuv36Z82K2I7HwjxzwaTsNUBPSAPVZ2lZerk7eRYMd8
JGB6aSPm/C0iIxMrv3BHb/MKI9VrrCF8dYtLrvMVLsBVxmbfr+UnKREZhUX8D2972p4CCQHY2sbK
0Lks7sVFVm6PxeoQ1tBBsXES6jK+T8i92F7CbFs3kuDMrRfp/6WQ6B44X75itVu3hK1CU0VRip7b
SnADBTUty0FKdMvNG1ouT2vGwbt9Z8jxPtZvDmte9wNTDeNJHZRxiYeN2rpFxgCN1/yndukqieer
y+kCh+SDds64mOwXGCxt7VWFE6wAfQQNtSJuboOZe0VeT7r1tt677Cu0HrJSUzExn/uXq8HZfmAX
3zL+jy2ykOkZCfpiyzNP1Igf5vIfApaxjwJH6ED7FiegF58Kaz2jh2MtqZzyK36XZWIkb07akuBH
N00om8Rt9xY44mRGgc/Q2fJZ/XUfxjQBhTl3HMCQZpw/71f+c7blej8xAQxPlVtvsdPY0K0ocCmR
aOIM6PiP3S/P65OGBCIjU3Lhu0jwMKUcVEkqV1z0yRRDfbMMyKP0OyUQM+AU7aAmWomFlWh6Sf55
M6jr+LIHpyb7Yt5qgpgl6haRQdQojKUXY2OTXjwoNy0eO1SjaLIfjhZ0Dce7Mx6uv/4xV2mxtEzH
ACcDwjWYLMdIef5xA6R8XMRB2UKbwWMgPmtuBMq7HVOQqMVkI+xOTjCgI2TPpPdiubUtJ7UPcwBZ
cUy6KGyh+t4THkXWlF3T0i5Vge89QcqWOURbFDLheplfWChd36qLYyGnBpVR6+URYs5jsZWGBUrF
RbMYwyJEOZIysGqw5UAML6ScbRydj6G92BGhet/mdD/NxYvV3QXl4asieOu8NFjUDqxzUA0SRv97
AqCUz19qzgo8y82ZQp3XbLa/WSSU7SYXViNSZ/0X7eAo4+KMZm5k4DrgUeMFKTZUM3/D2dUYB4lz
q70UyF1AeJyJH40ERUG5Q8aC/kgnpclmYwziRitpbd/c6jFDPKYSt0RSKaKDHAC7axUoMj+2vMAO
vknnt3kFiOGlVURSEfBRvFxvYzEOIyipvvN/dA+bCUmWK+OTA3ondqsL8CLJlvV4VaCfdwKrLZpj
YeYU+jCecP4teM8xQ928ouL3PzicAxn6XxPE6iyvng1MHXPA6GQGhKXWH/qPh2RaVu41uSfpyr4d
8jWeqa4zpw7RZXGtn02IhlNGDbENiH2+rTGBAN0uDrdyFJRZvGse0711eK8RJ37wk6zFRHWL358G
GjZj8h72jI+HvXPOF/R+cIuwvnskHatI5hM/yuGszsloov8FPvCavS+5vubKfWS+EKpF8a0nq6NV
kZRggEOkQGnoFwXRNV/J87BOnviVtV3Yu9YWS3AmkV28K5JsbU+64L72OCyK4wosSYXQ0AWZYV20
A61VNPfwqKQMTJaK2POKHArlMj8kRyTzkE8skp9uTLXUHgRxFocMBKbfIwv5RTMpmJ1AiN9sQ2Hf
HyuQNjm5bWpixcqJM6wbZq8jFut8pQGu3Fzx4p5X79+VwE+tui4u8KGnpSl+wx5qsQsPkhjfNKKT
54sWnYkmlzEsTec5m3hmIUWPLc2XdKPc0kpZrFtyFmezI7XaqlaIDrxLFTbvkJBHWthZ1d7tNhax
os9KA3bcqnwyncqjjijNyqSydn4EPtQBNhorKHBm2C3WXBgwFjHw4b9cbj1c4DNvjmwOFLSstcR0
arGcosB/dst0ratuMqfwoh9afU9I09cUPLYDcIZqUjR7Jx98TgQr+qat649tsuww9XHpFFK8dC7Y
yU7IQgJIHpFgUsg2mzgCq4bzRFKLQ1z2k7yI3hd/umjBbIhybX2+hcv1zr7SedlFrZk+mSd3lJRT
5rexFpggktbza1WvrQGZ0IDoeDZ7yAeJPrTIXGuSjMi0pdC1nDuSNETtyY+xagGXnDMLUmCRx/Vc
Dzk4ZYBY5f1TxPYh8Zb/jgOLJIX9pAa0NSLYEY12zn/vo7VEhdro5dUs4o8M5YYxJo1Tw1Zh2LR4
GrYzHjI7ukSvI/U1b38YrvdnEcz4HhooFHOhfjOrHmbnW7hdoRb+MLk/ehVeqOo3G4O3a0fWX9jb
cJxKb332Z7Uwd0kYDlYaliqR19IATZUNUFA2g0Eu1f+j71gEfZ8EMpfJioY/GJFjnJJdXzbrbNF6
V7WGnPvViIh6bPO9MuxSIshvZ3BfUZyZnsl02Ob435yzsGO9QP14Y+AiSamRYG6zQch7ol4LvMjU
3U8xZBF++Ph5BRQu+9byFSIMg07JpQNW3hOWTX4OJK7zsOnX09+4xhs+R8dJqHKFZpGhj1RpmY3B
5f1cBcQS4q7B1XBMINsHFDdytkNIA3qjzpYNES5OoTtgT5RcU0vIni6Uc1i9Ny7/ttQno4LciE5R
unHO8BK+cukMUdGr+0WerqoEfckpLXmIV2QeLhkg8ZQJJTlTF1iweBvb8V5sjwyPCvi3+0CHHhOz
+hEpDzAF2UP51Q7vUp38wAgfOanRPMWcUYrkgeKd+2cw/qhn6yYbt7nN4bd3b36ePBwBTAIdE/Zl
cyt54XHqzVWTZd9lY38aEsS3mDWmJjVUekaIxaVeoEofivqm0Txso/+utSJqXvtvjCejv2tEZmBi
nXG/Fg+42llFJlyUSo/qT+6ZXZkNcgvnwgmYeSmGfQkmrKluNv6vmcyNm5uIODy62WbSzarn4dbm
4q2rX2DaC8DeC4lzliCIOaDXnCGk4Q1wCKg+tzkcuceXsNa1CTb6bWiHDnIz3/CJo2oorDnX0wdt
7qcOnsrCMrSE6JGWWCPpx40IQaU/zmTCrFGHSE0Z9IuVolUqCLyItx3JOaQNphORwUWf3vt5Xn0D
3qNcuUd64X8FIh0aSr7DQ9/0/nYuSsKah0XOQbnStInB+zdZWfMArggiMl7+aR68vBHQZ3CznyST
QQqyLo6Kcl2/2WjsB3uVHg6sHfktZ38QPw8JBU+EPm04vA4FTFna1FqA1mXHJXlVn7XLPdasLdEW
Bz7PnlE1fzqkUamvp8rokQuDgBsVJxBm2CqIwZX7lEMWrGhUa3+QNSe6K3cztqlIr6ixCVVdDJZb
wLSsvUA5RaU21aoeC2PfOjUoB55wFDYo3uFi8W1k/1nhDYOuMprAsD8Iop8VAZLBxBZz2U7XEZGF
s+RK8ZlD9qTKww4LVJ1fkSIEtPN8AXmsZFup9aISe++Sg8JcQpdN1N4wRVu5kcETNfpqeGfuHluQ
7oxV7gFhN5TljXg2zTFZIEhMZBMoG0JvgXnUHC/I7S/4N1PZrP4A8jQfFAnVGbMeYcMFZPUIQcim
883LZQMX2dh0EZ9rDGp77iayN5lBh+yw5QrHjLYxaEOO9V2qlMy1Ktwem3z2GmS5Pt3Uz1NmPwJv
8pt0R5yaimq3ic+HilnkOsvuTgRdlm2vkMF0jm708oizw5M23hcKcbmEcw2NwvInMXOiwcsDn1Zn
lpxW9t7piFl/FSGks5GlkfLgpLvKDM1EfvlNCBs1V3hziIUD+qUz34Ca9hiJj4+T91b7b5wA04F5
i1j88UfrL7c8eGjYymlw1b0vL7xo+bfaIoEi3PT1gTbxLKC0k4Z3SwGJt2dFNMR+QHmHhdU6zqxW
IjOY7GoV4osVYy5lykK+iAKdZPMDOAKln6ae0gZhfayt9teEfOZ/VnDP2mLo1kXiO9/2fqb2abzk
G9sAYHpCuRMIGeEA5e60/g+p50H4juqPIoxdKAAMuZr5w7+zTzyPWvAVl3ulQJ9/SfY7y6ygOU/g
sqeMzirC6h4ZKKcJet00nfP7vCMe1nbOPA25NMw3BkdY7tCwRHcTQD2czoAPBaUV5HQ/Bz0f2eVo
76Wl8jtGl0E8eDi0T8kpOTiRLj7MBRJfqBdYF+4zc6v37Fy8KwnYLgu5B6PlisIyP5akU74wUXrr
ZN49eEpyNQb7gX61N4h4aWAuymNFA1Fv/siOdGAm/kX/q2TOzVHQLC9+yNjj4sc+XFrNPYqg79lv
AFbNOZsPWQrAQjaKq4AHVqUxB+dB6THetlMVRvoSoA3pZy06yC3vl+ikABHhvgzTDhzbfxJeZc56
mHmC3cJPWMNLPwX1QVVyOE6G3CZrwBfATMpYN3NXO9AJQtgF2V3Qu8hkBGlPSKltdRGIHxEdJPct
Ftny05LdFfo7nNRM+7h5ru3NOAxpVlvBES01YCyfMmO8kuaYMV+w88xh0Zcnuh5RRWyCy8lq6GwM
yEGc0cv3Vk4eN2ySkCJeS7NU2c6gQWSKOUnlqEbbjlls/OWRobINXikVdcgH8l1P4AzP6b77Z/m8
y68uA2v+Vc4c9RDiZ6tNNXAR7VK+B3V/0WtD4H78Z3N/kOWJy3pfkL2/wmJdA1ahjhPEuU7n/0sv
1RzCoYYnGTt7ZsVF3E4wGaSNYHniJ4xEODsMe1PKOr+wBtveUvERaYHUQr4hqSyiUCbbyhKadwl9
ESHw1i7DnQCDC3afQnHPxLPKoFxDAh+KHy0Wa4Xvaj/v6BwQ008yDmFQjjmUVlE0IxCUTZFlXFCF
o+DnbR3P3ffJmCbLQ0zPccF2TX6391QnQREsbdCXzBXZVAzlcblumFKJzbT9wr4Q6voFsmgzvghT
8OUzk1GhcjQIymTNG7uw3aJzkyVNdRoksMpO3Bxxy+AvXKDx5Mj30EDbGoRTlUFNMu0/7HBobc+y
tAZHkpavuCZwFDZ98T4pns2TIghsANam42SnTtkkloajcsz8evCrisbyGVeBqdQorrLJdLqvN60f
bd7btnX7dsTstXlVHPHWnsphOLEHWsyu53QaNdVvXcr77ceVLkDnkQZoBgRJZOBXuVQfjkq3C+CM
rKXHA9oEKxXAfpqxielnl1Dgp2oUpUidVYX7Lj2lYtP+Y323yJ5vriYiFPCeoTW8xsMUrTLEFlxD
n8nfa7C29D+Mo73zRrJiQ6Omj3nl6o0ruimKsXZANzjQHwZk9xU4SsyU7BcARhzLNxHjF3Bd4W5H
8HU1aDH4ol5y1xMOnOWX7IZ1sv0WAi9HQsTD7zTL3R+juiKmpxeByhEAxBZ15UIdYrXr8wB4by8k
VuCfBkDdZIWnFdjW8Uq0NMm2w3IgdSes5V3x8LsBmo8F0sVRCbvLgDjz7DGQXgqb46FM5fI8zt1T
zgzdP5DWeIcM2QeDgTJ9aR1HZ1z/RXsZK+cpf/bJAJDrP4ZE7P9a0g0+W+V9L1BFHXwhKDvg4GwO
25vYiB45GGA1PfxMnbRyTadevZbfWFdPzicOmefWDqEaHVPNuB4/rjk4VEtdJq1BQ5DdDa/to6u7
gosVUdPb27UI+8fPvrWQuQpL3pMFbQ8H9O6xWKxJLqBR7MSnIPKfwawJZ1ZF9J9cWTKYZUcaFAgf
+NKEERpnJ2O1ChwaenBM65FHCps5RF28qpB0HnL4Bv9tUOqO7Tyh0DnjJSUkGFuwk2vG6Svjyj/9
D9Ah4O+SFfsQguZGtE1FYfZGy4FuTRkAcayi54z1YpxAcvQoHw2WloeZvZMvEgGo/CL3jGxFoefk
seYfVK/VEJndZyXyQ6VmiClU3UkPpGF5bwympO6RiqIy4OgLKmqOR4Wxc6T4DVxq/1r4PZ2I77hF
SLniBhOldDbrS4aQG/VPF+hSzQr1kCtKEk9jNd8w1ml5ecmHKB02vVN2HTAF8Ac2TQaStLmSWJpL
KF/qX4SSb9DBFbbUutRd51lYAfcGk599zTDrUnAMihJIAaI4S5zEHODypuL8yBP3hj70Dr6aqXxM
X7keYlHt1OJxZD/5i93G9PPKmpeflR6l+/j1UgNwGSXnCZJtxSH5dByxOU3j4+xRiZ9N+QuHiIhy
g1lTJTMrznLAOgMZ1WYWLs6ezKzAgWBVV34DmJfAExJdI9hQO8Vur9oEafwWsMklhSEhwTyboglA
dulaGlkRFz/CxrJsE7IcIu7tIKmuLx2SMhpmhWKUSqwdpAUd6hUJ0weyp1YWzQ2RgoWd0KJQdFD9
G6hSpzQOVbQ21gTCAR2NGraie29vzqRRWQ8xdRisP2qMgQFZuJGiPOvxd8iSDtFx3FqRLghExWqi
inbq1qBNfgI3GkznSMdcXWxLVusLbhMMUI/NQr7MqVGdOEKHNxGNGBc1AR1l+X8rPK+eqUzuRd+C
dUS9epd9PbB6zqMxLCWaGrgkPt+uUMxgnpeOmovTUjo7wE32XLLHZ039aEJgTl8z3KSzlItCbmvx
9UZ81m4BZMIusaulr52QLON6gpRRSyMH/t+6dy2+NC2eoFsPIeqHnaGW2fIsSm2naNTWQcryg703
hZeNMf0smhXwRnTV6+sAT+eXo6icE84+5+B9q+TbJBoB0mDzx+e+bm5B31Uar93J4yXoKeEfZkce
zPQyEQQ3faW96TYkAoQg8Dlp3XFUTF6YT61HZ94DlI+WIvkX5BVOvePgitxIyoKqKMyDVPvaMM7d
D+wMrqvoisK3FsRhgdufnh/2VMxo97XXlB0vcIwkux9BdgYnPWCFSMJucnT2b6YAunt9eQhO8JcK
a1QXpkm+/yBDlQfOs9Ena8sKW78skwkeLlwlnG1rU1wSkOOMF3HBzYXNzkD0J9+b/LKOaPdHciQM
SrACjxcjXyQ2OBydmONCviEt8UJAaT+CUociLZAXc/5OviZMkCE6Fjd5it5KmSMbVOdjwnWHKp3F
Z2GJ0NNW0k38Zw6jE8TgmyCssvyRVRYurh4ZynZzmg+1I1B78W1OoBGtNH2jVMfvhRd1v+ZFF6h1
/QwkMjWhgy85gMfEoj3mOlZv/ey/uqJY60vSfjz3IIbicxljN3fJ+5+pfuor5DXqcSR9ASFT+EHN
i0f3dpYudWKM7sWlxTC12VlO/t7cQW1rqgmPq/KIpIYz7VLtWQZfwt/EsmPqU+W8OKePqjQrlMpf
plcK1LCCKYLsunYdkCfQe+uu35z8RrYXkH3t/Muovs9TUWR7xfWcQcCSu7mWiHxLZgw9HAR++WPJ
AHtTPS2/P1yQIvIGhPUnTeyKPDUH2hxG8rCydFpFonbTMDJXiAGFXKk4DwJ2FJ0vnWP0OLIJ8IhH
YPK9nlPaTbJP+FH/EZiE91DenRjN9Nec0MK0Jk8O0709rVCehqmV0lBxeRYnqk8OQRNqsyiQQfzV
dbDejUX2CQ6kRd8AmD5bVtMWtwM1uKCK4sbqpGSxTWyvQNMNkv3k1zRS+aN+PERZfnoxWD+V1u4b
cKBzjMRqWb4peckhceT2nCTIhChDqEa4DCv09dc0a8fozbh+b5y69CeILFjQSWGGeaWKZpq/PpMu
9+hU/Ma1WYVpEvchiypBvZbpsRupbaxKSxASepjRMVkfS5jfQ0G+kUWbKH0Usjt1VfRt8CVEqygM
LIJIKB3X+jopJbQtRToBUAr/uurNWMVafht73OyQKKumEQeQEs6alGx/CdxQGQ5FHRdyu64oFOCj
2jt7q3cH2yl+h9j2JHdvcjzUDj7xYfUYZJ5VHEPgDil0VK4n4E86wLmzPEDEG6UEG0CiQdAqNcID
fMKnAR5acP32zVROYfGxU2VXS4CPXY3rKKigcIN3O4VmyDrrEP7OaS53qjjmiCqbT/flSrC9HyIi
wx6mJxwPdzHfGfJh3mMwWP5SjP8kZV+g7jOSypgYpG2Snis3ZGb7H3PKsMfMfFWWzeoI4XNp2zmC
u72HwBV9uI8mG1y0A/CQxEiP9k1+GuFOeiYaLWJGjJdIZWd6RWt++wcPRXfavQxrl4QghjA3O5M1
vf9bDgSLtXg/3DJNQInOd5GwNPkhNaSR8PPODzCW11iYp+X1FB/hfU6+orXx1yjNU68iHGd9F6hC
HRcNTEhn75VctUhTeEi3Fpm4I3vFPpHM0y/U6b4mnkujpRmDD+kh20o44A9Z3l/MnoLrxEXv5o8K
ecLE5rmeuVqVKrHTwDdmX9QTe5cSwgd6hyLyWfh5t/3BSXSX1PA1Fscb5KEFttRrNoD197sLVePp
FcUYqQgq/N9D7RpSymcvwq/e2/KvuvS43qlZqvRDTyDWrLHdpB4zfdPG7m9ND9H2qJ6brXZNJzNW
JHCqc1gergnSzwFRSKdm9qWUJt1h2NGitE3z441fA8HbSzFEfiMTQwIzLjGfUbYLa4/aZo5aOIJt
6t7Civtn2e6wFtg3S2p/3sbKuU30+5ZAFpq1fmul1IU9x1969NaEFlMQoiC8/cnBFBZMV9q5+i5w
J5yKlgbLu5+t5A0cJmu9ki5es4ijmZHUBeY633710AFAw3SSl25GEjW0b+ZhvA8gDKKgDYpiLfe6
EWYVDMHcLApZP13TkFJYuC6mxtPoa8ahobjl7tPWIWZ9Mh56xFAUvX2aOOcpd/useBHOzNNi4Kfo
CDcuzqWdqWuwBbPALMhJ0F/h4uSSIcGS3s2gTp1IkWLX3ON1nd0TXVWnGPM8i2NomWa++m4Y5Xyz
692kvd/Dpvx5Zc3boiVVHRYtFhVdpvowbXk6OLw1vvTvnOfYlG8GlrbWZtQeGUBgeD1fFpnMA0JC
lSiKbcsneF7n72mgrRCSnmICUiqhKCLjTOdB5MyC2AHarGxbdKHGGY0l0+dc8xp5AqCux+V8134W
6cv45Fpa38zpJz7qMjObihegPzLYsx4kPyPUZG6GpsoBcWa2hMDf6yeUGBGlx7SWJm1GKznaXlsn
kiQnl18g2l3lI2iGZRapk+GcyCOMSNs5u33vx3M35RkuB/BLCGGQsv4EC540GCP8BU/QhoW3FK6J
9EoTHaVqxi9Ku/TE0w95qFXW7tWR3VQ94eeTka5lO2/N4TTEhZAvN/CXUgU4Oyw7Pc3Vv11wwZ4Q
3N25BJ/6nZKJat+2EAn2DQhoy076ia1mGXBjN4/sCnWyb9PGSCQvUHSFE9Zrt+0bGoOkFC+UGv7e
FJMoYfxAKmLe6yzHf13bkiM2x0SiMF8JtkeWYcigDFIlIrGoIJShZXw7RGXgOT+GE4hJEbuNyh9g
RbxnMmUEyAONcUPLg4ZFmcCz5foyJN4gpbCdgtHv6SMbepjs+eoPUEmaH+X0UnUedN9SxESEo2V5
jliHs01aIHDvnNl3GHfatcXkxzCJxknhPUCcKcYnrvqlPxN33HGfQgbaOUthViD2wU01pJso74jL
3GJ/JQM13jaw8UVbUqWUAVDaNHa1Kjpp68OR51tPQQ+vx07PS1vFH2HEbCeqz/RUFdsCz6RtDb2/
reUHaYO5Z4ZOyIo3WJV8Jj1R3YYgaPyLCRgN6r4VBsmt8x58ziAJcPJ2FyNcXLWBaBW595In2UHl
jCSHCPNe4o4p1wIHwmOhR0RnB3wNUeHe+LvkhH1Ag6cAz4/GNoned2mMbGbKLqvV4iKSj7rl5wiB
++YOY5mz8UdxP1OP0ZxkuDRJamwEOU/k6/uWvSbnlHdLq5HaLuZ5kFL8lx7ez9FfZQVk9uYSoYGs
btpm9peuS0fV929z3AP6q/FxLrr63k1MbmHQSHl/Wm9msW7q2bm1TOqaHermqWbBVqeSKtAa+hLK
x4tiasARIoOUkebO9Y6aLxlur7sgP+pSrekSkZRI0a/iu9HAWtwWKgcz+oHpz5FTa4rme/BQxJ55
20I7H3m6oTrrEtJX3zQs6aZukLj6mAWn9OTYbNbZJW0DsI9bBgsKIX6lKNuOvG7zWRD1gFMZ8oNp
/0+pjCT97r6UqYQd3UPA6Qw6RvBMVPFFyCfo2wRnEyLxCbKHbCwckEPJoK/EybSdURAdkISSAjp2
oEao23C1hfUg+gpMCdJ8Ey7Qp9gD2jyCkKbDnsK79Ubq6UGNl99ctdoLr4OSuKzQaFTD4krPrHS/
e/MNgmAsVjVJ66KaVMedj5sIa8lU2B395JIO9honVIKow3rQVbsUiaw9UJGn+1FDYvdq7laBj330
Mw4ZspJWOwNOLNhUXuur4fwbB9CrXOPr9X+z9szQIW0NIy4zs4NGwh0q0qhKqn/mIXKQkEOtQ6KX
R/NArGRu5iIrv3WJ78mgaUTrFwIPcxxUe4uF9pOq9ZnsGbYJCPL+S9DQ/qY/e4+CnFxXvo/ShrQy
4bNZw+XEQ7vD+hEYGB86oZ8jNb761gUA9zBqDE/2UAS5W2yrslMJXYfDvaIXbJpPijyLUHhIiRqi
J0vf46vry/5TpBBDQOTKg4FsQuQNZdWdoh+E9hCHNn6PEyQy0MAFM0EO5BMyLi9rziWEyxsO2Gjg
nc8rmciUwHWXORvT+isD61pk8HxsrQXKZd9jYWwzufCexJG+U2TlNrsIhraGjCJ/wBomXciIa8dU
fudIlLpIk7V8sBoTLZOELPVcBBRzuzEJDrgCBM2muN6BPNHmK8FHksCK3o/mFaSNN5NIjc7bq26d
+q0k70I6iCOY0h7LI1w/5x+B+BdNmg1tkuCObhP0Pcjuqd88xrGDw7HRt+g/c+aSJRWoKjiyujMH
rWweIDPwURQ2RJ98mCzEn3JJ7wrrXdTaJhI3ajRrF5cgI4PU6pnF65EKRHO+BMWNxYbrcKwbFPBZ
JccJUGKpM9fb3kSiHMAqkK+KdYd0joxXrCcQYGo/a/YFZJH3HQWpt5EAUp4Mca/XOW8AzXC2gyJO
IK0mI00zb6kBORwBRtVPE0KhT9c/nGMOe4KP/gB2LCXoFF9sWdiL80kR+oXMx5eDgIjzpZyAhJbh
dJ+/fe4Y9tl+RJ9VuiTl6zur2mKDX3EU4pEcUFMCVUQqptHBhllLivKoN3R38304tPy6ZjYCds83
I3roBZoxbXl1OzK/naoLnwk5Tze+jfaHnVfGVPstlnFArKaYmN+wTeartFQD4AeL2itw89uSwIwu
FQQ9n7goc2ek3xbCFFMmO9E17vsaTpU0Uk33uTQAD4PxFYG0pLlini8grVv6CYAFQNT+VfkCoDk1
lVG0fbevZvnIct11PXhMMsP7oAvD1w/02Xdip1wBF5xULQAq/eWNHtJkK7RdEL9NmO5MdN+ytpj5
hSO57/eTMOHDOLLLkX+8UOTtgbo9GEHly7lNJivoWXBX1udTrmR6wfGQivVhIzBYBDlIqE/RlVd4
/ElkUhgHVmC3JewQ+cFOe+nk/lRKfBvyo604tydqWz+4koxI7raHEAzgALX2HBzOD8Py/mDfOdUM
qS2FUeM1FbX0m9CxPJYjBGr+7Mi+aNVtKkkHjSidPQZ44aHqsGfT5EmRdorqQfzTqBxuvyJtPBsU
tM8KhwhLNKzH54RXLsF/awHNwcz0h8Dp/TC/ZYuxBdrvuexWRDpNnQa5P+9pFQD6ta9ixPXgu1g4
hU4l9Y1Bfbquw+qrqbccyWYXeoevBmWzE9o8b6e9qyBY+/Sf23lcsfgavGGA2NFYjzQTMN8s6PFm
8BwRDOm6fkXiQcBT5vs0W03TbOEzsVTuyIUofpFjZG5RyUQDxi8gZ714Yv+5sK2fbujJ/CcdcquE
U/on6tmiYYtiWCZeWEzHglcIY5gUtB2Tb2v6+cYnpD1vmEQ+k2OI6OVVerj+UEgIniqcxe7KSh1D
pE2LFD/yPFG3DBR5n3hJ5twGr22pFv1t8cAQcfRnopLmJ2tIsmImw5hm39l1tztDXeSmw9AN5Axa
bGxNQXjva2QewJDBSNXx9PBNzoVFXxHK3taHg9C0WZo79gqdBCu52WMxzdFEyQbMREHwn4MXYu2F
BD9EVSRZ1QpLmmwvGkd46YzOdKs4WkDBiMY9BTLrEBIS9CFlqcQPjoLgJtjZCO8PFg30+9Vs1KRh
Z2Jm7qDCHCdS5Esd9LL6JcPZeTMwF0ljjD6zQ6rdssEOqgC/QgyDd58ACa6279SCwKmkuIO6w/gX
qgtwUzuAull4/+DELR+9c4Pmy5MbN2iZU0G5XB0nrUlgbodmRUcbHerJzhQpl6XNcSChI1L10rrk
vCrusVaFwAFuNw7E7dveSKfmjAkATqlFnDor4KkTLsw7qHORDmiCab5undmZgXzng57t/+1G+Cu2
EetIz3ttPf4c4WA8mNiEjXqeh3wP1+E4Y/XgIbwjn30NSYcW19Qqd3FfnGLYyWj8P7QiR9QQH7ZB
ZkJg758pEeVVxF12J1XAKhpOjrzecWjGCz5ln0NTg0+ey/jvaR1tzDR6OqJIPTfzWJqPnQH4z8IZ
C21CZS3QcQL0G0WEnfbu0h8LnrRzJJKkfsWXLnzQfkJ28NLdaKqQOChXBfE1vAzPfMspAvL8BUEn
L/8YIFw38kOpUDCTNNU6kqJMpEQgebR1+HkZXBwStMZ16wCDWyZyef9XvjfZe2Hz5B/SQW9zjOby
9OR2TZqIoeiienhJTuwzn5/8U5U+z6GfxQql1k/tA/cMR1Ap+/avQeH+M1LZj3tDlgzZbst2Rt1e
lvK+iyNBbpOYgrP+HOrsPhT6vZ4wC2uGvAWyHNOooFgNEimjYvPYmkzGpjfGe7c6PPK5N63XJPjK
0BirTlW4s0rVags7YQ4wSiVpBxKebwEK7Drjl8Os5ezgQKYsWLTXt4bDkxsQg9E0V8ywIpBrcYZs
HIlBRFglmES4400+cx507To4hImgv4qcxbSYxtfErEXB87J8hfqGHfym11ZUyPocpm0eJPojUoCG
ZgM4TwLWoUY8HEpuDA05qWFMVJAw8hB7JgKYxIP/c950+mC/ibKBTL4Rle5DD8iVlPci1ahP/2fv
cTDjFpGqC9XBbI0GtWPCUq3B0atacb7dN5cFrKuZ7YaJoeCC484I51/vcS3Gct7IcTlmT84B9VIb
t0VLFgKLSocZqAVOwSv5gBu6U2dBR2qm+VLrkArxiB8FIx3+a26R2Rr6vbPtlG9ElsmYzK1WETqq
rHyiHGEDQFUdecCWB5H/gqxXYnuWXX++VWb3V9cYuRdaPpCFWSVpduyUuMp0Mo+t0OMiHBsWKuuA
g5RBx7t/HwOnH93yZYHEvww3hkOAFR+azVix4g5DvwxFxpSaVLfj+59wi3NuUvx8ulCnVK95c5yg
P+8CCIPxqySRhDekdFQfJsWLlKRK6UfWOv9h9goS4y+PeLfBJojFU7yRZBKX/ab6Kvzgk+DYhlEL
0oAhjVpQmUW6IRlcXl81dViGopAtLkwJzT/CGKPyx5T4ZKL5m6N/cFJ9cEqt88/njYNZUzSbR87I
B189GUW2R1Igrlg6HWsO5PashU8EZMIpgiIzY4CBjNcigdiA6hJWV6lVhV8lkHtoeoAZjMahJYOk
vpPtsHpUGXW78eAeZ17bd3uldOUaMjoZJDSGHSuMkXQwTfL6tHmJzVQUnQw5sjf/RyhnO55gaPM6
N3c2KrR8XDktb04jIfJgqN7ktn1EB8Dni/x7HizLqeavjlboJ/Qvi2X6r4Jh19CWqOv4fQXeRHRP
eT9qwmHj2gPt/NKnsBrWkWHPvW8U2dDYS+IrHmCVhyG2wgYiFmm2FCKgaQRvvx1o2GNIbxf5qXYR
FKyLIRYj0uAfSvsj/OEAHuPMjtMP8bRlMGEwJxKMYEdYtof5nrnT4DiH5Lat2oFTp5muYyx3dQLa
aEOnwlKYObkADjhw+hBebafrtQ0JSwqpLdF6yDWfp/rL/ao99DSw9kvEUoHgmKx5YHa9bjijovBz
Bu0IUZVrcDX7BCW+HUyTxocvRrI7mAfnQxpzMk3SjhsLp1P9KRm5iiHUNLkrEObatgmk4zZXnmgr
0aDOcmaD1qg/JNMGz3C/YjG4CrmyJQnT5hLSTbScr1Ok+zYuAdo0AMXGxyYTS8w7080/3qAazok1
/wNHgJWV5p0Ui242eosJPlwy7PQQJaVxRURNouSJEhMy7GQShLszc08r30HWT75Hzo6Q7GTX5yaF
FUF/9Bn4CU1DvRjCAgbrQpchPtCVFCt3evb5BxGRYX/zVueuTFSrYX+oyKaydk9UYKreWiNkg6xR
6snEoNEProtP1p9g04aoGffBzZPaUICoErmU6mtC4eDAP+QlJEBG9ZT229P32u7PEDPSZ2c0eivO
1QwOg0RhNFZqxKYoz05H5x23dQgPsBgQRHUkup5D1BswL+Qhg6sKkEs6DaFKPK6UW4iGPsfKXiP+
HirXB/B/Jh/G9ygLlkJfT6g9GakNuJgyylvCFMkl5DsTCekvP05Jb5zk7TbMOzfVfOm8KvEFUhMt
uKEI7eAKLJjYAhizRARy0qU30ffhxXbUthLwCUKPTPqjYjUv2AvTLcnTCOO8BaGTbjZ4OFeY0vd9
KUb2CTUjF82Y89AUSrnxwTmwDxExUWESIigOKLp3etLmk8uP9r7UEQanRTl4wH1QqXMVJQiRXnZR
qx3OPnqjar1b5LQQgG4eUj4Ju/iYsZJtU3mbmob/M4mMf/zlT07RefGduSdWGxrPGxIiaJNuksml
FMul3Mgy2y0TiLJ2Dcbdm8OTOJ5WpFFWBwl/ZUCVT/WTdRKFnIBZV56R4Y8feHTKYh4eippNOANV
KheH9oRwi7n/rycm9wSrZIYBelEVVZl5eYbV/CH+Xd8jj7e4HkFEh4f8yjyaXAt370N4emoGh7AZ
WJFlepvChU7UW8J1z33uz7mdcrvdPaUVuRkI7EvQq2CEKdNfBk9fmDCA3nNXQsHcBNXVeKfZWT/1
Q4fXERYVpKiTnXh4bqRx3+8ISuBI+md51g/iLdJXk7JiBzcwQMfGO/+pAvh6HJ46LrevMTEKEvVm
XCxcB3GYT4YZ8ebKDefw1AdllkP0urj34NGVhSaAtCOlAHsGGmvY6CT2VM+QiADoNXfJL/a1Hhon
tbbc8/LTJ5EMX3oMUJYg+HYTNudTCa1rM7ABy140qYtuKNBFXHgQh+5Ekw7diOgPt7IY9AowihBP
QTBVnOoYZxHjkzmRJYWVJVAMcrkYuMUoKXgZoDpHXZ6nsHc1oNDDkxbNcJtKILzChlcGjGyGuRMk
mMRpJoIM6MzCww+lvkSCDll0nySb5tRaBW9bPicMFXrGIKvXfH7RZUp6xItuwgET0R/3KMvINzLA
Ab+SWh3Aj4HTjF4DSgufIMSjZXxgzD+Wz5DHXBogzGv3hVQHRmBAbZcCVzCEMq6bAAbcxmc1gWSx
8dms0prkYUNfiZ2ZcRw15x7J1FLlc1MrQlotK5T8aAiuTLDc+Sas1fUTM8Qf/8f2vA5dzv23+q7b
DsoNWjTwYhCTw8GQ0JlHjGWrED/QsuQGB/NH8qF+fQwUO4GP8bl7qLT7QFGgBqpWfSrPUUFuHj23
g41dwYTDE+UAdxEVjyoiXYysiyHUzcw+OLRM5D76tEfFt/qbAmcgeVvQmVgiDBz4msJswi6mQ/gU
tR62s/tQeC5A1XbJMS9DYYP0YyIkU5fFlQzF4O7xbxM9hF2azgDq0Roh8q0TxhSYmBttgc3ZpYNq
FJCDEqBBLcR7IcU9yrz5x1thWVo4uow1hAWXorhP7i02MFcivjv9EtsatTUkruOsQUFOzsC4xdMA
M8Gg/tqAKs8yx7xnLBqoxVVtA7J8a9z5NLSBSrwloUc0kh0RkzaLh74YiKH0J0+YU0tYHZmrLPij
i4fDTmhwqdycuLudmAlXsOJBDov2PPiR96LavSZomyouk0RFCkecOCwzkYPnonS2RUaIBx4YL0Pn
F0YCeEb/tgK4eUwyYgWJCAti9lhl2wmEs/MHJVIYnl814Kj6PHT/n8SKl+ztBX4pA8xsGJvowPsQ
GJ0KUe7b/GScC+DYqy/R4SGg6jW/kAKw7q9J+pxdHOB9UK9r1MvbP4KgwhA5ylnZs95ylTniCfDH
MsSFZOsnZi3nj2tFri3Z9SSdztTWqGoWEiVrT6RZJDj6lr6ZlbzGLSaRzdV+YVhxF9IyxeIbFe3N
4VRSqu5k9nnlNIbfLQD/lDW6oCT3JwBisYSbRzDrzvE5huUTDDWpixh5l88EqW4YygDL1MFzT3Nk
QNreDL4/XSfCqI7XG2aI5mVwoqrQfdQ4+sQGEKwE6NbWoLIm47dZsC6XIDOiFdgLUxhYLF3QSkgX
4NxUHZKLJvtJygtXFc6N23r5entHB78SEn72r63l1VJ5dTLs8c6KZA2CD+DTkLNOemhchazqWIK5
pvS1+tcbblF7jRY+qOK6RoeVZ4BGP/TyxgpSKglJ/tCQRyNdG3cANJZh08pYWIsBslUO75iPbvz3
qRMfOhE4vyhI1LMmlzfdADWQ8n9Tfebj1KHeQtDs90EwmWD8d68vWosA8FsvW4dfoohUFqsc8XUM
tb9i42ih5VdLphzx2+VQePWzmgBxXfH+1ViPaOK8HMF9VKgdFp5uJJr97BZVSbRZD5hlfU2yIX1U
DObgolbnp+bao0TLlP60OnPFrNlyMyWGhm53RPG1MsySjb1lm4X9WoQ/T9ntvIVbQ+N5YB9oQLK3
iqdVuUoutL+KPi39a4GPnbdNeualjqQKqXnZlacjEI+p1AtlyFFlVnJ4NwC9dBbm8m55ZgLBNT5t
JXfSuD/2RUrJ3SyturrEWTtfBg9kxr6a39pU/xxIFr89aACjCOyIQQikhFpwUvha4u1ASvvn6akG
ui4uGiy8BbATaHMFgv/5B9ZLCVzAhZ5/1I1ZINd/UlcjQHp5Vw5+tjSwLS8z+AUKba2ghUrlhF6W
RZU+BiLNdT+jjOkC9wSBzfGxUGGChYeK21YLQuZXQThlUiy3HtX1UN01Al0+TqoojZ7RHs6w/i0Q
j9I6Z0Z9eJvW9oPEqORjg9QiTlcoTHPYLkhASdPoBVsKRiSuJon1oFe4j7C/q9gnVlpnsqteZN1M
sZJdFIvU7OCOf8hAo7QemDcmuFUntV8EwWayrW8sWYPNGmjoZDD/Xjg8jJglIZNQoqQeote3POrk
VXOqPuM3y7LbDSp8ZRgVmFRgpga39NjQK7pBeGH58m86curb88xnhcqLNvDhI0Dq41zBS4TmnvBg
DjRiiSzacfNfvyUpuA7hSNV1D+058v7G8Azu5iNCfZ3JLZacSETWjggY3HxmGY4NlRRvmt4bBFKH
GmbCvpjE93meC4go1OWKDy6i+qfsWEkrGnQ7dIrQ3AKJTRXZNh5lioTv5LC5Y3oNGqNuGsDDmqLW
vSfp8nPPP5cKvmYiCXN21sJIAE4Hnh22Ys08RjTNz8uoPTyf7IuXpRgitxAOWVIS30PZzVHJCQQ2
4DbIiHBye+YIzqzzFmwrdBBXPm25BEQ0y4Y3sg49Y7DtgLDdXbjjBqFsFpnf7hKoqUMhPEQQwVMP
thSvAuOVQ5Gb+FNA/LEE4B6pmhKhvD2pJ9TTcVPih0MpKQYKwRnECwA0VzTvKDjyDYjLY8l4Ng3t
nY8F+A2MplcpHUXXUAY9ExtAbF6WfTWOloOrPusbInd0bcU16KDE24UZN/S17Usvkf5juz/DP5Ng
atkOXHHaRG4H4B7ux5O34OIJGa9Ow4xXM6bfxJcGDGMJqEbO+QS14vflP6gc2zb0ArZW8H6RAlAl
/TjGM30vwIB3knAGNnMBZ6i/J54reeh4QhtMylHyqZxEAfvQEdKTVJp7EU5Kuv/ZamVF5eFJNp19
ox/nM8Sb3NHoon1vrNrBaoHZagG+0uRYrk0Y+b4NO1O1l7/GTSlRb0KPeUAvMZyAiIkEIFtIFsCK
LFx0e0ixtFpUheBOatoDLb+cuGzpmuM6lZtMHWBKlIZkRblXeSlvVRL3shiY7ljp7WgAuQ7VXInp
1bH6YqzSAwDM5wOq4bCbIUv8e/w63/cQUjMXZifJ5KgNI5BoHmm81fuwrB9fz8WFVV3AE4BNzJhc
wuMgNBlMVdDCyC4rH06cOmd89LJTi9YxplOfi1zk5XJ34TyguORZz66Ymhika79XIGIW/5c0BNrj
BOXJ+xDexZiNYWf2qx5xrVyIqVMwTvXjFJ9UjE104GwQPqdh+mza5E4p3qiPUtCFaR4PdT1OoJKe
3zzKKCq6xQzsOwgQ7mfq20LiHPDdA/s4kHD9ecgyr8jCQTh+ywrHpd3AKXpGvXdd/g1TD8DcARh+
i4WVifidMC26g7f+FxPj5B0gUxfiDFF5PNuRGaZ0SHQJvJwMX1vCKXqg5ld8jbBSz5IQaqiph786
tLk1kX2ArZ4K3UZa2I/SIs1W2jqaNjH3hpXYfXAzujZ6twa5fuFvzlHfFgWM4zli14f9V9ACvLoE
l0iMuiz32LWylDW6wXLLB+nlvWN0p/Nkve/XzGb+XZw6wWrMLjDfY7YLEsENd0vR6p7l5uIBGJBb
IviDAIpi11l1nadfBcpiR5XAuRjqNdSM9/MJEer2aN53axkz7Vw4xkPiOUnfwZ4nWWm4joGvLIqj
JFG7V1zEKAKXK3+5Vt9EPK9yGkOjobKDnnaawCYBTl2AU6PV1MNqpfoEDX62035kST6AYtm0Fp7O
mX+iA9imvRmd9k8W4r+gSAF98Imzp6NfY6EC5N+KCw+77PKNGFsPYgyQz5Y3TigrwAPvN1OeixNH
FwKVT+G0QqXG8lVrV0VMmCUlKpjNlWXOzNiJebhbSZOBp6z7UvZowTTXYiAWJg4D39dhF6hj0PA1
aV0ZopaIRQ9SQ6KTu+zcXQQwk8owjipjHWAgVief+bt5ZQ4V9/jxqXup4UsjTSGHteJEdHC1/smf
a0U0WBkmMdKMq0/cJvqWukmQwETDJstkYAO6CpCntEBBilPdhp9Nybh3939Bfhvo6CJ9Jo3rWQsk
wgGvDxdj63QWshi3TWXgaE+5ZbXJ/Dg3LqhmUdZz17RDJ3SegyhI0noRJiOJc1BviW1DVEd7uzD2
EXuN6puhtKwyILVp8a66/AEol/Taw7bwFHxblrSyNqRlwMagH3JaCpv/oBjma6+9cTkKL7fn1jeg
t9qCNMcNmWYTY09rqTXIbE5c0Ozao1b1epFzTuKmC32FfzVSRn5Jw1vyWITLiAgl8oAQ3HKm/zN6
nICeEzyBd2twWgUfT19V05bN5sy1yl87bUZgRz6xE1CsJiNwv1J9gL+27SneWk9VvZgWoS0u4QTl
VKg6IcvxWji/isGjW9WVD5Km1r7tYI0Neivew/aDrTVCt6P+aQRVLDZfpvmP6v3eGUJoUNXbTnSo
MWDWE/lx/b1hhsBlyqlce0iudXQdu0Vu+MIjRn5p/sTWJlLSs/ZntjWk285V+2qWGd9s9Mv8+NOh
8/eqLW2SasgUE39DI7hAW7vcgLSe1zdos/Iw66eGWrzNRuDtlOfmhoww++nmxzWZlYfJe+BWMMfP
3lNISpMuSkIhCrbLQkzCuONY3MPRm4qjwu31YwFL6bw6OtzSKAKUYpVIIQvr4iwnIT5d/VHRjNqe
qadg7lvQh8+kIGythU/GEAv+SqMjjSP8TlX/UHgFTGhRfHBct/dXq7Yx+IBxH91W+dWYXPtgWeDX
HItkPhCtG8JzBShp2MDkAXY97MnaT/b4px6N9ptnj0sx9Tm2HOl8WmwUtueBsT9f9/yMewPwGjw2
uwUoZHAVPCFKvvxUwPtxtAUp3njK+QYtKR+BFOOCjZBOWMNXmkb5o0abrpG9L7/ymD70fWL/R1Pv
XrHApigOfYWejllZMzpL65jtP9yiQZZSL9rRWBXtyiDUhbovgHyLwRMivsnz2HuqwH2ydZfzZqde
hTg6CX0vWZsGg7IFFMsE3vO6ZVEnU44GhaUFg8JHKVi2b8D+IY3NJOcOFYJmx5t4QqSaBmypFUDB
AE/HtZtQSBo5yb69lrsz4iFJbYgPLJsjfn3eBUJPwpICXp3aHPVPCveXvmuP5LOIW/essV+lDKfb
cLi/vCragu+Waf6XFCl7haBAUMkyKXMU5VsqlwJQ2jyxBEMT2HltqJCmJBeh7L+abtBreZMX4Ni6
I/d7ya23s3ahY3Tokct0FQNbxIG3RZcfWzg9L4t35pnTYkK9XvtQbcT1U8/fM2OzcpMVyors+ZAB
GaBehAt3hJYitv5E38pQKvu2HvMpTXB3BKWjFxaMejLI+W1nDmUmdBt6yL3alKo0Yf0M5vbdZp5J
h6a3YLQOvuGwM4xom6r00JxAz6auNklO5xQTt+5YS7zyLsrSOIBnroPIPcrEE/3W90/T7iounUWQ
VXtTjGd7Y/x+PlkeLMTCedqvRphSFvnxbdnP7dkfUtwxkHJIRXzhdHkdyWcbmb3XZy4YsfjBJhd9
GJ9YYcuBmYkSPXg8qol7FFeuCC8hqILxm4Kzjn5UlaYWKHpiqgpOvq2nGZ+Dq9xzSMPacbIdnPfL
pSlVBzPEy0peCSlyM49wN29oK3MXpya+yWRWkJIZ2sHx9EEWV12D69k9i6YiInupDCtgQJPDl0Y6
8WQCkpLbQ3e7GEE2zD1RmIYtoAqVlYU0Po2m9tsX1cBL7xt+x8GN+BEvzM82TpqU2tf5d+mJZN2J
Oe0Cj0wH+VaET5NcEU44VzBzvpFUHqo1s/2HdLpZjNvpdXYaAmqr4g4x7dqRNHXedFH8yBHZn6TK
ujECFJBNiclAY4WK+uzfDM0xR/2DN1VkhTRE12f/hgJaW5+C8SLoBpPcWP7nfrpydnPMYzMub4ov
+6uBF54MCmKAoAbr5j6VLFj/iHvf38/L0B5wzHehlgLmOJk3ZJAxPNVCRTnPf0MjAYIzT9EsczyZ
5HOkY/pxeDpR/uTghlz4UD1kPjC+3Qd56CcH6F1EASJc7PCRY80QaiMwSGfCU5HSdRuUNyemlBSx
dBjAa8QRJbxaIDJ6mp9ggPcJpERLAOkSb3eTOfXFmtbHtul42X/Rdw+HhM0SRSdVO8lxJkrz9Tj5
LS/aTuQnbYSy6WZ6B9YeCY6Uga/EG+IrEBLTaHTUdQT+J+/XuoHDIv8ZIXoHNbpD8VmgAa48ATJ1
4ByO3Kv9qXQZKJrcJBfjJpupQsGM4/iHflxTSbGQC/w0Z2riM/YWUBfMYQpm04FpcuzSj4oP+O2n
wi1hUJzhBL5E1KF7PgSOLZAdqN6khUgVc5BoK3YjAKPR/kD6o6Mble7juBi1mXR/UyqPSrXW7JmC
/j1kBCoX+70n/v3NAH699/gmPmbpycWcV4Yof9+wtX/iwfo9j4O0iUfQlWVFUdYr3VtKWBA39NeJ
bKp6Nv0zCU3UiH0N88kGpm4mfoO8IBpwDD0toz3ft1kO3NEGM+2Hcg9sdL7v9gVJ9B3sRJTAhVTL
9NSBFXVA67JDjAumGV5a5qvx3fE1A8sRw4uzYC39m0iOHEWeppXH3gNlYJAC1ogHjOHos656U0YT
Li9OoPHTwvoXOER2NRV5A9MmWHFgtSF4GZ7UNtqNCi2slm0bg5uEtpG2i7XVsTTXaeL8Ff/nFkGF
PkqjyKT1anlMUelo4j1flH0iTG5AdhzXo7397ShkvqErhO6KWRsoyc766+XPp9FCSyAw7EOpH6OM
PHCmKIM2hNKbMhJxXVediAWHW8Re3AanB88+KgNSgR8NoLKFzUNN19WgB/a6Y6Ao8uiohFhsaV/X
ZxkZWx++gjLlaiVwH7WzdXTZLFVUpSQYqdKfa775rFxt58Q14RC5KmWS6HvNQxrXMJVLQSjsaflA
5jmdQKgn/5+eWqYI7qh/q/eKUOY1ka6uG0SsoF+9zyRvgWjGwCDtOP1/OJTP4iKOZmx8vIqZLGFS
r8MqshDJyGAxFmyrzM3aVtRhT/2jxGu6ZJq2ojnEd7YZxI0gSOCNDD74lpDpmH3yGN1CEZHsXzNq
bGy2hCAiYq+bV3Nig3A+KvLVgtPzvlzKKz11uQ6XCcw+afyMDkbXXQVzn4QRLkDu4PB2Dvto9j/u
kPV3ylnvuhspn7lfR5KTpy+aZlW7o8OgrSWZWOgxVIfquPaz3fvfNI44m4J4BrgLVSqz3ku0vo+q
o47EUxQC26sAweXhBXMnPth9xiNUfugoqDBNNp0TEAmt0CtzNgMwZwrw2M+BFKpLeZgBfSKxekhI
7Abp7W47EIU5CfzqHzWyWx+XCp8HcMDCARBs4Tk1dZ+ZAn5tgew2KoPLC1O6w3jdJxQ8eVbQuZ5t
jtaMTT72ZfsNbn+C5aLJwepJCXbDBNClFy4PNSyFm94/wyj6H2hhkwWLCHWzTE+BzvH360nYp1+o
kMbCHGR5Uw+czIgC9iqnIhm+GqL2+1MWhXUQbcDUkmgz8fDHvJ3q6TOmhaxOki5co6onaGI/zrBS
VZ18Cih84uXlXNyvePwWApkBbKxQJIJNKP8YOZPpM9nIrHvQD1UmgnsiZyhoibTSWvH/6Vc96EGw
1TR3LMQZPBmcUbSd410pVQg0MaHC4ngGH3jgtVBsc5IfZvltbkp2ITkBKafvUY2oZ5wDmRWS6iIj
61olN1jUUY6FrRdTH+XxaILge8BBf6cW5eDbGb2d8R45xEsMTeRM2JwkF3eYjwedbu1UQ8iFTH/r
S0DRjGpi5Cb5Pk7R3oALhDNoD3wUw5JPnx4STQklI8TEmtUvPz+nLHtQzs/Ln4slh8FLGHfweLF5
moLsSClpEBmHGRl2Re9A06rFSLm9KQI1MHqDQLxsdvVh+iCrdAJyYjzZ9bUlmJa31In39+joU94c
kGNpeoNjlWVDGAhbdSycNn8beOI0j7XKerbKEkVEK2kLrjfno/3lb5LbVOXyBdTXjyV5g8zrjE8a
Qa84+m6n8EXhvh0zYGynpBl9TYKfv/NXWEzuaHG5vA7uGxASspBwFPyLYqCQ5GgEV3CerKYk82wX
Xvxa80m/lsub6RM89KUj2rOFQd5txucmRHuTmwbrxfcUr11MNbEIt8zQ/EO2jcYgci7p/QL+0d2a
4pprhjkPF3NXbCys0vE/d6pn0fQNdHjhrdSHFbMOgVVLrevURo4vLMBvvyReyoqSOPgHgn46pYXC
WbjpjwnCtKyU08ANTV/MMNhiZtupVJdWyywS/18W4Wo9ruMHLf4pKPKMtvbpQ4v1558ALFYjBB27
oMujdU5mumZvvD7yThMQ09jtGcUiKR9xaGMkJlkNdVSRfSA0znuoUVekE//sRSPkrjYoj0WVsLZ0
qPQGMJ48p/6QwHGNgPK2gBZHqPpIaD67rOSksifwss8SKV7PcHiS9mojo8u/vf6aARzbgdEx0rTP
7kxcSOtgKerQ3+DOLriadQob2w1MPcuZfsUq6h/CWH4+kP9+OagMGXdw17jSC/v33EASffEJBIzT
bEu/x4hg5Gm5Fd21VfoRBQGd9HQWgQA2hlr9kcl5U50Hkviho7Xm7t+3hsmB02nAa2eWdMmIGfVa
5TJNuDz8Tu+3KawKK//JtjuZdIM5VazJosj4bWf3FXI4mIxBBxDVsGVzJuSMGsQ9GmOEE8ZH+HCk
D4SDTeGWNUUh7H6xzuPF0bn9Om+L1CUbNInjqS/SFlG4fjiUbVOGLnlybAS+3z2zL0m7rqaHx+xJ
Zl7Z89gwQ5pahqpkmqDQ3j1+dCdpxRphY71R6Vle2NII9QBBHOtMTNcuhoVXEl7u63BYFgZzL0rn
B7bXd3UUNaY9ykZBX6iLDGefZ2jrmNQSWifS8kk6LHT7OMm+egvOSUUwukBxLO9CSeHDIZKzBGBo
0J9UdKTVz+BKvbu47IuO18u4ncr4B0E9PqxHf2+CVudAULfTlj1Qn7b5NvXlVDlHCwNFoh8kfFbE
SRO7J9UV90aU7bt4RmlySQWBAoTb73sWBz5uXI207AVkvkI8xZlt2U7oAs2csPBP947o3Ur/uYL7
M83j66AOq4GW43KhzQdRW9WtE2QG8AgKLA5rgjkNcN81XkDWpOmb54323a+kkSDDuWBbVTEyCRni
GnWKHpPSpgJcc03M/q4hcD/MJO3sUOih9dKR0xbJHMpWFvNsNcnCiaq57WjrezJz0uYrht+rgAUD
FgwiOXlaYKDJssnWT0pREdSSBQuROMgOobRI/TKy9dV4ujswVlV1cuBB9ewJsyP/OaZtUvt8oq6L
Q/k3q/KS8YkXxosW0CqRcz+k7tooKRzhOBS9q74sZq7D2NLid/z3v1NTrrdfjjHEmqqEMUAxfQkl
FpJ+k+ZQx1bX7T8dlZCMbeKinKuBjbDwb39lqi/F6ADNzZkrdtEL6Aq+NL49hKYhB2hHms0NsN0y
nn17nM0BVzOvo2BYWxCxCgRtNIjABX0BPRB/vnQ38rYqpXOXyYsmXLxofg6B41si3tG4MqCwsZj2
EvaRpmtwKD1MsQ/JCwKrgHn3HsJxVo4fySEixE9CbZ5V9AGzoHfuQ2hqqCJdb6mMgAar3LHLXBWF
xjtj5abuXL0DmNSHDY2Nc0SEO4diWFV9VbZRHvW6oEdMxC42fBYXE9ia188i6WYETJ2FddMkYLug
+1oUOhuVjp8ULS0s+MABcwNf6qxAyqKkZ09F+mJVvHSWtSsuq208lr8FcZDZYS/K5o36z0ON51TJ
cgO+H83TloproHZXLPW8q54zxUMfh6HLtdcGqaW8rjRkBXl3nFMOYLVliXReCnOL9taNO00gG7lh
tt5ycB6UOddTm12WmibtnQZaKnp/n3/qMts5unslEGLet6NFcMT5RV5wllA2Zrud+iGtZ05ImxOi
gANK7Gl0Egr1ihHv+G1J+bJyOxLNqyuSNEKNb8jBTFBzgkQqsHhKYERM9h29nVk/W1km/2v4R5oe
p+FBU8ljMflQ8eXCCqtH1ueACRkxYpXKTj6xi5aAwUZytca0J4Y5CvF3hVdgMu8rw76QhpYTUpad
FHPNg2AwIvjELI4otrUHikTg0s6OyBbxIzlsacd4emFioJuE+za9waXH9LGW2+/ALHwxbrl1yLOZ
kp/isVXB8iEJsIdMbHZ1SmT9+DwfvyOoQELgb24tvvEGS2I43Hyg6ePvM5DiRNAVzIH89+Gyny/E
NqllN6Mwnt9IDyfg9xjepv9PXjgATCSgbPmB8FL2a+KDxEUkghu5KzvBo8ugTR29bUWDo/iosfoY
uyXpEMJEIfQi1naPDZfCio2naeIHDo3ljXP0O/scjzaaNIuY0D/GZVDz+0znhXTl51F3Yh+dI7m7
GmEO349PNRgj+hCciHwu8I5hf+hXlAf+Zk1JactMwWeitnDA+w9J4Bg1xeQM1fir/RjZVxzF1Xpv
mihqQNmIaX441jJ6SV7fJGNoMMZPVhwUgLad9Yzr+nplVNh7ZrzGG8FfXvdJ86Wmzjp8TxUB6odk
jzIMEJBthf/LWE0NaTUwMGE/xvo3dmhexo9EpDY5EGBEkZsav6dNgRHJZ3BKv/3tCJRZLBLnHaiF
cC5PpiuLKETposngcgE9iWCWU2d33PAPThCrFuDPRI+EK3G/WvPg4e1XE6aCPWbkr49xDWAx1LOy
0SjhzhclziylFqCzMQCuBx0YMn2s1M5IVGhqt5OIwxKvBQIraF3MUZNA2LrQECeIHCxaioVJbR6g
nCitsnWx6OxGpJ8lpnEkGvTJ/WadAU9Ar1wI1Jsw/LwlwfvjQLNxwNpBB2czU8eg4d1gJsI7LOtP
lJug634hXEa48zDpYbjnXQxBCAe7G+oE7oIcRztjQh4BDNhf/OU1sZbx5niR2OEjd2U0H5Q5b9nv
yZC3yjVV6uOJp1tuaqtSleRucVi3kEqx2hPNMjABUjWjaYUYMZP7ypmgGlicSlDZLzpBdODrvUPs
awvb8BTdUj8EfIpklGZVfsyQbBTASF7AoupIgMoWqis2XcTMtry3/ghq9pjZbTmejFA38D/2YUg7
Z/7Y8w2RNAMrXw+0Mwh1GC449Vh0sLhAjCo2y5XXVOWgJoiqLDQYg7womXFdwOStJGDyNELqDRra
uWLNGkc1Ev2heF7iDqtV+EzjxSq5DtdFPijuKCfy+RnGx7zRK3IYN1MCeGy53iy+ZvoyNvYqALmx
msVZexE8yfsuMjs8glkC2GgUS1ZDxSWjSokoSVEGr+rECRjwfo3PRkEShxeSEzw+SqNNHMlduEtP
hqpoizKCy29s26moujvqyhbo0pFC0UxkyCy4mWBYDJ4mV6DG9vP/0pnXA8nzoUL2Wi0iL6PI7Do1
iBrmczAhtrvh/qxuCk2MuQb5E9bSPJ9AeLskAWKKBHm9M6oDogFXopd9HfrIP1E6s+9M1rCwF1R4
JY+b6N8ZNykLEtKF6dcMwQC/lurDsWolrJq0O2rkfEly/L3vnP4FDDBsEfx7ufzgEZcMM9mwDpvI
75goaYifM9MOsA0wjM/0PgNgh1Z0Va3FsoKTBD1jvdCs+34QbEPC3UDRRuBTs46anA2EtGEoViUI
vNasubEwSiggWPBLqlgndIhf7idzC7wyJtvfWLja9MBns+HGQ7WTdeWk5KSgIMoro+6LQQNYSVsq
nSL8qvzoOiPJ4EWAZ1XluaNnNM6wi6IA8CJje45PmTfzdLO6kAjWmy5hQtfnU0uzFrIk+XssR75Y
epQf7mUp82nlgTQCr3zefxQ9YTIPZPSazY0f5pbNt+jHoveLbtl2/TAHratbQdYsts6+wNr4B+oZ
S7xtKvcfnW/9Yak0kjAa8llLpytuTEiLNuDo7CK5uWDFEcw9MIttKDhnxk9VH6Zco1AqQvowg564
aHABQcmVh5ST63jTmEPIo9CQl55uniFdHolU/AkpSkFNY4dykoYKzcbu/5EjJF4bNm/C+aNWY6WL
Sb4czVdmQhyOFzNPutpNQC6yrkSStCMlb4zI/nAe3AB4QuUYaPuvBctdzh6UkD4cspmaFUd+WkW1
nBUWwewMqKfq7gqtBzAlAnIEAA/HsrBvuWrB6bUi/XNpjI/4M8YdVe0CFP7aHjNzaFCeV72kG+6q
mp7YFa4AYq05G4S7XOTGgSS43FkAx13sEnKkzxo7bu7HDhb/UpCzTiNKp7bOZxq87sjwudrRrhz1
oBjgb86nweBfEbw99+N92Rok8cxkOGTk1TeV7N6xL3ZSqbspiFqmhFPpXTyUECEEVu5zptcEASoj
otk3Jrvj7UmpKFHPmX4oTiNxWSZijhcALfx5pKLT1nYl6sHt8PMe62wEh+Gck+qtpS2lxTB2lElV
EPXLPA50JNZomM2jtHn73limuMVRsCoArjzlhPaOzoU3Qt5aWR2wQAty4TYRrmTFu8/xST95j1Nh
tXsyXO155Oa62zPkimB7A3GWW/UuLZEgawKG1o9i1RZDCind8fjki+aky8vWWW4e4VoI9JlPgMyQ
kEli0QARu/7QtTFoESzCQ0J+cR1E7jz4NJe9x+ynLAH2oGUL3bHjbBA2icoLZ1ZYfGnmJSjkYDPQ
aq6DHnzEpaBhNojPJh1Jc64D0hVsb6nNi2I4m4zcackpbGvYM1Z76UAdsCugvTtiWlYmhM0CBXIl
GPQEP5YRPrA8+CY/gVCpWQ7j16PSr1v+Ny/tTRGAnF6DxhmnMOlovTkDF0w+67OFxb2mDFZ3YW6v
U792OcKyiwlO8xc8yYQ/Xv5mNHGaQnjRkNoI4cotybNLoDmAy2TLRv7BlyIRXjRxt4SCID2Szpgi
CEGGI895BqbPGRkYgoZMMTtr7BuKa9k7FwXVyf/SnZYmur0fXowOGkfuMl0wE7mdgZkVHZJufCa4
KTMtTCwBPwkUUGJ9qtOpeRf8FZrTr+iOfPe4w2f23pfwzRzBKk+qQSyA56uhNW6xc4GzhOQzC2R9
LMtAmnc5US03e8mSKwnGBH4CHaWs+T7PCwyQIo9xC/pcxVmt2seJygdXRdMPUlC3GTBFT4JYt7D3
py/F55y2Vy+hZreH5NTWu3RY9uLNqKRavZjjRDbPqOUnkaHDHioZovjQ1vpudUN+M7htUQUziBTd
ZB6QZ1ko+Nk+j2mSC3MiWqkTO6mB1Pp870Mmmwv0BHtmnE1oD4gl72Wb3HPPwy+TCEtSAyEPvzqf
B9JPhqF59dE+IfbJpd4IHyZ7Ln0ePQ6XHWFeS4OY07rTHmTqIXIdUbn4o+gJgYeuEwLfbplwAm5+
KjHyYwy0hvDdl3FxV1OluxweUi+7bE9w0ZGmFtszbFCoRxync2NirRDJG90tAu9AngWudmD1X/5r
SBuRzZBKkdEfQDLQxej0ND7BoUNnRoSmf9QWA50CuQeJRTsnnNzE23g80AHKriXD+mX+HyhpRJU6
JSTKKaSF6AexR703MeCy1xGe+gZ9wAe4HGu4NDI3bdX10Uuv4W2WwSSte8tvTxmkmHUtqOGuuH2c
9tTFb26MK2y+m6bYJXf0dj2rkA0+BSUg9BfwEg3hDnWo0SxkIn78cO4Dtm/d3Md8fS3SfIuxeS80
scjdN6W77wTDpuzhuy7fRbPsyctdLTFlrtz8C5KPHdm1B1b917OCf8bBIUlkt39N5FhAPFoC1SuS
8c9/Fv/X/iE3VyDJBXLvyzdBgVTEQPRBRi589i+AffvjKyXdIBuc0j15Jvw4cp5LV65Ri+czTEw6
BujRtPgmKvmkjYrfvJU1d/YllNJDlkkKJhRk+nWhkaipBqAII7C5AlXefahJhcP15ukYuSDWMlF8
4kObT2u03lDwvT2ncJJ/rXyKVnwDW7usKxMaRhjjqtCyjQ8DhD2LkfbuflSlSeTsM0n3OY9QuYa9
tty8iSJmxfqVI7F6hnQY5PcgH/60cCHn1Dql3bNi5v88XZkrO+csBXJU39SZjLZuVB/egMS+N8Yp
SfXjHDvuFOZooN4sS/wQQv+uU04utWP0j5nKSvC0RZB8THNOirNRNS2+2BRGckUGJCoAGFOKMHAx
nRgKSQlrCtE4mNKUrESXBXeHL/5aCDgfDcdIV8QR+TBOhT+FigtUwUTnyBJyaHcnFmhuzraJDxat
hIbaVHlReUo83nyDyni6fyAsVYs5wzyM1C2W0OpRhGolABkt4cB/A0t+lfn0FEE4bOG0qWNVb6Kh
6OLe61nLprBT/TspMP1S6Pb7WGGyiwbXPIjec1C+OUGueThkaDMRjnqTKh1o1B4B2p16hoM/4EOS
yJXQCLakjobKiofqJcXXlsQYn919o+mtus2Gb42onId+2e0JzexLKZ3ZeSaCX+GAa/6C4R9nUjeJ
mFEjSKXswtTHPmBCAGrXP5U3sFkw/dF5SzV4hlPZONkTNemLoayiJAY3aRxK2iHoZKCnr3ET6mfd
S00DeYtdpvuXiRoNS6shw8S+gGxY8Nneinp47fHuC8R0o1kId18k2eiIfhNXCpGFKkHIPY0eyPR2
2DEEPdtXol7V+TimVuo4PZ0vbwIyKsvBvTvs9Cox9agHTcEa+pf6rxJ/WcBmHZ/Pz2kWZMY+9N9Z
2TZfyuMfjbsOf19Dv+l5nTcLcDewuZSFztyrVjeyPef+6JiZWeQ+KVGgts2VnMsot1rzVRWlRuqc
/NJeynkSOknUhvdErBfDwpuJiNbHG34nWlGBB7Y9pmKiL2+UWRYEKUT6yoTLo8hjZZ+boTTRl+m3
HwofzNMxsKGoakaEOa7eywwpbX3mU9+7iQAMrOBAqD+mfgQaEcs1vY+efdpdZ/hVxvPoao8+Q+Mb
JYgYIP1sqByicKQsEVGevACxD2z40unWFDYUiZ7B8uUBumvCc0C/7UUE3IYgZa08fiUQeayFYN/E
a7QYfxAK1UPjgqNd4nYpL1qKzSMOZg+HZYy5sdKVyN7ADDwiIkuj9/Ba/OeCUIQlzcpJazrUYPG2
4MzKR1SwlljwlbTTRWJZvSf8As/+iPVGVVdKUWPXJxdwcUqWwIQ6uDN51pMoWWBAEf8kr7DgCHMM
EtRLr/UhOFjbPOHP9pJtnvobqdCW8TXfbG7wxHkBiTTv9BX47CqJx9HLIhT4+0gLy7OoAWc9dT+F
rk4gc2mZLOVOD0SCjunHOUiji1GOaWEOZNP36KP5mkdgMJynFuUq3aUk+iiwkUZvXTpyIfEZGYQl
HV/b7zur9hwUxlRA+EPCd3ZJJ4MjMMPfIJhSfbecU4aPTJE2euG8BCZFNC/RIeApCtx9W7atJ+L/
nzi8QO/SQtslnHzyhpUFavM4MfElqKfD+9V83W8+kcKlpsCEG++lqP28HneWNiTKp9mpN4Cu4M8E
/KfPbkt+TL0HOFrBBdkP2WrTKcufyJfwxzNkeInOc2ef/4h0tqqFNaj5H+S3DEcwIcgCKsAc7hLR
OTh0UOt3ugeLr7Pth/BHXW4dhz+gca4Emmewp5PIZevCScWN/9yMG8pKzchysMPs5k7VtvkjXPME
B/HNtgwY/Ounw7vpVz2L2OuSvg6aKMjOSBS0HHfKNe3tpobBdDsM5cjt0iXd2vV5TBkxeeLzSyo5
yGT5mFCmR/6wbfRkwDA2c4M4qvyTb4V0gS8t+2Kto1Jcj6V5T4tZilOgmR7dstlomWEjOIAGrsoh
7mx4MuaI3L6TktVzanjhLPQtX5oTQLVdXO2PN6Eisfxt0K6Mpl2RtO8NmZ8HjyKwLOvaBb6mlC4o
PNQ5KKDbtmczcUMtBTHI/tcRSEOEIW5ns2gJtUBQw4rSkLiLetb06jqpVN1ilWxcLIvtwiPwfrRg
zNPFqjfFj+O6Ckw+y3rRloqoiE1W7+a6Svs1AGT1p7fdYgBXA/HGVpCbK9uLI8fOFCs12kiSOPsl
3c/sfeV4GNGuNHZnlk79dekxTXr0N1LdP/l3vFB4O01VRnHkl8l8JEXemUJaqvodIbE0Q2JtelBe
wRajJnZWb3v6k3F8/HbJGjLvH8cHV5r5X/blsNXkaMWRqSi8F1FH8TvSzD3BjB2/hda2fNosyk2S
AXGWzKyaGtxK68iBNuxgp6FrK03RPuZ5M03TRpfXUD1gTZonnJIwL79Qwcf4Ci26r2MndtEr1siP
JKNzE2cLqL9PVhUChEdmLthiM+U0OZqhHzxJgeeucwhBN6S9YvI0PBYZsy+NY91/kS8SchhYcbty
8dZDrEadD4YxQG3Iku7D8TPTwX2VP0UJAjmNjaHnfEm36A/R7YBwMEIASYSUrq+67F35dKqXqwNz
mhsmtTGKUYMeh5hFrLAqSIIl5jlvhWNXV9HPnMIoUGnpeVMwkdmY/Xu8R5kaLMyzM2Uqrc03t5zL
0rL5+f3wz7anQFIAiEZP7t0dOpMmfa9KCX2hSRmjk+ukCE03JShIU40WPAayDxd06W4GNWuBaFw8
JXDSX1W5IVHzWXwdoUJVOhRUoCQd4bUX7wc6iARkeHtCQpu7HsrJ0f+6C6tLcoboNx/HZpzm2Rh4
0mbK3EIVleFZIcpNNBnhXEf9oqg9S33KAsMtmPbAD0Ju/1TUjK8JnIS3HRLb8RcapCzj6H7ZGR8K
TO+rFPcDyy6EnkAXUj78cquz1RmPiB4f+CaR4ZfHW093/A8UF3GAOZMBtZ539jP6vFQOiV1LGnzb
yYYXwdR+Tb1LWy6AyGUN4G/seY0EoxfEtT7LCuBRgplV9+BBVQ7ToDbv1YVuRIk7SyuU2tFegvTX
CQSYAyGL6Uz7pdqhHE9kJDy+P8sDfif0z0iFKg/N2d6JRlKXdFItMQ9CZqmWykLPOMALJ1BI9RV6
5JgB302K385fKTk5pViLLsBfUF1iwFQmWDw2CGih8G2uq9UZXZkLhvkYYUzaHrL7yQIffkaK3kHD
rDqM7Vn4gWKsWcIPupqKeBVDqKPi9TNeQbXdrLsvJlgA1ywOj9j76A2SnJCNOm30tLXvoEFc6Awn
uT+3FpgzROE25BI/5YWUPZsliI2RfL1El4/tKNiikh6U0dlMtZMXVE8jnDA8jbaODPKJOKKj5WPn
Vv+dc4VrZ/3EKE4ZHMRzRFwt2FdRAZgXkv0n48Sn40/X0TyGWBrLDySHQosNFBAyGfa8oKW8nppr
S1ztigHPgVC/W/MPMSlVdtoqeVoV7Hesr05QkhF+xqeUkSyWc2qusUZosQbG6nl7gS49qqhEFga6
JFqgFsSNOjqHfMcPzyuhMVhM3+65+1zyPLBUgl+BV4sMFeWSILQ8Due06DJUimqbVJXAeg/p0Iwk
p5tetDaib0T6dbGnWngH3fRTDZVO0eM4xOX6fNwW0WK0/s0q7Zbfsq31vjXitvwoRojyZqsaoWPh
sAFro9gO2eaGu53jg/ehu2C+YzvZQTuYsIx7zWW2WLAtJxgNVYxbz2jay4cudg91tjQphBISXWlS
sNw1Xk3nVzfrcePAuWqj4UHJ95+ouPGDpS5xp7NixKHuH1RcX4WScs/b0/PSQn1/LoHerYRxvzqp
VYLoQoAhkgwvk0qtzoJNvQ7IgvCuO+ld7cnQw42c6ytzXcOHD3D5oEwuvif26puaBUDrXI8wKiQP
jJiHg7H6RMT7IDEIKc24F+dMgN82m79Y0yywBeicpOSWXizPd02ilqUGBpfTi6EZ59lmf+uDDrd1
EcHI2qPktpXRZcpZeBx187pbTgelpeG9/ptXgDo804nNRrSb2fpvpcUZSa1Ow0M+aSjD3GrNnx36
cd8l/NiE7X3cqMPeh5vrU0uHGVr52MmkfSmk2P26gaIyjrC8/Qlk6kzKaxFZGpaVWf7yO0dglkDN
snF4EPvw/ntq3DcmHV4tJ8H9IhKHuFm/lHobfK70PDWUgS304t4LEAO+2MRWWEQ4tFBlTRjctcZv
mGfivSH6fN26F30vn1nwnIDjAjhK4yUqrCvi312SzniSxG9hyMaCfxc0/W3p1QKITm9deEan2sHS
jrRM2Mx4tH5QIduWd/c7ekSaRnwwx5TfagLXeAHw1UW2icvkxrsEr3i8HHwrogLTEYoIOwUXQHyb
ipoWD5NU6cEAZ02f4I9YyAlS92H73ST7kz7arkqerFDbcxijMPFxzLdbd0zoeAU/WmfHFAebrtWP
Rmn7WRv5EVH6olgkJjTdF9GXBvWFz0DfMx/apgok040FTAgMuOiBvhJ/n8jy+54e3MZMqqO8jfly
CH37lzMmqzy/VXJKrM5CsFDF1LXx1vTSSquvdkSg3j41Y/4RqwIihUrU27g9xonbt+FcxvcbPa4s
UCsCE4i8F03G7/0urXSM8PiLzyA/mTXF+YE+7b2VA2168oPWlciwQclVqP+M0txGGJNhTD25U11K
8IAqnKRKpPeZ0PU3IagB/5SaMrk50fs6dKD12XeSnyZXC100gKsZjhVR/QWZboEFtPRXsnIbCNaV
H7SaRxic8Qg0BYdlOyIT5CcDR0QApyERTYslgzX9WGzOcWV4Hlw1oIo7ADegCpAvWyNhFngfLfAS
DMFfkhX5xC+nWQwxKIpLeLR40ovfXpw3C2AksNmGrnsTDnlzqzWwukcTTEbMqCY9iF3S7FOPVwal
QeTBMzw37jX6RXPcBlXLWrCLp5l4E56F9rO7eKlyaQx5qvXxPCpkevo/PzJnTSeyGMaZGeGfrj+6
BteQJg2iyBlE1kn9D0+pxzOmQSXqYCzeHVGcNfoRnYfZVBGngiqXk9dWbjQT7wRSFG4+yD4z/Oib
GJ79HAZAbGigp3buavTq4Y5ydZnSsktRIWatu2sSPBkQhP+uMZRfj+YHUek8ufe/3ymdrG0ByEeY
wtwS95MGcHXgBHsRptv5WN8cgheAWF5Z5AO1Qxfy53Xa00al8Gtxi3GjbPcC9XeaIi0QalijNOYs
rZkz3U0ANVmNrr3I3akVOiK4Ft652hCf8bkQS6j6JEebAcR0Jv58g90ggFCfs7mQj5MhXPWL2mug
t4RY81S9dYFwnYG38DHOHU3Gig1O0o3F1FMLRY80VdH/C6e75qq86PA+nh0sHa4WuqwNXQH2fdkH
QW0pK24X9sZvKSvgIknZ60upcCC5Ur0KeG/DPtwIS4PPhMTfxq1Lx+0leGweZ5LNNBrfYGB1srxi
BwiqEfWLRiiVYYSgslvuJL4ocUJI7IoLCCYe4eHwkNBh5v0jXrVpF8gT5cHtYqvAYcZwV1T4wTWo
mY1Wc5VukGh7ubi/5VUTELh/ALztgOcWSxNG5jOC/cV0EGqUl8hSKWHp1B9+vHe/FL3TLeUbbJY9
xGyjx72xSJhnoEiD7tAHIB1F7VOHVs+Nw4vEJRYS2sVgWi6PKVQ5wcJlxZ1vCi4iO32iqNcm/duc
yYor/uLOFbREpk0baPtElWRdcQTar5bdTbsYkzqyuV3lcctK4+/sX0ktP0mWvs6jMvgtCHP1w/xT
I52Y8T7MMfXMvrXXo8LWPir32RRzZAPzvZDrHC2xvPO7Cs3ckiwp2WGergCLGlw0y/tcmTowhe0a
iypb74/knxQAKhPmq2SckqETK2A1NnxE1EcQwpszWW/9Cz/5gFcUOYxOjidDPkxHmXbMTRt2hmQd
wD8HhjXhVW9h4oLk5PvMzrGbwjvOavNGrqyfcmj7sQXCnincxXKTtkI1gildQX4FBHyIwYYZmNXq
KpQSUSvCSYkxgL4x6/JOvP8QgymLSP27IjrLpvwpX2FJflTZ2cyyjrIIKKSmWYB6wTAD64ZE7Obx
m3e0W36pxYszPCgonRrhQfH33Os9wDNuw6z/opt6T4m5Lk0pEsTNQchYI97tFkjO0snysPv4wfCl
55YittyEW0ZYa7n8NVgSel7jRYBkf0wgn8ia6K6nyBfbUJHlmzYuNHI/ZqUwyj6kMBesTD7DVTOG
dRZKBZomfXwVK9kqsBoWqDoaSzTquxrmul6Zj1B0HcM29ErfKZfXLHh66JTNl8ND6eRTm96QIOF3
oz+oqZfuurHNwSpnXgQ+xyuB85Kk4J3LkOzZhZdm6JkGgipMY+fFSCCKAqEi2Fbm7Bb0uouL/Avf
GHMPkLiaj5Emi0pp+5ZB3KyPjvMj6vFCAJ3mXbr/DMo2w3QxGfYul3x3MatGzBDu8JoVTG1kuk75
T1zZzsSK0nag+QeGeIl/IukNqgFRMAbAgLT7QqgW6uKjbs9i+pURidc3vuB1ERpMp38bwxq/k3Vc
LtBz3bZ5meJrCbSa2Hdk9SFwbntwpm8xUBLLW7tQ2DBrgA2ItouOc/fAXgc7+CJViOqokfU2nqyu
FrZ95Gz8iY4r42RfddI2N9k6Hft0JhkRWJIfeeEpwtDCXHVFpk7Dwfp84ez2CylxZ5VsBHyxspQV
dPh83zW6X574asTRw/yW0Q3s8AlLpPeOiIURXreLPZZ5KzUe/hqYrUvu2KX+yR8yYLBSzUS0ds6s
FYYAKFHwA8DCfm1vtdVxDOxErRl6kOn795H05i60YpQMOAkaKBfVauc8ozSu89WmueWuV+tiu6g2
ccOGvXdvSLjMIEBpw/3w+x+OF9fP/cTO1JmOkVnG5he1VMSsKwpTNWteW7Gggl06KwQUrUHUK7ct
X1ujbzUYPPpPpSqXn6sxIGZfjRQcIEZL0acVgbTg1yYFg2rBUkgV9yeKmA+ztakxiemq2dObsZMv
nNMCGy11hl77hdU/s3q7WxuooFSZHE90buyUR7Rck9AVG54uEGir7z6qYElJgu3IfeuVAfQDpILO
F83I8rz4AiqonCNTkj+oJiHPAJokjuN1/f+OeUmllRlzUjfaugPJ+kvq3PEwT0ajv1My3z9jJNTP
bn4qLfi4XcNt3G78kLzeHC9x/1mbwAed2gyC6SxGdTMAkwYbt2+pV6B4ZHndo+rkG0qaH7Lp9WA5
EwNuKgfnhIzp7KXxgjI/ugFpDk32QSy5TIhi06hrU3m5waPCLNxkcrv3jxQGdiu3lU6Q4ZPajWcy
BDUGpgfykzOheHSrtO8cbHE1EfIlT6s/Vq5W/tchR/IAInwDmJVtFmdeuwHaGjLPpPVMzAaIAScV
hrcY8mjbcOmahFSb4QMk3eEocE+fOe25OTNrS8aBJTKsSgp+YpKwXdgr25PRbJhGZh8PgfEk9c5h
tXiyh3ewZOMdm7fj1roEXJUoM+HmxEaXL6MWg/HIfVdfQNTqxGRl3P6thceVAJKM7hTosa1RU9kM
TeVvfonJn1IBkNiBcPWgfUZWfAEeNKAGrpFtOLdxI7/6XouxtgMdbOG6AZoOqVKtWb7/vtI5sO7A
hd48JSHD/JQMu7yeClRypka5by7uq4xrZhHVc8kb75lJQ2+unIGfl59r8bfKfaD9ecdNBsTEBxf+
MS09UvkHxNgHGhiWVIrn7pNYUln1Zkq5IMUhTqJVvxhk378yA/377zhsD53uDqM71qZ7/Hziirj8
EvoVeH4STuiOLE8FRmB60AcAEerpPNZYuPWfPnGCWEs9+wQOUe+AmqSRmG/fr4kZ8CaD7jv/JBrL
E5/q/oWh6kghrSTEdwsu8InzazsBO3rxpkBA0NbhsJeuOEbo3O3wJlo6cB48rW2jigyIHqJaDfRT
7tX1fGrlhN+fIqtTv/iuOFQJ4Owv319PWXW/4GFNIyyq+eFaR5s+ltH88ZXZ8mqqIMru+eHF994Q
qhWUvO3r7DLE+7Umh8iZwUKcFN6Sk5/k0DLotqQbS6tdjMs/vTqdwvHzrPkIdUMcyGPoz2FBb0To
nxFvwVmuMHt52LH6iZByp/4G9cfSbd8O96mu+IBBP5uQbnLGDymtT/7YNLlclPxbmZ8OruAODYwr
NKgesS5duIETS8kRz/VnbYzEK99KcmUuvWE/yI8BQQyV32cU6SLcewbFC2zy4rI5ALvYXl2PB1//
IntpL25xH5I1vsfAEQK12AlldSbJRYR5dJEIt/V4LIczbnoYOGN1qIQ9m4Ti1Go5C0cJRS0aIVcB
HTKPuJjnnx+E+Y8xh9QpinjsE7eNDw443Hebh7nmRQuraD3ouYwedzxWWuAt1SrufYiInDD4FaMm
bs9iG5S8iz9ob1EQ4ATsra5SMtVZwpYjdHBhnrLaz2WkcI7zPldz1w+Osp/fK37vU2F1jtCDhU1V
XHWhbEjGj0JJ79Ll7y/w62OH4JFbttq9FJ36GgrP9vKoCqDtmA/smm51yJLL0AXL3JF5ipN/ekBq
UiRTHEHjDtybR/xvFaJH8YixoCagXJpow136eV96BGDRS2jfZFWGTc7cEuLOH3VOWS34tzMv7gin
RbyUB1vICvKx0dImcM7RFgPj0IAIfQ1cbWf0nsc6vB4Tui+RPpI/SRujXL/IS9eXwNopx0b24FV9
/0weotmDjbH92ku5BDg0hmlsxYKyvBwNcp7si+sq7kXJGk1ZlN6DcQ7jAwdB9K953MlARO5uiohz
0FhM16aKfsH5a0JR6g2K1DWWmHvuOM8k6UYg/o930eNJgfa/k8H8Zy/kxlzzpyn6Iygk6+yi2Jg6
UD6jtwBOtmREnvHDYepu0cwhvJfsYGn3/NmZLm60u5mQxPoJGPNrXaId+Gmx+eTVci6x2ckSawB2
ClDEC/dfOfb10npKfZNijVjL63QT5BEPTPq15sDgNzVM+Vk3y2x0PYW53ZwYXbalVigbkTxktc7a
7/aDCUDJo2LOiHKotNB6aE2JOgDRZBv2BgYMcmmyrNk+EAkVSe+9FwG+hSxq4KCk5TxyGr2U19YF
1qRIZ46XXCTh461blYHyjtw7PVf19blRy0uW1bD9MhUwqU06+ukKt+cWI51kO/+tZYkHZd09eU5V
PxHZUnPLJbzmF2d068zzjw7Iv+X8f7wIrpUfq5yy7MHmFWdMsG5c3o/lPXa3BaYJaLwcXQtL6TxC
1Sf3LZlVc1tn3IXhZdA2FwGNWBgokmJ8DaUzU2QMM897bdUl3KkWUEUtFCpO8XdPQf+Xoq4fbWsf
hwVRIJZ5X+iDSOQBfxV0+Q5v4J353n+U9hqUD3/hj6azJyXDSGm8OZdyh8A6EexBHVaqml2l5d+o
HAu52ojtIdHOH4yn5rEELoCBMTqAkFwWuLsYLHGw5i+3UmKAhhgkL0GRNR/7bWkWCgu2k8L60H+U
HEEATKBBbwSda1TjASqovkMT1OItmGQjbeGZF/0oEnLO2/g7LUaFTswQsKhfpkQQ+A1WvFTgtx9B
KvrEBoYRQROiiP7MKUXXbxCGP1s6Glb+wXrDVnE80Hwc4Q9MDpBNq1ShxxWLFGCOiAooN9eS4s4f
BGlx9/7JW8HJjfr+v2QODtKbyPbeVIjCa7uT0HT5Pe7FMjpQbRG2R8EZaZe49RU0czr+ofL07tFj
DKw6uydL/+WvW4SDJigVEZddlH1LYLMJpxpkJXmBM8HEsO8wywMf5HhaHheymvgtG2dkgmgE2xwc
BkTTOzZrv3wvVllyiOlf6q/FxfMsQq6x/YI/Pcgpa3fO3KL0YiRJS4brjMlBOH+AROjzXB3NQNJN
tUflLRRbWZ2QC/5BEplE3Lu0q6Sj75Cvr3Yo6L8C8//VcriQfzATlwuC4NkstEYElgP78OUj/MLH
mRVdTivlgDVE+CCNZKJmfk+zej8KkSOSZrjMGtlCEbH9tDIMgkLzmtei6EcxtB5ZKMO+KnOWrNlE
VM6EzMc9Ha9RQPNr/oa4RlDtjG+vnLSq6eCDA/sv6CwCiHWzg/JZvE7Mrxr0lFe63g8/uX0PAI0z
2HxNpYKRY5R3TgNuI8VZIIkswguyGXiWJ93SCPr5i+9juIZyWO5SHfCCwj4tzMphwk4ca+1NG6k0
vyGsLXL6lQn6Xrz6grkXSCvrOm+K5/hmaew2fAezSzWK400XERMyh5TTgHviXpU8mOphDQjyKa38
nG8gVYGLd+L23MwSuqELpHMRX4DSJ2j0MCRnctPx1FLlMlbh05CM9o8YekH8wf7YMrftNtQMoxBx
5ZWmPcAlUxPcT03Bt37KcTTEfZtKzQ5LaTytU9gcWfM22zBmr4Qk8GjQoyx7v5QHzEm2CfBLo4m5
kI2oRDHv/ArO4MtCS5ff3uQKLWrvtFpkCyrqr7xNJ9O3J1OTEcJXpj5bMm47Qy3DEr0fsafIDZ64
T6CRjmOunhIP9pOc9NK1fVG/27X+WKAZ3ZdjUftNJ1ZD14fwAdHqPA9uA1MV7uW07pPxC7ED8E1N
vPTEg1G/2RNGqavMuSrIc3885o2TjNbbDX+JwhAb6yV0o5T4nRj9WT6w+H82LzrCswYvlF41QQP1
6Ll0hm48a5LO9Ul0TlWwPDX3jfe1cNd7fF/RhdqLUxbVOrOeSYu77yXBWAPqePF93zFbycKaYrIk
vwLxBn7GD3poYn0dum/PdGn0T3fkmzhkVK+unBaJvAt1q0qllEdiHJBqDwiwSCkajgPfOhDln9E3
1FoQgeQANW4tmUOv3xhnv1E0hlFkuGTFeLfO+aizndlnp1UwRKJGsaiXiFbBahEZzXD10hufdRa9
cvrkmHBNxrdOsGbhBfg9zDAf85yU3nZCAPojC5Z2+jndvPzDLhLmGB0IJaQ9jJvsZUeZNYaZd9m6
I+edRKnxmmILA2SBentArovq09tCvlLC5Uv8R2RL74Hm5i6132gvo69mu+Fx+cNX9uYUZyNXbu4N
/6UT9RsLGQlnRHKUj9Pe05vPYIRxlkayJtOsr2R9nqj9fyCrNq12GPZxR8vZsPghrHWWYkCFSdLM
EW+MQ1z3xttLWQbPo0NC52wDrrGGYefOpuQdeKyS+TO/wpO4l8wirMtlgXATnVMnV3O5Bu9MJQ4Q
NrgxtOuILlADhkvUUfmB/Q+Drzs2xyEkxw+00yit6KasB62acH3jqw88TloHvbFzmPw0B5f97/0z
JTg/KxQHMfwYuB1yfEQ3vqeQ817k8y8o81GweOSgEVY/fgtC7AhceXBL05H8qbrQc7EgcgAeuIXC
3ye+dWEyxuuN320DbQrFrOavboefyTGGSwvWcSLtj4ygBkX7gC/VBcZMu90JgKvW4GNirIuBku8q
PqFu5PolPicQWiKywl7LMEaX2CDUXfRghpo0EMTJSE9ZnemI4NDuB03ax8QBv8QQdmEIkmvcOW+X
c4WevtkPn6GsJkIsUyQyRzAedmRtyb/XzZ6vptK++AiBOieo+q/li1e/iBfe3ttJn7l006Ga6BNy
K1JFi9zYNeiwXZ3J1h2xl9NIYyl73TCwQc2eZc5vrL8bMMj58KxsAIsgV4jjt8XOGCUpZE0ZwdiT
2tmfSJSYPLdXrgQy+/xc7X/KI1KVyjsnM3xit0IGXJMcZhghqAeVV4mCMHaqdHKSBlPZv6AjwG6n
aJLTodBjI724g4CIAuYslNS8nFS/gEn1im7vXbF/gpHMCF1ZZtbkP4/PQiYJpk3lMb8fgOyA9KnV
nJhNwroKY45LSxG5n00y30EaVCOVprP0khYo4dOjqPWUOJcszaN6nbWp6ZMtVEpAXPFRj4OIjVQz
fsNCbtlFOrQNsMS/ZZVIo18WP85JddBOsDpGeZD6zPeuKJDpRa/ys9pZGfEMErxDOx/msSu3ce/d
/Ld8N7UQaRQ3F9Rvxc+ok5tyCLa7K1zUm3Snf1dXsg2Xa8if5fNoFim77a7WQ3BFlsnxgYPdz1C8
ioy2qHtGNgjNYwpm9wvc4jhvPB0Bi5NqrQeKrjajcx+xI9LU2ImHvTi1g+xHT5PjYdA30UClEGjl
pEkCGF9zTYNs4uYg4KjihqXK0ytXO703QT2etcTrAy8wKAWaVmsTDvhcJNi1xr7oJ3sBRdjAHG0J
lMVaMtUIc1cmU5zeRjPMPRKVaY+FynB45Xft4NN6PsQJ3Rb6Nwtd/swQwRAMB1bzC6VncchCcyJM
VZDj+qYv2PeXfInoGK6E4IJxVk5qt1dyeI26YaZc7XlcfxRJKMwW3RwRwtKWwk6RbbMrNs+7LPxE
+f8tUGdXxztfugMlo2e/DAgdk1Ji9htdnQT8kv/kNGdtoIQZEOdBU9HxX23k4BgcJpQbmJGNdk80
izPTbBFqvkCJKtrL4O55pWTArUnhv3Jw6KRY4eLlKwim91vq6OTy/N94HBFs+Lzyr2/R10RJrPTR
rPFhPfqHlXsxoxVPpVIJK/gB6iEiEcoLS2XelYRUKvF340NBn/d5aKu2s5FlXU6M3ZyBk2/u2vy/
5tmQ2b3ShczDl1c3p4JViEeWOjlIzeWimX7D90u21V4u0us5JLX0TK2pOGrSJDFx/2n1HWAd+ujR
Zo9WfVd603kAo4G1AuJNjaLRUmhU/6CSlxkF0aJIzyLHLf8WiHIjZ3OfWlkMivq8zscSfv52mw4v
kwCvdg1upPNAHaBASOhLFGe6QTR5Xsu08oj+w29BaJJ0GuKwetfXqOjpOJjlQxGQRHjrV8HNmEmS
sgB9lnQtJQ2d2oPRgrMkO64MrDi8EdWi3MjRjJZdKtko3d+NIiEIKrAdu6cVuh7zqsmijFZamZM2
lWolgoP1I8wOlR2BqCvm17ybaOlsgI9LgHaaUj1iRxvwTnaw6I5J3+bFAl8IBdUl88cPDEwpQEAI
M+VLVXLJWKNboeWP5rdGTNgccNfRSfcz2ZmQdSJqtl9+h2Wddo9P65jE+h5VEAtNOCEyhu5uE9Y+
A8fI4yWuMvGFhPn+Njyb2GrxzlyUcP1TiIHUMCIlxuojqNjcU1HL59SWH7T3eObhrE3QLQo/owpc
/++q9Qii7RVb9dI+9GSOWUxX3lSqwXrimYQ2S4jazUoU7Wdeoa06esNR/1DEYSL5rEybUEjycr39
So8erbekF8RlCfGSdYePqDUFKq/BaITrv6roH1FaIBXRi/sC+ut1QESGAWEFJWkOJOL3suk+D8f9
ndRMXfGxT8BcGaMaImfDzNKJp6IR1y7V+oY8+XXYt3SB70/kXAkACdND7tLl31VnIbiTqe0Lg963
niTm2dIRAAOc3DlXbTrAvWNgyDmLAFSpSJaXBFVJhmVtJF8J6AxwgJ0vUC1FpxbSLu9+vyXM7zz0
ZxXph9ndTK88/WagJ2IwiHVnASsqD8zL0qcYNK941PRmNZ4JLJHM9qTJ2RUYNuq6WjdOaRmsb5TU
BTasmd/a5WFtFcTL3HUUeTdPUhly8fOinhQGTJ1wn5GSL68qKRnZnIrRl7HvUQin+gKGnKQVPRyw
xuodXlIAlC94ZtredlKodTInQTdbNl+hxXn+OadwOqtXDWlozbEHviBvqhhME5Wgnb3BrHKKDahy
dsA9ctYolvsRovX0uCgr4h+NwO9ncdRD30ngwLnhvzoM0ihmPg/e31fcX9TwS5Wli/oPIYvPTHXb
LgglUdvLmx6HL/fl23cBqioU/8+Ni6FST8+ZzyyXzNvqTj6cWeKnC4O8PcJN835VAnbgbvJA9poE
FUg0xG7B+Uy92SD5gCv2rnR5Jan9ntRm/s6eL/aVpZeo2D8hnYHGGjPMnvzTEVmBFuTjnhuibzVB
S3ufwgpJy291IQlNWWWszNPF+6c4+v/mhCyk/9EXdXr3FKvA8S8nKRfoXi2n31Emz0oveebeY+3e
rzyTA5xL7bVxVyY4Cck9yJ/YrLrl0B+xNxU4YLpPMvSkE7gfWnzU/8TaTXirMnuueY1pd2BZNp79
xjiQoQTkkbmJP2xdU8N2oy810xKD6FkCSEaCD5k3IhXUgyGFlBOnIt0+E9td4c20kJAIn7+5JXIZ
C12HNYtT2DgZ//BocNmBbYw6Ddnz3WjQPmA19Ray+DR1Ot28dL98MtzJqwfpSU7+S2I+NZy1OfGF
SPvX7Aqp0XW1xwjjSHV3qE09yJt8GHBnuV5ZmVgmdWEXLVvD8DyPl5R2BFGRnG4rWDFfZtJu+vEu
eL5N/yjSqNy6t3QeKfvXkP9zyD+abybP8u02J/oIOdbwKwZjLkRWI8jKhGLhZk/t3yNDMwozjEUT
TWkWvU08zIT0jiROR7PwSim3Vnzv0e4ysju5I80lVA1BgrswUBiUNEr7OrlOPUBDGFlzXPrwNcjX
e6aYaRR5SP96Q4QadWLd64O6AUXiIzQPBGOqaEGb4G5Q6lzJ3ZWcX9Ut94GeIpHjnPA51oDNmToM
PAvgIW/gqX9EY4DFVat5EuDr7IZY3Q+LFbEkS2hDkaUlLk6lPiiSvUsaXHCHG1ZD6EJqohY45rOu
A29yNT6+warOPp+2Wk2jfx/1i5YZXBW64udMFBjtaQn9oPuCDFA/YsdxT61/Sj/uSFkWd0OzZ9uE
aysOVmMrsW9M45jeTBdcAofSCEpkmweh30Wxh2DcCqs5lQ9uYP/esUeEFgyXvX/7u0H3ZY1IP2Jw
KnZszNsPHmHGBpeBOZqh76sqGpFTiVKfGuWtgU8LBwryG9yDQGYqX1cpuP7eBD34Mt3K0V/7JgUc
uV31VWSsJjnkSmVVInRB3m+xLzyqlmaIC8D9b35igSRahVj9iIauOwWR/8IYJwFMMyfvjv4xCoCh
PvH2RC12kCLrOLdYiRtTCBPY7XejhCTnzl1I0LcYp+3R1CPPWrx0Twwb9bZqLIiu26ZPk+nFbv4Z
+XnjLM0N1vpr8VDIfcXRNemuGAbjgAnOYl/tLwTXrXHYhV+HaoELr2I/MvCaAvbVmumA2xhuVfe7
5zZ8sTawCJq3QlvqjGDCknj5KkHjS7LcrfCR9aZkg6vW/cCQR6vm2F6fHOQKgjGkYwH29urLqlau
OFEogpovaTtqRT/zA9NW7hM8pb7U6Bp1g/5yZhnXgU9rl2MDLen+dSe5uzQHK68p+e9YpmFm3Ill
uLNiNgPKw2U+2HebxJajKHtXmnDboUkAd/5d4fLjzooqUeRG1mM+uThbh9982SEs4ODktwOFfx9b
OjAjAHLTtzq6OauuFDicFcCIUm1ZHmRh+9CBkZjyQ1TK/rTi0zaZnEV/u8KSIxasAi03j3en2Apl
G3v7DZefFeCTwCBnaqTV6GFx4Ct9GwUAHw3NLSawULsGlMZZ3nX6CCVG9ecyhEKCaTXDwoaF5+tU
i7rqF6Biy7etUe3CD5qdrF4rFAVN8AEUTBzurQNaRDzCmjihsSMVZqMkq4sreJP2XAiko/k+Nq1w
n79i6dIFkWIdmKrElPyi8AtL1H1klHZ4I0dwoDJFqBDLyipgFqnfLACqOONPucCHopIJPhjl9x0v
XxHSTPgYrHpZqfEeAeKVoPhtwJaN3PoQ2Yyc3yp35VR/8EE9+Q0p3auFIHiZlsaTLuIhMXfpsl2m
ep6++TlFCoQvTnIGkD2eZed46AAcoWa9SqoCwbwmuwA0vW2n5Ea+VXsZqx/6YYhfzJv6BBCPdXPV
qMfD0+mEsn1cYURUwd/DXjKwOSnbyWg2HK4Z5y8jfzCTiA+A4nnv42AoJlOYCISybRYwOmf/YOtv
vf2sjBu0vJZSSp7trtt/z2OTfidebMj0xKdLUsO7ZrsWmgFXXC001DJkaraAS01Xto9hrNW/Ua7T
Ri5iIkVgRqtwDMMCa4Odmqx+mtuv6zIb+CBYnOzQ+YK3fGzZyLX3NwHuFrvtUrzMvmmF+jRk+LbN
td5qmEOlkBmHiRsbxP5/BIqM92YDFMlwfNqBvOfzgeYQziyRLODZHgpsg0ODr0afm3ZitwSdlG3m
XOOQ44Zupik/XqNMuftcZoGxgTUe2GfT74taeoDPSedqDf2RQJi/JPV6wYJ7Cw8FqUNIjRJoGsQk
OxHmx9Vs6aZE3bkIyv2BTljTXvIB0v05V+ut7IZPC3zSeiy20904S3rkeVubL5lt3oe6xU53W2Lp
eWd6DS09rT/ihKp5sghUWufHZ1Unv2OVkj0rEMxiuv9wNvcSZ6UTZnuJcw+wdq4aDmw+QfF2I4Gt
Geaxc5NsfTC5zNYUab9CiBRMQ5Xv5tglczU6mzBEffmDSSBWYxbm5muirXB4x3v/g7lRYCjpvPt/
xGy5OOeofCVW+GAqryWW/GTTvvY9PDy8N2bXd2ZNMCZ9E1uH4vrSOoaoYAt2/yd0sX03wFHr5M1q
Llc2xv9Cmodkhq7Fnn5qV3c2Ef5l+lQkSssBiNKLpc1yBD0Ocqf2Vdfiah14xzkGczAm3AMKgau1
h838Nw4QHSDO9hpk9aTuvpx3LeZdBYBFN8wh2WPK7k11O/Odk8x9QIklz0dBTVd7NLaWQ9Yrwj9R
n9q/OymVlLpB6098Y4mp1mCI2A7WRxPJqBOiUP52jDz51MudBwVykkaV3SQs4bHXJKxzSjS3PUly
RL9Qk1oM7xZzDTRsDMqAUbAFbFBVOXb15fkknt6A8vlGRX0EoidIVQTSulWZIiCkAW6mmGyFQ/ng
IKDIdbWxHsl3bxxsRLUzyHVgQmcUN38vJJeEi9dMJNJd1HUlMOvnYK2oec/EVdvel/Jdtr340y37
iJZPGr53P7u5cROCZDJE9sUCrOXefT4BrqtRLkWCj+pktwJ2v7xGqf8jz4NeaWaAmTzrNOOPKICa
dIG8WTen1yb0TV38TSD7b/NLcMw6Vp9voRqV+3RlsQrydsk9LsxHFd97YOEOJhogB4cIL2VCejMv
uJubodIz75w1CkcW6AHhKUA+VGv3z+0Kt9l7EzrC65FjJu7g/gMjTDwNE/dyYS4ZiVb87pDIH8n9
dvsSZ4mTGY0+NojT6lDGbrTWwfT8N8CFDoh+H7+VOesidoypPRXifHVfTutvdJVVuo0VBEO/b3m4
7jy0v0hB1bzDAT0jW9gqpi6bJgtyLmG3mubdiuQ0bAYbLjRkMr/CGFfsrDgmIBLJmevsEIH1oyFJ
ROMbP+/LylJ1wCjoczf/LyHZuBvVh4mr8FL8ZFWKzgl3zI/xxsZJWBV/We5fa8Jogk8lFvhXllwl
Wz3QORRCdG+CsxbuyTzqCipwaepjpMuUHo56efadAtrew5YkfYpzJMEP6uKHcC1EzRAx72I05vqU
i5XZt1PZrwq050DnJpiZmub3ESX5FpxIFspxw5SJkoijwvsQhPnA9AugzqKZIbkeCiO7pMDSGk7H
VzVG8dLQQR90nIvr0dVxaDgiQEW0d0SWpxzs04ML9Asc/JaEhofT940qKPjzehlgFgzy30fCxmUl
G6ihrhGmxrn71lsIFMqAHaItRofkQcu5+sO0/7tWszRSxkofqU4YS8ScksaHdglbK1k9ca3AAlWR
SySR3NB3rylRO9xC+wHBDjeEnMm1h3ZxcXvSOsfp2P/WJHsCREv23XX8WF68oh7ExKiQ5kEoH63H
Tvi22eAQ6wHwB4GMLy8HzgLDy7C8zZx4PK8Wym3saZmAZ6KI8LHe6onOrYOXw1QACbU4ncUDINnW
EqoSqPqH+UDLYNavAforsMRPtTvJiDBQKXGN03UkyTJ7OJETGmtQ6OoHbmegl9jAC7+Kmks1q6fX
zzrgiz6ytSOAut0lJwt5pIdXM6OBIJQNSLp7o0ixZIKgcGhKAZ4JcOHLIvAMvudCsTukVQZIlibU
bv12tnOt8Ai9sIidasNpJVch9NuTGKVHwYnSnwSWz8W0Dt1DZpTVSliTHVnTKnkQdiaMMNI3V0rx
2jSL/sn6EjK3++c+WA8nshsrrrF5Bren48qtV6FxmIcXf0sE7Nn9xXL0cyiiWQRDGyKgQd4MzXAx
fXAg9yWv2JJg2Luo4NZaWQbWQE3lAhfE7Xefh5AUv4MUh8VtkKwnhig0linw4rQFSnPJAZctEci0
KkgUq/pBxY5BosxoDCcrEKVMajcEpCvaCqLiTwZEqsiGO0bp8YXVzJkPqm4ZGP0ziHtCPBp9ZICE
mjZz3YPBYIsJ12RMbQQ9fJdhXMAWn4YVavZtxkl8sQDUw3hs914DBEfaKAVLZM4hdwMq3/ZJEMdQ
rZYoXtto6e4KcSnwf9A/GIrsr969NDcoMxu/N+WYPKiGfwjfjfavSGVHrxpO4j0/T/+XFnHMvGEd
4NAH6T9My2G2QrKLyX8KwMcNjeJsA63oN4Nd3h+puJQGEowRdRAgEN1bQl4mOuT62EspU7IuY4Sq
sunZoTMiVnwR01V9wVaEE8phO2E2UkePAP2t1wpI/kmeIHzUP6D0MR7lIUVr80OYZJN8oxebXoGH
cHLCQtQb0hbt+4SChW0NCOL4ltvMY3GvveHa68YTJdGUpv3K6emrnTa9+KYCR2hxxe1VJY/FY61l
74w+27FWOddaJqofydshafqDN4WAL0ixmLzsN51L5GY2Zgq8T7/e8h4jZuSSA3Vp7M2IMqzDUxZ3
Qd0DkI9drI+AYHg01Zyue+35PpCGQ1khevPUMDtMuh+72YlveRJ690dX852njwLXJem1y19qBe0F
01jzZmgYk45Hv7mu2ucdwtxGfpVmEd4Mcn6M2EVj+hBk0ru8HHt4oPgB5CpNpA0KBFSTmko+1WM5
uyEERAH98eN7WLoYfifUXo7NfmLuWrbqJgnWqSfdH1U5aMXP/FNXo1APcVjtP3dJH71lkaawqVxy
2FbIqON+DIQswJ9FdBfo97XgAL8Us/We6kI+m2nlh6j2R1sJ/caL4h76mrcnnHkvsgL4OeR2OZKo
CTNEJW+bMeXmLvXbLatnuG3Z6FlYunAKktWZtSIoVtc1dpRFSt7ZnEIurWdPzhtB99rOSVwPsM6f
+t5F9j5xsvcid+t3Gu6YlPawvoeQJ5tUgWQel4S1LR0MB8+JTxcLOVHQ/hiapu6u+i05M7zObicC
3FnnrrsKu7E8axCIHXJBY8BwJ/7Ep8ZMgYc2aX0GiOiKOXeh/v+m6xCNkbzDEmz7gvQVco1IusPG
7zqSr9KAVnmGEHvpCB7EJZKspJOKO6ZlWwRuo/xPXFYQgGNqAHDas7h34qzKAZflsXI+HD77p4dU
5oXLQxZGV42KrgRnvYpAgRMbtMRw3X9KE1DTfMb6ddkEIavaQA+uhqK0bPBDP2/+zfb83mIFO8U4
0mGgbXmHEMyBwq5uBTBdDuCfTEdo5rexWgCSZJ850B3NxgS/hCTXSFRH8dpUCN4vGVWeDvXfvnYs
l3porUO3QBa+EervrFXqc3SPbSRVcqoAkW4SPiypzY3bYyKMid45tZ2+XmQ7JJUgecZZAP01ySUK
VjzqiugGJJBuPYVsYMwc+EX74rG2Bgt3MiVek92XrBGP2gvkslfJE7TAEMnUI2NxuEyPYF/cTP3m
DIsUy8DAp6d/JtnBxzmXdL/U+TLUYT4Qj02ll+yUg5UXuEzZIhK60TChJS6dDMiJw+/bN9tt9tXh
uyIoDOZalz8iqkzYFYq3ocMBOQzicI8T621usybL/5nk8m/fuprpyPaMpnHPy6TgwvqO8MRRWAvE
JRNkuJVZX+dWIz1/rZbSqfoj/A9gnnSUj1sM/sbYMaanOl0C3z+yTWYkWNJswg+8Q2tPxvZfgR5n
52j9uTdSlpBFPFaFCh+glzNPUKVSq2SrfIu+opEa9RJajV9R6sn3vcZ+P9DFHk1oUO5k6b5nRDao
Czq9M7/QBnF74qWje90SGTe2tqvgD5NPyoZTzdAulQlo5cy7fkDnt0K69VRG6N92Gy+GVXXqehEq
jlOm3UWXQlKgyldteDD5Vw1moaZctjm0XUJ7sKc0eaHhb5j2ffK/mNpIg/NBZXf9jOp0as4Kt+/9
ycbMh88KNduV/4TcC4822xHCNNDf3mZ1lJaUU+D5zkMZZT1vAjW+Ja4RJjFSd0BmjoAg9cviUWol
POlGq8zGUszZ6b5gu0LqNhBcaoKl9ZO0D3WRKlGHbFk95qUxgMgEzOirBTw+N9y4vDsL25D5LGnJ
JA8A+N3lFgH1q8z8U/2wbhEyzDnFVTgLFuVh5hqB4reTQNlMUUo6+eDSWN8vgjLq3qhRURUgjmc9
TkPKp7vJAWxq46K9UL1KZeLzGBKAGTp+Z4tFMSeKdOn9QVWZT/A7ctoTEnrwE/SMS0usIDDN4HaM
niUQaPbJXpVpEv080Pdy1jozUVaNKkP7ZfjmtDWwVMHKctYuvUAeV4vncNmuEqecoQN2t7954syk
xrdzzppE3ZfTKx4LjhuhOdsCeCCGVhjHHu9gPADAA4mcDBSUKZYMlNYoCBSiwHodFXRA5ARi2asZ
tJCAgj65d2Qfk4n11+kHzYE4aAcWfKr7I6yY9qV1kkFWOfwlMogtHE3aqsYfr5/74yu3cCCFoXrn
RO8WbaD7ZHJ8FhGTSLSgB9wt3nzhJoyQZPDKRVzY2IodCZllaVvf3k9BmF+68q0jZBj+NdVTwBTf
V2vN7QWMQJjlwgzsRBRTcCv4jBngEz/Gw8yn1ejMpwDTl3oxZS2gnuudgebxkcaSLknxNu2eQrgO
HYcEf5OBx4ldP1auJt4cdPOv4e+ZfQGb3yw5VSfiPmhcxBae2B32arO/j2sQICf5d+C4NvuCd/Vf
5qw2dJ9K1/7H8OIexyb9gjohhfENVmc1Oo471jhlAIJQbrGhNoukRz+yU+y4jOYi3KLRBLez2cSq
PrRL71hR7GHhtk7jcmEXTzV5UWautrPY03C8tTk7FLjj/rEZB0R6ZZDMeu0n/1puitS+QSU3f9gi
NNMxD+LQUTuRdwl4zSrye5piRZ2OGZP1QqZs6i40/hItaJdLub4J7zTmo2NMwRUcA7ZlT8ucF69X
J1Mg7+6xzSU1hEPo8ZupimNDq3bQHezWwLPtf66gymHIKzDiEqLvFRrOCsFoB2tSPhdO20WjCqcc
z54zZsF0gGv4YSGaHm+NpJKFXqwmngspDo5399O4Nd9IAYQGdxjQ+KlMwnx2kwybn8PfkY6VRhvB
qmp+4j1WLpawVeRZxlsXM2RYD4wz604mcJKko4K7f88B2MHrmdnhDHVIRK9zCg11BNUYarxBkHcu
UzWEJnS15NlSPDcSKegrDVxcsPvKZDJ+1dNiZoXSHHUx6SptMD8p/rIDLyOV708vmVpR4Tu+wrv5
UZOvP6PYsUYnPyJzpW8jReP7LChScS0M59B+YG9Ef/58bAyM2+fbjztp52kTEDpVQi4+QkEu3Fav
o3x59H/pda3udhjpr4Hnv9qu+CJA0POoo6lcSSFx4eYSSsp4dPD5qlzKnqvmIdCGWw7aikYV7r38
adp7xUro25O4RLGkR1oBIHvDR43iuJMN+NotSDTuV4Z4uP8V0/Ki2WI0hehoUCqIRTkTnxSkXCGJ
RTWc2xpYhk//Dju2PLTVyAzHq3JYLx2kHxsA6Tz6UbhX11nY2S0sp5Gt83Y9FKzM+5MtAYWQdHjX
zbZ1qmgB+pnevwlYwhhy22wLG9M+uXRJsDCoD6CG9J6OmZyfJQDy0mPkfpTg8fPDichyi6COLQIT
m9ZQe2skuBjARyPK82Y1ERViiW6wVTfHehTGsGbh2ocAjl4PFveQGVM5JsylkCw7zZyuYytpk76w
UdDVcZobpVsXwSr7Zv2M0DzR04v9Jpolnp2/mqnsnRHSnLu94be2hcveQOXdzwakCZIcUdLA8RhW
l2Z6z6WUdar+soI+5HfjTDUzt+Ou1kAio2cviZPqeUIgLK+LAdhS6fLDQZTkpoicGzAaC5ZLW5Yg
rVgWudbiW01Q4Lah93AFghnHDAWGbYtVXm4FTghHCyecGegiPgxe6xBthc7iOG9wJpVjShW9CaBy
HxsdqpMR0pqR5Yt3gvkNJywWqX6656G+RLKHpxoet1sK9Q/wbBN+FUvksPF0lX50xdPnvCSOnimy
/ohUX9yErTW7ZvLgrACBPgU22fXSzekKxUggjz1MnbnY4QzeQhAeysli46GJT59vfwTnyq2ZlPjp
lpyHVS9AT929Dno9JPob1pJFAP9x5Y8HOAPWgO2gmA0MaK+YrFcxYjJtWEw6Gy63unsA8fLLv7CA
A8+NL5imWLXPO0tGCuIgeflkPX1Ln6AEdyxAGhR5mwmU+4ZEBPqJP0dakipFgKYvB6y3CnJXid09
FdYG+svFc8nZW/fH1OItqEcpVanWtGHz7dXDgPVA5VlRNbL3by/2pgjcf1v8BpwjK5TKtGlUtXtA
5QtJ+Y1LgqwK8MYvGq463v/799cGrf73ktTHO0S2D5Tcm+iD+/xstueBQKjObKR/hQqQ3xzVeSaG
D+htQoKaQlr/3Bf3soGHfgfFZaTtI1PtHDLgWgjMlnoThQzPZdWcHgm6KF8ojCkxWz4NZsiOqxZo
853EgPJIxKdXoCsXLI4siiDDRr0QQH5lnXxngfDxpGtcE9rwmXFZwvbI+GNoC0Mh3SKF4UNXuBHj
Y4gECwcIyYT+4N/gfEpWJ19Azov6TjVdf6sfWwDgmOfwc1dzapP5gQuqi/HlNRlkbNhIKcjMU2rm
l6XExrpRk4UmxxlaOnO1bNtbwaYOf5jcePh4JREBHpJqDVSJ40eqpWkfTeZ0nQ4b5Job2YDKRAOG
pdkRCA/VVW1YZ8ann4cqyQ2Iq/cUi1hX7vdLmRe3Opv0jYSyXrOS+bEJLSLEMVhSt/57GvWCppJD
E6snf9iHg0/8dJZzAVq84ydeutlEXJyWdHmK7D4BpBGNihmp3U2yn338gPWkMnLfxJCKfz/Bj28u
X3Cp9D+dr/2Ij4CthaTLEuaF6CTNlJ7bFLcMaS2rExtlCjFtuusnxDncI2jwSwrVJwFp0UP88fqe
vcEWd2vdJu2mbsfawhVozJCSwZIEL56UJOc4zZDXAA+8x6M7CjlpiU3xdxbYqi9ItNVTd/hLCLHW
LwC/4TppEKNgU4JDOMbGaCK2aNKYiAStmG/LpGSpyIgqlOXUsq+Kf98Lz9x1J+tDbGSgWI3nFWbs
CBup+YI5I/m6FTf8aw8x+VyEGV15s9A9k4a/mmDN+bv1Ctu1vvlWSS5Dtyf2wa/4LVivpy+IEG8t
M6GQdB0jXSTJOryVlJwDT4gdUqiaqaUwPPg2TEsW7IyzpRET3+weFN/J4EnMuhjfdJKaiXbfKGY+
pT0t7TJ1nGTcCANaAdYrP91rPbXkxdGDyJFBO/vTKaPYXSWTSVe92CqGSqsl30sYzdTx743UY6jp
gDZxjM6xste7UsQajh7uInxy6JDeNmaMV7Rv843YodHHftK/AsXdoBWlb/o9ErZMAyeyFakPq9k1
GkHdp6MCTVD8j9CDSXhp61SXtMTnr29rIoiVHJ1nAyOuaVJA+PxZMCd22uUpCTIn99C8gvg4ADH0
snpvZCgnTRFIBvuOpzA87lyFEl4hQOOMpNV2LcuuqMiY4ZzxfGYz+pNDOzG8SPgfdgWNynQ54gcA
3PKHO7gc5DBhkH+HQkbHLa1BNErb2cWQC7bXUJUY1yy2nieSskD581lJsDph/DLwkOGuKyVryzun
QX2hXwguVGGkqEbZIt20Jxjcb9cvkOpUcnNB54YC+3SUk55FtM9JH1quAQpVIlUE2or7zxHy39Z7
lHNt3ZT+HqZJZ/EoJ+uXeLK0LUoMCVGKnIiAoWoUPvSA1pGBiHC7ZsEknhto86uLIEXE+4yjD6Yc
WJzliko0BBZcW/Dj7xINPjHktAt29IHBwPtQWmhvEtntCab1WdvsLEuHztTkA/kyELeaewI513pN
5dnaK4R6e20maMQKhS4HkdKXdSIRti8w+5sASVHVSmIiSiSUhqR0D+bP+4ecGU/FTVHUbUY6T6ez
DFPAKSTEe6Oe3JHI7pFrHnmafhoEk4LkkChLxlUnjrtI393axxo4PUjST62fJbZpS3kvHSKeNy6x
BEb3bzFYCubJpbq53VpVgFcuVjqdK1YB8s/PpF+dJil+OTIxTMO0BB8r4Us2IANs2A4Iy57XGinV
wM9IvOH9eN3PHB82j5WqV1HNt7sNhUbnHqNDn5U6nJVyu+dMZGxF8L5q5faU0cgfJ54f/6dncc4U
4NnCT3xpy7iJ8pPhyNJ7f7spXkfg1e2OrniN8r0I4APSjbb6KU34Jtylm1tE+z/yv7baTJegrcjU
0/h/+jrmdCm3YosD/z+pzAnLVNBRfq9Hrx5hFfnlZj3LVjlun3S45zqHQ4/bxjCkJSyZA4EfKqtu
iEMqnOLopIy8LF4jSUVr5CDAhZcJeeEYymmAHG3BNZ4XvdXrvdzMbBGlsEhDv/si/Omqh7W5LoqO
5UGdKjjEOory4hxZSBW+3nyJm/ayGEn8vx77/XsMaY6d6DjWOC0N56Wlp6WZFFFIHxhM1+MGYK5z
aa4squYUyDx3nav2KxxDS4RphSPxd3lXcv/34Z6bptHj3N0SYdfRfUN2tgMpVeN8xWtM3ezkeKdi
m0RrjXq8EzwjodhojBsBrlu5DmgNze5qZs5lQe+ap6bgXL74f98NpshVLu7KI/SAj4h45STWqC9W
9j+kWHHZwIOv4DJZ65zjs7bbBxFbxpJVAle9H5DOJLfYHp4k0qxjZOUCIDBx9fa8FUvqfO9G9Ryi
uHDML9Bt4LM8oYdXdUuQ41P5lu62bGL7DntOIJBFCG3+2hjx/mi2k+quWpyzIOpRwg9Zl4Bwjezo
gpkYbwb9q7VNP5DZ+sjatUUE0Pu9FbWEuZ1760JfxX0Pqf7dVFCzhj0dFGgaVf/Bw8tDPqTQLUFz
0ORA0Eq2smwJTjK9JXhM3SRSgr/lzIs/hfPCJ+O9TIViGUrTpo2uJKh3PPkBSBoBbdmW1rf5WT0w
0e2E7+pPGCOTKfYJKko+4M796bJyDea0sX1L4cSECX+zznKTVxzLTO7h4PErR57K3xqPLXw/ZTMf
WSLAtc5Ju1SOhou0SC4S7zTcN3rWnSClS6Qbo37lhsaYfW0AxT5RFT3PNNLafldc1K+vqu0bkMRf
5nhzm2MVAmRUpJweaYLTOARrqACTDlur3wB2/ofjpkb3fW4VzxwFcOUDdgQQjGrnBBLrdSoCE1vE
IFG46TyZ++J3CgLpqxyAhHkg6otIImMtI+jewh5jF1eq0fXlqAUOxPNR/lhVlvD46E53J3KKOII5
wOiylZkN7d8O3vgBxpqFEZ7J5hcK+IaHWzUfiqc1llK8ky6tou5Ii1+IboEfjEbhZw95eJQLSCmB
0mhC/zqTHXachrXfTwfImtfjCOhX85wi8m8RV3ZCNprG/KL4jr8hseVbQXNN57rK5t4/mT9pg/mW
P1N04AYZlZfi183FeQw62k8lAMd1o1eI4tkPtjq0bZFqWp6WbRPXJPO/EtzyChY23gvuQl9wJeW+
hD701QC+thNXZKYqJBJ8CX7P/3c9YHomg+sAdpjH+B9sFur5i5gJAOC5mRxpyv0hyY7GDuGiwcX6
SEXKxYAY09iaVGi0SW3rkt/FJ6CZAsNBUG934SUzFUnV85rwjTSes12baj00Kdkdijgz6p9HWPk1
MLGBl89a0d0+Pf6nX0UEZG7ndXwOnyJ/+T3+8GaglzB4r/2PosGpZrN8sIB6jnIw7m+A8X/iC4Lx
iXFsrcVMtTbQ4z2OO3/wtLX/Hmd1U18Jf1YpiKvPDuL/ArYDYz29wnb1fUNa0jj8HKDoaWu9eqvy
G3cy+8eIqv84tnb+jjSfx+AmBMUR1SFJtLRDCpOEZWQYxykCi03PSJXQIQPby/fQTuORsY9HSlaW
LGR0CWgses0F7LbCa02lcSmjbPreiiCHUEOD64dSIZx3P01kPyZPFXVS4i4KfViIbSDwNZ7L6Q9G
vN11EQp4lZYGS0N0FW3CtUVTFvVpdcsoTInbO56isRKJwwjsnXgXagHM7i1nmgp61iDKXd1wL+xc
Fi6Pf1d5EzTYcdbyuF6hEUDo0lo6niGQ4XQLd3dQAERLzQLvxaZ9Gavls1RxkBi20DgwdS5tz4CD
YTvEATtD3ySSHcQa2mH6Th7ZzZimJDGicrtKNz1Hm2MURuJPOLMl+qZZwZnLPeHzueTiVnq82Oj/
TQDVzna0uOr8K8uE8S8wa1JebZ3PGnhRDf7Gv0SkX4vk0RFBagKWfKzK4MwpEtjTkMWNLzX/BjtL
0h8xNY4n2DixlXy/Mw8EhMzk1LhCUF8eHUVeaKUUgeMkdTtyoyq8xPFxYOdrO0/5MtACZ9nnmXaU
tAm9LMH0wf+hod0GtyKU/FahVdbaHXT94KSVouTVETsaKBVv5dvjYoIIBBgq2nGS8htgBAfulpU4
prnSOniv0vJ0GOTRrUjGSl/wccmx8dFyynOY+/YrykLhZvWpfcJI6HG+FffMJo4UH7NBFKul+2Le
01CtIdRLis95/2l7xrmV8iMKbqA/xUTjDZNQvSNETYfreSkRyVFfq9rz70H81wZWE9WT6Kz1LkKO
rCkNdo2iynAZAMAy38ksxeoUU0pkc9QK0Qwo8gnjzy8jAjdb3ZZEKzy2vxgD/HZfLXkiCTyRhA8h
1c6StIN1/ZR5oasVA/U0aQR/mCLkSG1j6u8hRpUdJS8uYhsautequdFfXZ18ACCWGN5zQEPARvn+
lcOq0LUFUvLdTFUM+aM8LUQnsGfrG6uApvjD4J2+sQVAhl1+nqXGvafnEy0kR1MRmZaJdTWtYInv
KRb5V1+qa64ZUVGL3XPSvVZp4JBTU1F1nzYii2OmBBiJdIrxyvPe1gaQ5mIvQtoAiTilo/Gkfr91
3+sooglxikXF8VpxHqeFOjduUqod+cT4ygrzFHT2BfqyV5quIoFpq+KX6vca6uxTySkEBN9cxglk
3GcDudtoe+IVOA9EERUyvPa/y8zbYMUnWp60WM/YoU030wueVuW1aRkysNcL7Mz5a0uP01eFArn6
sthyVy6Rf8MK5RFdXi41x1l1H6Fy4PeIT6cdJ6jeEaQTeBunyvA4V193IAPkpG1pmXQuFAeb+9RB
Zr8qjc6sJEIf2QFajnT++OjcwIyLU9YzSMX1Ue/cucsjCS5CFuX640XU9Wgetrop3MTGSLzXRUpL
aKTzUgD2LKbF7EWOf6IzxlJZVXkWjP+LvfPEzpKyeO8MMPFbRI74VS/lUBOIYH8+0zzwFsXNnYAk
KPRH32rehqGOzqMZz0BmTklW0g195EeexIwFlhw498Ia5rRBi8Z5TZyzClBZHXPrYe4A3RUMYHJN
bAxIypGDLCrmiJfCwRtprX7cVP3SIkJR9zkAvFpmVjKYwsjUkn+GDykQof6RETMyrYtDbIdJCmAv
Tvdx+/IZOtPUDoZu8R70v9dm9kX5YXT1/Po9tysVbOmVbMx+o1js1ntsL/dRquBOqYgBRyhLGc7S
iAozxOwnjzKM+XSyHNhj1TOoNdsrbox1SBf+3XVKjVIkx3sNjiy0Hjc3m4wF/Jg8+vCPUsnrG683
QjuENCO2gXnL9HPUEarj9yiPLVV3eFV//JbWjmjEZNpIDiqunPOlK+lHzaKIWCLo344dNiXWnIzo
vFsK/ly72rdp1CAKxYdjzH70RFeU1+LULyBu0Bn+icHNeUPjPkpF7TxfAAZpx63ZDx+i5kdkgXOb
hntDNkaOfCWxkAOmU+nCpRK/udeKvMUQvDut+20TROh/LxBnrA1zilbeDQ4jYxQc9g+CEDnBwO2m
eklb50EzllFLwYbPzkP7DN0lNsyDds/ej8XS3ByMY3tA507NgPaYrhmNvxr8p1lguHppJxTA2BEY
fIUYzrZYbEsfxF9qZYE6bDnGQOf66koTaDW+RcNwc7tWFmWyvWOwkesIUEzmzClg5PRrCysJ6058
w6gHs3nB8vheeb27C10VIdw4n9QZBukmXD6LclcPLJxWRFlTG2KcyugkDhNp3EKW7JoO0MxpcXKw
C0Id5tCGhbVe6ADZjTFxCXSIroqvIvtvCmS9HCLKodaa+RTjlzL7ENzDR7GUyjnQ8L0PEPfFnSkc
dbLTA11c0Ue31n9mYlT14oAgtxE2WdSxRxn78UnOVhSCjZ5AsmYfdSYMYmy3DwmyMO8eFjNX6MKv
qG1oFPFVSTkHFYOwRUkZXeczJ7GiPMAh5e1jheMWPHrKLtgYxvpLVkqcw0P1zEIruJCC3mxhj44w
ihFo/zdIADHynB9oPp+cQvHhHJ+JDbBdzKKNnEEbqtLOhq/I6qUxtWdjDp3MDLb3y5b4FZZIL+/h
ewRUJIKZ4CKaFFAQvhggOTGy7/4ZahVhvIKMF1CEiNJKSQ0QTRAM2XY6rWS6fzaXAcr45Yo8PUMn
J6L3BInrwjxEkv0+g36DM9r1+PFQNH65HmH0RbQ4WCjuNXwq7dDjnnK0eXBr0mqPtn/V/o8WKxf9
GVs5/Cy+dTgbZBTAc7StzsD0+YPMuaEKcE7N3GtTg5+weZZRi9NQ6OJMO0JSryfKlIGr4dHm1grf
xcpVOSAPlop4Y7+Um4B32CCpdIQ4WoBez/of2sU0ZczvVgQfgfy586acPB7MjMnSVfT2juCwdK5a
X6hKl4xi6Imp5kE1KqvDpFo9ySG6wvnypXO6wHWfJ/RqFAE6a4Q0/kllodo08lJI05QBQN9jgw0G
ILspuSFvyiPQi7DYbO95f6kyW42D56Q0j0zNi1FOAiscyMn2wYL7Fib0lolaZrhJDJzn7SH/gBzh
61datrD7J1b7vUt41fT9ScfIUYG4f2DaXuiCy97fisCeyY35y2ratAHoz91cap7JLHT9TQQkYxw+
BsRThNoDCO0KTf/IBOjXkDbj04iz8C2OZoG+8HJn0bm/IAYOKJVUFodA+8re+IJnZvr6YZpPL/n3
5z2iIPSJPiAHW3kkRoUfk4oVjRTRqoiwj9wE7Uo8Pln8Y4BNCJGUjWdNUXraSCnPl70wk/kLy+rC
ZSEpmAMcAHuHVCz9b9GrX9Na+rMRnF4QDAy4Vu+O2ZTuXgygO+DeLSqFo8zjcpQRveXeyVT13SvP
0rJ/vEL71A5Z6bqMNW1H/4WYP/Vm4uyH/xXCRoB/y3w1uP3aPxppP9GyfympNZntUs+KS2uDtwnr
IS/Qx/zZuOnFK4koNiHlUU/LmbH/5cs/yXpuvS3BIKO6qby6JhUO/Vf3hu+CVYGubaC14gBjz1oD
mib9u7af7DRsSF6sRt0H0V0AbxAQEDzuRGkvuGqSponnaae3f6WBqpFhXisVgMt3NQv1at2PqQWR
gc7enPBeSDdfEzrwx3MoGhKQIrdDf06o/ebNO9FIzkaUETPQ1dloFQmm5pmVoC9Li118OS8GE2p/
G9Jq6qa7M3DpMVtrOAXJQsZJvLAtAg16Gvp2VhHfRKWz5iZl3DK6lQUnnvrh6hQ5UgCHMEsmw/Ba
NHih1Ix97mZWypxLGaF0IvpGEtKjRwOSZNcMcsHtwOuXuXNpYC3CWHWANXs54W57aHvzg0J00QLc
hMU6B6eH1c4jIWMxB3FC5rYkTNf/Lpq8x8z00XaRzxBBqPFAl/9FNofcZ2IlgzuWAeujCwalbnwy
6GjL6e8gZL1Q4O1yFXBRj6/6vhMZ/AJLpph4v0gs7gOC7RA9N64X/sLEDM411jnNXsTXznQXeytX
tCAlZIvSRhZyJab6CPYIWkDMtrCHC4IKph5oxmG9Qp87UH+dtu2PM8xYxmsrkCRGdIkDrJf2H70m
UmlmcBrTH9aHnZj3Sg+3zlBanPOH/1EQwyYsGN2HROTCkOyFJ/6dSD8DQ/r9E9LRCnrTvVRo+CL4
vkR68nBrJyTVodI7bICMZ3l6YfektAVGO+xMEKDvIfRroDKeJ3C8GISUoc4LvAltwH2fM2id7g5y
+j58cSD3goxYO2jD8+DlYCOocTCwyy8CuiBmxOYHU6jT0UCg0gySa6YsavYHDyiqFCnbuQG/moTz
HpJ4/qMfOhXPeDRQ4thPdUcUFjvwUp3LPEXsORiBj6bc0cDZoRDCmb6yKahE7iftCZIXh7ipgaBi
2jqJG7zhtBIHVPhtJAvFJmJVz7U7qaU6m+qCHmfn8Zp8IlLBIYioajZcsuS9vkkWInVu1P8KBqIJ
oLutOHnvchanq8nW00A6VfkvsoUkAp1Flar7hMIZrd4k8ToHVSq3DHFSFKD01cejlSrOMKt+PT7G
D+UTFna1bGbhHWXWj7TIqgYMxu6pC31MfpM7uB+K8S98VZRun1Pvulwl+fNxfh+ZeMKbXHbENV5a
CgaHBJF3T2rTh2UYiYcdYUAtQCcSiCK6AoEjg7bZN6clW9b51uEJdsrD6GsNis66beGkg+3ughwI
a0wE578wbzeuF50kLJn/4LWeQcHM/Kob4JO3DvnWViGsWtuL3bcI0BPLgcTTbKBDTDo9Njln4Azs
qWst9xshtD0KO3KKAZOyhebaAz/1sBVrGvpWJanOk9dlHMNKvItMD+h0Qjuon40h3tPyUj+ZHMGe
N8q9XOju+aa9HwbowRykx9/bVeutgCTtnf0tswvGI+VEteTldB1orZPaSX5qfldPtPFNPy5RKnj7
9xoYVLKaGQpt0mJCozE5ovli+a91kWHQYfEVAZSmZJvfrCd5GSAxACWoqtkWYbJa6BF26j6BH03B
k3selYiFHNYA96zLXQsN208PRTqfA1SWLcdn182kNLHwxonjad971kAF7Yx1g6SpaGnCi6EjgPW7
iZ4T/cq+ue5jJ8hke2N9MjIFn0iwBQ95Ou6MJa2ITYcq2oUyT7Vx0AfgBQEEMF31DCwy2P/tczxn
eSfr0loheOkPRbf5EqDsjQNkbUyorssy8u+8W3mTXG1dOw7dTVSVJyNNeEwlfyVULI6Vy8v+7jp/
XXlPh8u1Zc9ObdyHCqf7HyB9e7hE+M0eOo2hQriOrrH5EiJVUtGn80Wkz/K7R4eAYZxnzBvNUBkU
Ac7rm71YZdVm3nedpA4pBVgyKQKuxyhZu0agkvHOFnAKxes1d2Ptzzn7TUrPKvHiGoJrjSb6gV8w
odtG3p1ZRrdARcYaxRHPdSjoYI5+odaqtIm0wier/vILdpqUSbW9DsUXTTo6QaCuAvvqR62aoCI6
GUq964B1pbPXMvCMwtRJDxmsCUz36NB5rcS7xpO0onqxWBLxH5zIMlCa4uFoGuX0gSW2PZgeW9kX
aE2eKJ3bmA4bNJCzUoddX/PTESYy5U1s0XSNvmPdjrSeYXbPU0def4r6r6qTyVQa71NNiFgIhoH7
HjpyPU+uz4skwwCStJwtGy2EY/1a+wzn5C0BeO0GBs3sv4bO5dSFHz3BD7gTJkWWRx0mDlf5pONi
I8b0LTOWZlkgfQBfk78rBoPwhvLnJ1xU2AK4oW2iuf8V8dewnYkEWFRrxagFoFzWgYSlhDVDKGzM
W0v5Kn+ASelfpRq4c4oJOVjH2piR6JBBWczvN4UwWxOs+OU6jpIPY/CMdyiYmlgP0xW381UnGv4v
eQM+TCs+miHffLfrdYHZuX+2U+3XAoLSFOOleVuMpuhYzJCEYD0stFg1b38P4Xz5eYJKHiZnhuyB
eqLypbGUcASiKb9OTp1T7NijkocJM6HCR3PsIX/Cfjhbth5IO20HgRHrcVx62sCkuZTRuyQ8jaTx
5gO/uQE3Xd9lyed0vztYZbQ2PJp4qyxLaUyN1I9BE53U8UEHXKDNJkKtxMVbRbEgVqifPyGQV/f6
Xf9B4hk/582X9NC8fzpvXLHSYI7+MJMXQRzfvLnk0+T9fryAq0EFdCu+D+zf70oeqjqpwKjAYsPS
WCajds9jyRo/sYpfTz1cRBQnLK7RM8Tv7Fuhqt7JnRBVikzr78RkxvPY7vYA3g9mfm0Gvsv3vNyi
Dta420suWUCcp5T6ahejPZ/rGxAlscPLR5gl0y8t0ix/vPeDyXOji5KkNlieEeOJYdk8hKGWTBoy
kkoL4fwgFDLOVDGCYcWbe+5lAUnA9qEZ30D6s1+MsoRMjx95G328pihq60riqNtE7wdUd9pZwpnn
P4jaSPlbQ4f+JrY8hcZEx7fgROCLFVwTYrU6V1Acp2ED04vVyS/NLQ0Hmps+IBbshwT2F9geZCLy
kNNlkUJcGhE72ghbHlRb6B3RSW0kSANuO/H/hh+LppT1E88ao4s9qJ5o4387aTHt1SgfO2G8ZmBg
0ncpiVQUK/D86wxI1GWwFy4KBmaKCv7BMiv6hZxp8Ola+LrQcIp/NPwdrV7Gxxz/uNV1wPspVWLI
WPK1m42Yj2p9oaWD8u1gBdmajmMCbZbed7igwDnKnd7vI+Rvl/abRMmWkQ1t/y10Rz2Mf3cH2JDS
1U9k8zDpqv2820iXcj+/F+SQQVcjYVR5J7YaxHkIn+NT1CrjVxO8Bfs//uDwujrQh6GZJ3WjZgw/
rv+YnwMWFOUuiKlGhmQwBdQ6y3J+h34VoT8foea5WJXzz0m6bVm2EpYeQ8jIKBI96cmBfwzSyqce
kJeCREZS6ZDf+nZpqclHrkEe62G0Z1lk8a74K1asGKKCVRWf+2FKQxB+3aa50lLoIEwUkaSzJIcY
dzPEDLpehBVjmpy9uqeensRr7BIIfxF9VlV3IDVJ2LhL2N9InfRcTE1U9qxFAOZUmTBYI0q+6I9Q
WK/8RFyFFsp+WfY9U/Pfkz/YsiMF+b5tphQlu38/UeT8szyPuW4GXAQDFUU88WGBqA/7quGJIhY9
AChwBhsATsZIxIdhZLlt4C3fmWWM+bbW73mEKrzXjnYDis4piUDGv3nEXcQbt8YItPa6JpJ+GrZ7
yTu8ZHhQ+KjhvhSa8mygPiYWcJVg+pu9pJVXARpMLde1c8PQeISGgBgTv1cQ8Du7OrKR27WJO1B4
AFTIDHPPybJNYPtEOKluYH3WYY23EY2RpBaNAudpwfjQB8Ic7pes8k/FRy7LrhB+/ClRGOJML3Ea
pXcYMvTQrYxb5uWwF5uzmqtwkVp5DjRyIaiE0qwq5fw0PHxAOCAu71K/kdshyPs4S83Hb5dEKKGc
8xUCn2gt2L61nQkSz9R1XrE6nC9P9YGO1+llRKmFrYQd37UJ2+LFQi7WnxGxXuCSajhjspBXhIhM
L5Nvq66Ri6bauez0HmA/e9aMOAn4YnCl9DUlS9JfMK+i0gSW89r+7Yh2YqY8+0oBs4dFkMPwXL/g
H29XTDr1aVzt2AiwlOcIV3blsdB1Q42xtaccW1lwpDRNF5eyPlm4L1dfVDWTDr4IWJczufVqNZcV
HANkEI2LvsyNGNqVp9L+wJxU6xIG7aLXlNX5yzEFis9eo4rTWVGA20cN8xKU1+EUkBHy0K4y4XZl
lKZ/OaEz9pBplIVeB//978KjgISye8u+TtVgQqje478HSRPjI1HVi+h/fgJdTYf3lNCZutbRgCKN
KqDpcvv3OB57ILwkUW+gjf8dyTLVUA18AqL7X8jWzydJG88MmYaL9r6JZrnwjvzw5yEFGT9fLwN6
kLTHr/LFz3T4f68fi6gkwYw4vammcIh/4Yam04ZkCnZIAcTQyqQyeM3cxSP3qPxJ0xgNVPZM+wWR
C2+p9JjTTNXaWUcdN0eBZE0k6iVNpJJ55snJIpDxXbdCKXq7NoEjOkkl93qivWeQfithzoh1hbYg
J0nDFVXMoXXf2hJQcRlentVn4LuH0X54sG35QJZi4rDNht1awqs/zctxrz/BRrTczHSss1pbuyAs
/prjZNuZlKOZu7ej4zi1gOsiltjD/kkRz5WBCorv+U6WcTXfnVpHLNNc0q64Za7uOMJzR1pKuE/L
NYVMcGA+Rx7b1FLoFReRKmEFM5StuLdTKE8v0o9F0tFV4xd9ht2NJOOTKOimLkqnZ1qieLcuz7mF
ohkvt6rRpfGLvrgZLsLGazxDyuHhfU/Rj4N7dCSFkNr6PtyKk7M4m5Wx8h1Vtg6gFFp3VRO0VCme
ic6UxhAtnYtL7Fh4o9WPOBQ0lTSQioLZ68mtPNZ4N5fuzH1etgkgY/lAmdJApFUeNFPA9DUDusiO
ZlAG8EFD1Pj5CKnAScXFM2uBXzmTrn6XKOsglhZOkfkhNMkqH1kbFP4pY5OS72BbjJ09pxDTzFqe
B+NurQtSx3xl1yuW6mFLpxP7t3UXFurHrhlJHt2fXIFOCWZDk559i5rGloSRw7eNBlK2TvPdYXGW
J7I8WlbQW63lU1deEW3DAbOED2P00pgqGNSutaxfGl2vpjE7oGp4tM5QMDA7TPNIn3Qm4MT9PAD3
bULbiWU+bEMHFdgPIbIahkjB4g/GIhEjhOCbcskNe3sqUR24hh8w6HKIQMBNY2cx4sTEHiRVce3d
704nWx9SboaNJM81jna373iC8IeUOZ6yMobWYXq14ocQXZxWMH5XSC77v3e/a9WxnFkIW1DJI1JJ
W/7bUbimRZ/sIHzdh7oSUnQE/pbXHZilbUmrjiBPngjX3o2qjcHY9aCIYQ1KGZtx5+wPBjyoxJHq
0Bp7at6iWQ8qsW/QMVQT9H2bkSatV/zqFyp9WbNgdBLSrdCRiYB9hph4ND8fWOCaFvWfvLckAAwx
BjBsQhGCKmHVraVlmU34rVmJZvrX8GPEw5CeWCuRnuGrXNz0mQAX3v6264OceqapqPJ8fqmwWC0+
PijeUxtCxjQ69L7d316+7pe5P4eJJ1/u55mIdt0xKcqvM0418Mlj5GWHpfc8pixH8fAdPkEytGNS
F5GKb+WFihqVS2r61Wsk1tdDufpDX0eOvc3QAGKo/BQ8diKM6Z5vBN6u1gylI14Jh2DMXHUyFtHH
UrUgstSvD9RBmo+vTdqs0CB6V9rxjWs2rh9fUSxapsNh6x9fraklql5cxxHv8EXwa9f76qld5OD5
jATmfKW0hH0msc/GAHucHgq1T2kYDSv7V8ho+GccOB/0jVDmMOG2EAKolHWCu9ZH5Hq5e9GPlfgj
QeJ37IxkXwhIs5xNw4F+MwQUSCx9r5Gd9DRZ2qwxUa59w11/z6H0KMVXyWck3Bfzsp1R6RjOS2yF
Lnt1N1PmxO+v6wQDQXCHvIiyMlPFrYjCWg64uiD/PiO5zBDH2106/WM+dvDAUTLHF1PMQIxvm617
NL16Im3pAiEWjuf7X55AVBs/O9mFz3HLN/UrTqwbl3t3MUK2b2VuPYUCBizj1tJIPhrx7dI+5+CC
aHZBPRwNqJLe2vkeNWWWxWwEl55MJrSg7N4YSdmxka4SGMD3NG5FAThm2yaZ9pYK1y7L9Oag+k09
e1fwyUA54PQiXbjLgWDkaiFIlU1SHgof3mZFjdMwTXGlrJAHsNwWhUvmSGs6SIfF/HWqk+V3RyBj
FjNMsOR0fWqZoiQS88HGl+339SxNhtlrnv9m2FDEZd5hkph2++2shbjpEC4aDGqsPSESkkaSdRqT
1RlaMl2dMwtyeQuYbGtvEtWWYMSExZbVlt0FatbnY1hlXfxW36WzB8ijJ7r4Mdea6wpDW4H4mJC6
jGULOQI47CBR5N2to+xLv36mhT99xHRLtZvMk/cTDGlicECVS2xuH6MLJ0LyZgf6ezFUjQlsO/HN
g/aQFQYENRbt6/3UIYRPaRY5qCJRDbHi/vvWc+ndVY7jc09lA8FdB5Sb3yCHqy8M7II6lAJeVHet
8HRy4ac7j7pE+g4Wxt2SCH9CBzVV/iGBOo8BpPdCLNm7HxN9Annt7qSf2b+fc5XC/h/m6XQTK4UI
7t4TKTl/12PjoaQUWYLWL2N664LzHhdpEAtrXOYHsslHGhCOFYFebGh4OTkaj+PCB1rrPOBm7WnF
vgVDmGbHWjvrAWf1mz08SsrDcptnzelEW6fKF/44X4vtu8wv2ydnARpvBngGCPifxchw+JmfRblQ
QaVmMPiQ8Hjo/NIlfEDFHFhKJ7zmLa/Enq00b7zN0/HXrR7LO91vCh5yvdU9TTkBujqKVoD2PKHZ
eaAzWhpS0CMMfwGO8PfWPEF2Y05NGPO0L1BGEOco07tX2XDBHzpe6qAHERPfEa2g1V4TqOnG/I6t
TPSrMa0HYWCIeV9DVwThFkZVyWld0KkQV/jI4A1QUXvjUGVJ6q2B91gY0+n4o1B20OAyKUuvO8BN
KMLlkfHOJ/TsXe8ATEt/7UWBii6GDeaZIf028VFim1ZIsL2bzajPrCdB5u2xBfQ7QUZ7e835ZtBi
zDjN67zYSmLfRTyThdsW2W4T0Fz74Lon2L/7/p8tGQZUYrLJZ7cLmrDdcM4MdZZ53XOvLTjiUpF6
9QkcIJFWIIbZqSqd+8088WExmxNSXuMHTX2+pCOt+xRBChyITlt/ZEZowHtY9rVBQ2vZnl5h1TWa
nKr9rSLaULH9ofd/xvoIXEHOriZfqjIQ8iAza/sH5VseDtY6lmzxO0hQ3Km4wA4m/KGw7f2ioOln
c8x5xzeYlDXyvAKq+p8JIAUxT1ASTk9TRlu8SUbIQbQ2Q5Ba+9CsC/cDcUDbcCTAPArUM47LQ9/Y
KaYj4litqkrg2mhOMTRwwNN8sWcWAb7KZVyhHxmYgaXsXV8ukI8dbID7A0xbefbWd56ju4+0Gaqv
QkSqQMO9TQs3PiH22Wy0CZu4JM1UvtaOIambmb640Lp7Z7f4bq3Qx0n9s1u07qNj37g+nUvg2pIR
c+lzXKN0anuraiHakNilX11o27uFgfdNE9SD0Zz1yYf3T2B4GX1hT2pPZ+oLakF1CVSuQ6HleOh+
8AhPxxsGyu28gEyLled6xKV4wZeM01lGlMjRWxh8qUtmMVM86lM6C+oXsKFsdGQeLTTneBJHzylN
dfFDQeBE76oDHABM0d/nDmr2z0voC5M9R3g1GH63bEQCDDerS8G+nAFNrclaBrx0p/MOWWJl6ddq
f+GeJvo6Fi+Rtub5MoH5jtMU5Rs7faC5U4yFDrNcG4gMPobabI9Qif7fK9VwKwFPp72+t1mfFOYR
ErYP2fOgIVzGaSYRPyxEifLnpDQiwvHx7V3F6mo210RyXL7knhmLNn7xhyEyVxp9twqNyPvHoY/+
e5ASGbblikHYRaxzTHdfx0JuWZjVC9cCSQbDY0+mtADhiRdXHym+hZyPPS8KSAPtfK2LDq7yeAJ1
a/GedfHpewCAitMl3hxBmJMV7Jyh7o4ndWG6Es0CDdiwTsurg/T/JRlSOUiM+AesVfmIed2DpLNf
yhk9FCxADicpnpXo9OVE+6YQ3z+xjn+iB/PAS+jcHwKIlp1oewSBdqtvUz6//3VZa2CoblGl/H7J
kBwOwEgvABxvTbWpZ9yXxYfSAJV7RYF/iEqW43eHsnO4a0WcNo9FZPxTvAlmzc1LTqHT+yPElf+d
ViJ12SwZ/w2t+TAfvEJY2Bd4ugipq8H2PXU7RYm4tDHE3EBoqbEzeCZBVDqYAzImDeZ93h77g62c
/bhNwKHNp+a2IOia8jkkasX0DT9Fs3A+N0IBkkZ9GCd/MZHk+DI56ZkW4XyvoRlaCwHlrU1WjN5E
R10YZrsHf4zjSkZOwHdUoIXcMhGtRTDjEfYRBBIx32UoNIduJZ9LkIhX6kpVpi/OiaPCO6siG1+7
DYRg+NhxUvYHr35bvC0AcKD9/ZO3h2eP/c99E8JCdFuMemT7UwNq1r6ZYQBeZ+yNk25DColLq/qp
Hmp6i/nqZWiEkv2cCKKhho/pLBvOESVbW/UbOzOoVh6yKmbji2fyrkR7/Uj75ajiUzsSp5Gb+2el
BsH7AxYqLngQyren9Kh/XVngLck1qH960iGpmSn+nHNB0qvbqJYpTN8BLuq4Ss4pLvbb+EfIdT5p
51Ooubm7o9Qc1Glvvm4QZrzxR+3GU6BPB5ROLJ3kR6Tpo7LFYqfayDN5QVB+EUScuxY1Gc68RT/y
XGlBRpdZa8DqpzEIxoo2Rsj/LqA+wG1bsnj5uSCbMlO6UhHKeaxzRqgUW1EtEGevFgLeFCrmngjo
pwUtO99RjHaN1UxMkPV05E1lmZ7PzjApbrZTw7mbW3gi9ThXpReFBHbMBVfdKSRT42MruScnaK2+
YhjdfbzO2XjYJDySpb7/1/skVkztqk+BFm49zrjlgoXYh+I/ohoq86oOFCJ3wsg/3saFlhyuTrc7
aCuCzW58EjUHuy/OxKaWn7UQKz2aqWcO5aqxZ98neQFoOjOHITzHqBluOEAy4YLgNv1/gxZ7pOdn
1uQel0NlnZz3xV/SSzXrNYqRBUbX3b6zFpO2rbBbhMeBIYp9v5EcT7Fwtyw8n7svfmRry+yE10WC
1K83mK4KRTQXWyeOoAme/8Sk2iUJtjDhRZCn7jpRD8tL0B43lYm3A3xz8d8Eydwo8VQc7XIArb5b
gWidNt57ht3YCIPanZynhf4Qj1qQKVEwIRggWpz+iTH1VRftEh6rwMD4vOOMHuI900h3Y/SMDFgI
weYWXPXjVnVyal7Rsv4k83pia9qAYU7+XccsJ7jBo/8Ta6iyK+iKSOApmhtUf60CvgiXQCUzG8Vu
V8yiu8yLJiKUMHaRCVMfquAMUUeCvj2T5MV9vmkzhQyP9HPfGRA37pmcqfqNaT3ihXV1ZHTswD2A
h+1p4Scvg5vHR6ec81G2By99XKsvu7Rtkl73oJzBk8XihaICSWQLjYUNAxTEbkXfCh3Dxqv23lXX
W1ZP39oejsclxcaY3t+8bTzUMloIrj3nHXulOxnbNdU8m8gBWVR2FPwtInDln7dykRicXQ6hTv2Q
jYb1qoZGiQcYcA6kcyPGxXZQ21D/zrSSdUyUhK1WT1iuRsAiRf61EVJXMd3BhLdh7N7S8WmZX09M
jMJ4TNSyGRMBI+oM+7muDFylXS5VeK9TzL4w+CsJgJeRakTC7HZfHmhVWnQTidTAywmA01wnEa5b
suZIKLSWB6FGrelDvjXmPCSasuo1/NIiILWfFESSV4cXXBY7PIGwzv3bTkWWi2l+BS0x5WVDJdMS
RdpjtGBMZ0664Gcl8/gq7CgrU6FeKowRh0MgQliRUAQFfb+pXyrT2KqTGl2t1M0tdYuJoTvIuaSx
T3lVoawTyrxgc9P9MDVBNdf9bbQdg75uEFaq2KBrGMMtqt2o3cfx5DJi/HAIKeiZA3G3wkRPucQb
HJ3gYEsPlyMEbcjyTk+bwW28CgsCgb1y2tZwdQfms+z0ckSolR3fh9PlIt33oRex5vgRXF8haASL
1jyncKYIKVI0X0LyBrWaovqRd8hNZBWMg+UgrqP8jNaI70jqL+0zNDZsb0oZw35ehenD2IpmOABu
HYO5c5BbE/jJk7kgJIj7rEe8Sy7crkSTyRyvtyLmpICxjrxXWWQiIJJJLPsUCCxvuxfZ7a19Av3L
4hTEaphwjiR0zfrOGbguCeWcO0NTX5+tsiFhVl+U84U73L9B5qlM3a0WCyLy/g98H8Fd3OhNeu/t
Vywzw1mhqhN7gImUxGLGokqlysNTD5CkxZX0mrqWdGbecRTqWBDz80dS7+Y9cZETP8JIaxR7VOzn
smPUxZfb2RviNTKXPVJQAYbjk7jBS8JQPl2pjVON4Pe3/MotIApvVrISTVfCWn2p7R4slitEcq1B
OHReSiWFehWMF+1MqvL42zhCTiVeJnLdz0GKENZnnXM+CfTEO+D83WnULD2htcAcFl+WPVr7GgKR
KdaxKevAlb/izvp+GuKTqCDU76dZrvgPOMlL7ny74kryKgGf4tEVNaiIOPKr0vYkH3hLQdds4tM+
Q1/lFrduNVw37g35GdTUy7FAVJY0N75OR4XLj6zQu1lnvfvsNUHpdi3N0rL7n4tlNjg8RS7P/Tx0
OWWBRSFOIkQMxOZeM+6b4JKitSKVKSNGPdMKuHsmQmbaJOjadXcC1INtWmruTomzCBcNicvKUB2r
S6xtZtHnePSlr4+rdOkKfC6fSWCZ2XMu4Nfdd4xIl7ayxkdBhLBDOYddd/J+I9ZjwrUSKWC6Prjb
WWqoJTgWTLQouEJz7GB2SyK8kiDWXKDKptbQ6i62Jtjk4SYeay67wlz/xnfRC1gmFI9mfHIwEW1V
kxJ2vBCw47DjHMwBA//L1yOst8w3BELVSlrhZFvHai0avp2eqSi8d3Psv4346+bIwSuRRBnR3pEh
V0gVQlQFXYAUctYTqOGuBeRMacsW/3gb/VCnJ14Y/GKDixEEteQc6tgBpvBX4n3zF9nyScDfLMpZ
7SKFzAQYmFTgP2kAmc086PAdkTCPMkhfIFDWlWLJ/hj6Y8sj1Qc2rU1QClqtgz79f+CGONBCAbQ3
WuebzSN49wZx6ORWMWFJzdiwZEeJCThwWZj5cHT5Y7JICSFBx/FcpgZ0d7e8GNmhSf7g4i0Zi8c1
umacrEHt/XRhScgPazQ8l8yAU9p24efKDLJOD4hxdO4wfwG6DJM25MMTJmfCzdUR7ndICLw9c75+
oBFWGTtkD+YVke8AzCzzS++ZNA44VAqYEvZ18sv9OypEH/DgOwjGdvopGkWCzx2LPfLgQJpvmdIW
JN1/CGIywc3wAyn5zw7FARCkN30iQCuiF1hh+SjV0JatPGCYJW8gDlFrnkYDwet4i5i4KUhfhn5+
AAEAXn8zg9myxtAHPraw2+t8HfIPmeHExqp42iqu1/EWdlteZ7MGX3xEvWmGpqvEY/jO4iopx4WP
Plw0KXt+3W117Y0K1K245e1RBp4hIKrUgP45WtFX4jG49shv0OUlkmO6qgGZLqspUkShVL6SQlOB
2rwqCxOCjrbSRAbYjikwU3IaI9M3oWcPw/x6b7hNVOMnEGrSBgjdqXS6DHre22vMKrb18nijaPJ/
UJMCc+0/m2elQoEYsYvswwLqrRbhySaq+mu2EvQxgCYf7NlIn/6g4ZwJVwICfW0IK64+gXc9JedG
nj7815Y2yjoPywGHgbnS+eMB2PD2LlvhrlPQ8jyrdnAYP53G4f/U1WFLYEQrlbCcPQwpu+/gJpRO
AfB91qOygV/1u3ggUubFWJw2kl3jhwhmNlLC7Dh3dvtURVeqY/W+rJyfpqdEPzaZ+jN9o+6tbaVx
4KBHr2P/wI1MW0LP2fvWY+okX6RuKgitLWLRP7p92ea0Ybeo/GoRLYUjGgcUu4t2bmYzE1y4g37B
KpsrtDPXYPMMOFxByrGKLBCcMSVEI95i+FGry9lnZYV4gr3zXxInTedKWB8pAJswVqaDY4XTkpkt
Ss2w5K1lz+J1DYHMqbGFBIJzpW76MHDSg/wwO+qdDu8pKvjEvakmdjWW62LUoCUfiX7cnltZlXFj
6tCjAfPZS3glNCh9NwGeRstlxWLSKtERuZsWz6trYJvExKe7sw8SrPm0xCYt4EUTXt8GG1vunJlI
2bv3qozgWTjOcqJz6G8XXsZm1p1hGeQBA/hzd9iFZ491xmp/Kb2+6mSlhXSy+zxZouOjQ8OOEhyB
8rmGaMNwtihf/oORKorcsxjpGEHcotDhPJxZ5SLWqERJI3LFNRtJkm/8wfRSgEGauUu33xo1Vdsl
AWI2eIWuLoPMkk1i3U4rXh8EKhUTyCMrMHQ7VDWl1q06g7E+0Qv46GhGZoHWykUIhOo0ygjWQc/t
ds8fpQlYyFafKP937SJaOcatlB87V00jR9tbE3S1IW3/KEixXRGMHZ5DpmErVQh2Mvdw3vWN5aj4
0MxsyiDZ+DjYRRM0EAjK8wVtOMU7XbhyU5S4QfOM7qZmem+hK+zkmtWJQofqeY9rbj+c7qoUC8AM
l4PIrqEn/giz5F0gR4av2x9tCBXBSjG6p5q83/WyDriWCxzJtJSqQIiPM/D1EssdOjsbjMB4pSM1
s9xB0Q/d1aRGmeapi5j8SyAn9m9PH6UcIqvrbdCggMTcZd/WPptjqHtC1GPAxXZr3MCfzcBPMiq0
1EHvL9QbOq/S4OU40PpVGyVeYCDk2ZHS6YJ5v9QJeVL2B53UMGtz8uqfHmdQEG4PoLf8v0OMx+zZ
7vsXmJbvJyWHxMKbmycKzZDwyYI3ZQQQ6jUe5MOOFOpZJH9J6oSOfGpX0RQkwJy6O1vE9gWcY6da
qgp6BqvtLfqC19T8iS8QcsikhvAaGKjwK0VM9G0/8qSYWnLD6OwEb8a5ginIdzXZ2q+A03PD/WVD
bLH5+pp6aJbMTj+PwVtl6U1nJh3LQzMxp01F02IngSv7wojtPu/mjTMjucWEoXVv9C1Ken4pJp3F
E3xf1YuL9xOyDNVbhsZZVi0ZnQzAZY+BWsPinB7aj2FzNS61cIO0T/8cmSaNb/m2iMf+2zOeUlrr
afraJIIAbaZurQNC6yhbkImHorzsepf0QQe5WGf+YkSDmyuXfRHO2EtR1TaWimQ3oC/yGLMejFn1
cR9yaVVjmqQENQgV1rITga/oE2DtuNwd0LKWEAYPe4W9uifZv7dvRimcLI4r+lP7IDJ2LuUnu977
RHiY6SdW9KFKkSzea5meTOw1Xg9KY20UIaYsRkX3C2ctSJwdl9B2u5KzHNEvSu5BdRBXGSvnmjXE
w0g1su2YoH0hZSdoBPxEbADDDwbp1r0LqGdrpQQGAFkrb72tJ3CWzcHj5FmMzDqJBqkQiZ9Fkm8S
ymmZqEDKL1FFFa8oBqvHQrcLV4RMni67UjqeQmzExnlfzme4cuMRKCxJGrHpDA0UDO5+MGH45U82
kNmYHArtz+zRilSjCXUhPoGGlT9554CdP7EVdAWyB138HvP5eqvdLqoDfJEWvqpuapUbmN9Vc9rT
30hnw/B+4CaA/F8tZyUUv+nACGLGvYzEjjslXFt8dPv1IrP8duoJfoMck1SeKhKkzASKj6FfGWUf
WfCEFTeBhrn0j9xEoBGwjfXwlf0ubANh8X8QCkOBpoecwleQ07t+CZL8XYoV6ffnqYnOmWwq1hjY
cwdGCmg9OUs3Z3Z6nwcxjeECjwxX4jxN3a4sfGVnUwUqdW1EtT4ZiG4opXHWsnozzaA+sCjDX/pb
467kW7I1vRRxAKagjVeBDu6xEHOT6DISxFq8p8SfYMmtl0Dzj5HOBkr7okL1xteHKuZ17TFs8tXm
Wom1pJ/FrviuS5LwBeylcnPScPJJyrY+AduXrVT0oE1kwpGsj0Of3UHdjazLfjeHbhFl1RdrYwxg
NyN+37CJRsu30fJxIRL/oz4aj2L4yDerryNwMzUXIS5R/oOiIag4kZspc8g6q8F+MHJSTkZQqcJ7
HVkoDvGyL+v39luBOoWPCRSlaOiMigtK/5egzVtwY78h80w79bC8zC999QXbbqhbuVYwY61x5CXl
67iUDu9pmxyFw2TdY02LASwRb714PoxOhU9yfFli1BZmHdlJJCjQFaJ3o6uMEcrQaJ/n0LgK8LUB
uI+TCyORRNz390VrxZf3L5KNsSOstV+KMy7IFvPS/O49X/TxhzhRPEt91JXIU+Fgvd7/CuKKB33S
PdGSwyG143IczOajik8YVKmJIJnpnh70mhJ55oHUPyYnCe5oSUasC9+ZOigDIe7e5kG1WXgEyO7L
mHy6M/+8uIqyCq9o67jOd6r4b3Zt4bgK0DUYVcu5N12CELKyAhojwB9QmiLYMJo3cS2BjvdO2q1N
OcnnEcU03EVPNRNWavJVzw8jtV3yJp8sGMEJ+gYTtP9nXJH6us0JXCQSJGOdjnVybt2iD+9AlSOf
XXLpK6nElGYraUq3/xONPFTB0fnJ1gjmWXK8pHUB7t8ce2kYXLEJf7mTnPyJz//vfjQHCqHJEnLq
itC3vx9O+e6DWzzO2TfKRyrwekFHtD/STAsnjeKZQkTzFgCnUWK+9klu/I9SLelg+ybNlrxSxSap
RfqOMSNa5tyM7HdcxijOKJ94Hf76O178uO2OHByPsbB47LsUX97sbwz6WuIcRSdMZFI/38OZ5LNv
L6gOyHjL1RSePQltrdPYIVBgSz5tiVlb4szgyJKwBsMNZFKPbNXxlTFWC26FedBU2FU3o1G3cG88
3NL38i5v7GrnUuDmX90ApZh5qJC5W7gycv2ttuZLr9RaDr7rHndcS/le63W2Y34nVOGOZ4OSOAw/
gK2UvyQmOXmb5YfwqpGsUsr/PvLCR5iTmEuuGuJ2nMZO62CM3KJpSDxpLnSpMeeQqXQVr8eSayFd
2l/Xch3EywNa4vtJz56QRWXlXlMzT60zQHuCcglMflul7KkU7hmcCexYHwCPd2tU3Z3eyCIY5WrL
0IwKhA/kqVfnLZY1UH9yY2OlaMj4KRY4S+H8+WBk2GC1pn/mjsmICskHPwNo9tCE2KVLx/yxGhvb
wMUvpyD5w/eVwggCkn+FIHoQHMg4OHER0WSyvcvCkxRfF0lKohTmZ2QdwgFlyIGmVTQHjooTvwfa
+aKN9aM3rVphzBpIjVum1c+OdXHugYRKlcDv35YzF3MCzF0gedSpgJRYlQJKNJWOEPG/NWgw112o
2Pbz6+iAu/0a1gWjHEIxT3mT71uYH9hUNOh8gV8lf58XrvLCuROpMHwJPm599gkqUt1+sjULvwqD
osQL6yZk0iCNKXVPUHzdCNvKJAbFCBYBRsdvieKOpIpEVJ5N2HpzjJaQ3aUuCU/u4I/PIwrPMbmS
YcLsbW5l+Ojs6sf/MX0ymaTq1m/j/8/oGKXz0G3DlChnR1pSWn4b5a9zDS1G3H6zmjzO3SvY6c0G
hBSokA9Fqn/bnT6KE+Xz+gO8bMG8U1MYcrfy2rre58EkP8SKsaOostoGc4pu+fxACfNwS+Q2XX1w
i0A4D83oVSZ77/Vy+MLchmFffi3qc2CvViXpjYYHanmPPcfjJ/zyaXz7c6PzQryS916r6wwjez6i
lH58NutDobnR8ammTaEbMjSYGYmKtG1f1NEfiuKKleCgFyyH2ex10wNG+oBV9dV8RjTytmnkfYVk
YftoUJ48V8g9dcEaixccPKKEkacq+nHFryoDyTHadLnu0gVGguZO4I15NSHxTuT3EmY2CaHjpABR
SlZzfS7/RNkG8ARv0MopGq6flmWE9DyhbJDFZT0821rHt9+kGch9G0W1YKEKs+GpGp+rPPx4rdYO
65uJBa6iAGMWX369YES4xewj0ovCX6ewiQEjRgvjyMn1Lg6HY8DZJ8SID8jJMSj5remx59VOvCPT
8XScDguFlvjXqMcvYhqTQCFV5njk4Xs2FDP7DCfo7GICjdyaNmFscL0LyN4GYPJ5PmEHgtfrYUKU
BGg54RTRw9zHiVXfaDEU1w/VLZ/ZRrUMRZMWAxWq9oa9W426BEc6OwE5R/qZKBOihIBjfl5o3fQo
n9/J0cUZdJzm6AvTFd6l6d7GvGlBDBxV0z/WY7QdGgscDLeo8MJ2gmE6J2d73jcY1Wj/9rvHITOk
6TgV7YycJxlfx9RzGJNuFUEUmQSwutYGoy5Qp70SIt4qOvZsbGmzyA4F5cN8vNCeeJEprWoVzTvI
HARz81bqztorpRFdHEO1GECjC2fRvhqgNIpDonNIEPb+ImjXCSzZmrwkqmaeChMhc5xO137ZXE97
FLjMFGlzvrJKpILSmP/IRP6WfQT83z8Y2jEjmk3Q7x3S5xl7cYIh4wnmUFicHZPCSz03bU1/e5gA
bRnktGTbGfO65bTIL2QUZO8top+kIcENo5j8tEvLjWfKLtW5HBYjJ07osuV5AcwehFH15GgYJdKs
ElCFnMs62xfA5DnJnj7i8J2tFdq7mQhm4oplLhkOb4AcA9Yt0WRZZeMkVbsEijk1NX8UQUsUhu2K
XAb7IhEjuenIFc7CFtkJRA3O50lIBAeMDHcFFK7RGqmRxRbB5XZJfkv3Iwz8tWhoYxE6Kr0m2671
OKmMJTzdArdniquIykFswwuSxXbLDhpmPgFf9PrzODFvHF+14R37IrPtKR7EG8RpQsEtc8D24CxZ
5PsdhQajcvYBx9+YDfy/s4DuXqj2RFYTo3q69dZ8ZQqheOsRXBEIe7XlQ4roCIwHqMPHY2r2aZYQ
BlpdDOtUKcidyeqp5H2ANki/uTuFX06Mwwu4zMghmnqZpVk8FvESfFRtcn46c+ZJ27ZInJ5sBWph
kleaP1kL6rObP4G5vS9E4rEoHnmRUkMCPfkNx6a5qGDu5Q9McaA+D0AWbVTVTGY+HV50+ULitTom
tAz0OrDoyE0/eHRYYtDsZ21RG35rGa9q7pY8qARVD7PKZaZmCM39FnIGek1TyDvlasC3aFLX/l8t
lj1uFbrPny3Wcszxm4xO9mjM3eGS3Bnj28rPoAt99c1kgpuwnLrCdi+43rK+wbBluXDRpUGGspIC
MP3Wcjm83gNMM223YorI0sXbt1hfS8R3tk65EipYBiz7Xat4Y94G/bMGGQ5pTDNwKAMaYd4phe21
YcAisbzEFiKz8W7Pz8XtnM5p6EvKRm42ypADxEElfvagzUaXrAif9eU3wYoheH0ZPFJhPNPTGOkX
4G/5X0C8THC+nlQOj2xENIyuRqaeinETN2wNAVxWZThvXEzkUEjy9xNLccn1PAyaxlNYrjSoS0Kf
uCF4sP+SvEK1AOTyepkvO6VfAdPM0wOE0nAHTouUx1/EA8kGarzDceY+rPQPqO+sBo7Le7YzOjPM
r29fXwPSoHGd+2UPOaS14g9waIGcLDmES/1PpK9g1iQu6xO1I7xfat13Ak1gxt7yEN7tRJzVls3/
ZHhNYQay0RKbyhKku+I4xqXvRLPWwLZ1v4KDFOfTg7MF0ELX3mAeKD/orFf6qWofjwCOl8kkT8Lu
ucbofKieTUiDPuJnlAcCRmwWqHlAQ8tg+Z+T1C810v9OGR2v/3Ay65Aep8eop9/2qSz9+B7zaMFW
MBipPNzi3MQ4USRpG9KaXoWy+a2sUDzVX00d3unUetuQoR5FsyYTDfIG/7zkbjjp63thqKavVAcN
O1yA6iXqUWWAJqM55sADx2otd5PTwTWGcyQ6BjCtNJ4/ou8QHKy5KU0v+3WBzLtrUpwRbUHt2iq0
Yu/AdKqKLkfdRORaZrfvgMdnWPtMFKOP3XCNLmJ9K4ZfAYZJO493MnX6h1PNVHdQ1JlqUtJ0oxFD
ftHUzA/ZgrKm1WqLStL1JLKDOpofq8RLf2DYg4Y9LzyAlYGCD8qbh2HdbkZ1762KgKaVRCfd9Wow
x9N3+Ry7R39z7bYERsfXi3XXirhnI9MA42djsqn68O0jQAgcdd4eLiH9pjEKb7aXGnb+NFTkY6gT
PngqX/n09mXZzQ05YgiD306T43kWKtEA/miE7p1d3MrDIo7G7mZ1SzQTzcZxUNy4ikBza/9zEwjW
bWZLbSQGk5r2EvjiGAmKefi5GjUaJ3oYUQ1f0XeOZHi4jmuETJS2RC+f3Z/meiX4zQnjW4JLWy72
FRSD4T5CHs8CgFeLQqQ3FzZuSoFFVQKNzQl4/PZWiStpaPi8C2kjddn32jhmmNpbDRrUgVe4VeGs
t9N8NR9T/mnzcTaQQLspY0V53/pHbpWIBz2/cv0zfffT7rI8I9cETocnWp5hAR7Njj6FiVaYAu3D
kb1fHGYsWjnlTgSIv2sWEOngzluX3wEtMjweWGlJM4pQWU0zfwjJ+Wr7mcKPkkL+gmhmWJYzcCmJ
tLOv8EQ1/TUzz+qzI5EL0ipSO5VZigkXFp0nVPt5cPjd7Ajq5DGhRIjT+Lf+f+LTGCoINfZ0pG5u
dmm5Ptp0b3zzHTi/QLykF4+hY3xX6NMIPQyZbujpWQBGyEzeete55QfYDWYhsiufrGOGNepn0Foo
R9gpFFXZZGPwhK+XpEPB69ZV1WXeGorq13clH0jRxt+YdAv0/0Di4BAMUz5QSNER8gfG69KFhypp
/9I4cNylwgGAqirMjQKdyZKPtRiPN8hlSuwx7VRRyeWOBx9S1Pp9eBToygxfcIsCMe+en6BNPjx6
eGtgRn2Tx3Af/83iDHMnFEzyFsD0B4Xvfo5JqRTspztgr6Wb2TflTtdrDMNhoZev0MjlHr7BRgHj
MsJ45PG9sWZyZS7T2TyNPSApRSuPe5NnTuO3giTn3qXkuNM3UR319LMSNI+clcZDVMFyQnm7HCkh
UlVdMt8kZb0b6ZdYFjovwD2QuqyJlJc+BHbYO06ufHpuu1iKBocLCLnviaqyJXFWuCGkL4vKLFfe
nf+IUiVfELjlPGPAw5UtBFLwcy1L5ytDinGYiIXpHN6nd3qMhF5gCoc410sRHZWJ8ApH5nef42N3
hwMY8fn7TLDrO7c0jhfVCOMOoRQefxje5jztOXAnyQNlIYBkXozW387eRtgzHpfYwx9MbfctOuMA
k1U2VyIPppLXH5qJUeOqm2hGh5wIRvG16JpWiW/m7vbqBy5nZKIoO3M7mUbRA3S8qlqz5knPcRh5
Cfz3O32fPFz78qMwZMoWOM8Dibtmaiik5niVYkEgITrkZQ48+g/AB3KDrMt7UltaxGrAYlfvrxTh
oZncI9GX1UU+Pcv7POLDedeO2PdTpiLnb2kBkOlxcNSGQJX9BWpE8jyMYX99BVhDbzSBGrfW9SpB
9OYpAXeoSXnkKDdxBNmJOCYQAiymgP1nP+YmB76IYZ+8tUbbVn2/+R3BKFY67Vnmz+Xdlxbj1csD
dp7vJwoGrjuKBnMCIp4+P/nYzF/5QGdfzj+GpOSKT43t+vQ7Gpj/Mh9snj7gFZXZzzg+0weIQ2yH
l/uaeaEeHgO4UX3phcyYZnmLzX9nkL2M+3RIAGYwV9RhwgIJPoLuOBLvzXrnCmSudPlr9iV9aXPd
5/jj197Qqz0fdpRZom+DTaM2SgKEyKj2mtmpvmJKrFLnZVHExyCbQPD8h6bTsSz+hOqAAlUaUVX0
tbm/JscWxONaMdSIig0EyxuHeRHu0qQWs3jmcS5qDeAZEoawePGxo4SQEjpOe1VlXV8m/xiw8q9D
DUdAVnsEV1zq2zpRVopiYKWKD75C6ubU2q38ZGv3WNhbDxLLqXBBnPbgGMvD07XtmRnYMjrnAWsZ
3JnqPwYOlIchu5JSRTUpN/1q4xOykusIoXVbQd5SzZ2w6tNVYTM3d3ly7t7OmH2Q0Rt/iU0WT+ax
fQ1RRgveBcmMUWfVX3sJJFo5KM0CMnc0viVyZx4EO1CovP0GmZFIi++ZcbEPbQ0eLRBj6TUxlcAe
V8SK4TZTIdfMk3mNI04fp8o5eytBqnsL7D5XxVCj13dpEbPB0n3VSS7AAaKrmw13hU4a89K4BqlK
uy4r3Secn3mtZOrCkSXN7MMlPYVua/F1g0lLJCEVLAX9yE9O49XMEebNChFs1iNnihtCgiB+3l9s
u2HJRTWZOZ7vv9tbZxprqMwjUbrnfsBJYkIG5u8nVLFmWbupSfYj0+V5bYiaE90cDdt3CSUPP0M3
sQUv4njggb5hIhcXFcLA35W8kArzAxHgvKpKPRmuVZIT4MspY5NwTDFNSOjf0azVF9UwIuPBh70+
lO5c4WfApOyQniBelgpVKHFD5uDBOME/LAkOgm5h2p2zsRL+cN3wkTNnluW1728tob/DoIpw2Bhm
EInAVoDEuYy/oktksOYoAAdoIOBNT2kF9OiRjIBGShsWkslw9LzXqYWsBqG5dWZreQ/UnGUlbC5n
mzl3uDNycsjoOZn/U6cN3lUHEijC1ZuC+qbtzgLGNPkrCcOL+86gZvopAaGf6ZcNzGBuWRikGp9l
NO6HUWNh0DEhgaJ9223TjBP01y+S2cKm1RFnBVlrCZLYPtKtoSNxj3/D4t/6Hy2AojQnfK/7uC3k
kQbVhcEeuq1nnBl3L0eDqyjxtkR8fJHHvN9Li1HlL4vE+Pntg69Jm+JVyRGjwLkWewOHXnut4QdC
mhTU/q16rTqlAauEMoxNdCpZwozqUDi9dnWG+QzCtFIvxwafDxlvpQprcYdPZMUeGwAbrfk5nDmc
nEFMKamPZgQaRFQ57eH/dIK0euUNBCHPVgHFKXWNpmw4chlE8zvTyfT1C5O1vjdV9byBXBnT3eRn
Esuz77vxakHDXKyuTcZwXpOJlPyk0+0v/gYkArT3h7uvCbnqgkcRiWQCziTmk6c6z+fMDdEpmtoW
q4JvhNQeSpWHYaPqHPH/SYsFFzXui+FN3UNWDwrinTcQgx3q8D8H+GN63SWR1WFTcZRFYzn5GDCc
mYuHytmZt0RpU+MvilcK2UfaxuOCN28VKCKLYXOrcBJrSDhgUWeimWCgN40n3hgq4u5UzwKjodWl
Wn4AFKBnm0WIrqrI6KlaXy0SLHnnCaoEf5hke+y0hKe7vKVxTb2wkqIfOFEJmXUdoV1lOKLHXIaC
mMpXMK3ydIEXruoNZvCmmwZ2Ca3YyxKm46jVM7Jd0tp/psTuM798vbwSzbroHz7lWSRJpUVBQvZB
6+9Gn5HEZIVRFsjnZIzohyuczyVtjf/5uLsYk6yt7vRWnDFA6LXvwA/M8hPG6Qh2iVuWIBB3J8a2
3U8UUMl4v7dtK+a0ZKJUC7ZZTwB7/90r4508o4aAimQIjaxdkIPeHYVu8r3JueZhfHxyFWKtmS+X
zegcEo2+VJhGVWfod2Erjypy/i3hdPHu52GJ4Z4Qy6QQZ99Wzn4uz+L3vZT/j0/xRcyr8TM6zU5Z
Ys4bxnKPJIpx2XMIx84b4PU5i2SieaWbqFFlAT7klqOZdKtHdi8W38WPXEFIbN9hg/IzMu8Hvnq1
V9+HlC2+8E8e1kSxrfXUMRSFKfoK8jxlzRTL40/iusV35ObuiFk0hDnZPKaByvcXpXq7mf7hatBT
j9HzRDAKTvqIJFToU08nERW6cH3tFKUHZlXm4E4HO80V+nENSkf9gZDDdsDKga5ax4WaUEcK03Xk
GZ3J0Q6k5kNnz4ZqDjaBtPFiRmMEbp4zqNj7wxBxeqyDtW831OTMLfqkFeU0W7oXJ4/FQKyB1Yfj
gyUYpHMnymYMySKCvG+6blswgLj9TgNRajS5liCa4cGk9CFMIQPuC6yRWBqzl1TUI7wuxsxIxayB
lJ88D91/t6LXtH48FFCmekdn2JovCJRWjmzzKZYfGdR1oh6AhBdF+X58PYw4dBvTOdW78sGeX0SJ
EEP5YqNBamoF5lwx36D1cjXMSVrfzGhdhgXdfja7UaHSKbGeoYezAni+HLeJ1qScM2gLNB6fbBFa
MV/pSxzaCh2gTSl+TLYhv+p4byRBK8qFMuwKVkd05yoHog1AgANu0qX0ZIvaJomADtG0qeKfe1Sd
HzowLfnNbFJ7YoX9wLFJqr0GYv2QMDEbrBXBjyfdl4SA6VBOZmFIKSyU4oyJjoVtIUA2b62uAmNP
prHKII8Bf+EhS8xHzDSkOAaIL9IgKf8mUqZDaIvTGi3iYeLKnhw4wbe9d2G6+kvOMSrWz6ijbzT1
7WRIECdigUSNYztUv4acOVjPQXYBsWBqoEZlNViYHPdvg6b3JFm4EBYWZkKFsQG/jA9dSQ5m29uK
zRsYFoHWP0+kUodWAQpHcKbbaVwl2c54ALb+pcMd3nv02hMOJQKTb5Cl9flODUHGEiPC38QtShNK
1V8BJaCgMpV2lwhn8lTO1sCRQz6Cea31sDX2xreSMB+ysZXeqMqt2mwi2AK+kogAtWsaIVrhM1l6
sUXR9PVL+CU6+9zUBOq/er0DqJf0bYXVSGeiN+R83vgdUal4FYr6xYczXS2a3hlvO3Xbr7ZVInxN
IIc5JP0uXYFDNxgO17ULMeXXrtXarJskDHCuQDvOEoGgbCr1Q5xcVwydo8qE+6bOEbpLvVlrl2t9
KmpSp2I1sBlY0qV4NPN1DX0fh7l0Q8JJqKwFCPvkluTAm1SV9f1yY3OmMW2uIMEj6ZvFDN7D9atO
1d//+D2YTOTNfh81tAvLn/gQCaTnDuQteoV1/SsNovTUsR9OIGEDGZJA+dBPLVeI8AKtGsqDOuxs
ZbEbrrswjPWS6/7c14mdD2CzUrXljjTNUObtTAZZBIg5wtFy1E6KKSNqlqqLAgKe6dpw01ch1NRj
daTQ2SJCXlJT6FBmTyt+Jj6AITLCC+N8pqvjsjQCRnB7F60yjhugGvi6FHqc9Pq+PVMSlYG1KUf9
pr06NuravOg6274AhP49IXPYRxp8RFTfvrkp2zbjtq66ng6I2CTI+/GGXzzTABpAFP+BJ3Mao5T6
nIpc1SXmxJ8ii51VmLnDZ7jEFQoXVWSAp0LfoEc0LgGpTi7ugSSuwxmTWWAPuDFn6ec+gOZcLNb3
sNTUHDCwSVNi5obfUefG+M+wY3QzcdbT+wXOFulAqs8yb+Ybi4/HcAVcrNI9bP9wZEWXIfuZd6Ij
sY4N/+d00wEK2fS1D3zEngYsxmlnUsKov4GpchSpzlk6domYJNcCsrbQlhc34t8uUO4cJctHkXcF
nKgX0RgUG+zb8srMtCT3FOeqiuum2EBZ74Vdq4ucbtNJXSbhKtmk2g20/pmEhwPPFZ1874mgCfrl
n6+R902tsy6kVuJX1utK9gG3NBTsg8BBTwkam7YmZrX8XdNT6w4bDB0tOH8gUeR7jDNsdttJzoYI
4StQvfRJwj6qhdsMzwTQAeiYt6p7a5VV7lqeYZouYmawiYXgX8T8nNRoLil4oRNEcBfXVNND+YeP
5amItb2dQwsT/dWZAWe807NVNSRtJnsml8Wc3RB2Xz5LunpOr83v04y6WfLGFrdT9a1g2xcv9vw5
PXJ871wmzNOJSwZWQqyovwbBcLI8xr4x/GDSCNzquSpqfbNUDDac48vzj7zbqjlyhbgHnifkEzP2
V6ARXSucEQibbuJls+r6N4UMOXAphvDs4OLI6kV7h8FgKtWdEHYCwm8TiFIblgtCsZyUS4rPxe5q
zsNQnb+/9RTTpVA6varTTAvJA7CnvWduvA60/vBcdU76+iM6mFGO33+lq2RpyBOE2Qr9ebya6JYz
zmTkxo2YDZlCjN1L3hO1oxZD2aS+abuY9X7ITOApsBxMk7DS1ul+dVEzP/XRca/yk4qttE0pqTG7
AQgo1C9Luuu4bfOHMgY0F2MnXzNe66mB3v+orlDpFIBG6YWIwyl1319uJ0MLrM5+MTSFJjRw3sDu
xPV9q9YsDX1tN0SOJ8TMoqtYo6+nFlfF/xyRHYNxrwKRL1gjQKFnHYf9UtPUEq9YEhlKKF8OAVz+
QDEF7XDx+XoYpZhtyxzEjJJQz2n538hh8/rDL6JDLsMU7pmy7kwEE4HcUxFHdBYpENTHz5Y3J+Vh
/CYcOSKhT5YqJ+OwAgWVIdtMkROuasFaSKdDw08ZDKF3wlvgJifytVkIAniZ9xHAYARupSNGL5Fa
5z0yDly6+KRTb2KlHtH0/58m4jTFT7134y6pqvzXarOimP5BYFD4y1mCpIb1G78xYjF59OA6/NtE
Ah0RpVmnSbs2qowE66cJNv9XQRFps6I5vZJgh+HNHIeKE+zYIMElzWFun+XcdxlM9vUduYAAnTXL
ZyLjBnXhw+bO0P0tVNCV6sN4l63LVp4U+WGRGSjtCslDcw/9lf0wsg9KPItz+7T4OqL9TqFjvPWj
GlcoXSvbFwiV07spd4SUTgFaWDDvPqagTYcnrlVWHDlbaL3E+gSPOo0tTL9Tl+rLEi7kEBMqUP9g
7Z3PlHgaN2yRd0lkMipFXZDLOMrH440S/7JWSqxv4gf3eeZflOJR8kkTEUz5wc98b8YazahdJICL
L8lXwhdOmFPT7gqNj06wFYoQQMQurKHmausZRyAUdOcZHKbeFphxrKr/Mj5Bt/AWHSSTJXLqWv66
qM6KHA0URSEAZOGBUBKDXzFwBoYEQJ8deftrJLo8GEY1c5b57m+l33XL0FFuJKi1+W2vbbn8qwjD
K6Q8cswStgUmpjLHqXnD7k3jqWO7P6GEATBrrLyTKBFIZbY/cW4dDd+iWZ8SXwIChYiKZ0dnGdl8
4QK2KrcuogYc0yDEtCMdE6rnIu9GAOj7KzSvqVQjEgNpJaYeynkzEkFjPQ5dC/m6YZzsdNpZ6rjG
YjbQXn6FlOISUOl9vkTkZyFoBKM9k7gtaiBMNvMP9XhpvsIPPWNpjVfVerJWg2/MJaodvobuFQAv
uPYrTN1lJnyWPIzEX1UU+ZjGdfKcDtJtD0AwaJYvs9tTbVyZCH3CMd6k4uNQDyBMQm2o5JDQVN14
P4rUuSUA0MwoNSzUFWaJZa18Rag0RX2bqSjAiGv/Qwr7Oq2EnEkxTMufCxT8FEEzN6MLT2k5CqNe
33tXGu8JjMoa4r3BI3foRya1jeruHbiEJkTtCmHjyielWLc0GwcOsLaB9v/8rjIVsYxtBZ/8lgg6
QG6EuwCVVvp77qQuFPZY2K1CfmsuFE14V1I3H6x0uhZpFuq1aDMiGBOz8BMHHUXPxFbHPrsHDTs1
tOIc1qxXCzow6TawqzAv5Mwz0zDwg1AW8TIvZ0vjKoSMsrLIZ/jPoa5bvFGkNUmccFnmAego+olh
Cv2vCCI3zAL/95JThNbmuLIlNIOMcJpdQ5i1vSFOvVY1d5HQbiSmh5rG//PcM4EhJh1+Ox/7UmXv
ZhpsnoeYzEa4WxO1lVSzcaSZZNfQ9mHV0Tbnuw3H7zKI2ysdS8FLu6eTLP/td4a7xIc+uyzRFvr1
Bho3Sbr2/w1ARFWKOgDdtdZ82xcMrigHtVk+IOY9xyJjhSZI1nBzJrHvZqGxgPIl3/NTV2U17i+L
QDro7dCz7gBr6Og5kL8R5xHPFTDH9UGPAkqZGci5l5C8p5r4nx+Yj/G05oD0sTMm1XUSQdiI3GiZ
w8leupYu20trnXwy/H7Sa/nIIqCMTyJOKwY3I4EA0M0/DoBjT/f+ceHbnDqiHSTu4ta1Ol6LFecC
nNc2PFCME3/5yPnkCZF0NkrOtTOQ9hIuL5cdJt53mj2TQMIXhV3MOvQy2i8LkoSpvUwWm58OKoY0
IvPClb6SVeb1HT0kbwciqpVk9iY57+0yYBmnXisdoCbpOjxPUpFI5a/301d09YXnDcbSkfzWeewP
QlBXEm8rGIRXh3RVzVHUwK8w5tDZRg71ymOMsTE9Qn2Ps1pQqFblfpqhW9KUK02XzLlFhwwMqfwk
yObXdhQ9iduP4MNR90GymIkI0Fnve1U8Szmqmp4PbxNGXWUXks4ffJOOnVb3VUdgICSSoeIK5EHJ
Gj8KYhJtkGZZA7gxedjC1dyeW/fS12Jo2zQln1tcKd6XdjpmFzwVfW7QwAVKdsKklpmpfMzaoHO+
QJVFfpm+mFH11bq7Ol+hQYnzzhHo8rYNRAw2yn+VnId1lmKlEhnfBmupGTp96kQJCvSdf82urkII
lAQV5i5tOh8Kk2ah4I4+MMs11Wygua0pXTlpK0Ef05JsMK3PCfky9OHUdY1yBtNgyfWaapmL8rf0
nAGrHidM4cIw2jbzmTkEoy9V7qpDzp1AhQ7La9qB/wUsCL1B1skfI+ozXErxgIr7qgbXVLHqT2ay
1YZqFVFuKHb7K0V2zuIdEAMrPsnctq0sTZ/7HaNXJNC9C9XdOfcB9M3j7MHU760ikiVT1+cJYwWJ
lJZOLU51YvbpJ+PqwnJ26zcTt7JSl/e54CXxOZTh4BgXOoz9PhbaXshFHfIJ2CiIZY3szd/79AKk
X+4FxrPEzw6w8Y4aS+38IeMflOyLGW8f+e6ZlVKgaZwWrvUg/vC2GmmXrdJMHOk/aYvYPguNe5E9
lVTpAWdfiSPQkC1lb+lmS+J7SODwtSg1/FvWpRKQu5PCtE8TIjW+iZlwX+/Be2wLbD3crFJgNcUc
UuyZk/2IB9lWZKDPtbzuI1m41N1gkr/0qvDIAU+Eaq7udKMCnfReaFloRMHOZNas0aDSeW38buhk
qOSmlbLjVvuYcD/wPx/M26rdD3OBPPuBVxlKi4YoWKc/phRfOcuazXWixze5vgp3wGBRGNGl6Wz4
1D7OHAUgn8XuE5WvoVG4Kk/BGZiV1jYEgSvr8mElScIMInNHtOQ2ZQ1Av78ToCgoZr9fhXU6mofa
1//EvCBTX39XzaeZ0BUk1C2ec5WIjo1RIG3CSFQkd07zR3lZZcvNrF175viRpJnHHXHQedXIXIm9
v0VOqb9WT6ZmqnXHHaYl9qDJbsq9HggNG66cnCM9PXcu7UEuq/UtzZupA0xG/LNk7U6j40Ttxu3P
HRr8IffD11Ms5tDjPX7Ofm9QZlngFjgTmgzXKSPZ+seECATvtk36L8P6BoZi0ooo5ZVfIucnQDuo
YINZtOckXfKLIltJa/DZTo2g6z8vkM/efXUIrj4sIkafbgwcYLh4IRoJGFXsvR7fEW7xDX+gIJY6
DqGwmi2+duSjmPFahhQ/kXaLwFeIiGbQLrK92LnynFc5hwt6f0CghE8Yh+9gnpQRPYa9nhrv24r2
eARok9NaZLO96hTuB22idrg2yfWlBiAfdS2HhvwL2DfrLCLqjlQ8w5X9rbcL54uqfrtpL1y449DZ
PdlybuJLZ6DhEGfBj93M7+d5TWWUoEXlHBP5y6lbbEdJm3Uda3O4mR56M9yqarazQD9aq7ljVwDD
nQNnazJ20Ywnd0AzRUVVmwlOT4yZTmNen6Q8JUBUy/KENYKs7akBiEA8xyRdR+BQvtlX5g0eM0AO
vI6GIQ2nGqhM5g6vWUcVpvxbjtlsl/VjrsT4v6xWIOseT8mtk/zvGMGhr5GkDVvGFeMuYZwcO0Ej
H6LewmqX8XdA1ZlkoNwgYwXqCGFbBdw7FZE0k9OminAfvBt6QgUrpNTXVrmBIWYMPKvcA3XWxh6e
p40GZjSYxAY4SY1cvGyuvIxxHFfO6dzvsQa9lJXsNNovMFL550SCabBzlLudZBNSbw1N8/iIuhtf
FjYUUj/SI3YsYfqUwmLSCMZbc1W04Y/OvxukMxVHgNYOdds+zlw9oAAXGCzoaOeNP6TyXgBoNRQL
HawbFOBIkqDuN1b8ge6Rr2BRptRLhZ7jZUgIwfp/qKbTV0zV2zLLPythQmlr4eSYJbV+OcIi4+ID
2kKC9/2NW7SYeXBbIx2h743H2rZqUb8bB9zSfSl4TGGHi0qWAFTszwhvcbjh5QZSRQfbhpEq3L0u
ve6taIPmxjXhrAxccilIhCWiEpKBU7CQHd5mZG6z3RSSgRR+tSjmLGoxpdksLMyErvhbkMJGn2N2
WYvhXoQj8aFE5X0DuVCUccpHAYRw9NhxOYgjRx3/m5Z2eofAvE74rf/gtZBEJSb+iNQ24BRaK2ua
WZ+kZI4rCzRaIiUgxHi85DbQPAGKSRLfI+djnpZkmiWVFla0dAMjuqBPoy20xSm/g3GaVdikIRVq
peYo9PLkCdXotV+JaZkG7XETRrKmWU/vmcZn30KfZsgluXkC7A7WYmA6PN6HStD58wIbcPQn+DTP
57TJx/UtDJJ8XwFNCHpo8fatK6NNpGPl7HRyIdzlVk2eHBpqEE7NrOhTZfwzSIISueiE45DE5otF
ZYQLbi6NFcEnM40FdwR6WiA3PaNECPlf+1rNje3p/ymwdIbTLAxgsn5r9w4CzsvepEG9yl0D3Cvb
5DmhYQgNM1qdsPxITX1mJ1BKDznP+LT0oiDyyUaQuIEIdOhaJ/zdIL2lOJ19JUdfeLUqaNVxafsB
NB3q0+tca4xSU/ER//lTWXiub3HK7T7yO3rmhFok/fmK7JCnd+p8oxA2jfzx5i2Z5uN7247S5i2e
qxt4CmQabUbgJDSexPeD7X85C9/4lfoC+cEVos2jjbUW6l915YmHcdXWquNCTWWrMj1J/LZRrKoy
iSuTLfRZZK/f+ErBm8WfBt9UdRaB3bHgIvj6bS076eDJRtm5Mmh6rr9A+0wOOjdJbY0gGRqppsH7
jE6+vCFHAHE/SXEJ4LAZbnKgiPaej/p3wmjTsNibId383iNPKzizaVtTZYWFdbjuMusoqhyr4idv
TYys98LdcokP6fL5vSN2pp6LA3B3sWv8347c5nmXIXZgt0SzzvckuBb+i5o3T49fY46XLFCGxMIV
++p4E0K3JVhwMVHnZdPPMdGaLtHR9SdzqGx0MBorZks+VYFl0a+OxCTjhH0bPvCwcTWO3k6D4oGr
UJrgku2tJ+3r6z2VFvoV4IMzcCHGxVIPaAznLlc6MFHf6rISop2m0N5Kd68uDXDupqEI6KmTHmvH
SFsD0oHgfKKyQ69fVFDYj2uJ3WBDknaAo/Q0J9Bc1Ja/xyNLrFtPDkhAqWQUZbl2tuViUWLbncl3
+qcFi3ybenbKLTiBNIs+WBfpHDJL1+vfv5POsysDJPChWm6l4VcjsCbCn5m4uMwDWtts+Iiw6COU
HrdLPP0LebMJcHUCd6winzsmlI/0eOMRjxWhUG7FDI7kPXQCqD5rU9i22BmtJLykKQBQiU5NPMPj
NDgW43ZRrbncJPYChYe05kwcZCS+edVA5KQT3QdTusHbLEN6tMEbucXJyfn9YKPF1MJrrqg20hFP
ET49/+cdAnxOs4NfnShZ4+HzwE32J8xXq15FRo16UM9w6ZXu4W9OJRoy7wnb+QRL/ybs7p0oshnu
W/baPPAfKMHRRZYBLijf/pvSSn/YJCorZzdpk64ZE31yVafmQm4DZiO1uFGDWQr/Nis+6cIajH75
+bGZ5xShnhOQwULTRJcPSYXwCpO/Hak5EAfGNJJw7cji6m2njAyp26c1s5IK0TucFufHYpZ7Qbzt
WXZkkGmOOG3ghE1Tcq8x061+AnWZvlmZEgVSC01KhV61D3W1l1zAvstW3BIbetNhmWf5NduXkSnH
p5da8p849ro1Ma4Vb3+LH9UJoxp7rqJ1VR8IIOKcWRqHtTwghgxa2cf/QzVKc3sCniQjQboKHwEo
dI8kvcYBLDaHHnbRrfI1dRmnM8/gSkKX7x+B3xEKXp52PHi7a5QRf237k/p6OUlCgh084u4TYyAi
05NFN2DhY8Kuf4YzQlztA7/PEnCxccy0YLBdMD7QcFY0710Zq+aiZBAhLp5JYg7bXBK+9P3i3u2R
2QTxJCZJb4z2ppPVUfGXiEHPQFJEf51kMju5lCgZj6AwVN36mbcFxIba3Djf8Uro8i3c7MD464bT
iFRs8mE3E0KPWXZfjecoIs8wrRoMNDlq015jAgjV+kbh+7j620drEYuShkabdpI7PsHE5p95hGBk
/lqH5GyUEE6SKp6sLwq8z5xADDEdGzHY3Pd/5bXDCzk8y+cefpUnUAtv9AdREBXxNkOArWx1eOhO
ezv2bstkY4oP5R51oVMmCbEkgfhBO+sdwYOt3kx56NsxiwYt9F9k/5ItqtQCKjhZUUOa5leqLAH+
mWU5Cj6Q7aFXL8JXbUzsykYIIyoALsL3RsXZsESV1ibcs2dyMOm09Xfn9d+CpH95qUuYWpzKg2zk
HThiDKTsptcW7LNNGDXIpn4xXlvjGxAxOeqewEVQOdcT2cTmqsvGXl2ty/3mtpUNVp3pspaHeZOE
vEokfekU2+6nLGP1TR2ehqBAOd4E0RACxdBArjbl4FDsbCPTs/cZL3zzt7k8p/uHBMoUelSnWdsR
W5t867uihh4kRir4U/QX4KPPgSdA4fw38AY29kdehLKMwJBmfbvJkXWq7VmNwV8MQvQNxlmIcJ9v
rsKCNes9+dkMOAs2kDEAbS8+U9bVQt9PGzUjPVkynRJ2AnqOgv231NGJ3PUsk1Wk098mY1AptLCs
6JoGsjlzIbD6DnxpX2fPJfse6j9asisS4VTTz/IRxIU7U51pGEnfNkDfTQbvt7/rIfAfhrVdwdLd
g+ZnixoC2eioeNbs2vQkD0nZlwg60j6cEBczkks3vSrl07yXG7ChlMnX+l0/SFspeblUht/dIv8C
O66lBl6aAZqnrUmbN/oNRu3VsGKra8b/d689VDDui1YVty5jBeGrDGNHBu/pDDvn/WT+BBGhts5s
1WPR9GPKuK3OyCwLyJ6QyBmcNfYONas4CCBkyt4wDzPXm9pYOM90RhtyKhZUEwsQoGwaqCENtYwy
ea3Hw1+t6gfBjQqvCJS8jdGMjaIzDgS1ECQvvWIPtWH4jDPOWq6xCGOWE2CStuBc+eBgRBtDRwLd
g9D32bKoZTSMFtXxpdrhJlm1baCKqlZcW2kWF3tLxsjP9CJk7Cm09kXIVdZ164I4Zs11kspL5Xzm
gLLvEChv4UEPKQoDkqbHoyxOXlKUqKC5FNo9BXUTL+wefjwueE7pjNi5hEaB0HYK0PuHhznV6EdG
3CtnRAD1htm6w7PazEwNSpw97bsRSzeXYR9/R8nLjFEJMGoN57O6Aq3VIHluixm4lQ8pXTcDWDV7
TWRsqIL20hhAOKdeSMcmmY1exD3d9mFoevQTDMTLVuwr1T2vmEPK2k8w426XxqImb8EztBNkj41I
YcAP51E44BRF78DaOjBWUg38VSLZTuJXHmbdi2XYbMWEyYfoyUKos2PsgNmTsMundKyazexfREv4
D5zPrB50iBCqGXxMq3/fYzbf8aOe/SBH/PawL+tGqNEZ+Jqrjy8KMfm790FUEjTbmdcJHLvAzLw4
y7KLSUPCw/u7Zp9LD97mwZdyUq7nd6YFkVn77ZA++tbVmCxy5uhi9HQMStCFspdJvbEIp64tOZmB
BfLA3sEo/DK21pPdcbOrFqBkFDK3Bklrh7q0C4P19asXGjexOa8KG/HGbXFTQ8pBbVcY3rGL6987
MtKR8fpfWG478u8VzTM2sRhIYM5TAPnxghV6+vYAy6NJ97UqhCeojEzhL6nwZMZJ+TOi8Y/99dto
ND8h27kQRMnIPF1Bz4cH6AZJRQBkCpISIOIWCvil3BIJ7xDfemWBQsdRLFEblN5EBC/IV92ycF7v
7sVFvOk7YGwaPSBZhErfbqrwQiVh218NyRfJo+/G/iTpVhHE3eBtwAjcSWAVrcAcFRm9+Z17cMMR
Qgr3DFH9e/8ODwN51Hw4WczGtHO4UUj0Xh1I+7jZSP583hBWw4+WViczyaexzKEErwP20IapjZnk
dj66D89YUOebIhvciWoSeZ9sp6ywGqbcuDGz2xpZ3ubB8E5RqW59VpIyDSyhxzbWK+abg8jy5rnj
f5AnMbcDLTf0Ivi6A0a83BqojSe4ApVLiabWGAhDaovCOVCMZL4vTm41T7ArVu8pFrnyZ/9wsDqN
Thy7RJTBFy2lPfRmHShWPJI0HOOfR/j8e5t93+wVQJRCrHyxzhr37jw9lPjk+Y6qTosI7C7QHYC2
ViklRmnD0/WfAicsFOY6YMggx25EspamyzJBLjTguDcEJe9BYNGVXO3SwkY4aHMV+FJ7DKFSW+I1
ihWi9aKXY3M0l3JZ2rJ+R77QyerlPYQG4lABNQ7HEHpVynU/HHH2C+QgFgoz91CfgTkmxHlh0KbF
UqfF37K8Ev0ep5I6TbEBuRqXt55I4aRWnJf8ET6vV1PMKcVG0bqbPtkiwy8RxD/ZvzeYLgWwrqaK
vYEcAsjhKrjCHsj8bCAQ18GCIoPNEYxnGICjh/xMQFgIKkOf31iNKjBd82xiVzUVJaDCyBlkQ3mi
f32/+jAOgTb/qQLyJrGTedr/W/3wiAdE8EOV98GCMqYBbsl5QDKG0uxceBote33jC9QypyKvKj8L
wf7zeFQHne2iT+JmVdI7/xA0AAwJNLt4B6/6coqXcpoXFoANXhR9OgSjD5LkxvpyJygChRN/OmU+
0BhEx7KN1mD1aMAgu+t2G/iyElqxT6SsvDZljmRMXjOQ/ZJQUe8DMfeXkHqURZCtJFaQXk+wWJMQ
saQncMZVb5bFM6awQKuIBX+RAZ1cgFz4K96GbrOIHOKlLPaO9PCIViIo5H1+Y+uJnGa3U187eeCT
ePZ7TSvxaVg9V0+lOP1JNvNqFjq2jyZQNMDC9MPx+d9x83dqKct4ATpvEvIhYkbzpzDFPp+20mRP
IftehKQdDjnv5dARTB+lwYG9YY3F5+55sY9lFrAZefJwTtZ7O/hW5LBzKsY9Bo71068TgxRn5Fx4
s5d6k7snObXZg3/pgvyBWUUYmu9ARUKucww9EG86n4diJ00JrESg/JvhVqoa0Mv/d4re9RmEESCp
JfmVIHuqJ4eunje3YPVw77hnp7DpRa4szFXZnJc4FPVOEbBD6rvIZ/s6+YxxS2bbtHjS7E9d4+xX
/qZgzKV+9jHpCJFIGAfdrZRQ8cmCrE3XznrtL8dtie44xhDaGAuN5B4F7HKyX0GrHHgI0YTow7ak
DIOPNK5AhwJG5SSZSyJj8fCxpH5V5XT6ynnUeU3ORq8qGGya1GY5liCX67qEZl1xrT4iRuAM/uSM
zBvD1uSVuGctTAW7e2I5L7X+Yt3MQmrobgInKglZugmK4x87ThF+yDNDfAiYhELTn99OMDW49HZS
QNHiml41zcfZ3NoeI2280NZAPPP4U182XJy1BtdUeicgTtfGbSInEz5yIGEIY32UZAtKeTLAsQNU
K2GQ+o8jW/HHKu9zLSLDn0NGqXNQ1bDSd/2i3lUlkjkdWV2cq0rmNig8egYwGutrptflb7kAu7QU
3awu2jd4JsNvLH/CJ1OyUyZCGxZCekOaTA0AIgqgnQH2hM0jslXBgY0Qbvweg5tz0k/KvJkIh91Z
YcmftfZbqhRdA1daB/UpdkCPPnlyD6EnQEH55mfGEETvK8sf/ovQADZ+ULahIiixH/T3jbYtDnpB
nZn+fb5H4KErtBt9hE3rJkYX7xseaBIMVXOOkMyLq5yITmnLmNvEqckcE/nvRgpEis+ewSJqUF5f
xV3i90y3wnOGHq2+gp5G+KehKPLb9T81aoftXjploLYLodAaprF09lrxb7ROLzpfpfXneFSnc1BU
GeIXcP+PSzj6m5BaPED/pVfO2oAHv+9L2pP+PhdDY2J982n8xrRivPCAsmtKfrTlf8oBW+Y/RpBG
d9kjRZKG6LvxGu0kQnT2CXCU1CpdPUwnrexbEt1UxDUZLVEHC3maONrtR3q9S661dzGNSZlLR6q3
Glnz7Rmdu05d/NHuNZaAV7+X9lB7VcEMUV0OrrXQccK95l1ZkNN+DcWnaLLcBKCrVBzvJgPgZUpe
FxUH3qXysfddCLBXsO/8rnNUWTHR1zWG9NPXcsuougjbFhrQ/GqwnXBvGLOdctoFzcuEbbKKTRCX
PBuEwD7Bh8gSB0oqHyDbqELiDSLxr0T+io5l79RB9jVzCwE2prK1SaLG7mz6ckUksACPhc1qdizP
z9fvfxALy2rx0Hok0lQN97rs6p/zQNUElB2smHINyR09SdxOROET/SEUq6E4uBZg8X6/gdoyk7ns
fhHhoqKs5oZtmM2riPr3LtVKkqS/ubI3PzJFEDaHo9mupswibZMHw3XUs6ugP5yY+vAA6R9aDdoK
5k2zX+7j/i+2PI26unOrZA5NraggFqx+bB9e8mCxe3HJjPqyDnFliJPXCWfzSaVl6QuUwGaXh2D+
FfDc/vSeFeaV0ejLQX8KynMKbudH8BbZNEjIQpvWbMpBMbrG3rkHPlIJtx//NgYdbPLuU4HG4jNS
ntp6JFxBbGpisO5gixfxcbNpij2MqVbfehEWYx+4F0J99r5eVekMR51R/uy+nQUYx+romay0R7n5
mHFsPz0NbiVaZXIP6YpEnDgbJtc4uKRaffXgO8q9GFGISg3asb+QRT5+VXqbRGajwwC810O1HVPa
bj4Ynzl3NtKdi5QDiA9eb4jabHf6f1lpDqep1D+r8YZnYr4AcPZwMbaAXiFyiPeY6JivcEIFUr4R
4rs2uOoK9FOuwGJ6SpUUP4rMeIzQx4ngNqLgwO8NrWmtIYD7QQSV43mvlsbqD7zSsMiGeWZq02Vq
Ud/otTvfZKG6+kO7OcESvkjMf4cLsuJhpySdHMubCoX0+ZgFDo1asqgZrWEiQ0sjy9FkXFNTGkt3
zcX/Vy2TdWVMrrokN7uZ24yQeyvQY8y52QTokccw9xwCVc2s0nN84YR7rbq1soQ+ll6GPbumSm/H
gPruCj2UOQtRT7ZXSYznanE3plQ7Rk7jyqgSgFPMuCJwSUgWZzUYRc7UdnitlTBe+JyJ683ni8JL
03iXbnMVmeA+Dj3UexDWchW6irvXmCSSEKpaZ529dbFLLUgJOXkuN9j39pfXs20CI3PuBuCoNVdV
gGrDRDvk5AxOuFAyPWOUIvXf5ummK9zDUepQfClnEEDbxQycVVdo1S0FupBD07pSqWDK2CpM2FhA
8J2A+MN8iI4zrTJtC0mBxJB1f5Ua4PgwuaDQmeP+k3V2fy5tvkGWTDOz7r91xHJkTQXWWraAfLbD
xb7dQKtisHqZDZdqEuP/fIgkf+mqMnZcaWrAt09Yp4c5+UKrR25JZ3Oo/OA/8JesMSrMSHt8pNzJ
ZOCzZCHS9qC/ELRlJHJg3PlJ2AGTIvCUKfmdA+DQlSxGvnds3ZmODD28St/2ToUiTW6jG95AB3CW
HSKrr4L7frbKs7kJZgHEYDO4ukc8ok0CFKhTif8UPi/qIC5wAQrp3S8wBTyywBT/TL2Ci9sCnVAW
uzZkaFlvGwmGqxVHqfCYTr5ETZgb3Zz0r12EpX7+7ia3OD4wnOwooIK1cAYH3IzgfiiCnUxdTOyG
d4LokiJvnSAKZZmgQeDPaQ6hw7Dg48vudsJCFuKFoRWqVbdw/D/FCPF0F6WLd3dCIWjXGVFcXT+G
fCNNq7DzJPkIUnYHQx3HOYsjVicnjk6XiYCWG5KnVnGqUi1VKTQkEGOG0hck2n71HDMvX3sUxag6
Ob7lhfjFLrVZUJ5LXdYC9b8sOEAdEVQD9D0MrsQu+4BFmZq5ITgakPxubgRfK5yABE4eNaswHKur
MJD/YT2+VKyvfvpRtvx86CRkpy4AO0JZxY10+SAfUWDJ0rQNo2veodOKg9ouEKN2HzsBkjjbmhgH
jrW1O09nJGbon1NeIHcQsuWAHeYAONZzl0ur1iSJkubgR/xTUSzrCf1V13Y8GYWeAulbFz4FM7YZ
FJxJ95Bx1kRx39ABo/TuSgxoaQ6ygkot+WH2aHl7a8kN7OPvtIkAJyKg3cdMFkUaGVEuysUpPxoM
F/3mrILgT2F//TOtkUYvMka8WbO2KecKahUIdEwDNusDN8CyTDdISVAZYjohi+T5O6xUN+JUIHYs
GguDpVi9W1kyYDieu/mLN5GbsRMoWn4P2Ywg7rAnD+yd04zSZDOqjC2LFt6L6YUI+r5AGH2uRRXK
e4KLjKeQXPAneqr1muBjQvluI9SDbnabMh2s2UMU5IPT92VvZZhiVfeUwH9ijJL7ELPIEW7hRrOV
o+dYNcjcbHTJPuJfwnCHosLPdqXbjzNGt63GxW8pAqS1x0ljs05S7dSrnp8S1/EuEZs7GJj8xFuG
sI5Gj+4LCc5t0CaqTvTzmKZQJkGTbGICJsatyFvwAIMmpjrBiS2N5TKIsD2t2exCg+3zapPfPbHS
vqYse0eOS73xg4Q775q4MC0Ym9r2TYvyKQ90uyQFs7jZjIlzpb9J2+nknzvdzK81eFHT6NX6JA2o
guk+IqyJdtaxJRmTBgRx12pizXo0vsJDog4BwwsgKNgUIR+sXxF05IxMDAkRZCv2uk6DDFCzY0Fb
JyYZ3qQfZb9T5wpECDInKkTuvdzp0v47l9Wow+HC9cbCM3QQG+dIK4B0CZ5JN2iTxmJUohJqXVSC
REJGARr3dcQyacWB9x6igwrVBBlI0iMJ9sgCny41Scv+T9OUW1CBpfaI6g8Nugw/Iwnf/xrP0vH5
0s/fKhtUlalj1bMlfEiuyD9x4LIav5eDoeZzDUZ8FB/M7aE24bCK2fXW8kGCd3QdB6s7r5q0gboY
PP5VjKi+hBv4mH8RD/EBMEYbgzO3hRTMwJdnRsOMzQYd5liMVvzxGfPF8Cd6M+/MevBcuhQgrLv0
oV0pDrBmWmvV25bp8mHip3e+eonrqJQ0FhL7hVGJWAjGF8nkpuIii9tqiVUkfvqY3808RsATOtl5
9ev61/f56lXiAFFlgJH866TypsAIq8yyw+1Lue4UOYvunRs9XpG8mrqmkYSBV+t7hf3arUO2xzK9
R1cavD00rPVyhBReuuU3E1rxWCHlA9DfFQoALKN3imgDWwP5Vf1X/Sl8SR6w6iFdP0xDJMUuUpj5
ow2fAjT1H0N2U9MGVWWZE+B7xtBwNe3XK/gjRyKURsOeZTyxFBjwoTvcIInzS1dxh3ddx69/T6o4
W4Qsv0V0vX4dKN1wuEy/eBBspSkfi12DwiDLSmeIDdn7femPJGQxeb3c0Be6lrignvqKYdW/xljj
/0dCC8odFOBDiVWMx1oQeslv/kET57oleDgdr/mKVIAkSatix1tSVIdj87t4OFBDxSgqA8c4TpGB
qiy8RE6AY38spl+bonCHUqxYNZ5D0bjMS4uu5maFnwQ+5LWW5F8bjF3StHdk7CO2efM64IHF+Bdb
NNkWCnTGcrR+mrW/ZpDD/y/768lWk0rU0fN9/+OrwB1tkxOX6u4x8lohEKfP0ascQBT1wIaTiohq
BpEtbu1AyIL53Xnmwfzv9P9fCvC8g9mMZ76C8tEE4wJ4bCzxW1wrBZ8H+WUzbqnoq7xGyLHMqdfF
093B9spfInKhc/I1SbCixvn+pbWavS5K3V2voSpq9voJwi6HRFn42ylk//K6QjY/6jV/C+R+hzCj
V+3Q7D5CUNwVjbXfgf6wljuWMm8QAlj0V1LZawaxC9KThWMph8q7KmcQVL2/c6+taCh7hBaFOtIC
Z2y4PLKNJaORjoOWQCVaFplj9A/RRz7JS3ZpSkVaMqhPOANtG4WQErhkt/IrJYMgCSEMCQ2cnTnX
7euf9LF2ZQW5DQcy1vMS6k/An56dloHwKpqsNiWh5TuejuAm9WD3yFNHbHCD1bOvWHm+5BtrD+Qh
0Eja9mWeXjVjxlixq6NlOFZdxPIAo+fmmAi5fO4Qs9AgmioZN6U8NCt3OS1+0EyGhSNKNNp5sAD1
L7Cc+OGbFXsuTbctdRVoXd0ghqjO7h9RgOCLZohSiI/L5S+TxRUb5WXTm4jYl8LDcDz+AZmOTDqR
y449ipwStOfvuRUAvipam3SfHRZEkc0U1loIyWEPKV+DzMWVyCkU5l221OenAmlW+ma+yXxOmmMf
tzceEYhR1c1TVvGf/oxAUxB5ii0m5E3w+sYZWP99GvgQFVqJxL9xRZuuFvocYbg8tk4NQwI4c2ce
T2VmF/AyVTOosyk3lvjaQ0Eum83776gwc04Feli3j6Vkx3VxPCxWYgf05hejXkEZXpzURJ5Ts3o7
TlCTsrko9MrsKWKCBy17YfJg+xU4QXyHZhENIA8x4MeKN+gqB7cp9y4+VBcQUg5J6DeJO+wQrbxF
kDoen/ATs2iq1Ic8PxFsP5qJuxgNq0xXDs+uWO+Z7zSDnCxg59MtmPABY1CrDHCEYuVO4+PUg2zM
nkW/U9ahynZ8UrJKNP7yu6iSwUcjbVc2AKSWAy1M+GzQ/Diyr0skC8eddb4UBERm9vaZqHHoelkS
Sk+a4JfGb9HDIxvsCWRbYhlaJSkGcoYNo16UkRfkjJ9uKjQOciPoI6XSoVvvBsOUJFYfb3bt/bKr
6RL2TyY/Ma1ayWxZzKOwXbL+5sA3G3GjQDka5ht6CTwgWIQ6G32xe1OZFYqZUln4gD1y1GSJJ21G
9QbR319nN4bQOZk2kZ1nvbYrfX/0xqSWPTJAmP+DDOtnPamb9/lqtUGmg6IP2WvWwKTWWJAQVaMi
/3Nm4HJQ7Fo2HjJq7pk5C0m90lm8SqXvhwR9Rs9WMA6n26PXu3kxkXEAmu/w0J4QSp4nGecAr1Mf
t5hYLuUD4Z1Pak0iawYWBH1w7gdwDlXohg8kIJpPC2kQXm+V65TwnBZ2ju6BWslJPqMpEK7paXb3
Jb5VsUkT1lYwjpSNYoMXt/iH79tGTWAZKww3PyWrj82LiALiOoGalC0xEwRkKjAnearVLx38ToK1
s2eN1LhPu/wr7zjmX5jXzkcJcm00MBi5rWJ7UsCxUBHz5k1wqZ45CDbyMPLnyiwZOx2TZLuFMBiZ
fV3HtwD6LM3PKPxY50xcjioJ4k0ejSYUo7lr/3ocjuqWh4WLuoDGtL68A/qbSGRLWmu7fzRcyoWN
wbjKBr6UGtPqKEGsoUVjSSAN71RmCjt3Bsq3MrP15d47AqbxzDks21cbrV2DgJDw9+VetHEcX0Aa
NEgWCIduLtJC2npNVvMHRGkxCDTSUVGCdt4wG4VAGA905+ixe6DvssauZSM8wOpcGYATWA5s9DBX
cVyZm6cmw9yhZko6fnFtvGZFvQVzMC7bVOm0yIvagFnJyTwPSI4JT6XSzNOFXHP03UTLh6DKeL6/
8HCr5cMzByQK74LgsxYY4EflM1nmtVUTN+DJYXhb1ohxa/Yb/qFVskQyaIx/ORa8EU1oeFXSay/L
4kctp4u/zlb51CBKeRsXlT2Iv9sYxrUBI0fefSgcK6Xl83Fw4O6MGNhmNLmz74D9qbDwswanthwG
GcCKONMckyn3MBXz6Hok9t++OHz4pjkFAE8aBMQDTEAiMzIhcPoKoI3DjIkpZhUSG8Sm7EHpnjBd
MDgbJOtFoguQ6sek9D0fph1HfKG8ix8BjzRU3hsMcONq6xNAvKiXN6+0Cktppirve7Inp7prgihN
nctN2LJf/+drW83wg3ohSr58QWEasWokM9ViyMylScuVuSXtA0LnWtK/KIokFMhUqPXbNzU8In/P
dyHo/bMhVljmNgV+n7SeaqvAkmXWGiobRg8xPHcHo5Oz/iOF+CMgFCLTbA1bo5GR8U/IdxNitZ2u
UFTQFASg5M1a/hGLGmu7EP+3gsE8fJ5uJ7kUbVJz2QAo8+TE7FFM9y38IHpt+6Tw3BjxfKJ2JJ4d
OF0/iLVowY3nFzuqfCwmbn4AstMJnJzRWERpzcT3ezka3CmViPXplzDrBlSkwzjXuWPFmpjQYBHh
rvLOKSTafeFOn1Ptam3mRS4SEOO3JWOZym7K1qV/Yd5YyeM36iwx9+lLLzGOKdfjtQGjBQ9nqYeT
isUMThHBhDUxe0C9j3NrfkgkzQvDeSbmTPajNrfvDoOrNr7HPIYNi+HpMX+bBPorBc0cgqJTUDsk
lKiHztpDwUcphtVJeIeS/zh7KnErs7edElCLdfohtCnnrwpvk0OHoC40TznUYTQcP5ijxf1Gqp18
OVnjsIKM/eNbX62eseEcIInWYxdhZ6j7xqsYmLCDPvnOntxyjoIhFkPdyHBtqCikJGiCllImLqGg
rkyfas7wmOxC6ikkqWtLS5uscDKE8Shf1vlUtapm3gbDikSw9i9QPVD2gD2kRlNQGCfz/YEJdKrn
J8PK3xlUwp832qoQPMD0Fzg1XTSlOxh3LiA88Sh8M5SIrM1gHxGGM80/tk7e1GSh6pfKdZGtrsdE
GRAlXpbgkRnZ0L7KYPLlKl1NDOkNnYBYiPc3BNzxvj+L1q4EPMmJWauvtZOcYKOwHJZrCALV0mVr
4ZWn2GH9chuJN/IlQvXUkP2i0lQ/Je18IxFylbMbL2cPDPTnv6QIA1DEfr50VxQXhOEx/dXIInDq
Rxp48mDjNQmzvQ6XfTYDDgIBNzzfwamweu3J6FCcs1iu5WhmC2LorbZPQ+FJVGHQ3ByXumHG9KQO
uTIWz7JtXRPMHmJ2SqQ52ULohfdVprKMWVlhhKTiEpuzlLMj9KYW2esCQHkhCRjWOVXgaaZIyxLk
LpDeq3rgct6cWRpGVWv1ZKcw6LkV61cXaQlcKIQmN6mtSCyDc3ZGk9NK6wNvkpbwUrb4RldVU11k
jzziMW1ifL/Z8tgHzOefTo+WlN0ziOuUcbaodP/0LbztwYqYevOxpRMaPv3k3gUL4wPX/HP5mIPZ
j5X68iw9GDaF8b4v5Vclkebjyq2J9QeZXX6o4Y/f2421MuXoMJ7EQnf/R/a5nDXteEqlqitXxF3A
CFDeYSJrLkWraARZmRMqXRISatnhXmn6VUnNl+w7HK+fzM6qNso3Tn/HBIsG1uufmjmHmSyMrUU2
ihgcVC/8DZzxk40/9Q+TQv3SBrqcM5NeCXlJbqoyEdWfmcqmxLl2YtPSR+wKU49mbJA1ex6yeYPP
G/dunX2BGyz7fyQPqK7lq563QvKLx1Yal7UXvNXyEmQ2PqfdXruTsQJ/atwVdwNXHZYmkZAzr5Hd
z3Izs4w6ow+9yAZllL/o8LGTjE92Rc/i9XJ+fZf/Lqjqxrel+xeEoU8HJOz8gvrjni8aq83yzMMI
7ql1WmWxVD4a+xoDLgps8r1OCx4jpVelRwcP2hwB+dFd+8DeKHwwjJeS/iCl0lWbTaK90pPXN90z
0nI1fyZF1JziwQPS4j/xG12RegZjzBH01JRWUqYFHTG3hKfoA+avwKRSRR8RFZaXlEYr2u7frsp/
S3BgRCd2D9MRMUOn61fCguiPUIJHtwp9iGvxrUB2MSrcQgiH+obmhD8tMWvBOJ/+xdeQSiPxExw6
DYPPN4iFhivCW/wW5lGUH/pFnT/SbvC4ylLwMqONINfDDyXzqpIDJup1qWT5apxDWXCyF1uHZVRE
voFE850bT54lXP542jKVod9WhZ8wN6PaJpnGmbhM9jmI4dSqKZ0y1LTFOGqa+vrYBcmpvsWY5Fx8
MemGtk4gLazs7PDQiLD2y99QwSt9VKwUljGNCa4URPaCRdRcKrD41OS1DeXfUpVKEATIVWwwPQrk
TLDlQeuFn7YnY3foIJEKanS3kwQbz+iNBvtOHOhBNIK97+KcyoPcvKCuqIhUIhlumtBDwSqCZS+g
4RpdFV1PyT1PtkmJvII9/isWjEKjVwu6MZ9WsHdXrWJ3IleVcDEcb42Gs1By/AmHxQrj16GHHbFR
ag5ns6/NjmUtz3l+4QcfbeoiRuWCmgLxKysu5TwieKEN80f3shdX33ykc90vkhfG+N5zhsOIAQWj
iNJeW9xeNetkTV4Apt24KTRYsrumQjFlz3bHapBSD76WRTb204ObN8Gy0UucTHHUyqIJN91Wt8sh
g4Nury6eY837JT2/bsGvtOSrNfE6t0eZv3+vD3pFuKDz48IxX0db02P/PTA5MMriFAFzNmBynl6a
nALM0kc3DV6hxdZgujuiNHxi2/3AH1mNzROBabxWne4F1qIsmYqRmHzUDa/UNeaN8fMyNWtclwAn
+xvCyElODotPltQLMtPnj1ommWjMuNY2gzRKVkmckpB5jdl13sbHmpwG1DJclkuF36CqtmG27M2y
9hZj1WZx2M4W0mq3bPxziYaTR1sA61YaDit5gyW/bqmZSxegOYVb1RJChHzmxCSDW3ee0BEZdd0p
lBCnwfGoB4s8Sj8CB5tGJCF94NH2uP/DaBvibxsvRwB+MFsfm2V3v4v1sS2y1/jiobXtccp4BhPr
NuKCJVt0Lya/Hp/5JrKDTcJDy9V/Lh0xPa5jiOEWvw2WOyH/CGh9b/YWLZidIfdqMxxZ9vBdlde8
25C+9ZzRCo6rueVeEzxRaRBZrAo121wXVXZRvjAhMYbbTHABXF5Xyukc9Ypz9Tp5nZLfCaDg4uw5
hpcBxElNb2nCfZe1f3bJAjb70uX98U4eg+RjrO8FhDYWzT3M7PaBixUuuceyviyT1q7rrM/6vws+
PLwljhGfHjMamDGP6vIpDb/pwWZlVzihKW4JATQ9GnQkzqkHLxKRzediixnK14Ed2m9jt18MfvP3
C1OiKUdOyvZ8653J950+0VbyCVhSEjTGZv2z9qyv9892C2jg7sH6OhfVEtwkL2d4hRqoPu8VKMAh
CTioewABKoAC8SMzA4Cuf/CYy68Tp2nufBS6DrUYjqXwCGfyHkbN+y4D+RZVDcTKlhTMmOv84pBS
qpZzaf0QpjJPomSUgLQvrpVs2hU/tPyMXStfm5I+9zvn73+puGPpItfunaxqZV0k3N0/USOoZnu3
detvZEqd8PcP1kfX1QnZ/Q5v7m716iHBBXMBq9ddgN1GKJ0BFjQul5V3XHgt5C25wSM2jQaqkHxL
iE5cUYE0QOpQckKxJPHFXp/vLbQQ8JB6q/JulTvV1qRWU5pkxLnu+xuiDtnRyQFtyKBcT3x8xFrV
zK+ipebYFfy3Upr5hiHq7A2tOFJkPQsQv/ONPu/+8s4mEMVsPkXkmX9TxpIupAGrUrNm9W0sfkaY
p/6lEMx/cGdBP87ucAB/l41Yk+LjyFeeWMujJRjZ52m/ILE8fN2agIfBcq9IffqESLbaN6PWFBrq
Ua5iKa4Mz0QHVgetv2rur5KPSL7IYiCJolgL7exZa1IJAg6H1P4qEkIBKiClHfi2leKQAXJVZAbC
Bz7Q2zrKtLCvDsvZ7R8w+b6sKuliPIVq8dbJLD4IqVf8KOpIrVqW8yxq9LrC+Gmq/T1lS3WUr5kY
7UvFyDSo5ubY7jembNh/DzD39img+rieJxhyhupXzoVAAJHaTNE5XDwQA9eX12utlr1CCOjfwieR
3HcGzhxYo4bfljOHbsUt7q4IMg2e67+1tEgpbKN94eje48KwJ5LA8taNZCpaU9wunKDYC2W3MQVe
qwMkkx8rW88lsmU4jO6m8LDTaiigmx+xeNxp4DL+aftJUBaF5l2ShielDEutr9X5hqdx9my4la8g
ho95EuEenL8ttWs88pKBkqeXN+td68c+f+CXiPSgDV0KtSmcR84NaPD/fAcjEBlgQ2DA29FH2/jf
59YgzsdPVrs9cWeRG7CTK2OhOEKWRYk0deN7MFBzTkg+4KCNGnOJCpR51smd9k9cc3VjBO5FkRsO
VoCUsNMUD9YyKSsPhqAleeTdSvYMpDODL9auQ77tlgCGNOjPTLPvp+ja8L4nbcbbxIud9iwLj7Dy
5sldlgfCcAaRXWUIFCaE1YnoJ8bzzqBPdcVyNiFBizp9q4677uloEUNVwj8JDTb+hCk0awg/OfxN
xjAr+TlEDO+OP426FCiB1uc6ShoIOOsRdYL0xnXOUFfi/BGFNoOnpPFXpEfo+VmdZRFXvj1JX9dY
vu6W25GSKxV31svTuOkeMwA+zkHNDf0fC4WpfYnBucH/roqFXWmv57wjlECbxy40PEDBU5yZ+4ve
cMi/pikX5dKWOQKIsv24EOFuCGbPaLk8xVHkIYZsqKkl62H8AZf+K6g9WxXpF1GN4B0dtG9HWt7b
YXnKgqkb0xnj4vsRhmpNw4pBE+ElJMq5sZfyqXIbGIXotynxzYbgy8HXtCT/LM1VONKRAfkKhJKT
IZjn8aOTOZWJlr9LfY5wRcdyUIMA9iNMo/BDyF/uFSQxRS+iWT9cKYNhV4ky346hTdGjPN1igwqP
kgAqvvYOaHg2Rp10srRW7g85onuvtvYFv61pV+M+9wgZIikt1LXiT0QTlUXbBqhdmsT7vVuwzcCc
FLoqouBXPtNfAgn3gyHF3BbioKxf0o0npEw2+tVhJTB4Ggwqh+BYkDni6eKNCGWSD7vi0Va9NXQX
lG/v5GGbZUJe5/LtM0IFyeDZzOa36C9Ep0tuHJZClWek2YAhwq/stkyUj67NRj/u+JQ+Bj85ixny
YFDnL6ShmMdLnKkG2fUUZ/Pt612FnrI4uRGGDHQUW+iGRT7IAC5XJ6vIlQvPu5K1vusX3saUQkWw
c4CyopN+lxjIm/MeWdj2UsZ9BcfOARtz0P+KKUKDNnPAB5PkjLzMtSvfW14Fzvb91LC4IzvK/goF
57Fuv4dFfgttD9Uld+Wn2IPGrcPza9r1Dx+mz9akdw/B9N3nR9/U5UTwVvI69Hnrc1Jr0myxoGBv
q3UarX1mBdX1KAkMFBUWTw4pECqc9tlpcq8u9EnVxJpetrD6uACtdQjhf41Tyb3zSeARl4hICwrU
sKMuu+Nlzbk+4UTqpBJU24wW1lKqkoVgtOCjJ/ITx71xbS4eweSNKiU8llCHnYPndGIaDSUWQGnS
yCwHI8Kb9EkruPi9iS1cmYkc8uUHEKUXRZtEBorzGTxL/PU1zzUNw5i9yx0YZeLHg6l+HYagfkmn
3+wQeaJXM1DIR4ebAEO0OwmjXtFpK67tWus818BBvXLdl2HO4Pchv8nEzu792ubQAVKDzjAhQXYh
Ks5sjrpwcr68GkBbs6ot1Py+pqlDgBF1H2k9U+f0t46DtyWD7FjKN7SHpPdOP0hM6fa2Q1XcAkVn
2OJGj/FjoOcK0NFmcqKsse4ll0Zov0pXeUUHgVXG9XZAheSPvJolrmOBiuKU4F6Zyl9PudwNao01
dyTFcIDU4fDDMz8vy9tgVHxyAnfMsSp+UHQNJRzbOnHyn6CgntD6A5LS5qSyUbxXnokaIrRg0H1D
rlsjBcuUHMCNUGKAoEnQsTOtPB4EHalrzGv2hRClFvSbC6CGvL6xaIysqmktmVquu5WgwLETFlrn
X64scNVgyOZqMSQD4WV97Dpvf/wyEAafishlrRopRjOiJ9BiBgBkO9Dn910MqKa2hq/D/wStUBXI
fPE4NMgFuN/BHEc9FIhyATDIpDJ+y631HgZyhZ1ZYdF80jPJNgGCDeTDs/76uyD94MVS87Oyn3WQ
txNvg9He/FzlLm5QetHwEM/3HpIjZxprG9OHJcuGQsms70jhJBixY7/4oxErF0VLg0tfd++MKq/F
dQb7K3HMoYZ4SyjwBuhxAwHm3ZY4oT2izrenNx31j+o/r24GeUtqAf1yyDXPMUCe9mjUASdmcQ/5
fjr6AO+eLa52yqa71szxjw7475Hr40jVX3IpR6RXjFSuZ85Tt4DBO36IjoQBj8OhcvKNH5wb62be
1c/3MDDe7IdjYGWPQvEuw76BfkaFptQQ0tnBEGBA/hrC+OW7BSfaSWSVVjIfe97JOtV/GB9H1Vpm
IdDf89sHXaVFvjM2oYDaCiT84obiaLTR60KrcVX0rYm2piknw/zF3Zzalsz1Y+ETUotgd5UhEJhQ
UZHcyCtwPUcCG8C5L2kbX9pH8thCwWdTASLKYjah2CaO4/pobwdTIh7CR3Ld6KFrfOtMgxnVrZnr
NeKIFk8gzeaMbRqItXO+/HCIHxrz6tbKc6A7N9ONIpDUC1k7ffQWhWo5aWeXWbiidGVk3JVlU0W9
Q0H30KbfcxaakXRV03mUVQx/ilrAAFRszrUqSLs0hYltT0cCwTPGuHozyW02JHbN476ylNlshx1N
4EqiVTyKwdTC8EJBYJ6gqR7RinXlYdIJBWB2JjR5DfaNwG0u/W35czcaetiE1ILe/huXjYFf12ZB
ObFbl8yyzaYU7DqPP0e8dDDWsgUOvWVCpysqEfFN8EQ5JNrR7G16D/HyW2yQh966QidCi6AuVNcg
nwryoq8nHCHCUsLeTnvZxhzRvhmmk+XEm2eFaXemp+xXYZyestf8s33tV6AzWZU8zHbtILxpDlEz
QxjWq/Ppl0wYHNiz/j0HS9msLKRFKD1tI9Y3LTaGVAsqopKUlDPAiGMh2TRj4YAIQBWzvkTFy+HT
ESii0Btd7CFynECoqAWdpA4U4+G18zX/cg1xIVEoib+tJAOar9+dxVXi4y87nkTotPE7wJRRuHPH
VGQjGvnp1TDUgkFAfVFSAak1Mi1pD1Zi7X7m4E0CswiG6kTOLnz+ZaAtZ2o3VsJ/nrIeXg4CfUlD
kcE8ElzFvfCWy9UIZN8xMieGbpGvq3bij5sHfdTF6KHiicFPGfwXg8pGmBEn78Qcx+EJrLFDMu8U
W0p+e2Rm4MgtDZPDuGTYsLtWs+Ml0muw6cYgHLLsqovt7OtHOznU+0zIi8sWgB7SorDAvI2Io1r4
vzEM/4ie+CxkDBcLi3VhrDqDoWjlm2nC9gZDrRTljc8nQe3Ii994QDufS3DH7X2106D9HGB74gBQ
wUb0NtnuCvbhRMlFLUDMdIRVmNTcA0anNYz2N6gc0Ny4V73dX+94cHwVEmFbBoT5O0SB932L0HYv
Xh47gpkeBazuwmOoMh/wQeOFKCTso3UO0hQ10ZYuCjlFzNObpND9pIAiU3Iuo3JJJ46cv4BKHGUR
atl3DNd7wy/vMyBPDbdPIrkA+wSQXuFQ0G/GkTILP57S7kdIqtPM+Ep7MDwOMXCgz8VsvXHKk5gD
AZQV/xt2E2BT7eId5zboZ/zKOXIZeRsNIzwedIN4AdN3UEWaoHM1l3RJ7zsAIVA2W7EVRJ6Fuly5
ZE3WiSO88ou52fi4GPy1/QYfamZCT8xcSg7pvMYnOjIbjIi3pEhbyXhYAFXWkmQsroqAuv8eYi10
wwXOFgNIe97ffSCnK3ItWCcmUBg47Crzkgj3wAOGthc6ndLUW8byHe/pp31VEwsDQplm1Mg8swqG
Ou7p9Mdrse7jM9vwRwVuh0ZbYWlbkJnYM5o2qL7ZYly5QfctNHBBm723/NQ2KkMfMJ79VmyoGmkd
CIs4QIUFCJkXGNLMuzcKa9UACX4g7g3ApwZp6xL5qpvgjfpgyjOyQGlfcWFF/O3UC9u7tv8H5LQz
uAd51hBE//0jMQrB2l3hw7MtE5/nEUdAm8vNTqH5ePsK6LIELngPqdfYjSaBXB8qdaNAQp762mN5
M6/QMTrHv6+2R9U6TuW4Tz5qfQv4H1oV6MefuXM0jDWD8EdMQO1FaOdvQ6fbAWISo0aG0uCZr1QS
xp8TC7ZxEGcUcSw1ArdshHs3Ir4av1lzbN2bS6MbW/sH+OTSg7dTi2QVAwkRkZzyGx6Iqqf+HSad
WAM7VMD3Mw4dR2tqTBd8iYm7/hE6eTYtG+G16sI8MvN+T8Oz4ww23dCmCj6T00yAMYOjsUoLN7o6
1DMOfFKdyyxu0xwumv4BxWNb/ARWy5ugd1WfZL3gECfr5vFZ+RtOqqhXlkJk+k0aD218VwbYgSAL
EJd9gjZvhB8B+Qfh/Jf7OI/Hz4B7ZxGvH5VAHbsDtUOsz3RqKhRogYYQ5ahWa3MU4VjvBH0FO/WC
Y884nzWMsAcUud0Pm2AHZC7ToN4q3z4R995IFvxcjWXlEhKeVPw7ftNn4kTrjYjP2jWpzJl4KIkA
nq6Ei3wHgCo1Wluc3ZhgAhSzrKZoIR9LZxe3XlYLX5wYJQ/ixRX1F/mVq4ZwlHMYRjaHoKD2SMCn
ViYMz3sQ35429mPgEwFdJZemjt+14dMJDdtl+t4t6O/l2t+ibiJiMTCZu5i9nwhLoHZVMGncVYDO
Whz+Ro4XMhUC5KNcTuUHLZMqRnoDvDbc2Z0QKiiWH+piZjMWjjRVFr4JjN6YxCVu2LzWy2994Q1t
aS/vljAwjqOWxe+Z08yC88Fra6b1B8/03jt4oYFJbba2w/IzmBMl9/JUqcxmFvAg8tzHmOOWvlw9
OoByfR9+V/xzM68EfaQnTUxSvUb/OYcRF+/Ng8cluy3XLgkoqzygRFqQ2jEcW3o0PyM3PNS2AfIt
ApMYnXSGxIB19y4hDpIyyiSyti6cC6ZJRfNWPwCn4qlnxjIvKNbze6qvABw32dROnklAB2lTp9BP
tn74CgoENUAVuIbSto9pEW0S2BAw3rTjuI+LYsgn4Ru4wazF/1U8hEU6Z/MEJmncTbuI+SbGBZoU
rNMhTMvo0KbEAvefQi9yyGdsSUUH6gULLorvQHlVp/fmaS1jng6gVwSZ2MjzViRh71jRIw4gm5+X
t2lOxsrHzMHn2p9UTa/kZ575HhNVcwPPcSrOKbRNQkLLbdg3CrAf9Pmear2vq1iBGu+OlGWvazQZ
f3IDmXjS8X3g6A171kJyDGO+H/A7cRX7U5wBou4GtNFFbHwx8tGoXvD+lAAzWz7zxUvSsFbuwt8L
53lS7i6/36DG7QeXoIV4OY2DmF3Bx1Sfbs79GegVj09NalBQo00wm4fDGSyeALdQPlJIcqb1iDFJ
P4lKc/sJy9gXreE60+QOg/jhYRnDDBkES4KuInpypqwhFkclABj6eHxZ3T+K4Re5Q1rd2GIenHBr
UctcjL9P5cpr6zITu+OIkFzRDjrJSOYtGRUsxhP7YDgn79X/wiEauVzI/oUmL6n/sez7yL/dYZXd
uKaHO5vUdcwl/ZMbz3BSPZ3Cnemrjm2vsABOq8MtcCNZVKXWaOFrAIrUBWy7e6wRN3c0tyBHpcWg
3suXTRmJcmuhfrOf6pYrWvC6BC2sDVUSP/6/OWrJT+Jy1IEiBQFfxzMcbkkK6Zdze7wvZynVgPj6
54Zq/hrXWv6DxvQzwC98MxJRsDp0/UgEf4w8bunmnx54TKTzvfXmPxGLoGvTVSknvegI+rUSFele
DTh3VyTdXclrLcedUjGfLD2r5iMD5aOFqkf2VnQwfBNfQQ8Rlo7TZUKnTeWDw/a/kFMLbb783vvG
kj6TPGb91Y5/kUdp43GQxP1dqpAds3vsEU4hTpfmEMlHwittvOvuXQXfanaLkaZ8JvL3EapMite9
qLvlvtxi54GIYWQ1v7gxxBUWhU7Jso9HKn8HZZ1kToTsFQlMxukhXrTGnZCyrpo10NVz/6qHr/1b
FC6wfLI5jrmC9R90RHhNekvNByrtVXhv/gqTTq1O3tYKELjSZPcEhHUToC+h8nSmLNoMqh+ud9R3
x6FEbwXYO7ALdY7+I0ybzaH6k94zyc7eUSJ+kCMbIUl3Jzh/oUhRrA1SEhwJLCSoRZVLZA5eWHhK
7l/ifFTovKAAmGADjWinR4lqjq2qze7QwGydVwoyrdm4keMkWfyiDkw3JqmxRGACYp9/JvEV/+3s
d8mw/UfLV9K6D/G5w/fhrev0Pr7LLCKSVd1XzigByOF6C03Y8Zn3rI0Qffa77Qrx6rmJaTRZBK4j
x0FuDc3l+Ri8DAc1ctfcRgZrX9LlUcU9edoEOBt1mKGCMh3Urcf/9VUPXQOyje0z7YxMBJ/54oRH
sfyeQktgnwu6zdOy9T8a89EBmRJr1o0TMSwq1ZORUrSgBlzYHuhq0rOIPoZngSWfPkDSOqdKZnkt
avqupfzxhYay+Dqs/4AXVSwn1vjezS3o+sCmcORfjZlQ7IzPrlYdYAbJstRzf5Bgh2XcwhdS9hyf
AxtYDQwXHrEWi6BscEMoOWoTMjry69KPf3a0lU67O8wLoNjf5mTkdS1oU38HZgWnqzaIUesZVHM4
KkxQU3ILDimSgCbML8JBrn///8jjJuFm3Fpb5gQkceps3VWTF8JI5tchA4fuUAXWdZQ3ZQrpBugL
Nu+jMSxxhGKs4DriWigmD+3l6f/7mjQMxhQL8AI3gX/yGaw1y/BDs5xdGftrmvBBvsuhpgSPDIaJ
+fHPcCNFyR319famkswRLAcnM9SBvUV8BECH6VnsLaSn2tDm2DG3aLU2by6ZrhtkLyCxEG+vNDnV
nJJbrVBuNlzpL35pCGb3lD0ALvYMaVgYXPPtz9J4uJitfjloX/y7nn7r/uEvrEB2gFtc8rYkH8F6
Nf6T11Fsk3dDH3747UnS2JoqHOdFZDJrxLMsQWhW6PKJ9ms4BwzIY3yKkKfR5yaM3fdPEb1uck7M
fBBSaby6kCCxHVek6vcTOeAGNFZyn09LwJ3XmRmBAxNMF0nTks4sFOEDbIuFM4PK68QTiF1YAFrH
1gD9KBcb7tx1sf6WuqnrkB8B6/jIzrGL+weyCB18lnnVqcnIgbYPSEIq6GHHnNazRVpEQdTxRKAc
MaS3oUxxUU5scl/s2YjW9/ekUkjcNBJRnd2nQ/IpRsD1sDAy3OxVOg7wPK01YYvwLkcRI9hFG8zY
v4Zf6S04KSmMx/9OwOHkTiwFhgX7Ihwui6lk9RhrrSgQK8g0LCi5D3i/GjEGkpx1vSrUS5zkKncY
OwzGGs0ud56b0UvisIrBaqUFUv8VG/yw3X72yfujlrh3KmjYXbcCa1YAmwx/bDyYzJZ3XIH2K7CF
A/JK2DM5yFSvBBqGVLt/FPxNJYWyH/QXydBd/KoLibPYULK5Yd6YIZ3RpZxTyBv2PpKh/N+/BN5c
nj1KoeXTyTFtW9R9m/WnqsQLy7Xag1l47YO9ZLDqwHP17EWC777uI6xOyaVwNUk7zwBSiz9jvDF7
4S+7jMHvMjhrIjq9Y1XUXlNbrdjMmD9TGsjWlHbUEL9rcz0ehAobnj8IquUifcIhP+cpmS+d3UZ2
lW5hn0ZxnA6YUoJzNWhm3zBAb/qnqtz2NpqgaKtR0tpy8kYxyoq+x/J0lQW+AKoUZtXTMgdHk0hV
ET4KzRzCV2f0gdyabqFEDYQsCmKjrinbNRhgNus+Pao+Txv+95dFGVGSCmawLGupJE+JSp3AaaGf
PqaBtQqmDiQcjnwAtRvqsYp7O/5Epx60294BUcSyKeTKlkdqyCXJswcdPpOZqpcBYBG09SYs7PPo
8xmpkw05RNWotfhtRVOfo/Oi2BNaTnEoc0/hHm7v2P5TmKTlNhIum70G5xLZ9XY1Z50dc369vUUp
7Z7oyGvLCHEgCPE4X4jEZVTc9PAWpG9165SVg6FT/46ain3AJFQYe5DmGis8Bmcu4ee0rfYwRQVB
zboHd0l65ekj5iJGzpKm05uLj6d5+uxjznHZ4bPI80FUpSZ3tbuLHznPD+8GPgxI4q8pExTWkgXI
gtjsl5vbCHmyCJXcDozRRSX/T7Y89ySXTjfJdySaD8tadFpKu6ZA5fK8bbjgqbAq+CFxO/j4rmTZ
ZS8NCgI4lW7fGodRkk9EMwQ2bHmZHW6/9/DvK2w/5JeCvdL2Wdf7MFDvPO53/0qfNdOUjbg4Nks4
CadeohWS7RN759xCOJS84LwDIfqTAC5hMOjGZq9jHR9/kscjxFwXWQ/pN/qBMpVp5Rdi9UsIw3vD
YQzk4XZx1y40azX/6zfjVm92Ph10cVQgwuaE8VWS5yhbqRp42BtuY+apbB1ooAqV95tq2Lj+GjxT
MUTYruqiDe6mB2cbv/cCmXCfxnn2EY9rSRiC5BPeUAmNI54eNItwVCu27+j2+CGc1U8ZRjZw8H1p
CL55D4LdjaDKdPkvJRwO9wFpVkVcrI6LK4ci/NUgkWsz2dSzNygCiQhwjMIpJn4fOfYdxUBd9SNs
OovQguiegWC1fzuWWoKYMavUQq7hPQ8WqbyPPrNTJEjXEKJGL+Mgv2b/Fa2N9FvY1fZUHIriw+1g
lDEOCO8IX8jksudvDxANXQuKtUgJqcxceDwWhAh3YY29df+z5L9D4PaVXvJrjMLVUccT391mju+T
JHNCGOwGVaqSjBqMrQzW5S0IM7TvLw6VTQRUGO6qQyVMEclDaUCtnHIFGR9bMjWIfJUd/cZTkF62
ytMimH+Pwl5P+XcurcG7V6+i00A8ip8u5DR+uNON32e+7O0UOzBmN2JNNm4guJ7ZjBLQ49reZze7
Cp0u7p52FViggjqb2PDc46C46YVaCBdMcIRLUN6L92mpO+H2ISQZ0sl6O7iz88osNx4YinzgS3Dj
7fXfCAARnVHeJPT52akcmEI3BVfaTnhzNDvwmSNmc7vNsD6gHPon06cy7kFd/J2oRnMxg0ZPVX7U
9VIxYglvZQyGEucogCBeaQZ3yAIlbtVGY9qTo5x/itdiSM53HdrOR+u8uQwSPZqCDfzAfCD7SQcm
Wu+tzKyS6dcGlYV715nvsbqm+TumdzgQ0L5eXMp1yQjEBnCYyRWHSRqJ8TlGv/4vVUv2HrxB1TVf
RW3c6uGH6VEIERTAU3RXs4z3WBioc1PYSVd+9SUkIk4b3pzlbpzAEnlAh6vh5xDlzz0Rpp85Tc2j
XsRAOgQG2QPkjbxi2rgtuZganEDP1Sh7EC7Nsqgs4ELH9kdofifoRZQMSXfQIw6whsFjIkSzWx8h
LhH4HsUiLeMIeP40xZczJ3MUu0j7dz4+inEr560v1EIpfLIQSJaJeHIIa3CTisz1qObniykMSH8V
J/0f/jCq5y3CZrWj1AGRC+3XV3Rjpp6xEleHE+m8cRcIKBIQOM44I8tSXDjWopzhBr1047RCQDu5
afrSCCkEyzsDfdRpTLj2pGkhVLNVJyNgxgjaKGltFo9DwVxyKIu3Xpm/FjAP7Y9O7vglx+hrtvIh
GhUDl4Pk1pVtQzsOhTkaVt5AvqBRxgQvjAI54vUw6p2i+AFqPJmSUFuQLVa8Ex/5934pfj7xPncy
HvMIF5VZB1LCwvKKbW3J0wKIBE3z9PG6aWqtc5YwvZXLa4CTHZ6nFo6kt/dtMUsBX+UOWote9UAV
VdxKOk/iAD9UCVDaQLRLlYLDdwhpfwyS70iKEPiROJdCllPy0iJfylj/4/S9spZ2tL3jv5IJUbaV
XrPYvI0VStLgSZZE6Z0EglW9HpdsaWz2Us4HdDhfwpC697dp4fjMLayA3h6rC2V4zUrFKVYPsIZN
pJunNRqjussogySWYfdZycKqfU3GbkQMBon0LWOu/M+sWiM/lMsDDUfdaTGxzKTpp5UnKU0vqXZ/
da0WQ1d/ZBcRJwNs5Op4UkXLgRUv63HQn9pvyMBK0NmVXzrkTzi9cQUpPHzT2DN/gYt9XpRLhsGx
4vkMBiE8p3yriRWnKGfKW4tpQso5BDer9hl1mCzN9IPMYXzFsd8cqUEeCyN2Vz5dDJeRgHc8JRW6
/JVjzVt8wt1MqwYlJ+w+Dt2+2hihW4s6wpxoYnaf1PRJsojgi6BBMl7hCeX01CPw3yqbO7xqOOla
IaZxhTommgwYFrcb2JeRmg6lYuONEIgYKcxumaJkcRKvumW3NXhbLXsa8cRJ7sPMKgsndn0JUX/9
h/w/DmO9h1VGoMdihwI8TdtFD7cEjA+ikdZsy8WrJ9S5Uwsi5kcUhT83I/48F3lD+FBeBUb8UXTg
RbeoFD4503mHZg2vLaooyMA14Zeox8f2oyRKPQjOq4YZDPZrHpG9aUX0BYTKTwZMbKMc8WburjYo
u7s4jyhPgLL/nVocMjV2KdpHK0dKWPLRWFJUyVXmu/ziDo3R7PYFnnQlIWU3ENNV9TJsVQ66XeIr
PYlyLb2RHnLNM+rukOfOQTAyLZPvUiaVBZ9VTfra87IhoPy+oYlJ5s3vHo1yvmBjWOp0Fjd7fTtf
U7+jtngYzauhHx/lAVSG4bmzOFB/+xoGf29IM5zcB8LxexjPAhE/z9W1zJNgNkI0fo1Mnw1HrbyX
bHxcCLIV4jtCrtzFuuSHP7fWyCSZkv1OkKnTWsCyOuwS5/GoaxSjlVnxxnlVGkYj3x/SCxSOqKzC
v7UVPLXlqvivTqzwAlX71+d9IRLggfimrA0Suwg+65ItmwZ7eyg+9l16kxw/RfIA+7UtttuZHZYi
33HowxRh7QT1nB5qrUeeuNflnOEl2SFCy4SEd/rJtVfxSS8X1evghUVg1csu9Gvic9iNZCODq1WD
kbAAs6c1oiIEPoaEruZkYT+TZJMkehklVp74h19Llry4EKRUSaaIiRfbhs+FOMghjLw7+XqR5e2X
Ej7mDwNK0qYULaZN6gi4zinFxDdnz3QxemQwpj+1PmfElt3H4NfQVeIYaugBBV//UasJMC5foP3l
Q5h58p0jEGchO6xGrUHzPZhsJtXfbYfWv70XGe7q6/MpPg9MkLPzQcsNAPgz8jC2BIEW/Z5J9EyZ
Dn6co3ffBytJE85Q9XpWH9EfCiSXTaruhWN0PU3wGwV+WWxlqWOd3fRJKTX2OnRO+zrYxnlxksAu
gWpTNgiAjJU1QB/kYWyz9aTM0J6zVg5gLws4QTMPdIPzT32hRaP9+n5Hw4LYtzZpdezmbvsBfGu5
scFFT0O9zNQV33fHFt7go/M+fPNVwwWvoapfMm+fmqLzGaIICi1zH/PY6e32cdd4LqJBnGBsJaxk
g2AgwW3mLrncaoCMzRk3+XY1C6mZ6Ex7gpTxPK3pfi+1wtKVXWvj5NFLDupJo2HxOaeU/3Oc4p15
/ITvuMhgila0gICljV8R5T3X1AUQoOdxgqIA/j7CC/LA/Cn6NV4iPc4mzQp1pOGnk8GsUkcY5mC5
eq1qlUwU7ML+5sBfWN19KTboLYC0q7IoL8i2Hj7SON1LKrKr/vJWG1zXmAPQugmE8AYvg/SYWMLa
8y4oNHwj9ybaFs1kPrgSdK2biBm9CKgos0YlHfEkLQWQ/AocuKD0akFyc7epCylIhokQB6W59b65
w/sNZbNYgDbh0V7v3RnLU6al4NuVpIWTZCfQIi9x0/9JZiak10mdRL12wQS6qBdSh8Bep6vJLJyA
R3elLyTKDo0EsPlXQRq6oESxzxsYl+caDCp3A1sn7uncOaWBs8OHPSfE06KH7SWZKKCzGdQPbQiD
/r/FqP10jpXGAOlZyDfKOPrpq2/Go7tEiZJPIlrfOfi53siY1wxDDy77NWt2J6KzZxOCdS7mZcff
h/LaemrxQ+tfc8DZi99X0qrnw8xeirP7QpNR0TqwKOAkDFl92fZjGTsQKRHX5fnsQ+AKPyjRuHdg
qioCUbSk5lxr1FMjW1qodg0klt384Pqzq7tZCpp1g2+mO+mFjwYgt0VT82my5Nfj2JM9ZoKGdq0G
tsGx/lGdQmw1ctTB1W4sR+lId7Q7oyQMBj7jJDd8LI5Er/hbz1PJuu1TuD450E+crS+Y0sW9lS14
hwgKCktHF81iJL/c7iea2lC+AAGW2C9MXENqyrpUMUghxOTFRNW5Pj8wu6ndTf2b0RDheyBggDpK
oItUyvNDf2E205CJDqcc2qHtnquV8PUuB+eSuyseUQODWXBNjL4xGveBMg0+T8WCiPdBDYlWjeMa
Y1fu0XA4M3hGaiN5kmr1wAPMv/FG36zxTCvspYmokZX/ZKnsivteB82f3AA/9JJYIYfX0a/a6sp0
Vxcnvozyh+CsmVCQdLjd2h+y9Q3wvoITc4GodTClxLX5oGIrBYiDrIeqcKyasw5tBNG2HepEsZhV
MzCh/nip4qUv5ek/wVwmGd3C1BfwopBcNhY9UiJlOmE/YnTT6bu1o4OcjBaHIKEqdbxwm69Z1tGM
8MIGa8xMP17oWG2nKA6DYDOPoTTmazWI0li2ydRxWKWyf7ui1BAhjKAziNQT+qcPKUpsez29M4cP
/HtaTGGZLoN//pqqvip50PRrN+kniiIRcYq5NEGi0J+O1thu8VNaVFNrIJWXvfqhVG5KgFghpVLt
qGN7l0TSYqwzc4F25HFaQZV/gcpWBuWNGT1kkvm2fWKk39a3LkuOAdEOcEdZt4DxDLhmEsVWE+Mc
uxTSHZ47Azjd2xifd550c8q4epoQnt5MtqBMMtcHFcMhJvokCHLQmHjtNW67aARvq2pkKt/nXNpb
y0PQkLJR5Y0t8RXkhcWlvnTKf2f5iKx9NdTqwCQ5L81oaKO+rVdLh8qmVVyKRACjC7vBOBw9TKiB
hk1b4iXvViWPlSDRq+PaFHq1DaI2xVI4etJJk+LuBjT4KtwoNMipFhNzItrRzSmDk98ilt+Y6maJ
Wm94DkxUiZgf4Dgy8+Kv6McDRgr9nR9t0qJcIiqdUzMJQT8pPzpMLr+o4oyHNgPsuFNQLaLBOlYq
2Hr0Bifib2Bal/VsCzaRlcTCSYYpW11wzY1wr3rNnCjiCTOMQb0EV4dHmiDIM+MGDtdaYECn4JoG
0aSDlZCp+iQbzUGpbfan6BnNAfmnLDFwwlwCg/qwzWL4Ch5oSAlMGfvpv7WSicWOPSd4y6sr7Kvx
+XGY/iqGR6KPt74yKERJ66KkVDEt25NG47Ea5iDroxyKGdFQb/aS55g032XfqBEq1AJD6KK4m2te
Mmh9quz5NIJdal3LMtLEsD7NYIbEr7KJGlamGEmxr0HcYwzy5TODSFu0nxGXtyiWcf3HTqex+y3r
Cs8T26OA/smrngVuYF8Nk1gbjUZg3R+K34ngCxRg2SizrDoER1rt11amcuGNGoAF+H/VLaQDUFFo
h9lC1XgwtGevyo2QCWWJz0fEb6Yc5LsKcTPvFEiPie8D+rftEVNnBYLEZ0cZ1NXkA81fVTprw79O
5dbXM/q2E+IOOIfeIno5NocT3AsvaOh2u1/c4tGj2qbIXLdwQ/AX325At/8rh01k7PpphLBoLMJU
7HJ+nK7zXc0H5o8EIijoIdFDC957ShT4EfgHebvEpI1k//6kEj4TdDbG7F8Ei0N3gmlno12/7TBp
qSWSMQDot8gVkzmaPuSSWekefvcNswngh6+f14qr+sJeBGBrZYivRSUXj7dBrK/c53meatN1MOjn
KWUvKS/y19BqKjn74Q3DYo4giJJblj3Znnfca1+AwCFLZZc/l8pDv1c8nCQLs5jy050cMlhGEFSu
l+nwh1PDYX1TOXirTzW/5A8AXMNxjYcEQgmenUosvEbEMCvTtnsMsfAh4IBrqQKJtR2SQnMVn355
J9YLPyMdHGprVUtpS7Czsv+T3L7eJ7PcNyXH2pYhjXGWXDL6ojZ7LN6+AHyZtjt/3PSU/zWKLbKC
E0T07trqMHrUeqNtYCu7uaox98pXnl+HRqhQIKgkdxP6ea5i4abBpL11NptBHNF+QpUce9OhmHkP
87ssvDn/dEU4H1G5TSr7/38DD3jtvwVeKEVgUpVPG67Bq1a5ccWK52DAh4EniTRnIQPzKaxeW+kb
Mej7Zxdyj8SE9tR+yoSA6jJmoBNdTJmPFyVqZ6WW+Xi47M8sg8DCXJWowm+tn3L+IEEnq+frE1ew
MwHwDqy/1Oee5m3olvsKopL1vatF2P5sfsjRH6Qosj0iaHCh8hoQLwu+6z+C8wFzTtE5+BUA99iy
sl6/yWKeYOn2yNgjzh+DZip1WpGtrQWkhqMZUHbwgbpyUiA1chiN9Pr37RKkQ5/qxIs6NZcQAlZe
7rssuf3qJqEzuoA2HuE/t0vWRCCU+dCXIqmQj7/gz5mbB18Xi5aKS3GoZPhJB57iUR4YNnpA4aa5
rvBtBCrC3A/7jqMCBKfJvBC2UoqdOilhWXKrR8quXD9t25Q/4WoFh+CVEK4y665x+8IGagCDJ55m
GkrNEZG3YxTdP0GsAs+0RVqeTM8vulQEqNMWwzmoYy9Kc60J8PlUcJ/FZ8QuC0RigZw+/8AtKHQH
TpcCHBJaGxJ5uTWU9fw+2e3AqS1OiovqQ48dGwI/mHcXWYtSQYNjTelI3+PZoX5VZyDLADAHTMz7
1B1jjfgAvPWKEc6GqUuEfV8sZ1wvaPS+paelOT+zs3wHvl3CopOSZ1fUe/0rVUG13FRyynwtSBCn
JnciMIz4WC7HeaODekle+Fvfxu2E4AoqlbEUxIKR/kuHLNKY1vmhrDhZ+ScbTT8LEwIvnns8Ecvc
Ffd44ftYdo+CRbWAhI4avjVZCnTSXj8oO3aoMxHvudn3Y38bPtcQRVey3lfu/HwWmNqyWjJx5pl1
V2DSZrykxqMhHAdqwpddjNYnN2liT11V5lotpl/aUNK715T1iGvKi78yCcHZ7OJYIqH3Bqtx5PQe
xHrB6V9RRwJEt3w8fn68HiyCnT19P7XLJ5AB9ur0GTRs8Xhd2Ss9ozS9/b85io40aS0IAlwKPItN
//s/OINz+Vs1T8Fc+liaID1qDfb3AB+SuMp5oEJFCqoWyNKdyA7sC1v4HOe+CiFjQy4Elm04GGKe
KzrM1Sb9rUbKDcqBgVKymba7o5/9Z6ZhsOf56sAkOh9ajDcnqeiRN3vqTEp7d9sEnqgWTdx8xnQh
zAaQIDG4j83BX4J1Uco8RZUMX2cFDP9k48Ql00dq4+nJoXjOpebMJ6L7KvHb9b5xGV5urxFyOL9b
vmujObe4+ZKDebVD1DaZenx8802eZyU4Jb7TqpmqtpHWRjAYRb5cfQBTQZZ0EDRUnDQkf8AD6aLD
sZv05rghZ3oQGb6ihjBrCVjGhmtdP55R+k4ano7FtQEwHthPm1kJZP5IuVyO9r3My2xn2isxhCXI
0NXH8xKfez+Rg8jVTlalpHsgJj+PUlakjrNEJ3XPPmPquoX8EAnk8qnDGloWMYpcLSQvrwDKhJj/
5YpaU2pRcAsAnhFcUDaPCXiua/3+HPS5jMO1vOZ8op1SSS+7QaoWYcyHZdk22cboLnAbY4khAodi
DsD+qcae7P6XRXwExU/f73BFxSJL+B7CtSQzZhOm9WVjRf8iHUFo3YUtpmmBrUylrAC3UUyfn4VZ
ho20wp1+TzzBorag7D22HMLaw6iKOJriTo/PJRjwda4gEfXeIF+AMh5Mltnyy5gY7aqnu/Rf1irO
++4pg6NMQnhM+HCO3MvLGL9WoaX2fl+rfdzuGR8bl669a5xPH66ZryBSI/KQD+MzxhoM26pAPzoO
W75iVNSiotPQd2pb0AvrR6UW9AeeqI+XpcE+be2WfeFrHra0UzzKO++O9nj246v7GgM0U2g6Z0es
KisLS9DH4d9HDeiFr+2xXCyAHNsS7mvaHhUyks2CAiwysRe6gP9vSxIYFeddiajAGMR6T78KS56v
YGgbZO4hUQWKky8mWS5dWQdotP/P6snSPOoGGQSaEQqtv+CNqsL8c5YKT/2oSzeEWQ3zUKs0lKyb
SG7EUToGCPTiRtK4+yIRNAwhvFtQCTZBVdTa9v/1HuqC6rAt1B2uwdIVtvvEL6IaL475nVg5Lf5i
/MWPIQP0BPUflmw4L4l/CLHksGLoJGRv7woP9je5JovZiQYJnzUewfqR4iDcav1PQ+Cf0svQ2gI7
JHM7uZZN+/IUbT/Btb0o8/399mg8rThaFhgST3BCwG0QZ6CPlKGZE12PAYh9ezosiOrMybqgFqyE
lhCMh4c1xaP/8RvTd6fomKlIDQNrSIs8NEMz7d5lEJf+OfMytfWdUJEQ/TZjBUxmu+9S1Vue7pxh
ytB7LAIdwsz61gdzm0cA4Ytd5qPJ3F0NoJlO0GL56PlFLX4DJXEXwvvN63y8OSG1PKxpw+lwEM/v
PPJ/YEycHkQXCWaZcxzmL5Oxg+E2DhkBQpC/Rs/89xeGNm/6Rm8VCun9b/z/KdLOR1Kujx8aV3xr
bpCenQZFPNpXExHC0WaVxZ2OubBwvVkt9RHIqZsG7AreCwnC+KDx2z9uaQ2PNdHN/W9m+08cDgID
rZ8zmzpPwWCSGnjw7iHFsXPAFKVPU0oGdfOJICK6A7rhS23TuHMusTFwgoT8vfh5cccqoHDbA0pm
yCykQO7qmzaecXvgKQ3tTvXMmj5MtRPA8ohBZEH49v/mVu1YsSaH6flnSV2lNdrBmqRbUOM1qrAN
HO1dFF5itmY3WuZzvojUJrAfhlk5kFvFMRXrvkx7r5c+SztIgb8LllJd6TtRjyJ3jj8ZCk4Vr2+L
f/TQxb7f9uJ7hHTvB5SyO9AQMfh/az74KV0E0h2T9TSRvhQ7Sog/hSLCeQ+VZJaE++eBeaw4sB1d
IlL34aTPvVPQBmo2DDLqksZo8rDM53YrVRioRT0dXGxyJ4N7Yx647sT5tfVXZu3eOtv5QEblAHYf
3purdA7Uzjiv9ww8hI6Ra1a/Uvy/vkrdxATY1hMT18tlwscYRsM0rsPmQT0H34kzV13qj4licsOB
kC9O+jHKrafExDVUQnTrqrkAG/ifF3nzXGTuURerr3mONC5rSScDsSXQYm1Qvzu1/nfVnsyFs5wB
hHKR1f+ixsGsqeHSrtdJjYNzXdueWLh1HXpXVafPM/qIY0CkCgbOXAxSuSwPdfqZK8B5qvIhjUSA
Nv/IIAGhts9+oHuuWt07UG8TGysOHZbHRmrmfSR3t5ksG1/tsAEyGcHXgCuziPt3jcR74lRHCnbh
2MqFliLomSs8yfY5FsRGOIRINioEc/pdblEszP1fTa4rvZmQp9+0eICdcSCVtrV+HmTJvqZHR7R3
GEJ7zQSUs1pjahK6TcT8I5IEKuNc4zsKGn8b5A/qJX6/2TFZxzF+RpwlG+mnTJWVAAyC16KMI54g
GP96croETNIx2V3UODxfZscc4+O4FyqCbjGtgsic6thC9p5HyA+JNkG0gHaczE6sueV3sv2NDI/y
z1zqPpfrw+oB4IT4ubDdO7X7AoFY1PLQmJrBxO0QlKAzyEUXxgKaeT/mu6R0gtNljCqaO/pXiX3z
/zEsslKx+Vg/xAr4MzZFLaW66sbz6Wrg/AOdFzkmYvryLu48XoKFIc8RZvZIdTTmRaKam1poM/pC
71lgCfYpmeoC2WoxyCBhdKmr4mFvYafsxTMgb5yP5o30EjtHZ0TXaTByB9KlFdi+HZiy8lz/0DZk
dEjM4WOHjB1NU3wmqDSzBFcoyvDYgXwPnV6gxFFvhkp/IRKrHvzeC0Nomem2s+4qZoNmUqtueT2S
sRi3SGiCsvdq/US+3Ok7xaz/JsyeXlF9GX/vuZt9Zht7OgCVsKhf9iWhnLkmmb7cJF/vtKSlQcsL
Q+kL+B9SNon/LU/X2RTf8QauBwpQI39Wg4rYHHW4Cf3gQQmD0enrh9yZzbPlp6Jx0AiczB4D9OSP
JGOcod0W5QbO3vurQoslmW75MFybCI3drojOjmwE4IR7yfwQ1avckLTX/TVtoEISGLKQZ/yT6Zhb
5vbCXMkIHxpOfmceFTZ65ffC7TomdLZdLjkgud2SN6lYQcVKj4mwIXgRernZFQ0Qlayo2SBhUmY3
Tno0+zm2mKtIMatb7wemjHIZAlzwZzNlkGSu2tk5nwGP4ZZsdR+JH87x7vT9Dpaoi/PhEuJjHJZ7
lbj1jKETQLpze+Mg2Fxv8ykkoW71yktEbN7eGsUXj2w4eNd1thTZIbOCynXCAS6fLWOYi+VuM1aN
a5xx/o7nqJmXEvB/WqQ7LN3Xxurvv3S/b8BaGP41La0+WoxvBLDYvOzw242OAwTA6eKvBqTCz9xI
NwwuplE0su/s38FEf68RN2xLmBjrjhm1TIfKZeWVcXoejQPhv07swHHui9kFFXejxOECJ0+ax5tS
WyiaP+UsmZfrjCygp/sTchq99CzvJ1q3XQyh1Xi5AQrNvwSgILB65Cd2NJ+pz01Zw+swFiGw5Xv8
NIJFO4S/rl0136BgSpLDtovz7asztpHI0Wn7ZjbePgTC+jUjYV9tVs2ynl2jB3uiwzFnXPIESn1D
sPKTHqTUEkSfYHTTezINcWwXaCguHQ7zrB4ZO29fzliS/Vk5sMaMCko7Yu3z7sJ+EjkGVgMQXJGJ
oa+IGD+Hp5gvVquQqnSXAre/xwZ9WIgHsdLnrlWVA/ssGno0Wavkwq3OO7QXJCwa9/VQVUW5Dnq+
nc5mjPAP9n1JdAAy4cqOYrm1Zx7rWHF+ABtLs9gZyl3UK6XGUyqO25cHYGMUDWNhPQ9AGkaO5jAz
8tnkUbO2JQol8rONUmkNRxTPoL773MXQW/PpaWsps9AUJMSYy8QBUB+Tb6omLgnE5gLUnwVSg4oP
MI8fh1f+grGniRz+PO90bnZU/prHF1/6vkuMhSxjuCPsS2PWfQ4i8ccuu0TG8YlZk7gaE7vrm54X
p5gEpkKw04eAK31X05Oesuo5E9vwq7vpEuG2MhDLYR+RmQFZJdLut1KvqrVqGq/JR4B4+7Rk8jWj
AnmCZsJmD0ZbP9e7dKZfwJ9AeKMufRnaxVAddpup1QkhxVZpjTdEwb6OcxQc9pZreITojHQjJnfe
iw64msSz9MuyPZgEYMdSgKUxssh6MYJwpKjTHxxpvsNOnDIfqF6BQjD3uDgRuYWXNuDmw8Npw/rs
+8dAQkjiizQBIeiy5qTZvkOSNYwj2FDyO06d2evZzjVnheBx48+duwqj9+IOo99p3BxSEp5AW774
bDuOTBKJYhJ1JfkFe4L2Z/yIjkhhAhQX1uTeOAzO8qzo75BhuNdi041YNDfEqO6KSM+Uz8BR9UdV
w+Rb9lR3pqUefDE4O9AWYWcdW8Qsu6xZCHE33JW2x6/AbMEQvC8AJ3Tmn5oVrOgpqQpkI2UmYPuf
clDMS5/z09BI087X3vqMxYLszGSxmPLCYX2IHkcOYo1MBFz7rmuY1zFQD+UHXOhblT1odKF6TCex
0tXa6y81RgHXiMUBdHeEA4HUmSDCqqa4YcZ8MCjKO/2BLA1N4kLBlyRUnedlqP/6sf9ppCPTsf2q
gV7uTj5ZRV6aVsV2BNHbEpgYkWC/+OEbU1Yy3P6v2kLk7figbXV+sfcHVpfDCyZxspIqYXMNHoGt
PBTkC2Pg622iH9lFjf8vebnAPaeIkKZoXzkP0FPKf2auS9clzCKIrQmaAlzUsAztK6HPF8PANpe0
HkIDynhiOiN7o/2WtN/+Vuo53dLa0BXvAXnf9FP64aQVM6XMIn6Vr8MrkpM/drXd4hP+jmyD0v7c
h89zg2zkbCjuLcsIbb0TEq7gx0Hk4bh+9XDs2y8Irau7GJGFT5P+DOvqAF96XJUM+P40goThIP2x
KnvFTnJMnkJXHp9pT1jD/N5cPhPjmIIt9FulwJlOpQB7LgVHpJwnjhi9mjip5oxn8ws5b6i1VlwY
7QBw8k6nHXSh3GGaQcCMDOlSiW+9XU0cEF64ycwqX3zsCy1Nz+rQPNV8jyZADwMl2Ugzvazk/K3H
wEmaoBa1AwTSIWoTE1i4DmJceQGlaTIDvmUArCPrs5npIfUdeoz/jpA2YkxV8LvqHFQuuaPj+4gn
5PZH90u6e6WqJIF97eXFYtcTPABSti3e6Dz+H3/37HD+uha3dgGvYMQgrR5sEUcnJCXBqoRMwWo4
HRlnmQgddD/bpdyM1RmKotBhCsnFKCvxuyJ+3cc8jUgBErq7k2W/qqyt6+RX/uulEH3TrJldtAjr
3IflrAiOgdFJ+k8IWZxSAXT//74U52QFpPvvVkSFq3qdr9rGKJNhwA0/yVweO2gX52eAkknZ29gX
JcmuAd0pEaanCwN1IkHVNDE4jITuJqR0vqq5NmPSJzBpAQ/B+6Q9ZdVoakMb5tzH/KZOi9SytYQX
Dsu3soXWeO5f8dwwl/y7G6VmdGAEHOzbX8Dmb1DjFX8y+nYxj7eq0SxhZvwUTkvniOWEyHNG9LpC
dlt7lkg5T1jqpKIXeFvEAJMKRpJxA7nE/lHqGLTf7S8w/nnq1rGpy3Qxk8QN5WKzUsPKxxqN8coM
+s9VQSFIQiW5WeNdlomss8ObZV1lhtLrN70Q9oZrhp4I8f0mM+4n5qcLGnCr2niSESL/a6wyiirZ
U7eEw6H7wX8GyT+ZLGOz4O+GUtmUHT9WKXkV4VtHd7/GSUzhpXYRXCLWnN/6Cj87cjB1OAeWMpue
WtLyI0bT6L7fWCgWQ+g8ywF5QTjIC42dcnpIsG1o8lXWpcrEGjMjyg744WfZbpszyN/x5jzl3+Wu
VtaiPzVp+tbTIRiI5nXHW1G+i/ppW8nefa1w7NZGwobWZ4flo51rmRzLio+KcNEWPuC4z1OzU/5I
mV0sd6eFuGd9St25mD/IB6Y2y1t/hM/qhxIwVtdLCLnPflH2SqTg2PGiLRJ7PFGJwiJO1RGDCm5m
pmUmjAz8wz07yErqMPt2H1DRMgODbTMfARyd0+j2D/Ax+a3wspNR7NEB0kfHQXI7pZdaZSGMmm7U
g6217KjLRkkUh3RCdBiXKzPJQ/yUKEykwXLTJGVI32Rkt4fAkvaFCafyctqywWFRmZ99WtDfVNHv
fKlr5ylhNCsCf0oL7X4yh4CCQXocErDHnC9qxETVWE/Z0aB9Ixu7vJOhNXYrffg344F1lLMdMM6S
1H7jj+C9DcAyVBF9pCWSVVziYxcru74IqzU/TmxSu01QO0wPyExphj8sq0mcSRVL+aPEoq4QFF67
YSZqURmMVuBIi/zleomtP+mXHEZgAiJ4itQrzhuPo1uSF9CGS+PdvAHbW338wYYcXeBCLRwitsZW
t9XI9WJKnjEhln3REPJwhRtbPC5NZZ9yWZxquD3nSibnyWjH2T7PQ9JDj99nFbprgtFJWaSGCfmU
FegshiW3Smg6d54Pn/DW/LmRQ26h8xSxZ4s55Tv87GphdskePCuLztTcdZLVE63uNIErYPj38IDV
3mrb0vI/wr8t57rXC1C7kB36yGrzclQoHVxp+n93PX3T3x168hNz85KvgU92CtMrlBuTUA8GGAOf
23HplDD6KrhTBhApmhBOIlfrlcjklxSWlVzh1sIQFCKGxecpGiEbubhBA7KAVxTH1/fzKGLNFI+T
aSwiL6ixt7FcYamEQFZSfKzO4rksabwwsKHBymyaYuyvx/zVbuQ1oAnulZobQuJrFTTS3NG8N/DN
2S+36RNIFvgGbweOhKOxXWkkqjR4ZADQ0yoSK9STT8iJSjiUBs7K9ISxarjk11usFpWSM9kY2Fjo
an2s9ZZQIfgkaxLSWvO+sm7PdoX4YYkZi7vgHy2pL4BmEXt35Xz6s/7TAyGWBtnjAzVlit4HzERw
cdHoR3qWsBQGKTFKvfonnJtdpqooea9fWsycqdVjhXRhJt/kTfbdu7js1Qh8nYh/g1gaVvr4d2Ry
pRTe36rGZ9zTbgdpeFwIkAKux846yQXVV4k3bXLgVUtkx2qgb3GourH0EMRZAV/jfm4lHU9MVEpU
HjZph6DSrPVaqBp+uNsLkcjenB2OLDuF9naok80gCe83S5s9d3Sxbe9InIVHLKR7Q5PJC1y9qcpf
fSeZzgwBJTaWgO/Nr7Y7y3wVQtYRnyMkzAGhoMCBU0Hx3NK5u7Ss2Hwfuwymni9Oh0Ku+qv0k2lU
9tKBA2uZxpPE3xHSEi8sFM0ankUOpZ7JuxbtO6X0vgCvajXdA80TpykO/lUMx/KkoxFhiq0l6CJD
MrFNfxkAlzTiX8nROiaSUUx+JFd3VQF9L1ZCvY8tVvL0zTFTRNgnW4tyQMojj4au8pami8OhaXaF
Zteo95/nEPW97qqnl5tu1/GJ0i5lgi8z/fu0cxROA4K2pSbAQRAnX+VNv0G29W3jWImm2INrb5eJ
X7HG4+Bp2T6+k94pPdHq7w+DhvexByADvvpBf+YnkbxPc89ZqIbkiTZmvW0S+K6dEJvh56XJTkeQ
SIVfkrhT6foyUVZDi8tFn6bDFLgAGpcOaWTSV0juYmgmU1eHxGsuo7lBvXTE0OLxqaP7KOdeOgG9
nywYzPlqBSJVj56AwxuuhgO4Zd8xzqPQ5NDFhVizM3yIuvT9OvbC8rg0yl7z7zvrtDrZtrWx+Kw3
eV5rqIEQJd6ZGPTeOrB7PFPSRewJH4Xve3dqe84Q+BN+zFMEma5SYEGreidDPXG+uvRIPBU1+UgC
B+kQCNVu2hyixbHybQsXNTXU3MEmNrd9K0FgOfM3VNNKISzaBOe7MS9gVRhksjqlj4GxlWAsYiM3
tdU9WqbFxlt0GzMAe8lwcqaaJdD20PvnoRDAcWsx+46bz8oiIONEG5U+KXN5AzHtUzzTunrPu/u0
hZz7xafDtxS/CEuOEP9P8voQBa62xXXAZJ/N0tSfyNMyWqhSsiRL9y114HYCNhRk6I6QaxozFGad
3OyLqED/FxY1YbhhD6HP2C0j7vGOw5G/ekv0orTVBCHi5w2uZCF2U2jB+ISSI2fWkmp6cSNVPlIk
5HuzQZRq3lxTA/GCnZ4DXAMhoBREGVXU93tUl0l7rJEbe2AfV599tVIkZUEpr2PAafEpnn56K9gX
zbn4HQ8EEbPegjhbwZJMW6dYg55v5he5cSEELBW080vvl+0VjiJGdw3tnGy0R0lSu1DrnlDqvPVJ
WjcxmHpWuUw8cq1QXWrKEsFMXS6xh1g/GogHEm/gQI2nPT2zBmoOUYyxQLGauIH2kT+NVNt9mlxA
ZEFDeSYKs5mYtuMZGVwZQTWZG/I7qUshvQ7Zj0JRUURSy0sCh9I/+FqpP1scrGjvqcPPvXxDTBau
R6IBBRwydzzAlJGfCeWj2SsE8nkbW6rcAqMRcKF623LdCb2b7IS4iVGclNiPcLmGT4/FCWfIq8x1
o7AtTA9CskEG7Q+ok/y/l03f3xSpi9L09iItyv/9YE62jrXJH1qMkDVuXm8rPSO4Xw2KNPSGYi+r
AKlTkFnFp9oR3yuUfHhwZBTM18NV8CpmeaFNlJIu4V9gzT37JKhsnNn5ccg+HM0SDpl0SJhR9n8g
/F04CRiD9NF1MYYnJ8pytYVN+N16CbVX2aVhEpNAeD9P1TIhG9fE+PtozBFMBRq14INjydn+SGsE
X9ekGvl1sBzZjlLWNq8J8wkKYy3tewhct0+2QmbqA2ZjZRx3jzZYVl9n1dXOfG2VEpEYl8sEc6v1
bOLrCW46Ua6iTIwiFxqaPDkBFcfYHqkttaoJs/uHMiLfRKNEOdDo3kZjd5L1E3D2kvARiolA+h4T
8kgyPnng/iQCGyWA2YwYMJw0C7pASxaK7ynrf+5Eq6xoTMX6aQ4yi14htqlFvnZyy8gemaZ91iCt
yhB2A6PNN3L7E4QiiVh5tAyw8f+fzwibCgq3RTwJpEI8OarH0GK8HOaVsEabFuRQi4S9z2Nm2+YR
1YVfp28KTzueMHasDR7u+BFlSz9RAqIuxpfldQzRR3uzFtdrTrQKqriq43ow/HW5X6c5Kjz0uUw9
GcdtcaidvIvs/iErDTTqJATzjf3UR2oJreomqE0NbfdbZuMjdsJwa3zL+xh6OjOklgsW/W0JCwOK
1RUa/cZ94+tX+gDaMbVeJTFZehRpRTqQ0XHxnGxRMDYgBxnNnhKS4iOCLUiTWU69Z4jj8z5X4KOw
i8YvDehixeSq1nYKLNj562CnVBBtL8xWItcIIzP2tDiNoo5hDTiOJ3DRo59TDx7quD5DaLLXmf5S
Is6I4E2ZF8CzcK9d49QTrst9LBjuy6+LSBYhcBVLJou6oAyIwLY8Tkpsvvaod6mVTglnTnqb29I1
g/TJpNAJ6SvFkew+vE8ym0Fs87judZ973tQYnsZh0eqkJTBjaS+fg5YkMhOf5OjOBl9J9fEXOvqr
Z3dEKqkLLnOWbssDWH1qWMCU8z6XGDa5w4T8SlVQD3D4PGdlCer/aja0AFRu4z/uiW5mDM9meE5e
j1t/H8j7DM8P69vdhZizOmLAmWUCd8nSBvmLjvutZs10vxTRczxjZXl5Oxfxkusr3XsPLFD0BS74
oIJ/VPcpD64axBx/gAjLaMDKsSan14P/sP1sKrhJyzXr0XucPy0of63AdlpdBlO00V8pq7DeaeVo
5U7Hsak4yuEy0gzD/skeOUfkpXm9vzXtYXqjwx1FY2A8OJt9icoDuoZ56F7UzLYAU7pGziGlLqRL
pmvGKJeRVqTrfan3GYDzFMT9vKlfnbDUSVSW8FHuDo5Wl6um82Iwf6ESgbtZDF1hnd8lD3zwVcyD
6MpaRTSoyhjtGSN8sWw13Lh8zzuucNGqBxgZvufgU7qxpmR7g9abELoHmokehwAhElHrOklG+cES
0fJffXdgiMqYH/atHOJbsvElqkTjmFnag0DDs93QQIgR25HGkNs8TZyIMYYWKfVvuCnzp21YE1tF
FodlYSdpKNQV98MlB7IlWATYHM9VG53eYW0qi5z0i/Lu7EwCowo2FuzGfbgrbeGsDsEQMOAlp0HZ
9DYFi9evtlY50+R6iSK3yLXpwOz0y99CR2W2SJvuhETbo7FLQbIPpLLJ4xKvsd3xiIUQ58DzXoJR
idRrOsLplfxkUZvB/1yuVTapJqBKBCObJawgd5AfBj1PypvS/+N6Ia0tzM5pVoxDZ9UTgNZP1db2
A0qmDVx1MNuy//tjzucujJqnGRUGypxgqNaSWG+eVTP8O6CfSUiBw9o3zFx+D0b1IiT4kLQGpemu
H0apsEsIAb+oWjsuh3WfFRSGb0B6SXzC4tg1gQbWJBLgtY4OnT7HajxgHuNB5DAHlzfgnoe0QM5v
pu0GuraMn8vfC4ycaTq1cmSnVzxrTcv72UO6KDddIOGDL1+CrqdLriqwADVU7QMLhCVgty6icOci
FnsPfR8T4WDmoZnrZDzD/y8gIloixx2wY/6VhvcUKTkQXXUCFG3BfdDDYvu+fKkHN6cZMgsHkPUU
UwDiRj8MaCg5NQdIS7TutqK4qo3W2VQxOSGb9pSRYeUyGHIPqVA2MrAnPZw9Mt2eclOZE7YsONRO
yjxNNpMwaATLgEcNmaMxmHnNx+VDSy7/wuqxjirL6NYPRWRhR/oOThDBOlbOMS6hJNhsTA3YavHM
yUs7nz5IOqi4jkJPgcw6SLbUn5C99ynbSmj9E3SF/mLGvoU4FQD8ayAWXFjQ/uz5aKeCHPQcQIYo
kKS3ET4kCTQnxOjcax919QO/4u9UiCl/x4D4ShTo6JLF4PIFkHKUpz0bTXzchv5Acl0A67l/OBIk
tlDuHEMoZQzRym67kyU2+3uF/gzbkASn+yCfAWTjmacJb7EzMfelSOiQvK4AxNq1nRfb6nYif8dk
f4SKvxrafUJNI/if7K0vbs20UmyFu/gHqZh4H2tmZVTadoBwblkuJ9gUoQ95ktm+KLUoAaCfcUSo
rfYc10Ci5errSC4AQq+zCC6z2UAnN3mrTn4hEulgkvfsVbbA0YNJOSfsuUuJ5U5klb+9+zJb8E/w
/8p0cieccbnuc87SDg7zdT1IeVgrfZLuSnxCD0/eBjabdlYRFotmZHgisUkkakPVWoU8R+NJ1vIj
LzTp4Zib3MWjh+lkkMcT/XNfaxyMyyRhgDAYhyy05ZpArupJTKAOpEtT7AJKcsIcqLtZoIW0Vrpg
yaURYBgd5rXs4pG7kYSPl7bSRfAj2lKzgQvXGxJo4B+BooxPF6K9Q1/bkdSRepKI3oxiS2+T3S89
/iQkWVddodjlIDA1vWz16jHTmQBkp25P5elQRx1nvinHmcyV7bj6hzWd55XfQLJv5NMk/kIekEPf
jQkXJcCi4agQIkWZ/8lMVgsxCTM4+oV9wPkwWPV+FR1zoJu2azBo91QWIJRIPrSYw+ajxxrjPum1
GvAWfAs8jZsDrIA1/ckb3MXVnKzdxArbP8AP3szR+rrTRwbZVFAZ0ZO7ekasaxhkRp4dgE1Tt/ns
tw+UutiPQqkyLf5ogK5kdeSB04MgpS+Fv1G0FZaptpitfrGKUYtEtuw66DQY8uMlfVU6frg+MtH9
kXFQsEJT8u8/2HDWHj/kEsUcJUh6yACd7n1uTnpRI50m951/u3fdcgIgYDPqG+DDc2BFTdDH6loo
RnNUlBchnWXHPKMKFRb7Qx7JKsOxu2vpja6tZAxTVOsmOwh5PdGknmvLv5GxP1OiuMYKDwEF8gIZ
f9fbZ7bOM+c9uYwI9aElidRY0LF6XZkMmL12JLLldYPh+cmxwePbNP5jssrk6IbQ9xNHJkpuScGH
XQiv4jo16FSetbb5lqazFj1aNX/hBX+R5KDkoYMRMLTteSXsI9zWYEwJuIkk9P2s3wUf1VgzIpgr
Os1cGa3TzrwChBIuL6yhO+adc9rIpzTHwVLQgLnOnPA6WIR//F4/Cai+aESSHGdqofznbgM7UrvB
j1Ksv2Tt2QU5yqqWXiPyqzq/kkm5YcFz8/4HY/6KQ6/M4ttP7Fe1s4sDhYd6I4u9FsgHhW0VdaqQ
AV65QgwPo95tnY3nymb1pX75bqSCpDQLn2AYHrN28CTRqheOVW9hNrpC6crs0pl8z6BJLgCO9+kV
tDnT8WajcV5ngb6vquwSaSZXp1zwTGmEw7wyF7qMEAH82NdxWgAJCcRBqx/13rrp4hFPWuwg4QTv
0hdxL4ADObWEV69NA3aIwx0d+rUwoF0DErP1cQVz2QHQGBzb1H1ockj0WXV1owPjPpjSfZzHE8iJ
AAl7+43yLsIR6XJ/V+xZPWwlN3c89610ZYE8Lz01jKLk+G+CINo085A20mKvkFbLc46sYArSxFNS
yE0YYXbAOVLSB63exczHgdTYeB8LWaYqhw+Vzg+/anQx8DD3THyF0yuXwKDITdF+bjzUYE/TQBtD
m7UKrRbKUX5GTXHWTdGFd9YuPYXG62XTHw2ZoUoDPd2IUqnodDxlQTJAY4F3XYW1BmIqqx29F4Pn
OA7IJPKPY/RLZjpTgvTEuLyxYVTgt5cdJL6Oac3/cic5WEbNj+sq+xvkPBuXQPyDL3usX6VkdyZk
YN7brtL5ySOkiryveILDy/NnGaUa6CXoADImJJAhP7tC4TPa0ngBxRDU0OabgP+SRcOepGdRdRMG
jdWyPFarFKoYWhQxs/tN6pWK7skNz67Q6/QecVV3WM77xCucdEdip42nSbSCSu9p9IHDtUW0enEj
J+LOpRfesqDl4hFyzS4pz93TaTsF7/Kpgi9fyIij28GTEzsI1Zw+K01G2wcNicVb1VSXp+wiiA0q
Vii6caZA7qkpeeKWvmlXgVMI3JbHnvz3khVINAyKO8+KpB09eF5LULsY/4rQno27Qzy3pnpGY3WO
srtQ9ZQX1UmUgG3tsBULgGcj4wxOeTKpw+SYunigBhRqLDnfXsUFp5TBBcNCwVdmrP3wjVudvSUG
lg34Y+YNIyK+5xZf9iFrolpNqt2dAvhwrmJ0UiPF8BSwR58w2n1tdPUjyZCgczfxCoqqnfI1QXzU
zYaj+tjvJXbaJkkCzafoI8CDdMiWCdh8f47boCQXt+k6I7dtunL+douHXAH8z81ItlIzeP6oYLOd
iy2pwc8YxxtwTNa+6H8rdkkeCr9zJZbHflU6p54iprsq75O8R1vwUQm5XNFapXwsChJadY7zadxV
X/sfupszGPpsCSbeKAU5gg/33JEnm5uv2Ksx4TNVIqSmglc8b0aQUbIewZ0nrlxKIarSwS6hOP7+
1kE0YBcA87ZmXlR9clEI7ZRqD0azIUo2fd/IhPBjngMiLL78Qz+XX73bHUXSIp9xBEGuzE1yn4H6
dZKbvszC2h6VLDS470wncp21dz5JZxOiKfBgNpn3qNs4RvtNNDbDZrLG+D2bbt3Oc+6TutZpDaNQ
QuLqdVujHBLzx74oRzQj8/xnEz1DQveSw3yiMoI7Hvx1fCOdtjlZzgs6RTJuRsEIu3xplP97u2x4
3MT15Vc0QPNnxrKaSEruZczspH8FwEQvuJV1AXKk7sZEFEiokLfuIAr31C0dGiObTgt5JB6yzg6o
rUyRJ6peGl/UW7v+yfXHGOZpJvM0ozDohgPRfBsIfaDZFkSqfTy2vTqRp+dB9fXjaZiG6E2pVx/a
mZCLx3JZyNAy1R8nGFp5viRPnZdE0zS+62pXIkYEwUhCjn+xw+7z1hjDp8072QnTdKgLHBYtEYgI
gXwYhs3AIr1/BO56z1Bys2JosEZzqbqPjn+hmr1vnlfwnwN+YJb23N9eJlbyfekxPpt3BP1BEZK8
oK63sOoouRfQQ06pKTIZIeOQ7LQTZObpPCF6A5s47e5IMiQLJqYg+Td8G8s9p3TjSnS0fu0vDXU/
aJGWw0I4dVTKcxJHmqimX9qwKgZpDLaPuykpR25bB0i6OMEqUvNry2Tu4ChQO89KYe7sf4EgIgkN
tL3wIkPPCI1aNnsE5BZjePv5I1CP+wFpL3ZOZCWhYXkIZP/DhiQZwE+RiH+e9qyhQvHwUdmcodMx
TUqSThM2QWDj9JO77PzPqgLmN4vfa2wNLadIH9ya79Q2+w1yw0dngn/BZ27Zm5LMkzHxo4eEbIUK
lsW2SC8Lk7ZlFapzbdHJyKuYMzSdYp/zS3cmYehLrlix2oOss9SYTgjUii2uwBYFUYmYfvqUbDfO
G/HHEfBWEM2q2gGRonQMNzyAYLrbn41CMRvdnJ+QdQyv81hKezVsTQ9Sz1w0Wv7A9lqSsuZn7wOK
/KOkA5PdrtEwl4/03EIieull1hUcv0S688ssP1eK9NO74FsGu0KK4jRR0KNEeMS8V0HHNODcCzay
Im40dxBLZ1suGlvDxYjSZ5Et7L31l804kM7p/RyyuE6zpfRAHZlD4vA4SsEELScufq7cninSlH7b
qRDG2G1nqYVtm8Z+lFzMJybe+TifWPJrAqXsJoOaoA6fGN4yFuTP1g5AWBlLVptcTHea5AnJLR0P
itMcxJAlpoyhpFexX5HN0rsfHCAwMKfRBSVdU6PIOIF8WJJww5NIX8hr1quSKtD/oNq4Lh4pmuhk
p/UNkYpUJekGLNM91B6lP74lj3Cp12mmO7vkRdiujEh+ZyuBSdw2iGJ7Mxby0JaiHWx5WcjvNFb+
RxfoYgjteDPUrwdR3AfyfX3RtLQM0WBkE1X5JJMRcbBHemIOWjgVu3FM9ysJN7xe4jKQtg2b3E8K
bpPmzFODJ2REbUFpVrH30dtiE+Or9m2ptg4CUK9rhcL0jLMfNp7moHAjJaReM8/JH6RB6JP7S9tz
tsQuqsQZ1BMm2Tnrv8TLr1LS/jTwTv9mSSMWjhQIXJgYfLBKpyTojZv99mXi/mxBsKkqSm2MLF2/
tissBOy3UdXnnCquXRTkO3J1GDf+D0PWFX1FZDctbLud+4wS7Vn/q+qcJDax8p+S+m+Ef6B1qR1x
aSIAaV51kG0Kc2Fbjx6u425+NHiclg+RdAeXaWoUNWf3C19A4s1KPOb+/+7DVa+MBSeZg9Jp6phy
Xitw7AqZkB1Wmg0F2sjjOdpVDD4KtyP5Jfrfy0sSTmL6vXp/xz0WDCk2nPtrIbJ2dTXTGinPAs1q
21O9bfMzeWH/DEY8feGl894MU4GFFM5UIn0B0H4IEEufbbQGE2uwwRFYm/enDA3Tb9toHj0BssDv
6Xl2RkCbiJqGGuTdDpmDUO/IEQvVEYzVrk+/pNdqQXV6E9iyA4tun+ryqKtUVCfFCuMDGsijN7dk
6CJrfeXDLBeaOGlEVtcRpSK4r5/HFB1MBxRmpcTVZQgR5lhsenpgCR9ZjrglZsYNk69rW7SnWAtL
Uqf2uJlIsEOSgD5wZP7QXSKz01iRapcUb81upk8mwXzEoe0ZHAn52EiIY3AZRpmfYFB0e8bu3lAf
s+E19gWh7ivW6/h9UNJQ7IBWHqOeqSCqpMPqsDSKFYhDH9uFwSM59mvvYtqf0yG3zox56QUzj2Mj
8Rf15gIDxdYwhSXq6p56EwlyIWADI8ZWIjZS0pXvn4++cB4L4+MbccwuXgXEhmdxFBQ3iFAYe1iV
3H3H32EfEi4/4AFVKPB9KAGXRsuPzGbgXuiaXX/sTKp1tC30CmWRUNJRz0mXU7vXG827c+68jygz
U3CwkM7u7djBzMz4pipJggScFwUDtyxuG8fGKtNJUnKy/wUqDruz3NLEVKQjEu/POj4Oy1RcbSNO
kEHiWBCnDWANdjnec9uLipZHAv/HDwWZ7ceU11Hsuun/aUBeVo7t32qQhFQssYyoeTLHARLYTJ/n
vOX4m3Kq9lLpgYtS3FahE0zLHENejP2aTlRmAbx64YlYki86cPbPrawzghLR3HnltxR7xqK3esL8
Mqepr2nU9TAMeXPsvDjENItB7LVnbzFfPS4bjZnIp1DLzzW4v2sq1FGHT01XAhGP4jIHsldGG9rb
TsYpm9UhXKE4Jn5ClPGIpA3xvmpqwCRXDLZp3VUPBaajZTjTyws1YF9U7aarGjbPPQjOeGo8eEdJ
2mBb3QnedJBmPT2RdmwVsvN6nONENITp4d6rrzCexkR/uMr+KblJzqWiilW0gGbsB9HqWpoCh69g
/7+O/ffCskZAFKMrOSU0Gd/NPdB5W8i38VRyz15pXUtYrYSX5Fanl1kYIyc5cyHrqqRt/5zSusm4
yeQq9GtMVhuEcMozJQpWVWkX4rnxcZbYuoaXlhA0OEeuXVHfApaEuLbcTPTTxhmAzeLSF0FAN+UK
yM1nYpIUrvoUfmFwTOlKeo3Z5nZpFr9dRtNLe+cU7CxGRiznXjYtkD99Z1p1tWma3RROPL/ji4xF
x9dHqjQrCAdMd8PD9ND+4MECH24VhaT/b98TLUDBHEJ32jB1Z3G0I7f1ne8hLimQE0E1JB0u7Ogl
HA+UC4DejJ/qAi38WNMG8SHuYiU0b9VsN54yg6orK8JbQ3gwrhZyDvBCO4GK1lw1SOfrwKX5Us6f
IbdvAh3jnUU0yCS9xuRm3ynpDKbNr0wHRO3nRwmJMvhsbcVmJal05dUGAwbCur4NxeQFnVybn4he
vxcAdDL6Sh9xyQKV6qPVq/QXCfxvgoKp4yHDiXg4VEtfNfzL844ZR8yIrA92Dl2jc/7UklsIuy/K
83H8TQtjReSmdbHbMG0G2/TDizQupCr4yZKOGV7NCST1+0h61Fn51LuhtJ4zSvljPrvOUjVOGQ4E
SSzI4YEQYLshqSTFHDV2JYZRxSZ3daPAvajRx/H31xotCbKPME00g1WvB/LOKhxT5gfTFMMpg0uH
nx6JPwfPfns+Mon/3H82IM4mrfGp7Ez36S9C0GfIjrh/fDaf10t9EhFZa425ruakvuHXTHL1Vst/
cT2clNYNeyjjl9pW/CJpDpHr2uawFlpHW7SWWUAJcHNlIIg5JNb9pMog5Dx0Dv2tII122Jlj3pTk
+he5qnhC1XZVa8p1dvI3962nvMGDvP2ssy3qkVjRSr7R87hvrbcEh0XUgJobtALdTU4dt3gpWPQG
hZjXNaLJWGdlSFytVuUCDVQFTZsxDzO9plcZRZdswHIp6O7fSGC9PXFx/Y4AwAJALr4C7gr5S3Ir
5mDsjqyTh4DhdWiGrZJBw2p3CIyAYhf1cnVxCvokdDDGYgXiGoHPTSfDub9t+JzW3haPh5mJzsBu
sx4Ld0iehgzFVM4v4oaHoFNlr/lt4vg1oXgIpKDuL2ITA5/n7AKB7UIRE5CIRyPdMjtaOIis/Kmn
S4DYzs+9cYNg9kvQV93qXwu8ne4l0jyd0QQZ+CdGTcSB1QmkwJ+DlXBlWrCZq++o/qHAXpmHr6bw
wv3Jf9o70SXuZw8ya2OCohoy7RlhUdnDWOszgBvinrkwtD+chZNt/cyyYd6QdYfyETSY1vQOsfSA
vwNy+O5ourhN6o9GXvk/z4W+nihE5AiPXjPaVFPzrD2Mibd/5fMSda8ruo3XcoXmBc8MAbxuleBx
1+0eq2iUh2fc3HIA2H8srWy+E18Acmj+9ppSjnEfzMVwto+Zvz+mDfsu07H4wQ3BgvhdO6d5qOLg
s6mZWevoQCZ6ExT7AqBZIS3bIiUFTNYKISZs8y6S4CIgGduB9Fy+M53+yL4brCGaRuB/5Y2WAGmu
4HrpcRBbjUxpkDE+EknOsibG4hWiK/qBktRGg+7px0E4ptVaHRsNjUm9HuCuIBYvD34cafC4ga8j
5rTEy7OCIGDCKOzU5Z/IARhxcjpsRD+AT0GaRlSWWJck9G1MLJ684bIsfzUV4IugfEllWcyHm37d
EInM6ZPpMY4zx4q5lObfXEBY2yVGqOTH/YGrQ5IvCl8e/hknKZDOCCU9hh3gnPt4h7Mrb7/Yc2li
aO/lwPnj2ULj9TN4gIeaQTo5zkZuRUMuqA9RJAzYEeewQf4YJwKIBI08Zmc9p1wep3o13ThJP//a
4/y300rjPNNC+xxOc3lu3vFvF6Z7P9b26lEoWI7XcGISQs6T1WMc4mmP25E6Pni2+y9Rf2U/rUIU
YmdhBDCMfima68TmSfXtYvD3mKRk2ycuxIwt/vIbrfVa/jiyTQzNBTHt5ikxe7NmSboHtiHPQgNr
PUFWW1tutnMrr43RatUdkywThs81eR17YPbmANQI7XdHmkzzTgZ9FBAJvcVkrFQVtKa+9eCbik89
w+fgU6QlfIrbKBsogUFw47eTM28CL2LFcdYbCB6oZw/AdhKoNZr9rT0C4WfrVauSqt5Vm6HwRJN2
0KRXDVW6qFSAMYIasPc6gVoftcWaGUEbHWM4l02mB8KDgAGKRVKBuFKzMq1R0zE3DXoJYHC4dEqi
diiVLYVpiZO4eRFB4LA4z9mOhBURf2juzeQz8MqH+M2W5F9/GM07YhrmrE/Qj8hkvwALrfKEl3Uq
w/+ATJqYt5m5VKM312p2VWuZDK/EZhYePfKlZBb7zlPcCtQu153BjNI0wNlSxaTRiyQWWgVgix34
rOuon+3QbgywMlgOnQAP//U6GeMr8r4AiSTojz7obXzEnzg9SHoAu5hXO7e1KAc/5Lg79wbmBfWx
HDoEoC9SHkki98jOfo5hqhjshKJ6G+P8aM6xZwFV9/ukl+UdxvJ2f7x40pHmkuiY4lYp7XnN+icz
hCZOVrRfatge9ufXW3L8rOJzrIEK+YwRf8nglZwoj2UmbAB6jfcwCQvf09oLetke2yuE3khoYKm0
HvNbbyTcbu3NTz3Lfn6BisMkYtv34jpaaa3+ufrXIJdN28M93dxxlBtGROP0EASuIkabg43dlZRt
KU/jiCzk3ZppkkoSQa/YfGxHPeLB0l0qjOtWTwX3Z/AfXb9oK+5PWnmxzCSvHMhWJwwDMVbS6B7Y
0+4ZkpFQtyUjVCm3z610iI5aJXaIr78lNpybU4uGUb44tqHchiR/DLJGvLN/x3KhUgjy4xZ/zgL/
EJIZnaI9BzhRgmsx3qXK23KNnX+5j7TAjGLKnM383+/ol24HTQzSWxxcXe6i8ouL8CB6cUs7CQ+o
aulToRbZNIYzmAmyWWh/8T1mmxyvRAuL+23GM2PkMWyOBdz0w/EhdECfzYvEhZZmte4//NVTmXyL
wJhIpa/YwVvc0LC0UxpR2qIqBCoMq6CNWVD70WTFcqM+lj7wmVFjvFfFuNdx5xBB8eEtPmK39XCQ
z4PxWSy7p6XwLcYLU8YO8AZq/wyE+NSwS8PCyZlnD/2Q5VwbUIxt4uQZFmIFG9sXann1eUG57IU4
rNTaoe+t1sYaxVZydIpV7P4R+bjRgtEozYzJKtz2rm9EowuqNxETR+dS6Okr/zC0ObZIGYKeX4Ik
TVkvhw5y5FzULE5zf1apFq0dTG4WTJy8yyRxnAA+b/d0ht1d/1lKYbvAh6HXF5VnXaECUqxjqS4I
CRIne8YDbDGAFG99vvm/L4Bn/JChntF3qDO8gk5rRhbv0dB39diwsPS5FuAjQTKtHNC8sHe/02LC
GkAiRKizmH+BNsmjS16jsJNl5olwA0mhnxwPaduaEwKKszyIsf3u/96iZiGVoNK0m2NLs3VqOY+i
JJsrmA+pIK04e59hF2uf4GNgsNtg77R2JzuJLmzsZ5JVJSTRjVg8cNQtpJ5tfcd+iJ0513BnpANs
8iBzPR249ey5H0taghMPPjC+6/TeXS37tldNlmWMZ07zZ5JHV66GqVrr1HGP2V5bD+e+HYv1/atA
Nb9O1iiMpuWAlTpxRnvYBDe3pzHAfrSe1b1xKqdDQDRLfySzuLC+B1lW2RQ1QKnybG3peczcRPHu
WdfDaYGr64XNO7u6c0LUT+hX3V0RwSWiiC8/tk7Jc/Wee0A7uVQJbdSm9j3dyhcWtiSfbK3TCLhC
ntoBmmX1Y+6CAyE6KIjaFggaJ0avmSwRCgrB7a4RUpYV0vrQZLvjYYrksCTyzx44XHgzKldHBWib
XvWKtGzsGcWvir1URBaI3s7Dc1zlga2sBxPQWaJyHw9qF+wmRH9Be124NPWLhkCPy4xVqeCrN/iE
Mzn3rLq+B6RBmG7v77JWmSQyrAyGvAFJ/pV7JyioHVsVL4R+xbZiH3sVHZWlBKu3nem4+5UEdwei
dSR3ZYmHLGQRk1OPhCFt0j5LtU/Wiy5Za+f/ZzWw8+/qRJNYbzt4neRA7VqRMAoPXtcDs6EA7nzB
cs9vaqJz23mbQmwP2Bnor8GuRgFmsEzXF5TVdBYs6PicdxGC53mmOwHV4c+uToJx6wfZlxCpyl27
39C1/2YZcMhLIFt0dl2iIBltkpOzZjzgsrs/zC7vBxyWtsBoK6jjRSMpSjl0dPu0YZS5vNpq2DtY
xCzHW9b5BjdSLiGaTGMNYTtkO0l8c3cXLCuLxicToWHR/yV/4IZXaCvlMtxFlqprnDac8+UGLYxv
Oukoy/DCEDGeu7OtViR/TqXu/xoNBkE78SFkN/v5WNhEeR1QV5xV4JJtPErJcLfmeh0NYHLJXpcW
8A7k/nDNh2QxKDXOZPPvrY+w6HU3T9nvEzICb2L8w+yAtMFnWiwuQ/FttTrRss/nmnG7q8gSKLbw
etx9BQkjf5bI4VzUWhO7jbs6Wduk4dxP2qYsVjrE05uMPMm2deGMnaYZBjF7S2l541QDyy/sTxNz
3laaM1/JbaSrw574gsiNSPKo21/Blim5l7N2Qo1y5SMpRzzeNQ/Y91WsVYRgPu7e1rVsl+LuXOI4
i6dZssGX9R08P5yDUKxlGmW8n0BCNDnmbVugXmYCIEmfsy9m86AYUtvSofdrxhj+gCM7WPgAm5k1
LfAsQIXGPm5NN6jx0ytuEYH8pD46zERFXxnSaDbvQ/p9QQ2iV/OQDKoVTVq+6m9otpS4pLrqfq3l
OoK4CtRbfVMb4gOW0muX36+PpTcJ5B5+YD4tiv4KO9vttdN7q4reKRQKcaw3dS/6mcBPTdkYudPT
KCv2+FFsYGfwjcnp4tss80vXLDapvdAyM8qqQpnMoOK/Sqrj5lrwhRssOXDObqmDMy6TNQbFtbKQ
0fWz++Q7sb5Bk5eBLf7XplugtpbkI+cI6/yr8Dny1ITNnVVyg6Y8VvD1DSkWd4zGBCESsoJSW+U2
xCbfN7yDnAvQAst4wqi5a058t7tEp43AihavV/c4b7jREIrX6d3J2Fn/hwhNBfsjq5m3V+Dw7S1s
450OTVQ7tumbWVSlAGKbL69O99f+F0l1iPhNuJbINLz68AE84n/lmiuJUIdryKNvb6E35i12pTo5
eJDrXmJWBUq9bDmOsl7LlznsGvogJ/Itakbe5lLncBqB1XsafNdk4OKlxWOAl4wj534rAHx1Zltn
oAG8z06uadP094o0lg1q2XUpc+J8RO6FZWGs+rqQUcvTYdTi3RKNCIoMuIj7gGaILC3RWPpH2edA
XF7+UYu3jsS1M1lPuA+9XvMujjNSqxYWeFmMqQr3g7LZIm38c7Noqi5NCupzYCkNyP7o7Tl5ejp5
jANitCqG+m1x1AQT7zK5jfStVxOmS/WZ2vmnwRD/vgvCTBqgVOcwM03XhacyJxxaS0/lhlg9BWZb
4h+7h+ZFQFeVr2/vIBL4KNCKayw0w/uQ6ZzX2dhq+TJHwq9UWHePOvlUtLzY666s5EU4oHk1M3B4
OHOsbOjtoNeTrC2FyWhQNW/A/uVxnkng6mn/kCKtuJ1EK24vtZPvKw9N0/RJtfasOeSTcgwTXjFd
yD8G7NFAQenOgeR36AOkeMTxv6NcRYqJGVQemw5u4gNLtMqS1zR0BepTlIYLa7A02lvNkQJ7zFEX
0Z7kxtQgPVDvDpP93MnlQGv6lpbvwOVI87JzOJxj5E10saaQCnJoDowsCpADnO71xMWNV52PtQmi
9hMH7hzgDhwPc6YJDx5lBXSnKJRi4B4sA7JSEj4B5Ks+cmq+vFq0rAK4wUKgFA2GxyjFbzNMb30U
apck5eiipag5J3DuzyUq6zZ42Es2+/cWs5VnnsiEikYCuWDrpN7DHRa1yElMpxBa//xlTOrToMBB
scw2wx/fo315tOITxZohtSHkeH874aXtHa8U4bzUZHYSfADLlLd903SkamhLmC2ETmxcV1fyWFiz
82IOSkDMfs4ufDLHel6fRCQScWVxZvHHpdLLysWYo95IiR/c6S0DQFJZE7tg06JHRPHB4a/Iw9GF
QJjMNIC8IPwFQvmWzbF7DNEmSetHTEvSGPQFk6LCMEjGL5UeF0YNyqz/5Lx6Ot0C1WWYVTaHkx10
DAuJVqzqchOafLxEdjDefHo1SmWPIyOftmmlyRBw6iptJaq3ovCHIgN0WwZOt0Sja8bs0xWhn808
1SXs0tJ7GNAFj8DckvktpL5vTjIK3il+rhydCbki8prYOqAN/yO44RiW5wYEfTDzQjDMTmVheARq
IOE4u0uOFyEmooz64qcUMdVV8xZUsiYmIqy8O1YO+d7sHjGO8hJkyzkWJFa3QycRR/B/sJiLwXP8
nmwq3o2d5tiS1TvuTMNSyrGp/IsoZlNgcLhKklF43ABk8PyFfTYj0IGywIcK2WKEWYg87TcI+7nN
Fdb9/k2LvArP2cBfSAuShTZ2qoTg2Iv2VWWMZkTFqhVmLR62bEOC1o0T+SwQ0bMrEaODaI9B34Rj
ueNv2YSpOAaDjFn/+29z8WrCcdNCOpnawDo7ZVrquHskwVHAV5itdL8ofomGFBmF8tpTH2uH4CM/
yI6xW4AS7TvbF7Gm1Ty4w+SpmeosSU0y5FOjIzPyBec5loB1zaJvWf0aqkaaKLCM3WftEPsv1xZj
bNOmMtcOxRvBzL5NAAnbbnQhzuDKBCveoaFViakZ5pIBynpFiohKgCEjlQRoW6wmr5Vy0dYvLLT3
dLTndDbJr1RffwL1dAMvT8ADjpZobw38OVElPm5AaUon/y7a4Jxw59tKl9g38RByA6eA1POcX2kN
nA78XQyF7S2+35AK9g2eQ07nA5Srwm8qVtKILpsaZcv1Cac1TIHU+p+3IrTPZgsJi/b58OvYSVFn
tQIgEJl9jkt4UTcjjown2d/NbMsUhvnrKErJ//FPMOfimLTDqodI8ieLkmPO8N+cgBje73cDyI1J
hFgTfkjMxs3Wy6GTL3jOvDHsBARHK+qos34Lm3w4o0bcYjyd1jjBU+7Hop67QAqJKHQ3duk1hf6r
O77UlW2anqqKLmUsvIG+s+yURReLPTQ1D3a6qveJsEUiWXjzkbRYcwZ65X3WnzrZ2OlFOunWuzFE
EOpnJNOoeHzD7y8Sx+BZIZlpgirlfReBf2JGKeMSxU3bc5u8eoOyXIUGT8+12Cz2ACx20xYYg8kg
+rnJp6dVXDJP9mVquXqIqStKXqGb3GjBgsJpJ96NowqfxWEO36D87HE6q+uakXmze62M7+SyU9VG
THu6MXWxFVHbU5lgNIcOWrbF8rkvWUMHCoPhD4SrnlN701ItyvGkKDx51ZEdgQ/2q01DLe9MnOHA
dEKXCzJ9/WumREU/nDOnqw0dTnO5/ePGgkqqVpNWm16VCf9J6QTqUF8tsVSVMi6f4auxggVPwbr6
AHSeEV//vX4si1dkc1+dARMn0y6BYjkUW5hfghTs4kfN2NVvz7KUAZnEzY3W8kYWZP3bz0Bl1tqZ
OebYRKgWVjSOgV8bDAlxL7529dlBnXKL4Hw0HjTYQyWnz2ANpWoS6XMWX+LJubohYN60mPAnz3bm
s4t1AVrCJwBGos7Ms406pBlPq0jpvTYY4hNY6Sr4A4ExVhKrO5RT/1wOdh5E/eMxXk4vaFpxMcF7
iQT7iC9734oMpAeWZY2Q/1xPI7EOdyPlR7tzrJh9+TLvqZlnh6cKq1QvVuMF9+kkNhx5d8nKHErw
GFBZ4zViAadbY0oMFBd5HXvkoagppYazYGttNIwSdfJhJ5VmKWgiGGbu87l+HEKvp8aahrPAf/N6
URcLmef0l8x93ENMko/iLjYSUspE8qJNYI4mK9m6Rn1YC5KrlBFRNyypmam+irfr51xfIzd16ASa
zJJqUlH84vqUQAqkDZqB3AkSohLulKKXIoJSKQosEBJTH2kOvH7HxmEiwER6zDPOwgoN8uMToXaa
4sHASpV6HcUlUwIUarvzi31s1AEd847Z7bEOShBt5IK/UYXNEW+8tpaAPsojBmx7VKH8WDNJatKl
pv3gI4laul9jcw93NXmZpbyqNwbuFDz+IKYIrOvndiq6aJfIxy8xSEk+cSFwtIW72Jnu6mwMp1lD
I3ieCuZy2mwbTQhObfj2/JL28DBTbm3cs3sodtuTuOcizhgnNfLktn5uHRX0Zan9Zd3nw2nzjAUd
ujolU+VMDwr9Uzq0j0iXhMo+4K8jm4/jDQjxxKDeE1chNkP00PtKNyznbLCpmdPmXspbhAHv1E5F
ycMI3Bv0Qkk/BevVbzoAsuhrUrlwNrquc4AGeIq8ikoLjvtodIEYEB+ZrK6X11ywGo6nH+kuRkLd
GJtBRice3EDJv9hK8LSc1HhOCf3nWr6/bK7659AK6l3/UilQfHOMpQ+GJ6lTsqCziGraenfOSub1
kGFh7Bw5U2Ur9VEPX0lgHu01kaYGprW1rvRIxw7m5tSHRDcBSSxa/gzsHNSlGPz1AOaDXmnXIyYy
cA9rCRx9dwXCSJxwwdya9Eipou1lWORO+ma2gEOTs1tRZz899WP3iMcQtdkNLCES8rmtnzHm5IiZ
zcwOAraGodObeufKvCkodPtzSfQmDktkjqHuJiD4oUyG3rc5M3N8B0HdAkZxD4sdFTgEOu/wvhgR
xsh7h0O7wB5hkojbTs91G38K4sWgddwAvFAe+yf302JBdk5qmN8WSgqOHeGfMqHc0OFDPKkwXwin
WIdRRt2Ed2D40v74zl4M41T6j3iA7PIHuRFSVOHv8XioKSZwGSBNjTwUmmINlpc7XUJhZ9IwLNUR
TV6dimjvoXEmJnynH8yTpNbyrvVimtEtB/edlMr7TEHmToeRdyO68Mb+v3cfi+bhpwY8BleFgcOA
ZY6qgvxJK07bmT87g0QTqks6wWWDn61lq9WH779G1s4We1LrH+byruqKD35l0HmW9KG3QSKIUytK
Xs1sDU5Si/pUht6DP4aIREN1tk3CLKM1w89druA7Idx5/eVoGFJgQ5QuqgOjzqv4yJ/50tosVR44
qKdjVUBXBPdmjTRNHmc7tNLuRudct0kr3YCdFGD0Uys6k17SlFYWZ4MOZaJOc5j4cI++AgjloNXy
gHH76pQ2kVqBBQDMBP4Q5WCbNrZLZmqkpU1RYvKwvJVQZpmJUlP83gfZBjojF/5qRtr99HjNFn7T
9wSu4xZLqrA/JjJVSMTGKWlIpQR0+EH70vuRh+JxCWdwZgXeRePkhxrlakzSzHxSxneZu/fBKikW
5bQv5ckh8g6WTqPdKbhp3ie/Ri+ecLebbpixhRkpkPmj809jfurg/P3DPDX/OuiDlDaQEbXnaNHb
NfLe+GDbpHMRGnEi1O1bqjQpt1rKp2FWoZQmhQ9j89ZqVI+ALlivuIvUmZizsVcV25z1Ps37wZ/o
KOgz/VzQ1kkxzUyRyzMLh2BG97Ceq9+keZtgsbp5JBJUydJBkormhWuLPaWQprDwPuQwpH8JOoTm
GmJDugpa3SDY2KAJgmhJHnnV3R+SPXTzSsDpUUnp2Jl2EEtkh+KrTAYFojKJQ+dXCJTGt1QyKf7R
8iF24biu0BNFRjKuBGgUeA5oghHQfVvEUptIOUolrGTkm8m/69G4/yS9jMt1ek7p/JVmAGQzs0Tg
zEGeZ16YJC5KnoFtWq4+u5LKRZq4l2hLVDe5tDubHRfOCcPvKzxtdFaD9IbrE+GgSXGctXT7a5iT
/CG3OOWPz+t7YcF8ujvV3udwaLIMKgsPtwj5mQmDxZoDlwUZzJQ7DwHqEg3it/OGozqceWsdwYPX
F0su7ysKv1+UKZoIeMLZAbYWA8VCqH8nM0w5zQ1zSlVhJe5yxW63G5jQpshVkZIE2rqy2FpJ2plh
u6XDJpg6LpxCrxz2BwIpf5LJl6uf6WXA2aMj+h/TmTYCTDGc/jxYBvCAmZ8LANlA4zoQjpREuyfh
WxyRcJaLXycyus/I2bQkdViwae48IL0oOg+l33F2jsDNYJ7GgIxeFpv2VyBSREwHzLCwwiy+qqwM
o7aKWO88uee9iAcAWGhRN+vRijtzQLRuQv7Kajzr6DGwhZhhkrgXSNm0l1JEYFRIefequMrnOv1n
AFDf72hDIINYzSFZzMdgSsTZ8xrbk3M7PLH/pJ4r74W6k0lWvzixDcu1YHZwNXhm2tPK2UJ+DDgT
WNlsVsiejte7or8HvGPxkV2pxgDWzJDQcT4FheChvw6oMpzgSyMV6PiTtcKGliLvmgLNO3Z7Akc8
Igga8MqwNw6Qw8EqJ/+JDVyucS1sCJHpYMPXX2reYEz6GFewLpUwuc99gik45B3G2Co4bGkypg0X
UBLsH41lWzSn3W5U3rMmqhywUtLRtzv15Gj3/vx7YNUFXwe0lo+dtc+I/6FMiRkJ8KeCvBHP0leY
bIQT2e7jP9TdNJqAdHO2eY67rpgFSgL7l+eb+1U0bdnQv66X1HPtJZ5wLgcTV/Yw2qGHmZP6GbR7
G9EftyAS86tLnDTP53+gkHQBsdWxY68OjKqBObLkzpy2D2Dqib8EKEl9dztnMPaGvmGicBRXSlcW
VwLbJ4AH61w9uzvLedx4OPzqVzwaWFjAc3Szj7N4ArnPEfO74J2DiDt+eS7Qw5wr8yOueywiDEea
uQUQPM1vZbbvnUilUD9MW4ValcMszoImJY1pE8uZLWsDzjSw6Fg5NZx36JJM5E8VQIoymSvS+ejS
X6yS61CmUaYbUJP3hIYaMoyTbTxvS+QPG7Eap1wQXOsUUo0ti574M02OnkOlTfNlr+4p3jjaUbrE
q5bszlIZjZa5vz/j7yb3zyImebKvLmFj+9UAptD4vksyjHvOCRvP0NRaLktWuNkBXHHdaB+N/E9i
BTIKajYQ6EQOfoE9ak2H7LwZA6J5DzFjZ7QDdPZB8s1xPCER90bQHCC6m56qNakCbvdabKz06uf9
9Ba1ALnfjSb+6vG/WciROjwtodppHsxKtFapwizvSl/FUISWFWUfBkehh+maIemEu/j+U2a1pT4X
6wEgkPl0FrLA7ujH0T5CaS20g5e7tNBfuZFoJTFCukPMn2Y48SQlhryJGFXaMrx2AKT84cAZN9JP
S+wobiuNt+DE+BSTdXSgeWnCOa2/cPR0EhvMIWdMaMOHh6i58HLFYxwA9wQYJ1qeXRyS0AjdzLne
jpCdx8gXL8wL4259StCyq75dSfWl7XR2H7DxLzsJa3vIaCIuIEhWZ/Dxb+H6g7Kx3itHTFK3qdF2
WPYmE1SaUVTMErwV1Y01TjarpGNx1aoQscR81Yq0O6SFR+H2g5eDAuRuzaHS3ue55YUtM2BoMwez
AWh/uj+t6O9MGXC7qoegPIo1pGjxwtQv11f/2o6tyOuvcK9djO2QBZsdIGwca+hIU55iM9pp67bs
08BOClO9Yo0bytRWti64a1svdAfGng+IcnkNKhmFoxQGZZl11fbjaZrqr6ZPseqVf7EBxtXeBxnr
eqmlWT/zMb2o5wtg53Z+HeiGlPZyWhq6OUzOnHLgQ/7dGT87RWHF7QKAjwyVOFCe0l2JPF6FlePX
YhEOHqYVLWStdrQVu9Oa/rzn4vCcoE04rSdguY9C2vznI0aOlLoB4bAFnldtP+6z8R0ZvCz5wD0T
e5HTzV8DnOR0PIqNJ+GHfXT/CbmX64DOHjl4ubbX614ZW8ndAwRKtw+lUHeuwMEYgXZweYW5eGyj
P8zeaMAQ758NDC0kukZUbJxVfOoriHGI3Q+wU8W+5X1APQcqItDVKrDskGjkgSxbh3ey1hNAqw5t
6gARkIo5/QTnbxnlutiRgeEobaCDnrZnHRpBYdgZEHX/UuCuPa+Ouo+w6etKbsV2NE0yRamnyZuK
if78N2gEvx8OpaPsijW5Syu8GlZyL9IajLW1Tua5bBlRGc0QcV1aZpmfE8RN8RgENi9jTdJWr6mR
xX5ZbFNpjiXErhuukhbdW51bj+5U33dawBm2aUvbUB58kkBepMCdrg5Zd8SUxWDOGdPEP1hz+ovh
eIeJUzJ7Q9cT2GSHgjATHsuj0twpQbzDmiskMl1XR/dc0llF4XFvQs+tKTQuesw/Uz3QYUjYz6c0
iGmvH3A8xH9HKMh086P+osMfC5X4mhUo/VF4+6yC3dCLk7b8Cw0UOAGb6s+2VHWQtWSq5CB6m4ia
47AwJLcbWCJ0AeSqcdNGrNeTkcL3qI7KKxX2dzEe6nbumHPRpzp4esAiKq+rg4FdwCP8733+0QrS
Yb0CmkZSWHPVV21v7jaF4XkQ6YHl65f0kOhQ80rBmSnwVpAcoZ8dZ0KP7WP8ZHSG7T6DS7Dyqd6B
fFAi0rqpbycYcv9UyH/7XXag+RpwMqkaVgOD88PeEH1C9+sSvKIv1wmYX7wG7+5u3fPFB++WnNq1
qe5FzFT8NdyTdjvZg+WIkRb0BHiQJYDsWuFIkGVVjsiZ02YzqOIM9Hk5/S6NhqhNbZQsDUQta08D
kPMtJdLOwRXDpXLkrlmW48u9lMpOVCJUm9HCScjidUbujHjHe10quWz6Y5x3WLACWgKMwSTI31ud
Gl8Rg0bbW5EB+IEh16x2BqPnJtCu9hDERdjr5io/Rdqgp32M6obbViPtp0Rp7Xo9gFZEjZk2s2hU
XEk3b75xsVpSM+8OxcyQfKqK49faG6OmsUp+3a67x6gMDHacqJg6/SUvZ3AvYy/fVcyklrQmYbqH
hAZTG1vdan722fQgpr8i+GGcpoBLDJAG6367F1Xv5t4O9VM1FYV/YlDEq2kRbxqFlLtlpWSRx9qT
rEOttzmni5adDhfE+zzJj5wCOL1oZ+rowjFAc771CbZegEvK7/Y1+HILFrxuLjXHHl+KK4njvthA
Pksl9U7tDEHzBrhw3DYibrBYkdR5lDQl/+CxTpITXMCnyY8peM3HEjcxTUhkSXeLMY8ee3VdeVWc
0/fS4h3dHlqoqMyyadsWsHfjUnBZyXpworFsEjwoZOJ0ggvXHHTPMKLiHWuEp6uQMlZp08kBOfkb
PwGFMbUnB30mEWLhmORdMxJMiImw0zd4m0khHMpBdqkO77xwL4Mg47L1JyInE2Oj5C2RWZqd6aPs
7J37gVCf6zTv+V56nW3KN3aMrhg+UgNHgGbHqZmWef63U2MlJq7ilp5ngij2qMb48U/n0pV993MX
Va4fvWMK/884NNPazRB0h0Ui9bObNZBUQ1olauNJeBbogY5NZ+94SZNz24Jbok0rpkZcL7FgbbxR
OT0TZvgy2/d1cECE/+Tml/tM3e6fLm0saUCGFlIGYu9haLPizO0YrZ6bdJ6Ohx9x6rxOYeJjsUFW
9qfMcCQxbiYH0tcQQ5Rf25H/VmR4+o5JEbi3/QaX8Vfejv/XflR1WK2qArYvAYRBSrSGkUo3skRZ
yM1dF9j7jRbi++gpPnHgdyx3iDyrAgLlKIOYJNtpZV6Fj+31DSqUnJdaOyp1a0Ejexj8roucwa2z
xKXoO8bwTvXkEVo370Gq3ZpxoGVZgH0r9aKLUqIilBaika+BJVMRqRJ/+hr6voLVqcaKY1r6w7JN
79FdGHGxpamKkzfo+uSmGz8M+opkHg78OppzoWWlOnR3hfv3GSWFKzOBkfx9OMOYMshuoWdWdmFI
hsTqA15Vcua9VyYowkWrmKZLdDEO6ZPoltNERoiHUjN1n4qmUavdncvbI1hG4fWjlTT1rozckG+a
BEYakzUmoLc0RbY1Vrzx9ptAD6hRzP1yv4Vqj5X3fzpS8ZI5Nea+aUdBmUN++7BS8wNxfVLKDUDB
ZJuKvUkmBrScFk/uLtp61RDRgNWEBT4UwixMKr1G/YoKnbUz5R1VaJaHANi7UWQBNTbW1AcxRWya
sTm1ynHjGI2iLvE3//dgcBDGVBQl6bBRNaW7Eb8CCPXMpfNFZtih2GJqh70nZfmN9zS/6EPr7E6R
pwf9GX+7v4OQbhXbfdurRZLT055tlFmX6w2Gc+vnWfC3RZU5lKQGw59dVjEhdM+Bm1Pvt1XzCtI1
sBnQ/s7GKPdoG9hFIxpPvD/RH8UK+znTeUvX5/gFirsdvS5DSNAPYl8ctOUuLWUb+NW8TXIVfaW7
5pQ/hNeUtfAyMIxBYwGDmMAxaLYANE3qov8OW4jkFxuIKYGJHpvV5TOGemrvTgY5BwIXbKmgUVoP
7GAA/hHZ4DqKmTverDvitz70Of3ONYg4lQSBumVqYzWtNY8pqAKc3KP1GMveaAd/Vn0ras34cCJ4
iGzJBmn1ZStc3WB17jpcyKR0UVkEyd4PElHaSH0LZq6LZ9SOvHL0Pp89dM4At5k5BvfT3BJiuE95
CAJIM51rD9v5L4/9gXrOzWrE9XG1WVq6DrpQ/jMU4Q6HiV/4EC1gpkshdr2VztLdtPuv3pt0GCAM
lYl0MnV689owmPZ0Iy77IkN4Ca3pVgFEe8Hb2MCsXiMaXc5b4yvfy2M1bke5yMLUMbWu5SAKQtnX
VD6YXR33cvattQH7HMoaClAJqRFlwu16GEZFQ2B4u1AwXyRbr/lRCR6tU6ndKj4WzHm4YcSLo15E
c98dA7sEW9KR2RdwkWKQ8JWfvCwj2htNwTJW96OdiKp1AVghz+Jq0uBg/L5TnYSMVX2GQAFNW3ls
u09Mu5vBDIwuwdNADXdJp7DdAKmbMLTSWOgWWqya15NU2ju9BmJ3GJswSvmNML73Iws4zXpUrJkX
GRWfeEnse4vxNdlpHbIGbWykQIfpHlSQucs0gSML6OwspLX3RHLyinwM+EqKqtDESqZq99nv715q
M8DQFdLrw4DyaohZpe7ZAXyNYSVjyfj8BuCo3Ddibgy9ug1bU69O7zRxqQF2dLhP6CJGcjMX8TPy
tE3oWuQEbCpyVDxq/BeBZXYGSUNPgZOpG656FlirgbBUZxYMiT1x+wh/gsq8cPhrR4x8jjBM0ds1
JqXfFb3uLlSX6CODxVHwwvRth/nMeYd0b6D6GFS4S6d6WBe8IVs3quQN18mV7QMenqHvuWNoJA65
Q1p7GqcrVefj2n0PoAhXwURoZBOdiRqgrYdYAXjdm0ij3sCP2oJokiPAFD0Ei/cG8eq/rtPK6f0Z
iYloAz0OZhzvX7OgNdRxNS1I0QbsQ+Dxb0kizMIcCnraEEjeR/7gTkAs9/EYiUwHopheumk9twez
iTLdBs5ZbjTowEloqgurka9ya/AzWuLKZVHOPbiT1iYsLLQkDzbAs5dRJ1NY3GTIxrVh+cal5Wda
4XgAGTIGPtxYnW7qKu8emt4pEK6YyYGNkjDpEbtPZmWW42beHi5MJ0/RuGMU20B2fhyUSDnJZ5WI
82n64GIsI7DsTUUYWvEwj7xpS542BPgLdCeHOtJMkVEnNiOB2muidzdqeAlXFrtL9K6UPl9YqCfp
ynV1tCVM53nUeBBT6YT1KzcXgvgmp1qt8Co2xFow1GwDIcBcWNg3YpKaUsc1bglylCGhDt3fJC6E
12y6vYZyG0hxi6J5c6ADdY67/PULXE5Y/GZ5DtuYh3CuVw+kGY26HhuwrogwqRR842+SuWwPXWtT
HIUCnkCZcsIPI0MtHWGLHYBF6y3ocZWlOL2Lstuk2PE4FpQt5q6K8uPTnjH1A0AHYc3t8U4jB2fm
To0dLdiOcrx2F/fN3IfL/zBvH+rqgQlSfDOgCr++PZIMxWXh3fiPHzndkJ0E5Qqx1sAzreJW/S5T
mTfZdeRkzQBAoY9Z1jGOorJnSIVA9ZRyVMGhUzFiKU3WiqlUcKcOnWCmn/67EILyxDGls0ROp1Om
XmopAyS2QmTNAZXf7GBzmL9AElApK2RZQeh/i2ltN5ZTT8FlVVsZ8ZxA7sPmCOEv/VHE8PMpbd5W
nZeCpjJg919vHMSL/0it9vCrbB59dURR41ppK0pwPd0KZqYvp+eDts49VdPVcwICiWSekrtfS4hR
GOMVa1IsFXrUYYHUwn06JH2aSBgyl14vu3A4Xg2b+PbwtWqC1oUiOzyEFo4eI4+WyoGURJWBPZBC
VBZSYEj0mP/zuFr+PAW77opp+TVdwFJm6Ig7DipV8g0idzUm/32bBKiZcoeLtaX62zv78Bwtzylv
6MUhmY0pO52NEVlfQTUerL3QqzSrQAMsOdLLcUlUgCFTMAPKVLQztrQIHXQU1oHnluJz9XrQDmkq
NsgkIjgNViSDYhIsO0U6FmjsacqrUbhEQUeqLl6d8Ud7Blko9h3i9HWEFPTAGknhWd+Bo5MmTeII
wO72cCE8kTMS/JSIhU/KID23rEIDklPg2VdDWDfUD2NA9A1kJNlnSTcez3sQyig0/f6v8AvbW1RG
jn7Q7o0JBx3cpmf/4JLKrk6At1sspaLY0c8i5atdWf48gCgDKgf1ttF7IvwT2jwBj9znWZbLkSqq
FTT1WsvrBmX+opxJBI9qGF/Gw2hsJtbHa5QKsozMgnpNiSFnaTZQ3qrmm7LqpcPh0kPZqb37HtR6
QdM4kr0ms9Yb2bNhHHQn3cPoxRcaye8+Zo4G9dwaUWk2NG9O/YZ63AokWreNMmkF+sE1m5vj4eLL
P2mQ68fvLeNQCc35tWvhw9Aas2sGwnt1YjRV46YhzugVvCH/G7qhX6tDZ4Qa9fmaZ2/++BgG0XSi
gqssfUIF1uDzB4ps/VdGYpTPsY1H2dXsFrWdNvXnJ9pTLqio8K932jSzZdAG877Lx+qqm1b/2PJm
CmNLX4rokEzfzCkYZEPZNoN47CsIp+WM0qbuSyrGp5NCzFGkIMFI36OhREN0uoxcP5NGYkm1AeH6
3uwSwyzBdy0ASryeqNN7vvXBmqcjKlGiOEwphtF+XEHgNO7HauDj/BObzAWvuYpMstrzqLIoaBPm
FYI9dS3O5aIVsVWgYhfQWHOTV+aAFrhK3omfvRgfpTPs4HYqraDx2/zoHaF6oFvN262rkTCsdxUb
L+j670sD8ZggDtRnFhDYSNyabFbU/gE023rnbjxdI0H+5hIjL1Jg1KIdvQT29Eyaki32lbd6s37C
8ErnzdwdlL+Q97kT+smZlqXAKRtecMO2JyEIFHovIXGc/0u9HH+aIaxWPgq4FoRQHyoedjs5Ii/a
pxjXz5CHnfO7GV588j01SYGuzVrK+HruXtNR57EnuXCs1qFEy79vLfD9C0Kqni/xtVi3zFxzEloS
aUXSlp5q2Orj8BYC7fLLkih1dW03tEP1IG6txm2C/jFjFQhPNRwIEoLGQN+Owx5dx9XbqRqhw3l4
wu73c8tQAbSgLz2HVgXhQmzPpAMRxhmgq7qSoNjcs/wQg+/RozTHmzqUFM/k4MMNaab0fkoEFiI7
X4ScXOOU9LBLPy3tjGt4n4bM5Zv73KfQ3NYgdl8JsMszHHhZDMl55tZ9+/tROPy5k+tVoUdqXUEA
777GAGyKV4Re3OOZ23ZL5UyD/A0s8z2e4dftNlPgfJskxYmKhKyP2cVU3NZSX4CiEK6fxEOihgmD
qJUXKVm426QQa4RBDrlIrvvvjHeVa3zlzercNTNkAtIakpExPWFlSPJAKvSz1bXBK8pJSsDzChbJ
hoGkP7FtwHCoEj8W2zQhb3Fw2BKSMVvNkkZLWKcNf7t+UlAJzwkg9DjMAyeoaUV0Oy9ceTEQl5vK
MCGX2gQBFdOpYlT02YnlUoXAL2VAl33BuDEE9Jss4AUk28ftdmP7qusEcwkPVa72+IToGOEOv/Wc
CNh3hU5QIxIT3XOTS/AfuOOWrg2JiKNQzMTHmY5ztRWQt18w9yRbKzcuR4tsx7rbCavbGZvzdyB5
4L8Qyirkd9VdKyLnYgCWnoGiCXboGVpC4z9lYrVOjCi8nG39GLlpE1DV4iPulUMHH4ujssJIrGm8
QqofBRr2GhVlOUNlGWVBAh2RAaG2PX3MbrR1GXeEetY+VWvhppex4kcTmfhxt47SPTy1ysiRGlzh
uI4DlwBrQP1qkS0hXRrN3oEi0iJ4WBhctNpSZM5LzNOYnXDKVcBXxqJI19oCe/873L/y9OmlEBau
DGAz39P8U2tn0BENi+Jds76+2a0fGnB6+c35xyjzd9WFMC77axBCVN7TC76LcZxzOyyabebkx4t/
0uwK0q3LgX2+Jmstyr6KBAa/FbuaSFDXw9YyHzV5AbovLtmZq0oD758tyKcfnAM3IjNaBdD7Gl4m
U1oBCi1dLHVUJ0rUIoWV7gHgO97iry8IvqxnTXkOZ071q+WdFe274sZmMObkqvo/p4G5re/frvH3
gLnPtnU0y3tZsgtP4xseSODnYr24q3WFLEvSGZ2khB+45+JRrXlQL9BCCY8hLJ1GSe++O/xSsjRs
CImWf2mWPvbQO3dF110xbdGV/zJFC/TRhXnc8BHyUF44R9BiiCvb33AHRyxt41y5lGvImMr3St7H
owA4EoJ9w77oc1phjlALtSgS8mJezEGg/lVx2B6F83qoxVfs8sfXmUB1OsQ9FHpJBWjqbws+UDpb
fkXY3YpMVgnU3quKo52a0gdHAsbJnNVdW1OGFCO2dl2cUgGF7MzCrqouulrQDlawvKPf2XT349Fn
ISP5UfZ1Abwo1tPlwJdeZ1L8bNpSEm4BvziUcUVZiOMp9PcpRi9L5gDi0fd3t6mVWTG7W+mzGfEo
pQJh+AqHkvtKKZIvDUXsAkdMh9Sbf674JcTMgmrVgtPtstxZafEuXgp8zVTjf+G57KB2omcJ5cmL
lCMEe0I05iLLB5FinBMAIbfc3VFwNwY8963Jhzci9b6KWk0VbxR3yb01/AEvQXAAPA3mGAHjJqH0
TuEbIGmtDPRxEa3/viJ8m10d+0VfPhfPgjt/ShvbI5THa7Q28w1+HqIlGnjHjpVdTXsrJtazgNCk
nii4fJcL7lyCjmtl+s/4DAoxar4kV1H+NjIhuETiwkZXiBVeG4tb2Wj68+FyX1/pS9g8JBKYQ5kj
uEK0AgHRKeM6KrqImwAAcOWhKf5DUcAt3W3KMFLe64oiLQMxVSAOt4vsJgE2R7JJL/i+MDX+uQqd
qh6CzkAD5MOtQ+tRKybAFRzWd0G1oZBGfM3/yKwBTHq8VPxcHFGNj0mYWSVsl0QURQMcBX6d3TLH
mNtGuyaAVQL06oHGnInRGF2w0mxzWaafUEpi9cByLu9aNLYudYMZBi3lNIZppqowelZNzncuSiXX
gkRXYxRxAm9zBqSjKjNpSlCG1Qxj5gPvykVK3fGQEQyQrsq4b0XvzVp7eq6ywobL4ggFZH5srMQK
nnnRXGgAGhslWDhIJ7jcABB/fIU0vT6LYHxBMvouBUuz/zmD0vhXek2so8asXb3fAj5IKW/cCHlU
sPV8NJLFH7APGdo4WS/RspaE+eIr+ShNTwcZm2j5e7UYm6qdn89RonWX3z/tZ8tJNhVQ0dNLpGZt
76gZO8/kfEpz7xi4Qxg6poRsO7rFKyYc5oCB3FQR4/P9a0eQPX0JVpz3GsSXhID/aoLdA3tXzT9Q
mqazolKP4zzyZ5WGeUYp/A75tDkIk8FwhoclFeF1SGhz1owBIW4yrQtCSY7Xb2qCoBn/U5cV72Tl
n4mgTY1GeRq28ixf7ZpFbLGhq1w7KqqGZy4e9aqxE/4tUlO8/sHz57bdWKMY0m87acaAz7weTs7b
d7QfHhWX4fSJmU0bN2GHiOXMIdv8tsppb7JOs6I2dwkZcOZbpsxlkecOSQ5nlokdadi0Zfdn+MN2
ieyj5ijZwC0U5e5c5NbYD7GaISAM1az9q4oRwg9mD4on9MXwK+iNbaNRbUQlV2DVQ3qPY7wUikwh
pWB7iJTMSq6zpFoh1dewyluqa5tlU4WPjvrj7lwI5l4W4elpRyWArVsw921ss3NQxUM89BMbI79S
KaoO8UHqW2jSVtTC32z09RmMXYvlrgQb3R8MMm1P82rKdxh/NPIdIeUVzRSrGi1dyrTd+NlGwBOU
+No07Pv2CwOj+D8RmsGBDINgVYEIvz+O51hywuOP8z+S4y5e0vRVTb+JX5uJIayH3v1OsJqnkWHk
iwgbjacPu6CbbkxFlssD5wK/shH3C4A+obxPiRpLGIzBQBILYx0PAnkHp++OFIaMxF3zkVw1uMSQ
9Gk0iidPf9DZqs8LXJLctbIsZmdGDDuzin0W7DmmFDGvsQM9iky0QC7IPFWh3BN8fkN6IGsmGSjh
866i2DZBO9LbHxfzl3FNJryWnAFYuWTSNHLTJzMCQZSNgtp0+XF7uF66FAmsp6YJpc+HFX1dL2Ny
+kSgYb34KX6hG/vQ5zUKlufKtRL/H871A5CquSlhAY4CvsHAaHd5PFWMnvBZLv/ZXa1K4RC1pMFi
luU7MvVVq6/MWD56M7cl3PEJQzr+u5CgjrrDQILtQOuVQBZ3eEnSUT8Ti3LmRTW88Cr2Ne3VQ+wV
lJ199S+kT+vqHDa4qoAOXwOCSzDOWupwXv171R1MAQNVvQ3TibGBJVL4WwOog5XjmO+kCYA8r8EG
RyvWWV4K1N1sJziul8jRXk7+FUneu9fQwVa2pSnzSy2p1+MtDaegSL7zPofPpMKKD7Uy8QpsBu2m
XYI2h9WN8xJCJmqtqJaPh2EYl44ofdP+xt3690HVIlXzm8At4CPOrH/8hsLp1Twm+5v329tVHEEX
xg8FlLgO2orjSkdlm9wHXi2rEyHGZbQWAcVeZLuhJE57yOiYDSjRc4l9jdRPRzIsStK/iLJRABVh
99laP3JOo8Xsg6dfQoNcqoT4KAtfNMUjvgHPvQJiJzuyCTIcmXwFuz1dHmsIaDF7UiupmigDP0g0
+maCZ60TBDdKO8sO6HnXsJCOFV+Of/CSsNzF99brtsYdFpjEEQWlQcVe6mumuLku7pvHiOdc+uEl
qYFWcBrQn3BcrQMraWnXtmuI2DSa8kNIsgYtRjYN8oy5/mx0ANQM3bjJRhj6unU+L5mDPkVJb765
LANPOMke4TXSyY8faYFLHujQW+3TwJ8AIRXVyLKsUIuRX4f9RlxKr9v7E3LG2OgJMS059bbOOMAu
xPHrfbeaFnE/yES+22A1fpNVHIyDjTQh6MAJ1HK/NPLy8kYIVDOhAdyIwONQPARfFJY8pQahUbdA
zxjTb6TbeOxt1MW4rkE4UJ3WFX8vtkZBF4AzOkEZSFVJvjY+qYLwHqYBXtkbu/QUZyVnMq0Trxu4
oB5k0f7hx9TEOGQQDmJKDJoCa6gs304LlSkEKXKJYSwlwc6sEx1DCFPJSR7dZ730RJYluAjW74Va
u8n16f5UQCNat039o/a+w/vKlD9DCZhoeAPOrrKC0yJ/9qgkgrPXb/3it/2dQk17yqq1bqyDuTwE
sKPVj1swW3lb42SWYB1OQdfWVas4ZnBF2SaJTvgskAP6brhwUw3SPWdSvrw3Y0EbYj5ibKTAoZE3
4WGXuMpXJwsLljLo6A8I9YqQmYqeTIKs/0yVxBwTwBfoj4dFhK/84cdrYfBLx3Ns3J1prcPgnFYo
XVajMgbTP/uwzx9Xfiy9Zi/Js9MNMw8usVhIZqf9QgBszf64cvkXfTkT45bghy/D2bGld9HWFa42
0rYtFF6AEW774zmhnKGH75hXV05LbCujs6ouRnDA1IogfALad/VPomBOzPOjNRDIkb38JSevGtx1
rRDJB3NwiVXLCkkWawLiTa889urQxO548cBJ4xqf+UxwwtO6e/rxaDEL9ccqSiTrwAq5ubq7POfL
74thsveGEko1MJtO8TUkv72oKKpEF2FH9kNTMgZXvDlWjma0TUSwy24Z/w6sOvs/XYvR6J2a+iaD
jnRrdVHevqT/dMnnzICfKo+NflADJCVQxHAw4KU7MIxLB1M4cyQEt07+SB4dyXgv76LTmJwTqEoS
ZQ9A7X7UXhX9Gc5+s3BAC8lLp9ZaHD/QsJ9lLuNyIBeYaIyXLsS88eK7yNmljw5SuufyZhmeyyoM
V++USsaK45qvwp3EAbj+BR7jrQ08HcqEmoxah5brgHzgyOvroAGLCBgtLqAwn6nKLn+FZ21s/r6D
+HhVPWwdnwJ87gHcms78lHUPdtK7IyT1nbmrAJyX4aMkEcOYBIGdvQkP5b4th0yrdmkAt8++uPoF
9scR+jjPvmg4fcgkSvtXl7zDIVEBhCV2YKhK0M7YKFg9IxFs0MibLb6MXp1aos0bUSAjUnIDfe2m
mPXteTraWnoKokZl9XsjxMFmiqDawdtsod6JmPSa6JBfyH+cw4IQsbKYV67AJzutTc0qmzcwkJoT
UzLfdgP/MuA8vqlk0ALCVDxr/Aba4kTNAmeJLvaqBL6saUe0tEZTyb+eiophAcC5rCSPszWNo6YV
wrMtV6Z45hp25g9OKfuuIdNIxhC+427tOPxFkix8/+epXMIR63bf5+sUQzYrrvm2f6MiMfCaLebL
vQMW1bbKRCaaxGQLhp9BZnfxdCC6YRtSt73wcKFqzQqp24HCnpOV6/951o5m4lq7Lz++xRRm5Jgh
IGg237APXjqdRyMSHj0i661CwZMGyDaJAaavAiT5mapQ7vt2KBC+Y5/meKp6WDlQsU0DDhjz4EcD
6031AZ1UseH2RAZ3Jo8xdQeFT9ZpatA/lO0UULIPRvvC9Uy1+7RXmJe3kNSHQexLDVcvxCrxlvYX
vogVc/YbHscY1On/EQGgTv52xIpbNqQLwzmOv8GGdrK1tDz9X5nQN5fdlgdXLt075TYppVgTtxHE
p2hWOUR+cWd7OusLnR6p/z13gT3FKXFPM+8nqEXaX8JTpm4UIlrA1eBnjPnaz6XvKneYTuXJw7eh
8Kjiq9EDJi4qf1B0WI1+VhXjt8eLGmJFB1aMgHgbgWFNwIoZTTA7P2Oq7AbAhjzOp8CQm32MB28v
lEyUGUFVB7RKVUcbzDegFHnvShklyeqwCpJSGYDnnjudJVubpAPsAmfiv0B4J1xy0pSMKHOqIAkK
vWKIlXs97SaipGHx4vcF5ZBB4E1zIZfMpho/Ng6pvFqSX+JmpW5q4QhWw5prWmeM0o7tDrebQYoB
RF9FAgL71c2/w3oINlY14proT1Al78FobiFOhRgcQPYG5xxApb0GeYlpRQo9znvgtMR823MOwY2l
5Ddgow9a0ofnNGxKY30PFQFtjzLGdWsdV6+J57atmSRMNJxyTfIpK+NzO/uaxXL9ncZMhyiFtpnU
HiOJm0wUqyMzpqK+8qdA7dueV9hyHGfUXVEvOy+RWyKLAynwU4zdSO3uPuf/5epIOPcvEormYmoV
15Y7scsIskZIkNU/Vg/wN2aWk6YlxjJBX9Uc0YZD/hnP7APbfjlkVWLl4Uiyw5Unt/bfFw0k1IGu
hcLG2icG29wYmtenrQ1XOQsLXhXIrWN6QQPgmnOi7EpUoG8yHzMnIfNSQyakKzhEoN/7X9e1FoOm
P/3ZPNIBSoDSzZb+a8o+prmN2WiLedbkNsyV4YHZzWrDgHuRaDM7AWpN4eFHBiyw8vuQP4X0RSOa
TNTgmvvc+oe2RFlVrzf6BQIY7IvgK6y+wHIBPzZKBQfmgmxfQTyPdfa+0nrdeq/s7Vgi8DrhZ7Iw
mcZfctHv+ek1BBh+iTLhMhTN1KMPtL34xexNjIBFpQ3jZ5LI+0ldrxM3oDNdMTRaYmiw6R9dEnJU
YsjQWpwJoPhftTY0mcN1k1IzWTXP3FET5wnk70ArVCt0k5hz4rH3DL8RDYBlwjA0T7LLlSUgpFFQ
9+iB0kr2ObXtdRFdj0U8t0l9r77wQKIpvSiATsiPm7xfUD2wi+fHHD2R3ZLYHtJoNzZKHxJxNcNn
A7fgHVWdzQjeckC2eV73YH2Kclw/pktnCVmbY9KuxXOL5hkfCo7HWxoP+EnpRkia0MKQLEryjkuR
GQnW9VYLxUD144gED7ClVOl9qpXbJ5yI5VILkXojWtsTH9OaLVIBtrye6WjuA+TJHJnVoZPrXi3X
U3/HZXYaAipFyZZ7b7QE/B/hNL2mNPzH4+UcUc4VklptNqrfAdeKeS8/3FNW8EEfSWLnf3d4Uuk/
2LHQ9J0OP+eYb+QERzFTz1ve9ojF0dc69hvPuclbw+M45ovg24b9B/4voPb3BSfsCDM+1fiAzmwC
ehEN6xBbhslA3nd2k+whE+Y/6z7PH+MVR3Y3G1xL8G0xyuUfQlh01WlTwX5g7o48C07XKTX+AHHH
6FU6U1pOQNq6KNO2KHtqPH7EsDX+MuFI7kd53ZryT1myr11/qz2X1fG23TRAOdCgu0EwE4/9kr6U
63FRPkZ2UUl0jKAL6gjsab29/KSSv+WE8ecLOkpQBb5EAatHOlESDQacZgBUcpsZalNvhXUCYoFy
ytxWpEUMXP9dWYWBRRpjHQmc3Q1BSp4RUMIxH+fOt25Migo6za00AISuaUdpIxscOboat3kByXyr
53dUiDrvLFtc+vOmUo8Z+FiK9BCPNsae0so8jMV8rfBXB8ahjU1BEWtent0j8FHphwi0j8NN/Ey8
gACAeK+5IHskZzo9QYsdbnlHAzsIJIuqw3Y0+ST5VA5yfhjjdzBRJzzumsfifhDYlO04Xxanxvhm
adIOv3ka5fvggzqynzBeGc7ZQW763L8djHksEczkf2NhOgamQhpXK+Qa3wykWgQZ0EBm+ICJ1nny
f2u3X2VI2ub355gWY4rbi5OHwahSv0SFoN7jXKX+Ks9Dtbd18Kjh8syHcVvRKa1mINrH3MYRWmV5
LDacVMVqBAndS2IgYDYX5CDwVRM7wkuNOuJhXwQzKEkBgs/NHYT2r/pMOlbrPsqwFjEQsQK3oGRV
WUsC9Lj/rbT3ePrgyP4hOWcuH5CoQIeA0vDs1UbeAgoBIut8LNb5T8MhO0cX9dJH/7pc99wCSIS3
yb9/h7vZ9uhtsF0DiPlBxHvMtoEcX3tl5YAwloVD2vpuxz6PcQfiA7+3+tVjLajeqBEVDu+W42z7
Lh6fmhl3ZVrslRWojcp/JHj0B19TpFPpCjqlQFoCwLnpuNeEf+HVhehFvifZ0/vmliFjR6LIbBbF
cAiaQWGzpadadLK1crydHtvkc3XzBYAU8UuNYHn3JnvCJcUhOHBA8QDmt/Rv9I7rFuDyUnXbu3IY
4GMQMXvJGLDnjmjLSnfdwwJAtjgoOaa2F7XH6SZMP/Ae9Iu8boHxu8RUKuvUoO8IQFXJL1aZenQj
B2y8T61Zag2wKIijcODIahmphTO8o7MII2PjgEtdzTFTeRmd0BXP2lhcfRF8b1eSd5SJEdL2bXNJ
ie7+EwLkaCf+LjDSlxO+QzYEd9VYia7LsEpIpHu91HbSAVpBoHZ+VIxKseLM+OLnJ5ScDxC5nWAu
CPekglz0OrYeI4LDlehT/VhYsnqFfSF0dwNio0rpE4agsc89mdyuylfRqkqMnXbANzgecAtIzaOR
z/CtAJig3aCX9ngsyi65fjxw9qkFXOJOeCaR7RjiuiqRCxM8sPf2YV4ZTqzN4MYDNSnwMPLFrns/
zDC3Ik1m7zVsoaih8pa9igf7r9wciiaFpGjoEGLNkjkQDPhkcUegKNVfGOTZErQ71MP8r1VEOPLv
rNHnf8LyfzES148tTN36rOxjWLNm3wTRxDt6VihcZm7e0zCLiDqS6/RQobWN//bIHd6nffuo8VVb
+hF5Q4TNc2vR5XiGOshG9P0dqT5geHjYjcODolJCSCmXhZ2dZSgcWUYtPcARoPP2SOi4HTaYhXx8
iKD4Ez58hBSV3kFwTqOy572JvCM9bP3+BWAs94xOOZz/edUkDLL/W2wcR8AuzIRJDsdMYNK3eluS
KzIPCXjCYNvqyp/krpn8UgIwFcM7r63ox7Zj4kskR2cLgqWihwKMxyaqSfLf65Y5imTwTvJs6Cx5
Qu+N6bIMaKgcuDH4iXvf5HHavdqje6lqjxuAaYf90lnOkT+PaLwXIjrXVbJpgZ99ZA8iTalDkrJF
rXr3odV2zYuuD/JeBn8VeYqIKyXltBOAU/q69ligMKboDbOjkcRwWZIQk/EQKGDJrdMgC4Ig1jA+
8xNBKX1Yod9K//CQrxZY8cCGd+xTJUnR3ZqCd3cFhmTfrp/xNh8nEqmY1OfS3GObvzhUi8wMn/BC
hPjhocDkyLfVM9cPgnbM0pa3SZ90G/mujTX+fEWsf88cfO2mBnf7AIdk6Rg8EN9heqDWpIwyvS/q
si5e5xU5tFirFCE2K7dSAiTqs6ujQXPxZjWh4EWJO9L4GJ+l4ryqIWAIXHXri0L7L37/pe44OFIj
urX4GAxFkoDQ5pNQnjudLX3SgbZkcbp69DIqSUiLGeUJJU1jS7MBNEEWWF6P/Apar72+VdYuhbkJ
xCaBhjFnZ9LZH83aw36PO8+KbKd1PWj9lwmyj2BtQO3R7i1S00OZ0ev844QIXeuOVsci9WxmktAF
7LyYpwOYJHLTs64odYz0tKCymKkTf2BV4dBaVCSpMfbwXB6MCHPk3oyADdVqlwcdHp1pQCno5jLY
Nre4JLowvg70PWYDYwSWEhxO8cdd26IpGH0hoGhVUwtlIuewJ9bQzwMvuG9KYqHZ/6P5r7+wTCmf
eshvcA0opHjOTSqvIGCKjWBnq0NVchPuTncVL1xNy6xf8bqvFuwtlkJUs3GPEBBAjWs+4nvXj2Cx
3FLmrFMKU1IpEAomD6b2Rca84613UDzlB1EjDJ6r4qKV8I34G9K2eQVakp+PJyleksRDRCbE3kkP
qB1juO0ro0isaquYiKIZf9+rCLC7Cx4zu+N6UNaXKfMGnF6/fTe8J1IGhJZU2GgBu+KA7ioJDJjo
bE9H+wOv45W69ydM73b7EeUQhhcowSs9cOoNG2ln5ECgrgiltPc4utsMttSReb7/OZgePafUgtEB
7O5VlKp/OVIecqeA24txM+Bbtqif+th8wn+G3OFIJHjZ3bJPcGVTEfG5jOMA35sSaOR9auSkewCz
QbHIuXW5PemUBj/0k7nkJKaL/s+zRGp/lgnDXzmc4YB4VByABoCrOqAt/VfBJia3fs1ZynBkDVa5
qZteyFbaumf8t/bZ1olZtkamTQfUQjPpKv6NJ9IjAZdO17yVPLdWtUik+0UzNVAqW2thBfaSG17n
jzVZTA02fdxxNihyTQw6CgT/aEXgixlkZ4l60XsxqPy3b3cjr4FM6OGBjOVU8noSXTGoL8M10lcV
d/7cVUliWpN/BLF7neueMZFKJe3UDveU0bA/vpbK/Mls+5M7b7gFM9X/P/V0a+tuBGJHSuezne2w
ULOVhPn5qErv/cp6KDIWtb7Q2buPBUj8t8Op3XZ0xlEHoBDk9gxfxs2EfD9vQd5MsNXbfe8zqpSj
oVhpEak3LiRKQWmqwg51ynOh8ch6X93h8KH69rGQxmwfOMo7AzATpiakynU20cE193OpXweNjnge
jqt5X8QCcFR/8JXDz0u3UrsAGANRFt4h3G7rtBVIphxWQKRETitegUaZ8ac7bSkX7A3/orwt3Xo6
U7gyniOw3WNiNlLsMLO71UGSpNWoKnmqBDv6DpXX+5i8wXVp72cMU2jAvIF8tRWYQl7aKzz5jnxM
v+Vk1/QF4W8Vs08K7dodPGix52RQye8ghT0ic55NupHZ9WsQqgmlpXeH+ydsDGO0X05nZbebLrg2
0aNMYr/NFJWTgMRpnlQzHOqcPlaftrnMg1gDgL/B8YWLaPAuvJK1udyENbB5AF/Mt7XX+k/rTEQn
NBdi3ixdwNuiYCAuIletSKX7ftmITa94TS0AOLO83K3karJylDEW0qFSfxX0gtqW8sMMbqFkWJbw
KhFWjILo7+kyETxzc7QfWOTzbC0ZvbPw57WmSUZiRPDxkyQe3ZmdC1+Ruidal9Y7QbmNYMOLsA+u
U3zT0/8OsIt2IkqI6TunUOE9/Sr5vCcp4QwlXqAeRZA+M8VSi+4gSZPJxj7wRztzU3APOoOcjV8W
4DwYwssybGEvuJDP6rU0buVYI9aDvKaGD2dpQKiovIsluNOptaMQUA4ezu4bYkpP5PFivai4v24A
A2DkA7G46J6OrrqFFK5//ZGFmh6K+Gjp06Pz7UMxWFANOFVJquROXO5s6EfMdKTKr+DBIwy5tvJp
JDHcVMvq0pkf+CjPiSFimn95xOTouTmJA9ykgcOAfEB71od5SSPGB3d2pVYHA3CzJfxs3oAzeqYH
jy8aSW3muL4yoJWXQA90CjoyTlIAYjGZQmHblTT+UN96q5bJ9hrXIP/AbZw7qd4njF9PO/h8Q2Hv
arEY0VaPUJxILBK03ki9CUonfCE5GXunea2TTAtOpR4/nYXzcCO75rFNiWx9ba24hEP66nbJAawz
j5njaRh4khAmuDxs1WqMQUTk7Fl5IyvkRIKkXZVEQmdu4yK37w3FWPjATCiw7jGqSHhQLIQyjEgQ
n8FykyQDG605JJ58sj3qenk/8M7MzjYWjtti/dUh7bPTbS9+UDCsOhJ3xmBsYmRH+htoIwjsZQPB
v3JF9g1INU2hIOx+BPq+Xz3irYNCELlJbgvHZYt0OYuz+VicK6VohEV9rX1N2CZhk36E2RvQ/ev1
llG5CAGK4B08ix8jh5zcJ/dWVaTYV0bQ7z1NOU4yuQCHRgPGaMK6K/obSwMHgacnXjtZOP78hv1a
BHcHSW2RuG13GjdoapCZOMpGGKdKM50Mqrc9liN2yRjlRiW4Bb7uLB4cactBR/3y2BaiYkBCA4XY
QJWsdgTcILZgsC7PNPWMFjN3gTmK+OXj15btSBiUJtpZvrHxgrvzmmdUFF2NiVBcoZHxxqQb6yk9
pw09FXmzGIjRsuhr0UlPrQkqYZK7AH+oaQEhb04J/AQPNKr3gDP/ghEjZ/hHdPNM1ZP1HakxzvC5
sehO79YcUSDCcwHMlajIyuWPQmhpEYW14MiXttwzUcjTOvZn98W2oY9i4Hy340cHGOD7vquwU+7v
SrkYMAdni0VcGG9q79fKWRBbeLjqjHvn4S+JBjNeoZYb63G5bDT6VNFsF2Ge1Vkhddk1N91P6E+f
8iElLRtQA8n/WUpRVPjpo1Nivy6qdcCX+2BzD8J3vOewWIjQiZSG3B+IKtE5cPaA/kfYmreXercI
VNyOpRTtU+AhhN8eCOJjKG65P+QDr9C2L0jHOL+reF/J0M+3yRVzoU46TGJCkMJ6fXH7zbEBwuiw
mKKo1j3Qag7jb8Do8CutTtS0wDEfMwd8pzRVgc4ltkemcbNkUP28sk554ulRv3Ki1DMr8ZYne/Wq
OyhXzm/SKcZGFtCo5zZ0R4C0YIwysyd7fAmLEQ4eok+RHCKk3BlDQLwCWbsFH3eG2jYvLacvkcmy
Y/4C7diaZv5/KNu0C9zqFroNtqE2SMqRLmdH332C250jTzMnrcFl1htkij2ZBT+MoGJej3z4usO0
DsCpGtKtt4CXeRhxJfOe3pQdxK3HgPGY9I1g/+7ywo5I2LLv21cSzoaggvZurxElHyzuf0d/74eA
hTWKiI3wM9RI25tPAi95JT2Ochn69MLnOy4oyss/CEgWBPLPc9snowmyEQ9y+1duvUHqDcQsn64o
kd4ZxdQ4MZc6qMqnQmERXL694eNhplmAIKEinrwX7qx8W81nidkxDCnCjCyPtr07N0tCp7jiJrOd
cD6+0c+BlEtuNMe4GwVGYXlJofjLd3WN3PSt7oY0qqkjQnnAElTbkuhmm4arAgK07/2pVoW+8DMb
Qe4cbcT6XmXPnSq5vcZNdfODMGxLVAa0p44vbWgbiuQkHt9J3kYJ9CWIOJbXcRStsDWTVEW9XgwY
pW71JW1roh5BEzQa1ThVOlpWBG4ds4M3O8guWrX1+m2AvarY3jxNoHjk+uhLLPULKGT6sBtwjM9I
L6bVGJS/CW/POeWK5QhV2g4rEQPnVkJFNNgfUKTfRL6e0KPJ8VWyzD+IVNQLNvuydRsaITbZiWJ8
CCLMK/4KeRo4HaofWMDgH+k0itjLWrLGXpsn2LvkEwcPLrdnNolrWZNvi2sEiN/0LJWcjYxEyH48
pEXFKXNO9R6UNpsARoJUliPMbx9W0lUwBdYKUI4baDFaH1zuFn0rSxizQisPkGJv0VeNIeWNc93V
yBsw3HD4xQxvbaf5jBeg7gBBqYyrPoMVWa6Z5T+8xMXR+G/mKh7K1zgHMYBYUSrjvATtvUxOC1+n
4UaeuoZl2KAtOS9jbTh5NX6OUbw/wzS5YInggp4ILLTsLnckCzME6WmJ46lfc79LjcVumA6uPs56
vOWmFAXUEHlDUrjcAXvpP4z6qzsbr3+QhXeXh6oKuFj+3M7ZQDKfOk0RJhJA8PK6Ac8IhsfGLarO
gMZ4xwIH7/43IJeOD+iHvu7uTCfq6z1vLlNmCAdJGiTysXXg/1uSS/NllRDITV4CZK3tQoY9yaFE
W4mFtVlChZ8tW+do5Pd9IG87SwuAZQa58lLdEjE5/+xfGYzpXLBCV118ZNdIu/eUOw7dgJTo1Oxj
H+c/6zeupoGdmXMcGCsm887rm9/ZWjyVvRNwiI4QdT0fLP3wV50J/ZZWoFlZU64AEIN++CPsxS/Y
lxhtEGZcm7W4iaaBch68qSsqAQf+28rVEwyOH/TGwr6iIleIp2CqtEseOw/0FG3UC01YX7t5wSbQ
kBoNxq7RaCyx4yXdQYDMvlgFjiiF/8VU3JOBRV/XUnjEDOIa7R23yraeZx/TcQfeASJSSFdJd6qM
5/+mdJZ9LMPw8fhxFKh2BmDrY43UgR8RkCuYYdtAUnocz9D61p6w07nj+oPZ6Td6WdR//Htab4zT
ThJ2QeDH489TlyeN6rpvEvJFTUnAGZtergwN1p3FeVYmYz4MCG7pQ7T6UR/vU3UZ/wjBlwG9w6Zx
OOntLb48FisAB9VnUAnAB9QudlRLuX4c69I8tvdgGDPB4D+R1PnkcmPIu8bvLk959NrdJhcG8zTY
/zg6rC/gyVwcA8AUOriNtyFJsg2zBHGByGog2tBZFMmPTCyYCuFvPCZdb6D1tlfJcTaZfaJiUp+g
qXnUVgRaQqoezXEYk9rhCNQOyyCBIltMm+m4BG7pQtzjDVr2ln52oblIkU/axTRHt27Cw/bMukNb
Vd+sLe4HSp61/q+BDHrKpY9DuqcdCQqIGCC8YZ1pCDn7rXCj4j/5TXkqu69rQi4p1Tq+4cTjgftO
XmVRJilPvC7tlWlgLypK0SuJbCftis0FIZ+A3PgCc4nYG35nI1g/Ly+Rgm+AST2PP5LY2u2Md7r9
gZQOG4cDw9lV0KNaabKJ/F/drwZPAQRxV3NUMFUNaAwoINYbrzsLh1Endqp79Zgws9NvahgyJ/6S
gdAwjiy0VfH7tO6+6jMGw9jfMGvjqKKe04I7bQ4uDLXSC2gGbID6MV/sUGrFe3Iq0h4YkdJaaWtN
eqaZwQExHNbOgPlq3GrC+oXfGAthQEvTl1qTgmTNcz5Ctc/IwC5idOlHrO89jBIEy2BHJbkQUhaq
CMubwZTlET/SWqI6n5vvQAn9lDqbrDPQpQAremWaAjoVmywO98o8h3uP8Rbqbaq2vY7nhJZgHAst
/ohPFfjLTZrQjatb1vgR94SyDfSnnnt16/4YvhkYMSnbeRJaasTn3u+vBeYOKZ6kLhqtD8WX/ciA
qX/d5m4foEajXKljsM2EahNzDuCsUlTlj6vgrof/F7e6ACLzxKBLHVrJ1dCD0aDOjcFq3flb/ENY
DuuM1FchXFYLWRw395nyHiUTvZZdDLK+CwpkWRXcwwUZZM1YJA0Q5qEnIDN1U/s3AOvuo4Kb+/Zm
doijpboWvv1yv0luDiKLtGNyEsgYL04t9iptH60YhaJwFGIyxvTRxmuixm2frB6YzVTZOXzHpbAj
3cD094YArwqlH3/g1H0eJ/B1MRhYDnzSUVJvvgfYh2PWQK6Lp7dqLIGbZ1MJee4oE24ZGsuhqjFB
BW9LI8dDR0BetMRW798fe0UKsI85iAantcqgfh0JW/w4lxP1PetZWUJNzD60X6dJGlJXZMXeUNGL
3QsnlgaTzOYWtErTcBaBWNA0ZNR7qTJGaHAstbw8qgAl3PBz7mLH7kei+h0mSFRSzjt9SZ2RYSRn
6thRxo2eK5H1HZfPdKFu2HikdiLZ5iBrSani8U3eEwasuRoGdPUIVstv/Ke1tbgY4e0cxSRCbRbh
HqYwDcHTloK79xcpJZ7H9mXmJMwfBQtLscNRokWEbYbM8S7P5GCUJhP2Nm4Ab4Bi2U/V0hWkDVsJ
nZ7eM/22LIABHZK0CqvPWiYcf8hdk3kyyS8Zwo1Gv2M/TGA/koGyjBXyDQ6zSXSxA7DmNjNx84Ar
8Qcu7jNbRAsm4w8HtLReXotG2lI/chuE3bQxfAJNNgWNlurtkeP7xRAYX6HrvLT2D6WNcbSvW4Sh
2cUJl1zIWfBHrpcJurPGNJjOg02a7MrrI2Va60G7TMltKB9HOi7HRGCSY2sBVPYxFp3ELPorulFF
VmlONDXLn2JAEUFirPeOQV0udTg2dzfp+7Hh1/4i1PSz0lxS2U/nEY9H+qA+49YRrFDlOup3semR
sXy5bfqOC2LzeX9zmXfvzXJYKBcxExuQlzDLy1xHdL2u42OVTS6mtU4qa5GQGYrLJPsFF191Mxqw
bgElrErvu6dh54ntwEVKhJGfE82khCWMJCZsPcNrQU+VNZfMIW0J6n2vO7bNJpb2zGoxQBBtD4Kp
Jk7QTVd0gL48BumQecnl0R6zcUhKR/MpXoxBm6HtEj1BwopiBpwKuNa4BgDiIKYao2ahIAvIzoy0
Y5VZU2T4K7MEhMcspkHbd4/oilP0QksOxWy1dEFrgTqjutmuqj7U2uSwbCpUy9DMIXjfOrR6FkbT
+H/5Hc4hTCQAH8+IGIPyCSAdw2IFFeDdN+3qB/WM5zChR3JWXez9P/Uzcm6gsaBH4nQmrdKmQZdd
HUOUolJYOMWg2XD/3UoyBJV0BopZQMRsgRscjh5IpyWY5fvor1IDMhopzBARtgWuNzAZ/L9MfrL7
9BzwH4AlXQZKFhBxaELLoMflDO+K4xaFuT+aBPHjUrvM1KenelLX3jJLIZGauyR4d903t9R5sJbU
awtZhqbh36OLq4KQpdKnM1efII4gF3sg0MGVbsNL1JXRmZUoViHe015BNkIEQupk27tRdhKpqs2t
hq1y0HyGbxwFbJ1NlG/QDZJ/acWuUCfinksv3eDHsm5lE6Mzzup2CDOMcc9bVC1jbMZdkOsb5MSH
ng2YC/EvXOXqvKy+Z3llbrEXxpxrsMJ28nijaqq6z1dtecEI9PggbvnCEEuCufITbf0IZUks/dxz
LuLqALBwmFK8LMm/78WLt+Wu9oWOl96rDY37U29Ui8KzusYY1PG0JF6pyyrNNeQV2eZ2wUQ/9PVt
W/peqM9623GbgBt5Ed8qvqXj9WHvyGeQ04vR0MPjQmXxUhqyEsbgA/ijzAu5Ykw7wL9LvhFBRYu8
aaCNYJ39xuAC5z/d2D/L3gMNraj3PRd4miyuAbqZVETywnFW+ze5bcoeILmaj4qkrNy6A9j5G1zm
y//Xz+J4MAdtmPs+RWIsTwJ3zecHFUx4M8XB/VRdlJ5PU7pSHJUASmmtk+nbojnkK9T170joeohI
Cj8ThCzvHDbvXrjAM9tAg8a4WcwDaNEOM6ktENRIpdcU+9HUyKkDDCQkiDWSk1XVM0wOSLx6pBQP
QQy3/FoI565cUyjihHkElBc55QyE2Xg0UPHz8rtVe/dgswcz2swPrY6cNMsUG0FtTH0WjowJ0/UO
cfI4HY5A9Ap3kZ7rgbHiydOGeGihdwqqAEMnS6r0BS2VvuTjwSNZZUCqwb5j0O/ociZXYeyENAf/
z5uk2Flw6HhNNbqvt0cqJHaE1zeG7Fs/B2BHO9gSDc2BQDfwMpiNPUPYgQ62jWZcyQUKTBKeVSNq
O1KoHfeJZr275vRZ7myKI34FGNnZU+FiDARxF6ov5z9X9N//wle+YgUWeQLzX9uIWoJFalraEAzW
8QPm+gczNXalvpIGMbnUig7Ut7STkvoeebsDlj3VUneEaC7U97yxeWB0DDG618pVs9sxMN1Ta9PJ
D9h6keh8J1UNm5uD3+oWpzta6pRuW7fetis9xtVecLPPgZr4/bpc+O9y5nzev+JffXQ7d2083pNu
4nNOa6xVP+901bu+gGO/GyrLoa+nmWpk6kqHHvVx/00IA0zLr1w4LgAVeKwAbmHpuMAF2vGMAz85
t8pJxRlEP6ZZWA4iYLZeU04tNydOwMbd4qm+Pa3RXHh6HMfKvPgASFvYiI1jzwirvin6JCqbBKTc
SQfLck9iSm1J8/bVSb0O13WIgJ/wj6bPntBq10cQKvgDR6KE8k36NXnM0D/V7RAd+dxnusibonOn
rzUdtpsaeQkc7fvPDbfXjBTlV9WzbYQNOgcs1cX6Gz/1qY1OeUyAgV0w7odm7slKbI5I8fTYIQcI
z4i40STd6ztvo1qmAGQHsc9ZsPmHtT3SIxV7faklWq4SlcKhXtnOo1K2+Gvkt1yLPM0PFmr4Akar
D8K/w9zP8kNdpjqXzyDqOWu8y+/WJI5ldgbr22u3BeKyNUlRyHlPDTRetgDHSwNwaEDGHAyEbiyA
szS2qtkezmix5Hx2rKFz8UdFsIMv6hFaJbVTRxt1p1coU/Bn00MdaWL08IuHnGRWsbPzcU5MZsmA
gdUnES/KCdq0+j5n2k6ml5o/QJEXXDzLU6LloVhR71mOocNCNBw+vp/vmhi6fIN4JyevNponTrcQ
KKzD5HO4m7esY1U1tAr7Fe4ih4r3LhwAC3Epzt11KN63CQBqW5zRcmE2+L5dwKMJtGpkY60uNNVq
BM6bR/JRtcYCsOqJfLXKNJzFDjOS+LvoLDp6AwZnfXXOdGMo3C0XMFGrrx7TDFQ1VaWrV9Qp73+E
SKs0/tNyA4wKrPUTfn5B74B/Ekhjez6mJHhxxJG4H76hWYFqNdTgFYUjd7ousILYv4wY8ApNTWFV
AZSQOhXvQEBobGkDjCVKpqZnd2KdbjZYHH+Ire252hcwIY+Lrty2PPm7s9PdSLZQ92HY4ERhG5Rl
mBBdjYshGFIRHlH84eleojwhAgGK2EGPUfK/DD5HdBj68GmHy3n9W2mfroitRn4KbhkT8zApY8Kk
JIBa2xk5sf91k/ub+KNqLKJtUgNtlWUxol0snO1sEK4Z8bYrGr8QBN3GlAaCcf0xTcr/7lvxEScW
yzPQRnVjzv5YLrQoXyAiBP57bLe+/7y7+X4/dwY1fI75tcmO1KJOO5pH1d5FTtFtNAMBVCT9nDoh
swo0YKckQVWCckY0h0vukMgbe9H8Rq30oHwu1l7vHQBtGDE3ZyhB7lRwNJeEbC3qRaFVX/yCB5Kt
G1YNkWlM4VAYX+ExC2ZBE6+zkignmP7/yDo0ijZjVGqNU+yBG0kzTGe+qamVrZt+oAiX6Vz96hWH
JQi2Y5Zp1FJcVVVL27nKg5kKcTrMMx7rTF/hiO8Vqj/kmEE7P1FYcfCLRwXsVGijfnzbAyieffur
SLWoSwy1G6nsBO4Hsmcz7DvSJ7svx0MfsBIQGY22NKObDoc+J0XideIOIFVLe7Zoj37KS6P6uPUh
mauTFy5KS6WcTl2qsaxDc65SrifKd5bAcEYlVvy7C+ZFZKD0Zj6PizeEckyt0Lckg4WguQBLcgfr
McJ1wYTCyQtY9x3uqJS/tHWNZPULP/aDZ50e8+cOdM2di1HaDWw6c8kHxNxC5rIqcREYVaNzwqr3
Q4Deiwfmr60fDkLBgeEqyqVnu0RgPdsiY4hXizSlkr5UPCEwnjlX+Z9a8cfHyvDzBfpC6nLMJSEz
Twm6vYZJ0O3j+/QPDkuSoucgzgWK2UZemVAgOE9VapG9FBc4aTPYPU7evUQB2OVC5n6+9Ykyzw11
Wpk3ZbvM6rfUTWY1ylq/fU7P0pKROeRNSIp5NAuw5+HIZr6XmyJ3QJdGiUfx5gY6seiVwhQTRWQw
pJj/DFXPLGqoOOnBqImjKCIszKsnANuctxhd17br61HveEOtoGPgdWDNdMDtLvcODcbAPpf1UQnd
fnInYkQ1OQlIb/JT6GbfBtAehPPR15mQPqXHxg/LqOog63JF7XNN2eONXT8ZcIwXW69PMjffIk9M
olr4fwVqmuRPp+IjCl3YYKrmZ3QXxUPlwqKz1t+xFQOzQ5iXwv6yi0Ic93HJNdCRGG+U4GxRVBr0
s1RFV19ztdFqCBxWdruDIbs7+MTPGb+xl4Z3bsjws7UOeWJqsM2K3kPkYV5UvXTgpyh/vtHi7W85
xBxzBlTcQNq2tU1gfuiYpRuDOYSwpuk8Not6RZg2hS78KS/2cJaz15rIRFOzS6CZmS8aEghcKm+P
txEMKbPyEwWw/plzc3IseLHQI/voMGKLP1UOcQjbQ+7/mtWKbQIcHRCSNsuFHnoNx5y/M+jRR78t
9ZUzjJvLRsvRTRL2hgPgWfFrp5qq4s8IA4MuJ4Fwh3BiCaurYyksP56FNlW+h5EHJeFcnMvIVj+9
4iRbiHh+e83RC4hDTgmpE5NODdWWuqgr9mFJuonzeW4NYt1FxZ1vJwO0O5vZqKU6AigD7HatJCYL
jh/SuUYQzYr82ijraBKcoDNgMkyo7DhUM5XTP5Lj4ccgPLyw2ftLSfj9dY+3bhGKN7vHmxvMIreN
bXkM8SYn1iD7y0IYTWKvJQ3wobTQimNCmwLGV0lcRnVauIwEcZvaBdmvwJsjcrxuocU0F5PPXtwf
KRxXBy8t1FXp1O7AgHQazT1Nvg14gkdIvRdyOfyFeWFtGpVBeBilrFdlw7KFlUau3YsQP6DyD91l
OxsPOWfwqWxzzOC9NkzDJEkyYPdbWd1QkX/fRAxZSLrsHYxwxpUWyNYddN/SH2CTFCZQ4YCZoplp
IYmbcPFJsB/fq1j10vyl6jNLkT1gMdjkkur3OjmVNvHVL0eWBUvAF/H0D0PcbNtwSrBOJQ+tvivy
bSspfYv6Xf+1WtPyIyl8q1ooKaT+gP6TnCzIRCtOfBusm0RXsNTUXLe5daqS9/6rsgqQZlykPUV+
zpLhzJYo9WfP17ETx0jUaNx+uiR9KqhylGmUB1PEDZn+B5eeju8lBr6eWp1kzB4+c//+IgN4B9aC
mev9cNY/NuCKV0iFr7kxofdW8oLkOUKjIFD1zAcW+3uNqNt6C2kA1hYKcKFZZU5Oy75eppbu/OFO
5CCa3/f/I/OUUB51XfYTyN+N5czqNHqmrFbiyoLrTsAr8jHYg2dbrFlsHhGhxsqhVEcHq0IOMZGk
EpEC+WPHbt5eb1htgVDw54OacMVI9ubqw0+rdlB9EVHHWwK9rK1zJAnJ9ONrxF7QV/H56tvaf27Q
WlTWHj3nms/D/R3MHD9lgzHr8Hc0p5y+QIqnxNOyLjuKpk0Lm6NMYgrJVadiLA5jEiaAcg7K3wRd
4uGyYy6CGjZwRKD9zJBLg/z0ITSApjiw4kpI6xwj88m3snibMMqZCSHIbvye2nwqLhrLQ08R6Pxt
btDuygVdRIcaNjKm7cnuBeJXlD/mEZ1IzVI0WNOwXawoQrGiX2E3IATiswrcupPDTy/xJlbB7HCG
0ehtnhEl1KzGnCm6FktGZxn78rbHa8HiUk9R2JyWxk0vFqpMjLsVE0O9jN5ryoY41eLPQzSrY3CH
8Bx5E7GWFUzm5xqkm1aSDKg0x+32Zp73PAsUvODUd4drm2MRkkl84hz1ZSdW/RbEG+VSrax03Txw
7wg60CeB2mbYmqD9Syi2qBCoNz2IZg8jCjUAUTXggWhWx2nCnqCFYQO/UXNyks0pRJYPdXKr3Hoh
cglFEiZo2td70DLtjrDLZkjUMSjIQKwoA2KdCxkpXTZ0YOzhy41sPVequfyN1O4xRiBupax3fa8p
EQ3AgG191ZatOtbVy0z8ExXridAkZhR6aJvHLwWRhFcngcRBWHj24mVbeoo3O1zdbFwJUl/8FfHs
KzlQ+ezlat+pDyC8CtsW3+8uwzcy09hl8tuXK51R8GBttGs+v1APQhqIFcjMEma6OtbBGGZAgcwk
CqhtRuhpHrOizT9+x3PqR+GtJ1MISeWC6xn4PrA2D1cxxcnZ4FUwv+dgQejAcE5+nh+yWiF/HcZj
5LAsGo6JaLeVtcfNiH/FtgbBDXrn48Dy/8OWWp2njfrBwkgALDR0XcU2Gi7bc57710oYm5hc2Pe0
sW0to1JPpYc93pV1zj9iCU7WI481WdWqgGaDhcvwFf/4YgSsekwCiIIwNDnv6mN1fiSBqs0KwJOq
85Dpm0iJpXIe6jyVlxxajMeMqG5r/JLoiDX6dl8Pey2ZBCmiFxvLbC02KocQAX0N1hv4zoQBuFpr
nfyTQXVrukm5aZt5uvc1ua5wbmcXOVpnVuyePZ2/HnKSHc4nP/HOrF7J8ZJLCD3kyTLzkOv2wlsR
X5E3YEug0Cw0ypyfheknR+/cy5wY8BCOcISd8VzC18RIgOWRtiyi15/G80fqTsHu50eAPY2ehH7i
ge9VxXBULX8fB01v4CzTcAg5zh56yIImAj6RwnP1Lqsm5mgSXnpBDKf7LRwUbGBlbZ63f8S/0ZhO
kbbniiSBCmxI6uyzFJMPp0jo7w9+SVUGicdmpeK+HZg7e9p13sxh1duaghQoTOy9ssS4DqAiE07e
Zlp/pcTJAfXxiFsOc9/t5xkJrRA4GwPnEtxoJnYWfTwC+cxmuPJKntE+xavO0YaVTztVA1ykniwF
WsMN65ifuRXR2HXnzaOEr9IDfGIRWqXbMYENDhvXNb95Up82u8A45Q05Ut4rML3ScD78+Wr83m5B
TYIFkZt/ApQzvrgbMS8/xATDhHnR2hpgs6b0OUXyIctol7xe4x4wGxWJFwS7CaqooSgNbgzQPYkf
jOIpVRT22rI1PPsyAPOYVOXzscfVNk8Te0GoEiIGoFuAw17MY0ngzGFLgfioplcQ0vVqQ5UYY7BX
NjMVDopZsGbYRE3SbxApCJa7cquUZL6QQYX/NIqyH6Nhw5BPbfNgcglPkBNIpuLPdheCDsKyr2DY
fIEinRsRTo91oKTgP1Ojd6ZIWfTN/2pRIotxZYCVqSvosyV3l+tUFnybuQABPKjSasq1Y6eQCCue
ZuNylLWZt4ZVnTTOpWHImZT/tIpiR5katBoSi707LZ2dQqSTdf6eESnSL1MkWItopBpE5l3g88Jy
1E/J60fPFFnfHRHZt56bUyVG3KK9pjzNZRtFeJTmIZty1x/Ym64lQvxzpX4J7szRGAy1G6c+6W5T
jwFAFSchhkS+UUZ3b8qAHVR18PQYVEfq5IPjYuSPTu1Yb1TqnPuEiuz1xir9eLfl5O5OBqLZ9vl8
lqp3PT46J4WM/QAww5snqiCEw7RTwDi79FmtIpS5qSb/1/fQANz+KcDOwyKqHyFYd8WE/cAQTmb6
g9liB8PXpY+YP1VAJoQMx431YE5eSgvWoVqQatiifvC/+uT3t9ZpETM7x6EABVaLS0Zz6AH6IMyG
B8w02w/5rjuenv5JlHiE8VTHUU04T8WHx8xSSjvXe7QOPbNbRqcS6dLJ/ajzFOAl2Jy2hm47oYnf
3yfUr+EMKOBXdFeBjigaYMDQ75fvoPM2SANxREGK2AB5pTcBIhp7hZONORcIeSAvVJu24TK3w4oK
V8igJe+sKdpGegfHzHWbF/uinMJT1J1/NOf9heqQys1nDtp+uI6ZG6KYlsvPQ2E491FZt580Sdri
LcIVrarrlL0tYEbVaoD11RjCcQt+218eWZthTGdF3By3HZV99ucbkDQDv0dk9ToDVTQRHubZQATL
5Og/C/5QDUP2ZTpgnec0sRq3czzqbfG3OeKa4ygyZ4q9ej/XHk9+Oi49n/fq3cD3gHWZzMM1q/ny
mEXPpcrGLmmkS8dlvisd+aUWXXPI/MWu1RVrEU8uiEFC1bjb5QKG+GD2n+PlmrspCL3gcYMyVdKM
ZPjIqH3C+z9kKZbk0Bf7IobSooNdYlHbNx1+pAdN0S2YX2I6UJxtSQ2cGB7O0wKAo98ukZtJ1qr9
IuSJGOAyMuza/k7k+R2g6e+VDHCRNXccF5sLx0ssoVj1l14BFnXIyK3aDLxoHMeIRl+7SoGbAtbX
ari4CwEmTSmCfvL3s3RtzP523P0xhXnwgDdn0Co01NP3rpVYDap8LyYnC0Q3HITuOFEJG045ohMh
oLBIOs90fhXmYgZ74BSS7HFsz2otdkjkKw8x+iMtGNuF6UPd7tr/SStbiKkom3wRAxJlmCJqB14W
MSRyjmr5qoM0stINgnsscqSObgqvT6fIdSfyTaDr3p9i262Thrtj6LF0AP+CsarrZ327jqQNvah+
hR1UlWiwXCKVngeWcme5qNIkyNc/ZIu4AbWR8CajoJea73P4mzk/kTswYFuS3pSycFVRHO4erQ0U
acdeY2RmjUavP1i3NAlpU1K2+RtFpJMcXkfwwCgVDdzvKxVo3sYPdOoiCtKKRo9BGxJHMgKhjMa3
PgNKavWtKMrNj3lpNI92FubVFhLKBTQBuKJvGmuTd4IUjfDsmYv8r59Awdh/HWSXmAyp6YXR34Rw
O7Z6FPk59csl62a712xqmmy2wAwFZEkumYdl9xpc+9AWUaxeLxJM2yQB4pBMCx+hQf3y79iQ94gR
trU9CP6DiV9j3N+QuYs9EkZHRzM80+bMVUvk0vFTy6cjWBANAlscd9VBex4Wow7d4p8hxL901X+9
Pa4XnhucIgNEg7blVUUq9w6ApuiDkJyK+L4yQNVTxL9vbx2g23dNH677lESQUSBiCpcL0ChI09iv
RfmKsYkb/GfQEDgCuNJHfjaglFExqSfdSuQqmxCHo4WwrbpIPTO5mQdd7TxOr591wmxCL9ZWymXm
CLcqLDnbLJD2B6xhXDy4CboedGBeJ2d9ZWDbFsJwjMYkioFXlFM7Hjp2SDNGCqY6dsw0pMmLJkl0
375ODg6sqO4qXeO7fA7QIdQYX/gYpB7uXuxSfd2+I9gBz3rQkDWQuo7j7gii9sC1nw7NNdsOClb+
BBWhz8YW/gyyLj7xODNBT1sVKELbkQa/ycczJhmg/D+iqpbcpzpqzZjDdTNePJYx1FRGK8IO0YrY
j0SWsiVpotGNcsq431g/unQQyEZk2RvfrjvOjJvcNqWderpuLyCN74GvXLvqEHupimSQ7MdyDzMM
a3UrS26TFutdf2kFjHgYUcIqpbR3B/0KT0BWER++mBTtSrkt8ov4ZFgfC+KAK3Ps8QgqZBU8OFS7
LJXJPks6wejxXOBvBsqC4txEz5VLCSVVYXdi3qLjP3j0j4TH0cQwDypyNhg7ZHWoKyXzm122hSv7
VavozJ8rYO2od1oVvMT4m2VJQy1vY9o9or6Fp7yvJqx4VwL40TDpBhO32wNwez/XfJkOTeST9Z/C
h03uKPvOlX1kWZR7+dyoDUy84RN1CK9+m/d7VO62mkHXIpQi4M2ovVMnLXKMoFGktmL2ZSmelTdo
yGorQ/pIWMLYJNwCfQtQSffXsxlPA3PXT9hzsuB14K5a6na8H+jr6c4+has3bcQSJdnj6sIGE6cy
z3co/bD9IuYXSpJvcY8W3kHN9mgo/hyBTit6XJr0d7FmjCBktcrrfKTaiBYwA6agp34IDFYOddZI
ugCGldFcjjCS5NZJb6euotvABjXoKhfnluPA2IxxZWH11b4nGMuR/EwOYp8Grkcy4y+yJ6xDv/Jh
jZDm28naEJfhDVqd5zV573k4fV3SZU8iYHXYcsfQ7EDisc/P/4l9ii5XYmk1Ug5uu/ZND6ttV1Q7
wSTp+U/8LKcKs1NjvoE1wQIgAnvheTA/fl/5SePtH8eiEV3Tqonvz7pOsxuRt+08zEudZIbv8Kay
K845tBxk2rU0AnbfM4/lnaQku7/efnAw5du6pZCt4ADWuv4pJhjgI9n8Vc/jaw/jUuDfnvmlOmCI
hgAXlKKEYDNr+s+1XskNi/yICdojaNrdggLe9CTIcnzXNHi0JPNg2WPP9DKPpnp+0Wu3eI25Fiuw
3F3vAv1mGw0LMW/ee22+2BFA6lNXmM0Xq+iDw61pj/A6iQVbAhX9a7tfRVKer0RkRUUZb8a4+sld
4IdDDc4Er2xn7/jNp4X2842iI8cGiaKvXlfc1auiPnQjkLLdJzlN8Fbed+JDLrDu40FTI7AVzQ6k
YV4ZEhR8Fj5fX3zM5VQqiOtrn6KumLacf9fYkW6WI9nvdHRK12cHvCErz2NZwsjcjStKn/s3su9F
Eq9y1RgWXGH6aKP95jIlt9FYVI4H3q1GbS7KVCbOh9WNHY8pm1BAL0NCFoSJ9bEBZT7EP5qkVmr6
4G31FVdGRjVko9utZ7Svx0qLBK3xW771B6LOvGebENj71XJo5ZZq6Yfe8uRTvpOfy2kQtRHVCAak
YPKVpv6QQ2jY5l37fCGnG8RC8coBDJ7re0tR2504GpM3g+t1LQQVsUQUtAQ02Fd9mOxkcYhWjhut
bSrmR1IXbxgLgjLTOmFUSiIA4s67TjTGp3QdSIEJqJPqri212/8L0h2aHAFb3EwDwGTWkeUuVRDB
DzyAN24WnRttiSZtzdj7EumGKhG0ZDexuJMWwtWB8szy6gIPyq4GLD304KHzbJbD6z1saacXt1+q
lnDffQ0Ia2/dwAr7SJf4QZ5yG7aZHRdU5VUAb3JU+CdxYkp+muhfEB2etuy49ACCci3lgaETKn5Z
WyaDIUsvLVMNRLvpKRTg75286zJtGlQNAGW8jjpGG/nTtbt+XD85qnxGkQYTtIWbmTe93arWNgC3
CuCBILHSqmM00A/uCqetVYO0BbQB2BDFFBWOpUwzjHt+H+liqccD5swXyzSTWiXKKnkrdik1+DSz
9gBMoBy6Fc5Qyp7+0vOdTEwzXoSg15HbuZYOf4iaaiJfjrENPhH8wUZdpIgtbuCUN0hqsAV7TnuY
dxUaaLzYcQUCQwgZLPv0SnnPLHlfjbnswcf0r7sqQS6HpJp1zxZDXPCCZ9xjrMh9drOjko1xBkL7
RCdB+xJfZJgWjzB2bVH2Uwvzos9VTLK2Ymtqw3uraCZiNPaCEynfbISzbwfUqm/zE/LTpBnKdl0t
lBEWs5l/kHboFDKBZdez8JOgM9ugUtlTrp65rjjwQ1vTjtw/SQ3LcKCYThI+nNSG7IxnZ/sZv6bV
csZ51t6+KI55p96D9E2RcaK5dexJkFo41Fhwurfh8qq/9HiC3E/NCoRS6Qz4gdHO45Aoo0aXwycQ
KhVbD/skTZIqf5ipI2vdk1TaRACDEAkX4itDdNMOwkjLNAxklf9090wzVG03kP7nLkK9rKaVLlTS
rkcvFPQx9ZK+XRaNLFhgs3xKDSjjz8fQejlbw+RXwj2z7W+QNdmp16z7UIxppkHhiDe+lESlBPd6
2oLh++2mVjv/MfW1lWrMIfflx5v2aQwHgzbjOijxrYg883YBBJdeOvixxIBG6Zn30o9kcLHMik1+
8CHUO23XKOFn7uDPA6L4OnYeqkTxYuBbEV2qY3f0QS2+JuunzmLF/WRQ26eLQ+shec+tbPyygT5A
Z2sf9rJNyojtTkJBXs/XIvWR61arFYkLippJZUf3Y9OlGUvg11ka0jJC+BEbHKJoVkeay45Juc4K
zK1Ca84K1o794QtYrjHa2IgkvsVc5oea2AFk9c2wX7XFEdAvcCKxvAfn334EUKHDAPf+/UnMugoD
E0O/Fm0y+y+ku8Iv2axeB/jdsVXoTiXjkaCdVyup3Lo8JBVFHUqzDRlWsvLx7Bpbb76lixGKWN9Q
9czA+qhH4hQPyLnJMfCqgG1Pt1DfipNIzs2sIOHDPO0C3G1pKI5SDSrisrjW9SyYOomKaMYQCaeV
3hHD+WtrcOQhYEFQQr0AQCpfannqbpyw4WbVfI5lNPYRPblUDiaAtFcWEBrCM+hw4AUNAys7wwVD
sVqMU7D3bxZVCyhisa0wShW+dV/tNsiwzHtjAK/iZTycwjqYG1wz2/lURXdMCTmUwi1EbO4KaitK
PpeX9KOnDeINK5Z92MTizFs91brtiz/TJRbMiu8yrVZX3itcwJjwD9ruBkG/+B610GxbpRPWnqdD
JTl1nH4yG26AVcLpUB11EwsM1LUTJBOTb/lLjKIn3AnMxsFpg7yjGEces3eqPfF66oxFJvHXIMCD
Te/aaAZl9FkdVkMQuDSxNwpw53ABd8jzh1kuOEPYYB/bABYFCTNwzoFQ2oE9ZFjrg0Iwm+/5R4Eb
X97TcqbG0GiEjLSHapT8h5ltS0wN/Z5S9yEk4BSNW7gY29N+SAZSa+L9ojJ4ysyH3+W0kpju1ERt
iRAsoz8RuGdWkuH5WN1wD3rB3ToPflNbdxGq2IBc3dg3eJv1ePQmApnYD0G6Vdx9qtW2rCWQsQ6e
waO/iU1ffTRMZm6Uw2W2wevlnG6nN9jyXObDpsbUwuetWwfQr0kj+Hw8YaI6UDmBuLj3YIpgPfi8
PP7tVR2i3AfDTp3flQC9JENcxVB5b720jKy8CrDmCObo7eNIQ3jPdOEj4/WI3v9i8vWSvGVh/bJM
qAsbkslYX8cTPPtHrKR15beoxQiX2ZqZm9QFWH9VVN0U4Nqpf13qeBtOUYbECa8dmOWeBUIzu0Fb
fyzgWHicbnAX4rXBFWUOzgPX1g48QHQDyzofSWe47DzSWnFPs6gHX0ukfy0gEOvrdY60VS1q2pEk
AIqVsMV8IaAyeggaH1iBwdcrWF3aXHx7nzUQFVx2/oHMllTr0QRg7lhovJccWcL3HkUsTwIeFwxU
STUvguDRD2FAyLqW11eOBEw/gx2wkftGCpyju+91LaPYPp1Mw6qjeahj2xBbH9lYNMSMhlyV9mRp
i/wG7d2cRJhqQphT9mHVOjyM3rnwHkOrn1EKzUQTMDc3Chi/dIfof7z45aOPc2lcjLW124Qee8Ev
dxoer8EMGQOKdm8yrgGXCOQf9h+ZU5Yu46eF2n8EkDxQ8gUC2Ka+9WkRm+x4E4GFDrEaHN9AxCxY
G4JdH3xGRsQFVImqXAeMjlBb59OLiUV1xOCY+LFesWuheKNXmXYZwvHxMRzWOUnPz5Da4Y9afpjT
u4Zs76Rj/T09/8cZL8QLFMklSa8P8tLZT8Oc0dMGP2Ah+TfbBWV+NjYSw39ocj0l/umQpR8v/YVZ
GinycPL2E5dga7oytqH135pFVFsINt9dPlqUzmSTABgnfJhtJfqwni33osCCwLR+Nk6fMZaUlK60
UtJsTrvYPVEuUksjP4nWzQB8cD6kQXnfG/jTvlmjKwTXCPxFomt1GEBxTNnS48qtjqeY8starmTh
pxDrcuctKI4Wsv3/j705UMARRD+scYmOzy+n2ZRTKDi+eb/u3TIZ4tiEnOhHAv2Ykw9qE/k8LRcc
F56eyP7q9na3iL7sd75tA5wXLQbiRvfjnEYvJFkB+QoCc+bIFyzHoUYHxl9lfsXelSg9OfLztO3S
TyThgTCL/xvB+qOzksGdESBGRg/m1jL6yXjzj38oIYt999atM4RNcGbK/X98twT8Cy7bcRurEhmB
ZeoAnr6AuN7yDisnlTAraD8uQzgWFQ0SqiLgsrd070Fsc4MACbglCwSVb2jKCmONNb8WZd4Y4AEa
3VFIxbn9bvT4qK524ftrdW7Yr/PCJKpFS89ceFsmtSZFDa8DuAQVmIike1VMNYDu1XjNUGIHymyu
hkAuDNndXcDVN7GUW7ym224DiMtN66/wtvM12YDivZ0+868yM1E3Y1d+OWbwoBCQdnsTWpsyQ5j2
Ku/wTR6v8OpIOBcOch8D6AOgUjYZmAcIERmisw2Kxrtsi84mGF9mmgUYOizAEZOr73HpxFJ+tglX
CCuRHu92t19sb6tg8JadKO0MZBbkghQMRy7DXiiw9XMBdKJuukfYi21HeQJ+FNQvR5NyyFi/xEYY
Kbzrjsj5Cx8TT/U5bclsMOm23JHBIbR/97Qf8jPgXbDSbzSrz0faFR6gEoKKL/Z/CgiUeinfynCg
FGObpgA2jAvrnyh9e9+xrixwyy5355tFBHb8fKuGexpdZcHj9oqvN7HrX3uARnT8wNTfTfW2c+eq
LfdLWldEqsAsVQK5E6YaTnxvP3+XHIFknNDoLBGQlc2t6sBsMYZrRsyH6g6UUytb+ETBmQBDopuM
+723nGByUGzX+w1pJ5pBGT7gRinmu6Z75N37qVgWK4U6eYv7YEl7EEhmg1VS89F7UsL1rGKUfz7A
R9Bx0kpjjQDKU9LJgXi8wdycQGM+FFsU+A48SeKtIgdp0Jf9R5CKhF57MBS5PKAQl2fHP86tAFzp
+94yCWfSE6ePETLFVaTJdZXRVDdGd4tEPDrdx3UQcgdOiG5WVL9/Cp8SuVdrcTNYUTGtGn2J/7aR
Vw19ibNCd3WycpCmIXyxpAuD0KLEVk01GHdl27eIH8jlnngJwGceM9LqFdS1uBShvnXqN+1wReye
j/aFRE85HqZSoBTq8sUBYzQr8G3VeFLk7ri0zuAziIkPOlGQrK6FoIqBG3Y4V3qQEp0yYX6Td63+
HxfhW5JdkOaTjteXAEak/6uCmt2HVHNwVFjxvJPr21hMjF61vBhU2wUjZVs2T6bRdhao4dMiiXme
v95lfBxFxVtImndkj8+MP4XQOWh4JSPeL/TdZbcrOy+n2rr79tn0+PJjdGhR3f+1Co6e1QjUiA7B
NlMH5qhf1m21iIf+MT6ixGvFvrBOVLbcDiVyK+7GpVRCXV6JoW3aS7Oy5ShP525wAlLdhnrvfyHK
b7rCjccmuTlw3kjHhBC00wyO+9UYiaVP91Ecyw2gU4V58YTgy4kMpCCysXStLgFxBSslYFMbGdFC
epppKLsMa1jGmlLISQPBmlBUyKDMVEVjlCvNRis8oDqzSepFCgsL7cFQefapls7uV5BBYN0fEIv3
wvsTQ/Gn/wF5VaqiodKgi4mchGNnaeXBH9vbgkY9Q/Lk3wpSsziK1+2j9X7s9uwEjbLXk3jwFr97
lSN+TDd+G24/od3ZkiODEWFC6feQ+DOou3aMWvqvPpNNhGsVVI5L+aBH6Y+eyVt3gRTeu4VvIDvr
uiRqSc6KDiGXhp0+6J3L/P6qb6OPQD2gmaBv7j2zd6itrNKzC0LkoUvf3WwRMBAA43QSHxVXm+U5
nYU7OoyyR/hT4vXu8uUTTIH/kPgpylvTHyp/W5MQfV6JNxQYhrr5NsA8DdertP1z6k+xnYBJgl1b
Q+QBCzcHBHaJz1+rKlzONl1picO31g1XEx1c6+dvoUq+WUJtLnhBW8EadyP83Rngfl2EmN/K2GdU
Gbekl0UFGSOlxG5iKmIU6l2qREx7mh8ogTH8qqz/GSGlgdRlFcBQcof+A85u9DOC9Sv9Nl0Vnfcl
3VMhynYRUv52cCc413325EZ0fLzR8o1aWgxLuc6rBP0vxplRdjjOih3fgKs3eL/uCm3iquQJQNys
GmokKGnZYXrmwM5TLeVVZ/GZUBPLOdjeQoytsWcHvoh5idinQJgCPJBqgherRil3Ooz5CB+m8Efe
dVjvTpMGQS+2N2N9OR08klRxEfdf5/5eV08WvK2k3Z2CRqmDtnQDVqE2Y8pj4ZsqHi2KytNXL752
REC9ILEtkeHfaoy/DG5zIXMzPjsJhZAdXXFbWAsCiKEGqxNY2PqZOUKKp/mEzQUujG++2bB4+zBa
wo28dhsX8cWYw0yHpCY2vs5PwH9AXzjJgHaPb4wn8UHqrwDn53E/LlaWLMky5l3Ux/c3VWd8MhgA
weo6Lvp7ODgI6T2KcvcwG2Ce6y2KLqvJyZQtfOPdV79v3nX7XqudUySCEYzgR0TI3c0T0cMrOkGo
PTChjl4DJYZd+qAh4TorpVdUQEn9JJ3Lw8NyXymm6Y5JREbbUKd/UmCrBkq1ah7f7WEZedBiipW+
Tu7J1y/P9v8pAvumBcrp3p1CcMEFTJZiMWbRREf5sZmXwyv8unH+JIAfLencCMkLPNHKxxi6+OAr
IdRFL26ufrejcZy0UVYRmvcV9UJkC8hwfLBQSXr0CZba5PHfejD94RrENL3zFkxdwEINE/BNS98E
NNGU+WjuwllOgqEFvUqaMcOxYRbKzoLAmQn3e+x+mR7fe9NKet/zF3QXKeb5d5EXmHSbfOuRJCPD
dX2jwkjH+4S4bUV1s5EASaElkrZ/slz6IitWDUzRjsRWGQR0VNCzp5XWwrDJMaE8dWiUEZkIvAQ7
ECJXDBrbNjkdpwzJVNWvqs3TTRdSgyf8f+6aeZIJPLHiy85zvBLb3KcIlYxlFo9FOvxzjSHwn3CR
MYfB45hWHyvJPgXCaO5d7k5NrEHQK41iYdSU7Vgs8frBNVWe7A5Bz4kSpoZSgze7oFAOjQ/Rr2yG
7vi5OZr0J5C2DvGdJKkNEs0CDktWTDaU7rIoz6XokoNCa5ZJ2z8Pev57pVeJax+knzeSAJlB1J23
mRN6Nz1h3f3tw3fnoaYEyg2HRQsogP8eOJ5yAIIsPtXSH3OiVZl/BqFUVNcrc3vJhnHub2Vc4eUw
QlKPUjTRvG+89D/1dxlgsc2U4mzHZqkvwBwx8ssGYO1DpD7YiZCapixwDkr5jWFpQ6gmH0Ma6dzG
6z53KStACO33fNvFdHsoaXu2CwElMMBMX9oo7s1QrkdqY9D9niV54yXhweC0mqWrtaNVLAOASDI6
wR0mOgvxApu+xmFX5m7ZV9URFvtV66hRkBh5FJSCNsy3YFVvLxgjSZ4/0j17ezXovrD98mfaCnNs
oFC1OUfp8WJGRHON7l/8OTqif+C2kDapYNCSZeZZpB3j/hTaT8feIMNsSoF45VV7+voETT5je6sw
L9gYHO2j/wXSW5Uwb9iMbQcvGvCe6mrcWttCbTuZEunBXpfuFLMiGRjzWHIziVEYXMFjqDsBCxoJ
ULI8ryA3FPGBJ9jcItyjDHKe//F/DYjOwbhdE8q5E1sCTrSpgUf3OXiyUZY3pEJRFjUkIIlw6hIu
WrbTJAMqCazHgV3gd4cY0duhzgzVXyXLHeaY+mLajVt0SRdWAJZxPoheT6Ie6F2OmFB2ikWUdLo5
H9Y8hjlhMK4OtQep94TOb7katRtsP2i2B2DuqpR41PfHJCAxEtoD70I9gtSmRYr/IWEZf8xe8yU2
txxWhx4JmCNvydKEiCT1JttW0R7WjEfBJvC8cyghD/4RvR8tQZjOBUmMiCRsWD8ObkaWJaycNizD
QOUNa1nyalMzPAvvfqRG60OEJF2qvmFDkLU3GZtm777Zw4NVaJ7BL/GltgrAttWCA8RfLWrEvTvT
4CKNFvxgzfCug4PlflOPXdojeM5fIINvqUkA1Qwp39agh18e4uZ0VQiekTXrhi1DHoKFMJhJC+Hk
M3N3uel6n+r1s+YdGZYxnO/vuFcP9LeFygl9eq4ufB8b93LnRn9Uab160wqRfqSIEubu2OntCPH/
1LcATzdaGD/8yhCIfIB/Nr6unLCepOqfkg3HBvhbyn06iCnnb3NF7Oqy15V2FdFfa71wS7KfeXu0
h8UrhcJVnM6qfXXYyvWBBSx0QuYc2qpQ+ZsUmLBn9zL5vMAxkcZtznlCnE0jB3DnnjSZR73i6KNN
vFyqf+nGs6U74x5n7CjewZn/1insCHgT2pzKfb8M/Bup2h6PSGDrRl2bWd7QD/uzmx+Wta/IwTPe
lWgAfK+pMfgqm3uFhna8t20hVKdKYl/G41wkLCrYEDzxU44k9XcUR6RS45WIQ02QZg3Bs68xy5qn
RdlWhhrPRlucKoYzqrf0jqI6C9YQ477MRj1dUNM1Oba875hacT2nwIDizBQ21Ru5XB4HzPrq2iBn
gnzGXHyovXD9w7RUoQEB4KosRgcG8p085ptcjeidJ4+cs3y4T5+CKq6Mkhl2/aviNX6/HP+38sun
lJh/n1KDvOlA2rCyJgJcvGk57/gWVbulF/7nPTOP21FLBYFLCk+9+bNN01F/kmYxvm14O4h4mWGj
ocC9ytGQj/l1wIU5cSIaOdJnMrz6Ys+fLQX4KW6DHs7lRkhUUuzQ+fx3F1y+y0jiYJq6gEgX+38b
Qe9bSx0DDRrw2fMuHdssxe+zAwGKk/S7PwWFvsb9T4QWCHKYGWdF1JtV4IALSSIqsbnEJQhU8n0t
cKACj9cdhMmk8+2r4igdqspaKSfC7kXU7xYGOGhoMpCe/PuwHay6FjSEhA5+/8oT2NOtb1uDnUvg
hGbUiliDmkjjmmu8D6EP0ZODVjSu6MHJr8iQ6uftYg7kMBYkgzGP7O78Zduj8uQo3S+ik05amNmU
QoO+eQtOxStcerFAGYlSLyQXIw5wsilr5sA+N4X2TM4ogEgcce/qNYVfbKPy+Cf8IQ1IAsBwQPJq
Sm4VGDO/x/TgNJpEPun3AKn6lv5iNhFrockSiu0IxFtn95KTdIXQuPOHeV2LSCicRtnSaqD0b0jp
LslWLi4dIMJVA7r/X5uWmpdkGa7API+q8VlPwax5yIXGHCk53+2OWXKCsFUCJKw3wrrPSzVzzxBu
QBADgBEcHtycno6fmooQ02t752tnjhrI4Nzg5WKaXMaY0CFMkrkysxo+CxhCg38b8HZq2BN62r+U
3swnry+ExqfNjFn813QS6g3jMzte9tHgVaO7VbxrimExTcDipYRTG4PrRou8RwOZrnvnQJdA0f0z
KJjxySRGc4BAbpTd6h4iwxCk1FwmEZ3UqpqrpITd1qyHM8hoHnq12qdyaAASp/nFHCSbqZn6MGFa
sEnmHaC3JypwiwGXjW+yivxewJeoQCaSxGZ3LHuEfQzjdjUkUOdeMlXsaFREqfKgrqEWabaOK4KZ
0xoTo2zjKQnHdDdNw+wNu3cbpoyhqHV7FHBNArofe9o8fFWIUbwgbTDHZJNGR/MUZTUN0kFNbc06
UNCGsJTv+fhg++83Hd13vSchFghpIXmmBsNd7m7Qv1ocrNanlMNZMz4bbefDPvcEjZCqv0xWD0ns
n3GpGosMstibTX4J20d+kEXjA0EUnbJXScnMV5E9b3Faj5VoUKZlt33zssmRE652Z7KNBDwEE4Cr
ThJ28+8qD3gyRNlpkoxgq2E95cDS98W1Z0ec1/0hm7HvakO1S7nc3czQFG36M2Xyz13EOpXTDVRN
pv+k5UvhLBj8uqSrZNizyobV28TPRqwD8j6IZFWaJ38qRoGvibrUFNGQze0svGP9RNRkTMobDymZ
7Vn1t13RM1tmXXmS1sSQRv+ICSdduAg40Zot25RYWua49A6lzyaH95paqEiTVPv5nyzj8/olWTvv
mbG2PcNj/BtdzkIDwbLgUduOAwfKh0DlCaC/4Ujwff3LS5yXwufd+cATUcLQROHRsCSVNY1pySli
bLLoHUkdHUAjTIfdff01B6scEZlgBiQO13pFPvX1gcD0xQzP5f9S1ELgJ1GAvn6+DuyFYh3Z+9p3
vMjio6DUtt/4SxpQW73o+RORY3mLBm7dSx2iqlne5jQBYpaDO3vQZhbR3vECOFjM3vMSoV3peNL3
edtjHq2Nsz0TDdri7J8bXau+tfDh2sTVv5jkMk97kbhkZXo8st7fGuzBjVhWafP9oQp7Zy3qB8mI
1YG6GvzRTwckagQT716xx9/3j5Zal2PPU6JzX2HTMwHuKhp7HJZuA13Uq59HBGVf7HPITPr70sro
jqbwjXHnI3qsKQJm6QkAO+6CN+D28FZTn8fTaVoxMqEi8zzlcgC8qGU5Civ5/4FujksudOvCPGKg
bU4t/JhYgUZSfViuAqaM4tr8to+VSrzCANryPJhPBHkPlnmQGndqFe2lqUG7DVkINl/g0GgPb/bn
2JEcgT1AWX5MXUAMVQVS0oyWaXxZoB5HuoKOFpUZUXTCWDrwyHoxTGQfS+Qmf8bGqOmIIeaj1t8f
JJdn9kYgEKrrT68rf4mC5yAjaXR/lI6h4VdpSNRm8udcFL4j6sPvcPE5GVY04Fc23nvWev8atKE8
kToY5dz/Cs412IfkLO9uVsBLid4KG9xMwHkDnTrLi611VTL6YYFSP3TxO7ZpqVcZm5Xcc9W4zlvv
EgtbuIdJtJIBmQ/07jCpRhL9GdSzG8pEKr2TH53XNuE0GadgbSJeKZuruYvuh+T2XH+GobKXBnba
Dr8juLoJ1Swy/xtGKWaLyqld45qZPUW846G6EAGxNg3MiLwfUKPJghwkhMZZ7x0odkZd+ASCK+D5
vWX4bB1LNrQlFuJwTEomvLqJGWtlz9csuGIsxiOMfri8kQQ6gRdsNsgxSJWncxsOEnlimP4A9Kw6
eS+ugZ9zOA2JG1OFHir0dR43u0tLeF54Fn0dZT/zX1wuGMyfj2WAimC/2j+hT2bYHL+lF8CPtlmq
9TqX+iqs7JLz90fqh+Nmtxtbp3jOhVYT2FUWCthx0Cto7kk0Stn8AxelJgrNkzv76ugjG7Ajt5jb
k1qLIcL0V4+NoaU3rQYn6thegKZCCf4s/2ckWQvG/NNd+8YYgU1wdtcA7EDTF0MYd/gF+hFnVYju
hGE00okYBdJ0tpVMi9IKnwQAMzK3zqmIpfiskUwnKERjaJM1Vgj67fxthCowmFcl7xuRYVzwEJFO
OalXAKVHbwg6T1rMb43mUITxczHYvlrmIJqwPiBcl6yeQ5L04YQCem0tk9k2C+OXZHMrr6akSAuA
c/mr5I/ghfH0JF47OowL6g8XnQ23l873xlUH+Ci+qGq4UtRsRCFStU8GVd7+EZnA1JuIlMkjbxdP
fMcPUIs7PK43Cdkk3V3CfzrjIb5iUsI7SBMv7WgCosyv00nG//K4cPOITlaWTyTFL0NltIF4fKiA
FCdB8blH+4pbp31Hs6C46JZUlb0PYMrQttCF8+PLzKFlaaGTdnu5Rza0B/DjfxxmwQOTFJz7u6yQ
8n2GByrfv0gyuZIEcn2Ha4h/hpwljzcMmMLpSvxPFg+dIaZiHmvzolxXUDu5sSYyKNRNXplI4gnA
MGhmn6olT0aGE3P/dpo+OJxw4HmeKec2N6zyhDUnoQonRpNMAf4BU+WfXBlT7xfD83+g6pKNXE41
/cp02NhKGpfB5aZN9qkA3QUabzfMWpOBOhLhBILOmy+Md0O/wjBEHhhKNAMUIuVrbYXLoc8P88W7
mLPihC1DNr+DHsGZDVSX54X410OiTQlAoKetNDjeP9W/8FXT2rssA2/gT7QtzplNjz6d3DmjIVvH
wfWQ3+lDXNAjwpdeFWNkczl0+EJ1lsOMz06tqz6Sig8LYxKqkpmzfjkVvcZ9C7rk5T3In3qfSAN8
7+aUfRNvD0yije1vuDTP06mqU7ZlHSq1e1gQzuwNGLgpt6D4eTNVx+ngZeP6gHEfkmEi9lMFJEuq
hSZ+I81XMK43QvM0zz6RCRgieu5hfHCFVbi19d9FGgsfGSaxMn/QeIxC454UzH7CBQyexplLDoFt
TbWjiWYnUl9QI17rj26osgd071HEB+JC8+PUwgh5W8H2x5kV0D6gIzXvl61OWpr7b2y4omH+wB4g
3kVR4zXvzANvmJ/SLDY30IN9VP8ODARQA2y8pwmQVCQywPZglvNrXGiVB86esKmbyLKC5+uv3dzA
0O4ULhknuLELH8WwA7RywLVaIaN9U5V4NP568kKW6wOVuOfqNKF2fZRNRf1lp76OFpPmrW+rm3uZ
2CULDiLgqbkU3iTy8ntMeSmzuLZ6uRQuaW0t/ZKhN7gg0FQzRQa1cDvjS2hCXq9KHy1G8l3nrOV+
vqQ3v0Mm2MXeS3D0ppnhF8BwTPdxYhXdx6bjGxcVIq4FXtI6skpmNim41Gd9kOhhuyAVlfcSAhv8
o5+4/Iza2Mc45Ba12Mkly2lwNFwO95bKVDM+pnljdHpl8AfDtyj+3Ulz6EDoS2K+RPRFGgubleG/
0rrLf12baKdWkBJ+DZ3F7OubcymC34r/TKceCU9i+af5tZy9wPSjR9L+iUf6sO4DZiTlnkwrx+dG
Q/RAv4oi/sf7f1o1ntj4cY0i3fh+oPPQLV+oACa+NLW3z4TNR3r+pPehbvawkQwG/SgQP1Y2WhSE
8fHIcfw/n5trCBSUeR6DJFqZQz+o5opX1r3FGgU3iD7MLRzbpx8AyiUb/tGb/ZF2+UdRUVGQPO+k
ZlqsIt6c1+A/eCZxZ7zbz5rAjEtxIJYg8/yepc2sqMo92G1IkI+UbSM3A0Lf9G1fFMuK9Px/obIj
6rCGjMZcpPx2WqjVhFBVtT3dNmLho3246ZPOR3S9qKRJuBHQcaXtYIDY32cr9gVYevY83E80hL1j
hcJj9Kf1nxEDT0uF2LP9doaJI9qOsF6x/WUR/qjqO7Uk8vMYrvtViWk8m5UJsvrb3MNCcOjPo+5l
BWtKZabDz5Y1bar5IzZnSKjNH6wyENhcqmXBUlwnGI18fZzBfL+jEEUjfGVGWCzZtseFZ0DPUWjq
iEdyqik5A30wzvR6Qp/58bnCC++sD8+iV2CoWRA37EnfrsLOprbQX13dAB6KdjyTsdL4+FbRFr2d
NB2y/ug+//F/KJa+trtOQH+b4NQfarhdIXReotpgg8hyr+drSKms+ZWVcB9+gsrDq0UA4/w11QZ0
PM5cI226ogyk6vkKgGwP3SEcRQ9KgmwXy3bgxouDkShNZ2y3di9yZWzZugRJRJbgesZZg1k8rbjB
RIW7Ae9OTIPaXht7d8c4Lt2HFBbyuDyRD5jj2ySfvFH1v3E+v89g12cdKcFF2Se0lNVUk5s21OnJ
cpaHZ1mw9mVxsI/p40lzsB6gPF0o0uXof3peTnTnpunBS0SVXLQt3kgq5t4wmrWzO6MIkk8bpNNA
9OWJMH5RQL3snuk92SICnNI+QbspXfkFq/AIpoqlq8vCc1emS/YujHR9V3PEGYHzKue7WoV1Bksq
cJNUPK/e7DoswwHcWteMcgWJxUiVEdh6qmyc7nw+ofpRxVo/QzPe9dyh2JpdrEcVWxVkwsZQbC+z
ZwXg5/Fb9ZfyQzGyOROe15vSbJwYGCWF+1e9B3/kcgWjP0zU/9sw9A65U/njs6jhL2+IGEoUuiW9
J+pitLrXZTb2oFD60RjOljdnMpEfoeXxO0Ai5eWkmOj7YuQKYeE/mXlKg3h5A2qmbyWg6LR+XGXe
bUkvvVQaacZrnVj/PdBHOCqk/WbMhSbZeZHGhEfOmpW0PP0k+U4zqi5jBwv7j080W8C7AUjd9TXu
vlZWoZ+Okj3/wrrLIZLtcd0gZDDZ7QKdsZ+R4eGkAR9BAKceyAWkRH1RwCA/uUnkpzh0hikCEnLF
bgiRbNpQaMU+qAsOn4H1plXdkmX7puAjoo8rjW5K8ABQF1uG/RTDQR6CaLRt+3vOPyXePIxeUMxL
H2VYsZ7g0HpAWACaXe4XqMM2/sTCunhmt/WNWmJHOEf4qlXQyzIbcMG/SfWv5cUUQwHazCM2GeQZ
JvF8ZEoq58fr5NBKtTaK/JK7TD5VgrJrKs1e4VmstUNhw8mtv1DeXkOn6ZcOrKGCHU452UubDZ4c
tx3VPeVvOchVaZZqpNa/O/2WcjAjpSY7BgvH4v10qVn5rvsuew3MtITmGeVPl1GFmbXwb6qpHQs1
kNGxIL42w3tuHP9NhEoU9gy6GiBmQ4krJRGUdmQXgU7jEYrzXbnhKtB3qpwhUa7hMIYGnv/2XDJx
gdROtC0qm0tvaDuvPVHg6279dEV4tyhsNs6BogEo9Bq7kwyKPTgSgstPZ0e/TEpPMw8UOj7omM5C
BFBNeKw7OLUcAcw3/T696dXHs2N1+mn2ZvZimPRhucodKjKFE/a6dJQ1CQ2LJw4UinR0NNgMebb7
+cOCb4qHx5nxQBH6kw/8VeYQZUVyl/m/I2gOC4rR4OrVmO7ZHyyUAWGJdcE1p+GXtn0X6bH/TsD2
kZl6yBZE4LwwCdYFieBgGfHBd2avV1fk46zV724EjJpBFnc4mDNRgrOCjsZEHUzOpzIPZopyguPF
kH69/HVQFymOI35uuZ4xRYqt1a1R9xjPA7Kv3JxbbarJ9SqecCLMYiPYNNiRIQ4j007rz9p8cH8k
ZOMLlRXudF02xooBESGJLJxt1oIEPCr4fw8NgnB6iaDp7oDMma0W0b8cwlJzHIFFA9hlcES/QjvI
AoeEWzFiS1P6ejkrb/FA6wdMuIZ4rD74nGjtX9NslVlgv+Vf/Ioe1gd45R/PzDDxe3qIXHWWfR5R
gB2NvyLt/OJYffJXjfB8ZRiny4jGWbExWVUoFa+j3pprNQL5P8KKjxVCGXUogtZBFxszKNc7t9SN
9pixNlT6RwNszYC1RYltYxZeb0oHJnd9g/LsSm0VtHc5geXpHqCHD01QFuZfMW3mxpUkkcHe//0z
XAbAsEKVEdtvF7kZaVpj3rvRZbfR4+haN6bHuE3pNxavTXJraoeTqQ2WOOJ7pgS9r4KxxG1lz0rY
sfDl1g58yY6s0Bozho4mRnb/tyJZrrsNVxpiyTiTQxweARwDsThsBoniXV7DtVacJ+r1kP0htl4A
r8UAt/b2fNQlnHX1p2sv/DOlCUOgPOfm85J2kY0AxlattCqMbsWloeiWvawvVgwqL3qJWCl0vYIM
p5RvBatpRQhSbd+Kl4ijVlLniPiBtmzEDxfTJo8bIBu5rn8QPMOmXWSv+V+5SGm4Awji+3XlScWq
XPU4WzflCcA3Rwqt893Mj9x6KYtC13JvyVSoYPQJCZlZYtAFiyTI7cS/xwp8NeOj4e2F/cpP3bYY
9pwnhg7F6cPklGC48OkbUUE1vHB1nWMYSDjMp0cMssAKU47mXOdkUValksB9hCH7/41JrreUq9kJ
kcyVj8Npo+Tjh+sCGq1zGguPFCP3Sim7RHZX40gLdhXTlYrPk8P8dgRgN70VAnqu4L5m/6I5XGKA
dMG+yn1RvYu2De8fRsco/sKVFszSD69ZAYAdMPbGhoSGmUwnhCfNQld2VBdUYC9U0PywEC3L4pD/
EesjmrFkEFjWv9EolsTjo4F1leuIedMONhRZPsZFHrzRDq7HUTEVdMULgKWNG6HNeoD/GGITL6mT
hdZJEHyk2l+VYhu6bvkk15gxC259pdIvWq8BwrBAH/xx6bLgI6MesN+Q8209Bo/9o64MSAAyvLKv
mEq/6GdnwHCN3x7q3/FoYTvFlI79nVc3RsL7hyvgB/GAWJTXYNktryxz2sDqA93h9ktAh3XFk+ra
uE0O+ae59B+pZUh9OVFHDLx1kjNIsLaRdJ8k94qHPc7L4YZ6fXpqp866J5KcfLm14H3z+hiff98v
zeZy4VYRdJaqnxbKItY+sGcenqAqVme/48L73+7hM6D+gjVu4ZEmUaDYmEJpmxE5+hcNL8ObIpvv
YVHHybwIiwloGtipGCFCjwZh3MU6YUSzQXqKDY+OhOU6/8C1HAZoGyTnPf8OX1qnU3kELVOSqoZB
C/I92iHjL81am97XN7rqGimMeWXltDYbWftSQQlCk9HJ0aWrIvoJVVQodYnnh0gfEKqOAX0aw+yj
wvSg8wY8oYKk/gfIsQwp9IOhPgdddUlYjX1HkfN/9Q8vzs1idVPGdCKRN6zIlOi80Iu5fEwqec4J
lioQf9VDg1YoCSfAcPrMIRFVFg14wheRiEY63uAMJSrZaV46DPSy95M4ulqoiSsFiwCyodbADCFg
308PMaT7+80McF3JPMSD21j2RlJE/Q56jUHmnsPMGDPnGOB0JsskGJmTg76LRtgPQSdcdl9hzLJe
tstEyx5tGvR2/5EECAirQzSj115T2AId6PfaPvk7ZYqvlXIsOYXOc2WiZgRBNu+ZjtosAemue5d5
y/ZgHGTjlZVmo5gt4vJcsTGkrTsi+ZSSvZny99sbg58CYT1m0ohupOENy9yRK7+RFhcknq//bwbt
RHbXxoJLhOCbkmzAuaCkSn9f5GbK4eJLyJvm1r7La98vEpqqPcWW2J5Fy7m8uUFPn8oSt1WXiY8G
zDfbKyLLaKn/SQAy6A5CQ2gxARQzSzJs9W/ogkuICR5oYv1siXfIXQhZXb3lDmE118Xz1yM5QJfP
r15GO8Z0qLr2CX0foaUj2WdH3ilhKTzq0Xn73gkhC6qYRykM8s+vkRFnIiBfQIHBscXrKni3KRz/
AiGv3zbuEF7gkhXideJjdotYR/CG5Z5I+HsdAXMi/TfLGHL7xD/QZqkcLkKUUIKg9eh4gPws7Hfk
lQKdtA91hfSBJNKmiNbcg2onXD5XGad41MzttatF1sKhHIrquCn1K3eYqCt0Xu9+BDZIuQjsdghr
u3CYxWEVThPDDl/wu/79Ft+VSY9poPc+QEMhBwjuF17Va4wcQ2SKyt+py0NsQH1BYEhMgCsu0Jmg
6Pbrkn1hLuGN+QjUm8KmrK4usrfa2wTdjIvrh5UFzN4ZIOXV5d+CIqD04Dk1IgWczOUKhQqmnB8o
WVSuP2mO2XtTjU+mxaCFWdYErYZgZ5blJVBs+i07LhjMBFA6WewrtEK4wh3AMl5Twgf0f24ixv8O
Mt/SusS2Ayc4JDxp/5IsUZBU5MQrRzRmrukurY5eOo/9euZhhjhn1M2qwtmdyyz4CumJ93/95OsF
oCWtbXeLZcNm7ESlOf9K1zIeca322DbgqpOuJddie5Ih6+zYjvDVPDJUTFFW70YHnbDpc4PhihRS
dlVl+z+Q1IXJJ1POnGHdHZSzg301BjQ70P1fGlhRD7Ett2tcKYkzPlJqafC8ozAYjJh3lAh5FyGK
5TF83aJNHGsIX+mLI/XAyYrXN9RZYCdvfA/KuxXADO7jKLs3aLf+qT2SbwYRz3AeBFIuhE+y5N42
8IpfVaF6UKDEVFw7OcNMAR+L9cK58MTBzXlO0l79EY3TaD0VKskcZ9oiCJMAI1+Ft/mTYNlGuAwc
xPr79afod5VUH+8nUU/CvPB1rcTscmJ2cexiJ5hg+gkCdgCRMLTIjmcmwHSqaSoswZ/ZGEItsumo
PylO5zcGXiXpTAeqZqyTE93wbV0DVkGRbSmb9QJt+BJgGslRoRhepbP2xvoPEJq+Bx41qkSHhUJU
LwmR2sqsXOPgqxBVSsyyywXmFU9lwa7Y/TbncO587Bx7Nxx+NYHRlpaIokHndmRY7yf14FG7qkEj
9xSwvLgnehu45Y9XR1H+2YBO7oAKwxbWbv9FIluFRRExmhq+AhNu+mwDL4iL1ClfOI1ZV9rXCzbw
GMdfqVCavH6KcybzkcZ5GKBZTlLtgeUg7bG5i9O8zG6HUM8DnGnYxQTX9DBvCkH5R/6C5jBE/9Gp
l8EFQE/Emj5E7YiTpb+bXMtqKkwIjTdmhlpi4zrdnCpyYjnu7uAyqNMyWJPpGjCM+QV/+7EG2Sqn
URY84PLbIXOtqNfhC9vIVQNnI3pjvxTWK+PEeq/EU0hI4u5sMAT+JhaBjtYD4e+GCpvgUKcqRohP
Erej91+3SJPuNgX5s/N4Ut5hhkFFl9ag75hgPe3Q2VZ20ky2ZR+04GSHNycqV/9DHXnM8140gCLH
RwhqvL6eAlLMBO7klVPTp8pw0RXfSezR8H0IcJpQATflfr4OXrHSTzITrVsxhMNbGsgjYsU+mPlV
Utti18uuoYtkBE8wIIzRoFympoQm+EF0AShyWNP9gzF2TG6RjXFJwi2xXxZVyDnvsxXBA/GoGWRv
BYSqKWb4gdsi3M49hJpQ4XubBYsl5rgRv+Qj5HDDgvVjAfN+D8EHV4f+ZwCzUZONVGGtfjjWTxyK
y6MesPC+1D7KJ2faLnilJrfJwk8QfIIs4mRSOGiTKotuUFvem5kET+ax9pHH3eS75ZrXlojxmXw6
lD+bSFw4v3/zn5jmYHTPujXMUhUVEkHWkfO+0o8sbQXEbCopzhNw7+a+/8bL4VmquRYOlQ7ftWHB
YOj6kFTghdxPJdjZmRCotQD8GpjW9EiUWogLnKpeTYI7rVy71gY1Gwu+DVWSPQXAUrq5Tfyk4vXB
B4FrBK/rcxTlE/u3gNbgiAgDd2A52GMqEF01SII/SR3S+1GnZxOWPfEv4Z5/Bqdoxz3qX5b55huT
QGqQ7P9ZR8c5Y0dfC0RVhaT5onCbGqp3hdkDLH6yKwj+Zdkyw1sj3m+e0iS0FV4LfDxsovGAnWF4
7MQZYk0zujWardYFXnAvM2U0jTHWqmL13QRg33l+VRGzsreCkhIzd7tYOw0VJyms0ZZ+2qiuSSI5
bDF2qtAxZ86VaD0h314Y8GCHkeKlH/Q1shR2zKwxIFclPlJ0PA9EL8Hs3t18PXMmU8UrUfifwTCx
1coctiUDw/ga5EufPCi/ctOsO2awZZmfZC22FgIO6CWvymJzGuC+kUYVwNS/KMWxxcvAU7fO13Y5
pbHSwMzFhXOgWKstFd+5LGT5PgQIMS3/bj1a42ON/DfPSG9jkczxcICqfQVm+o7jo4CYMq4V4YjW
GtruvZPJFIFUE5prcpm/6odqELPkytFNeRS3dkqT30jSv59AbdrBzEyFefp42b+BYQD+MXRoTgbm
cMG6X4Q3JQf8lfkhB8XLkrq8XoudomHpv3KnYNlOI41ch0yL04QU5T+Iv1d0mBB6Y+N5cS/yBK0n
JivU5xRWnL3EuIcaHOoafX97yrb06Q93Ksjc5ZkGBbRLG+yZi/qhpPqftInwQ6Ld4Ia4b9eVh0en
8q12Fl5/+bNQdLC87qWvSvSPEqRcV0hJd8zaeH7zMZLB4va1cbXj+i2Yia/7ap/eZqbSzaFt/5zG
lSsAFaXafgHpXp6lYu9QvUJBz/sNGkGjiCsvcyzeRVNrjRqpdx69JHBEzV2dEpoVeqUtQp6feSp9
4huNP0xM578S8yOGg2YKNtBwNx79UIiIVpBlCvT0CDdN8juhGo0LgVEqYk41vaHFMjQQH9Fs3Zts
OKFE+6lusFB/f6pxqWlO7XIoRII/Ch6UQjmCqwjMuhaImi37AHVR7LxtpPdS30tcIZLVUx8yPU96
nXSWbylXz/gSOSeNXCLVKdwhdt7dZvDoKgkTlIr7l6wFZzk6EJy/xfbpLcFxzvSSwokYFUaeqTvI
UzEJJoWY4dEeGTZFbcLXZKKIJPMfJKnT2/FhMEduwb6Ktqizu5UUAGvgGAF8dnLMFcXTQwolDgf2
xGIIvfLPRSi6xyig0cPtCBWcq16ikPvP8h2DqasYhkhD89nNB/aEaHk3qN4oLMNhkJLy60O7+B9+
8ueit8qcVaL42C5Av1B4vZZPr5wQbpZzMIOHQbz6ckgA5cKRpOy5GqtJ2l5XfF9gpcbcRmDvzUkk
VxmR6IwlAHn7Zx9svXYeC3643UjFnMaJZoz7WGBiFnlcHK7MA4VCgepeOK2dFtCdQ8R4JKfSyZPW
bj+mlyKtJ95eZTa34RWtsQiKBuqEiIQKMFntb36D23Zp6j0K70sC0JGAVL+JZ964ii6lc2hrPs9m
+9YV0tSaUcV07UU2BVmr9zpKfQAO1UmDH4uJwsfL1sUEMTzQE7EiiKnUtwGq6Ur7mjk87z5/fBdg
1q5+n0Yxe1FsRt6lBCstmy/Pqc6sYEX2WRgds/6W+Fmd8wA8YJiwbDRWAp17ur1fIoc1h+sUw9uj
TwfqvyTUQ8Ypg7NXIaqNL5TyVQ9gQZVQOIrZrBhAwcSs6fIvO157XWkCpT/WXIX/HZXbkwzOlggp
TRO0rF6LW7JmF054cNolVimxI9QXQjLhRHY/bAUSS6CYU0iboHxBVhKZjmG+9U+f8mnkzBZV9EeW
TDTrZJVCNbScbWqsXVR4RlnBwF9FdvuUtg1g/g/iMfKEDoRS9x3d+781/9PnGwieOnNQHKG7vrwp
vmOIOWLUi9CTjcwQK6AbPYkVVmDLf5WnoX7plcEW8ixbv5a0m6jlgcfM4CC/mj3+Is7A4xNQqWw9
KP/9Xlfc+PmKiuACQvWa0BzUWQD3M7BUIwmyegU/UBYgIKbHqpSzRhnDO6TsEgEC5I5X6dkZicHF
bKhBRsTvLt+07haWGjk2AifKyjR8qE+A5cEpCgsgXwobH0zVIMM/Dfylxfwx1e++tebMy33fBBTv
0MuY1EEzfwIf3DMZsk9Kdy7dcoguUEfpfTcCMtujqHVriXTadKkBAHQi58rg/V+El3cMcdRmPa+v
Lpb+wx2z6hY5i6BYIDusyth32KjlQ2LWSWNzvVAahMwBXszuMVY6zFqhH6Ct3gFkRTqGO8RcM1GG
yx6tOckTyO+l6k1buhlnOKcEfNH0TrlXVW6OKKGUf8sDJk+46f2y+uGp/9xTi9ghxDIC+96NcOt0
c3amBg1zC/OSnPhiSoyKcFNzeV5orplqQXLa+zajvO3w6uOgqANPW5gPEFUK/AFrHEoVXwLw5dO5
BoNnu2l/zH3qXAZkZVrSqo5wz45HU3b8wgfA/h8X2sypJzhZYIrzwSN0vx4BCCpfyBxOcmyuKi4p
ZBRcta6HYJnuDw21GfY7nP5e/OaOwcCXCh0kmfSvukJyKxB8/HsN109HhOAnz4IeKrO6YMXmljJn
MnYKlXuqk8XlJiNvj3nAOwZk9PQGvJBKR1m7s2GVOIcpxbO7QstuCLBf+ASxFKYUY9Lp/Bi9WCvO
W7d7O29AGG5xQSOCiL/2lO26cDbB5tECXngZnbHr2FIJwwsK5iqztvyHRQZ+zUQ4nBmrtkvbfYt/
jju5pEcENUY0mE6vvQxgwaNh9yHOPnjq1KwKzGUcWGP2BGQCkttgkTbhjX2l4CZ9+ULuRitctEb1
iRzy5OFLU9eyfcI2YAx0GM7EdED6o83XTfB/yUYah8epyo7i1+j8pDqTDniu04iTrwJerq7tK4CC
UDN9DsEL0oWyO9Re/6QchAP5E3lHlTrWK5pHrwGkFUwAmS4SpAn6q6yckwQHBHH2TpZ6DzdTyk/q
VdmzooE3mdTraCFlP/SUUU3vEgMOeeJjm8tlimQjS5XnjHLaLuyBu4RofM9djGBohuTNhMeMaHnq
WRlelu0JGWaCqSEowhzcYMle4cTS0rCLj2/E9cx4tjFIgRz99DAJAykBBSHxPz5Xazgp89cQP0aQ
3N3Q9U+Ur47zptYlMGUcrqWUpR3rpvYQkXpqToB6ntuBf7nSgB7fpF1DN86NXIGkslYSiQK6dozO
cLHJrTRakPYFhdsDDg6nuLnYfp9XRAqeoYHS5LvOEZilUeXE7v6QkUNqowSxfTiaITeKvDm4eoyB
+AMbvo4Um1zEg39W3Ww/0wqJ47nnopwSj8cZfQYD9JlWiy5yB2a384/iErXyD+/C3eylHYFGw5ek
ltesfQPi9aKYgTXiAJykfK51o37diKsu8NYGVBHA+5o4wYCb9jOMDyQW0GyHxd1lKbBt+WN4bzbz
3kYDvUBK0YOWc15IeYn4Jw0UTXBHKTRakriqs/qLFHgkp2FUc/YxcmGPf/Xde8K4tU8udQ933BEC
1A+9ZqslrdGvxvALcRJ5V9lZGuOotuLry20Jz3z0jKSTXb7eGbdC72ba1pO6uGetrmp+ZLxqoVR9
sk5DEXyO9W4U6vWNHNwcmcGc9BxHOpa3RqPqhiqgliOzvgFHQ5ds9MVmySuArKNeJaejqbyRixLK
zMaQRWiufCVvP6JzhsLgC884nGkvJUZPAe7TAWI3iqh5BUcXxvRfpw3bYo24x/VCNi0D9nzeRv8a
itcS1eqMyal092beyrDZ2GXBVuQFmfRgxASQYAxqzTHnB9HFvc1md9/R6LtsBgDXnv8h5GPAHcTe
zNqIbFphki1q1oyjgNeMj9twWXV7xBtJp/Rf9k/w4DfYxnV5xE3LvpabNpT1o6bKolxKt1P1sZOY
Y6VDCcP7tTI2zya6ao8cXTci18y2i3iN9kp1qlQRcd/FXwCTOnWOlhz5/rkVbESmr4FKRnwzKk6h
dKM8AqU3glno5r0tgOTY+cUz5Cc3b9TS06PawqjIteWcEXTuGLbKznExf3QEaZARYbL/O9mb29Fp
BgorNkQYqN+l/ZCs+aLsr4dePIA+BFIclFP/w11Le+/zSGnFwp/LLpLXGp3ejk94Tr0miWV4DUSz
YG4/dKABB/xhO7qnes49rLHxGcE2TbzYVJhm2OK6ojSBkugbfOVPYh3852UMdF7AfSWq2otQFiyg
Gj/qDgY+4SIqbU45Ym1Emokw3e+wGAjxOZ6/2vxLiJDpr4qNV/tw2lRXAP0fpGuOyo/H2gV0YkuS
Q6SG+pG7DpKjuNvbl0UEDmMD/IVRuo92OvTvE/m/N4EPEqqsy8on5/K7QTaGLpzrF1O81YZNBt02
1715Xz2GvPhBahf9DuPeIdAA3Wr+3bbpgjFAXBN4hVDqlbe5qTgQeT+lqo/AEbYextua6eouxxfL
PrysETMhAUKVKOc9gyHpGfmdez9LlQvkvPNp/uyD7gQTD4UvQ+xEva5hC2cF4Lgo8eIL3lMqBTCy
zruhbb3z+Iji3e9Bpcb3rXxntGj8JWCvV9WTGXyWkDkhTn8eXkt5irp1TcWIPwPbkTJ4UNfQYMEk
jPXti/fzvmKaXD8cY739ykFgAmk9p4PDQfV7OjvZGdGpY0+5LUaWhHpdSIJ0Mf5n6itZMckRrcJ/
cdMdVYtvtXTAObkCPOK5ZFGOAs6njk40CoKtBZ4+bOdlZyQ/b/ZA/ZidJOR1l+IP39bMuc4sq2Q7
Ae1JRKPI3lEbn1sAjBK2ULKTnhgqsJERAqidn+v7f9slNlEodKP7suinJypXwQUy+KrrjfDzC5/u
G2QF5NmrBQHfYYZI7CMSdYosYNgKDrwSxh5Nez2CScsxLV8MIrx9pglhxIo5go0dy9Vg8mO6ulNc
7ssHm8xFJQi7HYBTZaYqBckGUg1mUOOfKDjU7I3obCzqf6DWUDUFPkjZ+LYKnFZKaym7nRnYzNqF
AW+3M4J81cRF4M+xLiK0b9tij+Njc6tYAl9pfvq73UVXIlCcm9fGr4BrbaNrS9PpoT47aKMgkRJT
+ZXUJw6iJynfeOjPqS7+xiu9T1JkR7MbVyXrZo1nmtmTD8/WpSk2KSdwo1Ela4KoSv47XKjzd1q2
K+he/QjVBM+L3pQ1EcRgFmTOWRsf8rhcnXZUxPiHM5JDCW+vaUWACk4d3Xsck69zMT2UBszH7mFW
TAAm1acoH0b4q4CHtqGXsZH8v/DR0kyfuPr7+poKJo3FfU34yX0CUl0cIbUrsTazWMBXjcdjVPOa
h1HF/5e+T2bOnq7XG5evHv5+F7edP/6QFLJulN6E0U+3XD9S9mg1DVl+FFYkTWLufI20DcUcBQUg
RDeurdhIRcHqyJYCelshDQ98qf8G/GOGN2kcasXgb1tWbWYLPUL7yHMixY9PrEBnEMqIaaM31LrO
3R0b/98L4rU4l7vSC78wjTWwD+Fkq5VqnHNvZBQ9jEQWh6juJl9g/S+YMrXEAP7ni8WK+rLCFXXl
tOnNtACi7I8zeaBIFPZYJ/8my+b2umlROxmEn96LLmb8nMI2LNzcI9OChERXC9/sjgYMefFZDJJp
ZuFc3AsMt+1quXeXVz80pDBDB66uGpD1+C8CTsS+tDakpKZye4G9xDO/wQ4kIoESrYu8Ek7CrZba
FJ8wLR9JdvGZVDxHWHNrF96t6uY48lmvltrioH2fF4h3ESTlXlaeymp/YeIZ9ofEM+k2/PdTPRQy
owfNgnhE+hYkP4iVOGs+A0WSQ0lG4336wxdX+WQUtXXEk3V4ALOF201czIUBsofRaWZq0KwC5dop
4OPksAh1IF6B+U4Infkfu2WFJjzQ4Ml3uRU+ubcRPBCdjdg/9oJkcVA849sADdg7t6Tuttlgphnk
vw/PhONl2dBig2swMjP4bmA1GiPpqh97AAdPkfq2fwnR+8VNOLKjZAxWPLspRPVYnjjNeHm3fHih
zLoI9TmVWTv9UZJTp5ZgwrxVoZq1ZzWeQV3pH9TSwfswJG22nKGcCZuxnCwYOMiacMSz5T5EbxV3
sOoJ3VFh4jvVyPJ7PEn/I7CSY/ePI2Ed2GF3gRoKx9kbmg7mxA3LRhMyDe2QHv+51XDjKOnGsXLe
njxFsvsEfIFpnbBWFdskUEmgDLti9Hgs9uuB1vjCLK8h9dUWZImc++HPNUPiZKs/7LN8aAwFbXy3
rVorl2RFMmfeTe6XzAIT03WiYXCq3Axb5bpy5nLPEcdcq1pksc/RgSvxpJs9S9PpLP/Wg+ZQ/3xp
aUnWXCVISaywQqLSynkOwgqliWY9UUQUVijGVaojqHiRZ0X6q+NEyFt/gLsAcuktw3yl5PIeInxy
WkIxj9It6jtEJKz330qjghWNG0mM1VNRA8ustPg/Z+iyeLLEO91YEQD4rnfIyWI763k5QcCSX5Hs
bdUCfKPlBlDjNkIZ9aagSR/+ATmdFg3IqXYg8vMvUHl1U7AAtRsEqYTpEJp02tPMxDq0UeHjHISZ
fGklwWdoOxcMOx0I8f450v1bEwDvVj5rFYU7wwy1Dhj35Dxd1Kc6HgdAsrYPyzVbdKwr7T0922kW
llzS/MqKhdISN5Oiw1iScuhlv70W6sxfz75BobuUKnQA22CxxoEIU3gFLj+7+0JOx0n9Dlc0fwvm
ZaG2m6OFjIsmuZhmIPRSxvl9YOsHLAwk91UPpoC7bwhLk71ENoVIOWfnrPiPjmMzQ8ouLAyB1h55
2Xd1dYVfMtHdeegffBczphOwsTu3kB/GNtEALBsxYuYLqAY826HZ5TZDIfSuoz3JR4sJ6zucTY7j
+pfORVbq1G9DTSKjGiIdlHxDFG+FxphMXOqF7greWHpyU8Pa+kkO9C3sHWqy+eO8PsggdnBJt9I5
QHwOlMSbeu2u2bSFYOjiSqdMWqJM2aPw9bfBioHZ9I2bDdCLKupq3gsMHbVTKZdA9lj1rcOgtjrl
P98hjLAa70E5VeG6jc45AOzrMguRBx10OSuqYoDCchlfvHaTYwqp6Kspw5lgRbl75HpLaODj4XPK
FfUOySYRQbB9k78wcbDkmuW9MOVtE0R5tJ5UekQZxb4VciKs5kCCER2zEQZc7oLXYnRQKFdUjVlz
pGQq7z3/RX2ImE1W3+xNIUcS8E87oIVMcUOP/ZmJRNxI8x4xraHsxVkQFbR75kxy72HLbhHUSADu
9gEitp9PlbAWeYPPRUWq1VAzdlHFQRw6V1G7gLHAO6o/Mq6aE262AcZjJYtnGwtNJ9Zq+BXsJ6n+
54lsdnWtuaOXp75h8oQLRDEOJiRoclLMwEVc+99X5hg3I6A04Yhu4zDQ0GyzqYtfUcnDxeq5CjXD
xNWooTZaEpngAl3cfI5A9epA9a0JFiYcppHWYT+pHVXQ0ro6sI2n/3ceCk/L2nLrXr7AzNaPLx2P
HbLw3l8T8ZPlNDm+bfOmirJK2pk9PgBeWNksWOT/gcJrcIYEl8dMHRInOjfuZff1sX9Y43JPsanU
wsVQahZhEBcmz6Jy8EOFFsaLy4Hmbq8eGyYfSXqNz268Cd9iZ+xpfTLd8j6ZdlQsw6NPKkJQODLi
t+0LUBploPvApvX5Kpzo9R0Au/8ZnNr3icDd1i6PwXFxwNDxFpaS6ftX1KiBVWuJr8E0KRNTkcyE
iCbK2zeECjWJw6kHdegm45imsYf+cLf+EceJCtn63fTo8gmu35GdgTyGL8Q68M0hCLAOYW5r2oa2
0WYjzfMpDBgocWkMuwmcvTRUD2rryNm4uSSkEZu1Lxnatsr7+XdEw78iR7ChEM5rY5oFEMQLwsfv
d0nxlqkq3XGl5OFx0WYgjcJk0ye+X8F/xT9i4MJVBox7XoCSKWraM3piqOvd0Q0Tw9m5aukTbQ2M
32BPmObQjKCfh/GOWbTGzeLUgHRLKejsKJak03USYH9atxXdZH2RdqRsCOwCGTXLa185PNYbamZJ
+UuhUIv8KJmSE++xjAPQnMrdLMKwajGy33BknA1SJXH2/AddOk/DB6ISpRNw8O+j0SEa+Hxm4mcl
t3HkdZwH02et74Kg9cl8tWjCxS4W5/tF3j2cs7DpvkW4VheXT5Qddo8np0VGNO1CRKF9HYuexouF
HJHv3RUGZJJtYS1YqtVzHdiw5mu4KHJECGwYz3mpMx0iIAlBcZdDpDrgV+D8ljzS1EOsNPX33FnX
2VwtpwRWyP2JG1Phy43tx106G2jdu++b6pqYcRRK9kxyWXI8c3GRl3it3aZmhqlRZxSPFN8MUGw6
vyRq4zp6at12nVaNUOxjOLX7OLSu6ijk+rShPQD11YIxNkT3NdWHggAd59nMCS3YpJotJM9t2I+x
PLeQS/IMAroA1HmsXHV39mZ/FabzGGJShBi8OAvfmqaIq/zGTmhSG2X0AOOMiQi4+pjEE2jwSzFM
fT79egjulnY/p4UhSGoxMUEBp12dKl3Ea9TqVdi0uTDVzil2jbU0vRHjGZu558gVtNQ62aTXpEIs
67igJDjwWil8nD7lFc+yxlcoBvRTCCE3k+q4XfLLTcN3Nioi1cleMRxkQEpuIKVBkEo8nc2gLH9G
W5tH1lyzr7OKrKCosZuTM4HfMoQtjLwkfpzTMkeeQyuM4WKMjqnNR1dDTEWWY9iQId+kFMD6jEVx
ccM/fOEmFHsuINfG3UChcNswbQENabwPYU1mje4unXt4AN1CgokUXJranx3UWkMvQd9yEbmHGedx
V7RnNJhxCvJs3HQPf91XZk0p5V3WMBV8wCOL5d/IWXe6Jk7IJsHJbg1ucNe8cQ2sBU5kbIeoUr5/
htUcFwvrdUAyQY7UMdkQEB7XQBe/zfMojjQU47AIyQrlEfftYBmwyc69L0xunqHf+myXjjBhfpdx
FnhsmUdvDmAUtBhi0BDExY43Y+LLmoFLZYXdLfDw+rZ9+K/ZbSHz7qs1qMLeqNyC9YMUreWFMuZ5
wBhBKK5psbIwN6h+EzKos1PKQAHD0/E/WfAYecvewsPm0Ce0MR4hrr6RxJFpVrU13E7JmHS8j2tB
5cv+UaW/UBlNYy4YLjSVrY1UiaGCcl7g8NqcCLePUz7VDvqGtEsSvAzx9pJkFdDyfqmGonMEzhQJ
U503VteafgpwyINiWgtaXBr/Ne7ygVFsDci5LXHLxpI2rJ5jOUMkIk7RvwDokqty9SVfJjK7W9OC
f74icecDpfypxtlSgxpn3b+VY1uNpI0BsRt6Ir3WBKRKlDEVubTpMQSJAX6G2BAMnUCimB+4qXJJ
X7Q9lbpy0LLvbMSbTUS29ewfN0ACwKgjYXoGJvvnAEPj2fA+c2BCEwT0N9Tsf0Q1lyKkESk6SN0g
ASgKttD4f39uWJ1kV3rPc+SyWWuNdWeiyq8HvUpNE/H4deCKGT7gmvVlqh9fa6LcsVaZWL9BybJh
aufDxpNWogQGNF38UjV9mVo3dKMo5hNqXasdYBSCsDSMZ5As2wrymvh5to0U31lII1MZI5b7Kuv5
VEZjtFNi4FpjQYBYBsAJtAC61qy3cv8lSm2UOQNt/Y4yT2ZSLyvgkTkNFK9vP4TeO7wCQFOkS1IK
38u3+T63LO1MrVjkkZi4yZkHSMU3wdRre1Vta3gGw7tWH+VON3cNCE+87fHOQRowGe1KsDxjYYuL
x8364sXdzq8OoY9Qd6jdm9+y+IHz9OzFfFjzUMwnPWmeTctF6Yc1jmhi8bDCe33E6Cx4pkJ4WW1S
cK4YAjlg76/hgMp3EnqARCHxUayRGwEmnZRu0MiYS6C8ReLa+kg1sJA3ByK0MiTaQ23qhzqM7Ltc
j8htLEcgGNOKjyg+CTUa2YP7xJOTKHPdNquE+plNug833YVz+pc/v0WMMjF27unQK2vgu/ZQwsGU
Wc78jsT+nOhhB7qZXk8wSZd6hwWyCK4Mp38lwGkDgw7XdHUGn0vCZ9aD3ovgBODyWYoZpz5tAamw
uKIPW7VCxf1zTx50k8PBQgyIHwjuqEsQfTAcMGKAdLAYSoe9/SHU2LOY8A9yhWDWAkDY6figcGNi
6yT7dAfJ5RY8Pc+7W+4Ny5oUZMRHHlgRsouKoc+YvjvndUo27ThI1ySql9/UYtaUa3xTg7deEVpi
ubgemTNDzJXQ0364HUQQKH8bRG5QND1a5bUfQcvlEmM1zFscqERqm0jIaHK1zYTkiS8yFBdPgen0
qj6yBBjKzm42H9z1iuLkGtbhElYjFgeL0cpmjIlF9d8NJoIqVajR7AyHfmFlkwxrWKFhe/q8zbEP
/mtLntM22q+JTFdQgdHbcl1JXjm4Qn7MEajcLIm7HUnJe+2rUqE2QkqWR0Cx6t4dOY4QkgPwbIVd
elINhI9ro5DLNRXsfB12rB0Dkr+dWCrC/CyAoVUHTKS2Xu0Himq/qhGOiIG3xviiZpIg9mzBp3Mw
+Gwa8ouToQ6fic1TzFXAvgu/lt+S2PimjFQ2/Lq6cOMIdCihuXA9UcOy0qA2bj/Tyc9PMF7qT3Ah
AcjMud7LFkFiyCC/uaMjuzMlpGek78BqLWvCJwU6OD/qE7VBIYGuhlOPk3NSdpHuiHJT/o5vnTBN
wvwTZ9rFCPURaSl7TpvZlsThIr+pcdpxLC3kkOSG9bKmWi8ifoalrIyZHfoU6WMlSZuDWKA+ljzI
qxugrw5GOZweC/hewcOzZZvEKDxMdJXAw3vB8yWRvwpGBIV4nBwyvN9K+Pur6FDM0Dk0vqw+Wvu2
ywuAejWpd/VcRhEOoXn8zXJ8FnFcW0H2L2qxaksP+L+44Vprk/kxyI1QKBIp2vyW96rZRPI+mJl2
9qOWb2ln/LoNHK7kvxRcAF1y5wkjgZliIR1Dn6WnaWq6TtWe59WJlhWdaKfJUISI9xkk44WyMfuh
ts1r30U9CswmNyHUs6XaygFXWYsDdVG0axHg8lwTOisLH55gq0G0xjoXygd/i+RzbazoQjMOjIpv
ZB3wtViZsSrOsICG4ok+tulwYSuRjlc1RXZzHC/AfyCxgw0lZ/S5NK3heTqki4alE0+A5AmiqEyL
VNLKv7Y/A30TAUHjtZKUPTYB2EwuwfqWq1GR9oKqQU9Ks0VAPiCQxfdP1ZMJQcGPTLK3GUIVyQdt
tsF+gRKhC2TQU5trgi3InTuT6kngBIQYl8JsyrtHgvevLO2kYv7/sO/t22fSD4kObwwPDNtkiGmY
E1N6fbsQYuO66t6CoUg5bkeSfFl+1pBoQ5J5mzjHuSVeoRW6LlbZThd3OPmw0cgnJWbDaxazMcdr
f4OwAyBfGuhnp8ZZem+NDwGS2WtMDVm6BlPeX1zhYanGuEHSltj90H9iBaVPEuYJO7xgNIALWAvn
D0hT5w9FRUM8dO9Pti1rBgRRiG6Fi/SG41qvjESpV06h5NOQUEarKtC2hSS4Wibq7dECbuKD4qQW
/QWdJeKAePj+EvjlpURHpW0K8Lh/dsmdsFLrH5OzBzZVQoRiMR63f2R4sdOE7xuJGwQtrQ/gYv7N
TYOyIJ2ITkcBbK+Jk+ibYLSvH+kqG1r4v55LZcCCDu/EeEzmU1mnINYq3I/q9mh8TKOCIp73OFEZ
Rki9eWrx/GJCzg4qrV7zDaGHn4O39W0QMr6ZDFf01yWQOXIZMAHj3Km3UJTxLferqo4+3Y+89v6b
bGIyV7OB/xQ8echRNiRdRYZyuLk8880jEjFUBY9WzftmS2yDVvsWdMBf/bN/xqg2B7C3ocUoTAP1
VsB/yKgt+Zq3JvwVJltzq/plvKTtild1ii1wbSJITv+d8Y+4unRhdJu+XC+MvYYRQtyOOrKbIdx8
SC1gtSRTH3G47Z+ZQjd6UYWNsjpH1u0LNUfiFOhA/U1XyjFuB/lcGF8S2duvGamfiTUWbmp5eUaz
iX1diaqR4z/DzHV1aqiK18/j4jAVMcDq9+MA9Q8Z4+91MgaBNCHgy4qr8TknAbe5nq+xiQe6Qg4c
BgT4s4gH6BYC3v3hRieIvw3w4D453LS85HG/Xcn6kbukKG5ZiMbUYT73kJfK8O51yitQwqW2tirL
m9Q9TCNrnxTw1WEH1dikOLhMw9BGmNt20IQUkiyGKPtVE3sE4HTlULAp0UzvHbcsvKSFTpFhGFJm
WwaHzQ983Allj5Oj2r8e4vCTH+/eZfGqQnI0SzC5xTL2SapJqUeGCGTjJL7o3Rl/dHzCzWFncrwT
gQUNTcgIJ1oXVKHtqKmqZeAwv0azT5uTlT79c5bt3B/tYPteH2gzSr97Z878piAkAzNc/cI0xMT/
8xusxedn88+5+YptLDRpfN0pEPbruLU+KGo5EDZT92mvPGxcFmvWnlgOBE8c1pv6O6s9aaqjf7Ii
2i1/am+ZUP5uOqy/DYTeStuPIGkjMZRQiltOmUxZheRN2SH3H58f4bxHekNDpMXYCpn5rIVjal/Z
CAcAalMrm3ElmPo/T3+qT9z+7Kbtx0dfvzpDRyNtd80BWVLMqUMruKhLFx3Bo3JXTJtbP+2e5CPE
y1cf1gT2HVUlLS3pHohRp48lDP/7s9ioD7CVfeHF6PtomJLcF/29jrDFDjyWvNf/hMs37NVDrHI3
HkWeZYeoqQAIGhZHQDdhRt6rtB07HIstJVmVk3Eiw7V2y16n4a6skIAvhHOnRQbCqUMi6hyFADSt
iMKg6g4zJF7EE/iP1UcTnX9SUC1Quxtbu7FPRhyZuCL3Q0uSRJf4jcus98b4E/urR//1yil5fS6p
jklToYn+P/zgf3U1i2i+aWR5SeEp/f+vc9wOtN43Keyuipe9TnNp54Tk0dfZifg32VIFTV5yYlvS
ZkBjvoZNXcuqsjcqhOGhcGt61TBx21NL/Tx4ruBTVc6wAiuVdUc/ahEnx1/raHfny8OLyHskLw5W
nn0UltVaVANsr0eUqQBQYlCilxyndLoheYvoUm8YU25ng584lKaxlZ3CIR4dLLHStW3Sc1JD0emx
XOuTg/cXKGZLIMTqiqpoFGLytGZQi4C0Gimbr82MxVyOUJWwu2gqUxmMSCMroogj576Mzt/Tb17x
3i7KG0wwVZmCkoPJjXbzvXLu6STKtxFDuDzo0RaG23jfKx8sZY9gx4dUid2COz53bIACutwUz8ox
Y3QIQ8auuhf2Nn94ox45kCme2cxQfifawWEzhmKVgXkDSC/kmV4LqKy66G4jautQldN2I6eKqlU1
U5JIkux617TErrZqbRaTGF+KoW5OKc7YRQ1JD9H6fU1azdkpzYPxJKI12YncSoBR8I5PoJB/wz28
PME/6AmmIFWKiWYLf2i4D1xY7DMji4FEuEovYgInv2S+ZQIxmgU94GIoeYtaYJ2g8zQo29fvG2O6
oT4mn6SgI37apWhmJAe19QeKOquE/5SMELFN+epFi9Jou+y8btdPgH86v4LrbAiMyw3ikoj3LZ7Y
z30yCSb9Okf2IDCGjdP3m/IBerQOYA1rTHD23gKNghCZa+gryE9M8nsUCCu33ZmY60rgaXUkw2ZD
ExnZIoJ2rkan1b+URHq3BT2WKTh1Bta863pL9QcaIVcJi3ZCAqZb0x71cN5e8Ivg7OJhSjUr4vGn
Ii3iVdvlGaoAkRGSXRHpKqgXsFHvsjoAIwwLmRxLn5ogcyB+frpVc+/Z2ITJvx2dZGtMe31IONEm
US4TiMZbQ0nMMO8OVKg4m8k9vlJDmMDJlbsTOYNJ3JrnR1Ie6kzLuWldevLTCy5+nqDADhnhwGGl
xeVTEaTWMcal3Y2zm9d7/XOM5j2kaVlBvfDnJTtyFAkbGh2Bql1VVzh5SE5EuxSYb7bKU1d1+t1x
Wo4/SkgSjxBrw/iABCa87f3WIN4fn8z4EO0EtsT1T1kOLNH8ZfUkAp0Vumnmc+yXwSs5+66iunIy
1Ee8476APqWdZy+y0+vDMGYIvLt/Ec8otSkJP5wDtvknUUYNRd4Vgr9v0HcCUmrwYAJAZCGOmn1T
r/9lKS2ktnM1zf7RxenStFKEwaX8lOfpfx0s6olAwx0vCOA2hXMyWTs5cCFodUjjnv7/TdZdven/
wC5G81kkDVgJ8ObWuBGzN+cGoYJYUXLFcj5eRYywAHASpjmV5Cpg9iIkmu7MYNCNDSVMEmy/EFnf
qWCjh4MQwbYdYt2gGJfQP2NBp+ux3OfWiWnjUDLeS5RI6dZqZuDqxmozSqF3j2Rlvu89jrXtnj1L
a0NCuCrfiSoV8aEDjU/bLXWYo+SKNjqImln/ZOYsajJ2iGqdhKD+GnKJfqn3J1dt7zoBf5IdKEPI
H6+tIzQaMqd+5BPDg4Iew9MlkD1x6omo0hBfVFIb8dP1rW6Dqqhc618U/MtsOa3svGj0R8/9mJyQ
7yvoijLG37Uc/iUZx5D9KAS2uLFRz3ileV6IQBo+rNaVdItcB/7r4IbTIImdH54avl3iXa/mLJ10
V461TmIWU31XqAr7TTfO+qZMZHY6UoOLdbR4fV9pKJZHlliDF8qkkWpV8HstMsKFZAqzxNm9lU4J
RWexEES3oUBzrdRXsagyfwLTN9HEFzbyTFnRQ7DRzsog0i9+uyEOcC1nSi5snhcamJs8LODH24mQ
/8qcZV+g8S66HkuyDSOyiyML7TEz4hOdGCLQrCXJmNzoEs7jzDdjKCJDgiI7QQrwuqCBthF4lOQy
oR9ysLA+DYB8wWcdEH/HYFHPQhJE4R8D4vd4MIFb18GAxKQIN3Y2Iu+G/UFvQ8tl3tR1LMqrNxNz
stwvLPD2mFjOttGPCz/D/2B3SDJa/kJ7stJgiWgoU1y01NHvjDR9Iy+Y5kJ4pRobRTA4Ti8FzLoO
MkAcjtGwTZaA80GA+9Enl5MoLKWtbM1NJ0uYYAwj8OQZ7SmKcacJF3KPJl7FKs0NAilHcaYN7iU2
bgAcU1QGETfbOh8VImmOSaTW4yt2rhMFAQMwqNyP05GGykrko07scg4N9ju9OAKberYrNLbvLhVQ
15MOK10msM6IYTz5Aj0bops3f1nEWayeg7MKcQjhf+oZOrKbwhtCFYOhl9vvn35ZsXXRoRps7dHM
Qs5TrqWQtXPbQiaYjLaXsvu7B/g8uAbxdQ3sS7CLujXnzULR63ra9vlliouVGLxU7koqobPv2Bhr
ExazusW918yMVL8SaVAkNQXsbNixJAwMHOjQb2lela1pfc7JFhdckrOM+cst8Zc/mqJlm0bYy7p3
+aDOuZvCiOYD0UtsjesA955ob3isYeETBi0y8pd9F+tnNI0bt2UuxZwbr4f51DjaCGzZ1odiAZwI
1LhiH0eDewY9aKy3zTbQN70ZH+ASLA3kHv3alZac6zyzeYZ67oKGEz3z/GsjkEG1oC5eZyusuWks
vZnctAWPT/Alxnq1aIqwdUgNbLvOx9UfYIQClBxoipa/SLRMxO4nHUdeX66YVBMBV+es0Z9jTcev
fd8y66e7GRreUIqK1/ykUvkch76kE//qfepRwGr+i81hdk8rYPtADwanITimnXQPy4kSkNfUW0ic
KGc/NPJj0tDH5QlI1Qfkttt3UbLiGrf6F6aKus9v3oiIchwxz4sTMQNxOUQUmmExKpeuJh8ADcaA
PKFHhSMgNPkvYrwK5hkGP3MnUTCiaLnB5r6wK7OzMCQNfwZmmn00Xzb9OH7z/bNi98aywYoKlVmF
1HcV58BC2upohR7r8WkNateUCS0iFGbPims7LZs3j+hl//6Ocp3pWClyE9vvC8goZREqafN3A/Ef
O7e/VPgeekhE6FjgqnRgTIEww3qDbPVBRBc8OI3WH/oSotZWrJwi5S3tvi+jECAbgePjwf7vZLgV
JRYWJt1OxaW+pcyAzeQX95Nv7ByYmq5KqP2iap9rLSb+SZT5jmdpA8dLztCNw5V79zpQQJImSFnP
AznKu3kNR8p7E4/caF3Q98vMkAEj/C8yeotua/g/o/FWyJUW1xkSfQv9DGBL8YWLNlFHQp/jQe3n
F+IzHXmhkmHCZuA5qnYtJ5vitU+P7KgqTR7w4QNjHKLrflg+gDEoz6ZMvV4XifOI/o2IixGnL3jO
eFZV9sxEaFOP2zHP7AfN+XemYFhksMdNg2wwmPCIvaaqvnEzqUsiVmugmPqnphwluWIx+5hA4DCA
LL1OJErsKXo4WHbN6KLlWXFoAMH2AGGFTP+9Udwttu40ydo/tenad0V4AEqogND8CvPtoyaII5cK
AV430EqX9jbBR3u7Qj2gwcsq9FWc1Jbl3FOp+VL6issA52ipOnd5ofC7J5QO1ecuCmkpLxQhN5Gb
QtnHXcg3mOm9Vhg9h0D9N34TuFTh4euj4/Qor1xUxJTzWJSd1NxxjVGmO3950jKtBpq7iEUZgNOb
MbVJ7DdrOJ6lCU3XsYBuepLDmE4YsrMZFQWm7IIOznzMTXO9g3AOLjXCm0MANz84H+1rqCaOcLgO
fmUxSD4U8N2m1rgP0LtkqSrBWSr6lo0x7uNTJHyzqebOt2uvDDauljyjVofZvaMneN10jVZAsZ9W
rz2vnlZdFn0iqBPZ/ZoQQP7QoicNaOc5e8bAW+qzOX0/u2hH0Yl7WUF3uJFRBxDp4pSRukiFX7l1
w3dCi/1gP/Z7VzpnC3CFmYkB1x4JS8/MWNvsMDMx6jbL+oP4Yd+/fNPMoc4yI2o3fwiBVCNeD0y/
vnQTHDokfG9GrJZHLwn1s3CZmRry4RaH66tHBE4Gqw4DrkCB0rInf5GRYxL1ElUsGGgNjDOWNKRo
xCFtwV4vx0UkknZjiikvwUAH0uUbsIKXuM6rns+q28+UFRbxWwdL+CBIn76jdMFxYOJt55f+OPsI
OEx0HYEJTz4eGMLl74u9pEmYsDO00QL63y6oJEA041ZytYG+4uRD7KT+FV+++MRFmkbzfThvuWLj
jn5Ndaf8CLFxgfI4nIgJKG6+jruvcMP5657aYr1iO7xkOlQyvQ8lm1RGKxfCVepeMImSvDNrND9F
tCBKJKHDtMcETG3HsbiqdnEUNFZo1DJVYGIhEAIS+wL8NK8bdMBVSmAyjfrhdqk4nRW7ixG0rK2t
Ol2U9zg/hUCABj/fKvdGb0LBhpzIdP3sMep2BEpJljYwN9c343ZBDDX2MbINkqSR0rHr8eu9HXPT
H+gkvOlAa+MtxxonL93zMyPSLmhBXAA19ijJYax+KFF0NOvcHnPL806aNsXeIqRKdT3aK+aHhEpz
IkXF1R/F5qi0DXIvmiDUuDQcFkb8uf3VKpRsv/OpzaLMCCo2qIE0EZkWK0cvHiyft5+y6U+1Nh+E
t/g71qhveXajxglQV5W7wvUSM5WjyEGD8Q2qo+12bXexfe2LoLIKlL40xeWe7D99H1Pwt98+iSxE
GFwm+z5Y/m5SDvCB4tuCeTHh1QmKD8T+Q4sItBNzkXIiZwgO2WYo75sxP+A9Kq06u7S0oaoF4TYX
TdT4mlsgrbKWxspiVj4nummJ4MvvlMXqr5NjIju8z6IQNevMMN9XhVrWRkhEu8ddfE5M0uAVVu1w
Z70ibERpG508hC6SktwMZgb77gy2JrsbtkFl1pkI00mVlQgcAGrXWEMMfR/Ge9FkHLpVyFkUpkQZ
mSiLJMSXl8Q2QX0WmB6NX8MJvdlB8c4rGDzjW5TB/YzCdlRajMJ3AiagGLUDsFBRtuYicxjfpKhi
nFFmWEoaQ0GTxFWpZqsWxyBFh2HwDAw/wRaAF3a6epLkExn5QXSMq/t7pojsq//qsINdCGSzynwL
oOO2Z6P0RThG+tBguFmYH1Yq9xpehuH5dYicDVZ8uLrSQq6/shIlJBN8pJi/HVBPkc1UN6Km5aGH
IuRBOWucIU685Un43ASxm4qDZy1NUiPX4MAHQEiQLyZ4iwswIt9rbHc8U5OwH4ozqeAwc0dg/qvo
rC0ABgK9N0MvAKQMGYH/rbY8YPfigX5Xlr/e6d0gCNknP3gXApXCNcDodFdegnj/6gemJUfUXcQV
lk5tKUrQznw6cwbt+MAG1dyAw8sQ4uqLkFM1/nC+nhWXLb3fcxKCoUn8lxtWILdTF5d3qBHRhsP8
kDdB7RVAAjfopoUo4/Capf9RPCHWB6XLmT917nHBpSO8N5+78dxhqMiY7acogJKmsK5QssPmeXxL
ZkuZwmhZ6OGbXEPnk2hqKhqWwkCcr9Xv57x1y6F+hXvoyynFI/uYJwYNezBEw5vaAllEDePaza49
JxS02llJGNSUoXaGlnImm6dWFua3J/aq6IfBn0qDKaY15a3w1TKpKos3SP9TXlRTO4qlLf/DrDLn
QZpJzDm2cXS0gGONnRgjjPGigiNn64GKxD1VocfI8tK1pnIeKsYDxVueCaixfeACe9KfwACve73q
3BaU0H5e63Hpzwa4f9cBBg/5MMDCz7Xkz2g3KZP/BaE3qnbCVVBF6sddpH8fbNa8EwY3ujJtaLRk
LPLBmZCitKCGxSt4MrIoDuALJ73JVe+Belcey1PG9rU8gVeG9txJKlVMFPFXoSulmMBir5Yyju0t
Jz/jBofxIzWLRzoTDS4YvTtPanExfAaJm7Als4zFAFkSYBCk0pg64VRXzr2H2Wom9OzCkCjbqE7z
u37/r3IvG4ric9qIc0LbCVBO/SEQ3u+uUTHTYSxItR7nRqPCxB1OwTBRdOkeDLTgJd3o5Qhhdmm5
aySFcxvFT+ZWdJdCXSu77VlwL4xNr7b2or4LA10829X6JvtQdDGJXnj++KeSUDCVWUrBwqTWwLaK
ivB1MfMfXnHGOBw1QXDxO1r1M2xXdzFH4G6OK9BP6ZkRsV/MAFfEOnuKOj396Re1vYLph4CF8erm
F0VkZceRa4lVQ4v6dA8ztSQpTtG6KEbGM7qbdWDnypx+ZZjpxX08KLY0dWAkuZ74ipv3F3W2PMJM
eNOZNhf55b4FY6boeXBezLVjnV5j6kvuayAL2X6aYIU56QMsDuJBtcOgEIN+X7CRUV/qv2A7h4U1
XkCsF48SZtrNrupbuSNEJN7FQS4cRZARLLsrImRx9hOg8neKaMbXPDZqlnj2flpMODlqlBYjNYbS
jh7sBAK7FVbFoevCNvXJg6FZB6kylXmZYIq2Uk7i+/dtfuphsPsAJVyoc/G9kPsqKrBH4sSEFOB8
Nm4DZmTK+w9HYYBpnlxGMEqWJKvJC230GH4CRnUr6Cx3xhV/ySrlI0VSLoMBb/lBL6dgmRkCyk4P
tUJESyd8H64haJK0/WC7sorqiJcJ9v/sVk48agIIrZ0Pwii8/rWO6Hde3TP6JjkNrEokZkHSe5bv
9B+n96t8EhWLzD/Qocq6iBRzqUWsR8mKj/kPgKTl7pJ00oshQR2ifIg58VI3v+KjsrV+azy7gDUE
V43cNXcj99+0f786dXaCSbw0c4mla7ZCaO/UERX0bZdMbIbNh3n5CyFiRNNGWaM3XG5xFcUpjarW
oD1Csj8L0ekjLQggBNzMtyxeoIbUe8s67363tv5LODYMAWSNCzNfjd3VdPnoQ+Qwjl29kuuuYdVL
V7Tqk9t4gCjrJ4GmVl270H94y0PpSPd17gDz+2xrM6FJ605EJ43A8ul9T9F4OL84Vqln/b/ARWYQ
j33ZiUaT2s9pCqcbmEY6yT0K7mgmEIbGiu6MCJm75ZA07gvBVn/C05ZDg8fupKGG9kPIFTwaLL6Z
Ezp/6AWKRdwa7b3/nkuida7nYGUVtLDhh8VK6qe04+4dOd6IM3jhw3obwNyzbkpsNFFFZIPB7BQk
osvXluMqQRU7TJI7wDIpFT+4c78971Eh9cqSYKMvQxVSgbXBFv12BuHlFG0cHElx27b3+4fOvo3W
UaFqkmafr+twO/VoTKkHUglF5hSr/Y2phqjbaJFTyx64s3sXIGm0KB2HAmj6xSK1o4Yw/xfTvJbU
b8GriXPWqn+0InI90ynPLog5K+w9bf5eshWJivuYlkgifo7koC+WHQ8AUKbGuhXMyu3Z8wNBJoNw
e3GplqEGgH1PEhCN/M3k5xdSboDXp1FeDR/Ms+36Vzidx4bHEYZ6oJmtW0OATOxQnbhnA3s9LmI3
Qkb1ZxUy1yJaFQa7sEeCANvCszP6nsoffn7QzVH8uKbIBXbr2wxP4XaHEEd8shHaT72taB01VrCS
g/ZC9jXWTFyW8vCvRLFszGay5WZfxl7c1tbxCgyvHQmNcfjFE4RWAXU5hpjUOx/QhmR9sr5HBurN
qw3kvknepCwWrkP2XlLHHZUirZcbeujiRBE6g1gzAEdDYRz45cSLa1gwuW66vIAUxS0ODXUu8wAT
41JQGAInxWG5l/MdZTRDOy45n4v51+/kdNfjTjYH4ntz4VB39XCZvvy04d0RR+YOe4SThPSVGUJ+
bVqhYlg0x+qs9l4G2r1QYaP1WbwX4vztPwxdNi/GXvgXnn+NzZDYzXAWLqjQa3I5eCUkeLyWIGI2
L072mc1IVBMAG4Yefu8VtrJ8AwYy7c+CceewRGvlA/JrnOhNzU11PU7OxopMguHAPIT5plXjVPss
9KLcJ1T/WE0k5R/yLCOiTokbvoFQ+cdHipaf2TJGGOGxEHzAw8BDxQbvzNcpq5iZnKw+DF+zjDUu
TufaQetGEejVB0n+wGupeeLwAGJ9i1DCa4b7lbuUeXt0K1Equh98Sx8N5B8rEtN6LyZc1cYR6/hW
vIn7mIDhFhx0quQ5rF6Sk688XEHy+EBDl5CPkDgGbIh3RZCNRI2mtUDjxYL91vw945N7oozheYit
b2GXIhFKJ/reFoilkrHp9HzRANYeLMGuqtDfYfEpn2iTZPQJzymwGdan5MtXqzE00iBrmRrqFwh0
IRG9aRlDGFU1jZN99vVyoSoz6lv9XK2yD0R7LjCooXGXUZdttb4jdrIJXL/2jKA4T5dsVqNJBS/f
x1g+iARUex04YlQFJzUF9DuO7h2DkkIVP0rKNZZqM9Y83G8KVbf0uCRPgtdECffKnmlq7Hc43/mg
oBCKwH/B+XEuK7EWSY2mtQAPtNKpkpRtsLuYrzL5Mqca+0v8bmS9OgiO3kihHWdnmSa8vynNVdT8
FWMipsbf4ZbrSrs75Ge1CBd/tSyNRQvu8l60kO2rLey7i6nwcUxC7LFsXIhHivjOhtTMBXAqa+7w
4Yf/N12T3ijlRvFywuyDnM5HsJnnP7PsNBZSAQ8OFjB+Qc/97Jo1yogf/sbgVsrf6eiq8EcUOqpO
mLglJMT5r3sC68ZsWjcFtVhhKPegYi7TrYlm3D5MCzTrfGbN7ODu0JmUZNzjHxzkkOZi3P4eWY71
uvUJOFK/u+VbHZIZrh1XKOoUD5Wr3nmpNjN/XCKBdt4n42xior8qyJNOmVssZSR42+vraPb6G/8K
lyk5QKqvyNbcjXsSvNnvqvLuNmHPuxcww1ATyRS5Vfa8VA/5BAiAI/3YLwlji/sXIJ8TRtzXBQvL
WBH5K1LvIicrELKB8hk/1Z+S1NGOkyme9sBcriHGEh6T/s9O9zVLLl+U16YgpEa4n42ESDeohmFM
1IDtJZODvhKwzF35YhCXdNdkLemqNow2lhDd4OYb/saN0E95PKpZpHIu06baXR6BFfw585MIeZP3
K03H5MgwafM0kUiwmDDKR1Zl/FwtmuXJZmaBRe3MDUFj4ptWu538oCm8GdQ6A/VQSJfRdG7O9E0I
I+09hfS5OTHg/VbG3LkOymBNRG+xwATUqosZwI+8G5GIld3cneGXNtgwvzL03pto/JHaQIE1WFsr
60yJ/JrlcXEWyjBd2jYkhROa23EqQ0i8yudzCeQfHsT2fkhr8RKTjquIYnoYWvBjWhfRUpJ0Md2r
z0ez+oMR7QPkg/ma9i2nnG+m3E//hDLocp5nGIi6sXwMV0ToQvpJn4+zkQ3wBOYbDvFCnkbvjiXC
d1MO2A36A2PV20ydsy/sXDPXsQL3798LRPlUC83IcQZHdr5towjBC8PQfcuTY5ltCC3gipCmFDAJ
6cyiT3fA1psw/OINZse+WcCU1XalOrpVEsXZYnVEzkl+Cna72B8TYHHWGDKSqskYbjqegbdWI6vo
K50XGTZ9BaVzMkmPhX6HPckbVfLc53XTVa/6ErrPaPzPvzQNYHLRzkW61n949bjXiv5oozoKTEXr
y0vK5tBqnQeujBxp3Aaii/JLE2iwxhLw8A1M+ddD/moX4AtjcXKMszPfr3o+HnoXHBlxfao3huO/
wRc7MFVyvXBMTlC9WDQMW0d4g35B8gcRau4B0UnF5YyVYoBHspq2QxhG+Y0LlH5qdpxpY00J4lDz
DNFdnRZBtURMT25PP0hlkmTRs6dpDvkGjQfElxAUWjc9Ax9B3hxc4rjt7ujNHHQu2RG+Fq57JzrP
UBYr5VGkEBUQDq+vPz3VuTgako+rKguoUJE1nIs8myjK4KGfgt3TFuZaFHVVkbA/I+/03jxrqXQ3
Z3j2+d+1HQI/HZH8SOon5ZKzLyvEnlCjLnc6XuRU1NKQ/DNuEjC2QVKryG2P/noYeT0syiBvaDzR
F9vHp8YawCgIj+FPTqHBB6A48POluaz81zDs5GtdajEZtvBOauHAG80qPFxKjrIWJkk5NPu8VSOZ
mVSxJs736YMcVwIJh5gtNlyTDdy2wQ5eJSyjb7H3CA4ZX2lOEJuTWxAZfdoyQFcQulaH8Te9rfXg
GdxGxmmagtGUh2TOSy8dktZisDKL5PRpUj+NjYHGSUYg81yZkBUPhHUSsIkemL1wLvqfp26M4LO0
9TZC53TYCLusoMZEi5zTfRDN2tWSdAfc6hoBOLGRQHZ7o7LnHgPQV0awumTEsySVsQUI+kKiI8FJ
LQkkDIuSL0Ik/pAEYg6N30/j5L1DT0i4fkdQfYQ/SIjAWhZvZgsvGr0cNlA3TDRZ3f8jnvBpG/v1
T+GL+lf9jEzPE33jktxr1JjKT2dBBTIj0tvMvHd9Ow+NV2zX4E2R65Xcn9ESPCZ9TWywYK3iUqSc
FeZfv+ZNybaUpcW3CguCwglK/vMjLNerqYpl9oQ5+cWDp3XWeJxJTh1iEf5f5NEr2Q2mB4op21vr
xkAtnCoR8Liqg7WI3Xy/RCov56HIALZZopkR761zm4ijgoYI2WR+5jtzf4ZegTdnkOLrYfx0tSXN
ZgLqIlMsJyf6605tVCbtzk1PV81KIY3wOXUT3uYVhDqD2nh0TcJC1WTz6kHxH9dWtG4WmjSUCS6f
Fjom3NxaeyIkhdkGMuBlm+LUfe0MZuewjKMjS9UA6YRpAgyY4FPFIeWXambUPpTs7C171DBi+MsQ
TZckPwyt/KUGkd2R3uJRQ61fmRgMjnJihTy/E2cLNp2QvIhPcMWkFzIHBaZCGBbdNAkskKGPLH0a
pRlcbJXqrB99LZREA5BaDNIrQDJpe0hCuWXPSSFj0dZDUoGiSQ9s4wucWZzZwq4dQVis7yFDIVN5
cjQEHjVoDDqNfMjlA9p3msx7IwqaBwrfcCAhx+CcLUaOM2+J/A8+qGR6eVm88qSHSja0lrRZ19fK
txX3G69DhFZAvo1I6TOuPAk8jCMRUUXfdTuM4108pFF6N156bNEXg4wpZa6pXur2cn/v5nqTzvQB
7XmhyoJSzFot7GvtRKNw/vtpDFOTuMdQFfCjtewNIWOAAtk64OI7jlSBaAven/5fkR8tykeBQ4YJ
sRpvfMgdH7gsEb8y5N/QorVxA5TUcYl+9lRFoJ14qYLiau/5PGZwLNADALqAwm7X37zoZM8VyLSc
QMSoQAAFEqL12BPBulDuzs1auuBRSi8Rdv3opKTWLqqtmhkpWmhqn0qTPm9TYPG3kjA6vc1RFaFD
Q05FdWwb79aBIkD6Fdkx+VuWi1Kdc7nGO460xWHNGTxfK8VkRj6MTadeGHK2VLovoxxfJr78YqQ2
bn2i3ecluR48KQE4yLKJ8eupQHQL75icsVhyVZPNxvWaZT23Fg0480ufstfbLQrf4HPxPkJfKrsf
magtDoJvWrbB446cNMzxmp5+DVYooJdd/gG4RNo+iF2jJGy4jm7TXeWps5CNpY4s8o/pJeayiat7
rYgvl9L9D7+XgvWR1GmlLJMVcmf8Ojp7+D5kF/cu7rsYaAQ2aK9h/pVDy2yhFXiYLSpKfp2wLU+J
Yb+NpZ3ip5RAsvQ/0guQ9CQ4ajj9K1+7IzWW6ksmySHoXxjDNeugkrCiUJPhRq/Ifpd/pPZ+co51
Quda9lVu/6EnguLSzhOTOUj1D64uASJeZ394JQgxEaeN5X+6A4FytXayM4wr4SzDJMf1Pj/ur3Yy
UefuajP0Q70cVFkJRm+Y6LddXZz/K8qd8nb8QVPKC36hVT2a8g/hvN63dxSk4aCKquVvFIr8koVF
ntrO8WB1Z9lXpNo9Fe9/PxHkSzzrKG5XrEWAyguMaQ30l8Jw2wbj5SqY0koaJ5tlQo9LbXgj2ikf
vZviPNWoBCSaC6D8+wEiY+l93nA2XfJ8Xy3ECqvuzFGu8rPrdhKHLdDqkhJECYiAtaevxrsTIWiF
1LpRV5e+hWzk+r2sASlN2A8GFuMwbI4ZATwOHtxgJ6USrNnIpn0PSsXodNszrvQj+MJe/EYFqD2Z
JlS/5iqEs773fQg1Ps1VbHcDzGp0Wd96/qUGrvE0lQik1HTX6ZyvIAHY7Zp/CRygaXhleHG8VYQM
60kwLTRs+Q1I3/i44wBs0GQk1JVOk+stB4r7buaLxY/hWfZLLUA6QE3iUb2JbvmTMo/QOJIl+8xj
WI5PacLPemDa68OTBILZaHV8pk/Lm/2xo1gtC0ER5+yUY4wHVFmyYr2iB2weDsaQVHPi6QbFOqRv
TAPZhAWZ2l5SZxDfhIKAnyjjr2mstKdDN5LeuBnrLQzhfAMWumxrGIepGQGLAmbWJd5dkablbT0L
pLIDqLOAEhpFRj7hy5c1v51ML0mlFum0AF3/nJUOl4x1mnpOdNgQ5inER8bKnLXDLCTui2IMlCgL
rFrLFIY8C/tyaRra8CkycruzsPyrDfP/U5x9BXATf1vjNftPdQ9rGQaTyvaX8Ce0sAKcHZQgQ+oA
mhWzV1wfiGcDTaOqD014aKfjhBnFbLqe+9QlMBou1eiWmqSXkPSej+KSZuVgZlPgsUp7EEB7x/zE
a+ijlxQoZBDqZYh87om2xrYNBw5Q4ZRQ6ZiNyR3WyTwlBR5OmE7uYHYVU2O5NUjqDP1RdcCGY/81
Fj3gMUUtlYL5jHBoxqGjED1y+00kHxZqlgV2r/Ohfihj8KwKyS8jBWH/5KPM/cPpZXGQBZNH9k7q
2hNhKsLEPijeDnyhdnM2ncxNB6h7vxQIOmyeoO7bm8O/tKMdyrSO7DsSk1/cfoEsFQiOo7an3ri8
5sQp8GAnRxDEBcoqHHwiJCtqVtAwIvWbiOWzTVTFCDkDCbNjYEKWhkEd3f7bpRHbRS8YjUtfu4CT
MZTh0XgcuArMR4c9sMxVFJ9QwTupmVcvv5yP34LK+Y3lGpfInKjf5F/n1wnCWyQ8DLe2rxQdwVbD
6gih/RcHTiUvjwI9thgrYH0uwCAHubufbdDLJFdr9+CjukSHGDfVtyVuYMhTYalwSOpCduZ1R+/B
xBAdLnx2YC2/N6JrbRgC+iYAotBIKmG2LFBg1/M/bdXdEDwveoOzGrCqb6WYr93XaMTr7MPk8xGr
rbqYSQiO/drGLBuwyo1csPmwXjbt5wXVhtv7nA906D6ZJoAL5745qZi0dxzltyO3i8PuKKDEJ3qy
+mMDl+rVlG4RbP/Dp7Z55MSHcqV38sKnZuLifzQ4Do3dIkfc54XPa39NzX5IcuKl6l4G3+jX9GKY
sYdeoCH4TKZkmYJ9OizWGCR64BTwprSYsAWSyKVfXO1qLRI3v0u+Q5KlGvb4pQJ2oEkxgzr9MpKl
k4KoocDof4TncW3lk12X3arwIyAtzKjjNsj3ZYoDd2e4VIIIL62WFs1hiXq4CwnUKUEiSlyWbgjs
3j2uYQQqwBNTIW2zAkkSdT8CWgPQGO5idP054wdbz4Zx97RDUi7IdxSciv0ogMsFHUhQOyDON9xZ
5VjyAdi6BtxdxP2/e3XryVxCfxKuVCRYnCNcJuW/mdDmyk0S2PVyLno0sdPS50Wh1EuRGdnzxK8S
0OutYkVj8MVE2MzLY8RcrOWTflydQothWiMLMSvPQWZRVz6UE9V1tjEwSUP9qu7uWOLxXRfAQHqb
G+/n4+XK3AIH7SHOc6gFPVAFnbz6b7bbRx0+lyEEi/5//tZ5UTdbR2d9AhdLaeHWDdXE5tuXvo1/
Eez9i2wYIHLq4KNtETZT+Yj5JrD+7SfgfeRYrYJXp8B6bsS+avxuLM6WyskF7jpkDc4Ubc90lUL0
yXj53BMs5ucijAQRpshMujczxJJM8Gzwlq9i5Y28hgvClRYoJvc0zBsVD6Cq4Zh2AcuPEmdi4vVk
HGXJea91tIXdph/0i//vjZ47GexxLuEotW8XwEBbcOlw3n+hk3NKiwCcGXW+fzLUHqBUOg/Wi4mS
sJu6Hvf+iR/JUFoN7iiIsfkKLcbw2ybO7wu6UMtz3aUwpAzeJu4cQMAzfgw9d1pgxqrFbxnhGqj8
Phn+XwjSNXCiDqyNUfOuuoFNW40065fIBGHguw1QoNBgT5z7L5hUv/mReyXkJtfl8ZsquzsL4RwH
tn9LzEgmhnmsn/aDGoVyrYI4247ZmURh0FcPdOwAJIbw+TNJ6cFz7v0rXSC5gqOMF7VFMDhhSEWE
PyB6/+sq4gJ63Am1hDD3A4J7fRXs9ZtjUVI3vco1FV0wXAdmktsQIUwWwTwY+aV/4bjByCb4LTCQ
YcF7y0BkMKW4zsGXRAkg0e66UOhWFUmygYveSrxj3ymBD72Y2nfxzPmUZZqGKHutMXe8MxmbB+rW
OMlLPRMVKB9013zopJlWGjHQ+6rEwfwrsKNaOwYmLh0D6MmRzvdRuyVxIHzNqzGf0NnmWNFNUHyP
zxoMbrH9YdI/Fa+rDZW9xFRUTwHC6v9SIXOuA7yOnuunOkP2fHxEa3Z4/PUFWMAjzOEfnx0Nx1rH
bvS/cRMwtvM1ZX2ET8MRttyTkMaOTvQbgrFlW33EvV7gJhGULieoCPhv+df1y/RdvvCY+/UlqKnK
Ey9CWl7IkTO4o6dxFP4j7hyhR1vc+CEB97XLH31hKE3QTxOsgiFRBL3XnrnHI03Bqqp2DzrANwoU
XoNMeiIomzjwKnyaolJ60q04fLdBFXKMh96c9sCPFP8P5OxAkzvmFIBcQnAOYRfEazlcQrNgh5hH
MHYPb8aoMDLaiBlzI7s/ripDgM6B4QNDWI67CxPY7i2wTdH0I5DEfwq50rOH4TF9LsbuXPQIgJ9z
Kpqy+9RCpM5SX7esCUA1S4lGG6m3ESEiBJVnd04sHXTtXPwHSMawGPaT+c2s7DlR4gpVAit8QKn0
tSY8tgGKKE50uMLEy6HpRHPavhMa8M674gMoOGzmsXNIXY4O7EQ/DlsavMmd/Kve3JjmTRPP1Hvh
nF64ao3JwZASa2NUXkGSG5fI6tNkdHcW4S7rLGG6H50C9/yQ0CiwQsfRUsiSFcaporuG1PilGB1H
2w94Pp+WQauxbw6Hgn5pE1Uvht07mchoWHM9OBn95qMH+MwRHHK3Q6YRbAWyqOjWG93t6xRQZFUu
rWv+t1fCpn0AtZz4MPsK4wQpQKfNLIZlMYa0oXK47HoAgMhTLjD4383F5SWrFNADK/AOTRagZGYZ
f1uuO9NlHcTs2Xwd4x2LrUCkS0UsW5e1tEBO8mPUKuutM4mh0XDS4JsOrYl53tVI4bQiAhXscWV4
kV30BW5xohQlO0IRhqZY9tlNVmHS7UbQiXi2ipeqyc7o+DZAVpNQl1nPbogzJu2y2nNSlFnfdmmM
CHsX5WSbkNsiwEkE07L/nn+nftlGMWswqAS7iuo49LzlEFoSW1gsb4GBfxwYittglPrwJeX6aeyw
d3afaJwaRcZebFmRvizIt9vQh2GRfH+ufrjCgmExldFRzSD0CDpGboiriEbW8imxEskZbUrWRixv
MfUEAofa6Tm+AtoBw7h4zoL0jQW+GSVBq4LRv8zwxarfsn5FLfpeBFkbUcOVK8w29AKDqBV3B2eB
OZcAbME0xQ/rajQgS0kCWO2T9ibfS0J1tOYMnRSX8lpR3ESpQzUL2ipqqbmcwh2fkHwqtDLqYMlb
GYMWW6jqQwJ02tSBnIwN3zYQXAX+QEjQBumKqn+2juja56Kloz12jKhpFLzx26EojmC/8ZJGh1U6
xH2F+/qESJjej9+WqY9Lg+VOkaoPppEKGxGl6aFIOyO/Mfyx2SrjoczYe+KHwSFxPsem4acD6cA1
zzVfodHu2jbFChIwy1ONEn3Px0T/k5NBmVVgHmIIxircj6dprKZa53TowhkDO/6QXTGd86/KvNbx
jTOauLiJWDHKJ7gQzUYLEDISdumuVm7XkyNSL9E1TA4ckdJmZDfsJS5w2TX+X+rXHZlupHBTstoj
H/SyxnyVMtUrLbT3fr8LCjZGt1mbU4rVLPICbD/Y94OAcy9N5DbOOF68sYIMjQ/FiEF0JUPdo+AO
C0TGut3M5zdQOPXwUp7F1OGSJrZHTrXmM2GCKtxxU/Qw2MQhtjDVCXqjRzxk2O4AvhSHv2DruSHR
p820PjyHF9WgjNOIKBvU/HfzGvMNNSafO36PsdE8myL0ySC9h9QKjYd75d1o0NQ1MGa7KkqRJpkT
Q1TNdOxkLR8gkvlXK+0yTsnEbqBxy/QlOMOwGKUoCcMFj8z46RAd90X7NVlmuB2We8TuUtFb16Dp
SNq4+0OJhu4yfV3buJFyw5s/1yKxoIK0Ir9rEpRGvhpXgM1SN0dOulpZMNbjFqFYzA0hD0lsyk0a
MotNmhI1dNL00FgN/CaVH1Is2ZO10WYTrKxi8Rq1hi/1DUqetBxk5tvsTu4sndwxLpd5/Pu041Co
b/D/VVPD2uEaSfaeaOjFQjxaqGZRB3eAbdc50MDE1sWCgj8/iUtQXrSCVP9QPAqyGIQESk8J1JmD
ImhZ3aBoWx2ZPI/qbqllXTuF1eU5qsq52VK8IihZtsjFofXcoM+/VIL39E0sOUcCrVMU8Gvz1uXy
0abph0B2XOU9Bjb5bNDVYXSa4vnG0bTRVh5D5w6OjOpgr9qm12btcw0zlqAO71TwBAgG8D5HMEhZ
QJwafPHuEaU91MxUAAxkCGFzGN5iGL+2w/BavqYQ5tALzZY2I9SnWgaffJ297gQL52gouFuazU5B
2aZRBgf4R2SqGGIgoCtHraUvptPEO5zAcBwys8ClB27dmPiqZ+3D7sDk5GHbq6LvoLzWLYybIvos
4apYw2xeB0oMKTomUTZAM+U4x8YbECjTxd8EGi341R+1NHSMCmvZ2bxV1C/pSELHKtm0EokCqlpQ
9ga2L/BQfeSQcst+AaJPUGUBz5ErX7zLN3hMmwUu6pFZZ7WTPTyvQTjA5CFwFlGAD4B2Q4AZbH4q
he3pN9rqmIm4mWv9iz3ahy/vMNd/hyedq+suERxiuqa8O8qKR1Vb0yR7bu0+BfcV4ARC4xJICaxA
/gMeP/DsozcPDMnjW1w7EWNDg+n+MUfrj6kq8hTUzOaAL0gorfuju0nm1UHM2Thh7HPz+/MW/SyK
UMyKd4Aoynaa1b9fSKuo3CkFnoTN+OHf8epwMe+jB0Pnn47X8h3sXIz1gUMfJP7mvrIAkrMhI4iQ
BWVtcY0EjC7r+o2qqxu5EI7EQXjLPQQX/hAOjTWukqQCsCA8GqVOPrPRwYYuslCDspEAPODUk5Jx
7VKLlOgM8k2Gd4TSOYlM3Yr7aAlydRGAl0r87hTogMu8qnjLm3WSQB5otuaOuhoz/0G73nDHDQzy
RcsQfwyO3yGP7H371ZZoBdQ6cxa/Yzd/XBxv/az8Clua7z7Zvl/LjxVaseMRKPwJp2SNNxBiFLyP
ZfEXv1UdRvC+U2oi9KCBzNfxuqapWfNGQ1+sYoHBMN03k+g4gOrtw8St7C7K0T7Ve4VZI0T1fAHl
OFUWHj6UIxOGGbuD7r/SL4ygjHkO+RDupHM0PV1ehF1Ps4ucGiZ4N2q25N4tkzoGg3dsDIIl0vYf
rt3z5NEVY5wZ4wR/AjMxw3tLg8gVPOdb6ZGLlrce9J3pWona0ovepA6N+TqCQPpx1uOHWSbT0+VP
DCBIjiP3lLc9/39v8+NxyP8b+X4B0aXxFeD/jakTsJIZeB1m5QjkLzZ41HK8Tnw0mZ4Ynav7SzTy
V3KTOs0Ax/kFYxk66mai7owjISB21u7CSR6FrdfSM0cUouoyR0Ks7ZpJt7LVL1ojScsv5w/T8e7u
tIeCuvUu9b2fyEzC0wELI6eyNLbZENIyBETQUDDrQRGnsUrP7TzWXyfVED1pyNOGwwJq0X7205aA
Jx5hlrGQWvIEbPGnCgx58xG8eojeHvxW0SvH2UP1uiyQqC4YKHcKGCX/mWv/qD4jjpaj/p7i9O5O
4X7iw1oluoJvdWyzaOpQvDTeMKQ6Ob2UUM3o8sIWXf/CqwxgJEYyn6tUFP+EhTRtjKJPIq5J3qqP
VMPw/VaAjTxytVkxwbkyaY/FeZ17FdTBOewGCrxRZQtbPh3P9jp/1JLRFSpDHva/54OL3PAyWBog
YvE9GFhqi1qLhwaRqjpyfYDku/7nbrjm4clD45RU/6pDlqkoxUl9YAlBzAsRl5q9kVKp2R8i0YJm
dunlwckX3Y3EDACmoxD65RGylGyZxWXXfYJAa+Kd9v8CGDVYa9EcX183cyqpIZWZNFIQA2b5yYxL
tWrMmiFVBs7jZHzumvNx8L+AheSdaNo/P3ePr3oQOUj/tU0GCpCHhwJ0u06D84OsHy2/vT3t/JCD
eV+OkSK5U+FjAUZ3SXDUXak1f+WhEZsLKX3kzEyXG0DSXONWesk8MeTmN6RZI0PEurnjWLVcIIAn
sbVi+890YBH5kPUo5JAiVvu71xJbFlhu8+8wM2bFJG6Vf0Nx28ZJzz8By1lyxUFIB11vAeJaRjvk
NS5bt6sKddrnmqY/i5P5WUxytY4VXNDM3Vk/kCvnW59oa7ULNmIZ2AeWjuvzCpbozhboPIcAHYJl
Q16dzL3LLtxR2fnlTYyXS3AKDRJz3+i+7EMes9mQDo/8WuQp81b1EXKJbw8IWW07v60a6PUzzm05
fyUdOEq6yogjAOMM0U3ZB4gsTQBpSQ/oC814xrswrVyJZ2cb8IlNkVqzp1+rXv+cFcRtTWvnMj4G
GN14KY3lvn0qMVaAgmWqd3oI8UIU2s9k+Mjpa2UO2rh7yYnTMjlwMWmo/VLgKoGwJlRSJnMIHoVq
pv9e+CSry5ZOzP6wCLiyKbFVIKCn6G717jfC4mhm8VwR9yGqHzEhEbohVDiwGz+mbFbJ96JEBFA8
1KmbNX8oHvU9rylUMp7TivZVaep3/y760wC5AFFAtz0X0RLkrH6O6js/tviMHeQDoblf1Cy6XLuP
DuI80LCBnL3YQF3bhDwHrkdM2sTslWp1gpog0y47Eegq+EZyvtOMM/ukon1mRqHl4DeUSjO8oHkQ
ZCCPyL2FoiCVjthamgdNGVsnxV98T+NTN72P9eS8id4JjDTdH/+wz7U+AL9ph1+tG6xiY0y9YvDP
HsYl2OliGWLAm6zE5hxIeRrv3dwmHu9hHifFhuaUCMoFa+Oe7TENcQ3CDGvVEtFflvtynnZpSuLX
rnZ9MZ+JXY6gSYhjDpQDZaGcnEbsKZqiCbOlAhpU+S8ovK2W50jBzm3K8IPW2IZktwOOgg6mwutt
rIRs6+r5bWLhvbHDEH1IoCnS1lck53tuXy5hWzgo1WAyeW99fNH8l15CmRL+magLHKmItvh5zJ/8
vtZ7Pg8Sc28+K0XWsmy+pfDpzGEDPxPU5NK2xdLDf/VtrFA6tPNDCQJs1lqNfVsF46MJAv0WtlVK
NS83GaEuI3pJXrZ7MX9UdgQ7KwL/wqYqAjXH2SWlesbX3wwYVU0qIhrYxOn/tAm31K66h9aSx3yb
7SGHB3qiM/mmwuFSD2JQn7eUJagDBzogtdGoGCeCx+l3jB/NBzqYlmJXs9g5lqp3Hkf/AG2D1Urv
Q6MZv8Tw8fevYFLnU3TcCnsG2CcEYQilZYw1KwT3cipApokIN6QAfNWJWgXKHsYtQWSzQqduV+Hi
KPyaFPfrT3tl/p0I6AygbO4ADI3TpTyFs/TnYBLxqFKF04gfH9izx1dg6+crLJV/gz8Xbr0mWz7b
hTUmHovxRWk/qdbbyFY5UbYai4ncNDwSCnqR28+N2MiMVY0g+dK7P2Gfw1r4Q2nSApXwxuq327s/
dAxK1tnDgZ7AqUJ0jMsQXmTiETANFgdvtoXtk3WJWvZrPrpV4+GST7enuJirVz811ZrRVN1qvt6S
7ltPIV/6UbPev2Kwr5g4pI+5W6184fE5NCOGXa+XSgJVq+R03dI+wvNj44Ks2Y9K50ZJk4OOD0O1
aC9jJvnE8Dqsw0uhJyt/Xe27+DD40xEfRwOEuO5LoYk0ylgIkb0UutF8VR//VgK2pLxmd+SW64GZ
dYF7UIH52ik2Uq1eTW3sbGC1418+712rrJvsI053YZq9XQhxDFHaoNvA6Cwa7cALqSW7WH/muaCR
9Ujk/sgNG+Y42bOhyvW7GIHQ2LB3eW0DrJ3EnCkTQeIfm7PwmPIpyy94jkeQGzpEsLgszYZX9lxL
IMWCPVsrI0QHUkFkDz8htDsExv3FbPa0/p50ioP84vYECIsDLRcAbZOHiYmaXx3fBa0w9sv3LCZo
PSGB4SnsA1c2v3QI+GegzbTJcyYU1qLzP6fXw0fZQJdANea6qDyCfY4G9c+2ndlZkEaAvdfRxboa
OFopEz3HylkXwX4i3H9uVMT1Tfqjau/UN7jU77kHt8v0Ig/cMBIr2ydmbLFWBPVXaDGtY7mkyxiM
tgWqxnoLX6ilAhH62Iu9zDVLlsHeIZJw/aqg2LSZeDVVfIzZ/v1vh2e1BcFnHwoySDpiP80Mzfey
lP6c6UpvEDcojo1Jro7fyygh/mc5Bn/SAAhs5Z2tmxZjPXL8nY0yPGD0F/gcj0OvNPVhEj1VWjv6
eXxLJWBIgoNY9o2Nz7cYMH/5ItdZWsh6xDeEUVmumgbAyYEaz5jcwt5Nl9d9COWB9CbKyeX0/IbH
ZrCQ+kuObCj8HMOnFUHJwKajayFsPtg+Zd5bCSFydupIo/YMX4/Cp/NxkMGmSdZQuY6dmnLTcvnH
1qunlveo23gGhbztvCi5exeL9YbfhFd5sCuiH0EWsppr//I0CZriXPGoPv8/m02sTPJ+ofHMzP61
FpQ+EkwL8UAuEhIxlE1p6Oyk55eWArBB67d8t0OPuZBiyiemvkLEO6mCPcNC37jFr51baKuhxAiT
rcQa2FBTBtwh82XgT8c3xAVuQkpaiV5vDoZhHIjjhOGpjtVtfmXFGY07M8CtN8vXMdE71NH31ee1
x8W6uLvfXt4wQ3UOFqzHmzuFgAuiHsP3/OBOvIcy0IBhRPbZKlY9QwFo2CZ4EAKwA2e9/IuTkdz2
WcHTaascldeaqfugaXuD1UyH3C0xVeB8pIDypSNoiGq2HSqfAX6s04yHs6h//R5slzgjkhcQdckp
tNPQkNgifJ+N1FyPm5l8PNQVynmRT/ow6yPFYCf7bRCVQrK1pZWSncHwUlJguMkCONRZQ48MI9XQ
+5z2tpfEFd4m1j/cZto7EJI2qEbYr4Z/gX07uSY6JCpSFVUahqaT+KuiIDmZO26rY0IvqL4UO3jJ
OZ8FLG3y4hMYAsBonNwBrtZwgc7TKCc839t7rZKW0Fpbe5V4nMVgPG2H2k1dV5TRAmZqTwtntRQM
xVzbjmODzJsECwCgbbUhntmN9+5qS8Q7JheiHDj815wBvnud+hV5dAeZApahpYlJOZR29mgTheFi
1doMQ0pL9wFOXFDCDgemC2wAUygl7cCSMTwJ6UNLUVfH7mqQjUrmX43Gh7OGLgfxN9yfwx9svfAX
n6WBsad9epYsQ20soKenXuBEM4fTfE7LoMvDhHyndVmCcXA0vqw4dA02SFvpJL3PMkY6TzPgleee
wRoy15b2eq92pOQChxERP3RyEzAaiTLjPO4/xovd+wb+cEWYLL26P+GVyfekI9TiidvjbWN3hUZ/
y9H2kHF5U187JE6d31OBxe5Sypf51c3GdVylakU8czMmhhapMM3GEk/hljwjlNUcOC2FUQPstxao
V/U95N5H6BH/UCSWtTtLAlDEG689yB2pSqEOYd3EwrtCUBqN+N2qrNSMl9Z9G0VPJ7BExq9obptq
ap7ymSq0UWcBVc9OPxNvq9eK72e/t+ltpi3X+dpFgrePR7NSaNXoupKslQk55n9POlHcgSmCKQVb
ydVs+X1JNk5bHlhqVtQBfc6ME/Nt7m2cPrtcMleHdMmXy1fwg47dL69Y+TQ8k70Qh0FhPATLV3yc
LlFesEE8IMSwAoy+tJuzDR2HwTZXEDWkM806/3+VoXsAbGY5RrSHF79/kU2h/PwQDAILpZCeQG1t
lkwrg3oqNq9CDF9t1DLFLvZ9LVr8UHUpODmXC+ojx86cOZGDNmANSKH5PDtPC9cZL4hykKuHIv0U
aaGvBhYtzGG9XIC0+KCOPSoGWO3/MdPnPK7tXYnrT3b1TehMyOgS4wCSjhxhdbhlNpH0cI0w5jT+
A/FF7UraKghJ69zR1RsLpkISFDfoqGMl3o8YTJfo6ntkq2JJzB3J52g2SWLB6F5NS/66fjfNWf9e
Riut5njV3wp3FM4EEYv4Q8HQmfjMcwKZcRjJ+nkTM7Os78+Xm+AW55T8rgnwyXRr929GKMr/hDjC
ODdT/epPTRG1EKaBSieoIr14pxFlcbJD0K8KTV+QRif7qDSTkSwlrdTVAfrk9hwazSGQHP6bPxtu
KoUyzPiF6lOAe09fPfgDQLX7NFcFprPATpTT8rzCpFa9SjTOaKCs3H8OuCkPUztqmHlydVm3+3lx
VoQwRSRJmKVOBC2Xq+utjHqSBIigLsktnXXhpIw0qzrzBc0U24ek4fHBPhNjqVFZuPm6xRcTMrAB
mQyHv2jIGr1u9juXE4AEgEjReR2Nsfnn2jodoje1hXeic/I3W0nxhdDG4EhmVwWNFL07gzIbqs7Z
6H3oPgpiAa+AHrjdmZ46fUKtALN/teENvNEsMCmjL/NCa4YSTpOGZb6hu7AVbnQOoe+cEjSpIQV5
qTaIKbgSjVx5/w41wgufKuBvhpuPzNNMDLzhz344BTB6npNwVQq5bbf591f9YXKCebktq22b9/U5
pymbZNCS/ZyTSnrSnucgAbvzk6hsiOX9KCH8y2qKAiHka3Y4pKgatVQ1dwtuyg3kplP8MmoRgpR6
YkKCmNNuNu1WCS9UBGJfR51YEI1rhQDckfi124u0e53xfCEog+FvN47kHRGbJRsESeP5oQU1Yltg
3YFMNQOAcmn1dw6bEEwXJ3aZUVY6Onj9ELjmj6voF1JO6bPyQD1lp20AbaXqxbskSmjyMi8zDhOm
h+76KFdJEzympFb0ZYv4G1RqwXNr9Tm1B4M5rH3hnXOZHzOdFRyCcOxxxSUZHFFSQ1ShhnWbQibj
IUEibQL8Bduwap0WOpG1N+sIndDK6b7XYKgfeLiTZgt5AzygkwahJlRNnDAKfK26FYHWe8whhAPc
YiZwdFC9q2NJCWtKevpsnxs6WOJnCJG/ttC9Ig5UJxrYaL4U5nGl90UJ0fGXWrpajtfR9vLO/tWV
BsWw1lv/nanqLjnMyn+jWPQCzlxmmDI77YtQdVejx9qteBL5jGcjj5VcY/BDjVBV+xDze0wfqE4v
sXxjBAWCpWcZrS7LdDXvIHvjSskCmfEM5WPdOta8DgbdVpwONSaSq9vIzAZN3iUBZ+5JLWVXpUb9
S0Y+ahhVvRnjW1yDdqhEHSG1y9YBrDDZ6skwK0QcVjDDD7G7tdRTeGiukOypk0+dGN9QBPIWn5AH
lBWevxHGEn2V7UeGVlFWguSOqOkPouVUStWHq9DTRSuETPRIgHtDkRfmyC84xiX1VOA/IB1iXBol
7N/QQJDDvUep3NzsfSOkEjISFPj33AYxSApC16IoulS1U0HprYZAFf9q5D/VKAzUM35mGEesdU4C
JEFN6sbr3ZI+isp1hiKPpQIBGTKzkJFgluvBPoYxwSRI8DHYYh56tLfRxmlPVEiUeATLn1WhvOZh
wrOahf5eybsLBDYqOXfmWTP570TlyKA9TbmEgaaD6SF0xx/5h6ihxOZtb7t8xeazBv+dH1hI1vEc
mn8w3770PmHmt9VH//voc7jZj0mg5Wepfr6CQcfikdC7YxsrvNHLTHEXElCit1ADLWk9CUTxnipr
tI9cX73JiTja8jLBvmDtudQ/3H0fSQMVL6BOLJktAnf2dIdf0ovlcbq0NhtK+3t3rxCEagWUiz+A
u9ImROUVvWtME4fq0F60EHtXhV7bPOVvlHzcVkZ2O1SWKPKkMhX48arPE7u3Oka/1cudBy/JG5UI
T2qSqpcoARFcPM6xeA+bVQ493+R1H7Z3RpYIms4cMs+37+vW5Z5qwfqv8OxFwWrkN49y3dgX9UzG
I43pVC1r2iDhXNMpiTJGcdzijjgv2Lh4Y/O9flNQlKPLTsGq6QWU/lHNYWQkJ2WgTmR9xuL250pS
eHwiEyGcTM5mxW8YS1VSbsof2g/QfsRepYAJmrbfAGfB2QExfrf/LLu4X/TQMnsadVIYqQ5de4k9
vdBYBsxPsZTyfQ7+tzez56yA6MXuuyltO91oS8VQNQzDRWiH8NK2+2Fg0uyDunYnmv+Xuf6KAtML
Rg9OWtCkEKAvNVJ0DGswtsoax7D6Chv4fRZMtkA2tPGruDh9/aGuMGeGXVFWQV3DUP21tGEKrhQt
r2Gv6ump9avSG8+C3Hh64AZnqsSy6BEu16C4n4x6AmuzL78tsz3/I9KIAYe/DsF1T3EIR5SOGVxm
R+lg4Pshz2G2aFhXmpZKAxGeK+w3pTVcDW7lGCZNH0IKTT3fGbpE1JfJ+njYs5/V3d2js/G+LCLI
YlGtovSzFwWOmaxrQEF7Zt8ru5CyOhzoVoFE16CQFTMW6+3OJdtoAcy2GVi7epsY2gm4Rc0RZysa
9IukV8W/L/kqlCZtHvlS3rtzc7AoqSkNEgLs9zZcNI+1VR/2X8+9EXILGUdMmN3+0aVHK/TtqjdV
1aDsy+NDvuiUVG33eCi5/RippICYMSzGAIU+i20+/olsEuIh5lfGv5mnLF7UY12NP9aATag9N2V5
c4u2HyQXT+SHTpLXb0BIlwPMMYpOh+Dt+iwU3b9/7pqHzn746WSV6Hb/aX4SYaXMoK6NJ3TmJXJ6
Fi/u6316ZO3e/juVLuiPSW71ar7aY25h9DI/j67l75yqMz5jjHCpKc+S/9H6wNOGMRNfl81Y3Bor
RfI85DgveGbD6C0/C9TXXiTSXNykGjthGyxJ25gSgHPd6xO3Sg6YD0LOdVaUAPc+/Jng6pkGieFo
MQC/CAotbltMGvMVlI7oSGJLXbC60AoNlRgYQM452OxP6qcxeMAdYuvOGEJdC0TT7VITKE/LNFM5
Pm9YWKIl0gR1Tu+1zBlclvFKSArwXWtkugjtWb66gaAh1O6AAn0jPiA+OgceWjwHJcLJT+fyWc6Q
lnQl55vZkGUmlsp3zu/ICXL3oV6/1fonemAgcJcqZub5LDn3guT+b8IBE1mmXIhBQkTqc5kXjAMH
Dspau+g9TjQW0oGJLD0vGq5O6BPVnVUaPxPh2uLkD8sSBOTUEco6koZVxsFbyrRUIl/nZvtIdv1x
1L8y/AM6Cr0r0Y3MYGwdNDi6MPAxXWXSmzrKSVjHrNiqXPjCryV6UWpqLN5M/9HaF/Jyatn48Qg8
e3nPrxbMVSKZh2G9y8k0dVRqVmP1Uy2U35jH1aQOr5zR5zN1tcf5X5wj4hoJvhh6AWOnIavCJBS/
X/ZNK0lnupfKyyS+jNxOkvzD0oVqvcfR1fE2x2vm49smeBzjIseXj33g8mrMjgpOr2HIJ99rqgOe
CxJo1iqB7a9z5wFnMzHST8vuYtzQ2yWvfP7rKnVIJ+FY+L+4Fz88MTBb52sLa3HJDB3LvAc6SUWw
pKJJb3du4n/ejAA3DuHeg0vZh40bd/PkVm1+AkpjCd0yGQNZS2ZRKb1Kuck1qkGkAzlebMlOREsd
JpmZl+lkOZOUGjKnawkB4H73meIxIS/b6WmGrmdXcDp+SNOuPbdklHz2NMj6yTKUfCcJOYLM1h9o
w8vBOqBwzU/WvTrmXvBbZxbjYdZ6YHysXgeyPHhvhvTLbJuhT8zKNnQnp/ugo8QD6nZXGreSr2rR
ioAbGpbO8eO4/KOdK6Q3WRDj2fiuH0e9IJW8U87Cd0fqCBf/V+b5IsN6VzE5Q/JnWKNsLNqxKcvj
i1vW6vfYku4nO0Spazv7OwIqvd4nClAJI0FGOnIfTgsMprkEfj/4KkiZ4/THFMHGEvNFcpixNHkv
D1ZHB8ozzXnPgb0E+RGqr6OY2o+NW66CQHOq3nFEuvYUXRmH7avFQpbwGjRLKkDnV8ni5t2cDn5a
ThQ2y9g3WdpqsXLoaPIIFNBxRPfQPtmv2lWUyrYzceubb3mpqPBVAc+YZphbLtIqmnpeLNKO0QdH
gZ/TTbI8axgmhKxl3PH+lQ7lz5kX3hSTORxYfKbnL+w0eYYaU+axnnkzZqSynvHvGRwKkrF5i9gK
NK4Rx1x1Eoe3DoKjWpkYWSEU7zBSfECFV8wa0tYYNsnxVnCrVMLBgoJMdTEOjgjnYcbUR6hNvJXn
E5lHSNy2qvvd59mHSr193PJ/0l8+xHpX8nHaX1zGaH23OOUTlSZ0CoweAL4ckcXFnM7AvQ/55cjW
cjTCjhnX6X3NDfHoGcfdR2Ci1+qYjsXjER6zCi4ywafSs+xIje2xFjuQYcUQREOz73vPKvJKN3Hy
lTT8tMW5c8k2MqzL8pG3+Cm+YpU8XyIQpC3BgE8WtrLnzsWI3SiJWvebJ/K2pGbSXeN+h39dDHpf
IztHqLif9jQCEuIlZLzw8+jlcB7VbtVwHYtsRwbJ+WWZkQu5IfBhGIt70Y7wtT4ZZEqlQzM5wZgG
56odaP3FAE3Eh49yRgWuwo15xpVsGWKckPJqG1VeYDMD8lKDXOtN4jOuVs6cbvuyg8rg5TpqqdiK
0hY8zmEfs1nW4vpshmQDfiF95qOwTyPCisdgM9XIVQM2gK5XwZWTxJnVMViRtpAF1bjpUwB4oFqY
ilZ1AsV2aDbMDBaJRXdYX2eMzDu3Zd4w1IqgdBj+KzYbja6/T1JthJaqLy8nIyn9W5v/XaaPVQ94
TJT6RSN0T2i+Z0xXuiGPmtBCxOIOfFz7afZAirIFRGk0COcXSoS0W71rqJoUEIyjpxT3RcIsSczO
D+fhjbET/r2aFg+3rVq26A/GUAMD8N9G1bTRMfjITcmr5ZrNU0FS6D0LzlBRVeqRNl0cTCwgt1Hb
PDVYslCHztW4SMMSyRlCRWLliEsf0RrtwIYVHHPSEhkP2ZcMgfwIlRS1M8/H4TxSvlzWwqO1rGYJ
iqTwiRrEmQQ2llgPBLE0yiRvns9n9bsKb5mX+BRVJSEREMxIGxYLsX227Vkt8sUafIudwFp2iBWr
Dp4lJKck4pk1OZgJUA9oMSq7ct2VuJmy+qinJONS/W9uD/4CiLEk8QHizfBASZ6RRDXAwfN5u7L1
HJtFieyDFTaHvJcgmRQJ3JaIqp3tiyfODfMarCv2rEq8Modwo3vs8ckFunNK02UlcBH11qprp5wP
4U4hza5xoV3k094HsNV6MP3d2b0d1z33n5QyzU1iQ1LtY0vnkB+B7sEXmFJWH6BUdAKerP0fZEpL
g1zRHsUNrq31s6RBJWLS1W4Y1v9o0Uz/KiZTzsNey8oxRixbuDgFTdgPjlNf4MIVdghd0jXkq/4R
2sNinE4kIvsJKV7GD0UkHgghs9wnd1fQol3S3ev0dD113dSD0U3a2hj0r+T3PYo1qszJM62K1IaQ
nWSwtiy240vwBZXdd56qLKvwXdUW+9r1l/7xVNqf4nYX9S1ZOVc0AkZfQ61cjcfCp0Ou54gnf0mh
QV/MUBdGnUHOKYqgdQXg1m5SxbcMA/aCcZ1TdzrGxrMdy6ApANhQolpYpl5TQozrskxJbin9rDwZ
vJzKRnbtMJuYTuSXSgaB4WOolHJh4b9BiRxo6YIdpk3UXM9pT6pESgeKJg0rmoHr36s3ogG0zwFt
wDuIJiBmPq4bB2cKwvtZEGiNPcyrmC7+3d2SRLIOaqMMYdeNireSdZOfZf5MIF0lcFZQqFRJPzLe
1iGbPDOTxp5wRSp6b3f0POwYCiyNPdCrjPl1WiU6kJ5I9ufnhMac32IKeuHU8WhK+SjFjP8lcAqi
F77u9gZX1oYbKtVF6nogcp7XTJVNgOAFdLkLXJN2HUYE6Izes43huUvoBVWLxnpvxdTDrbtIi/9H
TPzL8cw0E1CbHQQTnhdxI0U18otngcffLx5Kbw4bZsDP0FWlbON/fVyR3HmQcWcGGXSFWZ1715an
7Ttg+BVkT/exH5Xin7btNKouEfuwK7sF4Bh6kTPXFsm/rAVpFKf+qzucTjVWLYPlm1+K0h5Fe2EE
3t+fvlUTtF7D1nJl9oBEJjyP/S7I548bnZnsOpFj8zMH9/mvxkJkAt91aB2QzTJGzVGcR0zR2x65
xAFy4wo9H+a1cekhEci60+Av3b8zUXdL+O1i8rgFElz6J5K/h4DO4Y3Fo3qGu4rFqr4bG60yDKc0
sQVLDh8+pXroRUJI6D/MUOR+8cD/Zvslm43nbg852wm7aZJivSNiIuAM1dxubZDqDhn19pETe4vs
VqAWXak+HcGai3gzEbFNv2mzi79qp8AqlHsj33LhTFiHaVaNtDZdwNF57AqYgU6LdQzg/1YAxwHB
MhMoTtIvrtT5f0tu/ur69Ku+B04OFV5Fz5sP+IKA/AsERGzT30ho3RpVZzQAenTyLuRHHHG2CSgL
jD498NZMpmwpDvKTqGDbmdULsLxNFbmD2eXYTGXVLlnAzdoHwx2pIM0C4crSM+EUWRe8SnGiFpbm
sdfhdlSPxpzdi7CPpV9gcPeUsIBYIRucEARWKARNbY1A/imIpZVryG8TjKCY0UHK1ydvkh72Q4Fs
fW2AGHVlG1ewxCr4VChNLcIx9fBw1Xe8ADhBZH6KyMXisyLD+Q1orLCEviRybZvmK8xSkUqLr2jc
gILiagyqEm4pH8lqizu0DGXH9dDjOlliuMS0O4KSIB53mwqRvDlNoVmdzqgqp41CmQA2zhyRu49P
Kot4o0x8V89VxrEzNLok48fwB1IiL2cL8RJ04iLuQ/97q53YVwgsQ8SVlHDCHTMo8rQX3LG5TI57
LI0IW4fGYcbiH6nxoqp54+OkCTMyCvjt7PgTwfV75G2877SJv1rFSdIluV4lp2dBB8abgafZViI1
6nld/R17UWbf/9sD988gBuxrBzKxvegEECJP2y469kWCvcHQDfu7N5nItsZx5VMycisUPfDck23g
ZzsYl6HBDMOWPYOgVJa/0bdIHH5PN4OVHAAvhX4elSFpcQIioQ3eKq/Gv7ZIB+0v41hrpuESqMw/
oL8fuOgJQ4wj4rN5hmxZ1H98hGx7zwVjtxadpNxK3u6cvNrquG7/04Vm00rx9nhTy3IiLaS12fWU
WPLpE7qaYGROyVH5wxk7jp1/83VV7JAnJBIqRg7HLtgfPhc4s3s4wFDFqcSSJRyBAE4SWK7T5edW
EH4PxxbPNgBmLRrd5l6S7ng+I3BEWLaoCKHEBSe7LfS4TBhPp8A/HTmVYB4Coe0BIRfk7NIG4UU+
DIbm/sQvyIhxDi47lwySP3b31hQgjmFAwGiNkPgmo6noRASNuCQavLlwerbRCa5DTA5ZJi+4GZRG
iUaBYCr31nnF5m4br2r5CrNNCGjezelBjGv314FiBcKad2FBtwFAf6crYRztJa0rfJ0dwF6n8agN
ZRsMsznkSH81Q0da/0GMIW/NNbxahNnaFKVzGXRFy3KS04TTdrSRXq7lJv7q+bSCTY11EABWCkPD
nO6Y7Rzrb2Y1Z9/MJ7QUauQ9SkdNRSXIF31J6LOFQV3xCtAHrI979ZlTbJISEEuAROYx8paPw3FC
y0U0TsgetqgJ8Dgm+jd49jtynz2XMuijtegoGaet4jeCTkJSOUS0NKxGtozUF5j8pkwEI8OZQdb0
nvO8VmSs+a4FF/8jE2yZV5ZR5S3UGQtVOIz2t2TWeQPtIASNOa0c7eQs87BFja9R8nwz4g1D436+
8cdud8FIfHjebo9sUx18g9vQZBxoTtJQkxOd/AKszhB9P+sLbanxHEnUjcTzRa45L2JDPQXOnjB3
ai7MHJAceakgdBhKIGeo/Iw9sm4eeiLSgjlzBLyHk9wbePU5a0xrTPzFJhbzPDGhMjg+Q4El8UNS
aDhGvVknM1DQrYqD+eqfKcgA8KQOZNZUdKxcMbr9TTnP7ZrNo89MTDsx/Hhs40lKzDzlGKTf89gM
Rd9hsRK4Z439MX9XYdHzJstJmnswEESBFfuB0H/dmY3RTx4q4muCd9KZWXP0RMAt317bpgnYa+y4
0TJFsVw1TGGwOlQdlPc21J70cF2Toz4f8oXLv6qAV28Da/z9SUwf+grFvV0fSRgt/GfiwXmWpsR4
r5CaSwpHJlxAOiHT5FvjkjYl6crCGLbHh4zq5s+QBpwzEZ34oJAy0WJ6fPxdqZ/laMRkxMHX6Wxr
UxfBXwtdZQqWxfoAIZ5gN68ii9k/zWK1HZvPSz/Kg+BG6zhFITMIV0dyrt2LneFS4reBq7XwVvmV
jU6fIcQFlCBRbjVqmxkGTRvk6IaMwpBBEbkPkM8qUA6Sm4nF6272QZzbTgCqoEyBDpyrd+jbpAmy
zwcNXGs+P5VviVXK0M+pFcecpLZrb9y9ERLoqPfoe2x6VMajzyiORXk4lNzDRLer4PVFiI64WIak
8G/b/BOWkSemGi/augDCXf3yA3B8WXgNzaJ22ST7Z8OAErO0ajuNXFbeC+0iwsB49HEFIEsID0Rx
QbkLG5OS8gWr86sboZq+a2RH6IV8zzaNd0s8pktzQWsUECInXmTfcq9hGP9oEzV379he2me4MozP
/fuHVq5o0zUL6e3nbCJK2V0YBKev2pepjq49gX8bA8nKxw7RggO2974Hz7Vr1P2HPLWpYqVhCd98
f3Atc5sSIxhgUICobomjobTUYIFYecCfCkbJix5zYKY8XV7BwjvVhHeySGsaObwQobFEtthuHLhL
WixqfmWJ/K1A2JH1CDOgg9RjvDjvRo1SkjHtY1h6NnI1kWJacOFZtZ+4cPeRxCMb8BEkV3J4xY0T
ICKhn+uXKpcF/vJOmx6HKrnWIVykC04NhD7JRxlS0MyDr+dMFItzuXbyznnEc3rzT1LnL8RY8ezx
2jTfzoWFn84MxrC4QYIoKnqF72UrLLAiImhP5CutJO4poThXGewYJoTZJAHQOLK60L5iNh3/0Lmz
U9/GrG0SL13MypNW/oZY8dTvh0I4XrbW5c3tAhQd0tyVohhH2q9CshHbxDSe4+ku7nRV9XnfGGZx
aZHTTWpm3fNZfHA/kEW5V1TIy1/EM+BW28NLJbb452K0X4VfCrXi18Sif1yUYvVPeQIcw4FiA7qG
fACTfBdjB1+2Bi+ZX3EhIq+rgoaEBsc1aEqy5r7z8JTUVAlPBfST4ko+NGYj6A6VrpzmtGXSIhd3
mdP2FEJalLSkDGWEsWFa+hmzh9I7YWNL1v0vlo5/Q9ZO4APXbF9jU5L0xbkqWm/M8KhSC6yLSGiE
N2/bbKukpsMrQFJaX0FR4v6L2mNeyWVUa5HzU/1FGalPMLyQVzn33Uv26HMhFydQb9CfH8eTXUdt
BaBEcamLB+t/50eHqaG41QQHyucnQ/PeuqbJ+Qs6GDc19N2gEVsWdeUEi8xfi/sdfGEkrxtfZD+I
+yB60CeRnot8VDWxGweUjYAYg6wj+17DdrnSa1cb7FP+LhaxkDhD5SLJQsr9I1WTW+qoiRq1UqHQ
DACDd56Q0ZK5AcUQb81bell4pe508DgEVocqwrhu4aUKgsN42J7KactVX8WYUIVSyFJR5sJdn3ga
O3k7K67ntizkg6XThlX6BYNdS3OhCq9PRkohhjpDrKzVCIEJGnWSQXKKQH0a3wegMiKVgEGVygqH
X/emwV/SEblRhry/lSpHS1TAY6PbgWIGqd+I0/Oi4kzNAsTqme8YRUi1ur+FLBKspgn96hX2jsxZ
pCo8Ccd/3mro2eI4kZETKOtcGS5pTw4hfatTIzmiXHN4t7SxGlw/J2mEC8eUH3pm6i0fFFgGBJ7N
PaJ1myq/t2fRzufr6qPvjyzZL6Nq35vEFAiNknkdXqZU3TnBPCd/O9Ok0gUA60Kqls1Dm2Sj0EHr
MIdWrFgb3T4pRyhRwqO5ENvFNOazkANaraRw9bQmMTIDkWOA4GSfFw4jwHyYkSj36ZJM39q0ttxd
YI/IPZbyn8S0OUPOUNiqjuwNRsRKY3vQhQTqID3pp3CGzsJn4cVKd7XMUTL2srrDUvemy8RRsrfd
cTsxft+goWU/0ActR2/Bye+LU7hIY5ss+Pf2NHS/Y7hZoOY5XCzxKfmk3Vb+PbsjK4Y9ovv/zOaj
smHwzzVF2t0apCdZAZW9L2Ut6hp+t2axC5aKXfSLCEzMb3vMqyDlp4xcm7+/epKnns6OYxSVut8m
f554ob1CTbLs0D/qxmn6xzEEaXHf+xEIoso0OnPk60fCDgKudMz6nJQdCOLmUMvUXEgV7LaHra6v
eOpSu8A3gV/S/d/05ubiRwZwF7QS7lHvty4Mw7mz5szlLbXhMaHub+WFZPq25h6CWG5ZdL7wSThD
RyG013FtJbGsZ1QTUbjamqyuysWvKem8N5X/nEXeBXcUMebXwv7KGAHXr+PAEGMBk6G0uDpd9jeV
h35V5KpRo2VQA3SQO6G/Yp5gCKCsC3AF7iXxLNpd1L5omI3m/TfBdvlFQTZ2N2dgc3M7yOH141qI
268p2jn5erOmmeiuf8J83Yygl7Ivh6g1oD+Nfj9/b4V9tUa1UNqdyVwmeHN6Cf0u/4weuNGfVoMb
t/q4D08SlS4OWLBWWDl/HpNj1WmVSORscaMBlXu4QfSUeOQpUCEiDd8H4IhW219AWGtxpUgioAn4
bmsqcEY6CBkGwxVBRxwV1u2kut/t/TAgaAobg1MgUd+5LXJfDwDTIqWd+G8js3ZaVriLqJZ/e0jT
qPp3cUkXKqUCteua/gLCXaKectWHuhfuONU3b2iY9rptG1vPTVxes2txpE2Q3ibXnLlAY0mGG9k0
5Pw09FzVnqLnOFO6uHrh4plkfcBk7GBsjsdFaqiytXYUAAo8XxydyUKT0YlIeK+F4YwrFuUFvNcl
Bg5Y5O62CXRf9Nku3Tv0YRWSxya6JtnRLbyPd6spZhQQ4IGWIcDnNxhr+sXlBTIcUBZxTO8fGkSz
VswxXmEbzL9AQlDTCh2yc/McoLjuhtfaKm/ZTu9XMx6xFRYay0CFJ9ZFHLf4KsHwumbXl0zbgOr6
DKQcEXPOIzTUYeXKQDt+PTICqaV04JNZeBUY9euZmYkqSlMBtC7KNdt0ML1cNYoPMo1KuRv9beY/
A0zDRA4V0NE3Gg+V/R2pgxbMURi0ZyVuU3tQBH7yV5LSo628qMDbHPnZcsHK6Xe+Q+qeoA1Z6GHn
esVxsYwg6OCX4wX5zRVKlG4a2ZWeBQVAhpoqn5NLY5MXgyqRW4fyNLv5hHC7pjt2ZPyJfUbUHQ+o
FJ/VYRy3UPvJLF4MbawDvuE20OxFO7u9ZiEE64Rx7K3ZWtxW6aPtGx8K4PZiTlor5uHafLfGHI0u
9w0d3fwenmMdtn5tlZOGaOGD8DaHw7fEFt3ZpZg/TWF2KOoyHwwCGt/0cyx2i/7gqqq5DQex57WP
4IklMKxLjpNDntLePXTYgM8Isp7bJzYcmNOul0hjVLspbt3GASCtzvTtgWBk1nZMlvsNAbzcoVjc
OHovH4YAKDrtGJqktUavcKBlSodMQvmz7eBWm22YNTHJRjOsJmx4WjC+F4kNdrWaf6d1VUbpYUDW
FLeomf3QS4Pfw6JEay48X85zGeqVUaRdhOy7tDSmwmOf6v18CSQk+maw2kYFrDEYvZn2YuT1hMmq
s3yrPz6ntXmjF/GpipmOAM2HV5KvkvlSHnSDA0+sejP4M+7IcBmWtFjXM0qi4bR68M0GFpbFQh19
DkYC4KiQ+iKNje3Z2JQ3BhGKxv9usKSdlvlUW+5SMo05qlAAj1lFtYi8RqiMeSG9CWn6hey/UwWR
sRdAUkp8GgJS76hcvnzLT/RqyGaI9J8IhwRWdqCNH8SgNkhty/Y6rUPi+icK6QnhEYTAxcPPyyXl
QO7K5I6CMiWDesdQCo4nBnHx8el5jKvSXKJgksxRcn0alaGN7tvqzjFAkdSSFjQeczQa5uCe4XF+
I/tBz4tO9yerr9BnpziddYkmbx0i8avCf3qt3ZCWVtaHfAzYsON1m/Z6LFiQ507OudDgd2XMp8pf
uxmyBM0DZnjBJBWycP6+Y5bMcFKoqkyRiv0HVl4gNwgoW1yVqmC/LcdROsMqJ8kZIMBErqu+5J5N
vmuRM7diPKkQcNw1n/sXQ9zVB+TLpDJcP5pzwNG4bgp47wgtv/3rSlRs6aHI8hNzIIU/IMCNhwB1
hPi8zTID9jnuATv5arqO9pBTLQoskYocpWWx6lUCY2IxK4CmUQaOMnhO/7onnv5IkH/xloiDN6xL
9cxiZVVMxydV2qBPy77tLNbJzgPF+FDvD2Pf+pED/1KPVdhgOHmuOdUMqS8vkKljNSxvowQ8joyv
TnzZhd9l4UtKOB1cdZgoe93NXHZG9FIpu+XtSQ2oeCh7iBbD3hHkRlBf2x1thsUXUjLLaN6u2br8
RglzA8jJTJr21479IG7bYWTfN0rvmFnnPMzYbSTO44mUsSSdcplp7E4TpzD1OaZKnC77suMr9tYe
n4OUSXZV5saIAlkiyGIAkNFG6lxmaeI8XgArWJwpyICM3XJs6WdvrgXz+0FsKzoBt+4kJ9JnOQjD
MINPNEtV1G1QTtYzNC4Og/cXFdlspCQd1YxX70nSOwHx95YF5WjYNohvE9pvJlGFFh1bFOEuErY/
K4sooF1D4i+iGWppA0RrYyOlgUT4nmTZns6vv8mpIvgcoCG8CZ90KNf45Wgk3fQkvo3TXJwa2lw0
IAy0DX+/TsqPN6ky3ygVib7QYNFioQSp5cMqlCUS+LWyWsPi4RvR75Y3cRerii72477Px6P+uXtl
PasLnb4YovNcS/EPF+O5O3LoAA/Ss3ECveXiqy1vnu8CbuRlJOwjI6QvgwTmNIxc3e+53by8N/eX
8hf3huN6exIGm5VTXuNrQCG7nVsIK3tMgnKw2HEs/YOL2H+Sll3aIDmLTG9HKaBLHCNUISBey9SG
UVz3GJU9rE+eDY+evS2LVTKh7RruIVi2vFVk+KREzUeD8K/L4qdgxQ7c4FyMDRTxA66TI7wyr/k0
auMXATKjagVZ5wf/vycQ7mn+t1ctAjwIWDOo3ZSYWF/Sir7IQVzCclsDkCjluWdpjrh21tDl8LvA
jAybyHoU5Uf3NK2VUB26Dga1JGQ1iC6Woi76fc2Y0UjwzucMVNl+idSc6dH48NOf2iGRZfSbZbUp
F+9C6F9KEcsUwAE+rkr6spydiGqDmT/HHaZzmIyJmD/t8++23h7ZFkmHsbz5fvSknhHmDgzVmpRn
qftfUsgDMGrfzn5hQtkvTsCQYyjt3dX7/7WgGffSsalwWWdms+Z6KVI0CJ8IL8VMKJ+TTh8Z/RqO
RYqX6sihlzgUBqKDO+dCoeLrUEr4+CrkVVW7CX8PbtycwBjmlC8i+r08Ty88DQeoq9aNgeoKrCm5
MIBfKmVQ+oGb7qYpE3QFBrfSeDGflgHgoCUtFNLrAF7YvSwHtGJypp4pXiv/MbYxTGNp6PS1q265
c41aeYjMCsSMzS8YBO8zKNkW/6QuG9TsCFFW9i/Zj0MaBE0VXfPaG1faqVpe4qh7Ol67ueC6PgDL
adP/t8IKUqWyJ9TB4DOk5MVSZfmrrRP0LqJAMgdMQ1mxLxB3jxdtjBxNAgwlf2sBTRS09jnsapyL
G/8DL809AoD0pPGmJlk4Rh+sLST6SK4k/321yQnv6ucNyI85zZmbj6ztlSU40wj8DJ3LkFn6JApp
eWZ7Qid9BOHgfnn/aNGhzc8Oh+T7UfU9v7oSM1zoNMSI+Uy/RTiaUjbhPtarDbYDkGibAgurT+lO
gj6FHsno+jF5iAYAiXvWKXd5364K9md5K+F7dQfgMRhxr0UpjtJ14VjPJONF4JBNJNdlQU2Vzoea
e4aZ+Et8p8BIFTEeJvz+VGUvZIx3WDSxPM2vfL2aS/iJk+IuqqVJ5WjltzQ8njFo4QnmO346nOvR
6NTXKaRu8hZV3cgH7RuV/RXbrlfnUZdM0hjRAS3vI5Ya2bYNge15gL3KU1EZygmZynqSWtKVwC97
M9lGJijT6KBY+b93WdENVKNFqytIVx4BN2V9k2tpG1kRsLZwAEY9Qo5DSuJzr59h5XN9ThPPOxgU
kIuxwuG+MbUJno1O7agqCFV/Td6xGnfibRICy4SBUWR4ARrlPHrzhXsZ21iNyaResRiHXKW4xfWv
44BgdD/SKkSYsTWexGacbgGKLRkaJaFRGwCOsh2tUrS31llJEXiyweP6ecLTAnVxjWb3cx5dGGzg
EKS4pwHFmn3+DINywnhXuvJ1i3azS3mxro9D8kVSBCor9Gp1P7pNHw8PPMsjZ1wgp9+Vvs64a/r0
ZXS/TohUU0NN7ehv94nn2i396iWqU/vr0c9zgbMyCQOVuxwnOKDHzFbFMDp2s1bXUPAa9GfzHstz
6u1P+BIWyPlmZ8/6RJt5GFkc4nDZv1IyjuJZJGx5s5zgHFTZzgo96RZ6wAVp29b9roDrEQ4Dqn1z
quD8YR3vG0tAfjTrjMHD6isSP3wmXbF8F0YK/q6uMG0h3cmSirrhR2RoUK3/ny6GsicyjGjpP9lD
uzxdVU6mChnHop67EvJJuv/OR2SKMKyh2V6sOr+OxE8970Rq4D91Tq7jrhOJ6zhcLLdBD6PXW3jz
Zxt5TGalnxmAG3gJzzq/3TV9XUxgOXiQkg2kNkxplC3eWE3P8fOug3d9UYnzOKtZR3DsH7hB8HWV
1WRYTff5Uym8D0qmoISX577wf8gP2W8Eys1AaWNbCQeXFvDPcBHlcms4ckhRVH7984aZuUHucp2F
1U4sCgRk6iKPxYcS7jprvJkaTgT7szetEWEGcz/XOh7hK/4Nz7wpcOnQs2srxWoZmSoW0mzODZRX
G2Q2/D0iUNYb3kzcWJL0xuoMhAsfSYtpDCNFM3TAFLADQ7ymlCIDIzIp4EwLpouwIlmuJs4w8jCo
Jlgn7NGMqu/xYyfbXwtH4p11h9ni7IJaS/cuuYM+C/Aj11gWASfvaExyyv0vnPXanxMmPJQX+MGS
znvtTsZs0siVnSc0CS4VpZHAD02jRtuYOYacZwMjzGC+UNpGnjgjmpTfSOqLOmSnHb9A1qNKeS4d
Ih0WMF+6VcakVmR/zXXL61VZW0UzcotzuiJRO/tjynQjTmcGHjQP4aG4Do2D7PwvSeksVvYd1asN
OuFn0FDImc9G9OiuOkBBFyalLqiggROTjRRUYdfcHwkQN+iyR7pYGsvsqrUTnxQjVISGJUlaR/KA
pi8LUla/VACtzwQNTlty87jNlLv0UUx2pwPDYXcDY1BaJDSl9DRqYsTn6ZUCVSdCl1E/3Zx4rqB8
xQpT7HRN3Kq01aM/cMkuKyVQ5GJl8v93MExm5dcZUNSL2DN4ReoaztzGemuGCvpbNvacz3IIoOzc
tSuGYcm6buqQ28snG+8OeVnJND8WzSwZIHovzbRlgZJb2fUcOst1zGP6I2BwSuhKIQMxk6tdV0fi
EsHcJTbu6Ij9vsBgGv3jQez8WTEdbkNzuZWvttE3Yf47V3mu21mkrfbvF4yExA1zdTonK7pBzun7
0L3yilciAf1Pcfhh5yc+5727KwKWpjdk3Ey9eD1Dj4i0Od8ks2+Qckdf5pdeKM6zloFQ9L3Os5ln
ACHuGxLmbkzDQ2+iaO3N0DV8LFda/1GUJkrEOyRPjr0rAfP/KBI7vND6OsDCVkt8U+iDnqNAol0Z
xrh6NeZOIKj2Jc3UIKiNolU5RSUbnZV+2dtzCeFUqYHP+DVmuLqbh3w1szVXZDJnnMaIdupb0K7S
DmOV0pBnofNKmiI/nMc/XFKKiEYdK4IBMe5QyQM2dQuwVqhzT0e1R00gigEchKsLXFrr402IyWqH
ueg+Rvc6mqgN864wAPxfyddbkuWWhJBQHonY9upSVtDe2SkJwF0UohOlgAVxOBqpdkQcNe42mYQD
D6j/ZKJqcKauzXUlAaz3vRLUs/CM0QY/WjPRyVyZWHVbIWeE4sBAuTvi5OO2V3Alq+0BqbHFt4Mb
uSyvRwFxJSyabCxygeE/NY9/aKiQnxXsvJ6EceNXV2VsazwIIHmRuPZaZJ8gbTFykgGn5W8tsRF8
tVUL6oHF7ZU7soWBh7ZCrbBg1e2ym7ulnDJPW3eYohxxTWrdO5mh/Q8sP/9nKrf2QdhF63W9nRQr
HSTbpQo+9jDvO1TuOqzu28e9IKurhTmSEiXH2WfF1Q2T0B7G+aq8MkqDdNqPmrBaN+h0sxOmjjzB
sQZAFUE/MlxL6VL6nXBk2XVO4PBZOmyRu9bv77uWiPoRcCuAIDCLG1CCpC3uF7tdxK+iiyMn2YZJ
MgUBphuloJMDGlHC5sPjRBNrEShwYdW5ptwkUIVmrbgoN2HMbSxIU8EV+DDWLPjLFhFil1BCT1Bu
n9oQUusgLRVDu7TSuCP0M5/WwDKdFvaP9zC7271ktJEst0fDD2JKbBXmYJb+tjZQx2peDra9D/5S
2czmNVx1OzpA744vy7qpDEXhrKTn3RXyWVXZKhEOnl5/yxz9KffbmbN0NiNN1Xb59mCbhtZ1fiZQ
WBraXEyO6106cpHnEyH+nk2znnWOTJhUZV0dTW7HwDnOoo0bBOTD85M6EzePQxE0u9t/xdqTTuTW
bOUMDDcIjK3Y98ywa8kHvBEQxwjWbvZC3W5Mg6et2Bs/ItQBU8qf+MB1x4xjXKAroCKPQb0JlL19
7IoWLrKr/rBca/KIlL7ScD44mi9Y3IbOzAcNYcDhQTPlLNCRQgkrS37JlE+e2c3QJwPDVY/S18jJ
e+TwX9RPR9ahuG4zr83S1F/YoN6vM0mSQ/yhNlmiZFH2z9HpBEcN+kqPeD+a63LfFnkwGv3jgbr3
tTppRghAOJo45/ww4W5ayWL139IPTlSi3STWidWbHHFxm3tBZIU4/9xD+rJzxdZLUyRh55P6GNCt
1joBfEj+fYUKDh2Mdbo1wQHYcgxZe4hJtrwzPIX2zIh8lSBDrtq3t2mw+vCerkEWvE2Hxr87lxTN
Vc03Unf7EAYq8wgkfnpHQ6+sgL9o76UBYGhptIRUtPk0vCLky2S/U0M1MQWdAQu68P5idRPCVihL
o4O6ratCFPZkWT/SPcHttmQ0OGbnG3imR+O+/BNNOlfYamWXZQOdERKZEnUwoDHuSrBzY6xZVJRT
9seNFTFqg2Nfn/M9a4+nT7Amc8OJs7HCFfTOshrwwznjwwgpLyhC707HlxluWvHsT2C8m+d68TAX
YdtfOnaRegG4LK+0CR+yo+oddMaFdf1Oqa3HTiB8USR/lTLzaZunZmH2sQpaw+oFsE3/SrjXYL+E
ruZG/miGnbDshDiOh7dt9nFHRWrG6pjbX1uhNXLNPh/CEhMnF0aOC2pyVty0ngJ8hnrgltxbIvi3
1HdwtfnmLPNlfjLdwtwNczOmAUyNOyXH48k5HOKrp5txXxibZfKdxWuwsNcUJBOovDDHQAXa0IwE
GHfyCVeBLDRLxbjZ9uhjQYqHuXQlC+44bFONaBRWOgWmbl8VC8FjIQJdEkoo1H+5IMDTWxbBf1Ll
P1cK7V0j1tbU9gw9Kav5z3UuAK+JMb8YUdqyw2oX0U5eRnyaRs29sW/SfagQiwAVgwewLoOF/kWO
jPijFWjwuB+k3U/5DniFoZA/+dsr2ThaJ5L7UMcw5nCHSMc9PV+1gsMTR0pouS6WdnZdaGB2M4yH
vOAU9QbGtxkTeQpZE93TCg5UeKgTSij8n1vcm620YbofCsrBRt7WBLBUj4uFJjUH6I/Z01iGIIol
WFHN1rajvvzUPqTvea02DizTj4JVmMRTdmGCrJ9mOCzv2wL01PSGR7GE7kNZeHcTRZ28qR/59QpK
MhmwwJ8o9xpM2TAD1zDVNz+oKG95H8SIibwm7vnR0pfk3ujoCnwszTTCG24d+IzYlWsa1h4zsCcu
bqsSMmSALrhH3y9Muq2kopQbgkp8IG6tBLxJA6NUlPEvvfe/XmMA+MYXiBAqyG+opfPbohtxhSne
GO4o7Y6Rfjb46Cmyt8EsP+uNO5CkvsysDi3fLabusSDOJoHXpXE1blT+l2oalQ9ysWZh6UY2Umyl
xYNi9Hy5qMjONW65MItkFt/wg7vcj3SIMFWNU1FZCQrUjeWOl8filMyuV3NkCvgxljedazieL+xf
RO9e3afKMQcCh78lBIEN9BUsVv5T2n2eFhWqWWSR7Frc5+hK+KUDTQb79Em2ej8eQKEc0z/oHEU2
ncVNWh8eoBmJATevPh224NsQ1aS1hF+BbpgvIW9kF+ir2nwnQb3S8HgUzNxNuXZOOOuljGwKYkkG
Y7CvDkjpbn9fVJ8paI/FxAVyqV/qdZ6T3/oKKWGRPZ60OPQI1HhB8qORQcMCEn2biK8S15cbiMKU
qA2msdB7maTIZCVJyRalTobB+LRJ0Tdmyb89L26Q7GorfG2WrENQywDlMXH1LBuIuyIe8BNln8yh
NqNy1OQ0f15JIWbiYH+wleAgjPesmnQf0TAtDj8VHErP31YSUmk7tAe9etv6t8YO/EyUnJi8DAdM
kXllh66hJMNEdvU2mNnA5foQ6AhhR4iQfkSfhvdppSu0gXD+kT9ARG01KA33BvEtUw2jv1yKYWdG
NnudM2dsZBh8jRxVoVaQRmw8JDP11EM8vnNEPck+3cH+US7eHzRzwTb8aL7FYHky2QDcawU4Bp0F
qNF0qb1WOMeLWb+jSKmTDRozPBneVMEPZ2j4pisOIsdpWk51WvYEj7qKqyfix/4h9xrvUXS3mpJr
Fk/ilZY/o8ZZgIp7Yo32n97s+pMUXGpO7mqcNp5DN33X3gOsV1mbRt6gqKscpGSgMbwZXC+85HAS
xabOSXO8E6iYGCKl3bEhwcDxh5LJlHiH2bzQPij2V0/3mVg+ue8I+umd3Tg41ClSRYLE4snssc2t
Z7We1Swjij2Woa+OBfOFmGHFGomOrjta/nVUOOtCZ0EFGOlcFvkr8VO9av+50aVdOtO569PU7SBp
nsTdsQrSu6awl7yNDDYKEXsubiHgsOgmXJQVxCHesqrca/YFq1F6cZDpcJMi0aYkO4qI0477wJsT
DouwxH4gRh/rsyEOX+nFoQm4kQkLXV7wgRw6kK3UHDwKbuqDXnc6b3Jx8jBHqTnL5l8bgT9ToFYB
wImeXwa5FEIz+roVOdQniqnARS3C4tD/uoBviGNIT5s6NZJ5QaUHcCLQCILOFUFepRO2Kpv40fKT
otbmXrjdyyl9Vb5YstEHKgOTMQh0hbcIxahbGO5PNlI+qpB1uyAiJgix6SzUuUZvFpiydxSAAjAr
tfEybuehw7q+rp86bq3YBiCP8RktRS5AgpnmPr26ot+ajS68lnWitKbjDrOsPsUGZw4DGm2qY6yX
1TUXVk676HkUrZicVZxHryHVyv29zTaMbB/5M6xUIyWFUxY+x/jvqmcOUyHQU9JjYtQWKNO83Qln
HnGnHvVi2I5eEd/as7dcW6kLM6/UcyiD+2cmqvJL3MuaSNSiG3HeXdo42p2QNW2WN7XtOa55KcJ0
I7dI02fQrvjSfmqXcmCJSyzsF6W/vGLyqc8+YVQxBc8IM5zHPrBTHSIJrWtzHL/CWi7QoRpGjHMy
8cmEAPgEFDw7dtR06dnesXjO81PSRYOKw0t7m9vhvtIZw/T7bQ7q60nZ3ZzmjVYA+n9HC+i/r/05
M7u05njsh4ea/XAmIxQ2m08LhqB8xCGCk7phzmCEfrynbw07VKq2NEZhZD4gDjVQeum2EFTTj7Cg
VyoGe5UdglyhCTHHT3zljeyjvoYPVNqGLlovWMcSDRHsIpF7bKw+M16BaOTebgi6bUGhUyqnkFRM
bHq/A9IhFdEKSJnQC/beFenw4pmNxmtVBpPVBBt2+XPZPNv7Ud1dWNQtNGuN4uABb/dkbAYC02y6
teE3fbP/smQ3OvXPcaHFg2BycFMzT+ESs0IO+Zf6LFmedMF+x3SjHgPo1hccqZK7E5QRxRDuT2W6
5lRkytxYiJ+j6K7zRJ1RYH5Ty43ywukdaqlcgjvdMHnA2fejhgP6Qx/DtWocFl+neDPFliY1DnOI
ZdG59JUmABbO156+ZHgDsfJr/7kMWLzZ36bOXZUhKFjx8bvb48zZ/0l09RGEf4k9apo/wikXNVRa
4OcJG9BMNYmrJGWaxiS0T5TApaqXvnJWsfzXRS8kKr72h3mAxxDmMhZWE84gEVJL+IW+MQhO3HHI
dz58bqSwzUz8iXrfkCCLmdtlPY9BXAnPYH5ug0aZRAwiHed5BdHVkPruBUm2yOhE4b6yJsTnk6qm
P8SDI34HHO5UiDG8se1Z/bum9pWJ8IO1/Yn1f69+xXLZLa/jH5psYsT/sPzR2SYCXcNVEd/vpGf8
qSEr2flHQmD/7dvt8C8DqT8ZAbSs1YedxHlHJNIY8WcOm7F77aX35OBIKN9iXb8pvPx8Ttu7sR0X
Yl5QDqQiF08VCnXWb6XYJzftbMqdSgUL5KWbAjzVqrUl8BIZ67t3Eusl9tHBJbn/PgVLYj9BauSW
paZ/3IBMNhPL7zXNx5Yo8Pqoj2WFNy1oJ/sB9wampSvP/ro1L0dg30+cFnhkuPJOfOpg3eYycRV3
Zl+Xea3RnY3T3jQLayU5pajfE0a50MZ9SRL7YUT9DXYTafMP6wB9PUuU8emZQszY8YE/1Q7aTx+v
XqOk2zLaZ2dlkh9ylLAmAe9cEWqQyaFdvaUgpnaWKqUZpgm68jN/yskeIFZD+zTZlBTjigH45hw+
DEVOR3JoSxSSzyL9MiMY3T4/S0tbOmalGkDyBdA156AofFXBs+OxQQh4Ki/vKKsOcaKRU9OkD/OC
bd1sdXrZIluZsgFOW+bi9iR3R5SLtkEeNa/lAmrEzPDJYMLsK9HM82kjXoorI1e34E9kNNK0Du3z
+iWw4kfV3RKkS7oqcHmf3Afqb0oku2L6osb7WF6peckl4ZPcT+MYP+JCXi9XkL70P6vgRat2a+qH
EOPX1iDFBag65Xhp23QKGCkFhl8AYe3ISeZBcTuRrqt/FeTcFgTTw6vsA4KzkctKsCRBTgPD8q7K
CG4F9tQr5sL8Y/Rfz8uZkpyc1j079tidBjk7N+pzH1mvmRokrthaFto1sjbSJNmsnYTYwG91Wy72
VuIvLfcSkTOE0XNeawwCUuVExaus7TcSl7+cjLIQl+fgnJil1yZssNAVy1xklFixGtf2dFc+VO4w
APgyKVHxr+DVHuih+9GjiELDvV5K+KmN1KR9MzDXMVYEPVxh1KbQ6mwHmm3735zJbi9zwp8Vddjs
8Gh0XL03UFkt2jJT9IuXd8HyaYDf7QFn8grtIKPeD1IK08LesakrLsNpYbW7DU26ENRtzoyac7HB
3lMlvOVOiVp3rwUDLDS0duNd9wvujJFS8KFJv6n9LO5c70fD4WE3zSSXCIwVw/FlMoSNfJvUN7jc
tSlTHcavpS1k89sLH38al1ew+l8qkVC7mk2ZAWZThyWC49eiwOZ0OcZXTcyFdkz7HgTRAEhX3sgS
RQoqkPuyt3CUZWEDnuTrqWqgMqWKjebXwAhijY0I8Ts3kb/zg9rkeC5CDv0yTGjHyY9ZO6EI/Yaq
+/CS39cgufQkppDfyJpFnXqdPSg3RW9DLRuAPdUfEevlrUHVDEQ9nPGWUx9RMEu48Pbh90479UHj
J6NelBv2ShqAQNDDkcPUdcTbRrFFn8nPQO/etUlOD3WxAjWYgyS/xHAEUZqgl6YZxfzOAOWKPtVd
E3y41alSOjSZ/T9QMG0KYzoS1p1tl4lNxcjzypHRQf6z0l+3qnDCFx9fpqPC3V97fFogLX30WiV3
REQJ9OfpbJrJSiS+CEKYagRyZy1vJrXhtelWeTw8E8AjXqoaMhPWG0HDt/deAKqAp2cmmjY+k28N
YiCTpxg6wZ4JLaVlkalh3+1Z8g6A2EVIQT3528NIO8d7zlJvpyom/+u1o+Dl+BrJVraKkgT5rhOG
eXIuon/meEjIMk/MKWhi55i4gaTnlxopErVwHd7gPKEbTqFzHL9GyLw3r3SCQRNkc2mbNQzaLDKe
PptAoFudlupIyTSfiKNbizr1cUn13vH8c8ibE6nV3SWYqkeBOxwZQWJocFW9TmaIXaSnQjXE4rn9
JUxLDWcBalrtA6jvxPktFTH1xq4ngqFV0X9aeYaWVqj9ukjbXbx7T2NOvbSaH/CSFAiWS376yHN/
2r8ttyo29LByHu/b576BjXMk7XlFjMNsXkNzPs2Mv3q7oNMHy3AA25f7DzRRSrHM/rGhcoa9jl2S
lE/dF7H1ZWxncz7dFYOcwLKxSoxdnf+aWHAkvK62i6BvQWvqLuheQKxwoi6JiCGUUW6NY7TB86vn
tQVJo1deLHcWrlACpWeDlaFJdJe6Fcs1/3AGAshPGe9g+1xbifHktCkDIsHW0NV4Q9ngIbRGUC4L
3Gk+rrzt65FT3wSm+QlMHbmSd8f7bD7uNIpezwnJcP0GWY044sCiRWr7eMTPKgolkedGPVt6NCDA
9JOO7wT6Ki0oDbiIxGWVzFV6CQX5B9YM1U3oJmaXskdd+az8mAAefEFWQPsogeEOAENiFrgeTzgb
Y4fsaQmCnehgzb/du1vSgZpcFlzQJ0LEj4xwcRYPNIocKCmplwz0YyLh7bz9zlnOObwzT87KJC9c
gr5IlCMdAN8wQwBHl98kTJDciHqLZ2cOfRat+X7Ra7NYAkPg8u/PZTJJVcg/nrOwH/QBYuxEfWbT
xV86cuW6udHbmlHW2rjtXS7FOSKSJqHzWeYdSJuvuryZz2AyCnWBDvy1Up34D0cvB+9tToRWXvPG
r3ITP8+O6uWAUnYgNVk/UhS3TNLvH6ehNR7pwxoRTqzHWGdDvZ/9ND4EKQOA8heSvRpCN+pSWWoL
JWXNzt2J7mY2gWGx7Gc1DWM296zjaCdGzImd1vYCUcUNvWyf7ERu/JnuBX6hunKFo6LipcSpbX3m
cCLfG4fUQA6u3+AaKNaZFiO59zW1hfMRyCNcs7hYMoXPEeC9mdf2ILOk7akZ78mp8jyerbbXMOS1
0g/kod0VG18R3Jv5ecF6qDDVidfCXfd2zThJgGsqFe0/Mfu95eZPzI7yJJiW5uTxhsZl378KWa0N
9rkaPrMKLr2ID5Bh98YskvP0g5BAtetcIwfbRwVGMnX7qhV0P5ai712hSE1N09J8rhVcj2FwkPTy
YFvQWC42lQfF13gkg4wi0Y3dIP+CgPqY9Ap7VLYOTSBOb8bo6gk/+xtypBI5vUXqkdU3VdZcmK3v
bSxUZzrh8kqUhUbWxVzvNodSWPpy99l2IDN/pPwMFefkuBMpFJjNqgpcwx1QDeIwStakqino6nEJ
8hL9Qz3pMbMk1UOBxphlt7w6BfrC5XHDxgRPTzxPr2jodO3aLCUUgADH/jeUv/1qCxw0tc3HErzk
LIgqk26vp9zL8wZPyGFOJ57F1IQmXbDv/6Ym2snkKvYn+H5Uixv33D8+OKYLhzumO5XBgGiHKONf
itk6Z3B1bbWQHjLZFdze2A+sGdptMKvRTXJOUjfDMb15eF94z+I/tNTd+RD1nlik2Zj1Luma33sP
uOayynuPDpDrFDYe7E2wHXLwAUvfCShiy5AI9DJT112dFJeWdlSGlXRG65taTLO4dnkrIlrnzGSL
BHpF+lJE+PbWuPkref6e+7OLeOapR/MskXsOmZeBdD3FySQDk9aQAwtQLkD7VhdntR5fs9aws7q6
SMrMYD5VLNP84hG9F2LhFipcQrcs9apdRF47bumrcZUygnJFzUgXzOiAjANAscdOArkDlZJPviWv
3TJVXX2dhhPb7/VO+l9u1DMnHhTTfDBnYhWJsJfiO0F93WymVS8+yhfKraYnwWc30YaESQtyfnbS
fXoATJ5e69RcGxSbvsNArA98ej5VgX+NR87J3ID4+sPfy8i2a1c0ObTMr+YSAjbnCcgQa3pBiGre
I81lxbm+poJ5COJWaTWC/mbhvPzx9YkKhcaBENy9wW/5DHGEMlQyJoPNFvRzJeST98u7ZqxUwu0L
dwSZGbAhgvSoRoRXDgE3a4mnKUc1DdKQ0CMcdW9nlah9Z18SsmD2QHLtV7Y4zpw5TIbCCENfex5i
iU7E1g2ewnXpltD3fhhRmsyEt34dGFPh/CFVUJqwbRpVglQKQR9bwSRomX2Lw00xkXVYFhOYh6Nf
LtSyjlT38qwPVQx8+JcDTmRJIcVPKUyhlzum7xBy+gW6JMIFNhbeN27dh2gb1Pj+0QE+AbQsRWvl
Mp5HPqJmv8AIPaHwX8Lcwv/S+eTVEbIPDbWaktL7gxLpxG0MMYwJWMm3HTGZl+FTG2cMKpicudUx
S5dOkswTaG41Ns7m67z9CK2tRUMzsuVOkHalKOc0ADLywWB7YYKTr7lLQSR9JlVBx0h9evlRNIfb
ZXmNmPxZDrP4qUCOP1Chr1D47313Rt0Q9n8XtfAxjGveeFgdcq3wxIKGYCkT0/OGey3/ZgWP6H+4
fm8xw2IspUWsMWSy2+46f073R/iUtO/vLBQRNDhhryGKbg+uqKbFS5fcBWf2PKlLGQvAqzxQYBVU
XqnDJzGFooeh3Ya4AD1jQ92Mbm6dZ5odLO5dvI0AwA1gtSCkCeh5odNat3WC/UuJK7U+ciqBylOS
V0HSAId7ZnrqHHMS1jnHABuJaa4HKwVUf3UdHnEMYoUiurLypIKqyeNvrVLwVYIUfudGFmGSM2Zv
dTQPuowxHmVkVmoISZUxutehieJAgWRbRTVRKaV1/oleYnVU7X634qsCONZ35f7wOS8EEKo9bRQo
82RNQcFf3ME6Z7Xv8oqxbvhP4WUBhNIOjCJ7obv7prYXjgxfUImFyWjp3jyKZS6Dy+YaP+Df78WH
lrnmWO+d7OpCCLlQ6zfxslIyVgKxyIxxkmI7BMLzNbKfhb9uk7VfHodb1O8sYZ02y3o7zkwtyiAt
4TURJPD2NTwbhNHJnKeFOfZfo5X86+Uq38MsPgajKMZLscLIp7pkanKymcL1cNvNXSWEmE3HUGYN
EWbl80AKQZnTYerr/A8f4cjjBVnIs532GWUltC+n81xmQvXsq3jmNbbNpxDvTaSXwa88GTsnInyz
v+NIBCrxeHLT9w1Itrq6t08i3n2sNypCyCzZZYkzULzMzfzGOxUV1yxmU33MlIgu0G3bVgFY5lgO
2W/BPK92xY6LhkXAFkD7O/WCqL1nbiNVfFHcyCkKeHyet1xyrinRja2x8l3LPvdU4T+TB6MRtgR5
dEnS+N2j6ReS7TZr/pTkbkyCifejwsXEfvzYimKEyiq528inbNWHV/v1zV1J6quhXsXGOF/tew6X
+CZ5cvOzjvno+ktI5r5Xd1Wz+iYciAIzWtz+Iped4alQnetEmGV9IuRy5A70qIL1BRhk1USJrMy1
M3/UCA6YCMGexRXG2HjPxv4PEtP5yZ1fSnXjNBgY2cosw0r4TtTcdGCCRWBG67BPYRrLNMttQOBl
/JFF0CP5p7gu5zTqbGOWOXO2LtpZhFsah6iYjg7klYRZJFZQj/Tjpa4GYLTiUkJ6PXiJ2SzpdhyI
iMoxtE+ENFuXzOOqEALCTI5ScN2pei+1J6bR6+ECOkmgpFn5352FqkBHklNAeHmyRdAXS8+jqFNo
8tCH99oC4ulHXXa7GyY6g/reDN9FVFcg8/EtgvIG10iK8Iva3u55+KDb+KhvKYwIDhCndrs2u7HA
gMNwAThXHOXMvNvhASDMQlyu1tHPBpD0eY0JJOMAbq129ARX/lHILxhBczEfcGN9h3igBJXS6aA8
BMcD1FxllcWcpn7Cjt/c1IWXu34S3bH2VRwyQEQKq6RGXip53wXrZDtuD29Dnfmsnfa2+tHihhMJ
79fT9mCeAoZicbJLJqf4zkSQH1vmwkWSjce0ApB9FuPK/lFou5qmvqH3EvtSamD1wasBk7FT2s4A
WxMYsvPLcUDxJJZS9077ZfZ2oecQMwsvJj8JSTinmFJn7pLtFaQInxX2BEjtrkJ+cCWQrmBJyM0T
0raoORUZplkSvbfAftilSbqTWwnTBTeXTdoeM4qsIytjhg7OFG7d4v5T9QvpjfXG+eWyrF6MxeK7
wVsoaqU+1+jM6pYwwtBjjD8uCIXRo+I/BeqMMEXmSDHPkFRbfq/qQSMLSEKt0iZkiyjK1MOKjzG7
GHCtvV710D25z8hBNMm2DDcTmFtIEe7kHKriPvVMlMEUlIBjqbyL82R2a9BIAaNiGDUx5uDg+XRI
/hjjvJT/ZZbohJms/x0ko7rQ3ZsqoTXyUBmg9bOluUZ4w4gSI8ecH2MCImJZQePq7UcMw6QExWR5
IBO+l3PFoyql9Janov6/2sLRfXxLqAOmjH0UBQsuNQZ3LIMDL9eqtoXzYOsNnos/2lUYgDW8FWCi
9vbW6FJPDMh4SIz8EUc9dv1EKxXz9mVh7jgc8NwPFMy3k/ANXvnqsUolmBv4CeMM400+4EF524jj
xC+Ro3Wem8DRzmbQ3UxmgLw4GIchRfDGpEVMK7jkvC5xEvt62rNU80oH2sh4U5uSqspeKbKe31AU
/0PqXEluxgjbW45K+VcqyNuupDiKW0LLYWu1yw6F9vs1BIQS4ZavR8vkEBmekuB3flfPVvlH/io+
s3hvW8+C20sJK7/likcAV6q1YYcNSe38p3N2KvFt5LjJQQ2PuAoloZigAo/F0Z0RSBaQFQFaTDB2
tRMt0xCEXp+FSMr94plka8CjbGCwyr+AewPZZmdR+57+lz9sRiptvIF9feOYMAcH/ZGmpFwtGndU
ZmGG3hwX3TpW72fB5g7OmJFeEuHx9Ze+fvlZ4SGmDCmz2gUwE36jf0F2g/mTMdg+OIDupKjO4yoi
v5e4c/ONrUDUVH/p5KH51dvazkXoRXgcidl8qH6U1/JGmFgk8ZjiSkFtE/e3cudHqDBOUE1Jw1E1
D4qePS9DlXJVoZXpq4tllUtbT65V7NoWIsFU2ywJ4OniFvl/5q+7hi193oa+919Rg155n/LyqoED
RwcdmwwyfWN8+CmtWkNNd9d2ONtyKyoWr8K5mWrV9HxajUZGACIbzHwnXZV2tjm3Km5lVYdn4Wj+
58LPVX+Qn7UO9okLNTWGcBORb3tZWuyyrpBjdNG5quQb4ge8odKizCezlYnuVmfpEvb5FwGbdYy8
eJlpWprZC1PlcCJn2+4gXZNe0iO3eq/u4p2GjUKG7b2Xnb+pcZm3qmCA05s4hxDv4MMcv9OjzMKZ
pPtZNWtpmt/uQ38PuDqnddtEOdRkM5p/QyXAmZVy9Jcf8NNFzfmlT2TtmSVxJvea1y2pfwk0eYZj
jt/2n2mnocubnt0mDzjHIgH5dkl5LO/sH7/ldWu2YdAW2IZQph8EVzWMukyKLNIpjantnJoWRU1t
tkfdV3/F2aogV+xqdNB2Umcst7TzQo1BumLC9mV3+PHqaRLCyQvwyh46TlakcMZ/gohgVnpSEyKn
S3E2voz/rduAtqVBwRhs4WGBk+709otLPmVIp4Fw8gs6FI77Cplexb9yVYjQS57aS09h/Hyncf5D
6KHEzarhXEfQqQD2O3GJLyx+CPP+zqVQ7GsneWryh3SnbbnMrLrEtyozx1OAv98AhBS4TISDmi9I
9JoaST0Opx+hP6P8I283+EX/ZHPFkNEAyPIsprTyyrHCaMqW7UvDszZWZ1bsJkqXemYhUsePqHTD
nuGCCDqKQaw85M8ivW5WOGZdLgYpLARmET5++jxT2/vO2OR10kir0ezhqBNQcQafTYxhwKlebSrU
OlXQnuGmpbud79rSjceaO04cJOTesejWQOxAy/EFdXSN75CeQ+3LmUj7ttQjtFhTj8mfKF7IbtVK
vxA2mA4CQG4KUezOm3dYQ5LbwWsuljIAR4t/4Cqyk+zjsCJi7/DEcR3qPJAJVGziWSM8N2D7RiNa
CDpJ5y7HLqs2MKZ3LKP6Xv0qhBtzGQCRg1OVd/J+GIem8k+wMFHLV/3B+Jq0tpsFn73N7iM3+gmX
odg8w58jIQB+N4u2b6FqNUCiwURqVctpqANNAQhDGt0VhNfnKnMyue9DuxQlAOa874v0vqN8krJw
FMXm33SZ9CwVcBU1G7DSPdF3onzSZW8BxM6bwSVvVyp+y8CGbgxm2mg69jr/Rof4YB/N1LSAK/LZ
vAD5TPaiWQ0CFvIQd6I1y19zNKEOUS9PG2NsxiNYurhCFFiyQW1xHDb5efPIdz1QCDPrhxsttssJ
ziqR6oAci0rw0O1qf0/Yf5u4KwZfEVKzAD3EfFA2L1NcH6o+AL0acinIV+2pfom99VgQvduu0bdt
Ud3WYMsHlpcDoHOHGQhwvP2eDovDhaWH+jKF8qR/AB15SLpNV4EkJGn9EwiqBEXdZUjh/I91/uch
uPzYcnN3FDZDAzbWJ1I9FTN7wSzxRhKfODEAafsmnBBjDvn4yyNRCP7wgT5IKBR0im1noowpbtnV
8mAqVVZ7Fx4vbCwck0zeSGaXh1XpXvjEJw49gKtpHEZouW+oZK/JSvJL/DC5fbpWJZACYeMa3Iv/
zGYLiDzo8QZB7aWQIoga+pN8rFo1yEAl9D5Zi8/G4UBpwOPO4oDdSJmQd1XWkDpqmyPwcvFQonp+
4kcU3j0lb8rITpEI9Cd3vjXJ2Rtx2t2CHgdFuayOLKAQQnK7vmwIZhFTZ9oYbzyoHYfCoa21kZmj
pQ5c+03O7FDMFzZ9F5N90Z31GBFgTRb1nCHWWb0c0/1RWpDlQ0pA4AlDGwzYEeDyb0FBMoN4mMWQ
S8jTYJd9YJVqKN5JAp9eXs7c4z3zBiNLQEpvLtErUzeog1Uy9xuggrlu5UfEQfFrNL0O7N0ziXWq
dZB27JUXzx1vfjoM5rQXBiQoF2raeM6EX8hpYWpCcQnKHE9mwSgtQ33/sA4h6iHuvfP6snkA1GcK
zcZ95AYsdteYa65DoG03eVmjg43yP3zo0TIGJ7ym8IhTkZPrsgc9X/oiMiTnTZqaXryWSLRi1HaM
9f5xgugJFW7zIlScwM4HJNyoVOfcksikQGCtSXap5xuPcq4CjIz84hXCnDU69/XaHqSOHGeqyedz
MgkHNt2p1O/3XhL15uH1kDWY9z3/lf+SCYqUVzA0BG7HnzryX09Emot8O2xrbt4TvW62tvbIZeaz
EOXCB+gQqHO6n2jX+az7oxH16y8Md33+U9SLVe5zKHy+x/w0Bh2PPC/tzTMvtjvXZ78pf0WUEXCH
KbqdxpxXqZ+pHunVGostUl+pBuqFHMK99IStq464tSwbif3IvDKdNiN72J1jE1dnYATMWociR8ti
4zxf/JQ+dyxepxTc3uqwvZmReiNc+2RRxTwa1euHhxzxxKSn7520MYLMHVnHviXcKhMJ6d8p3/jD
D3n+jgokoOJ7JQ2aseCo8DHjZQa0I4sB0fCTBJ8U993m3tFfmprXkV+6YGa/SF8N0hvcOj9ayQoZ
m3xqUNLz+50M9xB1jgawB5Bgy+038I3CXYNaphX1RoLz1El1VXuuWQmPOKsTNVUXm+FhnZACdsuj
36Rrm8IcoNkD8WitiF0m55XYxAZp6n0ZGVjfFviPwyFTiUCLFnE7yvUIeVMBJZUtClOZx+rPswih
Rdlz5Jqs+ewHOxxExxqmgXqTAZ/8BouiYrkr3Y1g/QLu9mWLmdAUgFF0f/iH9yFNXHI44WR7bQwr
KS8RXJ8z9uJwMAqjlzzqsIxZJdCgDzw9DKagTc72gUqADSGbP6uEds70ZRkjYFlcx8SU8L/TYHOZ
gvrNHjGnQzH1hgmdutlMPzd2+rEPDnrOY9tjIxCvqs/su+l8o2ERTkr5wXbn9+qGgZAD8IO6mZsC
c3aGoKxy6rclnlR8VDmk25edq+BdEe45l63Y0YRPxHNVsBkzPN+n4hrDEdxLj0wCqWc9Q3bLE4Bp
CGQclHCsQbiaMheGzpFEvglLhmNQMyOe6RbAS5wLEYEoAbt3XQU9XusXnr38BfSvSXsd4txnINk+
byp6KL2GmZ76qt/3iXE3nwq16oFa5MRiNFl3Sad9fFNSI79JQ2VZODqcyaYONqiussFxdJOQdv9m
sXDpbVDmEGPauXyfEnGnyFajrng2lc6Vcih3wiPNFCG2CuhqyMKyb228h3NIPJRMwn/o71nc0ddi
0ob8E0U3yJOnCKCRAZaUbZnz0pfT55UFtOiuiylwF/hU0rvS/U5NSWFCtThKRK8JoLFojWn8JAHT
CGFw2YqIaVMxqxPMov0DzoWdbZYre7nUReXIqMl7m+5Vy6Wn3CKYp1A6w/uVuen0X9X0U5rVMX71
THjP7j7alE805UELz7yaRLFLOKGIXFk9+Ah3KcOIVuUxvlCwX7ZQhcFl7syFeYh7hWgIllGMNRwf
8PTBfF2tSM2OYWpd5fGyN8lkqbLkf8Po4r1MB1w8pupxjJkTSM1gPJntV8E8e9+igtFo49t1eVqe
HHMmSDU7OtJ3UOVNlbHNRoeF4GodGkxHXzIHdpoI5kK12wd/Bkh0uZO2D/tUDEL30AA6Vu+q2yUH
Sttpc0N5I4/eAQxlgAkunJrhFwg8RHBsxaDZb8TrJEohcXZwrf9OGNMjsyTlzWwJu81P8HaE3v7x
6kY1C4HlpfcCgGuvCxNjCyxlvvVi9LUZn4TnkU0JpqVOusSB+AATr8sosGYBxvdoXZd24UblbZmu
jA7wYwAKeuLdFhMkv1L46TQRKdkclvsaybV5jMBx7isP+61prrUU0NEAkQyX9XGBrR/+sloL2Vex
S+QuaQba7Uk+mAQ2yVWwptBkJszoLwsriI6yWnfDxsYfKbwkY2XL7yIEXpW7fhnxpGZG+zxvGzNc
Z5CuegEdgcPCGbqqDsahK6SQIpCWiDj7+bl/vgqiBipGFzuhXbmwaA4XAvjtFGyeP12eIomv0eaM
WSFXYG+05/HoHbU1Bb/PGWRW+S/OfkS4E34jPAO8hFfZEXLwsU3j30KHyNMspr0fC3hyivXu9/H/
WpWNXRNMU0hfMugq8V8YTMjrYVQdqqbhUsWSqgkb8cQmDcwH/b4j8gre1DTtLketWm1WWFi/n2dl
C0etM4M78HzwW1D6EsSAkZQH9yOO5b0Kym9RrxpOtgdXcG25X/O2nCoU6igVK3hbIZEq1ZH4thAi
0HCmxWQwB0njc9luIPK12xKGb0r2JA7XAhZs3hLeXXyfRQyUv7nBcGLdgqyhsVvklAqAtHvVQwGj
06fhbPAU+ciUOttjZj4cNOC8ECQ97ll13fbMxKNATZKs5kb9oMoTJ3d2B4WAbAX/hE3XHrJ7f7Hm
Xn7xurULv4lTpt7NfAHp8cR1Mco0t3kW03T8L8CWi0DNdROSBv/Qq9dl6XJJ5sswMjRl47ZbKzbK
dYQrTPEAil2vJSdZtmi54/4CwQWAZN4dNZ/v7z0e+dN/FqtZprikJSi447m55Qzr74VwXdFL4WpP
GikOEDgJvJhLRzewfODo2b1+5pBgdVKLEqe46hHELDJ1/IKKa78oYaCXZdCKDAa/4E6ue8RA1E96
cx4NdRonWGAlt7wGX0XNvDhVmn4hWJh4a2WGyyLfA3JU53iRlYNM0w3Twj6O3uXk5kKo5woMqZev
ey1xpdZrxCMcK+mIdplX4AIxfFOldzEvM+CgGlPSMZ1Oma5GSNd7RhFdFFC7s6m1E8wBRi7gAxsX
GCK0Rx+BgRTU1lflxS2NAMvebAi02Ew1cDasMko+5ooK6oUyngUVv0+iBRjysPLaKI10aBFHmhT+
9M9sHjpvnY1j1ygW84rzg1xj1drwsEWEz1jsjxBKvHEl1wsSMimwMo78ixaNPd+ng5iY4NeTpJHh
hueixJwmnGrqzya/cJwNautNRyeNg4V4FEvVEU7+xu4EnR0ARzBSPiJtBLykdT+G97CTjftop1Wr
hijhyNVUd2B9Gw6ozbDaBCMAJGT5/AQUUvcQf44w7/y1qK7z9dHXDxHhVoj/1stOsh02zvDl280e
DYUOUloIyRWFJspoey/5YOW6AgBiEqBDYUZlNtH3nGfbJP4zjUlFPTGwNFuBvMa/kADM5TJb4kEu
pM4H99n3HvK6MPZ3PJ5VeLHQClJXnEj3C4LGm/j3uqVMt6ZAkPKmbDJroYhc9TxIZ9cyEUpPG3V/
M7miEmu6DNxLdbFNdzLiMQhMlOUrDZkCqmYIC7G7Nbn8RpJjl2VHHUuznjnOKp4+EEIA4jkHyHFQ
8FackNhQaeeCBNFX8RCDBRqEotDvA7NMj82QbzA73KbCpmwfwxginkSbN8JNV122cbldXJUIKFJu
wbNvDM1exsQHBjPwZOsRado8ir6O8ZziR6E30kRhH6hJ6EdY7dYruQhl9dxhOwROqHBIDt6is1vJ
EVD3DSuWcg5XdNtKLpNEM7WzZYo6/RiuHh+wCeSZ4hv92VIaABB4KvXgbiunKe2c2omsQfTLo39T
RCMPyb+jW+1k/DWDzsAsHl35AZdxbfc4JxcnQ47nNLj0TogPSjmn3hqyO4ZEBZ8WXP1J0gANHrZs
+CwNslniI77SaqtwRY3Gzzk1vWzE+kuRMSAs9xnWZWo/qRE7+CvrDd+AEmaqJ75TvyG1oG3NdlZg
wQIeLWOwKnlT+2qXa1UQbF+6asfGAHh4eWk6P45noQycCw8ylYdPmfTvB4bIwFwJ/2TUM6k0lkHd
v4wJ7l77ZF4wXRR5Iqt9z5o/Fzscodw//vcsBsMJMSKSH0XdL7erKEmBJS/IKVMmz177Sn68W/M0
HLZuwAczzDeDdNgF8nc3IHHPh2aaepyOk8dkSBxXkSg2kMIK7Zctb5oZxRI4urP5c9ne0q5N3K4H
/CVLQfozHKDLPURUSra7BIkODqdYmD96Dfr3DTeinWi4XmEIlognUFgbafzVpFmHpUJcaOW1nOwD
9HTSqStk+JANEhsuzBuTJ6lPKPbhFXneJhYcnvM4e6yOz+c7XKErPZ8NKxpyX68POhdgmPMsu0dR
8BPsndd7Ft2kxMUfGuMZzESy0LYvH0qMuf/bTBWBd5M7/7RqSuYaXNNfAxrDcEy+CcuBDTAenBqy
N6110Vprzd/xaMr/ygbJb/R2wJ/mWC0wPM8Q4cOtLLwE5RlXaz/Cx9hQvlFl5yB0JIDEJfPspkjk
N/r+v2FoMW01Y0txuTsS0fGcX2ZV+YAPD4TNsec1iUrKVM1cHMW3A2BPaI3T5SL8Ox572/gMuPWE
8Y+Vqy8tswaQVfi3kcoicDIfK2h3bt56t3lK/gAflFAj2CRAeCPLwP4rPh7ACwm1KKdgSr0pJgUQ
6U2bgiqIwp877xIc1y0FI4TTs/17Wnnev7/WqvcF1E1rEkmR5OE2MB8gpwaBWbLuL9TNhu+n8Cpc
9TLruP8btciGejs7tGtc3Gm5q8eri9uhJ5zIQBHzcK/xcuVJcwr9DkWBlWAZmiNWgPReEig4RcvM
D3pDcgmipSCFbktpM4wONgkbqoWUmGt2U0GxDZVf9RS5Z8z1/E4XUTztvo8/yTNY0Xja0UwmzcVI
TV4lAD6vQfllCoK97vmLL14KUKdldbi3cGSKp2FAwC5idl+022LWbY5yXzE4BPIjVe/ZtRAViMu3
UTEQxMmhqHSz2nfEjHxZP2Nh/rTbi7pHcxcQq9OkybIJMVkXxCD59LTY71HoAZfjnoKH3BoQ3XVQ
Sr3Sszyo32hH7PWy7AeIRo+HhG3sc4DWzYSl1vXSXJgPdkRriyRx57WKcuGozyvi//3LHJWKCOH+
9Y0+A8sVZf/Zxu8SNuF0x6jyV40HaEGYLUfHjcaHZFvrCloaPUuzoOjIs5h0y322vFEHaRmcFU2z
58pm931sDZCugdG5HXwQWCEQYscidQNM5bAvkHMlPqbKYmyWDvVX+mp7cVNEj8vzopzotJHiqW/1
wf+rz9F9tnWwjaNik0XqO8T7Ix35zDls5rzbUtcTfGl8ESn19f6KsI0axoI3eW7IHCRr843vPrcp
fy2gvKVfM/0nP1akV/3EDkvWCw016olLtB/nkIfWgIpWPKQ1rvr4PyKJeIcy5w4uIdKIfuGjhssq
9XK96mO2BEGDZUoEWN53xd5/FxiDMIScuLD8pxPRk02pDD8z4z//FBQlc4kTgb2L2BDroQFVxzXq
ka+QNykEeQMWg5O+196nR1Af3Hothp87sdvYwGljXG9AdjkN5SHHI3BUPmO6Jpn1pG5Fq9CuqO9b
VVEqJq6yeUuvnaCawUvc4ufSzXoUhEovMrxDQpXT8FrBrUPVWiLJ7smH/8iS8PWNDHCxPVTI2+KF
zeh2KXUF0HlfRbfXZOlzBxIh1K4smiZvbfF3OtHWz/E6E2bE9kmQDvXf1DIiWsCQ5gbtPd/UDrlG
MzQeVL+SjfzMSyJLCaEZZOMg/6JLmS+bWaCI/NwRIb3OqazJhji57XdEpGxtb9rGJvqZCyFsjpQd
rbe148ods3YCRTrjxlMJeDrUNcAxkZjjcyPZLtAqzl9IuCKEz83Zj7FcW7X8ZUBKl8Y6ZQzADuly
AfwTQoaaHl1ASldNMjflnIZfAWFDUe2lRVezewGXY7DJT0u1cYMyuUgpdWpyqANRPGRpiIrdsNBt
Z44gaZtGRZ9VjqWkDI1C4B4zg407BRVAuCKWLw2F+ubRbXr8xAeZOZiKbr3niGUFQzJznXUIrrHL
I+Q8UmqbOearNisiUaGE3M1ZF4YWxwHePG3js9yJcLLKmcTfg6oVCnqHAWLhCmLkYyhM1/VPVTpI
T8OscEUjBEgQCy0B4WCQFPugG0iULfb86zAOll+0AUQBTxYAu3tEdQRry5LVTx7CFPuLhi8NX6XL
pLBz9Xb1jbmwBzZFGTzlmCf0HlJNdBCHBL49Kb6QUnv5oxoSDC3+IXpH5XweGbIxJoc/bAX6Dr2U
1kTZxJW1pBUx/yHaruQnLT4OhCgly1NLtpeaW/IJZnVpp4ZhN3hbrXM2+r01QpqXhDoe/oFEZN3Y
XPmgKMNRKgX/VyZdap8JUEMyIsd45wFMMrb2cw4es8t2PSSsC8WrAEjl//AIwIZ2ErDlsHCvBqpt
cSsP0eFsUPtszukgH/P2jWxtLO/2xpfGRqANi0zGO4Gf6vBi0rGmkjAoOqjJu+TzN/IPQfYSFvN9
SwOU7lYcZrOqawkbYwhgksExUBcIvz/7b1OtXNQfl0wWeHasVVesAIHFUUs23yrxLSAAOfb/TxVS
tc4BDwpdnndjCNvcbZ52DIlzhSrh4lCX7hRyMRRWjFdwtSJmcdc4JJQL2tzQYt+N07ijD26i0Ml3
lQ9ajuUhFoWHJ+e7lO0ds2/S09fmhhd+JVUMUeB3iPoDVefJ1Hx44evxLYMi/wDbOVcOCwttkWzO
ZV35SYqLKe3QNubuQWD1CmfKyOp5b/OjJmrgeQcv9g+ByloqiLVyJoApN9VOMDsr81O37+uOMLCC
UxrgIY4j3NRKDRCaiUdTsHlMZgC6P4w1SMBTbk0hePfgNg/L7LYdL5xBK+M3tqQNgkQt+Ovkz1/a
zCstmRA9kS+BLqbzTfoS1IIdVxAix/lXW1BQuHVP4neBGQQwlBUd3QCDeZtdok8zJW+4WrAPCppg
pzVvuSY4t+8eE1XnVKUcygma++kupZTOPcGoXQcWM6YYqaYSrO3D6atcr9knK0QWds/BVlaH+YXd
A5HgW2OnRl82pUyb5vsXgGbwtdPlHwArNDYCcIXIPcnzh+L9H+RMlwl4JAEA0kicB0M8ZQsUz53B
QH1RWnULRYJHYu3ZNE6vt30Z/vaA4RjRni7A1DLTIt98BMbVEujd63VGb82sCXDlNZbEPPHTYldQ
Cv00120L3OEMsCMvc+o8RXP7LXeo8USMScn20TB/SzqaNNAsKMrOuYU1Of4OW93OXLkPKYs7inkn
rgyXaTgz0UQjO4vRnxA+5HVAu41zb6NkBX7nSc+as8pUMUXaDrTEI0kCzjW6S14MhLMiPxGIT2r5
wmFZLquknLOQLdPOjVfQIgDEdTT7/k5oAWGjt9UeZtNSuW3345jBcDNQ7iYH3cVYKjWfTHXtigBB
ulPxkXErPHI1wmaLrQKUZVdHEQvGYiNb5EMX7aTnONETSPZaybuRgp7efv1TAMhP1J1Ew96hPj+C
pvb22adywrSA1EcFlpRrOBrtp6ChA4LpFevGlRqpcko8T1Ehlzz9ARzce59yRPdnTcrtduCmeJpP
sCDr1DMseex4ZaSSStblvu3eBYDsJKi68yOowVSgI/4PIZU68JuGJSjrHpgRT1yqDUMnlZuJ96uB
z40K3mLrLvK7F4h3IMR8oXUArWKvUv8rC5qlhJlcEgBXcHcs2W/D+XKgHnkxCadJRR7OkwPJD82x
8dhGnzMbxaAwxqW/dONOVVHapQnYCzYbkJRQot3SsRNRa+jcXSDfkA0+aLA/eblkTwmPpMXjimBT
AB9304iwWjMekJSW2Y7pkYqkloL0Zw5Cf4x0tX1cuYGIRzqrbMfOrNA96GDJoHF1ceOp0jGuaDgX
ku67emqD3fy1E9QADnYGW9Pdj4xQU8xby6QSOQsu2IdzHosF3xPzD34tdJFrS8nr8i0dLdLZyJLY
+NPyGslSF1QzaU6X6iVw2wsJuwHUxfPNwKahVv9HvOLJKJsoYXKQE45AcWIldo35EX6DWOhGL8oy
z/fE2fr0GeShGo9njzhYQzPy+EARFHlUg3MJYlL+xQ9s14r6fQ6FTDItLvJKQqe3nMMDRzaSMTv8
gcAJhztQ/S2Z/vLvj9OSBh6t3tDIVRvb0Wl1C55811HGn0H/9Si15GPGbmG4toj/RKhsudHfxFus
sOYknNwjEujhifcdlv1WgH6MI+Ie9cQ8v9lxkXraArN699b1CGfAemBcwD2x6P25LZjund+TBQnA
ZgsFE0CppqkNvR5u03L2aAobHgKJi/REwK5vUeeo6zcsVbv/ZuTSMJpXJsuWSgJYfnbdZAJjcTaO
UtKKGrdiuX1VXdCJxCjvcHCtEEpSQqTvFwVd3gC9Ydwu0lXiZ921Ui4r49K155nRcntASSPCubTB
3rMd8aUHMF0FTPEzBN5ZQ6YEnJ9q40pnuT4EtDBd+LkQrqWsLZFNjPV5CMfuriimUlXOl47fKuI0
HtW1EdAiDQjaSnKSgQK/j3KzeD0fxLLdY+IUR/9Qb5MJ8rW/sezkaW2mo7hoN84pR/4elD7L1tgx
ydKQ5Xj2H+n3cmGV2WGozbgEksHP3dmXVm7H6/aecKZP8QQrXpcc4wJnERpXm4kPPwcp3+/29BbN
VDNoNhJZOBsydS8OI99Xb/zbDG6KLVCi0LJoignHSfwsna1t06NK6ckDpAq+hVxhjbRmGM6pif6K
UkS42SJrTB8iZT/PDoMk8c4BagYg08/9hp3W+pKNx+cS/UevjuElhVW1lgqq5qeHFpYwIZEP+rk9
OqwAdWLENOhPDlIOQbctTxWyEUm4lSWkdvgWJURIVNLUDDDHyyFDI+s6Yehhf2/5VK4WyQ0ZCVgb
kmLrQ2GuLLn5Cak9W+0+c133XiUZlY9M3A4N7P/PaNPmPjKuWmeanooAipYu1UxznCx1BJ9aA7at
ynuFRCE8ZnueOQxxGVn25YRijY3MBiWBW29K6tstQbcODbvgUy1rn3MdZBd5RZzZgnnj8z+4lZRb
xFLpsw9c3Dfufi3Ed+Y80am38PtyQXSXimWBVzZRfsNj3+8Z0gwzPvS8ETST+74MvhKbvxI2U+q7
AZpTZOHl1XHiYvgp6VlIoWOPMg9wTO/9GrA+9Hre+SSpWEQ1XZeq2i0sn7cZVqvt4LPWoyBAUo6d
BedHPRwqRsl31NCAFCv8wI+Kq4CnZ3hcG2glYCHMV+ZJdhzoI7rvrEBfcnEm4sRwSJ+1SD5Z1XYa
y0kdfxn9eq0RA9R9tZ76D9vCe6O8TjV+axTremoA/xa8wpWCnxiR4xK4FkcWt4e8Oxs3IKgrvuQ4
BBcdMyVcO1LKzdK+TdAVrJihRiidULxkLISU62BmdQNaf306yaGOuxb05YUDqVMDRCB1Ypv71Lql
Aag0AAgbcbyQWx6b36lfUBd9s00l/yeVNBhF/e7bv43ZqoSdPNF7dX6VjMREUTSfI6LzdGehEWm6
XeE+cLcNQxZEqxVBYYcHacCt6Du0+lIy4lyQ6sHAbwdRHNBQrFcWg1Jm3sw6lwdBUeEK9DDlEBUg
a93BrC8+HtuGJfYdT7zVuzlFDBvglakyf/90hdpj83QIbvHQfcn+PCGCZHH0xGBsx3iPb0TdZ70I
NIvNB9o86ZNFBZS1xBE+sAM1JFHldFvWPOVVO0h7+5B6jDglZX8Il7pVNtcct/3XmY28lj7rDkGP
m/5n2VYsxwyF34c9b1hqQMdSMqc0cJTqRLJH4uV25IirqtQ4+2V3tQl5qdwwctkMpBkyiNCUJAer
2WMe6aOSroQsy8F0ATxRru9J32TwDDIiNFFE0wJnj0HItt+CUv2Li+4OOLQoOAbrw2vXIDYW+TGT
5eUo15d2T01mhy61xUFkCGk04uNiMdPqOKPNaF7Ws46CsY6tsngNdtpJ+G4c81NxlvxLnE1+F8/M
9jS+QQN5+ZhwK9titgiC9y0sKch4PrvInDfOJzs82Nzwu2MieRPOM3gc+tKOd+kUj8J80JI73b1t
TDDwkUvhYfAgUFS675TD1ujeScxhta0yOBtuzp3b3EDj8bqKTnd4U+UFo3+J9eitE1zOxvXi4LTJ
xU5sUEpJE4p9N1bhkbJ5hUuVK0sacpHA2OvyaI1B+8uOMBqK50cn7kCy7LhqHbILbToi2j4JEXA1
SXEX+5gw3GK++2FpsVKTT771OhJPjRFRO16+EAWcyXBXyS6JOEOae57zy2yYiPd43K0SiJB3TKaj
URf1IXN5o/0b5hD8dSKFmTGotq83j6LUN9VtrTuqjQk8j946YNuIScgx1XbfCgOPv2g/0oyCZ9Bm
4VMzj0GiBhXCs++DXuGExB8nL8v/ysrivrKNlAs40UO+s/YiOvkcSNYdaux33neO/L6PpkAEUne3
wWDhx73NJ3unVt2/CyHz1oVJAizaaaCjMnF4PaN/DsUWh8Dw1A6Aa0ZyYesOybgBNAxkaNe7UQQo
lOLToGGaMWrYHAFVSgI1mwiHKpOWeOWxSqNqe5CISEWprtaSQFnmm892zl0fvrd6q6ZgM8lwQdAc
ffzpbvwy2Y5GTuCy9wVAy2X7hl66Z9usnEJqfklESZ2yUdOBI15aW5U2Yua13stZnVrDuPoranet
Gn40bTtPDgOsDlvCWuiyxcAP1kqfKlURFwOvWnSsJE8g8Gktmkh6n570yXK8T5VnxY17ggdMEsKV
LOStPWVLZ6iz2nzjjdv9rD/3LxmyZQSUJjl+yAWl3Re9xYk6ELzupTHn+YJwcY3K9yGqQajE3Mim
oM4IjmTePr9+7p/C3sXc6INYFGwDZt6rPvyC7YF5YssugZhcNpkCc+0CB0KFHXK5mczsmybQLbH4
UmxmzumdtM9HhJ1s3N9vio4R7jLugyiWlbI0ttfJoKglOiYPzaQ1b7MO33mH0Ss7WvUC+5ib+tDE
sbA/DXIGg0czvvBT0U+HCkwvj7b0YoK/oGgUp1nCRPLB5cdu3wr6m73FhSxoKa2d/Ke1LW94SvyJ
l/xkIiqr+6qZq6SS4EzlQtAftp3IFmAdJDeyFjDwt3HZaamGbK+XaMz+oIoXfv4KIwB6WphSujwF
fuBFTnYp4BlHcYIstYdTxtGFLBFVTYkZSJPj6q3RL/SZC0cgxqh1mYPh0HdfcwrdLCjLeIXFeVeP
TCgY81r4rzK7+iLcGYf1VFHQsMrMuqrgQR5inSLmWUjzvBOmR5HZGnlv8oTswMSWGZNbtAI3tmEJ
doyrFkfK+LJju36GfVLTPfYtJ4ywkjnHxhUyPm79AHAQQ6btn48eQgCXV7GAuGchhinXjWA6EH/B
VLsFDImxPbOFPN8+bGZdB/RSvz72iR+nUECDv0uu8+me6xyXa6ND09/bwEyIapiupR01/KE9lxqp
btogew9d1nezvNcWBLmxplAdwjW6G7J/D14UQb/ivCT9ihKEi3EJzC/WYw4KFuWOVBMpKXZgh5wA
EcTyMa/1ohuPpvDW/GhJY36RgpFa54cbU0eADSYx01j4uZMjw7nRqYZ2BtYxwISnhh8Hs1IvQzMf
V25r1mVlxRvoSbEXbU52jSQaAgjLSjgw0nAuIwZ/39o+eueYC0s00aU0eyQPltO9POZNmdfbC8dG
reU/KCvHRCt9PbSlpLtDVjT+UzDV6V+zRb30zY50XFrZvHrhek5uMcrkTACwc6XTE66SvU63HU1D
FMvPYfQgnuIupObqZDxAc6mXf54bXW3H0Pcp7QfVHrwQZCtIdoASY8097p/wO78EbomHj318vHD7
Zv+aMHYt0RInsvDyewCvHK6hrXhr3M77FdQpCDto0zIuutFrNb9XYge9dTj9YbG0UA86FOidbD9w
HJY927M0aMht6hZXT8AQrM9DQB3Ei025Uhd9n8KuQjzC8l4S6S8KtAesy4vgPb7mzjRv3gAaDyIG
dOVUfDCy2uYXGrgWQUO0whi3OUmNuLDOc36ZfZaZZGdSA/tw4/TUZvLoQKL1xChBEXidGFQNUT9i
0UCTXB4QT3mmOPt9DSpDRzzWPSurvO+DERGrjygpSTangrtIlfi5YW2Q7JRVBvkVeFfXBxXHA45e
4ZdMvMAGN8I9xear8s9aa7t0nzyQ4D81zsMBnFGVl3Hoq+nUcXyloY56RUrSInrOQxuG8CQXDT5T
wTkFDmC0G6iG5QJKYbz9PrXjM3m+QDJv6JASFiEHFQsrBJEMBkCu+zMErJYMcPBmi6cM/pMHFL2c
DtqbKFfIYSKx9QOSGiq6r6SuB2Z+RDw+mZNWAWTK/ui3cyBXIQeBAEDekZJ7xSQHTDv8GiWiXSMh
UP4zeQAW5FHmM72dxyftnzxlXFWoymYOcm/Va719kiOP7SCIv3L0IEweukoGwgR9xSR9XyCPx8ax
mB4qt8TCWCgv9ZPOM9RdR9GtmXi3GFngruCPSDIptYzyyIycVB2v+9RnMYnPWW7Q3X/RqnV/aM1E
zxLpmXikW5qi10vjV9FZlL4a/YCHA+/cJAiBhaQIdqNouTSrbL+MHtf9mastfg1injOsqjdw5HIl
di+XfPqfvAWjGZKCpyFdPsy/9xbAI6xyUBi/Um1G6KEfOxOaqOhNr2vsozd9z9KMeLVqB93N12IJ
1joxy7U/tMOzW5Pw/MCNzZsvnkwnFfT25DWhr2SLhhc9kkILJ6z4XsELmO0nzjNbpK4dfDEEzlJo
O0ClBgbP63ltY1IxwG+GgBcGBlKgKk5AhriIV7sdw2Mxk+MDXgxBKv5fvUV6UKiwuQ9F3gbDvQ/+
IAcozhm3fU0uAikOXQRdJ1Mc/D/GeJ9pWtR5pO6tw0B4YxyqD+PIgSjDQ+GyCO1IwdZjPcj89U8i
rCixSARBzCr/MvnSIFa90qJh5yFX9RSi92GNp7L1Qa5N3XfeiTgCOTT3zaq+Cr93HGXh6SXtcTNn
RGlYrz9DFXNQ05aCWyw2kKIJ4Jbf4UW8oWT2pAAMyp53klGv14veuVuFucyHs3Dhynof+IopqKnw
meSlkrN5/AQppTvy74UKK3/rpzWKHhpl4d1hc3TC3E7CYpn4gERiYo7BmSKBIljzXQaSYWWAeyQ9
Qmyuue2/CEkQWrNIArHCATngqKgyV1fwqjOqULVkz9xdfRlNoe9Fh5ZSuiXWlJAvMv+9qxj+DQpj
G5AYDZjfMeNmAt+CUhMNjODiNP0o0vUo5UhU/z6NO3cUhFBzPM8hm6174HWvxgMSBVPgnU7fk7al
WA00cKgYgM89LzzQ82OIYIun/xg5sMeRpJE7qz/pphFxR0RV6smyEEq19drUfIMLJaXEDWRfFYdK
uXrT0wAVQlWClX0oO3FpFCVkg6JObMS6irhZfzXy0qf2jrMPzAYzCsyQiFcRZNzAfryHaMnrMNQ5
HvPtt3LwHX9VL+AJIKd5aVjEfwMthUkYM9vVR2KAveXmk+yyRi2CqkJy85/FX5XvoFEpWZdT/bVL
qqFiWFM6lVSK+RbRux3+E1qR1PKFiPkG4SVEEW8MfbQ07TbGsDkdROlEGxEU3nChxdzEwpAi8pIi
zoh2skFSSeHJlSZGGhHFIa9FilsKhnO0QAglseZlQPiZWiMJTGx/wBlIo4Z3U1zJM2W1cygbxwkd
7uiBZMFahCDGr5fPIvjPZDvdVFkw9cK2z2otyat3nl1TLGMLwyI1I7FEH4bOVizaSE7Ibvq896nt
0K4xueLDp6ULApXTvKHdAYnJarSmBirhyRyYohlVpccxd+leXew48xmKCoKyeJwTUqynQoR/IG0z
EkUtoUeqyjdQNgGyRKrFoPWOZZDwIE+/QlVF6k+9DBOSamnVc5zfIMnsR4cFotzcZX3CRbaIZdRi
Msc/o7xHXC7eJUmXhzsuxWKrcg4H+dLHytIybzyerkYf8nIbf2JYk+h2ELrqC2zUVco0ToZZSeYF
Q0GxMcJAxR5tNLGUHVle3yPZ1h3F4wnoqhbZrCVUCcQ0QkQsib6XbtpuClfabRkZBoBKo/tNLugt
LLNkPxrVNxMJ7KbMWyakL7GcgBEgA6Q+eho+MV+ERDHS9SZIS/o/4eTaCNY98Qawx+8RRdvBuW+t
d57L6w6S7tfANY6RuvqTJzZ0gKLiOp+Nhad8rfP/Y8tArMh9c7wjnlsTrTF+PzYMqUIlW8gP474a
ZmA6Sd+lrNFtCpJZM3fdNc/vUkAFdqD1v/ARhClLcpMa3i9ZL4ZCnngIAepM6bw0JIzP3Kvvm4ox
m2ZMUG2GAmym7DRO8F1kdrk3WobioX0PWs6eHLzgoVR8wt4U/lCzY8lkWX8tXZluyBLcKCFWbDnv
EGRpAZWxOdzzrEjh2tsqSMDIHY4QF6sFfBLVVAVzlxygs+WTW5CD9bp4kso8s+bxTnfq5ZZrQ5ej
N1rihADipau1hBkdg59bRr6IfIXPWpKnaFd+qoPhDJeZhCoAfKFP4DjZl/r3NPx6kqONSjw7QCFw
xMHLS3IazaT0+Ryb4GYu+uGL2kL9axPLOInlhhnym6H4kjfBU31FFjpTdHksh39wzfoBO4njwAf3
VccmzhsbHFUOWtMJXNbhVveBeJWraPT8Jr2ttK9mWeJIDhHVmADemZUCtyHj2IDkgfRwFeTY09tF
c/3Bt8+zIp+BWFsqEzQoarXC5exsKWBJ8YE54gDhfEf+grM+o4A9XOxAS6gxz4x5qfacs5QrTN34
VBc5BTHegdavZjNcgVFINGYtrxiELbYXeg3KOM4rBnUxtASvLpKpOgIz1Z+N9+vGoGmdOWvL7TCw
cwCH++GtXH5F+EkgCTkCCcK/eFP1Qrcs3eM5hdiSmD6464qR0gHKCp5Kkui62XzKS08/KXTAmmtW
54/WS/IypdA60D2QVK5choDaHXB2l3C9K+3Mpv7r8vAiEsuh0DaOfG5BrAswZieNP9asP7PQqmoA
pAj7HYRWnvvA10StoE6ZLuaXUNtsH/B+oPuz+8zefIhxzj/U723TRFNsH4E1PFbV0BcNnI4BhilS
5LgScYSiqrsPc/0dD5RfaDtUaGHZwtYUpdpLlB+TFrxTC6HYscU80cWXOKa4xKMVQVllVZ95I+li
hZbtMZfMXQ2LW62bl/RDysxBgLj9pa0cHG3r6S2pZjADXnm6nofQuhn+/EU06UzAuDhABtpyztxf
SJS00fbAwJO3IOYAZoYGoH0DYe9Ux2KbpSm174jVXDb54ht++f1Bx9MoqA6i1kdj/qc1LWZjXWE4
cWjr/+zKJGz457KhpKYzLcxQco8Gq+G0vxgGQz/Y2nw08pCSwjXdqejfmWvQKUln2tjRQ5N/HYhM
qh8ag7bJDERLzpwT0MkRxuRo4DqmId+KCsMxevmJnGW+ZfO48HON3WYi8GqTWbeG4fTG4yiuEnf2
KijbGyM8MkPi2kpzWp+ZAzLt3FCEyd18ZliBexod10q1QtjRA8li4yhvMj/Sew6z1Jt1f+Gk+mqV
cquNdGmqMka5eFcDuI/TPTwOyKBefrBfUJskl+wk9dpjfJap4dr/1UI6vckLZgeKdFQpSMx4vNy0
S7GaseoeJVBNBxprbGloU6fv5se7aDKkCX2fHYAnVPUH+qvNR7rkguIEU/ljWFB4ts6uJ52351Hh
ZNMz6ucDdxYISAlTr1eZxgPUfz2ApyJ+kQraJdV6eHm0SmSHE7C4R5DUkxWqJC/JC6+e4tj5+yPB
od+xeTmFCpxA407kOfsvqFBB/GISsMNo6yGqCGu8vPfyXxIVZFTsTicOQY6w45L1pAAyEUpgUXEJ
X0ccGJTk/rTCszaX/tMRdByci6PqUMO4xUG34wRMWVrvtkFWqYObdcG4H3D1X05DcmFr+a/WbuLa
0CoUwyC+xCYawwrdfQYA3W/l5k/f0yY50r2xtYN5JD+0GTKil+bRRa0giq5YVPZZxRtTs8jL7m7i
Sg5/eP2+AzfT4CjOzZ101aD4n2z8ieP8uVEcQvde4lE4QjOxJ6+NDJHA4eSILRPaYXH0UWAgCJTZ
fGE0I+sJ+mBUsy9enPJjAQrrgoKcihCbm7R5nb3cm1PHLhBthHEwhbudX2WOugp8LQC9DTIptsN2
H97k254C4AWTTrmmFkoLD41azeYTo7oAjhImvs5qCvffU/sxlEB9YMtdc4JyDb/MuIKCEIsJw9ry
tH1ljIcjkyAAowRXd4xx+SM7ZxK+EdTHSRaG5eHwZUWyQkeXklSV8UPTlEBaDqT30PJasJwS6EN7
AczOuHVmYZb3j4+qQ6kzxSyK38n+PW07hW0NMOR2bKGwoQbWIHohqtRVjHijva9yAX+tTLkcHgHJ
HtmL3b/0BrF40q9qT5KyiobuXv82pLyNR2a3HSTLOuKSqHojaV9+VlFk76LePGDFIZEHXsZQt8dK
x+DziB60v9+myMY4cABrT2Wdmc/GWVfuwm+p7kKGAecG1QIzmp7o34wLpMmvc7yLlP8dODHfGu/E
hKRsy6PYboeg923MIsWt5GaduYjyug7wOSh6iIXVQ5T0yQzIB0YdrjuTV99sLKAGO67IndOUy+cW
zfy0HAlwJXgyoBMu+2nCI6ccA3xY/x3ixWKGOfiV9EQKOChxUtdXVgtR861VU1t1SWlW+rf/Wy8k
5c57sYlqO2fOw1e/W2zycbl2aNee+vwPgRmFkVi8I9IJh41rykP8g5PIFDbqjLa78w+WwTPyKeeG
/Fx/Ub8cE1zI+OdXG+q0WEqm/HBLm/hRRZnjiOHLllYc72FfVg6Q9n8bJVJydxAvbjaAcc9YgKTf
AAGY7q8lixUEVsJyrP05h0jB/Us2TVioe6EbvBO0vRbY2a7VKbGShZsjYsxRXuMfHH3giARYoU2f
lu1cD9KLEhuLlbXRNENhygDeCZqS2ceV3mtmpNam+NIPyhVNbEFBl0GGFR6in+Df9A1HUaVOgD02
fHu0C18vvWjcNrCk6B0I3VWj2kwJIAqsRkUcTg/uAZersIjGM/jbKd9B8x8KL1GLhUk+ICok+VnP
BysWrAGyoIjIYwaC4bfTwT8QuH7350xCWmQAxhv/rSnomHeJI9K0hPn/DNW5joZbc8jLVulfxXdp
tFI5vf6xol8xcsIaJcKd4delKfYqrXX9YRgc7uxCZwuYtO2GyybyS0wZ0rRA21zpmmEQxchX+eUQ
lXW6wuwntppGvBZjj4HeioAYwxNbpk/ARrsVqFcBtu2D9k5GdEv4vJcRAYM8nfq78AslD0RdzUqt
g2ZNtbPAx2rCMlm5Gt547NfAp4OMrXVQBsV2alYvnuwCuSGJODQFddR69IMiZkIev8HRWg0tlCT0
z1ZB1h+0th6aprKY2ltLOg5kFDWB17m4d4ajppJDAZHyJsk5iYf7ei8yYeG6dIlhML2Xa9umOTeT
gb3Q/nbhlZpCrvr4quJYtVKxMLXPPw+WGF5Odo33EE/5wCeEyAHLr3zWllklYRjVS4MxpA2XmUCx
/yCEO1iM+rcsx5UpGkZUFTOsqzImHkzIv4JfhpHa7nAfZh91CkhGe+AdV3ziOQ9FODAcq41EARFi
vE31GHArYOZH6my1C0gm9WdDhbORuBHuwBddPz1nP7EyTbAGH4rUUXo1N0uUV+HohoBiT60e26TW
qmUri54gNbMsOkAxr+FlSjUC9vvIW4FB7rVt3BilRvV12HoRg8oTkRGjyXElXDOVFN2LLJIHWXSu
AeJni5L6RRwEZTA7A0PYd3cHlZWHQbNtGZyihmdvVYxrizwLwrv4Mz8CI4pBIrbww08UjSd6bsEo
lz3Jp43QiWLWsrNx9VR5/bff6vO5AiREDwQUDQJTfQCeZnXt40T8KKbZyFxnrcGsTBY1TOhaeMk5
DDFPhTvi0cInWGys94p9NiPept4CN4B6rGSxrxaX+nPJQKIcesoqAWm2U5nedmM2o6YDp8lgX3X8
/jf41xZW8bFv/QTepOMEPN7UmKFUdPKlw14laB2AM62Ls9uDn4Jkw8ku6MNFi6UX/yqWrEE1BDTL
uxr4Tt3+1wsSvXEvbtLrtzyUfaqofofmKdysNNSGJeKJnCtWsj9Pt8AvLOh+o1eW9/iVsnrRErwH
2v4NZ/y8znbwI0F8NepDLJgizV5xjFmzG/ccV9ABV/EtzUcifQqKdtfJtQCMlXtFVWu/Qa7eSae0
B81FkHU/owoDQBBZKhWTJhV2iDwq3UikPaPZpINMGVGF3gh8Fn6WNSXR5VcAfkGJUrnc+4Tn6t4Y
vOC6z9dW3p8trnMs95B2uRXwEqaa8E319FQY8zyk68hbEkk5B5sgBMuwg9SkcF59S6oVTDh8WzIF
HmlbhPwJJ68WF8Hte3b1BfBKVM+WTeh3SweD06hnN0TykA+BNuXZtV4rSRJn2ApCHVBampme6va6
4v5B36+1WfWvhMgw4TJzm28qT9uaZWcM9SZi1+MKJL6OUwTUZWxRkc8NsUvkVvi3Pk/AwD1iOXqd
fJ/PYHa1TxmYHuwygFpsP3oZslhy+BL8fxcg2K4GgLvWclTB+cMFf8SHuPVtKs0DBciI/BwloZlX
hooZRbnEGdhdS6SAYQ+wWAYDf1zBQscQI3xy4mdn+kpWu4TbUXRBcSrMo0Tgi7HF5JRT+1XPXViR
xMQOKFMH/tI9slqEqqTms1XbtnJS9L8M43RN6Vs1q8zyn/Etjxgu5MdLVhh/01CNKTkbPMP02aHO
2A4D+UvYMyg2MYRmOqkItX4FxYF7e9t0UxU5rqssNg2LfH4hIwPSjuS6k28TQf7dAI+VuaSOBTWp
32jNINNNqaoDe5Lv7LNRCZ/a1t6UxZw6W/rbU6tODOoIu9GRycY5vc4aAqs2VajQNM7wZokzethY
bIzfVpod8vKtYiGPRpPueWu+JGbcvAz+0U3cTvrr8DCamUyZamjtR/x5PooTqLmLx3sSxHpbvRzh
OZLl5JhXWqKoE2zw6XRslKTMe0lmhISkzAjydMGu/DvzEKvbU+uZJ/5FPg2nFyBsl2PFk2PhBwy+
a8219f+7r/fUgzxBP6GEe8PTOMNxjomrZs2eE68M8WXVpBQ8JUS8HKtio+ac+HrBli8diyDtBDVJ
fEKDSOD0Hz2yScteR1rHd/+J4jVrzPyzfE+ZEQyihORaxetj6HagXmwj03/iE+xPGUWZFCweHsfv
UkfzFjfTFwHvNK9FITyPhIvidQ5sxKI47pGz9dU0dPQZxK6Mu2p+iHTLQoaS+VfjII1y5yAgpOar
SKTfedIBp/+FZyair2pnbpsOtVydXO7KKYfgbLuI/BhZgeBR4HaOYzc0XfG4WxXgYjjLr6EGDJ+5
nruTy5J7ldOzTov/skSNFYZuaxGdEcMt9mtS6qX3gHl3msfGh+cTKVRHUhjro5ZNC5Q1KMvPVrUA
SDfSs+CdbSxBV2ZDrstMDgnzyr7B24JTtbbAZjGnKAHVW57qn+V/FJje7aG32Ik5ZxSJMC8i/9tM
vtQxd6SMVladMrkz6bEpiN/ab2RoBrGjAa9B5Q7Rk15XpUuPTjFU1gQy93dpk+bdqTtKmMsG2yWD
+kurfyJTtq+D08BNB2yu8KLD2qNw46vL0T12rJC/TAKcA8r03Pox182jsJ/JxDsV1/BzEvHc3qZA
uv7W1MckcB0aBOiGyCT7xeYq5lQYqMbDRTffzQNtyp2cK1t0CF897uEzsW9G89Fqgg5SHPl7XUlg
ZG6XSZQBUItTGJew0RtG2BcVpY9gS/wROcOF8ZkrH+vXTTPZNXSlmoplM7V1ctZGqI4tTf9jge88
b/0PB6lyI/rz5x0KzKgUysz3vH7xNpk95gnYt+jQnKsi1qJVBs0qX5RDV3sbHdqtIa+NC305jc2w
89hnvY5t7yUSRhlelI0F+uOcGCom32eek4TZBAwdhBzZ+PMcK1EZvl/0y3NBkhpoegzpoBbazVxv
zpcNUAa0gbzHgUQoSci2q5AqzbzZ8oS2lkIdMG2eA9B6ds9CykxVUBd0zbKl0goIRZRtuHmERuZ9
yvFuhyvxwn9chmr1c54s6e4QbDUbZMQF71vrpY0e+7X5ipkAWl3U4BFw+TGbUjeJvtidJ7Hib+/t
mkbKD76jIX1Oe41/RxhekFFMCccHANXqFQH8hvA9DdqqLpOLwFktfrf6RX+41WjAk3CoOOyZ4yaI
w0LCxiz4zg+CifTLR/A+sV7kbjroscgvOvXFLkjkF4yYrqZhvkoqCd+yJX1NO2XUBGxbAh+IWcSP
8zyYLrQ15BCzB028seJa+iMDb3CrxMa4NJ4pWXcaIqpkSA7KgxuqR8R3Q9Ws6Dz6uQCdbZzfM4Pk
x0uijVWGkDRP0nL1ET/MGzhTvYYpLGYgt+6gKnn0uqKvLPwDlzQjc1PEqkdCHDgVGAO+SFJ47fVa
GUL25KMtZ91tGjXLOQZqHTQptE/xvCayGpMeEXdc0K2X/w2daQMEbJr2ObtbtozKySZFelbOvkaC
WhGtZpzggREbh4etUqon7JbrdtNVZLdfsIW+PblF5nIDaXd9az1EtjNX+bpoEmrtVICycytkoy59
LbEUi5HZfss25vjBxbJ1e+4a4HC9q+fV4fBaSkQKlDcw0Z75wz+XFeDefo9SYQvHpMeZIG9XOSfo
GALfs+ePY5l9y1mbOMmka8N19VU1TBwLjH/kq7m5pXT1j25HKY4zUsCIUg6V2Ni32hl5niYnSclX
Vx+TDaQ1+QQux8p/QjuswkEiFc0r7sW+zg8cCJIVPWGNc7qulYpqPXNyoPIq6nCoaClYg1IOy+gJ
3XwULuzCrGrR6+pWz260Eeb2c88FUp1kX4JLRQ6H823c3H+/rMOGa8MA21HCdVyNChueCdEVZoh4
+zJtciEV29lrOinrt+UXXgkxWkb+asH5b6jJLkvNZJoSOp3/+hWv+9tMHMgSfbV7WrpFuyiouI0Z
17O48S20BQi8TyRUPQvdvATvCq1347QGfojE5dV9M61n1lsdi+HYo736/74yi5OVYxLMMu4DY+DY
MTPw8x2ncOSmmHyoAssrlDGcxZRpZkuLMExMxbkYQY2pC+B7fn9yKdjwcrHlnXcDOk71qhk48qAS
pL0FC6cq0TnJCRAKIxL7C/X/Sh45aqp0BLGTC12icCa3es7ruhRGVQWyO+hgZyZt33oBsUoNU5Cn
kC9aAUy0nUimYJS4G6BX0do6BQC6touiRWkOiGiMedkZ4YQPgKGE1pksdbyTAcWSCBcekFx3r/SU
xbWJvAyxn+hQcYJg4FTFid5Fp5I3OjSsSi9nBb1Y3JJRHvpwr3VMKFJ2cvkRlryxny3HoW36KOKL
yONu0r4rIETMYWdLU/HrtuPePrNg/4S3nthvuyPH8+JOU+5ylQ5/fzkY/HZOFSp6emX/krgUI+9b
nsm1PhvyLtSTA0QGsO+DVnA4mrqry9pgxmd9jVKG0Wmw7s34OeJz/v4wKR1iE9QK5yEf88LXN8Tm
V3h/A0ZfDZPwyq9yGJyJj47tndtRU6Lp4ONNLKehA+Y2XF0+aZJja1IFUDN0o88nIcNf73INVmx5
mfnbJE37Y87a2nIgXU67fMYdRUIkMZ8vWrTyIQr7UDMM/JnMjOiK13/pa4DxXNWyAgUX1Q/h3mTG
8Cp8OofNsoKNZPEGT4LAdNvz4XpRyTsTk3bII357D7Silzae9GlwacHKznTon6OXUpucnMwjBPYc
MncxvQgTMutvGcfpcAIBjBpYKVZwuydygWug9pNj9/HDr53vgnr1f9f38crNKEKKPa7ZYKKYUQjn
LFT147Saxae4jk9JrULiBIvkPs9jityw1RraTBeis7pvK4O6SoPkGoBb+grWx4DqN5QMuN2vm9Sc
eZVHIKubEp5m8PI32LywoaEQnOhj29TsKhEtMEBAqLRxnPPnvD1MjHBSSOzRPl5Oeqn1r1Be4bNh
VSpMkwU8iPUE29uTJWHZlRIkF2NHDquErQWM9oL8l2iHvXm1b90QDges1hAgA1yVmkEfsxcIVYAt
ce+R50dkqO/4Ap91Z2AS1tPCvEtv+HRom9f0fAoyqakGBn10OGZS8oNx/Q5B+qxmlbd15MyYFxo4
eLwi6MnG/pJ+6kZr55eoup6RHELZIkxMkOp+3gNrab29tGH8b2Og9C+Kwl1GYnyLvYDqjLj9TT43
CcKyVgT1STnYIfCXYsBK9ZCiP6U+mh95ZBmSYmIzlRsZDVS+JZ1r9CPjR7FA+mJwT/far7wo/ZLn
ivmKaMXgiLSZ3P6wZ9dNMeKBuKhbAKiVFZw5w2nrmR7SfLsxCtYCePTzHVL6HyR+IKbwAVPyyPV4
H4b4Amv+3ScX+5h+8N403ZF5ZhnbWmOpheYpuCRFjFnioYwLR1Y2AcTBA8YtPeqf5GSGq0jF05xn
9HhhrYNQseVDtavX1gCSIX6qacxxaebS6TIRwHw4pbPFlOt0GUnBSh2M5OL6ec2Zew+m1/hE6NNh
HWOlrqsbG5c6yUkQ6lkSBfYrLxAoLn0ziG/5DKqiyU0WTrm6XUhUGLQM0TdZDpj+0scxu+8pnIfN
K2AR2EkiAxl517xViV+w15jIc3EpoPoo60ERzNDs72X0sheaw5aGnAFIQgGHpZ981XhstLuaxS2N
G3W3vjH3LNDS07nCaTla3L6tRtp+ZEmfEHTAXF/34IMUUuz4PfxfhzZX97Y6p71Oaxy+lkAu3JiB
wvBM2WRauE12Z8kr75RZQ4095e849yBiYNGwGcfYJqD8tTwDUUv4E/uL3WT3fyJPbiXPUQN4dPvH
HzNrCIHq1ji9PWImDeVZRZkITRDRxglTjgaUrDMqA/5YPFAkP7O4TqCUh6COQ/oX1TxiMo02mk2R
gyHYNmfT1YekYxHbmQTvcyIJ8jvlYVmOGKx+IDFS+AqW7lN3HeL65tf3ezEKURKNUrWRLeUcqLtP
03qGISHyjrQLHvzIa72VmFAsI+o/kDZtq5Rdm10YsAj6vqkNq0akZ0j9IxXk2KPJu0b7+OrQcWNy
0quhGuZDywgG26pqg0KV3gTSdxjJQTnA5NMFDVFxz1vy8xix5dZ+i/hKwTT0GlnTPmlxQecQ30gp
yIsPVFHinnsK5Q5rZ6pWs/fmG3wNyC74zb1aD6cDKoZKiEjpFWaSuy35q4If2UKiYB7cQ630RFke
Ek53+xYkJldTQi0IgjfjESmcl3abTZyfsrHDGg9Z2wV8GLbkhq6pR0nP3BWiXhrEZIGMu5HTJDS3
WitPY4m5GTux/7/4wM3dEUP8Vp1S/bZ98rze0rjg5alNKW0ka21fXGuDxZTZ+BOClV9xMRMVGpDK
WHjcwiXeP+PTyMvwZaa9c7klwTt/u+xnNLrKrceR/HJbPKP52o8Owbu3UZ5TGOt+4mJovHoeVZ0e
IIJXgd1PvH9xPNq/yUgVVyRJSkyeh6n1fxsgg5bQXb70rqz7NE7YJj2jD2lB2d/HTV5lCJFpP4k9
ucWSqoXIKS37vRJiSBuifSGnX5ybQRYvgZ0QsTWLNiLF5U+ItaqTZ5khoqBzHJSJHb6I2z3i9Xrp
oARRhcYI43RF4ch6sbPPRSWYR6O+L5bGyKy77b9fyQPlk2iiNqyuGcNhPsfmhRF2cO7aztINBjlX
d7AkVRKAJGCkcGfIVr3swxJErg4D+EryXCprBy7mxgWg1+1gxyYJFSxZCNVG1RDFSSmhUPxnodEy
9qAgp+wQSM4+RShQHZW5BsryoOzhQgssjUZBCRvr5xNJhK3zhUFoQUYjNFAV+RpDSfcd6tWTTumO
gGaZao7WCOFsUEtFvwpkOI7ngdg6Cur58YPav3I8qyz2ud4+KrPLlKtkrPex+m2cpmklo1JEv8ge
2fXmso5lxq8pAz39EnwderHtbifhNYBqc7+KbBpylcoFONw57Fuhmxi6LlSwULgNLmiW7hO52IjZ
ip1FFSGik1XvynlEElP+m8hfsLpKNi0VY14qAYKiE/aTgjVa0tbjPS1/FLx6Rk8TWYwmBRmMnr6m
AGZkw4uuFTXpxKPhwiTFBlDQ9nPHYmTRCiIbGXTdgNk1WsKQt7qjglOD2mxpMg4J9NpcDG5x/lIe
araAslxfmc+/VXhmivnXEUIzO/IekrX40v6cPHL8/sKXlQuQROg/s03f09P2AnmLXyH1OHBDkPiZ
iF1G8WtgbYQEN7KrlCg5cPOauOrjY63YnbDmpn3BgnvoeT4foHEwPStpVll3Z8Xbv4Zmir07jS0g
pgPR6c0DVFwhuPyRmH8dLhi7kG5lDGMXrpGnSqaXMr2JrZMsgAd9vrZXO65K8X0aPOo0951n6brs
O96Pc0Rx2GgiVFXQVsxJiMqcC5p0LEW+7Z3LU2Hl+iLifQ+YX9zM+DbKIpeGvc5X5wWtjtnI0IqE
iFfvJT55Ni6qEDmqEB0atWrOtAgw1zkP403vxFMoNMSweTQT2GhlDJ3CGfGjuxKn2dQV5HPQc7j3
wFSPukFWmLV2l5rZHkx2mHCx/aKwZ75KuzdyYQ041alhHhm9T6ScoyJ1e4OWbzrmERRrB+PrB+YO
Y7BiwBg6qU9pfKRh1jgBFtomvn4HV5tvqiwdPIYTdlfYrm6tL5Hi0iOvzZj2lvt6yywh5RZC12JW
gh9BAFMpBC4y+goQsO7cTg+5J/P1NAMn2LMgUHA2nn5YOSpKC95mRtNiHMJCX3FNnR4MN7srUJsy
Jya/ouIbqXkUxgmSh/DFl87+a78V0boTUUQRf6VzMGbJxGqtOkAPSDwHKAgq28ApUkqsMuS/vK4T
uQHGzdw1FTDEVG7LpMQEjpqpqyPzCpYuU30U0aQuR+Hz4hbjTyDhldcM7KWK3XhqfOsaSJE7me1q
qwGrbGuB2xBtAs6j2rScCbkf+4SVqa1vjj2ICwP7gDKOh6TVdTex/ZJoQbuxhECfutn7v2+/Bm7K
QB9GfhEU+UzMAFBn1XUIheVWnvoikeKpYKxVyi/Y3cNHakbGZ3Vr70pRDas3p/2+1X0Nh6JXQ3/Y
Yi6WTVFjXiSQ6xFMK0eLSdVVlgPdAJE8kvv1RVftyDtADxCYVq79LAehNDG9QRBBmXmy/hzkHSuI
+G+4mC2YZLlSz3AqxMzvNxr+dljmASMhDwAIn1LqzG3EgxRfT+y4eNxQEv/lEnWX4NLe/EA6uH+2
/rFT0oFAQSTkhY8MxHc9ZmvvNWfz4B8KHBbNrEF3IPxYwLEIzDfFcvB7iuNY0riEhJ7AQFM9ZYa5
V86q/KSNrGqPq0pvyoY2aO1ayXB4BLgnvq5eGiIjJCjuGmdgIp7BGSNp4788magJY0EH7TvHf+jB
QSHaVjTwS081qWvqjNqNvmHsT2vFFtOJdo+bqBMS8UnvWX/B5H9SogP5oTGdoU0y2ISXnjXdV1lw
8aKvLOU2JCtdtnI7cuzMragH97h1a93xVUAoiE8aSC0NfJUDkPKQ3040TVpWwGTPPsTt2kuBDYaf
L+RZiOSOldBSjxECAz0G2zBoehcBaiuTvfJKYay+Rw2uyJWqbWTrUsocMUaZItbebzIWlMV9MR6J
mS0t8XoUza/oNyBPXYOWYutrTQApzj1DJys8f3dFuRzIOtXZLp4oDleXoeiMs2SRxvy7x5NBwjAU
56azJ5yn3jnBrImUwS/eodxE3YEP1E4hDMrzNQQGuEpRmNz9BmNatqlxku5U0xANrWJ9+4Olx0sf
jsWeIX7GyfS6rMVtJp+QtT1MPQhnX5jDzKzwbEjhl30cGlOQYQLREEC0RhmXAPwKZ9K01d2/dKfg
I3/o533Hd8KnMi9bkh3ZEOwAmcpzhCc9gg5TQ9sIG4OMgqMJdQT8tv+8T+H26SBTbQ7bE+HtOOtT
9Ire1BzBlYHbrcBTHNU6c8yrrfRHllR+hxq94bZcA9es69xmtW5sLw3HpeVS+ldv4lBIiYYrxPSp
Qow15KUkdClY0WDl45iCtGebeb3p5+TTLI07JlJscxGBGkiEOI0Cq9qXJ4JvBwFjRzEVEHcyP0MQ
Q//2ZzqJLuJ73ti/Ag+oQtPKp3v3DIJpJ0SL8dmNpR4d6zJywoLRY56l+nh6pfBDd6ptZbbmKuOT
D6Aey1V+zmlC5of6wI+7vLh4ZXQl87SnnhwH/N6rDtsk8sj1cgYY8om6L+Buf5aFJkQ6y8yCKydo
8wWSD6cBa8/22esdn7RdPTGMdmmq+KUQPUN2JTGBEMOqg/6cMvZzDYZ58ulWwQCD8QmoPSFmorXg
cKwqrQyEGNqknWP0xvVQI0PekMe8Zc3NIagMrijIWZBikjRSyhzRbRFUv1zMoULtofrtpBXUvRts
qpfMMgF+wVs3CVl5hqwHcqcediznfBx04TzWwrVlz2BzZwavgN2KKC3eE5p4MOuz7zQ1AfYvCkkD
9QyliqOHeOTYfaAjvsSMwAkqf5FraFcUWpLsAW5Qh1GP1kcPGQBErf1q+fQiu6HFVEZwi6+69Bwc
+1C9R87PdV0hWVXIsJj6kgET4HRqiea5OY7+e1hble9Vvc3nLNB64Axi80Y8Wm6fhefQEx6AUB55
vCU1fHghZuSizz1PdzbpVfoi/+U9Gg4KyeI0TdeDQSax8los+c4TClVhAVA6cPNOMIVhABTtSSmq
u5OjEQW9pH5a2NMIRRI320C7p/NtzEiK/5mV3mKdwLQqKDqvYEZR22LPFp1lbsIQXYF4fxG8ZDpJ
eKwjFcGLquDoVCP/m9cIHf+YMggtZspebQ835ARNOk5E9YEghwEzTjEEIGabFrSgHLGPL438dPF1
ZCTQ3F91kxAnEPqdgHLu2xzkd646twfIJGRqjVno/wlYKsWjn3hE5cqVVNVc1q8u8awTbfpYUXds
0OMMNtvgB5JHrIbEaLsEssyWt7D5Vf1oQ8eopV7bU60C/SUuP9HOqjsICRV4n6hFgsAro8e6UDPq
uUCj9q5+l1tVcNGeSQH8hPm6D7TRPry/ZtqP767FYhUWyGa6wJIJNBNJa2P31hq2LbTB78VbNJGE
6aTi7LkGTG/Mp8otVAzpZ6ct9ZdLfHFpluIg/mOC0wY7SwhMep0g+j20vGcB1ca2FXcQ/6Za/ezV
vEMc3R8OJ4IqPj2DK4iZBb8eq0iWWeQpa+w6F/4iTcWNccYnxC/KEqC6wPBP6GIpFndhI90LRqPR
OpHLGigOmKjLZVVcFUn4ZKOmltau+xbRGEoMe8ApZg78JuM2oXnTCPP5/j9ul/gDEMWyKbG0qWQ9
eiCSkNLzoLuS/jSL/r72cUBdz2jac3FZRe4sjy/Wd+zP2/74L1N8wpAFhInhDEkFzhgxQk//ZBdY
KH17dasg4Cu+qdNxIDqeNSYUQNViFCYGkqz+e8yxIUgnpZxTpGFysZck2RCuriL61ghQcpgU9mJI
MIKGllNFZFR9dI+vPyqND2cRnwzexN/0jtTVjHbSFDSotGObMUC4J25he0wLBaS/GWAqvEso99E2
6ix1ZVXitqFtg0MUpn7x5X07G2dRdGB2ir/M04pexHnB3sPK48e78YT+FCdma73gfL48P67f9RnC
5WIbYar+1XAbnsVA2ZnVVAxOdA1qX6UBh6ykG/Vyu+ePsoL00iwh68zLT0U6rMF0sFZTnclkwBjn
VRF8VT+SOQuAU2eLHkVY+8/5gvtyh64EGOVzMNLCpH04lpDPAd3Fy05nMbcYjmypVeA0Y/gd0qB7
U8Q2uRmgiCKvYu8VDtwzpHe9ENWR3ISDrKFrpnOF8Kakbhw5stWWJu751jhgNyk6IVeGgNd+BOau
f+n5SfzDxCzFnwAbTjXzK85hYQYd/dCWtCLeFvFpIxx2snxyLRGoLTqNhXVD/rsAeq8rjl0bwbTN
PDuz08rL8db453plpuPWQO0D1st2L+oHPB28X6MhIw5ys45BlUl2AI0iwgt43DaBIZvf6jNRAC58
ESdfwJ8erNYuObllV+WUCvVVqVvWVpa+UeQM564a1Tdi4D8Kxl+Y2T26ipE5SLn78VLZhfzG4+iI
kg0wzjWa7PHwFIZXcOgFmrLr3dBxZUOgBexnP7prilXGeBWjZARAvItSfgd4MACJPE/Xbrh54KuJ
wRIGxv+GNqziRBMbEgo+8cghzb6s2EJuUwKufhnmizFo5rrw3ZWjM/CqZiosJDjyUxWciRmCvXy2
RFTlJxPzuFFZD033LrQbpoKJxjyl7pzEDqfnQ+A2vjgZ2DdtpPuEf7gUmfsYtJ81hhM4nzQHgsGv
xxkS6gJcuNAr8S54NMcqJ+7Abd6UBVCHidQcWClIHvHZ6KtfAi8MyVICVEhqMfdLepnTFrLOl3Uj
KdE1h3cAZZ8/91m+6giezbZwYhV9XxuMVigoOAdaYSKbUB87nfu/zwb3lojz9lsczPJu3rW/X42o
ob1uAYABlyc/fVFYxU3lmyA0mDr5V7tBaXlbQt6w9rx1/nBMe1zvGZrPc7WUzqJ8llSMCfh8uSU8
wWm49qQBQKHKoLlUeettW1txrQkRVQBqzB5LfrxlCvejkg4zXZd/JS4zHU6man+bffgmIUx3Fmnc
fBq8rWH5mokIyPFaWwP8Haz585IKZotPfOq9lgits6T6yN+JuhCoMwi01HExlEOGwQKU36IC7ytg
9xzxcLtuCDkLLh9yk6jWPSdVKikLE/U1VDjOZU7KDf0oKnRX7osk+FXaMK9VGkm5701S77+DiuVU
Hy8rg3ziOFFBAOvzRR07Z9W2kNTACOLZQBiWxOvNJn6O3VeQsTpKjnNhUwWC29Vfvx+9dO0tIwIR
KZy+yHHpD8Zx3qa+0P7ACF6P/Npa7+1xKCW6pIrMXF56zCcWjz9iRFYryg+JUEExuzAJNIN+ae8k
RsQvJwj4IUYLRE5eqLHDSgN3wAaUayF2xiCzF+h0yMm9sDJdVsyBvkxwSS5hq1CVBaGQq37mFDAm
IZ9QINzmF5ZRo6Gr+7T4e8zMl8+3UubbAU4M6SVrAqMBqe10c+go1PjtBG7vxPNsO8/7gtL9m1hm
pKuGiWUrjLobos5DiGFmqLj37FjRjWPwZHXDNrHY/Chd2g+ZJB4YBf2IAiJYIOWqZa4nf39bTZ1o
YeHXmxAStCw8FCO06QoBjSpi+eYbzWORjl0I5wwh2UYQ8ObbdBpt69xkk72q/B1KgYbtUpaDnpFR
tDUCBv80vpkOVj6O5kpNDFZoDT2Un6Tbeyn0U2PJ3WJ7Q0JdgGVKjvzHIVbxaVM32CrSrU83HqAc
h2E4MQ+wAeCcYWWpkxwTqXzVSikjCCewYPtJ2VCj7sP9mjAXtWucu18kIWcDtHdnSLxqFEjH/t23
GsBzJL4IvR02siR3Jhj+Yy05/wPRFc898T9XqCbQCBwDlvAhV+pu4Ex3EN1NKK6biKte234I4+wC
k4COtO/4DBrFcdRTU49d6haXqWTduYQW4bViWpHDd2cvExmSb4gkVZh3Df8woNNUkWEQJgbJ8bmi
H8DLY6j9UmnPmBpELNf9bCgdhw1JuGN5v67IoNONa+MMP9vq9aleYLJ9mqBpRgS37Ys7dFZ1PVjb
lQSVbfJkm/C0JgWxV6iZ826xkF9lN/gbxBYixjgrRK/cSujsr5Ypuoo6SUYvjJ13KgqR17BIuUfr
EjPAUzCfgR/Tu/yKZBUltCeqUJzLvpssXlbpPBq19up4cP3oFlFcLtUXBn0MlwZPBGiQR1ld8kun
+nifzFFkiFZJ7YE95yvKFsOEPVoeDwN2HZkn6kqAJWTA5047MCZoqir5SOfGvEO95VbfVBvmtowF
nF3jcgMPDjdbXF5jbh1EyGzCHSGL82z1gPxZPY0y+HIpuv/R/tjjT6Rt10mfAFYZgKK1VW5ZIZqj
Ze5g/wLmUtZSoa5gpF2a/A67EePmAFbRk6Y4DkMMsDev7ZOPUZ6PTPGsm+FiUZeUOruZx+7vMpVV
JKs/UfHwTLEjIqjK07vzGq/JmwFayvur0grGJtc7nsFI1ikuKlEuaYbvO0dLsR9ptz8ZDUTAwDGR
oulg/lFLcwONgOuw1b1Gp21sGYIXL7CuaYgi7osjhrT0RXAHDaqmaTcjWKaIJ6k4xO4G4XWlaGIa
WvKzQvT3N5MFboWXkm7MqrcueM+vTYGwFLoktOOyPHKXoVjXScG5V2hnOhI3HMMPz3nKvmr15ooS
vVOnjUEdwH3QULgH67mjv4bBRGQxqHACyb/1sLwo3T0k2XxWpDvKVg9UyrkX91UrgIPUIe1YO9kb
17zWwimIsL2eTgCKiqCYM6X+mq4mQL+WTWA5e/wsM3FADH7wwkBZGvNaT5YC15o66Mcy1G99b99q
GZsg8cuIa7ju3r4+BRkRAVaVuuEnbaeYLTr9HiuNDNKqiVQPCPzizAfbhEf7rt8OHDfb65S5zBVp
Dxkkumml0QaHja+jXfa5UZKAgDEgo2jVhqb4u60fZvQIJoCoDEXSUTsYAIjy/q1DxEloZdn0A+bF
imk0sSaVWFIbYfFCYo+qBtOKKgSxsYeOrcXu3S5WJgr4OlC5EGQu9ogq6J0KFeGzljz1+VAOQjVM
ibXZ9P8srHOSRtLaeqsKTfJdyABmRxaU+Z8EzRya61jFiNaRcFk7i9+iS51ulNaR83RG+wcbE6w4
3LU1qIsdBpeKIT9GibhiALRu+VtnG5b/btrXcoZ47Pgsw89x0qD/D+wjuS7PjMbGhu58X0HFZqzM
hlchBnMSW2DvQJLk1ddcO2aKIqKGtE/Vru8s85tDUePOKPljGJWi4k1Cueks4yuT4n5Mg3+Sh8LL
2HI8ztlBQ+v/PMdUxG3eUXYx7YmdXrYJ6iSCJyhYxETzPahqTWd+WanFoPuqb1QyjlGnQ07lT52z
DbdhGNOeI7WWv1UzhkOrT1Z0poMFSyN0MBDlcMjvuwsFgFHGuyp4Cwop8CVlY6+Qe++di0J3ZYZO
kHiYelzlKK6uFnMtaogDM2uv4J8esn7ziGZ6N/No3rlja1Cg85CvqllwrZ9KhKchC38Bhx3BcnL8
UGMGiMPmMPj8xyebvDw/ZstlbKF0I/uDLjlbo8hysYoaqPS3mOS02lP6pVXIHR13GLripSWqZyOP
kQaX0xXblPaRUYQq3lkYQqG/0qkUWfpkfYIhIdSrYXPDu5wyRXmwzz5a1sxjSMvY1ZpmVG2/bNO0
yocry8XDYYLquBAIyaEOYx2Z8Oo/SC0fGvnbJuRFFnT7fuYYOY+K8Q3w1h6Z3xRuL4CV0SAI0dVK
HR0pYB6cbZeK7d+tT+pq6mVko/314ax+2x4J53qfibqwtn6XnSVfbGRi6H0H2eJbes2L0O3W1xBy
0T8Rl6bx5PJqL4jW1o4T5XB1Q6IUPCVdmwOqaoTDVxLlal6cIzG1XqrjCl/awVz0KnPnfDYCvAxs
caQn/XM9rtYsJaBwvpbt9bz0E8/EHCvosW5Cc2Bl01p/aQU4HS5oxv5XB3KlNede7GZDpbwsmkVH
2RO8o3vRiL5UTmGvo6c6JzavOnB5hY5mCQQL5S768KOnLX46c+4srd3FwKaUkaoOl+6Rfxw2ODFR
L0NM9sWTPzuNHJaGqzsGwhvqtztQmoq4NRUlRzs9wwADW2nNEHassNjjQiArJkCkKSc5wioXGevT
6o6OuyIMx+JyG1HFhx7Ku4VFQSn7yIXyQOQoozsWl0hINDbuz3QAbBlB4KTstWcObQQEFIeooxHb
HC3c0GwAv9DH02sp+H6e+y+JdD9GiAppcyrYvSOKPPsudIkNLpTpfU4C3jSZO2no1UXXf5hBS5QF
oCZbN+o696rjYJGEIPpHl56x/b7UGorujHXLM5xIQ6Ve0o2JDMSB08OcxE++6KkaeHjrji4y5LDj
dPSJa0L5nfSFq7Iv2KmVrdxP1Uv6LSLvb7dwv2ghbBr0BshxGitCjtzWoCKGGZxCmREhDbAMUTIN
TfIxlH7KViQx3PznLsfDqna/Qb+MHRMEXASJF+2yFeAdvquIaxt1HNcGZLxT7d1tUq1MRmPcIAko
vVtBSif2sO/AQrInblLGAHtluE1HNuEM6JxgFjdAhSylJLRhkNhXIrRwG9GNNx20g6qf0eX2crnk
QVqW9i7FuEgvfXuWnbttFF4Y/RXddNddq8iD37rrAL2GOd49Q0wwfVFr+L1zgRpBd4vCeXUMMtdP
s2wByKesc7OhJ2Fc6gxoU2EVmIVViQLHo7uG4SbV1362UqsmGahMvLzxPu0NmC57SbaVcpBbrXLy
w6hB6buU4lJrxZM47MG6Ap7kGetMBjtDvL9FK4J8KIh+7SoJWI/biWQgAXK+bZnRNP1D2Fq+C211
7G3hRdDwFBzvd1az0lesbIeBEqUiEUR78jGyest71/AN+eWyNMMt6u18SU7aNPp7FuSz1q2IcETL
QMZeYLvmEQvWThibXrXubbfKZWXUSiTEs1mRHP5akmLqlA+JlpvKLsVHRpAqYfEiTotZ7BwS9Yce
bCXwcPa9YeBv//e+8RuoI6ExPrSmy8tWWtuh3g/wdFBSXpozCaJTsZOEOXKBzN7kmrAZye53ziih
oE4ajGUA5pftAV7Efc4GuqGVhx7joLB7/BgqFEtM5QnO3ut6JX5N4hBb1+pLu4RZGQpsr65kyfiG
X/ZwbDvpq3jD0WkfzE27bikUIa4MMEvoCDxETEIPQR7l1K7JV9hqKbJ4IkkRDVGj/R7zLgrGQrnd
zc4npDY1jZpYjeRJXcX97wOuEsbzNIaCMs/ar8mdZc7WirYmxQIUyyA/1/xvLirIU6eqCVkyITfq
BOB8qnt+QSys8cj6iNWb1eO0Pg6ZPzNEEFcdZUQV0JvxBGgXbZohejqI4Xb4Nu5ydvpixiY6lsMb
CS7eUoa68sqvFXD19EYRbmpg6Iek1rIadR7/kx/+izRixJ3GKxSqxAZJdv69Sy+F7PHM3r1iGi1R
qM641FaFDxr2IwfEzW16X7xst4fC5WywP2XekZDKu6N5b0J4Pcj+cEdaB6O7tqG+YOaa7kaM0vis
uZ0UMFTbfbgDUxQuzHE3/56hsYPQhSyM9U63ENGYvUGbFsPPLusx0GNCXdIGcJcPVbYCz8bKgWhG
P640ERvXi1TmGjeV6Rr7JvRgW/Z4UAlAduWVKvMdIT7V1JtrneDNj0+Izf+jtOe+tfr3VLx+y0bI
lPwZ4axGJ2dJvcSjhwMSOPucnOjuUoO8pY1Wk6s0OowXaJcrjBHAF8CwKmstC4LxgQ9gCbCXVtLR
HDmsPbunHWAj42ZyaYTiE+qYbp5zTecLmi8WyUA8iiPxQij/kywuONvkhU9WaHAEZxSn5Zc+b8Ka
GUsAJxICwavecj83N1rQYfBYUqwjhYWASYBIUReCEfVz/gX1Dw6L+jIwuLODggKk5zMFbAU0lkdi
6thqRIgSA8msufgicET9PpMs12OXvh7FCG+d5pCEsX7JSkFAmyFxK1KZqQ2JKq13oL1zcF6mMjly
vVUHTv5b1cxlblHju5gwtYn2RyRO8OtcCLWH8v12EUBxD7FM8q96TxvL9rIUQl2u/PJABip1MsMV
ZQG0PWwTfFpWrPYupgJVgYuia/kKYk/BfFCklotUwGWXcXEnYm1dGQo1cz7qDWI4BfEYIqaDmB/x
Qm1gxjX/LM4N/B80Rvy2s9nUbt+78Uj5x7Ryr0Bby1aKZGMjwwAb5HRj/zGdTd4tYLPCkvYTA12f
7LSwDRlRjcFouMUlfiR2ZFqRgLL2Up8WEktHxP5MSTwRt6eFTQaLDZVbrZJDyr10ufUQC/031sPj
tj6mTXABzEpaYi78Ctwh7I7K2lfDHKadcv1YO9S/AskAihiXaMOJ7YKLSgdPuKpJ882hafvqI689
QFVAMy3CIURcP2SImiARf9wjeu01T2PkvFBA4OlSuTEMk9YPXk3IbEUxubYiGPhnL5At3N5kzjiw
d0UpyhJZaGKdoXl1wK4s7OYY2cczYQSpJgqNMEIm7OjKc35QYTVedi9tiTyoVrUZ5zplOOE+j24t
KDsHaP4uzOfM85n56qxTR7n+Xa5/PsvaYwy/LXbxq2SrtgCZ8d6U2jQD3Ju+pVeaEDYAkMh1xGr4
BJBQXm06lxp8KFOhPt2H96ceN5F8xxH0ObXmiIpQ676KFiolcwTnhlqQT1jjsPRI0SXxhGV1tXjv
7UxrqQycw0Twy8falyxUa9RitjHvqFnyoLQ2oIxFL+8UXPCgHJOP8bw3zD/zoDcafh5f/7cUApxD
iM3y16smcN3tGumjG7JA0TLQhTy7AfbaWByNwRjade/TR0OIOh3ZGYSrtvvO+ob9L+oscTdqaJd/
c9rNqYbKY8Dmi8CfbPIrLGDn8HVmwFX22E1czVXevHR/3KaQ0lUzPvJwhPVD+KBN1r/P5YhRWSJj
aFoAekMEfGJdGU8avdtmu8eLvZzFSITS5xZnIAjIMs1gyviDZGaDxlxVFOgn4KbEYFQF7KFg0b2Y
Hxags6a//+G/p1rhqA3tMRALyiJ9mvmkuMekEoUc3CwQadylzrcM/OQxBBqtYEmlndmrv+mQkUeI
lionPZD77/92Wj6m+LS+2bPh35GOjECUrcphxP+Ysqd0wO54Jk/bb+9+y3/MLU2Q0vcDZk9jRAMu
CtaOdQnvUiT1wQm61XGZNektmkCcg4U5N7aSt5j6hXCp+KmUa+TPmpEuC2gUK1XTbtXZXaieSqUY
/OGgwdk5pTbebsbvHBhJi/uHMKLfHOOTUuvX/OpFGk21YW1SO93x4gnlKxVHZe11vMSYybFxmgZs
CCjHrYelmiFklwEC9yyUtFUwVugK0TCJQiocyXPOgH+cMZCuonMvlnAQpSKm0TLHLwyzY2oEb/6C
A4WPaoqK18kkRoHTtMHJOY+pTcJkek8KOJmGLxHdBhFZq2WjreffkTEHRaAbMk9CSrTaIxkb2f56
KAA6LTeU/JNb82mFZVHQ0osVn41ieFJMjBA2l4XbWrIKIfYfA592TliVEHUB5kRKSnXEbeYMYnIC
js4Y8WG1zzUngvXr7Hbyi1JjB6fXn+lqZS09piR38xt1AD0OkhL9RhThGG/ZGRDOmzBZEawtIEbw
BR6LnbNjOo2QK4qzXpsnCnjTqlBiqJyW8OfQrD79sooFFhcXDOdkrIOf15maWtxTwh9QdLIJy2U/
z9yQ+Mxu6tw6gwjVPBZTjyT7yLQ6IEB1dqIyHDQjvv/q7lG8Q9XO3zpbJRmm0/FjG6gEv2ak63ZG
SbvpQ9E/cGADOtUZ2+fbHgCaGE4qS5PY/5uIJV+nhClkkEp4c/CRBqgx4vMq5sIW2oWKyiTLe49v
C+M+Jb4hflPVI10KW2d4Wa0bo4qS+B9SAowhk40GDzv88cyVJS3CK1aloeixUx9quw9TZWVm26So
1S/3iMjPsYIWZqKbBUslakI/Y+7SIuKbd8fp5ed2ooRLJtnRuDXoVRcU6sDXdV59Vdd9r+G2ligO
yG0RVGL7NJQoGuXqaL5VXkGPaXwAwAC1LB+XKkhqrR5PkoBjwDbR37DDBcqIOj9xkVwAlhetrXnt
kEB+9zSbNCFJ5bd178ypLHrAvPr9inbPX/n5Y+JyTogqF0irP+xDJdaCD1QF3h7AphPj+lawOeb8
iMqhPHU+pABtfnLADIfLOOyZR0xgqqvvjAtO3aYR3HknlsAxyOkYEpiOnVsK2J4SQYQGIxpwVOVG
3OkB6Q27AYRkrF/yYNezcqBQUW2Af7PtUuH7ZcRlfXMdDLrcaY+GFejiMJ2C1Lp7s6nH31gOxVhV
2OD93pQVcHQbXmWEXRN6w52YBAlony+1kHxpF5YXo74xkVyOmgaci8VBLt/0SwZ4ZNaTg99Vf33O
kAd1PK3MbaPfsSgBPzg9usdlyMyK1KJG2+5QYOBWho/ZxfkfljHFobPj+1aVK2HlvDjnxtqwgVcL
HaBwZKTqLe9hNUxqAHKX4izEBwiiUou9n4URAztORGUlvuL2ijiODCYOgAyfxHULOSXSdUNhiFHu
k6hzfDb7OnxbZVEgR7MjY9UDq0Z0RBb1oVt9r2a1rWS3ozUHHcAwcW/0T+oRK4qhj/qsaZQ/Sq5m
JFJyS/7xXspB8VaBjGUqYg/dno9gnieiVnqY3RfVP9gunPAB85Pw1Yxcfr5Z+2ZtdEwtbSJ1LGB9
CQmXQKCG3AO+FhEI8e2XvhcpPZ5vv8fxBvhnPthKUN5wWXZig9qwpH2QzYVmLz9fNfJoofg/i0xc
VG4uZ0m9GPiRRlu4/avOb8pLP5+OBF3agJC186eQdmWVYpis/rfH/ECfoqmjF5FX/NVxSC/kEU7q
ugpwgZTf9iwEMVljq1yLSQnL731cr9rN31pu6sVxiO/jWL22s41sH1BoyJLCuqbx4OlTD5TSayBo
LZMYU2pLaEl+XlfmCOwdoWoglMA1b52bpkyO09o6KlsVvE9CTiQOQI08/73rrxsGoHbY8BdKq7Dz
OwjH24xJD7bhxtHv13Wge3ieIFk01jxul11S10wWztBWfpZiz5Qcqckdlpa+Xq1EA39KakN8j0oS
lbVbpbv80QtFX7WkfKOYJX3csHqL0V6PussDTz7ZZjEkoINky5mEtLpOLot5HVWrcCpCC+oTBrt/
3edLDD50zi2FYQUM7u72e6tLwLB74niKEMN2mJZt18gCdKNEZwhVwzFVQILzHtTWxM5mO4YoP+/h
jaGCrkQVuODVeMFhgHNgdlAI1JW2iosLgSBh1UGIeT6b8Ol/+83bSTVbuycLaW6QO1ir2aiXlYfi
rshFKRvMzHPF+uaV4tPGRsm0v+yO1bIDJuGFK20sdrpQBtbgYxaNgjXEZ395rjCsYW7onciEDhpX
QvhuqcRTxekq5DaQvtAuDsCKfZoEju70ZRJwSIsEYgX3UEH0Rg1c3tMGy4ZYgQV2pAytxhh1V7Pj
MXwWCF4bJN6vfUV3GcYyX3UShn4kT1r/NKmr0bA8NjmeuzxdSv4jFpOaG9DyL7g7lqlceup6kHS4
SYyaAWp6KiWO67+to8dEhXK2tDaYtWqk26OybZWUN4JczCoYegaV0XGbxnAU8Z4l7sZnbEpo2c3h
zR9ppf73g5k81ruekprzTT/tpVCe6J566ISv8KhH5SpXpl5R+d1u6kVzqgzIrj+4758CkB389qLo
4n6qbV3YPlaTssvDbDEJ+7irLiSOIAwW6bYK4S3N0F1T0qk8VJuCKnfSQD51Pf5F4KJdheVMNNE/
YgvZxoJ6CqJg2ZYbrzwcNB+oSK7IApOMEAHMbvQblYENdZLWn2Kntv7ZTpaknj3Dx9SHv8abiRBM
I35xbI1Eqv23VrYbmlNweQr/SKP521UhILwhjnyzr6gRBfCKEMtJt7G9LinRot3YzK06V2m90dSg
z048oQWuYye6jlCGMYrNeJL5PXRTYJNyy+/v+wJ5o3XJwmxiQ8hbuEy+aSJREs45u7ee17YN/2ac
Wdw+blUBnLLoIn6SOpHKw+48MtJxR84gczJD+fY49EIy2pxJb6wy/npcpcOWTgji0154ZVy8IwFu
tF6B8NdlbBf9aj1VUYaj0JBlA0SasW8csw/vMZphdqfULh0OmZn8udOm6tpSk56y6BkMFNLdnkmJ
+yIXDu66Vqj+yE1Nvra1BQpueH25EPw5R35rgD3sepw7kXEUEgvQJDG8N6j0d13OUtStLWaKnoJT
s42qZOeFPUHHC4tC7NCPl2e3LrbXf4z/edQihbTIw5vOriCxlpzfogs6Jo0RB87ndIA44aMDjwTd
8D3Spk3d3HfY2vMPjW16QJqGQWPItC4g273MijwO/8abvUxE412YT9TP2SxqdQLvPX8FnEQlwENx
GZI9pKRfVPwbEKTjgS83xPfNAFT9H1DgF5Gwfq/D4Rj51eq5UnIEk8vv4g/uxhuHUVFIAxQ4hjvX
42wR+blo+CwUbGDT1Hy9lt4LgR+A+/b06TidHtY+8r7NCsUcGm31caqbGBlA4+pRa0I6NRIhXvW+
R8CGr3cMCzTGJY18CVRjf8l8uLkrUpzV1VWmalEb0iKpbY0CU8VhyDSfEJdhRQu9Wx1GbcDDSxz7
4Rme9fwyNPvAEy3Wqt0ZDho1xtnLK4iszm6Ve8LVqX4hWgM6jzuMbb7H6IexTzxQPLiU7PKZpZvd
6CyBxTdLTU5dFf53VhcIYYIMuIxh4fZnwKeIQ1SYt3+qaahOJ2iM6GvTFD31pUxRyzTnKHVKwpco
ADpPu+oD//PcZ/PMzfG9+I9v+H5dacbO/gXji3p1oxPM3g1IKS9A7944kFSzK4mRMye5l8EL53B7
IgRHosPsoSGjXnwhy0WdcWB3Sbs4vDbV4tN/+or84HyVLCLEnoirJyzkYjzUVQpea79YpgiaGrv7
Zi3Plwd+vRC+zlbBgHRnlE194o6P47vJUp7DET5SnYNKtTFPXfha+7ioyWzkLei+skGe2UV4Y1fg
Qj542Xc5seX7gUvqw8UXKxKP/1W3EqJ4x4R8/H5Go4vnLG6PXdCuFgRDhyiWsffRBLdfk+QH8qBc
uScFUeZc2o9UF6znPFA4ovqooV1Rgn1APQ6SWod+cE+cPUznUDMvUC2s4vPTD0/NRIf/7pMNjeN0
Q4vXW3uLal30VP2MYTqR2VUoULuYhreMkaP8I8aacTL93ZIMldPuTdjRqjW5bYDZrh2fWrRxeBRT
Z9himLLDUrMEi/VH5Flt+XiwvN3g1YxSFdJXYvfylOX3c1sS+Iua4wjZtR6JawiiyWBzb7h+nZy/
gkV4DE2sVV/U8ZvOdPpP/gJDvDzIAcMaQtd4+F96TQW+pMJ3GJwecjR4AvZSR4BFkGtLxAEJBS4a
TBVrnVutpHbDE+7Xh+vcTvmvfvaEwyPg/B3j6V7vvl+7MJvms3aQCM1hsp4YnupI7HYYSWnhDrnG
a0rxFabWbCXU924ugcVpudF63aqw/v8vALzh3E0VzRKEQ9v5f7eTCj8ZQZVzbVqHwNyk4iRTzZAp
C4wHjUa506SiZu6lc4ToDF/OWTObnS/iBDYCHEwIO42ABHumMYfK3ZOjIKwOnsOYYXpRuk7Ix4iL
fL1HhGm/gQ6EOvIDPCgf1A0K2eBZ7EwERyMwx13hgP9THJCZVE7gtmNzpujIiHcmoUlZZeJ3FaL1
3O+8ZWjZ1vs8S4T8bowH9dPByVkud3HfO6RZmk7SBDKNNsinnZ3wDnpxXaGFGCkoJ93tC1V2fwxU
Y0ZOvyXsx48pansDuhRHosi8/kiVBsC9nbRFAZ9Kx+aeche0nBGwkEriusvEfYTmfrWw5N+/tneS
Usq5sg8pLx4JGsRnGjzR3OZK/2hhFc0qRXwCE2spY/V87VSYKqSc7r9aUDUgmktkVnlkGDBbhPNO
pwbHvjAonNior/zDIuVIbMOjSZm0ITyuHBzgOKJnXPZU9CRSMcxEQxRBSAx/yS5BBmxG3W2au1Hl
LUG1t7r6Vmsjf+9PJ1OydChXpaTFLFzJqGh/PKBLSCGRX/psMEtY1CMzqzYHhf5cnWOABTn4bLdA
2HjmppA9Rhd7YsAgG6DuMEU6+JAxoj7TG9qLplP/vS/g59de8utHzPMYu8ldlW08ShqLH+hWxKI7
4IZ0e/kXA2bqblPWERKW7CNx2nDO0BXmozk7hr27oOgBITTxcpAplP/mWT7riJZ06Y0XTmHhKrgg
FbUJM6RcWo/6HoWHbNOl7CD+3Xet80J1JtRv2pTdTDKcGC0hs80ADuHOoPDRCR3plhwIdvaV00Zg
YPGvSfKBP1vJsSVHIPJ3yNSO30vxeCU7PiaC/4nkrwoqJP4ciwx6lf6BV+IVoMCkbZDa6kF2bEM8
uwr893KadsNY9HpB/s3uMX9dsR/d7PWwH8E6zpMkacrGkV+MER3Ks5JuT6gV+fN4jegXSfwG12TZ
Xaj42J2ZqG4HT6y3MuKXPm/uuVvl7sVQHM06llgLIM/jeAQjQV1cI2rMJnhrBCw+tHmhBN540Ch2
Ahjnz3EYV/2yB0gkl+fgWb3WjCG2mhfzO7UJNndh0cunrR79kYJExVXSnum4G1KTwZJgg1/xYkFi
qh671qFq3fc57rXLtiShl1PaeL5bZzd2wRSzvsXPr4H28f0Z/d/aEYlLvQglN4ROWd+Wd9sbQSXd
4iRHSShuJAL2fR7lcDav8NiDh9py3MqUbkqBAxZpbXVT7lUnSRA4ZvaiRNsNvVp+d8OMA7n49039
1Yrq0P0gufSpnpspLlkNolHVZEuoc1b63FZCcXrwoAvGwU1ryrhiOXV+pSJAue5tPu/wPBCsePyP
ulJSJ4ooZe0r74K+qV5+kpa2eKsDgD5BMTwhY1PBi7/ZqqhQMP0AoJSErFEtjbxjk7+j3VVQbBQI
oJa9m7idSz6HM8cQdBsmjFMkUpvM26wwEBMtpYu3hYPV4hoGhwEV7jJuP9XSZvBgHRptx2lNpw6y
p7sBym1Lszv3JIP1NY5ounIWyYwQWX6H56mo1x7YNpExLTWECBhddAvDaeb7U/FxkcVXTfts02W0
hRnNTHwWZuFwcW269niXdMDy3P13CisUvJ/y4/lX118xnY7ivssXofVZqz1qGpJyR/bCQQN5sLBw
6HB/Si41+exNBxehoxGXmEB6p0BAL5823v39U1t/KBlGM6c7Ka+SBYHU1rdYZ2MPjZo+PxBxYQjE
akz9LIDF3skFMc9XyrNUr00G7G3zEm6qSOeE3ARgHJSyvGLXBlXn/n+WA/2fyARokvWOnAK+/UCH
SG9OBO4VECMXlLTc5TsljXRTyltAOUyNiS8JtueCFSM0B/TmSFJP8BPQW+fUuW3dn1/VMg8sKDMW
7U0/2/r34N6uAUN2tZ0neiLepBo3jzJkufPq1yXnWDN1H7NhTI6SeuV8NRMNCLd5q48TW6XXXl24
YWoxU9s7yWeu2Q66d2Rh2g9qHuI5nX91xKsBi6OBSmfeUUv8vWdY9WY0/3lan1fXjJ3vXaJv/WVO
W/9G1JXtMoap71NHjO1irJf3xRXpvcrPjWSMboYbJod8JASQZ6pXYcb9Iz+4sGYqm/CpkNNj2ApI
+lJjiFAix75mAMHtCKjgP+pxwPZB5NV2epCBaeeyyWfzH4yrHYqLI9SApLAtovyu39ZgdxHDY0Dd
zE9d5iBtAABn13LY2//fRyIImhSUy1M44SQJ9KH8GtarOz9Bolz5LPN91dilJHuCaalmZu4nKrQ6
1+ipzTNptNbr+x1qcK2OnPRADFZT/0HrjIbDHutAM3CerpGgHHgQlcZAXHHvSF867NzldTgzxilw
tjrrgjLRtc6uXQhDHKR3s+fxEgT7M/0Bd1TQElk0DUR0QGd0DF4PnK777ID4SP2vU4x+fsaC9E0S
bAV+3l695K2dxzGpGYUBqPuhETaN+olmJ9eP450ns6As08D2oID2o6CPCbrs6hIZNyuE/pncKBkF
omIIOi5mTj5XSj5XNM5SMVFwAreKhmzVwD2f/MGaaV87ZazQcRYpY300JPQHoOybLKzTrH1iiUAD
4YAoobuL/urNQHkGpz/n61znKoI134yRbwbDXgKNEPVRfAkjRi3sYfv9TjyXaPopKpspFY3ao+G4
uGfCQOpir/0wGXNYN8JmcXXYuLvC3eETY+Xc+vzieVH9l6ruMEapjWeQ9qA3NU15YgtOUk/VzSGf
bD/ZI0nP23H9LWXEWgwcMZbwArb1+pPxSkaE0bkDyRadc+oEMe+poYV/QKSQJba+lEFMf1TN0jk2
9bp++VHEGDRbT82bOmnOQpa7VG7vsBASCUwchd/AsLPG9O3yM7FgcbH9ZcZ8ceEHJNmrTREuW0dZ
IUnZmh7M8sRz4RwIzaJ3JvNvLohwXb5gGdq1aXTmflq6Q/vvLUQCSBP9juyOzszJdeJ4SC4IqjyX
uf8fsNCmEOr2EkEJUfg+sVZOXmO+eWccGO7IWozAxnaxpJIrIN4dicEV4Nm4ZQhDgz0NvggrA+Gz
ZPV1zKtB0hn93S1b2htJyU6C3oy4falO5CqPQdb7Ay6crUA+cC1L04wMSWukaGlaBJJjPO75+vfI
13KxpN7Mlr2GSGhsBtO8fpSTvaSAy7wXv/UrTkZqVMInUixxUCc7Dfvgsz3Qf+mXCj+wt/Fse8GN
A+0UeyDBw8t2ixno4LRBSv8KZr4bTELICTz7YS1C9iKu5X+viU2sT++n8ETvZ31+Bd7MAGsnSMBN
RbTaJLXoE37UIey5KhQPVMgrIg4FBMsgUw4wpPPGfmXAa3nQ0j9L/xy3bcLP84Kr5HbbIN7yG5LT
aYIhpekUsOuJRquu2nRxrCLB31PCPYTFX35Cr3yGGqvFm27RD1BHfdpPS0gDV6g4YUlry1Z9nkg7
m3nkrgenNGRBYQrQZWW3H7qiu/Wx0WE7sPYGW65UsaC7dhBPCAERHAZ9F2v3fSDgDa7QU2SMO0NY
1VXfO7MVy3P0X/3rS8HKoYyABH0GoEXj03UMoE+9ReZb0hgFbnwNWSRULT0bsjgV3YvrfIUiegyj
5a8OwiVfhGhIzsw872/MGrnHOvRj1yc568jrEvpv77Hpagg0HduUkM3y07l05g79EzrASXvfFCmE
6VocycVtCUW6DkrG/idU9UstJTdFfLPbauO5Y8A6SMN6J0Ecw2PsWRFscZ7uTv7H0ZZ5PkXd6Vdc
dPpiisObKK+3eo6YIi6eZdY/0NjVuv1qHBNcYqKNHZTZZ9hgIk2Vzvd5dZi2LSM9LvUYubeo2NsH
onT1JjYnHufY1XBzWRka2UdfS+uk1M/zJ+U2VnFTZ4SPppKMlTDYubSmc+CDqjj3/ZqRbMWqhSjL
n152npprVKhoMnQLSzX81JF4/JTH7yq8l2pyOH3obc04GykQRCm+hixIHyIdnJiu9gqqKPxBaZXI
HhW47BVeTd74dtqZRnGLgoGTzHHKISiY6MKWX809Ka4Jm04IF30GjZ2hQqp7YyymC4ZtmMB1hXLH
+GlXdK4f5KybjxtS3IRDTjkUysST7s6k1Dr0Ew4LHZDLVJSoPPAStJIht5sOmJb0hdtggAj0Lnz+
kRZkOy7XJ+bf+SKUtrnKbF4X84lhNynCRqiXYPV00T1Zy5JmSs+33YHlK3jU+wlieNlQNq3t1Cbv
Mgjph4gxFQhg+W+XltvHa3ItAeSAkLl8yo+n0QisIg9+km1yZ8RWnOPR5rTKCNGdpS6YMZrU7shM
7kKZcQHneecCVO6m/7/Zgm4adWFVATd8HHOv7XbcloHk0Rz8yZ5xF825a+SUkUBklEwm0BbwwSxT
EBKDj3EhP1+z8QtHklYqhyYsyUQgeFM6/hwFkcVd1ZDGsEiCDLdSo79KxqRJbca8KuhaqtGq9Epm
kVlNC8bsLQieI2MScLSLX4z8U7cCWjvVIw/UBa8GGHh+eWr90tp5DKRhrNG1Hbg/p6bKj0U0HTY+
2YQft86DgfmAKNz482liMw9XKxD6h/TM76RTl7R73rJMen1XjDNDWS23MEhFA4BGZl6HYIcBJttk
jokphHrdWE4VbU9C8jB/8Q+3Z+4tWVW2mhpSPtfibnr/NRDTO2vGZWXZLphA6BlJMpYCuMoROZNZ
DZ16hD6inMUbrEPkLkYEdoGjCaqQKGH1oRvQT3zY3dXdO6aVRbf3D1s712xbR7cOhzZZ0nsITEIS
2gQzsxwpl/BU9neRrnVF6xyYq2J5/Z0umJT/UtFLRjhaHsjb5sqTI0G0pQnQDexBEikXVEZYMgFb
gmkrOIzSvaFefRT0xYxJLX3GHkd2IO3XbVQvRfOf8glvUdIbJTY+EBUNy7MrFKJaoZy0aj/QgLUr
NGo7LNA9fYYSDOzjmB/l7BP+8jina7aM3wuWbRnwjZgmcqYZV7LTsrJKEeJWdDgIptXyLnCm094n
PhnWb521CK22+jyIHlwmW0IcTKS5ZgQAZpADJk5JcntSCYt7O/HhfMxFype5ocC4fN934zD07pJd
MHI9P08FxC+qUsam0SNRhzRiYjTrlKXXr6l+4DPEPpNU+n0SMBpzP9NPNC9fJG1af3rFxl1INYll
5PA/Ui7Qz8hIiYj8sxbpwwFm62NaNf2wBEeNehmpRNSLlAefqAE+2jVpj+dQmQFPp0fKntEQR6DD
dZCDYxfE5vbJfrwf9886a9cYGkbw+Ypzr7xiMRhTKP0yK86znM5oQhJSDnwss1dN/+LsLsBYUXis
Vq3JNmt6o6iR2z/55JFL754z93AavYrX7ir/RszSApsHBRJuySujx7L2WoGO9dQNZ9Q452sui62a
3Q05QAONscuYnTzUn7eEwH4rs8/sXqhpbrvJnKJHncIy50XRBqYkQV4f7HZ4OkUVBkCvQT8wLVFs
81RrOTjD30qGjBhlsma2bAkp56TDdffo7MstW78Ijxgm0P0SQWA9XL+Z1Fd/9uUrWppdwEDVQ9UV
ZQdIAdKzMqsB90ZD3I7gR5sVfozGQ2R3bbuHDnxuhWOETF5WRX8XG9yZdv2yzUUaYOBfx1R3QLvo
kO/mXL+LBuur7553YwoSwE+kXnfYahoNNWrkGck+uEhpm77BNsClomXcoauM0XMG346g0FgIVHPE
L/NQFAw5tp7DOPuBOPxeOO0pb42biiFVgmnlLPylpK+Na5cZRYzobQPodvDXisFK1/8FVGksLqid
6HHAKSQq69dmXbcA6+uA8tnm5+BfC3bGgc+tep12DFV3+ndvUWI763ON7gxeBcwjnRkl8vgeNGUm
grcC38RlW0yc8Hl0nk3lVdiMTMgMHl2mRZLmGIu3iMaB6Jo90/yuWdAPiJ7zcrNCT34OgXm8laV5
NMSiI1ZlPEu+yGBgWNgVsv+km0+YsMfxmc5SD6cgnreBYYC9jxPBEhSEg7mV0iHGTglUgtVG1E51
fQWReqLhd9rYLcSrmhETEf3iV4YMwokW6J0+d9u94o+LRZEZopRot0hn5y8CSMVtfnfBtjqkG0gz
QfhrNzcggX33eTx/H8NZX9oAcNEQfLC2Z4dtRG9V40GjRqp+F75MlFt00KHleLt1uy/Gu2YBD6gK
XV/gHR/B4qh7EkB3GJMaKQLx2TjUU2jFdvkgp84oie4PNvd7esgSAaXA8tCerpGQqZe2h64DGqVL
9IQlUft5XJ6SMNrt9urJYLBvFXQeBfp1GyIvZKnnUqsZpwO5TcGB6YJc5IDK981nLq0kytdQy8mD
PgI/n2+ZRY0PbMEBAKolGh2pQwUMYfYR2yJgjPqA2pd5hXjyLacuExwhgIQB+rUODW8VJjuF8QMG
EBCRGS2y/jMizogTIqZG0XGDDh3AgmPWY5oRiYpkrmJanaGjnqltmrDVyFCI+iH81AMt6CfGVDv3
DKSNJxktAxNAHCIfEqlNo5OoBCO1Z0/x9zv/7ZFlyt3MPYM14k9B3O4j5RrtPHl+eGWeZhFOKMth
O2+couIDBuXIttdO83wR7fW1jgLExH7h98T59BnzuJHTW+yKEuCaJVgCtmJUTLEysje6BuXVGtka
A8yt5pD/VonRZzk62nkvMvoecf1L5JkiJ8NFCgDERKyh0aCKvdJQEguixldvEjxWjD1FsXqMTyh3
AOLkzQygOpbeUWj5IjroC7MXW4X7pd74wkj2N/W9YajBcX4vM0MEFgzUTK+RwaIx/pv0prDGcaf7
Su4Q8OOyU6tzu8AyZcR45u0T6FT/YqQ9ODJLmy/nO8PoXht+zedctZwFICV1m179w1jvsASGKn7L
wfUJC8T35O2Qqbxd6Wr0rQmTxUj05AmIUWMJZIqgtBeRzGO0EOOiCVmW7LLntyANRGfrpSPYZkWr
PTFbYMQdrMqHP3bFG0v14/F4ibIBgej386cyjIxWnnJfEsPICHUY9kl/OEL6fa/Szg0uG7OouRcC
kwOkWOr7/h3URQY2X4BLoPUeOqMcul3aFK2nzctvZa7GNGksnRnsCzRsx4zSQ6loA98GnfFdCX7t
7UiNSzQfAWqH4ld2NhjWGPKYaahIjR43rg/oWw66kXk/VfqAVdAh06WKl1l6parnsKOEXtF+XjZz
3wcNWJYLK1Wxf4+CWJQry5hQKugjhuGTKlaEjjbm8pL+2aY/+4DvIbgBV/1871r4VozwbjUs0obA
SCJllMu4YCqTHdkb7j0/1JqX97qK7CjfU8WfTmTc36asrV+S7RSv6DVsBhNFA+Qes/dXTnXBOdq9
EZDLDVONsWKNG8s/PvL4OxY4YirC91f7wErXd4engbZ9T1dRqDetNBJK++szLe2dTdSTqgno7ybJ
I1QLHnNB6g221Hfydq5uo+ZbKT/YwIcpohi0QMSy4uEjRgQ5uyoLL2eSpcVQMVEr7evBTlHBNMcj
teoZYM7ZP0lho4aoK8oKqcXzP61EgUHgE6YQu2tWrj7AahizW2nnNCYuLkOXjv8oL0m9D6Qp5Teb
vBsLbnu3ghr4gSwNDkze42w7jWN2XYZrOnenhhux6EnsmO9cEvM7I1rk17dRCotGUJ8AeFT8/Yoz
Ke9IJ5o0UrjjUeJik2LGAmoUdrd2SNKZkcBYE4W7L2t+DhKe2bgdJYuysJvaKvO3LG5jJ4Rxb4Uf
W7wt80Y5y7/KaDL408oTQDAjWeTRxv4C7ku3E5gPMgI89uIFRfyc/urcgHh43ZckBU6mBSe9Btiy
FNomnIQKFL60eAzusASD7U2Q6XQ+q3ZZdVaUipa/4pkNGGaYhHhDkS36aKvFC3REFJDOnKghAkKn
55upswE3ETVtVtcnjSPz6icRn9cml5RQ45hU9SsDVtuDfyeDs+9lq+kUsISGNAc5EsK/ecW+rw/W
3HsOTjLMXyIzrdA2ANPAnvnyjsK7w/KTxxmw/p5KljrVdy7oaJWDsjPWcef9uasuS/l1irnNr0px
9qAT6B2smgQnuHTD3kWo6TSpvNC3/XNzZ7LAPUa9suTX9+WeqDXVBIxREnS4mHpkm9zTzT/IP/he
E9No1QkUPLabcCkeyKTkreVun5n/Ek/y8hNC/DWI4DDXN9tYfr3RXeGMYAcE8XwgZkL43zVZtFLT
R0zSBNcsmyXl2mQnV5pDRBqu+Mv611Jhij9M/6eEVdMKUF58+maTIE28l0/3hUYLc+ZbXTiniVq6
w0m2K3wZi7xp2MglWQKQFQHOoN3PCAPHBE7FgEmkgmN6Tc9trG5vK9MAlYhjH/AbDV2KS1B7GO0W
Db0MryqMQE2NYJ8FmGOFAcv1hDVewiKeoBxJj8ArD2IyimQgGp4D3iYzTpry9yG0/jrKk3NkboVV
r+XPHQ61vzu44Yh9/q5tfR0KPO1EOuoJ8ncaGZsU64+HdCyx2Um6bi20Jm8rNBTAQ0RA6uDzOF7T
X6Ux+gzglUvtbFdXNSUbvl+96MM+8F69457iV/kHqjA4/RU0bAyVR/Lc7pybonEhbUXiHf1a2pGC
SYaiQtDC0tm78KbJAMd+2nWcKYpOaUs8+enFisTRSd3mQBcM3uwuVAg1NmUXQ8y7mAtW4CQlRJlW
cqSbSAp/aXcRJvbUl9HwNaNfeQRF3OVc898mbZB9498UqsBpYTsgVX9fUp9tEDX3g3rV6bkW/ri0
Fr67x53Fy4lc1tbzCZPcozl4v1/H3daFNdpNHACHsx7cdMdQQ+ro8P4bmrnH38FLy7aYGppsjS56
sAxP7OxDqWJP5gb2LV/TXhHNSlWYxIQ4Xr5POnFAIq2v73eR1KUcr83/00WHCSLrqwd7gjBLgnAw
xziVNrpX8btb+v2ll2i3wIu5wSYJPE2bDg1yOiW6oUI5NrV7qR0HYmlCp3xcr1wZmstKXnGBrXEf
GiucwdPHClh+spUN80DUrY/WVUJ730BtwXdX4E+59NjvluxkGWgHzIPxL4pyG20kQXPCEwmpCqbq
R8yffJEGSOtbO268c/leYLGqqUiOct39+0rlI5kkosFBlM/TG1wrXNTIgNk6LVIucVJwfJSfOqtT
L6cjJqRlv1XSsouMtC6h6igWWcXF2yy4US6P3RX3aXhykLfoNPx3xUr6YmMfB5fjNjdwNsjzEZEi
1UjIeJa1fpa9exg7x759uy3jEpqD+rFWGEDk/rzBl71D+ZK02qPrXVa4FlMQ2J/Byj1Ikp869Kb2
hjGVptCMUufgc/eF+g7c1lzCy+KByFh6uwqHarlwjJJmf+J3tYD2RFfT3elkqunWkbOUPLQMn8pB
IgbOgXx+pqtkbQ+5LT7Hm8uJXSG1t1sbhs7jIq1gZqYn/U7fWPKneJaPKY+fOL7a2ZT0J60wb2ev
1iWwIYR1fvr/5JbygvG1pP8lMm1wKPQbGbDJXEMidFeWxRyFlWIx/5EcPgBgaV+9Ya34rVzc2LQP
KHtt44kJJ59ktrvZnZta2UCLsiDcRQATv2zHBO35ynLKx9VuTTeeo1UjzfdEftA+GMNmzZpaawuj
VsW6/z8lUs8P5H1iYsxatMpTZ9FPeT/vH/ScEQ0jKTLu46oo9/xpOfrVkjojZpa0jZz97iKwvBo/
PS2RiDNzckdovY5GeZ+Ya7j44un3TOlmBS81Vztnis556ISN1TN7x+X8IceGboXmH0CU4ANT+keQ
yI2tSf6Jc8b9vjIGseeL0zQXe6zdlEs2zHFHUu843W2n++CSLJYTzGuPdBBxk/IpszymGcN1K+Ee
szURBy5Xp5XGOvahmRf3M3ShzkJLlxxfRE1CF/gmMlaYJcwLWou9aXppjydpjZkQLV0O2GEmDwBF
OKcHemSPDNCH2bMtK6TaDKFTC1j7wL3DqtuZAkxxztD8qBdxZxE4/Uv81ijzxgtI7GMOJLFMKXqz
+g0xpB6OgezsdRwaIdt25wXFYo3MYvHMv7luG/QPX2z4t8U0DJunP+RKciv7mVSPmrOynntwuISX
qV9NYalpNPoQuESuhcUIUKPgnoGPDgPEf9i/gCFNzmJ0aBe91Kcrv4k8r8PoRodg7p4ZiFiBZzH6
1M7B6uaQoDh9PeKBI1aIuWNBBosd9RQwkSF6Ey7mUwYawBZfszNqC47R9KserDcXLGv3Bwlw9z9x
V28+POoKRPCfnilq278Xk5yI5J1sB225SkDZ9d1HgqnMLtysQbFfT329ZkscbPSi45gJcdsZLQ6u
9ax5QJJ8TltI+t71JI+/Xn+ge9jG2l/Joz/kbyxgxveY50cRDuYE361yDgJrZcFT4qWhuly18e44
2bg5YJ1S98Ks/0tjMs5+fnua3+roXD16kfdCtKLF/NyuYAicaOgNjGvdh2in0fAnWu2JGYy4/usV
dNIeNbd9h1uoQ4zK3GCrz7t6hxqXLLlrwoPkgiAE3YZYkdOQrhADbO1xQaGNTxFxO/jkO9DgrvUh
ptgIZgpaQQqmP+fFEVDXtgvUtoBqTiRHqpd0+rO5KDep7hKznrat3M88SV0DDuAGHNiRp6zdtARs
hYv+tmQmgyJwO6u6lO6y4EB4c0s7HC3tC2LpiyAqAtndRN/c5ibQyHxriGsY2qzo5YJAsE9+ReBx
+pl2mbWwfYe7QHWzqMiCih/ch6w5cph6GL/gqbLIIoHUYH0qKJ+C9Q8bFI0OsNxO9mlnACFu/BOO
wum24igePa1UV3MP3O+u/RmtSlV1gkJ1ZKfphAQCoES/8n+1ParhtYbLzzMQg6X8Y5cmta8Jq2Bb
TLaTMxRXtRK4X1WPOS/qh3RUrsrLYAPjuHemg/WY/SLHd41O6xJWgx0MCwsENS4kR1WHxJy4+tN1
YTrh9x3AIU9jFWGTQxcaTGnAcXIR28/5YCfVOgNylgx/TpoK618+CRZxHJCwY9mitKoghcL4afo8
vIfG/duIkP2ui47mxSlQMppiExx92STJVJrFPB3Gg63Z/PLQLqizrkmcJM+0EB2at35H8jNp5+ap
rcSaDlnXixBbN1syO7u4BwvKqvaiRKBjQ+NnWH00WR6BwPFovZiIe8e+VRGBQbbcO7TOQoNGGyop
0swKI00ZharxyPSAgVT7HHRaJy0ZW7KgxRImbEbQaK0BcVUy7H02ZYgpmKePQmbNjX1FpgPh5mzY
zxoKlk5Wxc2HBf4aNNp4kULnlerSGE9AzJAq/0oXZY1a7pH2x8CjPhTxDxvpQYjj0/+UG5iB7xud
T3d9QjtFY5CRr9Pu30r4dBMaY4oQkEP1oN5AOU5FEXyTAg72+gu4NnRlXExBQZ1xtlXqj+OrEoix
KKtxL3VbenutkdbKZGI0jVMbQNWlnn4oOnZw5lFEF6ewIqFFTUHpCvKNGYRQadYfnPT3dMTadIec
NEQ8ZoaCdjYUghUZP7McfDQMw+UQBVvDuHaN9442tUOK0R7clhUSJF7Et0+qO5ex7hWvDwNpus+f
UwR9tdSHWLJ0qDu87hdp8LbBY5MIaMpq59s4MeqOPpCLCCeJtIvzMxeCuyTu23mmlRUBzLEiUUkZ
/4mxhfp+Ap+iV3PD/e5S2bvKtsp7G26NKA3IT9vpg9TK34gjBeA2+Ay/Wo8RlE9kibolKyyRRK4i
xTAL/gge9XgolDbeRLaF/WUH2u2p1hDqrsmownDMKryfuf4fYxBu347b/p3SrgSO8MY0/HTWlx3U
hHtXzrpVYZ6mpYwZMW5gvmYRNum/wqbu5zp34lJLT9IkTYzHjp7UvtgHQplHW7pyz9omY/zWBEkr
pCTtdgRZDfBc2b7iTU0tUj6S5cMW9poTLqnUtNcE/QMbiyozJXHXihhOHkKkCPCO073Y8DotFbBo
vnH52Q6vFXD0zpmYnXR6Dta/qNrA1c4TfxphWnLkq5jmJc2JvsacE10rlus6fPEzevoQr95JGJPF
yB2GW35/Dg7SH2enoXTENvQFkMbysss9PKTl7Nob5nQg4AFUpGBZx1xhY0/yTab3cSltU/EkZmxY
QjQf9DjBW5Qd/xFiuBaIM1UFX4QqpYVaaSZVk1mlfvnDN0/b6z1vM7B4h2vR3m7xzRMNtnsmdmK4
XlxqZRf2Ns8IHKGm6/Off/TZOiL+h078JeVB+52BWa2j08PRdCEnqaTbzkjHY+5mBBvAQWyAPdrd
1QpFqUDDao6SkkWQcYhp6EVjl5PAJV705MUg7KlpF1SW/CJnXaKRNykLKG9fmoVjt95VigGiE2JR
Snm59qJE/5UGZ/Q3TSWzWajhTCJQVuwWIPTRcitZFGSDcRSkIVFpMHQGexUdp3ES/fLtLGotKLLQ
fxJdHrKM9w71B8lQI0npV7JIMfgi3J2YmZrmZBIzAwfJmFRg0n7aAyZB4uUfTdM+jIdlMJUDLoYh
ul6aJZXn7JX7op47VffrYnjUkCzmM33D2R5/z//3IUzxzKbYFSEvd05CFoKhoP8XXzy1Cif4XkPB
evmesDU4G3OkxB8h7+iY2Y2RBBkuFWonrZSrSCT1jiueAxJRrvE7Mz7H2+OioVacH1hN4aHGo1Tu
UZwFoBuDXb0nT3Dekpy2bG+JzunrvkjBOu/w9UvPm/9ST2+BAvFIw/htWXrOlFKDSFRhF+8qQODj
yNXmbnC2pe1xVKgI8R0nYcb6YtkgGQEg2MTchlxTvFClEegrY+kDvHsvXzirigQPFLPnuPsRObzT
FVtQ7RIOELizm43XvtrviqzSN5tGGXYXDvxWmeb0ujWeiXkTKbp5KGhLkVRfzMuOj5g1HijzqrEM
q4wmwiBWey8oYZQor+QhC0wbCFTM3U/II4EVRYwJtgXwBGdgi9HciXJIapIX7UPlGrcjBctuDVB9
nrqUIGTlEqrpokh2A0V9Z5XK1tSBo7zgjmyA8/2dmkzIDX8zpBylqxdFetBfbmGvy5QakIzsphan
OnCb88SYqJLSty7ZfkNP/v6VpfpYoszcl5ukkwADq+43r7rlOGuTRmZSkBqzaUrOsRLHF+pfv38S
t0drWs32IkHQgHyEOqKnK4Upsn7n7nSU7DSUkYI0wQlU7vdL5O6bX8Usch89ek75M4G8ap6oejO8
skZJaCO7pgZlXTJ7iJo6bUdJmgCBirhcAE1HB+y0KWeizW3LlYkpyHWiL1I3sQakXhKOHikL3Qp5
C2odjrtw4N+2691hzNCWT9uF8PIRVWYVsnd5Wckm9a92ZZRAf6Pod6mM7lo/WIv4pIrFTVMHhErI
+I5I9A28+YTM8vRvqzgwWks5qPHdHZC1u8CmFu8GiUEcoTmB+LYOfHogwcFNY6N+8wXZqp2J1157
sfWnvJJSl41QWYLfnZmxx/LUIrK24Cxkd6gCK2eVkJiQyyV1nTBPN/ITcLERcNmZ0VgnFYHz/lao
bkGPD/kiI6BT7uGOPjApLA7dKK+6RL92WpJa78+cw5dCKhTcuMUT7LBFyCcSu9WK0fz7q1nzptHK
0zOgsdWEMaRoOQuXxjxYWZKVCuYfi4UkVdr14nEM8UTnoWTYnwPNkkCbZvhufdUCCcZe6nSJiGIm
OMkasRVtKJFnuPIioiEQ+KW/NFefPWjb/GqT530dxUotq2CdvK0c19iYVIQPdFN1m0LjBgjZGrfp
i+vZ+34oO0BiZM3mFagxrwwadpCNq7OcMvwieDnWhynUldtWgxSQyoRTFPZHmpM1ahH/nyRx3nNX
noc/nwNwMIh057jWk/GEIrAcZmRRBhuU/S3Jly2SKfUnvaNJ2TWVTt980RuL7VwwYblxhgkkAjNx
/FKbEVkIR/DFWes+C1lxfSz+xAN/SUtFRBu3OZXBPK18e+JODo9/Z74MEJLSI/hkrU8fXFdE6Vyl
fw716/zQTzUIF3WWwecywtKb5ve1RKr5zDJieOcSfzc+fr0sOimK7diPuAuoHsik51nQssVhGngX
jME8Ts2XsJb8Q3+newheuOB/WFQLURB1Yllcu6wxRuyIek0tvtR0bHBwqiuQQ7hk/9D/+UFJfzW6
OKS+OEmYgqjJ7mZFU2njh3fCAWpqerL+e5KBvtlfFIgFdJ6G43zfbN3d79LiEgVr9CButCCC1JiT
imHdNEjrxr+iTZB9bRrmgz5gaH7TZIMjjmwfxgIYEWoS9FFYXoBNzYI8GfxGT86DBL6GmNmrKlyS
36AUSMgozh8lMEMO8/jZHTHpuvNGXsLSmSHkd3V5Au85CfwHB6EGtel3WQsFPAgM3Tj6Ej5EN1UR
mZjt02Fcl7KNmH+8bkMJOFw00sFHjec6SXrhGbBsPx9pTx5t980DUKcCYsNGrpKVqu1KssGF59Eb
GjVK6BuiL/r2+9dYkev3MdDMG6NPHg2GHxdt2h3v2BWqu1hLBl21paV2xJZX7R4Ge7n65fUMOA0/
LUUNDAuaHfSO5JubLawShfhmuONTzNHNNfnA2NDn55KZu3pg+akYxfDAzTAEIn9z3X21NHmiXbwR
y7wxeuyyOujQl+NAUX93IgcQQ1e6id5pLZLGIZiPXOZgZp7fLYwC/uNYLi9BrqcXUPBId8b1UjvD
7rSa7wLKvbQxCmGf+eklcgPK1O4Ic0ugdpohreATwaJK7Wv5yUMPVZ8w4JrTn+wh1q5SpCSE6c5v
34Yi1qiyd2MolISJy0qmj/2YHSASNAV3BY56VaQas9l73VZkC4dx0WU6rO4pGHEG3QSZGJpFaNTB
crfZT016GorAGH8wIpAd8wEcYPanaXyciRXEwuWqRtX3ABZzBAT53pQB30FBWZwv+TEQXY6uITYa
aN/vw385E6PQHns7Y5RpqutGdczRxdWCiQKV79fewg+KHczx0pghlcO/D8NACqvcuSgHD29eBqQ9
8aPnuNKXtXJ/LX9UTG4fV2UQK351GuOpGolttkv3H371Mb13YSTy2RGCpCLw8iTGtJZbdi2rIeq1
bQbWDt1AZePhjPPG6/6Ie9bR17WTYHlX3nn9AsMSqtTGBWWNdN26TOwbs8d/ETIW8m5yb70FknEo
CG6yJImgOLPZjJmbGOL7W2hQxLhU3XQ7VwNJ9HpbYDMwcbIpfI2k5tNEQ2UEjPwsLDJRmzVELcrL
6fjIr5z+hTfV4ZuC1Bilw4DRwUHkRUhArzySYYp+8P0yBhncUnyu3TkBpSjpg/hew9lY4SP5tAtq
/ZQCDYAvKDyS3Oj6Tjip2Y6etbXJA1vAZfiIB0rDmEEaBBOmsYswGhJL3IrLkDYBQ2tctYl4OmK9
GqVSxaVYtISTllYJfXspkzK3p6VSHUUrno3sb+YUK62+0UV1MEsKW39aJi/Q7sw9Pyo588oAajzs
taAe5jjAa56ao97tZ59iZ0xzoBgzwfElUSMWfereCHFtACR7N33zY3DIuUyvt0abo7wqI1PKZ4ER
JL13af2mt1pUuK1tuY48ZAhA0IP9ij5NU4eJ9FaKIX/qYXca8DmCh73hFPa/DY9609OKrvbpyIN+
FLN00JFZIy97GF3hFpXM6d0SYiz8PZ3Nie+LWfdRR+Fb2LrjUb9twnHYwyrk+acqwQ+Xj80W+Qoc
lqadRAgs0gazH4B6RVIRM9WrSQqtcWcXIV1Xj8zxJMNHqDN2dl9Bpuh2dWapyjHEAr1uIJXoxwmJ
nvr9+fvBJNgAsiAcYnBm5XYK39NynkroNVrRcz8xrke0xdGQv8lk5SIRrH5kl4mSF5fT6O/LP7/M
QvnkzyIG+93KwmUTwKzddys19XTvWuKNDSSYz/uotUcS2eZjGLkDbeVb8Yktmg/vqsRdP6ZG19oX
+9QssBL0TZYJHhakKhMjTr1P0XGrSaPCy6ZbH6djGDHPbA1kcQ4OJiqP8PjioInxXSqx/U1ir9vU
wZ5AtKMMYA3e+V4qtWes3PhnnfQ4/dCIMglwOkXkpMp03WO+5Jhz1Qo7tWI3fBDBmzWMLLBimjLI
jk+hTHJbX4rXxmRdeC15YIILwRbxA1Og9SZYQdj5BlwW8gt2/7x9V73zoqN7CXWbVLfIY90Oa9LS
fPavotyZHFbmEnOQkAOgavP+i0gtJ/0qVhqXKy8b6LxyPh8rN+xOpG5sn8oZUJhO4+1oo1cDetu+
EtHwRFF7WDGoVHBqIBgCfchYxIoFQ15CrCZcZEk1xZ32JtRt8Vndh5ejbdUxuZyDWs6VnAL2k23d
vNUnDeBiMKE10Crm7LoNjMDtOCvwRwTSvUXyg48+f25pd9zfM7luEBYnlPLzuMfpWQsCN8stsH+l
uKdFuPCDH4snvMX2igCIwOOY4R0S6I6kxgxzL8k1ECMr+iktHSPbvEEr2XyyIstbbzJDqKnxpeuK
GOihoGcgb2/c0uYX9cZIH6z7p577ISXf9G1KHXJeKU7iqfGmo7J270IYGO9dtq7wsBBLeDJCi1hx
mc+SLOaYSL/clcY8fn9wLOR4tsoBmNGkGp3yCb8U3KTTvChOD4uxqm60vTcHnPRDbY3Q/n8/HGTO
ajhsAFIAsq/yq14DQWbsVG4fFy7omJufhoqq+ilc0xJT64STzRD1xzBrD5W1iEeMeaYAhgEaOpW+
oz2iATi+pT0ucRZZSGoe+GBgFPjfsXktVClKsQuY84aoG0ERDqgOUcYZANi9BPzvWyaLiuy/v3Re
JZGXGy3EtTHGMsVndzm4hx1q2cfEhP/mnr1weNWpbwgqpMuVN1GrftcHtMfrQTPwnXlWxSSMmaFF
9ObtFHKb2mkURsrgyks49TB/t8NE/Wg2ZFJs0BwrE2QTo/BzYwvoEEC5v24upXfoiQB9LUoXFmnO
07vWYnTATNuiYcQ9kfBlWTJt1AbeQWfsPfzQxlrkYdoASyhuSrIKBQA3D7tFuaHzL+f4ue4TX+V8
8qNdnrp3+OKQUjCQqBqYPbAZEpX946JCixZrNnxh0nmhSBlmvwG1stSLe48QY10eJhNYIcjmZRDm
4DzOoEy7jHMPq27HnChwke2ijb1jzUjurC3CT92NFNRefbbl6P+XsaTnyFEntwaVMQMTIQU/bAhj
fyeovRZOMBoYTlMaMQLbUAtP7I2Y0wHQdNPySLIJpYhpoindVwm8lGIafe3JHHMgy5ZF0jQ8Zj6k
hIdOOIUvu3SP4xRUOha0Pqs//lQoF7gcQg52pZVjR7zAajdN8vWFdx3zJZ8uvWE67Aa05yOeepCE
46puMw1XJDcJfWjhp+DF0byy6h1URg2/e8Fk9Dq6NJ3jKDY+3QItCNlZrLcxXI0kaNfQ4JeEQpxA
6PkQs4N+ZCsoxeMc1xSqMvMINZLhzm8INltV6voubSZVsaxrDX5Gl12k+IGGVsCh1TbRcv5hwEAQ
Lm/8nLzTcSRcXMcQ5G1/WLalVy0fXMqiuKJKwX8wHIrSISO/PrUlDr/8ZAXtZDKqDW3Ffr+S2NSi
v6MhHWzpJU9v04s4RNYOKhibRRLpJW5CfZ1dW0hVviYRFqG6oOiJgVXSa5nB0jKl8T0FUP/pnkpf
/qTmZTcJ5uiLu+ydDvXsCveGyA4h35TTe/MKa8m8eT6MdEhAyC30ZqVBpfrz4TUpiNtD6lz3op/k
kkWy/YIPpxRvdKGaHAymhAr/6LuDhsABZqoyuAQJ2CQxy56MhDN/+gjJuhhN/dzfj4XBM0z4603w
A37yaj/Dj+eCyGTVuIidzFQhV1SrVNFSHlmOZs/wuxn1YaYjBDiJcHVQ449xNk4CfJbRdnRlOCqu
KBqWpdeHTAGM2y1jEpYpclq+XgDBvPJiUBSRk4Sajr/8ID7G4o/qVhOpPY7wSk3Mth3m/I+XHDMt
eifRENLNZ6cp33T6QS1CYI382+lbjDOb7wF4b3pGn9Mq6G78e7qG8xSwcvyNySXwLTyCxY3aBpEp
E9IalvuhMCqzeuJRkiHKRK4Wr0XX3+6XzEgpCaWEF87L8YhwBLOI4gXDn/X2n42cR8+/NnAOs0Bw
vZ+FjgsAZEsJB2Ahg++q1Dw1xH60hbIvm9cexJp+7kIpTyDxX0OP58r/8f1SpYwk0H8/j/RmbAo2
zSsfYzn6QcXUHxHUgIWC/4D5IDjgapQSDWtNQ/8C2YFYPxEzZ0BdZ0+RMwxLUD8Azp5TQaH1oyHe
t3XRQxS/OPJykhCRBsxnYzZ2f+XGzWhHLSJe4X5Hnx1YcaBzVE9Fas5mTeK90oS1IV0SSUTvUg2G
iiZ7JAo/08F8tP4BHioYg6bLFDZESUWcYTuRTzrtlr1r+k812HUqQcmxxduHi1Q/m7hzaGLrGmFW
Uvxf78DOAoOCNwHT1gW9i9NlzaDBX3dFRS4BScu7SSoPX9OhBr5MTnmFHDUE/4WyUiaNxYx4zJqx
JXkDOCv0CGKzr79IFW43EjjUkMP4ltZ1rcNoePPdFmWZbdiVR5sdTfplYs6TItc06vp8VI4KQ7WG
t16ua8QbNh9s3sJ3ZHzEF87FZk1qh3q7e02g6KkzPq5V6aa0WP6pPUQoOPQKocrP9q5OG+l9iN0q
EHKinGJIcT6ZKpzyvbcYNJbo2RCDveN381fLxTlWC47oPreNr8Pkpk8x1WjfV7a6EtDLs0rCB59+
xLWFPkafw6zUu9mIXgBhtkM1KIoKEze7OIqXK7hQUEBuOInFfYrePVPlfKUPldd8+2onxSp0pRFc
+XoDMRSuuZJkHcRFIJJ15F0K5xshbTj+Telg9mFe79bGEJprdXzoX0THTjfiOA0mIzKKJDSuKtHe
bXLWGZieDwyiKMbWxpgs4wyNPXifgwg0F01yPoO5x50jCbD8w8ohdt8LNGq9ORs6W4kDYsi5qRde
YWpDt+Ygb6Ghh22Nmufng3L4gkhDB6JUOaVxD0jALwc4XSmwP1U5WEe5pUuyg7X00ZDgZ3O4ek3m
q/vD0PySixWhC/1TM4viPRwRhMe4vy/0nuUz0IRHWgaXocqvTGL7u2w8CHanzPusmHIIHfeQI2mU
dwYTHYkXCN5uOPUIA4LPS2pE5ACIii5XhjA1Hn9C35uFkZPnu8B3pz/Nd1W+j9WoVdEb4vjfwKm/
KfvOi+pzy4dYtLYA1P6sX2Hx4JJ8ymUlwOwv6nvKas7ZSl4ve24dGC99aopKpC2Ps0SGHQa4JsFN
w9vpleiJphCVqjVaQcYbGYiDkHy2nGDLFyVnTH9vEKLTJtuOYVaAatgWRfhCczsoBAunh4KgiexP
DyiH6SxH9sbqobf5rrSsk/HTXASTIhlbCcc5NLLiTlv3Pv+57XGxC2+Su5B42Xowdzjv3TMbPDG1
xT4084mZLQ709DKRqOL+F267mTZl6LWS/FdxuCC1EOLip4mvvh0SWg8YID5VMv4lgBxGXpj+J+Vy
oen5bLx/+cPeci/Mi7ioDmkaj9vajZVVjrgI2cntGjU+C8EkekqhGRaTBlf0Az6qDyrcdlbLDpSE
Lf6f3tqDy63PKP+yP1zdIB+WOF0fhWefudl/dYP5gasosLz7Mi23NCAxF5mD5bY9gP6nUXI8RfZ4
gWAQwcrbRmTDWZLlUeLH3UBcLxPmLav4UwASyQjbvnSYbd+7E21lW14X+sZuMe2Ut38IBFG15mOb
JVrInoPYI94LknaQEMfwPFjFQiD6FqEVRDW/+al931w7fz88vyEO1yldJh78grL8oi3ZvyGbPsYe
9mOTk9H0Kdwg8eL8vPbNcoOr+vWSMtG6lz+rtnNLuSgaUiLbkyzrKnC/WGcnWVsvCP+cWelZ8GwK
sZBMqROfQrmxOZvHyKS5FACfFz2CuH7dRO6Eh6FPjjqAbEpH27jEfLcKW6XsYDIEIVa4G2cLzrkO
4TQZq0YEM5I4o0fexAEhLqiKyXCC56YcPXh4uZKUBU7Udwzb2nV6JNb9GiKjQTDxc5TbHHNfjPTe
WgydCTurhhi6rZQqFX1QJ0JVXdXP7VMl1DlidocV8Zj5OIUngTWDWwYp9/PcRg4lRc7m1XKj8MS1
+kwh7IIe5GyKvcPpyhfkoJPuHmu0zRWz3AucoqneSjcS1jxO4v/jKJ97HDnOeoiulEWyasRittCN
Mk3DdUb525gODX7dwBN+Mtzh2Qap+YwDNNbXlED5UMC5qDIBbsfqj+gK30gl5hcLSC0GOHD6c8UL
W3GFXloLmHIGNCIYoXjCNidlHdXLlrFBK7Sg7h664HrTYHSnYTJUvwGL+FOwEM+pqBqzkMvsqfWm
AwXm5reRQy9X5FVJrmIFJo+xyyfu45/Fva1EIqk9gupx/Xq17BrhLik71Hmx86Rb/JXJ2JSBQtTw
Dvj8SziDfZwAlUPtC0ddKYhnL5Ys78LXXW6exD6+hNP6BAj/9CP7afHSRowCxZZI4aFJH9d/H+Og
Jie2m+RMRCryIegfgr98Kx3lK0U5/TTCgylc89KRim7wkKVFOn+l+SKTpISqeHUKUtIQeS85Lkvb
npiieTHgOfb5HfbvZxvu4qofj8raH6lRyNqq6lqufrfyKKqXGYZ/haI4kr+VegixHkESsC+po8rB
kFffypqko90zibpI/fWbrcWTlIEvjWEo9xuLLGl0V46FSj5N4hxG9/P2ZWrG0mGsO8f1MFCBqWfJ
ud19ZjiLqSdzY8dMsgHOB7L0LTWnN5UGI+06hZy+EG7y/5+gqLO9dhY+IyR0IeOzeyW22vUxn02J
UVe1iHrYEEA19NwWlqDL3hbtX82NakGGnlgjjK8I2HJAsheEpzHY7h0ghU3XOS9VFXgiMl0uF99O
L1Pv8X6VdrUjV5LWO/VcB3VeomLYXJYACa1Q8/AHKpUgRZOB5DSSlGqf/DQOFN6sv5VxG9nA59fd
FoORGFs1ZwF7E8EAstco4scg8Rx9MBojF1Wzd65dSEDJCOLmCFWwt1NMUJjI5PxqLLkhz+KQiCVB
j3h3Yw5e6bGgu1l1rm4XuONFY6uIGcO22A9kl6zcWK/RcTsYlm42hNjCNUh1E8Hkg0UM/3H/tiIG
fQaZ8a/xlMdZEVnlfLLKnr1hC+92Rkt9S+5ZNunOJVR7KSXLMexA9KGdRXQ/51DVjWtlWtZCw1yW
m1m74Uq1vjff9EjQ8764kBIOIBNOEmkOQLDeHNywdjwkXJkkKt+NNn481ijszpEMmws5q9vmtZ0k
90+l0z4KQKlTBcGUHj8nt8Kkz9Qqd/sGuyyePcCcho/gvZ7p79zE1HkZC60FhZmfFBtXGBNIwsbj
wjyXC46cyq9mmcBvI9xvOli6H3q1zhTDFFKv+9o5qfsPtc8ziMYfbwH7uVLIz09IoUOR2KyImP7u
o14z7OSHoXD8F+Olq1vrqhZP7VZqP9gzvmFk183bHk80jeyvi7psGL0qSqygvhw96pDjHFFHOXuC
ZgF+N60xte+KE9rfYQypn9oAUK2JmSP14AoPXts79Pwd4xYAZ35i0YJamx8XC7A8LYunH5JLIMwC
kErOVtTlKiG1jPZKUh7g/C+RiPWG6KTyuTiKfxtlNyXTZY23lhMQMWXYaDNxECnmJUQsBnMM6jHh
C4mGh96KwYZfWmPCsZfBcTgyGhEZ5XKC7keMe+oNlLLIxFRrZsrVrufbc9iPy3eLjKhjLFTH2/eh
vPMzEeuskk1AtX+rcgeLkvEOl1Ykreo/fGYWrEqh7HqSw/0d1a8KaTiJ7ooE5k1OySDnMzUuBiV8
FMHFs6liW/gBJ4pFrHRSk5gGB94OFCgPRiS4QZyXlR3lwrD08oq16dMeiB+P5TtEbGTbZ7oqEB8R
hi+vuRhA0BBnAWuaPIHa+cCZp2o2N0E2S5lKMnBrXaqIpYLn0G5Z9fNjk/tKYVwnsPrHJkGLGoF9
U3gIbEfh9osLWqWm91IGB8IbVx+qdw+HDtvVABkHXRaplfQvfnMvyj9ZYUBrfnWV92wYT7U5rL7L
g/gNB4A34CcgSujPzt/4TH5UZhZfTgkelQiPe/Ih8+0xH3or4EV2r8gAKpmam+o/8k5NMy06JOgf
d9yienXrQASNNJS8+pnvhcrRuyjPKFnYE0BpqWtXyfotznwy+EDIMrvvQ46+1blLqDfEr6+5ZGmi
jpODxFFTjStWTkoKZZ+g2ODsdnVa3JSz3BHd+7EAuXErLQw05RGbBktvFuOLKFjr4+dVgO6SQpe+
Eb70vnUhmRzSix20rf2XoP/Nu68g04MAhyEH5yUuXsisOYzwYdfaaZ3db4em/jQ18hZCCORVQhNT
zk8ABAAXHXf3egAW28gJfRfWvemFWm4+vRm8//vRuhj0FT59ys/XSmUyTDM600ipiKsfn6Fq4gkG
G6Ia3BWGeN+CzAjJgyyXD96azYhFmRPjaqoyYldsG/yZRu562cqnC/kJU+X0Kmok4WettZQvYe7e
J01NXQqP5916Ajgh+6qifIHzo94rfMz+wPXatp3iEEGKnz9fK+VXZVgDxZWIwLwsRJ9lkt65/P71
AeKqrFNB6aFm0IOZpiski2elOMykiturs3AV5ZhYIp3cq+nF+ka12CA5YrqgJ6RkM7P17zToLvxT
N0j13v1ioUE9Yn9QGRhXhoB1yhHmJIadRypIK3EyWMK8nat8IdBQ9zkLE7ZBbame9e61Qpo8MURR
PWc4goBkgAOgXLdwGd+slhhnKwhRTj+mPMLd5qGcQfCY1ldbiIsOtbeZZz7A7RHyXmmVgid2yoOL
rdidtwEh0nCg1Yhuaq285q0i2wYgVdF2bSF+m2PT9Qq3nkEPR0zDJxxdgZKjgadxWR5667MF/Gen
F2ob6If3w+EeVpXCdRHCOFa8QMcRlE4bJ9mis97QVkhvNuka7Msk0fyvoSKUr7leInmqZr53WGO+
PWPAPxUfJA9olBABE7muqxsg5xcRp+2tzCkNcErru6Zk/b5xtzXZ1Xwawtp3ZZVO+R8W731w8CJu
qqSUCOVqJSm475bLcIlGyegiGmkD8OdP2k9keSCHxCcz5yyp4fzE++9rj39gqjqS3dFmnIT1KfGq
XJfSa3oLxk7tteAilpKvEDzJZzQaICn4XRpXnHyvTPhRuDMm471IfjFFjQ7F+RfryoYw6iMFjofC
M2r85ek7dE9I1Py9QxcnRA6gitUZTeOvPYOZwtL+UAu2QDs76WqyGgAbNlWWqRhNDOKtMZ5RiuED
ze+5DNsTSURyDILOo94BiiVIifdMdluCe5OWVCbuzUGRfG2qWI3uONsi+qN2blijeNaEbnnfBqnx
GdD/SXoLbxI43azlmJyay3xyLeKMFDtiKFBwqTjOZ7mEOa8EYx7FZG2pwGxgfSg5pPyBsINFB/qR
YmED3FwboBGPAEWeHBYqCX5qz2cnebRs96Am6jgJbiNXgnB7qIJkiCp7k67Kqh2CWMWzBV8Cd9e8
y6s7AMNiWq9b9c2XRSvE0MvxZgdq9pkB7JFDQdJ+oicAc5jyXdhzJyXnhgRgvPqHLaRrJg56RF3J
jF5MwrFDjdrf8WaZiUFcBcwXS8mekdb/BYVIpHATKZIwj5BNyH6VAdAXvSzNih9MGa44+wAHZ5io
h1jEV9JJ/XqtLxJ3Mi/hgOeBlj+pw9paevslZv0fVZtk5BSre+oSUWUlUh6nOqtFREmfAnm6psOL
t1ZdG0DIQtoYmOw8OxLZP2PqWShsKoJbJpZV0C1vjtxrM/EG9mqp5mu4dsBKzFpHUnwD3VTAH2fV
334RfRmQBe2RawSPQX/nLBdeA0h3+JygO0kFbxQ/p32nAgekX/P40duSk4aPFKmjPKirSNTG9XXR
P+HFZZCqHkvQ0xcWMTNZEUJJ/TcLr1WxqnYpP3S9zyouTg3iZC8LRXj0MURxyOr/TklHqTBNERQ9
1/EK9if9Ew3iP2Y/4Ocn4WB53uAlHSeyguZDBhA85rVmGLpexEOWqZczxEA68dO91hORk3dlzDL6
nTTw61gh0BMjYTM9bw64wCAy2VEAQyqgCzNggpqTHunZ7EQcb7bGaAOlCvoyGV+46lCBpK/tU5b5
S+H88q21u2ogNB3NVg38y6+mYmD3JdxhQ/x1I/QiDtyigIdGL/+SYmcQALeuWy4dP1njSKxf7kDO
/IHvG05OHRdfuAGCnPNLwjCzh8G7oQvXNB/C+kUmwMIJ16TGaeEsuO5vx3HZdd56WhuqmVpc07NZ
Blr52zUbogMBov4SH8rP4JX2jEOEMJQ/FzPqfsrNv8yZE5d7Wu3c3HgeVECroSS1EC+4qBDupVje
FfeEL8ahLj/oJO5VWpv2olGC0zdZoRJS9VHHiYBLD39IC3FBADvl7OMYoOkG7H1aohe8BkGcbsqZ
Z9MTUCpQ3DyUYb0RjldCtkz+8EtOv4i2fng/L4wPuDczVcgFh7O6K5pCSxbgSwYU+AHvJxvHuWug
F05Jy33L7i1v1s43mE1u7/AuphWzGk07guxapVvbQGMm1gvzuegOYVRXwWhgv/Xt3FPfi5qlckPM
qjz4g7kWAKZe3ejay9tgHG8Nv162qIkKcqXsA27Ycb7FANyRHA9gZpdB1f+oXGPrM9jedYShESFa
sr9VufAA8Ar4WvDs38q8oNp82acKr4q8B+6G9hUlgyXAXMj3eK0Vf/HntmQ/5rG8W/Bv+pR9tgPQ
v0SYzGBYCrefwJuOYp2RlBQ6DJYwX2EpsSXE0j10ZCIfdhBkEhFYEiQlXsRcgVVHFtWddYlOr20A
G6rPdJVb8NqYTp79Z7Dv5WNoCFQPw+jEI912osqxGhDI51N852435K+l+jTpcEwkZd5bUCFOkUYk
zLu4zOn4Wr+vx0aZyVstHTfJPZfTTIe8qsx3eZnFOTupZeLITZrfKHVoVIMWeNKtccyG1GbOhYCC
mB5tPvkdkNYhjENbX5mkczXqKCH4wBm3yFRa1WYbA4PZACEBbZWv//5SBkQ4y8di84NhBatfzHVG
CCb7u1fdpuA0MYuh74rt3AZK8AiJnRF/J4XjyWKAFSTAVWfbuS0OUkYBAGYO1d8jP4f5pEmKZIlh
ykKkON69E4KF4+WjVtvH2jW65efRIqsNMguP6p3LikMujQUYD9m0y8Aa/tA9HegC5HCVjCNn7HrJ
yW0eBgwX0lRRikZeR4j4Cbnjf8D+Fl+bxeYjloRoyz9oeQxiyp9e17fKJXMfESLv1MgramdafsP0
kjcrL10dq7c3apAcsE6KET5WE3+D9x2eJaQO+jHVeqojMWs7GVNM6yghX4Q7kA67yU0zffR1I9YV
4tM7cGGd4dEZghSffka4QlxStEAKmo3xLTOK5GQf5REwSyYLYEAGtBsXBH8GN3hNiXq/wNgaIho1
o8kkEawWWyAG0zlLB543pPByjXDeQCNt8Ka3mxh3Z9yT5sXE+pYtmWyLDM81dO6wWTN5pgy2Nsjt
s7zXLyzH6Rcs88ziz/j5DfvQk6PIpMKM3RdJPcGMSW7fDM30W4p2I8DGsJGwyRtPcZv/QzXasXk7
Bq9MWqgZ/iAXIESPdv5HX4Ct6wM9jqgLNGNfx1Z87kUvaJOL5NPdkGO808ixY6X8UoaBTyazPpAq
BBmJu2NeUqhxt5rUkLJKAIal4uNkU4lS29N685pPWj+iFI21UnD6g38XMjNv1dnMtI/IJsy31sSr
+QcumHiL1IAsN2plW1DsBUqmb0p5awl9S7a6dJlVbBxflVQiIySBCqb4+VnhIQETia/Up5NhTk74
WHDitrr0LpPO0rhqPVxHCFPImoJ33cH0t+KrshBDU2cwa66PZfoZDf/g1vci4Qzn1kGwH71HY/P1
vFZV8j05WL7h+1yK/0e0mBk2RPWjp0fd7fMVnWRAqoW5rPBTmtMnzmw5jZwn9GIW+gAC0IQwRac0
N4R8ArehGadyELkv7t4R71PebE4i8Ncj7ZirLHdqRrzGwTp2A92Uw3QjJoeB1CutIB8zRXPcdGLA
v+Zf/P0stdYl5OSQCzpwPsRH9sGb2PwkzhoXaQ1bec4xDpOzg5h8xzT5Q3pRyhdlgxzlQqMjitnp
KdWStV2yuQOrop14u+jOxB9/iTWQjzAOwOj7Cpz7dYS+4cqZSOB2+4bTffuMv2gGgEIIg27efch5
kIKgSTlSk9+xRzDkvb02DrPMMlgtMkvdmc7wn6iD5MA9OUHtfiSbwbc5nxjh4HWTPaWQ1G6BAbUf
hZoAKlqR/QJQDEBjg9Ih+b1xv8VUKTgTcYNRrS283vUsMhQYIVJx6Lk/EfAoQ/OkuMBOtyHtahb2
m0kHqSk9PoIov7RRK01BcB6W8hGo4288vvEJiR2Ap7EqU9h3gWijpSqMhM74lOMeVfF4xZM2f09n
BFyjdXcJ/AKfSA+brLzTfMuFCe99ri5J7gAMJq4T+8RQwLhyT4tAwN+2Tv2CpwyBQRdVY8lZzPEW
Te+2xrvQ/5StxTHDZfigSfD1HJHVJ1lnPXx0OusFddhgUJRO4fD8EAInPusHfynMzE2QTyq5HNhB
ZoDwVc/EYlAw+e0ttJxUTiiMAqHVcDOCJHkW9hD7btA61oQ+oS8VSSun19KK3gvQdl/pFBGaSbl7
ru0NIRjhr74CUh8I0JcdRLIZViCMCiiUWFAtjjg2JrAu226vFBC4RbD2tLlHl0MPM+gXxoqVUKio
zaed1vWG2hh9DkP6Hwtqf6EohmP6Jv4e8ZEmjZ2dwFoi+eAcL8shIhVWdJdWkS9NFB1TjspzabMr
ZxaN1QezCC0cwz+lu3nCitxYq8rSj0O3UNdt5C9PJpfWOWYPX/xGSRJKPOO6nBT6m9Bmu4qUBXTl
miCHAu+4gFDnTM62smxFEcrBjBOk+5d8Tq08SNNyFRws682SUt+gkJzVUqfT7diTfu89EOlYgwTg
weaqWdRK3ntgzKN1ozMZ5fW7hSD7UQyTSIAoAWEV9/E6WjAvlTXiZ6BZSOYfg1vHwdw5e5SiDfmb
yZMThOzBsGu65YqinbbOr5q9paur0zk9SURUov8HHJKJdjmDkgmk9pWE9yeH//opA6tc2+esuB/5
nAs6cbHnBDbqrOROld+WcETQsxIg0KIM+nN93PD5k95rl0KJvjTkJoQG7gC+NwOUbZIw37N7M+T/
NukkySEdjxqLR8oHKX0RChnOjuHZflaeW52wsWpE5LB5Us1WP/H4Koxsp9nEpzMZtGgL+uhwy9hP
McrjpJiYcgqR+44z16EXyv3pxTuuh/MPsNXXC8d5JAK6vbBAbi7f8exVv979hZKZItN9z32i2q0t
AJA8/7KMUxBGVagXJ5qfs7RRGvwhs1xGKsquIptNE462Y/kXnFvnIsZ88unJC/YgfxJX8E2VgCa7
PR8RL8vLZJ/XhLYjW9GNbtyD3DfzvfCPlPnyr715Vrv0ajksgkZxpv+DKNmObnYT2N1zo6govRya
P3kHEJLBHS34EqO0B4Ua6CBSuufThjaoXYleXlbcloGlUSfaUwSJ2BaKQooE2zAWxpVcdhOYcAeo
elExocGhawLHg+qusDvjNxD+GieGTRA0vIMxBFeQLHp8ZYSs3fLltE7fYYNTDsoVYXTAl/3d76YW
ug2Wt4I3EdPXBMdKZIrGUrTT387KGwbanjBEkbHknwrCPaH+DGvmly2DFbPCPp/lW2Ph7jv4hpMD
fVEyCQCbn9QSzFbQrtwBjMTngecvLHHjcH2z9COXarmAm2cwlxTQqQUpzPZxw8UnKhYwjneoCbzo
IOxKPlGkIgE9EjeTodmSM5ML6C3FX3VPLqK2FfgZioMHqO0JSKxumNzzzHOYJnCWiYcHnI43vrGl
KhkbfW11ZqSPcI/g73YcRWBF8WSpAcVnW1AFXmJEf7O5tIOTCCG9JYjXnIKoZBoiyCvqra2zIS8t
S7D262K6LPmELdWWjhJV4p+UryhsIvQgWmkqtl/+6PVg7UNeEdTY+/Y+Do7huZiVRtKgwGB0VJRq
E+MBFmMqUigA3tqpWMbtl6n0A0EwOyLKODDQSGTYO+kAIgTHLmBD4ctIt0dXOadKTAD/FSV2QJON
x975CUXju87OPOGMmpQa+QQlilFRyIpBLIqffjlX9h/J3MfWH4MOgzOSykFCgLOikPMWquUyN5NX
eQBn2A31k6ZFFXpFkv0LjDMw13g2H/kR4eJMIlusp87++khXP4lhsEbCWkYKWcDIBB9g/G/ByypJ
Y3Hmb5IvjpTg7aQJZVKT0o2jXWLj3QMlm5ZF5qOIrDmaiGB0lYeBDOIX4sCHJWUHqzTGrqu+lifo
wYKhyM7cZkGr5kaibxoEvB03eR9u2JkOqIc19pIpH8F94fExNXNtxSGqOznNw4L5qjhLObfjBxEP
DZaDjmpynQda/ngJehgzc3r54Jqqt59jQxQBvrneYxc5ZDZWcnXHAC7RbogEtpPIaBRZp+CtPhmZ
3JtUrVCjfrvpy43sd3JUbZKASV40wstPvS5+EMfoVEgN7ZhFhv7YPnudKNbNS2qmQMtwxCNf0cWH
vnk4ryBB6f7pGH7l1zKgUIBznLJ8bxjOE4B7eS4/hPDjwEYiXCp43Yfe+TWeh6S9E1LxBazJYBsg
scqDU4pXZDu143FruzP4crt7Di/KXbQaSkAnOxYIAOsr9RpqmRYAcpzO9xV3m8dI+Zs8OoerchpB
R9gQWwuwdxLOOlNowGOCpYU6SfAF4Yo+M0FZr98bFoZ2QBkm8gvVLAmLFFGkqf1IJs+K2nQCpcFd
N0FjEotoi9uRmp38gmLlLFoMcsxKrPaEJOKtfTj36D84oAle+pZpjmwylx1/zA8wOFOYO5v3aEDe
Yjx0dJhPgmDtFO6S2Bc8/x1jR9B7uSAt0ok1+hTcQQTeM4qA8cuFtJ765ke5lkqTtM4A5lqdsor4
DjtISRZumjr5N6qOBw3aOAgDxnPlAHHUwFeUVweRtmrTGpx2aRUrrvz8Kx3QyC0ZyCBQacIEIGSu
yptSsdhp/vGk+Q9H4uBWEzpvZPLCR4gM5i7hteGz3Xc1D9nnOsaqh6OajdCejThlgOOf3ofJMKXH
nb/Q30kGnXiCI6n2PSxo4sACnRvli6Cer+zHsQrkzXlCLhC1Kw0+MQKcB5cge8fieJUG84VjEFQX
bxyO4MZKTtnGh5hcvjM6XH0MrEW2gzuapKwjO+d60/BnuYVWP+PWtR4jNQ8NiaiFE7jSSYUo3Msv
mM5dNgms3Ut3dIjrgi3V+AeEJr7NPtGVD9f7Mt4htdb2ZvX4/0anmGdhik05mDFpVV+q3NM4pjoh
mRsSOttXYy8TkA4dov5UBvI8ozhSY9frm+iMDq8zM7F054hDcjHR23vaZL81emgSHyewGkJH+HYP
SG6mX7eZl3/wujZcclvWuYWFQIe7TdJQYJI8xD4uc4aKNR+FIJ82y011nxspQerhCUFIfZDeDFci
AOSZy9ex503Eh0+iyQzsvxqGe2J9B5ctERprYIP5ktNvObfLt89rmDETcBmujPMva3hZKenJZZMg
+5TF9ZtRNgBMzuqX+Jvtki669c3xsf+inGHMDmLERYMP6J8aCsa5WwzAItWex1YUDMATQ1HIOa1U
V+u8b4qhTdlPb1Wi03kh7GHXUxSRvEEn9aCHfwfOb08YwwfiQCeka1tyOwWZ5tPDDl94c6GsoWCs
mFXIENgxdUF71cHQJIJyq/wcRyt6S8RChArvUSOobmn6up1NRWw1mGNfrf6JymDyq5MnynIxEa34
nVN00h7zKB33bUKiY6Q9Vii4jXYE3moG5T9peNytv5nMP0olT9fwoaQPt23hePY+RSLNOQd0G9Hc
NJ7Hfsd3yX20eWy4mfCIAnUJgG9VRgW0tkAv8g82X4magEauHl94P1OU0FZPqODQVNl2A/IdKw28
21sGoTzfDbw3KuFDVzfpj+n3EG24oAXZgQmEbkEd9BgdNk4QL+1f6GEoqMEXZqtyG5M5ghbYhAe7
0ThQ56nyTXgaQ5eCna0x3mK8oB7EHDzi8LfBaiBQrL8Z6Lu1g6FgChZOutrwaJapFwQtlip2H2X/
NxFruxGaHFWYi52Nv3cf7oAEybOCs3+6Hoxi35FrJG60QpSVH1p+1RUOAVb/0vNF1TT1B8LQmCwx
TMTjuArd9uzWRS+vU381GKLYPoX/nWYAXvzlCAzeCa3P+Dt2G1/Ty3szZDvw0FstUsX4xo7KTG/4
7ii5UrTRDt7r0Znycnx/ECB0c/5Ws8LFUMYoIJRefqC7W+sM3kTaOCiAJFr6zjZB9u2uFVG4NQRE
lGBsOfl4FwhnFqima3+bapfhEMF0kxOpUgGFrl6MshSsXIbH+Jiyuv8wPJMX2eajiZSd5supc07W
ucIGgmFYPuAltJ11gjdpFAciRs36zd6xqshcyry/qkdS32gz/mNMsNPehr9ITKl1iabe8u1Xw5Lz
od4G7ikg/AYlMZXCaCwS+JJZj5WeQ1Ek6jZWlKQ/bLvY8g+S023wIEiVLdsnf2f4+AeKcpC2a0GG
f5tWXe1kvC6GM3+wBDJYVXaxNRpQ2Ck2rqbCTxYhvdlqQZGc7LFouTpdFQiOFzRzP2UBW9W2ygNK
lfnG4VP+Qu8gxEV5Vo047Q93It3iNfNEXAPo9a9x/tgylxEpOWfFIViC3D8eySRaiuXg7WXHF0gF
goNukXBG//KqmCbx+xcu7pZWr7Pma7GfwwF65kSq858Gk4vpyISoSh4w/NZckFbFmzDe6YaU8KvU
XjrC7/q/vqNr+jI53uv4RlZjzF8gjDinujPBGiZ/Uek/Nn06mmXZeZpihNvSrL0CpME5Ylmfk47L
hgsceToHRJgfW1GMMkGBRlaH9+JVGsa8kBubbPMqJCAj9Ch7Q8S3rHSyen196/u6jW9E6gRT8l20
WNmihvZ6xqTv+A2F3kN15hqMD5Zgcsax6Ge5KuvmgqTmV1QloS+AAB13A2KtfsLPxLoMJJnQtClN
Q8gJAG7h1RBphpR2IU1F7OCxjfT8BJn+RVEG3VKWT7FQswz7XefZ9PGD/NKjBhn/im10ad/hBU+J
6sZU9cZzHl/BEl9I0UuWh8EGz5b5o/iqIs7KJty5daxa12WgIAOKTPvSwfZjlbVaku93i4gJMQOq
j8S6Zkazdp1InbK9kidS1manJ06taSr4qoevTYg4LxhrYS1qUtqo1R13aYVYzgVpCbm2qJrWJOHm
IHo952SHWemtzqE2QgmkmUa7K1rhGOyL5MsW+hOb/B0bef5g+WPKVQjIVxKiFmBiqqwweIjYq2ft
puUYqG7aNPb2W3cj1v3IiABWKTq+UjcTjj25p8BS3ScLA/oIMHU1n1fcjq8oqIA+E7BUjmuP3rL3
iRVtDBNFeVXcEJlJrbLJrqITc1kvICv8LjhyY0HpC8akZNSStgX/0/7eXsnBPlBh0K9AM/C6Lbp6
dqhXSjPJmKreLolmN+NTRR0vdFF/v5sJNnngOOoaNuyvrqOZe6CaxUg3Ug26Bu3m2lGedsvzQ0t2
EhKmxPV5doY/JrxUOAPPV+TUilpUTK/PAPgNSYSBHN7OMdRhXDdhYCagtFDN1fdBYZxZ0Yrn8e12
y2HNNzpv7J6+/phrBqkD6oJwF5tjQutTsH0IkL0+Q0bjuneRn2GCFX2e9T09jEU9m/x8zjdCESfq
7PyOw79Hm1YnQKqGO3HlFNg04hrjEFnzgp6VxqNO6FVizHG4dsxo3YcWWYKNvyWD/d4U1/vw7wEQ
Ky2LIoeu1hhTErQsexbb7I9F4sfEn+mAwG/m96Hy8WbskFkgODCL0X1zuyeIFK30Na4h4rUrYxj8
ebfOV6o9bCcywL8bt55LrnUppCacCwuYJIZI4ZB+3CvhEfhxYRn8TVXjKN0A1o/6swt8Dlsg13xu
QMx5dZt0Ciuy0nrjgsRpkVXA5nsfNmZXJFWkDuuCMKO6w15LAN3pOy3LOLBQSCYOK0WT1llD1wBC
BU+zZrVoNZGfGheS9q46kJ4Qh+eLfxwF84k5EhQp+3gHLZVRjf2oXd2lIoSsGt3NQgGoQS+jUaNh
ZGGKAgkvmtnF6z1N+iLGYPSHz80N29JW5y7Ito3INjgRSYuW9Y/dLckjYsLPkxm0TwA3NKltLmj7
dswBd7sTJpkepOQ7Ol5LSS08huaqcwTTf0o6HGXUtfCNXEsszx6iv7wo8MVheXZEsySzQF49W3HP
Src0bRvz859XrjGFVgoiYNc/y5ASiKisHqm4Hq1XdFxLTxz55p36vGZumhpFnQCvheiqEtEEa0NY
UCGgDMbf6uglXubUlL1y6bccb4/BoyzLSEL502Fmc4hlEUGrKUhLjXIasSl8/xSiRbv5jp0R0xNC
XVPB+s9+MZwD70fPekZTBNaDK21dE2Mfq05TSReeBGqp2KhuXzvP0BUnvl3+1MzAHe5stb5noUXZ
QD9IOsAeAgbrDeBjIQ1aWZAXxBbrSHYlWIuX75t+TRaOJSCprHT5RriFh+rtbWVsWNBcPAw7PwJ5
2xhuGAqlSKbz5FwvS98coD+uPxghnny2BsKBu1USXHyKj4TEEHLZGvFo6q1Ktdnu7MKuUDEtdhfW
/RyMj3hzrmqh3cjg4DlBvdRNL22BvekBNO/FdiqK8D1ZjtDIVIiDCaCxzLBeDdY/v5bvZYgz7rVH
xujidxF7vUgLDM3m87TRl5jGzxBKPoZcmV0+oKJZ8EvjR+QwOjn5iSYeKsw8DfvBixXutaKwhfCk
8OlXxWLG+kuJi6vGZHeJt8GbXVRIRccx9jQ1f3vl/NnTqpMZWJ2mS0SUvj3FzqdbsOP2gKdz6mb9
7aLaZMvWE0j9S2wtbKDbUr4sss26o2tmTexDOjw/Fj0w/lLgtK3c7cgZD2z6IO7ryMwxPkmeeyBB
dH2bJ73udYnCGKQyXstgZ1+K9qHQSTMtygE3zIxSy+H18Sz+VTiUBOLIL/jrK218c/+FZZ83nf9l
N31L+Td/gNtqzDzOZ+Xb/NrWETNZggwpyKHPVUCI3UmZUNNbaxdgWYWCGq3HeDBLNWNxDJhjY2W+
eD9/2oCvSkmFgXc9soj0quxKmP00ZGizIA9IZh5G62YRnH1/PbjWNJ/RfmQWXKvsvl/a3pRWztmi
bC5WXif/eEezy6PGd9sVx0qTSKo/V1rdtzss5zL0xZF9yOhoFcPKWLKLmybs859nZx2Bq9SpSaXO
Wu80XCIiOkPK8VTUXq5uQQKmVFNqlefW4lepDmJVEz9fDxBLEoyLAJzOKUQyoPUnrXGVnhAJTBHk
My3XFC5EfzVOgANrJoIivgOjun7LuhCZuCjQuBrWbMKI3GiDx2V3vk+rnBMcQv4cvZK5E7ZQSP8i
Yv+3B6690ZhHRAfJh8V36YI5R08stKdtOIyjB2AAjMvmPYRpckKqjseumHfoJvdWkpAvItBx3RPQ
iDY09qO7yMzqqSiu6iCFqOyPwcnxLdrcNrWI2TK+Z4C/KRwmiRwZi4n6yGoyzJDN9pM4dwyS4TLM
pRExydb/o03R1OID5DvQzV0Zc6ZfxuSfxNNdZEEDH1TjBm67Bhrkx9ZcX9slGyJ230BnZwH4b5rS
+byiUtoC2hj+DbdVoN3xo/EmP+wkauKhGdOjMeTBXej2opmscz0AeXbYjEgbv/LulTD0v4ugrkDy
WFDSuaURCJ1XS/8VIX+cxa6ZkDAWG2+C43aWwjYTl415GhtdSd4Mwio2cEiVO9YxuYtdiNW2zGY+
mvdk93DBw3bIco5cqTRuP9t96D7W6g/JprvLJWTFYNo7y3QlOgGxRJ7PQvZi//0sx0wNt3RWWiou
vvFHnb3AREbiXudM1WC+JNyhSd7YplbGPGBZuO5nIOEgdNaqmyXAWzKSGZCz+Y1WbX+TpLtUOOzS
EFMhk+vJUBVVPojnEMqwWrU2siUGVJtnKZF5ORx2B2uYOliE5Z4Pr290p1vwBbzb1AYJBonvcBom
d7ddYLQ/PF8iclq0iOC+DV7zSnZGJ+WLvtKFRhnSI1fSHi2JONTl1D0gp5XrJzL/vZHx5jze5/ci
t0+2Ta6drHJ6za2qtvNYnzgrL13egQykEFnZD6IT4I7rzWNI6mCL6dzmnE2IdbP4n9T53ox2dEPT
n4vAE80Cd/BEbUBrvOML/SQydBnoWfsb0/q9O5UQjf1bTjTB88SNzA3EjmBA7a5q2ywTYX6gTFkm
+gYLGelmxK4L3OPQ/OHEESnWfTTExL+MTzNB7n09SuZzXEGiqMumOuXDj0K0nLuLokGKw7hWSwrf
YBjFacdGvVYWWpaH4OPWyptkeNnY4bBnDuwr7tGpjpV2YKikZiuYNxYjPp9ENwIOpIe6w69+p0Qz
BxaEwWSrPa6W1ynO9Z3r8JKt97HVBvftW3yFUjKh6Uef8mO7xGBzv1c65hqGhMaUqKKeGzF7nhcg
FmkAdkVH3Sqy9baeWhHvGqsQbAieex0X6X/CIgDudQgBMwFbVoUenjIEM9tmCyMFeJ4211/bh8IG
P564Gxm0dB8x6CcFSpMYfDLqvqbKV53MjeR3STW52Gz2RXQh1/75KXUXhDPtNJD/MAz6y3/Ghmof
zadg7UmQuRofbYDCH88vtwxCBxwdjgA6UkVcHvu+nhpDu5aGQl6pVJldrpm8Ut+ziVOrkqj/bhfS
TJHHfvL6M23YtBzCVTpFJOEbfNMWM3FcDfz8idAVGW3qEdkYDnyzYBTUcDjRaSn/do7SF77ZMkvz
5VMUfZaTYp48Y8o0aje6868vbOHjV3mCA1Xijrh3aStHYEaIuGhHdawbh9WXtUs5e0H/qZ6rd89M
G+IfevCZgD0I5oCe6sRUEf/UhcDhgwwBmtKTkJ39IDaD8ozG0klyOEW5Q9zVFWrhl+2Lh6cCQJFC
SYsyDDIGAqVZZt+A2FYBtLqzZ0XpUgmG6yaLXOHefEOce6c24jejWNCi38JclNhWLwXWSjh1PzOO
mtLr2AJwYION16vlV7r5YowRmG6zFQk5p5Fy3WEAodc51T80QS53csOnRDI8+SfRJzfYmYUkT1ud
AellP9aeJjWbEkXort9VG3Z5VRObn40FWmp6h/1jvHrT1SAQg6EJzyI0HDQCRwnIg0qmuZbDAiE/
rffiFrAcv16TipVRBxMRB7eDPdKvteWNkXPGvdbcVHiEzjGnC3ayLMK3U20Z5x9Bcz+1t77j5WXb
VycDE+f0gu4kY4yG0Un2IYmbqABtqZYdaNVcsNW+I4eoKUOxHjEfjbTtli3bRHnkNqQS04/8wv7C
jVN0A+FVx34Q/IfwQah8NJakfMgkQ2jAE4wcVjF+wYZ9Nxlz4tW29/k3XGb67CAYHAyjOCEcbwzy
PTMg2w7g79M1WSc73HH1BxtVooTGd50cLNRz91EjPlk+PC+R+c5QxQmMkEogYnglx2BmSzpycsUd
QHhF0sA/lQan5M6od/4L+IAQe4XhYCmtUuCv3BomJ4CDU+fM9ZYGYuB+ILEmUBHtdXGzge0Tv9mr
Jar/KsqdQXaeD4hH7vz8p9zOVe0OwuYbHEdIY5LTYEeLzBX8D39tHOL+NeY6K7oL+7rRABUDGgp7
6QD5s3mrLgcv7jHJObVyDEHKrCyO5xHoBEXXsCqH3TNJ8PwZa8hVzAPPCM6boFEiGnagcVCDdtLq
Cswo01Lb3r3RNmb7JAcgW7i00He6BuHMlp8nlvckV6A5EyNyxcapk+OREi4CeoMNMtdI6zPqQ3en
X0Z0mAsF/dg30UP3gwtDLhg+6FM/fzROPNUFdXw5YFM3qkOl0wmfX/eRYRWyiOXBy9yaCGQEsUVV
AWdXSGkfHtSY0VShVywDOQB9zIw97yisz3tNis8M9rnttUBMsJM3If/Lie2MV+fUMuDyxob3uRc4
/A6qNYDyfc5Kk4sjXGotOTavI3ny7CkhJslyozqVR0PTLMYBBVTC1IEuV2C50AImkFi68/ha2Crh
NnquC58tl/SXc7Qr6qNLGurEXVbfQRE9CzKXQifY4B9yNiAXhN+4KYofx0DvGlmk73Qt2gc0s8lH
/JOu40rKymaepiXgPTIY+GWP5eTe2XzOx9F+ykOHs152eZAZv7Bldh0OjNvKpfj1JTg3EYqpaxhR
54a1TrpTxNoUd0lDSe9gzuRrNmED2n4hU/d85H8wCH0PO4bOFFHWeEDfm8ArzeObpE/n+nws1tv4
+EyCzKQ74e4CLGlxX/G1w+PVWVlVqQivEx/pBZ+1rABoAsQp5xo32itmfYRzGPCrbIn33woupjTK
1q2IMphFQZ52J0j8lC2l1ml4HanKwEQM2io/JcdvqchSrHFI9Anh5hHY79RDpX1WI39D5bD+JEk0
48zKYUNk87w/YKk/2vF+0JoQy2D34Up6j6/AyU+BC7Plt5qCLhX9UUVxZ8zl8DuPH5JS3x7oFDUQ
KaDTIT64uStw0OTH0HDpa57xDSaSqoD+/u+Wlwl/OQq2PHtTdDvxilM7p94TVpxZCq+Xjl9WnR3J
6KUOvSJsgj2vYK1tWCskmekJfwNwbS2F74QLce38nDxJFeaM5QqMcp7HSKE7EC0iTd5Yzop9otFI
WiQtZ8P6ah3GTZZamYtU8HOYOeTRW+OfRxnbnArIgLltnMd18MPmUKQEn5Z7IsAtGKBUe3Bzgatk
CTO0LsU5HptA3AxQkHHYf9pd6Cu0L8MolbIF3AxoQcdqRDQIHic8xWlbt22TYZacsr81BBEQ7LhO
C2SjTQXe4PS0sTP++eMk4P1KVhTRc5Sx5NnehlyCi9wMSTtxz3C8J9cJiuDEEgPbmVWLdurPWXxb
Arbn96I1OzIlowwsp+szWm/XpTTcUXMS+tfBDdX18Slo4Q7aw8HayeBMnEeXEKCiKsWTvsVq9l7T
m7YvLg1b56SWmkNotEvY+oGiGQB2BYdsHgPnq2hEIfiMsBkZ4jomvOUiHXqGKgspHGkxwMA/DhNi
2f6dvzLBf14gkdfmypHD+uvkSIpgOpacq6oEZ1mI98PgCduBtUAuZHGmPSaKy5GOz5R9uixMHJpM
acfYw1WBxwVOhgRkskyCDMY8utI2OsdzT0x0f0mW0CKiPlO3R9e0tMhKZnBZaGPiw6EkROD8GPVt
6I7O6Jd4+/T6t9SaejjU3Xsi1BgS9EixYFhjgEkxY19nkqbmkMVYIt7fNT5SamCu/mKaGpaK4D8c
ELW78iXaw1scG0TQ3xTCyQkshm1u3tWO05bN/IkKDUj6P6Sfs2g7RXng2ysuEv0q7qeyUV5WLRyo
Bc46U6S9hKRyKpcVS31G6HO++1/SHH1dmGIUzazJfU71/xM83nxcEuTC2L5c0tCh/LQmeYClMxAm
5sZTcF+bgNqAsV2YtbflZ4oNf5wtPjvaMIwFeH0qceGiIM89rOHPrn13jMOx/StAr9sae4m+vXIs
ZFAcz+5ZcikmqjK84AFQ1+3ub+cN+oFJGARRfx9R4IcBZ6z+VFyIEKQkisCZq6qhzZ0phN/wJOph
ntMHl9OJSvPS/7Nuy5NO29kkBaIMWA9REVBZc3Hz5t8ckjqq4SvCw5c2LYerFEkeXHDnjuUGjbEB
2JjxPf09RjRrVmL2gNMNxo5iMgrV69I4enj/rRO3BmdaWHPsKt5ohmk9dqkKTZppE/IFfcc9QyTX
OEWjcLWEpQaMpDoSoFLJh/psuuhzAxZ3+U3yQYDri8o+IiWgrQ6Wfn54SR/v/n0kdpyoEI46OKgq
Tt5dHeLYWTGeBAgsOUWVWGgIOvZWydCu2BWK1Py0VCBRODPfME37354CZQSumIiregYQ+jresRV5
IgVPgIdBbEJl/tPN+YEi8tIEzpzwGNjsFfwI0Ozo2QWekt5jCln0UGiuxEEG4h1xSUJnS5xX+v3l
FWl0ZgdC5Snzv7nSvqWmefe0es38Q/ARkdx7bj87lfKAgBlUK0AXK2TA0aIrVajaBhZn/+yLcQtW
YzxmMcLYWIJpTaJNjxTEJd6VDiPC+EfyoIK38qRVOJX5Hhm9/ehrsVlSVAjlaWSxw9JDo/qfVlay
XKgB0rNzGwxVdleDe8t8UDWIHMWFIxNI9FAuQ2f+bzPHKXy0qGSjN8Fbum6ExthuHjmPUx+K6ukU
nPzj8MeuO1dkybwqxOL1CAJ20JzUUtfsnil9jT9qCEJNVI3iZlss13rPL/gpW72NzNOKyY8zG3wi
+nKor6uxUjPGFryEXlpHBaDXfy53VrcJoPqeFWlEYkzD4K/hxVVHs7wDfJ5meJuArb0YGyBwG8Pv
GOpK8nlHG5kIerTLHlVHow0rzW2ywTmu7hXZX82hRX+yhO0SvehFJKht2y0GYzqRv0iIMW2BaWu1
ynFv9N+c4hGsvmv9+bo7RPlWezucTC4tBqL2kH497VE5nS3zkmbr1OIcrLYuueDTwSfiHdsmrtA7
VXQ9pXPk06tHPNhRtWNSlcRsGGTutRh/GrRrju2L/4OQ6x9pjHxBC8RitlQUwQ2hMubuDPf3ra/C
8kQVUQiO5OlLfb7mb4v3F2vtfuWBiAInLY6t+FjmV47nAyNqzQYizwHoyIGLc87fMEz7gAP2tvT9
Rucxz6DRgeZCZ79R8osbowpcVDfltlU4MR+jnXbx+H7Ce1DL2GW9yuS8QNhNMyxCCdr4WjGGOWz0
jpdf7XxrIsVGWuI5FASu7n2hmzqRwoxowdNqqLjKKIRmYoKqmTy63n0GrtMpfeIrgId9teSvH7GI
f646Nnl7M2b+HGKw0/te+DVupJ/SAPdD2FRZ3mCRyWtzRZipXhboYaEOPAi6RZZfUxk/tIESuCht
zS0x2uXlux6mCdf0mQPwRC2tb9qt6M2H/UMzOidWGXHbXJ8NUo4YeBx0qzgFdl2grryA5IdbUlr0
dBvw/orisk7LvySEOTfCIK5VR/aUz0t6bxyQ1gtzyueGshai9uFQqdYFVTUkT2kImwGhzIo7jcOI
YYaqHMH61Mox00I0LkrAJT15EjU4gWwvHwJjDhDN8rasjjOQWkpU7L6I78kF+dS47aforPwM1mFb
Xv71fMh6H7bxFoT3Kj02G5zCIg/7gdNBGzNRV35089K2N96k5N+PqiAFJnFx7v/9yqtBaX/S6Icc
6I59dxAPDBQ6EI09QZFWV41KO6Lek6Hlr88+twuzGkD6S3oy4E+KtEQj87HQFemVGIcd3QMolDUn
c/NNGwW9jxmAqHmB0hgkibX2z6RMbtHZ1bIPgOkwwu79of8K71Rp14FV1gT6mXNdkckIU1IZTK/s
3mhyn6XdqUqpGFjvApYXQtA5vnvna4zuLb1AoQH8OcbOwc4a7T2xbaGnV0WJ22oxgKtRKGH6hyhR
eW8Nc/i+IrSYFa+LWpsC73tZbiMhMrvLKPCPlZdoGgNVse0KO16BTk4pmW3u26SXJcZpEGblhSKx
HFzppAdJDDZbovhzSlv8G1SiBUd/hHjPGhe2X2HQL5iW2Ea9Z741sAuDOh3MmHqV5JIG1pbDc73I
d97kWmPgkq9c9ekrwwm95XeqQXhsMykO3unFBzKamV0BeSFWee0fHzQjA4trjJdh0QNYgOMOrDIx
0+CqU8ypxsIKDup45yZJSciNMaT9IHE2Iu0xsJ4/lbsX80GBUYn4gZjocukJuUfp0en2LwQq9VIc
uYT9mFEye3zhqhc6r5PkWLOQILeG/dtEBOagLElF5PLz3RnMAd3DG5C3C4W+xwF6JvKu/GbBYRPH
tR/vq4VtsrFJnAdWyfrmI8EIFvvT7bBA+4r6bnP/jfOCfBSmt4g3juf+PQv2lrANTIkW71AZFVX7
CG5MU3KPKX3N5cOYphJ8TB6k6KqWezBVBaStS0Zk6ZiKpO83JXu33SEhmr4Oa2v4uk2KXX+tN+AP
nsXKwfPmzNLL306NmIlqkzq58xA2zvxfAaodxQfmVMT422tLgUSeYBuNJSbC8DSV3vbcH7VnZDKE
sr9a8HEVm3TuL6EU/iGVd+qyyHsHAD0Ui2kb6pdu5OmnBw6deJCFZnOi1qWl60lGMIc5TGnq+QCM
ONKH7YeLhdESqp7zF13sOUlgvXAkwVR4RH3k2jQqxKHpNMgziPvrAy07eUlv9rrzx8oHPnIBVtUI
WSZtDlDWoDzUdOiSSlp/bkGKQhqoMb3UKbkLzlhdcS3PHfzxrpPQaaJsSqb4h+kMfp+546wEwqUx
c2NEDS0/bbDr2bwSxzG6uFMLrtMxLG1wVMK8X2JI9mB6dqIIPIClN2OaIPTotvvoXKY5Y19pwshv
dgzjFgxowHznw+lvqFi7bS6kzC/lyLlJSDVQLXVG9L3BAcEatYX/H8ix9ld401LatQGCydDH14y6
5s9L6iGzvNfRvS/+37zJ5iqtnXdMAQ0luchuliBgcTJTYMATGO53UqSwPL7ZxMPFQDs3XBSZWl4h
1Od3umAOIpOsBJ6oPezs9YtrGTFBmiLKQy0Iokozd4ckfPeyNLF3PIFRkPBkbLPNxs6ysTBwU61Y
PxYR5K8O+G2qq0AJomMtkbuCBDJq5etSNft0ygVxer3y/MXfnPoDAIALU61LuZVMzDpQYF//yCXz
YER6szEAk/apP/zTF/Pd93ortimz9sd5VV1z1rPAsaxlRJUp4B1D/i4oE6/IE3Q87fjh97bgwtU9
yBy22AggQKOf3AJwxHQckiGC4k3OfLEc8TcYxycOsAve/5laplPLAlM5jzNvMfgrdLUvxN9ymEXH
4dOvQ8MLxG3AQHAyjkEtELjP4jF1BP1EefM5wIUhET8cWR47OLmV2NAQPlw9SX5Oi/KEPyzdO5za
QtIiuBxCr/90GSEH3z5Bkz5MvBPq7W1EOu5Y+PS6yiai5B9vuGJY5KQYlPvSAVZVjDODYR409QQ7
V4PCpv0rZ5PTfFf0ZdptVYX+CXwaD5w45aOIXEv2Q/Ia8rbfHVMZzooIuBLCY3cq0hGwr57cD527
XIWko/TWwmtz2A/Pxe0AVxOxtn536mO45z6zpSZG2NeJRLHSAGDx+xHjTZEPZFR0clkdCBRq2wNd
vILIyUrkHw+bmHQrTxVyT84ofnEAm/0we7M+UYnPZ/aYMvrzZvp/YW+R+axCJjumYtnKFRVZkHw5
0MbhxLQPi7gRQFEAcZxznVpBEUuWrdObG6maw2XzmTN1rE4a5K/srs2hNntG+1pw4lb27r+xOeWj
1D7x/81Ys48HmgKWaCAHKGoGjVF3uUFuimzHKp60mOkHW/oQ5vrUV/SXksq00ZyP0du3tBViVBng
5R8PMt112etM02G+YN/Khdb4aS/G4MrnE0IX+oyOyhFxa5XL9dybRaikGgrFdvuL5Tx4rpTF8hCl
hyINWVF0ePXC/gQXoG19R72wz3vqa0rRlsY9DsPA3geNUnODpqDVEHAJX8ukwlkT9chbxwYDjHPp
JT4erqhCZmZ4QSRserds0990mTW2WgIFD1H9tw/WGvOIYTvwLM7VetdxcPHdOXtBpoR1JcAybXYI
SoUrAng2Xkc9YrO2Y7rLi/t+fZ8G1L9Wl9+MOGd1VasFSdm3yYyAD0xQZNr8FgL/AboSTuYzfP3w
NRNCHFPT2rTrv68KD011d8RYTeRQvEUVTEtZ4BjNQfKj8whYEO0fDVkLQgwOvn+YpxTnOUIl2QXB
eEK+mBimdHytks1AcFBdCwWGMJkJTKcs7+irZd3pf+WlFNPJ7YbT+vnwAf5jyj28+oDbFg+TICw0
7b77wcO0gml83++mX6fPBola5wPAis4ydclBsqMeHQOOzSx08U9DfCHlDNiKKb8G53si7WUT4ya1
cf/zPPu96VRBAKe6WIKeBfrvu4ds4l7meZLr/PwAQlnfLYACn2YfapSSppncjICZQo6NdPI5muMV
sbo11Bk/FJiraj9jn86PWoZZ0eoLa7ikTw+lqzMXOPVi/9B5vh9WX7kaoXcprdnfbXCHnBtXMRe9
CJ+PVMO1zbia6APzQdBrU2dfK0VhtVoJIHUR4XRX8HJtHkgMgCmcfGERnHiNafqqHp7AwaG+O/8q
jQ+0CRhy7bPj1yYtKJiVL9W1iI+/UbuYRcmih2YtNkF6ZXlb3QwXPyYdYY/NKhpNcOjpioIrCMYH
xmVd8jLYmW9B/eT+/2FMDgety6nfHkMt4xv70j/8TEFn3/hWrvtaD4dNAZedwtR8HhTsDMBgc8+m
7dx7OsepopDjeydSb+yogSzMrNkmx0th8yoGfCNn1n9KxQQMXWI/5V3Wn1PQhvSMuJko0ninb04k
6aPl8nTMKbrify3f5RAlcGBk3WjV0dENdvys1qsRch5yEGkasAAwwq17K6xxXL9d63qwaq+UVixa
tmsxAMwGkO0W3xmgqv7IdvANXwLcQOMU5jMCtfcbTeewCc0t2kh80bXP4mPtcbp6Sc/qLojZUUy1
fSLpuc/CcL508oZ35vv+T/G6YvIo8Fy/VO9kftEiUAjJXMJYQk01OsGPEqHktmm7bpsqQtWT1KXL
YklxV7AFJw6wDZd9xzco6j3e62ToSOtn37mkVu8yOLA42AXDRC8LxK/W37z37TGuDWjBCKa/RrhQ
D+BJlsQisQfrg8PejLFdAhMQ50CaxETgQhnONo351Ji8giOtvKPVQ9sW2qBCG7gLPwbaxZTRqFuR
cfV/+VU0YnF09SO2k5HlVtC+AYOPo9aYDGOdGyEDzicVJovo2bR9ViuNuhVeQ3HM5kECz0kiJk7z
tRYD2yqjIaYylRZrVmrjQXgonEb4dCTvm96NVSDKR7xvg345WHvUu/dJX2msWrydrRqPoKvRJbAh
l6H90Vo5wsNpY7/4K3jFjCJqaMDi1b6fmnOVHV9S5gYjz+EosEeHn4GFfrddpfsxlf6n0LX2QW1E
wPKhfbTJhZsfy4vPRuguE5Ox4DOQzxc1kPSasJfNEWoCGGEDyjyR+5qI75hoFXveRR06ZnhLEIFh
P/o549g2YjwSPnfs6eG9dYREz54ieS+NQ4wCtoQg1RD7wgJvwH9QZsA+iKPNKb8wRjXl7OrR8quK
cHIoHwjvw8+EtNW+3zwwoALNF+D/WWdkiXC+rJVGGmUjY07Zo00Be8I9fUe1VGELXGFWtatBUFzC
x7zPFwp7nrPA25BvrTV8dzOfu8LP8Uq/QGYtEOTBTJY5l3wmJaR77+8k10sYSkmQSpC2KHPGjItl
LQfdUHcHl1wkUWvWLxxT4UxPaGX4m6cU169UueDOhH6pVNnWizFJfHyHZ8yKqf3Ip53gh6E7iDM5
cmzCp1ELn1Sghslz4F/MgQF2P5TGBb+OfVVU7YOkBtaLsy0tF/2bg4pCvufprGA3y0fxI1WRYuXy
MLMIUd3yg7Kmbow37qKotTJtc2X5oH0Hj+5XUnFgdHiN8wxoGUmUWyqo7yTWcQNJbN/RLdsVBcCf
3RZ/9uZI7f92OTMmxaX1uHRjkqnzV5iAnKRtXT3biNgKWcftUfSaHbJYJLL2z4lv3I1MjefWFCdR
lQkjr0+6FyXAYtWbKzaKVhBbnkOuy762lopDBW1nZCK7NA1IabQKXDlmiYveDA4yxFFXC2XKoopH
QRuQFKvYORkA0vVi3R86MM9cVZBRO332Xjqjjt88ZESjM3rBCaxdoLc4oUlTLKqSuEGZl+QVYFw2
RMhlovHunmdRQdKt/8MnZaLHzTQxlCYmlM3z0xTuWvpsO7NPGk0U1Negx9KAHk4j/ThttcEddkoq
R/DwJhSm0eYQcJu7Xbx1/8cbmpQQ7ZO5EZ1GrrGEYlQpJE2r8uGxPm0EQFZKZMTPPTbPaFwvR/pe
ZD4WRdS2gUgxu8EUb0qZDz94jaDhCjECiHJPeG+ZpE6Ysg3pCBgxsMSnKpLesssfthGQd8+u5VKq
VFjG2a84Jxw7sXkQICG4M7PGFhoHbHIzYYN4vUjPj+fTot//YhN/jUm/vtv51ou4OmjnRuK9r3Fy
/tG/M3/5nrmGChPuMPzW95nyFAwW74wgvNeCLF+8JHXKbNyE41R0d31d/lXX4gfURTXhHESOIU59
lBOB3XbqIa4yLRdhxAt2OPXcJoH8kgmlhGV9D+WvpTs+nWqNHQir8z1P1Ws7T3mqPw3ICsP4Ihhu
r+uTELQgv8vr7R+OojMbOGCdOQhQFdiXFaeQNI7IDCvo53g+9M0KipGpFrgiBgNZbjcmfK3zeVp/
EMd59rl29SsWO3Po4jgSyJ+VNwIVzKXNaqsWtsUm1CT91Ql5L8gVW13dqdO7lqS5WGCQID//ydtL
r3+qTiXtwZ26s+m8GqBzNaE+GcoH5J3BPRguminXc65WKiSzHSzjQoNuLdlQOtVE+D8N6NS4ZlNI
KZsF+VNtJniavI/lD7XAz2250Qwjd+HcrbMrpYaC1wgVXNG6V2FP9ns5m4ycDo8qlnwSUvYHDb+W
SAWS6Qcm6AL/K50tE9kjsrwfQoS+C9wtvF5C7pKgrywSHuTmJTCPhNbk4ve7lxygjjKbHjfe7uzw
TOsOjeD5iM5Ew/vwjchd9N1ryXzctEjfOaNQbGqEX+bFv4ntlwrRDcjyDxgwfLIwphFaTTV8Z2zU
WnrzL3oeLaYtjo0XTl2fOo+9i3gjDhhPb1+rXy/afRtUZGCeP78HzhlovgsBSTXA0ARUq/816TOF
3Pk60hwq3ynZp6NqCHtl+yLBEODORMBzLVoI6eZQu4StcVKb0+xFqihfXynG1So+XYLXZDZ6Kysn
E6qJod7pyJfjk7BBZKtDiWhjm064Me/9vweaq1w7WtXzIQ9BkvV1xb3/JKLyUVcNSsOUZS9+qvqi
2bMRmN7s0XbqIrLmcD1TUh67EVORZ8trz26Q1rwVUund72bDZjpWtc2stBycPmFASO3Ioxs81Pc/
Y6Y/blyyhlQrhRpr4vWWqDfHjAretyMxdokz/8Di7cWZvIhZhEUBKNaYrQ1ItvyYpKldH1JQLxjw
ydiw7idoC9Dy30pwWlqSUFlBkX4q7QZpMKay/2JYJ3fLXQwvt8adEhB5gv/4ny0nLdl8NgcmGYtZ
RyFf8hEAEV0IBVj6Smgk/TvlxDedmEsmsvfO24OxQ8WEqLyLxsR8hr6CDW2ylAcUUP7bfBop+SVo
f0NZatblAx5AKF0ASFil0zJ9LHHDMIp3kD6XEN5CeGkwujSSziElBI/L4D+18eKoLU7V8po4hzbr
NG2iY0ypxVyvBgKso4BXleFcleaGhEbWXRq7YY11gedpegZeInh6ulLZ9goq7DW+qR1VpQsq7fth
OHdxhDLBy+/MCBye5T+V54XfcmJR6rtCalcBen7jzt4XF6bsHWnIRBXUbIuEnrLoE8VZeljuWV/D
Ln9c2pJpWstOrT1XzhYj380GogvlHW+rGg9DuKrWW3ZEmwiBonHU47pEJNtUPZm50xCB5AJ3k01N
+J0qlqm6UUBv3X1y9aZpZ53fHs471ZHd8xo+RCEJfYXgRZaPLt+tRKMMIrVyhfdaLBQZ73t/huzD
GCnaF5SdZ1dpe6UhMrFzYGFQtubfHTIT7fXJu/9eYH+ufpd2HK2GFulPhBoX+YSMqoYNz5YvoTWi
27uPjP4jh+ObAEr9bX1MfQs1UFg9nog4m+kFzqyLBNdvcGQ2SRyLJx3IFXsLt4ZmeMDcvHpnTvTG
Iue1AMNtQcJulkhXn+Kn4tv4j/gKX80ogbisDQkZz9zsGaT1xnNAXCmqqHeQ8h1O2p9RmyDn/H3a
L2tQHYlYvaxsjrDRsuaTR7FJJTcizjQm88VD4gZ3kX83ko3hcdPeZA6tunbjSKVR4pXn/x4/HmZA
kXv2otReTSBg3W6dabq4+hWUF0aSZjMI82A65b2T5nkS1Dn3FO1+ZJjgCpReXSpwxv7mtYeSk2f8
JumLwq74YzTarxRLauKS5mdsjWTn4PQUIDa1KjPffFaxouFFnLKPcYeN33hOEFVOwOzdaw4NN94n
+JwuXHrX/EuupMt46n830xeV7Y+RhYI5ZLdctPx6xVlpWjmpWHfDkenSvW2dSjWQrEhwNLLKNfny
aJWK9J0UH2WfT+kaw3vmCto6AXAwQTV/a7cvaWRv8+3gprCnTbSGpPQB1kMy6t2x85EamzFRfOd/
lNUvrAa3yccABbmFgcTn1lyToIiaQ+RhW3mPW7r+qXSk2ubSbXCNyL1ipRYgKxGCK0m1e6bQFnjd
DvM7uyTeVxvKYRT+m91uiz6oAXAsD7sJsy4X0sIMofBjcgjZj4Kd5OyWbOottHQj1TS1qmHpXNdb
Xp2aMCKorCZ+Jncstcx8Hw/AXLJeicV0NOkRIXgKr8s8IopCUbBOSKZTH0PTbAMm7g2eK6Go/XN5
OH9gGh4G6IXL4POci5MKtvOFPLsauBDZL2HKvutFIr1Zct5yFMucgMWPRq5cJBqBkPPBHdbQSu7f
07OqkZPFCi6ipYH7LiZgSUNCoiQcyhvMe8JAhspPW1Yw1/IBQXdXGtWReWc8xo3OevAcGOIZjtRq
bhQBk8sH9gqevnQ7Odc/FyUP2Q+lFEVRQHTVdUrRzfCUo8of07KqS933kMt9njHqTgqFPS9mMJxO
qkyyUJWhi1kJG2wZhLFVTNNCvfKhnN7TUGBYPQLUYJYBjKiyCjfEi0zlSg0XY8urrbXbhFLjwkGS
+Bm1o/FyC21RNrKK2fMYG++E8Li7BhGAzzOCQfY0CtiRdjNZcOF6CmC4DvbtkTzMqHuHxkN0TEbO
izdDXSAT2E86af9okMUEE9UEV9juW7JJLP9aq3L5wOIgD6DCNdCIzw3eYIE1tUHqcHL+vv5M2Ayz
KqFMeOMc8xPfIFgYE7kQAJM2KIuwyZWbIAWF/njSK372F/U1otnJfmT3poa/++ZkXbjb5EHSrjug
+T0/DdUK/el2JFSHM90F1Pm79FKngDM+GFcZTRaTSI++QJkhEVn6vmpR7T3J3fJjYLyjWv6Fp4YP
Y5Z4+kq2pKd1S8Ub2C9wKvy2Bx7asNqoj0BxfP0CzaGYhKLlCsAgd/BfA4rXF96y65iLC2xgXff9
MsPnBh09awz93MX0mwCnt3sMn/tGAb78XZROl/I7eP6hpeABLNyQoYSqV8RhviBICbMEV3Tnj+zv
jQ2YCpi4b5B+Cd3W71cWRtTStTDWE3cU3jSdteEY2OwPoUPrkI4G3HboSJPCrmQ8l/aBZZPGnDIe
mvllnldMOCgh+Cr1oKoO3lsyU1cXHJUz9TpXlBFTBdEfTPT2APgqjJjghVx8gi2V3s+BJwTCMTyx
jYwxWJU1BQzC/D/TyNrKjFScbg0U4U7l8nfmFiS2HjkNrLRVTh5N6bQNHnK03RBZgXt4h/XD5AIF
4YbUOpnj4ty3C3nqQlwS4hJP89lp2G9XDv05Rm1MBaI7fl5ETJMZbbt5bCLl6TfFsQ2oJCG13r3e
QzTUyrPGPMPWfW6CjcbNwClEQ4L2qu4/E153IVbLi3jgyh1c7/9B+4ANd0CSpW+y1yDrNjOiI2qB
QF2GULusk5olYWLz9J1W0r/97nl1+1QC3N+2EdlGYWsLlJUD7JFl3gdwP5iczzzJR7u9YJOvLJzQ
tQZF5w2O2wKOIEEbzzfeBLU4zhK73SEotiGPGSxHfMdO3SjNrBK2f7rwrcfQSzuNK9c3V4S2Xz7Z
T2RAGHvZlvfhbR0KYDRrYULibkd1I9QQrW6p469v8mLDBpn4w2hiiZq6lpOhCDeHLqh6AkaYKukN
I5AZkYvjA2Egt6P9p6dVqFsAjuATC4gVdBSBV2lpCoaPR9dH+116z35JRuZlBc3LdT09z+btkT+d
E2G6ggrYzdp90mDo8Yc8KkcwIPdlIl6tvWRN0kFjADvfGzSVMAU1MG5JVgWj2WkxNfKPU/wdYtIf
qgKtDKnBm4PacCifEE/BHjXgJarz6BSeZQnIWPE2MFolulYPpiqslBMt5ZkDeSNDNwfC+YxBnaxs
H97U85imXWJQUJfWHY0DIFghDFPGimyl8XjfRL2EuznTwmi9uOK1ZUXBzpLmTGQmgTk2Lv2pMlFy
iO2wEK/On1k3ilvATGbp0PCylDJma0CbAcKVEbz5C8sFLsKLw7iG7HvXKAIDBZhekwqox8oHvX3n
P76xCA69PRXvfXTNjdPvhHPxTqg0M9bRX32lAFQz2syfA1shXpAgrRzwJG1lp1vWVfwlgigxjvkD
pXujfn5hI3qrabzJX+hwEyYPHpPMELWMArq+ehhJTnWGu7fs9RqweOyDPkv0VI0Gaedyqz0ZtNrj
hl48hXY5CGkzvyHYdxdC902braSS+sru7vqY9lr3wHVK5XqpzXVpWK/3oKl+1Oxxc+L63WBYXPW3
J4hrC5Ek3VtXhZm1b3Kw/jf/Q0YloPxY93e4edgUjpIpSPR6hA0CDhbx0d+6I/fa/qjSL9fxCgBh
/w0ZLVOGHg1WqHvZFZKSHyPVQ8sfcaZSF/hNJBqHxFAO5EKgCNMbeF3Mtp9g+iaE6DnKxEEVjglh
uK9Nz3cuHW58jTO4vPWTwA8zA40HvZXvZ3L7zVRf7R+Y3DF8mb+lLipgQrDYkrA4qOtnD1ENnPHW
q48WDH9TEnvEueo7jxpXWop4pPb69YHuSFMygF3AfwHAeCHjdsgaUzI7a3NmfwPVFbgoWd4OpukI
b2WyoIDDg3FYX2TzMyK9Dm0HKkua83ASgiDXy7xVHgHv4bAUAlhEE3LJ5dixR14NS/dVGk8+Dr1b
oj0+jtRyzVielhMul4DzwGEc5BwkYiFNzB/72NvdoXVS+YpD0sOvZ0ketMIuy4bAg4wqCmowrLNz
KJiBbXTj5D2bxiemVTVkK/UlPIETB33a72LM9TWlUBaWS1DY3tNbKgXgxp9jf/Iqh0qobN+zdtqN
ZXT5OeiWJ49oU1sma/s/Z95QGT5JDy0hTpAW8dyiJpOSdE7q/fc/dRs4NFB3Uxcb4wCa8cq8Gix3
wg2t9xRnZEjGFyfKu/OZBTP5jjtmnLS8nj9XaZPSuWYxZgUuSLt6IaWlgbI15TJ/aSUxtEs6ZZd9
qEbKmJEItui7fUzYafqB5xLkZo2ZE1zXjD50mcYCrQWJzMm/QFu2FFYVwQJ8NnP5EYWF4Kedgd7p
+AgigMrv7QAkhSumOsPU/uAODsDMH1g/6YmyJSc13I1lreyEhFmPIL7+xArZj4cJWT8MXlQWmuFz
/u6Dgu+1PBnH5UzS7ZEPQ5f5udRSRLtETK/9PYT3urUL4sY1wH+UAWJBKv31pRH5/yDglXzSMpa0
A+CGapntgOyog2YK+joDDiWjYkE8p9eQepHkiOJQFCrXtlja2W+5s0eDLbkPPW+9RcyItoB73yKd
31oDmVCHMhx1H99nNQCpY6M6b+jBZ86Xf7htJIB/L/+mnugwwW7RsYOMKK/xvjoMV8nI7Epwr2Cc
V0oxzR10ixKLpZU+rN6SGtmRP4l3nAnLLZcEsLKKNMJe3c985DMh9VfpV6fEUbvsWf2zu8WJAcFf
Rr8MEnM8l+dW6b47WO0v7Oa6PpIbVhIvLYxvAK4Gm+3yyQ4TDq37sVZdozozKLmMj6H9Iv6yK+JB
ICtEvJAA4YPoHze642gG6LgoW3mqVlZWcP+7ltzIZadGcQUaEMHrxNgsDk3zIq6WHM/mQ5JXaTJa
B0flyLqtyNQkix8Md1irFs5WdSQkIxgDfy0g9Vcs7b2E1FfLRFrm+mmSzolGqmg+7XFJNBqMf3Yt
RfEXoFeHe6abaTeA8Eca70eUcBnlqMdgF/JUXYxhWP8bVxuEMla0bwaDFDpP/NKnn2i58Ns8kWgY
DvNke9dB+yzsQ6IymzyUuw/0I5UW8r4bcALssFBz8Wfm4I1dxNXSctlpDqWt0Vfy7FTcjZU4Tm8D
nrP+Ek20IOYTlL5YWCZd5yLgszeHKyVxvC19WNBaGyjZWdyg6pEyrkaVqWMxYt+fP96ESzMMG9Oh
EB/j0rRSVoOhtbH422PIPDlN1AUJdshv+3cgwoe+VUwDfUyO2N+fSxwnXvERhvx0ezbPxfvbLblR
KfuQiHwXdLMJEemjkI3myktqsZkcKJ2vEYKi6wS9SHiQO/5BQk7bWXju8EIQYxv8USwjGl3m+DUc
yQqVMUMHNviCQdu2HAqN+6XWUZ3yS5yVfdK59v4HVIy6nU+L1JBAC8EeLjoET7XfFvKshIBD4COW
a1rXpz98b0Z5oON2egViJL1Vxluqk6nadM2JYLLgqxWMjPGk8ViivTeAWmLFgyEvIgX80dm8iQTS
1f2/U9D9QLNEDesXyAXNNIKE0kFq0GBY4thM5KC9aeikOZ4/OxPImet41XZDP7i/1BZ6tDx9CZcG
CS3wFenCGfhjzyXIN1xubfyAhvHxepLGmnIhBd7f5EoCNpogZ7Olby5TgiiKDTLZGc2NMhiCGlqh
x2MRvN3Lmli5e/0nKFbDvksh9GK/8Dhq5g1JBdlKnNgQJzexAlfokG30lgn8HORXTJPCfFR9hmul
2+9PLgWdU2t9v8VKKdDBSS41wskQ1H2ZIevFTQ49Zd9MUw22fLAGNRdhIsKe24jmrhDIvjWZ+S12
AcREsDh6VSPDYwsLFYcKcFs9wpt3oiT4Ih24BiotJDlHzH8gPwEyZ0BNCSrmfVlIplqXhUSEKhPn
FvL/5ue8L7Bux6VazCuDIHHqQOPuhzb8SBmxoGS8+i58FE41vPE0lmYkNKhLDljlTGaMRP7VBy51
OxxturRP3GlFxSfOKOwaHTRPBKGu4YbQyl/jYr5IUujjTWNPodsW3Pum+uLCLvFiXQiQCqNLEg7b
BUpBV2mNp52stEM56JaKs0OxRxOA1dCVlARcV25eS+nvciFl/PU5JpYjdxiO7jUmIRVcxkBGNCHD
aCHb687nmp3pUiJCq7el01unYJaDy5MCZtYQ6idsIYLZxwC7T5kFRPviYHJifdysJgQSlGqGsyOA
hIw4jE9rmzYhnmSJzq4WdCuwBsl36NrePSzjBAsujGgHehrpp5RE5Fl4adb9R8BLqpasPBHjuoqH
7dGpBS+S+wIUCn+vh0BjI5Cnyt40XGRMy42xdGiph9lg5WLmHTTimE5rbWaKCAxa4qWpqjoe1HHC
wtT/8EvBnFZJ5tc4w5jld2Ku6Ai1ZrZ30kguBCp3KgMRRU5Tnuq6WyhBg8sC8gnu6NhtsGdoIrZm
4aavjpUDCS9WqMPpyv9dV+fuEm//DY9Hx8Yhh7rjDdgK61UcT0pbWKxLa7SwrKv3WCq+BLwQm0yE
DwNYLe6b2y2v+XSZis5IP/NQTp/d3s7U/4rp60F7CQ+J/R2b38Q/aClJiwVnF9oy4fOJVtnPTYNz
ne3L6m25s4FMb/ZVKNTNtgIpwZjaB9YF6NKBoaE1yNmtcwqX8QHks/vlSY819AfSDeGPX1kVe2Jk
SZEPaRnKa+a3h9AHLiF/YrEFk70lOwSHGb/2Qag6dM7y+r4S8Ga3fzAJgeybuAkLie/y7BL2Q10N
ZDbK2wUrD/5STflp/reN6cXIAxMxSZ7fIq+KjRDueUPBPlDThlEQASznAWdYsJ3znFD6RuQsSSGT
/FwUbOC8AyiLABlS83ogdv/ptfTHLaSlL25lMagzDE5Jq6T6wUUx/Fke8plBWLI7drsuWidxzKGI
cPftFsHq5mOd8i5diK40mJ4Vr/85y5YJNTQg4Hx195RWf6dV2kwzhxaMoUikFuhmr+qyy6k03Fgx
KH0q5ZavaLostHoDrV8CCCNKFiSCnCdpUwoPpFcPZx1TNQc1dWHge0SeYAqMCV+l5UlxjStJq499
1lWL+RBt1YtNQyHxUggHhdIhb9JacK8hxguww1yKYjaJDTcWP8HW2dUKHmVEon69QHIOvLrneshx
QD4VSmSPTZz1RBzONuaoayyvnaNm7tcjCTy5Icg5Hflmof4TiV7TcjVpcqslqXehvcDixvxBdwo9
wv3FL3YsMqDRuLCfcoSDxwau4cw1k+Sdczx1u7NxmNeMT37pDl8sDSIeu2pk2rTsHYBoQouZJmMt
o0m7skkitlywNm9ny5vhyg/emG4rNSs+4GNFrSnsorRLve9uMsLkEBeO8CHpMAAlENpMBFeh/MKW
h8GN2AqLQr7RnwQi/v0mHtdurPvbgM1jjUEzSKUnfqZSqMp3bKIDkhfY8LSn1KX30ivp/owep2Yb
Su5qt3xxHFg+35aevON+KyTdnz87/J7Umjt/OYp2quVPSxhXubM3RzucOgM1US0JzrQR4LdOvLUS
imGFGsHnPAhDx9ohcLaN0mblBdUqZSszahaH294qiL45WBX7Nv6TKSO7RtOW62x/Kyh1mPhLm5eZ
GZQcpid7n+Tl+FXrIfzKZ8ggZ5jHSXIG6UxtpMydseI7q4ZbAt087QVh/jmfQomnuWBQ56V6VX5H
W4cXYR5pJFRw1RQ4aMKZNUBEJNIK0c4/flrH79k0FeGa1bS3gCtyU00gO3bzEqf9aLXN+cOELT8s
G+tIx10rPcduG4wsL+X7txHmjR8FTFLGtgwEkNmODm3NRfSpEBLbE7ijkHXGwVjfn4yDAMwwBlmD
C2WU0LonqxbknaVp+FHqeg7bVAmQ6Myxt992GD9kbkv0vkrwaPk0H0RV+GKmtzXnTMRZh5zj5HFw
PZzGKf7yLpSRMx9ZMTNYBH+Rxc1yQDXV0ADzg7eH+O9his1IPnEuOrLLXnKiNM9tj8QpuQ7ixKU+
/fVWIAvSzSQMWMejES2xeUNKRGLsZlGT/9o1TIbJ/A3mGFbPKCdrV9l44PxZMqq2e4xaQT1JAO4U
26arkIBSLCGFctbkKBBvyDZQMR/2Qb7DyAEvG3GWhLEeD4mZPnrrFWd1KkBaE9/HZEu1F7uGiv0d
TgaEGPvid99eeHBgAcgf2IWHMWECHvj9AXN4zcyYUmgnFCEbwF/Nkc++g/CS1Fhddid7P6j1gmoa
jT6qqVHHvfAbatKqqzECehAaGADi2Bw2JUThd86RP01viThIavpEuO4QdZd9R9bNxsHug73sJJcc
K7ruAXVNOOpjzdJ7iD9H/2apU4lUGYohroNWrxJcJMcXC5qOAL/YgnyfPrKR2NIGheXzJa3xxHzL
TK+ZAAPCY+KFeqMgHTsgBlOvgI1RBOASaT647v5L6QoGRQTJipqPP3f9KlqmY6kiQcsvDSX7FujG
xA+z3yTUmLAyZ2rCMR1tEy7L77bLY98Ty8p+dCwTn+i1lCZp7cBQQ7XE/RKqIoiOU1GasFux+UTX
y69I/0uZO7I+ek9OnCzy6PksrqzvW9Reil7qnjapZOhZJX/IhxTxd18GVlsIui3hrHwPJ7wWT6ms
/s914LFGzqdqaT6x+bebBXj97Csd6dmrUj+VT/frlqZrc37o/lFnvo6Q1veY6GuqntbfQ5VT8Ygq
4Imng0RRZnoHjkTyqfELWGDAcdYUTGYWEMVfmIG4sTbX5HG9EJXeUDHI0rRtdJqbhjdqJAtIX6WC
IC8811PceFlPmn9vBwa4wQGRsn+CoIEHlGP5pQCguY5+lr+VDMb+A90yusy1wh+vxmxUdiGpxRjB
1iEwTB5+5xkl1+SvLKnUsI/CcV0RvRjESvZuggDlWn2TQbsZgcGN9e9OmZuLOHRWV5LQ8mQxV5Co
Qw3YjGbYBUoPBRnQHNiPvVReJzv8Ebz9T8QXi5Mn0WvQwvNdF9Z4Ao0A3H9GF9XBxNUZiYS0Dfyw
/MpcggC5TNfmvL4cCWNAmOZSb00ghTmAzxxGW8ldcNNkVtaeQeNLEQzB60c0ae5EZ8GnWlZ+rfNi
Ml4Wc5BRuNxPOYCVbKUS7Yl+gdMxSk6xqo83i3b6Seo075Oz120TsF40k2FBmWQSwmWEzldAXGtI
D3QdD0vS3p4SbvLxHw/ZNtD77IWPhHNFwWjBK26lUm8C+tEgikl3DaxSqmOCw4f7VioOPSc8Mnz7
Jyxux+AMJdtiBOhuIBwqQl/qhhCeqgSeP6lxLjLJmBzJ47uuNcfSP65IZuPeXhp7htk4gWiR0kmr
Z0ssNHqvpxXq5cbZj2xy7/Q4c/RxrM4u3F27HIIFknCWSSx05YeUUeAZi+y6AXXCwL402tJt8+xX
bWQHM/vndvxq4B/38jGpdBKcd4LxBaX7lDj3fciOOBwDY8T4es7QJQXeXWaMWt4Ttke9OKJp69va
GPtDZ0sNZV+oMfqn7focYeT0u2UPDvaJdkA2x7Z5fXyYSZyzG5tKcWt5TNdOZXXfinAOvJH3s1da
WhKR4PkBNPLrgWIrkZ0kT79ST2zw2IolGxppLQZY882AaBedkzO5jV9NsbeInlU1w6nut3C8awKV
PSb7Vnxx5NKNQTWxhFJvrNLOoclp9ec6ux6QiwdfhdmtekMAYH0K2+wfi1zQ2Xc1uZWWt/oYc7Ad
gKHJXVc4gZCqsEoy3PhWcp6cd2hmGFPmqQ4P/AlLeecPkPKgQLDZdk2ybNvtt0FD6rmJRL2nL+MO
vTyFECuKP55mUVDOE2PIMqWiQZwUJ2qJ7Xi6HK42kPyUXFJDWDcH/gVaeA1KXx22l+ERm3m6kxQG
zfT25DKJKKGx74HRLeYkbQdzG+Q1+1mLXESwDFErgPtUE9+RrREa0aPFVgvfRmqVYrHSZmI3fDLo
VIyrqjUg4kr8sMs2706AYrf+YocFJrKzVo0FM7+6f3TGIom3GdbJ5FsK+yXzKK8TYBJPfGKyJzXq
k6XtQ+6qlvdpylxq+cQtrs2z7tiAc/bK3KPCktEgEXfDuKvA9hiat1ItrN7BNBDdBYKIX7g6Y6zb
4ZoqHnuApY+YjKbtZzcKBB583wCNhQcLEQ71Xv9tfViUS9F7lCJmtF+apC+JDHO1BuaIykmhZv0T
kgYLqikKlCSnJifunOGf100UrquawZ/+OL2MRGGGiZmI4bDcfkICbEngAq6wphKyoWVFdndNI8+P
1POb4iqsqKtM9hzxb3DRfzER19uba0gRFDrGze4H4IgoyxkghNnSClTAy40N+RvdY+yCxozF9wj7
HfBZqX0RzlXXE78gUNiK24VvEV4HRCnOjnxhbsI4/8hA5dayxD7W/rbJRmU2KwNwCiHuI2BzXY8K
g58hjOSlfIINs2P1VlcALFtQSnBNtVSZOW4GHDwWEinaB5vaCn14zx7h1nr5Nae0ejhC2UCHNXM0
1eBud88pS2cqMEdAbh1QkUuOmVP+eIc+rNI9ssR0FvI2OoAKTjPGIY/yrgkGdMZYSRaeGGYFBvJq
1MMTrbQJIi9E/dpb0sJfwcTkwtOXuPZtwDPwzkLGwkLyeULUd6Q2QbCkx1SkQyhe+NEHtfdqzNLP
Uwti21bHVDuqAflZ/T2/iVNA35OihxX74GfQ/u8Z3qlqvvDpJ7lrShBd3SWGEj+WaWO5TjM+smr9
yt/1pQNfMiwdFFtgQpbVMwnQCy2VjQ7yh2gZ01dzR2hs5YMlj9cWAuYyfFtDT+GWpp+S/jgDBJMS
t4XCpZcbeSAm4hfzrBjCxuczXdGGntn0Kcaw1M/ZmlR1YtVgRfL8mOa/pBcQS+U/gIzC7BV3dZts
Ie6H2PRlGdNmK94I4kP+gPz3gBkp1U5Gj3eSZPnqew1cW1f4xFP8Zc2ATh9vpFVYbBw3ImlOHdn4
VxmRcCqOwyxkizLi/iIq7tgws9uZ7fo28KrEKLfgq4sCN1Lu5SdERNfDVwPx91SEFjOOzvLRjtjZ
w8aeD8DRAfKkNwNhvnK8c6DchaXUg4EXEfUue2gadnpwnYSaMLa9mJPWfIPzByekaVTEKK8ozLxc
M3N+CutxZINl72ywx80eVax8HthPgFkJud/wXoOZkHpEYIyIu0zxpYhfMOZeO3RoB9C6d1i9/mJP
sTvB6IDTX3S/JgNG71OkM4arKugfORJ8eKXPFJp+IUkptQfzuX/3Se8IzCsqBT18o4WIKwERQVDz
Ze0E/efuRU/N8a9n89Dm/5XXNaUiyCbSJ3LE3llY8xbfdS1ao4tyBl9vhflsev6IieuHM5K/+BEc
OJkw9rI7WfY5W38o24fWSTPSgfwgai1DsdzlxhHhYTkydejUv4rWCVQ9Z9m/kW7PPefHMd4+WisQ
iu2PxzbiuB3VkpI6LolpDSs9Grvrg7pM8zZSWNVgo6AnQl6PRVs+wCjttbRTg8ybSi570xxGYd6C
PL5xbMx0kiQZMMyfCBYyxJwkyj91ZfUX7ftONotdaisfb53y3bq2jQwwB+hNKkn6baaXcfJRQiRE
TxF+3Cho/p+tqI9C7iJ9JZm3ZI4SXgUJVHHpYO4krR1hUqp8PY+2bF72A8mWMKMkIuTVMrJxW+It
yc2ouSRzVvBkqfhiNkn19Vj7XUOeEE6MTkZeIYNL8MeE7C+NDR3gND+5c2hkAh2rze0oi1UTVHm+
C0TcaSdJXKqsgQTAgPkoHuf2VruOoNJiV9f5OprJXrd1eoeZtRMPqUBsbpFknwzBs13tt6zNDoTa
UB391xUF8HWG4/6ptzuUUZY+hAxzvMgUct+r82pIBvhByDJMFgEL/sXdHcsSVEsJEke76miUQOJ8
CQmzial0AHMPXF6eGHECp5B6hxYUqJivvzlc0juF2vyPnteV8kqxRI0Zf1RxYD9BXULRoIlLmZj8
aKB3f6x4T8Q2/bkSUiQNmvbfY15LK5qGKsuE3LkHCB+UFD2ph5tZ8bXOXXK8HRXSrgi8d+BrAQ7M
KZyiwDOQyP6GcsSZAF3ngTs6yaIwbgz2rxhjb64cXwjbTravxQcz2GjGxpPXJzFihRfsdCDha5qV
56XY+HkCF2H0SqkoXlCYaBWAUt+kN74417dTQS6q5lTf3teWjX0l28KxKX/DMXRQCarkt7A+04Rq
6epHFEJfIZ5awsg7Ctjou33k40uurbe6o1UA5q1AUtUnu817/aCAr/vrl4VtlsMqd1b40Xv0euyc
hbde+Nb6s1Iu+bdWTS8uyA1m4RSmqHaDX+WJo2usdsKnPZsPpvsJ/mHeRzc1A9tVv7+W6VL2koFh
/cg5jcRCRwgRSEkWMoFuNq0bcgXl2gKe1UaexZmlav+DRY0Q/udUNViWnMZmkx2ioALeP6EBgXbd
q3azYWQogVFYfpsf/5Mwt+oRsnChfbdiU0U15QeaySHbyMUdPqdEmZewlI4vv2JjnFdzbLGt4ICF
S+iLQnr6OKTVE1qyKHNgiQLEEwRYFCUvY9Fq15NOA5W9bM8Fn1ddqnU5+WwnOZ1tTUooNtocBt8F
F84bKJdqG6UC6G8MqZclvY1qZKZ5T0+IJ8XBuXnLiYJo+c9+PaYGPAbIsvVVBLy4+xrpuUA5tAW9
AqGGhneDp0MbAAtonk1F/RTcUV1pdWNYNYNJLS46ArYq1w9n1FlkeZH/saXW/eLs2Pdze0VBA+Fx
kp5eTU4TmO+POeNB3VhRFkn8yaVCjBfAeSeLhSxLVmIOpSmN2UdhVfS4OJ05e5TT+fZ9X+0Wb4F2
XvvnvizwV8DA6ajSabVMABplgICfH8fsY0Bs75FprpAAdXR/6Y5RJUdQaxSbO6THnS6cyso0lvCq
c0mBY4m9N+q9w4KWfSWXLqXqJJHUMYh82aQjSQ3IYqFvAvO4tdBN4QDzqS8qshCHTHNGpIp1r/JH
Cd9GMbOj17Ohm/LIHo2dKkmtYverSjS4CDVL11qhyH07QYtYF6GurQ9SIgIcWBOMaHuaqOcbcajE
RKJozZlOPSyDLtbXfbkcjM+rmHuv3Q2jsUOuMmraTjUbtIDuREsZs6qmgqqcIIVJ+/xHnE8npsBT
q5ex3YfVgGQrunUApMhuKH2iGpg78rJPahoG+orpFeGR3YDRo+8eL8Hc2lOoZjCW2D2/x1dxHGgt
FRvphrlIo94YEwhvTiHQgWxukiORy1DymPMy6tsmuAJ4SXFQLmpJMEXsEt0ouUDgmh7FFB5hvC2r
MtIKf8pfFrRzItRtF12N/q8MUdLdGbyXKDtVeVzG/n9ozGj2FSqw7RM4ov8+YQ0aAl0BOySQwvP8
DHpvcKqWvx7bqNwkcMoJHzJjd/kdDyZEK6skipTD1+v5KZ91VY5tKyT474vIY0uN+JzBee0DHHyT
f1IERP7gjSK6BgFN+wBuciEQt3BXHIwLADslJLE5Oe+xdCwFf7G4sxFhDNKf2AHFP4GoApGhfa58
7JIOIBozRIBjj2ilJnApnKcTAGTVnPtqy9KJuLUaTzi2DUK1j89quDcC1iK3bHohHrDvd0HhO6Ho
4qBqdnjS0hfx6Lbuf/QxwecRbCBqVY8pJOlbDFk1ZnAX4duxZAqgM0DXhIZhrPZTA7yyw6blhTCT
09ePguXwi48x3C8z60fay9gdTGkFOqteF4CvcHNTOtCT8h5ALFht4X9ibR6PZv4nZd8X/MWNHcan
UhhkOAni/98TvotYiwfv6Zw54P60k8gwdx5Sg8f02FU8Z8OswVQsHq+TlaHFVOpmYPN1tl2EX6ef
CyJKlca6jU9p3NY9gsJcFXaXlM9fvX+z3uRr1YyTHu+5OPAkImeXgkNJRfOjo2hc70hMYn0kGZUp
wEWonZHwb6lRPztXSjRvWTS+x0RWqswFiYiVbsPQ8u/+4RxA7Umy/ZJJtuMhn1XFEGW+v69lb+p8
JJt1aQBkRWYBSJUeJ+yAO5r7oLv08xwrPFlGy1sYXUE7OepXP6FKXQRkj9seGjObaZF15GjApWH0
qlpg5UaLUWx7CGzqP4lkRr6kCldYZm7kZP/QW7sTYt9RQzP1DFzTV0YoMltMIo9FppUroSyWxDtQ
8/IqguqTEAp95kDckk6N6I+7M/mJcjmCprcdXYvAcH5l8HD8Ww+95VrVkPPIHMSV2SYftj2ddagt
cQqvK02T2Fxh5+N0GysJTnrP3mnvDA7FCEtebfL2LmHrrtSWR3CJqTbfDxJSs+1M66MEAuRxuNJK
GbcGJXfPnZEHr0HodBNm4l0gyHU2n3RIvWPXzVBGaCg114iA1b3Cpf8pllw2UKzbCMFGp3bY0HbJ
11AsOSyiksUuSiVEJkVbT4lpL/UYl4RMZaBc9RJHbg6vTf7JYE57CmEQPIXioCoRQ+zw3Ub311Ay
sd/Uv/fhtaEL3qZ56kIOpVyNJ5Cc2JsPrvQ7w9qNz7JSzpZOzaLmi/WeiOnzeyq5yNiLOcer/8Il
Lcl72xil7eLB5w2oXEhEz9a9RgZMqgOFAQWkt7HJj55fInRIO5cE3wBq1/X9LfFgtg0XZ0cz5Btw
ulGw+goQcd4FXhlQkGGf6ct9orOZMCaaOni+ea4e4Y9FVNlU82dL7yRoMpOsBJ9HWSo0iVV/YX/o
F9M+stob721z57xGm+Ofk0mcR6vAdEYyjr1/Pc6thGra+wWldWcHU/ZdhZtAJlDSR3n16cxdgZp2
eumVWKbCwwMPc5tRDCYqauykxGiSCraPrN1pR97Sru2158hnDoA2JhbYCZavmYzFqf+fGfYRG0Ud
qkC8+Z9f+zcQbBT5Mafb+rtpSIlHRQ6LsrC0YuaiidQISTBn8nCi6kylpcD9gnkXm1FefwFHAhHh
w+roeqdBSmpAUXmBvjxsVgh1UI8cGEAlfe7MqclKUSTPRgPj0qjJJhYBQQtH9u9TTehFdqHlReqO
tXurSuTzgFR+kaBxIrR1WgNDq7gzyicodTcxDob2eqyccHbsNGr3E4BuQAI3DbUiQzxxeZeVWXpX
I5oVTjnjBQQo9yTuUMlKsVC2muMzHVkWn7xOuVMrSgBja7uC/uKixELqcSBeCH+PeskTLVz/cn0h
csf4CSxNYjwPh3cgvSCnopl7q9aICLFWVh8KlCdYEuH/H2JtDTJJYf9XZvjJil1V//7FoMk9D5Ez
kJYzmfBnJkbQtQetIO6oKVMKH4XBO4rQtDbo0+dKGSEOmldY3EQk2uqFIy0qzgJDve5SYAXUl23I
reXZL5BPjgHAUnv2fMI5b7fcGpzuLqHvngifwPDgZ1OfgrX7DcDqygztilEs2rSFqXCYs8fK47LE
OEXA0jnQe8v31mVpO849ZxF+mOXlqmNLkEzJdR4VTGkaxoN5u+nFSuQeAS3Z3fqHHGP6OGkE3i7E
qldzYuRTTI4KFXpEi9QJZ6sLl5UiDJgqp+TiHy1SAq0WwqWDfVIIqcFsuynni1WfimWeIYK/IfdE
TlEjU8bApQQkBlt4oUdu4h0P9OBxphTgArytDOyqFcYxuSPDbb4JxA03aCLHd3A3qdkhQCYmbCve
q3UL9zS3woUSW0ioWZA/U3luCNvOI77dBL5XruXO+V9EAXc8HcrMGS1ivqz1CwIhYFHJbRtnP+/V
Aa8KNylEV91t3WZJs898Bj0j8y7PLyQBtiGuaZNbfrTaQRtcZskXRugb0OF1/OT4HHzRxt1Mdsek
RO1UaXcJ5WmLix8buCkEFpruDZebznyorjKrKxsHMfHCVQfDVbdLkPPVR1+TZL6gXwg/W91L0NiE
nqXHor5LmyOk9xrbnfbQyXzvTgtzhbjEURVdmbMJLaiTl5V1QmAn0kFb6culDGLgTIwjj3voqIyN
ji3ZEhTzsmIsF2Ld13QDUZ97b2W+w3vadsoIzB41Zn+oq9ZV1tHWVVXiyjBQZw1PWf49J75lWhfB
4WyiAbCaDrR+eEy5Hm1NCgRJocrQHZDo6AKUgVjN3H8nPdbZB1tKFIGSCceTM41XhW9+DMx7Th1C
0EbtfjD1wnvyYPGK90WBKN/6rygimkzee2iORFJnttbvEndtjEojLu/rbpI1hCQUEV61T7k2Nd3m
YXr5lGKdQcPt/7DMtWhn5/sW30K7iLpXE7z22vNiB9mu5pDjipC9BiGToGJU7+H3qsd07DuLfSFD
l+sDgUjHnlJVCf6dZp+RYj0I0uGaHU7obl0W6ik35KIaTn026p+wL1EGW0pz3OfI65G7o1r0mwau
ZtiimW65GxgtgGT3MQXWslMKPAX5ic+B/IGLLMDqBzUzYZoz2Lw7cVajh03OA0hIALpqVASeN1rT
B7PwuGavaHgCEuG70wqjgUQ12295fVx9Y7BHuim7DtQt7Y/00z9v5vetETlibBOvi9WIERUHIvuE
hw5LL5Fg81fRZXvMbIEOBK1PNdeuUvh7GeJHe+WK6KCc+Y+fBeh1VdhIGHC5euJAVB1En0aSzB3H
ttL5/76b7ZCRWt8nsnatGYleikw6NGrnZR4Zf3Y+wI51yiUZsps6YQqNpIAK/Hsj56EgCFmAW5FW
Z+MZgHor4B7kgolDqk6ZT/KWxLZEDfJrA967ulT/J/1OxrwOM/bJj+BGc4Q70me7jpMJlWgubYKd
4BXshmlOEItlzKI0svwR5pn4z8RurTxNsaomAxHeAI7w/Dd89znGdnXjITr1Q5WXYGDS5NN41itl
37PAyNvshnLauAOLyET2JLqQt6lbi3K27nLLZHlLauXtov+pL1Tx+HOQ5+CWToYLo4/bCfI8w3zx
LDduHYx2Etj0LK3wsmWyuYQ8jv/NiV4nkJrCJHUcB4dKJH5QLhLER9AbOfjY1duYzb787AkTZMPy
yFgCKaJOGMLQ36N8U2WbF/XH2GWdJ86hGqJS+T95VOjFcU5fL5mxaY1ygmvOo5E5K7d9aOwDxX9n
YuWyiqlsB0O1VPSuyssT+RTeY21OrKOIeS5ohX6r8jpSH3NJMW1yCIz/jBT44GQxpuezNITscn44
qaQA/HORRxZYfnKnz4bgJ4fPNMbqpottdHpDV0GOWhGwIh5GGD1vh3Ibk+CHOMhDTjsDJ1INzLeF
0WaoGH+5j/XCSdZyscPaHRh3XXDkfQUb5ETGtoseitaaAXmg4aY/hg4CGC5O6Xf0ODMu5ZUw/yX+
iCYcdksr7qwqmilsyIt9yr8CrRrIhgD+FqNvrYPGw/B8hcuYMxyRssRQfNdV2wFJzzSxHEtVUyVJ
GLRiiG+g4z6T26MDYCcex7J2nY/1zrLcYal8Ehc97QMy/D3febRt+QpNXfIkFVKWPiogmpH0DwF2
RFke9hb3vj7jbTcsHP6cCLtznMDC4Ar3deeZYMOI5lU+XQOjaAq1Y5kE12zaqeqGiHn2AXMghqLE
qIJSL4b9bd7B3EJVjLebrkZ1qZJmsJtKXCooA9AssYOTVST3BUO88qNTBj/n0nmRTgEFLN6Qux/w
/Dcd4rPkp1tWFHaU3Li6WDoihZCEtUrQoWWXYWsFXfqMZCZSJVmIvBkDrdnGSRSMY7/ghjqN7XrH
vjpjHxtkxHG1PDPRazcTHZrzGMyACKUqEYy+M/3u8rB1sgZtXuggiab1LAHnnWCPKgSjUQe/B9RW
aSJ7qkS+9H8vLSllATjuk8ocWYZg0nlS6JQIRjd7j2VHG8c42R64YCtIixm//fcx5Rl7BBvSuySx
KT+R5G6YV61XVZTC3QQOTc1JVzq7pSIMYcQW2gNQ6ewmF+46DOTYKXmpHztr9jp9uo1kuhQ2C9c2
bYs5NDLG5tuRreOzR5SQ9/xSX0D+v9L1a27T8olwwVeHXpCMFMog++sypEdreYW0x+JWy99HCnCF
B8fLNWs+90HM+y5nmuLoZV7LDzpM0p9B0rSg9/gDChfxqgRWAWZCnlWW1Y2ceWRni3yk/1ETuaFY
TeoPzlGgQZqDKKTcmob4Jh18sOuaj4O0MA7aq3sFQUyztwJLewnypi7o9vu+3ZLNDEBHcSEdVNnv
UvhwXxnLKFUQlQMJyqQAl/kzXTkLPgRJ1KvG16OpVINyjGrL43vRz2w2L1kOsTVk3nY0SnGGB2rX
aAvziLJ7GZBG316+mhGTJmPP+ptyUfGvyKUwAbF6+S4FeUlQYppVpgj35hkHifpX3OMYA97qJEzf
HgTsFysklVF29ErBwT/tcwH4p4mFqZ5k4QOedXlrWaPwhXG3TKuYxaroWYI5zCdYpXjRt54Bg3Gs
vtDVSdhI9ohbjVRWAuLb8l+aie5HzH+MyBexU4Bk+DCR2AUoc13Zxomn5AdAvqeqJPdxOvNtCkX9
WhL8sD6dul3ip4UVE5r78qU5uYRWuJBkNQa8DzuclCOe7awg5pWNPPgU1PgY11tloCY3QEXc60NO
VtBPFISpZL3LfJVG9WkRIN50sv2/WFbW1kX/27UVWKmz1lfz3xPtAgkCJxfjDfeLcZJr9vp7Z4Lq
fCVHhObpJwx5jx3YZU4QPUMNQ8RflkNyLreJPeujKR3VaHvPh2d6H8xGn8p5JVKSfFIHmi0QNQMF
GfQKSfS6R8oLoahjj+rju24dRA8ULJzukjmFfSBPyCvMUPaz8/3E9E4FcrRB3XXqFk6L6EgHqW20
klHqrbp1TTaUwHpvn8N8b6pM/J9x5+NYc/XffenqWUkCYEau08d8m8xn9MJQRYhGDtlbgmECjmz+
dSdK9JWbLZh6s8SjnKtE7ONvHCFig735ADUGDTmVrioO8kby3asTbFoOUQxl6kRMEiLjgMdAZKya
NL04dwZ5guB/TAkHUrZ/hZRimlbet15scKEkclfMOMFaqc5s3d84Nn3cZHVNThRK58XX6YASjDk+
N9G5XttQNRvdiWCTa8e5zfdC0vLg3CrgbOymc6AiQri56+9tIgNsh+tzzQY/okBkPi407/l9/3LT
GywwE8ICF05ljtVyH4LqAJ1o6TeCDkdPrXTmW7Yd+OmtkVxWji3M7mtSBaKzmxFRdiF9wdvxI+9I
e6sB9/ZqOzD4Z+qz7AOCB3vIz7bNmbHfcRgQobspoJa7LJ4FkC5Dejn3QUtRr/D+4Y5FSFPERWTg
b45Qq9eq+vgu2Y4IjYUMiSMgnTVvRAj7wEGDMrdk+RAEjSg3ScO8nbLJSL2muX7h7eFnD81OtRiq
lhct28yycseP4v9m1LR7L5BfO5/rQes2IHERUd1CKSHzW7Oo6cFGx9rdIoPxXkJ7kgqeB2WJtOrE
9gepH2zY3YXaW4UMO6D5Xf3xiP5wvVWCcr0xyU0OPlAoY3bcpG0ABnvY1lSTF9IacnfAqUzZvkDN
gotS/6iBD3FjXPJNlnLmiP6pK46EIdiRw7cUpvnaMO7UWW3LvaE/6sFOuWorX3tnm/tSIdW3q7Rv
1SmOTVFl5xlii73Cn7ClKSe4E94unH0xF7cT2R8P3+3IuejIxuxC2qvAmaqZ17zQ+4UXszrqs2C2
m7m4yageQ7jhuvkjePAu1kg68qUf4jFijTGlnkSjre6kE9TIbCZ50in2sdD6KhGHCAbdcD7LfThb
2fOar06C+gKOhHBW3APDSSIfWg+n66o4TMtdvoDQMVhXAJaYP3/RaVZOdutt+zd5yW/p9tG0WLc+
KY1vlW/zDEp6rk70ftA9ZxwBjTJ/OLAFne3y/oPAyCka6U7or0hl7NfnfKKXM38GXt5PEz0fibTW
nnJIwnKrrBcDP4ZFKRBK50vvbXzKsILAYRqOLIWXcEgFwnJAfeBY/cWQC8VT+bnk962OU81sOZkQ
GlAn2mfNjfcgdp4jJwd19Kt/c/1dmLTq54v+oyKujdrEDJRNQINQ/ClFNH9cft20dGqLZegJlMd0
mdvffXsaf5O80ba+tNjkfrfSJHV0t/nZ1vH67JNzn10OSEM5CVbiD6urNFhTrWfDOPOIGmiZm3Ut
Nm1kKBkzGYVVldFkfNjbmpJ0e5HYrJlnn+9zwCvjGKgNL9ZeqMJNjszbI/DPhHAMPfGM4fyUgt9P
7mQ7LkgnASbW6BGPRavzY0v9hMAQkiSUG3wLB4gGmGpjZ/VOA/GQbbjmePwShTKSlO1n3LDYOA54
8xeltbjaQten86deauWa6UVFGnzYg30+lZ5EZmktRIICDrzyiRIQBgzQ9jhWtYDWGOBVhrEJ7xn0
SqOedqB/08d550+ygegnb30EF3bmBqcHkZBlaQHp8Y7he1pdvRLzvGX44C8t42Gq++Q6jLwtwWSX
EMTiMTysVkNpF/29ffbQsMZT/pBKF7WzmwIIgDpNNcBuuvArboB4m56HSEzbRnsZZrFDUtmkTwJr
mMilX8c3f1bcKCiJD2WrRMW7IipHy2cO+Q/vMUCdOK1E3h/7+Y2o6kx9/vCo3MdAqp7mqxHyhJ6A
MY1OOjScivXjxCt0IbHpyInyDm+SOS+8G2YoT/KAjacweym6QamNO14cZRb25fk8ptl0altIxNeG
5Xj9pgeEh1NQ033I1aLJ1F/ixAfeWRElH7z2I3mi8UfGV5OJ0vISy857590WpS6usO47gx0mPThC
vFKDRkChp7QKzDx09pr47SYFtuBMCdwDmhxh18JNXkposoYqERgTA0AxEy3MAfT0K3suayFUwzE8
56B22+DSzTqP6vP84TYUA9V+6KxLJnQf87GDreNqP+t27n/M44CTJ/7fKVROqGapiRj+ivcl61cA
CBAJWhLt34lu/cmbeyiDaAo182OM26aOMSji1RQEh5iqk1QAo722NpTGIFeQD0QGDTwaKXCKHyd5
smIZJYj8VZ0e8ksMPK/vXYOtjuM4CTVzCWxQbP1HakIwV51Ar3m/RWGc9iEy/8GwvUPdBM1lsX4b
77dTLbkleGYd55pbIFZtWWWAngi8iYLB2AyeS7yEqgX79QhF5fYGFh8mmz3VcXt2faIHScG7u65F
PdujU4q2Ku0Grqf/BdxqkrTU5yeJ9F5qIO11a+S4O6SRp4sIFdzQpf+9RIHIWKLlKZ0S0lo9TsEa
8fwWNbYz6qVAICAyJJ4biVPZv0rYEb5WpMvBF9pWEgc20aN7EM6fnYEDeNgZxvaLpSBSwaazCfW+
2X4q2a50mYb+b52JvLRUWsz4FWf994G0Q8CSsLOfvIKW4i7dV9PJ3Nu0bMzaySBW6IfFgobOwM3a
saKhqeC5LoyIKcMe/Bmx97WEAkwZwaC6mt5uMB0AzLKH3tMidGD5bIqySxAnwwZ5d/2VB5/mZiIS
Yx2zfLcDCHWOkPFaOaAltpY6DnAYV2OK1atuHMs++0zNxdB8WYvYB1WVlKXvcFgfyzrcPDUi5drX
pvQ4l6XMDGABDz3eJ/2odJ17MmMI5iCEuSycF/0mcTrejJX6hoiBNnpwzMokFGA5F8mJs8GA7fhi
cTAWiDMZSjfdrvkWopchm5ThYkbtQuB9z0/CNlKRwFBGjLG7r/LM2+S1s/Pmcbm93jupiIAO5SVL
Z821zXXMULnK1NRuXs+nwZIHq2rQcnBcwFC/73ACe1fUYsNk/kvno4XLfb+LWUqF1I1rhQS1ouJp
yAglFmBGLNBYjIZXRRb4NPOxSymibxGoqKXFwdw+cWoTG3cXXhLQiY7HcUFvhcOQWqNkT8p1bSm0
fr2oNVPQBvinG2mi1ryX7oLg2tOKKSakzfY+hx2OAxOG15zlhE15isF6fagg/GmvIIqMjy2yPiZQ
HU9GMD4WbeD07mXxAvYaM54++vc1aPJQrphbnheNzaFvfVABETuK1/9y8JkrjoSdkcxFOM3Po6Ue
iZbHRq4shuKIcp2+ZnJXH7Kx/WdQn79RROic/zvHA/zV2eOpRf4+eMdAZr2YU4/+MKG5Lt9qLeym
P2pUeSVWuo8bBIXXgqCOKqf7HgtPRk98jCI1iAXHZ5kt2FEeKZhvRDeCSq8pdECp0hEGMoX+CN2z
/yVsGwQaZ6vgdJ9Hw94XwPm0j0B3SOkZ6h6UpEQS0vviNBcjOaKVeuWNr9AkF8UagNmJ7ZxqvwDi
H7QuRJtkbPVdDyePEA5Mnv1PRmcjfJ4XewPEgp9N4eHsrtM9w3gSzbh5aOd3GiNcvvB4nmmz4nlF
uKTBse9HaaycVHXESyzMciFLYmOl4pq1C6sRiBu9wx6navwiN7y1zr8wju3NmP0QWY8mtCn26ZB7
r0at/meg2Hbh+IzCHqV3PpuNaa+keTK2KkJB8QXmfYRpsvO4cHM7yh8b9snaG8pCFqN8hx4BUDFN
5X6mn7coY9+BN4psysGlbzdo1e++WMgugoFbuaGD8RcfQ6ZWxmwIqaSZ1eYMHh9bWqqPVEOAz4yA
9GYRQwkMd1p20TePIpU+dZ9WCuDRNw9o4gKgYjAdG7WooQ994RCNIFdR1HuxBoDDH04TXgGGOIPQ
aYlSDEJYOURibe1F05EZMEZuN5loAk49bqYrLA/ARzDfZgA2Ob7xeVKmiaB51Pu6ImcThePTLLyr
32BmuFq+iO5eaA2WUoSqAWyDetvIRFjbNKASdLxkzLsepGkufliOt7ZNLL0zOhqtEUWPvULE404E
zFtt8OBVwUuq502eXe4kYQpKHdUhPQE1zh5pldfWusZd7JBl9JPgq5C0hZymBqUVev/lAuh2WyTk
8qZeoQ+MHai6r6ebgbbSSQDvGroitUKW+ol1VchC8iijAt6Ikm62p11eW+pBNWsyk8ECTWsWbeQl
CCxvx5YL3iL6GsWTE2YF0iE1BEHbgJLG4e6stAqnj9BOa+bygj7xsNfJMedrtQwcBO9SBeGMrGqo
mgzV2l2cReXyklT/hFISd1at9x9jB2BVutJCgwlVpkzyEEByiwye0XER46p+BeIraqItXJA0tZqM
eqvqRI2MKMz6krJna7GxHtFMZtbWJLhHKwt/eJGKjDEbTSdwYyZkAf2hthslt/M38QlX28ATO4aX
OuSU5e/yX7CK3HtDrBxuMGNXq/WpxnL86Spi28M+r3c8J0kpUUOesJAy+bZ9uQIrSgI/98zoHpLh
Xtox9aKt8i3G2m0FQPKgJl0YwkwpRafUKpSOOvYJ1KoI2IwzT8jWljZBp5BCmgG38H4kFoBd92/5
1W2Mm7ROdOTb9WPEE8PxBOWMI/b9NpJPKhDp9Rd3ZqzyNJIRzl5LiIR/OYrOGT8PAeAUK7fqfV/H
uTwFt6to8mGJDUoJznzuoAQw3puSLBJQev1kC5wQqYygM11F4PTJkbAJcgUClLQSqdj9f63Di2dA
kGi6cuWlv9OI3q0XXK6ZrLEDyuRdqakQswgBBG0tC11czGCUTSOa9UP3W/LOD+CE41179Tzd/qhV
O1tQb8CIt8MNqdwsb7k7l74TCiIv2xEZWn/2X4dy8Z782WsqZ/MhwQEU2cy/g3tpQD/ApQFx/6yF
BtrPsP3t7BtaPx4kMtxK9uQ9BKL1XSXQ2fBbIt6zfkkUXROqoQLYYNddPr3NLlUqXNp+pPpMlom8
7h352XorcREux4CWs7V0SECOf251ZswSG/vNeHlJC7BOzITxM29MPjQnHfEHfGtY1PuQ1vDwG28H
EYxAr6GljSkFYbgQY6If+4iOXoCVH65I4DqMQea02+aqaeud7BM+xOOKjbIBKqolhf+Fgxd06B1N
1tD7RbKLGCXwNkkwzL5zF13vw4CP4lQJhnTzDy7uB4T9Q6ovvdLCD3R5G1i8KwVBTFWi68tFqT3a
dVodMe7BpKzCvTqb0Yx5WdYxNAwHzuxja+irIha5WoGvD81IG4r4l3AGHqriYf/cdegU0MllKGwC
M3fgngN9gDxSx/jdLA9VSfa/i8vU+2oR2fLNw/mpT+oSSVxmsQnR4z3Tynu5WRUXpQFFPZ4SrXTs
kD63oNeC7wAz3P01OHOfn0whvHeKMGQyXNECVM9FbRtx5b/+jC4PoDSWPbaWwVksyCZLMuz6ylhX
yvrMk9PgYdEpGduqGq0wIJnZLIL2lyn/335AQz5SAuM4cL3Q+55T8cjUOZ1w2ja5ioGaNufpKijT
je8mooSFfxPPzOjSO8V1jJF2AI0znHJLccZsB+55NROabdENq6m7CR/FmDHERzZsa2sIhgt+qCqE
+Wmrpd2DUT7y1x+2yEl+XjCToqJPu/FTWH5L084DGRfYsIEIOx5zpIj9GRFB6qQSBkG+6TP7gO9Q
6KVSIdM0TU2q7Co0iKp1G2OcBuCWlTKR+WsAxHMpcDHWNuJqvjBpFd5Q0GjOwxXDuh69oUGGafBn
ngwIVqlSxIrDiWJ0Utz454nd1tAh5NybfR8paemuSbK/6ZcsWHuniDxQsmANj9LxFZl0dlp/em8J
89RDHaB3rYPvzn+5AMX7y6Y4z19dM3wsvAwMhmafMuZjZQgkhU9wLqf6HZx3e0QmwZ80Jg8CmAqj
jFNbAVUB596Ei2QumpxIAwz/8MW6UzkTnsugK+5oiNiMKSwC8OD08t3MQu+CedC5cwlloN87q+w0
LimIAdMKAI3tWpdjkOSoLE3uiPLg0M7yVMY0PiOqv8JE0Z/LUtRZOLhY28A/pi5T2Q7x9jdvFR/4
BUKrp06i50pfDM1Jq/9hMCvrbCqHFZeOKJnfrSmEy5TV5LXA6Cpg45XSiycGR+NMFILaG4Jz7TG9
8FNZdU8MXkZQlu+l0WDS72fP8VJBqmeCDFF/p7z3jKtrmpzFG/CQKI6NMKA8atpnIXElJczu8Q88
veVLeCaM4CqwcGt9SVQYFAbPUryEq/wMYpjl/OXtwVFXikDpm+hi32+5bbPkGc5l8pvfGoPmU+KV
Q6V0dop1t8vsQYI+xpUGhBZYM8T3Vsx5DJsr6a/6hPQqQ0BdNjSl5sDi2L7oboJenblJgwt6KRjW
emtgqM9uCETy0XllGZ97Fj4ODcEin/M/Gm/d7pKwgXpWOhz0xH0CMyMQYHmEoKJxp6/9VJVtEm2T
Cgi+EmFDnBnQ5RRZqFK8utdajck04J2/gl5bQbeZ3ZG+WRs6nkMJ8MoAHfodx9GtG27zqkMmablc
7T1Qqwczs3AOlT0bXavWakmB4W6THTh5u5JeBd6uF4huxQ169Ekb8tYxNYn0bmcw8KJ5WcyFRNie
UK5SjX0fdB8u+mW7VePdLQoe24p/YJ0WZI2MDPAOj5LlOc65hA/R7oZ+1Grlh8u2dhT/Y1QVMGeT
XgD85wPCAbyJkGEXxGAjGD7Oj5h6wbfYBdGYP0FMFJ/mNXonR1al7sTpBk5DIx2s5LoAl62zhZVA
Vkav8gdBaiZXmhAoPTVFd99m6mryMkyKz2AJeTJQBdplDbSXAw6SINuTIf4N979Lqmn/xcopEqLN
YBEFzZ4y06nAcXVZdvgz4+QiSdIYZIo+i8NeY9MdpQEVcMU3Fuy509sxBm8Hb6ns8KfhAQfkpv+r
BcWsXg2b5zEW16Z5QHLyooYisA5e7EF9NHjqjaviG9wC+idzEGW7BPLQCLFqQkmG/c266vExB0tq
rejQEh4sGQlDveLe0rl10xkZ1EKquW5mNODUI2GfXTKg9f4Ds/+cvkUXX9L04aZciS5sY+4oBRrI
TVvvS202K8pwLR5g1UG1yY2H1nDLE5Vg4bCAhnUWu0KEF9N9j34XEpAAAInPJtI/wjBalHgOI63W
VFVVqzEdHfkkVqFqId1lgJDL9vf3uYGw9h9qUWVEY2OHzc97mJdT8P4H5Dcx5UvXfrQGs9DmWsvn
lSz9gAJIUOk7cnwPPkd7gVH9pfYDTlJspZ3rh/2HU9sRVCp2wq+VCQssgfmLeumZY70YaThTgXux
1QoALG+U6UE1lzuMl77Su4khlI9Q8TErg1mGr/fIRx1kr0gbZRAIJNT306ufFXvsiOg9Nkq57lKs
P/4m+2WfiUZDUmXeLz06r1LCkh02CFXLpM2g7ZqSGd6dx5HRwKYv+3g72i1m8z3G4VD4HfBZxCec
swaE4aql8zK1AaGhlghysYjGro222RrZMyaN/aI7pNwlso8AEBhlTS1Tpojf7tVyOXdhGnQJD547
YPRv6VgwKeNTa1xtMlPOhOt+PQs+uh/6dAsfAznUMdUIZ8dUuqVejlQIGN6QfOf/sqxH8JJ7bZ7T
pqqy99p1I5uwDJQJBU/H8fa9+0Pqj9IwRxqD+t7K7TvzyUk5g3LuAr0sLtsnrGO+YH2ydBICgR0Y
V3aunIQYePnsgQs7ofS5Cy8zY70xpoSXrPImTuC57AQW5dkzr3rjAwKtWhch+eAFumDeVCbCbEmz
i0bl2gZUDNOnuwYe3WPv1Ce2gqG0fXNFdReqJ255fkpXkMDe/IfmcaK1mf2CHrEyjYOmJxKjOHWx
npsHbPXDwr+XUSqkjoVlbOyu4xJKa0EMX+ZXRfx4BXJUBV7HXFZWua34Z4vCyTLxnwpT8IElNvdf
rUHf61GLRg4VbaztsmiVQ8BM4AZwmZ8gv4dpJrfU3MqyD4qpKS2U/8+TZ1pfbAXhwnCm3qINnm/U
OC1kqaVcP7XkYduvUm6p2FPtgyuaZk4FMRnBrAWB5BY3mtUpgmz9wW73w5xMDBLaGU9XFiy+JZea
0z/WbSvmcI5hTUREBFS698SQyxhqqtD+f1kvf7zHSqBzgVRStHv3CKfmfIthbc14cnLXEoLx+Z3g
POJM65iUXcWczkqBYacHvYR4I5uAQwnV98qlgytBLUn/cFgc6g2aXOf9hNlU6YpR/jbVmAwPCJYx
9Hevk+ihRayVnIKgga5pnzjUl2sd5ai+mW5+2qIkat3WPM3i90VQaRC4mvCQ6+/e1maDZGBX0aZb
xyMN1GVchfbtHS5+IN05ebCKNwSLqn3IP7LRkrPWJudl8ggOH4qE8YyCEDiFbTc0jIPrw0HuNh5C
IV4XaEMKSFJmUlO9mk8LnT+YI5/6Hr+Ki8viyCc/q+ikfRSH7uwAqek8rpdb/EqP3AqMQKRfvxvm
9qgghgAU6M4X48HmrkBZvPmMdzanWZCihrsxObncGT/nZ3TlPercsT8cxrOY0bOv37RPssVcyC1i
BUYxgYxtexjzWUOpNJt91lYu1qq/pDMGM5uQNMLrhv5GO+4C3psjz//zSnjijGkO4mTgvU9qEdft
ykybolxXf3Nhc4zgwLYI9I0ugBNc3+A98RCT4TrBWc+FpMJDRRgQeJqKjx4mlvvgaZUYa7TGGUTu
6G5pBGrKCd1VPPN8JOMT5NHKYWcek7gbX64yEl7VxdKfifRpXdaFo6W+eP4tFbtv/WH+70bzZpYf
CTNB2UbewcHOeNIrdErEt1qO9F0t3ovu8oz3LDCs7E1yeNrM3xb0av5hzR83qhGBtA7X1hbdA41h
mLGuzSPD7RFvzQ43AKx+d/BaoznGoC0K7Bcjp5SdfSd2VWvL408z7lqlOa9Q5/DN5YHbU884kZkJ
MByUK0zQBCFFmuqEqFk8yOAa6xCtguc/XLuhsttLOw9hV1Yb+jmCcpApoxoEdZq19UgdNyafB6HT
toe2MlFDV57QFFbis/30bAzhiOEgQqd80pmOFoArN4JPO6SKB5Ajizw0pg8m99Azr7xyXcwPTIe+
gIL15u8ipPGby/4L/wCnPWmCHcoqf0lIfSsW9wO6IrkLpAFwAoJNPaSbl9tUsYsfQUlZPHuclaYU
8uuG1Y0A1J2p+qhYTW/JIBeK9c9NeCJtv7McGjz/JmuQIFI610bGn5PLeO6wGNz+IWP6VmF3soT6
+GN+0DdMVWuNxdSyIm9rLcAs48BdKobWDH+l6a/3csCxqLoWp2hhCuyzpFlZRL3HfpW7bbII1GFJ
2+e52Dg2TG4PDgVXZSK2N2Gx5uk8Meh1HB+hw2gQM01yPiGpauOS+IcOSChkCuzbPtxPnHXd74Ix
Zc960k5aGTyODNhHE/IJGCN6FOdwuv/Y+m4417XPPWgkrdV+B47KDKZM3uJoZ/rVbbq7sysRfPBY
C1NBDaO1itFs/xcTCz1q2Dc67Qk/BBPOtwb9ecOE27H3zV1IzLoc1wypgGNIJTZauKqqTT1ueiB5
usZRfrun5CCwC3VEgC+DKXOAOGUzN8Qc3gtwyXUApCtnVYSacuPLICiM5SbRLecoH3X+J7dVSScC
XtVQvsCB0geJmlXYr2rgLhS+s8CPnxcXJlezH0ZysgIXXodKBaZO2FjtA8ucWqRdCOnga7vm7STe
1FcwCI0L4UJ5HOy9RDI+Gz0CxKacVPcjXFyYvJlkqOhCJUnZNFMSfTOHT3tPtGgy3W/FEmF4wJPk
67er/gU7AzWQY2dE5Cus3aiNczM8CI2XzNzBpBzFad5DNTSerbPwjTK9BQao/WosFzDe6KNfspTS
+8tF+JoIIplJ2BdlcmhAWoEDPhu059Uv1mPoocz4hWaPib+ALgnB2fVpuOvTo4kd/2ZG9X3xvP9u
+zyxMeSYKBrgfndVMdDVfw/yOGNKmK+FHqkfAXdmXSsfaqGvJ405v5w9VpBqm2sTWK+O6U6puFOK
Tip6Z34BgNxVEOgoI8Wyb0b1qAA8SBCTOWJtgiLuImo77+lDfV/5CYPvAz5vTTrjzrvVXEMO9WL7
/WnfnJrdfcnTtXrRi2SUucIHI2fRzbyKAcanZHrz62m3bS/sf1EZWVVPqTchcIhiY3jlNYVO/s8z
13f6Hnu0OqaYp3Yq+gfRR3oBuwR+n68cKdDR/dXNMOvgc1XMsUbGgj49KlMo2ivJfR9XnMqd6EE8
e+H5ZsbTHe3zE9OAf7J8vyLjeubn5bjv3FXcAxPsoZeNiSXZ/8bdrcm7/TE7mHuCOrrP/Ae6DFsx
utOoCASrv+CkcoEUJapv5YEOBnqHANEAIYClvoJvUzW+EqNPEYBErdCNAQAUHajgeF+LPO9vdUxp
dlwGyvDPlSZOhptfRTVgxdwx03Gw2BQZYoPSmCW1n+6s0IKPF7tBRU+M9Red1O0GIkE202NLUaoI
ka2sbiQp8UbYP6X3Jk+PGnyguk1rv5HmM1V42XpaB5Lh3AHI2izOdls6fS+LXAMBf1GI1z1PtK/c
ne+myJ4HedkGJTpsbn5AOMV3zLsTmz+oGGMHcByu1ywxArmWgNgZgm3jCwZiVcrHSn2EXtr56c5C
kH0xsEJj32wNENVmuO6sbdK47nATLt07twsCjUzYvXlBPgoxcLnewKYuZeFVWw14A3zjxKIc0TH+
OoRv7F16l9L+RvLXoQNgMU+JUflpShZYBgRtGQq0jdqgljJNKMzMRbdu1Bdo0vKtWTfjEzRZW+sE
mf5ZQ0oTvW28afSdpd1xsi14GOB3RCSwa+j5W6pkBzIc/ZGyVOVLj/lXpCDusBBl+m57+Clrs0ud
FXZxPzODVU20/IW5zi+9md28tGSKO2E/3k8u9N1U7jl2Px2j6RIm70mDXGFMFooAM+0ZdfH6+Ss+
n7j3fgr7qypKgvM7ynmXpAjqQBwGNrjGB/ZDYNNFaO6xkDNQAK1Rk66RSLaUACiLKhrOYXKT2deT
GtIw2/a7/+NzFNgCBh6dTGDG6Pxnx+lzWcVwMgoZLGJ1h2sUePVGCYaDbphSge1KY0ls6kPURPKh
XDzjJ4uTd6aV7G8NBMab6mEREgtVLhum9zmFQxD1ou9UlxbnuR2h1yNum+fIvC5W9S10zcOLPbr9
7x0FpACzIGkaEoXqzmtWsFCmKm2qXhFYXO7vf2GcBkNAubqA6LtmdAOl0685uuN7xKOmYDqKwfTU
IdVa2Dhyo4oqJx0k5iTIRaHDYcbZ6E4WPB53YfrZLrBQAlJognwcWsKrQGywEhK1a/nopVwINn+9
gLkpeAjIt+S7i7jAamYWi20O/XPoXWTGeM1IBjFnnMoeM2odJqBkJni+ibXLqdX607dvjEkYTnRY
PzK/F+KHtwFymNZcu2NPwXVNP72Kh1VaCmqhPmLNJ0X1y849y2A90Z/2JB4ZM+KbSpeCDIZ20r5w
WndHbnD0NKYLamElAOvYMpljw1dJr817Yp4W0aPc9MhBlPI7hvQhp17idWgSCC3Z7T9Brhf1e8ub
2k0MGBsL64y7xCziYJqBf2/FJ/8rR8LBH9jD3H8uI9PjD4GNOle43HThacxXfWIIoiA3ZwZSB7T1
PGRfAskmY5tCWjEuslzitexMijOjzANDMoaBjvGg1UNuNybLUpS43pEUz0iHBb2xjQFZTOdHwp5c
mK1yB+HHUg4nUa9+Jg9kDiFrGm2Mk9ir8SBaWrpUpu4Da6DQh3QjdUs9/S0m5o4saXmaSHDzONL1
OMrDI/Bai4CuIHVwc3AkvCZBjH2NAtsApJgdBAPUNpdmNPqcwoc3W51GXO71+MzZwfk0dDXFKTRm
WrdwFs8cVKB32xOKJoZBnVONXg6JT4i22RwHn914v3hjxjhtgpj3cdpXiabyX+SGOG21kGb7ncp+
9wAyi3J12MbClteux+ILMqJ/0gsrBckv9PHq0ZdRO7b2P4BHr5TBJ890Ioe2ixjrw4oDYz3CgL0C
0Q1XHU4oBo1bqrUwFSzEb9b5tNy3Nr4BO7ttsmiPQw6+UInwLWmIVte2SI0zEQCpUACM1BbWbp3x
Z5jgKSW+7z3jZNY/Gmni7GLoNG2LrbpQcE4Bwr8Ri46BOCwD2cdHzA9yPd7LFSJGs4Fm14o2U4kV
cRG3xrpyVCYhX7Dcft4GKQfefwLqTorqpZz8EHu/vIn5pcS4WGpofs3FkeEdvTt/3UnuTXQkU0Cw
I7aPfMqmz8aVbZxAwvPdrsj7CgCX++GxGm0AgjRorKhHqqEy1CuVHPZkoRh/KbTU/a4e1IUg2CQJ
FSVzKvfa1aU6lXZqF4X/sFIzsipUjdoQ0S3rzhWCccizKnENne937VOZsBrSE9srXWgg5zDKu4U9
F8mefMb+0dyYs0iFmV3578GQhG8aGT17/OzKPVsTiBHzyFNCqyn9uKJWSbQgeW5iHczJVsFZyDdX
jeniYHzU4Zk8xtCJWcfT9TM2rsXAvSNpzIJzgClwDhy1Mu46bK8itnn/hCpSEjFtelk3UKhApYZo
5aAnyHO4BoLXtCkF5hyl18i8xg413wwlqqPp264i7VCNi59wdX6Bg8BHEfMoHewMNxxgIamCRKfw
KvGGsfreAhg2krJPJX9tiIfEHzuYFqP3KR8FzftMyq5HRXXe6e3TdfObVWq94n16Z5eRZLWm1byw
chvEw0Pz4KCc3M7jOiTl7E99tWgF/Ev4gHQxDr0jhW0obbeYXf95Z6rPMEBuNAhBNJgG3t9FGzkc
/itAWqDvaZ3HnsWjf+BkuCRM+adTMni2wIUQwe3iv0gL2/nXikcUxDOkQtEVahFCAOgIaC//8lOi
jPhjAp2wF+RMGfwi/sGmtwNbCBOKzJcvSZkjVblIhRousFslxfksYG7PmsVCdOaYVpOm+oPrpT/S
sfDOatbl3AcxEyUekJEF4NxHsOIrl8k1oFEjeSbCI2uOcBqns2yiLAiOfMj1CYDlOZ20RlCBb2e1
zkANrDxyEnalSBWuzyKR6ing+oN8ecY1peiiDZ9wQ7r/UyttOLNB7XpieaW1tQpkALZdWk9S2D/J
v9O8cR+lpYGMiYeLtdOEYEcZ7M2vP0IZq3ypEqzUABcTQcigcIt3qtzMHYThBNIF3R6en/ZWXE5f
lIMkRhXY+iiLBEAxiJcror8fHx7NxU3DO2GTySz06KiaKh2n1AnwUCNn+T2HTLDi335BFlV5ZD0Z
sAkzurtqiiONwDY7IDKvMjR7KtaPOa4FdrbLstWFmyEAzpTO4nr+dZ9n4KP+Dg2OYfsfih1dKic+
jDtpmvcDySOEvdPzCEeqB0VRhfRMWawo/rvULtUeY8EqD29/f+K+dXZTnpAWkjXgAoazdTcYEZIH
a8Nieu9Bk2TXGsbSHjPiB7kBXkOwIDKnDGjBAALz+O84bpPTt0WHC1a0teui6Jc1481ibk04PASU
uW6jtB1xiY8Q7fVKgqbtcPs6k+cAjzF/s4WMe2UVMJVYNOcCjYNlpcTGE0JXaCD7xTvE+NoorB6D
Uv37Qfdtv77iyN/12bDqOQUZRcoOs584d8E0AwCRAc1dZW/lNZwX8bSYtOUvxCCCzcnAndKd+rWs
JN6oxS/SByJvywDM5RVv5g0r8Wc5ZMVgLcqyoXObEDoyvgjdKfhFNkURn1Nb8p6WrlNE0lZPLjRy
U2r5CY7dWJ8JuEf3oUySZaSrJuQZKEzq1RVXu+zUoRdZ8CGoXx1NEy4rd8dArp+iiNgfjViKNB9z
o+FVpS+lwf2qJY10NodbKYhTWLWuEsT08BMLJhEvBiKz7Cy/9n37TrPUzgUS/FzZDRSv5YiMTlQg
qWPJk9ZChZ6SijiOZoiELNEMXSi36Sb8sVeCC/Nb+0skF4s5j72ubS+EUKt07cQPEpZNcWsWGktq
2S4urVMXFgdZASzHEBhSHjbSU2k2vkleXgKAjOyDTK6hcc03XnZ1fFlIdusmQgr4rrqntooplac1
hQhJEvcwH8/nRxxy1iOUhOudtH2gln4qyBJmunSj5tw+LGkRgAnhHSAjPDkv8v4Oo5gQ8Xs9sGv6
pnCXtanfvcjNsIxB1ddEzdpHWfFTpYWZb7fAPJ0PGKAYsTjjWtj8NsnbmjGd5aZ25ltJGawxoQHV
Ru9sNo2wOjCCNh9r78AjP1JW8AASjYoos77yRHyDV+DSqb+3DfFkxpn8CpL0IXZvy/x9v5m+MBxn
yOyOIthQfAy+YVM7hsrZ9ebk8/JfOaxYBB8vHqzN6B1GRIw4g/FeAiEQNtgFlp/uR4qE/GBZ5cn5
i/znWT+l5YoRyAWTPeeLSChJOOuZEWu5NetvLev3jC3Fd1iE9n4AcnnyLCkVpKi0BaM3L2fKlp9X
sG/SCHb/5IKI9/VKiZqn2THhUm1fArXvW1RPFFrsUv0ZCZEW8pkBlsJ+aEfceOLDe8tEgeqVel4x
ZLIjzYusQAWx8x6KmAwjsZf7Bxae0vNdQOUASqaTxiREctUBhp6UyPmwLOSbbw2LkQ/GJCjik3sR
5TZfRIDHzmxpcIK00+jRduVw3DUrrkj0A+dRDto4Icb5kRSyw+md1+eVGcIMUQdYbDrAZs95kBr2
xT2vFLE7m6YeFBvj7Eoq0ycQKP3Nlbj3ZUwsNzPNUjCjVsjr8RTtzxoiqvHJ1B850NXQuSWulbpA
8Bi+FJANYegza99VvhcapM3Q0KUI2HZTw0o+l1sudAcFU77glauBqqvijWU6OQo4Zug6H6HCjjuB
7hI+Axeo3oi/Ma94f/FOOA1wrflV4LosEkzGQsJvGZpj5Lq5sOfjh5vWN+G0iuTw36qX0pZRH9Mv
LU1QVC2GD+tUGNckUzxJ+FCJRIfbMuB8TN9y/dXgnMHetEdfQMMvHqjCx+MkxcWaOP11yfKZI6yo
TdoiEREwRkHB6BfLz0Kr/r/CxXB/tLZYb1J1m+U94WaXsjUUQYMnB6u8/TCJvlzUp9u3Btl3VVPB
Cg2gPRVs9QbdkzglUflUKI5KxZricGo278IL3lQwt1aqPcVxnFItoe9AXgheWiafcTjGeRn07koC
hjOotxjTX+2cFQxrRxs/EXFKXms0qNIO0TaY6Nek1I8nsCUZ/FUTcWl0rEbmAjb29BS2EH2dy0r4
9FZTiCUVimC3gJseTWf99vJnAXbLzR8UALOTJ7r8tjgjPHkctIJSaS4E4DO0NQwiuzLXRDqAthxi
TAaEIfg0XpV4YeH6VSwIVy+DTexQchyYvJ9ogGUCPcwUA5l5+LQeUGuGtT15BRdRQXEubAna8+TQ
jLxuKr9DNMxt4IpMqnSCtOB4Fhtn27BUL5H7lQsxwF9tBVDcs6gB/zlD2VbBRjmfRS0lS45p8zvL
kDKsOjALIE6O5vhbdUZ3c1cho9Ypb9yAUBb+GVgfymOY9zWpzm7T7VbWFnSTvushxYO3vgzekial
mIm8Huf2NJlRqge8LcHsoRzsdY408PC9RXiZDCHoPM6YM6Oxi0gLwd6/1M76TPcQZkMhiqtSXsDy
ULdRCbx/6lDmu97RlPcRVkC+tiSeV4aJSjISXRJGz1dCnIuwHNjriUvR+zjfH/y8icSxLrzYwPkJ
uwMdmXijY6cv0oP1LppfFV/sOdAnPLEVdQ4VsjxgGwHYUDZ1LUpJZ7E/IEvzd+J4I28KQIZoqNr6
n6ZN8rtrd3eYrhyGq+S5hrrdROL4Ze1eUwCUx2n+7tIf3xtg/BUA+/dH/uDHT26TOEWDB3v1P0am
+El1L/4E4lyvC59OAyTAUNe54lsWt8OHVDtGK/BI6exmtFd7mdOfbya4hp+DF34vhPtr9UqUv5ua
8Y+f8GF2NqeXIxtIG3nlBj0jZq1RmPYewjZ2SBLu58Guu7ccj/e+JTirXzxYXcsszCL2tFfvDZq1
ZIJ+aYIt1PKynFOtepRijjeVKMToGl6qIoquukj96UqWF6W3ORnVMIYapZQxgT3AIZ6CmEkYIWRF
MOPt6PeuJA8V5IzyGxweaSb5Su0eLlCisVxn1qFs56n3hmagSuvJjfObiUqtM0ihF+ljol4YWDz8
Pjjna36TNTJneAnAGc5+kNrb6Cn9jrWp/keO4wmVmeiBMuCSCJ+tAlz9HLTw3H6enUtUITr/lI2G
Uq653RJHOjKWDpPhqHtHhV1f7W8vP1cEbczyLErYJkrr175AXny+2tOcfoNvdouJ/jI7t7VQnsNR
/XLUu12WUdOlmrPQpZpUEJu/CYKacrjxhP6QFfpLWRcr71uiLGn1Saz82R8M0ji5VD8DZ4eZOdHN
Wgg2+ry+PA9lsDRNXQ/x2Dnnc1KvJtrwbPrDLveMvgi1w8Lwue8VR+u6eeDVF6LV9z4VtNncI0ac
hLW7U1I3UhpO4EbV7ZuJEZzFWxmH91b9mRDugip+FumfQFb8x+iHbPUDSIZ5RsTluRWeEGL6j0vL
GOceJSBEq2rKFqWcHP9FbPK2Ot/ruR6f2bTQ3/M3pzWt/4EVHIda2TLGWVrjFwgiAXaQJ9wVpe3A
dOkr9+NIQdnZmUp8WbuXC1eFeQXo4SK1ZLOe5VXZFeHOxjsZtcpY8KxBYvygEN2vR9M4L6o2PhDY
MHqZjK/NxiHzPSXQWaFkcDVZiFUpEFrzZQa38s57iCrJZYlfc4O3QdhtPCYp1XABL0iFZiugBJof
/O5bigqOOPeVzIv6+cW89YlFCO19OBj/dqQERbP/efGzxAHPkPkHyKGfX5Up4zUUOg3wP16MjI0O
xE5MgFc5vEYzNi0Ig5sVkEvt+dcQOX7ejYXfDW3N1+/YZ5pL4UP4n4B/3M0xxBdVWBmtVLj7eJ2B
/5YzrDyMQ/PLTMccNrGjD4qXT3bNvRFo9YnFo5TB29uXlrIJ8SombxJhFTuM9bjhFIixG5ndEm9y
94pHyWNbg32CFl43iSok73K2EgwTTp/iRhKgV8W/ore6CTMydUU+8iAAekS/lxEaOTYSZ6Q8Y4ua
qf9QPMTsD5iH3QrZWO7wYJj0+rrdodjSSxmZ1BhgU+LYz8UlL5EBMlRLgpvujF8tgI0doJcQnrgT
NOqWRMG7OS4RSbN9uc1CLo/EhoFWEU4SryxCBaaw6MCtUPUMPobYHXYAthMmOO+WBRbrJjWppjAR
kjVZJNDrDq2WdL4/CG2AM4a2MUGzKw7lWOzGO5CGkU38EgED+RUJi0c4xl/o55DDX4YSIbZeUgQA
FfVPNGArMUgYeGWW/o5Ro+IOvUIGRW2tdZ5N7D0Ar4GCQE3eGvk2nLqpM4YkH4hiaqinupUenXUv
qyl54H96FKkO5BWnRdDVc2rKhjxB7PmqvxAfZMfnHyfS1e/pjbticcP6UZA60rAh3NnoC5ZABloP
kf+5Mpuw5CB6vQbjhEVVnb9SbniLe3zO3vMVB5dpUPKxrFMJkrWO41d6TMKMkaScX1qtGQILOuOc
CpIEggGChIPQ0MAwoHxwJZCjHlP96P5VruFl/DIfBywvedB6a7nf/LzJrFoeH7zrL1nAsJxdt9N2
fqhPwPeVrJGPlaK801YzqxNzNCi7OPnuY7BuroKOIfRtKbB65OkO7cHXm18kivlDBEJt2DSKK9ds
WfkipLfvMM8oJPfbSKmp2Hgl2meM4TtAAfJcnv7a247kWBZWs5u4DVbdf1jKxAgXFN4VC+1PUW4K
5QcGy/BssFzyNqt1DyS9a2m6e7A/NVAmU89gS0pCjubKVh8lkqPKoDDrJ74g6s1IN8ZfP+4HiDjN
TMqv24lyqsTxgYLLmcCq+MGjMT5WA9yswpw+biGgi1tCCOkEjbq7WaAQ2MuKCnrHgkcWoCZKF8QK
Zorctlm7cXX0cz6ryvZsF7KTXymfE1/9bkFD7b9qaxxqDLaNt5+JmOb5OPFQzcpifnm9zTvoW5HQ
YTUC6TqAca5SKmA4GXIKIkfJTNYU4yF90qm3IJ9cFUpwQpo0i7jLZ1pv4+kRbav9RWO7dZh9Ac4q
u/mpxG6UBaNmeLSXl+pk+8tNk7/QQWlU6bHR/V8vcSU5ORdD8yVvmyFtQ8jt25cBfXKbWnSYJCaW
4X5jkZ60cEAkBDI0lxGNAU/UzwQ+y2VH6fPs9fqlHB7B2g8fc25oSHdysvZDicbEK8d5lCW4p3S9
aSEEbpi3CH5GM/14br3j1g/qtMasXSSzUP4lryyVlGNE02jyxt2VSGxBc3n+Mn8ovcTGphyXPMyg
KQltb/8Z+Nw3lMq1nedUHtEsu+bUjTGgJ5637syT3Lr3gFj3QuXfZ5opViHeA9ead8s+3EwHzyiE
ubteyDRxzJ1SR6l4bkiuxj6QnuP55aqwIcm992aIxMzQCC6xAFiK7LI4Okapu74f0TShYDBDBlAz
pmFey90YdjCSlOMZ6gyh14Uns3MImz468zybUuEgbWhKO7518ejqXQmfnD5JkF4izOb20uxgHgNz
mLWW4vmoHn5xKDur6zjqV9cIzEIUsm6Zib3oxarwiytHJ8BkWRvG49Gg9uGKlBtMpyPMsGwImjeG
ObrS44oXT9z9PtEtKyrrpacBFZfkfLoa2H0NBpOE1YvziFCNJ/wCS9FvijPhsUoCByJLLPrpypBk
MXF0atRT741zbIkAYzWPY4sGISAbmgJat50RZ7hMyTTJJoUkfDb5MWATZQCgwlEyvoJ0zHWHdyH+
i9Pc7zSaVtDjKtCpXUlj3c5uw1o8l1i8x6u9l3rmUlmwBv07JubrJ/3W9ojAyHCWwrGOJ1DeWBzt
cODb88cwUmp22zsedBb/ZLwLb964y6BAi/cjv1K8Sh4b7Rflsjzacq+l9CtTV2ujpZ/CxTeRx5Mq
22sLN/jsMJqck2w/UCGIdn6TT9lTOGsARESyJGKhyr6bHf4EGbXPU2wt0Ye14BcYx4DQMtEURJG0
8Yua9LJce/AiI/2vcCsgHzoA3Fcz9T+5ovgLKHaIm+QphlAvo4/adH81shBcgNgzPZGevCZp8CIZ
qLEsCHrsyavZsu1ycfrJam76tcaiLC/26jExVbzhHKtJPMTxlvaxpwDrYQPHSqzNXxYDHNVUYPXC
V8qdXmKPSpZztj0d8JeakYFQwSZT0pnIR3oYBkMvOnK5KP57/8YVjbpGPy1bbL5PEmDCSQSt0UpA
UqaPiAH6/hQdhJ1LQ/j4ynY889PZAwgEgpipBBDKYJRdz0Zp+nWPFJz6vJYmF/BgtPc+G548Adwb
yNlbQLvEdsc8Us0/F42QtAIqRYueSPOG4n+FvhmIhIvZETzVYO6s4GgOrkjvhPWhS71Wx35wjT1z
cmD23aVmxO6g+Wdk3o5PR1kiZt4Nm+LDPEtB3Zymei8q0aQyZHFkspreTxZKwkQUVExg9PO6PuiU
+YvGlKzGvZZ84sVFpR0KJmRYb59YaxugXHPSCzTlz4l9KNFW51kNjgXyXqRsIW3tNu3B7s3nQC0d
BpmOGCadaXIFkAa+efO5lcciDuA3NpmZH7LCrOafyn6n4VY3X1tHspshwBjD2vsZhkiNLobXeBlH
he9l6LKsQ0jtV/qzQdPaHvuQp+P3CH9LIGqDBJtFzGQodD58OiaLPIa1oqpeqFCQcnGuDkikyABH
ayn4O6it2itnKD7uyGdiEN+4/dEMYTPNAo7g8sR5XKNaAv6aM//mNYwMjMXYqGUlNSt4ykZd204d
QwwMhp41NUVr1wBE1p4Vyku/eRJ9XxQg2U6rJfTIFVdJXK+29CR72h6Ihw26tlZRvXg0B5c0ptcI
RtKboQ1rnYP/GhoCN/6vpv6jl1uU9Z1oGxjxy6kQ/yAylA7xL+m/1aPTcakNII+g/RN4qChQFMVF
Hv1ovHMJvKptm7Afm2VWffpvmtACrXE5x1y/LpAAofzbgsa6YUXQmWMcdZD8zi4NjdOT4z5xFIDM
2Isty/WncQuWkKZO071u9rfP9oeki+CorfPU8dgXj2cAVHZJ4wMtuFxI9b3q0Omo9QcqMLSfz5JY
1R+zjLhxi27k3aDna4azB51euDVZgiF/Bafe8HTKlXT2Q259ln1rLvzGUB7sAyB1++hbrrMF+B9U
rAuotX/9wznh9dSwgYILd/Y5Caq19w/h6tokyNGpG/VEMpEE+2hLNstIKheVqD3IDbFwKpM50yXS
Dhrl9Z/RtJWUVmCXrRaEtQ5YGHvHiRRtIxoEZ9QbiJl/SE9YRDgpfKhD9mSbv/ug9y3xLbY9Kpdk
qHN4TcNrIkzyiTR5AsBMPFOYWQy6+MYvaVNwWOa56yjNiSSlukakkXCRNMLz+RiPRCyPvlAMzqWl
etRdBq4hHEGptP1G7gU7075gS+egD4VrGpUwfQgZKOUi1+1CFV1ZXyavVm8aosSUecuwoUEIX8Ee
Iple7zGBHMVk8QMKdDMLj2soZWkGP/qhmm5l4PT5ijnEQh630iWfJQIOGg4iZ6zrCt4BSj1/Im5D
YXhhi8Rf7FYZhZyyJtIF/h6MSnmWO6QpvLZfZdzJ3QlzX1+4zmkuIqk/lNxy/caDx5+k127sYUOx
TQHnSIp9jY6r/3AkGRv9vx8i/tdXD1wVU+acbqgKCUmv+YGdrv/1QDc6u9ldZK6ME4ndoabCkRd7
eQ/PKapUZUjTWuu/f8NWbUv8ltFsv0UqLgdNt3edUe4etFL996rJTtrzQ3plcjLR9jDurONVZQCP
g5fRVHITlUTrccxGPsT6eqx/SWj8BlQBV4uX1AYyK+wrVGl3UNh1mURYxX+LOCbtbQwIxY5hKGNU
NpJHuIaeet+2wYmoh73FJfoy6uYdE+PdLDRXhoCsf5TcTIwrwLiZ86AQCZ5MqE0yGxG44rRA0NFV
NyDhTIY71LydMJGNkASjMY1ji5Ras+63jzKg6eVb3ckOWa7I3JJtfv9X1R5t8npU7nKbMMdJVha3
9TbGegHVKCNdYlppk5DdGqKsZ2aeQ3jNOoCybi2hj73U60o06Opiubc4LhgGaBOh1zka2WcZin53
2Vh8J2OCKPSGexq0HWV5kTuCHnDsJ0Urt9qlXQcvFV8fbVqctTfSQ0Jkt3/FjIMPrDSmDxgeJ/ru
ttETIVE5THoH8DXb5fFRZh8xhsEBv9Fvy9VxWYqzAV95xeYyCkcELZvZK0rzB+vW77Ynd+OL1I1N
si6RO9tY50wOVewjjr8WsozaG9wFJ/QDjVD6bcO6iAiapkT5t3hwq7rsd5gnXQT9NhE9eES9rXUd
31bHpGRrgxweOfGPUQ9BezWwKg2GfIih09xr1A47fiw/4+Q5mmsJTmQ19eXIL/0dWZoSR8rfiF+E
NGc3Z5zu1jjsuS4u87mpNlEeUyCO5FP9gCtMOz3uoFvZq2vSZLBvsRjxO/vNKZEY9MmZr2MOBY0L
Hgftefvj2icXxxRD0GcWq5/EEvO7JpdChkoAjHtGl8NKI97XSME+fgX21vE2DYoSQmTwO6N3nbq1
u35sE/zSNRjlvr/L6On9FZpHA+oP+yDbBXVSH+WvfiFMBpLfB34A4UyaFY/AhPcae8Krf4bKgarr
T4iPwuVxyoC3SC/Ly2opwVEnr8KXXfaJSyWF2u3cbtyEkte+HKwY9Hr/t9WpTofjyEHoTK88fvpz
YnkHn4U8y9yd6IBpZHaS+nLqvLE0FkMl4qUyIlWIGK8XE1hhwtBw7l/6lU60rifvczugIZmZPIfp
7ImeCG3XSmI2M6/4INenkWilcj4O/zeJC7djNTWIItBShOhxwKclbJF+DXiCme4yPbDLY3cWt7fC
HGC4ftOuMToquievfABgj3qs/dLn9DAlC8Y44TagsSx9/pExt9Upai1ZMzU2h19EohvgTgwZeKVS
78GOsEr18XwoiY8wwhhckAOZuHECCmnPBSUaSCioCzmDZlaTQJ06IiDt+gzsj6cW7xIZnfTnXwPt
JDDBpwshF1ByrhH5k0Zfft69bYVa5XrXQqziLG573qABFlLNr06u4/gKeIAHNAmJOuMwYEy+eRkq
BINpyoX6YI0QMOwMFoJuMKQjdvvw4FQFBemCD23rac7RTbZZ/1Tf8TBgfMluGTwzOz6LZEOWEL97
pmAXYQ/jg9qgHbXCxuEx99aXfNgmPr07IrSl44t3LPd1/r/O59WhvKEPX41kfWjwJFqgzKaQkcFB
rf7B7QqNm11fLNfH8LIc72PLITp24ZF+UK5bglcqXOHhU9oJF7AexOQYQBjZWNjPvRxs7SKaqjFs
H8/LqIBnNdR7tUfaw9fYRRUXHyjiuaRtKBYRMv64lcYj6Cf19bpvYi2fU81VcgcWNpALgZsrlfHp
eJrTm+y1q8AZBUs+csmo+zgriip7sTQD8zcifMPviDvzgNlE6VDjME+SzKYE4NxPTH7X8LBhsggm
zftcpd6oeQQM1FmQoA1MXW1y8vFARtV7K0EnPX37q8znGiFwPP64uzEASU4C5s0VsZ2OdFejH91p
ctsoVqoG9s5apquOGsCST/zrL31V55ZzAitUA6ANg5fDmVqSpnonkBUT4NArclRmZyXXvb3rZPVn
bL7H9GmuP8+kH1rJ0MscXVnGcWLy49A8deeXKK+Mp3z7O/Yr5zOEbDVC8KlXnbjLuqsNGXhfAWP/
knxCUan83ErUcQo8k+b+8RFMVhbGs6s440XUsr0TfWD5iJ/embPQ/+5zUmWMzanFbQBgpMFj4I9p
XG/XFrFt3CTwq/4RSQbyU1fyyEz8dUWbyROgFAcucqzT2krgdhqyG1Cl27w0/cdnCDN9u0tCgaCm
7+YcO7nZm+WtokHmvJ2MP8TNHZTd6c3wbDFcaR2ur7P3U8j689TvbbE5wwGfjdVasdHstoAclaMA
w3Xj7/H6SEFj0FjLbUgSlPfiMaEz3769ycp9EJ2oeIvFMtKqsUYa91iyaN7y7aU+JVGDp65TIq94
DBPD+yfPvSvKc0km+GXAbpWq5hzROoNBTBZ4yWZKmpdpWYPeZ6xDkqU2zoi6WKT+jjpxdvGg2A+l
WGDYEc0e3egExAarANDN1kIEpd6NsUeqIgy+VFg7pRsq25Wwem6QWFFYxLtuyhm/45zr/I6RamYn
ifZrjBo0asp+Yz1iMBYtpAmvh5aZBLOL8llDerJrcDjDhKYFvSsNFCl9AMU8n5Gq+//xGlhHdhiq
B/MAG9QweFyb+pgFu/gj2m27X9TjtX5ej5i+LV8UEshL68HF+h7t8Fzwsk5uIR0qSDlJyVOMAah9
LPB7w52yLUwfBCkDRs6+LylPuglRKSR84N4Oq/uiqouPSTU22d8tgURMoVGW6vMkkFWtK1BjMXYx
A3mVPnHIJA9W6NZiEtHlOnHeiKo56L9nX40KMJW92NOde8wOhtpnWUwlT7THmtiWnCrQBXJTvSCH
vBZicX17Zb0prkw1Rjq60HzaHZ1zaDsCDqbET71p+Dr6M/2PsO2tkfeJsPIuxoHY6WrDfcl6hh0B
32BbmP0RaXm2Lh4RT4mQu2zOBk0fxKGlqjZ+FIu5hWbYEyO3+yy8Bspu+hsW9jicLkzkbk0RY3CN
Ubk5mQ9vo8SzaGWwurz3nOxS4ncXfFNaj7jSfqLIZjuAHm4UY5hv82q7fXmY/F4JLp8TM+CzaPzM
8RIkCrJ+lRn83eFKne9i8Ev3zY+dTJeY8NGN5iizT9LybIpe1TiGo7t4zif3e4JPF/C1D3dkEhcq
4D0F+h8G2QEhDSiMlS1x7/DvS11t1iy9O7TnTKTyNwXFQJnAQSpJ4ehlKRYHJftXdN02Sf1Sx2Bs
dJ7XiniGFLDL3Wzk6y54Zv8bfinji1Zo+hgkdjykPSDe7szrS7F5DUEEk+ariHo4XaXeh/hH5umO
hcfRcJxM7PTE69Edug5O1bUrwL9/uytZeQ/WHhRPC1dHd47zHUKsokYv5GZ0x+OvUtB4GG6DiXWr
UNsgTC/MUJ1Gcs+cbLEDZ8b0dw2iAzGxaRofGZ0mUJAfDXBG/7msmLgzI3xqTXkH+4+UYTUPeWwC
NsBzoUN1zdNPzdMRMY6IqqoMV0LXfjVJ2Q9gP/LAAxE9bPZmcTFWFmDi9N1ECHPdS3ExWOAe++nz
11n2RLSDJ5W7GiEcWEJZ6jRiU46kDCAp32VsBM0WF5r2q9HSW+EOP0jUM+FIZhpT1oSOWLIaqAKg
BXIk+WZkJj/KDEGoqj1kAaWkn3bWCSwOBtcuAFpM7r1RpZoSFnJyMNw3E+A+AcKufbXzZPccPtDH
VTUnbd12Pi1eL8fmk58os8NTeWvcmVPT3AQAoRN33Gt0ppMAG0FnqUOMgk63lTJLdk+qn+G2kQbD
xdpKsOmtdCuGm5ikBjc2pWe6s9ZAsE3A1Or0RpFCMvH6S3WfRmHjTPVGrZophHFWuS1HIMjyE0Ec
SU917G2bN0DN8E39rzE6TuJoGZWak0IPs4GkUEPgkBcE1rrK1AXQ3ytt8lx0iYx5iMgxAc7xzSjl
zPNCCXd+MIzgrKb7s9h8IfzfR3yUaIZ85r1tRssmumronPuqZVDrHIppWVCqLguQD4Kob0CbMbyX
UhBufJ/7RXkTfiv8X7NQ9DuJQ/qqTMUi/piObkieCLFLM7SrYJBFkTSv2lR8TQxlB4lemJ2XdzV1
rQYyftdyi0+LPbeZYOdtlRT1Qqozs/Qlpx9PFn3jpFbuCmeYhrcGnS1ph69E+nod/vXH3D/tovRa
gUzC5g3qnRxta3DqcYLUcLWAYjXlx4EeJ2IT4B/tAdpjtF2jEVgiKoGQ8dSW2UNAuz0gMYew8hgX
jkHb/RsWhDukrR6lVJVEpR5n3LYzhkQSKTMklTiIgQJW/PjvsIaoggQWob0HO3HySNd/y5S2Yj7u
HnboZuUe+3WnxLgV1oGf6nltp7BrMK096wFEtyQnIRg4zvoXvet3Mlwysa1QWedJcm0mqur9jjrp
E+5Hl+0V34g3Ibmw1o5/olioSevbHqU8g6KM+lixaXweLa5HAnNJF32Ysvd13kJWgfDL/EyVY1JL
QtRshiyLTXcPZLVyKJYHMwyewajpMwLB4I2Pk+2MIr2D15X6sHbP1g8mNpn7l2ejb08NYuj36IRe
NDPVgfM5yKk5GL86vr4ZzeaeqaVwJ522otzNWjdNScEt5hGwv7WyC4VtG2U2FEB21jaAuFSN0JDD
7E/yzC1GEB3+APlSQPK5+5UrzSk375Y3Xwc3qAsJvozaPCUFhCwsyo3vUuleIusAEiB7783SPbag
2nl157cjThQm5KYjulPSJXRgaF0fkGXfpZxWJ3zMVWfergSrkLWOMQifQGQt8jRSN4oRJXBUKFER
dB0m+l/UC+xo8438Qe9EqlUz1PGhoPgDZnUC+SMX3Ka5I+yPedKPqwFsTzxgQr15kgvxxvuiR3Mj
N5pZPhpHKhpb3XOoAxRjKF8JdpL0vSvtiPhWsz7YAJ6xBuIDwxe+iPYxigvAsI/MeH1JMd5NsXAz
JaPN8QhdwZZEE3MONNAku8T1HAVKwuuXSB+ARKUOt3fIwCSqVGW2TtlkbWMvahUJ7R+ZtMLR7fON
9tBhAfBN202xRavzCmGoGer9/X1UWuq5LmZc8WOlmyfN9lmsXQ6syS4MttC7j1i2qUfsSvKlOE7A
2ONER8PzE8I38P+R9Z5bUDCOVNSbTFwS3mJ/p7cT7m/nwsjA8AflW95hMW0VhwlSjixIul1wR2L9
ak+Pmco329I1dHj9IawdP4HmNngT4pvTKSDBaRnndiQTLcFa1X+SoI6j02mCIm9kVAB2FVc3P90D
9H/es6NItgbB727ISzWb9uyJArfBHTK7kBRINeb1gGS3DQpwPvQ+Tt5gbdNnb6botbwtP2vX+/aA
bIXPzfSgafMEQGGc/WOIrZA8UzV9BfedVDNmHWf630fmSGSNRo5yRq7GQc/ZLXIH0Cpj/yJiT3KB
aa69hMx/eY9St138xJR3b27gCJ4MT1Ltkl32WlkkoN0OwqJIRvfu4dybNUELRbDJ3hZAmWGIo2iL
YKIZ6cO/CUzP6ZYJ801KecetUWnomQWxG59jxkwcJFM65BXa+pYo+62ltfnaW6NjYKm5SV0ogzjU
yE4x3/i/3Wuv7ROgeIjGIHlIKtTBIv9mijiLSmfMEnxS2mS5kO/OWW7zqs+K4Jla9GRDf2ZYIbu6
4NS0pM/+iY431kVbFpsPnJezZB83KTHwVfPaIabNyY8FkitydcbbCnJa+ZiOESmS6m3R0/9L71TH
KkS2iCGkAbwfdqOmmMOT6FeRLt6zTqwCHFxbMjeVtWw37r1RSe1uVpzSofGSqQ5pY829g1J7tgDb
Kpkcx7QXjCvMW8fT2vH+u8SmtTuFj0B0HGExsGUjdNxP66phKy7KinbyJOaHZEXS5jlwjUIyEfSG
dlCyFBwMOtIB7Fe3VfysQtonYFMxe/7+TK+8wCkZ0BFjptaYpVyNnOEqsa51uT4jzkbz+f64FPPb
XL+B6dau9FGBGjnh6NSI4XpYANOTLaAxTRyMxjioDn46YyvrPq7eOSIPBHrHnDDEzByoWY2Sl4GG
F7w5xyLrwFD8f1XYvJ4WX9DDO8AUn9aTzssltcnWdHhb5dwJuUnpFes/MddgMRW+TVjPqEBYJgNf
x6OLDmsuxY9cNEZ/wmOC473ODLV22OMHgBaFdN36goJgljJMJpeb7DyhpI89em/OV5fFfFVGHj2w
L32QEtw7WSZU1r63tsfb5epgdAOYccH5Sx3bRWkz1W0jU9qSbJFshY+ZILE0D2QSzGu4PoKNcYkI
xSa9n4wds6Mwryj1bPp4QhW49IBYP191PYUjGPUcfVnrBnMPOyQKtcC6lBqtX2AOZS/mNv4H+oAq
o1EIfJ+XfEozNlKkKu805108ul9AO8VIUl6CryIe8VKJA1i17qbpjP0vuYO5CsJs/OlF/3OPEeYm
PrrX007dLDfwxhd4l1G0laA1sr28w4tA3BElwFQvrvqMdEUbacZuQqGkA/2feRae2Fxvfn587W0W
eBg2Cqf3/Nb9BNOVRBVrckimV2KLi62lNq/AqkBLJlwB9t8ysfhr1AZACPe20BU9eSJ56qDWSBWY
rbzoOBwV4FNP3SrfECp6OOsG70+bYkAYAChjkJGO4iov0aee6Ze11q1VoOtuqLK/L83mleLvb3+m
UNDhrKfiCWGtqrCdU7KealHlk97y+KYmHWsh6dCRo2YkNanHq82LaWAkWHqrnRk/Pe656AlpJ1Cn
nxfDp9RWm5jOiuMsAE/ytvsTJn6WNvEMOfr87wgDC/ZOfBAYTq9/Nu7MwHTWuvImK1o0FsjrSLyc
jYXJMxRnw7dXETrNegQiProgkEAgoZMl6bbqCgbLK9mH7V49L5ey0wSHLworA1kVhz+oJ0M3NsyG
+pWiEgRSHbUI1nP5eC7zbdDKaWZyQG/N9iAKEyrV6O42j8/5V4tCgsJUgi9sRpFUs90YryuPXWH6
lcyvnhknNQIWgXjpPKuTgJ9vZXlovsKRwhxa5tr2mZ5T6iUX9FshytpP4jSnp3MpNq/VKymJt1l/
9qsaJJzFybtXU835kz4G6jFvozMkk0ypoQg6B5yup/N+SXF5oILV+60aBgtZ3QxdsqkRyeW9egpr
kuYCMKi5SONgEVoV/t0MUc2N5GKQJ6Ki7xjTcZXeyv3Ce1lxReUjctzJWXx3FZ0D6LCxBPIcUezd
/GGsfvIRCWPLA+7cZ+c48+yITbfAZlDRPSPX5kVAAws6GSDlWhdpfDEoIedDldS3CIGPqJuhkIaV
ta8Kb/z+dUKfFwuvcv8BM8qPcSzdgelpHuUzbeaiSq+ae2SnAqm1j0yE6yzqWEMq8+wq5XGW+oFy
B9rV2vmfQ6dpul6cccbnpLIc8pG253ehTzmY5GC3HQGmPKdpMEtBJABIsplO9qKNl1GfpbkyoIhQ
H5Bwfymij6OSGdHovX+eA82BXQgLaEmVBzVN2FOVwDpYEYgaExUUYZh/gNO8WuKVa7gGRyXvd/+7
xp1+RYNeWGaqGlL8I/FrIyBgz68gPf2pV2740oI2ZdJkulNW5JJxuueg+vr65hpv/jTlXxPCPv0u
tl5aKU+jtRYTUEBEneKSVGVLc/fV5m8ihN5GWmHv/e6rR2Gp+7ID8nlM/JVZkuctIVrk9bG289oy
Q4TozHbZahEiDQ1YdUFNIIMHT1dwzeOHiSzXHdY6i6BKm0nFumXM3r2TeMU/Lk2qIdfONcle6bMA
ShBubbdpXADfDqkyci1yqc9T+XIuoVODrf1IwkibhSVLK2ujG86cd6jb5eg5q8jVmgyoCF1l8gZt
QuxKGTKKHAJ2ktfLm4di0Z2WB4QybN4gv7YNsVPVrRLBxUdWdniiKXR7g4xufR5xQ3IxGP/RMH7T
JDs3Vm1DRAyRKNLXfJCLh9y2HLnKgJsHXV+OFlvKcij927c6vSvetGgkvsHrWed9INFX6plUbU1v
h/YxdIvCVKcDy6JlmSYPJnAbwFw9A5hbw8fYSRnAkbcprE62iQBKw/ki18+Yc+iivhVRDhv557aD
wfF7CHyvQdZarNbn2t53+8tLKriDjnQ4XQmx/H9BOHNW7xFVIRtpiqNgjl/CzBUu+3yr8f/CMmzp
hM82gVqQ1Yz2qhrIhx44FdHdybJAQC5XbKVtMHiDH6ecTxVMSqoDCgrL/qVZN4R3Al/VktCPhmZm
vebvmsXtFgjsO6FS7I5eQJUX22cKcTMqeOKE6qaEkAxVPRdN6PNDbRgIAtsDh3xSM694qfDHpXYP
BMROTzeVzMVTZMHRIkvSsARYQM76SKS6UkWF+wX6eTtLtm41ZLJwtBGCS28x8bA48zoR5x4+2nIu
NndOt21N2yvFQzQIl1NoiCThAOvcu//+vdgXbThEPgcPyhpCT6hC3XXz9ErGf3IKlJvN+3PxswAw
1/hJQ0MqnsxI3/jUN39QMMg5hNGPF1C40goJ3oezibhSCZrPx8bFK7rfZrBizogKLGk5XWy4UICm
N/hAZKbjhiVbKMq2DkmIO86sRkZ9BcImKZvsIUYRJK1ayqEIJj9QDIT8w8uUPFXGOebEkjLmEVF1
6Lv5oc36CZi3Qeu96wcO0B50tbh+2hJ9Xo/4dxMWCIeqODGzblXZruNWXVM3otvc239iO5biVITw
6yn4vR1gK6DGWmVL1FtmZ8oIbLR/4G7f8nJG1XBaxU8CbGUF6jSjtoNLiTBjqMVlY7lA0SmSaCE5
kw3dtsYhjKdVuwcHcJu2EfZ4QPyWRAquf+5MOZOWA14B3Ie4FiydirKY9lyZR5gt4ImtOThNb82r
Y7GT61aTnQ5PUaGhKNAAFE7Hw4IbildbzSDJjMjhtb8FMxSJeKe8SCr759NdTNXnWiH676SntUdj
inG+Ut6x5fkF/aUSaZfS7Lq0IYotG5/JCphIhQWAl76hbi6NGjDN39JOzS/WCPOy+3Q429wDCiiG
W+eRLSUPdkn3UpSd/mH0P1g9cDG+HYIQ3HpDkN1vKVIJogSB00HmEqNxo1bcEPdeamLxQWHFa5UR
4VxD5PZ3aPn1tjS17yEGE4ZDKOlYvvmdB92+5EInZipsa94pSQVBM3nYDT3EKCulEcEt8G7i8rsC
IWLVN4d21+9EcydPFzThgDQ8uedzevV9zySnMLH4vlyNQ0AzmCEMfrsHceA2j1J+chao8BeDNzKn
H+tmf+eJs4HLoWcfS3SYzv8DAd9sP7HG4D/VYXxXQUFgGiTIp3NJDPvwmzzuvRJEZM5g2yCPRNya
EuZ/sIZ+TnwWe+foFbvRNmJD79UO514hrVwbLNKj/7ZYjqKh09pPHsSnQpcupkpt2vr46cKmu2xz
lBAoslT8bnRW2VcQ05pM6ZEPCXNq1SOkU+67GyzJXkdrur2Z51dQMNSV4yCVdcuRH3YSkafOpQzy
x6blijlc701jwIYE6z7CyJiWeD+Dg3qzXWAYrHuhSYnPmHRP1Bw4AmHiPDFVAwj+mO+zjYvxW5sa
jLNuLN9W6n+p/TzE1QvRyimd+PONTS2m//eBWjHgdzYO0kpjP9BZoM1gs7lTFZeDiNhUIGDFn1W0
NM/YO32NUzhOES4tvdy0fXbHp3xsF7EFvQ11nZf4bfM5RbkXPXqWLqzfh9CvYL0bEITIgHaIu9Uu
EFVWrZdKtrWijwqsj6joGNMKZQ4h+k5GmTRyNjpVXzN9DklW8NxCGjSqQkvY2ILcsf3suoG7qmbv
clXJatkoQIkM6alTel9QLJ+EgloX3fvCEB+1axnfw9C6EkfKElO4IMcm9vcpaSFCndXA9+etL2ab
F6TpmQdegrTdnMChiHEo2UyZE7lB5BzDWBrwMfYJ+ezmZLcohS73KUq6luE5b4td22RZf7FzG2av
N1BH8R6bRHgU3zC9kQ8CD0kMy/zZCuFsbi7v0oXmn9RGKQv17ylGZxXUMEJTWouyAFePlp149QPf
3UovG/DYgUJLTH6iIPv5uUSdsTeLU9oZe7o6drU/miWaYVKAOTJ4mQlnIhpNbE9rVTxbPcdeRD2H
0/ZJRJZEtFf+jgAXByrZxMHACb9Pw6m1RQ6yBU6uJhoTfoeBMCL+p3InIjvda54S8Pcco2qCiMr7
FOIk2h03fCKZLfZ/ebNb/xL8GEDv4aZGZ5K5RIHwE2xET1q3HxSz6dasX8eYgaYHK5utAxZ3FU7n
HTLDVI1buA2P22XoQD+UHpZNbFXN0CIzva4Bukbz1vI6+eJJDjmSUaM6JFGRjET25HDIEj4JA6Ef
rjf9PmdXmWJ1izfqqINtMpih8noCkXzj49sU2/uI/xjTH3teKiTqjSNAqTki94YtQG+8L6sRon0j
L2T8cz0TkXZ3iidhXqBPaiuZBKXBW+j8+486q6WcYunemVXCY7WHMS59FZU9awcX/nEjf00lUG0I
PSSbAMmUrqwzaezbv8OGKhgT50PaNv2mVO6xJOt+pAhRXEP3Ff9zUD8C7BZKnzfAmw98IRLCS5tB
JRnV7MXSTItelfn3/FWK13ArySJL+zXz8MGU8WZRa6dQLayabSqH1Y9Vo+JIC0B9vcVM/8Y4PmeZ
YpQ02q/xbhtSDNomr6FSMrRN4nLUoaWgvJ1J0qBIwxkjBBIHtaA6r8hFT9x6OLEMSP3uQv3uHLk6
4nYCU9v93KRk8P+lh/4nCnEjCubvdc5zGlmEBucdXOHTZV9n/ppXFEFeqLjX3Nyo+QyjKbE0mFkc
2iwguwOju2e0JbXFcnumnXn80AtQNqFtsLB1Y+eO2dlvlUoJbZjfXQMAikzjfox6nFQNyF00A3ap
cqF6BIgYpiWeOSqxCKjAjJ6bSO0DGvSLRY6OKgjSEiLtncglgFc7ucA+lxxoLUlDcAjOzT2GX5dL
XUtRvk/LMCxPRSSZ4vd070QTn6I9XgNO3bE+2COT7L9Q23asuv6x+LUY7QGXZyxDP7YfZj7TxjH3
Gd1JcSkqoUDl21qo4qWu3JWom+Dkt8OwHxDena3oSEQ8SVoGxBDZUDMbwqdfCIkiHddATR0VRCJe
kmseGF3LCz4WsRHOiDsDAVifUX2dUWZqj7gmL44Zl6PpjS3zKMZDkglWjbPHhtIjBXo8DOp6ikMW
bPzjQdHQjGUAtSCM8UxIBK0UV5eax9NM2qh0e2+YGSAo+5hgJbjo+SfqbWeh8LyqFTqKj8gr5RJF
6+GutpptbZKBP9cmoHpp14Om+8H5cYbAtbdrrJsuMJfkCnW/P3iyPpJXhNd/NWuenf11u6FawKVg
8cJQKr1yXtx2JXKq7WxOXY+4JCUkomgQtD8Wie6DJeD20z3qJaVBXBD9InH1yqjdIoo9m47z51di
Da5YvkzZ5x69DpftqYOUC0DYAR1Ii7SNJFuk3sG+XDmBvPQF6J/SKqi3o20DoXm6dCy4AGwAwpRk
nM0Ub1D3G73wlfseIh6oUm+y0ODHi9HTLSiy4ap9YCNvptcCOwtjKdqfFQvYSxSaspiMuwmLoo3g
+iz5ZFTf+zmIxGz0u9AitAy7Ab/l0jwQAD0vqzLh2ISkVH1rmqf618dcBQt3In7nXKdpseQUEomH
K6+Wu8Aj8+GYe2BGYcT0OV5t2CDufeqE0tOyCpypmLa5KA6XFyJmqmMQqweFDtOf08QxF9ZBXnw6
HyTU3WjwSac8SYL1EPavl475a0ZP6ag/NhdIDbNb1KqylCzTKJpoTN/BDAoBRvpJDBLxC4XLAqx4
CtRAukn2sqzCnzHS3P2Rz82yQPvqLptuziP7bv2BXWCOFKwlNKTD4aeqGcpRbPy9IoT+S34EVWT1
1ajUV8zHfLCeZafVHVvaf/yw4TEOhNLm9CNqFWhZmRGpThdPR4QagCTJzHYFXBN1CiwsDPU4ZY+8
CbVCrWVAC2mpXtJRplUtHlCkF3R1UoYm4+1XE4HQFV6b0wa9CZRcg1kHsb7h7CA6cQFtr284gGbk
lQhs6VIOUjbSiNi18Dr/R3eRUDc/3Cbb2SBoWby7HXXsIIDAdoeUgskOxCzLQFNgt9dUBVvPhnyo
eOweYhiyubT3uopSu3sW0gvZELtkJ+2JwqZ+P8Uy0OCgrFZz6NRFAYJG5hgYfZcA/1HEUYqqeqNO
oCzx4j0Uwjl4ZEkRbQrUvu+HjaZkGDsbqmoP2p8gIvaO2DbjeNBQMLODOc38LNqmwruyJ6fLVQoE
hsJYEq0lSOUUSKBNPRZwlxRUeipy9p0r89DalmgEJi3Pmt2KqKoWpajRzAfC+ilzTTyik53KpiH9
C1tFk044jZabjIAUMwCdWRAfKQEsm6GKimH09waJSQvdyqe4L7nwn9mOflOHfXOh8cDgGZjwEsFR
sV8KvG60ItkDPtNtQYZtroq0ouw33kkUXqV1Bzf09pe7mbheGUGXJdHm871r9CZri/ztYMDFenR9
+1b6Gpe8aGvonYmhkwzFsZlhbEwrRs2App9/igsfhSVoUMUqxzTmuyxt5pIB17N2atZ5/xKPL5Ux
CM1DucTqKG6OJ64NjwXBz3HLmGKziN8TmM3PHFJl8pZitqLQz6vcQgiO3tHQV4HOnY+0PepoJxq/
BxdgZrOKqBdA0utO3xVFqUwpLtoum5FXbyDWNyOJ+ClUcpKHxceqX+aPBxrtEXLlLXzWdnoT76bk
JoXNl294rIUI5H345K0rT3AOwnq1A8S7DK/nrkYIACbmN/X9//yOKT9im16P6biJdoRSZnx8ijtU
QI1yWa17VqEoZWLOO1C64Hfq7AdwKyjClkruSHgfbaLvQ8+GJC7J/v/1Cf4TY4JcyFlZw3URYi+v
2WpFG/5oFQhkdFzkfFVrO0S2ABR6fKtN0ZsVgzBk66DGIz/jg7o6A2XGTeZiu3aJHY+aKKG1oO1y
7EYEUfTPlLR5cu2HRYLpcTqI2AK6CMqY9vrRoASUHron/gO/Vfkh6oO/PgjO49ewSbvffj42T//x
NvxYz7kF4nav8EcIExvS7fPsuqrqPGP4xdY6Dp/ROf9gBdif6H/tqm34YMzN79B6iQczHNpv57nv
Y6KjKRE4kmxjUOSw2LWLaUliyxZQEWxqAzeSiIEWEyEmj3P2W3Oo+YRqh2hIezQ76HIxW4MLnA82
VpwzOQvHb0O+OXHLrnmULZRCqGWIFQND44YsI4VIwd5GyvnBZ4I4th61/WPLkz5FUyDCHO9awS0v
1HA0RMAUUgzth5k0W2hy/cccUNL+/ADpNwGylqr8WLLyTXAcRkJprFQGq3h127WxErGFDG8tJiPr
cfTKFO3n3JT/6X1WLk6b6G4LZRNwdM+fpH65gFn5VTFCARg2CpI+LWCaIQFBhEIGt0/4rJppUVDN
TcrDuOfi/98zpBHXPfDhkxlKqSftUEjM7HCkTQcbGdf1GZsa5a9vHHaKX1ta9Lik7pRPTiLsA30d
sgB9FI6UavhMZk1FBRJNYreUshW003Dq9SulmXFXPACSYBQtT1kBIT251cshqs/6xbQbPm6q6uqp
J8y1pFH+Qi6NJeUhejpV/mUBLqOMHSNMHaMW5oGVIxJafa2rQRhcLsb/a/GZIWtCKcER8FwwgC+p
1V6+MrMMb1cNFJOFuHMjVgzWbVw7DDWBezIDOU87/SCc5teSjpFND9qL/H37pELG2QbjJQl6iYle
CpvDF/K+PhrBJlOonSO5o/U75tWPtzVEgbZnb/gtmqO5JoT3cz3lAXer098imeVEjznSlQTZLkzF
cQjq48CRZpqjEpjlkJ5VSOIcfEmX1CYNx9yXDtDyz9dDsrKYw0hyz6TY1PlW3r86KC2yKPKh6KkC
eyDMA+2ruv7ACXEzp6JkZTV1JG6lKnsp3t/1U11UuM/IIY0uxyOONiCbc59im0c0FC+yPzQ00RS4
UjjWdvvEvHNuUbPq900pf9BN0a1smWtG+CgyNHMEZYMVvcE9YZoSJQNnQcsdat2xENP0FTQJQFB5
gExTUo324eryK7ua3ikQypjlysV50L3R07OPZrjILEZAt7xdl2+tP/pCxWUbhE7u4V/TMrfTfApa
U0uw/d4l6/Qe6qCKrMHb1ztwfqMCFFYoywPby7QpF/E/xhdf9TZkJevpNKk7X+y2ZQ/Uubug0kBC
2jHqKzxtZJcxsPiEsM8xGI2y2FJtCS+0mwbm7hJ3V/7BxEpVvSMUJnNfXd4gEnAqTIy/IkAvKk0R
xcVVvvIS7LhQkoWHuOkpFDYdq+zHYX05y89o6NIC680ahiNLSp+CjTWGrykerY1GlKSE3SPKz52P
RaRKMRJUl0aJhGAimP6CHWSw7W159L2F40KzsDb9cpwfQHGmDnTZfqOVEYCv+YVYHCydI6sG+egO
dW4Bk0iiEuSwxolo3fcIo9oTXEsGbpLt0505MkacmXqJ928Llc3OxT15acNyo5Le0ot5yrvjpVXL
/uIg7StVrMMMxDpmPE4BgroQ4l1CxHF8HX2cUsJOFdaim0xfDBr6aTpjcABVifjTboQBWTMHYt+O
J7alNmLL2TffJHys1OnBE/gpSBh9I7MXdw6r1vhY416QgwXejP2tbdR50wZ9RwSrPENA5L57KB4Q
WMaJS1QA0sgWG/FUlbzhkuD8t+FjwKeeAcMf7LIKWW4cvPEfUdidO/cnPVJUnJAAxervPImwL59a
a6QJp6y/qsCw+QOvAtcwTxda3e+mCUwJiCFRGduOzLBAotcgbibQT0jgFDk1oqJxfpOe9M7MP5bm
rt+7X+hDZXbXSykmqJ71MTRwNHqW2wExi6QfltLdLCElGVn4xjaefIi36rtt9uz4catNVJbz9zWo
6B0Ex3tHKAMbmohdUc6T6IYsIoto0D6YbbX5T5iSdNc8Wq/uFwIfhE09p+wTY86dne9t7VyFj+49
8XfU1qC8irABNdEcUZZd2cz0YEHBBQGApHZuMDhKUq062SnTF3XiJOARbNAv4fl7cSjtB8TVZ8lU
3sTQe9FcgTgHWICiHolvAZisD40q5qK0GiBCt2UpxCwrfJLJ23/gDVpcaM9c31A5FE2mFzZqsVv/
b0VfIxv1EBmGLyziwm0+JzabZTO8R8vXli8xG8cHAA2pUW3FvSj7hMZTt+FPrLoNgY5TB/Fxnjxy
Es/sOAClmGp471P2BILHbicCAd5l/6X0LHPcODfnORAaV6PggPgM4sZM2LGq2M0q+lTNgDpI87Fv
H+sN4Kbci8mrJ2AhLMfQTHh413MqKbxgkYYojRGOV1eDDiC1SHEj7HaVS8+lNjQPagjpqVSfrBIq
5PyOnRkZFEBRo2LEZNvMsoL0p4KFxPsyVdm1W5w9GW2h2IXeniV90bI0Grm8jDTjKxThdTR8794V
vhBO7gAPrfLdgTih8Ddv2XoClUS64C5nAGr81TjdKXv6btQfEZhJWjEhwH27iB+EThiGZfBa/jFj
QWOhounhVM81lE2u1KKoEbiRsnTTGmxlOKyCBTJJT41PWCLTPJYjIV4o8zIuWxDjgty9erROU11s
zyCTPleVHKK06ot6jauBzGFnWHa3D1r+en5S8ep8AUtofpIJDqNNEgJUceI6yRO6h8mWcqxlgp7f
Gq0C7gQbcpwJjVf2y75J2LfEzyNlLgWDicIuNxjhtSlaP/Rn/lkDbNn3LB9MCGOHXTXew6xFDnFV
h1vkU8Z5j26QeI8AsC7/a4J6NyfNvro9TeSqJwMHnmw/NDfn1GvFgOQVMbXVFMp1iDi4GnWEJ6jy
9camJ9EG3cHgxeedHBZMMfJ0TFwq+3L0mmp//UMiLOJdTx3UAhc0tFSeVoqKEGI0jnvnFvv9ev+R
+3XxyZ8NzB8es7vt3x8+MlUCxujgQG8Qu8pksrEA8w0Z6xEykSIu8574p6I76qX/oabH6HupDX0q
GiINAMk39E4/mgB3n90hAsTGiZB41qMDEgKvh79ivq8dtEnVU5EtMH1xoupfKIpOd+wozmFhKGLE
sIWvU0xc9NsQEaj+riSSlQkZ7NECexZ+68G25Z46rnsRMtYJ9COee87Wr1iadltXwdiC1Zt1Lky4
UH5mCogjKJC5FsfP5j2h4mRlY2pPHTC3ChPtj02k0IQ4h9cP3v8dXTFKEfXdpRlz1yi4/UhWx9AL
cqGaWn0tzcQHVZDNECRw7DOz1dAx0kMufIBNA2741C9CwjRVTNUMMK8L6QfC6zz8EA2/srLxIUI8
JuExA4mlxv9uw4R3i4Z5H4E1Mui8W/G8TGpYKx9jQnN7sRg2/AylTImlZZ3T93CJiCxeb33RPJ0Y
Zab+g88lTsAsmNeniseKjhOaGcAfPZDwet+FisKTuO5D7qP/Mw2yl9wKEWFdOgh4b1EBzREEbNDz
OWCngVM8ZBkeX+vRjw2ENdrPDDou4akruMj/86R+h+MNUy0G54FtqH9MEtOhdmjbufQKs3vpgWaJ
r0ptHD4Liy9VH8Qea4ZtuqbkGjgl5KX5aQ2R36NdESq47F8hiAQ47PxT7HqS5gGXZZrBXNcyBqgq
pZtFy3iiFA8SqBDKgZmER3RkZmvXwtbL7YSwBZf82iR7JGU9hdPyeZ15g9yoN5Je441elafm5JqI
Z1Y2Mfoy+8Wuoqbqo0k8GMFEZzoxE/X+zqvBWrpH5+W7cFY7ZNDGiSLyZLNhMxh3RzaiLnTfBSzz
1NHuMvRfT1jnUsZT957D1+2sIxrtqlleUd9IscBDy+HfiZxRwAlo4djsA7TRk0nvSrHvAgBpRBfN
lE7kFz1LPWD5/d1hQ1in1zHuu/SAekt3uoAHhMAC52gxsYeM8QRs/6tmCMKLRojxc8fWILm8zcdt
0g0C2/HsY076qFxhNTjN5agj9lZ9PhHr5jrLrNsCmLCnEefuH3LHzEvAy0TDsfwvyCz1Q8bkbvRl
nuWppQA8vkLhPT0ayNZwGBjr5XPy4rbCgjtQIULGE5yXx7jAdrxOx5+n4MRMINq0owZ4p8MtagEV
CjH5TKcf2aOWGkEZackmlYax58fAqTiFqBnLRsvJxH54SmLxMboGUN9PBydKXRGL8VIgLZ6aiT2D
o1fGT0auN5CTneBF+fQU7kQldRp2g8m2yOV3KENiOGxjH9X6pb121Ch8/z6oI9pBwyyZH7CaOMDp
6dXEFq8YLtV1rDDOnCjj1o7vXRdR6aJP1U005SZvf6Oh3r//jPH39uNUK9KtFPWWEBYmnfT7oVpM
CPbSaoe8aGau31S6XcEUnLfR6YDqOIZHaBmIpGlsAiBKXqdatTYdyIfCm3cwGrFoJydaUpW/oAJp
yJtZll4gOUun41eestS/CJI4j9FNvP3GemiYyR1s5CP7Av5a2McR6fY5nJIwzx7ZNrmnQb0mun2J
Ev8OPlCH9UPZwpPPVbF3aRx/lV3oFlfXc3xq/o2U4mxTr1nB+Or6dKFPB/zavp1eLPUPWR6intRW
Nbl8QqWmy1M3Kg53ZfMf6DBVrwyc239JUQQjHzTQ++khPhR38wEf/XDv7Qw+LgL6VWIU1klRy1xg
2Gmt/omqasP20gCCboqwfhziPhFYnc+fdNfOygev5z827CGgEu0JxzLmS7mn3FK4R64gkbu9UAPa
5Kyc90hQi1LilSBcbqv5nFNfvmT3OQNAe4qCsjgEvoN95apJZfYKB3+eOM4wBBoIgqwteqZSV7Fv
e1bWJSP3NO1m3QRw7JdNOJrU6/enD7wxNlJaEPWNyhxNh2TysRk+VH5K4y+soplnVfrojmwRiqx4
wBF4MzizqJZCyroOKBb0rHjgXKJscEacPWP2Np8tWarzxWKQf3eUP2tyQNF0UX5hZq8tt1RlmZlT
jDF/JVguJRXAMJWG7e6KUQUDzhQAa/jy9X6ejSYVUkwXCPkbVcnLPI2ZqPJLbGid0X4aNPabOMnV
Rc3hRjcC0ZOC43Wxlpz0TIjy2jiS4KWIg0s4SH2wE2A/PgCSQkvNaRHRwM0eVSWyxL7udwQcJ6cn
W6KVQso4OX5bWnlD4+lfTcl9mMekdOzwbNen7nP1CcwVSW+nydN/6NqPjaFRH+vYTieW58g2KIpf
hSmlZLbMqVt59q/ahTu28B/pqsewrVy76AKIekl9OXg1crjjwUZ12m+VN4dDqSi/buh7UnHIaVbQ
lJtak4W6w0meMD/YddN7+EOQpzRlyfVSsKyMoa9lG1sHfUXe+5VvtGLz8xWAeae7r4T7cbfO93YI
7BEvZ+JtYmQuI9+Bpcy3BOUCSEJs9bCJjn7jLtUc+eHEv5LEyo2n9x2+h7fzGWd4Wb7vfBrGh4Ok
WBebQvMW0GWxJWX+jc/UCZtaVbdHG9QosqrnISY1Lm+uTg22BlB/e09YIZYx6OLnnTcrt2W92rR2
2zHzVNwHbat/C49rJv8BI2PsmmC6K74CKe7k0hJIp2tJqKNFzGKJbQHGv0T6xetFcTKWyqg9QLdz
RRgtbmmrrix6L6VhKkkh8yQQ/STXar90lADtpj5ywevELOCDrF+4F/+AxKn1BosKEtWojJVVtAfc
9dmOqiNQNPZmtYGEKeyS2tOBF2vJBVD3LI7SOR19cI4EazYyvkCO7wV6ULJQzRPOdHZkvsoqkBHU
UEOx6TaAMAYk/pnW2kii6Ct2N2nCtYNnYYC2DsZZy5dGhZmmowB1p8h12fjLWQYiVWPKy5+3QQyV
z35RXruetfm8XRKaz879oRKhQlFeK0lmvwHuVMbbNcBdf+pcY7ChWEZB+JGa/aIEi18qNxZmpLJI
m9271K/SZtQDkEKG9RvViVkObryAYCo9fqV6LEf7k5rq0kvHlIO4noIYjcyhBkSegOzB1FhYOqr+
r/LcDU6YpyMwPAfNWJkxocboKAevk+oGFZJpVaKaUpAT1eh07+KQtGNEpaws2GK3ORg+P4i/sUP5
UtpKnoZh+JYepc0XEwesq3ncvXNyyFUE1pipEv3DFlLPnqbNUrUWjLRdmVElfMxpAzRxOYOKhheG
mZtbyyagOoxmvZ3gByc6sF8wSRHfuNEdjp7YSxFblDcMcA3WBgovA7aeKLA/jLhvbqZdOCknAen9
prkNUERCsmXVzQks4FE3j1hVl9tgdIGO7uyZe8ERN4eg45bNG5x0UouDTRgz6+9UsA7tZLzkd1/O
MXoakxKbRTxo53l3p+VpjUyRmJjI0Oj5Yngum41fWmfHodEENAhXKXYvXDd0O+WfjXIs8cccs0n8
QnO+jQMeqtDRFtPS1hYgtQJpq/f4XrAK5t7nRsGMo3WAQ92wqAqXwrwfl1iIltiZC466keg8qcla
xrVZ58LPIRGALbvKrBIb37T5r/lQwhwdJuJiDNxczIknRGo3/HLLEsrh58wWlPhTfMR9AkFFLQi4
C48lsw0fCpgMYLx/aTMzWrol2BzIFy6qe8lahk7CHqZarbFxYPxOwPSYl3FJUBU9mY8m1gzec6yp
v83IOyXbbhFkwoN454Ch6S/A5qqu9hMJInOiDltTHrJKaWZOrNof/LV7LYv93ftYFSSMcta+cJgF
OUXRje25D5ypUGuNcKX4Tqjby6inPWJRllvjJTXi825cinJTYUW8zSwuDubyaRakLvFm0OyBIDe2
lw6R5gxLJXudDTAJrp9Es3kqRP21Fk2BKr/FRaZnpj/GhgNDCZTAVtoiD8fxZOXJRd2BFssWMoT9
6OvEbKyhhSovZXGzX4fD+71ztZcOVeZKb7xOb+GnKganMXcsLHhaEWLFv32OrEUqEys/jrwWRB3z
V+yFphaGk9J4QktSDi8EnIF5IXCZ6Nh51XeDnaMD8oS9FWzmbitrornRNngL83H6R8zyAb5qn/YP
dRNtBfKxtfNVxnxKMyyfrOlmDkSfBRUEGXlXGspryIyHsBArotVEt0Wb7jNGZl+SDP+igKWjfhen
hdbhpWTPVkZcwKjycnRJotplwtqvASf3h4qlVEIGHjVUu4kiFqja2pUO7TkQ71XxFqwG8/hHPz2o
fwADt3T0PHiHGzQhrXDWNLUmjUex4f16xVe+q5RcCVbVVajVco0SW41Vafc0yesuGbvPdSs18bx4
0ZsKIajZU4Z1S8kWavx/iBJ61LaS8BeKLXCKi0S/kOICaVDJ2HsBypYLgMk41dQJ0gIWgU5x3DrY
MOMehjxLy+qE9sIJ8tRb7RClubs0Ggn/FIgeREQQoFKSGNl3aavthxsoi1MqS32jQtnqK+cevWnn
RpJRaibVrSo5VnNqY+NzxSu1Uwp9fr5TtwzyyD+LE3RDXaw3A8FuWwfOYNY357IyOfn6jJv6bmt+
WhZ/KlPLQghaogiI6bExrH20FcjzzmldyHjRBNgD9zdtJGxrEMi59roO1Ta4G8C8WdiC23Hm60Qb
VocBwVzFgVy6NGRW6y53aP2Pxw/fBKkCaqzMRg0auUGTuUCxMzBpR+EiM8WlxqgkeFVhmCcZjtXl
jvT5HO7RBmj2KGT12liOtViYffVZw5Su+QgdMxDzuB9z4qDvR33DjsX1BYWbTVMx8rVELEUEBElD
XXooYXuugj6/EJWAn/X+zcsGElvmkrnookrTBwXvMopFFqztW4SpgdYzr3+MN2bqS3VRV66piDl8
5OnZJbs6gK5syJtJaiECOjSldxu6SUWfy89oLWYJ4Zi00qM0mJGWHaesVOQpQK/LL2ftUDm9D27I
NQDsYFMzBSL9pUhf2gLo1BgrSqgXmdewCZta9m4f1zZNRFDczBZ60F5KY1vlagf9MunnidGxHwJO
J0buiWB0316YRr2VCWYENPRfFBsqciq4R5UFViUS9EAbXO7SDFQZMjOh/9a1IhFEBFFzvN2CYDqT
pLbWzECkUx09Z9lQxqA0qofi03IritlxYOP7l1VNpsI5JYTUZNJysf5rFIbHEjjxc5aJytNGd72W
mXcSS6x5+Ii+ucwlSVCb6WGLTjkjXGhYQ+0d+2Dc0hKodqTU10KEjnqG3P5VMcNBwxxuIYdmCgWI
ZKt/ggn25/f82sXj14p9lOANrB0dfTfCcv6b70SNJVI0Hb3jBArzUjFUnhhURo4ZWpMJ/JdALxMp
w/G71vp4Cep8X1oJ2QRRmJLBrihdbQiyVUjOjl0QLq5qRw6tWRJg3JmQJs8gq7oUxDGiRr1E3o/E
cP7qUIm9Bz1w8O1pJwbg0lD57DATulVFbTPqgYVw64RVl8ih27Xu/oNa8WCrY7Vynoyc/SSelEVs
YS+NZjNIRbHMJkSfSEVAjTKDrUvlhqswQ4FBu6KR/QWSskG/5Uu16M7KkNBwQNbswTmULPsET+Q9
J9XEmsisB/kKXR28QGYl2zyoeSl93AfmCYRk2Wam9ZCnB21hbuvNN7XvAxTBa1eFpE1Ud6V2XJbl
2/qAvUGFBJgIwHvRCcfP9Hs62qKYxh1vd/ERJGagan7lHOr6xQdZV5ZuTMqhNg5VEGyC9N3QvaG8
B8uGHJ4mtICsNlz4XBpIvglF75KsATW1v1oUEtCn9iqtKWWMQ9dY5jW1IdM5bEUogCblvoRXRtO5
3ZcFQrJl2jDy2mO45sM7pp3TBsRvKScQKFfs2Ckcg5g7c0ndAJQrL5vcIIAC1X7cJ8CEAgGyUpRC
5kBwm486pghzZVLLAnN2cSdgDwEXFu/FGCVeuJ0IUGKdaR7GxAZyMFVY73RpEGy+U86NohD8Bq7v
X1iNyQrNnEhMk7DfJmRFZhpOl5g0oquukjuh1jMpVjiut9UgyqmDi4tjjNC+vfJ59c1h9rb9lZ/o
LEFerf8SsL2guAyY4ArQJZ3Zic25ns7AyoVEKJlQC0AsAR1i1LPSugwSYwCDdmg/wC00x7u+/hUy
Enfon5OPkREXikuYrdMWw00GbB6m083ecfPLZi3di8AHkkBkIDyoTCZRnXrlPFfB+CpU8Vp4Dt1l
rGUz/McP9Nm+b+eX8YJG1GtILplJ2zHAlbu6cCKPMCtUBaPHvoQOh85BKjerr0VIGN59VeP4KoYK
KbpRWbXVbNWsctbzguVMrK91WNDtIEOJLuOjFoDWXCzy82NSXyErTFwvA0PdaYdN77I0Cg5mB2r4
oo15ZJENWaO90d2zjEw/zcaofHmHSKcTHcnAInu24q2IiCmQRYmZ/VP3ZSl7wTF8FfdT1YYGozKM
pDozb4wtHYIg5PPQaEN3nBPXCtVj4GDQBU8lexj0K41M7Tz20EpSIJ69fMyyrJMfT3td341wX5ZC
/MFfnEq1IjtROFI96TVeu9eSCfSbUHvwYSjsuYNzBq57PeqAxto0bMuVN1DgTMw/ERBsfOAs/rWP
YDGO2W5LMMfdkDRSamUxfc710Qu9Kii30QHmAZfpg7heUExU8Avhf9ZfY2dzlrHOe31Re94FWynW
RVmP9mfAMXfnRe4jmMm+G9+5CTnNQ4gxljb7mTXCTzQrTx+m4Swl2gBrf30I8xmc3Adm5MZnmgH4
9w49rVmjaM2mwYK+p2VyMXYn7s9xPk5B4BKz+7DCQCZjiDliIFQpfF5KSMvNewYChcja1ZVbTQpQ
y1ZlY8uWQXkgBhNjZPZX95qwF7z5tmUPouoOXHUxUdYjL8tYBuyUBYxEbODXBsk40t0TjEr/svED
TkRgVAvvNVOO+FvdcFi4+yn2SRq4iL2tUIuvtDVSdPlhus6CNNK1gph52H/YVOrcICKnzQYExU8p
c56RUf1fbvtt2ohqlnSKaiMgyU92zYKlTnTzfn7shO7kkYPokCTgmFD+xMb12DbrDR9Y2OEaA0kU
fRFbm5fW2Q8o6tKZVbctYyIXK4l6jBBIS5O44MEneAkdvSHz0ZXx0KOx6JN6k9D7TwE4GnJ5xsr2
qWumfWYT1b7L6Ic5cxPnkic2+wafIdEMMRCWP74VByVf0bLXGUBnkP5CsjXCzk8wCSej/KpfbQcR
TdxsKszT22wx+lx0HG9UsBE7JnAQQHEGcbkRTFsqu6erYHGDy3b4WgcMxWbpbv20AMcyrpHyyD+6
ZwjlW05ZcgoebSsWlHxsFulT9eRtxBKhNy448MqVS6x9YeHXiAFgiKWv3Iv7QULhp/uljWTOS1Zo
7sL/sdiCXYWVJTv4tRnHeNfXj1FBJKKUg4MEFc5PosbK4M/Q2bGyU55uzqHijNlhQKamUACjcbcn
/1u82o2BGI3ceozse3rTihjoBNAep2jZowR+DEE7LnKaRYPky294UgRpYn5KSuqk2M8rxIMUSVl4
UIY9rz4kIDyLbhCPsH22d4kYDuqNdUVDJgaoLKtDPOVwP76gNf8tvxXEIfDsajdHBLAUFVX4eY6b
f4GtgRSX3Qok2IBiaeIUkAkmFr/jkwjisvwM3a9tuSkO8z18JZInqnTLYabK/JIYmmgqrRTVk0iX
NMeJSOyZ966bcCCYrbDwiCwe2El+6HjoGn68MhXFbufFduXse+7byubwnlTY3xsaYurcp/G3Mkor
eY4Ss/IQWUgaBrRUY6VXN/WAw83maFemfsa3nzbL/W0cdfD67jx9kpsUA+cNSlvxP/+kwuiQlLZM
HB+KuzNgJEf53d70Xn2dAd42nXRL/eZG3Kk7jPsL9WHDSszLJM9g9Ixp5U3WeUlvt96Qm5aJfNIB
0hPO+z3X2AnOEhVhq0blCzJERZmwvq2wqlEOxDQ6ASyvCU5H/ZGbn8dYoQUDVKbTT5SsYtbOAbJu
p/alzDubCrcKG3eH188v3kzByW4SzOl+S5FaXqm5AixzJQzeXL/cPjdRPHnRLpzv/W5/b2UoicMd
CnlXbOiOxsRyuIKwWP2kdoFpxF0ts37sE2n8Gyb+rOBY3/7IYbxWaFq3eaNNluQxVv8qWwjU/3YP
gTvY+v5XHvT/PleGKk+BeHK8hOtUeE9mpVn8mHDc6doHg5cUENKZydILRyE2zglJqc7t4b66aE5i
IU3IFGqN7fP21t8EbLKkbLir5Ppkf3iGvrXcJXyGNyK0J0zfrCXLdcw+H+qiA8iZlbQHG5JU7cqR
2hXDbAwvsKNGmd9hZc3lj0fpZ/Mvq7sRGRwDzf5PrL8El/TWJIuNpVMJTLJciiUA+Q61RrQExS+5
ECY6XLkfCD3BSXNl4yyTBL+3YMqsCpXAHOxpXwkv2in1ZsQgZsS7rSCHPD2FqBNXrOV3X4QnKVD6
HkG5PPauPANalyCslHwPa8BkAItq02YqsMKzAqpeu4CSHEdggNN6Dr2djVX+ZqRluGhJ9Ot7SM4b
EdJLHIGbPUvyvxrDySrzeKTSdjjHcYDnVLchqNSu92RV0XSCNKywpgsD2BkOiHVZrdWfUnunflm4
anl47tv1fujKi9WZwOTo9SOH//WsVqp+G6+se7rRt5fd6refEtRrueW5LbR5tt3gJzvpY2D7lF2R
SrqO2/ZMTmX07PjMA7zgxZuRs6I7iNiMinbOr6BRQPrJG2vkhPHwhP4UFPkthQLH7f9IhmgrQfDA
mA3r767ataHeuvi1QQc/TE+y7MMBD4M/WFz1DhgBHueYQa5jRrPHyGRZnLuChDopZSPBdzquVZBD
5gasmEVotuGvYtUkVAAhWSocddWXrt1HnijXzw8MY/CoFkH/7bEg6r2NikIe1rgf0PXiJ3dIzncg
3XUM51sKdAIO6S/W6F9dLdWL8iN1ELYD1x42uXI2g3z+Q9Hgylsirt1RMu31/F+b3EUNn9B9e3NW
n1FUxF3+gFJfiakjN2b2Qiq2uE4LELNPHVqXHPm29JKaPgDHtQ1kNfRll/AFHZ6DIooM5UmTjWFU
8Pg0DP1GO3t8Y4nyfgZmrd2uaZFkxjPg+ZC97ZmY1RJk/U9ofaZDUk0jwtaQoBsnT7cePnYk9HAX
wQWCxJghPWXk6vCzi0Hpa55Hv5xiUcHFkFwXog7ehvgFadyekSSQ7+OOVoV71Gk9rxcnu9QE8aK4
Pt4DjPECF8JuLpd1UsUzzY3f+O7ntsn2/FsBsp/+ArsOOSkTCY/ADDkRvPR/TdWRIW7saahpSJTs
WVbHuViILH5DsIH+HDrClGzDqoxZZndP4AZNwMY8ekn0AgmoXJQOheO+D1ELVKrjMcfm1iakszVg
u2Fjtnsj4pvoNJhDkFaBMxWTDSWgd08BQkZAyGTjhRxLvqAN1fLXa/MzhVzcIBKUFCBgCH5Adhaz
+ZdH8Vi4cKqPzaA24cfjPWfRai2/Wgkb+TH1+e5uEgggSReL5im+GHMNukodAgwwv6gTi6puktOO
zDjGtfrLRh37l9r29Zk0hLUlgbgknvZMcwnWJPSzx3qX3QPy6InsjL/ZTZDt52WtSi6bEGEiKaZS
MydgWqfoDMDDHwT9wjDn78wPmql8uXrsu2ndiyl+SGb3B+SosNLsM+O/iUhSm9Yq4B9zWvyqDub7
TmasQzf74/nvk+y+yyJOl79UvKzyXJQnv/Wh8yR1OkMCDA7TcvtXgFqMJiB20pq8mkl206RVqGhp
B2pMsAYGHq9NFyIML/K/odJxAHZBzsTY3gw5L556s+Atq1wgR+b6A6D9rnakWGkSuITp/YHgmykY
RwiHeW/ac1pnKeQP/Mm52CYQ3qmSctk2sTFG4VK+UFZUCNuOCpJ+RZritBkFGicu9lLdkCNnSnBt
Dgc2F/wqze+aFN4Rqrw5n1htuJ8fllxMjww2rQIluh1CrdprmW5K0WaG9tEmk4HsLSAtUKAtWn4z
1VUZIOWXuO2E2i2v0aiIZYg1W5dy5OuPwfV8QhdhrYHKnPNcXElIukcJljLIAlsQEq+Ae37AfLmJ
UilU9aB/JgrIW/HgvmTrlvr2wbFw9AMltRqsHk+lOEEVI+uKC0i0LIfG6UokOcLkifefnkTmFUu4
VX4Nx+lh2MGLhBGZ9Wo7zHYZkF2K0S78xBZ8IvyjmWy6q39+X9dJ/5Sd5c20qtJpZAMqI1DN1jjk
bR5WTqqhh5kCyhS/ASn2eevMIGXaU+YN8rNu3RzBVCFS2ipnN62FYpC5YnLZHAqR0/9sCvKmcI6C
G8jp8nOPl2e6MVpVhQhhP+TBoHd8ZG0aXe+hl1lVhzK6Wj2Ce1eSg/QZ/9WBpp7eVGQ3gAUUwcqh
scIw5LXdoGacVnfWUXzKxn4alnOuNt2ShKsIDNvA0Z7vRaedIhL1hdAPS0usHfjOLZHX9WDmh0C3
2MNBT1zn/JhODWnTnLtFcz+zhJEQlTcAlW/wkxuVzBRM/zXD+zkz/GHCZlC5n8DU0V6QnT3fS3q/
K+X/VfB+GCiHWYPhqC9NP/8Xa3Zr0Ur3q/XYjiATW8jHzeGZUOuakSH+TdNZuhZkwP/ItXw9fXWG
uDhBFcdWEzKPmB9eTi5KRwrXowkGe+iWB5DVo6s4m0F8njU26mv2MDg94ltm7m5L5qFPSGzZuZu6
yqouRkYYym5MeuGsAEj7S0w94jb7KZqE5CEt9qqCevLyh19GRMy5VnT/EuWhHZfKLbOmP8kFqcst
aPqUKN9XEmWbYO+7RbBFLlLewlUUOQAA1Zyfrg3uJN/mqEc8QEJ+5cRgHSjcIpKQRiAx5ZkZzYn4
anSXJf2ZskTGjedsflRbu4vcsIhE9Z0hanjV8UyR04/zlFRTx3pinsmA342Y6yNFeA4po92nYEOc
n6egprc92bX+H9dlnOj+CCqntXufGW+wfpAOA4MAb5pzqjDolVgxnZ/NN73LKALjnR2yYc4uiGVQ
hla7pAaV5mK8myzKt+bQQZc0Lb7He4VM37EyGgZUYTwBc3OtKvDg6htCWuJF7jyv9KHslW/j9jTx
T0b3jJnH+HveKtu0EQCqpuBe2gpeQVtdlbTp7Kr27rFfCvP24b5BK13qNyb+l+gf6RacKAiga8jR
Q2P6h/I58ry0Ve2s3J0q4F2H+sbEa40Wcb01NZRmPVzfYfOILNpYWjMyWjsMyHD4kVHe0xH8i4xs
FEHGpWbPd/IbdAHPwd/o3nqU4LM6xQxZUJZhDtgz/hzCL44B+hfuad/ur0WK1gqYeomIhjok5I9F
2ObPqi4QBLUuM1tvjUDSimNsucmSD1Ck73n0CRIuiuW5sTnkoyKLi7GQ7Nd/oKECgv7zGWS1G8F9
0pGQ4nHQK7U4MxEd3dKx53UUFFCrJqDRErUrukLFfZzsSvBHxoOH+fDpHh7kvnEyMmEm5RaLNJD8
A+isbCpva8SvAYzB8dk6mlNw12InDF7TGWf77LIUTmybk77xnggX0xCWl7axY36xpJxPctN5ts91
eSMnaqFDR+vFDoPJJZQ10ZQccJpMSjbMHfAz++2FTWJ0ldgEegvdZIehc4BRZI35aHPummRE5OSl
zT4oAAU8mXm3CP0Z27yD4tznhJ7KbPdyq6E0bx+TP5ZT6AmpE+5Y7On+9Hvh6oT38W/kN9vEPtfD
TvoFV0IblGB0XXcpA51Q8zZvqI70wNqnBbGybd/lftVP1yjcbd+vMVPs9yTyHuWUYkjkeUIHrH/k
kzGrg6RtsNO2ePePOyvQJ9VYTmwvtCtAuu71mdEC2KOYkhfOc5/HOFujbF2NqrgfGGfS8LLm9tEy
u1C2yWNMygrWl4hbxk+iqQ4QUesR5VpFdiLjvf7BUIELqCza3C7ZxamMZoC9ZvFNNRSiOoW6zX5m
+8PisZ6BwV1eLmyMid9uoUavL04aONRKBf+CQPJTJY7V766741JpatH/H+tLa4/EKbCxSn2uvvNF
gym6v6kdzxq4LsjCqdotTVEWj8gjE9Y6PUEYgWPwQlwRaD1WSNkx4pDpN4jiDV5oEJbpWdS7fOuK
stH4VY9MFYrHAlSuiiOa9KybA/vkeOlTeujRkbcmNjvjvncbW29aZ70L5LgEH565R/G605QaHx7q
4IUd3tCEepiSlFEa18ru2mtgH/Vv+Ml/5ZpMdLmgi4vzMW0Z5inB20Kxxc4k/5lmYnyaQ8cNASFv
Ksjp6n7oen+UgsYP9pORcCdME8x4rUxeKH287JUZ/G6FKtK0oYSL9dWY6SdLxaiQIETgtBfp8leq
53ibqZJX6z06I91C/DZTu4zB728AZxA9lz/Rx/q1rZWAKP34nhlOT8W8kEdMT0wGOPzvYY4YrUa8
jPfy9qEO9BrfvNP2vWtr+yFYO9apklN4qz/MbcCtj6LxR4HCSCiJyCUwWIu17SbuQjv/TRI1YVUa
0yuwUyCqZSST1NuGzJdQWTlFlgASqrvv/YmJMtzJvokW7KccJ7VkkACQKSktrl5PIZ6iGldSJSS5
2mYcM4gLzMzTsstwqDVFBsqWpWfw40Fu0CmJkWB0VB3R6RXv0Cg0dkfkcVjib5O0eVD8zOa5zGan
xjHRu6aqlNKKsuF2XGTGTk9bKdhdzajk6LCoEm6YksokuKSBy7DcagHHIhPj9RBkzuV0eplYfQxv
f7n5dapSr1KJWQ3YN6n3in/jG9skelzEF4Rmwaa/BW6Rg+nPFxKydplm1vYRQovFChD/Ihh2H0QA
/Mr2Yc8+paslnxfRPpQl73gcUz+9cjaNnbnCfQEbvITC6bFf0kWDurkDbVPjricU6dv3bFvejgal
vzjkwPPNgyVTTjRv6gzkvfNrXeKmtnDWy2nPBePOGSJtRreQEbjierCIOxoz2Cg3QKT/3bxdmbWR
j9/YDqvg2hMlm5zWKLuFMnFFz4LC0wo/uBNzNdBhJn3NR5szyuO3DrXJgMWC79p/NdWfiZEe0gKT
5IgvkLh9KmmL8m9+v5nuqDhdHU0u4u9DIRgtNY9HxXdhcq02R6IRraye3pMNUcmwi98ljr2YhXtF
Se2kLoxX19aI8dODMoxYFDcrlUoc+YCpPtLCFDzKe/kxpTB2E4q9xR8sTHlvkqdTyv4CBkCzUpdm
7f5q9m+eFSl+AWPCTik/0vRuH3BGxMypV+NNxgbHlTNfMNyxvt3y2Ig/S40w2uGIc9zf1N317m5Q
h04mWO8v6Uof48drt9Nmjnt3KlgC8eZMfRSKFw4wbTbEbITmHYI/iGuA5LWSL98iFBkInqYqbwZB
euSO4p/JoqP+7xaFQVRBoEXBf6ZMRI7WN/EXKvQ66r6p032JV+xYsCMhJ+BpW91e2YF/MhawDUVA
T8sWdc7UKMuG1OteowWKEfy+FFGsBNmUJI74mcoQyJppMjOkHh8qv7sOOKiSPuNqRwTlLVDrRD0j
pIAntOXPLfU3l9f38yE9DbsndbsO44ssadMYs1M33eBx2TJe0jTW2oiROjyjlfrg52X5IfvnYMmN
A1HvjzczSDirgsx6ZZgrZej1SIlZUyz0MpCtDDYVkj9xf+j/DZrjje3KwvLMubNl4+3qS89nlTQ5
JUdwhdHJUNK7LIDMfoUJJea/q5aTYjh1DgxDgE4wfKosiMGlzGOioDE6ZiNE5PontA4ZPoeVK4hz
BhJii5Ufg4SDeQIhoEIkAUzcWFTOdvP3pVysdsPLnnP+kvlmLqdBM/MouwAYWpGFIZaKc9gpC3Qd
82P8yw4BpLJdvK1tcNA9qRy2d5ge3ry/7hjXhMVtKmXw74Tsvop1ZDxO6uEGT0d2Kqyd5dm/ECYy
mYOXzysIHF0kET+e40W9szh6MSHJO9YMGtO4RefRuf+hYJPSR5RQVU61mccP5wKBTNMJoNrZNi5u
uavV3qWvKjIySChx6U2Px2OPLqVrYUdi+Dco6wE9rKPzonSYQ8cp4l1hMw7XjTliR1Sl8lcSbOXk
JRSVA4zQ+b/AK4nfcaDmYdMub6AwZeOrNK0lxFpjxq9KP7Bn+QLyuppv7Y5fL8msoinzFDLWwTg6
Z/qKKaVKxEdtnJNpIbCalcrDc2is40aXRR/cOGMjgab2DDhYSQaOno4Hiy3C9hfpVVbRmmMVA4q+
53BPPSQ55xFztuM5JnRcAZhXhNEcKOEAUDW+hxquAATAuiTAf33uobGEr1MEKI8ZjlYpk742WTpP
poVlOv9ulLqF8N2aZ7zhVyzlsfJWGAiQ2Wc5R8j4QCijSFl2NJ3ZZyswg2kg4BVJSUifbU55CWyp
RGXY3OZD8Ubm7bgdAgLDgW8ClbFfo9qckLZO54/AHKHACBaVyYGaH8xAJxmv42cQiIqzwJr1FrdN
9Hso8wn3MqusRn+7VMa+9K7NhqeBWIo+bDGLFgPulVBih/vypbrgJfvUXDYbZ/zlM/vbizxtlDTd
/oUxUmRvO1vHw5K+zs31AsbT5eHExvWKotjXIajPjADRiL3gKpII1TEhLrQXxhMQzVXZUeV0j3CE
v6eRrOmZ/aIJPKjtRjKD0c70Yf7SC3vEiP9mAQFmVhjVEQKcMK+2P5zrAeac/6ZcXn98g21t+jYm
Wj7jkKz4pYIZg9yQHJdvmKyCjHbcUsVIszMOuq+5dwHb46AAzobGvTgE+siskE9cDbyRGS11RWHO
0QNfhRCqxtWvSsPeWFrt9NQGQeHFVdCRiHSohBVK/UXks1zvZPmqwDBqMlzrwa26cCEq7KInEPPA
K1bHjEERHMatfUHJopYRr2djQtVqNFy5HoTNHAPTLziqXGGDv0fwKMXqdQzsB6bWLbquNyXNFnVi
YIf+aemzNiW+gaLwo2F5ofy8Ralzk8z5Ig7CfCNN9vYuAKHkU6iCg2Lbfbkraa0mNaYabazRr3An
VuKpCOwPfJe9MgVsSaw64jdNd6KvbWhJVroAIIXVNkXV3zYhQViqEtDdltFfrLEPf3I6K6eNf5cg
Ap51D1tahonuda2X2ni0DqSXaJkF04+FcIJyStecanbaHP5Rm6hFBG8nYQt1tvOgLH9vqQsg7skJ
QPZEmu2fcL4a2CAKLLWHBA6TPyak8UobzJRSZq2YCA5g9MaK7TIxWX+bhUDzqa1muMhg+o/78kkz
Fne/VWkl1E+J8cxcU7IW2knJretescSiLXdiyNXncDZtp9q3z1TU28w6H74BNjZ5tSpVDNn8gH+J
WjNAUYxnMFJ2gOAQcvZ0x1iZ+ff9BM+u893vRRrXv0o7QQC/reGgvTU9h/sH1upJz9DMbqmzDzDk
hc8lAzU1513rKxqpBMIop9VICm+O+l1b2A9aaIk/RqG68uyvt/4c1hxyBBGkf/eD3YUG4J4V2x2L
jDLgQ1bMQQMg6VMXwWcp+Modz/qrMykx5Aby+noiubsv9XjBlA3ld9eDvVFRlR8zfMubm/1+FiUm
lCLrY4G9s5C6MaTbBVk+uuk9KBAcoa+6YjqQ1Dc0MNQAC5YILbbTCsK5IQY8KQEWBRwBM/H8Usts
+tjhAXG/J2M9n32IvN+QUGkCI5xf1kCFHxIqzpo885iTpK2zhnis3UQtP7yXHscWqwWbu064hxF1
wtEVZUEfWyrFxRgsR0oA62Fuil/xgGH2QDbdKZAXKDxiAkepZHaqDkBsGO1lcXaF9q5Qa2ZFa8Ly
gByNKQYs4Q5zma2yGi1qG66kGKOD42jumICTjlRAgXOmHmZOjOlwSgFDR9ttzEHp+jBh2MffsWrd
xQC89AlMKaJtEBHDt4U+Fiq4konMUz2WCjtt+A9OirpHkGfYQ29VWHKcl0dvmZ2Pz+eRBawsl7Uk
mxkuUF9Kpri0n5xpaT43dZVy9x4VsmiYHd94FOzb0l2IbGSr7mcolz6Kn09a8+ws/tLh+Ctbvivf
CzZJy5UWpKeIyk28TSf8bMcqHeCsDQoOOFtZ2JsGAH8fc40bIdqoAEuKEQjBkUGCIYsVCFlVA0Ts
6MMhFsHBdF9vrPYXYaoRDU9I3IgxmeKKRmJXniKxh3ja5q2EToUGGCM92xUnZpzR6USGrpDivocJ
VRDILXZkz+MNgGwwvGUeiJnjZxUOOGlcm2lIU86i405LY6cxfYoq4dJKFZz63SWs8bd13OUWi5wQ
eryozE5DTykdmUcRhNyu48P9wLvJWQlSJexb3C9ZCfkEMfGM4o8tqB8+aMLNMPFNp2hAOwv3jhfU
8fAXq5x1bnEYWWGpzgNghWxkg/fliR3pd1OOMUHNC9wgVtuoHag7yvGJCEh14THuV0UUyN/7URy4
fgLznvDDcUmjLkFDFDMK/RCHCyh51U3f67LbLHA20MgG6tC6rF8hH9PsmP4WGfgvJ5OlDjFzOqFY
2xMDPnpQBS57reaLWRHjBUPBrDy1GVGZdKnAcMC31Kg1Y7OCC0Vg5ZH+m4+iOPu0YowrmhQGukPT
Y5PMhC9RDwgw+b1U8DZB4b/7RcMJoWa7wvffJ1fPhIYvyArODR/652k1mWSC53JmpKJUE1mKHOpO
cri5W9BUB2RGJtyB6iY8/wB3gbNtjhw4fyXl8P+y2z9dXRfNvZFnBeLmr7y+3OP07SeS5CZHZtQJ
lhkbwFAtTbApHbLZrpnIjuB2pq+OBWvAM36Y6c05xpRPBxsNETRqko7itTmYCP4c4pMJtrmj1mqM
xBTRRdM0Arm9iulDg5jUCttOj5KBzL/59lzSmIEmzfwTxiBVcA47DTPq6WIPeHj7ndEbJSfvSjNZ
E5srZpIqaTxAN1jfEBNTWMQcmQ6EoleXeSX73oBc/poGfSUajVuVTMI1TOURwzPH/D1cdvOPEMWH
Zj73nBhFBdXctuNHJwGRVy5T/qKCKgqJxe5P1cQXq1i513HIkG4hO8VLPQZg/ubTBd+v4SJcMP32
mONgxZAsVyHoAL9MPzCxoprBnDJQZIJZNZxDcWpYvltXlNTgPQMMfNaM5PB6GN0UuzLtMEVBN0jJ
+AJIq6wTDLUfA5QSQfJTgnXzD6Y4ObaVxw2y5HB2LBSA2IRnBfgfbFX+P9v8XAgGWAKTM6yyMEbP
tN5NLpQSEdEih+FwXKlIIzqdylCFHO3g0TvfDV3HkKHeamuXKdU3DqT6wv231sKYWTxNBcarnzY1
a8FUzj0GMbXRJ6cl3lC/19NPeil/nx+5xR8kjkND3p3Je3Lnc2RViWtnuLgFKHA/9g83WO9PWcMB
pN4UGy5Vto5HwehEVPutQAGqcktIXimBHeVZ4ceqhjBIPmH/7l+PsLM2tfLqhKLqnsm30v4S9FmO
l5ciVH01e8uwkOHOYO0BTl0Vr0kIRdzOMPz+BQhIKrPPSa/RcCsSmNbCA3twQNOWf6wFIKC3re5w
YePb212IuFgLpbt8Znsrvx+/grpdMK9AdbZDBMACoUJbGL/o6cq75XCv/lxu7rMWSocRK9lEtLt/
X2/iepOXV1re6rdbUlJ+fAi/RctYq2mkka7pVw3efqO/YfwX2kCvm1NWV61KW0/SZcQJIuWdpKqg
oac05kbxKQBs1vKmzcY1ZCRzOD8qDQE7ngzcXd3xgHerL4xlufg4swSf4YKVjnF+2sparO83FYAX
vvFzA5PQnrCQDcg3je3bo0BftPyZa5iogYCvDax/PXztPLmG9M1SE/MBHZEvbpoZGuTQPDUIZlvq
paVnTWy2vxbxvZhm5Wo+rA4Em9BMXF0CLN0L5en0DVV3k5qs5XgPvh7tSusEX+g1GGO7pjJeBsXJ
JliflgQtsJd5RWBWprRqw7rH5y0a5EN9EHzV76ohp8tU4FKGZpAw780eqYyV92manpEfPlKlYkuL
CUkEY6rTOLlXdpo2w4giiKRcSE91p7RAwtAyLG5VplyPFNSCG1Yf2C4zo/3c9Jfzwqf76WuLjoVL
kOHvqaRXhA3jTJ7sDCBp7bZj0qpYfIfBJ8mprq6R4XJTtpJlhf8KEuB+trd6QFDyUdSRyhJ6qfWv
Ztd7ThzW+d8WoQKbP/1dEGQQ8+nUSyo0NLdwSURh1FUs06BIW0oKh8EdTee8KFFFYeJorElsf9Fy
oGFudpqim3KvA5bmEDcSq9IACSybPIzMxcpUaDT8UQC2eqPzx2kwsPXWx5Qa9g59tw4qRCpawQFt
5yIrqvmEBXkgHh9+ntZyim5TCz7wXGv31Jdx+T/LZPbE3Pd5t0d8EPREfke7l6SkDFFMbCkQb1YP
5ahdZUvraZ7j4Yp7pOnzqXoAM+Q+Ik8BvH78+EVXQovEfSaCB+GCBdKllMA2NzOifpP4XKR51iJv
uox1sJmDIfU37bLtmVVEoUXXpD3R4NI+WL/C8Ek0ra2Wp6jz9YWUPoCxjUNrWvnz0h60Nqv/d4rh
XNLxMb35yYkbpmMtfbdBqcNwdkOWb/MpRb16z7dRzHlvGKVSOFM/N58taRWb/tWkb9i5kxlnEPam
xhkbRnaUioCxK2ANQpyTOlyTtUIfSzRVXVJdiRlCWYOjZ9TAo+o7HQwpmkFn5tl/jeg3Yhx3Jp1L
hVrtfqSBv77U6z9+kKnOtRh6FacKMTSP9L/z4M6CuqkPmNnAJjqeQQiSD40hWISc561YSX/HbvV/
nmTWMQPfWEMSf1BMRfcYeY7PDU+lQIP3QjPuDUmUtshPR7HWMQ3z2clOMO02kjD58iGA6FEszpGD
TvJjhMC6hwbsxCyKg2HXGHiXmeje/x3RGQCNddxZRg2cxssn0yz/c2fBy46ziLda7hB8dCO/9F5w
tUEY47+RRaRnPZeUTGFfAZOqRU3BJECPTZ+mTIR3DJZSMfUsGboqtung1eBj539JvHNrssdkAJYe
kYf3ZAyFn23vRPGMiU+skqHNZpK/9yk1qZPM7xBM/9ADKs/qq4Bkn1TvmB9DjMT43NWnIJFw+Ncd
5GC2qugKTCHgNhZCu4g8p0Eu0pLpmUMRJCBluR2D9U9GuJLxQvneO5PlMmznqQQlNIYuu8z8ycVm
vUZSwZEmCw4Gt+YeAklGUTXH5IVxveaJu4Vq87jx1chajyJuOVKRD4ZqIZjhZTYokOMEB7+9OwSQ
RGnOR5TL14yn+h8qd1IoNDZKD3LYkyDWRfPVulXF+dx9zu7FQof2aM/La+xKkPNxnmAfNuTC6cSN
mHk3FeYswGb0GHXmof2Vm8YyduMctr6sE+BIN36zIaZriQ1Jfl3RfJknHZFE/gMFyqhHQI0zgS/V
tNSREf0HSpcKtEgH0Rah9T7rLkMUho3+DqBDZobmZlpzPU03lHHh33GVB3Yp8SZL/XZTYPZXy0fT
WSGRkxm0Ir0SEO25CfgI/iQTYMGiIEr+bv3v5zzByUBMw4t27MHeu0NwhWUFkJd81SLCsQHQ1wD0
GKBNqEShlbW295xE/IBcUupu2ey3/8nuIDFjs5kGRKginE6XDL1d2OrSGPoxR2edqOylGRZmfkSx
+Fwt7CeFUY9ZehN1qWnFs1uc+J1H0wlbHYX3KaT90aHe4oqlTjTNRwaDT5w6CvOiPhmjq83hb/yx
l/wZ8rACMxRUh5B8FCtryzm7d3I3n2Cn8ivwsOcNon1EJ0CwmYzftpb+Mj0AN7w3u6zxVf48MEkf
ewQdPtWXG/NtUFu2wZYki3IGdIZ7Hq53aT60Z3VaQWIfteA0/N9QHWPwo0boFk1NislSjn0adLsT
Jw04+6JM6lF5HwIsvdfTX7NlrYP/YOLOWx00k2kxOt99n53PdCklrJhIPy9OtG6gtU0AysQHwFup
u9AYNQOvcdgMCyr9MnPBGETkl0rtJKLQG8K/1bj1h0gliLr1HZtvI4yXjpMbPhD3HzuDp5Ho6WSW
aOc+q0t6+OECYkMN5eOgD5Zt/7wjGOkPu00ws8KgfaSZArDYc7sXG3XwPQJQsi9iKtErCaB9hucQ
v31QKy+AS05ppLLrf3Cu2dKeNmOdZhB1V4M7uPa9SZkT5d7ySa1aRFzDal2fLMEpD8v/2jOnRPkJ
rK8RGyV1pZ6YFnZY0dr9O9w5zLoYyX+S1/DFPA3/UUQNvNcl0xpUTCkFEWOvZ2yj9Jdnn6FDh4PT
VjUDGCaOwREfOYRIWhGJfhgEO23+fBbMbEOJ5pKOVH+RcGQ68AVz5nAkof2hF4dzNYzV2Dl4j0Ps
Y3N4eMKrn85A8bsJeT0CYNG8NAKIf9sVT6elFRKjIHuB06EX27oYmGbjENEuViS6nSE1gMrGHYRV
JzU9gGnkHUNlpywufK4NGhFEfXbH9HGGo3FpXtZdCQZKPQZe+WeV/65ua4r9OwWmDPXQbGRyJ5zI
5qY8DZDHRxTBUeISd/MDij+LJ62HKUyuRU0e+ZuDy11atYgiBVeb79Vny8T5ZqlJbD2jqB+1Lfk3
RRVihEkP9MKlaWRZdDS6hcZ6CDvIqnvF0sLnwYR7Rmyy4aAZOOnZeE7JIFLEQiqGmRZwRcpbRYPD
5sauAGyiWncoyfMTkXKO3E3oERAwiG41X9YnEFt4i7FFmQKt4YMt/+GMKWSiyWLjvKH+fDbcCw/d
7zF7IxDh+qF0Oh5RmnqjMItfGydcw4XeriyEIpvNnPNEdupaY3lp2A/t73n4/TKCCt/QSVhIrQ+X
Y4xmYYxu1nAn/SCyKGBf71rlkEdd4ezrPSGa6O4x03JhuOfgIEMUX1K+LWgyMzMg8XzQQknp5Z50
Cax+LesA0lNpN0kG9Puj1ZUg9bdcL+rKq+tEiKS3hw4LNMJmoPLjetV85yzZzTJsaGVvNEJ+PHp3
hH1gMTdT3mQfGOosiN+jIlCzEs2ZjucGBf7nP7pNRuv0phvdMWp+xxXrZJNROAVqCxB6HNW7OWvd
Cp/gvtr1YZzwAp/mD+3/FCfZv3pPsBuv2h7QTnUGxYIm9oDjXt2vwyrKruc3L4Z9gRL49Eu3oRiL
sDEw7kvSC3dEpvrHLOtzFGWSKT20GWnXzVOH7etrlTijMjjfTcAVyGHCI2O2bqIlsz7GRtym1FsO
SHpePn5sWyfIfSelGbnRZf6u+p1nCTbr9bNwP2Xnm2H/YHfiKpcDnmkR7Mv+gx7GjfYqCqrbkpCv
jqcU9CAUVsx3y4JD5gC35+fCQDyWR7m5iesC1mTI1t02ubEMBwFMNhLDHiSrwpzAjd7Y60ZwjYXq
1P+M/ausRRqFA4d0mY7fHUw+P1TdZv1sNzz1gQ166wrw9+c7xB9fyAqAdFgQzgoX8TKkrJSwGpP7
q3r5mSMh5kxi+RvvoGPb/QMEqMk98BTiUUomeM+1IfCpiuNo8yEayDpRQoBcFs4GMGhqygRDS3qE
8yKKv10Z2zfzk2cx/M3sWp12DTOntVaEaMvpqZvoIrWBFSsO96dR/gJ2fU5N6fNWNxCkzWTF6Jk9
dVXrjGnISHQ3a082Rqe0+p5TTOArNjJ160xzEYVfHn6dqDrnNhxIpT9wjsJeJlejF65M6sFOat93
5WZAIl0Y2Zprevv/5IupF5sQ1skB7uDlCP55dSGgD4GTGT986eSdto+6CKn9bBI6uJB3hILcI2y1
DgWdiL7Sb2YErVQSOvlWw1rNDNtz2o3Dd0hx8kz7g6F3tzQ9s5PCODWn6RMJxkb3yCf5ayHudz3c
1+B07s3n/Uvv1ZYJzmlNz3oWYBvChrWk899IDySepz4vm9XaJOTvwS2mSnQxstpgGaIeU84wq7f8
YDcgQsFdk8Dz3EXbF4fQossfg0dcGhgdYC0kcrG2Z05X4kWQTKQUwkINmZi9t8llWE9TjmBsut7K
eZDIywM6lozzV1jPFeHzDe9Rs4n3Ec4u2y2zHwON11ytK+5HzlX/pEK6ZQpiPj3aIFXgrW/wgiJf
usVyYYDbp8Q53dAVz83qtShjHeWDSk8r3uckpuBmBvit49QcHIL5Hb0Bz81jH6sdgPiIyblnyCld
I38z92w7xvH2hT3e57t/FN2cMBN4vEOBCRfgbYn12APmO6Xt0IjtoqAAT9EuJzkbaWDsM5OkuEyD
edGPdTHszTZeplrAKX97iojv1wxt0/tIsJw1gtBiz3hTWGMUJBdGTTR4MRtjtu/4e7RCIdNfKjXx
sHYp3b4yNc4Wu6P6Oav0LP5PMr15OIEfMMctFLNCku5q1vQzb0jUr3YA+RS9PlOlamFKZ4vxmJqx
SLjh9oAtB2Oz5puG1Apc0IOH/DoBp6/4FJ5Dux1aLsZ32SEJvduS8bMRv0pQv/9qeUyy9QHMg37v
dbPHOkja3kO3ddjptdNGhg6SC+4TwaVKenbWfMXSnZBCVubVBKjkWofybXQL0BYzqmVxChjWXEWY
sRzuSIiPFGH89wuxAC+woIo/qiu/iAyFLI/G+k3AY9p2XqDEtIsmxFovlwuEYdH4/PGhGpwC9YcI
3ubChtbanAEN+cdiFDgh1UD6H38FYf9gHXBwYHxMOxEhcKV1kOYcqV9adig8vNOEacaDrOhQShsR
USD7w/+iaJfiUF3u28sjM2reM/km7ICmSn8/UyfpeBXmynms4ataRhwbB3r6zacld6s/w27MZiQR
MzqteQXQ1HFuNTGZXnp+nz+Id920gaJB15V89XdFQSddXX1EoXWv8THrfU8P02wrwoPwWBNLCBeh
ygnbfSYHwioEDYkVD1NUjntxvgOqScVzAgsTQ/yu8sJRuTYDekfY0+oy76mcvTPQY9auGWQ1cp4C
IjPqdvvcKRxp2AWQVVtES6eEaL35s7ljmpYla7mWzbdPuBFDlTk7UUuYhGFXXfHRXsJBQ5XDMbdB
lsTw+FNpiXrsD24VkCquJ99F4LSAhjK/CMIItetSYENkGPwivx6ThcE3isReoL7oQN2BfQ8Y5B0J
bq3AI5V34N0bMVtfzJyC4TkJORV5yVqzmG9FYdA33VjaI7bmr5tNRxHsanc8kORvw+Dxe5Xp7Lti
MC06iMhq8W3a7qVfH6lMfNVoCenEDI5DYA8Ok5w4e4YHjg3N8KyFt0ydratRQW0Fh2RL8h6FB+CU
KZNfIApHdpNnQb7EzH31MKiK25D7DWyyPqvRdvBJTvKNxo/9Ze7tIeXY/QWtB6ZI5V9vhlfG/n22
cbXFrx0AEcahVwoRJ091GIEQq7VBy1ZyrEDqMXt1dF/OV+UPiAaUtRGn/wrnALDRKG9wYTuvCC+u
f723kuoWApop576WHoKlogrwDBJ73sNpL3kMHDZfrJ1eTz0Ia10vSWcMiLVoaMTlajk9DyXtWSN9
broOzf7qaI+ar+9mCh3/Dr97Wae2FuDVk79pB0k0e4MyE40E04URt8HsXeJMTIgxeZqE36xcydYL
ILl/OAu3pUD66ek7u/Geg95QAlz4Oj32R5qOoRi4pgWKcHgGDhCmnaZcrutneyf1KQgRuQiyG/nx
bTBshZVoSyUXvLmfbP2917qe1IunmptXVevgjkk8xg4C0Tw3cNTWuJnI2zpvzGIfXMV0N5F/e3uh
TCh+q3UevuFpkBuaQ/qvCJdVY2fCx5AXeb83+Kx8Qf5nRHNhDxxXd8GJ6DMeiYuvcaJegYl9LerW
PThkSkPtvaSOJ07ijn2Mudpqjh1EThDqzv8OLa5j068GmI00CvgqX/Lv1h4x2ZCDLj8uzMeQlag8
vKX8cM4cC4kZplmg8GlxVFcHeyX7+tBEE35eC2sbF7excHV3yp57XQ2GHpt1SS6FBPy1M1Hc4H+/
xPp17tKEvW9lhj2idrs7TTymN/JfA0JJJ2uAj+44RVVPoZOSA1eQdehECkBTwGRXe6dPXq/JRQ02
ea8WAb+63o+7zSHJO6xBvyakSXzDUOU16ETwoyLM/D/WuCDfJD1glI8SVqtXHzQl74QUY2/33ylV
Sm3fXjDDoGLCwz/wyM6GEGyANHzykBL7fe4d8MVkQ9Ls3cGIChuhqPeWmwL3k9FciorwDpMAn8Dz
YtXShdoeFrkwq9FPHD2w8Gb5ASQNdhkVwgTS0ojAAKuZbYcDnR0+Zdwd1O3d8su5AvRQh9CCM1IA
oohvO0Bv5ovR/tcKxnQOSnLTlZc2cTiCDlq+FGbzWSGm15gGIMDmmWEC3TcSvscr07o82PXPekEA
OMEXBWkjuu+JxPR29/4U5sSXCBMsBjYAOttOzOdglaGo5a/a73bDaJXJbXs6s2HiD/eBkdmccC7H
9USEvUA3YphVFpzoRCnCLgtw2d2UI0KZwuBALg9tbzgJt53VWwp4r0d8GbNpyBvLS8V9/wA6rpuZ
ktMxjADt2fqjWqtJ9f/M9xPIS1uy1gmIFRyrU/NfFzWGwWoCb/1fCDEoEsT80RUwgpOA1+AK+3KN
fr9bYKsEuvb1+lWVT87YKKrh4qJDqU065ALtlA6Bj6VOF8i4ym0Ez11ss0UH1BJimibHfEZsYlfz
jDs8ks+vYffQrhGHSXDlgXR1cNHQ/Tp4BJPB2KzdgM4Gg82+dDdLfPytdPD/z2lqn2oRVJTA2Jqu
dTWOf1uTvyd8e3ACQbvVnd9J0kju1poB+Ltih9e3YUA/cSJAF7kZUQ+OYMDhDZwl3qRA/aUbTSwT
AeyjM8ll+Mk2n4zzrv5ixyJzYsr3PyBTMbQqqJSgD29oFSjPlyEuH6xU5zcSCAVCt4GG8yM8cc7w
EPMBDGjSKyk4aWrxQTf/HT6YcLiIMVn8xndTVwOqWlm8faUjwdjnWLX8USd8LzaRxaucd6tKZcw4
aCsEK3ZfgHqqMowqvbmMfnhQfRTBW7Rz9PJCX9+Zbls9CA70eYNrdxDXaMQxR8z4Rtx053XkbzoB
fUFjBAtnngb0hl+cRHIjpRhUE4KsAb8eYHu4JtzWIKk8NHj59HtByYuUbVWQp7qABqLqp3J/1fkU
qRJZdXZ8UOkXA5SnS736fWOggqax/ysCnWpxVxWonXsY4r5V9GZ6QDaurrRr5u7mwrLIKsa/g6l0
YM/Zzap31A//nPmNufYoYCn5weGj/tf3Uaza6vhyUE5Er4rUnMtx69Zjtg2/14LSN4BPspkl3X5h
LzVes7lPWe/NcYwl/cm3/BLAN5uMSj0F3Gp9tZfSzqZRHG3MC4Bsriu9PA4og0ateqroQM08jkaU
na2sTa7f4IdVwpYJ3nV5edWAQirp4wQ/ZaKxcH27EJMdrxVy8vPsGo8IamhCvP2/xzl5F4lIOLfg
qOimOOv93N6DFIhiStLbAIYBTDCG/wNFS0Q8hSbkpHnhZFBIM/csoJ1uvT5modQ7nzguQEpVV+Lj
T+HUpCbvukAaiSfjB2nCxxBqW7IPVtC3kskXye6keXJgf+RNC5K7cIdBpStXhJMZDNLKAPEmwDIF
C172uMhytqdwaCU8qKMyNnklJyHMw5kh4C1/vtxC1OiUERSA5IrClmEc/0nbZhG/NbdzJpFF/7Pl
NiamV6Y0I67rykjmn9Bi4o+x8Uv9ikLLhUeIcHIJXEjc9ohWHnHXbiVQVIJAiV0KTAPVXmBRdjAA
BUTBvYOpY0IXjHpAEQ2lPnvon/VN7EXOGVbFSBx9Mo7QJgXgcv5llYaHqUy0hm/iWNO/ZkEWrKqU
OJOraJuXbk0l7iQ34BdLyAo0EhLT474GXrrkwTx1IN1yLYuMKlkOHRZxeciqeluzavlRTSR/FUTa
4/5J/ih/v8zrdnsE1lPUBNa3ySM447weVCMH17BHGDftVLXvIH2mV4p6qlVv2qnT98LDREWyvMC7
ft9ZvzBoTO1y+goZfUNobcFpSrmRrubI7AcxtWbPZiQuLSdivmY1m6E8uuntd5/C0O22dtvgGU/h
yCATkbJueRpFVYVKSw3EXwOvhHeRw7hjznRFgytda55SpnXVji0qqE5mA+gbE7/ha4KueWcpNv7l
aDUy8QvaYLfP7TdvRnMjIaxlGpuALhqOiZRE7H7LLvvvv6HaZdzdN7tJoSGq+Kp8xk1rH2KbEzdI
h+BtggzbpVBr1TIU4mqCVmYAdV9ANTPNNd9nigh8A9zqmVGZoXbi6Vt5BT3dV8Y4UHx3m6TcPRfr
LEL6vtmml+WkeeCdht0uA3ELldKTbZUmUmO80hCV1/j6eAmMDKB4XpnOyfpW2Pn2M+AtqPpVOCEe
eYYevdg59f/KFrprkjknXjzdxmk6QyFFPsPlttNTnwFgGV6x+KvK31zr42Td+OpKGlzEz3RGw7/U
rMLWUU/sWAjwmACREygSBeOYz6BIjKWiHysw5pzyHMrhQakignu/YI4efXJtiZnp8qfe8qrDbLxd
J3ve6IaGRIytxxBOe4yM5m+S+hRyNDiioU8FoKVy4Vw4gOLtlxu2Kwsjqz2024qLU6VDQh9BJZ2R
FmY4J8/V5ztaqTCL6asI8QoSGKiLyCC81pWxBF8o9iYHDyXkAPUj40Fkhqmfb6vQ2XwIrF0/CtOF
SOM3JMUzIiFeH0rY+IKIPFTkW0ArvtbHdc0Yx2xSdPxL+uaxRzin+o9hpq88/QvbEK+T0rQSUkyk
r+OxIa3o3D9LfqcYYeokE8WnixsvMKKLNbpqBeRx8i3qnGAq+X8skpTsFZ3ZlFVn+m69gqWnT4NN
AZHhWGOpem/VUIwfV915/p1haBQRhCiGiUxd0PKctJ5wmcI1y4TUYojVTq/JdMtNN3v+apnyBhiT
2IfVECzR9q5IhxZreBgwX07h5/rCVPwn7iuueIBQukhd9V6TXXQrhxtulJsZYpbOZVR5/e41ZdyS
BuGF9+q5wsPxdyjyxXGRYfe5rQVWVMH/c9vchLqCOaLdiPf0l6fGhCX0xy4uebLOhMyLG+o5vZtI
qX9AKXSF9LbXUcrowvqvj/H7J0tBXGeYn2uaBKELd3NzCaMi7AQWk3NLfsxBFT5iJKYWBmVU0hbF
jh9ev/kqQRfj2Q+KwADAlpPlhoDqMvTEKA6JJ0JZ+M1ozRQB4gpM5f9vGx04vkugHFFVKBcfk6jF
MdaMdP+YsfN4qVp4fE8vT7z8SJJ7a0tB6HHJZjJr7WO0fQewc9MmIQrvvvCmvSqmGy95Rrw5KKwz
cKXoMENqUl/0T9PjzIeXlXH7cjWpYNonDv/8Zr66U9DlT3EG8YUjbTNCtf1Wx2zo81Ej9aZf0tnd
O1Dn5m3LDcdq6eOT+HH0LzYAgBurWjkZk40LDZZlwbotkPPJIdT1Q4WIOcAnPBXcQ/ZMQL6rL4zL
qWRdmTto/W6nC4+Ss/BuiD0GR9vVG77LmT8ilYlsRWfAmWoByrHHIQrljpNd3IYfnXNY3pK12yqo
ugTzdi4Npmf6EO42E45z4vZ596IvFUtcC0+7kgNHke2GzaQDvrp8Df2noyXpBLKJ6ZfscwSkdOjP
p67WsA5lKXJo5qzFgzLCivlo6gXIJ5UuySuuPQ/MPpCXmay91Qct/PBMmd/MhNlih7npUs96Kmfs
Hy5FCmS/IwA7/gY347mtDO1FBEpOqUQgRl+140aeJNtQR9mPCZ7sOihm7LTAt6vE2l1vnExY/Sdg
BbkvEL47i2+wT0UhNRUwog8SxhjTOI9COEzr/3qLc4vo+Uahxh4Hm4NIP59hyJg5McvJZsfVZ2St
3brtblkPdSyLZ/nr8RNZbcHx6mYgJT8bj0hROI9zt6lyDnTXd3l1ziu0zRQrz72Kb5sUuu3JtPsE
8v/N8j7diA+gygAC9mgPxmxLd+vfAuS6l9Jajy/QlH70q6jlGP/ncmyw1Yq/NrsrCqnoOPprThS/
KaNzg284PEZYqNmX667BQKAjWhba66rKXY77jkY16ZmW7iWmjwOHF8UuDRztAAuMQOUeOBurQPDH
gT9TdFgNFZ5ThvU69yBxWxFyq2OXkg6XlkwDoV6UiNOcHtcTu4mhGfAxt6CuVdgadIHFOgRCJk3S
mqvVNtRs83334Vr7hP5eNjhBBCksRiYMqHa8NPKoJfgS/Ky7/H6oNBD490xRbXfaZnovewdIhJox
ji2lmHKPEfJbcE2RDzIfmGzDuhm9JkK59i7GnyNN5f7NnyOyPp+cVp7CKgw58yXdkEzo1W0Qp+tQ
DjHEFm+XeteKzgNVg69ZlGyx6eJb3oVXSbS1GIOf9FpMTZH/3StlE3atkNwSeSqQL++UIgFaWWou
YxTUSbnWfn+ZBW/h0EW55zzPdEGitE5LjktQMolrAr5dgVzUQ9ENutoEqfOlrhlZrM84IuSpSZCZ
IdBgiNOEy+CO5IOu91ZJEbhfYjMMVeql4AKL/juOSDKFAAncLHnKyQ2fJMboP+XBI6qzRyW3XJZ+
SCVuKA04tZwcInZntxbk/nruWghEJIaNEEMKahxxCr2JlU3lbRvr72mwwcOg2iZOZ28w+Cx9Uspc
ZWUPFkSLRtxNi5wSsAv9zSKo177Z7WpImJGQVUe5+8uBnr73glQddWxc7dBsk2URLtff8lruzgPY
iflS8WjenVb+BzXR0HmZJtFy4WHPDdGlPQfzkfTtLfzKL4QHrdPZs0Godp9CFxrNykGqK4fH+4Rq
bCEAvLJpmxr0o2OYxWhex7j6YmxavU72naDkgWPHLNsIdnjCo7009j6j3+IE5axM82YxLmOdeVJ1
jGuv45MuoHs39D6ZC73+8C6UN5H2AsnMNc28YcKMgnhxwT3StKsb14U+qc2M8zVuaU/Ne08JzSSL
5kJWUqEUQccU7pAYOxqoJw67XbKX+CIg8dEeek5Kl0qQj4bxBvblMvzopPO2+SZRiGytG6DWrcYc
3UqKKS5VGSznuYZG0wBkQ7bNs6eE+mpLPDBzfccNAKP2u01lvWoD1nlT0WeW8KPJaygeTBKUl179
Dg8bzQIU6qDHlRbNtjY7iRrZwIzi3W+zUughyAUaown+vZPF6xeMAPIB/DSF2XSTgtFdl4RSroLf
cPJddEgiWYz5g3PUk50DrNy+xbQsJP7kcKDZ2nSdcEK8wxTRhVQImkNlgQ8xAPMKFCjRWujT8QZa
En2xB9bvPOOg5+ymk8R789ieatH2Xh0TsdOCo2M0XjBMHYX2Nt3Re3DrjN6OS46NaGt28zR1eiwU
17ZCCSA8mTImddy6fdT2d1dDobQW32wcFEzqstYocP6/jcXcaDp/xDckkSMin4Wd1fgNBMK5xng+
/HyaM7ErtCGi3qq90RoRxC46rxN9FeM9lDiYRbT4HeGzspnBvLdT4ltXZOvnCJCUiY3WI6vfCZRO
5uWFupHwBkPFFTu/w1zUqsIRwecFav/+5OjiyPzekjT62QuggXLu4HvXBeBZveGrKIyvRQpMVHT8
rNIrPw+3sthE8XR5JmogJTjf36bLs5zdht/ZNUy5wzpGNVqR/fDmSOepOv6q9Kuvo9ivQJhgFumR
zLfHVi+NqQ90sN1iZtDcEIdIeMa83b4shUZMZYrbVTC+AbwIf4azwzkvSYsRTOV++/jgMtvdFceu
sa8ko0GzDuWGYm6YLSbNjYJFLv4DxeQZtrRw0kA/AFhyyERuPPyPWOUemjdDZB49T/3n3vkLbRQp
cKN9EOPGlw21jXuCcIyinkOeuSBTQ42eFOdfwklwliNVZB9uEWhug48OWYXiUme29kIpESebv08/
w7JsoMKsyuSHpTs8OYAjak2x25Yr6J0LScLF51EheS5IMGMLxXkAfF9XDeGrXIFdYsi33a+SJ5nT
p28U7Y2HJ+5x6TtVTe3Kh5xZEetsE6084elE8EzhXK24oAmnffsmUxKO/1PEeXQp/BCqwG6x+AXk
bH4dz2n6ijREKjtxZcNloLGkgceXbP1/g4fKIGPuwgc4Jiyiu8iQdlwhiJOh7IK/vBjoW80mDYnW
LhiHZIewUbWjj5zmsK+q2laz6js9sJkbYrU7VICf92vejix5Mg8nLRPkEvhjGKJB3ZR6aO/vJO60
twWTBX/t9jAJu1fZOKkxxqKWjO1BWlcep4CZebwEJHvcVyxcAkVP6Fn4hWLw9AiefQegrHE0A7bi
VDq1IUD6u9JjJCHaC/av0zkQLhm1qh99BX8qCwts40ewpci2851NCZWBdocl7cW9iXTrvjgbJ+6K
j0jz7Ua1DpwBonGWgMSTBASTANMXvQkuZZqKVXj4392BSuSzyohF07tXI9q5XqASzZbbHCWB9FBp
10TYN8+kyCqxh7AlPk4KI/i804UJTT7jRaLnG37o6Eq27alOmOQRmnlgF+9x4+/cBeNy9UX9C/9C
KJtVverDgAGM24VGGAxxzz6ExlCm+csLCbUPeqELj8cwRxCWAHsFSMe2iF2hhIuJhviNx99OFRbP
fSO0U9haTzwjuYUN9t0Ukwvaq61eFHau7Rcx1B4jK3gca7quruH4VORrS12olPjGFT+HK3KHlUJT
X1kppYEPkJe7m0+QclPFOqs94He/pQHHxlJvSrsmiiUAmfFr9gSusp/aWzNgsQ8bKyM2My6N9dq7
60tg2BFPv2+GHhiMfklwOX8hDcWNEd7aTadmvzs2pfMOq71veQjaUGsjK/fjZamrnliK6Fz4D+Ti
tIUTlZ5fzJVig+nUW8UvHs7VWtXn/aalge1XB/MlGQz+6kk0T2yhYDjMVepNaWOXwrKG4a/wQPII
84nwNOi2hLIJZ00+IDoHHAqTsqY4ikj3nEtjWV7gTxqm1jbZf9Kw+pGv0ojxCp+iqq/e1+1asWT3
ShTB18EDfQzZ9jwIuJBQ3qhvvLMRcPrnQuXIQ8M27lon/NCjCSVpDJv3G3WlLsItkolPgMUUUeg2
VWkzuBvc1EkbE/tEDdHJvsJVWJEwyuSROX9JG+vvYeQfGaJWkBFS22y4VXTHmrKR4bVH1ntfRU4I
GV5hI0ZmEXvCQVa0fpwjS3iUaPDAANsDM4Cvi1Qp1pqoMFjC+Y2bszx2woYQ51GYZ299WFltKTLm
1X5vUbEM1OHHDpMIW9LV+7jfHnUmqXYBC+zCiXV3GlSSg6feTSEGOFDv0q6Xzz1bOUIXfj3IDXtR
QC/PNDgbFYGlH0NWfTBanXilHxDW7mzhV6J43VDnX8xb4F0BTuckF+/7O3+2h3bbiS+8TSGWEhgF
dQ95zxQS6z6y3OnhnV5hm7C0skfK/ZEjbN5SpkRah2roOyCW/UMR8+dq1HMfS6Hw7uz8SN+5AkNR
fagE3KeR/pk71OHo8rilHAr7eNXshdiuc7N6z+FYBqzgqpWj6ojnC2ONIo1ixnErWF/xybte+VNk
rkt4UmfKwTD8oKSHiYhA56Gw90xhH9H4FzQ3SNlbjJ42PrKtq3pQdYgtNxEbLX7ykXzC4yE5IY95
awRPU+fndqyJkyGX2t0djeu8f8eVcbnum6hlcaTXU5jgUJRhBrJ76JSf7c+TkAJn6Jivh5Xr6oE+
g41MSc9YpSvyj054/LykZuqumzj7bXxdN4iyniYcqY6uuYned+8T4z9oTKu2pGdwLpR2Kbt6YbCg
EbxcOXqRJL5nIrXfdZkQX/YbQSrqM4f0PajbdCpUegCRir7hARvF066arpNvrao6w7F8n2Kb3wND
edbNWx8Fu4MjefUBhylvY0HBi+Uu9pXorAYSsKSmunBBcdZruryTxqd+H70VjnPKTiLOtPmDY/KO
0rD4sjTPT7NhfHSd/z5NVPwAbLOWukB/xZvPSrcJVVNXKBQPUB0VdCHX8F3sa+ANJgElZ/D8Yo6/
tysBghht2ASheKb2eFZx9uOiFj0HeGdJdljkB3R9cLEnwT5Eu99h6zkglRDbYeFmsLc+PTfuRsZ9
ukWpchCBX21yWjwTVEhSM0RWtNgZIJw8lq7x4J8K59UX7BQ4/jSTEpNVVJcUtKSjC59spQlexIYG
HaU94hHWWld3cWv5oD/rZGphZDiXtgS9kmuGP12Ytia3lY+VlPbA1TQkvvRbB5QM9siTMULnM4/H
tc6e/X7/SPUFETWBNpZnGoYlsgOWAPg0qRxz0VDTXpYYbdBr/rn4PLX+gSy+KEsyeWt3jrPlqyfN
MgPgx4Y31kzx8ZBiXQG6a4tEvzWqIM1lDirfveyhK+yTNUbxf9mBjJ2blfae7ZBY/UItY27FpA+U
a+o8Frr357k/6wl95oF0Zr1KPJtSheiXCQWVk+FinJKemTlMupAfc2nw+QnxY+8eWVW9YLnFm3xc
aaAkVW89WCZZpJfOD+yetfwRjMPwPcrHMLMxd4Y62VT2m7E2W07X97xJmaff4ms33kV3ufLro3IH
jnZ2oKZVXLTMNr6xcswgJsVDjQyBEloFZqast1owy3xkGrX9GoVAheBzd9sYpZLIPx1//yxniXap
FAyKrBBkOxqcQsQ/ruvUip8Gdb5ZvybmUqIdn2naEjhWh2PzKT0arLptUEEYOi9p38Ckb4fej+4u
AOdsishhR/OukWSnApsltkzrgwus7BMGbd0v66/IFQuNjskcrmv3T7iLuKTzkErvYJI2gHNO0R/w
Yb3OvrTpHLO92fhqK+NAq7h31bKbi9YBpeJTqGkVnepvaaKmqI2rlHa84dqO/OfFXTnug7lCP4xq
pHLcryp9SXeeF6IecAPOw0VEn+lzfR1DEBx7sXERyPEKKn1kubGJLuysysS+c77bjZbZqI53mV2+
vGGYBKEfEiqC2MyTz/5H6Lx/DucOImh1deKuY2X5pv+RlLC7AqT+nMTLS3iRaFd05ggZMUkTvTQv
xvKL2CEeLsU0E5iXhUTIa0oPCkAs4AuHjOqtecoeFCOonWFuVDyKmHSRdl0HzwhWz1WN/bXO9FGc
i1Z4LkuU2nX2UhP109CgZ9VcbBWe5xBp85fyDGHKuVLC48RI+GtCAPABbdnTExha43YqVp/9M3kZ
Kix+u/kUbVHq0WdgpEVzQG0Bs09fkeSaRI3c95zCJmbYgeLb8xZp6QokYFoEtzQPao9OzKakWSDn
MJ507n449YMHSoGpXzIYkPbly9rLsnwk/VGfYeY9cI8wyMv/blpqXSzWhs2eiMoHcKhaxABE6EWP
ycXM7rOXcwC7wXzW24zoSbJlVEhuTyqbNjhZ1GEOKVRR7lliQycUPwBbRsdvBhLp1czO35yaH6oz
GWYeFaJrxFrEWfVx4ne/Z9lEoMyQ7F9/uqyungmnoHtmU9qX8ei38ZnwUyCQIsaUY0TmgqHBXE4Q
ZqTjGqEvohFwPGQ3W6w6BFC4zaEitXD5/GwRCDvtfpOwXWUcHFZKDEi5cIHdrFsnLpwCpe6z4K4+
RLD3ykjzMggWkAmW03j7sS0uvtmgS4dQ38PNmT1PfJ/ZmAhkYzDLEwShT/ssGyQR2+NCRU9f5VLN
TFSmzuTjTSFUmXsRH1xYNxFZXGiwwErFsdMA87X60cKR4eEU1uBvETlW/NZw0dIRHVjeVBTG6Cy8
IgwviAzTaTCE9u7WRpIyDObs8Mv/iupwOvbrsnMNTbT5CEmafp+049kktacUp/Si/ETFz7ojga0Y
uqxYZ+JX8aL21bEPDJwL2AuXE7zH7sDV8N26hHrC0WollucrX6Xm0e7fMVOxXS4v2i6sxgOILIB4
1fjewsrJ2pbTlOEyBNVnjnTqQf+Op8+WB4rxkIow/LyB5EweHEPakOrAgZMatVO8z/Hbis1hYWYz
uIkIID2f09QzO0tvmRbdx/mpHcFF0UYacX+42qCHJvxNe3lrT3kxnUU9DvKlFsN01/nxYEGOLQQ8
EHo4xpttfmqmQ2z55/JmdpeWuOI+BOO2keDD/Ma3N+rMJ/AuYKOWetLDVeBKkeObQ4Jb8UPGxhCa
1k01n4C7I2Y9+bclKoykhw/3NHeL0FEj7Vv3qocpnHZD4ynG5WQL9OtqckugxLsH8j1XXx40OAXr
3kcC6QAo8CucXSTmdSx1BLn4KtrJKS6QWsvw9sACNgjaMTO0M/TjcpK7QVbILBlgPo9azzneKdu/
E81BgB9w6N2kiSWBtjpCTK4xPMeAmsQYnn6QQxwxaW1XeaV6VP/0jR+QpSnK55IvnkbhPNGhgBja
7vRnGzQQBrVDIjPeZzWenEq5ZTgDlyc1nozTiY4kAJmDXQp9CkqlyYZlkwlATqNRz5wuNy85a6Gi
6jsil7qve/PMMve7EmqKWH6OhGSWAbLW6s+imKFphbJaV5xfUgk5LlInC00i46+Y18oLM/gPw/gN
+z42vfK56XRbCUjB8KpDMuKSEbho78P2LSuUFHiyxFwjBpLOAvFbhicd+sz3ziYE0M+e4kX0DKO/
wcXPY8Tg0fDl0C7ADQPSyYJlqOhGhIWRZ4+xpA+qO9Mlaxpw4jEGyVERad94HIoftnzTqlqeLLvZ
zJqc6Axgkk5nnKfSx/ZwCXHf2+UJyQIEtW0nN8LHxEQwcKCsusb4RH38Y18NufqhBoCdPfTrjjcQ
o3xiPiKcm2VOrTFrn9xo0cOPKyJSU+SWRq1IIlR+FtTQxySlVBnPnSMagRpHKBcio/PYmEPZ63LH
CS+Fqbj3QDfuwU6NOOJ1bREPxsCLZ7pW2KrqXyi3kJnW6pAS/68ii0pncUQnOks1BK+khvEqp6Cf
zKjFEYpNOu3/95QMS4k1naNoQkCGxllKYvFjFvO00dGEWIzB+Q/SWfXCZ4YRwMilqHxpJGaS0D4B
I7LaZieS6qPgM+nfld8UFl/vYT6uOKGWyhRBLZsjme9eOV6x0VbLwgln1puvc0prrgpDgBdDn/fZ
YH+KW4K/uVCsdHM6clbbpXND/urmvMdcg//Le9//6t451C9H9juUQP8355KZ9l438dJVGbY0qHnk
CB+W3eiEAbXTD2Y5eYt9ea/nCDaUKCQ/sQlwKF6hDWsUd+aIMZhVEBRAXXtrw1Ftsj5WdUVxDG/F
CZGk5YC5bBnPjOa4tGrbSVmmgFkLPlAdS+OWyPZ3LPYsWqQGzntIonQUWyUhj3sMDt4FUYC6k5wY
tuvMcPId6OnmS8KYHfrOh6uoq/lcbsNkU+Z+93SA5Yg4o3wF2Q/cNqKK+Dic+gnscyZk92Nte+/w
3pL6Z4hLS3YYrru2Ci0OytYAT6WXhPV0WTImK4qs/S5QSzkCV0Smqp2Rg+B2r4qtEJQ4Yva2kxvG
KgcmtSEGvZCwvQS+DAyXXoU3qbhL8UZ6JF9DaFszLqIo4BETB8IuFrCoeKiqcTj56Qs2tJSAOHC5
iAFPMSpS2z1+2SCkWyYcOJW29WqADs2/o66T9hbHnSeRRACIwz7qXqbBIqPlOJ5EAGKkLIu1csEi
UmFouU1EDZRP9znxGAQXg3fUDCtGCl0cDMleCRgIEFQ+snvrW/EoQct2XHsmZvc+Wo8Ymn7RfZwI
pvGpABQOc1OtNMG4GfLOoD3hFOAZLBsrsWz2//Zc/0VNjnJ+sqkAIPjuqQofoUYg++y/0XXd/1sq
CuaCaZjHO2guBVrVf0YlhvCpAGpLJEmSnAzyu2dzzNkJcS65XGu/FKSX/giDh3VN3bmvXvlDntB3
eZ2ENMWYL6X7AT6JOkeuqfTxR+MXXipUehwvnsif0uqvUcx6w9E2D7mMDk36Q3mUISnlsnnWltnp
U2xL1c+gChhigkahb3p4kYFfhs0VbnNM0L0ZRTxF45IM5UOV6KiMfX9IlIsbbTmqD0Be6HCSof90
9V615FuvH5kME6+IrhSimU9FIz/L0qeNpBaY1NLgXlO7zG4dRVykEtPKKK8Je+1/1AYLFXCUf6dM
sK3apM6X9ZKtyz+ihGYeHyHLo4JyPYZi24/rtfADuRyE92+BmdGcZb+e76wWtu40/CvzAxPmlwG9
X/kzB5+zdwWEdF6QEkHL58qybvjNfkbE4H/JX9QWmnH2cT2hKanxHWR63kjGDZFPWTGo51sFyu4t
+LHFatrSwVXLV1eFEfR1kR7ADjiizxoMBTqYgnWu/BFCAigh9Ptu9dbTKNCG342I9nq4Qm/XeqQj
jHyOzdwvx0Cl0pP4M6NT/60mWU4NEK1vB/jJPsqK0U0cLLEgY3BaGD8RoGFwe7LJRhdhq6Psnwg+
yVbgJIBN8T0OFu5ynYAsvDVKcqEu26ps+w/vdTePj+My528hnmQ1xbsEZteqEHOJYKbxUonMUMbQ
M8WamFWuDimrri8lDn5GEKsvk1nkS9g59skRXc/lLBKP9ELX3+dhhvWRcosKPNBIJgP/BQW2524x
shu3sn0DCHBLpfbF92Cvf96dbdhi9Wvv4XcDmM2giIkeNFRQHgxgUNB++1e7RFd9WJuPwCUTOIYN
/1643YcPV8YyUY0DhijowtmLYJ1pcmiQpa0AHS2IlcwoClv7osI1QWXDdPmBZV3s7C7Zzovafd0V
Es9WkLzERKehbuJxDNHcz9H7M8MnFHxKVd7C4Nc2wpuf3rrJ9MN8WGmGXjXXXmMwyWve7vg0w4Y6
EO/1AE8VhnCnMeGJJX6AoI04cjLrzo2DE30Y693uzPfvCIqI9dyU6YQe7fMb+Ex2nechQb1KvWis
dj67O1nz7Su/IlLYWwQZObfGm3WnS6M6j1JODzjnNL9n+UN4wHV6h1iAhpl0EswVahgqrPzbAnIy
pVYvK61TF2bL2VfxhVQUyHjxpUU+IcJQ3zBU1EIqO/1lbH7L21QecbqrxnHsn4UyI+e5wIhoZPMu
K7qKzhgdS55gYtfop+OxBPJQfHn6w4/uWNaQlibdGpe3lvdfMXKABwMpyCa/0bjDmPSiaok48tga
o15bslUezNnizfh489OOO3RUdYSMjjG2FdyYXWxhZR2j4Y5TNYcuLb2OgeVHkKTBnAr97ePCrFwq
kgDgNxU14m3IdPcYfxiflNG86hLtUh3O+vIXW4AwEuytVpfCSMiqTfQm4IoDcXLju0YwhN4ZGR4O
8GWaXX+ATDE5g/PyzjqcErLKOpIVFxaSq6cB6FLK6W6raBHHPEjIPKr7DS7ajCIXIu+vZUbXFC4z
RblOxN/QygvrgCf/840ZNPDHI7YTVsoiAGHDJnuE+3e1R+FoDaEph5yADg1o/px4HUcoXTzWuaws
xTWmcnzuK01tYjFPbim9uiiB6SdCmKQEn9AZucNAvbhzADwTf45RPzO42XxsGvk4Qy/uI4Byt4cF
H24mQOg8eH1+AD30JgkW0hQov0rdRHljZFY46UUnJqElms8ba8bpGArLAEDcUUmQhOzlDA2bvOIi
KkcqclaCGYhlN/H/2It5LZNvYDPecPVkIkeZi6nnFofoYtk/nZpYWDan1aA5DTfJf384kd/puprV
WQrKK9ZB8f2+Ik66BR+Bdd3RvwmyK6zwv0VyUrgMMj7FtVnz+dj/Tfvt+ddgoaGNdFNeVrCVqQt2
0Ossj0hewq7Rmz/UD3j8cHsetWMdEHCJE6bYRezuY22hoTRD5bPAXWvIKPBqzDecxia8i2cIsPz5
zZTq82+fszvMHINOfbLQEUI0I6I34hlpIBf+84NhE9xQyE1jYhqsNsrBGS8HSWuvUKMy65nleLMW
N+3X/pGU6MYIilb4r102W00FXPiDdgUJOz9eaHo5wjY6IHkQOJVhR/EcbUfM8g9RhwgpuFBErvkC
W5E6ubeb5JHYDJKr48x8X+zjwccAce3ZlW84B5aed2XGtKpAm8yO60L0hpc9dvwUJ/2SF5nNBi2y
zsSr0E5pl2oi1lNDjdOgzLDY3a0pwpr5rzrycKCH3v1BwtohBz0e6jJIiV7FeJ93sSheYBaF1hed
wJ19uQPG/tPBRikAspMgJh4Pg8XfYSHR98QY1NlVtMVun+m65ItWSNiSFdXvQ8xBJpnb5FSFa/12
8kYGA5Z8GGShHvq6xsxIlq6pB1V6Ek7XBEvgvugNwvuRhb+ilBDYXaWbz20IVMvWYNBW6l20HdDb
NCr6p0gVvyVW6Y4DEMzqtNJ/LZv1eyOFLa3vjqTK6KDLQdVKYSV5RrmrOCN7WuSLZyN+/aRP36KB
J6TZsZeVjBAPMu/gg2JVxsfaz0ln8L6kSMpIimOhk/8g96YmXuAB6NbBUD2fUCFs4Qi4DQ1VaK+s
8qPKm0RGPHsmz5FzDdu9Nks5i3Yez1KjtCa/xIAKhy+4jdkL9Y5B89xA5wcSkkXOblgkWkCtU21B
F43+qmW58MGx6tTldKgL6KzBWlEtvx3vOyjQOfyabyXLY4GQ9AyPYASEfm84CScRH1xqzKzbkmJa
sAmxK7KneBxyH+zYVjQcJdQTtnXXTP5MEJra6z+pN8WJtm3GygTuEKw9nGZmu8OtDxN7AGU1al5q
r9W9h2BLulrqE7evIi6vtsfeUwngQfvOUYSsSS0IJWIA8mx/fbzhchBYPEcYttuRgqcyHw1cekM2
pxObVhWTTlqZcBafkgPgBqBTybFC+nzH/nG21yY80vnk2xhHtTJQjS83c5NgQqAoVPzmGRu8Rf0U
aLKoeBwcBlt806OzrYoicfQb+NNZYtvtQN3WRBgD0Vtt7wKeYKmgzSDeBTV9iQOJASrVeWfQ8ywK
jbMUyi6yJVH3UYKO0t2WScEQKgG0N0SxV1rddVPSW55i8NVIfozCqEhWTOjhQidwrBZ1Tq9a93kM
G2JBfgbDL5VDl9DDke+PwsncBtU1jV0KKe82puKZ3U7Rb80qkJjYMo84xzRrtih7QHiEmnR4STOX
9FZyswom/6qwIjRE8iViFf0sKbTry5Z+tCqiUa6LzWbISjb3+qpxLSMUt+9awJpagP3V/zKGxXUH
ZGROJYeqmYk5Y5Mph+Lp2xBurFZrJxvhYhCcRhuArsT6IcGdVZj8zdOg3s6gLqk5/KMIYluUJxFK
NUaLzTAmoVD9/okEE4u03pBjY5ZayM6H0SdzZEuhL2Q2AjH3ro5utCxpvyUBBifymgyZfbwsojoB
rKaf/lrC/5i8v/SBUbMFQdSUugGWuKGdjqlQNS7tLZrjY04oDwk3hLiIRbp1ICvw7l+1FtbQFDJ4
gNXpgui4+tPJbSQlXV/7epJdgiXDZxaIAGEP0UhNZp/7CX78J5qKCF3+lK0c+/lQZkAZ5WoqSNwZ
VPaGxehYuc/yRXVbRLLV99cCNK4o6INxNsQSeFrc6whuRmOz4a93OnxQw7841+qlUOd7pdxUB2h3
3ygbfD3NxyNOB6sEWTKx427EQUbQWCj2MfkrF9Waj6CONlRmj7DuO27u5J1maMSNIYN6XswZwKZz
TN1o9sOdVn+RvXvXrep8jdRW5oI/yhq2mrwZfon5AuSu4ZRzF7asGIfKS4E+tnPT8bS5x5g1iuUC
cnR7KUtynfuN8tewPNjpnpFes2n4QlfZo2EhRxDkCi9aYF966t1qixHTkOuUFf1UN1fX8BzVd2A7
5WEfXe0Kf2ZhQGJYH2arxQQ6nyoA0LsYJbrpQrFENv3thWeIOAQMd7Vxi7+jmbLSQoCrxtaoinAF
MxFD9j/EvwMXxBVIbo4yJq9opPiN8ArS6MgubCMIHT4xMHV9V/9IPB2DxVZ9zLRbjhXLqoCgIFjT
TTHpIshOzivk2DMlyetkEFnda2/2z8q63anks120pOe7YictG/7lu/xD3K2XWnJJMMex5lZ2m5lt
e5ez0B/c2DmZtps62nnLzRbwmV0qJc2cZB1S9QpYAQi+YlPjsP8rkdMG0KYxJ0uYFcW3pNh/GIcH
emcIGmFpVpp9LMjUh0KgplmhnGM/rKt7MbDOeS5Svnw6ozAtPkVtHJitWqpe5H20L6+o61JhJf6Q
hERgoBbwQ8qvcKQT85XE9Q3Y6igyGabtDUAxpXVxcVnkz0K4zTE0XZ3t9A8Gh5GWMX+DP31urLkL
bMoZ0ludSi0b6jDRiSdisQeNDtViz/l8oYafH2GvJEKOx+ktvxiFR/ISWFMMhgzqAX+LODl/FP5D
v3udaQV3MSjfmSIl0s2tnoLYmWfZs8FFpOIC2DRzvPp2GwJ/wzG3C8jSdORElsC5KXWWbItw6m0o
IRHvaPAAnhMPMLLoiwlElD5P2TjEaKMT4jsdUOdVVRbWtqfaWjQz8xIFeryDbuoVj9kz5GoT6uLY
15YhRY/RMl5sxQZqaWIa97AXA+KWiJvsfuGcAdkpHUv1xf6v4XMvLDRPknjpy845L7XJbQl2O0NG
9VNDVl5dae62JyxEUvkIo7MGNyJKUOK0oiv5vRNw4J9L6gaRffUAnwRcJkV3STIR0oL2f1bJFTgj
ztBMjtda4Km8jo0jq4F8fcLhDZ+vUJy6obhQy6p3T0/B6wMZB95R8RflGni2JzLuFI+NKNnseUSd
0JO19l5N2dArYxvxWV8VSSuL/i3Hp2jDBipezN7IUR2L2F4wwb+UTVSMztk2TXjtRx3HLtdTbi++
hIWIX9IKZQxQErV39clMkL1w91zeGoMwDCUXeZ8UUfbZCRel1cUDnZt1zU6V1FmhIf4+MEc6C2ad
yNpVUMPRQu3Sq/Xf2zD5UaHLJC8SAwkBavZn92Z2FmIDvznlVZax7mNIetZ4oHejxMQdfZU74g+J
TeNMNGuZOPRaPTCA1XsoYjAL6P8XaRYhvePNkDT7D9MRdSp/dHoCeKefjKaaKGXBlVY1TWAD4K08
sErdo4lVMlGtTHXvsS0Tckgqs5vGjOJDx1vCtJQgZKnz6Os3qOTY+6KPOKOu1dVwkhJQbPilkd9l
c8q2KfbfV0GUK4g75RWQP0QhY1qs/mba/d2B69mf3MYd21gfJ9eQ9lG+FzWWc3p8wkmxSh5+PzEY
oloQDqxByQhI2UkIjqdrqYMskWgYfXoI0FpsnMEWFtQRbkhpX0KS7ev0AxtzvdQWw1BKzjisDky4
pE0Lwtj7BfmY44YVESzAi5vGmgMssvaOqS6S2DtHs5gVJvLweNTSxwZyd6wCRLJTDEDB7gwwJeJJ
gRGXxcgQNHfiaa+k2PoAXMogzaGHoySAy1jlJc1IYl2W9IqkjaOWiG8wqHEAbhhWnUZHUBsqluG6
RiI4qZJ6Qm88zxhiAg1fGda3ojQcjsKOb8OvW1c2P4u6ZhBTeKv9npt1b86Ci4g3rAH6myzfUuqp
CoLWwcQ+jsIQFLmh+blmYjCQ32FfGJ16jj/qbyjpuKsCK70KX2ek+6I6ov7YYu8xItJsyAkdbBgq
ze0LAUEQL0ZGyIp+pbdSsF0Gi/qDROH+8ymBbVeII9peePhQNkINbyLOZbrS3QimGGJ99YHARXHy
decxRYzkbdIPP+ou+lXGRvcHWenr6Wpme9MemtF+SVexresLeUihuH1P/yYglXh+Jr5W4BpbyDXi
kmYQxJU0IhqlQ179rU0sStJpPnKz7iV8ei8kBQj3xgp39l+/mWnxLxaCT/lsVn8Htjx7/Djr8+mp
KCcOdfEXw/ofUSVe8mzHkvQZdUsXfJ3NaDOISAEn01RS2gRhNYdiOzcxhnKqSPwTEHvzT1PVoUMA
v8uPyu7AqrQU3AwElj39fPv+Q268VETBKgV2Nq5Hh29mu81rfTWnBlkBosK66O8r8tJPWr9FAkQE
c12dG9dkiUObsuLqCPmffVaV5MSyuaNcWSOCt2tunYjtYD0uKo5tDk5AjiJr0Ef/A4ucE+mwGPtQ
ZCNHpQGVYhp5EHlzApSFewkILSGi3w00ONQNqYyzMijXdWQs0dUhzlwZsQ5azrjweLLejTR/yy/Z
yDDrbiAD6Pxr4SBVi9HcGQ8FjiVBZ6f8D8J05/7EynwEyQfH3OrF/8AqnPMBzxCG1gxQGbqm39qT
Iea4XmSwYxsIXNrE/Yr2T98S1hWt1tacO4aOmThWdDrJ+mR5f2vR4Wi37hWZhRg2rCNyIs5s67O5
/XSA1PJR23mMaiFnw1DhMg7NjGxHs2WSj6qnF+FrOXw1Ce9AQ5NqGeVx4muSCl2mIOhQPaUE4POf
ygjNhHvr7s9sv8u+wod0VGSYFWYTwkO8KbmDTLspUig60enhCRfuN2zQwUzWUYFy1YE29QXcesiS
a68aAxgCLyK9M1GZmbno4sdy0fye1LKxz4gzTPyF5SskRhUyVOmkrwhZTiVoTDibuw8jfWkdTZsa
5vhD1wmVdWwcPmGxe6K3olBhrZj5mA1kYhvhcnCmze8MRYZPIhq5Xt5vtpEMZ3Ql3gz0wFtGf1yj
xxVfP9D6/VBN3ICwvsFwsMXgOtt8xJ52DAOcOhH9ASE5C7Mg9ToELJUC6pRVOKrWWo+mp4rC9yO+
YW8OCB1IT/TMPsHtY1YoRnRTGLM9EVTu4+p/PzwHzAQTsLUX0JMji53L50OilF0hLIIyRF0zvT8P
SqaBCZuMr8nXxsCqcP1RsHl4oIEodTkACZ1WA96spDmcu5Y9lC+sLWyxmYbtPlrLy6aIhnoioWXm
gDc6h82Hyt2OWLTaAuw0XlT4tQ0JwQDIr5kR0WLfx2jqCIrgjZv+QIQ9M83yRhfOsbhx1UDih5up
XhyE32uWak3hzjbQ8V5/ZOAHX/qNn/18MwwM5hccMX97+nUX+Bcha3UUyGgYP0Pm6X3Vm/dbq3K1
8R/Dbcv5ezg41vO02nBnBliclQNGH+l2SAkT6RItEuWN9U8xDHFWMlI8nHuSbALSVQNwKdybZqfn
xwy/X1uDBFOw4G7PUVtjSBTV039OAbla5w4PHxHzrVovjcgE1qwR87HBWq/gXmwMI0lSUB/vrtyP
0FPZMt2B+lMrDc8b+D04/AthgRteCVeWhhAQOIB5n8EXf5uEiIztBm5BCLcfXJsGd6kmKP54Dnzl
0yMdu1Kp6/vjCGz95wlK7d04m2/NWC5uVRVYL5rTWEroBMbOQOZJcGkzlJM8jdSrTH/Ik92oPLDJ
beFOPGSnQ58B5CpIL1Hx/piwNKx8qQ055vzDOaISJbnq6O5LVSAJn4YU4oIcLYSvR44hbHsQRzZf
Zslu7Sfjs0Yne+5J+umw0F2/A3J9bIZNpKjB1UQIonCqUQkdtz1iVMfEp5wlURQJBwvHHSacDF1P
upOBnl34K5hJD+ZvZEFby3XOe964Sbux9KzEJBRwesEn11ijRIZxXMouhtCNbFo85xsgM17yODfC
9rshCbOxEmzDs7xTzkcmhInTQUDqD7d2vlphoS9Z4kYjji9H0ANXXd5UeSnJpc4fsAGj+spZ0Xnz
25N5XgKtQpYk+MrMOREMzc9empG9+mlUyiECI9ZrTBDgYny9/GzkM4uHlSea4ZCUP90j1b81V1IM
wPYn+1gmAMoAIVBfgH7QuXpluYRB2PDWOGOM1ZiTB/YKabYe0bYw3JxV5fmWv01Rsaa54b/DZrx+
vG7TDsaera9+b1FFduRZdpzfjn7MLIPjzwgCnL9TuHjGn8ICBMaBfC2SwZoDkifZOKWfNTF+7D7D
tKw52KhwzCqkWnhOHCBdqtdo5OmvnXucaBFcmEHGhWGsqdatv7RZIhF1yC6JO+zwJe+/Y+uxuOs7
5CSxrXcCUSCjNSfL0O58XIOX9tDExGPPAb5U7xQ29vdwsLWGbJ8rzZtjScFsjpDXapnYWHe/nDRr
xRh7GIaMM3dS/1QM52SqfPdAJH/uHm5ytrRtFychsgFiZVFRg7En2tSftC/NrZ5DBkcvdFnIt4iA
iKvAVDegLp6m8UpVtstkPPGJqUq/YKwIqocC2+FgRWD5Jj64zDdf9T91SyiuKmPd0g8by3VWaHwt
SFoNYRTeEP6hlPMcrssjgFELMcNhPR29yYM+3BqXg38G3J6lEG2NkChg7m2w4HSk6c7ZzamRojV1
y1HE0P21nQwI/TUn2zQ0n2fZ9LuWYPyJ6urGeQAMbB2R2QL4bZQ5rYbn/lRBsNt1pilFASQ3Gjwv
e82Jh8E/CgzTo1cO0GrEa8myowcrXIbYoiSS1qy2EaiAI84bx8pNaXXU0+tTYxe7Sc1TK8Hge2Xm
A84FjhtCku8/1rIduxqxXpXfzeMRAFE7X7Ta7qQaTK2J4C80ZLxhwDFTg3wvttqpPV/7i0rlGlXu
jrzzAsLBf24menBOHrVU5aiVVgCcH4pwcatHD0UDNBhhgxP7Ak4TBMunfbxJMc9ftyvUQITRct4L
Xe+tuAcKLLo0IhCbepUu4lFpLRG2bHF7isZf0wCY1nWPOvC9MMV6iliLjTp+bDuCVZ6NH5fU3i0X
+USPikYFLsP9ZRrdamhaTcUcEODbyJi63IumTvltEfSj1H7lFI6gWE1hZuMqc4U43yxxFQYLXgSv
J4vixUZa7Lkw5P9MeoqRExeqCRHQg84og0CdnDaVaGLuwNvTQ3PozXr7bW7StP+0AuXsvMsO9JM9
AJrJl/6HS812zExJGLp8Y4BiJFsBjcDVCz9rNXYbk3WjuN9jSpDCziINOSLjPI0ryvypkOvHLytb
hnIgNXHi+ONi1CysK9tltfKuUXjePN8d+BlD0xN2nfli/lmLSrL2lUPB5FGJ1yxJgsuOAUEaaDEX
/9KeSWCNjrFwk4/QlhEGGECGB9RYAAPX2Xgl2tlZQBMpCIQnr4BNl+92ZKp85vgMGEbyBbZJJfVl
RCp1EYOC6g9yed+8iDVNQQzmkK3Os9ZnW7i377OpANi3BWA5UkWkGQBik2OXhnaLzi8mnOSjKeKx
JT8YFfxtH6shl5ZXNDHLPHlien7IGdEgU/Ov3jLCvSV2p0e0+2ijreZTB5fQ4qAXVz0EDl3xBKDe
Ng63DmLDB1C8AG1T7S5kLyJWLNkGugxU82Fsy+8tIa2j0wRqN8+PxDqnfpGMkAnUNCh1uemRYBop
NBUrhexojd2gTeCXEk+mqbRYRqg6wEx5Ta4xCgByTfgqfWYHiEEYOwX6pArLLkAAralEPQkfzEbm
gOgs2qVyHCEtbAt7MW6vRcbYwgkfGv2odLKluj8fPOsc3wjPWsrNGtKgaP+sEWtEcHElpdf30lpC
2xWs2BGvpVmLsjFQbzfF/R0PTGfBCqnee+AUAfyY6aqbm/kTh/CfJMvVcurv/ChwrC0hRni6Us97
D07epSieyudZcIs+1piaaLRl9PDha69N/YFplbyrsdiSayv06oVu8AIDoGc8CbtYuBQMJkE8iYFU
dwWUgHp5LbRrInr+XSOmSS6P3hkDwTsX5sIlKVf62sXxM4MN3ZanM6eQ1NJgQQKB7ztBNOnp4t/4
heB4lu0lCFwWBYDPH9hJoRexJwjgJT9zKcBh7wAAT5Xi5TfrqDnQ2tLxOX6RCOY5NKdKoo5nhyX7
SavFaVQp9bqjMsILD/T8ZNyCF5I326Uv5Xw5JA0As0hgWoE9PTQEO6PQAz2nwMNtjQXdM7oxJn/y
uxsd+l8qql+dY7G/cEzvhKNohdfrYNqpbzFmSmivNhoA2fTCxsatxKGq5hgY6kMLaHNNh1xCxDK0
HDJVFr4rzFrJddzDgB9UtDl+wbMWAz4y+oQpTeKCQXAapaTfSMJGIEXezYvXDZBFbYrX/KZOMmQq
uZOqgqE2Ukk02FK69/ow9dIv+xB6PofsKwXSgPRq2N7xenIpSoHr1/15B+fMsTx300hEG+HKxxU1
RwAJ6Dzqr3HEuounbZZ6+CfSgEABVWBXncvpjut5KLsLJue+sFXF0f6yOYCkUXL9KAbyHpi+Co6U
qnTFmZAUNx5f2CO2BOaJtnY3/dP/iu2lFzkncXXThNMf9+hskIJcvhl+2AFYQ1Mdo0kPEKkNk1/n
eNLWaiB3skmpBZH9ITg9tlcd8cvH3Ii9BnkJ1m2EK32+QH6B17ogayf08tYk36ue4n7eZWeTkOcb
xiuKCuyH7AXCx7Y3iN1TWJnPV1Rulk7M16N2PhPcyHC3Xy/ER80d/qozUEXuxsR05h9n5tpO49bt
HCg8JCmK/kod6aPhGeVHcZAKWSFNQ+76hAnhotnJ/2FKIKZHiVRuIhcmdB0V+8L7g+moOnMSVODQ
/OmFlIuW9NGf/MKJ1OCYokPWgP7eCRIuswQdOjreHHj3vDTbydVHsTRlUMPStcO4DZJeJf066aON
2wGTqtURFmpXGcbEesRoX1O/ObyHyiEv9rbQ4AItAYCFJdAm6dkyJlUXuK6dxQwFKxyZzRkSNvGE
vbuER+y/pgGuV2zUo/YA5ZOwZ0KfqLfT03salT8St6C0Ry+eQEDq5JtSTySSRnr3IH75WvRVIpOW
pIJpSxTW8LmL1qbiABuzQGUhV/iiNtxE3IV0etQMfdBhiy4dFQrh4rqAzy0BCYhqfbbXc+6V1EyQ
WEvd+OceAyAdSIPhuHDQlf1WkP296XBiVltjdG/H+E9R7iIO/L/n+dMeI+to5tegg/eWJdIx3Z9Z
RL1LDUFm7b1r4LxUp7jVae4YkzI7P+n8V1I+GUISDpvRQQ3oeDjhPGHwUFV0g7TD6mtSLF71FEjP
+WN8jzeFjLTdQOgtR6mOFSU0nxoIEsrdNW8VezJN8WLhRWx42oyIbcu4R9/HDmctJUq5/3Obym00
JERScwuB4Sw8wdV+WIqPLZiTHPLZjhF/FBG3azoMnzMilSnghcqOVQGL3b51xoPbWWukLuqDkobc
CcgUXCMq5/oKhxilltQdnRCeR9w4dhgS8ICAKGDSwIDm+zfadhhabFMc3VjudCsu8hbBH7ssaPUU
94hJyFn20/PMfXxj3iz2hrPqkap4lfdrteXnMIXYbGnPiU06sEYo3PuELOIZxm1ivQFEtCIWDItw
FbPkK5hpjrSU9ekZmqxZpZDMbezlBzUPtIyPwUlohSwLpXFt1Q3jj2ztFgwBlkHtGdvRa2fERviL
mwuCPykfyZ2npXMF3L2coVPON/FjGBFxLYtKX+3jq5NixkkSmrNFZ8y6LN8lKPpDaG5DUUfCEmEN
k600RCefAHDNRYVv9izQxI0vSoTjljb1d1KWav8PlgWtFwChERBNOkJyk0RaqC2fITTfFrzl9A2r
jfACMdO7uY8S7ZyTCiqmbw+Sgo+igltrqbJpgXEw5ozI8QcTxTxlZ8z6M667rwNetAjpVfkAzS5h
DOeC1fnr8ycImuETMq9Y+INloQJtp3oegohol4HjOyk6DdYqmPf9NGtC4IYy4BkTMcOYWNclTFuk
OQ+xNw0D/1NsB094jiPFriOKwpVGzW/B5V8mfUPRqhUBc8gfBVcrFiVGaYTsb6ZfZa1FPc9UUejJ
5n21jBN+Sn02IHItpfbINe5pxPUH7GuzQakvLkThCRhlTcPN/5y356llhabSVlpgzTZBvM+kkutr
LW6154IKVKUccznMh5klWtGApn3hewAq0eRMYR9ySZMy3esdza4qQ+uC/wvXGS3Dv0MJuudLw313
YqTkM47ZPWnQzF2YvcFYbT98H54aCBGGG4ISyHUeAwbcxQLkU1mDYbTWwvfSYO3qYDlwA2Aa/AzH
+5s3Hx8jTXLVLERp+mKya4KWgHf3FN2MmgrNB4SuUnblgquHY9NlDsCeA7eWxyo08WceU6QkvVjO
A15zqWlLPcC3g7apDwOWC5b+yDN29/VtH804PFChbv1zcDwQ8Sa/Ew2telad4vusHsWmn+ersghQ
zXygMlgVwoy/D7nMeJswciW2tXR0RivsLfJklnBlKjE31DPl48e5uW6YqmqR2JvtuxLlWKrpTkFs
XAVm+h7SayGAsGIeLG3NMucyM7IVOfPUkHJ1o3yBHaBgDPIfQZMHs6GVSdACDawuZSHkxLAKnixw
wwRKikNBixv23zlZOsfFByUEhQhdnMpt8CHAmXkE4ZmLjQaDIgSBI3EBD/ulQCsJvjWtZnUV//hs
Alf7wejwMVVV5+dHKycvAVYI76p0gOYoXh/coj8TuVDOsUaksgtkQZgxugXStlvcxsP4cJx5qBtv
HjNt97BXjv1giBnq/F3QuCLHCeeXf6g5UDt4N0uXWb7yRU5ynSaZCHumuYNCxfZpetNFhWMlixaS
rZUChxA1goGd3f1a3KarsoXEOAvOH/BkflhMcNF6Sm06F0DnuhKAumLnvdLCsSwM1QoNk34UCTN5
JfKyQb+uPgyVxoWVnNPSsKw9Mxf37mtZ2PB6iR/X2/qDF7BkMqEsG2nSCe/M2YGMkdYMTkxXayjL
kfNKE8RozmH9q4mpzaS0ARo6SgNIOXgvHolOewR+ebWKa7UDwaQlWtovVMn16jCDjgyouZLfX+8+
pjktJZePwR5WdKoMPvd8L09jO8pY9ZyXp85nQAHC9WNEfI8KaNySKOva4aHOe42p96MSb1xh0hFk
txy/gBOwjkt5rw8SCjS9Fu5fb0WfXIHEb/OBxr86Eis68bceDMlyVwe0GhX2kA5idj+Ula221y6a
PambGJajqOT3P/Ec5hpYe0dsTEBL9wcz8fNTHbnFP6XvCXL0AYjmqWHDvil+IdP+V7d3f7B4x9rG
PLCI9rok/C3ol6YTnScsPaxvfpuUDXMO8kSUnRDAxGK+lJT8B65nfARRX0droigpzIdKrXIrHxLO
+rd8ld2mKMMaUPEj/PBdvY9kWLGmn6aTzaOXIal6N9J8jiWOhAjFFA91Q9qBIZtFcf1katCbHfmT
N7oY8wfhc/ct56E6F/HX+0zIvLDd7gMQAevlkXx+F35behZiXf2J96cRpeh1u05dlCbWfEZWuOuE
SZEzyWwqcYPyMzfYABIfkO/JGOnzqw6Sp/0hB4JdJd23pC15oQJJ9SfzlIOQzcMV/jksaAVPRaYi
fJyEk9x7V8lH6OKFdgObTtVVGziP8q9wVOUp3bSekuSBGd6atyU1Sypewv0Nb3fhqv9r86vhgYlz
sM/Xtu+rSFkO148qNiPhuFdIQKcQlKAj/ZweUo/OauV4M875Xvr2Es4XKmfJu0AZYS819LNhoKwi
G1sTqRGbkTWH/NkCkb9Qbs4vLN/6HaVJ6MAtCGvGLA2j7JdV7A5LcBmYgtTcPmSXRdEygSdcXMuc
CkJsqrUABNyZnXtZt33yqnaRGpckWxXL1maS/wdTXvgrUVzU8KkqPzpebnTJ/OMmCc8wSRCym1N5
T0SggsRVAAzbwPeD8AvzcKkG5Zd2UN/CSGxDswR2ntzPUrWrvBIk5VVH3TjVQufv99Q/YO2eM/7G
Nf6R9e1CB78cLp3R2oTnZ2qJmlizPNZBH9qrnoXKwGLBnCymmGmHkStjT2hDTAGknG3heskpadhJ
5xo68JUXg0FUQ8ut/+wOIcIrxb2PqhqRnLE8v/42MvSqWU//DYn4ehmtdXzTvbpP5moc9tYNxp03
SxHJp66buFvpkIp/UmKLLGk6ZgJyYkvb96AGfrnGa3WP8073eebdRbtBR2zeCkknecRy4QSiFWvJ
TLesb0SgzA0KbBg0wLMhQ+QDZPKtlrsVdV7S9TMGa3gJOvlRzGx6MFZOAhbMLK6p153+60p1XixS
f50P9129X7MphloelucRoR3iNIV8mcNSbanVWQcwJod652h4GwyEzKPbFbq+YbDz8wI5hC9tPUCM
1HgYyXKRrEQRTH3Ul1xMBmSQZSvJsC9qcMCss55noUBW1/tNAqIORiXLOGIrobcngtaQd0zdMUdg
Jza9Puv5Wq7XE74DxqKHgi1fl3iI+qinJ8wnsgpo7FjDDvSU/TT9fOIlqQeH+FWRc8Sf7R+Y2O/T
I+CojLCdQG/JLwamPfm5d5CwsFj8v0NT5KVL/3DYmAMx7yC+EmnlZsA1+OHWYKlN6pSMpu+ymNla
y1DVij1QPxmTITnBywYj+9Q6rqLiON7EnHHHrpmZpd3VS3h9OAW1K9CCp4d+HEyb0w5s/sgeWVPk
GbryTnRGnZ3ct0StF/fPHKVEY6jRI0HfUFgeJ5p9nsJKg6gMB6MUyfrM7lmmMXLf8PTdsloxjbSw
6ubCZLI0b9491h1rYesKPNG+CKeD/7pqQUknP2PYMVTmasL8Z+oJamL9zG+2um/an1JLjP8Y++jx
wxr76+/SrkdWoTUc2ehP4peeRgc3k+3TVAoW/D+HpzsUy+KWcUYsqMmGNXfxIuaX0GDZQjEnDi+I
EBZGLW71tofh7Bj2J8pQHeyLzVEJi+lxtrNVC8OS3JKzymtC92OG7gKpOqb+YA6ZAFyigoVGiDzm
oFi2nV9+eYiNe4qxoXdm8pArVaR5nhkVkwUjh4tVZvZ0CZJ8KKClUwJBe39F55z+yvZsy4znfzeh
D9xVcOHMw6Be7xQMsHTjk5adk/v355tnBsaotaASATRpjhDH1OS4RNVajF56fe4B+6HSZoBk/L8y
fmyMPpDLrKfTOFQIjQRgiSIRk3BVdiCpCQFrHdhAQMgeVlbjUOT3+hSbu4L+VVHL6SJG7iAg6sgL
4DaSDjt2gb3iuxIdQl0uhU19aEfZJbIPDbTc5OOKYMeTagj4FWSmwr/AXHWsVtptrzMwT8jOo9VR
YQCLR8li0/yuYvCxoZ4w0dCsau/wccnsopDA+cP0wxA+ZTxr77vMm8caQpgpfmm9SBwJFQ8uOxPT
zaCqqcB1hqDlQjupS0lOrF97rRBcWuLIyAD9XamwHXQOcPepk0Zy3IzLe8Uf0ToVmvEIOTQj8Yub
1C6Y6/ac4I89NUJ9cg3cywv3iXpNsZ2fB3c9DjLzQdkynvERs81hhaOjfHVGPBvZyqVR3lQyvoH+
yVeZYBmS8MNTXosqDZVqln5OxhR2ntA67R5Ui1gEr2jz5nrd32NceV618JmGZAErpXtMCFtkaQn2
IRAHInopRAx1vfrJkD/rlOWHkqs7oKLTIFfvKV8jg/WK9Zn3tkzHbdhJ9nrZ/KEuwiyOMRKh9wBo
S+v/OzOyiLyl9x1LSaiNMmB3g8Dh7noel/ibIXGvJPwC9nZyCI3L1hqkj+yWX53u9PhSCMjeltk7
D5zbUEd4Jntkr76L8MXqsJ5HJp8JFslbQRHsDwYF9n3WarbbhzGToPY4oveNkGaORlnNtkIQmZPk
7CJzwHmCeJBGUSM7ylTTCmqImyc6Ydk7Jz4UPukf0/ovCyNlqpDU3k7n5bpwGxJ5+hnfI6y3uyQz
vQDJPNXLFCT0rBJMjawxEIBcqaWoYT7NE/u+3HOFvRkTAnWvCKoKO3wQgP8mUr0kCLtsIesXx6xT
AAJh+tYqIPpMTDimgj+wUqRrPiQ2U1iKN8TbYC/YalRVAPSX/9aqHw4lD1koeCqyQ/k7O75hUC+S
Y/Qc9rbopwMLXzpcjjlk5JJBqQS0CW+4JJFHFbFA+nIScoKFpmJfdWW9KmWdDfBboNLVlYGnyzCc
gcj8WJ2en/43nUSf2DzfANC5A47nJf5QkwwRGw4HF6EXNnQDLVAPHiganIDlM55CjCkFivmMyI09
gYAV0SbcYE3szUnwThXZ2q/Oav4K+yqKec+CPhnAObcA6J7KlFsSRzmdmqm4THx4jokhkomJUQyJ
TE3sjUleDE4mLhOEBToPG9Yu9c3Ztr1iJVukGXWCujcH6qUeivvzonCj9cAlL6nMxLCWv4OOwqRB
6LGJTg6E1cAuAN78FR0Lqn4W8bo2+LE7qzpBNSCu735G86qgmwyPPL1Nk+UyHwSOte8Gj/FGFwd7
J+iqfOY7HRNWTSUZUXUHyQVyJjU+yWuVavp8d8dzZiIxOH3gWYvgrFlbxC/LVhkZcn609ayCqR+R
3hHGaFwwytLUYfkxSDWv2rbc8Yhif/bBMoxog2246FmxVlReN22FzlX5y2/nslIu2SMNdgJ4d569
Py0e6DSNmB7sD/Z99d3Src6nVyKpka2ke/RDm/mADQk12ZXq5tmoxoAfUB1cp//Jrg5iJdq+KQY9
koz+baSP1xuU58vfTXGB06uj1xj2Qrpoo7JumPOvRVphRPl+wEHvoCczJbUFeYF1ROBouUbkyJA1
6HfX1zxEFVr8sAed61fE9RQ/dYa73K24sZY8z1aGR6hhQmBdOCNE3f3DqEpIKfbYlkerMcci+gpl
Nm/qkC5z+q8TNMw2av0jSnDUEbBq5pxXKlAYzo8eNPMi7RqGLBlvQVd9wPEHqsclI69elIPurFv0
kSlEVyoqKdLQioEm+QzAgDU31RMj1l4Ozj8MsRkw5gZuNeect8iRdsOAMsOPQ9YGXXwS23/qatrX
jecwUGRjtgcc9BDfSynhEOgTYxQRh3CVmuWRVoHG+eSzFXSDPDXR944K1SPiq106htSxFrEn5GFu
cRz1NMHuQYLakAFi397YTEnsyBzYLZV1t5VHy/RTDqCxfT3EDy5QyBOJ2o3/rzYtjNdqJuOrPT5b
ZR5wI85Ln8QYRPPkg2h9m+6Z0WR62JI392fkrgDiSj6X+JbCNq7611ZFFadGnwApmqhZaP0T6Uwe
iJze2vKGMHCf5It7za8dE4c55dt4COdflI1VlSrGY27Q50erISDQ+O6Dbvj7vTaI6qkJ9WOpZShm
IaDcK+IrHMvwRrJDNkJEmzMf4eJEnxhul/IS5gw6/Fef5aCBkbVylIgtMPzOgWShvlV42fo6jQ+v
LuRANdPv3zEFlx20Sy3aJEJ/FKxwdh2Q7SDl2I8IFb1CG93o45y6ugPPjojx1xGgSeyqkUiN0s1b
+wTiTHOZS0bPL+prXPxwHXtXzfhgjFX0wgQjjd5paUtESKb/RSUa8h/rY1GQg/C0EoANbgIAuIKv
kTPIAAsW1qC50+CcfHZY57FOnvXuXh1eLYkYwVg4sVUifv6MVgqtBxneB9xw7xZfCuUe6qCiJhlB
Rf07OkzqY4Koeo7yI5JsbFf96grflE81rdcZJTBKcU9IZknQP3ZdD18FV/oTV8GHdWrBjBzG9ylh
NmlvtnAgMAUhI6gD6NXa1WvqQWrjERKJUx+lh1ymSnjl4Ob/m0OZuWodCOhtOhUeW1kyEK9zgu67
SdfOScMSSmf/4PSPHbzFOUlyLAlTxoqpSpe4pBd7MauVP+CnJ34vFMgNSn00fyH87iw57KajcUh3
SLIEna6f/BXLGRNVTY70vplcWBKDNzris1zhy72uzNbL8xjWPCjaorlpoMWvalL+dPVyPSbz44Bd
TXoNgbdPTlnw7SjvdxRm3k05OuZeRRGzuxsJr93uNQ2UqbdoPYstdSilAeIRdvr2Wvnnsj+39g8y
MMRReROgePtoIfZOqD/Sxo2GjxFbHgSTdV/bhS2jD/i+9wpZ+NCVl+z8o++3iZfJkeqvBZUzn1pg
LxCsuEg8fvHQYy7kFMQ/yls1U4lDVOqXkh56yRfErcx6MfCYtYmBUoZQgsJE+/s5JtBPyKU83xpS
HsTWoQKCg0EOwMRYhc72nZoJzkNLkA4Dz7t4VWsAvpKgg1hYvmHA2iJdR4tkAzegE5t0lrYm3eF7
HNKFPsgum/qe7o5C9ZKpTijpu51REE5cm1Vadkt1/3AjYXHi/gCt3Jgw2D3yywQphZeaDKtIAMV/
ElmfkIlLtbHpGFggR0s0qWS5tU9gMkfewBwDJpfFERKZ8+LzFHi+y1y1cPtpeDvAx82ftoyoq8Zg
rY479afxlqXKqE48zVoTl2nyZnE2LMvSaQd5giefzoo6IwbNeFOX/45T6yti0AJ9uOBJSwhqWd5K
spnqKfJec/Gj4fwWHMtBUwXIzAI+Cnh8gJ8pMy47IeTtwq96pnqAk5jAQwBRRf8LzWkiJvhOe3bK
mplnElrXvxj1apoWoSeCpmMDbtBrmcukPNH5FiLSjLYKix+xHCHVXLkmgk7uURNAPAUGJ6gqZMEp
LaNuEQVSamykpv5It0Q1teFjVeXOzHqpiYF1CkQuilnETxakuN0NBr5U9XsPr2lyij8FpQ/k4pMx
bTT38A0OKC6tomde0jlVpHO2SWVdNgAGmboQzOZQruOTxtUjI2GJbubGVok1AHs5+E1c7GL9OS8W
/GgiKLWkmGzXOU7Jie5qDkRC95lEV/Og7UctMdlf9YM6trWhxc+PPESPR9VsrqViYYCap7QT/+qj
KnKZDFhy4GOwd27sG1hn57ZIzgUB3gomUD5pNbxe19uWT9HHmpSqP1DPGXQWf8nOeSshv+9eSMC/
Z92maYY22Ylg6Oo1NhUTASs3mdxEkyVM4ta6h4xLRANaZ2SZiiOsIzlxhuJo0AL4/oqIAJuB9Nrs
qleH0+r33xCHhIdnNuueq0CWuaOghLg1c9wsljK0fcZYQ8QMPm7tV/iNGIiOR6+zhylRfegvPCME
sQXWX9+IS4uXKI0JeWMncCqghOrgVBU5S1bZIJi7IW7pZUqZAcKt5JHhBMsTZ3j7mihtKJA9BSxM
p1BRKK578A5Xfj2pwbkjlbuDyWpIUciP+wKAo4GJ2fjZwJ5+Pa/b6N97Gx538qBSuTW6lJ1W9WwY
w3MEy7/h6Oh2dkBLRJLy5zmf2KplaaCsKQaHcLma5Bxus5Ta51KoU/rVeJ61ItMKW/o+uBXioKpB
z69dO3RIlTz92GkLptAHCUtjExwrQCzz0gmJcrCiTFgbuL5ablIFE88u7yXAopb2lNaLwRFFB+Fk
yQRT/F23K2sbZz/KJ2qf6vnSRx5yIhZcHsEYaCwUcOK7+mBUaUQVv902VqfzL5SKbjp0TT7wx0v6
OnuHmQ38+XOFzENq7iYVSnI22IFQNY84TBtU+wBxVYf40YYgZK1pspQ9u3GvdoJaXSA6FZRtqrt7
z5lVsK2WuVs84kbavZZiIU3wIAB14M9DOONa+ehcpRJTkgKBdsWvsZQWmwa5qmmbsbz8ncklc8wZ
MXcdr+Fq8MZ32IE/E0YyoPu+/YWzWWlKkt9Sdyugi2Qk5jEecBUI8tkrO1aYcN03cEM8Te3DZZ/a
U6xYstjkJAkOWZN4HMAphcM2iSeVqy00WXC7M+4n6rLI4sXl6ht2BKGNAinipUcVkO66kZyK1uGD
4wWtEadVAE0vvsduiP0g1T7neSKuR331hFjjmGVqj0ydm1Fwa8Ce0TgWXmzgPxFlyajHEHsQHIId
pqnBbwuHBDZeabSftNxUBI/++JHG1r8hNIQ0uDPzur8E8Jbij5+ktXuC2P9v/vXoyHa0NR08jNNt
kiRdFAW8HLnRTx3qufZv7eTLNPEIfGDO4LhP6rxCb7IKpYZVXClYPKvzULRvMtE94pdOc1TB2Pw1
K0h3xfRd5Jz9RtS4rCEySNgENU8NA0L6FZ/bEl2hi3repbg4SwSKNlzD2SxUnjQA/Hz7NCqAr7Fe
Hgib/U2YLxhE/Efa9YKmps17DwXrcbVq/cJS07xG+ABzKqw7dmfl8425UABkvMNBH7W2cxBrWPuS
JFaNWVAB1Ou6InJCNjQX0/lxnvtmmZlObeiV4ys66Yn15PQQIEihnPZt+lM6yotSKaLaf936ke86
wGGVQ6Ogt5mRMHXGlH8j9XRikEITSCz4Y7iwG+0QBr8LE8dUEpFkdMvySuzSVXEwTI0GghwR3ov/
id7KUXL/YJsobNIeoSNL4yk8BphOqr9ulqql3E5475G0eSn6Iwu67VR2sjysc6Qdv7yx0pBw7zfx
aSRRtedtb6AkUF0T419EjwiRRU90W7EAmLxTsr6baSfZnQhvQdctlVE8tN30AGCqwhLNVSjnMuqm
QmxsSiWYek0vjeBliB4wNOUcj6q82+aoJNTTBmznyQf1rjOXqR+SSAobK1D5PDALNhHF9R5CzWgj
IQQeOUwLnHw8uHL97qlLGdRZ3UZgHBih9Yr+C0CbT+7+8jDXqG+hbel9c867z2WdTjwJvaVmbf6d
p0J1oEb2Uv96U+recj0vXeHfHjvOBT0KW8E5erGh5s5m2Vty4BhIjH95t4ISmeSdpisyEGOMVyy6
rX+gn7HcBz9lgpwxlj0/Q86GHAh+CjCpsUKNrFSbWdzDXuq0gOPzaH2mvmjqJqcJmVEfWezPIluZ
w6BNdcExzb5hOU7bQxkrLJpqCEF6CVAzqj+IZtVcK4Pl1ITSnrVUl6WCnm68QMvX5M9GDFigKlGb
NtZEmzGzBDuyaNUUaaLysQKRaxwJyf1r1ZI1xSVOTm2C8Aj2LBLkQeFsCkshVtNSTeSGsUdWx6tc
hMREWAGP38Ki0pKnvQPhKHcO8byrA88UrSetGa0qDGq3gogla8b3y2SJ0GpMgGBZzN7LQiy8rs9N
HZDjtg421VIg7x7SstQd02lh6/HotkrKXDnZzzu0WQ2o8CF+p4YWf+dsRXdZZ8mVJ5g0soYSmEXu
Cj0JMrueue5/sdHVRH9SwQtxtn6ZwC2TvARg8faJHH1mxeEywt9RE9Fju39cqv+7o+ZZnOoqMuk9
uYZMwyaJcjE2tkHxvhr4e9kB+gDYYDSi7TOYfO3fEu0D8NPr17u8Ao7GkjSbOh0z/ab1wvHmjjCI
vfl9ulaoMz83J5tWtVP0AuzToCBL6hUDmUmGKFTKkN5gSAyozDdsnfUiiRLAqXZ/doDRJDR6LpLc
1yHiKVutsTXXKeFQkld8COQAm+IzJ1J2zKTTfGY9flML970hs4EMhiBOfI2hjmMHdgf0cPQG+q5r
hLPCPrif/kukJ9dg0GrI+De1Vp8Hb4FOmyCCugeP3HdGjOAwQwBcYaB/ZpNTx4XKUf+nl+vDP6Ze
RhisZgeUdLOWptlVSlwJhRvpM8QWFgtOjHgKEtKb/wLMHz12Eks1VaqeKoLxDE0n+vWszlcWrZ8V
LKU0OxEsJUZh9ZDTwExUv0hm5pC11ICc7v/eSiVw/4thc4/V9bb7TG5UKXE87FR648d7pUC0W6wK
kxNQ2TpBnWde4pU/DeT4BdrFpfu6Ei2nw59ot/ajQA9Ibm0BAHOygc3JW0vtjn/riD8lzqZt0nJB
vGLpIZ1vXiOGofvAivh5q+5oHuuVRpOGQsTAZSWQk/A2HAegh9PVJajIjbqaZPT5pubho3Xravvh
SbZaAU8lxZMELu717GQPoqTpgDLAay+kVK8S5BQ59MdLSG3R1uIQUNg3nnKC4qTxlV5tmUjALue+
6c4hb90CS/JrLxSvlkAS4kBqTKAK/5LiC5JYd31yj+WbYXnWRhQljNlI2OMH6SeqOhzd3BXmx1Tk
QmU5ZQhm0QYZvOVNEV4bK7MVlHxJ1Ynijljt8sxfY+1m+vvhOIu86JCkJLmuv9KotCb6tccDHtvg
hH+HfJrV5rBl27Wcs9SXOGKSlVfrIcD28R6Qtt6Il1mU8glE6oZXsK3qPgcx1wOcQPwORrKT+Rao
sPZPD0cbJkXF97NTcKQrn5KIF/PlB3MO4HbKtzZmA9UkWW3EG1w1TMp6weyIsE03GaHZ6lMotrP6
AKzNht5KbV1nJiBC1/mzYe6vzvVQt1cvJqb8S4/l7ybLTdyY6EFkheD5bwDX9pzM7KSqdon4eTYS
zj/wQYBpbGbOCgaewo9ePgusdPJbOKPGjwyjDgzOY9UTgBTS4FtQsuwJ8pJJGEoiHB/nKnm14gVv
H0eY8FNgnnc02O8ejAtvPv42evCvyuuZ5LmUiSfQKJ1SoD4AplNkiLtz8JTwiLegXxrAFN2xDuGN
D9eolvwBS07DX+ZTF8guz7Ta7CPsFUZe0MM4XwkihOrc82H4/C4C2J0/2b8KV/YTyM8cG4OOcwAk
Zxr0ynVssR/olHRjh0BLO7AH1Y6I7JKguQ1zhRHNGCksGFEKiXV1Np41m27tWLEQXLFbU+HF7XIr
acgJyB1tdDCFGwod4hDkvHL/xsf97aVQznjbYwwrT9w0NOglGvFbSc67YVwqMXxGlF+EEry8WOWo
/CEwDHz+b/itdege9Rn5bKMGpQ8lYVUptnECqUypGroQCVSRBUKDBPRKfnDqzId6tnB9jbogDgRE
KQ6hlyaGrGmlmD7Qj62hj1xjd7G0vYFagARFQ+ODh9JBP7oguPFUKNU9yShNPG9XdL3yQNxpWISt
clMJDqlfsfipXYWo4QYxzWWfNMxMPQiYQsF4uWSfJrJA2AbxYg/t2hcLVsqjLdBUsxmqxO8UnjYZ
ieQX9JChfihXKYDirWPn3eT3HN6ycpOuEahB1olgmmfgwg0g/2taxkvZUJjJPJqD9J9/7plN+xSJ
+WncDV7eXDBLIsfwFXdAcSgxponcUs+JRAhgKu8K67wNxRuu6hDPvpf+AMFSjOGoCWd+NePZDV77
xsdEScsdspiw3JF/lCJLq2YrqMBB2aNS637YgBPFpVkhD2WjQpOtqKmePZhgxS7Cjp9N21YQiFoa
d4IM/4D7qPe8mSOagBqtLOzKol0DT9iDfRB20QCSHYOXHoYAT1kpQmfpXJ2dYa7HK4iD5vkLkCoT
cBEntXeSTVjjSfd1eiDs1X+M2iTrTMT/QtYcct5XJjoQ8PnwiFRV38Vlzklh9tZmWTL7lNhqiwfC
HC4Be5EtMHaE35V5P0refSV3AgrhRQDHsEHUxQJXaIylgiEtsrjiPFT2rQQZ61AdJAV85n8eBvEB
CT+ul3T/hbb6ueXOZ3JZqzMp50mafTCyMSzVgCNoPISzhwOrXD1RnZWIKDg89UJv5HVltdIfy1k8
sicIh3PMAKRvuEyUQDjL0BSCYwxPFdRUQ9oxNKciDn1B/8lBd0qw994b0Yu2hJWstf/J8MQ9EoR0
ulsmr1rvuovojVbd8ix8xE2zyOuqKe9gsbKcgWHUlPDCEdFauGz9/gCXzcUZCd8u5FvIzRG2345u
cQX5bV0lu7p2tk6EIbl/7mwW3jk0/wx/zb+gJmw4ES63JbajoH9nii4mNE5Db6LGuzmn2ES8uWMc
/pYMA8nNVZQ9WT7WLLngfd8rHyXWTsJxC/+J+UIkw60hBbMEPnjGi5Ifhvxfh2Uil67wmwUs4vGz
WbMkhyxZ5+Ie8p63FeBq8wc62Ta3NRBHPsQw+3doiL2euupEw4oamhS37lk4oLle6TFktZ8tOpt2
c3aUyDjFvldtinAQu8IOcah0GSz5QoSjhTeEhtAWiZabFNFiPs91XCtsOGkrLnJclDobjtE5e6Dd
kzZVMwI+arC+Kpg17WPyyuk2xlpDF5x3Zb8mAVTju1Jx3PQo0qOleY7rsdgef6W1dyoKjqJSLcxZ
H6ETbKVwCKNZb9MiP4Ewbo9oxa+Wvlrh/QBJFtIPLF3+C4aAvpGR1PPUOHmEYhblTeYPlL9+atIB
FnOuRPulJeP838ZUbUbMZFbcV9OHqP9iVkzkpg6aVlLMHKMZQBhQAV0E96Zcvz4pT0Srnp4Jzfem
13kfDU2T48+9/ammSJgaH3BXVk7yLZr9ZfgAp7Ilx5S2pcaiGi022DzkT/sV9PkT5eE5FAoked97
jbJhgxol8TQqRhTrBwSs/B0TA/oMrzdglF+3bFkqcfeoI1lVbvlOz8yA9YPjjKYss2WSFQ9ZsusD
GvjEw4eqUhSSHoDuc2w3Hy6SinUOjY7DUS68/urltOw3uWbZqzJZqru31BMm1OL7cXDBbdAPVO8+
F7t6Ecueot16qrInqsdEHYcYAMlo7grlT7CQuVEfdZUHAEwfz2/QiyeGTCZZP7sm7VwxB5LGQ1sK
6GsgHmgQt/h0DzAzdv4sHLyE3+bw170PWf1cxwYz3ZOsaBDcs+M5Ewk+PNSPHcO/cO+6ax4OCV7f
+MwfZmP3msJW2qzTvPVJhHtkhXyquFspO+OvCeZ407RsSwyOdnMtAFeICq4TXVaSXBDfW681jNbB
wvQh4XuWN2H/wlgdTiTkY0SCpV1/E7JS/iARoZIb/p1BxnX5QY+fG4HTKmUHwvok0zeFnap/PdCF
Dce27bAJ1ULRux8xjjYng8vwgQcO8cfDySK3y/FFq5TNvrDaXjvVGy7ey3OYziVEDtYeHV4LC/wq
ZVeVTPU4x9+RiC6LKxzD3LMIhhtwV91MbKaPTlYILClugwObePeskuvoqNe2o61XbpfkvH7OVyWW
NmUoMVbIUihwnHzLEveVczV3KqOnTYN5Jd0bVXNA93dqkXByLj2GN29QLqY21EsBVvJYpM53AcmH
46Mpwia4kA2KNLG30CsVSCAxEJWseUerewvypJ6e/lBjrpWKoQJTQZHqz2xUQGHXRZ8oprifMX44
ugh6BPoANLJ2//v9MPPK0qE8+vcTz4QicBteflCZnq7bpNFyRnty6ijWnJX2pt6bdcKodRYZ8ZYB
yeq16rdOvYDY0cC6r+ixgyuZZUnbd5S98BtFKHh2B+7XRQIQtV1Rwuak1C7VS4i0kRw+immPM/HK
O2Wy4PjYR6MjumnI6zbAIqA3f6T3s8xijq1VEYcRObmo2Xo4X2SJtzwzoPKXAwK35Ydf4npaEFg4
BzwOa2TA7b6alh2YczokwodHThC+JF3guDQvWh4ZF3omP/nacAKZQGrPpujXFM5ZGOydTJ+J8GQQ
EC7tEIsYB6mKqcUQdgljPrm8m3uji7ZEP+1+CbOZRIKrOpJctKcc3AmlqOKuWfrCPkswIYp1mqqP
9aVcJ1Uod0s+Wyrp9Aufch4CDdZVB8DZ9kPQRRS8sTUco5xV0MsBGBCegwmS9rVrCUhxKZ/MdUrp
t3SE6gmeIUakfQ/kzFaS1+Z5+a9Ayv/C1NGMR0FAz/9AHpa83t2CKd/qRMzT+fQIehDqOGjlD9RH
6cq+os/IkXmIWvPtIi5nHEo8tPLrv5IY0ugJZOKNaP7jv7j9DGdiEfdUDaePOskBfmA/3hF8xfep
BQAWPhfkn1Tcgv6t4PZM+NIWULXFtLIB1Oo1rbKXGnNXofGAgGg4rxtemMQ3yBKI7TZkigP6jSvN
nvOkD/FCWmk3kSP6077EOXC2dBBb6Q0EDJS1aDXjA1B9hy5XAeQTW9gHdc08WTGSpa0IHgXHokyc
Veu4ZxeK5R7mKnZoXZEMpDU8GLFtszv7t4uPBCJI+6jKDqNCoZtAQFgq3SpMRZLp98ptExIc0rfa
z4ZOvYX9vgvKiBOjAEVuovK8HkAJTCbeINrNa6Qq7vY1yxq5RT95sKkNx8Ym3NZCD8rMFM+bAGhN
uVRIvJcZpOe5AlXS6nRT8hO+tE7/uodOMiH0ZP4Fhv6afN4p4PqEZDq4Pzmb5RCA7Axr25LLs6tq
ZVcx9bk7ytm0lz3VehyddQoQ37JOH1Dj0/F+/ezMUgkfZMlx//vbmxn61lgfOsAolQCMfAq9GzzY
FaFAIw2UE7zhwNt6BKeRZZ7WgonBv+GUaj9zkzeHfbPRdJxRej1+670Bob/t/03zhV7ArSPyQTDt
8QeBNj7TYYymGIjlEOylTQ1OVSRz1uCMheC3S3/k/WfrMJleUGfCd+ngvchb3i/bbbN0b6LKxn2L
blcYlN+8BjIKkrHaCRdaFiD2EWofKgYZNLY9U7sihsv8tkbx4Mc7N/tXFpIRlvNxU+BDjdpC3Slj
SqTOWeghRgsw4yCMWaiNrs5ZszuUJrAeJJ04qQ9JtEPY7sqqlxMY9JwppPd/vwoF5W17j9iH8EAE
HwaI+jOWOdzYKhaQhWvZ9KWuLBvp66y7JRbar/HcA0lE8i5VjUo57Nmr5ps53ZkQRItCClwT0oyB
N0hb21BWpuFHcvn6lQUTnPkPlneRiKyCTd91u59FkT0qyL5u5Xnx2LnESRa/1c42A+7FoBHPLDkv
W/8ka1ypcq+CKGKujXaKGBGXLbP3VWC0grC+VeUQdzdZaSFS5h6HFz4G7lMivsRYtkmyq6dqAxzM
+RgT29IL4YTO2/Ip3fgOLfM3oFaDdzQYubzqAgoZ+cNAmheeit8QFHmMWiuYIHFja3jspF5YJFP3
2QRPz+P6Ao4P24J3EEDbfK76Wtsa4Gbq4qR8RDa2kx/UtlaD708X6qtTaGkUGcvq88iuvPujUCf5
54RJhfgKHSfAhdOe5b5AyE0vZrgAmE/6HJ4yMRQoXfsAnIZcPeSmQZbZWxyqN+pFWMqH+McFFQbp
JDv8UXI5eJpA2ijlr4W8o11837qD2yNUhHNewJpSOr9DS7n6uynEBRu67k1MsKqz2SHXigR1yh0m
GWqNUKyjr5kpgWSul8pdb/f5i/+wG6TZzo/Jzvp/iLFJVd4TZx1gkOIJ3ktxl3Uy1pzGtB3TzVC1
Fz/n+Ca3nyYV1f7QiykPGjo64pKDp2zyy7/SX6KK87MyWu2alnyBcDWs2UzgoLaQvZr0N66vBYBz
YZDj+cfFJNvFvgjeKFwhZd6QHv8nuknyekihYpAbYCk4Ytqs5PsWWuj6p8ufsbCfQjnkjEsNxQ0S
1Q6+2ZF6JYx89cvU11XMMwgRUj0NTepaTyq5vGrxKBle0phGphVdXA5c4czB/FKFux0GVZkMVfJu
QUruIFrPp2C++N3kaaPwcAzxR/FsmdBuzRRagNe0ihE7oXIj8D9Z5Qcr6jKu6Ys7ncgLIzwNzWdM
RQ/DwfKpbmJRqQu/1Xt7udiP4lSc12z1tGmRwZElzL0nEF51+GWr+gD0inStD3kdqRM+1gIYbxzE
bRSFXCD6Uzj2G/OrToTNf5sfO1rLw8q57rR+SDtU1nNv9v14ufWg7vwt8anT9/p235EjK5FVy7y/
m7xcOhOwxys8NIGO6cd4g2IBCv1lZ70+5oiZF7mtnwEDimbJ8fOWpp9l5PqOJ9gbClplg1XViQuy
3VFR0gVB9qWGupW0PvomRpSM3999+gG7Qmm69Mpez0zMKGQH2ADxiGlXA2yRq3/aQIbmgBL68Jqp
LI2Z+6MDe+lpg6c5sPIdXrrCGLM1HUuea6vASF/Mi9IUXfw1ImJXNFQiYPVUijhYy4Ppztv8tob3
WqJdGp1Pnx5EDVMHILKfbpDVU1r9zjVuHfQ7L+K0OHIepY90l5blEHsqvbvZxfYiXEmc5vBSHhdk
7S19pmLQ4/5xbUdVcuApvSE2TFv4q8ZbHyYdeQPjCnenRVl84q95uig224mXGuRb2OpmbLUXASEU
F5xaVcAGDC3woxghwPVffXMuGWcAFsrjuAF7cunOzq9CsSNyygD58VelkVjjJqZI+3lVwftev9KS
2IAmKEZg26HbUE6TQDnu+gqU5Wrtsp1iHRZh3j2/4Vsfli5ywe9ScKqaWIH0PQe5ciQHIqs3umId
cVpizF0RQ2J70jNZlzO0Tzyli80jQm7nVCxo2cZkCPvVKRFAAauQXNBe00uVoQWzapNafweMvauc
HQvfethIpaWUqEWY6X9oV/7y4/HMK0Mdh/r5bSwzAShUW47hRT7tZgE8a1uCih+cFrziYW9FnNp3
mAnb5PRBjpkT1nSpALQC+dDjTF6DNfjJVz1qQfhBYpfG6UfBbpz57vu1ftwmRd24bTA4knQtAj7r
ly/m6jvKw0ckfnBdns9WfowIZwfGAVZh/gt74F10rP5J2UIGMKbfV3+EBD76Z06yNYKRpF/JcN5d
hHAxh40i3Mj/16P3/HHQfiWEB8EIXfnwrS8DeSdjB0QhuKePxI84QQf5LzjpTzG+Lt45xT6W9MJZ
f6MPy7rwAr8kaAp+qySGZQwLIvbDVeIdTlCXqltlD2Abh0tL7HpkMYD+cvZ1j/KAwlA6ZoMJKeMy
A6p9RZkfKnDhbkscc1crzatmffOjhPvpvuWxevKtZdL4X0LOLdLhOLqpwblE/10DrNJmNT/YLwKI
PHtt0No7BTi4DXwp1Im+IBtE5oq1mJVLr23Puro/oaronINLJm4zgCcXIHqshOgusDsihSLgwYQH
9XPDUR7u4PW0sv7QtZBH08sBRMHaBQMbLWfQc4cUwnyELtIYqos6nqTaeHBKNfVK4S3Pyjch5INn
9H4NE8xOUsd2izUDqxeX0X6RhyD/+rkYcRLbAbGd8KF+gOdEDm+TbZ5LfmenXVIQtwOGjE2rnDjo
LOaiQyO9HGAwk6JiwHSt+YCncEsGRiQQZsSO58CFhtPFtEaNWnpsI9y9LYq1WeBcvJpNoCwk7Z74
kq9AXoGD+MUojLo9efeX0jZu7+pODFLpAR4myLgB+xPeb38PUrh38jYA2ok7LDa1j2zGLaX8weFY
QukycfLK/rSIipxV+LJQOQIslqaR50iIYUxTWRNkQXBXlw57vpAy1Vnysk5ViCBZF1iZ8ivHCwcg
K2VZiiGe6hL/XwwjzB4GT/mdT32mIUS0u7CHjsr3+9axrCIXhuNwK5D97KXWMWMHEEu8JPwpLgb9
NFUwjhBFm6wXZxhp0oS9o/B3pFYvpxNwUldNITmM/QRfvla4uW7qYTZpnUZKOedRI4JoXEzvic4T
VT9w+caJRSWAB0IhEHqJHAYDidQMjCy6pjW10A677BuBlz8mLElF+DTFbw936AkVrj/iJjqB+SdM
TkFdosA0RA8l06ixUcmeo1BcbiqyX6niEUQ5Pmn78HUGuuyk6BJEzjOJaytfMrRDw/E+KQ+ROD0Y
1V0GqGDv4sMrpjB0V0iSbmM4oS7qZcCrQPIwPVwzMSQcPA00vJwlki4bSNMUxUrhd8yh7URNiy+v
ZWoVy989QMZe2PVNxa2uPUSWderL6QH5Zu0s/bvIDuNdb5eEghZNporxRa1eSCFgsV+vPgStCbvu
r1ZXj7LV3+Up0q1Rp0qjGBMIVpSCl8ifbZcqB8LW/yt4p1e3cOh0ziE/P8II8Gq8wu0CpXAibP1A
JdzZw2SRUUmC0LO0i5qwXVFshdmL3pzvOYVswJLfrKjm5n0f9T1AqO+j1tSKTWbONtIfrjW5eTHr
td81dQ2rz93eo6Ig33RfI8T2Z9rSoRUktcnE0yNJhKgLYJ7gT3K8MRjNSn4dyatq+G9JMH4j+RWd
QrVp0utqvaohb0JkujwLI7h4W5tufT4yamRvqeKJV385hvIbg0LC2urMgbpgbiNTv6i+7Y1ZZrLj
pUC/PMoxXgA9wQyCOBv6ulJnLNw7yAfZm9DkCz4nJAl2VEksWiu3bbhiPGb39nllNFPGr0ZHG8gt
Ot+0L5lLLjiyPDHL56zxrQ0SSBf7d39EEq55sLXjgC47Rq4WutN4RRECUNX7ywWTwE7ckYn9PqUe
wQzt/m+zqDwVsaPcRExRyBoMYmAoyrpOw9RhPY1o1SpBEspQdwYOU3tfJT19TYzVwYlDV/pPaN5S
5JB7eLn6IVyvxqJzdZbL34f2qX2RbRH7l07DhT9qjfJTT1dtfudMHvT9IGmJPYdBeBRMC1L9SsgV
hdQWeMjO6B/wd1BiNanyvqCp5X3P5+/U84pgbIT4fXjdNV+tDct+WtI303Vto0JukVxL/j/McQOc
BHE83dWmX/K+RIDJUEsWMJOtE6OWeFCuzr0k6fOyy1is0125SBgK+i1GRwrX4xcHPb0rtEV8t71V
EMxcGrqJBrKM2XPC7XWqXr2vqFBmmLxUByHhD9t2gIhF8EwY0DUyoEbEFgIsrT2mF7YkP9gpjMpW
1E8gc4CSIb4coPA2FbQmrKZHzorNGHdT+4SBnCFkCBCrIUBe8p47vrVsQZVNKhVk2ABZMdJ3Miut
zuAxVCPqzlUF80BRB3vGeuIwj/tLZ3Q0H9h61M2wuLf/WBOffNLtOnKaoWoOIcH6Yf3vBlaNLi7x
1MtsK8GgMiicGMZwYXZVAVojPydT+AP9nyrPNnlmLBPOX6cRb3CPO3K+jZIu7kpz0OmBXxU9qyMI
LlKdyMXEbZvlgFCA1m5MkTW/sdwGS3kHzAsSicRoi57q37FoDMX/jyiiVHOhoKTwc7sX2oCuogeh
U380/WKppf2Au1tvqsW3CHl/a/Ffo4iNXprOejr0lG2Z9HKykphGyJdEj0SlQsOmPD0FxEkbY93d
sBfF+KRtmpvQIpvpCz5nCVPEPTCQm1Ke2YqzeAcZPCiBfvZcy4fskqF9R0LqaEnNT9NEym9FWllS
9VIfk4nCpYV3bTOj40SPWD0NqZTQj20lFzTuq15ZS4IYSqCuh8UC+Cue/6Lkh6b2ElkIMBLoqZwE
STFyrQlK3YvoH9Se0/4s1IpKue+dkrOeR/PKTHMxY9oxoQL/+pp2TPRZv7svIEacdgwu6tLZw5MH
/fUvWgVU6+AKB8jumSKEZFjT18UFUuJFbTTPErzI3nryO2+mYVMAAA4mzVf7cI0bDZcJLfIShKrS
8BVFJlo0c9JzAy5M4zUSbAsYx6Hn146ACgP1yuUZL6Xli4f4M22YbZsaDD9mnp6mW847UV8ACOT9
1v+Qkmg/eo+nxliDPFVBOOyaVyP6PuHKdTOJhUdLYdYOfhJt/77TXyxaUVIPXiLXgk1kV7z+/KYc
626LYC5LRSK0n2GkujMR8zGFyOuEgSvq+QsJJvmDpRMkQ4xvy5W5j2Gj7nVOJDNmTQP2f2/PvkMH
trIdCdKIcFJyfpuVI4URKeZv3FmpDCsPcHoBhzKxHVnhad595/yoA3oaZO8TRoD0SoGHsD6H82Qi
w3ofoBzxy8qHLM02pL2QR7ru9Lxkz4eEjxvME9aVOrn6jqLCxKzYOoz7zVkoSPhfTbG1+4BXxiga
rJUecFZPerWRq/Q74fDvh+3wM6K5i4C3zXFSUelXaIZVgnHa2ZGQW6lFQq1Ut1WkeLrm5MTdpoy0
B3S3J96oAF4aJmtaTAHNREN6vyjfPvknTk6fURVtXiSCic683J8Usfir7cDrO/FNQohWYgZcbsOh
qIhpfHJO3OpnlUjKuZUstubsylXu7DFOefbhELMKh5iSfNRK4EvWhT1c2vXvKuY/BG4Jz+YMiIcY
Yn1VWF43xGK80OnA0EMqlo9fCDthlKKBFWRr1mJiSqbKpEiAjq4JhDQRS6C1L5PA5INSwNDCWVrk
p1fdf5kvLn4Cxecvv190vtVrhdd7TCieN7tos3uyxqH8ZJYA2EiluAn1mg6ZzaO5Soat0HcoS0tD
7LlLLIg9qDf/O8ApeftyINSIlPFe6R6slahITyO9BwJIMesflzf9m2mpEJebVTSBghQdBn2l7O0n
Mxc3WQoXBA+HJFnsgzHXxxF2BGLuWzE00EUGimdgdgzMwQDu7DrEa2RZqHfW0j5xAIKEEBe/YofD
YT74HrfX9P3uh9R3kjCAimZjzDUqw2bwqLBzrO/Kdooe7jVLh1JtG1mSxRZsLGYeWfNeVto+1Uny
5s1U5oGNQwpqkdZPPHpmgxT99XhVGfIHVXD3hOZgurVZtapM8rVx0kbKdM6gkOkZrXRF2OliMO+y
t7pMoxxwbDZdq85ZZ3ubsWvievKiAGKdUs0Xd7v3/yiD+HjdxuVTsu0n9fLxChDYrI/FZ+oyTSax
/undReKagI4sLZqnfFFqgnn4IsasrEr4nESfqDXPakiAqGUFoPUiGGaSZDui/EzXKFGvrEH3m8wD
qXf4DZ0b0b5/YJG8WEz2C7MMXfv+Gat/fV95em+71ei8JqzdJr0gu4uiCOTrff/iXOjGxYYRwsdy
u949YQJDuL4ndvbEizv+uuFQs5/lyAfQelENxXVqoEcaoX9H3HSBeJfGvkf2ERDni/hdm8OyTqbM
C9p/DNHZFDmeOog/01LflZW/pxrPHeW2IlVVbGbJisRSBfxUjYk/5UEiUEGY5UryghIdYrW3zuw8
dGEl0/0k/aAW5t+A6rgrej1vTKMTzNwUUn13shRoQ+/Ym+9Wx/MvTlHtOLNqJHcakcnj3/XfM4Oy
CW26FiV5Yixz/u2xY5f1+0nOlSBLj3WTct2Zue30mq8yas7n+QogBlS6IOdsa682qF+/aUs4WENj
/f/qeAgWrVOxp3W/C6GlZTWhlIP+7sNRDYt7Lg1gVh985WoJORlOvNP93GRnqcB437TO4aD2PxBZ
xZIUQ06rSuH8mt9GgscDhXyoHFodg3GyhqWXML9udr7diUjr93vhchmM7d/A8jFSErsf9Cx1e7m9
C73EQfacXNMtIOdYWAogICWF3e281pKSZc56toAPhE50A9Qjzx+DiMn5CEEPu9jTKvz1RarpGc22
lCjKwLOyyqDk0owsXOJEKCw7RngIoo3eS8qndzcVX1W31UbCSDDvHZHth/Bmi1FV2qg/JCbf79Kc
g+/JXVzTdx9ojVkIvr3QfPjYn9DZQyU9WgaHPqVrgWGxcFhZML8H0pz6/jzMUNytP+yPurGXf/Ta
d+ciiB+gy/Mb70gcchbSpzg6gVENNTk23recpvLRrKO9mkqbLUidSYs42Qd4jkN0fTK3RcilUVcQ
gKwYcsvUtcelHdODEvsEQ1mMMdGBGf8AW/y0lr4sJJ/aHRgIrRI8+yloVMsZWJh5WLceO5i/e6mW
0mjAH7aw9dkYhkgERsYyqZaVNiyYsbuS1cJ+txTcyw9gX+4Pmj8WxNXH9LhpYaRxTSagGTVKbUqZ
Ie+I6cYDwOsquZ+KVlEue5DLW3u4g3KhwNVc8lw6HP1LMp8g1lbE/NbPTFm8qi+70bd6PESqD8yJ
EIvVRD6EH0KHeENXXAODbenFKMgilDBHTdZxQwlRwiqpGaVOYfxOpv4eFB1DW+TI/BxDwHCruGeI
ywplQQtrUjXkfrOYT2TVKdrG0brIRGFUGbh1Nj3OrTyq9jxZc4TStYBmcIwexaTmmFDeykxTnNM5
1224bn6Pe6s6HRjnLuBENdlkm8h+EiwTUqDcdInW9dRsI6mNw+xDbjon6tIPPRJosDjUzRJoFNyo
/HkdGw286x5vgdp0uGrB+GZjJmoghDuGe+wqxcHf8Nj6HXNqUoej8Q329FheQNB495yeGc2Uqtgp
DePsLr7/rqvWDsIEybFX0M047K8lO0s/u32X7faz4peFLHclG3gG/UviH5v1rK8y6F8dBRdoq8YT
uXojR9oo2Oi7AZ/ntojX4Yrw8nuX5Ez+J7fY+uorvLtMJ5wtEN2cqjrkz1BjSNjhYXfqCcUk+O8i
eXvCN21NlSLxEO660lS6UKmJMCcs0D2wo63dsqd9VM6MyCT/mxD5BTheuQKqd1lnpZaJw+PjBLNP
A6gtmBPII+1lwbxkiJWKbZ6zCblpEY+kwAMCKeOV42HEOK1fitSUYikWt3sS/Yf6egLi4vOH4oNi
oqAprovbWppKQ1RuO2ekOjZ7g+YL95b8zDmxmgUgu9qTVx1KOfV3MEZ1KGHqYEOTw464lJ0kPTi0
so5q2TkAznrk3PwkeS9+VpOFq72K380vTqRahdOAtDMvfKjt1lKCNg0LCbXqmDulez72Nubqo8ih
Etai7L6o1Y1OyiHx62mM369lcxh4jtOUL8pG1SCNoy5QQOVxprpN98t7IPkPZfTvU0z2UvnrafsW
thCpuv74JE9cMne22DZxMtSA0KTPUJ3SknUvX6lTNIF0pgW9sayGFpzXSCFZ72EgcEAre/AIhWwp
ZANr8Z4emuBVAVN22b1ybZSxEKLnvrABhLkm7cnT7Jbm8yfYkEPN2alSGagBB2I6smSUMXPNjtZ8
So70+fMRTw3mLh8Bq90ZPklN+SlyTB72hcxnHu5M2rMTlVAuBSZWkXEMZcXo60qqUp/ex/mBj2WI
prxThxh6eH4vDUNnwaolxybAg6UEiWozypQK2vR1O1bqWuesTkecvwkGZ9G+ryp0kgQgM5rlb8pq
Rz8BCRKMfpMCfT/SwWCCP5lzbJ8+YX6TTepSPuCCvA9B2Q5eDrcaz0FpshR0nRr6kXx1i08HrhqB
TgSbcdNXKYdQ2Gm9AKgSjwfJOCS1orJccdTJBMnXZMdN2fuGmEYYnvNEnrqFKcf3TgNX5aUwXHOC
lBspEsQwlEJ0uihwgAz9JahfUNMzPW03G9FKe3UlvuxGowB+9OhAECzRKZV0g3n3GhXzcAuN6cjh
hGcFCyKzwYmbU+DZvQeZkNywkvs7w+HQbBaY7WioJ/gT2iydMaetKliee7+/qG0KXD/HuaLtZYsM
spwEovYajeInW71aBPF2Q3gZV87ZS018V5+Y/tzzk1A1WcbA3btZ770huSXYc9GDijLEzibDn75g
T+IyaPhPWviOwdUhIPjvPkHjC8+tpUgj0cUJE3qqlJnpkHGbUG7xh4cHBGv0T+LEEd4eUtGZoPdt
YZ1dXQKrU0fLxEFHL0NjKWxLFFIZ7SjgD9nMh0KS1b0XKjdRHdROxVUhQj5K+7hptyZX3zx2KRTG
AOGbo6fITZSUSkfg5lF37wzb+5vTPPMWJkfOmfY/LJ3PWEmsKcEXuzCgInK6RQkQPegc2SlESgHO
xBbEusJ8lF3IYtW1m/pIYs994V2d2d7Q6VMc4/qisfehleWxCUoE09Do4Jn0jLjSF/Bs3KSGXmK5
EatutkMNl59j0gLUYRK/sf9/PfRz44CbAL2VTObG7DLIgVOhgyMSlDwjWim8PtUKxqtIpO3MG/ur
q7qG/FVN8sBHuoVf4lFdaygL8/YIhTdfrlC6+zQIlFeEdrTJRaR4oeoNxA8ULIhDGnYfRucRwfY4
benxuxnQl2/YDrd4fJSvb+nwMQzlQ/wJfdxuUU8gckVDLj4PZ5hReXJZbzTLZCSmCCIKp7TvWxba
ue/lgxlOkFoZLMah8FJYE9OJYKfmcgs/zJWBlkvjweuTd4F6KDaqrZ4gb17dYRJFY099ShRbfMe8
jCAAHVZiEI3isdWuHgQIgOopX2FBhf3oRaMmSM6tqAaYmMxIDVGNjvcaFS7M4MMByq5pZves1DyP
aQYXg2yhvrBLLsUSivVSLquoyHwh2BFLC7zJLZxYQ86E1lqTSK4Oy2DE17XPci6L6n7lrvcEUMwU
k73F3MoBO6+Hk/BnSJlp/zqqY8Z9BSRe5W42m1WY/mq1TjlFnLLVEI0NLfoTkxatsWBXl81obRpy
HqDCnrsx/inESajyJc7CAybLu7vB1YYpfaGzmzdkZh/eMhCTI9ad/Hyywa9S805IBhNvhfKdujNC
dYScqwCcwyhHvNEam9o8UBPl5sqIMkBZiFz81kuTkkJSrrsJoKEKDBhrsVrwGi4KcSpGFGmHm1+a
MjJM5ETcEFfa9ZIRht0VJN3QZAgKs78YD51jF8R7nJ5/VqI0vNsgqr8INPOmMDUXLUoi7zcFv4cR
ueVMzIjjwQEAteESeK4audcdXYECzhSagqqt8byvC/VSPUktcB80LsrX4rObqoML9UfE9g9rlHOn
Dw4VE5XTteCQZ6hH7G0lhkGiYZfo+Yus/FT5qwiTBM39IEKxIUMmBp/TIhZ+PsSgNZZUuuIOvRrw
X48l9rcEholswBeur+T/JUacONbRJrREMnc8tpdwbbne92wAy5qmQytPgsGDsGJfwD05AZDG3Pco
r2+8J6wJGOYClLlWMZ9CAAW8Hx5HpTIAfs5MOlN2ee1Rlrl2Eu4IOCPtilArezajJ3ZsUtMkX6/p
Xh6Zlw6Kb5VdKCrfD8JfqFoCoF3T2v+MvA/lGnA05aDAmD4NyQojsNXaiYpIO03t+aZJSOIkFMGG
UPqWq9eWgHj4F6zdZWQDMPpT3xGNzaa5nWkHlIk5VVL0BTBlWnz+X9vtqAUH+lQPK2owzy0mj9l0
ptc1w9+SKJLKErsnkbhDU5JHCH98UKywQHGhByjDW5Vu0jMfzRx3vl/mZuFT1jh6KOlLBShfqx1b
6+sHzVvfNcPNH6MspvcZpGSIn4PbIE6a9TD+jh+B2OeEfspTr2cgxZ6rN8uXNuYmzMlCmzwUixnf
h5nKiQ8SOtfuX541dHwDUaeH3WF0RLlcrtrR5k1l8UFWUjLvzs9zCX/3p93ilQrgipCtF6PAwM2i
DfjKiWr+Kk2pLX0LzBAiUCfCkLmEjjtjydaisKwaAfk52yFOhC764XtXrlDOpTmg/Q52tEw5ckL/
ZUY5/S2k4XE1m1Zb9lVHsV19jCK0Fi65aH9gjpDYMv6LcSd0rab/fZ3U++AJkzIRA8NBwkBhYmtO
ejaYewFwlcKzL6HHsyAZrRl7NJEODRx8k7Dtx70yY/OZbErOIsrHRkWSXFbvC4DYcFjDVA5tGh5U
+NyQ4cUwM6GCByN2l8XSRFok0wdRPFpbzKKU14NtOCnHhbxt21Oow7K6GbUQT23nSqYP4sbZO0OV
z52XDOiNuK3jJM+ZKUsXdAh+fQ2vYyB2eH6liBgwXHPqqaGdF0FwoX6GKUiEekJg79msnAg4I1bq
1kwOroem4LkEHaWNOL9PZz09X7tq+ibPNdy6QGKsfTENfVF164kBVQbrSwT/bmLLzFpGVjE4ZMgO
PwGXVR6nqth7Tm89wgLpn0RNEdNGyEuxf0nXfib49CJlpnYGzJAJ28WJzV7mCpBxlNsuyb4G90t1
AjoapLrt+cn0EHPlvZNDm10nNaW1LZlR2LNQCBQnUAoQtcAdBaV+dJpTMqY1IVAIwRaxyjO4tmUa
WA0GAy5zpa69yXmoRguKKfgqTQ3kFDoAGWXd8u4UqmG9C2PT8kiUC0o4kGjlB28es74lM5j1cNR6
ysvT1sLjXAbg0Dz3+h3316VoQFVLnDtnknXMuXo1VJg1M60SbmCLZ6LjK3PuCNdFC1RLqnsgkFCZ
97sB0RJNNuVzPgYflj5ifNxt9tDlDwqXtWT8tgnkuFdPlAoW8P48jt8H+pmrbTXq8ueVytntpVHj
yVcXGC0MXpDemL/SyWYr5+HeGmaeebX1FOLCdO+0kIE1Mgzw1246d4PnFQBFQGFUDaJyqpEi2/De
l0u2OwQRsX7FSxUh0+mM+gLD9dLn14JGNrwvxiu6s6aFzBzMwdpwzmhKudutIUl3b8Vpc8Z3CwPm
g63ZLjP6v0wFQ+sYrIboJzPVg4LBSIZzHoA1zYn1QL44l85JFHPvSy4DB+ePZtWzxydGuUdVK11a
HuK5i8OL2zhIOX29YiktJ8PlBoZAF0RfJiiRAcsu1+JjWowxid0xBU8l8n277JzyVVahlEIvKj6u
WVC1aul7nQOuceEB4FxvpvtdDYT8FwE5tlfpFdDygNK8ZPiVq54Dg51rtOoQ+ZmGkoqX3hYbvbQB
he6ftUsYElQDNZwMNs70buyEDtZJSqPmHygNJ78tHrXpGAgDlX3T0gwvs/hsHrWEdlSKhc3Ilf7V
KDGlEfSwThznTXchpfGdS0gDCxqFLMZkn5CQ5F9QGMbPfYwWzqv2G+1daTs8oscNkJQWvLR0oVbS
9+a1riREegLVF5W4QqrRrXkhPpbc65yn8xlqXS5CtZ/2UZdXcCDprNhVpScPythoROQlg4mes47e
iuqjRRDAzsww0AyHLffsL/lgS2hk4GG5R2T/Sg92wBdFxCIfbX/ZDNaY1plG2YeA8jagupwlFWTm
q/LNngl3HG94QJwilUJXtuKl54Wiln6mmYN/x2Rf+UkCoDR0IOvbDiqYsvpUspzHd5gmiPTy02Zi
EH2cwitJTHkieo7MrS9hGNyPgJmFRh3bVAoAgxcf8d2Rc4cIPbt48lELNa4KBu/etLAhvVJtdvAZ
f1JkSOSKtJ7kqx5LkX1ah0pkntw3IrlDLhWFAFfZapl5t53KVP1toYdHMZvTyc+3VsgDl6PBKeCn
9JJ+OPnDL7YRv5b+YUbZXOIhkJGo+h/8UeSmlMxqlsw96xVLLEpncT4sabQM13kpl6S1azyFdhZS
JeyzLNxdsHtKINRfXUQMvsKyIL18HIjxRUeYZrrrLGA7aBW1mgB2Ni3TrJKbsUyZeXaJH4PvhtnP
nJ60FAxjyDIXbgadXNOGzeCUB1eZcfltxVH291Wa2AxyZSNo+wGJArLMKCcJ48j+qbeR/hkowZJZ
VFSgSBjtHMNh7RsXN2enetSnMM0o/FKIQSZcghdjYk6PX1WiCvwXnTuK7odpmiSY/YdEP27e+0Z0
UpEaztSjWBkeDZLSRY9cqkelggtSgdULukpPshpzO/sFe9qry8wj4on1ZccvVYDDa8+ZSBIIZCzS
A/+nP+kWcbbCg9piPG34g/38pJQVNraccMtMVc6UMOaXg4qi7hSgMh8H35bmNyvP+4FpCQxbGqc0
BeZHhTF/lBGGNDulUMnF8fXLpH+uDdnt0OPyY/w6bO+mt97fawuDbmPqhCQJYtG4hLmYsuyh2fIp
xftolQxJ/5H2WCDfXhJfz1hiXRWoIvftUQSL2Z0902r0J6WUHQxoC45mP5NTaCGvYjrxd+yUnTc8
Q9UTsB5YsATgiAUjGX3fg/WED1PQSNK0PjKscl0MiliL6Mx/9FctpsA3y8dgPKHp8PKOu9bNPWk2
rnQYiSwPAnrWLaQT8+saPWyKfQ4RlTb1ZlK3Df39bK3WQZtiXb3FcgyZ1dEIGt9HHVwYwDVkZSNf
gR+uBl4bLFk21LTCtmTTmhqxZ99QTVBUKIl/y9nwSLVOsUczezU8SLjI3Z3gswDsa95opjKZiwc/
rLZdY6p/QHqlc9S9vj+7NqPbd8jR2q/g+e+aZ1XoiFcn+V5+JIwFlQisvwF72d3JUTa4iidHqGts
bLRz/OApSOTb2rlOEoyUFSkU9QEWotjAUYST15uM70wGwxVGliD13A2FNazt3FpZNJVeQVJAokCx
SB+5BSoE8E5DL45lrSOb1GsVRJII0c2U1rDI847pAz5yFHkO1hHh8TU/mnSavikrnyu/4QjkgUyB
Cnz6Ri1oxzJp2JO/ikAMIe7AZGFCd8MIfitzs/2YICoMhlmfexQFc8HPOUJEAY5RUZ2OjEgEP5gj
vyQEMh7mVuq95hWZw7IabfsdUbe677cadqU9KKBa97iHw2e1IbAm2dMIYZulUVL/I3faJNjJey4r
d4SB78+pfblGVsQoxUZ+k4Ah4xH7V+7Ok3sqRZeKzKG/NaEbffUe0zhks4dh2j3y+cpqYBT7HNbS
u2N2fg0noCIvqMbaj15CmFA0QMoz1n7w66HJBCWok55pchWRBlf8gbLHFK98fIdzFLC98cckTdHx
ocs2OM/RzhFH3i5QVNGRj8bDTGTpfI5GnClofb9BOeFHZM/Xs8+Q/NSsQp+peKdOlOWq5YSaOAf3
kzpJtvpd6Kq6qu/Fdt4OiLg064Vkj5P2yT/OAZ8ZzsGtuDdSMW7OgNmAHckARCEfzgqIKxXCbt1F
BmUvkEQ+pNCoUN53ecOWHRphi364EuB1xmq0HQ4yHBnLjqzwE8tUQd5MaVS6ayvI4RQHwLOKOGfR
6H1w7EbqDPYaOOur4x6qKQOpeW5vEIH0iQJBHVaeNynxLw2ZMGcQky/55cSQczsmn44qD46hX2gI
MZK3eLbj628cHS/I3pSigBa1iAhnwuqUVYEwY2AD7lVbF/wOwjcJzzjz3WZU8LuqdS6X/WXID4fo
rXJaFL5EUcfRUnPT2HTIbKKJ0Xls1g6fnTwapxn1m9DjcV+cTW70b5EX07bCY434qhibYoq2Z+jJ
SaxYqLXB/7ewwJEgQUm1sFCA7xM5Z9CxA8Bruu7bJloLwi7CG09M35yGdaYfkBYwpYni9jpF/7Zi
4yjFhChsTv40DNnw7/WfmRl6XtuMgZrKnpZjR80R/EJIxePmcBZ4dlz0SeRnrKUdw5i/YmlUuZaj
mgGkhuGnO4waZXekccfoAkT2PCjrq4neV7eQ3Ux50AJtziU2DjVjzXTnYP0TUQlwNYLSenbIvAPB
3TCoNCijTXcIjyfqoRL9x5Xd5rNcERGtmnkHybLHWCW2ELUNNbgX6TEgdVnmfPWg7GpW1sN7ErX9
GsaDsdwe9pxwto9oKGd5A6B0L5pvszFmhGLDdwOHMfXPV228dgoLpRSAtv+zOoIpRoYjRPx5A4vD
+b/MgGaExMaglwGf/6Frs9Yeu6nRfHvP/rkMAv8Eopht5c7qwthTyiuRMQjlmE/DvVcWUw8s/7Vz
i8ogSJs3dh/LYf52ula0xPPSEA3MbQ4T+bzlv3nIN46lzHrC3WBI+7hqoxRnnPeHyOMOMEOJ4tk+
M+Sqd6Xi/rEkOyts1UTqtW2aV6fvCE9alTWyMJB94w15/t3iYd0XVFeHYzF4BpUHpcQ8UAEHhgz7
wV7fyqD2gc++e+LdFdY9WCto70okFSf4tvaVKY9+KSzbWcFzLJNRjQgygyvghCn7E7yWZJekTG8x
+1zpfTtXUylPBt1HbOxX4S/JW/Ar2q508oTXDLYis3tINgvq5UN3uTnv0Et6+O58PAQ8lFKLocUE
Xh0iWEBBc2GBma42dB9ENvtPKmGkAVTtS/nbbscfyGb0TdfBntQTWQy98WfsK9JWCHaKT+Q3MihZ
tyiUCM4MD36MgcJKbHCQs2QUNPBIJSwlfZHfDAjhUQIhz6zE7wwDCwBrjO19Z+tn81HhuSn93Frt
vPnXFrtdeHwrJk9mtPd1RCYww3lTVWnxflC9hSym/+4JBru+R88sRZiDR9HuwMxan9V17zfaTqgq
VeGe/+EIOJNu6tpKIy8P1KVZ859E8hHo8hfoC7c53tH4d/UPyjpCfu2uT1v/s4Jvs5MXFJs6o0wQ
bX0GN5C7/sAd1aWy4fA1NL4U2fjNcrDr1fRJbcVyyVsiEW9i7lqcJnEzA7Uy3hl+H2MUY38bntgu
zRVi3avLaa924TZ9pwTUF83MCwG5RsRnQLcFdJaH69i2EHB4nLnwvLzktcR7wYUow3sXsASaqauk
gp6kfh6BapXWpVHOlFl3TYsmGB0iU9TIeHjcwpc7VO0typxFzZBEaWD00YFzdY1dh3SapqDcrqwA
nMnG31XCSob3elsWeA6cbXzjaQTkwO7Md7IWT0lzyAloelmPEP0eXg1FI8+HviPgYo2jE3dadT/Y
GmqNyofD8Z2lNpLnlsZsN9mK3WPc0Z7dpHwP2WPgRgwSHVDQT92ENZ3zynsa7voCCRDPKWd20zX9
AWGpQZbmfsXw9YV/v8dcgMltpCPgJzfOPwJt5m564nh0juXmJ9eEruGoylyKQ9eAPC418tdu6Rj5
RegRWKBbi5fZxgh26qL5TRBxFUhtnioOwjCW1ysvPR2Gfryge/A31Ojb7b7HmSkphsznM0wrbgqb
i15zX+iHj/dQNTKTQuyFVxCB7rBajj9szn/TER4O1Cmuc1xc+9LJnWaucgdRt9UWQdmxSFKKjArv
1CYQ/V842IpCNvMWPtZuTCsk46qW8fZVRz72EpF3LpCtvm4r4EuuZdDxv9ZsTxvP0axgGImL7jQE
NC1aZ0UBSLOD9eh1yFst0KYey5LbzaEHhA5gjXqiz+1t4xEe3N3+zOeMfthq2Qeb7tsDpb7fBF1O
bvMftcpLVn85oovoP8IhUw9980axmP7bM470iHv6EmJVVDUv9W7P2LzpGYi751ZFUS/uBClT2UTu
BmWm+/wfKIt4aka5R0oSVN5+mXwNDAiQ3ih4kbc2v90fnn3+SMIRFiqpibpkVABQ7dl8ThbkEi1f
CoPXOvkm2Z9M4ZFvtMq/2qCMw4GhoFM+tA0TJpw1eDK59FI11hUyPqnV5BYPiUhkjbgsoL/Zpboe
O+Rgfm1OXppm16ZvEV3iMVwwOTxbF+7eSHZFgonVq9zzLWb0jSbTH2nGlBjZ5kKjVgo359obeCk1
itwdZe0NcneMqKI9aPU5m4vYrduQU9lOnZ8iZRX+cXvPg33iRvbLdxgsdSMnZllq2x/77m2up4x1
sIkKPPGhSfvxbOGNkK094kUtrz0kX9aaWk4c97gTcPYAzVYzUmd94y2PM+I6n9o4q9NXHYR/I4Xv
YfEjPCffCnd3Xef2TfkBSRDQt/htfUHJQF7tjvyVBe9BCoEKlfRKPJFNXjeY23ZKOj0g7+mdgkOu
BSfh0PtyaQ6qkNtvBjPQHgW6Du6DbY4ABhwv6UfqQ+v6wveviJ5ov2xojfNeyPOdEYk+d8ItWgJl
RcDpw9moME+7WL7gn4zTU6dxCPYiR/ppdc5DYs0xsugFFzoTCLmCZXCftbH5nONx3ccaWuIlE9lD
l4igZZ2giKt2562ywBm+4jg8RWTcFsW3xt6hLoMcDV3ejGH8SQcq1wSSjFRhpDVJ747XFXrr17Ot
ndHYikiUg1O0vuKrgFvAnXzfyQpLLbVHRtMlHlsOemG/AgL5fKyujR34yh3Y3ETwID/w1Ou4mdOL
GEiEVEEXDOg2kEGO82xoDP+K4p6DjWKHALWCmhsQNA3iGYBAyRxERzimx0TpNDfq5rG/UkgMFMBD
oR5zBiTpfkv+vJSZ2xwxK3V41EmiodlspLO79GafRAUb+rnWyw/MLnUX2hNCDn8M9hBkfR3yZbfk
NQdNjueowaSQasOYL1s1M9SVg3M5T8iFhwzoHDlSeDOZb1uhoeQMOghNMQ/lvdgM95e1NBa0m8aQ
yaYqdjdu3q1XKIytnS+Ce6QBJ3ZQQo/BZnLmCZXU/mLWfeucEc5ZBzHYOCTrq+dx7sfDKla6iKDe
eM9559f5FOEQgiutb9mwigtpkZU4A3OXfguIfTjv8OkhkzYulyHd2CB4IuPK3pL5Bf51TTkGFpX1
bCy0zQhkwreOPabuJ//0Sqa8AeG/iivditO+0UGxfdRD7fqvPOw1K08p9CRPMcRq5R32x00JLPn3
ZidUl0FSn3OguO5+pKaoLuJrQqGa/meO3MZIhrwLngWFN6ign7DCqkAkVVhMLDrKGXagUoOdwSab
LXGOECjNr44Ro4ANWB8VBRq/T1YkWuj9Lq0yEg/KWoWTaING3LwZOcqj2ZumvDJAZlNgmTUu5ofC
u1ujsHVsILGkLF68tn7pCs4/ftmGlY3doDPHIBfcZMF6o6AG5ktVk9N4Vz3FUV7gxR6aGmSrFBbg
UdHuU9HDrQfx+XxSoG4J0U95P+p2PgXcgXiwHubML5KCFtMge6OcM2l+GSd0OPdwQGcWG0ku63Mn
vXJD0WlAKH5/XknHrBkY6UAMFw8lh6sqCadWcrQC+VPxyB3skWnSyPRE1CY6kQ3NuI4oR11OrqpK
WG/7It7cHueFkKGyUR5KrBeDDB5snHVjnTXPJ9VTzmayUHjjB/XR4Z2tk5gGy5moIQJp9jZUCVxl
FM1Wz9tYEO/InYVW/VFOZDQUljb5KJC42c2PTlHv8iRDc4AVZm46ZhWJV6YjtMDNFPWJaACezSQi
a9gqldJ+lWooSJRdvd/0fdKOecxfk1ZFeSxQumSOWYHyoEqiVDTxyCX7PJhynXkGP/JrHaCS5xQD
a1dcG7REi3Us/LrJQzz6SY60wVZAQtNLVhRAfb2Hu9KQpm2AQwE199Ktg+1uU09Tw49Ve3xlUaS4
xJ3aJpci4lm2qAbgAkSb8YrZ31VyC26nPCQsvjSAdlxgpDSWgdU9kiEzVWFkEhZpPa+OwSjFlV0n
e/XqihlZqXO0VxZMCek2FFtU/askvGXUL9YnFzfti1bAwFv7vSqEt95Qoh57VL45Dy+R12HlKhrL
3/HR3Dr/QE55t64cfODxA9vU/pxZiGDaLxdKi/l4JP50RKzmGWpcBK6sWPbnHxVWUolj17X6YCn9
NeK/rD4w5i98kz/K89qsdJ2OjJ+43JcmhTcxs5rmPdfCNFrs6cDEJnj7ONP40BGAWWv53TiTrOpE
hEnyin1ON2EDScPTB8rzs9tD+EHo67+CxZSFn5/tcJbue6LAq/SE4fB8t+1TxHjt1BEDiQbY5pQm
cTzIHIBmDxwx/w48ZNhjxbVyvQbKsstxO/L3PZVP3o+/X1V6r1PmwfFDGpccqTpOCVqEell1onkY
B+25lih0Hs5DkAkBuvx6r+pnG85rv3HxRFUhuPPm/jgbcT53eipYUd8ud1OR8D8vpV1MgJKXkPWM
KrMCiMQd/6ZdbAymJZXOclVrrqt9lTT3xNKvDSwDSYgQjVpF1X51wGH++4dK4x7ec25C9oK+l0BV
rZ+xTuCUttsJ8Y9A2s9/z/M44I8TCHUiVXdl1hPu++Q3YfDW9ddfPH2J6ogBYC+LzDrPffg4lghY
u6GePkdh+x5EY6DsODPxOkKP/dB0nX2qfM7U2r2g0Y598CQ8qMHinT6lQWznAeBAOhWzLpaWCLB4
zSjPLrKfZZ4h0NrUN548AXBC2n/NaDYRUCsCgs+oB7k+Qgj4S1DXtMuK7qhOA7phQgZTFzqFeloe
xCQpmTP8XGCwr5tyZAbfMhLi5IxJSRaUG+QTNASOyhIr96r1xtrsrXrnlKas1fXb6fJYFqJAS/7S
AgsrLBZxKSvPUm4pdmOBH1NPiFtT2AX3Adk4OlCl0UaYVJa2va80XF9D+5FttOE6jrWfrM7OU87e
bD6gulk+Xvuj1ikn4fppKRql+ZgFbVtjPKshMGwqbA/Ugigb4reM60vF4IShfn3ZFQQOGJLTyRc0
W4L0RZdALTyKzdZaviURWSOM75BMvRWh9WDlrNlYbbJQnDs34YTGTEVMoyor9MK7gJovlkxijIIJ
VHumk3cyVQQrEoUWblx+K+pvwP+wWvR8kw07KPCxCbT1978iC35CnO+fpA3PWLKvQw/9b0bCLn3e
t6eUkT+hf1O5j8BSfVxAEa9xzgrh1lkFaeyHc+FJOM+D1H3uwZERStwjiXA64JVE3khjtAJbjrLq
s59W/DmlrSerNgsqrVT7nT8ke3qQfgLIG/+fLqEXRWaSCC2AVH9VtgytNQyHapLhio0lOs3ogPb6
VU1BiJ9LmX9ooK19yjaZ+PfPDtTGJp7O/CtHdZsD1JWkdYCEXN9jmJ6cPB8DGIVyj/iXyJZ4OBiV
bb+UZe5WloVJm7U3f4aEWZ3/YMMeet1451lMu8jrvbJ2KD3sRBwohfBToBvf9arcvC6xh08JR98/
bOY7YGyCvCIpF3+K2Zi4USn2WO7q1U5wgOPhq7/9mNCdW8NZuIsTFriEXR9fRVzW4StB0i2HX1ES
QdZm9A/6ieAfjLKPUc8ZT4K791bvVFAalIBwuu0I/Csg5JnJhkEECIxNf59o/0A8HPf03srCQxnF
xFtW88s1h2HOL6s16vv3QONP9DbIulpSn81QDicfbA9E/sdXShDL/Xh7+3SdwdKbiaMgm+gEnU0c
b8uQ3Nq3ztKmW41CQWO4sHwh2fOYu5zNYIFR/LDGKxNNU8S0Bn8YG+epYnEiWs/dDX3SVPlVNPMm
BQ3+KAYA4wsY8yThRP0sUO4742GIYJbr2YYaFaA8/RR3sVq/1v5r1lnjEXSZUknDGb9wkv7xa2Iv
g5eQ4R+nSotXDnN1i6OKj3ZDGwkrtk1JCJGVrOPIHM4KzTDKVcID0vbbbM+oYfqh8l2y3Pje7Ar5
XUDIaRg4ZhggCkVbW4t8w6Rn2Xc5pulAFNr+W40BKb2ihmX7L20c6lD614BohEVMFxaZUo2l5CBd
d7RxLr/WDeKh3UgfaUw8letraLupMEMDIEirOlR/fHflwCeO3mqD2vigmAF20IvaJFY+6X5pGjHO
n0Z2SGeGvv7fGjqWHuHLc8AmgSzQZErWzeTZI2BqwUiWGVCRT3PuO+B7q+9g9/gUswCSIIODeyus
tmyeWNWeXISQLrW8Rx9E7KfOO0YSJWAtfDyd1nMhl/s72u+nnvjq+mjdzm2ULF0KBAlhQECDiKX3
DvBSgq6L/non7QTn72/4cWeEQ+i/+nvaCr1HRUhVoErNwWW0tPLmAib+x1sLkOpoNHVIZWbYx+ti
zePtG0rugqpeCWtDT7Je5f39NeQK66nvld9IN596+qr3AVA4NJSO099R+IoHREvw69Q+IUTtnESw
jZ34SUOT5+OmlNaMr9nOXFBFSai7qdtPtvhk1EolTF+qWEkCZmWR1CL+KwQZ3c0zlaPCpWyR3Q75
qTNIrY8Hlp9PfGTIHlFUqIl6u3rueKOrY5Ofq5IVDukPdtZNX3NO53MN0qwZcQ3dobrq3NuYDiDV
VZDQUDWZsomdgczVemceFs9xxnlMMsF4o//ZiBW6kgb9Q/O3kxqjxuHylsoxlLZU3WNYR8Pfb+nT
ALXvKbFZg75GrOFVX++lQUE8wKNBP2aYpbxPRb6sDm4QZfNCTKoUVSp1rDV6SpdadCacn+F4NXp/
S6FMPhWoS/Kvd5ff6abxVuC1Y7uxFJFD89s9igL9hNuix6vRELmbv2noLSnSJR97l0KzLISuiaah
oVqJdmVDV6kZN75h1Otov1L7sZYwXsJLuYFmphCQBBeqYcPsohGLgBFyQ/gc6gazzqyksisDch/E
eOzXARdX5njqLQK4XPkmmp104gv+O05DBTXlGqjSq6JlvtONMCwqVnY/mtGekl0aM/Hx9HVl5fCs
DBqeeq8VL8JG9lv+BQg4IoeEzkHpNeG7e5DP1Cq7lIAniYbNR/KB5VGDgcV7F+5v7B+3WWa4Qskn
/1iJaLrxvcTEZaq4yef9VroCsppT0ExXc7oUUrvZbbNPmp55RGl8etnsZItsA6Xs3ZKEOqY8n4Cv
fk6/DmpHL6+jcoMeexG2t4VK8A7nPCKBZb18iiCa7/ISzReep9djMx0hBekT4KZ9TJ9s+7tkk6/b
mtchR+Fl89YRxkVG0cluHtrZze95kEsoCcQuxpnU5k6eqjz58fNQa5cQ6XOu3ixfft5gMbxKqmlI
swjV9hi3RXwqgcoFqk2SlZuvV4kUwIWEF1x8yni3VuZPL40vp8h+ZWFTYGp6R0caHx8NQT9TsnRF
OBXdjfWv60NcROZL5+4qMX0VuUZFfygizZy7jyxQSOmc7m+LlLzAUrhbBTujZ+Klk2sj3+01FeYB
ZNsvv1gYe+8flV2dwsg+LX50x6FDTseh/dzkANWRIM6OMkYQLQHsBHgpAxv8d0qhE76Rl7TenSH/
S0ZEBMssWhCLpzN6XkMP67JCPalCqnZbJUvTkApGUp4cvGkA8YswqaEXMferHCKJs3fiADTKJv9g
ii5ypW3ff3wfFs7bKdoRuFjMDy5F9o4TofZafppsE8iDlXcEzaqmHqZrCsp6WGxVBWnU4W09F2sT
z+GN4orxiAuZWFMMU7RjmZwQ38as6KE1olRp+3wFx42yDuBb/fqOEZa8QQm3tZ2AX5U+GKLTXW5X
5fkY0Gmh5z0heOP4RhwEpDffioTbfLidnlGFJPfmbwvn1dZSbcmc6zM201Mx8Mv6kh6inLeaOOfl
3A9sbV04Ua+xhla+wV7OxcATuUcl+ewFXdtX+Au0c/iX+JUQiMo0wKXyZQXLXB8pHFRkOohO9578
g1KYB3S5LrMUd5ZZ+7Eez9pw8fMhadRoQCb+GAFji0K41gss47lASg2j6BWDl8XKTXhsT0FI13Pc
L9RR3XTkTumGKy4nPM1WrqWW0OZdxz56ZJCP1kh73524H0DHkzVk/Y9AygAJ1RgNIdNbQzDhH9Qs
kyuaMpQmzqWzJ07j1fnTxU1WCjqKDs3uzNxgw02UFuNAW8B9ZQqvj6G8HcWzL+c0YovM76+F9LFR
6o0fdokDp9pVu5pcYejdJIyTTJlyUgY37KuyrmQTLg+I6bDKrQHN9A+9RPVMJo23fvZfad7i06x9
PxabevwASBTWcGiRZY7qYucQrhkEnccQ0+LkEldnOudaoez8sf3sDbcz70Zd6yX3c1mWOne9BQvs
LiHP6SHzQxt/TRkDQpiC+568xIEFB9xEa3Jwy/eSttiwinP+AYJzUrAnk6p2hLSjzJPLHD1ejCzD
9Y+Q22pi4t0xIawR7cJGGNvv0gkbmaUO3Kon+bBRM6r6JWlM9qYt4FDQ0JTuW+BCESfV2DAq8tUh
UZsCsPanwSoftGyS3i3zmvBb5bVYFP9j4z1E2Eb3V0CmomQayBzyhc4W6uu+09flmInJblYsF5KA
Jap5/onLNFOQ0OkfQu/2GipR9PDQhBpOr99DV0WRSJg9A9tWHvd0HO539wu2do2wyfGZraswUvSq
1jzv/fCnIp8xINVHqwZ/2D6SKLlwV9VCsPhhNPetpWnZhrYBRw/FblQFd15bxkQwSOFkDTpgAMcc
IjtHPDIL/t2ndvCXLW7+/TWtKBDfm4qHUjFkm27iZTsCQ+YASfRZXnoSBHF1nf+iVC9PtLTDbYsz
EB4kJ3X/x+lITr5WWXuM1koOtJBRX2OUGPzM+Qg4mKxrc8Y6UEUM1Mca8PVLKIiIVIgYKZ6ndM/X
ZlKV0rQ3F/N2cUEPiaM0TsfhA1PKjMmVduV6uS/tdxRbR7eTg8KVWlvFH0heRg0iC4Uhesi5BCbW
DAj54BWtmfKu7ViepqAwofa4kNdnDFxsdR4lw6klvyRBnnsgM02Bqt6073bDREBAdk4YIkIrlLK8
gfr+SRNXx1K3aI6sU5NgFGCUZOD9QRA8A4xJyzE5cpsd3QZp0HZtGR2RDreOhhUfskp49R96z1TT
cl9/2wnWlx/bjKWSXnnLgRoOnW8iss9cY8hpZXeJY+vuhVszyF2gGfdW8cBca58KD4HiFKZRx1mO
sqQplultOmaN+6hiprzrvZZBheO2mpnKET9jYSDYytWSZB4slPJmVmL5oyaVFn5zCBJTG5CVXOXN
sXQrq493O21BFgFKdfmDZocPV1ICGM67OK8ovSsTpdBRr5y6cGSrIjJ5Joxj+9XPAjlsTOTfNr9l
utuWsNu+rT7aH1UIDsT7vuexPVbxTXQuklhzvrYIOa9Dqc9Ai2HfitBsnBT7fZJUBtd/eY3LpnRk
uYHHvI5+zGn/VqxZmyYzDe8IFkjuHp8QgzeANVzaH0zUDQc0YnTI9jqzrUXgI0hTWC30Miuok2D0
9Y+rmn77lPLfLelbKhxQwb10ZSOqfFzTGT/j3eMqyTtGErm3rYCJTqljrgfBe2XoH9RxZCIu9oEE
+MVU764+lYu0F+NCJhq1c4UhizwKlGieJgs7hHoaXG4y+Crkhk74DDjA5vxvPFWiQUK7oQl3QQLj
qZMFO9as+ODKFPEMtuGQyEcq4t698fKW43L1AshHCKIScj1rm+Lsoteo6L+eh/OVyTcmttc2tFvv
0iwwF7lx15DqM+0O5cLxEMufSXuGM+DH5KYviMIF8Q6kOYkaKVcsKwtzCEM93r65zSi587BTey59
ot9BeG4Gza7IVTlP10v997aqsP4dECbFpgecoYzGLXGDj/8UadUNcsqwbh0H+zcdhLSoOegR5brX
8Z0NeX+4YNobQX/Qjl0xj2cV8G0WQI2hrRZdaUi7sCp8btkKszZibEPVI433Mf5JhnWmm2djW3ec
yGu2/odcKwm+9CVxhc/3mwdhgv8T34FrcTGOWqC4wviHvmBZGEPBrtg959y09aAa09lINi1t0TZ1
LfUU5iGeUQBI8Gps3OlpfiO+MyZbV7sMjWo5hjWWy13fo6sCD1SqEhuKu2vYS8aHti7SeV21wrUH
DbIsd9fNyWEVqEHS7FmZ4b+OQqvI33ZFI1t6m7OcO3rjHVsLQrQOJLWGjDVMK+ZDeWg0O4Ucuwhh
bS0R/tLJYEkv1flifcweT3lQTu93zUr7806tOpOVcPxu3l4b243zUlhgHgn4Llnndv5stL3Xl5Or
D3agXjnwyUPfLOaMyd6ZONQSS/Px8tpnmQj4fqTIHO2a1FNtdN51RXhXC0dRy1+PgTyD+QFc9Q7U
WBabx+9Wfl8Vij+HQWaVWp3AiYbqI21l4pIU4u/hWFETMytzCPYezDv7xNYQIucg7bhkndwZCyWB
q+znZcJCoJ0/9/g+94LgTmWC4ywIHFHpujQ5xj7tuQmFmJ8QPvSn6vKz5PbxWRKvz0TDKtoPGH93
O997pX3LRTWM/6iBuGW4SA8T14JGeNxkuAu9BWmKKm2m7KWW1mlN00BIecHvgTFMRo5uViC53aQa
gNsGxjOl7ERwucEQkpAZdA5MUq7mlGikgdUQRi1TZ2goweS+k9Lru6jf3k3AYBz1Stgr7JvJKKut
RrzlLkckgZBPsUS7hxe7aJ3w7Kv9C/8MqNHr45WwpESIZEh2lr6Yk3j7wzem58qHmpNwklKmuIaQ
boOS9q1HkGjvEb9I0GQ5YiO+X610Zs2BbegiSmnNZqb9K6CCSOY8I7/eh2E5cJLBDOcwMsgowHsk
RefcEviZG2t4ECGzKAa8Fho9ptsPXv97bfZnIPG0x3gNooPqDZAd0Y6szzift3C3Q6MszNIKGYLZ
GwcwCuOTQBWTbhDETQ/3fbjLHLRsKlIs5ZRBiuzLrpm4FSLJnX5OzPIEY3tu2B1FNbcG4BddWN6D
TYt7YPUbxBLErxAILjSiwnQhxv3YM0MuQllyz0hfahj7Jxahm/vCmYrO5XmzRO2X+dhoJhhbdzkB
xVKAlWkyITBbnpd5aNLaLWvGlFOlwMt5bMsuKa008JuCRGewQqLERZWqZvMYoxsVVuYcJcAODKGJ
Qn2s2gOPot8cSZNZf7jL9RU4zFaAXwD68gP9VinjftkVwgE9FvDM/ft9H6cOyKdNsWgNh8/5sDjp
qiQq38ykvU0SBckVXhmMUL3s9mycgbq3C5lGsLsAbvjq00ITNojnvWbQPDvgordwTRDgI7em4eoH
q9X5t8GEOwxU7n2hp1oXywLRnmHY5+h6DPXfZN3NB5H6AmiXt59MK0VfnEWVHQEDmVc5S4Fn+9N+
7uB35zQKbqDjChALV8TkHw3yaLcoLHN2HWhkQMGHGz3Gsdl114mX2Bq46zzE0jixDbLZ73foXh2Y
EIFGnchN7XDpWcF/IQH5vrv7xGnW+Z8iK3UYLBywrL0zKVF515RccaF6wxVy8qJbxTjbvzBfmRy3
l2IG6XOTY0DjXiaS6+6+27Fr/IwLV28iNWG63VmuwVHdGOyfz9lxS5I3hZlTJ3cvLEyIzelqt9us
ASio5AFAJBUMHqd1kww9et3X2hNxgltHg7m3NZxOItBn8YiLg7eUVzzOmG7lRjj3hTCqMvKCVRMi
1i/tL7dipBrtY5F1FRoci0VAwf8J0JbLwHKhi18WrxcVsEPxyTUpa2nEGiHgcSscFwZz3qFm8nXm
IrcIH1VO/quEygw2rqh8/yqIJ4F12fTyvCrW73+R8Kqp0dgXg3WbWr8EOa+J5+sce3WvFrhjbufg
o0bsV1X5VzjwmvbhXGOtSSfXlYnwnssLdYIqYGI7zZcxc54Wl3emeWI/EcMTeTzGfYQFRfSqfMMG
J59XFOmRJBv2iGpsRO7eVZCedE+iTWEyZTkRgaDko/zFoBFU0qfL2e8IozcZ2mcbD/EjinzJ/b5+
6ZbAnxKPi/ynZE/1GTEq6befcgxqn5aayRzCZuu1Q2V1Kb0vbo1AqyymStzVQRWq693OHFQcQSUr
60HeGrU31IsRLjtpfeeERiWfUeWUbgtnNo+LEVmFF1DTpku2xi3+Otmt29Hj80c+ImN8KeRca5Oj
PVO43ZAXzBkragTPKwpYhYaXaQDcnATSGHuaHe18PVX1Df+ZpCzRrl1NtmYB+txY7/39g7GuzSFN
NG6AhvEy1K4fdd1cTMD79iA9R77D2Vod3R7/ZJTxJeTIRmqAINme+8Iu6mm8b+Zq3YFzverevVd2
USV+ckY7ec9Bmd7ZF1P71AvzovZRqxqVlOhrmrmkdtAHpL0dB9y8SHmiPrq82KfQ1jskTk17A3MI
SChyrKtyMzkbYJ+rVMulPZK4sA+w5XwEUjmWIhyfuviEmvk0B9llCUh/yt8GEo4/+8eLPE6XKQ9W
B6EljidDb998JpaVPsk68r4CJ0Iqr1PPZ4z4Fy3wLFnBb/pYb5Vkrt2LU81qR2y/RfWUDYRGsHJQ
otcP/Wj3SJctrn2TkUrskxQl7rpkoIBnQZw1ZoUF7t20NlBJzA21vOVfuxoAi5Hu8LKPXJIEtoBv
3jaNPGvTeueyab7bHOOoPx2oqOaJQb9Y+dCm10pef6Z4zNoYdWYNvc4BBEeEIqEzKuMnF4D4zjZc
GOgtic17qtItjaeyUF2+AfIMQWQreZHkml3uZNsYdf5YAV1FU9RaUEKBR5gDtTNhMpqb3xg7uJQX
bVN6u9pF65+kkZ8X7NJfhJaQo9hijhUB6VZvl7f0jhCIni/MXdkLFGe/28vWu36eNw4uAQ8AlGhf
xY8xKnHM3qiPPUxMi+tNvbwj5bL4NXRmCzR9Jv/HocloEnNhbRCrgRSGlFdfRCsokWn8gbvrUdC5
0zM0qllh8qokmSo3XW6R07SZw0tMf5TVKbhLEPwwNcib9KgoavoqDUStlScxB0c5Jxh6S8Vn1lfT
fGafyO0FKp2GkKwM+QVd+mboHZhmhOaszte/kAhDc0u8MIMJgf4hJRcw9ftVJOLQnwP6V3Tt0ObT
ZB06CklM0K2DhNGtDlGCz3D8bH60tmtQXY7KiK9yktCa6waPu7nkUC+/F5NVRtNfw63ClFSJClaB
HLovWX3N/CzcBZlEiZQPB6LumlbRbwhAYM0f/XVgasDafekgOKbu/SzSirBDyp6k1RAnuhkfaqne
Zm8h/ALF3DfK9eSpa9Q+AqJ04qodaIi5bSAPoOQpfHtuKriVvhUq9Nv4yqVIn6e0QZoLgitkU6Dm
FLJKP332XIlJQZalg5dDcjA+GKiH8aZsyiM3zLtIfPbbNk5OdKaxBoDQRdP+subxiE+bQ/uM+pqA
H7o9SDisn0TVfkSK47kFUVadjW4oYZjrQvID2AeSZNpLojBqW7odAwtH4soBgfCMD0kl/TbEq3rs
VFP6q0d6xMpLVqEe++QbyyeoCtSNzyA7ix5GGv+jCzPlaeLa9IrG69kBui2/s4tsZ8awI+l4uVhF
DJ+MaH3wLPCBcYliqTsdqvM/qnMdkXFZsHQVnPWIc8gYsDAhcKXHR81HPMcLlMwhkum3XIwOk5ge
X2k++5akF783VqDkMtd608Vd8o0czKG/iNfIj2rNm3kqBji/9Uh84I0v6usgG5fMBLRnzFfcUeyx
AYutB491A/7b2+DoY1nRF2aPtCw1X+L0mLfG8u4Ay8lhVTgA0m90LqGxNSFfBJLjNJyLdYhm5qZM
MwVw4aboqmxLsOK9tUtHXqVE2y5/TOKvvWZWYnenE12GfRHQnbxB92YTYDMYX71LBtDFXU2ELQwy
BhRmzHRrylERr7QqBuUrPXE5ENzPwRu6vsBhXND30RdQ3SBVaSH4SUbnmLQweiVFg0Bc+MzCvKfQ
lb5m5gn936R5GeJ0WbLxBt/q6nWfvLy/iQxJhEc4p0ITvabk3Cz8Q0AVTX4wqUADmtSlxdzFuR3p
bw/8JIb4HxuXkRdgbngDQIsW+z1SiRTd37EV0ggQ4m6hR5KJQbedqZJahM2hQJRJkAHFBgo347O8
w81JmC973kNEcM3GkUfz1ZeYCnUKIjVopgXivkf/CXjGXYfGtVcSY4GcnFHGm63OuFX1CkCTJIha
ci4QukrqSqi+lgVCdJtS/W86TCqzS47s8S0cSCYT0uxNrUkLzaX6QUyFDz8WMY+9LfvqGCQMZblp
NkQN4nTOgsl990omwmZMEHPgO4umFy0tbItl2t8qaJYq1GvalASWXY4ozfd9O2wP4KoZDCJsYHn/
gR4N8XPJyyMfYQE8h6VX7fgGZCPMEVo6JHn6fSGB9gmYrw9BQIYZ0PZRiecBO9/UnlC9SlYRA8MI
bhPOWANBtwjWE59SfHgFoMooiyw3NNgo21KeAP8bL4hVdeIdJp4WRODmvB3y611GF2U3mB5pgg39
DAuXaqNkTY5RZihEVqwbt1VjKct/IB3Nann1jcV28X8jjhunbT3pu/5F4QK9EYxB/fxxdQkZDTxO
YqrfvnHZyvfBtePNVj5R5ZDrgjAu1CABFUkLbD5RJNbOAbWv4kCpXBc5TCRgjVO2J3kEoUWyzMIH
LEg3ufeg2v7utyRczehbYr+g8hOTygoqQn2V0Oqx0mRyNzpjMlil/ie4DHZX7WoLHugRpA7LZShQ
/NaQ4CW4RbihkMFlFjU3J7/4fzjLolXP9itCHcVAAv40NWpbk+XjTxFPY2apc7sdDzcCQjffzCWi
NlS2vb5mrxXKe1aHxHATs1IeNlIwO5TcfeXxsdCPyogXOrQN5MZizxll2vVsCubnz8KnbBGs+g7f
lxHsbKhgCdU8D9Bu/WVJJ/YOhJPnjs2Pe9979kfVfa9M8e3efDasLqr0rarFejkQoIGX7AOS4Ax8
vV7bl6ehhq3WucKgaIzIAv6Gitn0we28eIB8bHjlRyB/0xz2vk+aFtk/w4VBCgmwzOEIxudVj1Yj
d12Pzz8K9fhNiTtGL0NE/piB0lmhD/WtUxelPwMqK6jPCTbGxsjRzeGjrr+svRI3SDVCHOdKfBk7
Rz1xdskOUCQdDaCTXK2kQdL1v8yNVEtokEiUgBd7p31lcJL2+yQuth6ONsPRfZLhFCFC9hGHl9Lw
0BKlFVCE/YZFxTyfu7rWmYFwUuhlcW2j+tWv9CjDApwv3HYAcAhWeN4+JFw2tUqIox03qnbJn8FN
ZDBNwcttVzn/4Vtg2B8ETyHjhw48uzkqO3/M1n59uO2uWKW33LyO9ZfBfvbZ89IuQjqnKsxSCnOf
VYaXDA27kB5I9n/OLONWxpHqyhfiVgxpmZIkdQZf9Q0KXRgjcJ4bt9J403Th28dfdC6yLeVaBJ6z
JeNGCfEtsoXBDdZwJmQ03dvFM1unmGEr4S6UWpTpl0dteXsUzA5EvckcYy9qnceuaVXPvw7sSedQ
K3LCDP0zZW+/y4iLs0M/Rsc8a8oMFLlv7pltEbfkBxEjazydxbcJIe1y8lKY3UIkRj44yw7YTExr
VbToQav7QOvvqEgoU/ExB8AkbfGfIEJCeYkGMzBXuoip3YTyF3FvYbF+wq2yLBFp/gn4emXgqfr0
/vXu4wlj0xhOTVdCU0FwwVCT4Tf0tuJKykBhUM3Z0tapbYXnl0Xt8KWWjZcUbU0E/O5PbUt1DXNA
RpIKF4HTJ9GZ9Zx1CJgo/haSBnJ/YhWIl4dYfMbc4DHgakpK5GDfCC9mk8E0qGb2E1fIHFE9ObWf
5fPOyek7ZTI8wwnMQTM/BKxJeiz44Gt1ZUnWptzFkVOlsl0o+bv3ROu3u5sloEYtrbfrDiT5VOqm
yr2mx2cJNE+MbKjEjWo+71Uk5+qm8TyWdVD5cd5mXoNlvqdZgfeIntSLO/ICX0ZCDLga3Ks7c3JB
EJr/qXLxKIS/GDppW2Yt45jiJhCDLs16hjO4b7fgEveUIi6e187uuIyazh+HmXpYo/AICeLqC6ex
AkrkgUPGHmJnCVo7PyLF9F2E2QfLt/Ftrhczvw7F1nDasP0Cmbh4gEERkDqZomeXaTf64+91eM18
CIt21Mr2i5+9lLOTHhwe3ome/U3nruKcSr6M/VihRQcgQgV9k1AxAI0XnA9p+MuBP1KWbg1q/Pg4
mST40dUMDQec3qUEwloq4D46vo/n2mHt/xGhl2UGRYp+yficRDtb0TG0X0283kb355M8aHfhCf8J
E7psIPW2kCoc9OhwPhNIPyNUqXaSzM+9poSSTzCP7HMVqUbKNZQ8H0WdEmakRspBwfeO62WGEwUt
26Jl5pk2J6ERS4YqZJRgSqHryjM3c2NH15Bvw/5j0QRX0y73CGVvxWNGjXfIuZ1rV8iSXsYz+LBU
YBQr+8OPBFzjLFX4pc6fqwD4b5LD3ZnWVKsQo7HMFdZBd87nOW1WcN3UGq3x+DQfk9s0TEHRc794
57HzDz/b9ye/1b/rz0AlPmmH/WeDCTn2gyNj50FW1pv7VGY0O4WhaGiIa0wtubmD9Xv9E2yXr3XK
0KJir8zlP5FwavuCBr8G9Fe40QPnH9xy5wwhSmcaEJ47Foe2bihj5sZxqctjNFF5X1f51HrcaHAP
bD+Q2hC4O1ArkQqBnqpYYaPUo54OkS+awWnsIfZQE1/jWi/iOj1gfjQ/UxaqroOSAw3BvgLMf4s5
RSyrdzXBBW4/Fg4Auk9y+ZulOx23UHI1H/KACJJVDEgY60hQxKdNp4umwnby86zfGbgzsB7IfitU
r5eRIrUyskiGyEHZSK1Tn3o11dSQ90mD1Zp0F7BSfdlhqKedbT6sunsor5Otv8j/MY+CRGNV47iH
Ashww8sNMnjA1Y9R0YMNxAAMAaUI5qo5nBsFjh+6DupwDrXd3DKyZjSiMI/0mI4R2A1rx3RZgO4u
NLgsYoO6Ars+7G1LoWr1FIQmd1qM6JUtEPo+XClxRwajDjx/Je2b6cy86JjV5zJkzG6MFt7jIqgW
TmkCpYlbJFyXooRAjD54Lp5oF3zzwCsWDny1oO8VPLZ/7iWVobu2ruua418Fup9f0PSDfJPvTCIA
bKxPld+yapuydzdfa0eWapIDcKo7nVkNyVFh2LLYssc9Ps4VcQdeO5+zR2xxLZe/Gov/HrqJkUa1
zLWzzrBjmC9L4kHAk8yrnhMHOr63tU2pLnWBfKg39wp1YcY//2n12RvDwbGWLrS/euTBm9jDKc7n
ma6Z/i5Mznp8IQhvuT8L953KFKFDzLc8nsCbrsWAn9N6NjKJffCwbd7MjfuD7miPChyB1TkuAcQB
X5e8c819jFpFN4l49tCVO4fMbC6WDsYdIrkN0fHiQz+rOxfSvCeIW+nUmztF9MkBkgwgRyCnXoQ7
USJwRwgt7LB9noBrRZcHPvXEy5FikmvgmIRdxbBKf9SUClke9mIuHj/o0nuwN8UWkSM61sarWfJo
I/qqgr0v+y4gqO1D+3BwTV63iD8mv3ELdwLmu1+Y3PsKYSF0qNn01fFZ5GveLlDAvmnCivYKn+6A
Splhe5IqTO1UEYDD4wADAVpJoDiP1gbCQrR9DLq06xUIWrDrdqygF1ffnsO66sYjnWNqtAfl0Yd5
iTWQ0AW35fA+hXhSVUt9wnt+iKH2SVOPlrO8BuPUBRs1fcAHkJ2zyDj4xhuvf+ccT0SQy8WI7e8+
kPB56qUSjh/OYtnxr5TR5cV5WI2DirNsQu77HIV0jwYlPN8P5qcR7DgQ10zR8vUj1gNJkVRZmlVJ
Yiy4CJBBM4xq+oXNnC7OtaAfnmLj8eaknFTk++ZR13fGV5iJTX7hJHzZuW1zKF8r1mrEXNQNlSHM
XUs1ygDV+4Bjdb4lk7glVn/1e5gkebq8+U5qJP1KFQkNplVC645AFPtFrwQgF0iB5wodQeI629oM
9BDhPGTnS7bbIu5elCC14n4UJc+gTaO/fX6IjaBr2YUOKCHBBUFYd5Casy3d+OeAEtNyK7s9JGlP
cY4ibGe884AHvX+u7rkzg9nXsKlXWC+T+Nobdn5EvIuDhtwrUtEGtpFs06zqbSKyNsP4nWIxEEO4
CV4mPD7XXiCs35fVrJaxs80sSEEWRpecWD5KOJc9lzHdT9upwGnrk4RfRVMh0yj+jajx20c8JzDj
oGxrjxuVqjv3xfIqfCpCQO5Z4zaN8RMJODXnaMiBMMnR2azAgUVYbfgCR7WoibHJ+Ett3Y7KLdoI
Iajb7HxVh/0099hnJir47eskfyFiHHW16Fb43OVeMhirbIdGdBdOejTmCkhw+glOPL6w0klkikg3
/sn/EE6xkOqMFOl1Ju+j4R/oF1XPINs6WDmpc5raKefnlY9Y4UUI7s2E9FuoQelVSzdIDjdX+WAQ
YO45I+x4G8SHjEtoz+EprgFrImUEkluDWkEsj8plm/eRAkCUUmM7bplRotlGrmZ1kOiJZkMa8laJ
LuUfsFcwAlQaZRPaSpL0gosjGmlMnLRu5N/kVqV470Xio7moG6B23fQ5/kw17liaxv5DIoCP2938
f01VLm8S19jsbZS8bd7MRyGwDz52xtKcfIz+qCANGLklpfMWXj74K3v5GR+bTHQL2qr0TiolMyhz
2RfJilkncP0A4HlLByR6luCaMrgNxWmxR/ZRT5JzjllqIpKkU8h2gMbR3mf18Gv55nuopekcrWvW
l/2zMB38DY9Wev21WZPYG01jnCjytItn6zBXCmp0jClQzcqiARYAcfQ0EjFb24afIyT3ISnCoTwq
+Yzgg49GVnugwhOCLdmexHmq6asv4JpYfCbhddq2DMKN6ZmrVp6uNtn9+gZCtMypaaMwTVgDuy6V
eCMB5brXnlk/ARqqKSUzDxaxVG2is48jD24G9QgduNeuo1Ec6/rCoNmwcMTF6be0KeWdV6QA9b9s
2lKKifSC7xERv9uBbZvBQec24c+zrjk786zRZ/najYmCgJ53HRvGQdaaCitbsbM7MTJRb7nb95Fg
gr7Xdr3BmylAnmLTHGWkZrHcBmTI8jsFC7xvYpZnfzHz8mwOMLnb5gE6Ux5hQh8Qb9+WHoqc1ESH
J++deB8cdkrcPI9uGwcl+/QKxIsnhJbaCkfLKvlrQ/zYq5pGH0hYktIwYPNnJlSbPBpu3XoRYIRr
Guk6WcDxr4UJx6+6wib4Fd7NUzDUlKGK3QRKqxP9HZiwKxHR1QFU/zHdnmC5dD2lLDRdAsY7Jzuu
aMBTeRZ8hvVIgQILcyuGw0YOBl5tb5YxJ6tjAxgP1acEHP1nXSlvYkcMr/DfBxFd1V5QpdXO+iyX
snxMlZAHLLW3liTBpmGCS84Ys8zFPMgKGXv5rRsnp6xZAGDJFKKYpaPLpLxa3vGTG8YuRqfwKWr6
GiC2CBQhWGviuWCZJO9KU7yRDZihKyx4FFmGQa/+5Oe5A9elaiGMZ33olICjQJUrs6EMaR7GcbFY
bIEaC642KnQQTKt5htrG2D9PwSxZvP/16uQn9gQn/Oi2QDlKJCXSrCLpFsqUqlxoJAkVDe4ltONV
aPgd8+KUseYACGYaR1+sf3Ybphlk8MDH6w+Fxq4Pic9/afROBRPlAQSLlXbO0nGWoHh1hfx4LroJ
e6VL/dVE769PhP44apgMnLpOOvjx6oRUYC8L990W+M85NxMNt+rYD7wCaEqjefTi3A+Vhs47SRWG
tGX7dRyEeHleX+N8ta0y9JrP1RcRcj74APxz9i+5ndBChCkHvHBXp7tdiRwHo15uYwca5DA2quGD
FQkIvobSo8QpD2qJRxXkDYTA5lFOCxoKqPhpoUy4G+icdbDquWCKjEej/E43QwS0/F1Fbwiv/rQs
3oOxrmncGVGIv5q/L4UEVQEvSEpLvqrHfLRh6B8zUiLmfSMIuhF0SqsrI/viRtERK4eRKlzZMjWr
Vy5Ev00XQ3/TTIkGGT0uDf6pG15Fy0EwFVrN2hc5SzwbrL9vBoLHwSkyl6uCHA4J5SQ2BARS7Gf6
996DRWZMJOyt+56QZv7uTV5fcGtCxGGbgx9psef1V9y6ZfvgGPtkT3PX090MkEOL7jf8hO2X6SAv
jobEcrLBFsMQQ+jUyemQMdRK+JMhuehWRKu7wb3Sm8iPI/5FRD/vQr8FO3dHtYdgitQfrmCnhQU8
t0gSRbGKi1Dn6qkVWnszB14vJs8d1IiNNVc7ZuT+uqe7Zwu93tVzAAHDVjjByjLasvqUP4QGbaST
MEQbAWWJsQ5UaR6eJmfzxpPa4GKiccdiKK6QTfNgYSZmib2aQJVkyBd2gu38H99DNIllt0j3xQKk
vIAmvq2Oe1iRT+xRiNkFlVBzRitR682RtNEZjdZbDnLCS44yun1KHUFkinwhOcyDf4DxX4HOqOsl
lnVd60AoxM/JgYJdIpNnQAvAMTW7vcE5Inrw/7GofYWW6omx8veX7IdhvjItpT/feRwuGM9lihLq
GqxujCKU+rH2KBXz5JxsAF4oqQvPQ599paOQOSz3TdkbBz2Zxik/EZQIjUSOwrYOSlsZyVMJfyjt
AFAiFLBWEznyUjXmxgmdm0GBrWxkHyfL1+/WExkw9xPRPoEaSeKLzw9r/8zqdqm3uXHHPkNd6eBe
9DUX8vhEbywetQ2nKJEWMNsoubeTcUfYvL009474bOyP87HlPX/UyLmC60XZQ0/smUuE6kBtzywA
ifKS+UIlMiUSlCuaPBr0oKmbC8ybJXZ1uRGixFOoTQK1gMKf9kcSAIGIAu9yXW6VkqQUstawPvS1
M4Gj3rA6P4+xWUyJWQ/bLVxBS9pM6+aXl1jL1u6dln7w1Q5S9aSZRfw24wTRJ3ZrLe+Oyep47Hlh
vMm2EL6J396JW4tTj1WokqGdy1GQyyZDrI/hfuJPqtnrwVgTA00wPpibkd/bkpKnMgkuvFPm0xtg
zKwT6EJ588XT3l3HwdulQQXza/FM3XNGdlUmbhdwz1YpX3NZfapycosFdy3EBg6Zihq92tnRTo6f
Hub0Q4gfiLKcUXeLvgDGl4rJr2rZoVRdX/eMMf8Yg7QdBGwvJLAEQBLNa7sgFVHPavCE3Ngip9Uy
FEodqLXrk86CKByNWiieWISwoUlLHTxbRvUsAEeZMAar0xxdqUeCq/hRp8x/K8gE14K4PI2Ap8ym
aa+o/qwZ/WO0ILj4YAwpHE4tMDyHnb14dL5xpzJYEOAP3hIG3eT28De/jRBP0VFhtGysuNjkzbpI
ntCr2FAmjlpKLh+Apu0LAB671O+U/1CG7Z7J5WUvzWKZj+YC4mx5faOZUgB93XV6oYMFSMhZd+Wf
awo94CayXCnGZaIUnMFqFUN/TafVqfRfOCJA/a//UjSqUpjtlDlM6aIP+C8ofONboFHvPA7R8hZ3
NH9jFxH8ZAfjclbHtmiExrLXbn075SI2E96Wl1Wt3iuiViT9+gBotDnWjYXCgDRfIj/EN/HIiSrU
86eCu3401wZI0/NJIXzR+JzKZLuvZbEWoxywpBtqBO8hYuaVy5mC+Fyf0eVHC0F4+UGoWnP7TO3I
2/dZFmPXTn4gxjwbX/hsoeRtnaGHKolqv2nT1mp9BznmfCf18RXbD9tzWiNZPFsP4NDqjUbE2vN9
SUTNqfdS2RluJzmiyDQYFjs20MWNDv1Unns60mxu5OLQepgjhqsxx8O5HqyGDGVK75aHz0Ui/X7X
Qr/ddJvZfWx+YRuYwH3JD6C2ScrUQIh3e9YxfpdQ3Dm8xfM727v8rh2qKTU2a/QkAzH1dq6yE+ag
6MpukAUxBpZYSQUTcGOrtC62ncXRitDN47qR2n2dinLxH0q1KFgvLsydNc4oBTu2PPB3DHNs9DAL
hD5Dz5e5Gii+CLx/kd/ByLf3+9N8zRHaLZ8APi0Kcru6z7hmFxVSV6D2W3lu6SSYhoK6qeKcto1t
dtopO8/RK5YKa2Uy4bb7se5CIw1aiajB3Iuzoesb39Nkl1Cp4G2sJ9huxGX4bSWaoE9UoM8EhJfq
KQCHAqLVWqes5+P6x4lWRIydgg6mkLVP+xVv7YJ88UiI3KX72nrqKmo8Da1TsoG3Q88yRolsCjRJ
FUYypMAd+rMcKxgr550KGKSGo4YJ7SVlJuydnZpjybgKRdf5LIxHp7QeKgy1Zhqwy2x6dNVR5gcq
F4KotJKlM09zQvZYb3h4B4qW7weB2XCTzMxVKO8mdYO6r2bdmqrtFEvA2sxLYHOlNyl+5R/o3p/u
A5Hn//F+OBQlbUQ4pnDbBf5udl2ZQvPZUb83IKFF13MT4TLFUaqNHw9Bjqv+JI1IJcxMnVXgEsbP
L/vq1hNVIHRPNNEEmS9YEGHbYLU5vRKCESbehLczrFp5iAhYZEgd1EW5cRiyvbtThyL3KpPK2V3h
aKofoZ4KkdRq1T0GvSvLHnBK1uukKXuFa1lycR9dsm4udZ8m5BNZJUZMP22lUHg+DnOZi8FmKLeT
yLlyAG3fgd+orBQxnr1rPTahtQPwaexW5mQwc4Z6zPvUelJSVFiYmpXjaQadgl8DoC8LKgukfD+E
NxiRjdN6AJGMmJTTo2/LjNpZ//eIirDjkAVy7iUmMqyAfZQAY+czdSjbsknnsG/0L5wikGkho/uz
da70wTTvG0HeiOCqBWQQ8k9YWnJsvu3dPeUxWe6B9NJMncT1s4WOCX1DXadVFO0NicQ5oGgkT4uZ
LSHx3sK/JmswbNXYPjuoWKn/U2Lt98EWLLvSZOeUA2ersoYpf2U25ro5F8FNZUNdZTQObCS6bfNC
/ADnsrE8kQRIL0/weQgfafsgQkKU6PaRchC5wVty5sfeEHid4psvadblF0MOWteV2Jc0yBfL4Os8
FvQTDssY9hzA84z9GLF63rUEttx5S2k8lb7Ivf218xtfYRQ0m/32GYy41zc3QcBxQOYYeT+8MY5t
rdBDUhxFe640Vr3tviZdmHXxogJlLg0rOJUWaNfjdDF9ZFbjHFft2WsBrv8+/GM5gNU/Vj3spbb1
yHYOkPI64wktikGHQFhptJJ7abX2NBDml0okFARFv/4uAADqbyWpckpYllPbuWM9r159ebN0kyEY
3eJ4hHFV5a7khRreXnIivRkq4XuzzeRRP3y02go9T/lJJTUyxzOAP1CIBcJVFB2Lp5nO0GQEWrgL
/tCOoE7e4wonPCy0IXT624ef3/1lVopXhhPHnA39AheXDnrPxmsaws0Pd1gVWd5c18ukleG5/L0j
+p6x6c01li1iy4SaUb9y2qieKJPYyrdffkNFahKfadvWYh5v7ERm30g87HshH4agFUzeq5LRKlXf
aMepkhxVXOMDHS+JsxbcuMrpL1OdXJa6WJCVEtkvEOX4N+Np0jOsrM3jm2DwLoIQd+aH3krs1dor
6K0/CFUwihZFhjkrKngkroQVv/EmeeU4MHFguZN/JtehLua+mvUUsV2SYM8t/70q/QqhIMPLbwcj
2079aZDq3/rUK2eU4ho8En6NrNW2mU9do70a/Zl+G+Di0LzODfjQAUXFVqHtdAtwIBbEKFGXYv21
vCOw7eyK2gWCfpT/pHMLQsFZOoSSUm6I0vt0eoOZhb/EkKRECF9UKvC1IvYBa6RWhLviFyArCuNU
JQaCp5ak8XacD/wp+sv0p04f5H1Z/95z7pxEwB6KNfrKKuWh/NVDrPs/6qnSvxRTCXHb2YsMTe+m
8mEi+Ln4JTP916R6uDq0KAuyp18gcdmaODop83cyIOp9Xkdc5vXaZnwOgE+nVCzVr5fUirxqQhoN
kXw20VTHk8TI74czD1plLJGzZwjSIONeZ6237v1FojbB63EdoyKbNlq0wPAH4yCVNshgu4npAJoE
OOwAJVQOW3BS1PzAxj3B5MrOOGV4Wol2d/GSNynnjoWbt110PkoWXfu6WOk2O3/gcwPBKuk3Qes7
MZY/QN7FfqmQPUTW8AzzVh+WMm1bFM1ngcoMJmS2ijep2ouMJ8qV/CLnRt6qIHttTg17Ph8ifovW
S3KnmsScdGNfWcPPB93ht93rHFpU8FqTKrNCrc52jPZl2uc4x3DwRpZ4MM+bDmnihTAso7AlXbsv
BI7AiXTqsLj2SGR2gZYcWOaLj3dKFSVHYJWpPjVhK9pozZmE4vN+2285PhOiv8v6EBh7IXlfKTwK
OpyL8cUx7VGbwQbiJFf8y3MUTgRZvOkYssJnKdaG0GZ6npUae8JefVYlJGtQ42GspMBPlomPRsew
/qDC748Y+mdWUyaoM5tbQDWxRiPTTkn0SiE7lfimkADhavcg7eSgLRoqT0EFrlAySyufjyWj12Cv
gDO//5hFvJCMR1i6ZH0ia+a+Siq/RnZjE4dkDA8nCdJNFV2tMR0KPnSovKkxVfmVG3xFw1vhf96C
UKQPkxYNuzwd5OIkwA5p0KX6Zw7DWMA5/KPRDlevW6Ih1WvGz6XyXHK0H1uMiJS4aV0V2ZSeBIcb
DgGOtI0Qytt9ryEhVJaQI/xzW5J3egwtW1mmTSKFM4sAwy1pl3w32vKhnZFiKvSsZ8fd7wIuBz7P
B4/P7jmoPlXcRQgTkz39xFaZ0hBR9fKhMlRN0EqX/hWkZLWxncySaXwMrXgzkA1U6De5WoqaXrVq
qnO6nyX+eDRMShNlbYBjQdRWiRFiaD57BeS7sFNlkomUrLutucSS0WKvTT5RUl9zkqSKbdDNXGMt
CmJHjuL1lURFrjQHGRsTbSjDdR57F+hnYiMDiymxL2C1tGDpNV6xDBg7nxcWYp8AjSko+9ZGi1rh
6sVzd7iwqsGF81rGACaozHDWpg+XKsdlPtnxtxsz+mipPkahIb31J3ikwxEr6+AO0jzua0neR7WH
JXKAWL/nXC0vXpvYfDGcQp43G39U8nffAfYz6ETE/XcBwhWpDzVKjlQEwCihCyYtERw3JsIO/Rvl
558iP57pqO16crK2dIV7gLlRjfkY04634O3Li6kDOe71Km08f5RYZPRuypB3f0DgQIUHzymRFhB9
BWBqmtKVECvwarPqjQDYy1NpenIBdPwBDy6EOWb7Q7wb05q/bUNhTcfU36soVU/uSXKlpU741ObH
B0NWKhHLQroNdmtSxHaeIEAc61yCzFn+JEXgYx0L1bp6ELskihsC7JvbuoD0IksJ74jTZvshrRE2
cPsEqLXuEI8VIZsi+xEdHdpDloN4Ova3MZtkmD6cp0m29UKvXsTAQXxys8lT9mIn2L1BPmc9DwGQ
Jc2358OxClayaZzhS+DKgfnKawz3puVHLvOcaJC1JPhH/3ZS8Qku9D4h2i+PxmpgUSnRmV7HuyqP
phtFVm7+GV99NBq/dqFUlfCQPt6vN0RUmRVP2VjmhJBf3MhvMUGmuRiTkgIKdAoBu5tSeP6rsSQG
3s9vJ9W3xQTbHU5B7HcQpeotO6trZZY2IN4aYxJGMnZ78RAX9v09rcgOtWlqeXRychHt2iWwieYw
G8HB/osMD9R15p6nIZ2TsQflbqG7FkusGDEun3Tz6MfPfumqPeQ8y+OQlVsccDJy6iEF6GQNx445
xfEy8eFZDrpm5N+lIbtV/Vh90Y782dA5X6pFlsQQlAEWUOeYeWYkjouHD+foJl0iDiIts9Wyebu7
hJVETEhrqud9PLkQFGvLMd+b04U/dgw+Og1JE6/Mmx0NbqPgBCDAVbAtczJJXRoKvPHM3nykKVmC
HFX+PHP+yVc/xpfXV0NxU5OjVcCbYB3HadPQeECI5Hq+FRBmjB0PYPA/5TJrzOcWFLc7M4M5Mpwz
g/iNytjia91u6x0Ur+TXTiJTpH+hYAF15QnbE6F48KxhsQuUL7UTQeltUTKJpAd1AU8F3Ai0zSZr
0IMdfNAUZ/e74XYxjLz6SiXhNopA3ZW07tgkeVg8WhH7yDCbwyLRzlaAMG0GeaDAi9ZK0ZSVpkvV
gi9e8voOji0/27Df8E5kk1Nc9YCjY5gIYNhHO3UJbkpdXLqFSR4nBPxrLYhOlPqYLrm09B3i3EE8
sMfKMyuwdt+vjJlHKcgmntak/2pAQP78qvQWzElsjiFQPzeVgeodMIUSJdXiERmZp2vh6jqfSw4F
gpqGm9Oq5A1TS7Psts7lkE8pP4C7HmFuRCWTaXjLhqdhFEpVi79wzmHAunTVu1zsYnbN64ONxGCM
H5F0lixDLotG24O7TcplTFpVkIURIc8CUfUT/eIEGbgd26AWUhcq4mSJ/FX2+82ASWibNZopEnw/
mEnFgVfxMJM0aWERsund+l6dKzYNYNNKawLGWRYhwIJJJbuPUTIJRjqD1pMk9ZeX7FEdVwEu0aZC
k/sbQu5eBbxaEJA+uM0PiBZKVqX8zH4G1rfqDgaQ5mG0t7fWJBC0Ypas4bWtHFFpAxgCGW81LwXS
hWgg0T8q/KdwqLgCgcayiqiX6SfZHwb0Rg3sdIl21/6zAZhao6eZSwtRfAT2Ny2i+T4pSmYVi4Sa
BwCdvtp8dQkv9NZ5MuoZPw4Rlt7eUhiU+CErIETInhLtNCJGe/onB44gejKZECg5Mzqpee+fO8uK
+ZvcqUh6dwomE7d21LHc3nxXgiADpwg5vEOE5SrYy+WCWcyA2oQiD28jj0KGjhMJ5FQ3NsO1ry20
+Ig4rc5X/5PEiZDIt9jT80p5u1IWwVW4aRGt2q19AVMOkh12Pdd1816xbF/tnPbr0waomdVgX28b
VRh6g82XTmucAWvgAVK7emMel42eLreRVgjylrBTET+xQOZjgY2Uu/Mdb9CBei/kGkLAdd6FhYFP
yEwR7k0gXYtBthr+ky+LhcRcYByY1VuGw0Q89gXgc8HJAwslNz8QFMxZ55qs1MY1dr+AvARxjz5H
1H/OsYfXJpGA1wv3K9JfM2gmmw6kfJYqF4J/gjwrcIJd/Ix41NO5Lx54AUl4VdK1SrG47FgpUAyx
PCKY1WA4SuEsFk9EgmS7ividHoAe7UKoYDFaHO7VylkWgKlZq0MypeCPlBAVnFDKO2+oQ60JwKNA
ttCRdpAICq4Fr47KZjQvcThmGO62doNkbyG9XHvC70kAwpiiQC9rsQeCHJThVHVdrPNz2gToqY/0
oRoOMmto54nhb6lODGQjicIMX3ejpT7gwe+yfW/dWPc8SIZSlC7gTLB5i+gANex6RsdtkYM3HAOz
wW24PtYye+QImg7IxstnKkKyGfk1p4hVb7JNEz1L/od13mGwsOyxXpyrBBOR+dMe3LSoBqQa7x5R
YtSYZiNUi4bXeWRc2RHBmNX9S5LljF6wmeTCoFP8gg/OpfZdAQHQ3oF3MtUd5vUAx9aU+2DKa72B
yt629VxjRYWFvg5v1THKSl1rrbTqlrxFT1H31viXe+MRaT5pPgUWZViyhmd5SSrDa9zwj7INtnwK
0m5fYfFgeaVtdivnhizp2VxXASlyAkNvLvb/oZKrBYUADLShyBbWIwaTqTiQ7G1OQk4To69dVcJX
mRZKFvjR7OBeYEiE6j8aTGwbR3xlw1AfmnjWtPSmkOq2WVQ8EGQtGHlnt/hpVb3TlFpF4960w/JA
IuFFe8AoUPACuvKMHIpnx+yRDr36GqsHoGSk2sFyIPrWAtt1Z7+sZSpEzMhGEeq+DMamQKmLZ1KI
scXfDMHiz1kcYCMpGtflp3pnGnz7tCx2raWgmBt1sFRZJuz9UKjVDtYiH2K+LEUQ5qgVCY4MUL9Y
eYc98DVU8nzycBB5WmEKo3TM7CryZUl8pGY04MZRo59bWyTt3UUZ/ddYFpzSZFRfYwSufWSSPOlm
L+ECk4tsoraMD7CtOgiD4ovdMBtxtkakdfC5Q1UZdJlFJhUnNzwxU6fgytVqHRo5e17K1p5fUSS5
Aug/egsbuG+VT5nch4+BvMeA0qX/0zX8AftyB84gNA8grS8r2s5tYBvAEWtv40DcKAq0P/C1mW8L
sLlRPj7wDnvyoB9+2wmDhYqjs3+TzzH9F4ssaIK+vt+xEq+pnXFc+zsY8iQlJU6BXwFOUncoX1mu
APeyrwguiPB0QqL25v3pn7AN3KIkLy6B0nJ95svigandFDEBNbdscNMP75EmZSvuUcMAP2E5eDYC
zmJxX7v9uJL12+z5FVW5WtVJW4P2Cs64abV83YandILjdAcTIqXt6pWD4wceLRDhJrtJsU1aphXk
NV+6bXJOI3NnR3uiEoiz/GVTJFnfvyQqY7cpRiH2/UizqWOu4q3bQRVXk5p8+n1rqEUoNzlaGPau
qe/Pk9iz2M97sMQpRSIOk7T8E11J49iy3qhwJyZyf3qe83qus0q6ZxaDZ6qn2mvhiqglNBbBemLe
Z2A0hev4I8TFevOlh9pidP2zv85ExpS0oWRhCTGAqQp0Wi89Ske8wcBKsXFNhzv0b9sWudaICDAC
g1vqKqv4R4mLErpIHkUjbCuLC6yhb+6VTezjOWV0SkvkT8hjtNDj+OcyNnsrp7INOFh95m/ibNO9
8DqB776XE8usnj0grqEAN/y0pMzydDK+nQ4BJ36gDXszB4mN9Coq1OH+HiDuCSJg7a5iFtADMKot
82pkFv0zAot42bqSCp+h4OTWExPRx9w9Oitw8Lxz0JAEYdX9cUPpF0wiT+ZVDtVhQIMvxM5gNHzY
5riaq59MbeJYovuq8krMHwFhH+AdFePTjNiR/AK0J8rCJMcV2cWrD8XYufbbvkaG3Ka2vUEhl12Y
MoMmVU2eVDGWPdAbxyyKqwntTviNMAmLPUQSPloptbmXQAsfuguOMZlmVxV4o9/k8s5cs9s6ZQGW
iO0fX/jId7XK2qQmIKGUeJkuxgJcjXw/4fJEMWCP2NRT7kW2yg/tMgoqiErHy+8xDtFa+8NlFCJQ
cs7AVZORMThbrtq7dfqms4nPE0utfgC42qvBDQDKufkjhwdK8rJc9+sGS9FX6h8NpEHVE8m/QwCs
LuTRPot7PP+bseR0dYNbE9IVI2g7Vkxlzc7WoiasKxKNr3IjIoe91tNJF5ogQG9WizSgK7uRb9DZ
owat7ahbrxw3L/lBO78sxIF37ue1ohErYgHchjGnVClwJ25GfZN8jnB9FK1U7sTknSqZ1E6/LTAO
tLyJqauMai4jWXU7KM2TuLKt9u0lXgGkXmDQaD+W9NVE+QyIH0ydmAJXwffr6ymz2EjWbzR2ZldH
W7uZpuQipftkOqo2UzXJ3Mo4vuk3WVOlcM+XhdG/pXc1y441PH5rH1in6sAqsaLtzp6IODB+RbE+
LIHASw7OCnHCpcSS5tj2RVMtzTMjn0R4VW7EOO/cWy2637vhEQFf8xPhlPlKFxKgSuHlj82Wqc78
x4s8469o2le5iAZcOKj1pRo7FpEQk8s9WjO6pmiNdIXHFkHPZnk1WHoPEoTD0mCUeOI6CHzzB8f7
jaXhyqJ72pXgiQ1oxIEr+oYmAX7oj1QjkaEdCfgQSaGURRdt+kxAmF3tEhQefQjPIFxywCy2eeT8
uuzYuOXY8aqq2OPSrL+0XDh3GTawP/oHyYLy0LVVqhcYsOfUbi35FfCY1AhdLkbAd/WqaSgv1SxS
DbpOmKQnv/sL/UQmXzletPn6RGjyQIlvsx72s4x7NFuXlVHjqf+n1e2AbTfX3q+acxE6qwRrIyLU
HsJitz0UXwirXHBJRMDxOxshqOgpZy1h41F+673CPGM9zHe4Mkl1TeME46Z3u18SflquMZCJIjUe
sFoqUkCWD21hCX6Ub/lFDrXC+ZbDiYbMSgiXXkvd5wEgrA5pspuMDwMeK7gUnX6Fj2R8HXQfWF/C
9pshvt+g/w19olNv5OCxWKwGL7iYTQugAI1NGgxDEb1btvrC3VYKLTUjhPRAe6YEjwCzM1K/CjL7
yP3NtT8ROYoeiWO2z8zG2ktmxSVj5/h7Ty1c/M3b7Hsr31hC6PzoTOSxnDSB+unr+2KXEc2eXrLS
PxwyyaM2+Rv5ielGMap8TBCp9sMyEboJQYpXrPV/OoDW2sJL4bU2sdpistG+FeIJBf8fy9CRw/L+
8P3Q30YvZcKWzMhOdTwwXd56xX9UHzlzAypgv+QjIhvEP6N13S+y/EUeN29tBdgfHkViTRloEZtJ
GNRCcQMCDm4PCt78A/TkxSDv0ZU4zJHh/Uav2fAN3fb+6giPio9m4TtaHENHMFNgxh38vQNEjeko
fTUFENHTzl4uoxmp6+XRF1/Woo96jtr5A0WT6oolMndS37/roB7HYptGIQB2TbHEx9YL0Klw6wi3
Twnq/l55kWtPoAYsN9wpvdX9qrEUOV84QKQwXrQexkeF/wBHrUPxSnAA+UodFTlH0lUyxhVftLQP
OgMDHYQ6tiTvE2CNrIuZU10rMpUfI1kfRyARDw1ZigXqYKepbzTnWQrvBNaXQI6jy69DvZvlv9eK
KxGeag4XnWVC1QmfIq1OvMTnWiffvuEGvioX0p8g88lYnuHs3lM3nNIS/myPBGzbMvnwmB/w764U
YcYG0P7WHw1XfQSdPClhG0/oGjFDay53w1ugtugNkDepFND4jWAqWYs0aDmTIwN/Sl9K3YvkFhg8
FE+uMv9bYXlwx4SvEr/PWMQ2NVvHIUAOgLET7WWARUi6AIzrxtp100S6qEHRmNo/gxf5Qeu4VoU6
7XxClQgCJn6JglNmM7yHqylnDD2gDOCursXn8qC88if6lnpgMUZG0YFbLAFl+yqMrib56PFXV/sp
J2mMzbAvNMbUR2bh4ey1kMl8/bdDTOo9+2TeMyaObsPaja8SJhJgU1FzlhP7fet8MFXdOYYYanM8
ooXrM5K5b2+0iLypw5/FZDCN/lMupVLrd73nNAOJYSTCV/fMuT49FcwJNjbdfZJQeab+I9Zi3Bk/
Dhd2PJ+MQj5DRXu+PwuTSGXTxtPze6lreL/x6il4suQDl/HTR1eBV2TjKz1jvnVqhlV49X2sflvg
hVCS2w5ryUaL/U/UpLQ359DS5XNkW3g8rPNQp4UmqkcSClascHN1yKNJw1AHGm9qQU1/rFZDpJMo
hmzZnyBbDgbuGOn99KuPjSPJdVihNYr53ZkAYpnvi4D2GCaOKtXAWq0DLBjOfa/qU7BtFsER4ZRC
7mlA7BT9dlQokK1q0rbA3e8NDKhpZnmNuE55WoCvLukchkrwZkAEoJcHwTjM7bDGe2CHl5oCtLGq
khnP9JQYLGi3aojgEySQqV25l7rSz5mwBFf3xdj/cFzOn4A/EEXP5aqio700YbqOtEF9yQ8hbKq+
qmpK3bedovr2fKUTHV8BWQZKvj6SkGTTPF6XH/YPzjKl+fqpwPJvUPTPjPf8fbTvdld4/9RIQ62l
GRMnpVJynGdSvSlSNRKXUo6xmxY4RR3HQoat2tJcA9T5AEABhR7XYOV8fveXnI0drU5a8UUzLRFs
/0UkR4d9I+efL4i3j20BUcmfVPY0047Xcnzzzk2gB+lWCkf2PgOgO8KLDkbQ8QnWai2KSCwd7IOg
SFtoxVzfkBRw6r7elcq/5By1ibXlG/r4Vt+euAKfJXCIfzYyCghJqArkY47KCOo+A8kmyZe5ru6d
L4Q/eLYg5MR2UARurEbzWwEW5LMUaI/JY1yXzlmJLp1zxA8JTvHVc2nhR7BRYRHAKSQuVwo4Nd7w
Td+iKtK25Tuj8sh9cYEzPW+9E4P7H4UucZKOlvkMZMx+Gcu7h6gn2E6UgWfQQB9urB9erZ6dtFf5
X9sKEQhJxDTnielyLSbUP2n2je7sGCuB0SC0A2sHitNsFjdX9t1bpfgrLhbiSJJbLO6OnDrs9Jre
TEI0vft+RW1YbI2N5vYhKm0Rg5gqKXfA6HGLGOHDFQXEyRBrPAEyQF2KR1IApG2giw7hfwWfUG0v
l8FcNcjp9w1ooI6j2PiiAwV8vMVofx6d8fi8sMo5YMcnqKwlOLAanTihcVyTel80dpdJTbPKNxml
0jjZt9Zxe29ssaUbpM9rxNjyp8JPnLpUDRaK4r3wDwdrNgjQxYn63NfI5+ofQXscTHKRGjWrducg
0FhbUdayxn8p56FWOxyn6g6lIpwYBZVSJ28fq5XewARSuJGbOkSjc8YV/pyARlrWmwW/4jI8cvEK
jCiDHwO/ODR7CJPAf+U352YpJZhhUbkilCQtCOrI4UMzvlagLwpYlM7Sih8pcXetCnery48lurup
ksG+3x63rt8Zj4wQ2kBZQB6FweHNrllNtOa40yPiJRKwdmIfi8zao4LY7Geg2lvKlpMl0Iq1Egyw
MuCx2/yz8nZ0AzNKWSGYx5NdK4wg5WeuJzUsU3IfMOfzFD2OFeMeqc34ItbIufym3Mc7+rdNaCGl
QrJbtgLnfJh3GMNx8itOm0rdBvwBplkWzEmV6QvjEEAmMSU4sib/ZX65N1Nz6kg6p7y496jrKAJw
MRk3o1/7VIVDS0Snf3FcMsfrpwqh6J8wPn38xN+Y7hgjGFTYDwkibj5/YrEozITWivYSrgr8S3qH
vsUjebGuOnIN8Wgd2W8PATqxHziTOy+mf4zppPT9MuyW43B0e6SpMhtH5ruS8lgkAfbg/wQryEe4
LT8Cdp7JR44VbYoZf5PA6lBgNVDYQIL73+6gSRqYT/hAk8HM8AOpBfRwAHSe7GiVt0+xvZdCG4Lb
tiURe9L27OI5nO1L9x1FRShjBA+w0bfBzPQuE1NdYkQ8ArLE6UvolHQcCwIkfbiPzK6Gdbn4JR4F
T1hGhIwRyyWOF/Ffje/eTHyn48lnotmbMV17rdC22zkTh9iJRiQX9JueIWdH0FYafgbOmMqbHOcx
WYVivS7dj3KMDh1cfUuQaBcRSOJzPdXJQB7y4oFXyJ6cVYN8a3KsHpGDyTdwN6VZLFV7n58sLwZW
H7F4wD6mIQ5k5gu64bcJ6fVBp9UtaNNviL3T0yX7efQLoPISVaAIUdvAbSHc/UKvhjEeR6D4xgKu
7TTY1yyLHQjpd6lK6M+0aD2lPj1ykVkgilKzTm36p0DieRg+TKEpRD/rzw10xvvYYpgA9bBR4KRT
W61q2m4S+sMa3oXYCs9QjJJLFXw5j09+bwyCzwLTbFPG5kV7F+oKzJnWWxw2LKkWn5yqWzGyIxDw
dsijLut1Wjvlza6cfO7dihonaklxdJYHEWzvT2cT4PIavWxTCKR/zlAf1GhgSY2QTl/acNPoZoRQ
tQiKA2FTTZoW3EKOLk3TC431JfgYd9FBCVrjZbsJQeU9JE6956VJTh+ZacHgPzKYbPGQnMd4CuSc
r74BuVydJX5D+kP+TLMzbYfW1rxESIuvUoPPHu1kHZwnsM5Uvdw9Yid8QufIQ5PRyUP91pSg/ljt
NfihDHUD+wVrwShEYCFLqY6OU7slMyEOY0J9Bf2p3cFc3HaHtni20/OX0iyJMSdptb0GgspnaIXj
EnnVxRwVqksTGtsf4sO2ZmFy4rp1b7EEU3NFt+aTPuXSkBsonWDYQa3okLDPeCB4A2zo25ersBad
lUZm4MxUbjlXJWNwjGbQXdGLbSvJ7Ib4wnS+abSsph15uXqMVxmHRhWpUHXHsmi1zsDSksOg88PB
7ZzmdDFOD1xa7vp1iJab53rqWpWGnFn4xvigVacSLkUjg9UV5gwA2baW2n8e5fbsbpih++HoQ2aq
rCUkK5UBjdSG7i5YBhcPkxhttZys2WuIRkBGOFJwiAmTII4Ttr5KZF6VFqUajTXlrkqIWNWPYQtK
8iv497aIKtqsoXC6KO+8H3lwb8FLKfCX/C6H9q5sUe2LF5rivX/xF5Y/dQqDALdSdXHqratSxBbw
DqdhlmBNTre2TnA2IeC6gQShbU4Oo//rNzthz+lSfWyAra1marAiQ9++TJgBtIVndU9UOKz9qJLV
KFWkbvqU3zYyLxbb/1r+B2Lpo0L+4R/iFgPouXT3JjRpdFjfAu8cimgrqb9aCNuEcJJnpBV9V8Dp
AaCnp4jBAQt1YXcHyfp/Vlf+OpQoC1kl/CLfzg5uBi4ifs+Y0NEnlmmWzL3DqxS7nyGls1UWYsNH
UN+J4mpEvgnA3apB3rAbJGqelViiLuw3r6E86CO/UWK7J0UuaKokrQENpmWYRsvyRCqr8mhayydF
ASBdq6Bow4IIbzRA3PSVV1arEYZHzM7mcDqNZDaeG7EkbBa+uAYdAFkUBtACJcoJLFjZ63xPdjul
WYmkp8coE2IwcMIfGN1hrkyJ6q+sXqJBMFv31B7BIsNOTJKICiInjPcaB7ArvC69fztzcCIPyf9Q
SB8D/QflZ0nvbSw5y/jDw9W3z2NPUxwyr8XB5cc5Ewptolwi5Gpo8xgAOEsSUMio+HfQoYy5QWSd
1if2K4BBU2D+/aMaTMB9nV3imEpZOeqMoOwg3gCV+eHcJcAzSI8CwID/ON5KHPa1OqO3R4HlVcEn
mQBfSlvds0h6IKL+ABn+tGnCLXvekDFZHMEtwfCK6IDLg19qGq32wLbW1pVXK1TEDZ5Dtn71jSKj
0FUvaVuKWtQ/pIHQu0sHLeGNNBwbLPPKLfFtJ/ujGHEZwEcJ1XIdA3xPY5zPgML30rtEElY+ONYA
DCm4suvig8f2VwrL15psDIlajA7hPRmmDdjOycrmhtA8NUSRIRf94m3cYSHJSXi+OOllWOwXilay
ugXa4x4/JTk8Gtdj01LQayeOwnL10+W6L5nW5eGjyUwgtFBTcpCVDMFFnDBO1U9n44L0IbRiHVPm
pTLlGThVVF+SIk30OFpeP1zH8edaMpL+reBXLxHFmTTyogXd3TjI5D/oHk1kdg/N2my0vsCK1wT7
mE1gyeYneSK0afK5ZxmtQ3Ub5aLLG16ncj9wMjCGuMa1zLmeTfoBGQiQ0dQXPTTpgCarLXVumkED
Ok9obZ4b46vudZPQE6fNzn2F8qNl47xe2Ju+HKiC+5SFhfpxVj2uLW8HcCKgk7nFewYNBtYrlQwg
G9IvTtcUF3q2al+tGsT30IXrxaQhMCr2fqOd84NssD58aorPKQM7DNB+ctyApcH6iRNSI5cnF1er
sJVEpbCtNv/IXwfA+79SXQAjk/5lqZ+RmnyDRGZTISCIClAcezKDcuH2Ak3D7akLtJBwNoRQnsd7
85F0Ar30rxZntN+zjpp4aPmkmr66Auqi4YXddFylkqES0iALJ8+4fWEMvJ4V1AxTbZgxtVHFKziA
10Pm3KODXuQY8qEX0Au5lobxADZLU8cw0YZJfHJ8Xc/PcqysXdwMD+jt71QY4vMsddjHjoVpyKzm
A9rGp0ImxGkziN61lO+wJ5+MqY8eIQ5aLbUMo4qDVOXCJTPoMQnabTiDfEYP81kSIi4aYhXouzlE
7OscaKaU0rhzNzkpTHR0Nv6gRzEElPyPChkQ6HIlcn36clp1vb/BbUmTWbCI7CEK9uqddAP9AuMf
Rd+fWDMS9vRCX545Oh9IBuDzLXQTvI0dzcnz2cxJov1IR3vnN8l1Kg3QVpE4cjo9yw97nBhqpLeA
jKh2tFub6mG28M8WAdzEJT4memhfw4Zwpz1hSzkpMeI587dRCn2gXHz0LzflFM7wzYVPuQPOdSWX
BlrEbBqZ/SJrxTQRHVXHiRIPx6d5G8BR3ghT3nmzHRGJlCprc2aXLlElHXq1/j7WFICAdKsB9ZTR
QnaLMGBoIAbdbgLFZglVoNskjPEtJD+ztv4LSPpOfbIawbxNaqdwjeumGaP+mBmviLIhDKN+c0Ms
owhG4n79zERp6EciYxNU3Shkdv9J+nG3FUHZKuDG5QSoL2eQbrOOv4Z1DNAXXfFd4yFwRC39YDOW
deVOQQ1YsWAhshQG5z+WEx3Yq2G2CJ1BMTM+5V4DaDfI8cZ7CrFz9Qzvx9INPviK9nQ+7/rozXuH
HEBNosDZIVMVcAuBSMahLrj27pf5bNeGEpuLoXBYfa4Rv2LZkYAWp4u8Nge2jXpr+C5T1KSFxNla
tvLj+ukXPhF/KJ7+KEd1sa8/HOIRuNaIVSgq7+y2M4tgLt+1MPue7YCcOfG8T4Dxi4CMvtatJt7O
w03dxQYVkO/Y/e0jBBIqPr9gFfTWjqVSpg+4xdjAW70vl7iIYuaZsZOC3v9Wc44/ob3Hyo90jr9M
t7RIzN7s3b2FFjzqAnJzU/p+BaMeCVTgwao5EVs1Y+usaD9/hepc7syJ0J6sQ/KyxEpjO5aqU6ra
ta6ArRnDS+PT5r9Uk4XIGoAcNPsrX/Iv61mKg38cY5HGxAitQr2gtw/0EJU3UCF5s1cTG+shaVJF
4TFlwYBwCFq9MinXzzJpDFnHvR6aqCFjtKmuaFvwUSjeP0CmSg2BUtgWQ0FBZuXvJ6OuGWh5ia3e
r5Acp52N7QD4B3J9y30cA8+IwEEzkodWyFL8i7+NAuOYY//tMK8FGfNQjIwWGqsS6KmrpGP4HLdz
Izr4pIl322yo5YT/bR41+KmDtZmuGKEdpLnk8JuvaAQ2UGdHyTx6RAfgcHEA/unMMAIKiDC/I3H5
D31+m5YAlHDWzJC9b+XW3wep0UjS7uNjuHJkNW8F+2m0aiQxNru8AcHXDETYmwN95An+00mebWlS
B2ARkGkVxVnZt6eutgnnyQpt7ALEVU/q9L35EWIFFEKzllxbeVumpabjTdItBU2ptszknltgnspS
T7sNFLc+DzizqaNBEw0BgeZjfi/42pw6YOGkBs28eWZ8XJgqTAwP2vUF7umGiwZ9Uzuy5gI8HGP5
T5hEN5/hN05veRNoxnyCe/HwNF1u542KUN0CudnoQIp8AyCBqF4xtZfOl/CpM5mAnnD5w+BRNEEo
mWZAAmRtfL+5HPE9QGMKIBICjnleDKszQxLvzwdyOzVk5D8ivd+GEMkWUOm+YrLrIK7THlrWnrZn
qNafDj2Of6+IFfGVwv7qgIzWLiK3zNVoKcIsSew1EExtCDcn8pKhKm8zT0XouIv1NiGkry8i/WrM
oW32F7F0/LQQ4hgrRRRutBxyUMaYBo7zmBMPNq9I4U1MJ6VhWtMcE9qc2c4ZA6FY/VuI0FYjNlDC
M6qS+rme8ghcd8t4PmKVzc1h+GQrWdSe4BLKwZ2+rpGT18yfIYhFkUw4mbb+tmPNYoHBsrC/Pk35
FKnDObbLfCvdvAZ1dhBupNFjm/04MkrtBdjsmCgLDMGL1p/v2rQWgPck52Tc9xTSAV1MQNX1eHT3
u2R3RACYtKV7TQxm986JJlxjKgkgSiHoBc6WhNZkznZZnkfAc+dC3gd4TcZbC4f02q70zCym97r9
G0uScdfMPkpBbTAX1WDToTnTAEK5gQTERavv54/93e4gcrTqMj7Ozoe3vGqjQjItlby0OwIJq7u9
QybrO4FqSowfB7Xc0PzZyZL6sv9JcbvEy7ezBSLNkSVU0CDL5mzbdc8ZPk85MdoXLwNA36e9rtWF
AQdcPnc7xfRcl61jfpcmFXz5TkHUEzseg3bbHtVI6vCa35Qldl1MOkWFYoYAFgcB9apvEefNhdAL
rd2e/AxZjXMiSIGbE5NB3gd+7p1JVRt2Z4F2qLCjBjHdxoXvGucBKf2o3rR88dZ5vtRGDoyuMwgm
8KQCY71S0iErlOpFuuFHdxNHLe0bu+QUV+GgAnw6QdYqgYlw5m0nkoCUfj5c658qSBLoawghmlfK
DjAftucALHkVynEpFzAWQcnB51QruimvP/N7DLH4KsVA3LrwzrsVVXbreGrk9WlB5lLWCSFbX+HQ
AaYlHThlnB6CQWlZ0uh7NOdhYzEOPWvd0STNfeFVW7l+qeklrnMBR4Cwf4dwUOMr8XXzIsdWqfQW
IN4i2bYzmdXUyoM2NN7ZEHJsnvqdDp0eGdpGsrm6ei5InIRnheblh0YqNSX8gxpGChrewJbqd5SJ
VbSvwREpADZn1z+dLeF3GQ0Ifl0Q5YOy7Mw4/XbQKJzoVY7iNQmj6+HB9OL1pF6Z2tZQC3X1LFT2
pJ0w8XKn0wPQlnqpfTyxCTo0+8Gc2pDVHr/hWaw5XdWHKG8hoMQNv/bdmTsYqiOyxlg3LWjx1DWI
3hpFCLEWP81d7pLwkBt0KwY+9CSraIfYn2VvRw7C6YQqlGAC1I6kK1UAey/VGyB/SSKee7SpvBWx
nKiw5djIqSmVlU3z5RiW5FuMNMqw4MfUTbr4F+kYxKZESX++XTvt2sim5oHPTo9I+s1P77Xl+8Pl
HRnbSN4r2aucmX6TDdcErbmwmQYdh7me9vS1IGbczBlTD6o299bKGgujr/xDgMIT3AL67nRoR5xM
Zf2v+DODrhy7Fnb884w6olwCMFqB1Jr7jzpkm1bForh9lBynbMBDJNhI+Q3cRt91b1+h7PIoY6DT
lR/Gd++ziNXmMpFlTLL2gqW7Fc9gFdqo04Y2+Ph/NpT4/tg+q3UvregBkEEqP+kio6IxF7KPkuV4
9JihjEpcW06+K1RuZWlFZ/wV4eklq5IoZyCjRlSFrWAl1c/oy5DPKCiHbu6CE1PVE//lWzGKkEux
sS0Tgb3yXWL8JDkKzjADA+hETJ25B0D5Wnu9uY0K8qoR4+fbP0iSJurRkE2wH4vQDbMxmPo1Taq1
Qib5frHU1uxYBCR2TS07gK3fVI7i4aSPFR5L9N0yVh8JmD0+ARladFiFSZfuxULvD4QKuT3Z0LV8
MdenRf7VmkjQdgihxCTqgA0ema6TqJoxXuL4ESyckwiwh9jIyFzsBGpCaFswKX1SKbvPjjzd54zY
FfgclXqN5+i3VsrSlWMn+jqMvCChfU5tXDpPlRiqzvRUisDr/mhhaLkKOM29WAR5u4o4LWiwJxnz
kasEQ42g0Bvs+JEgdCo82jrHspt2GxzggNV8BDFQa2T3LvAD4PKWcH896LUhBvs79cs4dAB1uVQl
mEg14a8IMQQgHkWBBhALwfJw7xMpm1zmmq/9V92N+B9bjauYZjQZS3UgRYsBLTNNlMp0Ljie8HOi
cX1HZc00wLGdSvKlipVdXH37t+zSB+C4kSsa6GItEs26j/1RGvtvS3/JEkr5KQW0vIDgL1cdwCcG
Ktn9POGJPnCfGcfhGUfK7bBS4pc3B95W42BQh0SNp3SzGwWY7owjG+5PFXZKl4tVDKgae82qnTiq
pgVUDlqajOGsqWUkIy2M1mxmPP60nMLILlo/FgajNYOQT6fUli0+mxXuEX+hI3MjGCwSjpESNhV/
I6Vx1/LNBG6Yxrj8GnnCRnqFET9UaOs6GwEpiCAqioYePm4VQMrZw4ocnuYEgyF/gtX6wc6y2MfH
0TLVowf1YBzstEcyu5HnH81lMrv+QTskXUpXKIYVIcDHA0+egTvk2CI3YFTY0mVYTyXkvCnv4aLb
5Hd+8fFT4h6Y3IkzYN4DqTh7OR55bEZgoshYnNumDFDh+MYGH+1vbufhFP2PdIcMgrXk+tJYAFih
7+UlHvhrWdJOQIUjm1a74S+63QNUwbOUfOEfMAKH9sGV6ft7G4SGvMZz66cPMxvQZk2ctJluImC6
VLJ3fkVdUc/1akfLzyDPuVOJDvt5x0ucLT8NfURXkMozIxXnIign3fzndLShEpI9pAU2QUFGggf4
WkqZTzwstKZHk3SjClNcwJYZKh1+VRdjOjpAUolVpJOLkmlOK2+WuXqq1CHCvLOybeke5ce/ckI7
RDIzIc4omfeDmBXu9iLZrThaK7ySQs0THaBFimXrEInz0YH8uIvGYxEwXU0y4DUiZekb9BkILU8I
O+IITKkwAq71GEe2wjc5bQKHiUvW3SEX54KKV7Ha2Ahiq3T77Pf5USr6ZGINH3e3G9uv8N7bWtrN
/QqfEaTloimlnZ0XTzlr5E5ZL7JPZllJIYkjILxwSQza3dpRDNsVBJaBUVl85AdWRlXX6xq+G9bc
X5NYqty4CSGu43jL/N9jQ/S/hWnGur3Yd//Fo9tSQCER4wpsRYOVtUzAdmfwKhGuvPHn+qgrozv8
8YtQ1nknBghc+31NN1rXqKATvw8eqgdwKihd0THr8VR/Vjx4WFAtGbe3bKSzjnzdXNUrJbpGy/ax
BGh9Sxhl9/RNqjWR8cCATPR+BYuNgaM8EUSKyT1Vnmtw4LwniXdQqMBZlGasUCBRmoFI1HI6+WyH
UKbXuirKex8XQl1Cnki4Xd6FRZhvjTZwWkoyeCqk4Ds150Lcxge/1+UrPuWGPt8eolZMwwVD2Pv2
NmMwfobB3t0s+wOYqB5qDpdQbtCYqd3zlv4IVramfrqLc3L23qSH1eU23DVHHPnVY52IdCQRwt4D
W8TXIlEdmRbZwov53UGa+KgJl0EfFbkx/veCf2YReSiqGWMAFyguT5YVfpgzGz2xbhmZTKIWhScz
8cHtLtR4bG35VAY8dJCBtwe+9HqxcDxMW9wGhFmERqlIKZBmVNiglG5z3akF0ytoYdvhVUY6FI9O
k9TqRQ3K0uICAotofXSMnEKmB8Z0DgP1UDpm7SHT3t/3jHHOAQqrN+9/lbB4yxGoPxkV1HKjVYI8
FqaQJzJqFhqhERxhu/aaRtI4b575r1Oj8XTWleBnO6my6l8Wi0y8fg34Yz43cGUZvMPFziwIEH/t
CqxQrSroMcYeh/WkGtkN/VooiQ3DSKhf9BReYsv1+U+gmRyTXyIcthtGW8iJB3fQ/1njDDWFWm0M
VqvyZHZ4k6vTDw8ittVuvC6MowdNrcsHX+dz+XMQK6ePO84ZUFrhK2G8OCYZ2VTm3F8h1P6dhMp9
lGFFPw/NBcv4ejDb4Lo5T3HkjmZOj6gbppikBEZ8mHoEu8TX82v1UZcccRa92Z/rjwDpfbeJDL+U
/x9DFDrhu86L4XQ23XVaIfc1ozAsdQ+GUV+kZAVlGelSy1gm0XYKecFG3r/MR2X5DNtLpiJJrSzn
0b7jHD9ZrAOjLk1S8H2/8qsKw+Sab0MmzZYBMPwAVl6pMPsSLXvr057tynP3oOXevKYROqX09OwC
ZfcBdl2WXXX9TsLk9x4tHDo9c/Fgsc0ouZlSIo9jN9vtA0EUJqqS7udiR/AMFi2sLUL8TNsm4dvO
es89SjonL351ZTSt8MzjYGdYMv0jK2IdMDYX4OsCFweI2Uuypr+asbjLSknCkqrCv9hZct7n0wEN
HYQT2+eTzLGNXQyoczs8Y65IDMNUyJrh4umgnq1caGYzER7uDoOW88L1IxBQ1aY5I5y857VFgJt9
hU5JPpqJJbE1z0ByNJZzzRIAr3DKfB0uicjmrk6hewxnSfMK+1mCC3qXr6+RJI1EL7Z4TuxzYULi
T9CS/G9Nw6DJ0DAjrsXDxzyUZvXL8DqtGvhekQ3vikHEUEpZkWRmS/n9vlG61BoBTbJ7aiMmTfXW
WS+epSdaZA8XafiBvBefXpc9feWean/2dA0lf/c5AiSRHWRL2vPwMv0oc4CpIr2IXuovUkU2Xzad
ZhELGDjCLB2sN3mBxx4RUXT672DdiDa/D3LL0VmDVBntXkpB7BCJRgsotF/K760UlV8SaqZtUsiR
laRHsVDvl/W4UTVqzOiKAqd2vXAmPXQ2317Jm8hN1OJPDtfYb0ZPWqTVVOVFJbt4yK4sDaSEzO3K
AactW/DEPqsF3p2u+MNztwVbpVuAAJ2H40ADIGhDSplQUk+e95jl02r3AB6PYtMumwNKXHS0Ylzd
uojXxpyL/H7QD5WkzDeepYEzzCKnhw/y4b+BTiE43VGgyXhu2fnlMbAClTi5FjMGLrppwVFxUfwm
DxBZ1xOcN+ztpHS9SaDmO+jkAbmhcYezbbXYqhU1W2f8YuaG492Rst1MIH/sqwdSrnmAX1dfOV/V
olOgZPxkQe4jC0GU+T0kRti80PJuuxh7+2gSCPeVbQNdOHmAqZx5kP1zpf/UKfe/6BbSDyNIj1PA
9qQGZuykY2zea70NaUELplasgox/zW6MUxUIF3uIEmF1KALburKgQv7r+3lM0iiLLa0SNatCgTQ2
773yrzcaIZ680P+uy6Cp92XlK7vh+9HiUrRf6Dm7W4nlMFy2W0UhDYD56Mm7bZMgJUypGTQRiG6n
fDawhoRPSBF99fOuJs5wRQSDt+/Zn9vSIuuNaOWsb4sT+53d6NRZDKve2oGo3Y0oeEJHGLFtDg9O
3aN5h9y6XAeR5bmz8ivSYIR3NQvqQ6ts8JI0sNFMfDT+eiWT0KLL3tW29sGAI+yZ6dO5nPmTHs0S
v8uKuf9GPxes4rxawlHYrAfavROoqSjckmgu8zZeSWtAl0EZeQiqNAK+SHJxnLe/kr+TxtfIXB4X
k5WpaEbNbwjcfnLFp9Epp8wIzdM8OihzZ8biirNyMunxCDyvz65zf8igCkHujoYEj+czjo7LQlbA
tfhUdNu+UghrMa2wbN5tFXlbTjcbc8shSz0ICNKFH6coTHP4CYF/yI+VceqjPph2ihOToYGoKPOB
TcEafGlZhC08sXXg7uZ1gnHMS9OpM8D86E1nStzPbQFCpuYsuH/QXLs/Eleqs/J1e1JeYTbd0ado
wtUhJ31QCsXGZUiTt3TRuG555fYb9LcVptWMGBqoTROjewcbzIcX3xB6qCOn/qIFq5nyfAOnjFfI
1htEbTGSTAlXQLCIuLKYo7n4m80ITdgChVQUmMVvAUSbW3phLx/zzrWd+1CnI39scbU4chDJQpQJ
+rrHANYzp0GO4qom1tx3mVEBqzO1L7WdCi5FKjSeU4kILfuBKkgcKpJ1UNVSVFQTWqj7BGou2Rcs
MAQUvOzfgKFMNuq48uAZ7dNIR+oEJhbn3gJkzifl/r31dm+gwESVbHJc2PvTav16pz+2hf2NlR6i
TEbUSX30TMCBljdsWNoJ5D8g7WfupRv4APh+nPcnNLNTwh65enGV+QBZJSGU7qoVRhQrPo61xbbS
QulkLLLhhrXtjCcMBzP9H48vog971a2Q3TJHMviOEOQk4uxRvGrtdpzY3a48yqQFqoePLtud0XIG
0LHRnw6EN75Zqq7iylt3ObhDVZcvLaSVZ/yj61ZI4hFt9oK7rhxZPxC/oIIVn0rEU2P8Gt7D8HZV
kC6zA6MZEn4bXpqLkwKcuouPMNCwu3dXtVkf+cmxp/l1QxsPU/lz/hIWVJ0UE54wuM/k2TKTk+Tw
AwLQyzEAxurcs9jtSqSJVSB6LZcEgW+yHJsE0Qohoqj+24CUnPkCycrVle8AJiH1X5c0/CAibeWK
T1BsJESnatGJQ01AS0c1zD3/aJgO0JK72CreZT+VX2XtdbzxIQ6xYYxrz/FZI97gCzD2Bs3XiUNM
Sb3Uo64DtWoT87L95/pFeoQ/IBnoJNl5Ob3zVfX5K7nAZcAUg8N2vkeMcM1qO4diDLRef7S0gITI
DKMZBscLGKYlTuKTb83QNXB1SLqqfzJsGYxuXrr4rvKmR3nQj4+yuoRVFAl+bkOQmppYfCwnxl+Q
FzYQw4elh3iSSB3x/cmPHWzqmaM3mV9KcemtQmxUkpGLoc9hXrdvbOqqIpCZRSqj0N1Wb6jgd4K5
lAeP8AGD/q2gSEnnZwVYkcVOGrheGrjtvyGhugaRGO/HH3vnE8Vtja633bC1hj6BPo5DmqTBOYk8
yxMC3DnhDo2G8+yd/XjmjWT60w5sb7WQBMwkFJBSypMy53vdzr0teR4vAWdfK5hnhknBQ0qS2DZ5
vEqLDrW73QH421McbZ/DbCqFhVaeFE1EHzW1+V4CvE8IkgTnFsb7Z2WPcWs3vgCME0ldcSFksqTR
FIQ6/pgSSd67omjbEIAwnV4imMzOy/aXuy63Tt3+6hXfk1qR2e93vLHsV5IuusuxwvvuQ16AtxNx
FQh5ZWG8s0it5hPKi9R+FWRxgjp/HUQwNUi/NA1RuQ7QoO1dGfCc/5AP/va+nVjyqWvMpxqjbioa
UOynrXxgXBQmxxN0+Q8ktWriNRRLd99WUD8dflrJGSxdPOeeNI6OONyRvfyam5DHWc2afR3Rjyru
sNritV+ehQSdjFW5cG15vL2+nADGbwD83Da86gaYDbjbT/e3wMzwJ21+TrAugd1ytcuu8JJ2isnu
h4dDBto/NZoITUCNnRa0WtWfHeeF6XtNL0mQ5ZUd6gqxkHHuR4mYcW07W55KKu+rM0TYPXKYxaW0
/Yti1YXvFnJAsSV7hswDtcUbGyIIZKh0oQKGls5rslYp/z4lwIEbKramH4BvigVmey4IcVYAGhoL
qANRCFp8jBncGlO5jxQ8lufIsrrR2+s9/640PRSLAAk6e438q5BYYsLaTrqNx348JBc0nYAzJ6JM
XQ3i8Io/GKZDj00owUnRSGukM7xInq9WRo1lEITnbk1DVe7ieaOCzAqKfm5GtHjLiscFobaBX22f
VX39iFSEGftUdT3p6AC+D4JbJEhUSadG1rHKNXeGiDLjC+oleDB+cyFT9FB5UGAYcayQeIYDLtXe
YxAgQqPiLN2AnDw6OA09yRMjpR5RxQFt6TDXk+c7WyCb0TGlvYgQcROb/1GSTdjqEKDjD/BOJ/Ak
SLNuAiEPzzp+NCtfKIrI4bJeRiYbwj7CCY/qVh4MExhjT8pMwhoFbwE0CRJOs0PXoj2fB+cviHfM
hMMLJzC63KBhcBu98ZsCxNDWx8tplf+SVYhZ/Lmwe5WRgvRTzqU7EbYEONGN9W0PmOKkXxasXuyr
AP2SaLO7ytDB+pUJZA7EoJ0rlUoX/MfVmjL+nPi5OzscUy7un1Cvx6irrIDRcSJZQYWcMB2umMMO
iSCxVmNHq910QsKaLD4B3LyjDsWkZoRT2dfWFiWDPUntrwoe9RJnaCQXHQ2hSx595HfNP4BY7gSm
Q/wRNBVp/CTf4yzXjB6bDFtMa8q4wzth2+KGUSi2keqpJ/S8njxb9i07VlZPdaq9U1cLqlmefmin
ilj2fuyAjrZ3vLLlOEqOqFYAuCKH6//Q4B0+DIGd352vE7SYCzYNXodlHjFxmIl/i+ANH4JoUddw
d4Sqwm9pLwLlIY0XeRWlI1PTGHyKnQ71XcVMtdXOHx2yq0WkvadpRSCsqJRXSUPw8WERqVkCaFK2
unt9Wnz0G/6h/wQLaGkOtjg1Q6cbtA0kJGBS66cFgz9Z2Ow95XIvN2NJ8HlRzor6a9lqkxYtIKOs
4C16a4LXIxSo1bnYiGqWtHmWA/d4GhYRlZi/CUlayRYlL0bA4bhGOHHmhajZgKKEwYPJeZQnk+Mk
LQSnKHZ2sMV6wkwwj0C2VGpf/TThDQQtixidyFQG+MhuDGYgyqZY2MfNygdyZvT4k2+Fjqxnf1Bv
5eGcNHe7MYxwJ3zMkSgiSUyiQnbO7mSkMHkoayepQw2XMVv8xoCyiO2OgoT0pDLgTo5QmWTjT6LM
T9kEMu8xBPdgWeH6GC0sLwLB2tb6EM482R+RHzQgxzxCM/vCHmcuG7LSpswpzZAJNiFs7DEy1Qq5
0sP/bCgjxAg7z0K9meAjtPrmw9W00T/Yqi2OPxVvklSR366suKs25e1RHHaoKM8QIvukosA1JRsO
reegbhK1jk/y9zVmQsq/KOIeqkueVEJZbxRbhk8X8GyE34e05sFvBTEAfd7rTSZzRIPCFWwsC15Y
dJjadERj1z7yr+RrqYZ/gjlxx7hB7Da5rmc5AjkKdQcXH5gA0EMtY6ddv3waC1lx9xZe4sg73oAc
Aso1om5oIAFs4rw7096mB3XkktOspr/1KOyQ3zyb257dOlKNfFSDIFs/PEO/s/Gyhg5KvSicXSjZ
rwEElkViSxj5Emh0T8f1n3lPJqQYmgP+gZPsLmRGFTI3JkRzgEn25B0Bzg0r4RZKmeJ4Kjw0P/CF
1nBt30a4qCWwJ3XRMxHFK0C70K41SO4V5wEwjb48PYmo9LecMNTKqs3QfRfmpOy78ZWMy+jczQI1
QmJrISZhB2DcwqiY1n3Zl4RnBWn7XcvBR6EqvdWv6Kq8xAKhW7Dqfn4o6/hyMoSdrS4wkG+6Fs5v
ogf84smQH+D+r9Zg2RZImbGKs5JkFJODxnX+ZFm7JVG3bGrfSr9eLeSgET+YudVO7w4nUNRlMcaB
3Zu+CBl+p4dBrGddvSR/yXMxsST9ax9RDKLp2HqZRTLiOXw95SmNQzhGhD0ub1qGjnbtT5rgs8kf
EB8fiXrNq6NVt9cxxef8HMM4cCsPy5spTjsYal7AFAQy9ctEv2ZDvIpy5qvr2Y7CqZEgbnUivzod
zIM5QNvyW/XvGqxSLb+y8osdeHe+sTmQZTNOED67/Bsb6juE6ihXO97riBywsYB8CELhVacIQOV7
qIt8Uy4JS8/pR6HmIAqxP2GAPGaNpaA62+0tUu3sjlI2cnnbCUvhU4ALpquudgFKZPIOb+f80rD+
TbvEN827l6PfOe/1P+PJ6BdDFypu5jJM4itH1Lf0RHBXQJjNIjdWD4/XneWIO6CX/0q34Eoyk5RJ
9jM3A3Hb8zp4P+FKJYV6Y8bd/OsR++Dd3hBb9lSmv/PEhbLcY+29mFYw2rCZKtGGJ2RmzGgqI9B7
zZOC6luDX0K0qHAxHASYFDTRRQSZo5vdcybCyXP/wqG0YriHnjKMNkH+0fl5gZbzMg/AgSjjeBYH
qLVjJwOQOTXSN+ahvsF8R8Wj+OO4fpBf/6IcuoVwBlLWWJUJYpgtI+YLKD5/jx4Y01cIlzWSvZ7E
smOCKIm7I2+riXTrqCESs22r0xTSrfrQaNhQwj8mrq5raWTqP1ZB0tKrr0pYXQmZjKpA6lWEJfdL
1KEpQouUwtuu+iT1KXumjRV2NicObXBSg8M7GdD6HYn5i+rKICJQVDvajHx5Xa8kgOfJW78FDvko
Jp8oCh5yDzWWO2v75pEUyXHBOfKHfzr4U9BV6OwnIFGf0heZdrawasvW2oN/RTIbz6jXo+NFOUp+
38ENSW//g/y46Py/OYMbsdMQMY8iY9ebIyH8XzY6JlCEcUIIW+kw9UTDfWIvuz75MElzTOoqTR5/
QNT2Yhv9/qSPb5Z4PYb4o14+U54tnILOdPhtX8hDeftAvSHsThROK8VJtgEaFS1n9cMojKJjEiDb
13WyWb10vY5zFqTwdfRwCC4QoyaJJU//pA6bS8ginUgJjPMoUAs9h9b0IpS/89ONdgWGICVu9A7m
45wIqX9uAsdIOxf+nhyK5ryJw76Yzccu5oPHvtcbqaZdJNUI3/BRu55KIKSECAto+sr8SB7DhzPt
+V7N7RoHLmweT1Z5XE6D5EAYOnhtLpVO8QIV3Zwf7G6qT1iSYtvvF3AU84Fg8ZBIl7v1EMImX7ok
O7gSlgvtmGgpDgj7xwsGP+GHHrTXG+CO2ZMwoDqxIx1GJkMvH5mUhO7Wjm/4lhyI2UqJHUhoscwH
D1HFFG5uDilFv7iH7qhDQfj6mOoECK0vYtb2XtWO5IB6vVoxox6Mi/Q6rFnbykaUuhoCNKF8u58m
ufRG3CY4CsYWkXAKamOXyqZk7VbYyHPk7eQqyB08+PjAwvIINm107WHgw2YjTNsEFd8ZqXLX+zN1
IXFSIB6TVDVX9rhXGRaOmLfH8mt5SjKykJyvZkEwVm3yBOCuUp1ZM6HXqj1JS+IHZ5eQqJTQSnox
QqvKr9J22YaqQq77dQP0F6lsj4wx7jtQ1eFPvIh6TLlLuPHDIRdzDwQVA2v6ToOSTZQ56s0O/DbC
wadqvkZx+OSbM0oWyBpDf+76rMSP7HacuiDVakYlJX4P/4qeuLvufSYX3sJar2h8KtGxBNcwo5Ws
kwCxPBKaj3OH164A+JJOBO8/HODrUGzR0LdQoWRSV+/EoLk0azc+MislBFW32tje+F50mLSPkqVm
KishFg/wOzjDihrd58nejGV7vMdtUU+/3zCnU4cthqDEIllprzHboUaZiBUAYCpGwasgz144YWp5
1BOs5yALqMEdEq/c7wna2DotnDkAdy/U76sQZgn0ldJq/IH15krXzgeW47hiq1A+3urw0IjrjmXh
MRucPejHW1ZoVDT0IXhw0C7lDnfhHWyWinO4sqs6UZPg/teMpwPDtajtg+fJ0FRoD7mApKTuHMCv
10jMaP+q+23i4AUtevgC2ZO7FsQNJA8beYADPWwOsodhPy3jwKZnqwM05CAfl4qGg/TgqjafDkju
ZitdbIsh9TsLjPbhgnzR9L8JHcc+ttQnVgzLwDEezRRQ2WXWaFk7j7Qsl+LG6nzL3hacTywhL8aN
z456xCCW6vgmv5x++Ov0WJzOResTvBANFjZnCi8yOhsVE7bCU0imG7k1KeLEULYLhUlr8k5+2oii
etVQkQFDkk1t1A7quOIXmz3haVajG9/blWsE9FjTlv2uPIG7llDWu+IMizBVpI4ijki4kJdnX5dp
BwF/WsZP71uEJNzMOAg9qV1tvbw06+4lq4qpDCgvUxLiq++dYOyQIkkv2KhBDSpLS1EN9GHJ2rI0
NCrzhTK9yoFFmdvSr/752hRkbXJAI9oruz4mv14VpdSAvu7BY9NbUxpjfsIxA4rrl4DBhRdGR7dM
1z1Xy8hxaBo6w5gsuUxx6DCcw50bkVqUSzaXJB3FDczeW18bxKwWe476PrMbjnxZJb40coJBvqyp
6GDHv2myqNLQGiMJjAK+VIi0TFqLXeuTDr38mKfsDdglXdsIUZ6LoWk3YNA6K1QArT/biq9tLfyK
mRzOXPqnLJsoQ3WBeeGEJL/WxozgB0Nd+95p/6E3A5bejxStnaFukX3t0YBTCaVQuTbxDe/Iyn/k
5FG+aFeAsH6MPxahHCdyAyZ84n8UedCqclnuAbik4dvSOjlk1HYT1EsmEqjFH1zj32+f8mVX2nku
AOigu632LSP5UmA8Tqglo+Sx/Z6q1KNS1B5umkDo/jlo2N/bLV3gzrWcq5TOOxStuQMnUJWm3mE7
m8t7YGfbs118qGCUhFZ8kJs+uWj6b4PEAL6k4m5bsQOxHnkdujo0+2QO1oQnIoHXnfvQz1sHd6qD
yPF9SSMQIP2I8qJI7yEKpztNGGasmgOh+CcfmDEC69CSHVFAlGGmcWv80vvNcZhrVhmEPIEexXTL
T4/Uge7AbJYJfI+++NtH8o3VlIo3Nsw3RHwoIOD2OxHI+SD003vA7tKLI7w6EjwHKY4eEajhQhdi
3EYvkW0S0cP9okqTUL+tU6shky+Ask/nPoyOjHDP7tFYqGxZmauwHsQzWLWNTLA8sMSI8c+dx03i
CV+9gqNCwm9DydVmTgiQ2m+c4IceTbfvCz67q7NUjiRvWLCVIWO9Gd2nPU5r0zN/Yy36+4ruLoeI
tUI4JRIizYuVzJS8G4B3TzZ0l8H6VCc/B6tzqRRhMgM7rqle53OFsHVRLTRu7lgCnA+NyAAtOeFw
chYUi710VOcssxYKtNPcHoyzAJTmX0LzZOLkjomaRnyFgOlsM/982q3RKDpq6bZ4sPJSUAOgWcMT
0nsXUbRdbgiaDwHXKYJoKERk3zK9Welt2d6I7NugxPHOTanlKOsrjFyrcajL0UL9IoJTZJY1C1n4
WqmApqM5R7eDv9syXOcFDIYNjYYho8E4NCSrzi7XAAU9+Kv8DTAZqyTSiuYdt/31T9Q/ucGHv826
UBDl35FZasQwZkM1Ad7O+T7BEL3iGv2uFtQWpBwTbMKEKXQj7FNzBrxMiqNVFEifQfn0l/By2l90
Y4FmWlng7TgczZB7uOFKyZTCp/JQv72GtvewHb36tbDqIoFmUClNtKk0Mc09opAB36w6CAA7nmKL
NVSo4KkmcIwZNV+Klv4a/zbVnrgItscLv1KlfEpAy4KSncdVdCPHKEL3QbKkZKBiZaxCdOhESZwm
epvfweYz3yYA2N2fXtkEqsSR9MbfWFmJf8FKHtiboXROJgGYt60aDGbIx+ICfzFQTVdKUVOnAuqr
Ga/Ze5Zd/UE709Wzyue63zEaLWboBNWvgV344jCTevZm+y/IDgS+jkWB1NTrlJgygrYZ9jytyV1u
dsxE8KX7SjEVIaExqgxzc5J4kSqd2yMiuNSTd970uMS6Fxe8FP/5Yd43H4XCtc5mLxpKQen3JTGM
KYYygVPNCnkRZuQH4r6u20lhzqLx/jaEglboJTFXSsSGRDXcJPNEJj++6dFn+lDIqQO+KLGSp1cW
gAcfh6KRcKQfnBk91YgfZzNuMUZsR34S3vhmzgCZLcEAqN61ebg7WPN8Hm1iyb5haOwVwTlNX83X
d8rv8B3yoom4EVlvKb//Rvcjovd5+xdUEBIkX6Sm64P0zbqLt/yP59NS1lEagX4RqSfpWbrR5RnP
TZuDxZ7nPWUboUkiF3H/BIGn7l8uKdb2hszZg6510WHbyH66tP1/Tx/ViJ04purlDTJQpsAQhnua
uYSVAufe/vVxeXKvyXiO4UHujPQoobGXMj//VygpO5xhrpZpVzakFwwmPahdJN0JF6h4FK/CztxU
R4u0KtGXTNcsrk2zoJGWj6QYxHUqHjj5x8D8iI/1QfmanFFl/q+r3TB49jXdG5mtDZGhIipfLIDs
NAKKFctTvP9yUlw2IiN3pfWZ08Y62fuDPLX6pRFxX9t1XjPU/6fh6OcbA9o9qfn43I+nbcYnnSeR
6l0HS7xe6JtLoHKFzZMwbcFOYSkZKL9HwH2fl9wpOBoQazIfEofN9bAeW/Pits3QC8Fg2oLYe/WY
vqyCt/5ea21qnb4ND1lQz3Qh+BnGljxIblRfPVYP/9rAOizx6fnKXuPdwWcEgoPvFYHwsZYWNrFm
5O49JMB/y8ZC5mp/YLLR+UMRQDGF8MJZxoR61lOm/mdy6AJg7vqhmhMlRTFElCxOTv9avPvE/UjP
YhzexRpbiQrRagCB5e142e7HcmX5im7l/dJJwmpn8S4GZKFSCbIPu92d5bWJoHYedkb89XCOhJ0T
I9TJQRKSLeKMKCAEma/DB4acH3zP+jogPisltRIvmISeuBAyHQL1EQ2EU01ACBYCeMbwAPCeRT6d
3PFMiOAUBL2+aOd9O1mwj/0eCd4xH92BcAvlji8TU8zffHBexE8pu7B+i0eBHi/8W31a7wN7uLsF
jlASTZgWJ6WQQ2JM83d5Y0lB0+vdlcsQ8Q2ntWbqaOBjs9Rx+bUumfcUOqvloYt4m/zpXSXv02y2
y5/gzzrm0huDjR31yn1V90TPpD4mIrOjgz7FVWtaQpFkozYkWWwRM5pgPiN8TIeGqnBfBYaVcdEG
2/n+3e4A8buw+oM1AKq3qltV74UzBKyDZI2v+6eJ86YMrguTza4OV9AQfKqQoy+2nZlR1fzadX52
D11DRsyIuxFZ1LT5cPfPygZagG1imeMVucNgGlRNY5h47iSSVorg/3jZae65WfKKqtS3GxV0VFzE
7rR8wDFyVPS30sGySd4+kKCW8LRlMgode6RVTWj5UiWEn6GCWY14pUO5ebo2RiBaNCteW95Koc9E
eKEtJlPXX7Sc+W48xUJgi3sw8Z5135vfiy2Fm4wBwircpvNZUYQld5lERK90Z7Ed54ATiogRpByy
Y7wVxC+BAZc++gbIrn5ptPqLtF6fF8GuPUBhG2ru7eVPoTnTluRP67EU0TEFSHizAjiWQH/5fqsu
zR1ZesTfCDkVFJZpKsCV8T0yiXlHGpQI5RJKkY72OQ4L6KZWzxmuDLtJ8bMVixZmb1ou00/C/jao
sxxL+A6Q8CDw2BwMbp+CcoSLTlqVTDj12jV4f/6Gf12rMR5L1dvLbxa+gbYrb9obuXbrqaLXTzH0
kYbPH89csD6wEnkTX1Z7xtJvyiwgStGzJCJsWYrOzf5CExYKs6ARBKJz8G5QOJ6Mvua9DAA90GUa
ezych6EBQ9DtKsAFGi6APPP8Bm91uQ7d4zWA03NZDeSj7i74dbpNeYBGMQURsPcRMnjf+f6DAVOa
Vmh4198lfDaWKnZTXAIXGYKZVZDMBOjzLQTq3BiTCzCoq5Jie/sdcYPWuJ+JO/X/cHNRHnkwwI3t
OgNR/uTNrw+HQUVMFraiv69FdMp04un0RLH1o/qsVkgRfLaUDHPqZPJjWtwEhGyXh00Vb0vktzv2
sAhwmPB+L4+q7Zng8HqYspme6Yb98XZad+nr9sGlCB3Wn4iRjz0HrdFCf/F+NCiwPfom85miknVB
kdYxpnBmDu39aLHgPP2zz/tf6O+VP60tUGRuIgBrkN3dfNULoRqFuI1KPKL6yHrt6ms2Hp3vS8Er
7RjJFNItS094rPCnlDf/5tPz9pQqWdx9u06Pqv+KXV24B9nJwGtyZQ7HH6Yeo18yLm6dYNcd0CAC
EfvKqJHtp8QjT+p+C8gqHzYnVbWwKYPPfdUc6E/7ohut0ThuaSU1hxXgxlS5HnE7N/AlBgvKZooD
BmNqxiNhuC3LyEQvRUmjralVbA5xUts1GLuMAqd0BDadYJHXswtTZqY/P5I1oLkESZL7qdoHdnnq
TcRFh+kfgJOaOc5mKlyeATRISd2XRr3vEd5PNTswyu1bNclArfZtIQmThu6f2hxgzHeiPyZ+F0ic
ftosvIwPX+cg0w0RLSXIfGhJyVUlUxcJcChxlShr8fc0jN6+1jtwZhfLABAZ0n10fHee8Nh/HQks
VAlVMWolXONMRn7k/B5EQdLSTCA7LhzIB2UXrHrli3ZbTlW9O+7I6SUpPnjsE8eXOevYmBTNqIAA
tTmHcmkZVMW/p29xP/CL0WEziMLisKKz/LYGY7Db5sxDS2VoEEUjPAH8RlM3VF8DTRzLXAgYDWOW
n+Z4MOfdqEdoLQ6pTI24pv+0tBjpk8za6LFftRRsV+hRq4/9Ls4bZ/ISjn64EIuHdq8JxFXPdfbH
Gu9gljX2nCK9pOfC4E7MkdO0C+iByvdangfNeKG2CZPOeWVFk1+rjE/dbshj5f/fMTXTj9LckImL
k/Z0eSF8fIbxjlBhZdiNRssED3Mj76Or5TS/bvfAD/+Ngu7i3Jyo3cEFfDu9CKHgPA8QLDTC1mWd
+3/MlDMSEbrE9H/1PU6QhfAmaN3yEwQrXlg2RaktCbGslmIqFaVJy9qi/TA48OssGSeCDoYaITzv
mEVe+lls8Luum75Sz7oiMjZQ9Hm83jddIPyOAWxS7EQqO/vfcVgLMxEaQo88zdrXPC0U+wy+koSm
vr/mwvPQ7aB+bxne6FvXgbq20wVl/CWYJuV1Psk/IhjGWrBpws2GU1l4a3mZBJiWiAivVfv2npCd
q5k67bsQwmEHgSzx5XOSwsq6b1ZscI/BVhXPFWGOemKMWthEnXNkIbPCFJG4BsRoY7Y1oets1Mdk
HaVhHQ/NbtTOOJwDJWQ0dB3BmBGf/c4z4JDMphwwbisWBp3D629/PfBf+atQtwXygcnno3zciI1X
aJg83np1kp1AtfcDG9jcbT5V+oTYHqq1MI1Iir4AmJ1XKGfmptaIaDvmi1EHsmmYyBWZb1lUwDp1
+vrk6LX1qHnaL7ZNdmD/wKK7W6iheLCF9ZxqUp0ttItMKf0bz1jn8wBgkArwrR4Vk28ZSwWiqM84
wOOsbN/zxdAOTOKh/gk5TBL3Ue7DgaQJ9FjG9te0qM9d+Kj1cnJLvGWv4h8Y63+w+q1Q1ZLSg09M
6gqLoj3SljHLxyC9WHm69W/AMscNtUcLSLRkQ1Ungw1XS/jYRru68sV/PyC+yvlRMa7zAinLWC+O
FJuRpMmdah+m5TF2MxPbDmyv505y7Qtf53P0KT7EcDcNXDEELHJ0Hfc7T3oTKH6DRc/AmEgT1Hyc
ZXmuGzGnfH0EQEJxM7ohKcn+7RmXRJyrYFskuirZdEuhhM67bMI+352BDkM5x7zQL974saMtZUju
/I2XwBTPI96B/JBbXymE5cUdWN/jb8Bi8mu/3m/y9+nouEggqcGDHt3z0HWW/v1lRPJ+tPOyP3cy
XQMkeHPGVJaOKwtS6uELJi91I6R23Py9ZTTa3y3LVw2uQXExW7yucUpenqvcme7XseTaAzMyEmTk
nmpXmF73MB1fV8S9VB3OAd/yw3FRZJ0IUYqo5qnDjbpY9BS0kha5ItQFsfQTlnX9H88TZZolHmBM
BgQuzZMKWCoq9WdReJdIKfJPkGjCeaAkz6u6xSr6yJqonPQHHZ3cqBB2YiXwJj1ZWIJ8AgVX0Jx9
h1PnnNIQxvvFpM4ZL/3zPgdjlFkDV8rakELnJmJvTm316WdnxJEryvMF3IR9xrp87emSOPNrSdSc
dfb0djNACveGAmA0q0UdiHqp5j7KmRxXxTRA0k+9JkdJfupeZI+I3YtVVxgExk/jQn8QB3TzEPsy
zO96VAqITdXaljmbmBKsXT20a30F+3a1tczR3yXky2cUK0YeOIBu8hlbPVFO6NAVAxfvqfqa3dbn
yEGXR1A+0CmsvX0xlaVyoyEvCef1Y2EcxIZQg1N2+0OJoHhcXhVA073X330mfv/ULAOWAsEpr6ZZ
45caKBTQXFczVoa2einH5O5GSv5qGiN1DEpLcPvaZ5aWiJQjBRxWvIfd5e+u4KNTY0w9p4QIzBns
cCazU8oaBZd+b3ysJS3wb/sOkBfn+7ZoAoxjuXZxK1WOjTr42bzrx0mGKhSqSbTlv9pISYGQfUIo
mjpxdd0keclrUkhoim8GHlxKV2Vgvk7WzHUlMiCkxvzrhJx7qQrp1w0g4H5e8Eew/jYtlZoIU7JH
v+XMx0sFeW0lHuvaTiEoZNT+Ed8nLGOFPHPH0lXyTRLa69eAsRlExLZ+3Am8XJ145AK6XS+BOQWF
eZsEjA52fpLuhWVJS3RutkZfHZ4jVh1DZfWtQWObbZvKas8iBwA4oBUZCOsr5EfUxXYilDELBdof
/nM/EdHp45HBAk4N3PU8CgO0r8j6K1oJwi4vp2JaPtPmWBbOpgvg8pv2Y9zD2siWRFMxOcHM0QfO
ftY7TRK27yxhu8lDxo1XiSK9ozQAPk9j8g/I8LVjKQadFL4y98LsB8m+jX/CBpmYP3dekIZo4eag
ErD+Ky1uiiowA0qon56J0SUoVj3yX1FTEjO5s6ZDZFHS9W0RX5qCfay7McnDhketUO4TvOpKTOK1
TAf+VUb2JSgWLHWJvxi+2Dqs8w+fm7Kt4LfHtQJkVv3J4gC1AoZXOJriLQDdBF0HJypeUCR2WoYW
kBWJ0eVNbd6s8XibJ+3Rw/YEHtOXJ9Sp6vfPQPkG5/CikxUud8L11GJ6IK5uLKcUzol51ddgF89e
rPgFs+E/03VJ+xUgRFbBbqKz6uuyaJZXDA/o7f+Tgn8brEKTtFCG75ZzA2qzOxFDqrBkWsVV+35Y
+s4b7cV6s9bCCwo5q7urPOhm7X0jL3deMsOYwA8sjbN29DIlSRgocCyqgDUXBlzGYYi1afoCF6Wb
HweP/yfcK18eXmXuJOIeJtxLC0VR1gp5BkPC3bErcwbIqzLYU2vse4AV6UtopHRp/tnoXDDrlBDL
9AK5ZRPA3yP8ufA8vofm5Cb43MHn/zrha1GWcSecZ8uKyvK8TYxR629KcfTjUSbuwlWuUkycTFLt
TtJMrL0CMSB3PzN514NDrGPxN9ryOzQI550l+DjxXPN6pn5WqGp2PpHZvHFSNxPb7RIzMwgXKKLJ
Q/NywQk8aIlkshGvnql7Xem5fULZSlU6AcQIReDq6NDklfvD2tsE73w1HymwqV1BXKHmMUe54Ye+
NiLrCZUJKiy2Dr/ILz1JkoskZ0UxvruTXJRwL4fjgJef9/fy5W5Jysf6ukY8IOvIu1rDiEUqTD7P
/GEQeyztGbeJP+4UGaT5lmexrZUFEtCH4ErsissL1YUGBSz3LrnRBXNClQMaQhWFwdqrtRUvVx9m
G375XfdMnpkZ2QqrbwTEthvL6+Oxu9e1yqhiPH1cLd/JHchvHYQDacbAXX2VH+FOrVQu3BHi0VPG
jBCWMqwZRvnl/aktuvI182jq8iGbvi1VyGFQJbCwbIPlySpi4wULbiV056zZzzXQ4IZsXxWT44SF
P+T0EcLghtdzndcieukVWHVFpAKm0B+EbGJirrk65Kto9kAXXn6zc9rFaK4USHjl+e92YS9kk5lT
L/I5cBSo+u+RDANtpqtAs9shZwg0EC/ohqUsjUrHPLR7GZODRZ9LJ74fX5CivW28yhn72x5l+9ty
H72U4wZQrm+p0I+IAV8z5S8KZ6kHAZZkYINj1d9Zqzys5tx72FSIkP0RT0f7qgKUOLiLo/2Mfwc4
1wRYAdcO4mMIIbMfyXRfc+QETBHdNX5QfIZVG22/SLk/TPvYWrHWITFLa63AWdG3MrYlnl0IBI8/
EdtOgQ78iHKfLigsO3fo15y8P//qyyc39tdErp1/zyE7x0FfVJfg7rQNVqbrJYS33IN5UMDpjooC
aHFm/w0V9iQRUT4rN+FkNJk7K7u9XkdZU8nQ5/Hnc1fadWx7Iwwtf1IuIFKIFTaqgvqfj/1xHD1m
ffIrI5jGfFCM0hMPHa0H4ZFTE+VgE2Ank/vPDeId9yh6+i6qaJf+DbcqWyOFQY2uh8f0f8MJ3JtO
NeovxXXgC7FX6B0TXa4EcpAelWwdvskb+RQdZIEfnIzqlWgnIiHgPXCqqQRE+1TFvBfoLRbGQeDq
4rfSYYo4zyDeLuYyrFCBzac8faZ1bfD3q1WMsObPY9S54087nkwbU8FojvwCK+xMT+mq7S4ufy9e
59BKlyW81CVFbREASy1Cl8SwM0NMrAo/px0IQVSsbokqLennBynDmDBFg3/DCF723KvivulllXha
sQDpJ5Qy1FYfAv6T+WxNguWOJMwWP0th/gsehOToLsQ2U3brTt9JQ5dbofpiER65dQfj4u977h3b
lqMOoeWbUXgOhUWRLXCkREaOop7psDpzs6M6nwJAw4/7YfAx4XCgZAfoj6u2LC6yeLDsfaJGgoDB
IVyX+zqw3VrrI64tc4gShNYZaNNsR4mPpPykNOTY1uOr9lEcKYtldKILVsvLCd1vWUr+mO70+JqC
IKNZrMvg2CmNJrJwwAq89YtqedWbCB+tFxuJfp6cqPYEYYns4dlTg+QriVdqXUz5WXCAFruuvH9o
pJZmfQbf5R8TlAFx99OfezfLkHsUJbONZWTsX5qTYaA1SfqCVTO0IuXbZU96qP+3A93Sy6Bn/iHp
n+KGzwsOxMCNEvpwtyV1j2RYtc1/fJ0tb7HuBZi9ag3SPcYB4rznC1GYj8XQK8Xy1Z5sg7AXeKG9
1svXwEhGbujeLLw/a8EZ3xAExUHX9dsnhivLpSV2LFL5I6inwTs/UnDp0/tkxKWHkmX6y2GQl5I+
CcE2Ed6k8tx4ulffEFt2chVMmRQE+RjcSJME+XsRT0Ofqty9km/dSAbqvLkA434DIAhEcGkbpG2C
8B/1zWlP8QZ1a4wbsI9PjNcF/uPoaSHmM/tzyEhXbYnW6N2pW64TgsPTnlIpUm9N10hC+IbZ3eGN
bV2XIYEWWuirFyJwKVwf/J+tdMsvMtpI7XF8amYVFbCCfrK8uKFFpp5xGviZ9Db+beODZ/UWDsmV
2qg1CRhPj7noIwtwirftPRbTKDAYs2F1OK3z+3/iVZ8j5iMvs7awNNV11UYXRl7Bv2CO0FYWWgIz
758dLJzqjf9Bv8OHzuZpbhGY8BMHvblK/T05LrSs433we3hdbTF831KQIshOZiIUTJwmhyyH7Hlk
XaQb385kncS5YI97V+VUe/VgrJuJOJ+vqBmUudADOayNwEHhwq30dzgAO3zkiLtHBoiualtpZYOt
kfSyPrRFimKji2tA9on/ZOY2Zn1Yc38WTjN3Dln8QlpjzXb/kGB8CvQsCXSTRaakMNBP1/RTora/
72h2gSkyvceVh6oieelUYbj9hWktK2G9LAYimYLt+oJGjDsuPXDCvFtw5RtHlnspsGshG+6RkS8g
oQ3sIwksjIv8wcFtEB5Y285q6hjZw2FVWrNiF3nkAuQGoFnLIto/NsYmyK+5G1gNuLabvCUxproz
QEph2wKgGxICW5dgcuAAcf7WtAGZbnpORUrr7Gz76eIvPgOUgpzpU1q8R5cKPSsKZgcUFCtqAZxv
IxEsJCkNLJFi6ikkDWuxD/5PwPZaSVAco/u8rIVJNpn4Trnw3RV5TE9JzEK368K3mG1ZTiFwfEub
06vZIDA5cl2kfl3c1RKDPFyjrhN3ta0sJ2O1QIMV/ybbhtSAdsn8+bxPxqELBYy5g6yczzs8HF2g
O7xdu9jMXyH3TskpyYRKcZD6gBu0VuWwlTslKiudjGHb/cqx/4utwgmpJqjW+LUBCcZBkvfpyUWC
6B+qjItF+hBM3WhMaQg5owp8yrSgMzkld3KMWPfQH9jnglaFxrpj+76JjV+fsl23ZkbOSQePKozd
WZ1S97A4VIs7H/modmKkOKMWyBBSzZC39gH0IjkJ1rESr7LpdW48GmNxO6rr2T1rrH57idJQwoHq
AG95Q4Ti3fdETc99TYLO/g8PNhTqo+FiqaH9+SDYa3WqLmGKTsBAR6GwdP5i6sLvshsF9s/HAnYO
psmPccmdMgbfFLgZ8m49LDIqkvOVM5qFVJspihNNkiOT21FCb9tLCb+7sTjLjI3L3VP24nA6YlYp
A/kX3Fid4cg8ok4qXTEKBz6ZyIidZaj+eZuc7x1ph6PIlDYFRK1PwT8ulMbPzaBhjfkmP7n/rQdg
TkiNWvGjdlQDs9UZbG+EQbiSw99nin/WHVnycHGx60U2GS57QQbB3mytcYN0KhXbGAt6nmF2eA4U
uv8V4zkSQ/2ttPffNU2GDN7Ks+txVyKRylvVvv4qSoZnJ6gMXR3KcqFwutxga1pK15+tXLmQJPtt
iDsA3EBiRfuq9Ho5wb/RjPlhd/vqvKqu1ZXPE/3PAf2kRSXjHNWzRo4c7e0U2k8ggwyiVAq71a2n
bxt/rtg4Z0FXMWfr3GYIv3yKV2rbLFAZNa5yToRSwgaraiMJhP2FQZ8tOjRJwGb4rCPENGNZ6AP4
i/OZHGVX2HgcBa1VJ9v8ROsg2/hTowQzIzMiXXWBiwCDL0bcO4lOOUz84+Sl5tG8EIC1r5adZek/
D17l40PuX+svO4640eiLN0KXbhYVDzEe/SormS6kc7r30OFUH1dzafY6W3dA5qOURaGAaynLK65j
IWQDq/ccjJocYCs7NMfoAa3L2jIXsP1hN1ZrNV0KA0M7ZcuFXVV/0n/YaZ1xp5NLvYolgKKe2cGI
7/rlLiAHbPBlICwP2XOFL3OkU//sdeWiZ0bsvnfWxI919sFPHvnBMS3hNYky6ZN0lPL3d27Mtv7v
yHwAwbNHHSRIPRX1vaIMFp46o/pSToMRC/xSblGSigeoT2wMdW0GeyFZrRFU3O9tUlTv3Ish1xqb
Cj0irvCIF0W0Y386+qixV5VWNBH65Pc5w81BzU9XcaEPH2tGJ/M0ELHdPwCO9PAq4/wJ0+IWFhCH
El0H9BgC7k9kHbVskZmEbx55J+Rq5bphMPV75KyBywIFUXNWNuJLtNEKK9ncMxgAPcro8P3wguCA
mnb0v5MNXAF6luFWVsrTEI88FDecVmKwVCwOK92OlCrJDTxUP3KGCF0NLyJag/Kyc1SoAzKdCI90
eNiI7Z7d00b6TKwihgo3uT0+g/3aJCFF+oYneKqivoFvk7WkjWEBa6Jkr1AXspKCCncIe01eUglN
pwe9SrQAYOtgOxJygmnk2sMJc/Xqphy9iaeS2YBvye+o6K1iGAKk3O+9b7Zzx2nfR2gAfL6I4q60
EhDizgGEV74rRpOI/5ARKdcY/RBB2cfK0FQFZ77y8x17Vs8anDNpICT2m0Kf2uT7qoqtt0ZzX1Bp
/WFDtGWqGDPd93X3yWS++jFKEw86ICQrRfx21OzmJZBVuYKRy7h8/pUx5/9Ep0Nf4h+nZNykzvXW
Ow4ou0M5OGzs3tKOKI53pk3j9uRejJnOXuHNLpJH5YjJYOjqYR3AqhcYXybW2TG5x2mnNfT0gazx
Y1w4Y/TsI8CXnovQEXthPFf6TJVaGgrlY3mrQsdvp/qPBriGfpZ1yxnN+2ed2hLUF6MevVOjJEyx
8xYyVW4602zegeFPPoWyVHm6hzut2DBuZQEEQ+I2jWt+dcqzXKQdXoOSLK0dOgCkbKUlwnbKS39P
4iJ5bLaOZDIsKf5ar0bNU2ChRfc3UB3E1nPA9iU6CNV1Vb9P5cjZXiRsWaqbK52goFY4nwvfqLj4
wXmIOIK2NEci52w4rfMv8Iagy4D+8qtCqqt0tk1PCWpCajf69fSFcRIMjUpBZaHUIqF1FdfLiYK2
mJsjjYoUFiyOz/V88P4Hc/Cv2k0iOGvmQPad4TZUnhdGbtPwwNLlm/IF3QpS4uiWpvNTv0KkzMYK
esjtKN9uBzT3n4OyDmekd1hFGYJrny8E4x4RGBZImK10I7I1WXGzkTY6F7XCLzS09lmXJ57u5F0c
kkVcLJl65slj2IoXAm6hD4Ds3TmuW16713GmnvcKa/xy0lcd8oCOj/MmT+2pHkbohLxPhiZ3obW/
F3AJvPbR+BjWHkbJecej2ex8I24u6x6m79FKMrcmQJ4BmMa/t3YqPX12VjXZIqGezqyoglfBYkGW
Fd9InGkXUrDxRMYEA3EDH1fsYvoEVGjgDUmOdj//OhymM2+hD6Fps1YJN/rihcBWDEfyweua3khT
ohZkTNS0Nxvo+kxJbgO+3x67tNnFADYji4LpYVDdmWJuC7WdcOD894BK8gZHncI8G0X2je3Aq4Fy
j+wFbs9etULVeVACk/r4Hhn2wEajnVNCeHtgfp3fEZGsoCLauUcDrQpikOWByA+cfUAdpV20zH7n
Wcb1whxbLaq4fvpYnLC5ZNV+hd4cdlz8Z+7WqJF5t/RZZf9lacIYJXAwqas/OZeRl3KhLVH+J1ak
tncrSPbeWLv1/Sa22fZVQJXDkk7Cj5X3z4xx3CJnXKV4MZRRDJ7LAg9VYkX0wuNmStprqVCZems9
MZKZ9BRgIPVmFMiAcE883WXF8wZ00KbidUzHAXg1DxqaIlZ+T/s100kKyGgHT3aS8aYW7hTu/FGp
tjolZooDol4djTlEClkGt7FFObEweP/Bfziih5N5R57PAjxV+t9kAuuS5U/3SH2Wf/lDUrrizHs5
wOU6d6sajwAFpHEoyMpV4cTC86huz5ALzVAtvDGaEQJSdlB7+a2/lbLzd/ca9XOeP8PTjoZ2+SPU
tUVNVq+ok58NKvL4cl7kSlbq6FM9J7TyHG6aIP0bUq82Fbmv3lNf/jDctYjb4oRoM5z/rL2FzAtv
/GBFbMBMmCv7+tqlLQ7FVpHzXORIVsm5PB029/m03h/CflWDV9j5AJn5QBRVPM21Lcu2WwM4pAzJ
mlzEKea7Fwo2yRVQF0aaEPY/LeBuwM6qZa1THOr9izc6hGEKGS8sydCDo8p/P90lXYVxELVWbjDy
D5Xy/Cig3iEaFkp9Mmm4YrxhgQsesvt0R/0sQ2TiHuqM+c5eoZDBqI2jpBrq43XN8KhPwaSKYEJv
m6GY8/Ok/7GQUjmC7zVcnakxAs4Pyn2L6uxf/F4w388G1nf7mTEhnYZRStSGx3lr6lItzv5Bnzpe
YVkwn2oNAv9bO/8I348UkJWjcVpp76EsaCS14pQlzF1kmr4SYVHR3ZPajMaOR83Y7N+rGFNtAjlg
jbi+HB0vbnqugd0iRStT8Ot2Ig4vEYRhx+vG2rHcuJDOAYzpMk7GCJz9o0J5FdvBNeGQhd6HFQBC
1A1EPX6cCT1gzhMkmfkT8LMTIxAf0OWHIbZd17k7Wi3+TaVSAl8Hxx72OXyMgiViNQzQ32SlIqIB
jIi8YfkJ8wTRw7ezDkgI5ZhZaj4MUOc8cFTq3tvIaENUsF6AyAQ2C5mNacorEx4JCjKXrDiKA3Mh
l16TWOLVWlfKDrn5BhPeXu5nDWbS2hquhH/eW3zuhFe4RGEFGqgzeCmYpbXdQnMEvKHGcOgISNFA
V3qIxzisGklCgP5yG9BzUjzQODkWfqLyEy/F4gt3oDJXp/L+IIJGT3lTPeK1o6LH5oFj+ZYicI+8
wvU+520+PjicFR2j7BcxwLkjX5wgBEak7ENf/gEFi44efW9vBKe1ISo7SosTDFc/C4C+0Uzex6ID
tOC6OcjQ2CALkZiFnBbEP+07JLG53qi9vbKfk2g4fnfOWhp2GXXORqtJsKqNaX8RqP5hUFVYNudN
blM5eXqHBh9YJl1rarmH/+6rZ6HWxGENSzU3gzm4GYbb5nORZ7cLURrn9GadOQOoT9spOlTy0iyz
JRrveYNRgDKQDECHL/s9lDfKbjOsEoSacLj23e8WkwY1yUYADD+IVorURSmQw/dKj7QYZHkyYYtI
lcmeOHH7jz6/fPZABRrSq30c0MgTDk9Xi0PbZxN3EKvqSVUDJwA8PrV3yD/INFMFytSnkwaDCTG2
nqOVwMGV2OsjE6KUNIRLRUDEbFbGxGK4zUCyk4GQEDZGSgxl21zYSQZeVUmNgYR3rYRenfqH+ONx
/zOipsNrfqO+8+159e8fzoEK94q+Sp7Ahk6NqFawEc6ADTqy6vFhkrlYrU69ILr84Ka2qhV2AI3E
LfmLDRpB+YKGQR8KfL1MEIwydgPixapW+fPPEoFHxQSbXlsMC9ZSCJxW2BUtY6HYQ4USys31z37t
UjQKtQCfw3ISgktsazTnJDbW4+0xjRovV9ENpUSunhlILZq22xi2kBRS4RDmVJgVugRP/1XAAvYD
Se6ZDnmg9qFfxNvG56+omdcvNE4A59SICOxwPRHHVDYifk2Nqnj48BlkSAheCSq82ABpg/kfXR6x
wqUsn5T8kqWdOrAuaHs6/EYIHuVii3OhldcyJAUKcliwBpNv4OV2DDfm2mVGsUGdUfB5QvL82pkJ
KuoDPWnXoLc8YVkf5GvKjs3CYzEm1hkH8JuLV18Pk+6tMUPhew3ZtvTq9FWw5hMpw9h2xik99Vv7
mXQ3cURvtb8DKAkJGhQ2JdJLVr5YYPmIhJ5QNTvb+q77V5Hkit9xkPmDfdiwqzj1F3+XXHX9BVpF
QIbY5k/FxUA44LrpLRluXOIQYNHBw2GRG6g8nj7nTSPM88QbCtlHipxMfArkMDu9DTsQThRzwIjm
DYA5YbSsVeXAUHm7VKsWsv33WQB41vY/B3h5D5WjgC9dn0aYQiXZzyHltvYlNvyTMIp9FfxU3tA9
Paa6Z7LOvsctqINwx7WTEXdZEpHdB3ZddB3ZX8wGeYabJhRLXC02EEd0eU6+RZzCkctTTtjqtJMF
v0+rPs15n4dhDKmDdb2gLrlDkrnarTyyaWbJSvxC0V1TZBR49g02QUHFmO5pjIQ+xyIOizo/4Imm
IIsHAgi7/MXhJVM7nFaXhWhYogViLnzqLI2POw+n+gLPhZ4go75mrcG6Eid17eCYIw5gGZyRSDOD
C9Q2MnT2/q+u3oYaEekmRz8hHe0EtwYOq0/XS/p3DGIfQkCp5avRiRKyRiljROVWGAVI9Vb6hCOV
vCO9Z50bjZAsJU43X9jZOYZDNiGFUSV478LWlvUUxSf7hlbEZq5j0Y6lsKtfJtcszVJmIqtOkdXO
2YabndVqY1EpV3R6jtqzkbHUxGLxfh1o451B2MKwNJwYffeqaRqeivJfBO2ueNSR1H1OUyJiVncs
LB6rTUMtYVQA8ZmVoQi6+wYWSBKJqSkeGjndkUa+ZDxFSb3JK5/bqU9xzskj3DEM06WMCAsiC9L3
uJbkiz9R1nV7lpViIQUDu2hj+1fqsu4i3VOuQAJ/4uZj8uNT0WPgzqjH/lDI9dC+EC15cgB14cuX
PlVUsGozzAj/EyypkScOi/gELf0O02vgrxe8s1rTKZv3wrxj2LzH1LIbFMXUkV6xiVsUDb2/UOqc
I6sSh82+JrMWmDuOBUwE5d3/EtaEF1gG2JJK5z7RY1QOnByNVXheuRaojJLv2s1exFBCbiSbd/PE
jt2eEhs1An9QtSYlMNvNW7nlrW91p1j+0PLWcpE4XR/rjWh/Rsgy8Dvy4ASzF0ql17n1776PFxrQ
FPVw+0+HnO1S4THuicVfsLZgA1HL62aHqn544/DngG2muYq6Ml5KjCgjJ0VRvPf2VnrzX0TN2dUd
kgh8xllJCeCdMK/PK2oVZ0Sn4e8ELO7IADP5UzmjmI0QmiZq7gr9hEjd/Dxw/KlIUJvxf3w6C7R4
gL0j1newYDnvVncmwciurEeXAJpNRoznbHQOvlDLovrWtEdbG7j9vySg8VvARZ/r56QenGJrXcvG
IYiCd7cGD9HBTR8WHYuEYS+Zpbyn8ImpfaT1ezYxbNPMAa6J1VUR7+Qba/X4GktNSFssUrjWlz/P
c13/j2wEpfdnpaifjkmY/eq0GGhmSgBwDl6NhIgk0RYtPGDZ0prtLuowB1jmRXVdu3v70DyPaIRP
HWJklaFMoxf0qp/oAvewKW871Lw0EtsdcEKsyW3VxVKHnyD+QaakDzOgqwabr81yd7nqiKzI+v/A
xxaQU3MTz3+yAPu78hFVjtd5A68+VXD9dErHxVPO5PdVjEqsVKyzdbn1EFnwgSjHBcJBDvUOlLYa
Gm6lvhpFnbA1LoHcWYKlqiUsqX/k80cHkjBKgun1poFEJ01jEWh/0I28Ur4Iv2UvoH/72DoINj8c
QnF5Xf3cW9+lhLRCtAQcZlI9Hncgfs0QzQtNhCDCRKD5Kzr7wzb2YvxY4AqxT6+D1cAoYSy5vAc/
18C8ZRSKZLjj5EFZtf/CsDYr4mxfEr+mqsICxi4S93SlFHsbkokWT9Jl6mjNnq2sxVboPl2MreUV
zpQeJXXbYzyCsJZxfqS5DW2KA/Kel9p9lPxgV/b26q5Pl1nXd+DpkYBo6nbsQTmnVEwZA7KFGAlh
O9vM1E88GYNBtnpVoc3SVXH/oYtNBrm7OnnxfUxkPovwgqQSHQjRj7er9P7rjY/Dk6CFoe7hG/ui
Bug+kHBWbJwy4Fj5O8JYrQJI8ISEsg+gehuu/mcB4JnIR7c/gGfLPdVQLKu1UK8CIhEkZsS0MDpA
OTH80lUjetPRMUlhWAMvCT6nt7YznW/d2nq6iDzn32g0VQMr+Hx+y+zStI/lG7vfSfsNY+lj4yE6
8b/csr0jnZldZmOEl57Ip2V0wyVoDuMTKKhVSRHkAABQXbbbr26IB9OK3yQ2+HygUo/ITOJtCuj/
fvW4Hw2miSxehyDhIC+EWcnqLKX8hBHl2rgSACneRnLqXRTUc6dH6THHTOUlIbdHBe8QfKdQMSuL
5unrn+8/ZbKC00ploe3sN+Km1sWABRw/NJWTVfUOAVIUD/7tyANV+xBcWv+942n9tlDodGYH9ptC
lP2pV5nN7J6wCtS6cUo+SaOGJAC8GMKxFi9XAgjv66IE4KDEtNupfB8zOr0B9MQoYUIiF+Y68Dug
Tw47m095KPgqtMcnPFwTIyC4cukJa8u1cUuBa2nbwEL58jbX+tveNyzKhnUmyQrFa1B/Rx9FbenG
jvMI28XFzmh0mJupxErntJumjdMeucUkzt2uGFktH2zBSzpMrxdykWbEfRg3B77Ey05rfok7Fyw/
I+/4kI80fLPZOVAhc1cuG5gnm7iRvBDSxJU3JLUXRqFMfRt+IvdBkRhAi2gL9Le1xtCTM6ccQb8L
7urwRVZl/tEjh+g8UhhuUaW4veHAtKrrAPuzc6eq2wFotL3J0JgdlUuFqqqWAVS23YzgwwHANJNT
d2XWjSRgDZeK1Ql+J+UOlX/eDdtNjX6k/8jsMSXt2H5csPkVVlimj6IsTwQPkU2O+tMXwZBY4VdC
N8juTlUKRbVQ/UIPSFcdBSjL33drdM8gh9BOHVj+X8ea5zH/7L3/8h1sgd4osWAS3SYXVUCXg5kP
ewVI608dwT01NFspWGFNDlSEeNgb0VOq5LDSPb9R7X1K8pOkbz7eoLKsZWLSJigR6CBlqrr8mi8H
7jzWjqw7oXWfcdL4sRQphcH+xWr6Sg8Ys5uOxC54wlCWsUJN9qvEoLcX8UHE2b3HCuWwoM4k/4cR
gfvqUVaPDb2v806oJflMPIoD9+ed1Zy8wDLul7e4aVxFqXe3P+duCkFQC+HMbNIqEeHqkLaIOGyV
GKlnFvXBO/3CbOP1wHILetHb7WchaSzYhSgnqvm53I0cTSCovlJMOOu6zjKqmRZGLwSjyfsc4S2h
gso91FgHnWQSglNRE6GM73KPBBS7OCpqcWWduUhY68R2qbOlrP2b2YLbVShtMcIw+1CCHx+8OXpl
ptcXzzRFo2AAETy6LhWY5KV+CApF8AkTNb40CoHO3TPKQTfPIWkfkb70BF5BJ2N0/OKcklBEnkPZ
KUILBKuCfJr4XPMDq9Y1LRDI/7pQX21sCjtGggdeEIxZW5uwQV3TW27lHiq2iXvr3zfZNpz7Bczb
oJh2/UTgezE/IWD8wGw3mXn3I0olnmmDtYwnnV5rbLRvBDxV812RJimTZo4aPV8neFG2noXh1c7c
3tb2Dn0jU7wJxlSR1T5hsqWHiB2PJYgYgxIl5ib1KTbsbKuP7yVmsZVqqgoaQK8kuDChFs8Ptb8b
dieJbDklIh0d1bQOiahjxFmlHljgA0NAgOxQxpj8g0qsYOICD2BN8/c5HtPwcUkFhdBMm+mxpiUz
FMBF07J5k7JXTshCGeVZt5f2LwjCi7SMWdG7aInGjJCxhZF54H1nWqTne+JS5k5RfDTBkbYVq2yU
Qn9vEdtCQxlbSulRr+BMzXdYE2l6BrVe96ZM6a9vt5pCuMdMCTXM0CddFsxhbLmV6n+9H852ZueM
WTHzCAI1zIOUFWCWexNc+ReAOgCeUUVheX8h0zGk7leqx9dH0JHhJZiqLxfqph70Bm0PYi/POWgo
SHsyn71y6rvZiD2MZpnd3L4tdFsCZu0CwFwp4sqqH/OmBWl2BKXjDOe+snxppr6P1RB2CwaZtXXc
uneKiXExemlTLHKiHklIwxPobz9UtzUQS8nfFQVrocEDbuaPcpDg3513HIt3O0E3I2MQplNfFLxA
sBrqj3gICJ1ahTMZWsBX9v9KQYAbevrjxWFx7WihXNCTHT1YATdLBFXEXtJiOQLGhMtUcqSiwSSR
upsKQbMHxgORqs3rRXut178DkME69zXU5ptSu5vC26wosS41L6oQmi1PBlHwlHz8xZjaOwFpEGUS
aFq63O9QbiXpRJ8LuILgaYQQBUVKbUnjsYRvYDlU+Ohx5Yar8fK0eBPLOWhA8NYrq5g6WZ3fH76Q
Qa9tiOBsPjbunTCmcz3yhqEo737/gW/7Y+bo6X79F5R5MkCDKui/gzCJcPEO12RkzgC17Z3l29sf
ECnbXXVUgPgmnSDzxsHptReCpLNdwPGhGvDuhe4s62ML04RUMHQpaqcqIsC0F3jfJv/8Xrqj6g63
7kPjsmMXbzpMS8H8SQC74hJcZrA1/TQeU+s1CYvueKXSTB4SmOKdnBtjHDCghzHHU4PbuTVrX6H3
3wpitWB4WvOgjFfR9v7eZUMP96TqZjwfRlEbKcUVNuGjhTZo53lki6Aqc0MIX3yZ4CNbjoDo9I3L
Lq/svZdgxU6RauYQZwrwX09deQnLKfS4u9EhKkKME2G007G65NUDPMbuOw3T2jVQSGdZ2rR8WPaf
vA3GVtDswkNMxI9A2HydMUn3eUH6NHWeJT1a3jzHNCc+2XJACt046aditJcjyR/K2oe2U77A9pVh
iDMp7cc/AEv37UlhzcnYP2PT595QSV1+U3ho+8YJk4L3UDuWVy2/o5YiVbuOu5eOB7zcweUGliOu
3YKfbY5/Gv5idOHtLBz5aAyk5BHMg7dFkP4ZtFad+GuP7gZwzTxGFCghC4y14a7WqWNVoqnvpdFo
Cm0ovS4EQwIhcH3dNJMoEZYZYyFGrCTgH5U5Y7NPYx2Hltd15lzqf1ofkrYKRAJ+liXXiKX0496E
2R6fgtZOnceFY4vrS5pcdSKwSfPQ8MK2/gM2aoGL/m6e/5n348WDwz5ISq74CLberoEQ/mMPvWLi
IJt+RGcoS+mZrL+JBuodkmH7Va0/lIgAMp5h0l1UJdy9iO//exI2zBMPn6X4392cpqZcdN3uqUL/
EjDVpy1BXGrGv3EXszkD210DM2mALUIreK6ASAQJ4WJuXDGcuYAcoTNHsybLxV5sjiuZ1zIQrxRf
g7LnNq+eWUAhyH1xF8rfcECqgS+DNw0Ln8ZHzbeSuHSb0bfoeryLSVzMdbhaqmbpQVq4i6XwXcOZ
6WuOkTlJG4cEe4zZFsxjvRWdgCGahziZI5TCv25Zl8YTTW/dGKmvxIE//19pQQxPWjfYCzjOFYKA
muWQKIV1lRnNP8vwHJ744w1ydJ0Scx1cD1bkPOQb5Jn9QGJpLVbtzLlgN4SaRge43DHE8/1GYFJt
D9RlUetJemmFqz9/UCeJC4Ne8J/6rnwHimXobqNoV997tf2Uurw5fyx/Ofg2t8Hz43BlM2HDZZSg
dTZ0OaXIWxdJmv1SLPRGDSV5OpUJgqPzub6VzBMUsaWyyXSDGjl2N0tYxsFBNpm/yMHdIHktmmk0
9bFtHX3Gr920N3bpp8eR9XnC8hNHwSn8tQ3joY/V645t4v2+qqszCH8HhYogTgOY2+HSijAgxJGM
yCWZZJ3UnhItcFBHVMdUYD0pHsD1+DhHXLlWgOGJhx+pU6hj8bC3fHT1otlogYY6QATWtS0ZhdWP
K4HaeGCfYXqPBvgWrBlujeZYBrpCb660cIE/lW8V70QcozrksPgPkw4KGztsP3toVznF2yMLOmcx
hvLbTiMBh6qvWbqluz3NJ7J+fdGylghrt/ZWWegWjVVdIgIQ83KbgsVfPwNz8a/+5U2ooCgw92s0
/c6v/GUlh5Q80ZfhdiKD18C2YwC/wXTbcILFxSntgFT30ttUtauG7cn4zqmNA7nhC433rwQr+3d/
frsyXxoPpa8DKk5gL/xIgPvErnbOs+Y+aN8EQgAW9d5HWUsVj4tMzly5gfiylUhLfrfNBafy3AMq
LEvWyQO7EuToJyeesaRUqL9tbGIxticSTD0lZfDpFj69/FfcdpzO5v43ks4bzzqtnVDr/+wQnIuo
uUR9fpIelmAPhYvijvxMAz7JnEpHMkKwhwDY6j3iFy9P4Z7Yd6O++cF9MG9j6t053lMv2/aXYJBB
jxKwfWdI8nuLOcqOSEGPrQuk62Y4V1jivHtLh+6TL7ndk7PnCU6N6E+ZdeINuYjcGoIBCHuXP7Dk
9Yf8cKtd3StRpyZ76qZDc1nUv2GVMerLc1Ri7Cegnkh+jcVy0QzrOcoXIDGZg8Q2F0uyEfRAemSq
P2ULwl691LLPtO/vJ2HjapT7yLPyw7SzNidxYtp1oo4CHp/g0GdZYGekoPYFZlONH2Cvuf4p2ULj
03z0B5AXNGtVoKwPzhxQeHSe5JTJqgcwrAESoJPGVoaXWEUmfi8VFTVuTN+onBhfw6CUQDgutv50
aY9oauEl0/QtZHQ91WBbmfnmksh4LE6PTW/QH/rTNgN15WeYgLe9LGopxvigdAvVMjW03l2asdxH
aSHrJ9x9Cb1E+vEGeRTWafbmeZOvq95Ulxu88SIFnPWwed0+UsINxfliCdvSXzfJ5KwrW+IW9H8u
SEVJ2XSVJ8ta8w3pZy223w+p+sCXgfShih1J/y3k3084YIu7G3/gnJ5Cq2+N68PaRUndWuf8s7T3
Z6jArMK+kBFSpo2jRyM5mbX6wyIeS+OCuoqbETwbIN86baSar8ddSbMmdV2s++dCJGxHX+g5YpvT
i/2U+9Z9TIo7/gq0FXlnuO8y3GinxnVNeBQqKbuV9alpE0MGZ1BUsT7ncM2taXdrDjAykhkRcsWe
KU+sRJukqaUA7HlIAjNYOIt7D8DspwM1YagNLhZ9bPMH6HMi45oRLmz2m63ECT5BxIggZ0CHkOFg
xmiF36gk05PudTasJlS0gUp/Xf4ObL8r1FrVol2xYVlH1eRBfdsgPOCHlBpQiDVG8Ev9H5vBB2jw
GVbXOCcf5q0VdI+CYFHUnjftbCKa5YF6iram1REYayFOAxb87k3y0L39inSL6kFHAob05L1nmdgN
8YW9qPNWbc57JGs3Qp1v/7zYoZEeVhdrdUMxnEMRLUA849uJlvSDjPcC+jbSfRWkaMpCN7Ly0V20
RTIW3IH6wccFZYHmN/qU549t0dT3Yj7NGsQkEYyAGGShhoKYgpPJ2GIFC3btmP9JVmJGbs+XdRRu
rHBxZ2ze9pQk7tPuiog3gwrivLIKBTlGCNPvWApuYGNOLfGGMCVgPBP7pmdxKmhvRuT1Ld7rtI5I
/yFFc/d6yONSgLwYsESEIUEyfEpgZWx58LVYCgPqjM9FWmAYXSjOhRbkIQ3KLtSzpYXcsFfkMSg4
YawOf/mUQhQ9c5Axp8r6j30BDMiyY+N1Tz4wlDa1GO+FaA4vnzZ54dQRHJOnh7xbA46uQyjLcHOX
9nP9nCCBuWcfuDOl+O5rfKIECuvRqKqS7Pza+WFOKurYAHGUBZLncq2+rUHM5n5H8LZ9qDH2BB+e
ffOTOaEKjiwp62W6jJJdEHhIxnSAi8SKbsQvJY9kQZOeVBenN1F0rxMgUX/I6SH1C5tBOd/OfgX7
2LD8BXmsBH1onl7GyWlztdAcjnQkDKj36TrG1ji0L85YPCK9ujqk8ym+xX3brv9kI13DPpPXzzRZ
wzjSKUkFXAsHnWtih7tN4kSn/kR0Pp17eTSth0b0zxgpB9hl5B3UoLoxGr90Q9Kjoqa8sqUT+pa/
HtOtAQJWwFnG6ArTkmQe4w2VZ6vf5hURvwqpZ41kGx4mgkX1ALGnyJo74kOcrkS1TS+d3l8gGPEv
7rpvm/cBwUuN+10Lw7eYlg2xO1eL+sNLqwbwp+PyIPTdP4td1LGHcUAGHkufC/AYxy1QtNTNXqC0
ZsP9p8Vm34ah6E57fXGC3s7Ddb4M/ApeMyfvrhhQeu48jyFmtY1hvvj8WkG9heCJ+z+fxTA4NL4j
BGgp30wqxdHnMwQ9jgbwcGg4fFT70QEWWIHHf1EfmyMvYIXbtR/AtOSm6fMqj+EjjjJHn4t/DmVa
FGXLmQFJsUPt9e7arwxWOP8Bzhwe49w4CjG03nE6tzwwT121bEnsMeO1RQINw/yDPADxnDInbhJd
QBqjaVun4cGWvvUYVLcJQoJoOwgUxHewaguZ3JfcsuCSn19blLx2Vi9W0L6yQSkgeiXkku41FuRZ
QXzQ8neLiF9DkwIuMa0Yab1UZaY9q28i6mqO+GG3e0lFa3MY4tofm8T0+kpphOm0yqhplQIES13q
kONqWLGa9I5vThC69NbmuN5tNfBswWuvDhMeZv8CE7OkU6V1pbrJ4g50lXfCQTiwEJmKoRx3/EOC
NLSRw2TfKItgHN2b+gGThwbQdATMgKrf1OvdMnQNt+hfDl8RE9Fa5pwqX5+aBaHhJro8rO4wkVvs
PeDd+cNdiDkU7suYFrg0cVCrutEPsJZE6AntlQJeCSHGwMp5jLjqCblAyt1PZvilGVQ/3XCeohcJ
xolxfsFMqiGW5UvAmQ9KFD4f0q38BeW5E3EahSTuPjUVijif2vmFXGMLbmLj8HOzqgxB2z9hSe6Y
7JMDjOw6GiS4x0+F4S/jJfGHza1sIT7oAE9+mZyvlfJc+k1KHs3ucLi7WWlhWx7deTO+7wjPwH/U
a+ecra3ro6+nu1GR5AKhQ0YestFs08Qm6QoLoenE+Df184CiEJ1O0t+PQCxruDfEdcvmDmfftUoT
JtUmJx6N110qsf0jwWvJDNwS5cKWBxF7uxVZxR5XpFgyatLplRVAcmzZZXXXZsMfeT7IJR0g9XlE
UpPCUjvxx9uAw3js7BOuNQcbhH+/zRSqlFhNGV4gCPv8FDom4jpJRwt9ZMgC3nJhFHs7Nckww1NS
SREaHelMZpuH4sF9kmWmA6M4ZWui3a4T7KiNmfo5M9cY6uKDIoj7yn1sF/Tndh6rs7/IwGJw1zCh
P94M7D+y8tKsUL5xvcT1U0EDS5KOKIJR1r7TaOMc1LU3dBgmK7G1hA6zpa0jz6KfskVy7O1FLzJQ
oeFCbndI1KWERIylFpImLe3hCzdNwU6WiGauCY6q8zq8NnD3dNUidcOGia7+gsxPCUyYdbLcsGEA
oCbq/Xb/6Psp1P0Drd26yBcUPpMSOBX/T4M7d33qowKNxURQh2FZrNi5LQoUHKNuKrTtIJ3KZkBY
WnJqu2XAiXav8KCdIjuM2BdSwD/RD3FBfkq0Qi/Hj4trkyqW9epfx+VZRAZOardvVjb7wJ3FwFW2
RR3C1GlWxhODSLRi+1LwIj3ceTjZ6K5ZVhAgdahOnUR1fyomFPRV+WyImbLVvdcn78boXDYYbxdN
IMhetYH+KpY8NdU59hWUQFAb4QQnmaDTSCfdEFp5/XR6uWRwrPYhORm+9Syx6p5nZeFl1kbMSpSA
MOf4fVFL5PAMsMaiJ6+kkHCmfWMAAMYwDmgJIp05Gu9x71d8PjB0qsz2nqRJYUP4kguCqsiKUe7w
1ZpmHBUrnbQ9jwWdEu21IPo07k/FFrnu0Hx787FLBFYt6iQr7bkIHVmHqXunKmJgLCeYX8cQs3Ml
2UVYChjdiTzmm7lBCZrbJO5zRjO/r+UbQdsTepAHfS3xVaw0EYpmjxiaxgPr/QpKH1X/gVR57q6e
J8cTUKyAYfTIGL90xdRoae1mxmnWH48rL5iZoNOaRaMWZ5gTRcy3USHTJQAd14qFaSwhPA0qEgfG
skfhL4+svLJFG+DkT1NM4K9PIxirccE31R3uG2v5Q2wtkZay7an2AlLmDgDXa9TUKNZ5pvm/dQI8
r7FpaZlF2BtqDcEWxR4TC99hhW7+qH8uZj3CBV6ZbUA6hKwYDcJS2GXrm4J52EbqaULvFgvoq5mJ
fOpI+DXQFDyaL7P4jwZSDDMsZpO0CFa+vCSt4qRfUDvGkCLaX3ZP5NUm7aeIk7araTodKhVqvxGs
BP1faia+WLix5Z7/tSO8gnuWbVvdRXhhoxKivrOB4fr/bBoau6Jg2zNNOmrVzMFnjh9QtwE9eDPX
eBzbskWfz/DRf95Oam3Es6enGgmtd11D+FOYRjJbbP82F1cxc7xNmF6lgCooAFIqDHJXBZiFLMle
PdJxF9sK8MRUXUPp1y3HFo3HfZc8Z5ZZgHXWhNhs/aV184oDuIXqP7EAmMIVATN2TaAIjaysdTvi
fI6MXjbo/ZUNPzUKJJ0/2xUXeQYVSokmJcj+pkcHCZTg41T1sh9tCRtcEaMtpneNbQ8p3N2Q3Xyk
d8ORDR4agMaJDCk032wgsX+0QOPdTZviEe2CFmZQmh+RcaupzdG0N79IRWEqb+z7EU7rZ60NbUM9
eZWamhw5dnsuJ8DjKOnY80dTToxtlSXlXfW1e/b1rR1MfrctZmQ4jndTexLpxvGZxM+G3A6vM+8+
g98+Stt9kNn4R5u1ggTHZPi2ze9TQN5ZM2tWTU2F3rk4DQe+xbMuiOFkE5n+dzXgCY3nIkc+y+FH
BUbjiBrU848lmIqyQrbAUydWrImRuZqP5Pao5ETvGW4MxipoydmJtTCgTKyCfRbii2zefdebIuTF
nF/9go3sLxz/gqqE0DJs4fc6m5kIhIJB954KITuozorI9VbVwhjuRv7GZj4sG/OaaMsex2y5KPL2
GZEVtrKCM+g56bm4iVCCWD5RVGATfNuPGYdU1SBGru7CL77Y7qt7JO/485dEwtui9IhmKkwl6c0s
qV9nIwhtg+5hbtaAKrWVbm9nHloCRTkpATMEeUpRVGomCXyOqbg4QDT9NOqin7jGBaG4eKfEE41Z
TNBtefGPOF4r1s4hGj1plH3jhsJyaa+ESWmXkmNNvDrOqp4UGZPH5y3+l5fXOZ6h3BFtn+K5hbu9
X4rn/84p//3IrFb33iUAF9zzKtFfqsMBzkWoCORGD0p+C9WcDoliDvcNmGwnYp7FsFg/O3ZxGw+C
5/3UB1arlrTTS5gz1UnTl5hS9BrjPK9e0uHB84Vlsim3cJWYzIhN2R73wDoih+Wyu9UhR5bgiNHc
yVE7Wqmhj6pCA3p0iMuc+zmAIX5V7LjQXxrkUicHaeJjV/8Noxf62HDCYPkh3dKL9OCGVt5F3vLD
4YGj0QNheCQblYc8qEM62p2vIzS8Fj9TmSE5ChgdO+NzDakMCugWEs2lhZ0Ur2LjBnj+ryi+N2xJ
Bjk/jRbfyMdBhHBFqtI8HN7cSSc0xGWVEZbi/GkgFcT+d89LADKFyrQ/FtrJxc9eLICiogIKJ7WE
+HryTdfM8YvdX8oT8OVtXOguCd4OF57QjeyIdX0o4GbaQMHbzy0neJRO9wWERH1nzvpTgOoq3dae
bAeMoustmlRIiqVco23hXosMogH2xxHzi/NdeDqGuJ97AtwRNhjMryTdSPLRr54UpZVKCSCYPw5X
iRAyf+jhMyPdmvcdtdSlAKyfBmsUHHvF9Ae+efQASSEk3GFqtAcAwsCrouvmlmeIxhI95OFcuJld
haVGugn1mDiF96EjeM5iAlOYY+dcy1IE+o9V9aufPXhcIuDzKAJGkU3CkPfkf2eItAXKHDzR+UVr
ajL3CpjBFbeLLDRalfEFUXS+PDC10mbZaEMxjPizq96lMQmroY0uEwm7oXojopwKqhK5Z5oe+GD6
FhG8KfgxfOHUU6MDMTcnA4YEt1uqgKWPfhFe46P+3HruSXAvp6G4nSKWy9oXxIFQaPKJD865wnhG
F77BS80NefzNzMfCICH2umCkw4b4cn3V7nTv2k+nI7GzY73Czonoew//Ia7o7FFStA+XrKzxF/aa
ZotMlZ1RoiKsazRqD+tsU2aBk1nSQzLFyAzbnA+Yt4NNO/tR6192fcfm59+LblskJQyzoSqShfOw
EV8pd3fIlnhW7maajHPJO0wFiNO9sSCn7IyCW0LC7EnmLhkOyqBTn4j4EiyVM0STTGXoc/FKC409
qqEQ+JdiVohzfZEv7DuGQ8Luh9lsQi4CAtXCwwVZLDL66zqeU8iEr+1lrCBiw9EfWuz7bMRzAzPu
D2N2ZqCVtLNxP+K3EwaC01gkNCcON1/1O+oyldJ3ncEtniu7guEG583dwy93si9wE2W2NaidbiCV
1SpyGPwxz86FsSVLki6dc+RTa71SaaWGHfb+tYc+hydFhbAQyuXOAW1k5G3R1SgV00LbJ+MD6ESv
ollFWfxpbZ+WBo7lIOMXN5xXQBkVBoR3n1LEZVzXEDZ77fQcSFlSYtN54D2puFcEHlLqvx6B2bV2
SfOE+A4TKw5+FLa0NyoAdzA2ItyP51TU86LUIPO8Vn18RPr0NBVWYdhgRMjmk9MkQV6ftR9i6/Wn
8Cyc0kHM/HUMhA7U8/2s/Uc28Xeb2x4YW8Poqo3Jb36EYHvnOMHDGE2gKqfHY998df6BGrH5l6lu
Lz/q8SBggZZVqigLXoMqL7suyJ3gOMTqlsw12m3TfSHzFFqbuvKroSIjpBOj8sIg0l74cEGchnpk
Lo4KFUryd4S9DO8na+Xf43hbYlWh/BZDyOiIxU+yNLuyr/vuekjBA3s69TTT0x3nz0aGJjciX8yD
WoCP52LyP9hTbYANSAbQuipSqTI2B9VbKqnRyTWKiE1ol2DomGYI14hHX3/VM6cpmD/dRyUhpRmN
E+Fa60CTiOr+I9UW5+Cmp+//uVCBdRUNAB7GXS+5Qw8XrmgNKtC41T6/bRZbrOE6PpHgPem+Sv0n
oL3oZFHXMGMkZm3OR/Faqn1sumtt3Pk7npRKvTCWh0E1OSO0iVzYcMpgJBx4Z4UO1RDpdSv5HsPi
RRO32pUfQs774duTIKp33Wi8A+UFQoPtMPJgkDOQbP51UGJ+KNbtdOAjzykFlCeOlUOlPPMl5aeM
RANl1ISssZMYqKORV5QIfblCols6q3TFZaxnQB+R09jB3P+uB1mpSzAF/wdL8jpbcLB5Kd1fA2RO
tldv8ixLPYeV33nMq9SZm1Wtujmnf/zz81TAUPcv7T2QvUR0tqVEdjfIH0w3vj2jTl1+N7jKQL5A
3c5AG7BA9P/lpJTXmho3NgCVHeRWYh+obHiEyO30PVTMt17oN4LZQF4FsEnqLxooZZww8TixybyN
QlN5xxcT3KCFYomi2vi0JJQBnUhiX4duNJCXPGdnsuBI8A4xRbHaDU915nwuYMjbSPjvWSueytQ4
xUo/shZ4W2SjEt/66sB66Q5GKJHEgs9vnnAnp0fcHM8MDRm6ABcipws8V1cqk1M1rpQXBe9eP9/w
iip9neuZckHlaYTGQaAEKVSfZSMo9EW3u2VKyjY7CzKDZiITeIJUNfZo+kyuX/+UM/6KvQ/G43Lg
j438mnV0bSx/I7cDJLWTb5cow1m0mWP/PPr1hnIFUouHmN++zqXQbWQ6U5E7d9qwevTplo1mzVL7
7SbvKtLxO/W4OUjpdQoKLEddEBB17j8di0y/2cMXS/zcHupq8ref3PsEG1b1wB35X2bQILTloQ3w
tQ3xtxnmM4lDUO2OTbacHSnEZV0fnrxxwAS5P3+STZcpcy/q1a3bcEx1oFLF8p8L4UwFjDntZ15Z
pv+1Xp6FkN50p2VgyhQvsbT13jOInLC93KqDMUv1p/y859fKdjhCgs/4hBDugK742GmgvYF9WbK6
KuQ+wVy50RqXZ4aPLZeTJjpF+s9D+eUsJf1NeOiVKaNu8wZiEsRjNt9rfdvDFETfxUeAmXAViSRh
uMp6QfqflDkPiB/bKVIuWCqRDL7X5UZjpqamkJ7AmGj9uH6ztnd+HCDS+SreyBbuFEpeEyhsBwp8
0WUUJWLbGajRLeffJyWBu/dJXs3BJOyxqLQDM22fT5YZyI8G4HJRpTTlus5WblkmWiiUOG30i8Za
pDBVapYuxLs0lH1Wjm78Wdwn2TRZQ4KN3IqMAEAA2pYKwRDHZgnwfXIENooRfPwj/mF9+Ma+R+vj
Rm1XiCE6ZQzAXb9MqxFhxBq9uFBq7nNgz9wOHP7VagHHgnMtwfE1QR8P+BaD35J4lrhOz70FoQOM
2y29X3lzojhVqME/pgzRKIchEwcUbzwhWf/wXaQPmrqxgqTv3/1fuC1FJ2KAmi2ay8hvJtahgSxC
yf43UZ7Z9tJZCQzLHMPGSd2UyKbKBpcQ1CcaDaA8m8WVQpgfTGVjpv9h1ayUyW2xBqpPvgiD9fEw
XwGqikstLR5yMeQFA+v2alICOeeKFtKrgXSrpYY7cXkIwe+5XTWV4r3SOh5TtGllVy4eqSzX7COr
l++BzdKKssj01FAgilcGGZQGRN9jqHhUzPVywUMcb6DS/Mi/cazKHDvccSX/bQ2DEEr1D+x98LQg
dEqViHiP03GSX4YVBkLSThgdKG1yMIiGX9UJpbeFRyJwDMXCK8Cqg5TxSLrVKMU1r0w6eL/KyYEw
jMsfhEQNhGT+7wH3cMUa6kgKsYv9wBFBIl5N9sHpOrcPwihDe2mvzbxE9WHZJ7VMem/acsAYtyzx
eT8DDcgUjGyZ/s3vbw/ZibvpRGHseC27OwEpywJ6NOoYzGB9Nmtn0Ye7MztNqyguVQ2+X3LJm1ol
vzuctMnAMjw6dAf+atd1BWeKs4+vOKNgTu07pQCgfdiPuuQcX5AlDkPWrvUtp2cfaOJh64zOQI0w
6wg7p2pSXVUKruucbRcZ77+TgZ1XDfS6siuGjf07xv9psIgH2/91CqwP7+dLIKaDNWNzEp7xl12l
BiTEFYoP1uUtewBj+Ve+Xo24SQhiSGoclTaumGjchpdzFhqlr3sMuz8TOTMWF6g1HCgHWEAh40mK
ddmfhEs0SGJSKWtqUHslAuD7jGOtx1tEWoo6Jr0uUMCBEOv7AnmG+ct4TxY3z7Lat9tgUnjFQD/P
WgftGMpPYKtDdwHIGgEAJfssRLeqKRQGtQDiu9qRs+0o4KiKcPfWqWxuFpII3IBhpv5WDAPg7q2K
7n7qawOJU+0cy5Z1d6Ws7DPmcpigBSfZ0q+02ROFEIAz77WNXS1/5XP4VWAW7RN2k5o/TDW4JBo1
IRmhnn31M78SgIxAcGLh7EMyAITgcPe9EMdbap2GJ16KMZMaU0AvFoZpkZ3EzGZZMsRrYHquf5+5
FTYvxvkPVRc+sjbjUj91bix5flW63M9Ggm8/K9+SxgZMgkEDvjBSuX4q8JJh/whoJkz++TjoeHxP
1j8qLu8sYlJLb8dkGFRoDShxXViVQoMpaSNrbCnBi4ogiAzqAW8zLEUd1SZtb+QSMZfoZmJOsABf
XLuQEgrb2xuxzGkJHpv7b6rmBN9+GnmlkZf48z8YJI8jsknuKFW1TJ4hYf90iumZiL/kkHvsO4z4
dt1bCqYKCN2s845amI4Z+vJp7Si1JLKZE7tN9vvRglIEnPex28nR/+wxwhrdzp89rJD8rlOQddGr
1ne3OfZCeYm4cp9I2BwfMVqF/7uVKToy2Zx1BaAjYq+ttYpb9oup7N1u1E+/gRNi9ArpE0Zmd8eX
ItHMQTtBqMhGQgEkg3e/vGQMC7CHynui5qfrZg5jqWkkX9cuIhxzdptOSucAlRjg9/Ynb+HJHHVI
fVgR0boJ9r7LXWJkITRNRr9327ZjUIPPDd1BKQxeEx393vJqrxFvq06tV8zwOtaCxf2K+jnW52oa
E59BCvIwn0CrWe7EvbdLw2+GWlBXUrBrwth8ZVd5lgZz6D3YVE8NA+8RU7MeigrrIdLxBBx4MzY+
RhbqteHl0+qksVXCBT75P5NhYyTETCeAGXKjV7cjYEI8PlnvRaJR/L8XX5ddsldS1c42JiTzpS+n
FyHo9GH32aQsYg5wwFKVFf+HEUspdFc2/WIwg0X5EZSd8DhI0UxIfVrHYmeh/e3+O1vUzuRPMq0W
mXXsihsAzUev5hKHH6/wbu7/nTPFWQD/cTp4BHSpESwzV+iJTd/gvSMrU/Evi4wzyUBjO5uvDqrC
xRWMIYe31dTxrtqyItMtZwCxNXD5HtBKk2/e1T6cmQPLy6Ro2TqFhgaUJesl+Pt4mD8wK0rErIWi
PVUoUi58AseATD2G3XA41CTS9KHVnG1G8+xIvfPiHrtlgpB3casUNz+kFqPpt3p8MvQT8dLCFm2b
NP4QZL7y6mCCgbtUL2ZhcHX5JZyD2+rFQg/h2HCKf68xNH6I2SQajrXGI9VQ/Zt5CdbHXAX7/UYv
DWpeEpJ8mgjL+06hhCuA9PpjThlZFuF3zqkNfLLyQIzOxDy1FuM5hx48rvaPrTHD+vUUwoIljycr
2Z5QUzWidSp1p1jMyitnl/nnVmIwhIoousHVG92CYApm9qQFexInVb1z7Jc/uuV/vy9NiRZAlyiA
lsRQsMlVsQXh8PieNX5YadoiJ5ckcdR0Nya+3n4mIIPOL5PfSFFyStvr1DXY5NYV+23JWEvmC9q7
NdPikh9U482qognmupYoL1cHbexCM/idAlLbqwwA4feoz7q+wow4OzBoIAab2ijac5xv17I8gAJG
HXVDNYQdzNwuDbxBTrJyxKKX+7q8hFUq3nWWQ1cfEBiT+gobO1ux2kzkI41regK641+1jZ1JfXBK
9K4V0GdozJHdUJ+4V0uWtFKp8MGRPbwSF/hwYQfjpYJn1lpPg/20WK5fJTwF9voYjsqPvmw3ERpX
jB5J00lmgK85aWRMW81BHBiGRyt2O+zuIKco7vbGQeTWg+a3agQ3Kzxldko2ys/7KbJfMOgnzYN1
mCEHR4aHgLUXtHe4voMLr5UIckraYNC5e3k00XnSFDil6Fy6nhgzqnGzco5D0eWqdazJpy94v215
yFOVV0trbh0sYBI0bC97bH4gFLQFZjedxnfGhpB7UJWKnj6XHoev+6RkcaDH2SeYLLGX41OXuAE9
g+exJZKWMoSyKEIwPzwbobm8yxhmzOgQS2u0DyP6svGIwgD9ks0hzXqr/Mp8iG68IyTxMdA7xUYJ
HhcgXYPkanqpvhgbza+W4m0dPAxu/69igY8KC+P5HPqSo2wZXbHI4inO7jMdwZD5HUfd1NTlSg2R
PY3vKDyd4c0AePRwaysdv6zbp4H4GmZsLDRaEeu4EXZAbrQOlWj69iYGQpkbvZDYDdnifo28+Odx
gXL3WDFCU4mx2mxst1DjJ/djk47os98+Go22lla6VLCXv3HdtBNwpPI/2OLwdRF9KRlKfivYyI4L
ucEoEZJ6nB9VdXfG/7lMVt++r7JwGor72qhoiszPkyfuV7ASVG42DQGCjOf+X539B/KOafJloLgu
FynUAp1FiEJC4qz0pJy+6nsz9Vq/Sj6q8IYSejJXHwCQF3ok3PV4cMKh2JyLRaOw6ouFarCuvly5
ibBbong+8/m0G27Okt7jhE52N3iO4leUWLUUJGMwYzgU76ofZsUg9JgAI8TDKaAuIvtMwV0vhya8
Rns30GGdL6xCm30HhtAutgrsO4ba6NDuwGRsszaJqL+kPz1qETs5G6psgy5OJncYkR0nLrxiMb8X
qa/YkRZv/ExBEZdF5/7hNTCE7YrF0TewLz3e7wcRkBjI75xljPGUxMdKGO/rADHW92jAKA5EbO62
75MkFYrXEV513pu1PjSrIfSVdLTLO3B4fLi6vxCLATGxvEKDnrkfukrS0UlCgRMEucqQKGKVfZGf
b/1sswbROPjOdRgUW6py/hLGSdmlNGkuZHUmgUbGhGDJ77ysAU78vB4y6cCaMjBRLHcyy8OYE6OB
/t6lNlQu11G/E8Q6kLqpcoL+oTPXv7A5/kjsNVd+bAtXjCug05v3oTem9d9JB9JJkFHNL3C8rtkR
AI5s1O1C8N/KsFOr30jBYqbUhIoiBOOA4c2Hy5OC1HlDpk9r+AXVVwBVtpXHkRjMTl3IGZyjfJ8S
tk2MKt4fjIxiKA0hzwC2hiRa0vciAPY2cU7HTQeerl+zMHW9rBNIbijCempHO+b5ygOYN+YtLQey
SiTGcVT4bVt1i6T1qxZ066IFlXWjMllGuM2yK61ZfL9ZCtl3RIM4PurJe4u2pUgn+qF6ieL1zaLa
P3ueXRNcQM9tSVrK97JJ02R4aYSMrxcLuAG1ugy4yRLCu55p7kbW5wH1FbSmMXGOeZrFsebWLWxL
u/XbEhfchqeomk1jl1P8LjVMS0pwmMn6NKPuTdZLLCdLAmYSV2hb3Kvyt7q8sPhk/RXobbPYb1Z3
KsyKvnkBmE6VUQGZjk1cnInxfkZ/r+3TiWk5OvY0iTZN6XzyUaMlIYzjAhq59OuOdLk9LJR8gUs2
pJtJnzW/6NyVwvLM65AKytzOISlRdSbZMtzCjlHjinjnrEmzfjneYhvsBxgDn7KN8dFYqsG7q0ov
GXAVqcdpj6/3v6qYarwEkNWEZrQTCySqtJh8RqL/PK+f9tHHrMWXeYERIagRE9yd3VLlV0zAa9PT
tvwIzFOi30aIsqHEz1gTchQqUGQ493cUXY0QBykWTSsc3zCAeBEB3y8urL6b737GDMt4/5IJmW/L
aORPg/7MIPl8CIVjfQTD0Qbn1TgY76GJt1m7nRAmwRWhDHNbQSj3RTu/A1fVVnZOoHssPAsnCSpX
g7BuT+3tf/cl3AAtQQnfUGPKBM7fyidyIqGPePo8NzWdG4huYPsKyfGJ5focwc0OtLRVCmPXloSN
ivlemcbceFz/zp0kJlTfj2Zbq969MJsD4UcHV+qvSg4bmdBBo5gFhW0VJnynjQNU7BwfcGQJ7ibT
9fFXCWBRu9qahr3qCJLLKkBPAcj6yjOZpDxQM1QRomfxD9kmEp/PNN+TYK/VHSPc45IRUKJQ06HS
1PvRjJsOLKt5602f8lMP/NOaQEmTq7qSTXa0At4VlcX9gm2163ThARVoSA0e8OTbpxgs6qvQG+yJ
hiuUna5/9LXZ5+DKrvfy6auafCliHN2W7kIAE7QHVwuKQMDDXhw8WFKWBLOY6ToobInN31Ackt7A
l0qzz1Bl8s0Lni5mhZ32FUNsrvR9e7pJ0Uj8SPIgHFiJ5hlSEU/xvphAFFo79SUCjwkyzeK5OYdI
78jcX/8cVECrM04RsT6rC4EA6PdIw6elCz2jwKjXgTfcFWi4zP05UwYTS1oZFemMFk2fHkkRwlFX
Lt56lO2dv9tUnudZ99vV6FYgcfHZjF5tDN/yVW/eccVrZIGoDI51CVRWrPB/982kp1QIvE3zuvLG
/3vGxaaJCkdhlEWFVht1Sl85VQENYuBMbJXdOM7YjsleFt3HafI2wOIbjQbc9u/+xo5nBwag8LyZ
iOD6xqJmdb+9b7nnsQszYp/+m6JHU01FQUTTDgD7PXMlwxvAXzH0JsRpa2XRoSmrWxhSjG14YVDR
tJJ3zqUJjtNZZnx1GA3vbM0GwkJnzxtaAzwjWCpfZQr76Apt8XMxNTC+vSbsvmPiqfkjagPjgujY
Lhdz5cHXKbpOqsS5akub0/6fAuGAP1izPnODT1P7gIicLwYi4azWu/9zd21Gu//SDNTK8yngrWfo
ohks+UYsU/MtdRIqrAHzV6GIX9259GlPdsFnmFkeGlku3xQ5X1mXHWgt5dI0/bozusxAhA5Lotmm
ku+CWaJbfMPI6qLi0Sx86AXetRd3ywF86J77XVyt9D05pp31kUgBHLFuBXNf35NaX6Y/MEimQS6w
NWq2SQCu4ZL8l/ZGf7FsGT0lOKnjsqMkKPyz4fwgZma4HlBRGvoWe/mZg7qbktreMRluJRFA0mNx
1VafBtkpLSg79hFd9dsef4aDy6RcQR4v8LURP+INEDpvTu90vuXhw71Wkf6eQE5jaiXlIjHxYhQ8
YczTuE8jV24ytgBe5mzj4fNwyUXCjpUcDmcNrD3d0Hi+/+G79kz35+/hdghH5xwbBIdNbH2nih3H
P0umbwko9rfgzap164uPx+kNdSFDSXtpEU0mGpkc/H2PkprusdjDdepUvjdoYBnkk8vzZyJeTAnh
l2X3QN2xHiVsBFGqLjnX51SWarMRrKy+90ksGn6MkykfjvWYviScOlapoBThI/wjUwCLt8J53gh9
kldTz1HRiiPBVs5m/BiMLzsuK0t7Hri+4dkXdLSr9/flscqQTgldWWxjYCy/SWiyrlovHrcjDJDX
Tykuwjlm4A1QajojK0RvxQuIZ61vw8F4eWxbtwPGolXGFCmVxDU67157HoY5jHaZ81RUbqo5NU5r
FrA6nWLyxEN3mJsnAJgOqbL5sHmtUYrDxCBbBl8ht4L7YQomkS7fJCopit6Ji7RsFllcvwDdQx7F
QSyb301saMQ6opfQIzoS3BFsRwFcV5W3juFYb4K8Z1Kx1Nr8ZtmohBQRHIllNk9xP1jNg3Aelq4B
jYXMQnp2bWgFfD1oXf++RZqn3hk1nH+dD6YePalc/k9hOASFuaHxHqhZmzEv8ff4i0d7jb68ZeB+
KK9Kyk/dVgY0af5Eo89vXfQXs4xxczdayPpBoRne2aGAJQpeGLdW7JQde0tudLAbxrNFywMgb2jQ
rDPO4eGX+ig9M6pohIIb0gZxo0Fvun6ZYoYvgRX5FpGnwacGmldqt/oqnfUUnhGHZLizD6WWIUXe
qsTW+spl0Dr7KVOrvXgQIyAMR0ZPL8zC6NeZ12E7xZCmU1HbI/+DkpnKWbEBTdVCYqASEHuLAV19
i+HAJnNITqs0rtIKYQY/1BZRwNEn2qFC7M3W3CvG2z4zwYRLwWzSNOHeIMuE6oqKAmzttVMBY8EI
TtqBUwz3TJpb5PIN4yn04a7D5bqYoqLL53p5HYA7j/4X9KkeLRK8b7MHbHlGwNRirHN9/9z+e6lw
ctlJBaSBPemEnOCytllWCWOo8htE7SGIIpydZR3naQptxG47QWPeqcAGVyszBpfaJpIYaNpY6oTo
ljxPXxrnRy9kyxpF7DfGsVUUC16mTp7ZPqoqPzCUlo9rFGdU4E6jU6KrHlnUUmvIUYCMNr4uKfEu
PQfemvWgXdJmppPCoCWhzEhdyvSHqnnDzx46u2nHU9eSNmqORHi7EXmot+B3WVbcAXRw4Cnz5g5j
fdXoHKJHpQFOqufzqZPCdOlFlyhdkObXSe/h2VuoPgKqlg0wEWwkte3EQXoOEr+0doNgQbpi9H/N
1RAml/Qf3G9grOTRExPygj57S7TXsDNYiYZxg24gvFVv6Q3xJniHHtYyCtrClT2A4QyM6V7aTnCy
AbD8n9TSatDc1lKnD1OMLZ4f7dH1OGDQ6sREm5d8gvej8qpB3bKPc+hDaTU1Ru3nf/jfcrD7AGpW
89sc0evGq+yWgY5yTbFFTcK9uJSH3xy69oxF/G/5YadjGGMzXNY8MTIBRVCFtCUV5ThEgoNdKi67
AzfwG1iXy2/bgegaBm+WFOlO6Oq12SKks8SUPM+mCrucwn1TFl9Bq6fSJbmYfqXhP51VZe2GF5NX
ZxhQ7R9mejE89RS4LmLZMqKGlxKBSJB32nUzNstaNpl6yzcExp+npC59KLliVOiJpihMrQ+plbx7
ljoX17qrfKs2VK+oKxZWOzDRRqsyjhphGh9hZiw5dsCGQ6/uQMVr/ns2ZRGhQcw5ka9w0JSPeqDB
ATbEPrUCUab0SjUtmpY/n/fUH229yKD9dZE1Z8x+okj23ukiZPbKW+hLUDhQSCFXs9Y+hKMovHFa
Fk7EUJ7JcrbkgfdZGB34CZkA3xRzmf9qaSt5YVPxBgqO6dTP+kCoo0J8OX7azR/phnIA7r2bND8K
j/KhYg6FsaHClBxDtMJQbdWeUvZop81NA+bx0ox/8V3hDLxAR79iE3FTMYakxAUMEpIZbevn4QRa
6kU1RH1FjyGQGxSuC/O32DxNopzViwQwG6GJEaGjSQLu4aaQLFhLmWFNvDTfyoZyJQGS7NbC2QFG
YIZhhqXaZbU9SpDAc6apWY1bLIU3sybsJmJHTwr++li18LK0NvgTSMj0R+ASiCxAGB1Gqh6t7ete
yhgwsiAzm06DMIayyUfNYvVaNHaD8IgdDtiUCCIivhViHP1fczUvXk9kZJHznLITDweG3QeHT+ZG
TVSE6MBNDKKjT67nu3/AjvmBqXC+IyOLN0IzTWAtcZMcD9hOLhV7clkBVRXB7vwqdklc/olTwIfZ
UjwZkLgyhJ02ogG0HKENHtWmmg0Mu8Y5T8nzjzNJt0LpeXsFa0KKvu7qHHhAyTzMSerXtCfkR9D1
yDhNDesAZSN67KrV60zeGS3zcfiE/ARnIGI4edcpvt1xGNAOkLcKZntiq2At91bEhFwZK8hrm0o+
c8Rinmi2EPu/Ezz9HfT7yqo+q3QunsS4dFiP8kN4VxutNvhGzSnmsWxyLjGvTsaP5DEMeoi+exW0
6tt50st+Yrsxj69khaJOSNQ0WIV/v8GFb7bsWfM5UQPh3G/z7qSKPh4hj0ADT6j6KbZYGHF8Hc7S
7/Hx8H3CpzxhPqF5rNWFARY2t23jZJbjNBYxaFsR6wFlQCU9kLlIlZUHfk5trKcTS+UKkYaSVWme
wrSQan/hrMe6kEQdZJq8tml7FMks0AFrxVrt7BmwrI3cbFEsw5h0/AwTFOvfMVmUrNDGNQLqMcHt
3w74TsqyoBBs6HvgX1fMvhUhRSSDiYzW5/1rIGHyw4hBd/lcanLJqP5KASD18szIoHVgEtyA2Syq
54mInOliNykKK1+ecSiGe3ia7ti+qK4wtHvsSWtVJQ3xTHfVn0fblwlYFQz/I0kYreg9RTDgWrvz
wqgrN/fo1VeKrv/IoXD3mC96ftlE3C6UfohhvJaSdZEEpaGjmOniuwrz7B4OM2ERgSBmCaFK7b37
DkNcgdpVNwgg6ka7HQaJdp4ovecnSyrdZwLJN9WyTMr7lTAFRzChMfO4Xa5Yf1yZOi0eNPLyTWIl
05ptLXcSSYBm03q8pCYHU1oIpGQLMvh+DCjhYgkklNgNmLi3khzn/euiDT+LkEHPf16DD3UGk1pw
3Y5BoGUO/3mcsYIo8FeinKTp+EKrux7LdsjUuFNOsVa11VHFkaXAqPfIOgPZOOJxIe2D92v2IHFy
FnIwp/lqXQ+dY5eAc2ZwF4jyRw6srkcfqh/Rlx28gKARnjfzPjdkHEKvlitr3jx6W9a054BF9QPx
h/PdkqIMd0KFA6XgnRcJMC09qx/pBredv+oaVUCXggn6pIkz4fJxrJNpid/CBhItphaqCE1dC99d
3Hm8Fsz37t9EjNDx2hrpn+0N7FnWRF+lXc5PTc3ynfOmhK7XUh+MfBR94Qh0zTpaRgHnXgIgdrca
7zCV6FnSg6aG8mtjYFuB/yrhPLhjk1MiVzGlZzCvOWoBughcpww5Q15EjFfgu+iWxgGVvh2vb6qa
FZRtYB0bHD95su6aUVFI8JA83tWuL1tmCC2z2TeqZRbHWCOe35NcgPhyhuNv8pLo3iWMg/KboY0r
6wj0QK7NCVYXpdB6QyhjkAys0M6dOwnAu6EHVUoZ17x7rGsL3lH6TxSVE6q0UxqEw83sw0ncafdG
FhmW3NLEHH1wNsEQB2euisraL9z1FpYS1TDYLQpeegaJdngEZ+gxezspdYbgT0STRMp0tycuwc2p
Od0L4iS8NP03LoJ7q0TCBT/RG81sc0qIi2tOUlaRhYz0QqGIDp6rhute7e1pPiTuYoNAJpTIqMWP
n/coijOXnvnUcqlyjtjY0NkmPNlB+3jUUcVlW5h3bCkvMzuRr82wIyVpmgfwfwcOKAnpw7HkXlV5
7Ki9/AAz7XryEMAZRDXJqVQ0cRg0blKy+johb44izWALUnhZrbkwcDqCsOvQDQTR/u8HIlFaJEzS
WLR06mshQ3xFzboQ7lMpDkbP95gId++I3l8hSLr66RJ6vrO6TT8NPNWfQzHdbW2nUo6j1XGC192Z
zFEzB8CUGFDgRvvX+J14rBulCPLkyfzXaG5NYS6P76jNP5G8ibjxymneoouvnBjg9zlDT8K5iD4s
Yy6JvffZnVjl0c8BkMt4raYnXg7zltDEXU1T9xLN91TZ9MGOoqTmL0kJA9AfliN693CnkepUNZU6
sHB7frBlbwJtWsU9Wg/JbyY3FyNG28gKZotMx5Yt8yD2CXiaV4lzsyJMboKKMQNit7wkyvPZrCYB
o70kgK3P8yii5IiI80mFAJcWIJMOhJCohiN/MIZxevMxMc8mwf4nb6mkMRpxGIh+yhDvcyDcAJwM
+ReU7jZohw1jmKoYJCwE1bgc6DYrfSZ7MQ6zPecfRTyc0CNj7DEvPYANuQHeOuQdqskK9ROqv3/z
dWr3qrBxyNAHyaP4Y6sgRB+B/TXdOlqHoUMSiKsFZtmgcH2DlO1rkUu2zQHaVRCB7/KhtYGv1lpU
GvO/ehaKWyc6ZQ9T03r8sNAvlS74OaOa+v7igjzhu44xAMxZt2Fa2/iB6/QSaNyGLLr8ij0nI6lZ
WmQaL3CncE2ZTKCiHxjTbd7I/ztLSKz7S5RUhVoeyZ4QwodrcYwIkRorjJCiKI5WeqSZz8GI1iIT
elj0yw45JGwrv+VwzF2AgXfOFuljScB2JL4po6DgdrRPRDcVSGEvR5gNcdYuWH4mQ2brQkFjHJic
jDuQzhQVxKdguLBSgllOveXjaFPdLMJaxxa0FGar/UB3XPBzj5t9w2qi7uDhA3TnLI6E100+8FMl
/ACR9ePTWUpBczly8E1PjT7YJpOm+fXyNCcilRbtSlyxrVN5lgGWt1dgd32oKePbqfhe0/ncdJOA
4xPPMpC+00XTHsNZrlJryaox+ys//xQVMoVlaS2zCpuSpY268f8xzWvu8RAxFDGYkuhu+z698zha
1giMFvuSTRZQD2r1PKkRYrrDMcAbvUIF/Ro2dM1b7xSKV49wCCXtTK5yzuBJK/tV3THLRMiZKpz4
JbcnJbMqiUdcCy4pWMy38dMCOCY/FRd+pL3m05KNTrKYiwTwm5h/EWC+ONxu06TOMT6WTFUtPYIm
SaEWEoaYTcHBmqp7HZV8IbKimSRUBozb0jkbLtjvTP6hdOX1+Jp1DwOKK5z+uXzv+lCGhE3xSP7+
cFWukNreFleHgacPz1LsA4+0X1CmxuOHOc5n1JXXQLdK8WM7dy1/F5PLR89HubDQC4S44vyTkEti
pz7QJVC6AkWvCLn2Z7QQE7NCNQqCSeKr8K+BD1i3ubmHMoED5+p2bVLUgMpNJp8n6ZS2aY+Y4L5G
bhw7FRNxIxbaZlLopvm2mzNKey7OstRIIgM52fXTdwYAHPI3Sbc2MffQ9cSQKfWTuoNfVOACW1iy
WguEYWTCCj5/8tjdTJSLkgpoRb+d1+CA83OIVy+j8NQUbMRTWLnq5L9y0w57Cf4qYRpRBUK7w4O5
tZ/IhklOqqsdIhZLbDAhGpqA2Kqy+3ioIks9Eaij0YphRC/56rMtrEO7Fy2f8bVzd0/rwuGOhHSG
JYrsZBdkuH+X5nZsnsjYKwZHHg1kzn2r1iPl0IUx9gkefSHwIiezSUXNcaAixu9xK/FrA9H09j38
0Krape1TprqQkfItizI8tPP76R86tiJP/G/Qq9VyEhdISCpmGtVGibNw6kpJVYEkhkwYTgidZAH9
IrNSTc3HMm/fEm0KV/y0I/OEjhpTR9PXz0S8o2DbTXvHqz7l1fxnNg7ASQ9guYJHpvIwUMkR8v8+
NPwmjxFZi9WD2TLEkPqITExBjtXDw8UjmoQyUZ+JMNMMPcO3NXgmVn660q9uIFrxFYfN8SBnqbeS
8iKY/G+VYFajTfb1XSw1lqSnxkJHCafBCidGwrC1Sm7EwuCzWirU1Ef1I8kio5UEYALwJdi5WHs+
bY5fG4VoKV+K0Kyv4LN8m7PHKEZ7W6boFZIQfLafvkZH5h1KZe0yYBQJKLKGKpOEozNRgjCOM1o2
OaU8WlpcLEGZHk5zaCfjDbfhr6xSGD++WJMhZPs3TwRM68PtT4bOJnOfgkGXT0sulERz8Z03lTkX
h2+o2Bx719RuC8tg7zfBXfYZO756C7jRZ91Jl2SiQ9/1jLJEgGiZp9b27R7DCCIFxtLl6PDnBqa/
obyFR+pHad1uUvVdTZJE/MqWXbGEcjZHlOfTW1LtqlV01f8TW1wVjbpfnmcwz5BeQrF3c6SXBSzB
Y1ORs+qryb/rSxjm9WwPykX1/UBh7LQDPEVTdaD8MKl3yDtXDFxkHoq8hy/EPlrIKnmkqiIOzvIC
RdjRWExtrEZimZVzYvmmcXLcDcbBY1wsiEGbl7zTipp79dox+pWAk0XIn2LRI7I+nJemzo/H+dVR
H1Ge/6x4kkKg/kUmxEZlhw1nrwNdnB0hnxneFAbHNipZiqMYuKogc5H9zNRiqOjaBqTdFDtMKp1E
LnM9Hc5Iz+cF4kc8Q6qUIlJKDB57JpN13bb2yDAMAXS6UlPlxZjlQTJtJg5GskUpGp8piFBBe73i
KYi+PMb9zMPsP+sqd6BWhI/5Ls78NDrT2vVYsiug0PRMXcNz5fb588PXcyo6Y5MPHrL7I3g8ai4t
sqTMlaRTJW+YUfQpmexydtDnEjLGR2jrbZ0Ykh/y4ktoLmDPkFrPyRJY1GBF/ZZAf/jhdy3gtKxl
yEzivyY8reYBDPsgVRWiZNC6UWbX4nbdEUKIPEgM6x05lcxihZaEbmzM0OjI3ajuXM3rYZmPscpn
CPSVY7Czi+5MVJXhvkK/1xyIDkY3cG7A5arY/RdUkfjmQDGRb51fsAutKQZ2jP2quQHygyLAY7IY
3VXalvQdtjt/qbPBQWdyn7Y2R7Ht3hdJ/hFAudDZGbnAZ6BwzD/ut4iuCvbCcg1qc/d/Vb7XzSL5
6UJb0gjmweoYUhgPDew+wXU1CCIBd9Z/7SftKs8u6tWWBtUVhAuDqdouzqUPUvB1OJp/eUWNhhjI
bCYjakhDKWTiIZm6iYfbI194ktEbOTqawdDxlZQHSBvmFLgpRqS2C1wanOHrv8ER+wXC6j+V63kA
6/Ihx4ApkAm8XpAWRD3dlRkKuZ57wCx0f+oYZBfgzipBsTdlu6nAb/ljZxJ+TWnAMZ0KY3GPUjyF
/7Z9WldKY+UChnnadN7NsOgsl8QH7590kdtOEDzwbl4gKnFZfW7eznIGQpq+BMD83zJw064wWdwR
RRwaDEzSMgyqLq8aRoGbMv7P3jP8t6FQ3XhGhdniIT9y9HxXK0X7+3CRR0uUEhap/6ZieI9cwk6n
WugLnkpjklf91HZTZw723HjzKL4jFVJz10ufudbj+hR4DrKFCR08nvGRxsekxvHdBZfHqikYR/D5
kLky04rOdrEeXeBPLQnkVSor9L/r+vq8gfbYdxmEPrEpzhePgZ/e3MQcXovoO3QuMou9yn6NzPQ1
llJjTLimw80ozOIxHPFuJHQh6QzFcQhjOupxNqLc6IrAqJnO0x/XrmGCXntxY35Rjd70dkyozJGM
ViXGBOgG9OSXaYwoSExFNNXsPZ1c48HCab1jYS5GiVmGQKCO8E+5DwNwHf8+xrZ8a5R4T9NLHmXt
V59NyV+49Ju3o6+LYXFcmcUBuSN0hfa0wNnWqEX0a5rQBIO9DXDUeEf0IUKbW4IAW4kjl3N8dkPy
iG/MEUmt3EBy0VY5nnwB10kFjhbHnRKT4AmSKHSYB0fzMrJCAzI4Pz2Sk1tWKJhHFZXmNid3oQkN
u69tbSpX/lqcR8kE7vyeHBtaC2hq+3CKhd/H8TK7YpBxtrl/h0cdMQNzrM4EJKy045uHdpERxN8M
+D86Inzu32+BvCe5T7MmmOhPljVy7eb67aX4FhLDtTGy1R96easAniE24XD4gLhzmp2c79FrB0qa
Zy0P7HbPTyX+HlAX8Aw4slxXJM13az3h46psnwnTqs4l6G5hqwOWuvoKhPPEcC7sMiP6fhTVudjj
qx7PQchtyRSs60XdctviE6ONNCfmcI9b2jhZdeUAVoieBVTwCmuE6n08+S5qKrsfaYx9Pqr43gSx
6xYTpEWxKVQeCeUENHcdtWoJ/EGS75MJegztYhVN/5jWFu3M6Mre8tTma97cKUSVzBLcKF1+FYQ1
JoRuZVt2D6VI7pLkvq9YMuFPAZRs/DLmA+cAiXT8mPk6Gs8o/hLdTPFs4g25o4qCzFNYwr38Gu8/
/kYA12/2NshHz2Rr0r/r0Y+0LtJPXRV4jQwSPpew4kqclquMKYhdyjckcG2igYdiNRZTclO3aDHS
yFKMIxLZhH+LUDMOntmNbF2UnRDjKookXwvkipUpMxRE4I413VgCXiLw2nTuly5Yn/T28ygbmBbU
FwWv66lws06IUh6sjgYicmvLiL1VsF4U1JvX9jaqU9IetxXvKCzx6plK2UY4Kt7j8cbPpD4gZz4s
GkyMpDTD3tIoIqM9WkK6kf/5p2+M31ihzIDecxYlAZo/AhParxho1q0R4naqulCau2lMtZ/nr7JW
w9G4DrqleP5w3W68Fxz83q9bHaOyNXBMBnKdAK98h7+LbozqX5OByjfSUepQOcug+FUWJyfIJZ8C
cXlgrHI6ZjAjVb74Vd82kj13SBh/kVnj9/DNzpXSbtxcJuEBMP2sQPm9wrjGAuYM2SHwE+OWotua
TsPbtXY6AbXvEiv2f77uWL25P7LXck9FUS8pqS1cz7DAof5j0/SD0+yLXPp1nT1Av3nq7VGkLGb4
J9Iooba0omw3n7xfORZEMFHuINIGatEkmk2Ek4jUYr921PeREVB6WsS1SgRnsQpVdVah8v5Ww9Fg
484mt9KCkrMPmPcEHSXhmYiJz/874hIdfq/JKJAWCvsfBsqNpG9d2250g5rqeAyUO++9cem1xqDS
wy6PlHYDW5BvnMoGg5CajSz09uru/6O5Iy4rFwS0ipuDcD61xAdRy5R/pjZWvAXQ8ZW2WQXWSvUp
fR4peEDxW4tX6yJrBzZLYQvOvGr9XW1+jD57P5sww/f1UgMGL6aMzAyq0ni4abqDIgtx+Q32ZnD2
+UMVo95+lVKx7FeHCGsGLNHMbg/vm41WII4J20X4br3YbaQvXBpsuEjxn/ZKQITDlRM+wB76Ku+d
Bq1QbAw056AZ3G7YHu3VF8lVMJIEIpJBKRhYO6x+O9dRMLOVqR7RC9zmtJSwv6KUv4fYW85MlKDX
OEmzF/Q8odfefpXcNQdYhZTUlhITn34bmX0wL/vElMIs9W5GwctjeTzdRVZ+qeVxRuVaQPLAhalY
9uR85sGUBI1ZYFobttjej1t976x2Qqe2qZqyIgwzopo4vUkVxl0zosAp012nEoDyvznci1tCFo2O
Q7icvT7wozss9vi7SKWxrGKoV15xvPfuq6r/sbDrvfdG3AsvOWUJ1b76TUodN5gdrpE64lC/yIwS
9QF8ayhtJ7F4v5JcIiMo5TZ7AAHKBLdiwdF5U9WchSywttaoAqjBnQHRGvmgucWwVdUDZbrTY5Ql
dkP++8tK45Fedt3xDH8NnHmPohIMuMaB5QMP9Ydc8XwOgPzPCKmG+OpOGG73F5/1SPbHjesBXVK6
S5Co9qtjQNX92mD+f7TfemslwXWni3C7NkLxOLG0uiGdT0TLNQwq+7jowuEnxj1OH6oQpAHYdVbp
+axwLDGmCTdUlM+w01SuU+3V3bI1uICdKO4HNq4zvRIs4zDhb9iMOo464TjT2UmPw2bKdbLUnG57
1idnlTbbBkVSpRL43x0LkxmFB8pKBYSsrgZDi4/KFzVT7G+vWCA81+hAspt8woNPftD7/8FLhZAT
fVTk/vAxtjzjhJDYL6BuLMnCm/oZPOlsOtX6CLmC9r1xZUbWBlhA75B2Ng8EC/+m0Pu48mpPSzHD
vbLDRf9sCla68BUZtzGeOz4Tx8994cwBLJWP54Rkz8VtsZBnP0AtRlUnitJBLpnbl04DzDeijF3S
jskfMM9DW1hcc+noCHdzpbnOX5ilqqp+yqstZeqWoTNImpWqvp4M46RR2mxEvJGXQdo2DrWmORiR
NlcPQJsePb5tHCzIW9EYKyuWhoPsIHByfMvMh/GnF6jxLzdJ2Drxcu5MIXhUc+UvTHdtv0euyx2J
+7BFPXcrajIyfgLtU3pNM96VZClTEVsFKb4HpCNaz/vxl4mTH3s7dN7EGRzu+avVRYiTcuCxlr5F
nY9jzrQ+X/palzsRNcxsKux+aQc0cScPFpcBQx+eGvhpnegn1YElE5KCzrsBVoNqIeE5vlBEorWs
Z2PbHAB+XpwmJwQxQLJpA5WaO3CmEriMZBJ4UKa0gjrb2DpPZUmG2dBH0ch+MVXImWv/Ewe3pm6w
CLqaqIdZyxCHJeYDlYLHTJfvNUJL+79QOpPmgVZRsnSdiYlpbFPUJ7yFFEZ3TQLV4OA9aS0pIXIV
o0qOxAjGih7bB3+D+UhiS/rbZgrlIexrtffdH212sf2cePhtLyR6EplgBGsTvsoU5jHjlYTwwgLi
+uaJceM9m4XVScwp/8TKcMPcsBCQHHDu+g/orZ3HTw9/QOdrKrBQLd4LnNn0+YrKn3Is0jyNhEHt
FkStBAgzVMq6A+QnHUiffa2Gzu1AfdLLCw5mibGXa/bJH0lfcefiT3PxBksx4sP/3XwL0fC1Emkn
Y7MQ3UBnAwQXCCrNJeTTsQxUElamp4IkA3p5RpTkiZBva9RB873dqsefP5NrJ2hxZ+VAb52o7Q1B
WeVsv8re/GuXLptGCOL+KZ+KSHcWTvRLqn/W3b5OsTg1aVvQVmRe+yx0qUjkCh6Sb51vkLQWKfcK
9KaJM+2cqai6QMGLXzrqVxGvYIp1Ax1sSJ5JXOolfi4Fm5vYFmz3e3CJvdIRDdB5ZIi2jUkx05ux
LJn8epVXbqu1u3lKvuRmsbbtt0aiWNd/4yVO7BPnTfDJ6TnOPQk1CQbgONHhCwlLFqCUTSRRukmU
nADiqdgxh/pAZp6Pm79mWJz31YXmoWo9PrFrd+gJ3V8CMpywcelpuTtMyQTMCVcsu9rjw+Fc/AY5
fuMHk+xFVrHUci1g9r70m6eKMJ9ixglYsq6s5FlvhH9MHU6+/sJC+OFQ8OCwh06gyT5p8Q551oiE
1mi+NHC6L9w6yW2KKA8Vq1e8dGFSubirBFsf9xzRdjgEQQFU3WNh/d0ZYZQEKSn/DEd/e1a6PAmy
26luxlzB/IVfYlFY1NyMR3iDu9EFsRdyoz6Jglggy6uGq7PjEOwc+F8ptB6rpSSlOFB9EwY2FMu4
3BAWRMPRYii128vPzr2kZc94OhB1877A9h8ULM+QL1dAFC9La/fbaGwYyFsckQNZX2ZxCYCAFdJC
wiQa+lKHJuyIOVtOffn2kut98vekkhWzuRW3r0SO5RSnwAZbjwb6ntWV9707WKTI5R+Vz66nsyaO
Dhrvi4nOEINKlNnqPFthSirR+G7OyTsw7sCGLtBM45bCYtWyFOciRR7hc0GlIlTPYrcrZz7sx+Cy
wZVYCzrl7RXoG75QTcSwLR6Css1Hx57jdSIiRtLjDtGjHTMRI2WMosk8AkLiKYp7C4JFxQBVTD0h
oBkhgFJsH9kp4N8mfUGtoDwjfrvMSZrmyfK4k5hlGSi6pm+h40Z1uBdwUiS977cbgZyMuXmC9cVH
J8F8HSFs11gEdSJX9ugwbgMcVi1NXY0/fl6xiADPKDoVtlQwrplz8sak0qj3i2RlE/YAPcV3crt8
HUsHFCudHG+PGA0Wt0EVMr+dWPv1Vfx5obHT9PHd8lwu3Xsi6gfpX1G4hXFsizUNJilyLYfHax8m
qAjZ5AOak/m+DbStQ3gPhB544gOxnOCjnv6u9K+Z4A9RJJ0XWTXdnuI/NFgyQ+nwPCLB1+YangBh
3XdKx0hgkap/D6WMptnftUTFgE7iemudkujxkTAAlTZRapr2kyydsWvEDR4548rn2/ATM9uiVs14
F6SPrQaEGD+aeLU7C1/8eTZt25UJJMVmVZIiU9I9Y/VE7iP3YNsjIN/SUZNhXaCwMRg7IUxZj4H3
ecRP2yiUCKNUvsqGgPL4z5u5J+KBBFhafDSszWOrRDHqsV7DF7p/JSbACorzkZre2aVr9xMvXqkS
UIBCsP3OHxtTN2bPh8t/R6LZ5FcfA426oLpbkPLurREcrrd7MCmtJPnRTy9GlOYT4Los6amxKdFA
2vBd/AgRqtvfEnmnmD+xyGLo0f975iFu8jE01KC4F2hiVipy5kSNetAqQP1CL7oEaRh3DAhNJ9lQ
DerrgtL/13winwpS5CXb/HeyMpBOl974PRjHVSGHasZn+3VKJEByz7sycPu0ll3B4KFxlKiwlhxY
AlxD2RgYOb4OFJYFJMrZN4Au77OaQRihHnIFeYB6o2Ycx7mrS8hHHuVuT5XpiTgbwUTsYDARF/to
lrfDAZpJJRyYg70kIScR+n97mX31RjyQ6vwpyl2zhdJH5ni8eGDBLkVAbyla2BYS8WWpAnaiyeRI
tCpphrEBCkZLMYalYmikQrDxYgHF79wRGWTKvJD3gH0qAVlFE+aB944kmxHlEz2lAOuOM8tZNe5a
VG9nzW/dE6Muna6a2MSh3y+07qKrtTUPWqTOlhax1pMJtfD5/8XCsXHhjDJ421oGSEPu2vJalk2V
sGYkeM1jMqmUUMYsiJzKSJZChsBqz144hfsrJeWxqBv18BfwfS0QMQv6Xc5Hre4fho60e519q44+
lDC4dEWj8CgNbwsq+YgNgHTlPAwdxiPaZbj6RlhN24mj0MbUMiZOIR++V5ooIEUMrbexlOfqp8Px
wv4LOhB76nqDg9CCjtrfdR1o1sqUWOOqfn/3aKiVo7luOxWn+qfk1zGV2rZYUlZcUIdHQqFQPyjB
k0nAEBxlEckFqaZU6i8Q8hGuS/TKEjvnKIi/n3xJkZAQpiXT9xwAOwpWY0RDPz3vsNP9+U70E0ZI
BCAV5FFsOk4wMpXas+aJMf8YMdZpZMQ9IvKNTEfwpWKSyqp3nrZMJ/iDeNzd9In4eBbB8+s35MbV
jAeSYOmqLR8SfOdxGsRwLWBwI8LFsdcc2o/fvKPYEf7LheetLwlg7e842cFaOxxq6rSyyhII4pYf
oWMkpHPAUWiqGwmKWUqPBfDc4lA0+TpA9ddnbAg2qG7Bl1WKSXrqjdvBYKZ19tD/qc4JZ4fX8vwD
iPD+1/xOVOsdQtqaa6JWPaUcnnmtOyJgRYHEUCUqNwuIzf36iTmTgcHxrMmI6ZYDQQYgKcyJyQau
FGIU+bVIKKpZlMtK/fcFW+f75fAzqdxzy2mgPkKVo+NsfFExpbaSA0kvkFe3pSvDA4resOmCfZRg
XIirdUXw1Nlu4aGz5qk7jTsAYEKBpjnsYf8sT3AAmUGG37N2A8IwY+ZIdaE67NV00WRt1JhzaWrA
uswntgpF8xwjZGq4roZFMZ8yvcS1pIsKQNP5U4Xcc0U3EqpV81bdsCblTDqCYTIjMpM+lrq3x7bv
ZV0exsjuCwGAPE+ljF/Vo1WOwMAuOxq/EcCHTrN+YzfVEf8c9W6xczp8AcLbtKtECwQAbLq/Ei3i
yTm5zaaXiM9896YAbA72vDFGa+jbdyLBUgsjhdF1OtvAEW7W/mUS7gxrf3OXALBk7uMdU9nf+BM1
ZL98dxvsn7w0ScQL4zKZ9fLNmKeFs5iCQiYNMjjySYMA6jAbz5e797eWjPcKqzYXJeTLfkGEIME9
uPNEdr6aazqs1rTgYtAy+92QHdYs2bV7fmtPV1M3XhuNUsUsEywnT3yBFNAbnQ3ArNFq/pk3g78r
NoQmrs79hmnYbfWi8LSmvPcCxY+gkLvkM81YG3dL77s4TjuSUmvdcRMFwn3Gk4rRWMV4thCrgVyF
SQiBb52m3SrbZkTfrSqzWANo49UUUagHNYmm9qGqPOdZWkVw8eaS7wVOZun2lKDrOM9t2HqNZC1b
R9McqK8+SWIFZbBti9V2xKW1FTMEnSe6KRfv/VwY2r4Bld7GXiBKKiL75rC6voni9nos9qDs2UpW
0MFgdISoGW83dNul1K/dkc9xSD+e2SWMaCTaby7YF6CMM4krTS0TpaSck3RerspR9opmZJS3+uu5
J94IwlFfsN0vXGW/HtN4hiiX5JfxvweHUWUpbEILx1Zsp5iGdQ9Fs/oPClJ8MfRY9NEE4UfSaSfv
z9IezfFsv10hw/C1zAyFZJroKcJdhnuSoe3PPR66+brL7M+YTwJzSuFuxQESczR9St01bFD4Echn
/4E6NtWP/+NLBhjtjhOqURkZLLL6LnIJpfjotqugkVHmiV7eAUqq8HSP0fDKh7r0aWwo0jHrQaNP
DXTL/AfmkTcs65gkJ6IhiEqkUJq2rMMsGBoIe22eRSFo9aCnIbPhGsYCfVTVDueABkE6zJ7fSIYA
mtuqlH4zzoFn2mDmzhbv45e5p3tpC5/td893B4jontIZDOjSuM65EbhJYXGV1irgRmqkf161mwnJ
RtDbM8AFbeiVTOrR6qsTFEllGDI9et7Sc5XCt7xcMAZAXU9k55s6Q8oYK9/Co/i9hgiUu9EPCYn2
AW7Dp7bILKVt3kirTypHMNq/ifZyVDMGBrk8wlpfDKyIWOh0sQKK5BhBRKmpbdeqQXuv13L/IjW7
LTkyDnDEhtWvRxUASxjNjl/nCnU7bTlwOErURlOh+vmQC+UuUjm4GougnO1qWrFu1qDxAn42NKrL
4sf8MOEn/HWsR+daAJKCyyL6rydTIj7NndNu8hZODGp4Yg4LQ79CmbCRFq9qwtxqcPy+QUEpVf17
NMuvzmbfdFLGMIwGip2qp6eBSEy+JsjP7g40+41ySJtueeeeXwKiLqsCWfyXbssuuz1fM3cnAJ0q
WT8Nv3fScIz+TVn3hZQwfYkwPa0ci36z5BnyGlPvqMRsLX0u5t4lBK8lDrN6MG5KookHG47atdaQ
Mzan9VEC7LYS4HQxsmsdx/hf/ewShSGjtbfmSGBgnBHQNqtQFpI79iun7XAjl+bGejXrz91yOPW+
sAhRxxYMJJrqdRLlqa2Dyh6rOIm0x2IRgM0x5+UZvDsRXsurD9BGbMcaHagV/Y2ZUtIftfSRZ3UJ
fnperjVEpEq+k9dcqK5GaipqLD0uFMRTcPj5+HqNDiEps2tf2ahh/JhY7oNd6TL6hNwbXV6ZI5qY
MsioGz4mf+Q8sPzDhgsoWeA9OQG9kPvtmLpRx3oG94mc7ZpP4BI4SzSzyf4wAZqHiiM753yjSBq3
MlFX6DnHtyvXnQx8SUAKoAVzBu8Md4dvvmFcLKKKr2vfk2hjVdYhqXH+nbMhd3IdzJ5CEkG2A0B8
NXULo0w0PAcO48IHsYX3gUkNcETYEGTg+r8MfSqWBflZ0DGP6gSH+Ex6jeul2hpU4dIJBVnBQldO
DEnW8b0nW0rOjhoD+lRw5cU/HP36UNEIwpnTCvywZJXKi5yvyt3ZlqStsFMoBpgzT9PdnBQGyQrq
i1MlyMbGRW/VOFCEwhukIDpDhIYuf5ohu/LGSz4m0IiTdfZ8JovCgAh8n7iXXxJVFPiAbPDhDXb0
7/LJ0Cdht9mcQfvML0qwgy6ssTPtw1uUQCDzMsmUbtWK7CVlRa/45zI0f5pwJXIIKCmSz/jvB8tC
3PEyHX1+4AINHrsNaDTJOIHQ1VvySzt4HcaB0MFXxmGjRkzGL0O847d5SJXI4h0LUYtsbIgzbQ8m
v3cNOIOd6rl06jk0tMil0e26THwMm0TsQkj7L9MHO8mkgvY5kqPqCFVaZ1PVDHJXPAXRw7rCPk8N
BY93jBkGPxlyUdUwrVeRa5vuofIHjDDJgYvDoSiINTf+QW6bR3BWRWlfKrBPHmCSPa92U1qsxNF6
Pws2tFAJFYgvRNbKxzb837D8IpAWutcuEPeRsXnX0FtAOyt4HHpyyUSLDBy9zI1d74o2rpkJE26Y
uXXWQmsvcK2iOzjlBqVoZE1P0gX89F8CUDREvN0qr/r+BDyVAOniy7/lVTPkTntzm4u5XxOa1C4s
gEQEE2AF99TqqEo4xKuDyVMwWiNezn/yZktkDs9KbNkZxtTRwJ8b1OqC4NiXN7fDr2enBnOUMw/6
hb+QEnXWM8j/pLColKnYJyXXvyuzmuohU0PEv/+OdmPpNHKNgRndnyVlFnN7ty4NrscF7HLRtc10
baKB77LLlk2VluXCHo4FOW50V5Nyi4ZUic8eCUmrO/W8R0lOHFo8uMHAEMFuDHjoFD+9Il0YRB2Y
TYCsRt3oNlE+K5Mp0+NLb0iHE0L5TuqYgcKica7xCRhW8UJ3/QGf2tAlVh4G5gNhpQUxOmRt9pHz
EwqFVwaTCMpxtL1bkLRa1jjkE7Q2+x1RIsdWNaBvtC/mvnFWYtPaUUK8KrGuPCbuonp05l2JDr2h
UrvXBODrLpUzfwvX5CZpncQ6XRxh6dk0WEBzE8Gd3Ba0qw0ZQsJV31ElmGscChaRuVnTTM6T7Uph
z5nV8LqKH2PuPgDf+yDVaELv7qEwu+iMziPLF/VJjzlVF4syvjxMnfH1GDvW+L9wlA9o3anumk88
gXC7ND8mL4Ch261tex+wztOPowOUG9CAZkdyUvrnRrpBp77ScrEJnPw9UUMGuZZ9XKM3oRHQRXaH
u+uN1gWbsPn0ZVECh3T+Fh9wYhTIMTiA0j9JKluvSu+Sm2ogsqB65ify+wKzkj+1PtmrC4dSkjLE
YCl8FR8xStaIY0LURwGTvjNMdZR1ZYy7JWy1NYq2uVGEyuFK15cyGwRvUw4QDPeUzu6wx5f//ok9
d+IT+rsqSHThn2eMEmqUVloTYyiRw8DsuQtPtHpO5v05WBwTaF3w8WgOeU5d7rm9ll03trsRe10g
w2AaOUC5JFDsbekeckfK6XiSzkPEJ9WFtHo0QZ6gFH/JpN6+AAxGEl8yMjmbvKBtXa2/H51ObmJG
n+Uscv3GZZlVb1YkjICmyyMepXjh5L1gx2pKQpTOVo66amRfmeoTt7knN/7s4g0s+iaFUtT2Z/zU
9YIAUGiCn4wPa86M41x9G/Guuoo35IGHdkqAo0BAZCRRYgkh4XiUwIG3+yPdJUaBgjxrP2qnhQpt
9put/GdFjmzsx4g5idDRKmmKJVIM4F+JAyuqGO7ZLAoFM89gJTViJj4WET1asFggdeyF1D6E5PVi
qVpDQbhi2ufktc1BiaLL+que0yQKM5YXBZtIb0IZbp7eBcjaYKJBmSrmY0SElgJKqebnSjAjIA7b
KrnZvAZTEFitzqdaWII0h3Rgzd/rlzrc0U1cs8Qnc2IYTnyUlwIKLxHwKjfySJbHw3zl8Oig3j9M
Ck10zrb1cVpXECzPOX5nk2rb4KRUyVqbnNMZjIcUfEnbPn3Sq1+beG4xKuMO4DJGscuD2vLoLJ/k
7wudS+fVs2NE1LRD2SO5xNPZ3uJXa8kguHtFV67LTWFR6uri2JG53cNc5oLfxI/I2Yga328uMQcA
smV6G15uMaYGnRpKurah41m2HhxIUt5Iw/Q+LQsMRcUbSVIxuyJmgNUymP8HlSxnPOWToG4AxpE9
hxQj1OtKeqkSFdNmf9oj4o+y0aSj9SMnRM2LN9pUlFosnVcRQkfk3VN/inumk2JKuf2+cDAjwwAv
/ze3sN4g2xyipnmm6qPzcev+boqsVAU/XndLAu2P5F92zKWwrbWl9AhKrvts6wZHkrQ2QmBU1gnb
wxeP80sX1idDHAZboqSHmEplj8DWvyoH45gUvA/Y8q0iopO7yq8vstDzUrspEYRrgEwHPio9cmW2
taxbNTutRGNhNQCjYMOvXsJ0Fsv5Ck8oKxZGPt+TmROxUJhFwrf5ehhm6tmsrazojI0Nz4WFLosJ
is42IKiTxSZHIlJSPY/3zOAJkya208/nZFLnB//JdS+FOs/+eUb65VfMNA4fs9zV/YMQqU37lpb5
rquv+W1v67jnpjXtmBBtx8M584QR0CX6aVZ0jHWDkrgPo1rXTBP+SHJ9Glw0XO5VrB3UImMcRQkZ
xeOIMIwVty9uTwlVwY/kp4tMlyRUafZAHFpu2Acrj5lhAcS/nqwwe0CMyfAK81mZZXt5TzvmTJM3
fNROkyQyIMrw2HN/9R+EiB/Co9h+mVMqfLbkTLAF50KobCKDuICEnedNI1UGLpakZ6HcJrod9oJM
SpMOvwIp5phSCcxyQPKHz/tcLhDb1fU29gCT/Vt1YNzi6G2D0ASTCyyeakVTLNchCs1RBUNjG3i3
gVQKJg+qQDlYhBP1UV2Jf60J7tCxeB8MIYGhuCayGW+1w/Ruh6kMu+kqBz26UgCfB/629ZvjD8V7
0UE6oaKm/Xm3Yc7AmpuvoqZsnSYeaI0B5Sl5Tp18tiSJJ1cGry6sqUosPm+alDbsN9BM5FSsQFvy
SFTP/3u1s2YN3pugEw6JQuRqlsuBCUJo3Dyb4iuRcIBGCp4ui3lFSJhjogsUgHSbBIn6L/h1inLS
eKr9l9qSzo5FaCMJlpgI8CG//kWWMSPAwYIrtr4QRNH2cenEtTMWTZew8kn4z9H34GF0+bru0RBC
CwkSHQA5mI88Ty4EwYhC1M/a8ULRVX9atTm2zqy+w7n8fIRDkPN9ghCUxl3kvhnfaSEvBHuTHOiG
8JQlJjvklcKN9QmeN1C4Za4XyQDJu5362gKOGWEY8n0oM2XECwoGwfXdKMAsY+rqH4i/cpsCqx6r
1CZFSMwCIsbIZI5XDi2TywRdaiKvKdKDhTE2BNCbqVnXj8fqWYK/6JT2aPnWUF7moHnC5eIyRho1
vIMOqmzBENqzZpd0Mz0GMfm22Jjp3KmJ9uqs7obq69EcRHSqTLxL7zEColCxfsH0XyiA2tVPWRLn
C0b9kDZIUyKy9W/p8bea8neZtERmLvxUeH7QnF06GF1D6gCf2sj1ltKhKYfal/yG6xKWG9yLX+Sh
uscgt0/ez/2bL2mRw61gOuPl7u1lZ6X2vOhDvwvMlpNkuNLcnwmM6S+iOqWSyTiAUq+Xta/ayOvA
XawaMMhl4nzWf5htWE431VLN2XqGeGibPBmlsPplPKhspUBH3+CJmDkbhOfO4MC6x5TdsW5YIZ5+
fvNyhL6nP57vJvHwHDSXE5TgOZFGXSF8cW/v12fHlwWPkt/oKhySjQda9mvGQvZ5Xr0z2wCY+4gN
gNuDl34FOAukfXVwQCgOw/VOLm8BxjkPLGUQoIgBY47umSFsvGkx0EXqZ0JMthDpt53jDrBxxE8E
NtOUU79fMW7lqE79BQ7VsAZyB0gLLORVsSw7yDa5z8hblKekh1CavhjKm0CavFRNmjmBUKYJXgwA
bkIVLqXLz4WRB+Mcdt31jR9Z0QUfhCI/G80KW+pwlcEYEmRZr7k/GSVqEu21jsv6TCPtquvemxH6
pVlTx5UYZwgXbMtyln9q2Z231lBRzJp1anJNcx+boa5aKGrou8q4Ik7aOjJdeTt13j4Er9EYAs3f
vwNhLhTjWPqbqq0R0uyVkqg/K6TwFIGooOpd8jyyHh3wN77hCKh4ASDaMQ63IU5yFg4D9PtIOTue
Z7TIeMVVOL2TAdYCXM7wHivf6kmZHDpgHbBt2OuYro6vBScOWFZu9FdVwHBWQ/bFf6nK2dh0CUbc
yPnDTMSf/kot/WdnrtISUOXQ7Xtm/M69tmtr45+UcpT2U2J/k7bqQ7WUu9OE87U5dAxhrgFw2cu1
Y/p1MkLgQi3FC5xOnwlpbEytx8+bBvcrP/RJWDfistZyJAb04v9cLhbzWwx55x3065Z2/jhT//8S
Ol29884WnVzciBJm0rjiSns3aORGIFHNvVXtXK1JFZsvtmDVpI71B+frZ9XiudJym+0Z33aaec6M
OeD19kepfIRuMhMuLHr8RPx6g8SLHs9SPqZufPL1YhXsCHp9VztReHyJDILX8e2jf9Ix6RryCZf2
EkdwTbZcOYCFz6g5iMXCmOfj++ouORPfBSzECGeRqDv1LtYafcBsjmNJxJ8BRSyLwqDF9D3I9oR/
CFiYHR+XZjdzo9Ciwvzwah7Gj3rclMlhqTh3BOLZiDq6bl5d6DtcHA84tzuDEi5Adjt68ljsH5HW
e0RLK+FZXENQLsAwyBy5drQg08RqaEOfoSym1nnT4/twc7Hyl+BcoX4V4FYmPTJlwjImgM2EuMQB
/XCJxLu2w7zSH6Xe+uefNJDGrQ19QmS80Z4LWwRdhCXXyyShiNfX0ksn6pZMlbJuWtiTuyk3PJ0o
+zmoIhfHD5n8vdY4nyXLWmONBhcLhrbpDSwvKBuBZx2LwPT1FhGB3VT02GCt5D9IifNLmWBzpK2I
g/yS6wvR7wL+bl3xeIqTn4008/h9QoskXHJ6wwHjBz+/aIWHHFHPYl5ICBa66JwSv+z7ejT7tIuq
g1yEL9VOh06xBwbyLiscYEgo/HXF/QZLrZEpQVoyWJvDUAqepWXdOfAixa4e0KT7l3Ldnd9qAr1y
3gL0Sswx1T04/lgDcJKs5+idI9Ao1KOuJ2kRgtuO+PdfZNowd0GbmxnT5EbYObimepsc4fhTg9Ht
BR4kIneAPb93lOhV22XEVZgZFGvIEgusOjUmn2dQI6xwd9l0vaDk4qmuBlVey5Wt066+bYrejP6o
cqkFSdarUDAtXNOaM5HKCvF6+xB3E0R5vD3n4M11oVT5bqxZBHlt0f7ae1Wqu5SBWS95btUqk/rX
6W0lHPGwK0dbSptbQ6SziwYJCc1+HPNWVlswk2/lZC3d1erlAE0Q1OA7cTysLOud8/4vk0Vgkxru
sAoUjyKleI2Jl6MGH09YXFRc1QtN0sNCUfZTqiD9DBqHPEeylS4PUeAe5YAypJJciVliy7fqUmYW
8a5TrFi/JXmT5haD3kLgtmJET9SydNHvdsnFSXx0PSziXkRalyoJJ/o4JV0pbpnPuOtaGr0hfoDW
fokiO6R6hgzJegPKlZuNYWnrw+9c1boVzRCppw1sN8R49s8MLsBWNLoQApLvVEK7sb1VvDLchrcv
FNwCVwXJecx5AYyXx5KAqwyr7/RvW62F98qwH54E4aGsWuVLWDvXXuR9X83xvKgISDIzz8syakrz
Akm5YASRt1HM4cVkw6RzD1Pc6oX3UPsvJGOZyiKkrXoI/0ILlnIAuG5Y9CgNCJbj4Rm7N36XqmSe
WA58lr0Wd+mYijWvYsJ2V6IK8DuF8MiyX3vqxoEsPexjImciPt0P4YLdK7CuQr0Rl2DfIhdOcXGe
N4knCZiydIaHDWz7VzTRfXhSG8TlT6nHx35PRVPgeTAYs7WvTMbMLmJnkhD8j7dJTQLRHm6+CSP/
ny9mgxs8T9jVxQI20kXzX0L0VsUWV6u30BYkmdi7kBdrzkkW+1CwCvQx9yhf+FekhKehjHkBLEHj
lOghqm3jJtMNlwS86ZA/KTM25iiyDyGesjuYfDUuKvOeekAaGM9STZebszd8eYTOsrT55JhrM8gc
elDo9jG2ACrh2IQyzjbCIVePgIyUrd0Q9mbdpnzuxYY0uF2HFIB+jboFGFgySVVB+O4P5MEIzen2
GTJ1kblG/RDavdOhsF/y2OLfAeGRFy2M4ICpgnuEcfkGUhoD0GqsJocXjmFA5PZhbVK0gSxhis0L
4p9Kc4qJy1rzEhqtfBNhU0AY/lSCi+vKGic5/zjBOZot48Q1Z93wTSr3PTKNzbaRJXU+pjxWHCfe
D6HbtrQZOYmQkceq2lFFGijkh3N4aU9N/pcWMsOt4TgdEBxhWcG4DSKFnchtiUlNlwbKY3Nvx6jZ
6X4BHgBGd9zUqdWBFI2Jpm2bVeXFLnjDw/D0Un9j1m87ARKQ3i+d+VkPdOy8mOZ4sF8+cb2EDCNm
IdjJPcJV0LkL1U4PwYUyLdlb/7GTDfwvtwG/QsXFWTujNew4RcLUCZpIPTOZon+XgcNMD5prbZn9
9mgHJdkZxF60ry/NRHLph/yBM1lsw9nX1d2vm+0zr+u2H59Mvai9ngEHDenZgTufpRUJMZH8HGcg
2RqUQ3LklJ1tAaW46lXvsxdWv8/tFyC+DVuW1THutoJQ5tY3mbvfAw1nCHNntc1dbqL3Ugousqi+
xU/gDz9pSakOozL+mVWfhsp0FrX14BXB+oOPqV2RQVj2EluqXIYCw6tyNPkJzIWm/AukUHKbm/VA
CDg6fLU+ej/03gTEgZD3vX17utZkHdAQvWzQErwKx2KBJ+FbC5dQQninirufOkAu4LZrIrwIZ34C
/vMH2/zj/XV5ycFAETDQQaPeYar4ZHzfRZAUA31X2VHpaPqepddXO8oZN2+t77Scq/EmXRX2x9Sf
3SYju7xcHTiwZ0Avq+x6JQg3UCPG5Hq2STEqETvRlHqJR9uUpmADTH+zdWhcg0udLu+N9r6dwkLE
jpGEjLyyG6uEzsGlHZQsFU4yreBPwKw3mC3WktT2IiYhcuwBcSUBJSkGzT2NmEMj1BNlX/GXPjPg
lpNas7M3EzhN1ba4K/E0Nul42nhPUtFQwAejh9cPiBSROQSVnEAmxYPjusmvGlzcilY4LlNeOtfV
ojSX77C8mr5Dfh3E9IQkBq/Rn9Oa8icAtR5dYo1tuDYX8KdTLJCIZSpnCLd45GLjHKlwczdZvLT1
lB4NLm4ot6Zz4V69PWGhr1mygfnMjnrxe0VKz2cOkPSQOkyzVOWINjP9OrHDCUzsUTQWh7+fLfyX
tkYpqcah3Sl4r2mDyvcdY5AFuWKDKOJxrfi5/e588LmFj46OfwIVl0wvrCEZ6tFViM+mNn3cG3RT
ExfUZmkpP+JCMqIVLPgrra26xym9EE0fWWZfrHFw0Kkzvlbq8CZhp+iB44YOTTjse6bd1eDbwp0r
ZU8VxV0GwNmJZzanjMGIdnlL01VqKlOBJjzeSC7Z7yToGGogLunHhijGBLRpapZAgPAPawqkR8B4
ZLnYOK9DFMs4lmW53SNK0HA7CpM+OEa3wIhGfnG3+7ENFaoIvMmgBz7DXa5aDskev4b6wQq5JseW
J6wOYs2UyIx++Mu5H3m4OX2MughlY9fiFzeVdKW5bpgQik5ZDHZ1P1drArl7Ilt6MTBRyUaqRJAz
WdUfmjrEVWY0DwYnBY0SPkcVZeTU6lSnTAt+uQSuRQSMHULQKXgMhtR+PbGGiCxsRMkJUDHTN3+L
fGWpOp4JHxBGZz+DJHgSwTWNicmJJp9h30/baDVfUF739r22gj33ExBAz6BlUbAvZYrbKmag97nu
tigvrzVO1uYYBaWfWS1egTPzP1Cz+Y6fbxtpSUEkmDxtUxVNrkRL/SWCuKB910K3c7zKDEZ7kVts
KPJVx+SK0leI5BJ4Ntz9nYWedCC1FSRWcQU7Kb9idUAhicJThldyOqXAL00Lio4MWinw1v4Mu0Ht
3h9qqBswjVNZJhtQQ+rZgiLuP8W74AGWoZWwZ4fFRoykLt2Z2l5k3uXQ8qKYbJTpsEtL1mAF/OQI
5e1m0MFABmhIe9PKXF2+HaPpe5s3lcNv6tcQ8rUfWJLIBbLGXIvzpgLZRZF6owSaT7l3/ZwFsmuX
h7g6LHoylpRrHz7+U70SZInyrqy5LmgpvnhrGDM+eLfZOfd+qGCqAgVlsEU2IBo2/so5l+qxyv5P
sXsY2WTExaA8OiH5nAfoLtkJEYZytTydaIrXIn37FNv3XUJh8KdTKCuHx/5ngsxrA+HGYSmlaEwo
olIFUROQtLiXFQdL17IpPUgNqNaUb6hKgfR5WuXEUDwkQ/x+dFmBhpCyyIXwUzRUpGBKi2lYMlP8
Vuy3H5EVH6PbR2AwuDnrFAzRsnsVvArULgQJFrqClq8To/N1psWTrFooP07F3WyxaxUgfb1UgIHK
EppZcvVJo8iIk1Nt2k5RNjkdmjKg3fQpYElpjjEDZNXKjJiIg70U2Qpn9n7WJ1NEdWGGuFJi4GFC
xaMyafnA8DXI0BYzcVB+2DDZ1Ub4DJmVIL8mWh2U9wElcGj3Em/3cbOhe3RSRPDqR7yaILqjPJfr
o8oyBsSYc9dfdxe1s7A2vcx4sWt3VvnThZT4Pez12UyhzpzvGGKLynm5f8igAnPYDa0749ZCe3el
iYrBN0bAllqE8x0lPOT9kZc/uiB68JJg7dSY6DIdHw8OsBpLiprPL/VCkBMrKyDcq1OcUmiNPco/
yJvoEJeOooyFo8DGkfk/tJCDA25EgQG4luHXAkCB+u9+cQFIINbY/8RtAsECQCxOfcgZKapQqBrj
DL5lpa5Bq8x1sWsvLWoBDkVUkMDEJ5BCeM+drWwWCgnvJ63pNm0XhOf3Rbp2UDDvs4JUZe3rxdAR
u7A7njEelb+/bHEJNgRmtnV8Z0umJ+JzDKK2esMl2vDdjPIORnVai9HDmnqohxQP27g5B7+R3nfB
fxo+QRxC3f2dqD5rU2D4h6crr+eGyDeuE4VX/dJgSYHG4Y31lS4MGC/JTvkXDYjhcWSck2+0MmmI
jx+51mgeyrmFzBkiMMp9oWel+Dm6GvrI/tWB6jqEu3x2XCeJ1FaNDRv8Yng1CNv3wQfsdYdoSFY4
vDQyVHEyALOtrVfg2Uup6Lql8TWuhhcrq7a3HmUrowFFmudRaPZ36FYtX7DCh/R4ypO6hEaUSQvi
BQdHNnO6wuXqxQrEh9Fmz2xFI2UCJ5/qYcIVpVZQRAmc+NpOQXigJi2ae9aq/xeGyHBePZQ48io9
rWCDEyackZZj+bDM2nlUeH47KWkaqKugKZpDdSFP0m9RkFtmhJ8O7Tulwfr2JSH9WJBUcQqZasog
kZnlbU6Ci8EIaXDVJR9rotAq5N6P1YUCdRHro9fbNeXRU2QbH8JzKLbjsFFhfEp0B/h/ENSJuNnS
i59UvDl3guLZhc7Mhgo3q5qUhSCdO+fbVP/LJC574z9a0ObhumicNtM/wZc1EK6Id2BQ6N7Ns6RJ
0Le1vUBUYuDlS8z6TmBL5iDuMzfrxICfBC2fCsYVtrvuAqiRAU4XWacF4qd2Uhq4SEpktKKHNr6P
Iaftsm9yrW7ihmxhQ34dUFfWEcw2/JN1ipRDrC0RoaCqiBvAFDm2gnMs7YBtQGI43AkP65zrDQnt
LLb7/HR9RiOHkQU+yMU5CF55THgSJL/Jh4C/iplF7/bySVGenOsQZG62hpZlTVCASz2+pdeNUsro
haUYIKCqmGHmPB/xSD/zNT66DoSal9OEwq5qNkqCygwtRgyWvx4DwhPNjRQ58E2vMHX+FcafxLl8
sqwjNhpztPqwqQgEM4FOUnFa1KLTjMM+XaS/i03aBDaoI0zzNzW7FefroO/N0LJVHVp8ekk43gA0
clzca5aURMPFu3w6OeA+m5EKZqismqbb5VNGQzYCMenBpn/5nnujULeZbv+W0E/uvTa9qX8LZ5J2
0PKDuOJunNAVVkMMOdh15FEw2FGT0LOzKgnBiog91CkEnd/rNF7RRija9vJC4gTfjq8OFLnkR0Ax
b2ZLg3+5x5FWofGXkU9iBUltyXuzYPzActHIb79ItBx+xTfsyO80sLedHyrofzrak3Vgt1o67lQ/
otoQIl5TuyBMn8NBLfKR/1iIFW2jq8wHoNUYkMr+zui7sJ/hJdf2YFUAZ/Xp2q4hdklyWC8yKXtH
j1dQMyqeqfVj+Maf9W592q8IdT8RemRtpAuxszl+IFA9HsN6xLgHpvjhq00WrQlaNnrdJWvQbOJK
hz2k0E160rh3RKZ/jkWORr0SjwVI9PgKCxe4Jqa6Ywu0WBdp8YpBmukmFqfz5TiMunFwBfPOuqUi
Vn0+4vyOrp7TSslcBGAwvD/bvzIjCfYkggGkbxNNRJUKnt+5Y70/bdb1ZhaIjqCSvNc9sgBQAHF2
vGo2VjYgAfIavZ6OSIVyTdBI8QifHzKL7MYhLGY592rx0TQ3oEdUDmAX7ntPVnnIPl0mKbSqr5ei
LvAikM3mUb3OPM6MONGsTUlcNd7iqCROx/3Q93RoFDUbPGXN/UlkJWS83bhuLWkD/I0adE6pcIay
JYGBpdAF3PTgPwbMrGJdbMWyLkiDRhoS4wSClliZgG4DX7MexOVm/pqviIkHGiASEzp3FPnfqfwh
7GMC73LhIRMaT4rSRu9tLeEFPaMV/hIRl8jkaWZrzUf2NKb2Jc8KZ6bYLFHo7Jnfy42PotekemqD
5ZS2X+vjeHM0v054SP/etY39nWTZhSKZ3p0ykL1AgILH/fZdP2L2K1U4sG1m05ogju44sdQae9a5
98GmCjmsJvlbNHx2PEgZrHUHQfhdpT4Ccxi62l947+VQtXhkaiAh74MrJzcr6flsWI/8+1u+M8dh
vwEaeebUm+wVJzS5LasNyx0aMSNpnwVt/J1zU8k3cB8VrT0RWrNuYDq53W8Uard5jWupWxo0f0Qg
/g1AX++3KXZgdG4qwzIMYP4T4cX99rH/t5yy75IQZnO0fCwztzh2j44AjXxAa6md8qhMdt7EdbCY
kGtzJUSZ+Lyel+FHp9nwyU49uWEpAg/MqhnCpOOk1aeNlHdhqwVYh/mjmejFvsyM8Ah8KW1JPnIr
PhfJ3jx67Bpd+UcsF39VQ2Va3O2iGxLT4rD99ewrLYzhaoWC9nO3/l0WNM7hP3d8clwl61F+qhhQ
4vpKyz7pJXWOKjUyKbGO54D3IssP8Sv0nLZb5TvM5Z/ffMMs7SmM/JpJaFP/mYPSXxfeRYpTnbQ5
hkDwz0KdUrWxFqVqJWF5LA07RyFhlsQi0HZoQKpD+08GYdsbci5PO+xheil/sNOEhPidJ+IjGqQn
dnczUnJtk/BebljfWEupqPPRvfDE5/HOJcuXn1wlstg5pEohtHg28Tx028/62T1vNmPh5eq4aLSJ
A1GihwUtWsYiNK06ikXDRtUopeYbuILGNjxcNPY3h5kT1wFptjBpx8z5TfrjhFVhEZ8WJciHkxB7
zs5aEVEiYO7xhoQ3MSftuPdOQutJ+pCHq3y+8zlDQR43RNZbS5oi8G1IjLm8Lzx66bvImwet2Q+X
KTg/xTPs0UFlGh0CrH8IXNBI4xuEg9HGOqaZqE6gECVIw9brdL4r6Cla3cO5EDe/bjKRU2icEbr0
nYZVpvX2do6wGfvcGYLd2kBB4gZJq5ShJRsBblwXDk1DysaXGJgh9Twf8BVvZqOx/AwXEqsI7lEE
G/vm/xrLy9k87EqGNxyXH9oHQu6gpvXqBqnKAzhq0xKdZKioMVkkkJbVf5oeZZ6URg+179kd0++U
m7CHgHL8ua/kmTAOyyvDWLvsRrHX0ozNmZjWpNAh5474DxVWP3ISbRwy2mUq6J8iKAzLce15sJOk
2vMm4lKf7y3dkYs5EDhJt7HcXOMdoMR7xY9Fm22bXFBI5dN2WOX5rZoijSGlGEPFVzXla8sksqej
51EUusxYheeRuQnCV2Mdwuw1BUIwzKyovIPlszthgQLF6dwgczXHy4TE/DwQXwszXwPnrLtieeML
OESfLp3LoM2JsWFlNCFe1e4zn0Pn6x+c6i54XewKwfklH8d6kmD/R6COT14VM3+mPTD2dhLEOUkX
ij3Kwduym5ybd+6IWUrH0SUn3Ru6Tz8diDWT8VZhBRDRweHTzdXTpGBcxK9xsL0E7LSn5DKFe6mA
xG9BtmotYRH7m/szcWzb4eeYOIP2sLN/9tfrM14J6IW0rRH2cEcf+JQ5YuZzKXTjG7FNC+dG/983
8E82He/49nN6ZqzizbRCFtmdZQiyj9nvdMiEOY+v5FdG9VYi/yy3lAfhk5uo1+txd/4OXZMQ+uKF
pP+Xin71idn2t2+DAuUvcb9WQrHzfWUltcT7hULGfO+MDwa+GVYUUuUaiDtk9H+dLpkSeptm3CDe
3c2lC7+vAGu9jSIm7AzlpiPDjGQgCiLxe1qAuimHwX5W73KmQVGiQdP9bSh/bnrIsSow9/RkA9Ty
bFl+yNLxbthURTqGPrM4GuWNUu/RDxt9dym+qqZTWYazqsGmIwCQqq61AUULM0UYMyZambP96H2Q
JkpnB3qAU/WDBmi5Y0Tu/C0HZtFbCK3jWMg5jXq3Udk0WXJsZtJt1UbbLyQJoMb50skYrAbVx9Rt
lCk6SuqURfYumTzF/8II6hvCWKNjTvzwrZAee922Jq5hl9321efvddS8M7hmrhJubyytO1uL1jND
dMB/B37p57mNYgGQLU2rBaD+07WJjNIbcLBnYf5IKJVe8+7DGQS6ckPqEELqx3RelMSztJ8qfjo0
70Z4D36pPVOGx4OsBzkuyhoEqrhUpzu2UbBKURaw5fwGA8cl5ZLIwFRMrKwTex8RveiIXkMNOfKy
7DA+V21oznws2PU/SoY0Kzt6dOjNycE8b7P36MpYK/HmF5LoBj2p/DBCRYKpQt5JRzUJG+OXI3lL
r/evoli9T7H8Jzat/VVUaw9ic2Nd/HeVPIaCMdXP/aewg5b0afh/esQ6NTiC1f2krm74ZLSTN7bD
ebpcR91lYdBJ4V/It2T2CSxmR/wKpHz0L7WcgoL8u49MJ0lmjvHVVIhwkkTyF9x2k3AG9RhJ7XMT
x5ficFhh9Zdboyd+cJ9i/YVSv27G8Zsu2QExquOyZbDzQYMTNTzavvQHy9Rq4mn/C8NZ59Ug2lG5
1ozintMgvX0VVmBLg2oRvZDVTolbyTNYLA4yeZb+/orm9YXlu3B2u9A+AOjQXD/NwVMhHXlXf1sE
dk8q3P7WT69fAz0+3Cg8ePU/AHcldlyzaSoEFLXSCo82PgnH/Lgm2to3CDFq/hZfIDyDJTY22kI6
UEQ37gRhi8U5nRN9l00Yky5r/+XLBi8KzpPIEwvjXi4UYmJyAIryUsg7Zf/IBLdcH4BrRX+Vvyaz
SEbbAv+mNhDH3aXAEss+F/uJ5huRnYTb0fe0TLKmOkrfs4CIJk8RZhXVV+afZcPsjwSfypWYfojW
c3ASfQFxLmaJGcrWIzj+kkV4nfLpC7SV0nRlAHyHKIzSfBbyXDYfX9bS4viyoRbtH70eRsZqHHqX
iW7YEtnsUAkjWxX7nUnuQzPCm4VpdElEKe7Gy9yUB4jeimiZgmICDrW5U2ePukLpBezqQ5m5R817
R7I62kuuft0Np5xJZiI5XZPDFtlygmiN+M34f7DRgoNZVlWnD+zkgmgc512LomBF3X/enf+qZtBb
GZmGrjl1+FTaPpJfvoalVz8tV0kdpdULGF0gEWD8ztrK9FToeGLbwsLIn1LfKnsbuCQm/YUdTWfE
TDwAeHUE2SMe8ZMwlJRt1oGe7dQjy9oSB9nGCit2kcTIHzejyXZetQI5fH463mf1PkfTxQJPpKTj
eInczzNn7Kh3OgAchnbC+rjT2Ueun0Io7YyM2wRiYi1Rx86Ia+uExDZgkqO0bERFUfeSTDSrG3q1
cz1CVaG24x8ELzTWgbBLvtB2Gyl8JdbWwbIM/PB6hxZKICk0QPZaXWCJqrGo/LoqWKdmX6kOVcPf
ceHFmtCvNlMIBgijPNtscHFo+xhXSSOz/vNQyatRi6uMWK7OJ/4dJgZdNyyX96ZxqkZasGX1OayC
Q2u2cHU6Gfr3bsZFkTdUWByCBWJiOwZBXyYxSx6Yi71JIy1YFq8DzOBUUHvw/MJOXpixjiv31bPn
05Nhn9MOowtuXqZj3YKso0HMVM+tRILQmjvsWqm8mJ5sCdUkwGiXcTbceh3LOlfwXNPETjChwE81
+lAkG0KYPqzZfUt+eFaca39G4mIH0uNzdTrzx1sfUvgtYHuOGnNFAM2mm5z/LmE84RI9ab77WLIX
kOChkWQd1bBo1ulXUGnRqxGITNsgWLmfpAthcj3SpzeYvr2OHLO8HkROUDeVjGHP0gdhyOIL31vf
nTarhZSVCz9mlOMVUNrs11ISgN8VQa/ZWW+A2ircQFqrqtdMdLeTvDRJyZawP7LsBmT0qSH0yrii
AtskEoXVWVDnP0eAy5ERfseDr7NxFfmeYwFqQSo20riKJ5b/PrGfX0vjpomu9ljxBp0JVEamGOa0
ZGb22lfusl/Mz/v/h5XzlWJYVYb8AMBrFWEKp0JFjCZ5UArOeZBmqmEnlfT5EhZW3rvy1WakHWaE
Tote5PWwqEcCQZS8SFBa/oJS7mdZDSV0WVWs5OZyaAGKkMMSX7xX9j8ZwVsc3olegAkeHQ/eW0X/
jmxiZxoPKu7w7efhLHnmOAuMA+17B4MsGZMGjI3yZMGbb1q/XHtKhxNHRpRH4eKpq76cUAOILN7W
824ZsIpEMaw9A/XnCf8mo6SvQAaFpMRUpxGzscpJ/cuQzVdKgQ/DXv4JFX9U36Fe3EM+cJzyNU/R
XUZAYfqJP9uMN8zrJpw1hutUn8of7S04FsFESyQfrj1VidVqcAQzM6nFXamX+l5Vmo+GdbtzZ7Yh
PvtDddqkDnRaDeQRiHi/7w9sPo4EdxYvIMQxtJMsz1SQgrEB2j8PW1+TIQKsRCGuyZE/0kVS740R
kUu9oZ6zDVvOM5luql+wpDsK5ydkuactEvcseTqOlLPL/cTkpGLuimCQBPn4gE52T/G4bwyu4026
j1URFc+lAHNSsiMvXI2MEFoH/D+OeZEMBADUE+vfn0Ct/QZHMC4dPWsMdLd6b2AHrNmZEBrkIlJT
wvwPckQB7Hyb1ZxBmc9yhzsMPr5XsKZIyZQH5dB+o1CrUasp45bg5rplUuajZPqpx0OOxRaE/fPd
pozZ5fzp8ZCSmtHtHcTj6AOOv4fKFa/dmfrOsiTEdZvOOVuowyZDv7Noq0+UdjHvtcegLCEe+Fsz
DSV6G47w5TGuf5y1HQivQW2crz3oW/TT/jcui2fb9E+7X+Ss9pLzknD3sIoJGWYs/Fle5Vl6Y3RU
aACgbKAMLv63cXTiu5svX7HIiYELgsLHT48GHyzEhLtp3blQt+KpKpQ/54txNJfrAxVyT4g3hXTi
YYT0S0bFS3+eMz43VrAcEsFV+iyv8YFhgoDAnojIJmwd70DZBmoHx/agTgF6A361CrxYKrVBnfvl
mqEHjbiDs9q4Me7+pMT8hgCiaMc4/0fGFRtnuZttWXaUG5DtcEx+Gv9YxJYaTUB0Mbm3o+9tX3Nn
JLSvOEpupK1vyVukn8b2z1pak+23C7PqdlvBgeYJ9ntIp6THvhOuL2JAnqoqgONhSnTqkh9mnGiy
1UGb5bLtdlBmwf832/JeDMPA7EjZ/Sh+RmQu67BOqLFlplXm5S/7y6fUKWLnda2imC6oG1Z10D49
M40IMBbwOJMuLSHIwPDnVUPQF7/bPsjqUHPYhp5ruKrcHqGmUrQNL3Cs+JfW9Ygp2O+PRcbDYQnt
lscVbT8MaSAhdNrpsApfng2+H6xKkS0QDu2lpKRjbn9ct3M7Nzz3+zVvLbOqG2fsrpJttIKgYSVm
yJatkHrmGMmOyNoWhIDo2ABM2MPcSM415ddsiAGOcRb9h2DWB8RVLGgQKFNO6BnirXUbsStnPqq8
/advMmtcLvT1mTdLdXijdNYQfKyfYNHv9dplwddQGu1LOyOonW2D+8BNyPnG5WnzrmTACQROBpVe
nh/XUoskpDu0VZWkJVrq+ZY8uPRoOxo1hXIAKHqQOeclv/tOQlXh5C8HqHDkOHi1voWDhNwbkJPC
Tt/P6AXoEqqch7JxrzY2h+7fg3Wv3LfsYXvyTwfozwcr3URgaXwMFt7VZnBeBNNyxOvzChEmOxr4
9lD2e4+dITc7H56MrHivbUAdmCbLx0y+c+Z/gjCEn+uP2xcnwKRF+ZKeXHrv7OxRncMCTQajz4LB
TEF5efJFs26+MjIyHduTCA1D3IZxOneUUSBCwr9EHQYZO8RfyRFs+m7DJi5HhAeYpKi2gC1yN5zo
YZorXNMUegSg7baPQbrqry76qiortVq58P1kJwp+JdlwWp6SV4y1NatGN34usZs/cOLqOMk6zsrk
zh5r6m0p5b9jwHe0VGTp9G4sbpaFiEVUFzrbQflcQeZh3qkKpmB1xCL8z2Jvkkjl3IU0NamNOWVJ
ClLSRuvTt1XdMqrPNpPLogMB/dE00gQNcd9vsTWkeXGhPXylYIzTewQIEcyp7y1xaYTgRo0yskIq
ts1f8/Wmw/ZNwCCSap8KHW5w+1oOfRscQ5+730lbm4c6MAfkjZ2mrCVV0tJFTNd34okC49GANn1J
NNxdOcvNRli9aZmcB3oh1/q4SzNbLykDeQgwl7ddFpA6d4etpg9D1HClTvBrtRfde6bFSjFA9CJb
nxZsRgYB0UqvdNSHeSYt703P9x2zgvAiYpWoQ9AiFZcYE/0S0sMSCkOv5EhZQ1er8LtumMhJFdQ+
rYwVP4bSt7qXT8AAeFzBxSQ72mzllc8b7Pllih3AadXyxeRNxRAPG4gK/eVZrdmf/gTsvZrP3ADl
Rt+Wts42WISr78OKHCth4OyJB5eBs0+GKAtWgtrf3apgJJg4v+ljKBl3ZHePrlxhuHAO6vmW/HXg
zNamtlpFc3N305+WK18tI4Qi6ZEIy8flrtDeDlnjre79rGiJIv2o+7AHGVsQqC0aFzB2ejcmRAMJ
UxmEt/tEYVVib80M0ZwuT05mf+W49sVh91nzXQ0uS86qmo7ORWSCqc5+9nXujvd8FgAGrr+N7zi9
cRKNEFh8tYoS7fWqCLVvPOxdprlbrJxFLS/Zl8E3arVyDxW79/S6+BOOF/PTsLwFpXMwBANApJFP
J0xrvNHXJP+DqD0FN3f41Lg7olxxHY5bYeunGuNd8q0CrgLlfZvFTTawMCaz20qf8h0KHoHyt4Cj
vIS4yYt6rg0B49rxjS0odq2m70OzpQDYPCJ/uh0qSdD1YJ3TijpN3/3hdVg3kuuZ+9HZuFkX1bhe
kxO6x5fT2EE1PxAz4P6MRN/y4tJn+UVElV5uLyhZrKDARY/CwKl3+yptOg/R7IJ9lEMjp8T7IZwN
GSXLKPg4g6LnMeFGncb7IcRULHvwYaABl58nbe1B4iZZ8UcpHzpVToflwFcQ44N9dIOgqgGUBW7s
Wqw0FGyHfnqlXFxDd7+alZTARaJvXaN5YDrnp/RUBMOuhBGofyqJByIP6E2N/Gg0yImqkzpcVcRM
TsbI8KylaHoN/ZNXjODAP6KZiPWrOdojWmyC7UuY1utTDI2c1XiRcZsQVLIUILyG101xFHKsCBRg
+9qpwZk7gnFO0GsShNEpW2sQa5O5chqggBSJrY4HKY1H48tL3VUKPXSwyFl6lhaucx4AzRg5VlL3
xX2H0pVTZvmbmjR6BZxDvdG3ZTpyzz/62dcKpVqKVL/UZ56KSdEOcNRcw3XIoWCIY4aYVYzUx+yd
7ylo9VDazxwKlTCExTaR3tWdKmdR3Uai7hfl0vWO0v5u/TdqQoxbREv1PAq8JkS2oBkP0vBHdtjU
L23yl9Xby8eoYSsrQhy6HjOyf0DDLS0C5Pgs51yC8wWMq05FF3AB5gLwqytk83tNRAs/BE5xK2JA
PADYrrH8p5PcV5EzP4rw1w/lBIc/FkZ1/WpVo6zbEaDQS32Gj9eCJF9WHg4KydzusemIDdUdJ2yT
Jq5on7frK0JD6AW0uG/rbjY3H/r588i2E76zzDBGd0HSHcvt3ts93MNXHVRj24xxHT7DR+65qOwA
UoA6huBSwYpgC5+rJvZ1bAl/dIE0boJlTmMdbFpPpMAQGl6uBXdldimWE+qQtFTIIMZNkTpFRdLd
YYrJEgSTvifqGfbax5vvdy8/V2m5JcPrq9wyE1Of0+KltMJNJSZir3iRsNpa0uLnkHURRQnKYirs
k2y/A6LKogzNuihtUDY0iB6EvuvPonOA2ze/PFQC6dK5r54k1FCQiH40C5ImFQg8V+UdsENm/eZI
AD5tJe3mMY3P8dcFpwk7AWTuBmvMEmLqvoZ3b920eCi8FuD5aHee1gtQbVjxBuOVU0qc15YZa5c6
ApSiVYVMW3zck6G2+W8Dlk/X52LBbX6J0bHDxNS0+VhzabAqZijMlmT1Ud5wD1QeCrjW845u57Ok
B81lBf5QhxcAwYdJj8Hy7R3u+031tdeeevbTKfQOfDWM+AwW6TN9VuPr+zdDjCOBcsSjhd1LIEHa
LI/sdNPE9aU9PxYLUCOPIyeIFLFiJ8UViq3fAx3/5IBbBh8Iqdbhq0PJNA/MlbprgsLd+V3jPehF
HdQPAF4XkDGAKPcO9uNewkjw/VHuJXMwvUlBwvffQeYLeZ5luZyrnqkWJ5+a24XOeoU0MMr1GdVD
ELApP7bbJjmvjBGVTFOpkqgxy6kvyVqW8hoO7oziANzzXn9r7Ip5AdhHKCdAgVU+JX+9K14490uk
qmYd+s44/38K6OkhrseWpVOvqPHTluYD1sPaQuoXSGftIcNInHA8vJ2/YvV35Ue+9WcPJRnn71Ln
t/LFwCes8aQisUIHvMYGlxOoIww1PuhxcDlqmazN9/uazNFB+jsC6cDsad6ACjSt9VuL1yFOPSzz
rG4TJB1hrvbBXPHAwLj14Za/EdK+ivtOk1BZL1Bw8weG40dHwSleWiNnLnukDS4DuTEsszkpQ3/Q
Wc7lK0XeO3F2WX6V6DRE/fXb22p5smCVLko+9+/pLHppAWplA7bZXBxgxMj7Jwzj+InoOOiz6EvP
T5wvSIlnlZn5XFVvItcqcdTNm1YSlnTuTrpJU57oyqDxT5uCAS0HP5KuoP4JDzQEVKp5ZVDuKyQz
sEmG779tN1JT49PSOW/6OPaoEPKc59Gg49Hl0vAlstPDyaEzJQIhHyBbzmHxJ9W4ONiA42z0FVDp
Fi1l9Oj9e8/nCYn+SGbV3XyuKUbqrOmP21GWuSl3YO0S/rqnEf0vvgIfa2In4izOcnHg1lKXou56
pEWs5WhK//3I+TWf16QiiLybFz1RpdwwQ1eaUvwa9f/OsSNG7f/6yxWTSiLtyEDvBn7T65laZDx/
et2bXFClOrtjvI3gsVB9X1ah1t7BgLvF6T9PGgMzwCstY7MK6mwh78uXnE/Cgck1GVBjpv+B+Fo6
QRnViFap5S0Qu90rAP27dwF6KeNl4GVIb/pzymJZoCBj3U6jlH+IGukid81ZJmSceV2Mqoofa9no
3YICwz0itFssQ0Qi0t4vwuD64eT0wrIkX+rq/WyG6Oe40ol3MzKi3SIYLtib9lXB3akmsnDqDekT
+VK3asyTItZVlZ6NKS5VJtSjnQ2tku0ir2Ge3Qqmla7p4CRMwQbInZEyFY5UC5qsCuf/H04UGGGt
Q3BB0Fef6QhSaXXAWZ10eqrsszixclcNzLeDUt6YZRl+vnVqB9IRUfbVcSn61TLwTpy8RC7QR/ud
GuPAg9saN4GKOoTHaEgkB5js83zNvO7E6ahMyB420JtLH2YVVPiINFQEgU2rCLMbkJ0PrLw023ZZ
BlVFXjeSo7r4/tmUIulvQPLIw/Ahm3pem8ulMHtZTxGPWdQPJdDJSkKb+m5A4uZK2XoyYqc+rZby
i/G5MANfUu/5dTMuxfAFQA250WKavv1QdJGjb+eBcuzYNFw33Boru2O/Hy/Wlic2NRrCWFiijAWs
3C/7HyoZf8O2OSKc4qnCjjgyw2fZqoiT9jMOw6uuucgx+0LfphPlVtUMrharzs5zyTncC5/lpyRV
fqju4S2P+itrdEfBkKGL0fm3M+DqB36MZF+fsatoEuiOL1TFlPqWUrl3WYgWR8wjon2uEdZES1ND
BogIQVMJ8qIuhwG/an8gLnPUtyW1ixfe0vXCgOhKwDGp5pmumC5tq34mNUcX8UhEco0cg/Pmt2e5
D0db61i1vpyoDLa9q9o+aNuklbIoFAuEvCRN+UkIWFcY+iWEHFkbf6NjhBWKPjS9yBTEsizS8WGO
vt0/ivLUDquLPapSzLIVW1Bw7TP1guXC9AN4lfKB6zcjRfyEFVUp2IHwkfTR1rOIZn5oAUyQ7Rho
F05tNLUYfc2rCOSl5cDSfJMQHelgVRhIaUiwz51Abs0LgvMBHDLzv+DdjDV0etlbYUpvn4TcVWN7
ss7rGE0ph2QcoolExRAkZyPh9H04Q7StTFKxjC3mBJi+eIs1aPY3gsRMpR0hUJSRBrWWEOpcH14L
cgVcH7BjtloknGDdkLp0GRQinLjnMjlO8lklfCzMk29UJwroivhzK2jffjTaydI1e09NPniTN9Dl
m7eBM0bGwG1k58PrG7U+ocnLbNk9QI7K95+/vEGbciQr0PdDyobXtiub8gpyu3eL/qVFAzUTXmvf
hCKnVxMxTXYsma0nTXpzigzUkh0nZ+3OmP4jl2gODF3F9vXLAiAaUm7r4L93UaMUwAc1GV02AU3W
ExWVqTWFQPPJWqWS8u+EfKghkosLTZuk8ZsCvAIciV3OlXQabcBCUQnCp8q4XqDkhrja91OjEjKk
5h/iz2G/xLxNOpi4lxGunvRJ8tS5XUEd4vQKj6dG1J4oSd7mkJcuHSCdgIzMUVoipoPChdLtB/HB
3gaHFefLeu/fK0EtDNtbrmvgP51s0FFOu+6zr2c61R2LZ7BXVl9SvQATuHp23eo7a7yy+u9UiIc7
gzi33t9MxJWuXmFmcpBNxBmaDqSmff8wFZ7r3FKQXklNbUerY97+8LifwxIqbDOQHcoHp5YGVXFj
BaN70PILUnttORcl5SOJ9kIJhuF/C78AjrqpMn4gHhbFlLHgNIvVmj3jQGQkqb0vwdVtSFKa8TCq
nO1G6beg1xZ0o5+JnwwiHJSNFNbqUyFm3qAgDzbm+3eXByrghXAxyIeRDPtfM5SLly1QozC2QQJ0
6UBJpVMfYgHWW4TVFryO6/KGzs6wrpCzsy+1/cCphq+x+K2me86zSfIY88AVdPvZaaZI4Gu5p3Vu
E8fFh2VCPQR7Kfxa2TcyapuNwVVVZ9JXKu9hwJnRSDkPxtDcK+QWYRpmONft0LIKKnvariFKzC/g
oueTDaNLoFp8e5jr1f0/QLy1UcVnbu3XwPuVTC0nBF+QPkSXoya8pz0jlqELzSSWBXJTAF7apLun
nVBlqr+sRESE8J1jLUhjMSDWVip4Ef/UehwfNG4qkDwNkPxT9BfShuIPNsncAUAKWbrJVcFeL8/Y
DW1JNCjNgKO+4GzdEX1djhWB7UKRX1+44F9BDUq/et/XzRt7dkU9KK9wSKa8XxP6mmiiQvVOv2Tl
hq4UhKQ3EPeqpAioMzudrwf6VymmTxqi9k54TpFB83bFO+m0hgGA6c3f5+NEUbDJCG7Iq2Xs8SNs
9Qp08fQ6cnHd+LYmUWVc+MzjWsYtW3h19OTa46O2NA3GUwKIp7Y9gwa3a/+nS7z1hVMF/EwWtAuY
MSLVoFhcA1/pwlgU9nffoZvmVWeegUe7iwWTfJHR7sKcCN7iODRX/E0Jkzj7TlrVPYZLc1W/GXaE
ADIVXtOiZHcNQOpXE6mWlG9cJfhVqpgJ4jdBtGMCvPqa9n+SEUat3h4UV6iz9hdlt0/9JIfGlx1z
5ULO6/Pgw0HmHEFT2n45+t8OPM5po5uGiAUJXTwGSmrpl0KWJKE3EDoeMnxsVFcbDp1vyfq2J82/
pkQLnxF4C+umkOp9u+VFSX3NFrZvIncuOkdmEgOIryyxL+MZXUnF75nHS7mapM86om4GVbakzoqI
jDo3lePHUFGRnnMCRsiY4fn8Qxr/8thxP6gCyfwfrdF30F/+NITeUe9G5VT+VFeQXr8S1P/WTt2a
NEHukuYODQ8R1ccLSXZELnubaZQqJI4zFnxmbau0nUfBqdCCaRaly8WKslicoGk68tHTsW3bnLMJ
TLZibO/1T0KmF8izC4lTxk+/GtGwIR2G8AUlnb2mTO8eY/p4Z7Bo9kGVKolaixdOoTlJT4MrHaZ6
vwFplsgAFqp6sXqKpw6f0va0igE+jj2n0+WoMltByKrp4asuAmybKjqwY4MV3J0cjHyYykbO2wZK
79wN+39qrK9OvoM8xU6O3FlEh+763GZ9s4nYZqHdgkGzFutjwO4GphnEPtgXMrKuHROlrZOogRQ1
e7maPnlDv7Dxt66hw7fQBrYVM60Pqs/ANOJJPW6P+6OjqxEct5+XjxWOvYu8m5Q/g83qtJrDigT1
cyPWLIGm164/BvO5fHu1zVnwAa3NgiI39QL6pTQz0wBAxwT9NMggP0zJnPjYPxUwTY0upbQD4YMG
WeV5+Ck4yZ+XMyHS2Jbp1Z+TW6Xb6Al4EOEa8peiKFc+O7v0aef5WlBKCfi+mkKJ+N30WVt1BnQD
7EtuGbLfI+leZm4ErxqPey4704qX1fQ655kxcQXf7CVE2vFxkWKlKKtB+9lvLLNordgRjFZFy8J2
WbFjkSI1BnEJYu0dYZAlSSDJo/OUN5fZuvSWY3bRK3eNUxj3OJ9ZJGwFiSp85TLOxP1LSYFLy3V+
4BbR/LZrcKVGnyBr1nlnUWuHbUNJKF8FhplRPccd9fb+6TW62TYOgCqYjX5mANtqA/8ha8w6W5ud
pyn5XvEvff1KrPVvDazojjVoEsbY6uX91Ou+KSztHfbj5rC1FU2kkfXMj8C9X/b+o0ZZzE2djbxb
oxk4s7A5oS4UBdf2q9qMjfeyrYHrPe+eNQHjBGD2cLaDSp2efnA4gcUfyGQdV29mnUJqWHgw4RMV
UrLa8kbC6S2ZUqjfRrqkM8AQ5+1BMpIi+y11H9lw1oZjzmwvYcU1Fp16rVBx5sng7S8swBJzBAoI
AcMIV5jLI6dog2T3h8xMF5sWghNtaefV9PtkrBUEvhj1XV1/AYlHuSKlFt8QvvUM2jb3M8wHKmH8
fhmJHOBaKJ5TTLbbSZs66V6kgDx1CWWAqFSTvUaRwbQqGPsbtb4HQj4vQRUCaGGegkZtWqMiZnPS
XG0QilrvRoWEhdK3LiX6/YNTJ2qwu2mwGYtb1wmntpJAqn4EIQ/uZZhMiopGRSOCK3t6qcpXivTL
uGTEhqmkGeBoqbiCUWFIFZ/pLq/M1L1O5bnw8RTV/GxLmnVPuxKilGWtf8PfzQKiXGrMebcYeN6h
WLPMRqj8Vqfexw+SFR9Q6160AM6FlwCn95TZ3R87z+7uH+XkyYcd1Z0ZvrMEuIbLknZyYqacYTBD
hLqRaO1gEl+9b3cp8p9qZXniHODNmRH3/9llCxpl2ldGgHTMN+RGVr/fETVR+VdEUXOqO4RvLxCd
+SlAOGObCvvTkT0tO5gO15iPk23psjhfztDchGcpfx0BT7MQqDVJZo1E5dnVixx9McjaKTCi0Q47
hoEXvrai2c4dBWivxk22hoLVQl8L8lHn3e97oQ1sEGQMFLu03MLMm1lBPjGnTKB2ZFLChCs+SKQb
vPMsUes8+hhtOiWepiRmWk5+0qIgyjhm9hHywj2gUE/YsZK/UVPe2bUuQPZHqQ2X00NL7/KcBgX/
bBuGr6uvUjMn5iZQFTcXeoRitcdJ36IAAK62PnABfdnw9R1GapPeJrnALzITyQrJil8hTjoYo2L6
rsnfr8KtoKRtADkqlzieoDLy60edpMVqx0u1wU3zFSCokDZzk19qJVslopbtjKS2VJV/tGxsXe0+
wJWOXYFtnx03h32tMSnJ0hyQWSMChKD69xnDx/aQRGYFSCGCc1JTiNlAFeWO5r6t19iCo1hZAXSn
tG0WcDlhd/vChHQ3YD+CYrhOqBySHyT0bQdInBVE8/DCLY9fpDEufZ/1MSoXztTgj/7M4N4DC6kM
IH9o74UlGC29kjisyryOsaJikb9l5qmR7B9uyQdsrlTIt2KsXRff9rfEcP7qE48x5eVRxbX5I3uv
acOxN6ZnHl3KOyKB49Qxg+sEKdhPyVDktlnNiUIAI5yYaP05sOJTK5qIGGxfC70I2QIX537j+NAx
F3piHScV4ApT0MWI77HvPKYSgNltUr9EoRAk+mpDoBqYPqpvGCMFLPsqfrpFz+HU46I2403qHvuu
eUadigWgXkdMiz4JmgP0tfMf7Xwok8Ep3Pqt10D6dGmtOYJzLwxByIE1QrF0taeh3DiitDdczWgS
SkYQSlie/gxIBw/0HDGC0eTq85VBlKlt+uNcGMRnP+oTJrxFRHPyIr8JG3s32Y6S+iDPfQQruD2Q
kQNhBO+7omh6pkFakXssvTCHPMXB0++MaZUyaRbbtvJuqs0/PZo3TaTV0eTOuA1Hry0aqyEhOw6/
YbyYl5i3qj3RDt64ySXy+c3Aw2ADOk5rMkYXQjPvG/+Nm3eQP+KYa16qWUcMFoTTEjk7f/fZnO6G
XF6EJH051Q5PlIf/4JvYy5SGw0MbJ2NRnVW2nVmoi2jrs8+mDnvbqIh+n0KRK2nZylMD6pcm4PLz
RPejR/igujGjmNDoIgTaXkbfg+EjXS2SwGEQpezobzSIkp02QjaaDz7f4BGL5xWVK3rIuFCLmRcs
NambRv+evQ0/h1VK1M6FYHN7bbnzEWVvqJQOd0BmkqqzK7pM3JUlu+bhb5CFPpXxgueAt2fggeVZ
9Fxy5gZK/cL5FyRCKYLI4bihIyjRo/QY9kNPWjGpgZNtEcisrtAMuUKBOTBMu5avQffJjP9JlNgU
L+oDpPCt0din6/N1dD1hGcmJEWR0hln61vt7nmR5tUjanAI6CW6hVckajYFiRIFCL4mN0E4x+81V
fj3jrGnQP7HG5wjLZhIIwTwTauCNoawZVakAku8BKF75r6w6yaYwwe7LFX1aTwJ0Oe18lqGxVM4J
/uAtdnxjf4rGtyL5ex7AHBFrgtZheGT74PGiqvcNk4JB2GP/Lnk+Sm84OPjsvLB2kxLByX/aGOyS
3gtx7rYALdMTKk5f1GYnUJXBsuvHaDyDf5y6oVuSRzUImjuVE5RP55GyMpnO5hvlNSA6oqjWavui
8wTXuXJQIgmxe8th+sfQuxDTpfgMUcqJDqOdBTmsx6RsFSh24YK3LXO4uknaVczKGVZsSaxj8VUs
Pr7zv/LSGFLGq8QBFSR53VmW8RpdcXresBAKpWtyJ63pCJ1oOWaR79O/i4PwXvkSw8uHVJutZM6H
cbqxdtTduB0rWAc3X8TUNkyQ6Xowr59zYq/HesnH676vSe3pupOgUTrBQdi2VMepfYIeUkOryfBK
LpicjR+J/kwp3/QrqoBEYQmJXj9qy24gNJ5MsimLsljSI7ESC/xtKg5G1roAlpCU9oB9YM/4iP+L
8rJrgkD9FFud/Y6Sd943dqQZ9YmMV6Ko9OQkfo8fILA2LsEqF5PUg66ZE5IJrSwL7ziTEKvyMsPN
fsXse5obuxUudCQqMoePkoLbHp+iPUAqX8KfGzf948WBj/pEya/Gc1c8QlLTAqq5j7ThTHR2UOeg
9n3e/9swuxl93pVJf2/KleUnzYC+B0AsC9luXuCSXPLbS42BROV9pAJfrpyq6OaWuWcVLNS1fsf5
ZNEwsrlbztl8x9n/yVOHMdD6cHZ2eDTe/7buU58M3QVbl5+n0GQhmgMiFb/gAbSv6Jo7Q7H708ej
WuNND8lKI5TwtghBC4TXMMeEEK9w09O/VbUBxznkcHDOTfLQlg8xxpODkyBarveo/Jp+NWUeqAaH
IWxiRl1WAFYGQUgYhwZQ4+CogLgDZ0KOVIpszZzwtCelfmwG5jEF7xIXGDqJz8k4R40OpEWAZfjs
sOBn3YgaWrzN+RnaQfxuB0LLKaNsZZtuT/G4+ji/48G20UNqDP5kXJuB9s4DCM1P4f69cqz47+IL
0r27nuAh7AkzIrUlydI5OE68dzxdW6m3iVtwpdNhaausz6j4cp2PoRPbOE1wc3HaH8J656W62kCF
sU9tD+RrpV4jMbihvm4ZTjM1oMf4c/+8MbH6GO6skHrQvtiNWlFB3+xHMfklb8B7/ZAgfrcvvBB8
ERZpwxfgNAofIiFHmJhcHQkPDfzY5pQ0KyWF2E20EKn7Io5tX3MF8c9fwv+wXv4W3aAn/8RA91uR
cs6cndGsCxCmKKAGlxE9ki/98u97N8Lf1M3BFUfCwjXiyOhFmHgKGu9rtyg54YETwqYsnmktwFz+
PlWx7b6c/KsHuNTcWqM6hnAaqnMSHKmhUOt29NeHiQ6zjYDdjTwfNC47N2JJEPDhS0joSu+cyqRJ
czjbV7KQy6w/qTqKo6SLoP/ZF3yQzyuPVJdlipFkoLrnzWU+T4OYqZNa62R6v/HWM5QVZi50am6r
/e/C/KhogNxV2/SNNdjRpQDkO5G/rfUWszjoe82/wwU9lzjQbOnF++TihB3IVNd2wHOgmqNz4Xe3
PFnfGwG9mrwD4kTsGF+Y6XhMoKB/JGW04oCySLD+01fqtM4dLruXkj7V1QH9NUlMrlcTrRz9XOZX
xtHnVL0U/NBo9lc1ECUbOVgOpKs3Y4GTp8Pmunti8rZsGAuoXLR5JBIuLe1+3WP4fLP1QSkSVd2V
dF3Kk+QRspSlrKKjr3hcmBJsqcVZ+upt3pM4FrnfxNfuv+1y40Y6HjeUSEsXzSI5URc+VNHG2BQh
Ayuerjz8nkIVjL4yL9aS7BmhfR73EVHTfcmB+D+puit3OebKd72Kxu3slNRdu28TYv4p0lvfuHgS
YlM+tA5PipYJHIqIwoYjlzqRBR+Hd1QyrIeTC1VevvhLhkavMWi5+3HwL/ZABx6AG6YQtOkn1aOM
gzFYDAxdTMCKdzBHW3FtY3eSVk5Kuxam7z4Dm87I7gg3EoCMAFPLpJF/CTgsFIqfIWhQaDh9xalo
vG4qc8u0S1YwdtdT7Vkm/fjIs/tn9D2nQTX/8HSTp1fP7vcfo+ybfxGzOpe6zj6I40/sgMNYYjFV
BJtPpMEt0L5ziM3gjBDAI2JU+kNw+ek8zqFb54DtGoZAWhr569428SmiTdW7YrgrP6PUe94z+DZI
xwqDeQE4RX2pntU8bY4d5UyY2pEQiKn1bxIVhsQTq/h0ceyyhmC6KnkaPIie30i9HVkxnXn4sNSN
a9FrcsfKmu44IWmOaimvOib/BzUenoh5jvnS6UAniaecdMW1Q3Yms2iEsAD0ZZPQ9HPJbS5GYfU0
7PWUEfCUSXofxIlHCG1a5UzaS17d+W7zOEVZmHzp8XkL8YoqPojyCp6ta12p+4HJ8O+P+xhj94bE
XytRfUI5vXKCHwkXHehQOxiaB6jOeCvOjW+BUtBFeZcYwSGpCw4ZQOYqNbkYEDjWM+ScdRf4pe66
zqbJsKmWsJlyA7E/rvO9HtYaTp5XxX9HDj8yvkzUpxbZ2CCGUVwseOu8XtgB4+yxQpT3C8zL1TNx
LeOCc7fEmxsL+4vzK4H/HAQYZIIzD9l8pHBCE1QQLt0Ab8V5ABtb07U96fLreYN/N0CNfJpbtkuJ
1IItgpyF2UqiK86Sx+y96UMzzKBNRl+vpa0rCzgIq/GIZfIGPUl6+2WpdEi4dnbX4gAmB/oeuu4H
lnZPstvkoAcQIsiI1mXOzAkcvMxrRZoZZ6WK4GVN1H2zacKPYsSXjCOZ2yWuhBvUc0+tF1M/apg6
bQ8PJnarisOeG1B9YcnH4GtoGLf/CIJlpaXbcI/yq3OKMLK9Nq50dGJpXrqAKPOnO406NgWtHK9l
eqeSiK0+ZKMfcXpY2q8tCjhvSWmegVLYfavUkF6cmfzo8AkvE9t56pHxDkDkIZMqVMpf2HpvUnST
+BJohURNum8VLtb8okJ2TwIaSUtpisn/e4hSezkcjcwVGa4cVk7mAeELBV8ckkck3IEqAn1cQz+3
81i1P/dfzgEQA6T30v7KjiwPBnCu+kFNH6q4dJSrP+HKTmR4LJpb8clbDUGKrgFPVD6YA89t/3gO
pK1YkCX2H+yTfYqf09S7qX295GSNLcpsRYDQT3lV6SShRiI7tyQ9bBbv67AV/i/BxKDUB5bqx+ux
K58u19XJVWqX5qiN76K9ibpWpog/nlV3aWtL64eFW4/h5t4Q/LHaQcC1DKeRLwY/wRtrs4l4aMcY
ug1gFY4W/f54NDmuu03UmFSjxlQlGIhuHBcOVhCaGdWq7Jmgj3BDK657V0KuAMbulQC26Tunjbav
Lmq7yVguQFn9w2d2PC5suPjAEZzfInQSwolGfaFWdLJLqKEa+FFszxVwYynWiwYmdKM5MJgEmZn/
TlGQHYQ3hlevo/1bnQfKZl4zVR2GlCZ5cKGe9sqnh+3bsIimyYSXS7OkqfC+C03AoEoF1Ad1RmDu
oMOgfQ3Oxm4x3YUyrFS5CZTng55tFyML3el8UfLjJFVFi0mGxBI3neiApEiSvdhDm9jmlhE3KsSg
Jw0hPi1TUvWBky57jxZUwlZL7nIFRAbDTMikPlUmvnFRhKhqyg0OVkQAHUUxQ2hZDE66ZEc8NImH
QStRCKPJ/0wBsLfCTeoJtlXvJz6S6+p6G1UWAuwbVRWCqTIb2ZI7mH9OVaWr7KSRx62qySi/1sI8
m5ZB4CbFgmbW4bSpEjS/kFH89faAYNz51Yvz1J9V3+VRFrSNIAB8M4UokJTWXeymp+JXPA6ESJl8
V3daqGnjGeLZghhGx5UMDO83JUHUpAyEu0cSSufcSUr339vm2MFOrouD/13ut2q7PCCaz/zaJ57P
LKOdeq0fBU7QvddFwjWu2OcJdDICqiDc7IY0rPr8vYvtSv/svEZnsLmjSQWoOA5IKsrn2UD0lMOl
8nQD4sR1TGskpqYm2xfDjOOzGnNVIfhM2eHd+dekgTHTlRzA+KFtz68kUWUDAt8qniRQVPmFP5Fh
vRhddk++2Xi9+Rlro0+4Z4o40qs/CaJutQXYkH1bezGDLoETpauJSL6P6ZFs/7kNPYy04K3fa/ue
k+uSCf7vyiy0eEm1PGX5WAqRoBJFdpQ8cxkCV4ao6iYZUleJ5mQixvvj1y5+jNk0STndUsVbfgmi
2/ca8N27tDdRLwIc088Oi9d/iYz6exmnodADwmrjFR538bZUbEzQHBKEaTPiuTcGRFDndqFI2rep
7/YBR9jBVjf2yx/oJgcl7EM6fe3tN6IvdX4O73SYquuy0WcxB0zKvPt17bE99nMHnoXDwGRVYJCf
x5eeoEM6bm+HCxbtlFr0wRpVq9nFLh7kqGbvhdV9WibX0jSq0mv/+5ZxeXc6pHBXpsdEgy7eQxmS
7zEsZZT2Bq0v8c8a5RwD+IsZwp2yppyaVjwTLR0+NBnYfvZihn3N2mPa9mxKOPlOjEcg47aSBMqM
eCK1PmW6Sv9FayoxWZPsoU0X5ZgYKRaw2NVE1hkRrySs1jh6w/Vp+agu+3qRXoRdVhitVdeWVGhE
HJQ2b3VbroMSpDta0F7EAiEOIA8m7hbKajqV/XAmzsKS3yBU9yV0dTMFj3mO67a2UPt2djVy1RYK
goE+fcVGxrVLHnOXOhYstKhwmY3NO/WQYTx2ovvcIqM0T+bOPCvX7HXYzBr5Nem7OcGCCN8ZhGxG
hE84/vjbX0hgC1ZM1gww/bXK8Kn+bCCPDU6XZ1ntpR74FhY4ECM+0EPf8HDK8WHXgTHFF73hzspp
I1Vr+GzUqCrcof1N+kdtamHwmuXHGjXwTOGnRxB4eWHG1P4FNpgP9gDU4UGrjZ7zZWgvjmh6f2Lf
BGSonttLByJhLI+X5gaIlgbLo+3yjY/lNIupvghhjz/LQfGF2wG/tv+f4Y0qAhz/D39eTlmet9e0
EBH5WiU+BDmSPjsbytsfThGEd7gLsyrB++HNFr1dfW3x17gvOlNId7viA2rDxVXqDIkkgrSuznpK
Be2wMUPlxy9L4keCEe6dkMhFZEhUi/AFgc/GVFxGvy9acY4PGkXCQ5mcnbxxlyM25GNuQQ7wYgAM
EjvMu1WIpVzCZgh566U2K6ng0Czm/AbbZwBJ0feC26taekjjnfUUBCNfMsFOTaQJSNF1nRZuF4ZR
+Cjp99Ny6FzTzzQEUuru5LBwQ17AuImppQa7WCsUB8TYHwWL10OEEKUKsaR8xBGzPAn1KlNJmgG9
50rG68xk02GZTCMxhS/r/V6R4MZOYp+u16TXASGrhgdYYSBQ5jleXm1lK54AvZzTjt+5m3gNlY9s
niUdz3fMuVsnBSpNX6HCeCICW9pzEriHHWyqscHUNJmULRXMovjZZPZ4qAnKAaMP7sjYKt6feacL
aIUJ+FahSqkOUsswqeU4ub5gNUGlutIq8IRtqP443FlF/L6s11ibGJIOAB3I1BoaMrm1l4F5b8IK
SSApcOI9bhksOGEMmGeBAhKfVGo02xaEoY0DZLYIVWcpBKR5D7ixfRJRzFDe0zIG0vaRmGN2hgWw
v7ZD4JMdJ05uMCyILWOe8uKsKHfjUVpnU6snN4joIjCVp8NUS6c6lYilnV5vlMN/dDVqOpu64kwf
aOtY1p8kUULapI2E0tvT6gjn8GlWVL3AEvAGwNgnds8U6PlGpRsiC5igFHZlNGKJthwwpBhiDDk2
TIWI1Vszy1emPKpoRowI3RvhbhAZ9f4OjcsNh2LjE60clKv6oBkbNY7eb3N8RlJr/GQzGAStgqs8
Iyquy5zF6P23hdsqPNbcfl0qodPsGRdlV5k4TJqKZBNqq/TkrbiKpnk+rnFhBrrDBcq7uZnin4vj
HNQ4cWUeYlGg8DAqLePxvzH/r8KCR4gS8/jfeqnmIKv7KUeUCsx3kr4nmmc6R3PMT2hV9SmZPeuO
+ZdPjhVSgTEBmR9wRYGgfdie2TRXdzBquux70gNZNS3F+UCGWlgG8uiFEt+xpXWPrEuWAHjv8xlf
DWaj10n7w9Ifsc4mUVe+XGkEIYnjaE7bVMNVfqBoy5sM0uPGuFIGfNAaJToGCt3o6eMur4fnUWXe
A9XNrAbRM6Uyhz7QOGdvcHJ3p24bQDWiG5oESF8JdgxgxZPwaPVlBCifxn1LxfC8mfVRXbF8YXFN
tOPVxUBOtCq56op/9xZFTeW+7ruIm3Mok9N/ozxrttZ44EBjMnRY0/p2TtNCA1aIA+wU+OM8jYkh
Offt+zBoo85nP/Zx0lkFwLCYscfxgPabaJTXJ2LpWyPhQf3SAboofPqOgHW0Vuj9HuHQowKbBLkE
GkM8r9CTGNPiBgVm9ta6ekbd3pCLFdOMjPu02aXrcNYHVSwUK0hgXqkCA34t4vixqFJc6+Qzi/PX
L/GiZ2p1BXehm306oPkJTh2CdryI+Qg/oJ6CrC/fEJBwXzynN+QBk4nATngJmFUokMQ1JmjuudQG
YvGb+O0oZjmoT5Y9AOAGbZr7oHxxdTf0n09NZDp72zeaFdZbd5a5tNz1NW3WwOGmss1PZAU4abKA
adMVLUFXENkWQfrJ3uVTMiH11sCTiumxtyHRkGCEGPYr8xmUqFPT6pqu0b/+W2SHAMOpxPVBzs1j
Xwmgz+r+BM5NCA8UNsgNSr2zqmkARZtlM2wLDzGU0ndMnFm33sshwHeUDe71UWUnydejbzNrzXJ8
Lg5ZWqtWoVPo/lplkMYCLQLzmb7ChpEwkR5Ra0uZ9OphKeYqPhZ4TTDoh1huZs5NEuMNLiv2/cHK
22RwDelGm7AwjY/5oN/bYiLozKzDVXN+nKyiNP64RdEgtfkk+TczIU8eosZdA7jWpXVoTsPkiRiK
MsuAPeF/LBlaKxx5jyuUVnWLTLVdIt4DYgX6MysUHKFIU8d8yvlIXqdO4nW0+CF5QSav2sVLq5FW
RyMRk96+W/P6+FGCcz+2d0370ddxlAhcN+YhO+5GmIJe35KedkpQw91DCaa9DPDMgLXwdilBCTBg
CdML2VBnHumOLyJAp7Q8rmsX9QVjjSU7ElHqBjTFTIpuRT3U2AlEaDPS9MBYVHIUMBdvJaNNhg+o
nKnU2pOiaBVWfsP3XUZ9iTZSJiQwyeFbz3TVIYDn7cxNKPIqwTjtBZbJdJ1KztL3qOL5+hKiRZL7
u6H52v0gWYR+XDAeyvp1aS5wgKn3qKgNpxU2Yli6NV1WFz+rklK9Bp/Uqr7SjayJy/wdn7BgcXjI
3KbZgp8v+B1H6omMkj0YaBo3ivXC+iGfK6Y5A49wjfaBvEcTJojSpCbRPEoLpDwZMHzzx14j8HSQ
u8rvsu7JTkYRrRssHTWxe/LF69x11+XiHWhRvqZmYTnTMMkBrZZqnMh9bYbqoOQXcALpBKJL5s07
DvjUZ6apMOWWmT4pPR6uHOyypBNo50V2Zlk170Oq5aCzWuheHIG9xgxD5HyapXn3xAQwLuI2SYbX
zjJ7u90U8ahRzZCzjEky/GPy84uzN+88Wa8VFTfIK7sq2knN/VQfyTcYekAiD23jqgVOwApzEKkr
T3KDTlgjsJU1ND9mGi9NiKUzYTa8UNUVEMHwrQbaaAJ764OEXRpdVJ3br1ytjsEaDFD8I7fbkfgi
AV4g6OEE50z9/M3YBUSNQjH/5nzpUwdu5Ek8i1T0ISJ9gFpkaKRtrRIPmIlRSY7/xGG2HjmVdQV/
qr0GZlR1vCAEBWOrRAC0Cb3UuTVo+hzwHfRQM4A1LOw8EC/Zz3e0HmVsukBP8WRvWMKBze5ChCIe
7VfgeOd6hcI3EggPRTpHfk7WL2ZNXWYQoGSTkANG/bFUq4clJq/rC8B6n2awBUIs6NOWtfcv5Afu
d8BVdoTBcQg4puDN4jLnkpRcZx79HOYXEeO6feWaxExDmBVkJanRSd5aXGEC0NmetQceB2eplkXA
9nqTRXkLq76YEk+OCfVwCEFCSKQxhH9O+6kxHBW5hv6dWVujMgl/uFPw1eFKxThtgQT2pAlgAozX
QCqAb7fYdd5dA77n3iAmBYuW5FbZX+mvSR3+M/6GlniHXIR9gIBnELBNaGQbkyohgC+qPOpXohiq
8F7UbZ4e2OpQXF81JdJ5meBnO6hUSXGTbKrgwTALxTLEBmv5TIz5GvpltptxfimBOvZ03nrbucre
e7toAZcRX1B9U7HVP/ScwQ6da1x2Dpm8RHkPAf6spMiUjg8G9zFQvcS7uQp0l3kJXdHT9r2yF6fi
HyFjaQkoLPfl3ARPENzaVDr7PCQtAL/ZPcEpa8onS7OPEpxT3OzM1M6wfKdQnd8nHba2NA5nCDVf
nvlNALKfmsmbAZHRfLoGlLoMi+C5uNNrSVivrkWKjPrK7LAHK41BLHzQdnLTfeaI+aS3NqGPkPVb
ov3PztbHyTrWfP35F7gz/cKAEIgKTPAGKgVeTeFfyRPsyV3iN0FGwM3ZPP+98NPjebKC55MMRUNn
kiOQGBXr2Vxs+K42LhvgrA8Pgw1iy01/z75xFYvl3xqTyL/5dvkzoPTeDbz8dvdPwRT5rIMSdcH4
1xq9dKLuOTjh/YKQ3lZlcdmhoTDHvAm37hwMM0LtJw4bGht8ZAcW5ZL/nZjb1tqkiVA9JLjYFflN
aLth2ca31n5P1Y5Z8BALAvGFaGLDUTS+AlBjb0c+RLE5NiynJAkp+yJNdapx3ISyGp2btCON9Vj2
vErVC+zoAlU1hQy5c8ncSvv37JhAhLh7m4j0IRq2r/0WYHWiwz6903swHzr7EPpimQqP8/nPC1ks
sDYCOeSbblITgGMCbQlqGcz2VrZujL1hAVE+QOdviRAdjnj/ZfVRWBbn60868yfRogsVfVBn6nXC
5QynTgMGkg3gGcuTuUo5myfDryjHFym7RX5xy9SkvWB5ux8L2zZ9VVzDN+zk1dTdvIkWspSKLP+p
voX8EGC+V4l3G/0fgKUbo2mU6a8xkVN5mPPtU0rMKByh02xzuwtvujGWUJ8pWn8CqsioaCED+uYT
oHyLa+ak8cxYjFXYpLlhn8PxAtF4nRyg1IgjIMXTUb+9HAbrfNzFSCWvCccKVmXysyMJVNTGk63R
LY3chb/Vz68P5AHqQVr7hzGrZuvdPqIH3K+eK/nt0mqklf6A8HDUJlrwN/x/EJCxJNE1+5HZtZYk
TCzcrYZZTJrFrG+shbsYcFc3a8nJZ+sETv5oqr+7BIm96JXsObGuvTNluY4fPWvJtuLVd5UD3pBC
ikisG0UIpthefiHIdrX3ghuIPuQsTrVC4OgXbT7FUAcHLuBGBaWfAaVRmOP4pJHBmEJzCS64wEww
w5DTm/hraOH/jze3svpKpUI9sQXFGHpMzCaT2aG54X1cod3LWrm4VdZRkkw0aC9szlA38ayNEsmT
APPdfRmj1cIxbq3t3mZaYSDXNNZmc9xwU/rlRoAoNlz2DIDNt/sZK1G3dohgTkGWe8G1FZ8d6493
rfG5DedBMoHTkn0zPgsg3b/eUgzfJZbWD/qooTFQYhn6KSdw834QNN7hN9m9iKRItobNJRLi6Fyo
SZCXInQ/jPD/jc1nl4YTzJj9pPmsSjuJ675ADpz0G8mGI79WSCypd9DjkYurQHSZzQGKGVxNYe+u
jqsZJpWSi9q/CoE/80AGU5lUfaOCLXZmQUeZ1sYCQBRst8xJ18nOZ0awiMQvBm331icvGnEQEBeQ
PF8wLaz9NeZ4o0Yx1eDipAN95lKA1qV4WEmhplcQh0mhE2h+/WzHq5u32CiJePGPpIY421ENns6N
3Q4dzxsCPBHsK4W9FPqVOjQHWHHbwj1zUQSBFx5chPMkcKqYRrlInS9Qc/l9tDivf4xC/quw0wiX
4V2xc7jFIwsQte9t0VVRdw8PCqAp7VKGZw5dlaIF3B67+w6moudJx4bj0C/zYeeRpK5oVu+oK7HT
Srec/KSEPBn09ZF14VIA/omN8kJDZndcEv3VViNMI/oKX25JVCTOv7aQs52SShtAIqw/0gidUIA7
woTWT6pTSXKGfU6p0AVbm0HoNg8VmrFf2FkTI82TDfd9MK9hNqmIn5EVn6uJbDzbBxyH1HUEHPhl
OghVq0hi3K6/ORnf3srqrT+Dn2avUkGnLtBsPFrxwGtDrpQAiQioGlQ6EjMeJ4Dp9PYaTJPh6olh
fxk/ri3ovDlY9uzR5BgUNjcPkdobRqJvFK5FCjjVLpmMzLC9Hf00zFsIoAfFYGtlyaKsTSON1w9O
xFlPzXrlfmzSxKCcilUnVl1GgUr74+KK1SFCEP226EKT9prphW3yry38JJ5r9uktaOkbgXhe9EH9
Y4xCV2xc+uHZXD3Qr9U4kNYuvexKDLyxyhH1yqeFx5Q1PtL1xIFbrz22XLqoVVgoBzYJ+07KTTH6
0Wm+a6Ud+lcuswv43L389cvawZSnrTYdYuuIeI42hO2EzVzNvofY+CBtiTWrRC2TU8n1BIzl65+1
bXClXI7a5VlRITXZpPCDQgu3sSZdufc1kA0xJgsy4U7K8Rxi7HbkZOEvZ//SXUVsHkWAwFhbc1fD
aLJU5+sH7+pcscHwVn99yhpJ04BelC8xpHk6xoCxja/BB2lQYEvGAZ07Dg95DpLwg7eyBOnXk0XO
3MYHerA7HzPe+S0OQL/rF+qKz2+5gKhsc9tiOSbgRE0By4hcdoKk3uyKLtChmzQ3yk3KAJLOCFzX
vhnDOYvppF1xMxuL6J+JvI9re9G4TJCGkr2DsdRDR1CHyBNV3nGqnhfzRUQ17YzKDxlJIFHk3tKN
pSXKj4cf6VdP4C5aCrmhkrcWOPz/bXNaFl3eQCIU/NFbCPoteyP+NGKJQThhAPvSkA8g1ymCP+pb
VTPdTPlrBPlUfvM1PjW5mp3fgPR4/UljO7iECNwyfyo+VKm1vLWyvz2pXVEXCbr5JPOhekADfCVV
mnPBm2Mbv9Sm3TzczX3Vph3XmFRPvBDmk4G+EAWAIcOjcoz8BWtPc8AsniiWeoA0qPqqCG+FzVZP
qFaDxgc8oqbjdSvJPOKP7JmKvKUtDCBsIBv9APbLQ2uVKM0oEjMptWkaZOYXVpRLHNdiSOhPlb97
QNK/AuyTmnUO8qtc7/UC/EipyP5SfVbzGzcsE7A8zWnZqLHYMOGVSb5j7tpu9A+d31proP6eUsM9
0mBJFWSXTM/AWE2D/uQx56o4SPHriKe0UUtATdO1FTvwHOqjBO/XAwD/wJbzY6IzZ3Reej3bgahf
3OKzO/ivJDHutG8QlNXBPDCpRSSFTLh1f3MxN57ghcciZ0IZkdZTIq8QG4XSHH8MGyAMSX0knNyJ
/eL1lypj+vFvtIMHZTIeuePr/v28SIOmB6mHr6R+8sioAsIjF9A4cO02WcjzVItGshS9xeIIYnkt
pavBQMZ8kHaYWCCWhuy8ZuEGsadp0UtVoe1SuuSubtdmTLG2BwQMARlfow709L8c7FyZsRKsgHED
jpWAWvPdyE5V+k9D5ZEaiYVENswcXEEInn1T/Rp7Jxt6rl2gNze+p7WvoZBtpVcRTCtWhsMWXL15
5jyuiIypdCaRuyWPJ2MQzXcn1U2MxsGjNGIjpAgFJ4vKh3QOkpl3t5i3bQRzfANURZlUqd222CPO
RhxZdq0N/1mUFg8KpNxCfLgNGF/G02i0nJejnHIAY2YPwpC8jfbJgmeC0VyZAlcr4zTCEAySUyIw
hBjVlCRX4Fr1atcKcw1gvbozd8nlQUFF6t0Un9tpQBC9k071WJuUJWx6/rULiCCTHykR2iCilRE1
gNOF1z2jHmrMjDiF3dP40I1v1j0ZT9G++ApDHIRlvEbDM02dXnVhwYHONHvbREf0tBmuR+MVIRMh
BuqHdJ/8KPFEVjQ5E8anVx2WJO1nL9bsu3C2v7ql4WTYU/mrIQNLOPW5q1KdTx6hp5B/B351FGx5
z3RkYM1bmtAVJb9NS7DjavWxlGnkSCUH8hGdStmG0YgkMU0i3zbVOhljLefbCISEjkQuP9lvrbh2
GvFelojBWDZ+Bp/f9R9wNH3BAWyvV1EWpRdsr9u26ZxA/JdE4JLW9Pt2HzUOORLKbrqD5O8hOgOV
vFtLd26eeX0v1NTMZFWwh+bXk6xHMwCsIJt/nx+1TbyxxpPEhBAwkCK9oTJRU7oFzfEvZcZjrGW3
bhN5rLUQm3STvDEJj9CLJ9zXW7LTayWtbMEmdcGuyt/GN92r0tG0QiB93yicPH3ARp9QYi0Umvlt
vE44OWBuGD64Py3Jm21K63OWojfoLRnWNXBsSNP0pXzoCC6dEToLNuQhOwdwnKRSfhOcsu5SABLZ
CQ16Qb0o0pdYLnyAy49HbqF35sB2ZKX5YESGuDk/R+StyMx9hI1hUwtNo1joSME8NpIV4hTUOWfE
xqwnlvZdK1XWktYV6E3gESUI/Kt7qisrYTbwma9j4hFEFpbFDgQNsYRoufG9oEBDgN0514Yza7Ob
pyemkx1qVOWWnDwK+YOdcN+81uYdFn7qi1psLEELVUMnCKMfkb9rThc0pq34m7wVOcqPtqp6B4E8
qXPtNrBgUfB9rAry3s99R/octi59A9Qf4oovp/ZnFlHB+HPs4ql94K5FmnI7009s5tNSz1uJsQEZ
L75pAPzbC/yg/nM4cIINHvnx6yJLJq2ytt9Fi3hb1j5/kmaIRX3VsVwotF+JyNDcjO+sG8iu49zX
a5nmMMr2gMTKtcmr0h+SLOsw/gY7e089X+mzM8RD+H7DLnbfXjxHnQM9gfyaKm0GfQhHsLYyg8UR
TYGkjZJ0pvxoUfQ8q8nvA0oE30ZH3XPX0BRGxSLaL/c670dlznqwjKkNaXZSl96ueC0PsmiDQeOt
m4DFCtFSE6ZxTtaMFWu+f5wMQI8fg77sBLPUmbL/9nTcPKTEW195TSD6rJD2HEeO8rlHCZ5/VXb/
oI/yxZ3FPJJBh9GDv8HtC6fv5JxOFdHNiAoJtfiOqgW/R2KABtESlOTj+rMQFpT1lPDifsCzjcIK
BVcGHzQLarjVOihi+NSIBMuN/fe1j2Jku0n0QISVk5+ddGydMTyE9zmL4tuqZLKnnWJXi895FexB
E8UGEWKmzFsL7KHrTQWqNtH+MoPznJhMcXLD1zKT5kiApbCHJAqPrh57iSIJiweUJA9g2mb+wKJB
mqQNLe4DTvLc9Alu0eX0Qt0cM9j9sQpGGwHJwtLHTyykJdLJJwuB9DHCBR1sjsaZ4aUl9cKCA6Ll
oXyPpZJv4LyCvNXplf3EhVNE6cFFhvR0XGXeItbk2jbBrPaeve1WLiZ1lACrtribfAKG8qgfPW5t
5/BNSHm4VkdtObMJaw8H/BSY6B6dPb1ZveEyevui5ly7qjQ+NDm0EYRzCSC4ShenrY7GLaock6aa
26zyN5Sh4LVg8O8bmvrZq5wHuFOqgHMsd/olE5wyURJ9JQ0bKXqeC4H4nY/Cf4uCT++HE3emto8l
Pk7RFQ+CJy23KbbOyu3dk2TDm2BcMwoaKfCrKQZekkB1/PLnjU7fUHViBGwAw048rNfkO1BLHFFx
dZ2+w2qgbocthfnnoqx1qkUGasIJ5Yf0HOVrB/faf2Knp9tog0BjXpxuVdMLmSskxuP9T7o677Yt
LhjOjPo0IOaX3mBKCvl2GlrfkJ73ZFZY7FfND0KYrI7I3voJ7zBwP1DAp9J9/5cPvgzWWM/4Y24n
/htDqIcet2wx/OA+nGcBAHew7/mEwBaAod7W8Zmji2Hh7Qt2WXrOvvOcBWWqgH6bCk/+6lAm0JLT
9aCL218tEpZAJFjDRiiipHCDcp6HFnJ+mZdlKdMBJ959Gkf3X3s+CaCvCinaB3i7QFg+gs5OiM4C
ZTgss4fBbarVPYMpz8AGCAFzKKbfZlSTvQbUG/siGIAUxquEm08XpKrwC2/U3HrCaYWicSepWDmA
MlcGR0y0zCFdDWrXMfQSax4y+jnpY6zgWAL9msBPYf/2lMpDdtv5UoTCMdRmlp1qgPGddvoHVYp7
RcTb20OuaRi7EFs3FJpVHbQm+xJY+yKJxlEPpvZuJVrcSNWWzMMDWokM5eKsdEDLHSb0UkA/vYyM
iwS55eE9YvmHAkgBEIgvIXzLPqXk7tzdcC0N+XFcF20x+SgiiVrySYxjrSPauIy9jZTlfsQZU77D
eBRPOT0a2zMkLkUwQVkJJjVbPR7LD9BlngLCaOX+dKCXvIf+PKVY1JL05A1aPAzGjCVXRkFCAYPW
Y24cL5BCx9EU2vXS5ETFG/V+iaBd0kSzRoulNmE7WbfIj+YQGhbYmt7wjSyAizKN+a0QhIsrQB0G
5H9MB19vpAXS3I1k6EXOQL1Fys/EpYg5fCs8LNsjiciZ7P22QynNVdTYApa0xMVNTkoQKSgH9/gC
y9tQYL3Vi9XlGzKIXJOtHhTuHnhIc127VA0WHvzGoJNn+wvTgWxzV/5+cZHKpdnrV224xHCpD+ht
UmtnuCcWC4v39HU3kbG8X7a3OTQszPSCuKfxzx4WG5b8yg+I1GdJ4mLEzQg/09XB3mEftqUTfTTk
kOQCFUT3XlOs9i6aypL7FwPbKLR/IGvolz1LX6VeYA2YttgL0W0GZxcwSVKsLD7Jl5Wa/SnPDEIc
dhzab0copXPYSKcz7oPc5rTTKYtQBVmoMXdobxJ3Cr6PvQconhii6SsY9kDfSrwYFQLgRGbpv0FT
PRw2x0uZ/TOhDNmXOpnXbIpFQ6BJPsG8oAmabiIt9lqbEo2CTdWi3jeZ/HJJvlRZ2QAMNt1TLxph
zeDiP5qKRLtoBH2aVz8Tt7ShKY84VTktumn4Q+yAqc2ck8rvQZxJbf+ONXQgzSLXASyf0QPhm8hk
BVJfIFCuGgJtIP2d9ofcogCKSSe19qSKcd2YEyCMBuqYLyEVh+wYQhnbVWTzDGQwe5MXFEWKjdrw
d0KnViDSGWzwJYY0MVWnQu4eiCsYZ+LhZNo3bi1fjlUr48w+b/L84Yr+Zn453ukbAhBGPCs6x/qd
C+YqWa/uILB1xhOXLdo1wpyNMex1RcLrOllwxUBE1FRi9n9sCD3rofkXrULus2ybfC8GAw6rPFEA
VTEI1SfhQxkRCAoUwNlwQp5b5rQq+gfWZhBl059NPrNSo61dmU1Nkd1yAwyTb9upEl6VctbXTpit
S3Qpdtan1BpY5pZBWI+L07GXgyCsrFrljzCW7o95u8v5JpCGpLywOMEI9N9sBuA943yxA7lh8Wei
eBTuejcEbyIpE9SfBod7cha1nF1DwspTu3+8GoeSfpwQWBpk9VZP131qsgUJCSdWJL7XBD8cUP5v
99F3Ozmmk1kxynawyFxBoGEXBrQSjZmV+LS+R+YlO5Ncpmdm0cnM7DXPYoi9iOYTyvXAox8voGNW
kTQgVPZ030Em/W1HsV9rTRaRZJ6n/ryBqZQnOFoX77yfyeSFRRD5Go1WS4XvIr1gdBqekEwWmGvf
uYv0kJ2e0+ZebqPJMxSUrIzwjVMKib8R790yboZUgxHaB/oc4wbUVXZIGV+FWnzQP5PleHQx0io5
sWuQkQrT70X9jGjv1L4ZZmngGT6YPtpRtgmzEKXijJLtOpbquytFGi40MS24MQ3Mur2HRsaUCtnf
JgFyUVpZKv0ZBL4HjQwpgcXSoO/li/v6n89eoojgr1QNpVTSTjlPK0TFuCzyG60fnxhffFRVLVsm
OsUFiKzk8Lw89BhtDlWd7QlzeLFpeQuDnsCNJSKmX2U4gafoXBXilIRwxbgNzgFzfpTjWnKpx5Kq
4finA1xyRdXNZovv1Unp1jIa7RrkVxIyTSmUqgwx/w1ssTLDLLmV/ONfdgI4mIVomUMe/yzenM2q
DOQ8ur8egcewCJ6zHxmW14Pjs3TByZiX8Ofh2+gf6vhTQTtnFxgCkQL89tXckQaeDj5Gg2rj2CmZ
+crdR/dLNlTbmby78oQsygU4P9QgUh0EO0uyOHlWOBwW8rwGSsRaogEUg50GObTotD3SmnxHM0Vv
9OZCbM39kt3312JjPUOf8NezxgX9K8m9exH+RZ+6B7yMJAXNoia0cExfMGIy3QDKbTZElkgzGk+G
TKxPuGVVHwxVWxKLTYWs883EdTPi5pYmoCzX5Xtv/jZG0FC6tKwR5fdqSW7sdUlqrXVtntMIQlVY
1CWfatBJMOzCvT1b34ryPSYuwSlFy0YBKIbULYrUvDG8W5+ZlYubul4j4VbE5HGyT/0cc4MO6jh/
PZyelyF7qqT4kpzTzj4TLfzihnLJsTmmWVrhoOUZV8bSLVnxEXvg1TOtf5O8F6X07MpGhDlb1BG5
1Og7ZXthQ2/MTKfORtJIewPIxyrEpRAK5YEq7DXCpBR1S68bZWuuF491rmMhXIvd64Yiy1eK+HBb
2pBBzUG2uF0kOAB69yqtufWI6KYfSAc8Ne7fICKdZpFqO++gNJs5bsntqr9V19Utg1UDvmVTpzYl
zr0j87VRiAPK2sLdQWMsY7eLR3XdsxTIOKVNaxVakc+tld/CgvQlzvyJ7gTGN1N0jX0lDYfL34dH
tBkQGRf8Rbou6Y9313CvtnbOQLUt77aFVfQixiAE8KpjFhT1gQZoJaLj0fChxEepy4YlFwmae5Fl
DCnOdVHMtMWVSBFPx3ppGeYleMWDv09n2qUAyQ2HIXBtcoXNXKmCxqgnVuWBbCsLR0k/2vd7sdpe
rHvx6g5fgKRcZii1m0qZhILLDp/uefNYF14GorqSQ0Spc66uzzUcnnYlxewDYpmB1PQ35LiEBen0
piADHHwINk5OvkBi77/VSsA/fJf6JV3V3Sl9EMcM54CgjDCZ8TtA3D6kKRHBqBBSHtAEesPPsoYa
BsifKKWu3JSQVsT8jphoJszXGNOPEggjumoPlZnqSu7glN4cqt2RE8OpBPvq39zEeQ1pIvQJaI98
eOVaM+PTrb3yEoykd5qbEmlKz2hbd1hSouX/O+yOncdiVIm5Ded2RF9myJUU5p0/y1sQvjxN0kby
tdzaBsX9al7+/jHbIWSnbAoPyFebHHitJQOLoeKcRbaxMHfAq267bGoJB9HFldrUv6fOEcTDniHe
KCf4m7wyWvPT5pW/iPkJvMnZyJ+e+sNv8aSHWA10/Cf2gS5sha4KH2o0prsi4I6Zb1uUyeMhi5SZ
G/0Er5sfH5Qt1SKa+1mRVoDwQitXadkzaA0asbspfgyWH1EoReA8wOkXbo8yhXZjvaKTEY7qpDyb
+UTc2shQIegyDBsb7IEb6qz5BrJqE5+vFA+BdZ8BtfKTWYOVE++28xOYplK2q647irT9uBqCEL6u
z6Wrye8H3RWfcz9bwFMKMKbbjE/04vglXWQdK42ppeGLjEmUGv+MST0c85xGsaBMinwC6WKc3Oh2
ItefjUvdVKOkLwH0Axfs18FotDB28BJ2D5PQET3STmHE7SBi/d0rDdQrNjU/0DYpbcVHBmWxlzY8
TtyGhYfYEiiOKvL4khlj6C37Encv1rqS8bMmN8bSDFaEXggQ0wBnUCB/uDlRsGR7ga2mK0FCXFCZ
942qNxg/2O3cMyKwksZFhWkJcYBlldM9fNlXdEwzamR5zgBskvILPsuswF+ZfZCEW8E1C+YTc3HR
MGYN/omo2i61fTeDNQCGBB+qVC+vYxwTuH0vcmLndGzRYjR99poiQ5wmcs/eju07loFzJMYPojJM
sirAOKLU71HTcfxvZHqVgxUMf1/WkAdqee5CWWwLtwHQMc6KEADu/aY/18DEkW74OH4m5MNvkxNj
1fWPxIhdOKu6dJlSWIg2nmFuHECcw6W3847Q7gKO3GJWCZLg7s2odNohGOoKorfaucqSYkMnKp7d
9SWA18HS9xoh17hgxNJtoJVoj2k77E9l3U7+bS76gcwE51rGDwrVApD2U0sSKY6aToqpZQalFbuI
2D/CKcTJqJlMhgcf42zdgFWRkf2wP/1fzWQrsJ3Jwjc+YHpFqDYhY6969rjf8MHwRETOXpjZD+hc
LUyAsVmmUM9SgmB7GoJ0p/0ki7hRMiz5cVTvjgE+WimmRgvNpDiZM2VV+Qkls720ONMzUHgELYic
SoYMhNOvtmapAokLfCuVhWUg9c8FP1c+y/08sdjJdpajo1Btu9g5tkmX2ut/PXY59mVlKjEGPyf2
HRt45ycynJ6G7BEPg+vzqDK/606Lh6GUF15HOSqgE9fWpC+phI660x3wfW82l59PUZLwcUO4fcy1
EpNIj+hbISf8iESVGopIfWNngT5zsjXbog84SIzZRQMsocSWM+sTzNBMFVnF9AvuLpPGoh/PVDbF
NkmjxvBJJWl6LLEWY+cV0CjInh1wCSl8SSOSYNQUMBmN/xqv96E7IxuMrBOsrZg20n7sxJ38mq99
K/fRYKkDmFn+xYYDZrs41Y2P5osy6gnl+xh6vUgwiqKgxojGZXnWCyIgw4aJJ6FGR++VdVRXpuoV
1X0mH6lJ1xy1UiwUJThFj8r5WeshzJeT+k95N0ObnVbKDeVFKx7W9NpH2GHqEvR6SJgFBnRtKKnf
PcmW+H/mdYITd2P7PWTpLIKA5saxjMDyjKlkT8VizTv2mYjKVss61aUqGRapdy0Zc1aCsgudC6lF
B6I7CRS14SluGyUHnWFvL7sK5AEIKmr0fDK3OfGKnXzV2Vt5x8YlraHGmsfBdXth8HtIY2rarWlp
pDpJlOsDPnrxgZfgYtNEtnRRXIpvWbb/8yCEd/YimE4LK4S3zOKHR5WnXtepRAi/SrFypoP+FUVH
ixRwQKPflM38yESeGSKR6P4npnBfE5iLW5H7vogoKVDVEHp64NudKvnTGy/eH9/F4yDvyxA8WKAk
wh2WVKJUFFw/0NeFaj7kNE5eItl71KAoNNIAZqViZRn6kERkvHmMX8ZBa8UdRv4gzT9YICXhr/LR
oh2nTrEIUCCFula7YIzGFj/jzDJ6EbxH2Tsyrr1Hmj9S23e3EPu8FySzuvyfvAn5gsAFQT26RiDX
jOe3/qqDxiNDVN9genld3Rn4/6nqhA2GgVwUuk365KTHBSk8v8w3BpVIsz0RJHBUvLIAQ28JC01h
/1KoPpWsBhdanfo2xR4c6DRu8GgEgu333B6vAJ4m8Uq6ISNNTIh0i/z6k9Pbzk2tSdFSntGMeUcT
29TJF8VrAyw9VdLQEwLXTXsh4gNvwFXUzc8lsk0j5/iu3fihgjQYvLa6XEWOUNwdwSbMdBRBKWHJ
wX2iCyyea3OfPL+pwAv78zWjZmcEDvv2Ct5XQ4hemsIn/1KXJtHOy+uWMXSyyCrRc2kMOfrzxUmT
oWkOKneMgVVydyCvz+GV2AimHz+ac8h7fcM/Yi8WkKBlO5Uzi08ZbHtvh6joDrpa4s0QvPIOVdzv
533Sea4+JnR63JWs087niOlijpC8n2e3EeQhz7269ULoW2O+kI8yDzayRawd89KI+X7B0GcqEFGC
qhMYvTUzdGiwYDhtTYx2mpBsP2jEYIEMB2Cst+kJqirtT/0/5SGAqry1JqikI4eRWoMeHtphfy67
z7B/dl8LKwCDL8IvazK64keCkRNAMNWEE21gw7ZMne+Na2eCPO7Sbqp0ncqKIf8uLjH//5QVjokD
f2Lw4NPkr0lGGFAyMTH2qZ/eFFzGYwghZI+Zr9BHMLFbPqxvlEVBhbq4qZAPgLPf1wLIzx3QSj9j
5UuuPtjKqYLh+ny3rRmsO4rTCmtPb5a5N4Afrw7Otk22fsArktxxxodhawHkY0bkGT5Rq9TJ/Asm
YA14s5PNjRboHnDaYZkmd0LVPcMv1gLSGdgOwkodjFZXWC7WsSUGKZcVAIzioJUgB/WkS6r3zRST
7TP4V03nktbraisozwVx4Wvj7dQryvU9/aH1yTqU5EYT6sNS6MCSuxRCuArVv2Nub4bWuBl/Z2Kp
BcWvy2Q7+mG0baLPTLcYQAD8azeN22919tEZM6f7VsjkJqRApExHNRPz+GgMyI4ijs0Spi1L1q7N
phYqhuDPTYh0tSEJ7wEWSEsddyP/rggpQyAjMf02LGTvdHsVGWS2q5+aF++PHMl8FQvWJnyVuOM3
pbUqhdZqEe4hA/X06H0ew6LjorLTZ5/VNmuIprbxzTPDqRBMWT8ADgMJZVF4vl3o5mn2KHO2B1XF
/6AIv3eO+7XxXFl2hm5iEyOJqRmhVd0Nc5zYJ5tn56yXe1cGA2wjo4E7TIovmKr/f5oS9ZMz45kw
e4xPyvG4CnRul73iPGtWxVKTqpg2HoUsHV7uYQZtEZMHD0QRkS89pnenhriHfD+jOtkQqDkUyCld
sR+T4PiFQPxXapskIOxKeohZqWT0JXN4FXmWHMG6MbwVvynG+A5W4AS03yLJQlMsFabiV7eegWPr
1HTyui0ta6S6W5GKLyWF7VfeBzCxwC38vpiffhu1jYNs1b6TwbCbra3JceKQky7hLtoIk+tsFf6l
jrHA0RSB0J3fEknijDgP2erY53PfhbweWAUl1FoQ+SoGyLwRKh5HPEH+0jfD+Ibm09QPS6GsrmQM
L8U+g/n2VYdR4ajZM2xTfm2In00kZSq3wTiSHuBiM7Im01vLfAeyj4RNO7V1h+YVQxiLNMwkmFaz
4GORaheP10Q66k61K5fEeNkjF6eFUDzwYTxve2fFe5NGZX9CEeeo5mruU10710aDr964OYkGzq1K
kSjjhEKnUnYGNaIXOTrr1V4xCf2/YCRXuy5JkOkrR4ctYULzTnkNK1TYy8Oc1P1JNCdGLgZTXvHV
fTaU/wmfzeXb7marlh+90ecGsKCyzyFgQ2AU2/qdKrFMRPgo2JL5a0VTwBGzNJmjw2acrCepisAx
ks2NKMEy3Ed+Lx4LN1UcwvQTRkh/Mi+ZYFNCGaulGlExcuWYLY2Sl3ItKurd/0HRWD5q3CivZ9ig
Vz6XHORsUyGQBLKuCgZ5tugqxuvvYW3jmV+hDFwiJrgly6aJQ3ENWwocqsfm42itBDyErct/W24U
X+1zQu7pnwZna7rkCWE12VHuy6+XY8KDWjGt5jYb5yA/8B05J5QblhHHFLCBGjlK3uovj6fTOnPC
SCYTcE/P/2Zan2NXC32yvNvrt9QnJmq50Y+eHDhXf4phQ9O0gSn0fOR8VLjYIqtDYYcKWRktLbHI
A1miiCdIpOG4hoRSgwKhh6OCbFYX/GEC/tdwsoPMpRv8sSdgHKQ6tu4UB+PKwQb6RV5He735uuhg
M0rtiVkkZbp0fRpsv6TJOgsvbH07yXFHGwH3vuqy0BSgCXj99WyEWdheXZzm1FxhXUujOe8/mYAm
hSSaSF3mlCkM2xUINvqGUWikpDOb83bQWe3/2Uyoyzrq3+231A5TS5hGYRKizQ3xh37BLav10CYY
xhh3iunQnzx0WtDPu2Ai2D+lXtertqMqI8wPKWki916nw3lPkzDbaFCZPUK/fAbGlUeja2dFOk72
HdwM6eVLDWk0KQNvp6T3jOHTpj3zSePvZaGwjcZUm9tR/N1g/Hc/BDFv5k15IHG5WvJvpDuOCwoc
B2cUvZsyhFs0T7WupVKpRaEcUs/gS0GTs6cIzJdQVQ5+YIzO8RK17b3pWuLbk0r9XXJTOEC5IrLM
ZCTDhRcpvZKHZ5uUegJ9fCQ0T75zau1Bst9sWlomo8DXspFx2E6hZ01w/flKZw3gTMk+9MrKLyOK
Z8OTBgKkFKu0wm2f53ckDlaQacpv4K3y3+2dOq09knpYefnUumntYpTRvdgMbJRwaaIDOBuftSMA
62VvuumbV3URedoXCC0+ud7eLUC8T7KLOGngxeu05ZJIKWCWhMONU7PXkGtqeyTtGIHDm0vXtF7y
UjkD4eN2P4j6tkhVKu2jT3i3UBAj5Sf0YHWudXCs/WIlpmH2TLY+ELOO9Ak/1APPXK2Xtxy6miBE
K/DoN9jUQiJVjzQHOxYv5n71b9do0giKuTuY4f9LN3K23PfP75CvlWTkNYWU5i/5IStpHg0j7N+6
Vb3rYHEDavX20MoZkDCVgHCcA3dZih1qTs3tpG+cLpbH0rtMNuyacgQRFizW+viOnzAp5NaLadk2
AEDSPbrpIx3ZOsykTEfiCcdfzwtD86kXPXYjL2nXF9B9bctVhCU7O9g2516xC24Q/yknhbxTBe/F
5VJMwX5JL6DoL+LMde8BEh4p5qkOcw1uhgHCSotgcstzW3bU1o896Sc5Z/XFzsq7rrp+Jk69NN+O
usAOy9OddFXta8XLbba3Kr72R3gJh9IRvxqUQJB5Z67QjPgzPOzeC6Ypt9h00H0qmghmw0Rktvti
Ek3ZiDcro7Y3nUXoL3KLHZLWFle502p0uPGr0qkeXtHkftuTlvLYCpOiyvq4rP/aDovZTGyFpgVE
J/SjU3Y8o0bkjpMl0XSz8qlygplSwKruwKaYZduXSLHV75+sg0zLifrKuaeGZ9lytGFXzXfdHxSx
wmWOljj4XEWZdRDQVI9X/PhI3Em6pdIQqUGPfuNW8j32A+4cLi1UNtAkuVrk8jXEv3TYjMbfeHft
MM3bixTRJr/Ez4TpKeg2iuP3d7u+HdJND7mgGz1FxUKy2bZwjySevvP+KFTgASYh2s3BYqvyMP+3
gRDLT6KUAkNy0l5KEPwZzF01UPT/Yhr205w/MPawjFFUpykkKB9oAm2GvS26ab0ugjMoDZ9yqIET
Xn4KlPCYVtQzWqOVtxpwLNyrkL8da+ZdInmiV/hACWLhDAzVs9tWFfHDNnGJDAXjZyL18ZtOOIzc
/wiFzuON1P6T9/DE0rvfHWJiWS84RMwXDx8ZJVlzugFTB+QivNDbvv6ASKdqoZzfkEABcOl7Vf1g
Q2twrE08fE5EOhi0dd3NU2v0o5bCOCOUCL6hv7zJdFuJR/R1VCFF3Qk3ggGnDu3xXV7cIKX2SZ8m
C57bGU6VbN7VMuCIu1LQoJ+KXKuYmNfhRHVaywN8gybhy0ZdnOXySPsY8QlzX6NmYmFyQBN1Ovzd
pQXXtacyqMCRCBBePRTPYR+5uuOo1vN3Japl2ZQaQzFLgVa+GvzAoOGJM5I7B3iGk/P2uOXWNDlv
9gCnOoZTX93O7UCfNjtdSyKZSdxrAOzeHPOX7GzdJzCsbI4Kj4Dj1/NS0c2dexH58nKk2Te2PIYG
ZVDi+CTUCtGBmTvoWzF/nDO6BIymKRxVHknJ2o2HGQyfS64PDu4H5HRaagymtGuZCi7SmsFwSSc/
AmCqvzJkvppvRMpvg6MmDTbciBJsawq9i2Lj8fTG2XHP+Hebp3xF+lwE9tZP3a77TOGxGgrJyEHU
vYMwCGdOzhyow3s8pJbLw0G3WZimWG/Iy9os9IRqcQWdvYStXYahlEYtiDhZoeoMK0fiUMiZoZSc
J2julOgU92I9qcJOhqvfgEex1f1sHj+ZT3LU835DElMx134vgpmZaDeETYNFdHJ4aRubc7X/6caJ
WEeOvAVNst2DSaAtr3JhHH130hV8x+p7iPfThxzWphrzp9sYC2m4fo973y/aKZRIVwwMtA0M4lUw
Bm83sRvMxeMaiRDzUDlwgahIXVDEHUjHCbIr511RbXqv4G+HfK/qVMSBlNvRsTkHjBk5135l1ZLw
zRuDV5PB/Ema0BueYc11yCMk5/gq7FqB/AuYl38BfK5Dpcpnj+Yp9o/9DibQglep+lFV3TQbC1CP
rYxGGcqrHaayf7ejsCWqBRS5Ewh6JNLyWYGVN009S0h8oXfjp3KOwpykqMj/lGVUs5KYDgpBhBwh
fO1BXyHYMU5UR7qavBuahkHqe4gHkULfzN6T+rf7Pzl3O5JDnY/KAwy1a4CtduPBabs/FqecTVSF
TopmDR2KyBmbyRYr2FEs3qxxWu9rHnq/t3eCC9YjRvPoe7GJQ+fSy/0IxJxgiBvvdENFnbwPohio
7XStisILlQ5VcOS6BT+E+peasY0PT0b7UTX5wNXzGupDiRyu8q2bugnRsZu89pa9014xddDnG6fL
HtaOxaMrilEpLWJamOxfSHaUXA4VjDxLpjZ+jOasPr8+gxrPmne0VAxeUD88PuHgcGDPboPM2uLA
mYTcADBNsvdaQ9/2BE2wot9QtVvqZ+1lpL9aLrljliDktW7QFpY6QhZIe41IISy3FZ4ir+pmg5XY
nU3A8IbFlWPqyjPVtQdUEETZmm+C30S9YjHiTERbORE86s2tHNtRYBkyAx8IfK7TnEdtxkJJaJHH
eYcRUJDFD+kd394Mh2AbAgnEa445Mcsr1aCVcAUPjf5gGeUvybt9hUReiEAiF7MNisMSZ+zrvm09
moqBe+AYygndU1Mz2uNZ7hnOILbo9p5nWhru7BqNDO0biarod90uWvxF7tSuZSp4mWO0Ork8pmdK
123CFfhNcI1cHWtEGlxV/rSso2LDcPkEbJJW2t06TP+Mpnm9VADOhFRoFgDCfVqVKxFto1HBgsF7
10AL8ppPOs4iJ+TrDCIvIy7t7d8h+EGlk1Y9dqudO9LNg7vVv5+X0h/4a7W71gQu70metVkqhCkx
T0lKLf02+vS6eaZl/dMLeCmKt8rqUeVyuT9fPovmxfIwlN+9YokKHlJmACl7LrgFOopybGX7CmXX
PKs6pZIZOyV1tbAyCtMBJy1AGJrRRLy/NCEJKNJpAW5UP1LhCP9OWrjBvGlRmxxqf+gLtWSIpsFm
02CZ+ehFYZaxxG0Mr37JbVYowVt/Uk4RnPI3Yi+OR3+E03xVqtTAyfP+MHldYw9qoZku+trAyJeU
sP8ZF9Q3zed3eUixW0ArOxVnH2jzmmjLadynlrw6Wfum3JYIwBG72Atrv2QpSXPn86hh7LVOSgki
vR0ka4Jw87ub2b/GFHmLA6oquIMzNuHuqJj1qOoY2Vaz20ohBpqwlSrK3F4UD7Y8YQU0S5KVN+gZ
oWuFFW/I0b4erN5VHZkRP4HTCt2fJH1BNj8XRPDDfxCfa6U0YWli/nbKvcNwcJ1jzv28QVxVzOdI
6zE7D1jgbE8I7NYQnEGDzOjqDiEQVRIcqrT05Fe2BN/7Eb/T+UqRMzyvubqWzQ7dnrDuT8nR7+St
I99bgsNq4p764/3Dp+euG8e48TUg2TdXEhGsW6F1LF45xThGyDKT+vdfXziTu9eBmbfnYeIeQGL8
l2f+7Xx+XZPW3Os0PRzLekXMBKc1qDX9TjHpnARX014L+u/DHHrk0exVMynpHxADYp4EK5W6QT57
V5nI/gD6yHmVrdr5oKvjJ08eFnoQf/Q+8HnS7qp3J0TcASbtxueFGTZV0ZMQRJvTi/WXNsjqa4Ak
7lc6uNbt4mBjbsIw/SOIUZct27fhOEB2VnW0k30zhjKVjLZdiKg5myywNwzZXNFM6gfTg02Qch8Y
dtMejtHzU89336tmvnWZoTuxtDMGwr8lVD4Zz7h5IgA7V5zkWgklg0khb5tKLZAj7qvhcgBvcJDc
rZLnfCrvV6C0kUgmFNxktFHgAk6w8fplj3KlAPOLElBO5k2UgWViIUBwBn4DrWYetK8MmhP2HqeY
mecjzfERk3kxrjZ/Hnd9yq/PPdlkK6rIocTNWre/YZDaPxbvn9dM/vZW4W12Y6kx0+i18EHg9G9K
vo2HUl01oW0I5XIvYGulfWLWevjHabYthzm21tNUpJMN9B9X48RBldiKtbJKOVi/Z9wzESOTNqE0
LdDDFN7Hi+d3bsPCK18xx8IQn8tEybNG49XaSjd1alWgVvqGfncoCAzQhZKbvuXAJG7BD9N8jejH
4dpoMsXM9xryg3tQLztTeZE5cfX+x08pJVg84xVcHQzJZjcDWDLpkbnxRXnOjGNDXAd42sCM1RUh
LerALZ+QF7kMRdpZMYYfKDUo2SZqQcpHqrICum6YL2J9KkLi4iIYUXpHUdkfrO6KV1splV4AgryA
kmE1x3RRsEZyJw33aKK0KorlTUxU8bR9cSdtFQiXWHMVf0sS564lWWeuUXKVg6tyMd5nHclWTmx5
Qi/HTB17oIN8bap2GkWD+C2fAQTViHZWeekcHXnsVQKDRqiX0t330MyK62jTyG86oIqYyrBxLSoS
qiFLEvCt7zqaygXelCF4BGl4qUzRSdDOK38hXKnpPT8NgyIIk5bDQHhIjPJFfFFcsbYnVky6Ej70
M2bRrpd9GNo2cQ1m4qlJTqtnbrs8i9Koccb2q7ZAq0uX4jRLgXhaJGOg1NlaFnxxjMdkcFVEAkR3
QTIbJQ/SrkXAQ+1SaPOlLZV4GldkIATiAk6i5YHGbrfXZTSP47Fmm8g4o+YQStCXLEZMYNneWT8d
oSM87L1qOPpx2lQIj5cP561iaxJqlh28me7F7blKnH1j46AydBOiAHg8mmshr9NHIfY8eNbWu/um
iN2395AP8NKgkekLvaHKn7JNfoI0y6/4bNfjQ21IIOaKxcxZOHLn3+8uR3iahLN6IyNU//9CVGXe
jnnhSgPXFfFzcbutbdg5VSKpuEaOHtAE3KTnfK/Lg0UsXxLnc3JppbhE2ccP0oOEfP42VgwRk85k
zUP1tigxN73Psk7hcm8Yis3ojKwR+RZ2piY8wet+Mlc5TQ31xD4DasLXNT+WLskfddiEpwegjSk8
qUwPYDdbwSXOLhSIGSVmvStwiWHVKckwRQ0ztuKhyY0jPbcWoiaahEPBk2JtHVLy6g2pZNZutje0
ykL9DH3stTlNOlGm52W5mxnY6onXLk+zNirmLI77a/dl85DarCQ76WphU+qfPJxdT90tVkmzsE5t
NcPdOH2+yCb9azjJMf39TATh3qMi4gTn1DI7y5Ulu7dXqMiZXKq8EJwlGYoP9Od9dhT7LvTy1G6P
bXHgNj4tZkbZcYupRH+oMg9L3N067XqVy7zNlRSl4lwWEZEgQ32OHQDvGUy+kfClOjpRme7X3DOt
HMPweRA3PXVs0kouZg0XHb2DSwkj9jF1xd+YnskHhLfIpW6IpOBjJ505+2KqzpiIwRiKVA1eNADQ
Hz/9PKFtb1X+fxgmIkAjFVwBucOsBnCCwhG2/9TxYNFUQkH0+FOuywXjbORydU1n7F+DDybGM3ER
DeEuqSshfyaf9otIfSGGcFkxlp7RHSTAaJdDR7rfMcJbmC2Vf+h+Dz/z7FEKqbiRMLFZHcr/IrT0
Zt+eJ9/r/eQDfR4zprCnVPBaA7IjQUuyra5ovRPSgBzHMGImbOlahkwC+C78LLQPu8WOb7LAmXZv
9gzgYewhyKdsBjEDl416lTgUT7matgzkubT95aiJKnRDfWdXS1R5QN3gh34Uw1KdRvd0Ro4Z9BoQ
GDxkwKkuoTCT9+b1vFk2DvoTitrKEqGLsEs412isL9P/2/mMr1oYsViphREB87XtePvm7sMX6GCt
gF1FVGdos3HvkGgnmemV7Q/3yUiD8vRxW6fB8P33BCyTbi7gxbwDFPPDwtSEGGyamtqu4JXKsJiE
EgGsjJY7zYY21/96QytAdaTXBLaCZFqv6QFs11TrSlf/H5jwS3r/aZYp6qy+Q4rMjT7Ekg/AErZE
akbDdQB9dJK5I2ZqmqdnzN7Gzh4da9x5AsDZj2hbGn6qsCjT/pr/Y5GxGxGYKJPUY5TDRARiPVQN
KPqgNq+PwrhHPntXjdbfd5eZDdnjeE0zSTKkxpvQOXOO7pzHm0uHLKSwfOu8qAo4dyq+UVUtal1j
OEpnPCJBuk3YzkzuYA900dqdS2xpmMVHnr1kX+Io48GQOtqUHy5n9sop8Z8QfaSmD9QXE14fTHGo
SR3e5scXDLxfhJAFp2N2Qp6VoUzX+2kNLXeQIEWsegNbYT9iT3jqdtPdbQfYEJ4QnJd82V4FxDYN
oM9CqwvZfypkRN7zhu4TxCU27yvCk9SsIEDzilmpkUbs2Can0tW0S7y+k8bSp8kII2g74P8xlYQS
plFT+jhK64lbqF3ijThQ1ie4Q7MHyb60HZ5EuFAw2OHHGaZQd5Pa5aXkLMQ0fulZBkgPzsBLrYBc
NBky0VV8KkBDFSBiQjMoEeW4pvjK6GUzytYrrkdzRFZDAS5Cx8YwtJpStkUg4VIlxWGPwy1leq75
kq/BeI823ieuaEjFPCvcN5cf/15CEuz44g/mXZY4ffLNJjqLhan5bQPESyEzzE9TIM+Dke3lFcgn
hTjDxiyabBcfwascDGrdtt2WsT1J82pqpA2ytyfMHQGK5+pWR9cfvyJkoD3Q99UaK8NS8pN/zuIT
CK7tLXY2ZPxTbIudRWuA7aimZbnFmJUYAttuhICA3eYzfyY4PrveA+Uildm9K+JaBXt25fknmsbw
1m0keTABVGQCn2eBsuAytS9RFORxY4eXX3cgRKRBnqiB2sM7y8w0SDSoqFs8XofqqSgFxfgrg8lL
n+zW1y81IkcNjhMAse10kVM0RDNX8kSYMDseGLq6gz3PvjdEZu5yYbE7gLmsW03IHhnkub27aW3+
T5pFrW76om0rluLyfK2kw5hXPwZ/1Zd6q+orGntsCTDLqE7+okbkz+rAYauDM+jwOHBEVMQSX7Xx
ThjJE8EeS6Ta/GutsZW8m54UgkC/F7FDuMCapP1p4TG7C5Brqo5KnKt/rQPrV8kP6NwPEoDzgpmE
qU6gASu4aLPgZkGz6mZPgEW4EDsZ2OT9q4gGru8a8RRMGeU84B//U/86FWYoJv2+QZA2uOuNDSMH
UVzOB4MFLz47VmS9Imc7UYDsI6JgloASvZcKqrJjopxfidU3EN0kwkgXtoOE7HXrgEo9Ocokrha4
+0qay2TUgQ8Rd/eBGURsKoHoaxa/mUA8uHvY0VxlL16J5HuTxM1k5LvTGjVctkSDWYPXyquucd8W
Y+8Cl9vmsyxWCyAtQ5KA14g99whJBpdNSCUzFmeNTOX8hgO0Ztz+PVNmp19er9O1PFCBe3S4pNWL
Seccvp2rVjsCU+IRMqh2MHPHnowA30qmfwrVq9Ro4uZEICCDiQ4Xooq9okRpiULdoXQHbh2lGHCa
VwUoHYxFlW7Xj3W7UyV7pLPbOu5Jvi/4Z/rQaq8SCE6K5vHNqfqUBCST9yQHiqdC/vFU46+m/fAZ
nZ8pJz93kML1HVN6h9iqZva6RSLCBlXQQw3ngcWped2gBwIT+KF7gt3kuHQwz9c89xArCAUbNPcU
iRlq2O0KEgxHD/M+ue+n/qOpbOxtiY9XLDiqvBDIq1PSw+o37nq9Miu92V7foKPZkBsKYa3/gSPC
DWdMP5aE2kGQmYgrcw+dqfRw/qzcBdEOviKzNxiSCKJHtnq8khI2PPeOpuEhaVShpwSunSXOdHMv
LMjGtTq77A92tP26folySqgd3NwWlT76mCYwTYGiYJCwkceFhdREFMaG3n+DF+uaHO1My20Dt6iT
FWlDLD5t0bO7A+H+9ds6ps0LwhCldrbJvrqkPtefOS2za+QGcFGb1EZnxppAaauVkOg9GsFuJcrc
zhkYv69wihcLcxcMfdlvtBqqdLa6LVwipKsiu9d171BuFxMTyeef58M6i7umEt4z21TSe3m6gdQl
CXAucUfjYp2V71oeZ0Pw4casn8/XX7IHQKZ8eMsC/XG8T9BJS08soCjwjIJLcyeLaktCI28dwKL2
etAZnYpta0BLqDtPla0HDLblCGOsl9P5+6UJTgAHMSijtwe1j/d4VbgPk4xnWBawNAaOIs9uL4OP
jtUb7Zr74g0ENZg1v+wwOZAIeBVrk195prXOJFafr1bu22qoZI3VKFBfvsrQMfNpcK3Gunq3lD7r
NOll77MrVzOJusCtwzKPHHL5PbzEB1Zk8JE5AySlqYQkgtpAgWUNQ+TBZdHiBN7eElR0+UxVVIk/
mZ26lwllMO4urVBaCHWI6ha5wusycxZXle5y+SfA7WUAN3MswQTSQcWRq4H2Qvs0QAitxvElR9VU
zCvEAXRuV8kvPasYeEVOD1giWaF4Ug38WFqCEdzoWQ0Yv5jG+GteY6hZer8IcwtQxwvucnef/AAg
Zev3pDpc5wumi1UFmu3TqIUhACxzfUa+1IwnBnzWdzby81L8Xkla/0sj5X+HPiuOCoDGXPtIb1UE
za7VeG02q/1JA1lQBkLumsUs8JxHkIfU5jdj5rg+IQ2RG4uW52wfhrGdDOC71CK86Oyn0PSUgZPD
jtYeHFQ3hvPUjQFSnb+O8AH88c+4n3fpvjFamaUk3aRi70Aw6XIOC0kgu0WLnY28/BRog/Ac3YuI
b8UTLhjFkq58wBm6Sf2c9BaWe6XOwwhqhEZgN3XhxMHRVfC4D8mYkL/P4T4VTgbqd2VIG8vSJqFb
eMZNl0WcaLLSNHNBNESU4z5gZVM0TcVb44icy3+6FQlOYfymFBkElCRWUT+5JjOEucG62HZrNP8t
wGxm9k6Dx0m+44z3K9HKtVjsqFt7YyHFxl74XJ2go2M7sjlbNe5Td8HCRt+KFMu7pYf1c9WlD+bY
a1p1GWZ1Vxpf0oWn8aKbIxbPnULv3JyMXnhalq0GNdD6CM/4v9XAi2r1NxLOL1Jm//lWx+6QDfbA
hDxbCUIYTnQJJr3+QuuSDz9NuOgLWxlNH/SJl9AKwX2DP2FvB6Xx1wXL54IyQiwNaIh3OpQhQ3Ui
oaWgrlZy3Lrw6aQgkua5QVtCKQ51JvodbVIASrWhQ8kngxP0kYu55BgGCLnhFautduzdW5/kE+7c
SgJwa7yAmhwwHC/1WHlMZQR6kU4hhuiwRbSewE6nUPBWTkezq82SXQyJucDEMlDgxLQukErO6BSE
3Q1xc0O/YvnNzg+o6c1zFJp4lRvN8nyBSKbsIQYcBmh8jpk9Q65eTTh3CyRNUdwxRK27bSyGrpP2
0YnVsy8LgrKKMb5GV9B/QgtjE0vupd/1JJxl7kkQe9f2doUxWhcHDtwD5Kfo3ZAHDtphsdQ7NEVT
7+DNbg9sKiak9KBiF86rKyn5igLt9SL5exCD/1iu5qbmtJRv22dIk7FCctOcis90cvFkFoCbn9d1
rq+8yD0er7jjY8/oTDznxhZ7whAU/EMvA0sC6w+SbFYFEb7TQ/l6kmIZ0G1jRlzPpZ+oUhd9flx4
JT4A/NjB+Zm6uOBeSh4MY9rFInEwkGJFWM+uyRV9MJMIpKbM6YIJZiy8g+Y+BjJI+ICGmOfTMKT3
OyAqa8ORxij9aUAjPaMiNUL032gwD6NvBk5/RpNkVVISQoZW6ng9d8zW0Ht97/N671O+/H/2es5U
7OLqcfBDLapUWSRf30PXsgtBCl1H4ZVeIxFbWiDoC2fILrlUgpkv5NgvdmPSx2E1MjMVLOqivDO5
hkFYfRj8Q61IOhB9UtmsHr5ChdA2twe2mu2jSalFZ2juLfe8USESxF64Z8nnIm5F5CkPKAVuLVqt
w7NsCavJum1pZz3QC1XqjiARnuAjZygs9jiD+SRPOflhCJY0iaFEyP4vFSuuZOM+Y2G9FxchWox1
VUe4zJtIVBWz7QUe7W4HfYPlADM7aXgP2aXpk23h774mvZAUno1gGusR5JNNPDLWiueqRWeKf/3W
Cc5NPbwKxHdRbr1L4Jl4s+YypD0NtCdulNDf4grPXeUcyMI74UillZ06Tv66YIKwyIgeo5YbUdjJ
E0QuZYrMaBLx4GWfZ0FX3xEtUtLqRcjeSeQjiB2F5L1kP8hTJNxadYZv+zxGE1c/DkU1qwjsH+S3
ETuvQb8+GM5+Oyajup1y4IqvWn1uLTKh2Lv/twvGidfhtk0SvVytqRhw3dVTyiJUvKbbSM6e4qCl
t8kDOhg+xpuh423/+vt1+gsADFWbF0im2XMPWNvJ8SYq0Kh8XWcukOsu+6YpHB4WOFCr47ntlB4V
WQgeVDXYlsChOstuJFNRMUaZlyCbB04rt+SJuFRjnL56jmULo/Zl+JHRd75sD0I3Ba3q58gky7IF
JICedh+O2gUR6JeEP7NSZVWD8aZQyyovxreiDlVBnIir3U31poZljQS+ZBmVD9LAN31Mm8hYQuOi
mzVbHGIMRIzval38a7J5On8tG7oMakGnfMESLosTY9RPt1UQJyCDy/rqAQG0dn6TvF9nbpz7jb6t
+/VJZwOBMjdXwEIuWl0/ILAdNDNp9oDFE327QO965RzdEvM6OwvmsADfqku5gFm+AhNco+DXEklg
hv96fxQpHxh9kgu9NybhLFwOCwHfq562vpjf1zNWsuUbxxgR1AO9NHT5/H0hqXldtQHezH6CF4UK
kjRbGBmQ4QHfhpTrB/ZHW2KcG/lDYmB2OMoqSUa5XKECWgb2WFhYC6hVyVSCMv7SIK2pa9hu8Jm6
PxSTCYNx/kccQWFY4HBBgtoSwYdoKu8PaY3zhTBGQ6+viMAQ7+xsMECN5zpzivFOP8HklFSlyWOt
a6AZaVgWg7gOxP5RLL3ECYi1jtpYNW1Y3NjT1ApKfKZIHlBep+8yZarnl8zJVBiIOKO8u54F6Y1t
DGEXlegviLkrFWzLVkFH7P+sO+GZxhkPaKKKliksP06HxaeHjDz/DTwmvaQClIYN6ALpdjNJwL0Q
oO195s/0+jwtzR4+aZt5jNfrmkpTm/BxckMG5bDfL4JdHGlPjJFgPcwfQo3Liu8B4KijrkfNH84B
hpJfidMoNmENjvM4iwO4ehfX/pSUgRNTihtgfXnwt0GZmVab73jkzmCTrKq3jZmrlevx0e403QMG
dPnqvXe7gO4EGgmaZWDsNRR/VvyeVVsCQMNnkpF6AH6RLtvGZP7A5DUmD6sJBgJO7pvbkg01dJcv
vxLUno0WwkQD2J8+yevy6yD4oQ2PktuQYAgquBDt/Y3JYi+zD4pG6DmNlYCt5eo9+ULLk4sRBh+U
Q5WitSdKP/LBycQJ2CBla5Zz3RwRQmnqmMk2lbhPfjfTHwzEMMVf0D28jsyxgj+vHnZe/Sb0otaD
YogRGW84m61tyYgngroCZz9XIQjJlk7CnsNJExnb8CsQ/HJpBUNhwvPggZmRTWmId34fFSuZFziC
VVZP/wCQYcsKsSADv/khd88lgJqsQGhUw44SlVVE356DVqO0EnF7FfNPq8TJra/V+FyS0uLspJNL
cuwBMp6mqSnySUfbYsDa7Gs8dK0ySWHzaom0CehE/m9VlDKuQbRha2R6WszlrHpzYhZsGzKBiynO
+ISmBHSl2LqxJxr1+Xj57x0Ama7je58KT27oDpSRgXxRQETw0WOJ+/WejCLxc6rRTQGbwiNGCmdA
Vdl9fLC2DZRMukFAzCZjbGnDpvvatFVijOIUq/FX8YHvbReA9TFL7hWgfWR7qWMT4J9u/ayX4gvW
q94UptsjPPm+RmMJhAuGXdbX7ZQ4T3QFKencH2iWAZO2uk3anFsY+knWACEhxtd0uFK//or8SoYc
1UUjvyLEdfUxZz2e0wf2bi4apz9ir7P3tm9hHAQnkYGNIsoLpFD9uelU4Z/5pEI+MCwNkJ1o8zYA
tzTMQSx/PgFMuzVLOkGeilsCpeF9ixuJTphJIquEMIbrrg6DI67nYy4sLmTOHRGR733rhVtch/NK
s/RmFh7sDINVW0A3SCzs/olSyjvmcCTa2Hwui88hZ66pV4z1lhopURYfW+fr7Rl5GM5U7xaaOUUH
gX4g1cJ6O334bsH+7ACEEJ6OQH9Tey1n4l7DkuaH9UvfqG/dB9QShFxitSVnCHDDtwoITBDsoUzY
E6fsy0b9p242YysQBIYq8RNJcsIrU3rDqmv0EW24C0ahOznPPleI8qEb6h3hzD0ZW7LiNAtrHEsE
ZARLkwSy2HJP1pFMnDRXVNDenkh3ztcTvGHAp+a8unjU6DfYF3z5vLwZGe9cHte81AfSkWKpUYpw
wC5jx0xYFbeHV9WF7ho2qKcIGjuCwOUQO+jyps9dxoW+mGkiF3mQ1hFiWQjzXpgS9mASGg10T7YF
dO+8EcNJh6HcXZ5dITy8BFXkUb+eO1vU0HxBAPr6pLqudfNEDDeUJKQnvNzEQG7sDANpsy+sQ67B
YrGYdX+f2mgCetfqdeMcP96DqUQ17QPBl32gRdWL4whzZanGwYlib1DGvjwmHpkUmTuUZACn9NnX
+981dewqKk3cEE/M81g3SYdudpoPO4uX8BYGaDFHf9Pe0GHv8UF/AI+ZQFs9u0A9vHHDS9pUq9Ew
geMmzvTplNtsoZXgTyK3cjbU2lPysvgLD5AfTliTIyiq9M1eDKKMlynqDocIZn2L7JnHe3kNOQYz
nYEHovGelJ8ofRvW4TfSPfWMJdLYiIhiC9mdtJmkyVcWS4xch5Hz2yHneUjCVL8d59ltA2bsLfkZ
dRa41V7QXSJKKFiMJ8pmoLxGsbJT+nNpeh3s90qT7egxJoL0mf900hI9aozZOu4oGnDmFoQgdLA0
XobyZOorf99Al9XYYUAUAHv5yTtNHpTUVEysf5hmwWvZ7iLw4lBgtJK7AYd7kXqy6o4swaBtQ382
sgZuPykxrESQNQkQblAW+BdkK8CzRtZfvhycGYmf/N6KAEqY2ic+9JN6/vkeFNE24+yBekjAabEW
4/7jdicULDMKgMRMVCFhODDiFc+4kzszHTp6cVc6NTmpA2e6KRgyQABWrauq1QGgAsqBMtrfm2e/
P3+j+XTcJOjIVtpxlMtMBu6R+9eh3GTRQrcGMzQkNZh7mg07fHWneV3LfLULe17B+Rjt3sGQm0kE
70fuIMMKNWx3ULy6bV72wXmMplNyEinCIx8EthTRRC9RRImiIVbICj6guKRFkwNjtR3CAaiYI3Jx
T8Z1MINnaFs1+oz02FSw36fzNOYbMQC66xmXsUC5NRAfruD0dsbZRmsbih9Tmu5xrvthDIsjSE6n
6KdHlOyIRm/UK2lZtwr0uT8Id/vI9iXtdFsxrcQxI4qzcpjYT4Kp4cxVmlsupuamooqgXWCA7A+V
6ANrzVke5mWzzng6C0i9Ddj7qDL8e2hRN3YY95W+qgYzGodMfC/SiYBpU3xRCR3xdC7ICKVUyrf8
24hEWH1+nD3P0a8HALKR6Bjr+7N2D5yoPvHg8XTmKUar+O+uclBmqWFMAnUHZnLMz7W1EXVmx2HB
Rcb6w6kF12863pUYYHB2obSKgr6dCWIIEvRb6itwvCC/rF6cYfU8FEtk+nziBeHu1Lqkij5bg7xo
OpFVsR4vZTO4+C955CUsM7KSW4XVifAU+I1GnsQm7q8ir8IRXPacztIn2FMiYOCeO4mVvdRqjrmg
SqJb3ygnHUMeM80xrvT1SXQ36jZouicn6w62/8+iPraAcOAtyVJQE2SRw48Y6L167sjNfUjLXt2J
rv4jQifc9zxqSMbn8p15pCwqgQxf+tdls10H0XmR2F7lZiO10/nfTE2UBn7wLqAIhDrpA0rlN4LA
Q1axBnf1acWk/6FXq9eOXOJ/p/EGHC2woUjm5rSCrd2Rqq8bbIZ0KN5Zvc2gbn0POcfLZc8R25nt
ya4m1sqIVAd8duSEo7RGNu+A3ZMfZqz/ZTzq/E8RYRSkAnBIxMF4TZkx2+pvrZ6cygQ1VcMtiwrT
1RGZsDQq9i5DhoMkYvfZZEAIBeCMLREsFJcowh7cdlfAbvi2AXzyJpnCAIYz+lCb+sFeJH6bNCCP
W3vPiIT6CbSJLH+JIfFjJMdjZoPkNNEDtj0q4wzlE0WjsUDf7NQwY5CA+X6+7H7Qyt7dHNEmDh7R
BpoF/wN+KVRFMeUTbUFqxXIfQ7K5HwC5abloXf5xlaz1+Jvf8Zr7avyyapffx+AfLIl2kvXGZpQp
JUoeKrvLKrHs6VT9yFvIEY77luBFaJzGrI22YRU2AvpJ0NtPsVHWY33N5HTRZUopVAkc0bp1T9Wo
qhyfjPfoOg/JUnd/qerNOgY//xW2TaFuG1Wt7S4ifh414gNP4wZZlvP9m/Ca2WBcKTkj79s8WtCo
fM2o28o4eDSkjEtzTz22iAFC4TScQkhMHbxpXZt3e1qCJjwn1Ku2FYqFojS6jyZBMBHDbnC1VQ6G
N1wvUK99j9R04UJc/OaqbKezhVkQV6kIYr+n8k1F0cz56knBADYRAPorE0mSo/7ce/oZ4zgRelo5
hZdv3+FqdDAITtR5t9mZ6rpYSKWLaRHYthLoA7rn5qTt1R5Op5E4gsacOKSiLNY+G7glW4bvxA5/
sf/sMDvqxmbkhI5TVV38NoK6BHwovCCa0V98GDg4KNCNflEPkSCCi35Z/+kzsMoqEEZPq/zaVbP9
89cgwk3LtKdhEUa5X8rUT7mKBRHlb8e7kXJx9ql6S6yuZy+BUVfYrAKdC1+4hjWtip2s5EJLb3Ij
7xZ4Zd93tXctcoTpPEjrI8ey7kIvjIHFZeejfZA5+KvJO+O8f3f4sAm6Ckd2wtdTCU6h8ZkEuA5d
ZTvLNHSNs6Wsa1VFAgbs9lhOmG0k15HRwN4JClVrMJQ8ULitOs0mUuhlM3ddj6piEVONhjS4nyyH
2FsjbY+UreKlzIXHWP2rXFVteZ40XW32b7K5D/vdN8JlbvGxYi8Z1c7Qnit7jkYSeN7OFBTK2N+J
UxlvksF75i6SSGcw7cAtbKR1DLaq522oagdM6WVcsk7QA4IX7cx2QEWwU3d/+2KSCTsZTNU8pSdu
hNucVMXG/PACbuyRRuswif0qqS6/h60XfTSp00IGiuQKcjRfl77HpZNyohKppOQT+ifKkfCROjVt
tFCYDHLnDp+PBLUBFLg2obRjMuBcuZrTAz36hlx48WTHojfh4jARdCfIG8D19iob+0bsSfz0Wdzg
vgVgzF+XlBF1Wc5vXeLskfzDFwNUCeZC2cwQjCZK7UqrHjH0WUebtXvI+cbs+LSIJO8f5Edyx8D+
EqORe1OzQY/EzuG89gs4yRYvQm6mMFOkLajMqwengH6FHIDFZ7FF8+1m9p2rbfcCiHYWplUqeNQb
1B+PeheOTrC/NzFEoWOeb/RF5WcJ74KyeLzmZu4h52pFAb0kTklLe9JGZSLAT1QkOFGFVD47gYse
N8ZD9xWRi0zeZyLxbz9RwlT9KhLHFyJG/Qx4QtTPsfMzUA90kQq0ShqZyx2NWm9ZQ4s/qYxC/UT7
n98wTbFsu8o5jyPcJ9PGAnuL4D1LUZbFheVaX1A/p13iwpdXMNMUtzZXTxBMxkTrSvNmaTl4rdL/
MQICDCpGpZsojpZRKP8zaF6yItJX6wApJjmHBTIAShYjETO2h431g1UYCq2zN2gpb4Wov2mgtGpa
qausuCq/zQvtLzkSln5L2LO7pL53tsb6PtbGkwV5IB8TTw5Fvv0b2XS44MMBjE69bbK213/a09nE
10wIFE0gatKdWVvxwuK85LKX1++Gg1oBeeYI3v5xuxNqcalXHoDxn9E5TaBEOKxHjVZXwDHi85ek
Kh8ANnjIoHXaSQKApeX/8U+DPNmgc5p/vWDxa4LFdOQ1VWonyszlcnoX4HuWG3zivEKizfRyNt9a
vB1hdD5QLIn0kfxwTMimBuiHEXQPYgnkhKqcdcldM9BIwKS89y1vPRMiz6CXuCAlNYyl5nnFqnue
ABQNVjsNojrF0WXdSEFtZ7fEXas9vfxKIJauRsPPUAqqR0psxmWpar2pR2+o1Lc8KghrFYU6qOUl
mhKtHnpxMtHxf+Pvgb9shRdlxoV/fuKLW6X3HYsGF9TFj1uDp3ODViEQ5TRP5bnlMxkQxLMsKJxB
nMvHr1lu9KtBlZ1IlKYEpGTohGop88TxTwqMlkhLpgA1/zX9hc0/g0DAGDyi0qsdsQoDcKuo8QBL
6VMA70xecjWwqzoc6V2JfQxj3JVf0zhgGtp4htc54dnQ7gSKGnRHbwL+0ZkFvU++M5Mw7ukcWKP0
4AOWfabuBU0u/DMWZKDwzEDYGL8CeZ/OAbjiC/KP4IMZ5nLspGnCQBPkn/v6neViTlVu6QJ4kmRt
3ZDSiaDtd0b8Ah2oOudENhNLhA+djIXrUfFjyN+XbGyx7W7PE2Y3nQ8GYcxmimqdvmht/7e4cdII
qYw77tiX6qJlyrLsMU43LuIuB6Ld99FmE6YbFUdAePr+oV+gNCQ8HRhZxTBmlGYdrvua731EnrA2
OaRTjIekEkzo3naCrfSSIsiOwOQT4ilCEqfGzvjIYxlA29TclVCFopvfK5yqGYrxwILuKQk0qUbK
iH+42IGpX+/+mJzZYjzf2v3etwFw83ZRigIlQmkQyYPuDlBGY60loC1Qo7IRNdt3XvR8Mq0vSaLD
27xCX/yCKO1113/NE2CAdTW9mTpnJxMoOaMMJ66CPML4nlSu1fiu5CXZbSalpQxtjM9SOg7zvSvj
GTQtHSnYCikTsYMCmqCw/jslCcy6AjvZtmpl9ThaYhich1RViB8JhcxuNAnXqXGI9RpDa0fR5L7F
EZ48P18NkBDJlObjUiau0oh7bfiMjdKUNotvnQF53+kW6De+94RTNH8zvpoTX0r12cCy/Vt/wMxW
6yWFGi+rQqC5fdm37QozbosSJkh754/QdEZzXOM2kujeMAhYygTRdPqW9u93AcrtstJhfjwc8Neg
jJbHxeZoRodNve1CxsVlEd9ymy0+HELzzZ95Gkn2Pmy6grMrSRKe7pFSAyW6NQM2h45B12DrD+YT
MSoJIdo0qynCHGr3s0QOu7IHCB5Svw6A4IdQcA6QcRqR13X5SKoJVuPUNUFl33TamMgQ1fvhN0ja
kOAfuKJEw52tGOyu8HYEd8t2uPCt95BGX2dfRGngscaHJFPCfebqFG5/e8Ix+jU/N538cw9jVaM7
7MwlGwt1hKvnXXn0PBZAtMuIe6IXgXSK/27v9dUxbEpjpJly51gfHc8rCWuzeBTrQ4qiElol0+W4
MWvOUbQw7tUcPxOkCoWc8H7wO02jzEeLjf2ej7J2d7gP2toacFyVP66u5HpIEqbCGtqwvnIdbikP
OQ60ZrUhnmp35TFe1BLKrBX3tO8UqdUTvw8GIPj40S09y6IcSTmxutI6PXK9b3G4gNZ7AugyyZLW
mC2L4JllFQWqr17YPlQZQnLCco+pnqxhA/5XjtKewmnYlHzdTbeQ8Xi0Uk7uJ2c2jU1ufrPCVPvA
R7UtN93QbvTcIk8jjs9GC8LjsXwCKvcHQRwmQ+aVatU4LsH2vEjbIwhpHxD3L+Tfssg70vBvevY3
W8d/vzyN5IEZKy4bqO+7vw+qTgeecepHmTu0Emq9r6Jlg5+DQodolAH7usZv2bKNEhsq2eVi3YjZ
Kb+BPYOXPvC+625sho1wtH16Qa6Yz+TjhyLLqP1lh/UOCOIMAFTgOJ4eQkloWK9I25Yrhg5aSjLa
LNjhbVIigAUaIbLTVXe9GWhgoYvMfAGpLj1avP66x26lmTziF/ggBWa24kSElcURHl11z5Yu9SXk
nqiwzWW92bNfq14XHiu8RgiQ5s/ol9sinHdm97hCsrh5HjY5ShGWLGUsofpsLFXRDhteEn8SYfX7
RwRGs80nySnSxY/ijUOoPmPVTLQeZVukSussD7eaRzcv29wkqgzHPoTzvXTqbNivxFswaXLRSZYf
pjmLTddyDm72LF659Lk2JzlI/4wEJsb+BCbzjn8Pu/QOEyCsZnpJyh2F++c3rFNaDqrM7K50aYK2
f8y7XynSE9Rf0Q4kpI/EJBSiTO6Ku+wBMrU4/2eElhhiYdni56nGKwlk8O5N69UoD5Qvi/k2IpWf
jI7h/4A2wk/7DnXOrzigxSl+UUoTSehst3J8bMvZgou1qe3XyT5807hlCPLCHea7RzX/mGek9cZ9
0gBSqj8BalMyXoIuIu85cUgpj8RC1mDycu3YM/fXu9jrYpdTzPanSILJCH1HKYsQxqJanOJAXosV
engsOkOLHvyeYeckRp3/JPJ1uy3c2sIKl5+FYadwA5UVUhXw6whus5JRyVnw0i8asDL/gdz4pZKx
W9ZgbNvCLmYzI1B8FOox5sqPxH6QRpkWlGnBPKe+O5dmq6wPyl1Q1St1kpMkVCV8yQjxKcdbVaqi
GcqOoUsMeM9xpCHMphkXCtFrVgbCOfyIKQfFVu/vD3vExRJPk4fnD1shpU48bAkFpiKi7aoiZ6Zt
Pnte90DudtyovBe2gxdMDa0gQgFIQ/A+2P/2o/n0xEVSDKdOCFHntdsT6u3hJpOqFH/RKYMGJSJB
Y0eZzJqNe8oy0xnUk1mHjhN8688mU1PcuNjzKBt/01tGOtJbiMST7IbcIlVi5/lOGsPnaOxC3kep
0CRrKM59TWh21h6JPf0JI7bxjEVk+k3frq0cCp4/f22c36CWBKxX8yxBTxwq0GYY8Te3YWqwyuSJ
T2NRjG3540CfQ7UDBpTa6LHCAMhTLeO4qHEuZPwkB+yEqRp9E0T+/6bgT7SvPszCM/8ct0lZiI6U
kQdOS/P60ev7JOyBddCbEmegZx0NcefyLondRRPP7EBevia5vwp8reQA8R7wQ878CGn+8PpcloTk
lxexBdUKacgiuahoyK+gKpfX2rmsloQhbz+9imGa7AesaG/6Acpe1dFzBeNgSJ85X/k3106prOYt
aQE0GBOkVbXmCSNR6DpVVzU5wqhz15kCvJIzAJykW0TMFDsWVdcyU8xHwb5JAOhtAflzX6AsaDY3
sPBKNRXtRQCHtmscRqngG0lAZW4qfROJNckBNM/CwAzt48GqO/bshFWrZIQOsteV4a0iAfqmJhhH
XvW4kVCakto/RNqkP+Td1YVf2fMkFLDsmW1qCP6s/ztqeke+lb3RH3gUYVn0hxgU/lk72dg0UX19
gcieWrdHb84twmlwtEYb/mhg09hRZ8KozzXZuuC5y4mojygI2wPyytI7xbZ5jLsyH/0Nhe0jJFGD
h2w/NkQVUF2icIWy2a7ZHrN5107+a2FQTBB01zDpcAVyYNcnsgdzGfMlEaa+bCmJmRblzaal0YoO
bdbKbvt+ny+wi0zjtnj8e6ZEcysHotQYDDhEArC8qnNLZeQBlEa9dJFHaU8nubt+DmLRmeYTvFGU
tJLsovELK/lMVUV/KByDYlka0TVBACCWXp7+WvXPzq/Tijh7yiKVVWiB9eBHKC4pY/4/Rm+MZ2nK
LcHrVvTYTszXEVSO0oV9uzdKNn5hrw54f3b8Q0dq0xXWuDfBT25OqwYAdGq2uFT+5fXHXSqsUb6d
vE2nmtSJcZ7R9uODFOU6Tam2rA04dfZk4V5r9+8IZ+u9xe4GZqbJrP1A1MqllJuWTlH62pTHSEVV
SOS5JBHW4nj+8rmt8AkIDvMQ99Yx+m7tQj9GiHZlXJLwpkt/1kv+wqw1A5emdeWx5VwygKuh8RJj
nT3csjfFW5TLr9yePwQqQMbnqDHSUNq8JmXlPnqyhtY3fY+S28BAjK9feLhOilsrm6vw0ZGq4yYF
ImcyB3GNsiwwqIQRaDpB3UT8FDfR97ZoW+h1QI6ABQQ9zykeNZdX7gfl7P2RuT0Pyy2okRo3OCR+
8dkX86yvjCs24uyW/DkaZUyFmHUmvGezXf8mOAna6VEaMUMti5bgMerw22iQ96K8vk/2+69B1ylh
YgoC3PTmMJwcogkeFK9DP9VIzCV5iBoaF++A1j19mjBO2qhwAsiYo7iDzDf0eqKGcQZRH/f5VUag
ziJNM2b8iNtzTpujNl1kxApL5hjoDqm68X9gy3dpTZftb0mUFjZ6h+/yej4NAowHiheYVmRstAhK
d7Dbaok+bBdAkOdM9Dp1Il7qxVzCBQYBLGHAD+5TmUzbWSKRBL5xnf4tWNglk/ZJZqPxWdRghk84
xc9s5MMFuaTfoWRdslspM84MxsuH8BpYH5DGVfNVYOq7YYGobvtVoYpjckqtjEwgn7GbLVomoQeS
Tbeh+tmH8iD2ClRf6WkIG26+FFZmPO9HHIEMyS/gt7G/WJSgLrn4/IUvOmdhIIIl4vwld6b427eU
aRLttEZMNpcuJLvRF0+MLUVSHQ3mZVc+C6Mrd/5RHGQxiROS9dCd9IkFHAgdbBbtDSXuB6meYSFy
poNsDMjgzypltEk/1OfZeD1VXPL0Ek+WyfyBaX0M+r6+inaALOMagYtcVO/dJdDb6yoYEngDjoo/
Qjynkl8Mjp9qmaOm6y38gOgI64hxqZb6sT4jUxdv6PvOuIYFaiQYCvq27k9n01beuEmTn2RFSB5Z
oWPSX9q/9s9JWEopYrNQLidCIR/+nC2bSuu2EKijIkEApqa61D3x7c5KTfgEYJgS16MGARcuHBXp
x3gR9hw9kxh5zbRfdQRQopyYImJRh4NQujZjmpmQ8LDvr6hI5+8moiKwfJFLDSBJ+wTKRVtGV+A/
/LH3vKi9zCn5rtrXslkG9Z8fcTDrRMN1G94wBzORfqA4UjyTxndkD61tTIoIkb5WcGcsJgogwGVK
B1L1/OyJqMA113/5Kwnx1XJzJiyAMNxkq7Eubakf20CCJlUOy5lyf4UAPbTQeDlHsJNttg+pS/aQ
5z6mncFKnQXuLiQQvZedPmCtBX0PGWZN5WGycCWOld+nQlYCETpJ6ewmg9mGtwoNYSpL2kJGcyBv
p03GJvbjkC23ARcia55qrpXZqoLZJXStVo0iEi7o0yUKUlAQS1PIW8RuRk82lTDDLlj6BZWU8C0Z
JeWtM4u/asYVvu1pPw49EQ3bJKcU3Zz03203b63PDXbUQPNwaZpzDkObfhro2txZTPXLLigl56iu
ohbBpzFocKQJFdqiLIyDTf2CEtH94+bVmjJVwZfSZRkIFASL4S3r8fwxhXoEuAZua+xFiyl8lkub
BaHR8E7RWwTbJizXLZDPp6mWK9SxT0Ase05rNzt8bLP19ZXX4mXlq6FT3pXdFbhpUf+KD0Fff/jL
miJGnrTff7YyDHvbQAVxl1+ZnjL968RU2BlOiLSKdpXz2ZaPw3cuZzuOECTzDLl/NmGVcCHLYqIR
55iODmGzp/qAMi1vEO6jrOOjL55C4RCVJbMltIAsLpOoduQMomFcJs6Uh1FUFiDrKbvkwvTkuHz0
T03CKVTbI/9XK7bAeSNIHIy0mEL2vV59iKpGBZGutdnO4ESdCCFoYGi19Nj348FZCeZYok2kNiLr
YkB0/r1+/kqJWWcioRFzjlJf96i0XaZ1iCFWfcH2qmNVqi7zZ2tFjXyYQZ/K4HkiEsris2sxAlRO
NTi0hc+1wg+TBI/q9USE3HdzM+hdYH1vqNVSDD61060z4bgJJp0N/c34h6UxfHqC1CHEQv3MGAy1
opXGTkqznwksLj5f4Ek08NZtu1KdWv5Gicim3L9K/k9ZgXE65UZkihTtyP/asXjUJiPgsSAfXjNu
WPEFV5ynGUB8/2c9FauBohteK0AktKmI5ER3V0xs1EPQp/1pEg+cbCG6Z9jL+20IxQ7KJTK2y6/M
hFX/VzzFffBx7QGmzUYN2YodBvtXutAT8GcOgjFQFs5gmoBGU8co9kXG1mHWFRuohOQ59U4UClrB
wuIyAL2i4Ys5+NbAQQ13YPxp/384A8MbIdzBrNZjsRSx0vqVl3tF85AvosJ49duIG6r/E4fyxu84
4j+nirPc6TI225BPUu2EfKU/VK1DXGs5yVomnl7/rVDP9yzOk7mX1Bmz3M1w/d5oSOaUNdBVjbsJ
zpd34iKwEta8nMnMvb4kOXDtxABGLQPcS23s/mxdeH0w9jlN+6jaiA2wkBXiiPAxbtaL5l2Cvjfm
2mpNwUMzu+lqN9khbiY3iBxsOY8XwdsdxODNJkwOBB8zrRKK2o/hoRpnFbQIpnbFMqZ1Z4R94T+N
3yMQgPyWHkV2XmvFfjmNbWbd92i/nZJLwEnfek/WyV2E9LemOl1N3IkAMhGRYTGOFjs08bv5xMVN
bi9zncZTerAz8YxYJFjZw6cyS46y9nGXDuNzv+hnrrfnrGnIg/2Y/q50y6kPCejM7cE5z2cQuaIT
FY9RQoMLaB82t7ZyN3IsANIguf2qTG5y0r8MUVjwIC/NRphPjMxsb9iAUy4eyiyw1aZsmPd1v/eZ
OLN8OWFnXfNeeCsmd9cOzHetwqxtFpUQ1Kiio8R6Gyd7ebeNYpEda+tvjAWInvsdn4+MFywR1ywx
vCMv5x+HsCYkAFPufZ/ld9fQhDu1cxs5FHsrJdtKxZTJ0pB9NfSnu5SzYuaFQttvAskA0I8NefQs
Uo5LUxAbU3q7zY58bjOgV3VRoTVs29rumPJA0U9ad8l5kYJMhHrYNk9v+vrR8U5ImK994Ku72myX
vOxOr9rWkoPdY58Eok21m6ZtwhHeDE1x3ik+FViwZqiKLGEYQDVJfeLsS3e3nzw06U1/cQ9oapCr
CBdneowgHQIXF/f9Nf/398o0qUAwBTu2yhYwih7+r+2G8gcTIm7Kvn3SRqb2N6H1w/37cmp51w9a
w6Ow2gU40zckU7b0m2YR2B9XcTQDXBhq7/CHzamL4Szk6uLcGJt7NXVgUuuRYFULoLXKx0kvb0Ws
NA4UJ4f3vJUFiPQQ6eZviSzGsym6cvnNKIBW4v+spbGO2zhEQpGKLPTu9q1GlAJ/lTVx+LS8sw4H
9SxW21Y8QtAHBgF51h6zuzUv7106J4n7GeHWMDpUfbU2PFXBjRklj5XufmPqPKMyaWVV7Olmmybl
6OD3TDfjc91y3D2+Ov/Gf/nS4CQahLEmSCbihEec9W/QgSi2zAYsNrHsbEZgDwavX1TDTntJaojK
/Lq5C5kIPDSLXTU3nDHIta+1rSYeF4TTjK1qiT3PcRdlsTEuKTMCfHtz1XIugrPcaGCrYan2IcgW
ZFUA7iz5EpvOOD0HQ9b5R3RrXCPE+gwUZm2iZxBtzfjtD/ZTYf9yK3lO2wSddyAH8VkrVD9se+DS
XhriumRc7IdIRQ0W7hlQStYiACgfmvfGOSFcakwNgDXhu3OA6GejvpdDu4y5UqibnL/Nuqy865jM
NjfxZGXgei/etuZmDP6NiBNehhD1ToiGVbaDn7AxpGfPTXkDviRsZtYjMaQqaifc+m1v8VfBK1AH
mmbZULS6yhCexB8DN/2x4Rqdz+I0ZSt2fDqpeV4QMjebqWGBOjViu+wa/3XoSpJJQ0L/WSnW9tGa
IwR3+yN0PFm0RvBwlY4sJiDH/7ySI51XWo9p7qLdj4d9MR0lQDVk8m2BPQrMuxhkY+Imm3le5i11
JtxHHsBh8QHNpSIjx/fVtTPNdDPqq7coVFfsRirBqJzLhZps+x6BAUK1GLpMpGernwF/wivNi4lr
2rsnIzwwLx3X8lrUUPK3MRVr0JcFuinwEy10aI5v1xDD+/+M3x8v8xmTldoZn7/KKgK5neJf+gIJ
et/7dCoRBIrHhNocIRBRecFP9q5P/B3bs3XLGAZ097nUU9Nw3u8ZvQgglPxggU9wd+5tupUOEaSR
3rdn+4+256l9VKWzd9oqT7erTxzRTUMfmRcZM3LmyfwQlp7CXwCLGEFMwVrrobt7nHzj0mFwMHdA
FhlzhGG6SDs9rjvgtymqvvl0kEQ7+SAN4nJdoVtkaiWzvTcHCkNH4s2w3A/3VM/bEg+S6FYVCkGz
jbFKusWK+J5SAAiwCEwn/b3XZIZZ7OoCGXAur6cJh03oETwVpMR5FUbUH9IOdMFrmGvP/AKSeP4I
6iDakKOuSTIDosZwkKxHAiLzaTXFFQjuik/dr/+uBMQZl4wenNhN3jlKOJQvktStCmGV7eZ/pqTq
WE6AASdq7f0NtCOe228JUYI0pO+GGOIJ/7/4TKwU+2VEoGQly91ykwizSByV8LulbJNuAofAFRLC
5S6RJDUl5PbGI+SpZvCW19bUBW4rsraLElimpCjGCgtzgU0Li2N8sqRxI6V5HG4VPKJlREbVIiZO
Eh6ndnjHw1bHwp2zKZsHR2I8MmCueSRdKCa2gznmGHKXdOtN55hU0oJGwZilfmSVj8opa4P7XcdL
kkmZk5ADeo48BbqrL6tW9JotoqVlcxVfBE2VtZ53KWWNZKsN3zmtO3uFNc+Y1P2N41wIwyNkquS/
6CXazTehA6jtMyI/Y3MEqft4wuMQrlgo105R3hLK84nmh44pHRS7k3vBrmtKDx9bVWhAMPFdYwk6
6E57H4jhRt2Nh3IyN8ObjEZCCOSczi1uYBtexXiBUOUODQWAxMuw4PP9c6pb1S1xBSoCZg32rIGT
Qqsrmrh3Yv/TIqcGlvsZEiPNQs3UJr3W43JIAr2m6wqfSHecSeH0w/IPT28AphnBHCgzj6jrMbaN
Unx4aF0kQXlSRbZrXNBQcNxsrlXO3+gVzf0zGTfLfOseW8XS2rY5AvThOhkqckICcmvqZL5oPEjm
SWuieoH8n8YyGywXyMNzp2SNnG/pvtXN46JQM3eDbV/yEQABqXZSprvUHsv38Vh9TctBgXUSgmOr
zP7qQJEb0yjEVko3Bw4qkbOSOEDVXJ1ipkXfXlwpl/T26O1SqXwxDsklZgWuELhkJX/xCauIj5yk
6kaRNVXyvQzPykd5QvnlbQROjN5yztoU0D6F6PvaDv/JNCR5eA9ZBE5Z9Pc3qZFmRu6GGHqreXJ4
wE7u3nddCicncqPLU6XkZ01Veu7ej2+PRTTeCuJ8KChwlrp7RK1FWjB4d5eavrkOLQeCUKMOiAKh
+S+Pa4SO82GLV7mEgryGIKrFRGOYmqqZd7CudpsP/QAgBa2Wa4mTnmuPW/pix2LnAfK1GbABY+tf
fvUd4am1xd29z0MB2KNw34v3LtBtJudX+m6xio0uynfQPIFAPVH0ipGCmHqV63WOAZA6jyLidfDQ
D0seQn1ZG/HvsGousO78t3FH04F4ob6cQPp+PO84WXxoyS0snVe6zCaWQMXvBiM7PkiBs3A6z6zb
ezrQYSu1J3mmf47CKKwriESTcPnYoe4r1JKa6ewRFpdfGZZXr9DH+SAGMQveuTQAwUoiLzS/atFN
s1KkIkMHadTvNv+i6L78Tqj+EQ7OvaQ+sIBAhaFCfRewygT55jB+J2jRZkPEPfhYnn3BsXNBf6P5
ljy6+GOVuo/0YAR/pFr1gxw7vxTkj/LENuHXeoR4/ZSjcU1cJwdzHB3/GawTeva0OGIHZUgyWQhU
TbGj9qNcidqFQ8NKhhQ8Ix5vy3MaMgbV90V+XVr4zq+AdZpCCpfmBvXEHa6AjB7jftJGFofGuWHo
L+ZvJAqo7IaQLEyZSPsJ4y2QKBSZLaM/mLgzvM0eCpzfS5c72ucT4AZ+eVaukSHOnYanui3F+/8v
r0QPUuK7B8TZ68lt7P13UAhuBzsadnLObBfuDpWUsVhzgsbgwP7mPy2PEHD5UhRmZRr77KO3qo+K
C/q5Y6c01jO4zhAiFMLg4pJesfJz8jLRecO3efIc61kfAT/dHI8Zfam9Gg5a0OJkC8Z+WTnqMAbA
VynQhIBcVEfKwNDbNJlpfA96Z2upllXQSrHk27IWYvMN3p9hkRERRANjlFwKP19j+vTSvhTUYCKy
pb6g5oyq4tliceqlyA/51g7AsdeCouA1UX656iNlXPR/nYjOJe0qRx77WbgZ8d+olg6j7wq7ykp0
O5lxD2ZwJxY8n136+aUUY8oHxzCB2dffMq3qX5VzvhMnMCmnCUIa8cMlixNmvU3cco+DW8W5Vehq
O9XF2P24SkCJhraVGl13BAX99mX+JPPOi87ktMpgSfBt4LnTZa5lkKXE5Iy/XYogwstpjLgAG5io
4evRcoedsLZ2/06MLwHJ4qEB3VmAHNNtkPG7yVmV7XXJOE6iVZy3evQBWgS23oDZKhIEDhUjiKsd
sJmuilvRU9Jq4NcO4zm2kD/bzE4zjem619xf7OkRmlXikwMCOPqhlXgaFbZdr9Ywqulx0qS+iD3B
NLnofz9DR7T+H2kDFc/Oyi6RJHRzLJs9rs1dK18kl+ZN1negg5yScxLcV+XmEBf0hedaDgbKQW6Y
8p2Jx9f/+MjfZzDu/CJEhM6WGPpSSRJyr8H+Xxx1hmeAFfM0IvVW9NBVq3NssnXrALz4I60QN41U
Jv7SZZJrLzJAoaB9VTWoP84LKjpD937GCYA69wCn3h9Xn0D/sXgEjGWoyixeaswVPWJkawV3p/HJ
xJYoDSWWSvpdi/4VtBFPmcKV2fC+knpVTb6+huumzqtG9qhF5GXWqmKlX1K1XFLmFYEmQAC/dam1
IIfbeGP2QNFeWRRjknhz54NPWHfXF30I0eXD/H2wG/rQ2rKX/rF/E5bFGtX7f0pPF48bUGQNthX8
FSFnD6CePG4JtQMaItHMJ+0u6F0jtbtK246N+5UuBnpPYFyZZxEB7stBPx3MnZUnL9Oi2psPLA1e
oQ5U99vqoKE5P4K50Ek9CEx8xmvgUujo2YqYGguxh2qlqCcs5CEodM/9kXw+l3WTpm71gHSKp0DO
HZDvdJyF6YursrnZ+xQfCGPqUj778tAvcKHMH60LjVDA/n1dVLMZD15UBFu6hLABJeJmIii831lI
S/ELgZhdJQlvhO68T1kpsEnh/yu8vC3cBbyaaxd5hYICWihBZOWh+xORJxDJS8qP7oeorGwGwGcF
kbiGPVsbci8WCJecUQ49VBpxGgrhf7LmG6bqkNmAkDjg1pFpdFcXzdLQv8/fsufsAXWxfC+APnAB
XHrrFCpLJ6iFwbgiTtR9I6/qzvP7+1Pmr/D0vbBz+e5p2m5AS8CWB5uzUS5xEK4bFXUN9c7ksveY
HrglNQVp2ckXeTBoIwRB8YUfdXuwuDow7lOTxWsRHlrW34y3hTtIbkGniSq7FfAV3fz5xbARJ+bZ
XTW7fdx86b+1jM9TENnFGOx9Ohh1VxJXptq7YwV+IuP4b/gptVdkWC3r6zmW/GYyMkQtFvbrmo2L
V0aqnXvoo5W47/ok5MqWjEJezAXzijjxvyiY6JhHaAPtQmM3z9dLEB/1lLD4Kxvs4dCfVrFTDRrg
EALy64hdK7PPE+5jI1OwggBmUjO7QQezjzvCOgW1upq1ABa49gHBtnFRn12HkwYmHIBKaRbkMzch
chaVTTnUqgFGfW4yDNu6VXaH8Z9Uf3bAyqLzZ0S6aMG2SVaO6lNy79NFhXNv59JnAH0iDPiz7g5l
YCCe21UVV43RrX6c2dRRBYAKmT7Lyt0/sb1cM3puco/wocgYajukyRNniWLGsQ/MqdWU420uRt9g
gOlJNg8FMQfMMXAvG2fzGf5mFh6GK11RUm+5o7QlWeiFIqI6ob14fsuMqCRlb9Jct/NSn4ksXhbb
l1u+c6URZxdDPnmt0isoap2Yv9VO9SJ63n06JgpttrBymBVHbJno/spQpTD8H8EBiQgbHCPVCgyC
I5FbYMi2SjKGCZTmZ+GX7/B16/TgKRf0OY5DDSfDJn6eXfaBKTLF6eJZ0Gj37Sm4rXy8kfchkQKY
qfpaI98anMEQgJiS6hnvSHzi5JsUFXyLdiNaiBSD31AvOoEXrrHlxo5uUWp+MJkZ+8f4lPyzGwFe
a+gTfnr0Yv55t24+B/wYLexcPutEn5F18YfyDqdLnb+cILxa2aF2O9isTpL1jIJK+G2T3x/8ix19
Ut3qJMQs9RJ4aGpI+Bmy20R/AqfWKOSJD8Em0GB5AmOD2fQra1LNORaQgC9zgECfZoDCn+NMt+Nx
CL33Mwmkt0zyP8wDgYkbumWRrFk0TED2xXedgrpZX4qOApIDjYx+t+aAy4VhnwHHPkTm1rVID//Y
3V03oyDhcVvHG3A9qSVYU+nYVOQd2v05IuiUHtlqgCFamkhyIu7vWklIWSuCx4lX1B/hSnuw9u16
FJTm6KUGGsuLwFImGryzS0H6Cd4A39Bbps60m9I0DS8PVtJ8BsgOaUXBJwo5VrxxQ4A1bPXx84dd
zeNM7QjJiQQaYfETWhTtkWywGClitbRs9qSFCmqeE49RZ87lGIhNr8BG4GN3dsd9lo4Opp7N3jjH
BPfhAUWr4fHC764aQbalBp754CTFzoCPOX17Fs2FrRFMni0PPGlvRcK9PQY8ZFP/COejX7yHAwP1
8tRNrGB//67hM8O96LxaAWmWVM5wL6IdYFIDVcJOa9QJlJ4wUso5JOYR6+ZR2FNKEtFPWVaVcC/o
W6GU/x7qp1cx9urMRmImWZdy2pWgmI39UoKOFFugH5mpxFsO+iR5+o1izAMo+Yr5xJFbGsxCD0OU
lDL3x9QZd+aGONouRQsw4t+qp3ALeFusmaePM91BF49ZfIYWbZb6HtfuWhOtYuQtPUFSTw9AVeae
EvCwphkrGOWElOpOabZZPCbGEBlPVMpORtq/MV07553DDmSxamvwjCWzzDE1XM/+mAHav5w4lNzd
JkW/Hdyr5c89kXwt08IQyFSl/PDUPhBehhYAcMtDidYSDtyS5mXHfWNLWw3vEcZLb1388y5nWbuK
d4SM7d5tv38pRtWpKCE82mqkSRnHfbIkpInjpPTHt/ZHM5AlWtyXZ7fZAWuDyuLNlcN5ycbuL0nI
b0++RwxMmkDSOD57kySfJT5g0InI591yKuHQajUxfB7zHQ3oOUId2Y3VJHu8i8MUha97woosiaeA
b3BoW/nCAduiOxktj2Q2q/yznhrKt3OokgPDCHqiEe1O8QoGQCqXU/rtPO31GcQ5vad+Mcxr3xeK
Z7vlicedTny6vB/xz6KhRiSQjW3Q9Ro6qg/wNEaRoQo4lNXXC1Bid75AoLRB4YUcFtR33du8GMxd
RHr3Tcs0LrvxHUof+VTChHn0UsmKXBYlsH/cHlv0GZk5NXRdECWyk8yv/JR5SOXVu4mw0sLhpCk2
fYN4sRufNupKpdOK7fCYqbnuJeBxNLLrEVPUYukbr4g/927FwSDUDaS5YjWSv4y8/KZZGYXKn11p
uf56Y/DMkumI99DFTQEyeUERUZQpq6FNdk3m849QWw2yQcBsiu6tqdteLYQ94duxt1aI9XTWTDdy
HWl10/NuDKs3xL3/LB2lX35cfG2jz1wuK7n5DgPRrg9HJmarrg/4mlYoPrhEGTwAy8D4SIyj2vyP
gKtkv/MHItuHYODWzqRFr/Bz6DyyPA274QWtnhIch+IOJj7G1JPqyf8jI4/T897UEESSxNYQsfgV
gpCZZb3jeLP7bgFafOYsAal6rggqiSATruo0bD6ovACK5EZDAtU1mdwNFSts0uajtirTdZDHBtj0
cy2T+ZqkXq6if1qFwgHf1+mZjmK21FLEUxbMY0qyQ0w656LeObinSINypOUB6vTHC4HJQG+05Jef
SzAe3qHI2kBtYcr6hV9YOnBgirqGKwa75un7S5Uq6pSc/xzp/CzzB+BXHeVM2rtXK8vZeG0XQ6bD
mGy4HyIJIpNSras8FB62uYpMiOYEBU72yxWdpNf+xEDZugPavclhVr2diLtTas767p9oira89oXe
jxeYfii/gtFTHHyYl91PsT01KMtBSzTh/fj6lKHdrJ9/vPh9fwMuTLGYLFc6nI0guD6pLyU4zNJI
dDMoWexefZcVrSqYfOlI3UGY118wvfInyDwawzjYKNt/4tfRZgR6Za+RWS7gRH7PXk2fE/HJ+TYQ
sSxl9MPckxy8imsapuQZzYeSIaJZLDuNO4q5EAol0wWaxy6rYA5YbwRhmsdj1W2y8kiLya7r97hw
U457AIa0cQOAVgsBHqSwt3tbeOQs2He1n8G42B5Tf/nyEnldoiEYI5eRDI0n2rlrImaQcM6pCAI+
mkQZhMZsBu5rEi4y0U6cSscd3fR0GzFVn9TWXLZGP/ZPjtMWg3Z88mxgwYY0rU9A1nZ8m1AH7BJ4
8fw9KhORl4HJp2q7kDpz1q+ZzoqLY6dVw5ZgKy5g5qA3qrjle/9xlZMrpuUFTrGzcbk/xi/3mbz8
/70+MpZIbR1/1gjo5rOF3Q24rpDZW+DCDRUAYM6SuzfTzx2ZotW2FJsAPWdR9MDAnaZ4xFhZ1Sqx
6YozMJelxGB56XeLfeLTI2fkbliIe+ANSq0qm1PIRvvJATkfBtFaoNLRujBE/pjRIxrDUt0y8CV+
Zo7pNrlQcDIeVwMLJq/LgsnGTLU5Vkdgqkdq3IXSBwCMFmzw8V5vpesDL+/ykjO1RmCHq8edb5fd
bTS3QrKPOOaR9cIIVN7Iy7kCfWnzesLMVbzclFkp5vd8GaF5gDW9VZFGOsYf8zfWyqx6AbJ5nat8
dOzYMrpMtuZSEqAMllt+vuTJO+gp/Af8OWcBUbNh/FaBQ8KOGKf0zoea6KNw0SfeI2f9J9HmwaU1
LKm67fYtjvfVgPqIa7nS3/lNU8ixYrcFdgH3XVlB1MBCeACyphO0853Q0uZcGpbyzS8luEk+54Pb
9H9cQA8st0K7hr8Kd4t6Me2ev6Y0S1fBF9za5/8Xdquf6oAwdVArOxRnnk6ZNgmep/PWC/ZBMv09
D506CADAhGtdtwRdcLnJ5IDM/RDkhqqFSPh6Ko5cccmUZjEHxScuSx9v1+WFnZb90pz234DkTcsI
umyaowEdYLUzs2fzesn7yGncFltE77vZrkEnyhDwzjDCJV+VOoJZhZAsUSLnzL1UK+G7UmatoYYp
E6t6ycJUpWKBBXLl8R85RqHF1idkdro694SxV6j+76XW98hMOFGZ1JUvzGJDdqat193gUH1EHheB
El5TksW+Qt32SJLyOHbkny7jQcWXMdNjEdFWgRL2VvLE1dCzGtVpmqTeoQG9GHwv0LxNMmYQrgbC
GYmy8DUprRRVmCF80pK5/y0SdpWfS1PeH05dlvovPzf5/t73AqVNQ742s/yf53aGuzeJusScu8gJ
IothbEQDgQdsawnzQT+edbFmwtoEfJacE4ppJFiiIfCSPOAW3Pj+Ca7HXwGNTFUV05meX8EKQ5XA
WIsm0U1vwMogTfP/RXVWUWa7+uDSWjn80Fjx91ZKs/4+mOLxaL87NV4pH2UTieHlNli52ufytMZ/
2ebqRJDO+pq1aaYncI02nsbydUT6PFDK4pQVDIqXRwMfpeYBrjey87zbHPym8yUhaIm1nTfFQgnk
90mERR1bJ799AUg/4CPdpWqbPqt++qEE2xzAHmVn5QLLx454tRCabY7DDLcBHLuaYCwePEWjKkI3
N3DgKbuuQ5kqpNE48MXSRWKihB+9/45DY4LrJWjK2Pe0qj1BIjbp04LAY4CRJquvSb4xaib02zMD
ht+5uIk0z5PzZ5L2fVzxcp22IAi2Sibw69uknFNH2wLSl23YS/lO2nslkEw/CbD+rlrweUKHqfFB
Tm8TjDksr+q8L9D6a4jD2YUQKms7h4FTjtA4dzr13E05joPwQIylT2IbrFyxHcaHj8hdmgmUTe5Z
1QDo09aQNm1vLe+olhRWxD0IluoLnIG3RkwBBP9CaKVTbDA3tRBgY8HeZwcapqDIKW/MkRbTUmW8
olz9fu8EnxJ6hGNh6KT320u6bkwE66MGLQnsPntVCsp4r4filLqKi+sGw5krk9l2yx5TSD/uxaCe
W+E5yQ6LaJlDqkcusdjRePpZqatFipEd1/RP3i5dheOIeE0iSZfYL8Q2eQKqauwUl5oamP/6Z/9M
lFco6L4ogkKYDvCjtk/bHAz+ryZ50fC5iV60b+SSHOs2GesYegNopjzTrj+R718KA+w+xiVdZPHN
YpLUoTqEN8JIU8KUhKNMDGq5RlGP0LGORvhelA7IMPuN/JS26GIJRJAEKjz6vlfTjr+JDhgqBIlr
0+ABSlG0ZCKFA81hJbMZiq4DtbpdtrWy3pRbDzQ/6Uq9e7GNKCraX0qOLGooG7ld3IbCbTHAfm4n
SLOwQLieieemETIRKEg4YUezWvfBCcvhfztGnHDRvj5ux+SHOTwI6mKMhynPZJbiCyxIFkvuCum8
PHnaKga2jawyh2uqea+vHp1iCvN127YeNRapu1xdTBldLOtnzdBj++PB690/vUg7OCnM3MwvewgC
a8K7dUgYrlvrHKnnJPSLrqFklAzaD1kVOxgAjQ8NjX5oyX+m4wK2SmHEqeNJeyd7NfD8lCpKiiGr
/uXeh2WtrAmejz8of1ouT0GrcKdGJhMnazbM5P/tIde2MRVpErZz4+wshwALJcz3EZva6/5LxLnH
NS+JTfgnwOyQqLZdfO4q/LEXr1Mb57cesAZQoiX6OdgZV2NP4PdQj0ReksLx858pHgYZ4s5C2sA5
BPfi89zZZGEnO0TLoQjH/qYVpLhdHhs8M50lAmZ28yCkU93mvT2fyjqJ7/CRhCd34Y87VFm9jGiW
/MnaRhbfS/Jl2iq0ETLKofgG8liA/RJ+wC6ZV4AEr9GX7RB5mG8tWHdzbiBZfEAqPqrwiATMUiN0
2aivY902m6O7PiL59AMzLLlZiYbHPTTyrdArsZGJHuLeUrqCE/b5gouQXqxT95LsufkZgBFX3xqK
wvorig0hGsZj9Ip4aJRL4VKq11TJGv5iglEithBftv5dEVkwOSHt5xQTLHDCJxIXDUgcYj6CXUT2
r28HM/wcEuyx3CZqm7cvbLDPa5/SIunO/o2EHryHfxLtJUbaVPXgQjrjnlX8ExOKvVjiM1/XvauQ
f2NQ36Ms1P3IntbTNxB+WCGIREi23g9i403hMZMupRcZQzHAQIAqpK1IzOgnteDMNDYjTV1c+heK
CTjiDBUSYSMF9ALD8g+h4hP08tFaMOs2dsp84pCXmaFqhfRMwqIrtrxqC2jdv2PzzbQi5J79GoMb
XeQ9qDRP0N6Euc8cGYSGls8BYy+lId+q00ZYn5GyRJRwbuVU1VLOvEYaSiwzFpDL9t+wgxt5knJz
lwE7D2Iwl9q4quHoO1xvvjRHyIb4Bu/s2bvi7iAzcSlCcozyxb8nA+S15LcdZ9CxPYt6FOfkHhhL
NtuaLasUJ7rLghlVSseQNzX8erEY4dn6BsKTxsDbHKc3SnUttd6REHv/WXUATeIZ9Q+th8ZW26EK
OkX8vHiR72i3PNgIqk0AeINMmGO4l0is2N0b7SKAhz8+xrozyapLIxYWOEcdYK/7UMB2WUdSs3wi
zx6FHc9SM82vFd4/N1xhMa6QDCKSY23TUsgIEGjPuAZBnphOxjugr9yYBp+Ohr+ZBszoD3MliWr1
nRof4lj9pJCom/mng0AMynnH9CCpTYWYq0eIyngB72rxI2H71QdkvpVEgnbMg0JLU48JDjVFAaaJ
0zvqty+SfG0fUU4HJ2Q1zd8OKBsiSIuj1It2dJwTnKSKxY3dHOqn47D3DRmFp8Tlss6BVDAeh9Gp
1lKVsqyiJl59NHnGXQuVv9ZG9rmVm5ffbgQl6bXJaZp7yEKHCN+EzIXFdYmeJRRXwQeINapil3D9
YbDjFEgQGitwRHqYoMLJt9JRXLc6YUmYYanSvoBG1CnKbnynXbK+EA3l+yTZprg0RJ8m5ijM5M0T
h784Vr2FOL/f9BRTaYokeKXsPflCE+5r3nkfwIC3ID/VpM2pYyvyNKC8kzr20f5zQrS1+uY8D3ba
oS+epEhR6qiG8D3cTLGBPo4c3gKrveLvgOklC4mFLRKuqXqGCxU3/gaOPk6WN2cZU9ppoSidr5dw
vd6FJUqtkXL8h/LSJVUs0tHQEK1EE+G2XnMlxOOUqFkS9VOO/tEYFC2Uw0EZfVn6xeizHfb+o10H
IuU1HZvT5el/veVsAe75NeeyV79tLJIiFp+fByPgjm/N6jTJoc+Bx7Eb0I9WsqnLk01D+t2RWwkX
2Re9TI5f/RcewaGuKETBos9n62vIbxsHV5sjRwMjupJ0xHo71EdyD/qVsoGdzZgAJxTHzx1Smcyy
tuFuycToFS55WG+N+d5uUsvDaxKGFMNb0/9uu4JwMAUQgvKQiv+cIovykfrjchPacpIXBUOqCthW
6pyMbq033oYYDM/WBFDI6qHtRfLoqsGsF5aAqFqE01CnuN46kW2+eydPNxNno7OeGbhgP+eor7zv
+QRVpvn9wCrXV3Ty4vazikpoTQqQE3o9VxV22mdnlH4UImqxedNWanpuPq++wzgBpXola/qqPzfS
boBLqA6gS+lJHIMrL4WIt2Lv4wvG7vryGJeB99oDrEDFi2Il2UPXNsgBtikIdWLOUFY4AAhtiERj
xigcdzqBnw365VHw43CXY7ZNRR5gS+a4DKpTh7G3ARyUH56vUCo7nqByqz/FOn7+UfTtn3QI777h
Y9w5l2aJ09GVXA1JZBjVNVh5a9IEnmhw6ibMvvGwnqda12rNx2AFQu41JJR34pG4pjZdQdxbYBg8
O09VCu3b9JXdkuoKp8w225Ua4bBOKjG3EWdDpwKHjpZQ2MKcMkyXp+x1YrMNz9pN+XgXUTOJqe8U
7xMfwOvNTBc5Q0j42wA3R8Tzj97tyU16iQPsuD/4sTTiFEN4g9mq7FHY4K7LnVlE/eVKYJHli2AJ
LGoX0Vn+iyd+egppr01GNBAqDJOQnGdjLIu5li9UkdyLVbc9oftFvEcYlLrh1L8+OZwTioOjYyA4
/7HeiIDjERwfZ2ofVJ2noTvWPym87QTTBdUPJzSwmCLp3XSzFSzjQN4zjaWnD+JiTCSan4Ptb5K6
bw17D5YYb9tII/nSZguzmzlb2pJ7pvKL7JugPt3iw4faljiUzplJAwubVMSLMmrIMjKHqjMgb6l3
4X04tr9NJui0jWD8e49x6Cw1vMPFihJ0Pam1Fc7f/L7xNPdUFQCh4SUy+LbpKkMyfTrJAUaLBEyW
EHVVSN04K9/e0pkbIUQ3t5enxrrCeOzncmgRqAicoQkLbhCsk6wHEqEi87vNcaYvRdiy2vxqyrzR
vWMRIVn1ADNh7aiPI26nwQvWJel836ml8m5d07kwqiJpqfr6zNqqMUtXxT4pfCE8jScNoHBSl1az
tTz7LCMKY6iwPbd1UJrvk2hYJWbI5+AfRVkZsxnxj5pVHRAXgdixF39H/YHrgjPFOZXGAShOi9YI
qGi5SeIONWJpht5BQqblDiI6CM9WuEfDF0shJipong4HU9hysV5auv5M6mAeCWpBXzSFlKaIu1b5
Uu1Lda56WSU5tKS4NYpKjL08Q5qBIDV6vhlHHbJgbSis701sUbHNfe7WrxZlBMZQbsgfBJlsMAMl
WldhyER7KQMNFCj5NeMNu6iHCyQi0h1W3NTbsw0EALp1H4NA6YJ40wpGnZSGJLZs21XcAhI6XD97
sucHxhVi2oahwxwwNcwf9aYCVxdfimzXci6K2yj7OS8+0v7Rxpcsg6vIwC0eRflckMHmEDVodR9o
hHhpgBfm+RfntAdI4gTjAlVxBMAm5S519IiMSb9nmYVbZneaaAhr1DUbFpfO8dJSnYBoYkR0rZxz
zhoP8/k2vh05XD0GAZCcFbOj7JzybSb5o01HDo7+HJC62Ri12w0zyXpsCXCZ5Crwdv30UuAdBX9o
Z1npxIg0xtUyyWsdW32lxu9D1vW05TS5BTSszArkIi7NAZbD61quflms0kWWQ9D2ySfAVUJ+BzOu
PmN/qKBKsET68ikK83ehhDi+uYxxmGmZcHxg3yFZUpdSY7fIG+BU5HJAAwlXErSk6aBo7T4VuCHW
w264mbDnCFgaZkVHLmiC591TeMib+DRcvuan6UygsZeceGlYvj46Jn6Jfw4uFSJTEZdjgSrKB8j6
RQPL/cx0cI1BFplFIZgeXtzMZA5CWnAqxMC7vR6JosAB/U0MUOYAIW64DPX56gqoQ3lXHjFeOSQF
+Kn2bgm88aYHDdxQX0tDrJVL//L0KBXyjSbgy8FOLNRia7Rzw1vl1e8R9+kLiSnvmw+jCvO4BRgV
O1Nm3zKSRJi5glizPm5+hQka8V94T8b/9+jhdebWlDkKf/7yW9GjXil92DyU7Q/gey90cE5Zej7K
KOuDj6z/MghcJXozIlOopUWkXrlbS24NTGqtVHXlIMQfRRinT4dqmkkkHZRQrKx7x1c292vbU1P2
RvPFc1YgUdNvYHaQeaExucIht46b1gu0z+Nc5DSEeNGTOCD2pcmSC+jTR6N8yrjo34jiAMwyi1XP
terhFF3MgeV1uXYFOJGir4DJlzUL2zsJK2RluLaT/wVOeHlEJfyIYNr1WNY2SK1qHEo7HwpWh05f
onFRXs05ZwuWgBRD3aOJ7K00DkaHRPFs6tC4T48MYYzBxLr7Vqwa+R1Ssh9yt3Ihmr6lH9KJLSsD
SN8DWuBh7yN58HreK0Y6/l41jbQ1k98hRp+H8+Y9NOlGk0QcnRhoTQYB1hs9eqF0cs6i6uS36gEG
d+BhgfZV2wJ5+snOcKp8l6dwntgauJtVDihi1+9cYPCp/LU9le7fY+/Nw1I68d1mJ4mHNyTASosw
ikhUBgr1QxkwEnFiELjDDS0I3bnoNZM/UhdPkXqN2xy+OPE/cUoDqosb1LmI8dFo0hheAqI5x5x1
vBKbfjjUpYTC7AYcvNU8nQYOwySMAF7ruIAKN7QI0LZVrg8JMrbmRz8y7ODejvCWiwotqriPFwVb
3tzEv4bkDqauexrcnF2VaWmPw1IgySdgs7rycU1A+Q8x1Cbs24/0Yljyi2Y1AbLXDm2cTq3qo1PV
6NupBAbs2GmkbYxye90TRtt2sLXj9p0+McVDHcuTE1t+y6a3lPIU/Bk2KP9hhRKg9BpKg5QRcZ8o
uoHcrr8pFcNJruuVk4OWxZwjlPVwSWYCLJxsRlz96sCcTAWy41423XF7mPwPibdhqp+VpDCYdl8X
YeLMV2wQVGMlY6H0x1A6aNT6tUfeTKFpnF580NCp/QFVaJm6c6TabHxyPZpzISjmxRdWU+I9GXKI
Q7ZI4inGjAOqXKqXo1u4g4fUhXwfiP2uqJF1xUjSUaUPOXx9PyBBnhtUOusTCEN0BytXI1TnBfTn
qvka3/3l2otXAfv99T330VaXbAxaJpDnoNwuLFrq96antvbGWoQYHn85ZoHfZRrwRsqvKNVyQQfe
Zd+g3q6zqS6ReHxJsmKiorhx75jSFI1ZG+4K1cQ8RLlxK/Jd/Kjy1FA0fIBc2B8Bgwv0j9PF0ckS
yWH65sRYCY1QSlclY4Q/5yhxI3RyNul0i+uqz1df3dN94mGKkf+hgfUNYa2qDwRCF64hhM2dMe+L
nc/NeO5Vt1QZhzkv1LvJwMHEkJobd161rrwiV7izS/DGmL+0PFODkdKMMQJVPoAEoQ55509Ap5P9
qb/vo80x5Htil5LeQbSBh+G1Hy0RYGtQfJDHb3DoNBGcmObTJ0++eiBQJlalScv606rOqScu2SAL
GdwdDCGNs4+rrVwg2R2+MaBrL7VtLdTnEvOptOHvK9TmNXciKDPl3cLmY6iH3wv2Dyp27JTdwuxN
pW96JdqioZM/Dd880vpNH3ehytbdKgbKLoAOtvbI4Hl3oMJEPGMr/OPjFwEYGn7nbFQ+Eh7iEsRL
UMv6mSEQiBfWdQpFCq9VTQm8X/Ar5Wox+aWkU7e3SgsIxvvJy6VBrwdHBLl64u/SldbCXtm7aumD
mH2mbJCtPTuWrmaB8rxb+vUI8haVQ2noNXBjEL/Jgy93fVIyX+GaYOgvOnYPVqoor0hjNcO9LGcq
Nwnb5UifjdKa4oZJuKzoh0wesnvlQTgcWHbZjpHM4DpEzAIIt3X4Uo0Vmu21aXj79X9XTvOsIAyv
NYnsqwMQZg9wufwMD9/IISwc7GMgaw+t+bgQhQwlcoEzocBDw/rbdHyCUW1uqQOp3Rm4Bg4lNRAU
d772Yxgwed/bYII6x8OtG2zYkjelXBP5gVWwztSprbM9JyHi+C2E8X2oGfkuWqXuBgt/K9wlFGry
twiQOwtp+7BXAQIyU0V/beOrSVE1L8QH6TJwufaWoRXrW9sT+tTUaUQp9GYo0FQARCUYcz4KE/JW
01l/Q2mThLiUtadij52xbjWlBWBjaiQmPjq/jFeXHnyzkGrewbe9aFCD11A6ReoaseWVwsy5Iros
SRtYqGfhpqJSczm0Z+DZr1SafFNcS6p8Xdu8PHMCODvn5czJ1gHJBJNBm+JpdfcaqdZfrnlpoFsV
ajWgpW23MUWC07kxvtnOCH2PPcm7memYcwg1tFgCAkXYBhhwhrpl4prsbBPwa9orYI0Bp2qs3eGD
EXfUuRhXPp9YdSt/2YbzujBNqqeaaI8SEWO3drvUw11FMS+s4p0U3c+2IJP3Igeeh2A5aWnnAK/R
0/7SXBcLvwsWoKKTcSFcUNpvYTSl4rjig0vYONy7Hk0zZU2vHcpNHnH1EZKe450domLYLxhQrnUr
1k/YY83R1j/Q7/yPeSB7QrtUblMWAFJUsPhjasbps4qTMOS88jnmJnyPvacxRF8Lm7c5bnQNWWaP
SC/ppIOJWNBvPnpUJn2Vboz3a9LfaSWofz5HPrcUsPFwKl3mabo614TpC3pbCGu9tQozOo1SzFTk
/0mgxtw3xzhatORLTH4/sJbAPJBxERI4rFOpIycA1X4/C3bRbMdXk/5luRxObRIceJ6gUbgdIjIf
EH7TpSRiliFtOiqAF6AUFVF8H0MQDDc2j5IQXWqAESVTyhnA2DNNPz6Bk+q+fvhbko/uUcE9WMjs
nG3fTgbi+dmHZ+m7+jyAZcl4v6qM6Mn/HdBkEuNdaPwXPUSbvuQ1Iq1+XgVF+BinNZlgCXvqk0aD
gHxRKcJ9PgF8YJCwfZ1CFXLOiqp1gUWrdZsfjwg4BogoUcP32jDKd/EEpP7Z17KPRCxwqNQfOGf8
7p7GeRwMOHPuu60yTZN0XILxQ+3P+fh8L1CWxewtSBdJ4IOi+lDoRK27g8uRCtJBiEivY+bfaVED
NgT9E9AnDRkh69KfrKOd+8pGPGhxlJshrcsxv4Z+egSDCDnGRCqw1E4+Ml6VzXjy0Q6C/cuSu4SS
zarn7cfLcqFu4qfPHn4CFSSj2TS5/DlucDofvhxc9lqxrtLGnDXidl4z8Cdi8dYsi5dG0f38OrDs
aYn/g42qqfKkb5lmgZrHxC0dnXhsQT95XKL9dX/n2fEmdMCP0y7jCjVsTDUru4M8xTjfSQao780C
/Gt0kX3DDqxxzY5KujBUarahdNqQbVErwwRHsJgVq25OIXtPClNpj4h4dUtgGFGW1Ll6mu4Lg138
dQzPRUSJxtOmTpcItXjrwyf89dCGeO5j4htTlq0ac/mSj8aSFulLC2O2POrBRomE7FOWYih9J1UA
xfJ1H7h52ybLinvy/aTbSUbmwvYb5iMy7jYMilvH13zSg4ZHoHeg3w6LHjiQ7gYxnO6LYVY2XwB3
iNatVS0PhvP1hNmIbk9p+cfkcopXtdcUDobccqYSF+gzDH6YknZmehk2mnexjLK6SEnLt8MwdOIH
OzNoYoRI06mOwuTCkbN+4BjgmCbEyVrUSXW5QEG0wtXgESUP5FSswceWLxBJa6989xhPkRApSH+E
rP1+5DynELfqz6VIsnVJYOQgeQn06Mb9uwTdEb8c0J46zDDVO5TlhuoY+dAkim68bDEdSY5KTBlS
r9w+36Gx/Xza0jlGJ1xmVhLGXFBs4aSNckGeCNqjGqi+k6C61J4KniXBpFwshtFrKtkj2nV5Ur+f
rAruN/HwiRiMNBkjg7xFDKaQvVVmTUE/KTdJc7kRJiX5tdsAsCRBSOlBFk2T3zyVJivNTJkVcARF
e4LR66WS9ohmtM+vrOfAPo/PLA+SoiGp8LsWdOGsEP4K+Q6g66hDLq3BqSyvY8FlQ3m3zz/8AlWv
Oy7058DcWsuzSh/QBSL1IYRN0bM9LAXxXuYZAEb000Q+w2tf8TBQM6pw0wa1uJ+GJARrbQSSZBdT
lrZX46Wh5t5gaZY7COWdnkW+kTCJNT32aBvIE11aS1hMXAHR1vsPd9V2MKytVqEpTBjDGpYUt93N
upjiAdnzbskwPR3SY7hx0LANz3gut6iJGsuzMhIrdRbJI5xioGVHyvfrMjq48+CUXiKy9cJj9be9
Nzli+h2GB/qx9IJwkTutZaz4Go5dHZMTilbMvgaL6HjECrBG0XGOYXpB2okmk4ucryT3mnPKZIha
Bw3iCHRDvme6n0tdso/K3/OfIp6vLv8G3/w3CelVv+z2E8Czq03jAqhUTZarG09FI/pedrqRjmTP
h0jj01c8HReRB68m0/kSEqO8gx/i8zcEJDkwVVYrt72RooNC/hF8UgavDfoKmuAJMi+DZsrDUL1O
pBClwAVt8hIGboiJllbxASk8VljXCkoyIF8RbWC8LF94BgobrgzNd1vkimGs+taPdj716YlL6gFf
i39CdJdRNbVApVhD217IwxQJ94AnQc0FveUyB3+bfIZi3Jn+mAxqo0eir5Kq9YxRSubZniUiWuce
VKV4tQ3nXl2owTuodlRygSdP+F1cE0pXnzmziZkSiXxFRp9Tek6TeVKTQZfZ80Tn8dgmT8n99QBJ
MVpUrHC/SWc4Eemq+BrVN7Zq61xYOpQ/GG31OIx73HLGw03E+9G8WKXGT+MWHpxpGn0qX6MxGn7Y
zxI57v2prNZ+Cy0EYL9VnkcAuZxAtyRpN1/5XUwKIXhmGIcEFH06qW9VAOac+jda0depR4fwLqgm
0HrY19ew4tGo58PRICbvo51v5KLzKrqvGSD39JAVf1t8LzSpUkFp6u7fGpU5XKKBh980dwLZNdH2
kkJgPhW+Il3DFoufxjmpKiGCVn/JWLA40Hgjfrq+Fa7eGkg6w6LhkVpBI6hXAeDDa205BJESsO7D
1pGqdQU74hc4CTzMss8J6eUHltu3ZtLkOdu9Y5TrOTClGCksqO9ruvNcJq5pJR5dObj3+/ocn/kx
6n6pl0ZbV9MmWoyGExxMlMEVP1KI5VvEZPsTmC8kOqvagKjkmfKVOqSb4Py1UiByzffGTXJ3HO3z
3La/C7m3OUj0Fd76SeBIMg9wDCamhq2r3xFW26FCmLWDYRm/ZDwJt4LZL5tBdOFIYOLRSeu7fhOY
ZMXLY9Zcp+nTPNF23ZSeNYX8271bhTwm819M97Rc5B/+0yIL1t7qs4DOR9piuWnPcUUZiqqLieun
jji8ZqW6nyNUxVY5KnvhOzSEMYc9e4ATY3SVd02VbNDGZJkI9l9DNaWuqiXL5tgPMYhp7pSVXL9y
/0d1WLhKwZKJkEcmsZsWJTSymeJoHhw6pd2h5gnS0s5a0TGS7akrvm/E2NBq2KuwZF/UfN/Oo0qW
RHb3SBgyqc4beWWvdZXamFZs/9DtkA3fiZeN19e8as14DwODebyu6sn2tnpv+/BBKVj9Kweduv4D
nBn/LafY7cpRhey0svgfidPshhKroZ27Xe/9g/V2LLFzunuKvgy34HHSCGabkNv3CsuQpFpoWbs8
EXtVZAiqBjTL++MeBDls1XioSUjwIJ8tkyrBCYS1Z31mqZsb6w87Tn/vAD9kUg3flR/nP7+c+X8B
a/N4U9N5V7CwRRoY53Tz/p1wBdl9if9syf6rn8eC7wG/VhdGI8R7O5hnng9FLmj+AYI+HUbdh7DX
Dz9f8+jF9fwJIDwkglyG4Le6nWdGby6JpS83zHTKb+Y3kyk222KswXHqjyELOnZjzscpSUXFSDdv
maYjN6xQSO9hPHYA5O0wM+qUor11cJWay6tghiD/LuKpZ8av40xqNRDY9EKnJlX6lUzhmaKhykEX
mwlxf8EIyj2uB4K/00T2qwD3qZ+20O5/GWIeXWvC3CmGlhfGkompt7agN5QXj4jgQgKSxDIs9ERi
vG/9MuCpQI+X4U9PMEB7UWhpO3A9cy6kldeyUUEG/KufmWVCfDQTtFOLd4e6a9/y8i4cL+AYw83p
XdQP8SceGdoCOv62hG1hfFJFhUn+QYktQqD3sAiXVXOSxq/KQ2JVYy+2Re90NKzbwpNUBAyLQUgR
tI49LXyAQbxorc/Lnn1mY20GD5TYcJtZnIKomefaHM/siHHJ9BVFhwHdfJrm/kqFASzv37hVas9e
/ptPK0vdbDgOCcSqP8l8k+iReOaI+syHFu5tNm7LXXOnLfkwmsVYd3RAfEF4XgtbCbUoonwpbgOq
GzdYvj65OocEILoeC5RLa/wH6g897RPQ/8p/s9pPJqBYW393gyFOtIPESPN3hypKTO4JyoZmLMO8
rAQ5hejuXvohS/2S2CaCM79dspA2AKTCC+rV0/+Ig0TEDmvhamvBX0X3qBTVDzCN4J3w9yFh3dqQ
bvF1GNuortTO5UDrBYPgnEcwiIesG0Qf9BftewQwUkKuqJcNE9j7KbD99eIIxFkWWzVrBpLWreAN
6k4rnMIY+e+YEp1ApNaweStAcbLmd/kMLXFKwSddIB2c3bLO3TscWGLleEKm16Gbtmr3yjYF6P+g
6HPTzFRkkWWp7IwFo4BuA6ZMwbyRT9B7giEEqGEikP2A4DKKQRDXex38GpBdh9wisVzlvSr+AuAP
jHliCsjSIO3cCwa319YJpw==
`pragma protect end_protected

// 
