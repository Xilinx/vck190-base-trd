/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa", key_block
WnUYD0g6/qDSYmWHmuZSsLHluSdi9+myTeKuKMxZY1YiclF8fPuiqftouQOib18cBMrk+rhxXYqY
YxxEMkXifSggXUrW22+E+kt/etsSl4zJseXz6n9xUwZYg3xlqNjifu0w0ji98CtnXurauen1JNyx
O3YJAh7IDwn6xZR3LTGYOPxMj1rA3ndIEld9FoiPlSfzRSRuhh7ozr80Ea1y9ZyRdn6UvlSGNFWa
K+qWQ9v0fQI5P76f/h7qmdvfXu9BKunBkypsT5BoGjV+yipSZpdDPJFuKi8ZALQ4AfQwwQQ4W9Ow
ic2MhxBJty6sWw08okzuCC7DdaVW8+sh3E0SQA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="GeeiI2S+0qmTuse/FWjb6tqEZItAqGIcIYeurwykgk8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52624)
`pragma protect data_block
1KvCHb5eogwPJFXkT9BIC4Gf7nRFLA43UIfGTemoaERoVudbSjAfbNUb6m30Uqxx3NV6vEZVXLxU
NjV39axCxUjWByYwmwFeknoITG+yxwTIjztNTg82E72X5ByXSlMk1/fW5BXco5sHtHMisHmtoo8F
D5p0hsEg4Q5SAhV2MH2nI2akcNRoEOWC8LZjGfiCp/SCdWG5D8KzaVinGN2RkIemI1gorJ7WnTkd
Y/VlvKf80VkqTYzcQt/ivjz6GnvnwLkYKtRw9LAU+EkOq43F0FsfKVivdaWWJN02PlIDFdVgf6m+
/ETF3QC2PzTKeSAiLhrRywr/+I9zt3Y7nRwTnwXaf10wxKtsER5z4Bb3VmCkiGnpgZK1SS5oyLWr
DMlzn1Ade86tQTJvkAarc6PhJc+9KIAHgR0ESPgeG6MeVe2tOjxZBaBc6QJP6WXX+aOI+HnkxX20
u0sswKS7IYwQGyyPptEUgsyia81E3lHPqlaKxVThG01wAm6hfe31psmfkQ4eSL0SlARZQWJjJ7g0
ai+VC/ZkLBLA9pj7XrX9DKD36cjjUAj0Po97KccqWaLXMaRUXNotrTTkp2nLKbjn0ANbWz+uNR46
rH4dOkFjLx+PTYsbataEeVocbHaNeKKAlKRxqBF06t/ERH+Xuavvm1MfNhTKZy3IwCIct/IOyBBT
E7WpupHK6NaB3Ui5NFsRw08an0z6MgExr81qFl+dF4veLDKjFHed3V0snfBOXWKw2Q5XXpprmuqh
L/QvtiODIH0pySE1xn9ao9scBHWntpZ7vt0CdJVQObw9T2UEZ1TntmzH372SA8Qbo8LHmX0uXXjj
QYsbgAZTgLIUJiVZgulyUz62ILn+/b9avt4k00g6GxP26HHYPCUkI8L0p9wvVmfk1zD1QWSuUhJx
52m3z/C8ZVV8GbjMmP7OcXxlz0oW1zDehZtJJzhxmRgPbz8/4tPtMMU8/ifHOzcLa2TNgWWtaXBn
uU4vI0GUUZcRaUld+mzeBpZXrBhm0Tt2TVjxJL4HZFZXz9khAnnppqf2Mfoqt/APATw0j0HPqY5G
R7ya1CEQwrlrgwnzB3wApWv9FZY+gcPM6OL1zvIYteRwRTnpM6c84ARstrfLI4jZ4Gw1/0ed3bH5
fr3gJ/gIiQi9fC/ezwYAtYC+YqvTnla01D4OJnZLf0JBC2fXxceifyf62h4A4ziDAIK/AI0/m2eZ
onTfcQc0rWU848JCA6gUfTsyiGGFRPXZxNHpP1NkszIKnnIQ70keYSzVP1DXC8LwqglIUx0WzF2p
62Ho0sMXmPLv/DULh/Z1upmuThJe8HouHz3Mep9tHN3d8jGBB5mQCx3USEkJYUM58wQXGZgJxurw
/wMEFpMcKK3N8N7Jw/w3Oi9WptCTqNF3MZStcsRBaStPCM5hF11Tw/CQgCKvvLy+ONDjPaejYYQi
ICWBV/day1qchvCk0nzw1BflwMIDBKlkXejmV7r44wOYiFvf2p1/JkZB8CFFOUOQvT7YrbFF01iC
2Qd+Pb129B1rqcl0g0tUWPogTeysjJGTUN9LiK2SosRy+d44FaGklsfIqpnnOQLxouK081D87rI0
vV6ixOelOLjWrzaFu66l49/iGp8oBb5p6rlsXs02AJ3TGLYrz+6l45lhLQ73+MikVLNBo5iMIPny
jVuNCZXmHQ3NdHXfDTdPqHyN8nERJAdmjREhG0pcOixIgbe50z1qRkG2z92onHbOJgKjhjGvQAjr
V9qUwg7qt4dlX1wJYST4Dubp01K00IA7pqiZ9xZ18bz9UaNcqiwEACpMPrehfa8l6mIxxTjUB5jp
xqt7YXFiGod4fekd3oQfOUt5I7htebZqcjEfxXczl4sJFp2wWTxgqTgLQ5OTyzEDcRO8qaWLeh6S
L0eqcitQs9PaN5RA+Y6TQS8P0Dy1bFDIZsvLgu+EHNVMiDoFfvtBbIAzQu5p/JRfTn8CVqPBkU3C
tAzHNROMVE9Iwwqg4NHFg1vbrYNbeKmjKzGEkx8qgYPLXPsbd1mwuY3Rug8Yw0v29wrQNrGRqoet
Idtl+O7gknRLSj8EOPhgzzh3R/qHjHHopaaRIf7L89FJJ/Qn5tv3oJHPlPVS7/E9TbgJIrxUTo4f
2g0ScD8qbxa3XirnzVm6A+TvA1Rcv6IIJfZeeUN5MGC00LIqK1zHpx1eR5VoudbrzagT+QqoQJ91
l5vQHEQ+Ep4JOCpaZH/o9J6/3VS1kMSsMaif4IQWxPlFD2uw9wrn/JoqwoAdPoeuScG/RjS8K6EW
G5dXVqcwEoH+F8nMRGodBZLw1FLdyYMWLydMwHJo1fEuQx4W0xxCNcuybG14nIYReWxoaBQ9p12j
QeOukjrW51PNk6JnyDRxdaOOuBEcT2MyjH/xmhvmDWlhty4hwUFOc5sRBWlO+xrI43oDpcDnXKbZ
IgNwzTgtkMlPvxDOFJsveMrz1X2PXLMCSbyQC4GQB/7jVVx7stBIuYAH85RgjExAL4sfM0roxYc8
6j8Hmuhr1sWuD/HtKB1V/w31Zhp+cgZZlZH/t7D5WtG5qtAP8H6SWPdOQ1l2hz5P1rR7yNJU7NFv
q0r2GPWKVlvu+YTBQJmRPbuZU0k3ewAtQZhn59z3X8/RVmFqMriHrR7/TWZuee91BjI6h+7SyCdi
oKaTtIHrwRkUdBrBF9UV0fBxZR6m/nXb5PtHCzLuyZ5R5m6f1jrSL1/L31r2f9kd3nWrMUmu32XQ
PC7dSpJNER4w0HiENxDCW0iPAUL86JMi9RBAvUEy/vkaVPLwsy+zeV/7x/m2t/t06ktRJ/ddx9MR
G86Ksd8l/wL6OW1jmRhH4Mp7TPXs1NHy+Tlu0dxyTOjtq99BPBPAVyBJLO1DxkN1NXecTNnQkFra
sTEoKgb4+6PeYKV4jU0lf3OFuxm72ks7Xbj0Rj7qfASgGgDpX2nndFTEMQKgDpstnEyRclZa5c5F
0TzI4rAkmL9Y3+aKoRk/atOEelr/6CEQ9acQ5CRQqMrmFZ7cSk6p+QpPMvp8xSj2Fq8BAO46E112
od3QhEe79t75Zxc1RNI/G1p0Y2/BAgU0Eg6IhFxs8995rXOYeMMBpnUluczcOCyvB7tUN45CnUvH
J5Wu1DYnS2P4eP02ZmxbPW/gLVYlBjt4JsybDIMVNX+uFKKRuJu4lcYkCwZVnBET6Xtj80HtkpwZ
4kfVx+InSdko2odv1fiTDdYJwhfZFFbb7ovwFvs9qDXAczW//epa//Hc5eGxz2K4eaw8dT0j1Dsg
JoRbGnKdkLQpsmcbEN4P1T8afQ6mcTbNsxeG+UnclfEcMBsKQ+grNXP2Z35HgHvFdSpxYEbRpbqt
4TT/g7RPc9O1pt5o4sqwF3exliL6OvxPJ5zM8ZsHE+diYZ7aFkpVOaN/nflI497VlelkXZ440I2C
3bQ+QfrGm7IRslE3ubmrvw3vh4vBa7UwmIbU03zf8DhKikt7bPLfYsB19fF4PJ7wIHoL0kdG9mdz
EwSzZkkQdCZhpMRa5BNVIGYIxSDVP4OSiZqBXfs3MbnwxGLpQzSqeV1q7IST7TrQxh5HnHVAb+4A
dIF8trPuxzfv2jYfREov3D6KsQMoAnJ0DWFIZyvGTzIIEQu3hgR8Y7ugB411hUaWcatmIgu9UuPt
k6SnxkjyTnyZyBXWLTUu6ixurtjY/VXCI+0gnyQHMCK/fBjEFCE+XbUdLZQvWx07eamzsaK+1nI2
KSBUPAm4KnRCKUoyvZ7S8dOl5BZ+2wcwQQPLlDS4U81Tat9fTY54BUXMcHCM8mvuljS2KEWIXoYy
ioJaiw1kG0+c/els+Vtu+scmqn6mtNxucBzFUxote1pq1jd4+eEcXihk0CNan6e719hhlFaKi3X6
ZkgCT52v/P6EktX4kymLu8NCHYbmMsVxzlzDbYEvcDqEbRc+ojndL0tgeu7PTQ6X2I8YbxqQEs2M
VDl4SjUasenG2AGOpLgPqswew83Gs8E73RoDL8B6TEL3cOqZuRuV954jxQ/Z4wgEn0mVNHYB06VD
lgW+L6VVCcoZ1URil8Z5QtME8JzSrnM4qdQRWmy5zBjuwsKA6k5qV5DjzyMiXSan/HRBQp0tUN5i
xYFBOs/LiRxmlP+rp/2Q2/+NE+r3rfrZh3GVeQkOPi/xzA9WvVwrT0l2hVqEi3WDqIUtMXEeVEE6
E1UBxpbZbKGKL62QGvHrKdl3T0qDqEIToT/gVpyyw0DIEHvsTRCpqMxDrsELS3A8Pgv/SgtXuN07
/evMPQ/yHUMjxF/FMT0Gg7aW+hqpzxtT3E32Rk6XCkO/U9Zpk///K6aO+MwId+GyUd70CURjfLVs
BABeUC1BK9Jd52Bsnny2OiqDVutz65xLIykxLxmJz5OAd6hRQsuGH6QxAnyVuop8qqe6YTegao5+
J3UxKGrquCYdlrLFeaaKk2mSUgVpOq6RUaFzMDjJrNl0Dl5EZ7RU069Xr1Kkppk/bBBlSmH1YRtE
ti3ruSu40z1ccMX18/GVQJVrdXUycQyGqgWIjjOajP/1KrkQ96RzOslKl/YKXIfEjGu72QVU5d2R
7/5Mm9AOUzIn7eFHYAGIdpbrZJiIBEvd/aFZ67zNIssmDkMoH77uSDGu4oS1Ty1lc7qMe8mzv66r
RexKX0INw8ByG4D7qZ/15ocpUgH6mDItH+K1+YWXbEaf6biRUj+DxdQ7EuyQPX8QkgseEk3sIXd9
sRZgnS9yd00Cg7SSpq+tzOQ9632k6EMCMAXmQe926rNg6aThMcEcUpBLzW0wJ6waJdWNS9CUVq5X
cXTlSbmUOu9BKEqixR2nUfCXG6I3WziJXGTdTQG+WNIYNC79QR0zErBy5ZD5iok5iK91j2tTPE3F
qCPx+/FCg6t+Ffjki4Wk6T+rL/A3b5BXYwxdd03ROKX+qtid4TyYEc+00ZLMihlDcd4qc3DG2mRI
tGVstU94Y/0QGxRgJ61tFR9NVlGarKIYYeyB62879Ih2giXdijMYcvlVn23r4OcFhpNoq/hQVmbD
iSLrYpeSErCkb0wtiKfOQfSiKIVKN9hQl7o4yHWtV4mkb0hHQH661V2183zFYQv8+pAv+6eOL2Qe
EBUO3thnn40SJxInuy7P9bSUQAqxAwItxrjPpcVvh11+OiCTi5tO3t1zlatkOU/WyAK+2dVVwsZZ
epSEPRewl6ZlHfnAxOv6ZMaNRLmRAdQgHYk0Cps3t28bCnWAnfGKFAHFa2rU+PMDrc+NHnsCPUk1
YZTowP7hpaa6EftDjHlYNlS8H7ld9lVBWPQiDBH1/a9C3xtD0Z5Fk6J8QkGsccvZC2kxBrfa9RZF
AOcjfCoirSFiUXc3frKEaZVurT8kMkxLVXWTZ0YYnSDB8NAjn+FQltoHH0Q2e5GlFIthRe1d18Dy
QG0kchIeeyHjK5fd/WrqTB0akOwgIMWpkt7zqDonUp1KoWpImCzF0rewGmcuOomxSz6qmoCaMlCN
TPywrO+IgA4sOjPszAekII0H4W0NdTupIjuAuKaxDauAmHI4o834+goUBUZ0gJRhDF12mItbId6Y
gcT5ap/KieYtXMnwe0cUsRKkiMsuUryaMqFRYONV7dgEHBE7qMXbbIlentDk+I2N7QA4/1ML5DXK
VmoTaOTuDfOR9SHm7BrMmhLTUfmII8nOOsZD43vD4+2fnp605WORypckMFUQsrTbIE14MLV5aXaZ
m0DTAqHig+ENL6s9Ls6QSIPM7K2xK7f95E2JwZVybdHWZBoVsXRhpeT3fxYN7I2+wH5JvSTIp851
SYVlsSWhjnf5qB04syz69si1fX8oXk3PiPMfQIvjbKuSFTYajuaXbkENqI0/LUULX8BLkD576Lyu
EsP3nAZh/KK+yJSqybnkGUoJu+PEQ9PAT1ZLnTUFy8/zLKX5q+eTxHBguV9i60vaYJybaDiPjHdk
k1q2Pr20hvd7Gtg+KAKd+48BPnchujHpQQiECnPAzbVRuSthEVOurfpy3tSM61gZcSDppWHpe0m0
iwhwppMn/AeF92qU7AQQWk/cU+FcwRTwwNaN+Khg9FJOubiiIqw+pLk6obx85DGauS90n+NeuoYF
t7Aygnd1pUrXnNdeEMVUgkfnl+4iGS65c1WhM0F4O5seZwrbK50NAqvy8P8BcDiPZVvobPmQDoKP
qK+LWGf80a4pSHYMRx4CyrMIv+z8uUqBgQFOZTnhVtVHYV9hana6DKSyFvFlxLrLR/0BGZ9UKQ6Z
4CF8l7tz84yqqJC73wVZP0wqnIOorahClGX8+QJ6F9xojxtlvGwh37gMv2g4qK8ujhV0WQNxwNtw
2fuvkyMSShZllNHr9Dsc8SDCGDJFQ7kv3UwbXViSACw/WQmTtSDATXTK/xBayGiwP5Z23QaB8ITC
PRxtQ7Fb5NDlzNTEouAn+aoRxm+3c5hDstB4te840Ah0+WH9bkcW4yBmbo12dnKTiyc9EcSS7K6s
BkDDkIofWXhiVInRIom+nlDgnyugi9YP8cZVFbGrGU1/TCsLArGEWQvhYtx6vKFHWoJOhXb7MfxF
QT6pn0iYih1Bxgu1+NKb/E5dgDR2wlUjCf5cYdrfEIdJJ3WG00+squkfX244KU9AZuH9OQ6mC+BZ
TnIrMfbPlIiJTn/ejJOycG/KLmdLS23ckm+bH88Lc308ednGsdzbb/hUD/wY4UzD0FxFwXeoK4Uz
wW5cuX7RB4n6qeMIEh9hw0uTpCZDJDnhm0uSWuNKhmrAzwvDscpwdjnI8XlpuDZgfrjRzWYEyXg8
IrUe4TWL4rTWL98TQJQlMq94ClZENB3eWJSC1ppZ07Vseqb5LSODXlTY5WUUrI3nMATsIHnEjpCB
B6LcFaMBfrLObNbjA5BjGU7Q1r1dR4MuTy3bqSNx/JN+dNYbPlnEYNi8oZ5KM6hpclYyiBHWi0sc
+jG597c9r4/aFrTWPCyhEQkYbvtDwzsfQGvSPpZP0UneaZTjTw8pCwh8tCp0R+uri91qaQYhsW1E
4xAoGFPxngxuiD6pQA8TPn6bLsrG93AS/LAui6eHNQJam4RzODaHXwGcnSC9Q4ZkHOv67c6hyT6p
3zOFeu6+L5+3nJgZAplxGUQuJO4AfFujw1ngsCNPCUd3hnopzn66tvv2RqCag/Qb3qVZsjCG4tX3
aaDsdHvhTI5p+1lx+KYH1JKx7hv9cqTJMSXV8SVU4h8yxyGh9dErpmmhJBQcxDsRQMGUQCxV7Hjn
RFUUqgXHYYAkmZLXnHI0+LGK4n5naYVoa46ovntBeaCViNoFGOTL5B5iQOqVcrnoA2goGicZ5qk1
lK8CkYdnAU1tnE92mrnoJMa2EVUZE4bCt3TbbCTDUxh2KssyC+QjAOyxkNK78d5oiyGpvpVdxYRO
xr/pWLda7FF7HPZCcYmA8ZcU10Y6ZFv/0ke0MGj4z40O72P8dg3BR6WosutNlxij+9vHQNWV4SP/
QH0ZCv6pmWvxS0Apg/dwnU6nTfvoGFwccVr453JHaA0pzXP3J+bfywG4G2GutJIwI37tNe/D9Kji
+CvcSTiOSMX0a+7qxsmSIF6m62IMqMWtQAvkH2WN8sUBm3W6jnVM7lC9s4lAYN/HQnUeFoEzTKEn
GGa+ElHuMZ4SdRHt8mBHruma1A5WRA8kY1a2qbMKMcLzaq4DWI62kHkBPtVopRJAiHiYEeAjX1yi
SS6HSOR5LgBIwYTteZtCI+JH4UgKeNrXnzj7FhALaCEuaEJHKLhEMikmX2KfCTF7ivHyA/oX9vjK
/iEpkXdIsEuFLSdoKwg1FHkSP7nst7SzeNWgoazrr2mqmwnkMuAecgfvGk2E1Eg7W4Drd/1822Q7
BvUlqGmDocJfvSjCpXxXPYZtcD5SSRk4oEbrlNO2mDQ+5r4i8daLgGByPpGd00sfsJpEuus0enq/
YzHW79JfM10lP83BEHWzjsm0BEH1K5J5q9mv93KxN3RzLczuZ9of/ojLpgy0F7XphKGPoc0d3JLF
0OaCRuBt6F28zwGpNnImP0aMF6NKh6aNpIKt0m0VaYuuFvFlQkdAdN1HSFK4l+Xli17GC1kAWuCv
fILiV6SAzub1mBU27ZJjp63Slda8+CTw5PeoWou7F8P31WdhiU80G5H6+47pj6uxa0fSOoujBWqs
jZZFy/haKbund7Gkaaiqgqycj4nnpt1fbzSyG8+FXELt7FeEI2LNwYZxvTEAxbfHJYbVZWXVSl0X
WzxIBGN9n7g11/kFyVa3B818lNeXFRULazPqQR4cuvFOH5NUfeSqHbEL3S+oMz4HOW/hZcHfwR9q
/ZBHgkrsCG4lpUb30mozsSlAXX8DyGu1+zDM0QVsiBdx8WdcaRRKZcnrEFFfCg4w5icwP5ic0CvU
8SPfSo7JoYxnB65+frXVhJfoxyLluy9G3+l9mVRgYpAB26+PZdh4BNYu6krw9WrNihx+nm+RSKV3
oDuyiRqRbWt8vO8KaHzl/+gyU+X66j2S4gGI4BPehANU/itOQalSAUK2zdAF7kNUbl2zV3wqobLq
BTifBqnVO7hBrfCKxce+eRNT4bQ1wLdm/1Hfs8uMANZSeN1kBUt2kBuotLYEER51hD0mu59WIe6E
fzYwwLXPQNSkv3UbZQXD/wjIRDPqDpOFl79MFlZTby03XLhu56O3TpsrH1uxLN1BRuX6aujADAU/
L0ngQJkPoKXTfvD6A18jCjujc2bhCmtTnAgekXptxTCNlkvGt396rykj3v5NctQixrIOqWOfLRY4
2/sdJR33VEjLjZlqSg8/RAcGnig40pZT6COfzoMRQHEilncIo0Y3Iyeq81c6CYS5XcnGKwdV5nwB
5NygXul2LxlJcYYOanU7+uiUa8b1ibRXFKbVaqXerypcpyVu3DUK0MvGQjvr2k0scAx8Qmt0k2Dd
avKv0oWHmccFLQ/QrmdreD/w1vRWohD8AuTp8mgJwQnyP587Bzu+g/mUQ3nSTVvYNB3QlIKna34Q
zL+Tl/730rYrUwJMXP/7pReRDc0/8Q3Zc2Ibz7IR0q8FlGdRezr2mKsBydAEnk97WYc+gTa9i+Tk
P92vPFM1dohzRBYjwCA+GK0tx8Gwe0mCKIjxbM08JUrVIZqOVTMpp1DdSuHqrs37z37SrifTIGm3
hpr6+DPL46qKMEw6iFK1iHEDFFTNmJRlifU1W0QV3Pe7v8Ik/DT+IzHVVAnU3wUR3+aZDoaGG97D
xknlNtH9Z8YSNkbO2mHvmH8+MYbck1FroTQazlSw/+o8GExOJiSNkcOnkhaDAhb3iACJ3burBomV
vQH6V2mwJuMGIvXTkrLaNPA8+i0l/8giy16rFLTva3pGijU2xUSwjbpL7BIvZ1In9ie2RvVxy19H
BSTkIOuWZFJ9akkGDrefAvKJ1jwxBNG57s4Z8a3t0DNBpGLQNmcG1yipss1EfYYy5ENvTS38h6U/
EeDtV99o/lAVSTAk7EXLsRFXYOP1o+vSxzkLyBp483AwzVYMTYr+aHV8GAk1Q8USFLfGGWI14PXN
4oy2rKJ8fmnnrDo6Fy6VsQTcYjMLFryRRWAMxRRe43P0YgG2aKet1EgQXZ8tPzpNavWpeHFTY2Xo
i3Om1GpzA7O7E237QE5sB2cmb4N2VJhzg+7WOeimqgdjwx7TJR5xWZ7PIXA182HncOQosLJMq9wz
j2q4P2IOuLUO5yFcPW+W+kbHPswzTm742V3/3dYvgEQviOTlcOhy/Q3UdnPn6zA/X+RewcsEeDYq
ujXqwvv5GxWLYkUuRdBz7ih71wcUPWFNJC48SpSr9lI0K0HbfNGxpgzzUqAcnpB1mjpwABr3RsLV
gBfscVuOd1tKyKcUs5nbq/WA4FOktPs0OPXqtLKhtJ1pjLmqJ8NJ88csJpYC6qL1GA7sSqDmkaC8
CnJsXaSqdsXQLY+WcNPYg6cf3M481aZOP0IYVVly7mB0vtzDqPFb8JLLiw8zL9DXSobay2ItqqjC
/IBYa4mNn6OBfMv48mnbDETlntFM6dRPfs9R0+KxUJUjIMZbdhx8BtnE4L1ZRhhUhcF9RfC5kXCy
fyWb4oLcMCgNS0Fgqzzo8RsJOcV2nnhsiQaxjcdmhETiJKNUQp4d3tk4mWsAwSJoWeF0WvP/6LrA
TXpHvl2+IECJT4w4I+fgIoTIzhrnm8HLuMICclIguTbEkgVPtUmaQyFEFw+OkfnfpFtVFYO5wxxz
YZRXZT3R/JTaFD3XZ43vDyHBMbLaf9XYjC/QQ0N8FaXpkOUZEi1cIbArs0oELZs7s/UUfCnBqABO
CGD50ElpSz/gN8DCSFDLcMhzGSp8Jh4jrIac+zB1fd90XZg+rpj1wNylg07g2Wn1tHgRSsApvxjI
wZLXR4IkMoKY9b87rUqPQivXq551ws1hUicHPdosCkAmWwcb7c5EqNBE/vg8yrrzvw7kcWwF0CpR
qxDyVDuelQKYb8vu5ETp/7ezB0vxJrvq9cUMFhOYUTE0hAlenz5MFuSO/sBpfsyMRlzKL58vD72Q
lpNhwd6p5779ZEyqw49eSTq9walSU0eIcLnEH1logIHMJQUyVl547lWIciet95gh4ZwLBhHdhzmp
+9fzg8+3/DL9UHBLUCLJ/gVH+malnqK6J/gMu0SGiPXo83yQMxMcfN0GG6mmnTkAOdIL4qex9SA6
3IWBsNX/2jdhPK5A9yMRxf0sKr8drBDM4RjgkmBZp1CqH49+jigqPvHSgbC1eR9wmmNB6nTO8wKV
2cJyOp4jdaYKhrW94F118eHzrzBDXJu7IJp0ADWJxnYVmeCfXd7y+9lFslOquHmwwzOhuxUySeJL
JjntOrY369uN+Gs7Oq1VNQBY6CYK/P/NU5HFyIvVVUTympBQf9JjaX038BtmDE1Jw/6Z9KuZnF0E
jpniLANzwIbhteCi9t28uZQ/NWSWIGQme2uViTQKhxewHMArVRBBahdmHlZX7mtH7S5LUizjSX2y
3YnfejCjJc9LReO69IZcbyKqbE6FIAXlfNqA3VbRSDqp836LcwwgrjAvgrPR5Jzf4u/YBxQzyfKv
IBM6YQ3d3OhOXr/5kaUKxNhPRAj2qqluhblbFsY/WkrAxel45B4EsEpP/SJpaLK7akDqD8vvepKO
1vG2BSR6VHDzfK9nOG2CGVy7KiMAvW3ljWOk6qIoRgHKDEWCQl58sDiRvP2SxK0QAVcs6JfbpVkj
Bm2iR1otzALLv+OIYQqP9nhy56l/UUXW1pmGMMpmXWCVAbm6UWBoaQ3AirCpeuX7iwetl/gg6ROV
32ITFsDux0pvJlcCOgxfpQV4T89gK8S/z9O0D4vPZi+lU1HBS2bc1AGOo0b3I7mxw/fufMJm6dZH
PvpbdR9RdLfI/AoPB4kDcL4ldcPPWqcgNff5Z3A0YnQuRfb9mYZqPieGeHN+76dBR9W6RxlA8OiB
12NYQkfBwbFUR0/++wIk6baFSVRexWTKkSeLqhsz9iniVFakTlA+zWiGUaOJzxuatQB8BihiJ4iw
bGDanHLlabESHqZ4QIlO3T5zXyPgGr1cXrRBIKsb/d0593E6ESozWG89n+gKtv91gkBRZqXHyp5n
uKLN2YTDbLDUC3dZSeEQxmMLpl74I0FpfWW2Wx6W3YdhamXJNzlGVM3XBuyBnvA4if91fY0wSzq4
BEj3C+qEQTJJbd72dWYncFO0Sv2DHcySw1uEs+Vsgn0Jtcrr2uokbSPGiZX/HZuihuCU1e6boHA0
nEtqiw38JQ/wj7DqI2ai44LVY+ElZn2E30MqEeW1X4wqcxTf3oBD5YA7VrgHoQJKiP5P57jY89J9
34nQj6LMygx5Ln4DSPi6vVZbk9gVel/HI450BWb56b1zsxlHma0LPYKJjvKCHUpAt8U+5moaEJLs
sPfd5f+OsISLUQkAm9v3LzVnRzrBi91H3lRMPr5cFSO8uxWAkFYztdVPZ13x1l5BQSJ+WNVsC94Y
Z2iHRVaQioeeDBm9w378r/8UB+ydLynU8+yL5HHJzk/DOXRtnmkRjBtqFZytW7r1EEzFpLqZkW+2
4yIfl1qjKxxF49lS8MwxKzibGqUr35bEzgft8LB3YtA1RDKXWaMiff7L+qZ59TNhlVH69RQzHpel
tn3hI0/GdOJkOFCy5Tkl0sIADjcPxEsCP4khdZeDy65B8EzPj+RYGFBFXS/eii+FYvvEqlxfblLR
9pnBAIZtwQmuYw6Z/Wgy3Fb77EX3HM+Pi9qBTa43cOsEymcPLsJ+lFLAUMei9j+I3+U9pFsJC7+p
taUIhAazQ7omSDUghkx2RnXq507y/49Hyyv+9PPBYTOLx7vVjEqYKyeriFIMFKa8epfdqDOxMWec
uwUoXkDvWakRAA28LlHK+jK7R4mh/ufKERijpUQh9JzAo2hjg6JMkdJpTLw/+SA+r0DrKLUVvTuO
Shuo5z4F33HzdkXdDkOrOI2TDb2Z3tIK/c5+zX2xTkVcpdd7w5m7jjDR+nfdyeCiUCE4y32W4g0N
lU4+ru8KSAca+05QKw95+KcRTaKnByd8hnjg6B919opg5d/5oFehEoQq7mN6FSbnfRGTICSiAagi
/x2Q89xsHBz15xzyyyEUC/Xyl58GpvjCT8HPnNTW5cG3uchOkPYSuyEN9ZrCmlv7vqlHxtq9Cgih
VmmH8A79grFx/an0L+kLcyrtHn/D8rJXshv1M+ruYyE7SdFRWhBXkShkHnnqlTCyuTY7Y65RY/vI
TxW6eLikPUTz5iOnbXGPNv7OBGDhMWeAHL1wVQ5+W2CgV33B+JZ9xfQj4ov9yPV1Rxxdn8QG1sR0
GA4JEEoPQ9eGBQOyVI8TxnTXy5Rfop9JqVTZCnmbKa30RjvbgmUSx30mBMVvBFoq0FxJ0g4+ViB6
7nq2nnbfDmV20xUeMPK9Cl8PaVlBA96UuN3yEQf7Nn+Qq/sC6FyFfXFA1Y73BtWokkSRirHFrYQf
Nyw7JHnbJDF9m+X+vzaUZ2KzCqVMhAYm35sCB4swnT2zUWmeZmtO1X/nyYN3uV4lfRh88U2I4RSN
+W+MU/Pq/WU8ieh8oBmPDYfJJQZ+0Sx4XmsA+pvhtd/zO7z+bkFVREOBJgHdlRUh2CtBPPjeXRjn
XEAnTubGVoI0a6bX1cul4ufjXrioUNzH3sEhUIJc6KfERfVXngqKU4AZvM+C4TEo2/Dl6PXTvH7p
iabuIdK6aO7ZOGNfwII+4zAbH0x/ziNWoD0nwdq5p4M8LdcTQDT0j0DWg0mpUnDv+jTL67SHdrEz
nF0qLHgD9MfAEyzOsgV113puNxazBujee+ym3p2XvHxpeN53CCGDkj60Y0Zc7QJvSN/Zb7AXO+h1
lSE0u9NIqy++8Q9d3orsYKSFx+cijhHZ3BK+RJFoAmlCC3vjLhtqsb0KPT3xdZHbiIJlQBwuhvmt
DSHsAPvaeD5JC/wlnYjjoJGpJTINryDvCHN7mFVa8CmJ6V/bocxXl3N5m2QOsWovM6JIeKqCUQ5R
HklR4apEmahdYf4Qt9U7+ETomzTypmREtuKMRXaNbxz4wIb0pGhh88rBdgC/cuEg5v7MZ0jq5Z2M
dYdcx1I39LroZWTW/fR/WC1HabTJrEZr1MiPG0LjmeMlrivC2cMRBG4S+n5c8GzEFDeplJtpckFD
4T4LIzTzS3FBukwldPXk9BPofm8ASdMQFxx0H/3Lvu1tsqQafwcdNZto5qTTHLMuQGMM+yB6r0Nb
IJUdVzfh3mvKaSXEpITplR+pDuZU3QnX0Nrhhbd69/i3FiwRV8SDA2AJu0EczGpelVVgnOrDpNnH
qmcbTJBoGCMbCQGnnh4185KFJTBLlkIcotxBqkzQWUE8P6YmZDoljaXLnIRXdft8iXKKbS5eFWmD
o4lDs3szgt+MkN6h4Ab5n7fR936LQYKexXnPd49XGwg0g+R6GMJrrZ51h36Qr2lri9+z3+leFXMs
3j7cUQHWxnQoDPdzToCrUSGXgkBlEWv3fYV/blGM4bN6iC6AiHL2lIbUUBZa7m+jlDiuPqiPTMHo
wA/HD07BZFLUWNPR+G/to1+b15/DhBDdWpEPc85oGOzoYKPjmyrFR2Mcq+pkYpP4uvx/CWp3FjnG
fXP9EjiXxQ/6X7j+4Y0OKXzmwDp6Y/HxRursuD+FOkb8qymxShbu3iid0ji11GfW9lqJ/unQTF7e
Al54CMr8eDdPYmUUfiTYrVRK50AG9ygbfekFj0mAAQeWqB1BFzdXFuTxQa2AUxtj0dhJ1vCFt4SG
+lTOSg0O55QsmBVEkpFFjLYgFiO+9dWx+/G67LNxTjIMEaiBc0bE4FHxap4FXJTHMfasmbPLgnwe
mTYXECGzbtKYcld6xSSYLPnbKpXFcHFPaAG+XR7udE0voF10zBHyMf//flwumIUKUsji5CaNvBEn
2qo/6gLSgxxD07az9VkqsCQNkQKm7HNEj6yE7hO4CZ/1D1i2V7nQ5p5b2MEIQqRWgNk8ktkEZYHq
uu6785s42xdWZREJdiEq+Zz7McuYM9pRkCirOH7JueHMBNBDe6p9Fx9tBU6KVE3VbaoJkhI25Gda
J7QQyKk0eDMyfhg4nwse60uRaBTUj/QAv3XlUkGAp2tc+mayU92uQlpEz6UW3lkdaexk9EqYL8S/
LgSpBTOQrNb78oE3yKMxToHcP7KEVjYp5RfaldOwbp6i5D+kfxXZx3zT+idEUQTmhlDdKD9K2G4O
n8yky1v3UzyXXSoaY44LuJJtmrn1rHDyxPEGpU3kFpKtKewFSC0qpwaYIBJVo/WM2d7DfL7DqhvV
ms/LuDR6CtcWfCjx5W4fsgt07dEUbBBtvudSocqzpyzpWKcFyMpVPZu+dSJgz0cS6+LqjpF9gvjz
szXAwrzRUqhL7XadpGZNn69svG7fiAiC+il/TF6+cwrU50AYBP5RZmN0pQgmuI/LLfSeWtGgqysS
gK+UPyNpeEN9Gpeuiq3RDuObVmuhbCwISomz/7QalzkHTT8ZkMrrIVwUChrawTmp1HXlxaDmNOXs
8dZg+SrfMIRRu2GbYsy8yYIDrSsTmHNMHdkApgsr8lnxFqHe0nDC9iDrwJWJnT+Vekvlp4DUBL5X
OvncbrygCaombhDAg+G0HdMOiR6vWpmgzxIK3D4AJnWoWIveP5XsAYe7zG3VBUfLrH80se8E84Wk
UHpifeppSwKcsmlys9xmGAk16TRf9Ct2NLwp+/aXRWTmXzNtRLTS0cpBDyDohorDPT+NtCxhW3C/
BeOTMiq/UyBTxYCBEcknl/+Ip+MK9k4OPTww7UjQj2n21o+oaTES0fvEGpVv26Wgqteq5s1q7Gib
Xdhz2vIpRBe8U0B6OqfdabchUTdRbbP/irrZoPMRgbGN3HtLGuA502hmvOTZVddoEpv/JaZxJFRU
M6Hrt+BfGHRtmK6hGEY0yNEBEkWct4K6z3/UsCI+cBsH+n2jYKmj/v1qqgTghtet9qlbrDZehrHR
xHoupXsB0yc2pQ0Hey4ZTUxrhCL0HcTuYNuztLDDzPS34rhzdi6yuMdK4namrmcdZUqDhf+J54WX
aa5+6VlK5zdDh/Cv7aglf8indWvwvl6YpAhoXMYy325YcbfDf/HaLmXOrGInW5tfu6Qh3/sgWcPH
YIGw+ly8WgkbhfWLm70JYleOWX8PcgiR6b41BHdbdtJQ4vsmRMeP5ob5EfkpBhMolSDSGdiTh5br
WqKuuvOUyiMP5166FrfHwkq0HnGTn7kUZyWMizmIhum6HhNw7suhbEmkAwuHFfJqUZdeggrR0oIU
0wUl/cakQjYJlimlSvcVt/XgvEwLA0qeQT1reco3+LFDSG1h9v5lKrrfawCNLLVewDH1FZ9+3Lg5
lsEBWCbFLOoytJdPf+cWwRZvyCH5EHPhSTiYc2brbuXcwU/PPupmuHK2xdJyQ0S+eiDMZBm9YqAI
BrOd3UwOK7imDz/L8DkjPM3ymu4bKIzJHlCRg4jIpMV1EFYYXPvU+6O+hUQSzl8BkC6aQxWrPkEy
sRBxdu2/l/UdJvB1OystiR9Id+yNR3l6ADBX6qEu2srQmFIqqvzjrW7uXUoGVLfaAITkTmjufPDy
rxSpubm4mc4ubmKg0Q1gmD87oMJJObHoPNS5YRGzvWWTjoLlrI52eEgj6TiKfB1MCZKHvXMEAQ0v
qvjWnDwvys1fPuBMU3uHAyaBYHxhE1njYN4hzCzq5rWZQ4LdkGFzhx1fqktbgCKBheurX4ChGmom
ogm/4KF//QMGpNNadO0wNlW791q6wo7/Npc4u2LxmVENSv2V7e5gbivo+qTHubM3CmQaUnz54+QN
cHqJUZfSjgIySRKTEEU78qaYHPY8nebqnFByX10kcl83aZYbuuTlfaTnzrhl6OR2vadk7Ck1aTvF
YeBZ3jSjZ9Dt5zg9NFEcgqAH9BurrSJNo+UFV+YkoD38CimEzOB3qj8Ll/BwRGn01VVfzXDEXboA
7+7KqSIrkcDQrHPek0iXwXs4+8eTGJ25QP1+e8YL6fRTO8WSKNiDaTyGghK3xyCntXewMgRprOse
CaON7KNGwPYlRPs/XrPVT2eAMOswRuaaGmIYjMJp0DBVjehOmzjHkSaKNt9NIrY3mHlkDKX4XtYS
3tkoiGvFiU88gbhbhYGEIXtXkzbdwlBLjJKNvSjx6+Fl8qg06r53ZSd87zNe7xS8VQHeFWes1M1z
O2+WvUTBmsEPje3U6Ag2tlt71Ok31Nze84QNFM6oHf9bcKN0l90Wlgy5vWJSj1OgWuZvHb7QOPqF
be4fdNTJFOx/BvCi8pPlZN3KoxuiFSTHF67M/WmHyqEoCJFvpMEQVGwkZTKCV/1Swn9box9qJk6B
oKZQeCum1fKMAVOFWKk+oIRu81ZkFohUADy5JMeI2xjit535GXKrzwYtSqZhNd/rBt/sIPq1Ps5G
z8gGn6QK5W+CGpcPrHN/p6m9edg2GhRWIVOamNFEz0xL6UIeHhxjQq8QO4UeKM2gOhNlieS24nnR
K9lWqZVobDf9RoWON6IB+PBhj032Ksq2NMlv9EdW4qxbs/pelFrVknrefwlfwbQXOKdkBX2r1Bar
0AgJ2BNrG80XTv9+DGgTNbqGZlCkryB63KWojfpog0qwoFtWQfb+bdijuy8A54PUUVbDTeSCCbhm
8oIrJCi6tZGY4JHylzg0gloiOhNTU7vgmZJKhoxzjbYidX6MAGfXjqBoZnlILLnHjQn5caerywkj
JAlpjofFMGtvQjEpC3ja7FwEDi+dswxvfH7zv/g8Az00RwbfBF8eb8KFt11D3LAIXFhZppPGh7EQ
Az0fOeJ5RKdIc+4IOzwKt0Hsmx+sxjJKXEK4C+K9EJfetA7XbSAmKkE/4xNGPyKiMDDFcEmS3FwO
vKeLRNB6F3tCC/5ntemB/Bc2ExA48OAyK+FFOLUNgA3zy0KG10uXDzv4qgiBQH2dLHmWoNVmrLbX
2UUJoT8zmymWcGI7WNM1bFXgnPtrZ5xPI4jfmjF15kD+oZb++qfJ4Yr1kECPEFr4+LB342RJGGZF
ALB36SLs2UtsY212G9BKdIqVkAIwRZh10fZ1GBCUugWA6NcQ82Bn/lNJkbgW4zQx25MHSvMTpsv+
wFGBVBy8RhjoD5pUiYvH/QuRqkYWEATb10gq7AWQaPnWer3tDUoXy999T0Wh0J/Qo5a8WEayxzUB
fPmnKVX5wlmfooxeLjgnxckDTvpxyoVJluiMutfshXLPJp2Dp4Cfoct1ftJXCAGdzxJWacs9uZ7h
iiSwjMB/wgZ5hUqjFohMh/Sa3REC0pr91zRNpPYrGNeKVaYdrRtBFM6tlVZIrUHcN7UKKuMC31wG
nANj6l87ont4n4E9MwAr2rd7VguYMzS5zdIQLu9qQmw4HqFZ66EBdflY/pJvhiJ2a6MzWhD/BfOG
NpZSWMziTcXDxciNt56xn+hPWLJDX5jvjwPmHa1G8Ga+4ZR47AkYlW2N6cAHWeKqRCk7QhxKsR1C
GzDV5CuoX257yEG946P5cJy4MY6cxB4ckazvEgn6R4SEKnfHwpeixjBTycoyRAn9P8KtgZKG+YhG
RqMONLddbH22NBt6O0UBv6SHE9/L9371OgYTrOCTbWd7CM1KAQHwkD46ZYTBUt+uKqWxa68YxU+1
Gjukgi8soMoCWANZtaUKiqOVZiKXxULKt9mQuKn9TfLg2lP1Ho58cdsAJxQw/eel/YM9CthLpg0b
D2O2Ud42hr6wXEPDN+IBwyX4ZvWizQLsl8z0scjqls+2i8WKBALdhPT7ZE7SMmkldldbi2lne3fF
Sv22uBoOC8vGQNSpdFW7yBOagomnRrSIumyqxX05AaGVEtRfFkL7bV5Jvm8jY6rIgilzswXjmZmh
KU+HYvlfbN/vlzoZQFKU+eUmXc623X02Kv4wHQA7yZPs/Dp6lVkZ3ipZcCw1Qy9g3BAcSD0AhOtl
aSw8m8brbfd6pp3R2k256jZelzDulEoiKmMy1wTRwWtn6d/ilxSBN5KSYDsB0MR8dmcfCMnHhR54
f22OtRe9qP4PLEWI4ntTSMKykU+O/ioiv8wnBXdfpQDRkA1NO/PjrmOUvz+D4x1fkAcIJuDb88S5
IhwEgZ23SxXc2X/CnAPRcV1NA3MliHPO7cwvaSgpDqYk437fW/I+l0x29DsXpvt6KLP8BC0fzvBl
3G7PfopwuYiKSO2fJFKbidqucaEd582/2vB6lSlTOd+yjqmCyCfmsvsqJEt/CGrmECwoxV+BsCBz
DX/I4YAmIcG1xothU9n26hugcbGdmFZB6tafkCp3Buf3ALB3MIgNK25gag25qmrLoXzdhN0vQE0x
sDuX+941+vQJ8p7uhDUPiu3h0SaMu0DTUCG576ANyCu3qTq8tnhiD0XqrT7Tk4RCPGoa6EE8uhjK
4YfSNVflhq+q2H8FU2ao68ZUtUkmt+4fnD4mIYawCM+ZsU5wIgFNKxC+iWgoMPIBMBHUfS3lhDjd
SzmWJp490KZaMPbwkz+f1f7TaPkVt4JQYz/CZoEww7SejVT+8WpZ7Y12lum0OSM9DGWXaO5LtHrD
CLHKy0wtHrHvHPhjk8j9MAbsLSKMpGCYuV3nIo52u5OQqFd5cUSM6HKGcCP5G0Ipurfw36VAzd8b
i1lBYNCoMmtPmkKaDeuUQdlBXdMDbWAjZWEJfb5p6YwmtraP+oRgYK+pduGUudeGiSg35aCCUzvs
TXoDhdc/c/JZRRkqpkeQmmocQ6WhdMxMrC2E0cMDqAFpUCu5AVXODaXvJat/Z/GBj3XihWAqMTH6
Lu40ljvQQcURwTIKZzD0JMOItCNYVKwbsvegHdJbPVGFBcplT8hNQM9/yhdLoDewH0BSFhu0isVr
WyVEi51DvGw1HkCcuGOmg5D967IdQ+kwQRhnLC/bwEcu1Y6UAXpdAkE04F25HlagDoSi+iNTTGf3
r+Xx2SCjwurC51ccS9pLIesayJiFUle0Uq2x1R5WlagidSPuPA+wJlFTKq9NDwOr9vDUIHTsp+R2
gsT0l6qlR+q+8nTPjw5u4Xu17VKcnTYDdZg9JfBBBP5Tzby5g+hvdz9DBVd0AL43NCd7GsS1Ncej
gyCd4DUy0whIwDGwHwftLDtf9pXiMnsh+eIFjnyABYR5B4Q1FzY2GPHENkjTUK7ZGMu4nxY0cziU
L1K8kKy1M1HZ8khtai/+xoTzN8DG/ZfRVFyTPtxoXftZaq2/Df7Jh1RJ4pU5NOBN6v01SeLCKQqf
9iNoQkibDJlGgGqJHjDVqJmggAYEFhSCD6L8hTGXkV4uYNnyfqzdwzxOMX9XJoZwJOLgcUutA0fk
HDAu44c2AqnRQSYpV/13kuuQu3OYoseUsFb0jKQ0g14o2CaEzc+omdUNNYYCJd+1K09/1Yy49sG7
HJh2qmL4r21Rb9K6MdwZ/SEI+SHTyl3OeYXK4Vx3Fa5Q7dnRSCyrubthiaK86A0jKO1pn35JeWcQ
/gWgeFvpOi3jYB86TvOsJoOht6F+h5Uet0xbl9CZibb0cGlmnykJnwga6gJ0hsYYDXIPp4JKpqwB
zc/QD9VAwU+Sg+7twu/ayFgfUmImvSi59U2ypvJKuuLAgtYbaJJ0ByJLcGrQhp9D6PTNe2vFT98R
mtiiiZtWRVIGXISctU+RYvrzKHfI9RmLXuYhOPenX0jOa+/nJlQTVC6Rk1Z9h9F7wppdsne5ixsd
YqQTRuC1YD6fF3Qv5X+jDmqjNGoIgJTM0GIr7LYqhh5UDzqOnBW4apUS0INko40ibmE02vwQju3c
jn5S/qfnqKAQsqgWOcNKbReFKRktAt5qHHKWSL3iX2fvhmJwzEJRZ6u2W9BmsLuU5qJIONJlOiEU
JEMxa3bWLEhMezY3J4pumhyN7RYbgBNj4ZqFpaMjJ6euYK9fvQFZHLn3EaSGlOXaghbwcbMQgeux
FLmgXUTlQfBc5937IhOifMojX0x2z8lO64xzL8dGCVZXpPpj92ayBG5XjsJjyHNCS3s8ExDPowUe
I5Z7UCJZppzhKupN8v28l3WQzXxzIjiZ8cWBkz+6nJTnXzN74amOgbEf+CzWD0uebPhMiSdol0cP
bCnqepSE0ayfIo19eJHuS4E76eeWlbvXE4tppoEpZ2q/qUl5bcYobKJCyHujKZkpCmHoKCslDEYr
ouugoOtd/HHeDZZUn3/CFgmJTEWVyor7IwMs+SgURAlFQgVaB27ZeI2F0FxLGLUnGlumEBdoSBaI
7hEi5JFf62hU3smoPOE73Z/FU8AO3Gsh9qUu66tIf41Z8B2jIwoNuzPSOgvlmaEdnHqTFKyLkqD0
hxVOD6fA7DCFOplhB9R55nPKXfUPcuhhKs/WRf/0rcMkzsWYZG4nax20Vvmd1HolmdgJ19dgnm3d
1i3gvxq77zRuE+UvTYtIsmMMl7RG4nLV3SSg1USKAmnQdTwoNm/3VnUpjsPveTloqbFshnrMQoFm
xkf2atkNEdTjagGHLU1NueEq5oJcxjOxd3RTv8srFIOkzt5FDDeywpXDMAA+h1LQyH82OG3M9lyw
t8iPzTsCZLWOhWakB7SvFc5tL34wS50sf6xLHq1BwkOuQTxiuTqjvTNSwWPVrHJmVoAlCJStjOpO
qLDRbsHebwcdk5zdndkWwo6S8A21nyJ1Gw5db3pAdfr87BJE7YYLp3LI9JxAXhRVDh1ePYsiyoiw
IoH3HCTlHMnGVvuaYjxg5P4WmP6AyFgkg1R6yy2rjJy2b1yI3goMsO3yWfzp38eE6pHlJbfGfYss
OEpNoxPo5gw/Ud+gHEf+QBotew763e8J/c5D+yCtPQrs3BhL2BW4x2eVoQ6oMiiUbZOWCF7E62G1
3rB582Q+kSl3sAt6RWZ9/JOMpcOPsqZb2IJgI/S7LOtAd+TN/Fl4k+CEMdUMIwiqtgA8d5POrCD3
Y2U5VtPYEyULbEa/abi5ZwgdSvGRG2bz5BIJ+tFTgLIOOWJalHidmYateBjdLrsMNrlf1GuiVTr8
tmFTBVF7GIpDVYNJxkcTcq3TDWN2b4bmCkPAGqB0QloGXaf4jjz52/vRDm61ncHSUj7BRx2xN5vu
cVF/U32vr4piYToTTkTl8ofXt9YQlUKNpfvsQwJUS6yv0wlPpFps2ooTJC1gKoIyoyAv9BiSwgm9
OynMTANCWoYppkUlO1ihXChjA02YrpBLXPNsUa5zAwKPYfiMjn46Qk4fhrv/91QjedBJr2eDEYHN
iyQ+FyG0VXr/ff+El0/tsCjKZXlFeWykoyZZS/kC8rybO59XwRVDnIrSCEI0SJy54ggsKY/nw/6w
J8uCTlKtIYSIHHI6my7fHogKDxvyH4+ImsTYeYRM/o2DWysjmw2Pw3mPIEZptZvpRzbagkpcs4wd
O1NgNvRAKfecJwDouYrlDyBvW+dDtjD8oPsUNdOAZX0GFETJ3nXp6SzjxOsTxCTYkU6NUTmjQSE8
dVuf0IYPQ3iAPwUWNxQLURribePWP3YlxRB4LaZd/gCba1CLO0xcxGZsei83jM5RwcOiVvH+NuCe
81odJ3U+V23T996kVchbkcH9y80pN4FVix0Y3VW9GiglJr3kCZbgATWFKqoEvGwZTEGUmD6UcY5x
JJZpcj9dNQZU4g0KQLlSd4EkeuksIB8Pa8N/I6dhwdlDDHQTivK1jzr+NERYjdQ0QjwObO5hYM/x
SzVuwdZN68gqnhG6hAXNideajlZNp3dGxOSllP9AetXu2FWu7rLLQ2LheiTcRkBS5A+AhA6OK/qK
CNVnq5RSpwkdyocgZV4bmbDhk/vRuVOos2w8bt8zxSs1dZdjRQ7Fu5cqwJdti8kaj8jAP/mpsHul
fYXpO1P/WHDqDKzVt0OKhQYgBqwFjsKxIun5wlGJFnbptcuV4FTMIID1IQd0BxOcYsH1pfpymZuv
Ue7GIKNjxruzw2yjlistr1xx2rqEOQZkNN9gn3OTY63wOjNpXSAlScwPFjIUg6vlD2QuvMyhjsk1
Hko0IuKeZ7Z5bUSyN9OmZ0gwQ+dznf0k+/LGHHzfUpQDPibTHsWOpWP2zDf4lQDFNNxQcdx47HbX
5iRyTHngn+cMeoD7kpjoY/7eDfmKZoiEWd453vMXaIkMb1wOrI1rxTdJdXn8H1TvgeXGahiZMvq3
uIkHmu12QP1JS8oGxq1y3rowu1gegvJgDsfIGXyr3YSs4VQY2hWu5u/hbX3YBSGsSkiSbRyeK3NQ
6DPNPqiR3jymqwoMshxLsq2d3taFJBQl4XDlczqPBGQeInkS1b/caCw6nyQLhUEHG8uiYs+BFBjL
hl7oEezu+BHxSOjhYYHFRjstAAHW108FLSdkRlBymnlde4MOgWC8bb3cWdaW/PIScig1ajPieUXC
Zo3zs4j+Nqi1ZRiJuvcE+WQjGgwyySMFCPRHDoCZBUarK6s1wl2N5JvQ+HpaA8o5QI69a/tp9frc
kQKIFwnQDZhzmTj2E9ANKvxRVyKpClBIpCdYrKPFnTAAWnec4jLikJ2del81oRxoPovMiCKerPDG
0XYTIZYM9yWcErzd0wnsMHZHbSLBHjhXReekjaHy1W41VrWqV57abF6zrJb64GzahV9I8HvbjpCr
BQOmW0U/Jvk8Mkvt2dR1lE4nkl+fvCvpgn9s6c8SDsgoZWPZTOgRdc4LZXr++NKYQPObO9vTXxCu
YhwU/5+ZzyUqe+ru6pEMcPDnpAzTtQ0o8Fxl4xia6HU68yQQz06lVDJ3Bj1FPviAr2Y6c+Vmxf5Q
C/Vwbv/T/qhA54FbrfatDFQcb4ySoopmopHlIno4KrIZEJic6IboJaB01n3wZmFVtUUMrx8U26jC
guN+UW3zTH4NbtQJ18CJ1hNYP4BH4YL5bdtHEpu5idDMlRUciEOPzhPPUr2FZ7N/dO7V0gBg4DKs
WoLQI0xi+p8gFHr84pHBPr1kIwi4GragjhhvpLkN+/FzsDxZcou/gx77mFmXsb4FmqTZ4ZSzUwW1
4QFWL60glY84O7eJgqUgwSq5nOXYSX6cWLBh7FOykGALCFoDyShpM2YIcZ68NaSZHfbmUywk8Enu
wWMS63XNxWufPHxdeUOLyfGisTSLD0AGIvgYz+raupmO3FODAkrKztlH6f4tFiVdn4R/MSg/Z46d
4AEC7XU7V0vk6/SohRWn4r/IvlnaslvQlY9cIhD6iudwjPTCxM3UzYQ2RCH7ng58X+e8c1UKBDJa
RB9iLvj/4KAPvDy/rcf7WpmU1jTeIyYextHaWfm3m75/+jYlwGKk1YUaBzD0BqjiPKtWe2XdJorN
dxJSwcM8wQENxpSlhHNjuGKVeiokc65w+KeS0AMKKonc8Nz+aVhLPnKIeY9/UblymuT74wyK5Ut8
2kK21hKS0XLHer5c76qDjzhCCNveMu28PP5DFRx/CSpK2npE76jTzVTvv9S6BRrxXfZD8o+XMuJa
wCcz2rBQkfF6+vUOEIRRbXjjqDSDk5izEBkf0wqUDW5A3+xIDGK8upBHF99+hn4QJX9sayWTb61G
fUkW9OOxiFgYcKr2RoC+xBggmfpZTwsj/DH1skAf0Bugb1XhmEbMbNeq6WX2Ij718CUZfB8hYCYe
4tG3i2f+gL/im2/d4VjiONpDhd+XVpfq3r0XpiQIrzJUqIHO7XSQMUKypSdBo1ICwjAF55iSCwO2
XO7wTwc/S2Lz1OKImWz8SFsUKe1ar2/nDSSmNgaw6mlTBE98Ybvd1WQ8BjHRdb8Gsa4TLtgZb5sz
PONcN27hw7dQO75Z6aQzm84imZuRskLfQLrmpPRSH3GIFucaDN8LTn2V/WVUeBU8vyBivWPlUrzs
Ci39tMAWXKCZ17L98P9BsIdz4RRsNtDPNhqab21RzhryBfR+f1KrtWKwUN7h29MmHFA5+QU64gXl
SQ/TTtpxOUHeuTGPSubl4XYOiBD0QdBf5ED/Au/kicxLFUE/k6/4lzTK5zLmp2/kPdrd/Oq++4dh
TnPvj0youg1q17a7RuWc/RWDRaEAXB32sg8fPkiO/t+yqi+cwDL2PtrZ/8JuTzq+ZGHM7hBgMi5Q
AO1UBrTzB+Qfotc5sqE53tzWgk8H97FWW8dCU9MqvNfxhDtwryXJxn9p8PfvQeM58vni7xdTvzx8
1oSACpOoqavkfcm6OpMSemB/qkPiiRjd2OcMaAx68XJTSRBybROnOx9A/LDPOw4AiCJ08L+1r1/H
u+7OaNv0uACuUu/yhlY6tEuDAZX+wn3BSk1VhjcE4rHLtuR8rOeG8KaJTDC4KQ3fJF6stMYodzq4
wonKksh8oiyVeAVa1cDamLhhjhS45kWqe6H2ZqtdfJH4JzkvpXaVZnBXhKpWvb+k2beEs/Cj+q3+
cET/AfMljKfCk2F2frVyjj86aQ6+WcwXPUUx2t3B1Pp1UYXbcNc0H+faEvSYg+e4lpNz+WGl1Pyo
V5iJacZp7vDCXW6pWFhgI4TXrqlfbz0uLXbsUzTiC56GVjMG9+FJHQbZxdwrY7bY9WR3BvfJSdwE
hVS5tKtozaew3MUL2/1vedvTVZSFa0x15tocmpPUISXDNe4tAeI3Dtx2TH290APq6de/KCpJmHX2
dABGIMX5ULA10ZxsKFrh7FF10fjNlmLMB8WZqmzm+EYPkK+TKeFy5Uzx319zfPeTjF1h31uit7KK
zuJ8dlPM3me7wrBB6UW9YuHSGiDfVk4w3x5MObOlE0jaYGCScZheXd4C3zvN8t4kgW6CAaYozEJL
Kt3jCRF7ML94zuJpF7NpcMr9o0q2THnLdS92vlLtyHiymwnfOLXPiRn8gkV2X8cJXE01npfy38td
6X4P7KoZDdV9ayTP8i83A18lrtYFlg03Wl4mstM1gNeb8pecs3j06mCPPc+df88h4Bi34RwihDji
zb6g9yWPurEvM6FIpqc5udfnINPzkqk3Ks9XelH6nAPi+SB6+rSDt0QcBfPmjEqcXy+t0LEWBRB0
YYf6pJQQnl6rvmWldBgcyF9u2MrjIr9xiz+x5T2uuwurQCcIZTMuoE6ij+3Ialj3GLo4afoxgfrJ
EK6L+z+MA0Q5jSJzmMYUEOBKAZ0GnouwzwaBnQNyTsOAjePTCZfy8oRuvcx1PVafm7wg2JghavlW
CvaRT8eAsrDroRICTd9PXpGafZZqQiU0iUE5KXlb8UzzLzpE7ACmr8axohwfMgFCp8VV7M2h63HO
tcaCyj+M0f0jajDW++PU6BxWm+teZ0nr1pO7xhIgFQysUuhR9qEL1fHTXX/9B5IeIDeEhvHGqJVf
4x+yVZghI9EYRxANUHccPS/qWQIMQPiL4r3bae2MGj6cU9Z9qAPZlWPsBq5pzkrCbo5BPXveyo7Y
KGclgIqMwMPt+U4g6Wof8GbJJP0dUNAZKQKZweu1LGgbEEqr/m1wOf4FGdg5fhpl8dugVxVNh2PM
khKWNHna/wh58/VwesOawCRx+FyWXmIlud18/nGNzBLxRfIYhipjfX2oUD4EzwmE1s/C9IVT+URy
PYtzbLl6BYw9s7XNpmNUXP3xPXP0KhbzS8Yk3sUB7QgGdTaIlrmDeQfuap5MWGqs1DOlLVD8nt0N
LiFpWkWitcAoEtkTkcLeKmObFcz/1HGpiaemKSVFbhtUbDVSv5OYeLIPFGzGYnJyIwV7yH9kcpd7
EV4mImnTsRjHHCrmpAA70IAgVEcpiFtepmketvmO3qLwDxH84DqtJ6pXkGUwJfUXL6LiO8Hjlm9h
NHWqvQPrmmE/LbfvuizbutQYMsOdMrL91cU5C/z7JsOstGwORdiVLwmeL8AKXpWcJGJ7LPyDEtLU
hjjDSxa22Cul0ub+uc+MJgJQ3ppgLdufVxQ0K+6xUgSF1gqMnhCgpPPk+LDOFv8++C4Xx9gD3AyP
HYBNCgAfm6MLT4Xe/5VYZRGmIvsCXBONS9IPcZ0v7VPYGgpI5998c76V1hMI/QhD28THBAlTXBW6
0OdIvsvLIYHhvPmXdX7t0+cygtZ2MG4vvBYVKRgZvi9wcdym3pogH2DMqdYeiVyT2AQ5wS8lyz/0
6VdpcYZMwW2Ixo3Bhi2cve/3saLOXYxLPdDj4DRX/ZuqHDgBGC+o3LWd7DDaGHcHjtlGY5rg/zxQ
xMmZvc7qziwnl1JNFaIBEyzFRGmuj77MdITKj8EqIqg3kRygElb+bOrD11sX/jpsUJVeC5LT3Lus
HWvl2LVND5zCHeY/KRTvZ5Br5Hx8JIZkEyMgJsUCenZWtJ4IjvJiLG+WeywDx/Nz5osSYQREtg1m
p4clwCXQ+81to2In5W63K7KHmGD9o3WdGDibW7gABfJVyCxNeqdjKfcjk1vpB1ddzGPpGxLlZfce
WhfMkAwBcxPZIk8TNiSh9ZXP9oOY3CMRBfcy/aeQLqwd9xQHz9lfCOtFdNGBIR7MmGWDWut6akuJ
6cG/Od6uEBdqRGUYiZt45Dyoz5WKn37WNh6C+ZNBlAteBDWsiZxFepcu0iJWO/DCVDucqc+QuneZ
0IP6ugKJqdChohrsgd/RbO+IWrYGIFfPEO+yGt4OpLed/GwDWwx7DKyPD/71heXYYHBexyTTDx0N
U5TjhQJMfK765kpErx4ntZ2gIhT5DR8w0r7soppieDORZtK8GuV/8inLy2pzhGgC1vxFKsFdIAHf
Z/UZyihhjzNqVg6OwucjZbRw+q2i5rAAuH69KSwjAka8nEMFEWcnY5NwF/JmnhH0x0hvhFaC/OCj
zpa8U00VB/uSatzQMfIH/Bstp8eBbr7etvG2PQL8JauOJZ9EiUXBmYdS6AeWmEfV4FJJSUTv1sps
qcaihpd2wH7Sfk8fB1mMdquETyxQi0o+iDCcgW2csJlqWGw6dntTJ4KEG9SmEUkqpTM/fm8s7dTu
IvMxXDzAWzzahZqkYCh9zVdKBhZR9OSLP2IJ6UHbfq3kSzv47Ysa//NnVca27hj6ntRkyCpzd02q
9yHbD83I4xI69IKdYDw1uxgVoPbUYlpOBxwPBFcXxFXmwNI5dWjR/XHdmDA1z+y2Y1h7zeRCt+NW
YJ4l/HgeCpKhJzuUn5h9vAlrvzb/WDVliDyeVaIa7MQkqb0tgRshIBOkf6pLBh0SmtHQ9MLRvfoR
q1JBauQBuM6tpb2AD/r8s8NzW+ySgerGjNGbPsovRNfDzNmb9ZltV3JLi1Gw1oa19ggUmd9SQ3k3
+A3z42njwUMynnoIgkIFqMSBrmaHX6+z1NdenwpItJIUhYZFscmheJ7WwXSymNLObJ+RAlBRwqpA
UZ6MEXlXkopQ71wFO9pZmzN1QFYLmmIJJZXCj0L24y2Pm8lAGb2FagpRA6RwQYTV4kBWmIFTy3uz
Yw1g1yQt+oOO09zIBzFBK3bAYcGGvFtX6Tz2QIvf5jARRTsNcv+ZOmkbroU2u3X2wPh89TOi+bOq
gRPjV+zKjprZiXQ96o3pn5EowAgl48lI3VId2FOsHTZphVDu/Ic42RitW2/rKjnhMcyWJ+IZr/AR
smzmN4aEp0o+gZyLwvt3hZJQfKcbAmwc1z7uU/mNrZbZHGRbUTXqHrk/8jeD0zozfpwlzfiV3oNF
5XCzlHXPH+yAOK8xB5nz1iVDZH7zqE5f+aXy3DJAJIQgzYXrcT03HzfGH9PL6gLGeJI4UyNobd5t
eRaJDyn6m2yziKDvWaWyKm9L+Z8no2z4EmF0ivqMkWGRF6Y5ex4NdjFSS2AqK6WTxWLwRA1J2lIl
SqGXrPGjP8Jt6uJF352xZG4rn4k1T6ShYQ5xpg7ICJlzy8UPW7hFuVCPdG9UPv8IAZ0GUDqoA/6C
3BXOsBwP1Ouy5pGldpeBKxn3PcyolBSYT6V5+2luBs70KSOcGvT5AqLSmE9c5dCm2LUHXwP2/e9B
oJfLZUbfYhwjTwPGgFcARsu6hhaALEbs1b7hjkGNA6J+WUQCEzR39bJjCzbbg3RJo3ndsAceR9XR
IZKq/iyfcqDUoFvvZ8wwjuTgM4MdaLizcRvUMyh/J0BZKVUa8A9j4UMAVGTFKmPoaFoctxUywrSi
bU7Rs6o+RIBTYISVThw5Ymri+Z40gyMUj3d1C5e6oPK7gKQLm78Sn3YdCVTa1pLnqwscIF4GvIaQ
cCrhn5tgRRQF3EsRx8NviZvblgIM+Ly9zEWZrwoUXjBZ4OHuF1iL3CMuSbZ1ub91/hTKA7y8PXy3
QSiXP5tdOg/iqhQiw+z1Lda1tILhLofGxPeduQ4W67aqEyUrFT39hXHjjoOK+y54+mrvbdDcXgbB
v3DsWaBkgy+uZdh9pxzrZtGuVcZL+zksNl7StaiThSl9MffKobf52b6F07FmGQn/9XEKbQjlSJPa
+QPVDx/S4qoJg9fwsMTTaOuwYjAD0SZB0+qu6JhJPgtLU0VelIzMJ7AfrLf8twlbc4ceMC+JETgF
j9nP7GoD2e+hktzGIriK/o9ND1hEIcanFlYnI6Ux2DHNkRVVAiA9x76mm4EN++ulTTksA9uHbLJR
i431IkwEOmxuyyfHCaLhcSDXCIVkuAhnyEjNXSxZT0AgFUmZBA1nfmXGr6a/kCCtVC9zzdNwpcsp
j3C6hBmHC3c0w20/QtdoeGTs+wq/QJ1AjB9e9y9AnDMQPHIGRoEdDx+b1vA1eG6z6F9gXP1KdfDI
Cry2JLSdUlN8UL/AxgHBc7MoHMNeXrTtxfyZLcTZI8V2wEUvbRNTU4yTD3/9jnv2Zy9kKrmMBO3r
6RXTrCfcfqjr3MdtC1qUCqG5MuZeDuXluHCO1LOT0KPNEm5xkR0IYbXjTJ/xAPi+rAa6nVHyFaWM
Mgu6s+O6AAXJz5GZHavTebFfNycGoDfM3xq0y73BS84ZIuFJPtKmKyxKy7zF7tsYJMH3HYXq30r+
oDMWeO2nm112xIf9y8HANV+qouFjMnaB/cwJdx6/ON+IbjpAQ9LGOqMbdvUHT9mDb/HeUwPtr6VM
jw/WxD7I4kuzcXCfMuk+kf50TKaV8+dFYvvNyXND06qc7w/TmKhOMzTChXKq1NhbGuL8Cljpbe5y
BKY3cfZUWnt6kITMbVj1WloJjCaesN9BDdMxLKXJ8TfgCwrLZOP0NPd9P9YPJMo6EUMgFJMOdnFV
0VOm3ge0Mkmg9VHBeVJiwOTgX+CvlasiATXq+Lmy1cadZ9rXogJZ9JHrhUciFTPAk6JzWpTL9wSZ
v3W+/+c/1UnuCroYMhD8CyISr8bQEUC2qT67g5rotlYAgLqBE/lb+4YHA1LnpoOBLSeTBxYva+Ft
xj9g7ISQ+/8VRXDqnNvZsVYVC1tHjZdpG3kroqDnZLwfEJt93i1f6kuCKY9D2v4YmVbiiPEDUFZK
VnEnHpKjxGsgNx1R01rB+aPb50wH9fo9gOXVfMb4HdWvgWGN7OAEcoo1hZfAf4I3261RI7R2NGcQ
T9kLXbT2iHxAcxJznbaejEmrLFXGZJBXVKvfhfOtaL+BdZVHoSc6gO8nYzH+7zs8RWLpnycBpc9t
bYaidBsBFLXKBTwy7xAoLxXUw2f4rcccau/Y5ddunRfIcoFD430gZc42l7b/k7g5hURvFZtVZ3n4
DfRQ8MFW/pQkaiXlRo8DZsoGzRiukv1pfudaK3xDAMBZ02eb1kN4RwqeF4N5/GfQ+EibgwA5lK9H
tY04dgAM6A9OYo+v3+rQBfEqcGw8H3l24tLb7DSBrO7ikb7QV/06GED6UrCKGKfq609rd1ZcLjQE
OVCaVAUg5amLFiSyJ8bO8VsBl+ZEFRLS1fFhPGLoDk70AqwoTjoTz9CAnfqhNDB/1b/2rOdjfxL5
r1dvmXUi4l688QTv07XAPKaXgMxHIapuiJrihRrZ9ly/0LzakbaWsW5eyD3uPTts3p1TZIySxCJ/
wqUrjcEBDJiyQkX8wkb6h4TG042yY09NTWU3e7qhsLQunGS2tuU1naGIjo1WJmdpN21SMakaiygU
uixLd4D3ZRsGlV/JO8gCTSgrpzz34+m1oh3/I6yx9f3X0nqKbc8HbCTyNJ0QP8Lbg2Q2fGaH978d
5G6pLhKBmSSCD+k8BGuAL024O4kyV/O/tkczZsNJV5fg124BPouBgSW49oCsf6PpePBtVDmvdXp/
8J0xBN7w6mpdBhq07Dg5oh/xBuucTIuyHUcOhTSqU4EgOT6KjFTtKmhwe9d59j0TXAJyzCcQwQdE
l1V3qQHMHh4TPK6ZqWmvhQNtu41axb5sxkrUTY0+hRfVgZqVXbPANAc2jkG6jXH1m6N4bQnE8IDp
rBl64p0PlgmWFeuO6jBv23Dyf+Hb42fqPnjpc89hdbETOhpf9+XLJ2sZxgcz8RKPuvJU4EWQzfnY
D7KSLpIzxTDzSZRNe9MegKRtqwUrA/AQdF3PeU59u/brcm8r+9AJQ2nbB+4wvb69truicsNUWqti
w1AFqSslRgA+zGXbNPh5UM0kVWFWGO/8cELunoWeprNmTMpDk2JgxQCq/v6Z/xSqvkjeq52XLkR4
HbOixXh9gOXQvFvmiC4iH6TZqpPhKZBIJHvHra7PQXw1sSl7h0RSHXxlVwvbRSiP/8EINSiwOWVJ
EFccxhyQUAvva1SMV0Tmm8E30qTlx8fHM0fl6gPdAnum67SCUz1GKvvmJEra1qnSrToPyrSICIL9
b7VtyfFBqqa+XDtbYCnM3/+TztyJxrEnOj6lXHLf6DQVmKcbKcyGx3xx3nTqq3mvbC39UvEF1TLX
oHU8fJHbiasfMM9bif3ryPBAqbAwsDO2ewhaL/IClQXRzxtq53hVkGuSI2y2qcn+JrLH5N5s/Eby
tR/JcHUf/eX2El/038cV5BIYmsYqtmXCvUFySu2Q+OqaOYbreCOsgWfIYGX6dk7GyyF1ortf3ucw
7rZICAhG1ywhuh308JbcKpqbKqkAKvZYe9ZGLMDhqGv3rQxsiRmXIsKjrioWwuZUnpSNmQTEVB6h
3hpWFJAu4Z4rdzQvnigxwaswevcKznl8t3NlC29b2RjCZxyihkDwZz4mCrrhrSuG/YagwN9l2W2H
ihyKG2JB+58JoG2zG9ihlaFrjSAm0R9N8FsShsbSj1KrLmP2Ue/HaHSbFt7QHY8ywjb/u/lhlB7X
yCET68RVkNMmg/Thtfw7JylojNqZXnZCFBxD3ReBTHaZzuWZJvVyGgXXTzgu+Q3jGPy1vLWGjxU1
xVzYgdsO81rsZS8/owv28I2yvZCEM5/xB27Pr2ODvfGLLEWnk/OwZ1Uit6y+puhtOqK9oZx616h+
1fUSX8LTLpCFa0osgwPz2up4yOXl2RS4uCLi6tPPYC9lViYiRhWFxpqPfU1Esxj+ekQJOpK9rdvr
BKu5Zw56SXvfyUqK5SRKK3wpRg/hCcDDMVkKO/wXGpDFOSxN6mBOQTn+cfO9S4MahyMUxcFO7BaT
3bYC7wTS3yJpKSrKBnzJm3JNcp0VPpuzEE+S3wMGRHUrGQ6gJcm/h2N9B5qlwouZVKQZhJf4r9T4
oL4K7n6ZvxgEg2ETthcWwovbaFe4CPZljwvrbvjzQFgef4qIlAP0Fmr//U96LwGhkMIqHG1USq5L
R1+pk5YcxIXoeRjRo4XDoe91We6OOU3BZfKMuV8+SJNkb5Qo3gcjy/OmEdnVmz9ZFMMQXHFKqETY
+FaZdMevExhPTPRAldxh1VOD1uxSZw+/q3JxAvPcvWHJcRC9z+CITv7kyq+w/t8yWORy+dwiDRkK
qT9ztP/ZwxkbUofK6f+wMJlSHNTEQJHTOVXwnxjIDlRiH2ddUbeZtG3ZSNNlyYvzbkLFugEvMcjW
/IcG+J4/Pow3CM1rJ7Kji0oxhwIPFu/NACu7wEhXymKP8ledmfU7INMTDq8uLsvDlf+LPMBqQgR1
TSPLSX5AbKbIVCnwflhoIp969MsCzWyUDdB5ZTdzWqPgECmACXgzyTNT2AE1Ynzek8mJTlIIw366
F/NZDsg+xZAnEbmSJtP0lg3XvF5jtuLVHjIKI5Qa1mk8x+kr0VOSblHjFHLVMOrxwHHAMZfVIm19
iSrX8Ze3I0pcEjgZN+CIBYnQqp1mtwYMlXue6mAHsykRHQSBz0i3yvnYdjPQFU0mgZi1WQJu8GG1
5eZKnpo8wI+sRKbTOh4wCe1oLt1kIx3M9R0UZjPqcYV060PoktoU5VfR+mEUGjOLdHqvEIciDg8t
6HY0jjkpGiW+hH9ac9CAlIsQ7x9FTrY8yGaPJw90XMGqniggjsGSG79lhRfLAhHIF+rZu0obvXMw
1AYf3JztugWGoJtx7vsQTVusa2JzhYhj3RgcsImdm5nFK5YxjkN1MDBfyEhKWZ2XfCe5cwAJpA48
wzEoKA1nT4g84HBopk4756Jar5jTYFTmtOuZBWleCTaj+WPENRJX3KH9+HNIBYtDedIYNlf1xYhu
WMl4kzyRajThMc+fbZryWQxB8WQX6n9YlKluoaLihKXjyVVNfuT01+5y1HagCdramOof3vUxORnd
g2Y4bovCwBcus0xVLrNMz53+OsH2ZoObFoDpF5HSzl/vDmO3MHkD0ZbEqI9dsI1drsFEeQtkpptG
VQ1KBGzGQo8k0uWavuHuvptiSLWnFGv15yHoctxz/Qz53vpOgR+TUwIAL0Bb2k9zsA4ra0g81kVJ
cYN9ov5f/9c7kby320j3yxv9kGyswUw7nsl8nlqsFFs6Rew+oxaKcSMD4Pg4FeCq5404DpRBJylk
ivMWx/puC6M9teKqlpMYXO9bN9Wg9QGQpko6H/UbPG1lB0vNcAq5D/D3MaJxA9a0xcepYiWtFUrs
FuUrv3ujAeyI6URrcjTDitvo1amWtLFOBcNglnZIUDqxAvA3kVO3oipctOHaLa7aaBF3ekk/D72W
jXJw4fuLQDx2gziMuhKEmpKpcbuHzr3PWfOTrJ7nEEw4y8UQ0sk3TJkuScmANvnxMiH4FnxuCLbh
94mfYNaBCB9kzoZ7D2y+QC9J5SlUKQJqOmHzpv2EygFj2ey9n3wcuGFTQ+TqphRmduDh0LHSTBiY
Xmt1wHKGKa5Ia5pchdt2fOXm0URgBROR4cni9Mg0d+K8pKw67ajavRg3pHeZll/MLvHzq0COtTXQ
1zAiViA8Fq6TOi1ivXnwitaVULunm/qEl5siiuBJb6mHSPLecnHvAG5DNhqcQ1Lhkk+6o8JE/Nob
3DAhI3hJjmBtfHINL3lU+LHYunQ2GnIkZUGMn8nXE6apgo1mrJnQXk3/MBoBr/DHeV0YKz70b1nH
MFE0JDxTRltZLlKNzq2ZSiCqJK+800h0E75FD9nyp7RhsqPAMrQa07/XNmllmu8HzrtJC3LMwSdh
ItcowyugduQ65ZrreA7TedXy2fArJXf9IBIpj+hOQvdEpOoLPMbkwHH0AgNIt4ukx8Rmi4Gyk/yf
KGppeyb3Gh71RKq3mjnQ9+IVTDmaLskfwHf+gq8gXvnezwsvLwskRELCsTbshTLAQsl3LTRd5sln
+p0d9aIOXI0C5KSMcWnVjHbLOSN4WxthllZdfSjCvKpRv4v02lysMdB5q2GmVcdpoM1sYbxD6Hm/
lQebnfmcbZgUCu+CCatigRguQIPZTgdhFCv7UyAicfH3nYBe7khNfDKJFro5ii967jd+BvHUqlhC
b1mGQJmXEVXPsyUEt5GO1qPxBDPCzXTdo3MBt8xLZuKLXaA9tHLymTExLqwDpLNXVu+FP+L3LARS
nsyI1oBnIekIPAel4nGEdmb077+M9FDWIe7zRS+I/VQ7OdR8AyhM4mE6DqSn8maawMWpD3xbpCgr
BZnSAfeGOubCWN0ZUMtohWZuDshTMLO6gzwxJMTif+61+gK/dFuRwzA2uGtIjKlNBHMPCRO/7S/R
VqyQfDTzBikeBH9ANlLJlDi3az6KfDdGho38szjbnfMYKiqmV4cH6eabiF75M9Zp8v0SpGh+CQoI
BUFvI4z924no0CdSWGC7z7FIqPJu85v2HfUEU1sZDee4IfeiIY7CDTRzM1P+Luc71gktSxqKWHoj
Ti1zt98Z1uq3aazs5DuaRswoTV2clKYekz7/BQHFQOyU3NQD7zAThDou25oyMANTYnuzgt4WsKxc
W5uW5B4VyNbDHJ7skkFd038Q387pxacfwBIgg915X4uvmo1w9+6xmmMrky+OmUvRD7DzxiHCGXml
e2S+OJOuqytswCOXSOWiu5uVgEsQZ/G7bETaSOQCOtb8KDRXvtjHoOW7DH7TI88suV+j13SeSr9e
oqO/dHOjPUpFhaP7R/dKIbYU1IHTiIxisoxjgjWxsQMbIyYohoEycqZzJYUeB/ZDmuLOlbD5r00O
eW3nld7MJ/Ivgywn8URQysc9EnA+LlXblfBREODBxHSyXSnCeLi+VfyZhMa8lfoxLoTjY0Tp5S1C
T8HGg0GU8FaVtdfv3Ju72DPsUDTz/s+HY3QAI9f+6Wykc9T/JT4+IW9+LpmfXfXul2PlYYK7ztQC
o/MuKmUbpN5AJYSQQ/9qOgvKmukBL39UoG+HWxi8lawofrrNqJk0nLw/FEwJbv4dEN0fXDNIZh2Q
gtrbJjtf4x99Oa4XOv5JCMO9kwGoGIgS+UoO+ZxMMAtWmQa/8lIdXGu9qW0zmiVRYawnezaSIO4x
a36q7rh4cwD5ExJaO+3NRB1LwQiivTBKKul96SUE2ZdDAryeA5YOVMXVpIQLLqTjXiMn1m2nre30
xx9Xa9FB2VcJwM524U2NfIeWx2CyydxhZXZKk/1to2ftQwSenzpUTAB1TFjsSGP/elCrqjRH/3yt
g+/mxiwpiit2+kz2+TERGalm/jPVCseaW7mqo14HbxMzgLHICDy8ifdwIbxDkxgucdq5+ZyLIbr8
OVRKmbhIZc18WF0XlfMRCm8RWbSvpwAxmxOwKf0M6RMVvKvHNV1TWyyStPuXSVIGAm0+VAqYKPyg
KrpP+n0tweAY11MOyLubq+TTyNrlL0F42dAT2k6pVb0rtKOoAUybH2lfpGCJcrzgPwSnlVLnS7PD
oXmiaEhmWkJFwEpkiXfhOd6LZ4vnBno1/XAha0JWBjAItcENPLe3E94OIXE/KzjuJRtGo1TKNhv4
1dhSQfnPyFGbls5FX8DB7SmYZI1ABLb806q4sJ1ckfqBNAsf5UGyf64XRN3ytOyEKTGwPSsxW8sn
WsS5QsNPd4Kthq272/Sa2nfwWYyylg6BNeNi+jj6ZmK+4lqmU0exBs47rVaVDM2SF2cn93TWYvCw
v+XX13MVjsrO5tDYNBxzH8PxK9KBhSjGCifwpuRiNzY/AgzvmKplu4mvdKzcpkKg/WZhGFGM4ViP
+wSXh+5u4BpcwHEWwNtGQlSr9aY/eQ80zWZTY4BHlonWFPXxikBvfjpfD03DqrapUG5tq6jl4w4Q
WmeRWapP//ChC2Me0AgZcfxLvyYXKjKPMA1IFd4oT0aKqP0r7jETk/O1EXPPNXmVUGop4qNqN85i
scadhwT1VEKala4lgh8msG0W5wpfarGyHivDrfQzxDympVLVi+vYN9vnQc8LAdvHiiwQ16EeQtmC
j8cA/KOTS1EEXO/JuNWVVCSes8eK6D/fI1eFOoKVsGoKB1QnzqlBmu7g8Iwo3VYxALZSgjjU3DWf
Z2NVqOIpO6MuEV1mpCsgDXZR2KJUNFUdYFWXizyL13t2iw7o4liBPTsf6s/jK+UaNYAzyeP9P0CA
xGjhjUOtLUiGGbE4d1Eh4GarWnsoiemM9FDVbJ9CEfyXVRS+ydYDJwIad/MCM0pXEzNwIh1MxSTo
4zpr0S00ITr2AU8uEOdpvjLBfZzEPf5PjClorpPm5jVcHg/4OqlVwq/AdvTYC57p8CQy5Hc4z12X
5V+NwAgcob+AGe+T7TXz3RMOlmf/mz36k+4PczZRLOubVKHLtlGP1m6TNzGFhIZTmNYghiLPZK4Y
FrSqQy5w9umUYB4qEhCTAN8hwV87ULat64fEv9ZrLSJ/6PaADnir/9s2gKFtwS4D3z9Pm3jI5Nlu
cmdLKhWk93KT9N469awiXLjTf8nw1u6Tm/x4+E0QRDXFskBTQQanBtH74L1KfD5lVIRekJZPhM13
CbgRGzgY9AWSU3vQ+RYwRSRuTQN4V7x1I6uJdRKU9SOTdMboif/SXC++SPe8fP7fhIgH0mQyreXH
kVen0zcoO9nw42ZnAEYu7NffH4jju0nbmXMwDaYmZlMlu1GvoAuFEf72ABfKJR3/zW6DO1TWSV/Z
/qXHq8rxd0sPQFbU+vAK/BwUDlDFe2wlM40lhG/12Ha/TFchY3mIi4ExN+btkAfOWUhq/MP5+5Sa
6aXIo/Xoc+7s62MFBOPrzsLKGjtyByryuEazjm5DqDgbhNPvS91aLyu4j5KWZqRhxeJRfrye/ZV8
phbwhEg1Kd8KThpciP98RSyyCx5lEBKGPSAuRPjxy2o88p0i5zJuGkFnbaiOdcKF3S7vPwXoUFON
UwA74uIj9Rr22K1B5LbNoQd1WIvmSVuSi2x5bl9MSPn86dcGoH6irqQbAcCJUMhPTUvlSD62ttKl
pCyChcLYexgJZEkl49QSZ5O/G3JsvYxt/TTZCfm5rsFv0KW0S2F+ghYq8DN4jkbJZW8GC4+zj3z4
wbQng2teqKGNt7ZhTPcz3s2LfJn24PAfATkHpvTmDPz9JFmKdgQ4RKO6uI7Th2eFcqrYGxH+JXTY
4m78Hk5C1Zl1J5Wt7F8m6bhe2vyLdDjb03r+TPa10omQDkGsuLH8uVGvk+6B/QHMFx0Gl945HEbv
Gv0QOvsMCC8iYWxgrcBFSU9Ij9CLmpsjdRE8wFxe537qfTDnZSnLe8tew+/gdNN+76N1hmd0U5Um
5kJe8ak8IDECBjTsb+9dPWE3a6B3a+EuaUvFrGNB9U0M2BXV6qb885GK7Tel4JsZEsenfHTWQsYW
k8N3lkL+pSw6BF7VnHFl4/SUVkBmDYbvhvHnV5hvpKnJgruGkhu5eSsS1cW+j8r6Ph7qHZAJD85Y
4Zk/IInQhAjHfJPLv282ao0gP0wjmOSYKsDrdhEHlOnACVXbrSnHLL265ZPpGfjdk502930259Pr
+IKskbvwbBf8oqlFZK+tsFbFkWw1teVIGLjqMeFAqMqvQKf2aFLO1K4LzL/dsPQ4V30376gebmsq
I/PV4h7nLjevJCqc7VlD8H4to0cPs4xtCIYNaVbaHW/y2UxROOUY9WzagdyGUUHc3DSWhR72JUl2
v1fL239uf9fWoT/UeJxiIxknjWtn1DnWCsB/GxISYsWVhK9Z2Ql2zCOG4EDeMsQFM39/Tr7oe9n9
Qp3Gw30aYGYQO3PJPW5QbRU9Pgc3RGgHevpyS2HNanRywaT7tHpMPmPdqI4umijvzrn+YSEFkzL5
kY6O0HcbwnBlU51Is3aXZqbIvofxlLdE4Dymk3GEEHu1LYJItS/s12uM+gSHMA5lYOychf+TySwa
DXEQJUnckWJQ3gCXNmz0N0434EuDXJtpVrCNW+9CI7JDdl39w81VGOyRMeJFWKkdFq/BmHoAwhaV
HUbXX4wCwQa8mmffzPxxE9k55MgybF4eZq3EEnZsNyWBelSqz+/QJY9wZ6FHwFkz/Y5w6u+Nifcv
LNtoUOilXwTAyZLRjgfD7mT94QvFVfVF2C5FwL5VD+xGDTClKt3e3H9xM5bEe67mRJEkVupcEDkY
I0VuBQ3JKz0faR4xrtB4FHBDIexrk1keC7BBm6w55VBNAmgcRdZtM8lC6SPBodlkNgk8hrTnTLEd
QtJo6i3G5q9RyQeKnV3ww/hAkaMLaW1kuVPhOMM/y1/QCiE1Iw+lHLTS+8nuPNLp/2chc+O7XuZG
90/uSty2H4KtPopWQyed0b4YMnvOqtunhwNYpK9ttGJrRA8t973tIUwBdSiZxcCe9TCFSo85El5c
MemknyrFRxHXWPKZnxXPBUzmOjAbD395E1//zlVtU1U+JV30UYKFXJKLfF4C1/1RkqeQRB3+aey4
5iN/AmDcDXvuvIN4ANRn0sqETzfZ/KLrt/m8H6UE4H9SMsFeO19uIKL0/071AbHvHTLA5AgZU42w
dinYyw4reGEFUIB9faw8ODITgbPJeUVJV6NitT3AURRretRCsJ+W1k00lgW/I9Oqg3RhAThylYrh
FSY106Sfvh/Mb/y4+XyPkZOrF7WyWxNi0HQ7mnk65N5a4tFMEu1gwfZgYlWOibszLNcaMkEP5y3P
3EpAXDsIY29RCohUy+0DzKRmlJo3Kb/06jmUa4pk+eYzDyRJ/asTnBpVARzXlbyEH2Cgb+qXIjra
DYxwXJ7YOBNfs1uZ2owhuToP5pQ+nDab6qzNemV+DdTbXM89Xzb+eJYKoKOE3D8/GEtog6lQknfo
wrYag8yPj15f2TMv5yionoyUYcnfPZjA+LtQ3zqJkPZpSn08cbawUk+2QyDr44G2hNaN7YI5+Moe
1vra6dbaWVin5vUeqUtapQIHZ8XEMk33fjL4uyc00DlV2MwJcxGkyTg18EnpTdIaGHA1X1YUl+8E
rDb/ANCtTn/gBbFMx9WxE6MpESULr4R3oa2gokBL5WxsI71iUAeBh/Tnvm4CpoB1EL29847SAdbe
RDLofaG5YF0LIvHESndGcho9E6RuPDe2HP/lfYqlcVcdYBeHAxJHbTjNQrW/PSOLy1pZ3lKJdb2m
DFH37pLS92RHla0rYXozZDD7n7hvMt83twSpBKS60H8J58TIqjjBNtHiNkICZfCFl4NLvTlJCX1h
VKYp0sHDRL9qbGyk0sm+qe21uEMeje9uvlQPkA/J67moImMYSiZWRryDt89oc60g2pOPBLmiFd70
nKdPjDeGEckgg9Gb7Ih164cJMQOgTAFO8xkpOzbxLM7OHc8iZ05qQsAaBKoOTBEjKFdNS3Idk0Yl
NLuxQlgHwauEvv1q8QIqAZ7+jL6HjeoGG2OHh1ooLw9Zfn6brvXV3bQTKY/JWS3Ak5k3/RJ648BR
2dg8tMeI/WhbtPlzsSL/BzNBLbtCkJV1y2oGFYelYw30emWmsk618IlayoTkkuZ4c3HT830YlMaK
+W9pdlgXXHmMzxI11VnSX8hxGek+0WmvrnJNqjXQq1ZRLNQKol9YkGvZ/NmDY9An0RdRs1NWH5Xf
f2FgVEhnssu29n2/r4A15JrygllkPgQOPsOk/4dFgqI1iqrwyKAzJ/WVk7Cy7KoXfTvJQpNLbpwI
O7OFqbp/iyr31cX6P17t5+J3xTn973sdTFZNhwnt9rdcgpv/BdatQ9eLtXxKQeiHsZ0C0H9gNRJX
E0e+pwmQ6K7NPUrbTgPWLNsVUosaTMGB3V9mLerQeYlfNLtdvIqnR7E3FgQeXODnVPkgtkuMUqZj
W7Fi71YGHUJxsjSZPdQf44NS5R0uCPL8PrGrxoD9DQ4Il4AbpGxSQNOJXLJm5e0jU4snr+4BDxaL
GKhLQncYOJODOOGmhCAQas6uHQaAN4+Wjbqh4ScHgJhmFR73tFrCywDJ3VNkyLAmbe2/XFvsGiiv
kLBYOBbd4QrLdx187aCBKyC7gcdsQVaqYiBZ+nx8exZ2f+q6El/05mFvNyBszAYvfY8hoVwXRC72
FMFWFNVVdARNOOLHSI4TX2KED6KKtfLgTMOi/dJBy1SwfiNnl6xPk3OWO18T24heTuhFATghBMok
2fARB1SAJD82mdLcfy5oJ3QFhkBg0tHRIqc3ngz+kIp2ifzOPUtCDdg46aVfkh7PeP89apm7gShi
XaxcbIjLFXRDT2nc4g7zQlTq17GAJLldeVzzZNmNCl/15cTEVsrE0QAvFsL4yJGmc49pqYCy0RTo
KELuhdX7sIptA3K1+at+KDoq4drm6OccPX0lIqwOK2D+tDTMq+1EHm9CnG5icVEzoEMi6mssF775
PUuAfGTf1DMPW2eDu5XNOp2nw5Cdvhot75/hQDZttYzQNrHfC1rik6Tbj1S62E4Iuw3q566aiI/B
F/KxlDx0tGiljwSYuOF268PKDEWQlL9+CPnsLAF/fNjECpPO+YM9Av6vb1A1EEZgWG2UPqtSHkE3
jyiRD41O5tSVC9toSF31lE9+czHpnJNm2Z5Z7gAaMmdcB1mXYSVS9c8QpwP6zT3khscgZoJ25IBo
/mfhx/elvSKkWQvH/PcdSRcaqZkmVXOVvp/GKbpBjN9JkyyohX0c1IofEhJk7TP6maAVisjYqulO
VfdoWGqu2U1v8cYGEZDgTfPUGIwt5m9qCNySrr8PQpDWl8pqLT4Txx8+Lzl71HAZVY4F9L2ZP5ER
bKYz6Cx1T+PbsaeIc0kyxZlcwHRv1juBFeIhcrSigp6M47p9FqNyWHIZePbSNGWpaawcLJyyyy4X
xHbpwHfXAnbdK0PDhL35RH2tPk83pw3co102CpGosa7V8ffrZHZ+xCWE4ysuZFFO6kzgl1IyFZ0d
kABzVzjLh1/NthfczhviWmsfvGR4+6YcYJpX28U2XFPr5pc2vV8+Z/lRqqslnCOX4q3gDp3dsZZw
6M0kerQ22JS2rlihqIlW6kK6KVpTZehlxNJ94EB69R5Nrrw336yK7i5dpZa+WUqran5EsapjeZgs
OgP1vMXj6kraigGEXhV9VSrG0cwUWIuM4wEmQWDQG/xXCN1BsXVYm2VnQi4hEwMbM9zy87Lxn0hz
nlB+xWreATFI6Eh9jAgUum94RYEEzxvr8HxYS/giOjxsdUSeQ1gPR/2R+JX6Erdt5H9yUlJ5WWpC
gu3D7S3qP4HZ8Lm7HtbWiw2yf9EoS8qhKxJVLfcEFbhpyyAPfS0sMM+R5EVVvU6XNMs14l3m89Af
CgDtI9iH40EvmQ0x84HUUdkqjd0n4FQ7/saTTDJWGKBhqJcaXrSLwabjSPJwu9QyrHuPN9A3KvQt
Y7HPWdaNacqUkHDhKqFd7urPOHeCSzh0s95crnJezT3AfuDEAWJyCqa1pjXRujypbOWr41nU+LWe
B9yXjyJ8IXIK24h5DdPqiC9JkkHTRjDWG6qBVitpu1df+WISQqGNa6MnvPijdOXlyO1FmbsjHXtj
X08PDqK5sHqoF3UlKr156FVbc5S6RBqVEUgdR7V+C7XGV9GDv/y8diNmJSUa6ScMu25ZJ4RAl2t/
a7PbcCrhrADx/Vob1022plKiDD0SnMLA+7KUibVhLtW/DxGicyVH4r+xUPx764OXHnniG8BMlk+r
IvjvT17U0HCh2v8jNRt6caXK9OS237CXKBWd54bDp+AiWAhljXaTy9MLu6tB+UITpOv62+K19XzN
XoUmpaHtx94IBEzxFR8+JSQYzld1j+VdgEtVzhEkfoXRyMz6/+9EYvxAJej0RbNtryQNdirhxcgG
aCEA77jCfVZPZSG+mhXiiP2+38QN3WwpeFb+d5BxdpwwObEyJp9XR6W7b//QnZr4YFVWcyF0f9Xk
xgZKUtrYRgSIHD0Sl/D0d3/vj16G8Wf59s9A0uTaf197QRzZsq/raOV+0dYg0kLE0/6fVZhQKtlX
XeKQNPfYx9vvMvC/OSVExsSwdJ6SEcdfCORFAw7aCK1ZTuGlQG6UBbrbg1CZI4p5fRM/IDUYCsLk
oYXR34fZUiAoAGiAQRpOk+YWZtcdHW8liLXWMhTotcojAhWWU8VCUJTRRVxxJyaoR4v1j4os2t84
Qu37GQM0QnpCDkTdoAaftzazaFzq+D2H0NZhqbm/aTI6hMxQFb5N3EewtLjJNpkpkDxfnArsI1VA
xySMygxs3kMa5bqxyvd/iA7EXvME34dHLyFdm48ddkYC8pytzB8AoE06MavHkguWaYgaZLGFlOuR
7ElWU5m8JUd97QSHff05mcO13JEhVqr8MIF+L2wTL6PTMUthTUl4x2WOMP3+gBUdWQ3Q1aN0Mfpm
Gw/SvS9pYeJ8Wp6zM7BkMvIn6GIyaRcete4ULKd8hfmxf1IQLkHVA5nFZyvF8S7lRFRBMSnS+LTc
roL6VA3zidKgnnElha+nXDdHDw1ipFL/qGf40JJAckBtjgEtFbbALMHY3OmF5WYozzCimNTIJdi/
OVsM+Kta+I1ZUrSgesqXTeWf7/oWKCgz3VUnJJCTxUWL75QvHXMACmCaP5khxFG3Cb8np10wgdZP
3hdPBbl+/Mw1/l2q5f92EyavoXH3b+ymhzPoR/HwQHazLjyNc4Vinmp9X16FFNtpaiBSh3YEfQEL
n8atW5Ti1oC0IWVV2evtKrplDuHFCGWT5Ar+YzxQnKGfsv+PKlkSetVbjHuCIKH9+huhVVlNDNZs
O9l6mkWL8Oju+9gpFoDaxSGmRC8pBcp+fpGHhVTBESNZi8xa1gc6UdlpxukQV59nLjZ5aILTcH0V
cQi13iB7do89EtpKMMB6MjJjSStXhaH3MTYVGi9ct6YAlnEW1v1kGWgxpFUaLKjuEVhKNUFsNMLO
uTBD0u+7qstXkYFK1yQsZOP1u7cJ/dmKhUtUmi00NjEs0OMs1KjeF2SIRpVd/HubR03okEgDagAV
uQJyBbRj6x7oVwHAM8hM0Sq76PLyBf6aXrcdUOHQHldlo7JTieo8PwhW+P84fkiEjWBUQUk8CIYV
OAJgjCEIk1qRlWPx9kJVzZukm3ZPaiarVJrEXiYfFHcwWStdIUzp/W1XC7mivQxnWW9zvXtLT9Wo
RYCn55tXWeB6mmAJVq0gH5W+Ra/qz0hJ8ygPo8PccfKiX5Wo3zRIPvyPnpnBPIY7+0AeulDsw/II
5BpsNuOfwT9z4ZYUnmxlz8I8j0ZocPW4pxddlOc9fE3lIhESyjIh47+withUNwTLJiMpoDnX0bS/
Zr3Dc3NeOh2fGAgiAqBy/6pA3r53OOHQyyMKMWXPfVkcGYfHiMJnTb9qZzATDLaN16eezppCqxto
VzEZfwPV+XTeXyDJaseSfxwNhxDOYkvWChYw+KKRinNNVPHjePumwUmfrxZJvCfdhaea1VLMl+Ev
AnHr7MmFoEyrNW3b+Zj4wk2CLmE/AfUXkSprNXKxPSy4e08imy5l6QHgLQ74bSTRjWEOm0Ne8QAo
41jxI7fZwdklouQc7o0YuorT63KEuTjcwRIwF/bIy9DUFCnsNb/8vPVbEVmMaeTjC8bYiIJzvBzM
uUkD629agtYvjg1bac2kXJb/HJe5VQqJ5BR9ILkKtoVXi0C0kPXSrx2TspYJkstYog8cVCK/WA04
tOlmZjsEn7ZizF3jIHevZzL8BH77LOZSLHAw4EFNG4ln722lXpQjed3k2fphHBV+jNmValfjyZFZ
zf3J33Oa3nHZzQf1zSeyVz5ZbsOlJBj2NytA8bMk/a5xZ6PY3TX5+/s+pRGQXNk5XfvJmVPRK0ub
c6Ljkp4lP33uki3u2pOpzYKz4yfUvBTcXC3DGr1pV5wyRP8G+Pa/cr6j+ITPjNzECtLtGwsRPtBE
LK3LsXvUQMcjI0DdcqtdLqO2IiXgw2epgazT8OBXymALbQ5MWOY62tPUtXUl2CPUtAZwKNCO9xgR
3+ffhaWPBUI0JqrWMvBOX6x2rekzhhqfNhHfTHo2Z6ONNGwFobR/8wH77j2abhUce6dsVs6pGoEl
qSrf4+VAdsPmpHT9RYXikeNg3tmvus5HJYZxRXT44/wovz1xZ2tw0z47SCtntcXn5wcTpXk6r/NX
IlpRLLp5NSVHoWmIR52jsYbQK8ZZj35ElMSOYhGV444q4pdVuAYB+3KaLILU1pB332bOs2xOIB3+
oVfLlbGZdFHb0NDKonqEA/5FYgBMCVzUDII9l2qE5fTVlexDtqK+dx3wxdfnDEpPd46WpaB6rAvN
iT2NHQ2DGJ7rlrJjKgkRnHGsFYt9u97FQ/bqLOIVXyIcITKpGpxlGEK8Uf7oY/KHrNoCt0t+lcqo
mMkrKdPk67T7u9GcZELD9yH78vlYVbk0GAlvanYbxnr9lglop7tTtdPYjvPt/2hy3n/v0tD6C9Nf
W435q1NRZI/xluxMlfBI7eCWZVETp2ZkRtVgxXfmgnRWioIOEJs3M7Xp2h06aZFFDEaw9OGLoC1D
cg0O84igZ3RSyvLR7lLOCU769RWBQ5dQpvcuNcF3IXB3gkaopIOfrjdojL0rd4ou/EnLlyWMco1X
jbqRi8P+xb0SvPhU8XetmKmwRb14HiV9tI7XX+KfNjRFsJ4/ck0ibKVeLWkWd66Wl6q8ApDcK0Pk
Hco0T30/d5/LnyXaulo0jXNmtDlVbN/UCUuW4iamT/8vr5CuFojCe+h86f66yxTuNgnMXYuLUHzo
eLh9kjwUIMSVg2+gZ+Drq0Xxpbi1DcnxwFTpkjb7/en3qLzqlIzDA5+qLudxsBLTQvuJipLtYkXJ
EfjgYw4qM1izLsoyGzJGXfeWVNPRjp9/NfwN+uBmlP3GvsMy+5R5HoV5s6ZIGP4it09njbMwcwP1
+BThWL2coEtak16/R7ia6FI0wRUJjA/7wCT4RctJt5Uv7oypVL6huZxlhQXNrNh87yeX66IBBr6v
V152N/oM4G+1iKnTRSQFt5EKoYCsNWtFrWBby04w20MvsQIuo1yCU58wXzvE1brq/9B0P32ehVnY
3NpqeeBmTrfzJlsfzea9kbV1u3cMLjRlIzhSr7WEajaaL0UOQ9V+AqrqEQPOdCLZ+h/9fpdX+g30
yELXbI2KCDxet1jLTDXzf7RdcHuciBaAoGtM6T/1l930dI88xIW2JLG5RXWd450gbzSI8JgBBt08
duTSSCAX2keQc0njXpDNhYrQbXkKafmBjjv5JLJhEMOJdWKgxOysRpO5jekR0hbDpyik76kNVmpW
y1OpsrLCZXyZhKc6na1zjZfcZq45HdjUSsJZICOno7FACsKD660briYw8jyZyr6NyusH+aq8VxJV
v6AKsXv2dUvrjDmVxrr3uLXUtJ1p9J1Fx0BHw6JUV6OPawBOoAYB7dN80EnV5RPwaEFAAXrr7DKj
YCodHUk4F+FRLwjWujoS+aY1DalLjh0mCprSPbWjoTbR8dgZdkgBahOCrjFVpbDVTVfJgubtlfrp
LfD/IjEGEYnLSCFifV4OjfJjVYlbCa3SuOdD0T0/BUdcHGPlvHzaE0Y2fhcH8XGg0XRifFL9b7EV
zdvldPxHwRCof3y0pjjmF9uKmt//mOo0CoVLEoy2aT8Kn4HzzER5pQ9/pMG7gM561abgBrDisJ9D
lE0w585/Ed78/8dtmJ5xXF6jmKxZFPG6jfu7JBfVedUeDRvwB26Y71L5E1kuIuKVnNLLN0IBecU4
eDER6+koW3jvlGhnzAGToe+olsMoQb6bfGJsKP3gS+DnCG9R4B8ZRhboOhoX3mWOZn3FmpyrKwOf
bpBPEhI0qvHUmFO5AoQQ57nGmXn+DLtxRt67U7BEkKzJMHxKhcXnNsMiWeTszXyfcWcSPYHjGolL
saYjV41BN2DtsiPjPL9a3HR5oHPT5f8l/wK74ysNqCbkE0KneYzZPl97h6FjQc26LDI7tyv2ifw5
5b3vpBL7NxTq/QiXnD19V1BbZEn3wM7FFXWHPjiAexGn1vcxJqQFv0dFJKT3l/vIUG9JkEblanYD
buM9WounM5EmhXB9PbGeyPnq/rY8qSttzZipGtWBqvZ5pRvhmBUwMIEgLzULZFDkK5j3/R+2uqGc
0pAoTF9LXmPrM3L9ri1qDU3QjMLB8Wv2/2lNds5K162rDjs0HhS3Jx783tRtnIs2YSv+1PdJI0kn
7EPXB68q4bYdiZGygBMa8W22Gd/VsbSvaW2Kxdd1og2NWIjwJw6nsK/zRyxbqwTB6NqDf9vKuKpD
d2tupv2AKKknG7nPkqXzbWfyocVoarubO71I9S+qUK/IJLWE8ykxc4qm8hveO5OoIS0mhJgQZlKg
KcrpNLn+G1Zk7r3Zoiy894oCZMeLJiJFKHV2p9qwXhPaQn+5KeAZZR3X7HNhnf6XykmUg/FXHNBk
gxngw+pwHu0Fo7OdEobuKpDhqJ6Rbvik2r3ddM8GPf5OS8Qxlj/DDYqAWSpvIiqtqY/odednUDsb
wlb5bKvpUhVxdc5kVaVVmuvcgU2GDvUZeC1g7eOanwyjdccA1VcTGosW5MOl1n9sX5krBe6oRQbm
zLRA+eWolDG9KBArs/4vnxXEVP5UJld5K3Gf9igxLsV/nau39jsNdjC5ZQFOIhZibsD3MNbau+dC
Xb7jGipZ19drFe+uCkbY2LmqB6/Azjwjfjjq+m5PTF6/PLaexxnj7V8bBWjwKcatUYJQTh/9j1kk
V7qdkDlQY6JwF2yeSSXbutnIBnKdEYQK2bJXuwtQrhutoQU/75riB8y7V7spZ+NdMucCK5egR5en
r5eJrwSQbHEQy9cohIwWXNThW4SwzSqfSZVc5+37pWZJJ7Nqx7deklL+H2pgelR/KTRX92R6/JWE
ZtRv72loZ009I3QZRKSbWTFRsYkKqyMe+dfi45TjpFG9lIghgIZqW31L9x8erQFpyb2JevoIj4PB
leJwwr2iCYnwfqOPz1dheRLsUEQn1thcYR0+LDcb6AeFyrCBkvIr2puBssvHnttahzO5CpQdTQhc
XSEUXDNhdHCtp+6KCQSAXpY05QOfOeJxR1MLcSifK3pt9yncy13VvgGGaWGw5wpy4WDUWAdA23vw
g4w7JaO315OdATBHmpjuTtsl2Q7aAEVg6RTfuhbHDdOXj3w3v8dHLRTMk1j0kToTLLWg5P3rTugs
OONgUvmosWsjw5NA8Cw3fizqQwIVtJavlKoYr9onH03n0S95O+FRyy/16XC4pwD66k+upHAlqUlS
LC/8jgqjrkFWH7FZ+ixq66VaVF8huuoOIZ2VCUvyPC3pyNoQWevN7yI2m6ggkLz8VYzjNJUnERsG
FVXvwkAC+eMLfWxHsTPjpPrHZ5O8M0xVZ4kmbJ+mw+OoMRjXWbf0AxCZJwlIgjVn49C3GwjPG8KX
Dv9zMfHgpj1VZjbqNrb5dCxzkNBZNp6ezdtCWyCV+L+VSzi0dbP4XhQbrsUV8uTlf5Ily04LjAg0
mmD4o3s1CK4Uskj1H5K14ij/mS7eRDbQyPQO8UGGsgiYAdsthSvDnICWTUqBSpFfqdfktvCIQ8Ra
/2wI+Y64e49O856J2hunDfYD1roc7ae5rOUkbs/wl5pwHiKZjwdwlmqQh4Nnq1vYvxzOJh6C5iDc
rLKXvM6+oHtG7KUAMw9vClCYX4hY3wh/XJsyX7tkhMqIywMhkPKhf6W+bsb3vLD50RNHtJ60lOpF
va9+ld57ZlYXknIiAlvhg7kM3fQ4cg9ZRynv9C0Cq+IZDjGsT97f9wtK0rxivflwL2B7jaHbLe0A
aPG/n8DpLyhjsDD6Hcf77v8YcVc47tljY1VHUFHblUzHRcSWNxlfotA9Q7T9P2+UIieiNagHt/Dt
R1VvOO7ogrwA7neoZxgFphTz0G31TT2juZlkqID3wES3NJbawmxiZHd+wxYqBRi07KEIXm/0O9sj
ogt+ACgLOE/AKoepT/jWgOaJhvb4CnhlLq5Q66Xuz0DG/NXnTzskJEFbUCwB5CnwLBiAa7lnMH82
7jjEegp/zw50R5j8RRKYMFJ/JAiq4TMVic+e9HW+b6vq6NmonGFyd9HpHoR0ymyJtq/PJ1WDzNAm
TCQ5hrIW/dOWU1G+DOhQCUuSB4ZnSLR/1BxcGKz6s3TGShechT9h++5SIzAEO6J9uXxZjlc2O0OB
iJtZ7gHoyGaAig59vTVkm2VaC8eLTqzvoZLtkuJkV/GC6X22wSWxRDsic+7smH0m9GkSMhpD1hE4
/8nzE+kLNblc0qKPKHdJMkNmwnTYpIc6Zlr9wbyGl9MJzBqE9WeuB1yTWp+NUXzNAfsfyz49Zy2g
Gbr5qJDTa1RhVd4cQkuu++A2/X43jagpkhwSmnqnvxrTmFzjwj5NlYmBGd2kpRKJ+wKvJmggyw6x
db0/bbi/vXPwzUNZIsQgBVeKZk2JdtWWuF9YYswBHhsbIPM4fVEctLZ2dRknvmbqaaxV8hhN8r93
q/FqP2GfIgLOOdbL68KuFZ9YL2ihcZaLv4YLVJWfFW7umBpi+EFB+sZTLzx0/5mMhb4znQ3KQCXE
ZCGEqnWoPWuR/8Lu4apv62SqPTdEgfUpwKJJ/59sxucw9P/0Yk1PijaQmoYw25dAYqVDNFcAxFS+
syrBm8oo4YoxBQVuCaSRCBXAUHpW0bCuLjlxkuWEcM3Czswqkkhn+99xFN9hL0RU8bHsU2q2Q37S
BgcYsdohKjTqt3YvaCM3qTCaZ+hcK3Xa1CYQ9lswu7LVMpQdoma6LhpsVz2wMuZAzbmGc3mlwuc5
Bt1HOE1E6q3JcQBzKq0VV1cX6KyiYngER5KiLV35f5WvQbW59rPlfTNtJOj+WfuPtVRA6KZen91m
Dd+2Rp909jSf1CXn2dOkQ4XvVQg9kKWMp6LbZhDIn+ZWYmFXCGOLje/fegBKUFu6KqlDH2WNjYNN
iYPb7wBEHYBTVd7W3BbZmQalYr79wgO1R/Sb1LUyYo2SR8PiPYaobZeYc+nIKZ+9tuGI7SpaOvGU
bNnE1/qUBNQ0oFId3DoEHvJuxktzwSxF9oSZWjFYqI3CydExxQn7G9oQ8UOF0zB6AmPt/n5r6zqa
GZeg6MLRHayONHZH8yZOpAC/R/KV2P9xe2QCD4fZc7ojCURG8OiG2QDGQViAoB3v5HW37xNB+fyY
gensdc8UY4699TUIPqXrfa1uGbSoFeQ+LCTZvEDE6rGvpDQYyrgV7Gu0LeiDSjVzmqozt8z37IqD
gcQPvHtD4xUdlb0laOJB1M3YKX/oH89jWqb7Lb/jGgrAC/xW/Z12BR/4Uwcpb2bwBRztpM0L9dCA
+bPij8VhSUwemH5W55ElvEAZD1PoqapX5ScV0gADFDkwGNchYe2PDZHor+qJ1pS5hjnZCSBYK+YE
yHbqWTJfU0H9Uu/3FlIbJA+jp4OK36ptaFRqn1z8v4a4HRO/8plv66aRbRrGQXjwL8xZG62WqoIH
z5yE//vn4oFKERit0EWytT75EGkYp86zR9/eKwEFYvRWZ0Wz1p2A3VQQPdwnVvzuXx0BH1mPg8mF
vRwnmN0878ASWksuggYZ3awdcqUyBjXohNV5/GYd7l/A21nW00nIbNT9yUmp9P7gyotrovFDNXjN
qdwC8QwWQUfNch7IxSb8/vgds1BxQQPjVEQPkG4w0xgnEYhBrOIAOmZCS54qp5xR6HxmnWGGjhMY
4AHYjb2FY4d9qz8hnyQQwH8JLEM2uCe4dnjqyKIyt9s3G8YvoSmXXF6tJveoB3Y8y4b/pisiBlku
5buon2n2a6q+l+UGrWh4ol5a4RBQrhwuSs9byqP0/JolTcTiW4VNYj29HpeZD8H9eZ6R+nxJgON7
KesLL3MHv5pghBMSzR4BlohyCp0p3HmuCQrPfoPMLj4RZS/u+HWsFeNbRvMTZAnfo4dKvA3/jYNW
L8B49YEhNKLNkE/UzpHpOJBJBTBg4JVKaAIK+xRWIJbZqS2+/3y44VSpAdMWgZNydiu394Y5og/Y
68Qnm1WNaz+pWWSGLPP3/2tJvf1BrNf9uSvZMDzYcZSgTCo4FstxuoX4sIQUha8qKjYV9ybiwpBA
xVfxgsGOzsp6saFRZBlEUcFBNZc77n8+BCG+TDTv5+ry5VYNsi3TTQwHla1LixCBVFtbaFxFdw5Z
9KnifrDTs71cM3KgDEaOEO6e7vNA8Da9nB0idFRztZ4N0UzS+YZX9rxvEx92Sb0x35iZ614YorKT
dr8WlxGxGWsSDvzt6NBZLh/Oy2smor879ebKr1uCzY6rRebn7JHUU/GtDEFlUsAEjT6cug4rnguz
PxpwoxmAOx3fVyLQTG8MBbPpRaOgNi85BFJiWNDgId3tlqyek2GB0Q/PdWWhkRX2n1i3nh6LcwRd
ChcVLlbeg238mzl4jTZ43l7FHB2LlBe4S7/ERRREOfC64wx8suK60tmHGP++thGEan3u60zgT9FG
IviEOPBRfERdqMdHHr+rO0ocVTvdKKkbs6D5La1yyec/57huyBQTLx3JzMnWKo7CcKj3Aw0tJsoi
OLeapCS39N+Ld3idchuDuSh/qXa6WILOsjN9FjsfR+ffHgyr4RMbbb9/fWJ5HRUEi5ysFCX7Y1es
Epttr0FExcvVWhS8/mtsX6EX4k3C/ciN2xDQvh8DLl27nJk1M1VPehROQOkD7vhTelAgKtRBfAGf
G+1ofqZdtz2JO1YdEbQ/Rkb9jL7lrb6ZQx0AbmK3Qa1m9TUljzsgeIBecKgvuPpjqRe3JiXJJa6v
cCS23GcTTOi17aiYBa3scwfLyRUsLKTMmELpiBNRs3x3s0EDaZLkR72woPNaVbKo6eBixKj82kUU
IIHSh93KUAyFABfuZb1qY+f7i//SwY54GrabLojwibtCJAbQX9CTLchEWoDlmJCHcuAiXVd7kYUK
+R+1gfcBdRD0jEL4V7eaYDhjS08dv2aiLD0quLzTPFXbOvQgBN0t2Z6bD0j85NHtZQPc465/ma+m
DjdvH3SosKZrUe+Up+cg2GoXbsAmeNE9gVFNT+AjkGemUmCIvq3NU6kT3McI85zdJGx9qJon+hCN
4mRazLbNrtPc+/uKcbWXcMd1q4myveP+1eV8APayVi9sb9TIGysGUl4CdGHyFclb/BAShUIXV4Au
ooUSfdf9bcvLV7cqD4C5fDhsUIAN2OqATidemC+OHc/4foXY7GHLaQknCfZvC7QPD9t65SmCUw96
QV6maEV2anUG65n2qALPyHMLb7O+Ebhs0pUo1fBCooVQ7erpXXtoQ4IThyfej/Mu5UmtlcfLmvsN
VsFcSIX/YHpkYPmabw97cKYoI16zkad+MawR4uqUYK23FO0xSX6mCLViRfISlEGoaU3nuy3LpIC+
OkTYzrt6wwIthY2kuJYTHtV8aochknhmW0WKYw3VDZrAlO4vB1rOGSVnSmTDGHHWAFdDDw3UHYqj
3RVWJ/xHaLkQDWgSTDI+kyPyRWxBGI/jr32Fzq+d0nXHWKgTYB/qO4Ex9TIh5wOPgMqtSFr0mmwS
Vm5hG69qkJ0IQnvJyK6upQiHxc3Ad50ruZ5H+HNdHJ7FLG9X3J1mRRot9p39Hb1/Z3uenujUWWCY
S0d5AOqKqsFSivR6Y18TiKPo+22ibv0aUVLB5ea356a/m8vnFrimJAoh5Ql1EaeTKLrPpBG0/6tW
Ds0dgrnn/sKAB+5hQqTX3fn2bK+ATsJEZhxrswBVV+zJ4GJkY+5PIKPB60Yz3YsXoGz7ZMyblmOY
uminPZFgUk9Y35JWrkG9PE7ty9QgpUHK0lHWGwaL1BTqbBRABdlRlQNLT06RnS/2lrq2AOUulAZs
Bgko+Ao/DVlJbCXMYjOSSil+XdzHsm1rw/ZuojrAxwxXu6y55oQUauZD6rDJKBCyJxRvYiNdFwU6
/JBoWTVU56joni50TYBBI548gdtDkU0lagEMggfj/uhg1Blq3In/8k9JE5TlZ9T1SYF6FEXjzP9t
jJRMX8ssYgcyUjIbxMRI430ZkFzRvzJtZh7Rt7KY74zfIl1QgRxt9v1n8SeQnckEWsC1cH06nVlL
XfBL5moZ00/NQb5TTv2tsZitRBQGFjRIZFgzI55MKXu9apSkApINEZ15fUCNw5UliRmru55A0V9E
dwE4zbZ1RIYSnyLmqlvnOetjyzxE5YrS5kzKdV80EQV/46EF2++UIjR65MffqpX4M8YajqYjvr05
6BpE5vr0ikydOVjSy21w+TuX9Ey6inWFZo5dcUuYZIFY2s+7dlY2BloNm+mAjelmY/L/Jxlp15DA
sUEU48mFLKhQ/duRiu4D6V3EAr/KC24qdmxes+UKY1SwXB8iXCxlPQ04ZEdOa2Hwpj9q4UAMewdm
h9YFVBEnpN8WMocCm8DPLfIpr78WZGD/SPm+J9dZWvoNAF2CR1m2ol93qUEa4LHPSZKMSkRI1RZr
FuBrqaYYdcjsn7n69V1gnrdmbFFCv/2270iYgRFHV4OHCubsiKPSjaJkgTs8G41Giopv1k/cgwL1
A7NPX3Az3FW2UtoJxPszEeEc9b14tXMr8sOfiLzZo+8n5KQLuA4rYgP895C7fQQQ/N5BA1P4Jf4W
c2FN0ra3CZAmg5or2ZH+dC+H4ZgVf3MqrOiG2MQWYUqxeDBzUtW1uQEaBQbsTxSsMx32qb9CST03
UwJgqG2elCF9c1yIFgqRnSvwolSGEDw4T/hpvLEI0kSnw6+fFrmY9ISg8NYp8+G2EWew82q9OoxC
/n5m9OY4fKaWSCWJGuUgoYHLmrBEMTnZ9g0Q8DHhclzFoBg/0Vht+9Mu3coqbnjSnc3YRQ7LHt62
rAN0ZEv8S9NIB6ZqIUfd08afGTlIpsLjrGLuOhaezwVhhZF83zS9o+EDbCngoMUTOWKTFq8EHXNL
7C9+Scvm1k9GvwQ5ly1+/3nVqj79exv8KNjdOejhlMmEmchE6wrQWCAjCWdxMsK9r2dCYkWGOvRf
nevIBDb4NaaMk+maCz0x3WYKs8hGgvqZ3YdEQoZqsaq43FSCLdaOBwglWr/8zGbuUuWv9C1BBWon
IOy8RC98w1ggvHYGDgSl75mOMYKa9thgCcYUCQmJSyETyIIDqkqHCRWzgKE0L2HBFFGBS25gWOMS
T7cROlmf88GUq3fPyozid3k/VcayEtY+aH8skOq9GAnH0yLlOEoZ/Ise8H1SNNOifQN2o8SrywIC
dJPY3MG2mlrTm6dyEjNLkp5AA2TZVTYS4Nz4SnImEVfmV8DhQ56Hm4MZkw5f8+EsbKuOyHo7jQta
02qKWioJIfODaditlqREg87vOtVuTsVX0mC01fMQz1rO9sbgTc8k1CYFl53l8jP9CLH/N2iS0N2h
dk6se6F617bxb5UvbUyGRiqfl7MpA16XCK2BtEn6UQH5UKfhtw85A8IPz5eopEP5kScJRXbV9hDh
KdqnkU9EbbjnXesHGBtbc+fcumBZXNxiw4fokjNurzeKo1eYqWUFVNTJi67mP1KDV/lmg7Kn60uc
lFuaEMFGdKRj7JjpaKE5oH5odAJHn0ggc6fd+nh6EeewsY8wqDOUsW151PaaxnjJ4mHkdLQTkeAn
lqZlrZjjBqqg7NqGiWJ0ATUVahqdnL3TpvgGicZd4mBW7mYbhdV1xpqHsjgWpDhwcdjJv/jGFbCL
1KtFB/5DgpFAVMl43VoLHHFYS+7Z8wz9gAbbBd5T2DTjYjKdA57V1K5gQPRM1XQ8YJ0J8ZVPo3ts
x72UqakS0hed80P64NeO9t3Tiq3SuE9KWd1HE8pQF9ABOlOaMG5BrwygdfF/Ccu3nG+0trPZ1Emd
GPXQnimE7Zopl1ZObU93Ehbt5/TVIqmwJdDmCnwoJiZ7TbF1Du6no+U0H0FDnnlRLGidsHIcbnP4
q+XWaknkzNyrNgySzyO8cwwFMMdlDzB6VZIUjLrecho8qSRkz1PvzZrewrlMpUBTcv7TTAqmON9E
xHwgu0MgQQPkq37XG7jrMiLKhdfNXQAH79jGwilGeRZ8mhLoe+Bx8ur/HOVcweALmQLCHUTg7uOu
ND+B1koNBVAHkWTfXMeBtYWQPG6lkuvU6E8Bza/0gZuiFvkV3pN284tg75auagUECLqc3cNuWYQI
vm8AeOthCTnddHYL4YcN0wcoORPd7NZkK0DI7/6wZYv4A+5Q+7jfsojD7TSMDYhyMfTHM15mzovW
iPoIK4HcQfmPt1/ieMBQ+zZU/nj/aTznVu6TkqdMf9etGWQO9Jc3OXmclJcBaNJjIgBu6C9/PwMt
63KmhrHNsNlzgpbM7fNTl3TzmOQ3I4fY1xY9T52keJ4cu5UcHXy2d5gxkcpnGMNPzSU9qmqGS6y+
83pTkPS6pituCMxUaF01hZFHFMnR/rPnA77mHzeGK2XhhPhBsllNgYks5lu87t2rTIeGIJHDglZm
ImHDLHSipZ/pelagchhjqsbUEbhA8mBdDoruVBecWgUnfP1Wz3gvuGnhJxJBd6gUxv4owU1U4XLh
jdXqzqn8eCzNZi6qLdTM0jDTMdQBomHCqYGzRPl44Szyu/xobGu0EzMyzuF8yxWynYujhRNaUMN7
T+Z3mYnw/POj+K27RcMxOkEgZgi+8OsYIXFN4R2YayWuRevXpGdrDrH5djSj9KPDgzBq18AIkXnC
X1q+RYYUFVLwPFRooRBuiSGpOVt6lXGKZJPXiVyzOfNC3NHi+v9XGjSNSCr4PUOGdxCfDyReNGvv
O3Hx6Tgd5ARmZ8ihRLcMGTPcjNVW4qg+oaSVa1y4rTcnMNCe08DVBPM1h1htMc98AWr2zDzDY2Gg
FKD4WMc0PN7/+M6eaJwdzQNsBYPVI9ptKrhLEE3qIJlEfnKpSxJzJbaU1ZhiFdH0vdLqC+L/MuZh
KFJycVsvtsqSWhalW/jebxgC/5hAr7AB+na61MebvYwS0ZqH62HoP2qXIllLo6pimhIuBDMqFqDE
Z0LjOb47FzWSwwcedNXJI/wBnGAZXFQnkllvaomAgVUvRSAqwQokrY8Ai+SE4ZWIDe0QvRR8sTb4
hM1ky789TCAGpFWvwcEsAJdBriv7ok8M5yHiqxi7nyTFneOcbkzdmR4bKiDomoGJKv9XM1d++C3I
+aZ6UEHDEAMQ68xXlKM+LJLZy7+P30mzTK0wKfIi2GOJS6xxMe23mQ/gmBLU6S4a/lqxEOpEWzrJ
cyjfPglujKZT6KGlQK0Cg1yTVzGp7YNmxIYOXNLTGvbMnhy9HhYZoRS3TYknA1jEqiStBH5Xn2/k
TvHMMCgsd/AUAlX1/EtRYq3IeQ6DsMgFbD++zgA7xL4Gqjrhp7AF2LjZU777tCVH3EOv0alSOoYt
Y4PHaAYJTbq1VtCyxHkQnB+HhHtnazuqYmadASs8E1+07sAGslnfQoOlwvClO8OwpG7ub1rqn11s
BgU47xHnEMC8jXe9JQSta+YGxqgnCWmNc6kYWCDiKyyrY9ZdNh1g3NS86jKBtU2LhtHTAMgnFLrJ
ut7IIZ1QjDiSB4ZUCQgCHQeccKKL+B2yn6y5cU2ltJbL/8fbk7DXuYCtwIA1k6p7rpY6atULdGx7
C3Mve1//08a6Q7jcjm59hr9M5O8rHsH/HB99xIpwdIGxgH/TO2ZKZRwpTl6eHX/gugeZC7bP+NSY
0avj8XUB/hBxAg0KEXLC3CDgLpJ7Tci2fIwNT5tZRTR3XuW7eZWof8V+9psEKUctZ5Z1XmxftLpn
a78kCwygkCdso7rnLsow23M+PQfKbi3t9dMwXOGucUb1TL+LHtsnYzj5VGbH4g3il5F8SONoqY7m
dTf9BBxpIRLkmDHTxaEyd3AKFHC/lFD0Pf1cDqScB3sve4oWkAoh7wIXGkglcRJZTE+nvVwXBrcl
pqYCdgP9sMRb/xYWAoi6insGoUiR2ekplIIRajN+Hx+XmdklDGntUejxlcMtX9mXLONEZz1yNJCz
4Wrllp+Ic6j0PrKQLlLCygyUe3j5czIcSjlP47SgQKowrYskVyahw9ouwaNFt+nQFNGBU55cdK3C
6J7omy3u/6ndF2sK/YUctAlfasWJp0V5/p6eN0pvBrxfl0TdTIFedHHF3MJzvzFV40ZEQQIiD8Ex
dcIXFZTHofU4G0exo+XA4Q7rpcK3Rsd0SpZykV4XD3STghVZwWE9GE/7Vm0EeA8CjgiQY3TWnwAH
GWF4YkodjY36bbd11QKYviX8CXfjyLfqFtSGXgUKQFw8Yxk9gYyMfh7+YNiI8wAA+pf2N30rIlR0
tfLWvZYXkbJBzG53bPU9TBQdmAaNyYf6K7csEVZuTl7cMntctoUylUzCSPrPZNtKMglZVO3pQXr1
kJ1KTST2tr1F3hBiFK273/DBDMhAfR2JenoE9CW+JJD5+4uzx0CgzSETtiyRdObgaCxDXGtQ6pkr
i0SH6YdRLTiKhRyZbvJcZX/4/OpZ2eAnyFWEzu7sS4fduqPuTQfnbkE2dIe3mC0mlgxxDACgfyNj
HJycPNTZEqHBELUij/OwEFQVhAUL8fLUHGavFW7gscFlY+MW0kciPkUfjaARz33A5iEwEGPD4fvp
A5GkfqvyrHYQRpozqfgm8tltgMVkjIV2HF0kagDAbu6JjDoB8lyl21xlv0LB2V1rD+sfZCuhaTFa
h01a3h4M/XDxR62Ctbp1SkWDbncRJVA9Hd2KM5elHRW6H34QzBfwfPM2KtB0aj0t5kcHXR4RlZ5x
G4hwu5+8vnG2UqeNYXkfWdpXKMszhJMuSj3Bk+fOzC4BdHI2+K97ocynBJSZEvJmrLG/IvM181Cb
ERu8fvLU/yOjrlmaw/wGXLq1fdQz5OeCCMVirxOjVlmPldeQNizROUp5NYHjkazZBxf7igRWzUu9
UNbZ55lVoJ4mVW4/Qx7d/1xX33rFjX+f/UV44YgKGIy9eXMxHVR6nwcvF2JSjxssDIWawsfEcSXE
1Rgajk9Cq1bfuZ6IUlW/nRG04VYqIXuP4YBa2YXXk0bBnQurcQePOZjhlssk4JIiDNhn+RagUrVk
gP6caORymCaMoSMc1gyIjnCbTjkPKbAsLEXjLJv3E8r4aYekaW7POmsbCfEzahPAQN9X/3sFBbXc
kLGJ7kBM54lBstAFK8cp2gKln60/g6nZhzddqbEQF6hVlrX+PwpiNT4cDR0JgiYnDdmd60jK8247
m7vEAA8j8zgxKRTw7ZRalTFvdBE+Tvx934rWVek+Q0G/0kBPkCwco+tgW5KD2GyER16yH7P0jZLc
Zr8ArzjxXggOA2JfCelZ5CZkx2aDyDJ9a44qbx5c5hzgwadPUhOu/CzA/oVRuIiwlzkIe4xtBxnm
zWbj0s7AxuuL29VpoFy4Q7Td8xHnQbgQspPpMgRiFO5nQ4tt3JxyJGEDEHCYjSq9LPoP+yyI8/zR
aozaTXdCevVEuy8ju/hPU6N9DZmJHKrZSuNMgJfjCvS+zymyfEVwv0joAapFoBzmV49LR7OXubKU
tYIfpBz0WFrKJCkjrb9s+j0QBBtjYdJORmDK69h4zJHsDIgel2eFTqojYqDoXZDh2kWHR1z0lLQC
TSNuXWICobJ0qsE0jRjxoQ5hTMzq2QiOnSiXPUMgLnQqE0Jq+I+WIi3AQNR/InrWHDYBxKq1+IL8
eM+tK9V5+IJJF9yLWXj/fbIx6DXSy8qNX+9DfboEarBo5yu6xrY6ySZfZArOeO1JR8x/9LyutHeL
vFWeRDBTL+bVng2qqISmFKse/wAAHoDdFd3Yb6oyk7NtsTg3n8TzpNfiz0vEexYPrymtmcmYBR1H
qnhoRCoAvHky3sPTz2vCmgO+e+Tnnrt6wo5DfvTey/tfpKVMhw8lpQn8U9u/+U9MGPidi8KiVroB
xO2ZZYOHSeS9pDmsmbUxe7IeYByHtDTdEiHiKeh3z94TmKZtWLmBgC5wrOWIhWP4m59JLyDfN0DH
6ZHAA07QBTRj8DP2z4b+OGe9em/Okl7QpkauwJzG13xmnkw6JKtreiQl/TbGF07jpgVnedjx7uq4
Zzkq/Yh8rXZ+Vpx7F+2Dxfl0gZgN6UibjFztQgRi7WWHuXYKN7usxP9LRmr4ytpYLbhgLKOCnQ6o
0pGgLxK0yBsDRboX1LT2LKGw/R5sFJEnArLf50qtuMafZTLHI+i4dYxdEqEvxENfViFFQuhI/cDn
fJfmIJeGR90JICUdbw96Qtq1m3eb/URkN8tjQzJA/C0aN+5ubfaw2hp8luMlvR1f29rfFEb0oaSd
NeSCRVEIB7267EelzYMtlS7LvbZHifb+j0yGwbJtP9HzGmgdEyw05y3a+x9aS4Inc9kGm1M5pzcN
5cZadCpRg22RRubZBrfDoPwbI1AEFcwGSu2a++zAQr/Fea7F2w3UP4tKAD66Ukp9GVxNpjVq5DaT
hGz5XVJQc6dmLW6Y0ag4NwGhRUhpFXHLKoJI1mIMsPrzL6MjCAcUy3AcYjQo/LD3E5nCAZQ4iuQC
DBtcT5SjnEb7fKKc8gqTzWLe8K4/flKWO6okiAUhCs+SyfKOizQiFLj2Gd5lQQdRH5VxjHvLLjJG
/XGX6cQmHutQOi7GMDn8GPmImACwf+xb5DzEclPN1owWFMYbaEFUf23qBkqIfPlfjoglgZZpgEnG
kdgQidLIekeBGUBAV+CFGT3BXkDWxD48IZruNEf174l6Je5J4f8tX0DuQqAU0onCyikbL/a+v2+e
GCyIFaYdYl72vVQHSK+Mf6FkHcaIVtOiMXUGYduS3+KyH6JfabSSbU2ba1Sk6VuWVVxU60D1hsTy
+CueQFKm4hmMI0qSOIm4tXo5ECMoqKpNlaQoAIwARbOgYQJy5iaufiW5V5eQikfK4mw3IQHpld3P
5qchBB/f332lCcCiBqg+0sHJ3mitzpTixmMFR2/LPtIz7cx3ImyPdqBJwMntbgmswKTWZZvG6eTE
WuIoVo1B8U/MWm3hw8c4dk0JaZSACHXrn0b5cTs2dGO/Ov4kjq7+ypuhJo5l4eN6GXRIHPjiPQDw
D1KLznTNaYVdQRQgGUvUgFflXxxFz/hh5giTqWPxkAYy/sa1O72xZhBG5JX0tLjFPz9X9/ifa9Ce
ArCqO1X3c30fpFRrcI0VGHm7q+Ac4HmXjlKjmSv2IMjIdw4FNk8Q/Z7marnBZ0/zItMOHGrbdY79
bq9C56GSm8kZMo59YP9Uk5zE3p0giR30GMQBxfWBKQu5BErwArpnoiwJyYWwlydL3DJhsBZwmk16
zLHJBJ0bZYArkSmM+5KdCHuYT9gpuhwoMaXwVK75FbKNxyHog+GmrFDBbSu2DYfNgS6XGU3iRFG5
nXEgkTC28kM7LVaJ9sJfgw4Ab5fxNNAHtHPCxiHOnWmNK6lYoST2IHbt5BNPhH0rrp04J2teENYW
V6d19n0p3RzqZof9tVGgZ4Kh2NdCVDmbyt2Iy4wQYMIecArBTN4QGR04rPrN5ZsrZRs0PyY6YJPA
/ChvhKjBNaN9c0Q55NV7EDicEGoCIzD4VMpR2+G40UwVodZd0zFY7SFXRAqN53xnmmHnDQXOnKem
NBFRwDjCGpM7UeoWeC/ixzPt5NuSU8ykWCQNL0yLKAwEaIk/bqo2vb96eL1yCf+UPnaTyQJuFsVt
msEwltoFQNIZu+KG/RzVORAydQh92912cRYpE0ETrSSoGRN5GknjyLMuzOhne1zNj0I/hfSXe4Ve
n1WuY8tkX03OqXbA3UgyOH+y9YiNetTkDrgxbL9zGk0XiBDSkHk7wAt5z7lS9ZmJ7H+LAVmugoru
9cwnrvKjxW3QnAgSwu5fTNzf6VEQdLS9zBMBdoZyL/OsaidExHfqIAfccn33i1Ly5avQmBrbZmuu
cJaG+wt2NPt6OZUM58LSopMkFX5fPPVzZ0no1kpKovBFhITYCQVdRxCTT0dYkc+0LwtHUyOvyr1Z
6cX5LSJJowc75xtv+6jLc2zld9VfgryPWud9Lmo5Ea2Bu/ZoAIJ6qQK4dH9m4V/fg2btUF9uygsy
fvjcrpRgAl1+acu4btPgDs+ILKbANvV4fEhA8Ui075lJMu/qB6Nfy+EZVFkT+fV4uSt9aQAiwD8W
u27bkH0AO5WbVJy23rFJvMo5hniO0D1SIcrRM2mr38vFBLnzlprJFtKUtG9YMcqU/7Dc+44lPr3P
qrbRO3twtsPaxhhi+pvAoZtsxWrTlzDQu49ke9V3OnZUIolzM6JkhwXFgyEncotC6ZQCzarB5+iG
W21SLR5T1M3ew/cZKCL0IORh56IG7IwlhvngN8djlN9mnJvT84Dor36uRsLnvw8T8OAAG1vcjztk
Ky+MeD/iKfKJRXoTPc5iuTpAl/iJEFejG32ve35TVyX07VsXyjhRmr0V+eWq9ylIqC184DMHYJp5
EDGn8OygTFwh2sE/9+VopBixflOvPhueVXFPhbX4SSmzvVNO6uKXEGFt2WBeEvxLxK1kiJlCAbno
LQBAmkGlU30uA0gRMNT5KgLo3HW516cdLf51mitICC6bSXcth7dSfKAkWBLYbNW0coE7l80jcqAE
bQmCdhki9smCp1kQlXKWzaGuZWF+2dAAyOuqz3iJKf06ksHIPPB0b3KYSWTWjTYFWB2cDsuZkRId
O9/0YaivgWbTizODZtANFcQnEOCC8ksWEtLa6rz3dGjGbreOtwlWlz/c6NxPoag1aVGmb7RX5cI0
AMjvMR4f7qWHV4/ec88flXkcvwq5wt5j7mpfVPRcTxxTyz9hKh9vtgNlRPX3aFimGR8G1mrf0t4O
J64qnMohI+UV4f1+ZI7YmjvfDlPITO8pUuMa7hkp7T7MLZWylfbc+46SToRj8yKvctVsrFM5rV6+
mvBBPjsPbMnyk6lxNSYrENOZKWboWPlg6J6Xn4qR7M4tSh3KXVJRw0hMkgUq990fnW/NBNMD5s6+
HQrDNU1wNrS1lL9HOoAVJMzSTZ0b6y7TuNcXvTs6+OImYXvRR1/qCiQ4NZ45doQ0opI8x0iewu7s
oK1nTM7UAqzglrHVu3dWIAmIJWBzQAiUdGKp3pQGbaWlg9Gg3f0LEZk9zkNqsLzPtvOk8IEtkU3d
R+GyAAUSLK5WIl8gZM0iGI/yBcJqqbkS+4MXAQ0PobGNOm0H8Vpc+Y9jqdrADClPYPEhFA6ZtMlY
DxQT9w4hI+dfqfKpY0AtfnZjy6gz3MfwfOnoSSX2MwjEkeJoyaxgi3WXmUAoUYRF2nNA/Ykm4mUV
oxfv7Np3Lh7dtQJbeEcd3mwkASFE2QPlopLD3ObNlesclbXEmUFcY1xtIO02pD5vwtBUS+dF5df7
FhM8pvecvVoTCf5h4xoIXP+7hH0K/srY3DOOCrvSKH+dhb2SsbgaFs3kgRkfmowq1xkIBJyDa9VV
A2l2whVgWxkqP6/in9TaU1IeCVT/u33erBeHFWle1MdqAw8o0l1sZdtrmtOA3rhovJnQUhPXUrG9
wrHmmkFQ4vRU3HMLamOCrwerjSnUSrp3HarRyw4+OvOpBM7SAkaTrymey21xCZcvCdeLm+Bb8uDq
mf7/dvk7hjVf6tRmGpolPDdpm4BAq0Ri2Ho16wwR5Knfi20FSPtzIkbsW8Apu2v4Maih5LuH18ww
crutBD98/Fk86Lc2cEaGM2/+eGD0fjgHJ5qjkTQXYRSPGpk1x3GS76KarB9R0GFONAZeXr7/u7FS
tB2nyP8DDtsXnBdy/ZKHho7+43gFHCAHf4+n9HwKwV8o3YwIaRFyw7Zm97DAK6U07Yzp4axO/67Q
FYXYonXs6uwc7RKM/RLN4sJTLPs8vMiIsTQcZJkAZiUM++TI5pmO1++H4GbHGKEkiFyCaDMBO9Gj
W92g+wD2i2CqnnNW2qDJMl4SyxmSMHIdXLlB9/zfNLLBJtsC/RBYbknIQshf48sTQ2dIKFng8UNF
oGM/yzGdO7ojKTVzzOOy/HwrSLUEcXAnsDywJXc2cZuR8bTt43ukaf9hFRPjAsVXbzc3qtHvCRsY
TdiWJ8eG269MKg2uAKAFFyFWxkPcsMTVUBb9l8oG4gc8DQU5XkAxyCJZEPPRanjBs7Z8IC37+4lW
jJGIMWswIVR8ap1ylUD63FF3tzWzlIIkRvQK5rpai9MVG1Dcv3P1HVEvbn/rwIl96HPtWBK2v1NW
astSF/cAZMpubqE9cWrdr1wRgIjTBlLhPqOUhTZypdkrCXETOGMMTjZSNiEQmuCStCdC99PdLswW
AdHcZgex3/KcRdqbATTbvKFNxc8tUI5IsxTyD9OFLXTLDStk4UJTIcQ9EatABL+NR5KHoH5DLFGZ
XO2awbREwBBng8H6bKB7SmWapl1Z3YyMA2mHUxl+P61TS9ZAl8jVlLobeVVyXWX1xIYgzSJKYvaC
CSB6tGFeTCBqsRFIxahGyOrPpgwHYE/ahU6am2M5tG/kmI1wdMPKC1tvfrt5SWdqKIph4xuL/Jib
noj+lEIdXKmewHJnG5J5/im6hS2CAvne00MDTPDG6R/AXT74qR/MI4ksQXv5NdY1bcY2j40FSW+v
jxhQmuWA47R4MTPH15TP0COP6bznU0siDYCy2kigMdt6yLtM4FKsbngdLgi643DqtFzcyRS6hZa5
k2xiwZxzNQAt3VhjCA8UUhCKuU2SLdEBWqg02+vM4x8E1JT+Qhwy8Q+lpQud+QwApvesfS03RcEa
QC2EylPVJrAom1W//y6ipXufWqSvO3urOLCCycCFCJDyk2GBouzeYXN66A+Zs8fjjBrXp00UziX9
BcAzBC45V/HxwiSGwN+M2XY0nfurPheRDntWZkoAbz8X+FSl3jXc5/VFuM/5RNZF9leztaJKag5m
7O+joNy8vrQOF4QiUIuD2KdX22SBMuzbji6gDnJB9Elb4OiwtCion7VtGZcxDntnSZpXp8Y7RuFx
KtQn0A3SUFJF1oWHSobxP5uArB0uBeJz0bMX/8vWoQiuS14lFTh7A9iq3UGYcFHkkgJbvvShsaRS
vPfCZSsyC49bEpqqgT0ENf4BJsyXmiMpzAwV9+KP2azM0jmaLIxrc9XsDP40tB9ohC0/G/IMZLL5
GmV/G8ukKG99DYXoDfzo7d1bIGcelgZjBc2Z8eU9rsaWOapUWPpZm1xY9q0Zbgwj8G0PSpXUtI+1
lF0wkXD0lNivVLEBHK3Huf0quC1F3yQ3r7UdtTUdnVRBTVJF4zQInPY23gK07Wso5phUAj/gXYeS
k+hDGgJwKdQ+S7HGwLEecFL/Q0pfgsNnFDkrENTzD7epmtISfiiLmjWzrr2+/U82+Uv99UipkguE
DYQVkcfh2vVrCg7sOn0oeoRBRRbm4qyCSZbDNkjklpeTwqROO6jrRw+JTMnIjrb0x7XOuPZ6Yj7u
mtRvDTE6IfKkevWQsqTQoiPWw05+ilYHdnqd7fL4KxBUrc7buenkz7gIatF+3k4soa7Ss1BVLKBI
6WS10WeD1kRAI5uOdgVknFMgpCP51LV/AFVMsE4VVQAQDhyitZZ0+N4677ZqSZwcXZ6FF0Jn7fi1
B5/hDDJBbz6zcPRXhmx0p+qIhBEjO7ak745+9z+D0JdLjQGewPLMx0cc5uqqaVxSgBxpE7x3T3UL
l6WxwdOhJlbHpSCG28g6tJcItdKoy4QMmFxwFhbbXI2f7DZpDR2OCzm6fHzvufxvNgP83WKE2I91
WTEIw01S5CECIQSeY6PGBRrW2VglZPxUbSsBIINcGnSXegMQ6q6c69W8oL05KFr1fpv/mxSfzgQi
Z1PmsX53xYcMKjTw+XDN9DZLTAIuMy7xVGxBieU0g8oTypSi50gjKajewlWM4yjU/9uAgqfXTgJs
jx3YvB3+bFoUFFkNgl5VztDwaxbCKwyQUaizpHTZsTnCF5988blRgoBtHjRzqjMJUfUSpVQd0/3t
6cY8GKnYjzwmVLBiahZ1x/rHkr1uvvnsf3VFE52lpyachV2wdO79JM1OIESuaN4Dgk9jwD9K4DZq
yWgFqI/3/9QeDx03PCIpoPsgOpN4CAkYXvqjUt4iQQyV5D2K3SdK9J4KsjAZ+wHZ6ZHW6whTDGfB
rVSyrJu6twKuQNezZSjYqJNssgu9V5kvUmgZjdbBafyxkIETtI6gUhXDJcpNo9Ivr1x1NqbTwMY0
mTbIMui5eGBB9j8ePMpTBf3F1zlOQFqqaSxfAsjg942EdCjiRtUnpu8KV2AnyJ4blScklweUNTzV
I1doZo3MwpN6y4p/zebBIGYQy9nCZHtigbBaVoo5DdHL5+8fuDRbn8C3tIjB8Z4Fcne0PtFs8jkL
CuBKuT6kHrOaZGkqFVdh7QUHqxEZ9McmqSoh9cJuzrRcwqfsif8Vcya+uk//QX99fl8uL++33K8t
KlQFmTy9oPieC9PvVkAadTQygK4rF70cpEDiTG7nb/mAj6woAQ1xUgl2GequDYBfWZLjpGwxusdZ
NZpVib4dqXdjlfhQo4tm/XPcC47fx/OQY5fbNd6AoVbCSnxYdSgEUgRlbI5zh2KjAHek0am2Z0tG
Smct8JBWc7kDHFaTXQr3diq7Ju3PO2AfNVutouy8xBPNydxX2VhenJ1jrPHGC2NFFr6QbtxXF+l5
L2sLdftBoD8VJGKZ3/+6THfI0PzJVhjGblUD7RoCaHdGF+MniDOoTMN2tq4fFepSbVi5wAdjmat0
mt+Svssp7kGH6iUbBahHWftidM8upGoNiAcca8KfA3eIRqRUKt16kIUbvKylDTfzZhgcFW47jaRD
dLEUCWK34hqKhAFAeHHG+GGdE89TvPuoQZeWCflisVKgh+EErRrGQNegoMUEtDwIPCKXTy2UjnDe
+Jm3QK6jSR8wVAnV3wZChZtD07CL/MqJWS1GQnOy19CiyTIvbZ0C2TNEKW1dy7Y/0k5lBGOZk6G0
0WZc7GPhoTSkfHYLXdAJn5o/RR8tnJl9Ypoi39MsrNkCmw8aqtpry81PRHlKiVEJ1WDKKjmPdl0y
Gefye+y0nHQ+Qs8DNiRbxvXdORnLdb1Nsxezvgr9Cx02N7NTo/9uSzM4GhCeErG0VAxtv2vJD6DH
97OzuYsb3MroDMJR6TqcO5HeeOjOlxvMbNWgCuIDbmNB4Gw9487LYCbb/5ou3i6bfKKOXCVO/Vlr
gMHbHWAwzQecuCRsgnjbZ0jAJ372GAzTC4iXt7xMJI5rzzQllqDkp9k48BH0eGVd78Sd7s4v0SWJ
SLkbEIvTWx5hMeeKK3F3R7rmUG8veB28tn/OXkDArY5ETeu95TRKhL/8c3wLwu58WNw+Q+HXbZtl
DCg1Vsj1xJoaNYhfnn7yJjadOZG5zmLrS9Cbu7ZPau2P7XN7X/lPqpr9958HL2LZVb0s6wEXrsJE
2T8ytTiUQaZWZYR7/yGRmwj9amAvj8QfQUO6zmFlyvnJ+bJ8+VAVr7AR7pkh9JkP/MtLbAd37Xti
eFowg/BPXaMJovTJ5c1qhRrXy33faev22KsaTrxCtdde1qXkxxZe9vif/PfGyiJZVF38t0DBwzgl
7ZAT5jS/VGpU1Hq5M/XzjVynW0Pj6wHDVBIMSevhg5kbxqrQAOtKX29cGnybwIHHbEbuyVmI5c4d
B0zdi7GN3J9jn+GRfnBWEiNAuNhBR6VXufmP6t2renYzPgOyIsrYh4H+kLwH/k5lofes5wbe/drs
c9ek6Cb24rMbLsQItR9pA8t8tmEmVp9373+pXKZyEyewxxG+/34PUQcFWGSjnasfhmDDdzCCai3V
rGLHfzSRzoBIpzWT+7maG1LkePMsMQP8aW+mxNh6LF8gETsJRyLM60FHk1khSg6D6BxqlLEZzxoD
0OQ3dr77N3bTtpdcIWt+eIQVMeuiChu3062o/Oex4j1NWcaz6jHFtT6Q7atlRr/DtUFpuy5B5tDl
nkhyQMJGoYsj7sq4FVA6bj0auGDUh9DuDDWqN+wIZBuwO55knjAsYQrXXPjLLjcOzf/STUs9qPGr
upH82szI2Z9yLlHu/T1wBrMhDq2WSoKE5xydZD/WVU53yzLbbZufVEBpuBejL4m8dY856DW8mR8J
OBzEf3W7rGlEA2/m1t+1Gg/Tf6C8rNtudYfdMf5+nvKlnuEnFg+KjT/hPIHtlIs5Bxt6Suxymf/P
fxhwhgZ1ReTmJBmPtNeN7KuMZuJD6Hdws/o9rAigf3BLtfQPx66X8dbrpuGGpPn92CBhKfXvgUka
h1xruAkt8JVT2ird2wOmryIeym43Ho6FI5BC7CqTKNK8r08Anco2TBsmAp7FJcAu0cvVWgm/ntpK
GyqNmYHf+p3VO+x44J4GiBR4kgtdm0LnpDj8eyN9OsV6HI6xNQZyGzg08sYz397EJpF767+A/eJK
M2jlFuyUKGgq5j7msUQM5hUIJrvSGUOMLBsKdVCDHSXuBSTna5B1YUnrfmZmko5aD9ANibTTfVvN
qtvKcKGng3jcQWkFCzEBm0v6tRMSIubV+XB7YShiHeGe2czKtsiqpLxWjeXgDS7aO56aKHnnkXm3
5xZKXI80rp5Dwnjzx3HwEpRlu8IduNVZQwi7AZ2F7XQ1Pp837ydDVXXl7LVo1dzLRoDSD9OyBSVs
hfta/VqoUsuoS6e8lEuF9PdR14NZHMQ1W7yyT7XQWNslrSdUlwMACY8I4LtfvZZiuTGs63j0ilsU
xf1mPgejFix7zsCv07WLht1obU6ILshrHPSoKE7p7X8uMC3NUEshjwr8w6lNCrFzuqMsIZxiFIcv
rRUEuellabdfptSyISTlI6vJgp+7vNOi1UoqGdiv40bGnUsBnlwtuYOrFNm3X1/X5/ZctuhfuJDy
ggCZ6E6ERwLYvBMpu56GOrp0oSI6fUMr4P53mKqjwGfWldLM+l/BdHti2bhQWKqWoy1Uv/oXMsOs
fzViw0ZLoaHJY9tOdRSRnpJ0cGOx7Z6Npy0jzDRCOBKTA5fjKbSCpA5nnFpIoedqt6sjFLdmngK7
ZNYj1vqFFbcrTgX6NWPVUSAgxNL6DMHH3VPVPg74aS179zpFb04uNCuJMlyvSA7hFCghnSobN5g0
48zRlsIUYCX0fMmknxoUKxDBEtmiWF9sXPx3dsfLV00C7ZfZv4UJfhIn628U+wFyiqACJIFWiyhx
ZWxJQKsH//NnhBpZ+DM+s/p6xoF51KX09AVkXNVC6qRy63oZIjFvmA880HNfQyDt0td6AuZeaY+M
NARvm6KDefYCLxlAAQ3bM5Zob2WIeTzBHNNoqy2b1lKvabf4TgrtwcIFB9qZPFSiZ678rF0NkKew
xjGH2aDSicVvxSyu2KXb+u7INnGKiIRKP3gUPncJpxFCn8TKUCk9X1P7jxT/vi6Nr3yCT+okicSM
d7+DjBtx3uHmNyOYnksRpc9Dmd41rOU209kElvqr6jpLaQio2OohE5qCeXARp5bBtTuJtCqFaQch
MROWdvSLyuvPY3vTF8Lzifp05UiuYMT5I9YQuH0YEm7mgSQp3S5oQr07XvwF5B6v9tLqb9ybe7wn
HOKzTtJrYwVnCHpcMacyf/uo2URa+tt/uJMejDZK1DedZgzv7JjWkwaOckPMweN0IQHdIBePKBep
N7T/UM0j8jBmZhqWdWqwNF/cMwpNdBsOHe/BOXINg/BxxsRZ+VANU3dYAcnu26AcJD/sL/ehdlUi
/iu51g4tys9atJF3lrGaaAPO3Z7pvkkuL5qpi5hoATu8q+bDvSR2mW6RTYJSoapwUJwi1VyobO3Q
o8pcxNAsTcfMWstRxDLwVd9e/hYnSwr0SROC9iLLfH/FVRxmMsGGGLwhwg+x7inj6SbftrGEiuAR
wYG4Mep7gTuvUHVrV1aSEOaIbrffLA6EU9RPdWpVvl6D+F1FKZmJ2LyY05z/xsjl5OkluHBcvEds
gboPyJolHu4DjPFvsT6QGVrdTBPKBLuYmBrphRRYMnEiHldK6g68I8crNWBBLFwb9oo37qRxSWO9
/C3YmhqGlQiT/D5yutshzOmcm8tQ+1Fo9K38qKgPiuNHyB03qMBsaR04SiI0w4Biz2cS1mP0T6xg
hDIiOVLqoAZL7vZ46A8MVfbL3ZFL7SYIptyZvBzvjQqE1KXpaZXxaC8m2CGd20nsXoSVKzkiD5Nx
0SpVjyFTuNmqB5++CtG1qsEERJ2Z0RR2g0ArXORqOzuAnNDLLFfTGWHKNR6G2BO263bfUi/m9UUR
x7mLNB7ntHQMgzi52rz6iTaoHMb3PowkVdzGedAzvmjEjRNjL+497X1EgCTB+RJ+pcSaU/+XjJ4L
lD5l1Q0WBLj5ISEER4FasRjzRPIKZPq638JIj+3+9yh+FcyP0YB28YKuiHUAYuLv8BcZ1XWt9CsN
4c6nWFOWNlhp2PoyCh0sO1ZLieQySWaAu20YRTpEExyZ8IS2hBT7JwQEc4Dx7g79Gz9Qh5ZhvD6s
r3HEPgCNvbCNVrVffav65woGDwq+Ei4q2Jm1iPSURqj0Pcuj2E9pN1y0+KQRiI175Pkt6oqRUz9B
82vYj+a9GCPK2jwlZcmqPEPOQjlgPkW3Cb1RydHg/0QPrfyE0k5NCvjPMzT1YR9LJsOX0/4NLxca
onSiBTVHqli/s1Hb7UJwhw9W5b/WfkrRv/hxYaOvbYlZuFJ/P/OPtanfCEiDXl7+jgk8QnN08YRO
Gr/RNyDv9Ptin9EkLEG7yFktV5cJ6Pof8wo9YFDtE4aMW7fLc1Ip4qBVETR6Jk2KGYWZWYw1/4go
YDBEnRvhYn2fUluz6EmhKaR1wr+RVaVacqW7XVX595XiR7xCXJK2OHp8fRst67T7zdyB9GuBIde4
+tq2b/E980f3s2xx19xtlHDbWqgdLRl1sd2jtEpPxF/ScoD0nim4IqdBzWlqy9U0/QBi3tDvLrYX
4WXArmlnSaaAG07RdNBG1rqVYhyoV4ml7//CUMejbkIUEdSPIwg5QSP9TO9SNNEBMZO7taoT0pvD
UaLWJ54xN8zJ8k+P9i+Ohy83yuFf2L0ALZyj/OoW/XGDVMrpf0Tx5omOfR4u+ipZsWeYW70hYr1g
JOFOxzmqo0PpiOXDUyUOA1xsZWvk0q9Bkpgw84hxpLjcmEgWZKeqErnFGuxGSYxFB930mlxGLIaj
pRvvGwV0Z/bwWD+ccwZ6MOPRXsXC6CPfe+dFItp3PelXmPLGgyb8HwVwV5leUBDttfXjf/Pn6vNl
TgdBwrK+dETYQJxcJ8Unr620IEvQ58EFMdMINhFLOf9dJoKsMDBJT0IemdECsxIi1K+1ysUVl1HF
5KXg0eapigVDyIn47yUgsr3JG9Z5YoGPUHTQybr8YqMFqFc5DCHVocHgE9q8oCv8bSj22reaepMm
YW6c8p49ApCecujc/DpTWwiYoiBMPQpHASd1Y4SmOETdpD0Z0OdwtPqCYfsYNqhI7pfcBfhJnjMk
40EVjcFO1XKcT4Yllts7zZ9t1RlE96AL1AH4R/VF/Czlj3UvR8UwVnEidXvW15dj4qKyGSj0ACV4
CM4aXcaH0MUZLybiQJ/OrLtGa7IxUstP7ZCAYgfSjCDsTBpoWkw9xlbKmu9ekmI0vCun9gxxmWDW
qwGRZMguSr5vu3UYmrpZBd6bf/DwRvhjkmHgh07bTeMi38+EaxWyZadla8RdfUfKxvZdQ3xq7e+p
iTqurBNxwZx5L1AqOwXXf2XX9+IUBHHh0dQQV8LBP6XXiq25Vy/qclDyu16JRgSIIBIweIMPCZxG
8S4xIIPjXDIad6hfG1wLQ2V0ViKZLGLRdoK6RusTfIFVK8uAq/huR88nJ9r+EiI26L0vCNlufn/1
NkxisuuSJx2Gii9Oze9C+D10HyhnlZc0eqRmd2hJ5ov3xDHPKeVd0iUNGsxXx6OF7h/48XgxMp7L
XproAhaXrBC3JmjDRSMws7ZM0vIkcoonrlhcUr5whRzW1yxL3WbN55/EWEfZ8X56qAfG4k2unpsn
Dru56UiKON3l3DcsEjzvLrF0DbZ5WdHRY1Kupsgx6vzFB2qOlelWQj2oYJ6zd1KLAi7mC1Frefzn
N9hsLY+p11MDZ9ml7BD+xIc5W7igsi19tF8F27nK6slgKvrFLragEQQCpnkMcDwRksKWI67FHW/4
JKgt4C6c+QbfW/b8MQ5P8bmJLBoqrxWIgMOYLIhiC0syvbdaGQBvJWBFf4BNboPFR4BOlHSQgB2Z
OsxxTUst/VFaZge42Y0dphywol8B93TbEFha/+4Nb/4m7Uxf+HQr72BBhkFHW+k+i2PyqpCVgR6U
qhBEM3a/Y9ZSE8RvCdzNNPszkgRtS4fbv6Oyc7DcispelQJorxraXnQgsrKmvRQXKt7VUI54hxqc
qPElWuqX1aEYC2otOg6xLGL6RgOGw6xZDG+yRv5765q+XfwNHk8HQ6F3bGDTGoykuBcPBeaK+3qm
1BLGdgZdyefmhMEVOLOWmxinNss1qknE++aoimx8p855D/OJaH0yQICT9swmaDT3ptdOcRFAwh24
8RbG7myMevcYcZD6Ww==
`pragma protect end_protected

// 
