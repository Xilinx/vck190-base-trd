/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
l4gSYexUXlM7ifAaBP6t2MLRFhQaRe7Sma+zo2L28DiA8DDFN158h0/DaBr1OsRaQKqTpiBWurc1
Kc+8TD5uaOBbdGAOqQnBtAA+GhRIwIir9IbLuxBMnT/JmOaK4MUYPqvoRzrgYyXFE5yrJmMkU220
b8Arh6+dyt3Bh0bC5r9kA89v3D+ja9uQnY/8oodAq0Q20j5GmOBNL7A1mEvLof/A0UYhDRCv3pRO
FKF8KrYOR3RN8PBeGCM1EFnr+wW3J99nOfKe+v5+if1arByO/0BxWK1JYTBdcxntFYOrk/8juzWe
cyuQA25yLLNZSsEfw7pTdA4YqggvIwnYX+4CfA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="nooMg7GjkDsMTPG3DLODBuXednbZgjpzUjgowzton6E="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5744)
`pragma protect data_block
OIw4y6hn7TeoR9JbrM9EZG93j6zNO5CVH0E+kkHwpSOuqKw5wj0viHtXx0d8bnGqz2fxNpQof4yf
asDO04vTg+bjR0A0xWIRXz7gWUqM3bUgcKM60FbaSQlOKV9tsBPD75ev04QDiNRSkgQHla5eGl/Z
yBvaSCg5N6YU62ckuuNfemTu6ve19uMrtjD1VtviueTiIcifEe5OOJSjS0PSfxH82wRcJFIGprSY
rP945zZ02D+q6LTNxHGjlVr1u/yYba+5jKgyHXhbDh2259HITHLB0cKuBCCPLmUo2a1uhiKhaZW7
6uFNsI/rGIFoA5xIZIbaANTmxmrJkkGrvZiYMWULEi4WMk0I7KwUVbaLlepfORQ1jHTbKJp2VF3U
qGq8Gass9K/TwNTmPA6fn5lFRK/DmtexqfpX68vwjeb/3jkuYmNifCaWeclIZxrNqb7wTklAd8Bd
CN7knvO18aci3ldduvf55hTLTVn2XVh4ZmF8MlOGeclyhMZlydoI8VMC5BOI9pMs+ZH25c3iWnbg
Nuo3m5P/0w7iccX2eKqN7ror5ItMpi5ioDvs5UiCCZRbIOCo53fdnZv4Nusj/rhKnddkCKte7GH0
2A/a2LB5DNn1fRvpz2Lqu4oiuQ87b79Ka6vJHmYamWZzVVuPzL9tOjw3KhmWjTMbPhquQrj0obGa
cz9cnyqd9t8+0kwwxwwcEo7DgoIddK0rRSuezSA2xOYUlT1yneMofhUAk4PVWi3oXp4UdUHC1T9W
VHJjXsjPV/SR7nI88zBUVAr084NTg1lGFAsAXhwRu6OALoBJKIoIo987DVhasIKKg+9D9wUjFSsU
6yeG7i3Hv7ZzmeWeoNWkN6sP4nLyAAG5RbksstGL2rbUk1oMNLuJJsuotW1L0hDEzncKIAT2rRO3
MPSEdQ4/vBlSgDCGcodSzR/qoAXDYWTF4xtetN3rMTABDQbWL1hDfdEjgxIRD8vFBIzPujYVGBzD
ETG808eo8ZIq9vIQaMV5C+GoIJVzFC49ycCdqwap7HAkfWtxnv/ydAclI0bYyCDEHW62JGZlIUTB
AoE2yTP674vGn2oxb1499bZlp8+rYn+zxl2aCg2cRSpGKfgM9efxJH44vX9+K/5F3gfMprYSZBBa
Sl5NxQYjqV9VTtrqZFWehwEztSKzwkH1Av72GzXvbNFHj/GvAkKW+mfjxOqmTZ/TmsfTFOhvn42G
EOF1NehOrGlfTJXLHyJVBlFxsncFrpnK3BfrbCY6JJEXAKll41cy/h8R4kWfsDgsBCAwTwgE9T6z
YXjJqVFvd8obJR5uCF5O4umLCnsNwTdqfMi+X6o42XhmGvjldfmgZqtWcjOS+HARdJW3ZaFd+CwT
6gKqyIsUmEoF82x3+sq7uvtOy63qCvZ+QslBCYCQotvqaAK/YdQ3afcD//mFJ2ySZjhKRarfD1Ow
bWB1U14OHYI5hbXrlbCO9nH1Q9qTyzvFDjx8yTVrmn3rVPatY5F1l/CACXUlvf/BRpx49twl2OUt
Lw2S30JQdofsp8w9/4xVGwaL/shOiPayGsgbj2IWgr4/NLgBAvyNLFvDx5pNMcKupMRXV7AbdzfN
JQJ6RoBn4ZgDeMNdHX+nD2TVizVA6zgT9JY1h/7snRKQ2f/jizJ6Mz4J9qN/bzJWV/FU40FR0ybL
Kuajo4spk3v+lwI04IfWTE8SixWU8aD8VgWdc5HaFjba+3uH8JAunB6AEuj58ZvcsSf5rsNaHEiM
NriQbCWl59TGeP9mfd0VXR7Caamfe0z7Eme6SPhi/B1m4IraAom6GygKW4+FLUndknuHcWr78MNy
5lt/gOOKnK773eUSBAQpzxKo1toUSlIdobPI8ILOChMtLB8ReZHCy0x7n11znzWSkYOUgohxYyro
T8BssIXe2P9MHycImgN5xeJq8SUhc0erPGqnsXsae/QGhyJs//pTIHZlEfd4vRIyPVcR0p4ckWA1
mCxTAWOaUDY3fPlBcp+EHOlos94zgSN6Hx50SaTMHbiKmvtKV/IvhXEAhW66/8dQxlop9WZIUBvp
gSwl4ROBA2Ko+1/sczQ/IXro3hUWM+WMK9eH9zKm8C+mlxnkZSdL8Vgl3m3LdlDeDXDzNVkpbzdO
EE6cSBNnINBOnAbVXA/2aB6Y7/GPcqPpx4XIpcYJcMxXDteUlqdu/f8hWDm0TSbquTroufI1QE7C
PpXCcR+kdeei0eq0fFFkj4T17aJrO8KaaFKznlhdJ9cvkHrIyRMkcjOSraywCfRw0EiGOA5GjWSg
H1x6JQAabdaHSoprNzoeKjxorTQKeDFyJVgp1AOioyAOnBecsknl607LxbjhbdUxCOhFrosxo4hH
czYatHvZpeATMIuZqGutIJsFXYtFlYPIIvrMo0yS+CJITVp/1J9IseY/mDigx7kM21NUBsy2ilX8
zJBzHaW0wU/wp2nfwQuIxB6pAZ42ey/+yDABnBkskNwZewyI2HEEE8NwnWZJc84CXzAxaFjmvBji
OXu9WvPcfMGRKrezBq9a8pbTD2KE8MuXdKj1NI1cC/VtWUBK1YAKSorWS+7/caiM8KieY9oFr8ge
tu301d6nmHsvImO1DkZf16RZ83ojF5EgouMZYj4NwHZNvJs6WokPRag80x5IaSUspgC+Q9ElkpB+
b7fq7WINTNqBsG4tY/irjXlZfhVu9g5rfxt1//Tob4XfMmv2dFVWJOK+SjhBdYETXt76DxDjsVXl
ef/Z6sr670fE1MknnCwTgTRZ6RqJ8Xgj9jtVrfuvwYc1sGJmZmZhkXixevJ8BYUD3ZkUbGSCAxaR
PKPkPNRGfPAvfw28hrxWkOI+qhdFsiEk1d+IU7O4g34/DiVLqqvug20KGCZYvNflbYk4TZUG5Rcw
nwzZ2oCTd+YtrDLRt9kEt38/eRtIT1DCP89Iyxcctdl7CGjbNu+GWEdrGhUpZcrG/3K81vWGZLT0
PjVkzqlt377g1I/A8IfIELVo2gVGjn6d6pX1cN+5K9Fc9Qw2NmZ2mY8Qfzs/tNEVyg4cTS0Oee+H
IL2kmQKQayBuEB65Pu2MxtKmffdVrbr10nSadPK/ThLfPvUpLWoyisM5B7/pjYhTH9Yq5l7SFy3z
/8v6UAcTbqkhxm9aUBD2RsPQgMaJuuEYR0520RoUuoloIHzGJfx307A6D4X0TRuLiYhak0Cqc9lB
2ukI6MVXKe3KX5XOtu/Zw25my7DBxFcqgwPxoYgn35zPhmW1OD9/P0j/fuuRRnvuprKeK3+JyXjz
dlhq9OOauaGU1tAVhMZTVbIqTu8GmKBqqvOufRRIOD1+2jURs/yPOjSwVVuDDkB2ExlscE/yStNZ
JbCivHApHnkafgYQgoa11nSCg6m3rb6NR4x2EI8rwpipxqiJ9ATon0D2LK/CpXsawSUmWjnm2gwQ
frHeFNnL0yX+JDjM6jSwJHRxC4ycM2xffiKKZ+7HYeAZTgCDgQXEKrMa/GX8C6r9lcdzDudJI7iw
Man0omMCumcxb3hmHD7EUTioh+x4Pf3srqymuO2K6qYah9rR2VnYqv2OQqV00HuLTlBdWypNSwNa
2gda8oKDCbgBB+NfcEr2zh7UXv/UoAj8tYoMO5Sp+V+QJCjLQO25IniXDPgvvaz7eiaYGpsMSBQl
U4QXjv5JvldNSmrTODlUq4fFkyH6Wjfe2FGUcke/FD5fQNm0R10nHRZ6KrLR4ApftNb3c6Oy2Yo8
+GV8+NPfkD9U1mvRC3JIw3/7gSkh6r8FyeHPJpZ2bSjY8Rv+o1PbfEMnXiOZtqKK5ZCGK1hknFpb
Lv63qjvodVbSKKjX5jr+HpzlhJg839Bcd5s9CFByMs33D4ZOmu4Y4AiVf5Nfxz9HLV+BTUPBMzRE
IHkMjqd9MR6qG9G5sUUpkgR1KdhQhnCaBRmomnb9Ibw4/Fmw387BhM5qNJ8FDMuPWZNUok0qhZ4A
r5gtI5KKwO0qkgTHKiEOsyq36Fq1BGrAfuZWPUcaC7G4pofmchxpr6gNKQ+0ya7fpUi+zuRxrx7K
FQsXQ2L7CHkLsg5pKue0l0D8SXqSHRP7PeDiNaYZlFqA1Tn5J/zvCQ08f3cTSNhcJUuToSQo77SM
CrYCJ28OrWFYdmRgm0GbvcZe+WM7+kv2TgYcDDNa4lkYRgP+HpRLKaCz9SJtlPw2L1Qij+O1zFeo
3Q59LypKp1HWRD+e7uUOOnPRyhYK3PLX5HJbcd0OQw3ddnZwAXKy9Huv0InJUGjaztXzOICCgxfJ
ug1ZpWwDhov744cERufQjKe8uA5OGFzBdNP+pEBmD1033nnToZ7szIXrae3If0GvGShxoNAiuIQq
YfpvjLrm7LYJqwbZ20PaWJE1W62EWDm7XOvF4WdKJHwS28NI69ZbuP/HqNkHxTyKcw0V1w8qRJL4
hXlgX9xpyi8BTDJAu4F9u1OTk4YPQzbTpgKSuO18OWPDqzyxw0l2gnEBQLhs8FZiTUxQ0zzfQqIC
E9MYgnTZHUcLHlpqJYdmTpav6NP8x9BtuNIzfp3GVt4JwwmMnubWv54fkvEJCa6mVI59h483fSuP
PKcFrnDoP/+0UjHC3naaL8D9tLa0qg2YCwu5zzGxqukhA7Et4JnJRqPWX7QOtwsv1UohG/1F3qIR
ggi6Qyc8/xz8Rcr4Lml8NtM5ob/P4RhCABqfZT1YnaOhJmGiM2RFlbCteqnThhDd6u+sh4k2fpoF
IrAfjPJm4HAhJR3kHUDQdzc78WGNCRKpg8l0rUZhSxW9kl6BSPL+rZsIp3eg+/nPAoFGBDpp9mBl
X0uvPiVMh/g4GimzkZ/u8xBroS7eocgz1mPr/CVHzFNmk2t6UTD3SCNhirqttilI1Mrh+5+s4w2Z
eE+bRA5thFIergISJ8qKyVONeC6i/AAuHkunew/m8AV12W2Qm5mq7kO8fAxTj3eCjgZbVNJH+5zq
hABtXHwMIJNph43LRMMgMWw0aPqmcR9cfk6sAissGdFsH70rCBI6xtrGVQn+tG25CosVvVoAGS52
v2MxOY9RjQU/Py0f0MMTGHcVXcz4llW2NrVBs0ooVcrkN6GYDoAWZMcWY4lQBF948JbF6QgOPisM
z5Kp86jp0mKYRi0b+VqhRVm9LQaJjjNeZXwiUxpIVeYn96eLjJDwslHKZGS5LYhVb4JLherjr3Pi
xLyv7HaRb1XBUCWyxduyAzfZBkUkhnnisJHy4/feUmSFGcvonxGBIyKUr/XqRSKMv0+hSdGHs1eG
5I/IRWxiihi5PrIpkKY5ojcvficn1Z8bQYm1tNAQC6t0cLbHfo4cWfNvLoraqoQLEEbfNC+Jcg21
ydJGRH64KNhuzq/el81fFjxkiSjAKa98xso9EQOBqFqP7eL9k7ZU3BOkLb4obyWSMNDFrmMqwvCo
/5uCj9Abo75LqLBqPq9ROMiTGphalsRZ9waJP5b8wCG+LqUR4yE9IAjExaYXsXkR7syQYWTd4Wjn
UMe90SSNLOSymK2erqw1L+zbf1FZxxPkGghrYYtmzBAYkSnxBO97NYBlg8pYpwwg7XZYTSf8LgVr
CcjCxtW8rdTxeIBZpKXxvYNOe4wXn+VG8Pgz4bHIww5edrsb9FrNflPzHn3b358y52u1k4mJZqkp
aRTKgtujbk4n25L9K59PFWOYGwje7+s2XLQuwKUAQTzEAPQCaVExkD7V8bDtXCAo6gk7VL1AzbDV
6a4ydvxZELi9alzKwaY/leM2IH0WJxBbh2060FA2Tdb6DOJNn2OI5l0qIONB6NUZYy+uzFierxJV
4kK61IysxTUucoDmxkfvVa9oIJzVdS0SdkbjD8uGLGaJ6GjYk/z+/LySyvf1Iu2vLvzjqgZakb4i
cA1/OTxYVusyc6nP+mgDtkb/CxsK+oOLJ6wBH55hanJTEYLhYLWs+v9viqd+iuCnvKCL+gyFDLsM
jPbgI9vRo+OV9oiExIbJwBmromv1zoXM5NQP1BTlg3dkTNH9++SlA8t4s5B1wVkX03h4BVeVXzRj
siTyflE5jma9mCwiKkWj+xpfBJzFmCN/qPZOYkryD+DZjnE6HkOX+Gil6DV+aHrJjqDSwR1WdaRH
/8u6rz+/SVWfU2Dwr8KHDPqovgThPhZeRk7pYSURwF17CQRl0d4FWpQ9qljiWFBvhqec6FlL2oeD
SdUraTprECARF1Xj9jB3CpexV0/6akHywuO7f2tgD5p5roH5Pljh10zAyD9ygg4gQbh8H+pfhMRn
XMhwZLjhwi7pzqKjTdSCz2Jg/3qoPLqLgqN9LADKKkhpZhzhvlR7weYqCSt4eAlBfClahvIEEVHU
N/d/apL3HEBxHNDFYLJhAHyHQixW1cpw8NTg8f+zqtF/gw2QHazNPMJnBwO/Lj46RhIUJTB+vRKi
jAMdqruPx7+EkECy3tb5AAIoeLbg4FhSHj0ljNJPqBGMOhTYiBLUc7ZXh5cETOMHDkvMRryHJpYO
XINDUKdY0mvZeR12h2k1926wKa/+XhZWjf4Pb3W4EWwAEreebJwZoJdkKqBqkcMxQ5fkGMjf8GED
A/awYaplpRH4aNNUCWCNwFl2DUY/MTB3VpdiQj/xLE8vF5e4icqLfG1tSn5L3A5wT1WOmhVNDZP3
6clbQNipBm0d1i1lm5rrusf2+pDdiXcKldLooNp4pv3C/mzysOJ/G6Lgr2fVEgCesG0vTN8RW+GI
C4U7pz3d8LQfSiD0anT59A07wvV3/HX/+wptm1HyaogT3fq0UlW6ZytOIEugzEsOCHhRBtJOpWM8
H6sQTmLX5pIkAUH4SMbcuvrA3WLSaodg4kultqxS7MvRPS0pselNRWKxPQkJGERsmGQOPCfQnq/a
+xOOjJxTtWjTUkh77RqFhatgCSzgByb1HVwRP23Hsi/WVCWdqSRUpPxzuPvdzGNbFiyaoYMxpcos
EdKHXdaZissLafKNO6vABuwNef9IRopwXP9u+uVshbdiGG47RGbqgrAgMKnWG3gx6JKl2Nu+DqSI
pMGKZKRc+XcHwidkYp0MR/Kk8usubkXAcpt1YhMC1J7fdfyAjmCy96ocxuRl6t5SqoWM4D9q33Gy
ujFEfeDVLyWCwsM0Ij1xk5JrbOPfW9BvmfSmyrtoGJae3Tx47ElsrCNXHoc9Zd/+G0nMjnXpa997
tQ765qnyC9VQ7lb0OSe1ihhQw00CfNgfOWtDcV98trh1qS9TogIgI0tcuy8PEJx6zxwZGDpW/O/G
s2IolKdHpb3vg+oXNuI5P0q91fwuTJISjwwn4rr3qqxTWhr2TX1Y6ILsiUxSTXiisv/oMAmKKKjW
L07Bo3aHcCbhQX2knziKfP6nb+KI7HVottPDCmPlNNDT7f1Y9nfsmYuq04RLCp5mOUbN/B7sBwxk
d/iupdePjQ6mNnshf4ISOCv2Bbsouxaq32gGQnr0nggstxSgg2VGt/mXyzK6yikjSzzcb2qgLoFk
4fI0gocHqDoKzM8Q8Q/HcM8mDymwrrhXBLS6yXO+e5sIWz+eBZ44vA1v4KdlRGEQIOXDWMSChxJE
j/OatMPfYdZmV6YKmUWxaC2gSt4YT1V2bj5ZL0DH1q1Gb2Q6r7f2ARSOz0cda+IjoCocvXz26oKv
pxe/FhfOTPjL7LBoBc0ocD/qQ0zQNh53iPsAAhYTHRNDJf1bpMr9HnFF2sk=
`pragma protect end_protected

// 
