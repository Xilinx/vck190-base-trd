/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Fgcvq9yodAEyu7zsWWZ7LwHLqer2uRdIROgj+b6me/wmyj6mu+r4+a1EPBMoGlf2Rxb0wqrGm/yl
7FT0a+0gf6RIUa901Ug60cEq5l3MsNjnNX0EuQ9QHnbWnPHO5sk3W38XYr3s1DoIymcMyzWSb3j7
DAgt+R0iGXGbLJHe2UuAgwrybNhjpWacbybFOYZoLu5Z50wmOHt3p6J+gVbTwfuHK/f+KnS4VtSD
EJxx9+hQNEvkukNe5IcvkATvsJ495o97/SdF6+o/UvTHUZ0m3la3MPtrbbqjxbRc5d/SBaUYwJ/0
DSKgI3IBXs0nO4MGwCQX4Cy0xa1KtNy17Uqy4A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="YyF30NSJW4xBU1bz6CmJ7uDDg1utz4oEiyNQAWYk7H4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1502352)
`pragma protect data_block
3JkMrY1IEAXvStruy6C+3tbJ3jNnihUPe6ljwKZ2ndLjBQkndXEvL6OVkXT81QL0jDCXXcb4sHMs
X7DbJ0JBOsvxw7VR+QSytPxxIa+8fywUmFL3abV728c/12585Yklv9MAC6qFi0fbRLpbDrIxaReX
H9Tbf0dS6adbYE6SRLdvmJy/ehXmWT1M7F/DaHtZp6ON0pHUSy21dUUrmBSZvia2iA9cicU194wC
gLuYjeD3Q1/2fgfsuSedU/XtvcOwE7WsTdZrphIInZerxOwku66wqqmxLZTvnh+bfBySSMHaSMr8
fUOG1W8w88ER1d+GfmFjt7+HmKuvNr4giRSmdCwc2JS/bzrs3+6pyfhFNVlk5s1D+OzqQozHzMxr
EeNJXXrrSCmZJauPs9sp/6gJXIdXMRDUhllUyxNciF1voiR+AP/Pkc2VxkJi1/Gf/6e+UBW/GStc
nBllmyYDt1BPzUOiHF/gnILpfCi29wBTkRGiJH4k5kIM/v1YQRoPJW7AZDsbJO6Fr5tAfaBXwJbG
L8uuk3ZiXTauYQzVuYn5W8DiQRuMEIJhd1HPh0hGXMvv2/8Pfd3udKPk+WJu5bz1Fs3+g1NBIVLU
F3y+UHkrwGu9ZnA/J1FgU+zjlcOe/9SFfHyICEovzleqpBDwINCbgB0sYND+3xFW7H8DRtjbdzAJ
3acJEwr9+E8KyVhBnUM+BNeNa3x7w2nAWOUVs2lmuoMVHerD/BgeJJALSyuSI+QYkOvrs8Wua5X3
xUurF73zQiAdYTbVzPfErlKQXREZpgtl0ySJ/14g3FvZDV5RelTVtz3O8z4ePdwMb31MaqVIllO8
8w0dsUL1VdtzhHiShqRRK4qJWfiFap7BMy+No6PPp7TQd3fdu9CxAK6UJcaZrkZNtPRBeFr/wJtX
ee0gfUFsQUocz7+IXLPXAmpSxymQSF9VvoWwre5H5ZOVI+uvLMpl7TNKetdJCrExuoHSjGmcRO87
llkkUWIkTnMTN9jiEvJcjqnhqqMRRFyk0OqplTQB/RAVWWnDzD4G5RBwrxrxDSf5laBdT91+I8VF
oQND+1gQI4Wyd2ZEC10FjKGImHAy/KWzwt0M0X+qCLASIc/oSZdWaTjMvlkGdIdNCTsaiFUWbVsr
M4xomxAAPV9w9Pf6xTCgYdVScOWv2grjanure0HTCAJWqNq0CzininXZ58+oBCr7MDjfCkwJQ3ft
KUN+O3FwxLm19OESPAVRSzeBR02Q+fAAUxBjMAzRIY7M3OnzW8ofpW+7kmjTPxTMO3tlO3m9knFX
HSwUhm556r3Kl+msXbuWXL9kziqfnN7xe22PdqfE528ZpiGXQPFJ7D5/szJ7ZcE5A2vAT3i3B/dO
dLuWyR66ug+9iVxf5SIGMDBAzoT6KFUQabFtIiE6kvohJ7AswisHj5mYFAHySJBNaEGEPl7QOqQ8
UKo1qGD9y+FJZBWFMBPFQR8+35YqbHOZl+AWl+kNyslRtL/Kp4JugTgBXmmrrs03O9Dx3KmDrPdf
lGhdVgzvAADmPd+XAjYpSPn5QwPYLn9NuIyTsRmLgIwGzMGHQWIP4qkv3jqa4uA/iU7X9Wpmn9V4
BQhIAmKcoUovRjESnx6QmsRQdO4vtrEtroWzcWU+PX6q3M8Ojtg4bssPEqqKsGB/CCQk9XXbc49R
cvdDqZ2KbZmj9EDvVfNdKTKUCVUmj3XwxX5h5YFDyqdtIeO3lqy1sqRkyqtCAGnskekBDeBn2tBu
txYvoWBxWada1eHaqnvZP1eh00rn1m/VXF4R+e/lHrakg1EqYnGCFWEW2xgPgbYRf9VJjZiFJ5l6
ibi/RDBomkPU3r9uX7Vo4VlgYkrzo3Elxalv5TLrn4cWHxmWSVzjrjkfbbteIqd5P3HbZa00hCYq
kvxE0btgny4Lgr3UMS6OU7akmRcVT5t65Ucg19DPJVMwTfjBRdnHv+i7OqAOK9Pn831NQjgbb3LE
Wdhmw4fX46Y47mA/eqcu4O0G7EgGJWG7qC4u9RXKLjO6AQYEsfhAvHzAzwut2h+wkpOEhM2nkgzQ
yYGwu6UQKTe6zPi3+58JaYStfmItl095NP6WhBgjPz6q3yYnijYa8tHc0duq/ITb2Cb/wlrB1o/6
ckZFGQc84ZkseD4+ZUAStO9pcBoveicdr4IHw/Lp+l2teM0Nuaoqs16jfY8vCk+3Ag8vhPrTLm8S
95nWeEzpNrhVrrArpQve4uvrdaQqh9hafxuSAwXSAsfcR/B3bgV0tgPsygS8QYkW8KyjJz1rFnBd
KYArG7YfFNncFJW9zYWZNepPUm/2SGNoBq3ejxeUBmkXYNnGIh1Qe/kaa2BgpGspOLus7MWdt1ay
4kWIndCNBbaC/oJdsVDFClov5+/Zq5WGDFoyGDVtqAZT1GExTj+pDgocZOIaAVJIMlbv4UIV1lgq
MtnWlhQOjClfTsPOgoJUzX60v/sIp+hqWjSgaluJz8wq4s0Sk/48n6N2Hg99EIcA+3pra3Br6Cak
GiFFzcCPen9rMLhMAqkCo81LvJa0xfiwRF50zLeggueCEmjdZNbc8Kjz1xnCbg5ng9QvrrhtWiWi
Am9vcZJZS7+0XAiKg+9StJ23cvzSllPpsCev5ry7mUFhhd+ZPScJbDhm64eT3ZinQqwG1uwsBLxh
zlrqB4/wp6KFCs1bHqhltgDPNVjtTLv9ETsnnfgEfajwUl/U5fOAlxseDtcqOVuDzUZaUQGWeHS9
Naor5UdWDWQd9As86/Ux1L7z7T+RsG95jwLMuQMwgG0DmN0uXHeR2hKu1wochWCeDtXu16E0aTxh
ChleeY7A1kX9UeU1MVUaCXmkua8GrUVggd01BdfczXYZI2gls8HbTFMJ/66nWaPCEerXCSzGr4OF
OtYG01hzWd2NgorWCvckpmIxyICEJeQSHnw+xJTicT50RNrj/GI9d7zyiOMNwjw3/316w78veFA9
sDorqz3eDpG/eazZJ6h8lCZ3IJ1hS+0km/CX2iDSf8LOApXWwei9YEJ2E8tQjpFnbsgxwkd5ZU15
3HwPTC5a0el/6IWbTfmEp1L8Oki9ogJyl5Q9NZUNK4OqAbGF7pFahQvbPTLBEDhLKxCZV9KwKSGQ
H0+nz0fqTBjxrvR/WntqxUtF3A9nuYwSPHyfEjaDorGSq37OUp+dnvld58rfW8P/cp0dVeB6Ku1k
F2IDKdDSneMa3w3TGK1fZr6iEVJULiXBJEKGZORPWVPgJygT23RcTEBGCyvc7kWMki3s5ao6jNuj
GYw7zBWt9127rDTlC1DPixbg+Nuf2wSnKC39Eejbe/P66BEVB0pINuigzWN3OqNGrXa8+ab0GaPH
iIv3+WwwUfk6JqtMaTuZoPqybQy+Yd83YlGRCbl6xGEc1wSC9OuOrya/TSfLeK+ttWwm5VmghRu4
kVhVHrVE8renTZ7iC5RKwfdqIX6hbadKbzWqkHJ3T/pO4nLf+9HUo6Q8gLmfrvyt+FWRumGnLqEF
AW1C0EN0GbeMtCPS93zvOt++VWXR2Jy7lePsgc2WaCQueGq7EE4FUhYNAY5xjdzplC5XCoRcTjHN
pmXXtl7a0h2eNDM8amd73CVT8XmD3ZvPZUOVfHuiAEnFFD3FmlDlx2uNA/xpZhvM+joKmp5gWDj0
3JKem+njP6OGG3+56OKH4hGggorsFObx4X3MlPdRd0XRPS22pXNs6lvnm0W5SZTwkA7oFNQ1uEu6
17ZDekPQfDsR7hxQ0sw3GTXUZ7/4ITEO2FBX+iSuEC6H2To6CoFqyxxFSgTUPqfoPkt/RmQaHcx0
9TRiiuSwyy8RaKKCy35rwuY3S9DVXY/qwgoR1ryvZ+fQkPaQg0JuPCCV5pEdv/p635H4Li1FqtLv
Q0oRTqWCGXsHcpYkLPX85+SUb7BEmxy4ZV4XSsxv2Lkbqq39W4XNA+I2vVP980V0c8GXaC6GTww4
k/UqmPvIMg9GrkSZjrtPF+Jo+9F9kKd8HB/wVYWX8Y+XkbZVczT3OUNtOsbWi26E5inlFetgzVv1
6ireaDhL5+aYn1Z4DSl7eY5LUBUhhdNl9RuSoNvvVOFoN8n7kVd0Z8ha7XYRcvAzEflkFvr510Wf
zkCzfJ4+XOq1UjC6MXKYApe+dpaQ5tsMcW8yYENFIaYIbQfI5ylY74heKzVGadz/iySu7gqGh1xb
aM0bSw6//fLIRNgwRH3h7tfjka7cwBG5EfDF6m8bZkVyTIbWoFgmKpZoJTU1cuAMLD+y1vzzJRcO
RUwLkmL+H+zrWtRhatd1REQeZP4HgqJCXU9Ku7B9Wyek+r9BYZ9yYfydxlj+1LHp1HHkzMefqVSj
QHfA3F111sbTGW3x12BEcQinjXocz9ThI0nWfBFiCQqCGZSziGa3nfwN3gHj8vTb/7F7HH5wObOk
/Tl6v76e139QXKhTfLtDMtmvf/SVVxpf+BqwL1sfJkgNatUpHKonWT90rJPZi7TjNsRcuy62STfr
rNtF+zQb7zARuMoUaIqUTpaf5f39Y+8x4CVKAzNOB9j75EnTPRi73o4Lp/jsGefEiZDKVoeLpSuF
Z1N9itKywtE8qiEFQGvABxhySaPCY/QisqrW99qRXYPOg1Brk4dwWUIwjrFnuxKWFDWn91RREguv
qTfq1gXoTANPctWvRLHfpXRgLPbVT6nXV4JH6MrX6Y4SCpjzeT8EnoW3CFpTjnf8pYlJuP6gIhXN
DE0OEqkm/gUy5i2QXrbXgV+n2V8jHKoxO10joLQpiU+xjk5PoIrtwLwMfaGgKLDHkDISabd0G3Xp
z4LBaWsaDTQZbRrhb2zX3lOUfIxQac5Igu+qLTUqDu8jegbEFj7P4yRYWrCLcQjDQHKqbgTeh9PE
jmqUxBa6ysTfONJ3z8XfyxIfUX0bd463LN72reprNHUwjWOmXwb7HHz4g86OMDYslaIlCoXgbLuq
ZzFpSlpSzt75UUZWd/NkSkWNr8YnVRffyPBGp+hIjRoUqHjroLmKyawEdh3/ZqY6tdrw5K8XexfC
3auaJGdWffcJWP9BdK6wpLx97k9gp1S2E9QdlOD9uJifaI/of/OMe9Q+HscagzmgjXSwx6PSU4IC
Jdgz4GorpKieDJrtQaZiolWuBw1o/pKTtWKPcaZRcIa4s+ys44/R5TmuFrAHBoc1AdYzwO8fth/Y
e9TmlHkVL8duYyzpSk/Ru2gOtWB/KhQb5sTXVm2/vYZmhX116m7G3ilBfMDCXdRU5v3EtoegmpC5
rwkyofJPf/PAEXBJQgb/h6VAEWLsxGPa/bkJRyqLRzr22NVMoepO1Fi32DikNpUHhjKavudrpQuP
m+0W/tnmbl0NsnlipdwboCcawVZ0Erm8W+mQL27EaJcDSsqH4rXmx9KSHW7TXPJ2/bvnxBftjgR9
SjRf7kxZ7NZc6cR3GryuEtb3+HBQAXQRSZaVSJCvz1WpCiA6ETwN0devKks9y5+Ub44GCkanhs/J
gHOAjUCTDQnXfOv/BZELWRrL+Kg14SJgX/o4aLxYdaath17rFmLWycSX7Oz4VBFf9z6fZHwY5Q3T
f/rIJtjhZXlRj2DwtDBnvIeeJDckJpnlmLhqX4ohvO4hSnAXHT7DFoCVFYk5utgYQ1LdC5EoYQM8
Ys4tM0cNHLbSQAzAKLCqh/0pGxS5HPgxxLbxlYL2Y5L32hnhZn4OeVL0M8Qkv/Ei1pso+rLn285M
maPudGB9Ea+ovg/N8l8lYjhpqbbbatebl2H0BD2VDE2Ri4acujNjAAVqH82TfzP+3zhDW0Pbx70k
wn3VP6HbmsXB5JNwQPZZb+NEtKSZ4jrW3Fm+iIpzzi3UtANZMeIIg3psr7sl2GTvtDPAD3yqDSfw
K15fcA+pR5SHuXogxD/ZzJcmRAuJIFPDMpH1sAyfvjvhXd81Ye8cXv/DSfKloRsBwzPCQmlnwPNn
/PYyZzXDYrKVgV8E10zzv3R/wDz2635fdAQO+1hdpY5t5fG+8A4DoVuiDfALKK7eC1vmoUFmVJ/o
CA4hAKCriASKqxYwuFvdE74V1vWv8okr0ZIBoDvK4nTRmnbrFHy3ACG+igSv/usy5TLqnP1J/kex
uK6cJKMjTMJa52rJPWv4Qlr9sjKJB6bwC3AWG2OIAKYpzQaSTipjFmhjg3euXKgHte/vpFR692KY
VclF2gvDNNyDAc0Wq36tXYi2NYFG7EJFpns8rMsVj532jxB9rykPyD7I4/nRVJdVg1Xfkd0fxVwO
7YvWSsPw7fDIz81IJFI5ws+UR++1lPT6L0OKT3bPnDZKNkLD42otNDKLl6IYnzjHl/vAv9sxCXdA
mP7safM7CLvsCqvqBGqp1lpJrFwR/CrpBC4d96vy9gKOa4n+DOAwtNZfZz8I7Gj9uikU3Io3prYo
QTAtRBNCi4HYfOlBGhfK4774de3gLZygGbXGC7mdTtEpGaVVHYTL14mpjlrrENkcyhI4d+AthhOx
2R+sulrKQiFPfwNsGOs5LNbaXG2UqFTp3nfEGFwxP4VWIxBD7hNKLkI+E8a+H60d6xPeJajG7Gov
nd5yheEReYyG1dr0kO+qUIzHsb/mCDT8SBY5MDBTt63gk3gqyh3lOJRU118jMXQQtiaMQC0epsSY
rdUhMG/WFHQ24GQoZLrpXXfl5FHqiBG7AMU0R0CH49IoEaGDGAuaST6PB4yl6RUguN5cqSCqkOKK
tqM55jZvWyJ4DddiP2cTgJlRovN1STJY2uYkh7LgKvHmak1TKwtRcXGs1e/kXTOdjcBO+Yz4tF15
Iik3qqQhaBa+H5Y4FnELFpOSTrm1kmJZlIROOBAyjoH2pNZL6ePLEVSJ0aeAJl7/i16s8mCenEaW
PaUvalYRl0wHWdwhseIJXCKycgD1nsBLWF5+o+ConVUqGAa5XqsA6r/JbNMz7GrURDAVXAfhKuym
PcwQgkjxSDvX0gWacmUWRwcCosnznJL2Zenm+ft4+x2nN91PcXuPQEAkqC394ufbHIUwvBjGH1xX
iNo402NoZgPKAN+Ad/LG0uIevthZO84/YiXxCEwVIYNjHzksZmRipAGt/+8iZnLdVjA/zCDqBlYt
1iCq/NItpuUyPOLY6T1fh+l5zc6unWR+X4Vx5HlFr42fWAwk1kNOAfZdG7D+9gXIkxZOMeJZEIkP
DJ0VUO0LF2bcaKf3vdpe1DOFqi4DfrhwIwXOAYV/znAe89rNXXfzYaD+y/5+FR+S8YCtqIaa53lf
bq7SdDkzq9nIBND4TKEcct0pmrfDc88mqcdg5qSNY5gRxb+ceETq6Bnaxrzexr35yyQvKdBi0vWa
+RqgeB7xlUxI+yNKbyyW5A2RsOzf/wK8tAQY5xuyCL3DfjPaFZmZ3tWMKFkGkA+z8u1nvm/ZKb4c
JIY2XLPi/rWDYAllsQ0YfoP1f3hZsD2e6sGetzkYXBhU+5KF72V4t9+gc0XUp7OttFsmFNSUs6bR
RC4Jb26FiYJXSg69zz0JmI9gqVoTS5I2hTmk7j1XD73NtEbQ1ZSX1KX96vHb6tqR98ZDBvlx+jPF
m+y69JdeAAzagxaXRVm4SosfnYw6nZGJCQ673iJv71yuT51sBJYAwfI14kytXoqTDf/mOSYV9vWf
xWMbYi015Tu8B2UYAyZDv5/PLgS3SUfRXQKk5ztWdNzQHKBtDsmz1e4sBV99zHHwDvfX5ueOaoAL
qKiO3g7FhsPB6dLmZqifuAHZMsmBJ1Xt+Z0s3G43lAaiw+NS1hMjFrEY2fkGlh3rH6fnw+NLhEWy
6+rjQB7A4Fex+NOQezfcqFW6FDq9L4acM5hn1JnLQoynlUs9aSdXLW3WDeCc6AlJ+EpfmQjz3pLH
/uXjwZB5yDsgpR1Tq1weQgCbXekOb13iNVqQ6fbOih8KJ+WGaDnuVrq2vnPYCw2b6xZkbHCCsvCf
lIoiJtHpG2ylvusiaSbJm5yetHBTh4M8xE68vUOHw4luOYTGE8QowlZgr1hmxHYKKG/YeTQKNBFx
0ShJRVqw7vJJ6XtPDvB1JWyoICV7EImkbzywmlAI46NGNtFeZU6RuFluohxuj/nNCQnaEyYUdoPL
PuGTKc6oaGwtDWB+7Wjk1FiB6njdnSGCvPTqtidVpUNZAYwklTx3weV8PC1+v7IeaVQCRkwJS8/4
2enxtUy8qWx966yrY8nDw2ZDD39wp7XUBtoUXwkvyuaBLipXQWaAhTH5mnO8Unryfnzlg5a60q1s
qNW9y6+Se/gdOtAGi1lJm6+hLdJgP0DBL0SZuVi0V/5MAu3dP8bvh+THPQXh9J0TrGiHaSWRgrho
WU9t6vG10WanOX+tTF/dQI6IWRnPYRRg+LNi7HNHRFY5jS0ka5Dw5tVO4c9TKWg8GOdSeoq+j7rc
UoQSTGyn0JegNc7rdGgUVGxe84AXrjp/Ac5+WTk+wraRw9XtG5WcPpEC6LmODhTY0o/aFRfWf8qM
iDGlyWhOw5mkrehr+nvXpIb2Xt4L9xgOzm4+CPHXdY7mhPb2QP5mHWN9kYUFxq9bkWN/pxk27UP7
8XZDot+jeCbxNZZBaS/n8k10hTokxvdoSTvS7DCuatw9hTf4Aiu6iQjQAfbi9VsJj51zlhpAL22g
5yDXxLsQwllrKQrI+DXWF0oRvo1ZOxCCA9nU5OY/ebJPFhB/NnFvMu+mDdD4lFcmxpoMtEZ8WHdG
2zxSUgS37jV2qGrAYTdMVsL+jEmN9mPsQoIs0DhVT/g/AoN1Pt7C28r/UtbF2vUNHhRqagkbHCJg
ZDaeOXQ2xouVAIbWPTgpaKHGRxHFwZlzP0cskBNYwOKVAT1ANlHnM5Er0TMqVou6tm1J3hMuSuiy
VzMlp3YIOri+drxzJ5kjot6jJrCkReVpMfXVU/VmiLMXmAIYPeuw0dKccd3lTMpqLzUSni38coYw
6uKsrKbOizCLQFk+al2S0K3rHo1xdPpJrafwj14woA3WwZRbv7hFS8uCdAgBUH3G9/LQ816uQb6n
BTwm6slwmHfZZCnE1aP5rTSRlEHtOAJTv094us/QhAVxGcFsgRXiJ+kO3skbDHeKUP5Jmc+1tWIY
tW/ykHGRWJ7jg3nW38c55e09hUFs80hdVxjvsYofs4hUYCBpiMBGtYiHREzdh6c9K9hN57QRFKDS
El6bMdgxLF5ri//67T6u82yGKdvilcyCD8rwQW3OOfE+7ziig+Bbd7g96OyyV0L5MA/DTTiwtfYm
YYFZvVKdz9LMiaDb92ApxTdItPnLCQBkfMzjicfVrzjvMX5tiB0EqWlBIPT6jWMFFtgDBWYAuZe+
UG2hvQtn1uLB46SRYpF/zmK1jKpda/4p1yq9ecJgQ4b4QVSoyh2q7nysZgQQa1Lozwurty0qQXQz
+UN38oCflTNTBktXSMMDt9xHpndpsBW+/IIarPo1pF/pHShaSeU+iBqeZc9ddNEyT53Iz2z8+FiA
Pswp6TDkhCgztL8jdMOefhd/DsHSKDh1HxsZjmBdnuMJ+VAuOPJJTOev5RSQxjL1WrwNvHz/CN9w
P/uI0whjby+kSoIAvQBQGDNhlsgJ41X+a0RBkpRI44WpbLa0m1TzLYkMJrLYayEWx5BcY9N2s/K5
nlmLUTcYuEMjyGrNjH+FIA8eHvKCQB+XIuPFjgcb5jhe1cXssA3fUwzbVawqQ0bkRbzpfywoOEqJ
/1Wih96QetNu+dfNeiwRjeX9wFoT8gVt+C4SBNWSYOd2R1mPga09aOcIYWFFDU1jf3d9BEj7Lo6f
LeynxZ3QST2giSReJSm69mMvcIJgERxZFgd3D0vytNuwEMsWjOI4T0EVQGGQkiC9l1hzbYGFfGRn
/sRqFfZzLGAK3IBwjM2H0yB2grs2mJRhVwrtwbVBLFocjX52RcSNBz9BcpraTGIF1CYuueQ/5kc8
M4SmLXJa20d/O9jFj3Iu3VYtlDuAeY5pjG5YRJUvTAQqo8JEqdzF1QnefQ+Kvd0H0tJjgzvKkdQq
LaSTPywjdfXVaXat4eyrB9HtjZAThNC8SDbmwJLCY6GzQYiI9VmzIugKP9HFPK88oWB7L0VgTAsq
sQt3nu+FsRmi+JqNVmFp9Y+UHrndcjELTNec7k/MEkXqucMiz12ex3sUh2byrHEz3h58Ud17j369
zTKPMeEZiopBYN8R2BO3RHy/zHI5vOANeiw1hCHDnDjVX38w/jPgS6oM5Z/Kpweh2kKCyOZTXOMl
Tp/SRg1p4bH4IHmkhuNhNm0aVbqm5iT448pazPx+JIGQcG2kXt7heKdVwiOk7F4whmZrIKp9BHQl
grw5trxmyMrB0T7dZ42wdSWiOk05/rEJQu0zRCB0FqVizFknx49Wiru2Vn9C/S1LgQN/f5aSXRf4
eVx4aN6BBbAkDrKIFth1tM70VlMtulm/9HRBZLMXaHoKTbjpXVkVO34RN2PhxHMOoe1jagqefcF9
KPao+Xq7fLEX3Z/bipRxx17WHeNKbgpJvgxyexdZT8SJa1CzUP18MQn/0EuYfIicx/BCcDdQJKpD
omcTM7kI6TxWMPd04z6FCp+UPqZcxSmpfYsYJ4ppkzh8TIyYQAFSirID5uLaonL154qEGrYCn0Ko
8e8G6G2S6zETf/Op2+WWq+RN7pcn9yNJv/Rvk4ER5kMNDQ89kGS7gRE4ffw3MVpDwgOGiQkxuJAd
f3mvHgQvff211F8ToeXHtOqJwOXL5git+P402rbWlFiuGJZo8I4m8wzazOLM6yW1hw50NZAFwdaX
oeo3NZZi7NXEmJVbTwze5/ZjWQdnwnpmkQMtK5bBaykEyY8Ai/qD+ciVjhzvhUZ/8LzboYev4r8i
55ImvLRFrt+zrtJzreyumG2i17r+YZZ2oz1vQ6nPVFtqbRBlxWF/VXSKgXqa1gbkA6Uo/Oxj8Mov
6qQ6RFYYZ/a7KVGQ1tN+our3XKR17ubJULZqLO1rT2OWSu4817Vk7YTO9y6KfBuzA/grrMqinP5a
Er78u5fXs/3Ol+ETYoTcyI6xWOBGaLLNpNNKPdERfj1z5c18J/wgcLgcVwuGUvktgNWiYRFrtUbF
SNHUHNAotAi1CDkrZLFZyQrQks7GMjUzspuxJYaJRBw38t/+jpoBB4g5SIE7/40wsiMQfUyIcVac
2tYiHVp8hnFgFYQIfjVhg9IEpaQOFwyRSbe0ucA6MthtQeKRr1ZyUBm4gvzD84XkllCws5lTpXTB
IdfFNDa4gD0sc4i3v4RTwBDODcVFrEBQzhh4rVvr9xO7NQS0lwvVJWSss+iR/i0eqnrkNwyPqbhj
mAU675yMy2skOVpdnlFFT7VlAYLx7nEa/HXv5+TEqf/y10cMrMpvok5795fpK6xwo3HK0sFPvbub
fzNx7sETRO/mVetty2d3pNWlS41iasn893R8AgtxzK7t7K6k3pDU/VM0+CV4pus6WLOBvB1b4aNw
rL++3Ql9+s56RwtISPWpEKPhhdGG+VDj/Up2nLXV8Uo6dnXriUfFLpuN5l4gYpLtPB/CmZCh0X7x
8wX2X3KV/pR5bDCy/4gQTxAkZUQPluMCYO1QUt34UG+xwe/x2Iybg9GRNgoYETsQZmEro8m5EMc7
/3jPZrF88rSt4/hxRhfSuAxBA/BoQga1u0XsOQYmHqOK2bzw4780qvB52caJeR8FZW65t4z8J5UW
nTaf7zYt7hp/ous+ahuxc5UbTiBh397SAGvxNUSNvHFdxWE2RiheafssyK4GB9CqTt+TLl3ikOoI
5j1wug9D6BHkiaMosR8nIfPyOEYrrF82i2NhCiH8DH0YSCIX6xOpL2c1fMBOGadys/E3X1DpDOky
Qnau9ksZJV23iYrlrsm+3EuR4H31o2Ri0Re5GzUH9iPyJ3CLM5+6raf92f035l5irP/JrrGzp7ZY
fY9nOoj3dvOdN6UgqBDntSl4h5Fb9R0vIoUINCTCkSE+qOOT3Ghc+MW1R5MMVnsDh0Dljy1pvSG+
NMenejfAOizoz/KeCIh1c6iDx94wf/A+TLWfpqHixIerNi10Gf8n4XGQdH59d8wkBa5D8/4k+DCt
OTarzI28sShkcZfZWJ5YvneQXDUkTGeh2jVjId52Eyp+cR0R/PTWoBhjHaxXbVlR07aoSTJT/fyX
dVrLp1+cWN/HTAAtaLjdsat3ojh8egGAIc5VEqlzdoExgDoV7Wllbz0QKdleZBn771VYThDpaaZy
FG11FLgOGWEssgFnm0w88U8i3ACE2FxXShMcBoWCmlql/+QsfmQm7CduD7azYcxzNHAX3QFRrIkf
yX7fUou46Y+G67baEki6pllwM95phKJlPTuG1k3dub/nZ8kX7byhl6Wi5Cezz4H2iat1TbaRV//e
LZl65N/obT5ody2lwNLFCwXpE/RqO6uzgTNINT8YQWYjKU8zNSTNVKGkZBRB3DDLiN0mM+DW+8po
rcF8u62Xmddg0vJkGgOYpo/OeVDcc6jxDNcUHoegzBSJenHXJEaT3nQKZO6lQZ6pmJhl6/JJCUHv
frkbAW3Vuc+VgUJpxlj7k2gugqzFdu0KWjRMno+pI7/ZNGoqDxQtwUbgX3th5ayBOdTg1b6hauxW
qQe/KzinFMCDxJ0uXAx6Ruqbheu1oqOWd9JBeIi5L9JQQaxVz417Cs9MJ5HIiwH4eI2YPsbYSie4
C4af1a4nDXY7yV8MRL40A56pdj3dHPGQ+UliV//IhZAHjmi+cjKqrTP4kl2SIGWL5O0L5W4PfGi/
eoK1q5rf/ulamHdz9QsSTyrQ9G4JIHbG5jbNlL4EVUYbI1wTjrKVRpP+qkAwx0A4+ccB7MJrmi7a
+estzO6YU51lyHpArisGQBMToEJlH8TuGOWVFFcMDs1kck0zaoXNhsldnOMh7OcuqwfmjvvfVmuU
+Cmjl5rDh6qs6LKfu0Q9LBsVTROhGnpXiq9zOmeFhfrK7pcwnFgtoiL3L3CZBP8nIYcXsbcluTIV
WFIbregYimgw81Yv4CANVMk1VBcHMoq2Yprq0aLXqE3P2w0do10esa7aWpS7/tazZKUIjPSCg20E
RVEzsJeu2iKFaO1EDNCUb17tQCRtM3MSmen2WWPaAEMP7L4wTV/3GndIJAr/dXDDXpXzKTWxW69S
BZvNmanc6kyQA+xJokKH30cx2UyY4P7O+dfJr/3ufQx0IiOFSCGddv9cZEN/S6scsqNQjfact9D/
mfBKb6T8D+kY4v3UYoaffF+bvxgNBNmE+chJ5HyRFdlKjxm/Jy+3OfATXDh5Wj+yrCj3rG7rai1A
rcy7xgIEjGdQ7gNBLHIQyJu/6OM74teR2j3TqrlNMlN2LvVwd3U2VWU51WwhZ8e77JyhHghdQLvg
rAlmZmUu8CiPQbTZfGm4hzBaVHrpyEVNrfyxoc91hiayxzKwk5Y4NIzinlSw+cvOxKhF80u9zpVr
xN6+xKmOdtYnNGsqNQaKNCxMLBJrzOZQT4texSxZtP5qeLH++8S9J73KUVHi4zrnO4Dko3ocLBfx
ZL9vvd14cF/D8OuDgXXvCs6R+aQpVQZI5hDhvPpXnxhzOz25i0ZboJIOY6qoS7b6pDadhPCK3tHH
D+N7qzePi0bnaWJOpHY4RFvoqonhXBGbNXFa1UZNerba1kpmuX2+irUlF2a16fXS023pdYX8iQr9
mOkVcWaXij4p3UzOWD9MeLacYPL4DjoI63eCl62+wTFyUd6wFIHHUMI4PrWlI7LNLvdMwdhgbMa6
hhX5eez9ECDTo99+0o+hv4wvGVs1aVu6XiCl4AqbFBJz25WJMJrfjofk5G/VOuRkIkHFvlhcvB8P
DyDdombT1kgeZWe6PDSMIdpsI4KIlhrfgSw0X7hhY96ACD2UoWeE5UlJ6K9oTL2bEF9EIrBwLf+L
w8XdKQdRW4M8FRsGjbnN+NWiMpWOg1kgo9w8o2qWeUX+MPwgPUzpznuArPyJlRkNygU1Y1sN2DzJ
sea4uJnkW7zOHRMz0v0AFxcknHeCJ2oObD1HnGuwC5Dl0GHGoZkEhUHSYg/pc7TVP88oJuzDU2lt
iQLOGz2Gpv/i7TuHktM7nuVMmSO3KPGEHNfcezaj9PGvZySlz0dycAHGSYBQ1zZY8Fyh2pq0oCUK
FJUpxT3+j9Ict+PgDNJL7+TvKXNxMIdwHuhAKcKmgN+eXKKwP6Vp+hutm8ULuGrvTvG9a63VuJNW
PbFm8uX5zUz37vSh7bjcg5MkRK4HuSOx7o35SmJm1mwLSb7+zoYmldq60/MCMCtgCJILw7o1Cwxm
6Fs3kD8Jt6YakvNZBr55K+Z8F7aO6rh147VDqXO4ql5Y/04119i/1GhUHJhhEuwG9mvhqjV4EYj3
MsIMSaRYXYoIiuCxIk8Jc8ZPRjcJPs2vAYXunjE4E6jwxM0sfXsdljhhVCkQAJVi6XJEu3ntyzgo
Lh1Wstkll6uHAHZuKJlFqc6gJVK/LqVllrmJppwIBe+Y8FKGemhtj1b6pUWw/EqozYXglE14ShWu
m1R93i4NH0pTwVPgEH0bJwH5Qvj+N0hThgUY5qsDjftc7mWgkAikBjSZa9+Zv3NiteNSw1C01W6Z
J3DC45I/qOZPYZrt+muatblZnYfWGheZzOOqeoogFobWAnnQle/3oKgaS0kQ69gLfwS6oVOcl9UU
nKw1P9PzMwsjphqlAcXGa8OgkGN9jz9hVC9/4MAXS7C1NdbKcqYWVaHiyJFIYT5I2WT0CUBvSNtX
WPKiYIAcaoC9ZaDkpCGPkenai+8+dyglx6gjsU7uA9S0XT8E+q8l3jZnN2JYrW29iejkImW2BiSP
/Y0POuQp4Yca3+sLLKjlh24CiNSsANz6al4Q+jKHQyExRjCdgORzXH0Y9t7x8zpMnUQdk7pn8aOF
myAtCOdQuW+ux8Ti5E5HGtqTRyGA7N7+ljYXbxQRvgAQvfzHyzYPv4Gk5Wdui4KvBvj88IKRBLAN
JbKW2vwrWk4cJuUkZICFBQhwhZV74YTil0IbXxv1iFoqgv2XcgJo0kX4DJPNEN5ejTkBl4t3hAod
M/5fjzLzp6A21q8zOrgXl8zQkssVZ07CIrBiFHI1r8NzxZHlRt0zwS23dvue4ZL2Mjicr9OTdGGY
z+f5qJtgre0Wc1HKu/+jou7FiHydC010GP7klEN3kpHNQ/tqYk83Shgy0rgWxObLdaIUjl1r8yPm
gYslYzstIN+0AINrKGoEvzmSXPq0YZnP2T/gFxmx5GTyM4ylv/0oOLs47xERpZUKNeVzoWkyAPPv
bdJBPJH3YK6x4U01yloW8tjZHc/+F0MPlWtoUdDr6c2FkawnWZkhrVIH6mVzS4VmKOKpJthhE2zt
8jjiWmif/Orrv/ZxHQv3UPy9Mj+3xtzOHigsVLeGTnqP7spdNd+/84WfzzSwq2b0X8wTa9LyElpc
B1MYwCEbh3PH/yXBs/pYTpTVQA+weG2QuN4dbg2RcheMka6BHilPRK8jMwW1JAjjFe43GD+E9unc
1oeHP8vXSnYpAe+OBUKpY9TAAAqSwFyg/HwEWRgmqq6g4rG7vTrxWqFOjjrz7udvJ+IUgYTwnZ2h
Ugy9ES+HgY9xlZbhkSkhm64nUgPC0mQd8YSZdNk/+c9kPLNB5GiDpKaGzoXTh0yBGCzZvQkJ+SfM
MvKWe7xuf7PPFzWLLkuUyN4Reo9dWNUa0pLtIe5dCXjewVUjWiWcQCSR9Ebo8ZO0PvAvGZqlkYpP
SqY6A+9wqf2Pogb2U1/glTTfy1FDTmgLCKZlGSShfe3oTlWNhmgA/IMZuhFcBjWylEXohQk5BYDF
FykyhhZnfENpnKvJ9yzJIh4oGXVrfvUn/qv2R+daIdnk4veO8cCGNf/p5puWdl6gJm9RjboI+rT1
KnbQbLM8dFXb4TJ/NcAiLFpPLj76l4i8UKQzUr7KMFnVb9ZrslMOQG7E+YGoLpPweAwdtznO6Tqf
GnzQxvYj6NrKnM8z3myjrjjYtBUAIlmgmsOW7Zng/CMnuj4aUnXDLGAVVp17VNtU3WrE+jDpEFAC
vn+LAE39nfnZMWL0vhnfrKEgnhZ54XGnqcc4XWKrb2ZkVSjbuBxyHP3j4vF3aI3MrB+jb24CMoxy
Dst5ZohcWaqpfD4P+heLF2mJDpkP4Y2hMo9Vd2BWWzYytg5xzHX1pL46gKpDspaBISuHzPoMXvsK
kYiTQUhsXYwmBEXzqGVVsbyWD+FnA/2vc2+jSRJ+Or5QX999k0vAs/iZL98Twkqvw9PCUbbFdcc2
PWmOe8C46zT2yc/CbrxRHNQXczyKQaZhvqUz8iSJWg5hgBKSrP8kmI4xU9a9hvA5U5A6DGALsT6u
eg5Xc93MSKrieo5njTZlGLswUb1KmctNt0K3yqBoA5tBGC8Oa/LbxyyF5AhSs/UYGC0BympGK9eE
XQbRS7OJvEHzlmuDeFtwzJOr80XeyxpkWn6viHUEZOgXzaFFGSQRuQ8ycjjLiOR9HTAqdIIURUAs
rugX1/E2JRknSPQXjYB4uC1EZ0iq51qcfSiLsrgM5CfRREtM9xxP1F3BTgnbWg8uEZhNn3kU06ec
Apqzprb5aZjKr5v1efMciYgeuPtVytS52Asdltll461jWNCm4WFIDFBln4/WZn2TOFMWUknYt23N
hVPlhYLP8zTuWyR6wHCTVxnCOAavFhgdX1Ra2dvS7/WkJQ3YG1zTDk7bUfoQiS1lX8vf1ar+m0k6
2BfT6qM4OMbvHJAb5++TXLN/6bX67ZHiyddXi0vWyrqLi1jcKb8SbbnB6O7ru5Mepcg9WLgvC7pp
wIKNd9ITXPeNc2M/OoDBOD+49WYTXSzZJoCflPjPoO9cTzqmcuATQv6IffJoUSWghphxdE+9/VYK
IAl0Mvhe9ouQ57By4gESN6SqvSIanL2fQ3x3z0f/dvFa6iHDpLKpbMLHj/hojTObvg/xWwFuc+1p
/X1WO6gFmQR1pQqGzl4q2UVN81k3GDcGI/hRe+pilhE2GleooFygt9Tl5lBOeJb2U0RN8sekMPNv
jpm0fpz9V6jX96qZK4JH+t17W2gmOYvB7pXcIT24lNLFmQHXFSIji5eYORFJHIvn4JRgerVWVEtH
UUO+hNpLot94qbP+76ct2ibKVYPqtHaHN4mTm70fvpgMMMZ1O++7CaasQbcN/8rw+v5LX5QYiFVh
rv9A3k1AUwqFzeWBVtKXM334rFcmQq8Wk9+R4Br/q1AZYN6Ejh/R6XKwm7eXbk+vQzxpymBuqgvy
2X3jsvpdtiCOJIqi1/OQRzatUSsx69psR/nyETbxTVaMy5NSxzVdEtU7xzsJgYEnbXmVOKzequS7
YXkNdQ2jasdRZmifjhhQRUU+hqL6O6dtRHCsDuuXj8WLYD6SRjR9pqMyf+gt6Q3NNUwEmfy2UY6W
WxETTKeXYeGivr6mqswajtu/5wGE5WdWXf2KNBaF27oKZ2eyWMaqTTtx+DlAPbURSJqxEnpJbO39
j6/AVrOLxTbZJ6IH4Q3y3Xq3X5zZxpyNQx9vGa2C+se1rfvpmfMl1yOXCpY2l2zpF0vLXXxGbJNG
IDJbLb+YQaMrXGdy7E5Ynv6LVQ1UEltB3pywTLIC4dYq98g97zSBB7jb5vo1VNaEWuxBYGOHyejh
+geijIU7AMKMBeVGIAOWp3vgucTfoa84BqFxxAI9WpT9iXb5asN0oH20hNbLHGkwefYDDh3cAe+3
LG7gNcVZfpLctn7PJxaKXxgLQ29kSuyUjzfi9au6wf2+9b7N1HdzilbpCaUtYfjv9YOfK3pXnF6B
zEXpeaExr85e8E7BNg91gpMT09HVlXHDwHW0HJ7bi0CIboY3z5FealKoYT/H6YpEFUQ8Z6cfK4Qw
LB6rNuVHmSH433DwF14g1upaqupOjuaSz8EGXyPj81+KeOFQjj7NIlpzk96lPCMI0mKT1hPEvyMC
Q4iKWU4/jyd7uVgrJSmZg8v4ptF85ZlM/iicPMMwjiXTax1MFQVlorrOi+/V8JrGSmpgnnKnYOXa
9q/7hy8XFn2cO2wjeBVCSaB+ebLHSro3XJ0iM+Y/GXKR994HSmmG4nUSpDOFmGRHCOxg7M0Uxo0y
uqZOlYZm/AK0VtG5G2IJE4IenL/JZCnPTz/n1jhu/2HwSKfHkgoXOjT7lv8qhKWYkfyT5FihTxvH
WNdchvUzRi7+3A7VZS8qcuFNVDbJYYuKEWiEY+S0ZdFRrFh3/j8N40+pWK+GOkGCDxCdQLvv1dTT
u88bBaQE4bOk3v3O7D8aZL2K7NLSVYX6aT9mxKK0K1pNKjVWVM54ml2zK4xTsbDg/OhBfHVRluh1
IoQTwAGBwVTNf89Pg3noeGzFI2bsO8hggIRt3bi7UK12UJ9R1V5WuUwmLR4VptUlAbCQPi24BYgr
1OGGualR3SCW9eY7ia5iyeMmxgHb2fCqTQGjDDCyutZIKKvYtbJs6Lpst8S5XEjfQKo0vcByMh/R
oRA5hAIP4q0fnm358i7vWAGk7i+V2aaAcWR5MoWtfqN9OlfCvvoIVWzb2I1O19ZCSgDAkruC+iHF
rbf0aauKatLYd9At/V3N4A6iDzrfQmpZBVcKCHWEV1RveDarqV+GbG4b37XQoYKk8u00OPtwcXs3
egNOOguUUQbqiH7J4i2HFAlQ64quWTgQlZdb0laAT8EWKktsPPNo19/aNnVU6rL2FCp8YQRvw6bU
Tvl1rsp1g/RGBbetfGO3mw4eY02O5usvEYtwZBXxc7knP+YJJIDsL9fJGLl4bwPQjScWNauGO93L
ncRKTOeMOG6ZI0zufTua3lThYJaWSsbbv5tGBTcw6TzQmzpMAVtRlN73AXunT7A4amjTuxzUB7U2
7ZB4aziptuzei89glOnxYcPRoetzs82aJI8d7GU+JxaOPVIo7loQV+qKbtbJU8d1iJTPH9j7Azs9
qigbW0aV3xfUBn/oFKVHlsrmgYR+3kG3aRvXONK/CKt/LF499ep30Ry/URDburHzigaP5kMDj3LT
u4IF4n7RNvQ5urHj4PBwe4cns9Il6Lzl0w6iCGshyzY6Xd9tiqpS150bwrjzWOx7B4k4wHuBLBTH
ATo7in+iEyY+3FGXAgrI9QHMcAn/cl4veEWW40nCIv1RJyi6iyHLFslxklnxHDK4FKzSEruImeYT
sFye+MYgFKLMouf9i5WxVc31vDj2u7nqjpuNobZIu0tdHOlrEyyechANEgLp51/y8wpzFsR9WzEu
4UU6vZ/Fc2tch9FiQCUqOM6fVcbIUVbNIPZrsOtJTZ1tRd1SxU2m72UmmCq7W/Yr0X5G+ESja5wh
F2N22HCkiAQrtHCmhN9q/SRb5r9ZL3l3XVAcjGc3WXS1fWSd3jw2wna/D7ByAY/fwVL/D83LqyJP
foswspKXEoNyTCkdLQX+72yPvgh5tr/5CCuuF7yHWUWtlbE1ZTubsqVF+mNipSBNlHq+ii3mibIA
TDDrUyp0hbO9noOs7F5mWWUXKiZg4EHBpn4RFpavwdLw05Y/PlWb4z7ykEmBAuXpgSDFk8qsrVLr
pCuW0sjFpIht1GxUON4DBNjziw2n/1YBfUdipAGwl3ppjAZrTMtAUpxDsgD0pD9nYXIc7/vo11v/
YGL63x7enSte8JiN/KY+04PzwiM7QLXPb778xEqBS8mL9FcW1lxqPjQZQ/SsXTwVU0JKVIvqp5Rr
2QDkN4+XbyTNTXrbhMy/K/H8xGfZloP5LDWIfIPoZJfzdJOwvtDXfhnec4wBD2Ww+/FLiHAYQmVr
Nn5QyYd/9a2YnLqGjgFOctZiuNtaQ6PDTOgvBr8OWOECFwcQlDXswbfsXrLTs/A4Lnh2L7dtMCVI
1OJ+mxICyRw4NHJCvNGp3sAx+Kbv6fEKV6q+yRB8H0TWzv3SakBLunJevBG7EY3QpUaF+SIS0bFV
MqEI8OrTJQq63+j7EmLpS8a+Z+ubwLJjzTooC08qPf3uCXTfCYoGRulCIwOKgfdbuIpqJ9lmzITP
TaKRvGWylfvt+AOivdrgyPoqTPtB9lFieyxspchWnBL6JWiNaBNyO1tKN7VPePSAe3i+HV6LLQWe
A9Mzk79oTwDFchkVdJR17n6Pmq1jGHAc7cjFKOsgUXWdmZw/A01mWxnHr79jgJFgIQMe0yW9Yq9J
njE5OJNGMsrl5O2iFc4zjqdXg8LHMY+YjKMu8PgaKNaQwgtTMFntzOsExIiLJZ204QsaOuHdFera
m1XhGbv8YNhewghKgweW3i5qJt5Mg7Ak8+J2f+tG1WpV2vIrieNtQOQVQuZuSzr1wcNUQwvQPAlX
POQ3J8Dt7uIGLVPB6qHaCzzVJkDMXTcM6ga/TSsy5l+NGgWGI/wDsmxejcofhCxLaZxyNC+1ehT5
4tUNtlGKkbfS4qvea+kgIuHk9uVUnlLEIsJxe5NUNjHmc5Q/ywiqjIPP+wszMOjxIWiVWCFOW16O
VpaHAZwXV9u0KWCxGwy9wHg3i7mHxOuB/9956uf2Qf1/yrSpO28tmIqHsY5n90iAv179A9sBw96X
0AMB17RT/3cchLBiMbmmaU2Fv2uoMMfdxGoCXAWLEbvRDOCcStS6iXjip2NVPNgwIlrI7ymsK3hc
aWpxjR/C0sO9J4rWzX34H4B29mIa52JLtPn9/rrQVaemLgbZgu4F4SacDT8NX3ntFBTkkyelanyF
W0DshFRSxVAc6TeBAq3IP9/ExdkxGhCklKv6QT4p8WWiC0MYLk3f5o1CqLHUjQQqOeAQ+9La3PmH
s8bvyFZJNcECCQKC9j8nWszPaAXkenQET5Eu6rWyscmNExpNqT68nAssyVIcG32fKr/t1fwzcapo
E6lw3EDWyIJWx67xw5r2XfziQcIZuHyVyQ4vifxumr4MTZJCvAWZpxCfPv7sXKTwjm6s4KW7W3gu
jAjN5ADMr4xm++O+sWc/osGihWqYKdPuxm+SpyYd9BsxRmTDrC+Ibt2dWus+PKgtj09QFn8s1V64
t/w+4A0yqDSjE3Wt3s9cH5htDThrEtZ8duLuEykEh6GmWrsZa4mnq2I4PHChchlRfoiVmrBRxOGY
laEmbqTxnZczmRwk+fNGZPrh8yAz76l3WCal3HdiHPSS7tCPk9VuPAywqtUFwmV51UZFvueEhpD2
zePOfDTVuIoTVn9LqUrGynJh2p2iEHL3XucRU4dkDEmkUtw5ppYxehawIp0+pSBswiqEndlXjMuh
S8tEsO+r2voN5N92tdx0IMTpGuBEoOF3LfsskdxrBSPDpbe6iX2bzm2Z0cqXpRY1Mx3fNr3Umt2+
0iPLXwr0N2Ep1L/zZAKd9liCn/o8SKz8Zxtw8tQYrqRyFu9HNmhi/972gJdyi0kfys845Xf+FT/D
Ii8pqR1RVkWBiBwuNf0ROadoUMSLtgzQCH/lckr03iPGSo1GP8wn1smmF9ZSCmTWXwcTIlOpqkVa
BsA4CnmY79032fJEMwYJiNpgGesyPiDJhw8+PQt7dAFqja1kSICLDbCrOiWcnYw7NquvQVl8Q1k2
g2B2Hvtp91BHai9/kXuAJpzIJ/ZqtHGqoNJwMnsyFbn5UR21ov5GFdj958/6nXpJfCNUru3NiRWa
t7HTL0gFIV8hAGbbA0tqQhQ1hCwmfF43GOeOIQVlq8XMPiIzEGAgmaxjdLQ7e9PVuJ+UMMvc9NXi
4Dd4IFwTsdbHNSmLdGvm55ukTAhu1815qNpicoWJrFrn7VL8O9pUPXmEvGv1Uaw7K7Gq18DTS2dU
uulAO2qisWa6Xe130M7pesYG480VAtxO2rdJSjj/eJIYOCtqJuBrl8c6GTzdNnCXqj9LXt31S8pN
9kcFPLyhKixA+NGEehTrXrgu+/j3ZcJGffWVZKtlJoYKPiU2Xh/Znqug8wRcyG21SjfXnlND/FWv
oT6HFtLGvmqw7L8zP/PHd6lFQV4fR9JfZ9aaUtZhbC+357ygo1eDWuh+HDuBMfcFm8vGSMwhO6Ot
SnlE+iDVoRZCSbdK7SieBCQs6vOvRmJs1GgpC3GbMHOlqmZw7VyDUdrm896Eoe19gkH2PI47LRL4
200Hil1RGBZGfvHFpW79gJv5NVh0vNALoiQ4d12GpHGzDGdduQKuKGcvcMmKTy4EVcu5PTP9AQfO
St4ESEFAmFOuD8UdgL7trSn1c51RwLbmBuzOkNWhxnCPgrZC90KkpZUD5W4ki1AraXUS+2PV1Gha
5/G0B0rtQufYSrO1zRg0wlFKnFftRyfIk3MQe44S3kJrK94o5N8iKsyfQCIpl2SL+Rtbz1MPuWb2
1C8F1A3onOwVXKMN9ErCzOvXLVf1zEgCEGw6ywKqp34tL/FOBrFZTxNRmahTB8n6Vm4DyJl9NYVv
1HeJeScKtsF3KNpxTflzOVO1id5aH8SzrSWouRIl3d/8gYY8lRlmgEfT5nt0TtWM2Z2MY1cMZuSZ
BjhlDv3jNz+6tCCLv+aBFGxvc2/FrQabnobf/B0K4G+LIfizFPlKVTXVzODYH6Bm/RKUmMIShOb0
FkCXZ5Uie4ON7yr0+rj7tJU4zuEJIZpRUBgeqK2cgNSwgD3RSCS+BiDnwpHzsPCgoIxC9TAhS7rw
ZDqy/BCq526ufueC8hnC4nXNjUr+GNmBgF+xkz+SD7swl6dx3X1WC/ejn4K5o+CaULeCGeODF76q
rRwqmIChvrACKgI4ZoeL+GxEA7Nkk7VbljPxy2swL6FK3lyt0d+3aw25zlp+zrBTMNQgrXknbJ9E
PnOt/CiYo81yGdI7iDfWXE/5hHhNIcgU/4aeaUVyLzH9aDNDUFH/koWMFduZIGqUnqemlL1dVjDC
Lpl2ro13uAmGk9GlRzNFDlq3zborMP08089fktz6mix/zFI+arB2jQoNveMdPpiuf0KWrpZM51yD
FMXOTQDF3QladdNTVjzfIyQ5hL87YEQu5IITyyfzhyeqcGSeA5oH0Dnurmmr/ZC9J5I/ZMg/qChu
KVfNtVCqFp2Wk6FUdRQwcR1glQkTv6o5wbFPaVuppj3QqWc240OMksR1mWip4UAN50Heh+faJX4w
87zbJjcGrxWuADSF3Z0XtC1qfmqGprnE7uDAxT9VPF5va68wXD7n2P4dJiWqUg4OL0VW8f4C64kE
64+D8xCabJLWoX1fPf0iRbPG1BPTS09tE3XRJPCMUVTinnZACHiDo6vZSRkt7RwkhZ7k4fVZPFAn
AJtZ/a0LjvOm9nNInR64d+RbKwgVmm4kNX0xEppE1XZOTFKTXbmCHBUViy0/7UVZ7/fSjYL67kzf
1CltacJ7p3re+YwBaZBnZ9A+Y8mCiGkCdFcWbOM1f4eZKS2xbDNOWsBPbOXdjCSM88fc4p5duXY4
NqKdlWdMtiUBUR4J0Htyj5jt0FZMyzSZelaHb3MJTTD7eyL7dht2atovmXdGr6VWV5eo0eynFT2s
4Iem5xEb4ASmUIwkC2FLHkGnY4XZ9wNDIO2KbrkE0J71sP87bTgzZ7m6H7oiEAwTtcxo1czWI2F3
ZeJm+cMqGvo+pODpdKkrC282Ih6YlFRlMmUskZA2PUsbMGRmNc6A2dfm9Y6cenBLRggYvJfiN2iq
mkZNPoLePSlPxF5a34RsRWLM07cJqy5pVcu94exBboXLRf1QLTOq02AmGBpsOuQaCyI5kolCamxY
F4HRT+dtVls/iBKgCW2TAGGP5LLR4E5Eo0q1XS/anlxgrJHTB3Trk12iY6IybY0f3ZEXaPOqHIgT
DMLH6noxqUqoPqE0vGQy0MQ+6D5v9A0NP9/5uiAzx0ADdkXpQl/lAj2YAQWyFTOvMuL3iQyGyMri
c9+JcNW5S0tU9VNYQ4mRTg9JjQx4q15tKb6hvMIlxAkXs2IyeN/b9gPLC8OyEhnnP2nbZhfwCNIr
mq3lZpl36bfVmPt340DE/LT+kpYVitN3UB1UstJ1OcMcXiOHBDgHkQyKwdG6Oa2H/xyG2EPMO7Xl
qy6Za0pQcVOzX2Om0LkilDzlDHkZhqvsETkjN0FQW1bGRUx6e9TXsOUVlPep2zZGGpxkhBk4y/pn
qgedGTCXEJLR/n3bpyn3fMmrt/RHCB7nWuR1hj81birlBaec3SsyO9PaMYc9GtgGJAGzaOrcKQRx
bUq2GkHM1oADViMnzE2G0E6vL+P3uZOvIw9iK96KrNU3lu4m8cLyOjeyf+k8KtdfLUb6zJPSR+rp
+p999U5oiupPp4Ljwl78j+pL+4NDbxGWA7gGrdoTrIlTfTzGMlo9kHgJ08woqbnomhcZBl1TSKBv
mJRtuztYHWUskc+LtuK5CWZuW94F93/vGq57EvlpiKUxSsPlvrXI+J5bjtP0QenQg/KQCL6GUbX9
4ghjvPubZeURNvtYkCniz4EXXd2E+X5s+BpMOZQjmWVLIFMeLJ2AKxp3Xj3+VOVJTtdvrH+nqN9f
sr7uZriyxwrQTG1Sp8DKHq+xR7k4g0nfGKDNRJ0/i6DFJzYD2wwLnvIwdiki+tyV3fZtFfkmvsMc
hNy+vUCGR2VoF6OrQgBg14EonRZFyptl5rUUHfqJeSlNSo0qKMHWEHZPiBa9p3og6eUAO3W/H1Mj
YJ55ZcB/PtkaAWZ8CS/JAEAH9Cq7XT8C7B1QiVWUcpEbPiLHxx3nw9woJELpQX+iEgaozVZLL0HU
C6VQHSW/yjc3u+7ha/86WgO0Na7nXE37tJ94XL9T1yOlM4BGyiOL2BRyCSSgxRCiEH2WqTjBYf9s
VX68cOVuvEiaV/047pEkILuA4aO7kFgNYZe72bQm/iQ8j3SlrBoaVYwZQWWh5KKkHYmlOUxFz1kw
ImeqF4guE4LyZBSjhSNvyFOGRZ/QEsMpvhWRQO7a4U0kLGqVaNJoIKZtTigDWe0w2Rj3+Al5HzHo
EyTzs+sW09dsjQXVYfkgt2EGJYBaZgcu3j75A6P18zx5UxDK4hfdQHeJ26EzEwkc1O4MUbskSksf
t4iQocUP7NeXBycFgJrVOAejbaX0cJNRn4+a3Pb1BEkbb44t00GwloVRrGJsJTca/0ZzQCXs4r++
aPWNqQGT/OjOYZtwsYnZ4a9QHryeYIiVs7/xPqQ6n1TxYx6+NnN9JuaAV8P2A0RjjYMD4P6zmweI
li9Gmz0jXt/JnIFK9i3XkCLr6ruXQwS6OeM1zrEXJ+W0ATf5og5ESnN/Nvt9xyJ2XrvbR3DBI3pu
ctHn5MHX4QOwHOgGnitE1yHiukaSeAjRDkrX9qkoS4fbThIPlKX5J477eR5zmkj1jTZned/sGt+s
kHSnGNPCT/5DG1MGRuz2lQAHCkKaOgIXWsEFlmGMjCaFBYWlyEtN2HssHKlWSyac7ARdvAVrRVY5
iEE39l5ZwzSy0SY6LbG2xJLfvbNs5v7bHVlBdar7oxCN1R+OeMhcZq9g3MTSTQM6D5ITSha8EJwa
Sg6YkQ7Z0/PZcUuJ94WIl9BmsHypooPdvDdNKJOzxkGrPAuDKJy0XAm0sgRaA2+P07uhP4UGRYSS
/yFNmf6b/NrFuyC/aCV9/ch/HuUAFXxznzH4tgwxFrOTuX9xRkq0sA+KyT69SH3yeoyTFqP0tXfv
j6nOKWjI3EjNcriTb36/y26YBdfh+LuoeSAXpTGl+BI3SwOHKeigA3DGkavQ9pHeLLWwyTtMscVS
jYs6hLogWjfFXSJ/u4NrnQgIUTXu3+yg8aZOfWE7u39GPmdo9jw6M0FtYJXfrY4iJrz+2FC00uVE
MOoiJx6PFnAsqOXcb28dnHsJ3bbUWsx3g5NZjGfSh2SUlg9bvTkdhOroU0loaxpgTDS3lI0xc67F
Trw/49Yfq8bCesEjof87/Tu9MJHBgTRMTYGiqEFEcdgxSeTuR5/9Nj6/enbN6LSWeaF9EHXqc4oq
RdL5H2eBlnuJEjqfLta3Jq9ej5EzBLkofoaFH24IgC1SakrXgqaPVy6PcuC5vR8S1ung0IXpKh5f
zV5jiJZro7S2871+D4qgOEui/OJU94imf9ARX4vwLPZa3EGvbxYDVJ0vk7DM5OUn8KqMjSxxQ7kV
qCAd9uJ4dXnYmzlhzcUNga98bZY/W442zbqmahPWMZr6rciIt03B/ZzM0JKTB6+4J6YcvqjJKjGA
SKd5caBSyvpg0o28xZC+4gYVa1gyLiqOUAlwVVq15/7aSY2Wp4yohOoW6IelAWkMP2H0hvjL5oxS
aivlbxjWqSN4/TkTtRQrCKG1LtRlUnhwKn2ISUavCN5LbAnoDijBWDSvVtc32Z28YSWXrHXFPi5/
2n93nj42XzI2RgYXRfum3li4qR/PP4gvO7+/a+ejh3JkIM3f8dBWUiNZuuP0TQDwFny+avO4SkPL
oaxoeC4NQTfQu3L37ogUBMFuv27wcuQvAtq8hj9tKgBTk62U/6YVkr5LxH1Ibgj7RDgHmcq0FZ9Z
FY5cz1EQy3bpp7MftKO0g65UnTFxLOFnqBJtocr0sLU09Ee2rfqYhlxIZOgtND6ifmU46yAowQlb
k/0Zawkc/VfVz4RNSupzWWFl2RgYiraHKSEyXcGh4F8N5OclZ93nfKRvb2wX5yk/VAg0J+nX/3Zo
VW3Ho8yUq2/a7Ek0tNdyZ2S7TS0Slyz9bB1qk1B1OQ40npFU+3Rq4XK6Fy03DsFSEdQzYZhV634B
C+cWfZaRSR5+p6j8FvRYanmpl07Wl9NIIOi2TOW0Pexlfpg3J9ZOfC6n111+3tcUIoq1M5tPQcbn
Sl7IKxH3ohNkqkcQHuYwiIHFPNiOFZVuiEya/MU1OTJ7j9UxHIOJIijBYNJIPto2kgqkP7TR3Ke9
m4D3ZvE0XlygUjuTGxHLLmV5i5m5Lwo0RRWtmfjKYLUd7FvKjrLNW5nSiFvTniBPQnyavBqMn9cL
kbcc81miSbZyPGs3BN6Y/+fxSpmIQ/SWXD0G1FqNlQepsx9jG3i4rojpi0iduK7LtBjCdEJakb+i
KxAObiqUkZ4iu2ZndKabx3EwEMnJdMoMgOw5xy1Ythde1JoWZR5Fxi/MDBOfm+rGbhh7xOrAnN7D
B4LkIOI6GNZ9/NBFnu9unpMrdQbqiYc4ykIh5eoU+S/IZlblLrE3s3BB5coL8DZ6ej83f/A0dxBq
17eME0pPnqKyemcoI8ZfXKsmOvYogpogwQw6PkXlBKoS2YGyKKTvl9YzC9qJX7CceNHk0qloKr6M
wm6p8foe+WzogPYP9V6KusuIcD2WN1UWjkEimg72eKCOHnele6+KryTA17s6AGk6KCJtokIxhDED
PhwpCHiwmGfcg59hPXXsQfZX0m4hGjX4WCJRYEXJNZb/27DQk7ShIPocQ52vcW/7s60OBD+xj60X
13fqMfti60eSEVI/5E8HlvKl5CuI4iu/zOLbG7YSiT0LLkgmi3hPoGdrr0cJ1ESgsZ0qqst53NQp
5/yPrnOX6eSQXnvSHUsimSamu6JET8iJF5xbyX4PJ9l3YhQrk1R2PC+tKU3lRUTEhqQTMGJNsyJn
Gs1mFujq/v94dM89cdzSXU72YwZnCaqPNOINLh1a9E+npSd9+hTY1Ct8/JIq+e+A7pQweaW0gMni
5RcBfmFPJnVLGcsDFnofpJt7agqZ8w46YLudurImSJ318IKcieStFRlVoSh7tGbn2kfmI1AW+4EQ
tRlLCH7VOFeoazW3rc5l3SAfqX2GwyWFh3FCvfq2jxV8XbbxdScaHQJrZ0ffJP/15ij5/jrsGatR
phsU+jhIKfCJ64Ule13qflotbyBFiP3kf6BQYU9a9WBQH6fdZNbST8Jt1ZgcNgHfybafBGUPnQyR
jK0AGGMZBJXbhvRaZ6aFMq012JGMxdsMxlyrfRuKTlel3Khs9LAdYmzpRVPAjtf2l6Q8+dOqjr/o
Oehb+yfl+5vUrO2tbJlgWFVTur1t2nG4FLoBusSNkngRJgOu5oKGMEs/qfbshXahzPPeKxw1sPO+
QDlSNFDfyQOzi9+VZCp55vd471BSmZZrrZ8gfHtT93zCGHtg3LwHXXocgKJMO4KUlQ0EOSA51pZ4
4LnHcr0F+1oIBD/2A/errWfcph+N7RsRO8jNRzvZ3FPktqOStGBsVEEqQRDpVCaZinkLoLmbBQxz
amMF0goHKw9cZFgI1/YNITquQFvvljZ0m8/XSec5AlYKmvGG4DBB7LHhEhrLNEgQ8TJsYwyMona6
82rKpIoor/RHrANKpJVFvMjujGCNkhLro0NgF4k/gAtPZm9suah5sgVFrhOBG5Ns98T0A9l2Fra0
UqQhgOuJhDHBKw5yrG94s91ZD4rxgoX4pDzBfJYGtX6KUilGVwo3NCdLoSXXLWdGkQUmEA0/88I7
rfYHqgnmZqBfYvx5d89zH5qBEKprlXFyqExE0VtRnsIIbOtsa+3+uyfYGsuEqTv714t/OM6NYOzx
EyoW+FzPL2gCYZq87Z9TWhF2+kLR/CqDeNMRTD8tJRuYFH1uxKP4o5nP/HFN2HGsaskmWhvZAiH7
X0nZ9GgSxv9hzWzINkp2PlCXgcBz7EzzMWFzfd/nPmYq9yJHroUbNSTm5DBm/SzcBrhhNcZ4EEu9
Gx+MpaE6bbSS/cAQVr1yrc8ZhF6ml0GVYU13at7zMRglq9EjcrsyUzgHndqYjtw541vy/tTysjCQ
GbW+HEveQEAmeGbnUK0mNlj66O+jNoNmradz7nn+6rUH5tFelkr4NQw1m3Ai4cIIcmurztxWBvWR
K8I6D/96O6PBV5TZwK2jXVGD1A+Z/49PY5UF+/DR3+PDAOmwJqS+g+ndt2lunWkf1IWlsDeuJMbg
Z9DW/L2+WAvUFY8KZR3P0RKQVz2FQ4Qjlh9Ik+5kKNqM2Sh3j6jdCf02f+4kHiBiOOvpKaYYjFnc
kMMNaKJN+XHSeu+rfCeIYxrVI73+2afQ0Tv3QGFWGrTtBPQrOZhcAOeaINfXyiGJ6XrPn4SWyKfX
QK9UkzJJvrwiP/18/uRGf7mrvF49BSHjwr+WjRC4Adhx4E5JVETSQ45q7T/TP73kt5EFY/RnkJfn
bFyM32eRYt4q8+PtuuXwWOQElo1Elur6KhdkUy6/pFmKztuZldPZ9xTNeygHnLoobn7ylg0SjGQK
t6TyRip94aoFbLH3vzJFoGmZF0jaVNAHE963aXndntppd7IEBuIYZRW8FYJqlYIGT7BBoiNr71/S
Z4KcE1+eXhRu5vE6PooxbfHACzncJX1lFkO920eLsT/w2vAwq9Vxo81YT1PIbec1BkzRjrvx/+VU
gs8eopQVGJ/QUpJuKL4+MRuLO5Y4rjngyfZgPVYFbac8SYpder9mSxWbtE96TPD0/Yjy9NJQBz9g
Q58etNJAsukFoUN4oqQFyQwLpWorVqbCgf6R7U1gb/q38jHfpsuWDTJfiMTbrE4uB5uYTZjzMUHP
PSviaj4MDlhY5HWweaULMQH4ARKTsVMjnVgBuYNffMV8U3RAOVf8G3r53813AT/QlShwFb6NjXrN
PiCNyu6nG/dh5+1Ft/vQpAbIjEaNWbFi8Z8SJsn30I7w3lOFFRLkgTjtrn40ANTNJhlFkEn2cqBz
bii+sDDfMq/HD2+F7/OFmnXn2cL6Lc7ndYcpVl5cxJaz9L5EuDYBjMfCYD/+OWnbMzK5ybzMXFOC
KudfKdls23Ma5Qpa8nSdBWJH0AN0ySgktz/EgSE4j0loBPj8CwpRbl+ni6DqmyWiY05pjtnuzzg7
647MGZFg3cEjUoPm+YNKsqWbb9QtJWbNx0AUERYwCiK7/fmlMu67or2tlaMlsVe8gxm9Uk+arZGo
puCTjannv9j3Ylb6MM5wDxG1mdIMmcEGfVdj6rPmq+h8xnXs0Lxg2/9nudjTblwL4XtkqmGOfv9a
72YypANV+KBMnK/0ncL/GNWmaQk5aObFQw8Xcjf+2QOO87OvfoUeL5rft0IbKg5df8DPfnIPSrBM
y5RTHYTk1P3fpQ2GTZLu/GXWBklnmZh3K19AGteYDlOi9NVBsSwkvSDJJOjOZPe9WYyiDr0tNz1M
w80d4AsPMDLkgqnj/O/yM7HK0a1g2TEyl9s7z47AOYlWS/x8dDeTwaAViK8B/afWIG+81ySZnqBV
Y3ZM5yvl9xp+0UkLb80FR4kKo4xGD2Mp4D/FL/Uy/sGXKpo0M81ZukKVhQ+gtcMHGlNpa+JZQwup
XPbvdfLrOFljSdJbMx7Kna+0eB/u3gGw3u5h62KoLtNZ7QOx+FRyGS77vD2zH43RNIgdpUSXPoBf
9uAYuiuaEn7M9tqSXjsLu76nWCZOdtormQ5KgJuU9x7kN2+5E92ctJIRz9dle8ehS5QEgF6bDBTF
tstuA9fPnHdpRZfwCg+Mw+jXrO7XfmQG2Ew7w3N1Lwoiomgao8UcYFQcsXUGAmz3pwy1mL/x9Z8q
Qx6r0O57EarnUxdRoq710eiUeGoyr2k+o9hq3xU9XvLisITxTPk7eFFlqhE5ZDORXEtvsrzjkEeP
5yly5b+iqQYSYhwBcTyrFDY1FAJFAAX8pZiW/wWvd9RT1aXHERu20Qr2NGIz+/5Rpguf1qJgHT1j
3a+EIm2eaAtEIQmxpj1ViLlB/h+Ha+q2qjMFVV7OP32IQNaVYhI7UnoO+BcRQFabWuHjpZdNQU+n
A0tZ9WP9dgujI91UblVUJGvO4Xzsh4e/U5+54fCKPMZ12B6OfnvfOCJZVIkrZmsd0FAbbKlcx8GY
tDjj2degmktD8eqvZrG2mFmfDZuThY35BQ2mU+/ePQ6u3PKQ/95PBREAYpxxRJMPw+35hEoMQ8RF
l5XlLSsni+TCI+U+myYrAoYiRLKyUQjhm6GrA68i0zZClrC/74vbsvcSk7IRyzCwp1wHc9MyLvMm
yos+j4Ujjyey/wBpGPe2dWoqt8mPM1RLxv+FJ0oW8noTq22MnjoHz2LVAA7ycNLpyjr7pAVmXgMH
HtLgRvTBAPt3UihjMBILZnZmm08LW3m0CY6JWKVvDRXUaSVYtLH05awz1hhy574dQmCAPxWHOS5g
DwmO8tDkNkbZAiPwOfep47ivpM3HXHgEkLL7CyHSrCoZ4xLC1s+2oZF94Vjulbo5O93xIlFYxk+q
NscFQSNav9p0rdLEVElThxvnv1tY3Sw+CyxUDKumnk8ZFfBdGEQfPKekV9K0i/7U4wDk7bUVbF/G
3HIpr866juNVXlitcFYVCIae8rOFklTPvpaJ74NJBlkmlzzDiDiqNqjGsjNvuEUXS8rWISDWX1FF
bRFLydEc446KSq6d98l9RUH/jd+cTWuvVLH4hgkM/aeYFvj/JwHjA8nk+nCI6+aIM7jGUoXDGB0U
N1id2eYYChEciZIagqAbFxTPBlqf2QkrfWdif8UVXppj6ouog3QxmntdE1QLB6H9KXFem3EkXBpX
2XkAmNQPaQ267/KWFA8MFRRaTgDDl/5aRMOsOdqnGQG8DaQdhXFIg/8M45nkxGxteSEreMyMeMXI
9Rbyj8wXcpb3ACVTstK1+6WPOpWUmUHUhmEjLFPjF82C8iLgZHMxvk9tNvxcWI0TxBXaQ9s90YfP
SOMu+hSityPMJqf7Zbc/B3llx3gyPrVnIvjNf0POnH+iiZFNxpBi6zg6s5aYxoaqt7KMU0UeYu6w
+xlR1bNbpLcSkyvEem4noZZDncT5wtDjxmSKUVhy5oDkmbSzhJ07r+sY5YfXxZ0sY4X9WDK0k2fr
mxo8gBb2eIKjTheOcJE4fgVcpIVqdPspiNfaS+IBdtZh2pOg5H20k3LH8Zir74q1NkxG4Pm3r039
48eKCTJpb+MCTi8S6x5VlxeIZ8Rcrfb9770PSgnR7vip3gKASxvrR6nkWa7FX9/mYgOH5jikoHqW
2Lyd9Ab4pH9LkItYReWsVssFLKJSWHzYsSkYH53EexiEjfaFJx0Yc/DaCtGkPnnUw9Q8mxIL28IQ
y9d2dV2rLyS/qpW3ta7Ojoo3Pi3/EbwZMJtLBvbQjLs73L/DdI7kNakZLwO/SNWNsvSZPBzMivJI
ZJmiYanxk5seUUgw8nyZRhWjFbyl5hmQFXnYU9T9XZclc6mj3X24PlajsEJLMvzsCbXWO8dLIPD6
zfw+0Z8SZPj1rWcWxe7TacxcGiYBQpPsyy2lPipz3H87LoRPg4ag/3PFTIprGjg1jWXNEEUiiEPM
Alp8pq2x3l0AsIjTtGa+OdGKA39A3/q59WUqEoj/+dPBxQmeEn4T0Au8RCa4HAoKhDPZNCMrZKGc
hRYJ4uM3VUNkJIQIKjocnAXcfaHkxSFkQvgncUfrZt5TmOGMWkqofD1sljlEdPUZ5oeilphUcKW8
HX6Eqw7OBXOF92MdsDI+w6nAHpv6EDI66oihx6EiL6+VnlweqCi1HWmPAIHr9vR3kVEQfesVhhKA
1Eanloy6z51aGbSk5c40n2C8Lz7b+BnQut5eygWSN8YAoL7tit0Y29QUdE5vuFMpsRmxOL37jwu/
F9/z53DEUzisx9odJ3zLZhGSTc0gvW+uqKWQzLKAEr6wE1SKE27Yje0/7lZVHHzSAz2ovk879v3l
f02OBc9U2YcyfhyPx3uRtXZjuFs9H065I8QsAx381IWkYgpz1khr+zwtoh5fjID7U2OfmWL25/mZ
k4vSwzsh8wiWInBnBUM1ibHBN3r7Jhbi2+Yp2JneiAgxeVoh84u163U66dvOlYh3qgL53Rz5XDqJ
ZDtFEj5MPOBllF6E7Qjc27xNePoefBfdaWpjgJIasf+6/VlChRjusZUJY2B4tjcRrcgOhBcofUb/
BSapQ8bfpN1apCZE/6SQYlrYl7HA1TtNDG8yWQBUfKS6fifSNFksOAbDy6Kv1NcRyvxYIcOLp/y7
nnHJ4djkuKSe05nId9V8FCMXxEJbSLt/t000BVNU93h5rnQM/pH0TFKEOtfW/4CG/khU38LHTo4x
xiL9qKjtQmyu/CI2dAYWWNHIGuVza52lItY56W/ar3Sun24SK+vUc2qmIjemmiJOT3gGYedXMHe+
25xXzco1hG8ezULdfX+F0poBGFHwGrRKMFJXYV+d9KBNkzQFvZ1REpf0d5SoSy/Mfk/VfuZIpYpd
6+mEHp5hy/NUePMcbTUuRRtuwGwnOf0aicY9jjBxKjzUlESC7qJm7cmE76KswMCKQeOobM5qYsdy
KJ5UwcGLDBwZINNwTTuum7kVuigN0IZ/3aoCsDSXZA6aKDD3SEcgFnuZztbQkvbpDAZvMnWHgLdw
K9TehoUfdtMbFHiC06KRuIt5kPgBUwDLGXWFoFEAbIt+Rm4eE09/bbs6MgA7eiUX88j/zRxzRCT6
8cnT3C/boVEG8bax1lxT0p/cgg0arSPcJqLN93hbaJz/B6hqE3jBCI2nZAwzLw72JiCkpa/8wZ3W
+rsrsABRGEjv/WQV48uxLKET8fpp7JgcdNwRgKh9bY3HwdjDTId6h5nDgMor+UBchTSqFrpDc4jL
iR2BcECHs38BSXnPc7W8YxR6LPwRaad5JyU5meLXJJWfgit1BKN5lm6aHxnGQ6nHkMLRewoankTC
pZeE2Vmci0QGLTvVe9XtiYaw3dx7jalX7PEBVTrnM1f8KC1evKsynNUzEPLae9h8ya55CKrGgp2F
mlLKhOeE/83ZiwJ8A9OP9TEWJo43P5v2aO7eVI2sh639SubzlGMQ0YQwQU7nFtucFxbG5nUfxOKz
3uaH4v3+0A82b1uldfOWL1Hq0A4r0IBwIpA6I9xVj38TnKRnz7CzAlavtCxpu3c3Z/kkVUEpDqfd
5NYzdiN+cqdug0GNPDpPglbMU2jcq056NRY1/H/LkUvtVYdq7wf9aUtxn3Gor3YzL1KQhj95Ix0M
Y2vcbKGLLai1v2FbBmid8dGY136F5Lc+DHAP2AdIHB+8FWPkKpwsq74Tm5ZalwnsV0K2tDEsmLzU
R4ASr3Fem0usv+HhV9enqANoaTZVnmT8KSU3HB4xROT+tfR6unTVaqjVWd1dZ56sT0DP/dy6owQA
6hiCMHiJxEvJxmvXSIjy8Ij0VDZiX6BDjaHKdfgMTp6ORtTPDON1Y3acylE2yD0x0Unw4ahuF9GF
kARqkHNqv456SJcv2XugSoC39NUqR4nkciagi3JxXujaBxnFG+hQHuOWAbKV2n4PPpKLj7q0P31F
A6xhFD53ZntmPPdq60nxbxGNBxvEdp+9ZzoavA093kYTOSezOLKIJsG76oSGFY8QIfavdAagLzPd
H5QdgXLa9lCLEMl9h8eBBl5c5Ki4CIT7YuVQRyuXf1qStqYOhJmOSB4QgcdtgIYS9srtW7+yvUrU
mvJhmSLu9Rw/HQKMX/BTAy2oLLwPMCMSibgalIlmz+KJb/efou0Xs7xOK/rxpxyeYr6ZAu0QKXor
Mlg5p9UPj/pTV+ftIvdYdMS2wIaMQZVFbptn362v24LQTjCeDq53AjBzUlS5aG4PPtuK7egCuvRx
E/YTuSW2l9JubGTcMI3aKNgHKKOHqnIWypliIh42qlnLZHTZaVQnI/y91w1ViYBnZNlQ8qvkHLB7
X6dGuXKOBMT5Op/qsR+9ZT+aFsDp47CYlJNpTB44Je0WJ4JRFOk6NF0ju8C3JAWHCl9oJnlFVVkB
oEk/JyyPzkHc20Q2hGsvGwHmW1qGBT5s9TdNTiKcfJiRG8fkMSvgjCMiEVDPdyR+/26n7bg4w5ji
5buyA/q9bQv9LoIpQJylHdGZbUERW7La/M3wVnxNHki+mlrR8IGrqEq+1J25vA/pxB1N/TQ6KHOy
lpwgYbpw80/RhwczmvvUH/O2JFoIu17YhTnugM/Uc4vMicROgCyf6YTr4vFAQPUSyLQiQXZwtDAa
5ucDLmYnczo/FJAASTrIwJJwr0SuI7mMqGQ6a4eRjTgRLYXeySy2R/pGOk9O/DRl/l5InLrY/P7b
XG+e8UR6QbkVkfi8QTFEClBB+421hXHgbXUiRYuEZmtj2uNzezcZ2MzodXJM1WuiuPRtb3GuZDDy
oL5BLZfrur2VnNfKoTjfB1iuQu+xpOZ9WWnwyXH25dTA/tRQY7T957GzyBDV+PkrUeO7yE26E7qV
D6M7fHUXvZZHn6qubPtLoaDJ49NVRPKdDnT7cum9OwcNHgvnE/2zctkLf41nmVTalPKmQWoEeF55
tdw9jy/6zBJ0V4z5NYOPwp+wavprSZpdYJ+vrsKsoPnFj94sFpepwdv8xPzPmP4FiBN7K6T9IU4W
igNkviGWqRzkha/HE2MyLMgbYeldMZ/lY+O8EYIv+YBmDbXcbPKtRxiZYY9eAkRFGb8gb5vO11kD
q3WfbxKV+gmJtIWb85f0QXX+KVeWuqgjxIh++y6iplCItwDA1Jpb14r89mOu+gNg5/thH41TbFiA
VD9ju4rjWFcP6dOXnQAdwXkAbkipqWkNy7u1z14hhmW0uZwgz4LR+vFG5Erx9TLie2L7XEr7ytIJ
M4DYTMRdkFR3l83evx3YQtIzVFRR/vUsfxhSa6skSQDd8d5i6KBq8pTNG355OUnclk+kJGORaAue
TVHJxCAa6+yTHaXKf4pXItTWzNanHBVxWIbvU5c90JHz0jw0q83NnuYw8Mm9qIWDTcV60OARYhPF
pfjfAHZjy5KjqSCNQIxWySZ6AFWx10noe6Fm6uEdU494UO5Se6aZz/kY/wDeGaTpnu9jBzG/qxSL
0CZgFoaRmJmwlsOWE/ivqhU7FYpCyS5SAyAgd99Ra/5kBph4ercL/xLMlonRWW8RZ546Lt0YuYiF
y753HHwNKjqfFDRniUQkhJTVg1GROyq49D+mtJFxE/lu29bZDYq2Im+f0RvAcxUDFPTXFbpFKSVk
scTcHM9NVh2bx4CNQYHkNLUgDeXqWz+u2Qn4YBp1wsTGltAx2+TLuG8yzUW0px6IlS73TXZqHNgL
oYk6b1OiUeNWi2pBsIGJzUA2vn7BXaXPJYB6XbMGXpONLXQB15sGwT1fGmmNVKIXvkOuuQ62V4lF
xnbU4tCuFKQGIKr2Vv0ZIYpD6b9Nb1TSKscKn7jwDosCIaODjULvQEBwOZMNeygMgougQS8Yb0XS
goSQZulB8g621VfYs/uxSI3g5CqoAdn1LG2y7hSbiD0kJIqL+BBkqQXSNsLreACSiT2qsufNh+BQ
ZhaR8byK6lf5EUaHKviZadJRDVZajAHR8w60mZGYYoKXG7YkyhCNacVPU3CB+co//+VPkDs7Cfxu
Drm5LLPf9a16/92qJm5WxXIAWEzPx2ZZcKgQsaYOk0acXQFBUhqN6GMaKHqQBSD5vEtNeg6jjSlt
QIFT8sof8wbLdT5A8l7ItntyxoZFNfvL/v6Z4PdrYkRChopvDPaz6+X3cr6Ni7aWpcuY/ksr+v/A
Yqj2Z7aRMyCfTZGaI7OREYGCa0asTZai4uWl2+jmiab2q2OwoMB5lHmc2ufea7AHJVRl+yXMVrXH
cLrnVsyZewaYGPV+YVIxJhvGz8Nj6Ip4rpE237SOXdTQTmgES6UJij97VGDiUWvdnAMsK4TmqjVC
XnQCuA2zSKpf2MdOk5rRTR7yQtslD0N1zPJEvpJ8z9aME1Aic/lHwtODU3vpEYgz1Xk0o4tUoBYX
3A9lhGpl+RgioTcLXYrUegrj8CAGgc/hfeilKhxU85Bvp+LRAedkAvN45qLyipC1o0uJUdkQVAb/
lPbsSgpbOJzQejirreB1REJSJHRXmU4FJaKzDcyLUZCmon3NC2G6VYpTWHv0NkF9z4hoZs8SGxEt
PI5tDDCgHyncHj6OpudN7QgAX6p/j+K5sIcpcafhI6xm6RBWuKD6SrLcA3Pw6fd9pUWzdFPkO2B6
ORNORwhQOxOopHdGNNQUxvjlvKFRftREm02uyR4Y2s8cd4RpicN1TZnDqxzc/Fz1q2aE/00/U5MR
9SDreYCFOO17UAlnOQyoGV4Ufpk4gIBSvmSXP9EctVBbokDKqlNQQ+tWoIHX0DRIlNoDlR4dJTKg
XiFm6GEuLk/bHpPRb1aG3Eb7mwEbpdUTULKPmcOILjmg4oMJljZdNGM8rmIvq9B2cA4RhTG6rMUV
CQ7tJpNQ9Rc8Rgk8mzhLY//tBrZKkW20t65W8h8a87bLP6Xqx2hwNsQTlLBrBWom28RINj0BOymB
KOOIOWW7ahZbAFy03y6za9oI9Hu03WBHfbO0m2q9E9M6VQKHHvbcn1/YEnUWkm+Qoyu5/c/5XRRj
Ym9g9dvp2ZVKBfrJPYT895uaYZf88qhjjrEbY2iwupWHbnIaNvbkEA2E8cD6uD9yv3DXCn9OyAZW
iElMXd3jb3vWZLKwUAL478EKpXv/a/uvHCcS41ce5TLI26NTJgi0RDQYHOI8IMb8dUHyERouhf25
XQumhysIeE6Py/oCFAdk0JPmUus86m4NpFmIcf0IMkhKpEUJxLdqjTmuWNcF3UkxsPxqIxrIMyPb
pQ+xa+i1774SiegZm6VPqBWQaxrfJ8oJ+uVKnsy7lPGDL54GTLjYKe0Okgi/FUy34q2ycly0eqsr
zX+o2aKmI4JLkBQFo31sEE5LG65AGUhAJw10NnQZgZPDB1/RQ/CmAxqDsrY/NoJ8Cmb/GufTF30O
PgAgQcEeKeSne8wcxGwntrq+Yjozankovboi4BxMrlVpR755vi2Jag/uxc9VCkbFkexd0zOGv7mZ
g/udgobnzSUYRPt80117NRVVumoyArs08Zableq8dn24/zLXw1U0pRMgArJxS6uo4Z3VFrKb506l
A0Uq9fT9MxAx3+3MNgM8tV9RJJvFtWPSw1j84YReNkJFg93U7+L+7+v3wXiXeDNW5I8uCMwy8Ncq
HcqjnRaxRYALoC3RTKQWt1K11QX230n9qfCD2aEGEeuqnlg9Jvej1I1xcPC/S91kn2osn8unA+vK
p2K33Cc6ad5yC8TDaBFm5n8mKW3G6qdcgrAVQTFXhbDg7iREyAInDXKn40TUVSPAg4gA6goCR4pb
wtRtGPf1bGjWiVNkXh6Gcg+Py5777ouOzg5B2WItkCNWMLvueNziXVEStWBH1i6zzI5EkDA/y6aG
N/lLXuJppXj0aKHvEoViTE/Haj4vUQujMQg3hpLQwsYK6qjhYljMEGwkB4u/fsaoOTGQg73fUQeZ
v75MZJcWds6ByaMCBJvI365CkYcuac3Nk9wm68UoTaUQS40XrO5doxZMrYFcMDytlhLCr3VQ+psP
6nSdJ5imjQrHpqRoi7tG7PTVWewRU/dwlR3Ab3V7bHCmvbCCFyRCs9aHPP/9G1jQdWqdr3R8SHp5
kYwge56bQrSGtWJ7rhRztrdyVbTOtOa4/hzZWzkt0LTaz607ccaqEPwPY/L6OVnzJ457OXe39rt4
58Kl2K33Phl7hQsZj1QDXAG2H7IvsHTUbx5TN6OS8ErHpTENYnMgbXNc+VNoRDa0tGuan1vWzact
fy1OWK1kdtjn2z8e2k81mMpw3n/hZbGiPqGpftFzqYkqaYLLO2bUklBTworGLmqgoyiObGd7CPUu
YPY+CNQ8PG7sH9ht/wfkXlblpTmoBY+fECLSifmBmPklnycc4K2YIrZ2ijQ5JrDzIOAVVWl0gRZU
LOvFLkErLdcr4vVjjrzJB0baLfWIYfWCn+L1YGg5vQTGm9AD+xXZEF5jcvXnCgYsO3PI4I7jifQG
FZfigOGljWJQEkx25b+2whONDDYdZ72Jlboazqu+/5epeDcPJCo0Rh8H6B/OG0mYF3jNN6JpQbV9
kqDwx/e/GLbE0iuRRldYM1bNgF4m8nqbxJBnJ0oDcVdh8ddDPlFw0o7wU3kM9xwp7ad3Xc5UMOip
JQVKL1DCQM3MccqH3lcvYaRTMBvJwUYamWDvMFOXCTRBXgjZoIDY8IBziqsHxw9nZCq+yp8yHHg6
TnEr0x3LFYhII98xAi3wupfR11IKoFp/Ipexam4KO1HDne+O+M5Nv+8lepfrLbIu0FGjXzjEIfvC
sL4aQFPtj0hfEDW3AniDZkcXeV2OElHIDjKhI7WNJ6sZDhH+1xnOzNX9OMKrrPO+kgmtl9wf1ph/
AnohIc80tFVHAK3gZwfO3kga6RKmnvyfNOxagM7UBRqo+1akzOw0B7kZhKfKnMkVstfz0lZG3zdh
nUjUoLRAcsgL7oyJafp85atzFHHTrHnlqrv9gJM6IMssRj/9lDRnAEJdT1BT/bpQORuKT7BFBu0v
32vgHvhBEl8zqkS1Rc9tYrmCP8dgnoolW0kmuBXCgxhUIW2ytvdu/C8GaglrzhxMOLhcJ/S8FELh
CUgNXLqlEBHVzOn5CQLf4nnwSFL1bxaVL4GI3kH3m8ve9TIdq+tZ3OEnR15yufxYlBE8W813qv+w
1NVRFCJVAdt85W/Cn1aoMHaN7txvG+x4+GVGZkx22QyMakF4rjB4YDXo8QM7RNlwxbC5um5sumbe
9a7QeXbh344n9LoIlQti1pCHw9+Sn0Y8wSXbtJGCzteNQcyHOoAGzPbBljttL811DV7bUItR0s/w
esZ6Rzy3s+i+C8IdT4DsRInqVtlUEl+rW1PCVuEPWXp0FnHT19ka/NBo0hnAVrYlzHRBTDY6WArk
rgurnCygpiht6PoDqJNovqm32XOWAiG24yCIIrvi+sSLurxJxptj3QRExIm95fsfH4GTh0yctdVJ
atYL7TmJfVuuG561nfGz6fnP1uudAxV6r5hs8FlD+SgJE41Y2quzj/bAiLVdEXfAXh0nQySWUMU3
uaNc9apoHY5cgV5NSIWDe34dY7q7F2QU2TiGI/0Ii8OK2zWfHlfy56O+RwZU10VSVlNXb6hkcdU4
M7NIkbUVmabcWx7xKbW5aVGlShn88tnUoT7T1r/rrzQEG4SLdSD5WIiM2z4rxBliJh66swfKMWhK
koFPtUsT8wN0X3Dtm0L0UYgH5/2brcdWbIVTN6OHBzBg+aqOsrNJOk+v3ni2d6GahGmAYZFr4Dls
S0LPqw/Zwnm1/TvxpDzBKpMHokIQj/ULp6bKeFF0C+NXqKvFNTYcn3tF2bBt3eMBmSWjW4t5sSXf
H4KEsmb0M25YkIq+AdqTR/GBotDy+qpem/Q6ExW83p5XYwlHSSKrvTO8GaCDUXREJzl/7g55fxwG
ELxARBN/JdufIQ+7sCa23SyBkuGSg/RQkU3JKmzXXyoo+lexthg9KSPJ4504H6RGIKHSDB+tB+Kw
shFhaXtq5QvFKa7zBmIwLlqhQgxXmJDOfO+eXkxfpdaprAQzoQ7GV+D5Zk90Pz6L3eNsgbJOGfZV
t5e5ZWS8Dq61D/I5XISAtdbcvXhadoI9stU1mVmSaZNvAMJONCforhIwa0ou74jt6u5SAvwhujbO
Yw4JYPLxxkTi8mf48Je5eVJOfE42XGhR2ChVa+ePBx6a1Kj/EOL0cAwgio+lmyMSpEN1eQCZrAix
57aTOnvJo5FE+iupIlD3vjZxJ2gAnXmYuSkkX7IlKgwjeeiVjIb07qbdjl6cOnmniOclOpyLanqw
rdgyjfF9xy6WUjoLCESe6Ag+NILgobZ2VvVr96Apz0PNnj453WHi/eQQlO9j3mbqrjHKvoC7NXdz
skrMsRw4gGckv/G8COqR8DNhviMJlrYip/2ZwMLNg4GQ+4Mkai8PIyeBnZdgOcJlt9FgFbD/E/u5
eyG6nJ/o1vJCjqLQFrF90gUjh7seTdeHtq5oReVCBva0lddL+HYHehbzNfkdVzVQQUcRwSZTVo9+
08jByFj7qvOFRCGttdTFz4xqgeYJQAiBBiuAFXlZSio4SZPkKtXqk9fPgReefjqUjrw83yEOpzQ/
yB1dvl4d1XEfi2xkN00e7CFiKVQgxRyVXQRqFl2FemkJJR8HpppDrL0HLcDpRz1Z3Xs5MR2wePUG
2Nv3VapBmGp3bquKlXkMcRAIuNroQe/y0Y5ckpP1GMbVMM81U2/Z3eE8JQzJ8OdROg8DdoA5xcK0
+jsYdObWuzuNarfmtSCuWzA3jiljk//4p1joG8kAH7HM3QL0LzKYETMqODQ7Emca1QnStGnv1EUN
vD7XxAk9YSuk0jP1xtv4Zr2rKHxE4ataMCChRyKFRaOluIklOnToYqy5ALem1CmG4ItueIsu+oGg
es1ihmoyiQY1CGV7gSi9r0zxWNNLD19CNwoSJRuJpH543UO42d9P5Lt17j6afZrK+xf6Yu86SFpW
6WPfMep8TentbuASgbmtfyqGmyqNsXOIOKqbp/2WEaokmSaB6ks2nuzhcJdPpDpBbDhPSIkLiSO8
bhnGW77P1udvv49tb5dp+M3MoFmO7Sgyv9byBRcrpeFY3GhjcAROiZSut2t0BosnXRT/bKzU1s/N
L8+zaGossslYZkgU07V2kcZdBi820TQJILR79//aAObNJ3Ax2Kj8kwy4jaDlEG/CThgzhA5r5HWU
VKDxtp6Z/I+jolfCVnEfDpwxuyCRVuqt+qVkYuBtI6VVtKTmg09n5mxI4u4aYOOqp4P/BWHiC10Z
m2q8LTAh4neWhpa886PMHIitPI/k/FQf3qcLqbWZv3tHaynztcdLa4VIoLs7cUCJXaaQk8vc3kZ7
9sbhXKmKPmOgqDcqKowZ1g/Kc48LY5sF+vqlQ3g7C0mt24SvZ+FcRlQAHTcPJq38/FQTb1rvmIL0
iqmhRy/4ktRqYbjKlSIBZNIIWPpx31kSWZW+Ga5KJ6Fc6pmCkFMuj9xbqAl3Pdikh6V+B/e/aeoU
fHtv0d/t3V/fjC5qigloG9QQ4WZxFIo9+egk19QLOmHbtwO38WMDFGKTqg8s9vv1twzRkXAXoyxP
mMpl9ZwC/MI+lhzqzCCITzTAvJkgVr10UVJZJoXD5+C4hmwof17Fiv0MjUcWIIYdpottLHBZSRFm
LF51cMixE8tHgB7WrbjAWbwqsSit20UURjQPZrKeh5F2GazZHAgOVSHrRhenwcO6EtN15jE0QItg
g59VRmFHcwdvBbLOnek/X8kDcTXSeiaSj9r2ioHvktWIyxpsOjXBlgmpL+FbplOO38QTtDFrKCQ5
C2K6LKX5aDdnJtg2xz/GSOcYW3oXoFxqK6lsUtyQLFSZ03OP/7qC7sdqTUCZ6N+Q/+Gt8KO/7bjA
CSX3y4NWUlNyO8RkzrTgcqYjBuztonSKnRYSCTRi1ShN4+vFZfdibFVRiY3m6vksR+to93rlSahu
FwpyLMxcH8bbKK7AAeJvTlGqozvYZ7wSeeLBdJON/vVLAaK8avWUEZGkkmpnmBjIy0etTPS6jcXP
qb/CpdBfgiUeTNUgIh+rQ7dYR46SVKLS5wb2X6OUUwUKKzBSB2V7R7Tva0pbUevTfV7JWS/Xe75p
XcEHYyGG+2Lx1/0iST7WUqiiAnvP5HFWCImYOvKVG0HJ/QziJ4hjbqawFWQBeZ5HogNa0uunP2B1
1bWfO0Mvs07FMD6RWnV+KE5YZW30HUwJuZ4kammJxS//0C5o3qX7LVD5P00olC4tTcoDsVoGlRra
oT8cFyCsfVDKZZVeCXtPYQ1/w70WX6Kz8sJg0K0fSnYld6mf1WOFQ25Yz6X4mdhr5DZCVzR6aBZA
Yb/VxcZTh5JiaB1EZCLvnoLsPA1t8k/SUgtDlYcd0tiHxQuNkJgAAV3w8WtA9kClpOv3/L+ZRoQx
yrvL/MhUOLauQJ9jks8u3Rr+KonJgaV5NVzoNkyVrXM7NukzWAdaQ+VC5zWSjOpR2xcfMbNGoc4e
5h6ThSucGCh/XzWjOfTmaQ0qb3HvydnNtkNnGMLSm6xgNRytH4Ns4LjWk0ENiXOIIFgVT2rcD6G3
QiKRPEx7SKCYUZle7BPj81pggyERegVz334tf4Bv/oPsbws1X09siI6BdRVxUR8kcCr1cUlmJLhA
69du0wKZgRJe+g0l2hwziZ0x8SrJZ0itZscMS9H9OpODidC/+z2OFJTBvp3CxaXsZ7qOsh6oeMue
6wbZgM6xCcI4RPou/CvNN4d3VB80oLV1Y8o1UycD4DOvaRQrrAKCO4LJf9aykHvK6OA/OYjqjL6o
z1LuNvuRfPKvr05qxMq6gbhI4TFE8jNAkPOeQyazlsfmgY9fGu/C+B352ZLwGHaIhEvhw7wWaeON
MYrnKmK6yl43Dpa0rQeOatd5lgfoI0DqYI4fXCVOwuwpYBstNvL9Jlf9vL8enVN6Ojhy6so2cRYi
qXBHcgFMc6vUsFSHOYzCVoFNcWA243QEnyntplepdB2NNBb6gFUBVx095G8dm1D4L+Mdun63+jgq
E2wQhPgi7rU8E0IpDIvbTws5zPw2HO3prUt7unx0MviRxcQHOPgslzSxXF+LuQRo7wClooIgJ5Ut
DOp5evgPOX98GQdfDg10Nh+uIXA0Yx5CwLFNSSXYbFYUQ+/7sIB5RNUND+zMzT3wKvUj3Vb7IqHU
b0sslIVWWZEvszH5LRqFAyUH3sNQwD/BK8SF7N6BvtUoLZdEqQnSc+JNacjg6RJdKLLmloYWo5CA
7CVb/t6fBimFddD7EmtjIAs1j8vP6DEb3AqM9kRs/hRKq4OmKh7n5kFvCxjn2qniXhEmsK8iWZeD
AD9NdPtMiX2lI9u3vriUqbG2benBPePxAWpRgq5tVuQC8ikEwiLyZIH+J31KlROqddLC8dSy8prA
KXOgSzsCEeLd8BNH6D2+UZnTNl/ZXYIBviUfPKtKSNmzPxrnIaHnbaDg3iHsYje5Jd4map6coux2
WHvRJ3gVy5DQwT9XazWcoFzBZT71lP4r/MXg5dA3dh7O1HqxjI6GbeTFn4LVKild4FfCb/9f96zM
dm58vVSAuEeIANt/4HbBenjFZhTixZ+aXNFqZJFi1EjAuHcznCU+MLeR8frn58EuRM2iC3t7RDQK
NlU6b0rgoS52+qpTgM0UOs21p/NZziLAWm3diVRUEbPckomBKRpymntQu/ZFTQnGgw0UkhP5avaD
+wOVjAU4TYWvMX72Vhw1NhGQjCHjBlBzxmljcvNcqFFtrdG2jwBBe3OcwUFTerQmUI+U0IlYpYgo
vKxDtUJT/cfYtPf0ylo/wbG+ZNs//0EseD3sD9iZR4Fg8np/Tho6QhvwtzXVs/pcYF5Tqcy9lORI
WCRWUVAGQmJYlYJ1JW7v/z7H2lErJRj4pK/9jNHgtpK+fXJc7ux666zt+oRSNM8A07QTyVathNzZ
KGFWyuHbG7022MkPEabztZuNgnAbPWbjC4uEXc+BsvW5KTOayy/GA6evncSVzhKL9ndL/7FaLE3T
K58ULMZ3fTRrN6udKglY6icHg6Gh2HK0lsYsYXoG1slVd/u+sv0GTSjoXisGGnJJhj7JFbDnuX2r
zG6GKDDm12Sq+BiXdVDK277pINRiKuR3v8Lojz1COmHGBAc1+OrQ/1apMd/xris+EbmwW3QdREN1
HR5j2BLd4Ey9jx2BwJBS4LDhXyAy7WUELu9qgtc7pQm/6wXsL37fUZQbsgZ9GxmYpr2fbebe4OHX
kSfZArbdKj2Sqq7fAeYRQFdQQm53ZEQ10lN3qAzVNsuU/EQf2zu1916PmVvXi2lcvA8LGclJdFzn
Z3VjNLWI9Yukz2lc+2P9SwX0hZ0KWveucsBKtLd0PK4fyb2sgHAEsPFMH+iHDcwiCOm7Eg6DTb7B
BRH4cbzMDfMnc3Wvqkowl2MvyD66FLl4G2ZBvoPKLFU9a989xLOAEgKcnHC+9GGJu9YnJujHiJq5
j82xbrdIoRMpNe4m5sYbPyIPsOgDMwp+n6CjAKhR0wKZMtK7PtXs2ZDphsaA6Lfod4VvP98cl2LE
ijPodYS7nLLqeNwhDVkx4wwe077kG40+q4O7czzpjghn8QsiknTOnk8PVeVdC+mR5sdfN7d063D4
tNtO1Ncd+daB6DnkixaPQfkohpPVh+vTTMM7bdkTUr4BBAuAjzEI5fZWMp0gr/nOl+MWRdo3iRvt
oY0MrsyBN8l1p/XdJ0WlJxmer6dtdTZRn6/Q7gQCHo60VYlz/EPQp6RTOlAVjiIXARnxd2/gqIjf
Swkicn58n2PUxQ7ht1hrnqz6c6NFtZwOknNBM0GE8Nq0FdSxpu9yA5E3v9EYKaTr6Pcy65govCrs
nKdxC0xOgDxib6XxodwCZn8BpsLVXJD/GyZ0q0qOcC/3QOP/8xdgs6+KXwyf3Z4LtVaD7zu2HXYf
OVjuj6IezceVQaoTfc65Ax+RbmmSOoTJ8S1fLesXfvR9FJtWWrFpDUfFgKrZT6+c05zwDc3SzPNX
UTq7rrdqBFPYmZrdBkmdWEFYkf99WmF9CInlwTClk8y1/WcWARK/qQfLfnyNOjDpomJG3WnYO+Cw
DwIqTZq8VN5gKrd1BGDNEev6Yibz0kyzbFoSZbkcqKxN4zhB+y7OLt/kCaPyNz/nQzWFGEXP0dFH
PpUIPTjKM9l5QoVLRxZ2bZe4oSFj3Al0XzsJIFozw3kXQ1htlLRCuJKoa4YmUaieO7lVlD7hFo6r
O43ndH5CqCLUsykdqgsV1I9HrvenAzMPmNVxeyH5mYkcEikA1ve+W3iU7rtcGn9J6HVUpxNycMWB
5oOk6iZoaMBk0g9ACnYAQC0yBCpitumgeEMQ2pbT3G5yF+YxVmWLXGbR4/66sVw8FHistp6hBdXZ
tbgiTVtcn+GqkSIp+080skv108NjROav50OeqlLXqgCqqVZ7RIZOiy2aT2vAaB0xQRupbMArwekb
cXm+PsEaMMo8eFeEh2zwGJxMdUI1TxWKheVuaEhoWA2qqlWnVS0ElZjOGEnS3HeNI919MPWu39kw
+BnqkRpR+3P775fV9crJa6Z3GXaJqvcg9F9VERhsZ0o7ZxcyVUlgyKMmOI3sJ5LUrzp4ORf9MrNc
zq5ac+WqFSJfpeDbvgRHAGcfJ96LnkgaTP7mmaEyIfjQoNCtQZv75VunMLC2jyI8JTcq37cbK0ER
Hu8JsBO5LdKLyD9JCEuKPrhNcLUIquLlHrACkKffEdQM9bHkrRC8zPpEu5KTrCHliHW/P0yzQ7zA
seoNKvAAv8XExydQvkvGf80zQq2YJR2z6s17O4BnpCAchqtGMS+/6XRwhSp8y5bQSUZbAxym5QtI
VhqeCe8xsKbAD2sZ3eYDfcGShEQOEPlI2Z4BpwIJjRs09jkGHJjHJ+LTygtWk/z4S2yrBMe29xLC
TWU4KKt9QGHquJU7clTGDlDTHopmaaQ+eD2A83Cir3BN2tOqkw5Hyz6Rd3Zdgpv/SRWW5rKEIFjs
7szR9SmhZgkW9D32x1/Zb8ZQsMmv0BmGdJIfcePGnCz3OmGX3rgksUul/TNgbxUQXChTjP/zePqh
tA7TJU/EY+2HPgOfE2sD30xD691hBELXC6R+Ff1W9j7n02CWQGlq09QqUHYbWWZvz+EnNLIjNsBY
6wy2L7WG06sIE1Z0tFqi+F3VxalBF9JIZMqAKL+wrzhpZf9wKQ7ktpBxWxj8Ttah5euZycbxswm+
UK463KiEIf29Kl1gbLOvzbDjyUwSwKNboSr/cle1mN+zZRipBcOhg67tMsLscPlHUmdwWOBP0K/+
3oFKhTRItUYbVDCyURiPOIHiPlPP7T6cIZaQCZuX+tlXdPK96v6y3b7USHWNFlCO3haj8OmafCOl
OqPoEemENMYbvF3hBdsL/K8ur2TWNXdiKhVXJpCQkP5cR3tyejQnalHsGXlzI/vXOwE0hxCHr8qN
tcNfom9KGLNPo1XUEhhNMCX0L+u+aCVZLOmZQY+KqoRVkGVMtA0D0lQUDuZfQ2BWmyVNA/hfdQW2
d7V9qqlU4NMFw3J5ele4wN0TjQCg5f2IBdBY4+tnDSR1mAP1GY+uzIx2mvt3vDxkr4i7lVLV0TyF
GGsxHwD8is4l4oqJ9VoZCU4xAmCKQGGQVVnt05XYilU0CC77N7nCwWp9fGQaV2NB6kalIPsHnwB/
0ZwwC8Qc0/Ikvy6pG9WWwPz1J7CRWwJne1pLsy6ievP2YvQnNYkr8i3uIEO2IXHgzMbvDkHyz/j0
+SAbYcIykN/QpDmYw45sFrkvqOD8gMwm+Di0c4w3lGQG8vXH2bwWSItfkkPh1tcbgwhpVPQuvbNr
+7qS/T06ZcFDVNUHeIY3UnIkE0wtc2pbPKyINLX5m8ObecqeL+4bsaKf+lbI4zJp3m1iPgNqjzNv
SIEOh5WnZdDQYOY+rzJAX/za+b0XHhVMgH4B1xLb/G4JEnpGZa+ionVgm0Q52WwpeyEX4ci6xyLN
Q8JGHCgttssIZ5tTnwfVwvLSyYLU5/2GWtM+nNa7laa7V4E7fdvR2hHZ95JcRrlFXF0WQPlhuJtj
noDTnC8GDUVOBHRCh3VJIekzGdXuMroRq7cltTFpxt9NX61ytpZTdCZLV3mXAX/CntatCNpTwHe+
+rT/9ClDt619WDqcyQY7IfFV5a+rv+MU7X0F3m7wS8zQ1CcsKc2xzOiVoIUrhUfYgp/aLRX02YhT
IdEzqau0NOSrt7eM7IyMyRxP2mVmnnHpGyZklr2iH2f0WfuCp8isOE72vW230JHT0uVE7y3s295x
cLxHU+GeQZzA+Pg22/1xt3TMmQ+NqZp3/qMouNJqbAvRw6WOAUR1PLe4JJ/aH5ODC2Ap8mn9bhZS
pbj9Z60Qia0mhW3hS759GRNTlNH8omO+hHz6+XyfxqCxRF9Y1ebFclnu4STHQ/Fw2nIrzfCsG7jo
ZLgST0G/5ApObyTnf8260zKCobMcvH3zMVFjlq6B3orsDsz/TajKT0nxpK4yUv0yskd5z3txYl/V
hi92SwvWxwb2+iaIPuS7HgK/xRWlgXS4ISO7koHKHJgBQluv8owpzvP/HW+KxmfIDWcdSWXL3WVQ
FaS654IbXVvpmqqKT0NCiUXVYIZkGID3ehjmPLeFE6QnheKm2JRMhTwIPVuHi/ymGJbhAdfMjwWB
cABljK2NZmbQzy/px8w2PkJsAvZl7IFbYt8qfxJJNPJ2jqJcFZSbBLfQWok4p+RRGmryVkRNZK4t
5M11hgeT/LLzK4llJjr/Aq/QK3Sirq3X97fynjjOEXYG6VQNoknafqN39fQcEW5Nt6SwtLIeI/03
z/rfKcC/rJm2URTd6xMicfs4V9Zgj0XyC8YvtmGYHtON0eGhGKMZBFejR8Pp0ZYruaoG5FgOKZHs
dwUGaN2Lw8bxgFiYEXdrkKgh2zKiemF8wF5OA0uNvB3HYm/pnJBjommPhYBjflGdvNeKAK0YOiTn
6L+SFMigS36R7QLNtutHXjgtu8GBj+JRIZawCLqkLGuYnXwwVlTX/EpJbdBiwc6foKfuuN3tDXRg
FwGlrXSdZBoSo7Vmkl1rgzxFLgn3f5kbx5Ero7TDswgB8wtJu88tOIpQNQFwtLaV1SiDhYRbs595
SKzhW5+nyFB+RLx+SW9GE+HYqUdYs3VMJmogZeGmBfg4gPF53DqWpCr7eSEbG7zBwmfcREGP9Gux
dVDGC4n4Dosh8kgA+8kr0qRuYfAhLRGbUTTzmN3txSuqa0LK5y8CtIcTjvnjF5t/l92PclPh9hnt
2NEO5Pony/0mXXuiPe8MoBEnDHk0kt++ME+2/kfMSIKMZ+r2HukvGIeWSt3ndQhEuM135DR7fneo
uFWoJ60AX44o4mEc//8acLhDT5halO969wx8GzKO9PUCJRAjrDOpWVfqFlppaSzY3jwcwjCQHSrJ
4dPyD5wQFcm04UbcmGvFwGW2RUJVUY+rw/VWlwYjbcSDqkhrRkPAaS18YvhBGWNEmDVDwhh72gEP
gor8i9wquh9iLcp4Tt1ecKb4hzyL9V/9QecTVPVSf+cQvUBrJQpJlWit/N7B/sxUr4Sp6eQloZ+y
l7FDfwlUZkVctsNFUZ/O/TfeN6XqE62FPb6BwE041EuvcEWpnG4Fy4OWWqmReRKkGfFMDh+hwHhR
yWR2IOOYdqhrNTWo3gRpkSCU1f/Ch2oTO1dCRXKzZv6l97Y5W/z9rKPX1kKhqkaeMRIzpS3Yi3HD
Xi9388jd9tBpRkixNrCeMUb9orsA13zYCQ0AgX+viU7IowmcDh4ebtzIVtLw7p0RKkgVqhSUj3pv
50RvOm4smk8TjVZ+S7FLqW3sa8TsLBjvC9soSWFyNhJm6QotIz/rltygxeK2QFv5VMOXPJb+/RGE
ewv2STni1y29w2BMH1su5JC0u/dPN2ujXenizKEcFjijAx0JZnVSHrK9isEsKUw9knD5ArJLWjEl
F3pxjmcwa+7f4lEJDYyHHvSG4XlQhmzGKpwyi9yc78nMjkOcdc7inhaa+ErGvB1UEEpqlkZOOeH9
RfwT1U1vCSHemH5zOSfZ+96hEAcg0Zx0o3UdYQhgHloOtM9/3Tik3P7H91JhNcLBHLr4vzT7kovK
FV9XyqmVh4jOdEAzSOFCjoVbCNKs3WJCsbgG8bv8JaudRlvZHi8Lh3mAn/CmasoQbMNzi5zuZf5O
EC/YEP4DYmtLElaxzmbJUC7U6hQToQBNiR1rqZyAFSGXSNEJb6CwdJE53y1wFOh5rueSuFMKPFyJ
d9Nj88Gh2tjhjxncrd7gWHVxl14XLf0/zau4hfXheO+/3EbObBIm3XWJaM4Q/rvBRaD/JyS8j7Rr
uYSfu+b/Mfd+eKwZGe7bR1ccwac01pvYWyoGA3HgCK7AglG1nY6Or4mU7OBgE1Jsz9JIv23Lsfpe
31nFNBY04C/SL7o1WQD1dy+8NRJvdm/JHQvT+qfiLWyysOOG88nmfzEaaZgOb6PUiAzsd6wvkgjB
zNmU4d1sNJex9DrHed3t5e4qVOS6oTe9dYVfbXb+hYJUNEow00YNHwxYlsywswTGstd1AjGuzT6O
qloag8UTFVpvtVWlzoELOSqifh6ObbkBNyEZEUw+63oCqrTF5uCcOwwg+3k7VcppCORpy3eK9sPP
kTOqJWeG6N7cbuNbHWRJgTERXpLktkvDFwnNu1VX++t7PKvCQiYor4lVoFY0BZ8aeKJ7f1umYBJo
AzOEpw9AzIeFKRxmZOPnxvC31P2oncEL23s3+idz/9KcTTV88Z88XUagNE4Zi8FQ8DayR+vdZYGb
WNSxReHB8AUJi6wN6qBuV0Q7Xy6o/Bv980RSx2WRkDzY93wF1yzJ+s1MQF6lj1Cy/diBu3ZEJczp
lXI01LtHu0R2Rm6kuwuKcOJ6/a9bdgN2DRWCiaSKz13qpBYhj0qTCs3wagPMHj+3kUjoYRiyrfOB
oNwoDxg+driD8lJUtJUo5AKkAPEN9SPGvpAaz6Q6jZKXkBxWJU5+vZ+OO/wxlTUjuprp/Sinj8+0
GlXVwXkfVOv2jHprMLraNoTtE+1V7HnnnChyInhAAqsck8bHKu1zS19FCIG3Ey1JmNOceLcEMPCV
JYTd2IE1swwXF6p4j5On4XECJmZ/SMTTLtM9rr+1GTc/BBHRr/Q+J3snVIA9stFlCCwFe9ZMqyW4
6wDO6qms1ZBHZDdSHeyC1anqyeTEt0x4ujr80+OkSlrbEAjkwrQY5XSmXMQs3FobuLdnHQpF6Upu
6L36ynkdLJemgwPdVnpTOIgwB71nIF+ZSzq1jwmDv2cwTb3HiUBKWdzgElpKkNyOZ8+IWS+WFnPB
0XY+j+GL/tTEzBhTgFEDAPU4/GbNSF9XH/s6EGMYxIMApgfp1xG3dMGk/mFWIirq+mHcIDtU+jIJ
6k5BPifAGoFdV9sGSPD9nxCyJ+Yw4bySwC/pZ1KNZ61xlwgGMOgkQ5lrXEHIOl/MbrKwo/N9jJoO
QMuMvTm1pp13yzDWnQ7/mt3K0aUjkHz9xgCn2cNKEsjZFO6B6T5PHi9bgqYFXx+TmXDk0iQM4neo
8e6IP3NBNet8ctBbww/bDCxpEeccTPr0xnkqt31j5F2h5VMivlfiziCIzWU5s9SOTU+shhiTt7Op
bab/w0NyzGoA3fEN4REeK2GB8rvrQ/gJglZeymMK7qltoeYU3aigCMMucNOJDC0JnRrh+eDHECEf
Gjj3wyiOX3WJQrIrduoajgHJhiVvPx6xnMVl/HZ6laxBrhuuyy71VmlJ/9H7oRgy4uqyirWKh6ud
MiiVag2eXeBCnFDCkxBODrEmPNJi7KjU4ltwJoFYbc/eiTZPl2GTh4U18R++aQkR4BhTTN62lG0n
EgqR8LF+t1KeBAJvO/mxmtK02l8liqsPM5kSGwnGxgDohXcfQ4oTqPcQ0l78CdCHZWfzvFPSCd69
MO8M/o/dKIsuWNS6HtkbmIN01qMp9VEL+AaFpgReyebHnA4fX8BlOZkEdeh/es1FeL3S+6lzLWUx
HzJpSNnsTiKaBiGkURrK+QDiXXhC+YXxEoxeZLKb2Vcgi6Lqpdbk59PJxAr7Os3NiBmdSNjZaaCV
KNZiZFC1LIh9vyDu2GggxHbkuLpudBYUhimzJATwyfHbDUbQ1E1jbPPFV6G9bchmpTSKOJw4DWPV
vZqYHKWaOVK6+qzHWASdpjgb4M09OaTpqZu2tWthmmdWAOcCtu+XW/lc+kgOVrR0hdZ7GQTvKdo2
B3hqrizJRbMjOcNTUHc3zCAd52tlD15zADO36J0kUuuS7IRoOLBwT4W7k9HAS3kYwe1CfbeXBUx9
YR2YiXm1mWkLW/FrsLCYt11xiSjzXO744dU+ZHAkRqLvYVi5emIISYNhfXW4+5lRCXEnCwi9ur5a
ywaBnjlRR7Uk615NzMSRsjqS4cxg96r49mu+XSkuQPyMfanFQR6S+C6JLHdRHh9dQe9Gngy1qbZj
/EkDpbdT8tXyedQbINAuCYKTIkD1Ev8BpwSWNF4cQq0MwKMBhD2/+Ij3U5fgidcdtOrqKSlxBmX6
Ws+9xeKQ7aUx1+Il/pyiY/JdLuEtJ6XEuolE1Tl6um+ErCRH7e3PD1gFxKHwui9sReCr9WbEniri
DOi6nArETKutA4KBnqOmbtdkM2xmrU5STuWNg4t3InA/8eYjcd569qEe+Av7WkmZR/OBGoGHOtP2
rcm0PsrAfmX+pjqLoxc21b3k1uUoWTo8l8WrHhbm+1TPah7yZFqGvnZv8ZJGyI+hemU2TwlrJ3HE
7q+TzQYwexdzymg7L5aMJ+ZY20azVc1wM0s44rC6KdfwqnCaFhEx+OVVyUGtT87DbLZJTrXiLbL1
ISc/ZC8ULyM7SdqVvlk9qeeu4GeGlP5UeUMdBUE7evhwnsDZjh48++uK6Wqg0AQfuTC/z6hY2aZI
1v78XbudlNzJn95LTMQycW7vRlUAg6vK9pRIN3xZ4/ucD328Lq/msiEV6F3k5ov89UmPN1VFoNSn
3fuDxhoLduHjZe76WbtzUF1ZcfM3/RMM+r+/DJrqaOx9Xqm+AB8LnwlvytBXWZEUI3jZDrrxtCLy
bXT6M1QF7vT5s7tdIJ7+cpdnJax0c2k6tO0rQSN2CMgH2ubCH+GHnNr28unJA1Vk5m9lunhadDlP
ZYFvatoqPIicAsSiK07lsNPk8xy7T2U3PJfs+TRzU5DRkrJgBljFm/zlzkVrgEQKopP1TCe8B8bX
t4iOSwVOQ7njhMS4s9yqQtk/s1mlHsP9ihADMr214oEiTg6r7WVoTONcc/YILGOWVe0X+Ml6V0+G
c1LWfLkY3FNxj3SOP8h2BxKQslFcDiVDkoTw+hlBjgItN3Q2vZCWjcuSuYCScB2XePVctRztgqmQ
gsMqIoCjCAgpSrukUc2briAFCuMtONM8z2RQiy9z7RFwq2vYJ5gDD+ZVNyRd3A+BY89BW2qB6Fpa
CRuRBtVekbVuRmZxOwtZunKvxwFIrCJm8gzbBgo+qP4kFk6xMF4HlHSsIVCJzskoqSvTI0VIGcM0
Hb3SZLk3IvZBn+NhMOe6r0y26y7rDreWmTdLmrpgSv34P9vx5r7AIsSiyCJfyxWB7GLrQIJNoZKN
uMPt9gTYTSXsCBpIN0Q1zxYKQClJWUBXe/EOlMSZAWhU5MgPOm4r9otXqn2qzKO9Azh83merYaDH
s3UQ1ZOTsOXgTXuuwbWuAoFWNElWMkO/sRE4rCQMur6wDOeH0/ucDB/2QdpdipkOUlLH/F2c6Ypd
wGbpMMQldUgZ8gCEUu7kHqryL+q7xZ8cz6W0x4MfTqtyeGYd7pJ37mS9Wy7gl0zUnKNEYFVio65y
9FBqOXzln+p7YJEPubBtyDYwE9f5s4NPrCYYHxqe2xwv2d6jzRCOfNJLp2lM5fz4xutkdwtUfbNZ
ryKuFm+nlGGYBXV+5oVI+TRuSWIehkijs3yXh1oT6doHQCqXI+xb6qNv9n2k7psFjunjNTGpFgtH
Ij0B3SFxMQGgINmWn0s/Yf2F95+U1mfmsX8q1KjyRcQfxBYwFFmZoSLfDNrLpQFgMTc1ED7W/+KP
5Ys/BZ3TIUHoYwbRN6EO/O++ajEE/rB5OYnqWD5nN71bi3ijDfSMEBKATl72ZZYS5y8wLaQkKO6t
jJZ5H04o+Gd3Ur1jbf3rBR5XAyPkrufJB9sr2Bcaj54ef7YNgpqNVrRq9BDZNgxs1vyB7gOoZRIl
+wj8AJ584QJXLYT1EbJKLGXeRabUbyh7QYRIf2PIQcWJ+dMnTKH9Tzln7DGnUxWacbDVsdvV3qHw
OfdudYWYXZVUKXQ5OPzkzuhbiNV9R5EFmJA4nXRcxFjH538vMUl4xrJujySPVgHi5J7N/iTCLix3
gW1zCUm12fOc0CqXSkiazvWbv9ZSDbJ/zFy+0e4VrHzeWTro/FywLyau1iSUT0u+Bh5du2k/xzV+
4OXTAcASOxJCueKqiW6GywL/VV6tLBSKXVT00EyunCuZwIe6NTTIgL8fn0HjLdWk+qKXZmd53fLQ
h2P7rjFuf4YNGvdIcFacgIi9207magvW3fChFRah6lUZhdpjHe19QDkw/OAfzv6mXwRJ3ZkJGucO
F3VqhthLI7Le/MG+KwFIUDowXUNHmyXJwg4YyaFaVm6Z0q71dVc9lvs25VwAO3YtocNEDgoeBUub
SUiMZTUtjxij3NDxNR1wLQ1qr5btUdGZPiFTq/xnjyo19eHNHuFFPARA7Z/0nd01OBSa47J3l+U0
mtw1elMFtl1xEGZe5SvqbGP760ZchztGoG9oIiWjP754JXZEX6hnOAsMIH2re1ZLeSzFoAV+u1XT
AIRaDppHP7zhcQQMxQ1Ksio1HEaggT0zNFZ9mruUS90Kp4dlgLdaWwrF9RLJBzeJZXzKjrZDC5bV
3OkK8VXRSas6ZaPzCOqg7R6WJ2Qg4Sws7v4HVhFV/GE48j2Xh3n3bk59koaLlSVA/fWEuFmFLp39
zb3T5bmfCX0goJTiftvG1qRRP+KsifFXCfGuRNFsIYAu2lMBcjzahhntubMM6e8KxEtjyAAefL+2
ah+KhQhICGbmnCLRssQ6eb2Z95d4QH7Abb5/a4M2feS9dI6FQh4C+26l2/JvOTnq1gLUfA5/mQGy
/vpwuHJueJ2EiXlGKzzQnFfXVEU3wFXm571M/q4XfmzlqOXV+4ukKlR8byGOExKJqUqpwSsh9qGV
S0esSNVMmB9AWULXHBueZexvOhd0Cow4XujwBYq0KtYULmtVPzju70hRFzqgmo07kGSTKauZXLSu
1rCOZTUggav2OLEa9DOEj4vZdvOg8aP3/51CkSNPaJTO6ys5J02RrrKBqr7+sMG22d8jIsYYdvI/
AJJzUUeqxlHbwRpw+Vyc0tQKztsVAcVVVMp527BG+5nBGo4yv0xGWSeZi+mWOLNmgLYEuuyetJI/
Y22F9vH87ShPdQpgN0ZYIUBoCtzys458n2TrmdDAD7mtmMPpFu6wm1+tH+we/PrGf1zfFyT7A8RK
xBUeWu8lT2tarTuGxMAxuSd48zt9Y6gNL0EfjAy1Ze+HoXpDZGQ/PVM+v4m6brOAKccURJTZ6DIu
ZpGzsjfZNlPSYfCvy89yy4Jys7eeVHUhhqiOriHXhLdX5NIJs0YkXADchvHs3veFncFKBmFZJPR1
0Le9zkZsAd1BF8OTN50ZdWJqApk0SCAYEdx0J9j1+5hI2YNJo2n+NdQv1/IJT8v3E/MvTBOJ6JRr
6u42xpKF5EFSB85EcGREqqY7MEloys87EaE/mi8yxFiC4tw+Vip7/fa/CcXHvqqRx7Yofbrv5PCV
m8jozvLRkU+eh+TQnopqAbGFC18aV6zNm5VJA8I8QDgHJBMPsgmtmaq/UhK2w52Q6WC3tA5jd1r+
A72SxdAJAOW3fhy7iW0oONY4AOUb9XSJOAxVRFFPmWaHS8jfvxztSSqAgOEgaBJ2sRKd00ChrJ97
4TDPC1HQRQt31js9/SVJhfaHk935OsgZY1nX0ncHudtsdVng57or+BehOKHuK5GhEwAkCaDGk7Kj
RUBZMupKXW15O30lnT1N1WQyLhJOwjdEl2Ag5pSqnuO03gq9Pz8ow4nrArnNGeSGWr1KXd2Iuq1J
UTync+9Lims+0gfcrwsJkm7FGdjPqUDYddzbXx7ymfS5HYZLDh4ecSys5z08Y2UUEvdlQ3fAMae/
RkxZpKG+z9ZdhCApcOcRkFKuEqq23NDX5JxjckgNH61LyJ2ZNIer0Cs9aPhvQ25eistw133QLEdF
xmf0lBSnjCu5uQ9djCzu9wILJyD2wyATJc8v2PPWZlfQF3/A5wHfFyNgWWny1fvr193QieI/EJur
l2ZuiHc9I5DlJAIYJT+45tkaN+okNniGI9JDgbbVmhJtNpiD5hdnbO3euiIRFCpjEquZQoSQ/s9y
sBGfN6BscjlPa0EX+QmXl6QOtpmgo46Cj9VYG8drQo7GCd+rTGVOQv+6Dck31eGc69XGX3XZ4OHF
5GmTHR87P6ZMVFpuV9LXd9Ai9v5M2WHwdA9x5vQJA5uoK4Samjozqj42zm6tzWo0vrpbvpwufP0n
w7wubx/V2xvED7S115eQjeqg5dRjA0grW5O8BeMeH4hFfD6i43E/EAzlD6bsJtHTFyi+mWU9gh32
3jGjMW3bKM/7hTyR2tARgFsUkJ7Tg1AnjWqay1ad/e7LBvbQYEL0lR8Hbs/IBw/bOYLBMEPJny7r
0D8jNJ5C1VifvZCUCTQbcsstK0tAl6ioaRgMIuPQ8bBNzC42unMPDYl1WErC4+csLQ4NV43NZrdD
v6kyGTKbMyD77gmbIu+hwRIXD66ORSuDJbTFmD2dF2VYhqj7qJdfRrhh+vFADlfxVSMArPalo5JT
VEhFw5+gKZcKC6fzN3cMH4MxtT0lVuNsmOG9Oa7A8NXTwLMJAnDdrGZ7qcZmoejhpVG7Rbek8P+T
cJsgKj0QK2tEu0RexCUckluMmkq4gU8TtaOeXfSt6xCCooF4OQ33QWd6sv9FD2gW2QHIO7Jgp0LR
1ToHp2ygl5szifTRR7BtGdKDk81BkyOonMTWMqnBjIQE9KqcwbN/IiN9BlMD0+Wvyw6ssndISZb6
9aLpNuiTatTUHk6uGBZpfkkWBNhrnmym85TZgmwlFL3t4rcudlo+GAQvzJU2yv7bKJ2w5NyJ0ZFd
+r1nGmiGb3nn3mjhUttDexnX8kFBNTx4Pa2uMSFnDAX3RAY2FzCzb8CvmzaYJkEK9EXUSquq52JE
1k5LX51Wy8wp1493j3gBHRu0bPWRayBKH+1NSRzm7Bm7eFhGf8Nsl4+u1pY5t3wMpcuyu66wWP//
yVkXB1pK974CQNN9KWdfBt/EdWMX1n5udnIKuLHJL1cI0ka/LPeTbOdUubAcDfbrh5lZEfHpfqfu
VM16M5PbJPH3e4dOzL+G340Ohv7UBPEocJwxECLjtN1kI2QQwXexesbn6WjXmsCdQPg7kjNkdtJN
h3kFz/BoJNAgS7ihLzWhc2jZk0NsK0P2G5KNvJmLYizdlcJ/UPPYBk2c4d+/bYJe31t5dbkDMBYq
KmMta8jdKvHA6PXd8PxwNHTEbO0T4uSaqckuFaGkUEj5/snB9XsViRIe7OUWOYfw/BRgBHfr78z2
onVp+CRjEsg7p5JWYlJMCgP7zX036k+QHZ0EFESd0Kl44iBU2e/QfpXCEm8DtWTP6KjRJYGlzSOe
eJdR8XjJTZTRJRPwxDa2IuaR9Qbs+PBL7afrViQjR2Cg3cHsVPOObNXELVgn+8tz44vSjjwVqImc
aEBC3IoJtasyVkHhqJEUBDhpiJBhn4vee0UOZfcUBQW3xG8i54j9KpttN6oJa+wiIgU+BjbRDacS
+iyueMoUGJr09RgK/LNO5Ot+doB/VGhizRD8NFC8uMiXQmjcLiAV5MJ7oYLqcCKH1EFKQRL8yJfa
cd+40JZUaqWaLWQ3V9ZDjoRjHz6mcDKMZ7fnvFK/pGDeZ+ypT+Xdq//8SXSLZkOa7GT3OkbRXXhn
ZEK7Match8i6tv6fUDPg0PSAPT7MXDrMHRpucKKlYAsRbReGy1NQZoPJpc7P/wQoHsiZDzAeU0WV
6eK70MJY89oFTdXQPePh+owg//pYytgOBV7q+dhEENcS6qxNhLavrHD/33wJqVdFQlxM0iF0f0qD
HXd+kmBys6f06I30ZRYu9ZZEIBdNlSSLNqb6lm7LRcZz2xyEaD7a/5HxdZi/IgpfRlCtO3QIIAM/
JF2ueo/fQGTXv7ivaKMkj2ksupKqNFSiurduj31ZcG2sTqCBMARj9dHfiG8wbL7JWmV+urNT1+Ck
h/3tb42cD3hBww9AOuBVVeMkqvUdk7bjAxYgSsfBZ76gTSqsWcSjjhhS4r5OjXM76BKs1Z2Hs2tR
xPpC1GY5zjxtuyT1VYnQwQYr/V//ChKo/etOcqgJXBBHe1tJ5riOEyZpTDhqpJUUGV/sLMqqkcYB
FD+uTlSlTw2PHby4l4TmEalbvgNDoIQiq1P1dmLziTA7sNWb4x32Oc1hBSeKIW+8bGfu5VAYj8Jk
Y3OjmhrLCUlYMh2cgamzEjTjTQed1FkXXvW+iSzfHHdtlxOjNe0zHKORLu2QkfnjDzMsFVlWwBp4
iAvcTAdWjqb3iACE8CNp/jQZXDH6QyzbVA96hg/FVsH6Y3DPZO0lm4kVh9j9MHZ1GdzI+Lv+FSfu
WErIWYusw2n3VQeCmeo9fONnSIr7osC2LyjCzzZw5PEjYNnibDwSV8FTBRIk2KBzDpVekqndiH30
Wkg0yiLyJOngCqXQ2koCxlTH8pSr4ybG3qytiz/zb7D4nSjJeS9a6vp2tE/DcQ8/xnD+9PUM86Au
7u03HFdd+jwHOnY1Y8Wsl2ehBb/5ZizNq/OFwaWq05VzO1xa6S6eJiIZvkamZHJ359HJkj1IPaEV
oAM7P8vc4jrP3VCH8LnyvWRhmqqIRZPrvLOspbzypVORx0NXxP0vB9CU+PBOycPCGWxjAOnOACxZ
FWMHdU0ECUKx/fCS2Xoi+K8k4UlzpAwZsMLSm/HKqcWQFY9R1RQ/FTwhNdxveyJ5IHfGsQfKREFD
9MSQh88IZoXnQAb9qiG2Vev61yd/VkL4XJiI7E/O/e2EOQvvszDKqR241v1fiQz7pw7QbM0fkTkN
p0tIJNNa7g6JZ0oRCr7zT3q7KzfpcoD2xwNx+Tc49BPImHH1TH5614/8E3qe8msnN6tUdkWy99Mz
SZUCwAITI/YnPJPDq2CP8LbVUYYI40NrOleMJkiY+7AfGX2qE+wIop3kKGUsZHUdzt/dVEBx1zXC
SGKILbKYm5nLBhhcs6skn3s5fIohvSBHXgkejH8JOH9dTG5o7tTJJX8pp5MVP9Ky8iA6nTnd6AA+
dXbULiRA2WV83VerprCwRmW7uk0TTW22RYxDSTUs2aFWydhmmqiLbgUXepz3K3A9fHZXEQQ3vHr4
nRK8ErLpeR+yt44H8uqhwoRJ4HyF3mrEU/iKKdWSP1I56fF69DvVcD5LOXrg1k3xm3OvQwPg1N1s
OCd1DPwtQu4TFKwTRe3PgG4G1qm3ziip20Umv+MiZNOTw5gHno9kJ583aXnmHTEOYVaPnostaRVb
aGwBgYBoCwuqRmVLMXJFF7A2HtyQD9G1Q9o5rU29gu4F0pG9ELlGiKgplw6IuUTxDovP/OJChVrj
pmOUAJ5Axzhfjgs62nhASqa7FWsta+twiIjn9aPN65GA9Kfp/uVdndwN7BnMjk/8sPrKtl2910vB
5vZ9wqrexQLFYJsFSz0SAN/AdiHafBQv7Z2zd6q57C2oPR/TV9A0n0GADyG4SecaoxJOkAvpqY5M
GA5WVz61OIX027nLU2i63+P2P2vqQW+CyWlOSDaM9aLKDqPEkFBZkP1s+zmnH0mOdijXhKehIlxQ
npm3cOw2dBvPymKOVkBstYY0g1xZelJMby0ZBXSzGbWbyWsTHAQ1X2hcaM6FJEbWNgtaPZc760vl
ibMjwdh4mojyumN5RkTCUQQA7cpUHW7g7V4WZc/AhKhDS++9iPs5xEKOaijHsSPxomyQAtElOjQe
tOushdohYjBQH2ogLtfR97FrhMRCPPu03B2JsULjGPij/v4YiWw/jfX6a+lOCBk8G818KjI+k36c
dZILWij/RZM7lodjsds5ZoRog/L+YVaI2hN+WlNOA28wref6u6v75DBxewBhOkJmUB7hqnFMOPfG
XjB5iwLiy6xB2x1ebyVbwj2DJCj12CluHk6HwqsLN88foZYUmkorVsn6oEs4hFmk9riQptuHvcJF
lzzMhQ10pT1iLa9NjoyE7UA4G8xFeSVeQgZSGEUGMqXaOITsPFFrmeo7e+2l7AgI5UPd637U0eEd
QlEF22ISnFmmN3rYKMyYBdLwNtmNlVdmM1EeUKmgbjZ93fbeouugVUIirkxulQcTs4vsKIWggHiV
oLE5zPOFe3LCb9acdYC1xq/yRjKYfR84vfPJDXT7AADnSOzlSR/VAGu5h7hm7VNTYqxEObuXnlKC
VfMC2eS0wIxZ44aSgZ+beguMQ1YS+KSrf52TjYQoYRpSTwdlSLrWR7akzc5h0T6Xu98zRIJRgx3h
20RWb8m6yz3hTvAWrwFo/czsYhbJfXn/SnSPQSUWTi9DCQS3Mg8e2SDTDykISIB/ZTDxlSOtkUlU
JXNnxNlwDi5+mh0PfQtLV+VzDMw/hnlzmpsgE8RmcUx48UefrGF9aZ94vrNFOGyzL8Kz3M3DU86w
Q2W303+nLtp+pZxNpgZmtzZupEp4wopjPNOOoaQMoA5KvYxu88L11Zc3Oosk5Se8whM9VfRYDxQY
LBOPawEtPdnASqVBMtcMN1Rx64l6IJpJBwWKdxttazu25UBPEB9+mE/G8j8GFBrzlO40CdjWPxuM
evvo4VGS18MGtuX6AaR4Az1gdfh3tCpHw9FguaxXqDuSI5T7+8zfZ/IvGjdqFzfI0IDGPxasqYWn
zSHzEwv8RF4rWiukS2Sg+f/nADW8P0OyrcbxAqDuLZWi4oBFfPIke+xyxUMQVOvGIHUDdzBoomk8
5p/AfaDxCOneKpUxv1k/HT7DCOFy4WDZ1IRentn8BGd1Lg8hM50g2PGzUp4KfZmnaajeNBE6fyim
2Yygk+m2vlFXd9lHD3i1yK2PtgVNd2J0csXfCkPM0VWLDZ36O7jOsQHtk9pr/x3s+Lawif/coYfv
u51GHvIo/S44wikpkk9xMuD8RB0/W116BVjhSU+5em+nz6iBCywSGlteJrquPjhIgNKA3lBO8212
2k04S61y5HLTcl4We17kyKfSRVGemG4ln5gjW1dZ+g39jb2LlZQanDv8JJW+1EpRmk18et3OfJ2c
Ynf5Ji7mzV2pcS4gnmdJoF7LdonYkY8fK22WiG7XYxzz+nOiLuDt9To+mn22rbsLnDhK9xuz2TJy
8KIHBo6UGALdVbmaUISNh79fGKVNhzZe4ZUilu/wkbuEUlWWJRo6IkK6FvS8vfn/AxAphUKbRL8M
/DAzWhIE+XhmqXiNcH/0wdqDuGqgkEOarW3J4DKB4vtFBK+TfgDoQVKYwD0QY37tbhQfiO55f/Qv
zq7/sPgc70Bz81V+mDf4d2mRn9UCk1XKUNiTwjx4SXI9tqzcpIJA28crC/eOjYE98JqNE99/2bcv
vwXPVNuwHG4SwMQkd+Ll2d5iZndbnQHMPpjJYFZBDMypckbGmC2fLVU3qLfCI1iCCfsP+uWE5BXC
kyw/W2QbvKLBbUzyA+R4WDmzMtFcBjHhOGDlKVvpLsGptuvJ1cb2kSm1L75obcfVeXyq3KlqRKJt
tbVSskRllJWGRfp6/NOj6yLDJdqTlouwQrsIkh5JUDdKmH2z5AmYmPeg5EG8f6VxWxMaSEi+xvI8
jtYOsYZh6QBK8D8uwoML4InOYw0vRdomohXXQiA7Pd1xY+jycWU7LdTePzgF2CgRAsanN19sv+Kl
+1mKJLd0nSpALHn7jZLuJO0BCYuf8rKDlORYV3+t100eU7fporU+J3lzv0ChatU5gd2s8y6NtDdI
r4CtsZJAkA6w1u285Xo1+oWxa8sitXq5/7peulOEmE/lrPcr3ssMar/RDurqutNqfd05J9RbmEQp
0yH5d86OUImLE6Ti9103q2uMkCjKqdnHe1S1rc904fpyXu8Aes1hwuUx5Uzh9xdX85KHJB+ph8zX
nrwNKEivje4eDFByj5kJXBa41SlckRtCB2LX3cKzSTeZHNxOvRue/eYVziyxiwV9rna/U5FNukGe
uDpIuOjOvvtlTeUnHYNJjX4qAy9uQGupSLcyCu9Z6Z6tdwG75Q8CGlwzHqKx7EuFYB5gqT4DLnug
0Iyldc/4ycCsptSNqztPL4j06lcnvomlSFsIdb+Xp3PmI6sGUM0z+MS2VZgXxmrkJROnt5OqjPvU
sBYDu0TwL3B2AErqG4j3k1euSDrvZIo4yLi0UFsT3S+sINZBx05wU+oKIB3Ozs5IINxv2B13JJJ6
eNoTf+JymqwpajztI2VOrl4U3M0LDbxd4butw/g4ozfist+yUPl7fRrgHNHAB2j/8WFoPmFZgira
ATq4xuArFqc65N/IoPsEao3jCCRD95rOtxB8vU6WommSYZjaEnHkL8D0pxrauC4gt1coAn+WCH+Y
HbMz4tVDqiOndZ05dONCI+WFK7J4yrJ8YNpeDVBZFu3nv7fp/tdfNR0NdqUuXFhDu7oqQfA/5+5k
BcBL7zqy1nxJfeV03wk/WMED0wadMnm74/GNhx6KZmZcBgjfr1K4Np2a9E6YTBcaqzy/0++JRh7x
J/+2JEflsejEAFlRqtKnF5yqO9YDe2YdfaLcepFkCUg5obzhCj+AgNcPdjBfo2SYJe4c0eSfdBm5
q0F//z+ifNbjhHsWx6StcWaWpufssDl9XtSrj+4lNNSfwwwvEpGb/If5K8rATgi3GAbfbd6PJH/Q
IAU2zb7v6d0J6/xrZXw2WtiFlxdZiVyXQ/iGLhcsj9nqWxp9Us0pp5VvB0CVbMpsExJ2Y69F7d/o
OrcTVfXJeoaxJWV+dg4sFSV6TXdgRmcnSYrIiYZKsl6CYhVrztb8ulzb7ziKY1h9SoQLf5E1VsFC
zTcvZG3wlyoH7ZDFwdgJMPEwksfTxjwWTaf5mHpQ9jrqIzO+Vq5oa+Dxsk2MZl2J9K6x/tFjn6cu
3L6puG5zRAlW9oO9IjqFuC4n0TjHbDbMmO+iCaZX3+IMmUwquBK1wBkLIAKmJVApkP612zEE3uOp
BB5xkEZknXCgjfIK4abgE2j/c3QpWB6bGnsRamcQ3a1KpQ2PvMwOVttjL5/D34hJudn0QGoKwH0b
ClLoqV+LG5FPEl2W1eByR90fl5XQSgI5uqMQM5IImI79iTzdJIbGTPGZGsLlGd/bG9I05zfQbOFW
SvYkSMNMDsH9pABAzuWgO+U2CBlyE2STODcw8eti9SyEeEd2/XB4W4DvEsvNCjojvtKNkOREM+8y
D2cszLU9fJkzf4qe9kx/OHo4HdXgYMRduzolRCpci2MJ9S0akEeGScIgDAcejmkMaU6GWutbQwyf
BAdHc8jDcXQyLz00IySvUw3WdxO8pKNddvFT+AT8HCDgaX2k9Xq77uC3SKh3Nsy8JyTKsr+psVQh
llfOOdQosT0TwuC0ojRSG7cAlptrFqe5yVf0L2bmcUrMFcnyhgI27KZDrVruxIfoRI+cIx++RSK2
wPM5aYpI1IzjMR+g4cK13FvluZze6kp/UT7+30TpTTGHVL8po9/r8uFD7MHxvNiZwAtXI86avs2B
Q42xmjcNxMebpRxrVZzNBWDW1mvH4OjYrM5a9DnuU4l51u4kowQ4fRECxHCoeMEFQmpPqsCZUnH9
Ginc604bHsxy6QdGb7zUuNl5bBBy/QSTSw9Cot44zLzpyn641N8pQNgDIBolFFQ10jr82SkYCh+y
F+nAYOTINqve4sKAddUa0HQ5VKYsREzsdtmYER/1qfnNap923susEyRVFnQWhrpLoUqVNpVTX9Ta
Mo48C4kTtI1OU9iElsc6DYkro07rtBrkSpCimP1ia22UnmQgts+17F78YJ6TaEj7rN6GX6NsK9RF
H4Afph4nEfDJ0n11B96/19s/kZ6Q1kMWqaYhMKMbyMPspu0Mk9LH+cg4kpufYp1IMEjsk/KElmNK
Ngnzmf//4mrUR2NgJ8ACrF2UFRsDFBOrOpwwtOniB0efLmdq4ddlUnbaiKOihhRYxSqX1a+Iyp7c
ljG6QjSBN74F8IbWcyoXAGmAsC9Bwd1vKfZv79f85LrA1etK1hSji8lWP2O6Z7gRfITAJkdgJrXr
JZ2b2fjRkMdHG9IcJUdDIVbrJ7XdD2nYWnqGUnGaGhAU5wk18vbaSt6dEGgsxlTqHr0D1z4f/oJw
vlbVY8U1tpTWcSaltiin8rYKyGSAUDk39d+MYw8rhXeQ3iaPwFhAyEehnGDz8Q+roNlqU7EJseIg
X0eb36HsQqXVK/kAIw0M/OLexF9GGOkpUHeHjJhUnAo7jGWdwa4KndZFpTKsaYSyORD+OOC3Payr
3fEfPQlM1d4ZfAGZAF0WrAav71uM8rDng9FQq/61Qob2HQJjLHhcldFD4sLzoIxTD5hmpdjjKAhl
b+aItE4RD5FWLq8v89pIziQUAJtifxFvGy0KHSWfXXmKJKAB+DEDcR7zumoHAcbapdC7Qp6DgGhz
dxAOx2JT51gCfuih52PyhokBeK/RcwHlJjWAJ9Q5boKcqP12ujsBupgD65pK6Efb7f6Lk7m0KP4j
Z5uC+HGBi+uJHD0Mi/U045mwq9ur3zBvEO8V15zK9gDrnd469xEs63S+g/ctStJuqm62EKNJdahS
+Z9jiPMA39uiRt54FMzGNbh7clj8iylxzlOIwzGO/M0MXLOHEizXZFbluzwdFWFwRASDmm8pR/ir
1QsP3jEAjfcA/rh50ZQIpmEvsHxZ+33Nh30tWvn987VOBb/7MS2+mdNFzrD5Iv2SzZygKqdJ2w7I
wf7djFGzr/pxwCUbvyCsD9rVGtaqUeHehn11WrvEDP4WQI291h8CTlKsHJ+4+BirDtCSKylJOVta
M4IEb9LD0z30YPhfoNkehbVKNzphxi1LMtidc1bTEzqi1VEawvsCVwtmrHjv0qA8AtHAWXri0pL4
2N2vr3YTISW9M0C9f0KMVv6T/KWpxqFxGd2HWCz8Re4kG135xysx7InxirRzhldQZ4e2vmggqCHc
EwNNjfv5O/LAjLZcK/sZwghvFE1BfjVUD+ElPW8V3ekJlSGli+6xrtxkjqsTd0Wbt5JS4HJJedBl
jDlanfWNwyCb0YXy1Vj+jvemMF0nRMERIQP5G+DxuoO9qeeE7VgCa+ZkqItmXKjUZ5QF5VpfILJK
VkyW23CFyisM8gz7+rTfUCXK/XgHxduYx5VbqnMU/xHRJ66GUVulM2Vl82kvICxCogmQCEPFGbur
eefSukBL8wG3gHFL9BApg3+GaY1YNEq1eRBUefnMFJ0lQkcPZrBy9V/ghb6BPoqaUgQEO6viCp2H
O00QGpX0HiSVTEkdjiVhbETaeV4WfIiTEd1/wkBd5jtP3YysVTPWBgSsQHRRKwoqL8ENtDbjzPA1
WQ90KBggn2YFxrgzfLipnixOJyNcuI/49HXT9+6nOtzivNtbFJKkuco+rac1ZoU6zJH4drneZMsm
aLZSZOYWiZfYWLdDSJfTX1rUyx+KOqWs+LIf0RBwmmY0R24DdlSP4ZQ/fMOuaEyicxS8TxqiAOAv
B9nGVYvXqCIrB/mv6yseqxyVMvh6xoer+JYIja9lbuopM0ufTIFRFJXUCM4+K3cnuyC5ePkb9ibf
R/Ok9sZBHr3JB2h1g07/69NMZ+j83uVJAZNtXQaS663gpKHdpcRcaAXaVt24v5fpe0CSXv3m3YSM
+STwhe4L5IsMGzKbqMNBP0y0sp+uJ3hNPytwTiwVsJ7/b9/tAqT/JMzxHUiCGL1RY/KdNuLGzLUm
ZYWPOQmPcJ6VTlABC68ucUAfg7Agq5Asx/jJx49Z3TkMsO0tnA3+N4tNuCoB/UatlAGXStH18MuL
rR1vg/a3nTRqUIdHj/haM1MjGZdVSruHG+R+zIYaNHyhQ9UqpRJsGZWVLNG4nGCa/rEIcRE+aGzA
libq2LoIo7DXqfY4lRtaJ6J8jDBHJ6u1/KGhmJ549J7A+Wf8OgChuleArYkIK/30G14bVY469yOD
1wMsMACn+AliwEKUucKl7c59S4/7xXvubT8EOTLjyliA47fSL0rXVvZtmgwJj9Lu2/Z46eb1I1jq
2QX65/xgRgZTCbNtwE7WjcVyyBAc4vjBS1YBtTi9ldUWZVd0fgCKuaxhO8pea6XyUmA6j9yNlp8I
Sp9vG8fZaleXjXZoZg7ziiHef2G75RiwYqv0rMmOtsf93ZCw+20Bq1BSLl9b9ch8sHggS+IPyeUc
DFCTBNWuug5E5ZrCteLQ6kYuxGQO+GiDZmuvgiZMnPbHgXeDgzfWkE5MgWRykSoxNVQBiDmOEn8w
/qUkyTt91uTi6pOBw9MJ8iKHHatEKKVploswVyZhz2PpmCnbwJDXRSzyke0Xyg7MVwSB/NEOnMnu
wDUSpko05rtp98YynVwXjAL68MKvoi2MVx83J2hgSozatWbsl9l3g5Ptadi7KNxea3DVIWR18hy7
t4+baTDORfF/izFXb4+Z2BnO4nG5rxR01g/blxgtxhKeW8zci8y+CpaO/ZkweHqY4UG059rfJK2p
wLPxCozLSl7Gu/qzjRxQzjK9W6dQ9JZ5YRXaGWo//yFAKSbSsggi7n79YOreZ2KHmLzysD7NWbxt
D9smOmJz5UBSoozora4WDEAn6+1yGult075/xElIzd2Sd/oEcvtY0dpT7jAp0ILA/AwAohJVnGuJ
1pd1DivCv/XeUt2cwqWsvMNfbRmtAyIzDHe/tt4jPDgs5/AdPhc6yPbi1xKQfYkLTP3QlvF9B/8h
wNfJ7kBWHrZ+ZQHpLu47tS3hE/TqAzbCb0T/+zglKheq0p1SpeZiimbJGNw4GEIP/O7bD//HyxHM
u5C7I5pRDaym5Tfgd+ekB9We9wFOo03VJS5BRoMzSSuEadoreIlCJIY76EYvfeyZ7FdNpTeiVpk4
SAc2zBSg/E4M3yYiLlwmUMORurj4Y86MK79NVB6EvOQCD8pNNfe2yG+hKmBKZeuRncy663cxyJqx
X8Mjp5hpDreIzyLXJVfpw5rh5Agpt1RZZ9/iNyen7dKNNld3+EwRL/ZNCJK7lw9hjF42obEy1+ZI
J3YUumTheJ1tTqA9Rna33i0pF8HEqCIWTKIcWiPSMY8MPoJdDcWdcvO9HkqK6ZtiDDtwXQvO3uk7
ZTPR3nycmvWW6K+hb7mf2XUb9W8vA6cRovvpVwuxRk8KuF2ZmMPQ5Mf3eK8Y0iOpcVuvt3ZWt+XW
iMjKules6LNaQM8+OQH6NKbT0WZalOXrPUbIa8Orj4jqoafPi4FFNpSaXBUmSjOfbvdJkhPHgk1O
656iQz7qLnY2HBM2+JoRWtvwduGx8zgz+MG3C34e2hEhV0KyJps1TPTDnavMZt3aAjHuU3+o7+ai
RaphJlCJ85oDyf58OEW2PFS4tNw6lbXv4FR+o2yfvDgaMCVOCF6QqFr7NaHPVR7vnC4NGugVlDbX
SZ+uQodQtt11EabWzUobUQj8AvK3QuU1cSX/C9O3Zq5AYyeC/UlFQjeDjUV5iDunuK1/uo++Snjj
eryxah5qJpbzRl6Yh42D8pakVaUuaF9qNJM90bKGz8eDYt+E1L+Q6FfeIHVGHaQLW5Hsc2buj6gn
mqj2gjma66i3pLHb8BC2wGWLAwOny2Jk/KXkVMCC4mmnaxswd+yuba46MDeeRCtD6dVLamzobj2n
iYgMvYde0N8LzAe07Zdl6oeFNOWt9BDuGoZ6ulArIlWEvRyPJwV+KJF1ajF3QNDpQ5ZrryUpjsBg
iEyVEcAyLyVLcCulZwcrkitZt2QXpUAf3Hz0SR/Vrvz2Elfl7MgvjtTh+IIE0wrRTzvaf21c+9ER
SZEYY3T5gQO2SwdUmd3MX0QrYaRiRr/6GOXDyCdhhvPdbtLuUjQlaP+4XZ6VQtCw+/EBI0RKuZu2
hl7c11zAvX9Of3AIfu6yqDv/6YnLcHRz5FgMb9X6ap5F4+4eo1uUoyMTk97vqEndsfc5Jaqbk4g4
0u7QHXjsEfcuyjFlPChrjcYKgYMP6xNy9eMYMaRZTyCHePuMl2Grmujl/nfdDnXByUJNwplBdGxV
8vzXKFuMDjjRTXjjQHS4XKxZFDbI30QwNezfbLA86kN8qw4QgJ5UitURO+xXCh/MOgx1a/Spyees
+Q9b2FDD3y7nNoKxYN8KoZ38t8flZhQLif8pDMeEwAEayf5EAy5bPdDoTzWDf+yUgCA3lUyG3aCc
fw2kol4XvhL7z41t+9w/dbUvhbX4keO+uFmp088P4B4mb5XuntJ8DeSBaFlpH4NtCjTEoklPrF4v
hCScpu6N3H/ICpPdul4WvJZT6nls1EqGeddYzssd/pcbYLeCi8Ah8fNO77phCpfFr3hUR0SQPKyx
6lW47NMtyYCuZHICW7AX6zks4z6uFg5N1HieAHMXWb7n9tiynTJCQxe9vHLegjC5SMGIXFT9Fd1e
z1fAD6PAXdGaW7FDI7CCgEkLW9NXZkITqAs7xh0qF41duWMb5csyaFvvntx76zfRw3UWMuGCnCOl
+uVmh1/Nc8QHV7TYixHt7Rr4+6GXcc9P/Cl3YrE76NGHR3nFvWazIYQJ1p+JMh+ioXhEtJJdtw9L
pTBCdJwuiv9nSUWaKK+Y3hHfVnu1h/0zufVtG/wiK+Qy2qbdsXJNMxs4RX2pqnH9u3soGA7Evk9F
sA4IFzo3hEaanbfR0npGlWSyuXo4/Y99qRhmeYHz2Uq9DH5P9LtEQ+7zjr3fk73SHD26CmwvmvRR
mOsyS4UFyRFH7kIGxGUEzUg1kUIaasBWLblq6YZEvJk2O9+CnikN1Q0EnpLjMEnIlR2bIlna4RJf
EO7Vxi2K5ToCOVhRmcoKW2bwMW6AfpLdLxErCPiBOYWQh5q6hyQzBMtUghTLabEUEcvTXQXMcgu6
xUmvnKEAjNghXQ0D7lGQqJ1su+BQYJ2FqSExXPeIRMqiPPHn6BPknHrTnOwGH4fXFdxYMDVrwofE
Bjk7iKYqpaS9orLXO9yQz9pA1NSBGthIwOxzfgw2nDa/wUJDPoA5Dr1+y5OxKvK+zD7OVdVsDtPx
8TC+4RsxuE20ovYPjK3Yf+0dkQpN9oT8r1gKN/MvI3XpaPrSlJeUtXCOuqjZ0zMt0eYOSI7o+eye
zaNwMpCmFscgwT9YPEc5zFY5prf7WBvPOI849n8Q2xnNc+Q6HcxqVQiRUmuMdw5rR3V/9G+FlW6X
dNoZ8v8/ZO8TxhO7ZVfjeBG0eWHqeR1FSVAc+KRUIvn4MEEbvrtZMptoOaOEV49P8f2zJC1r7Ch/
lAK0OWSnz3IKWB7Oo9sMc1CTA/JbzFiFPqzJdAHkryRcxWBMye3OjpbhI3kICc9fHypbakN5zrcW
/RzGTIOGqR3arUZ9yxDjgTz7lHtgrareWtbN5WZ6X9jJBFzflJcS5NMFe2gT0frWzc/Yr1DNDke1
A2hUyIhPYq5QDKGBLtI8BLJA9rsdGuvMjibWrr8rzWXYRDEuCWVVsg/7qv0jfX7Ne1mUrGisoWvN
zFynMeVuUtIc+urlCAKadW/bXbZcaW8qxYosXCsIQbeeuf5l9QSKrq+SVARnx1UELk/t8JoajJ/J
hiRyXvJ6qnFjWOlBN8VIEIjQH6cgtMkCBLDCNLtJ07eOxdcnHzxV2nkA1NMHodFbI7q7d4zHGL/P
RcrmYeCf7djJkzluRgGtiJiQa1jS3abKp7nEbg7fo4TAqfr15164P3UJX6aXs9mHSb7wMJxIPYhq
q2FPJN1UHRQvF9ns2nDPq8rbjkDZMT4s/cTuLGUtC/yZPAsryRLoPqE9qkMbgRrbtFU9QPaV8BVE
isuA1gVgOLnvBz2VuV2luu5r9beL7RiSqn8Sp02iI96SmZhynZ1WLBK96W5G5kCLq1U/0WCRsPvS
Z7xIERFCputCj1+h8b/zFKh5drdAlTEC34IkUIZ/l6BWBV1wOCpAOhqhmc1tZbyK6vLUu8mZFlcl
H6fOQEnHpJQSkisgKYxo2Owu3OON7tnCL358SFyvkuy6olR91V6A2tshTQnUUmCAIvSHi+F6aXF1
z54H4kvUFa3dc7hjJ9dNUqWhUca/rGGKTStl778vZS1ZxSZYo80/iVkPNNakfzxlA0crT1SPkuU+
EwnyTkFgDjk80/OQWjCPhM86jVu7w4O7aiGLTmO0VmvROK0QJ87/EnEvLfJAsvdpDAVtTlgFqiNx
PSYw4FFVJsEyGgfQneSPLykwkIwW+gjOuU53sQslLzchxNUART5j82VRa7JsrvkOmrEE5xD9Iei6
4DrFam/Uhp/Fr0aWPhcfhuXUvDytRBlVXRWGh4NeOJLCbXH2serWFI6n2sU0iy1/9EeCUqXFotLo
2cahKMa6UF6oG8JmIIKbaE9r7juZSgUwtM0uwF65Rv+ZhdmPif1aWuNhFaBs6ikbN1zGPdgQqDZf
kmrvMmwlMDh/7JG44+04Am31DucpoUpZxD4462gShrL0lMM/rxGWQU6AkfzGIt4DcyvlsBAF2oAJ
ZGKXrRXjYwLnvTaQh+p5eWkWyyDJLR+oXaINlDagaLNYDo8rOmjNppG9F5Z+SVxBuoLQ5Il9l5rK
qL7roGS/d0xcjBRRauTNWpFmNGogMTx2w2Xlpto/UUdpO2qAUN1bBNhEmcyzUwIeikZDRTUfkaEg
C7r+Puuikmw1Hf+8tj7qm9Bg8F3LWWSqe8yUxR7JOwZ4TqgKDGiJks282WBsjmmkCdFj5VytCs5y
ByOLhRaZjM3CmSn3pM6OkJn41ut9MwL0kg0JhnUXCaal4P0so0ksKkNvSSJKTpzL4QPVf9jhZXBa
0JypQ+T/UVRSUlQqvcqBvOloKzo8mWg2SWVnZ4pYvAe0PLG9GiW0JFJI05VWo8XJp9L7phDIf+FM
658/o1uOXEtkfSXdyxyms8kLFXScAyRW60iho4bFpdz9PLcJNVmeEyXj4Hw4Y992kfORIkLJXb2y
U68IkPYBHgSz9/ltxXpdDc3PrROEyRGXWVwcv8AzfRUURE9K1Xz4xQipIlaHthLTACTtyalPpz+S
ac+egU/GbYMhd+OZ4yaC6VNQQi4kNPDmrhH4wNWNrKwldg7E7YQKptKKprtcB9JiyQm2/U8oMlWT
6MBOqYgiIznQRAmBkQI+aJRTil2vyLG66c6Wfd/rONk2dr0af6CoXrx7aQL93ZhXcLhX15Lx8G6l
vpZfJxIPUXZ026Rq3Ykis22Z1UiH4n1lIzUr0PyZ14+3Y7MhrXJrYpLRh/j/KJjiAe4GdTIpiQIG
gsdQVYgkRLrxH+wP6IeR3Hjs9s3kZRZNctZmMGjGFB0sHdG916lf9UpCbhDEUNt8QVTx6FRZvcUc
XUF/QMiYRXWxSUHSztIHQNHuP1S1qpx5u92mvNf802kCxsGQ91U06REEQ1ENdLLeOLwo+FsKo5ce
9mjBJ7IkX27bJAcHAHFMDIsg4p6vkwgXhKGeNeEsmMZhetFrsjDbVKp4TlGyHmpyseGH8xM7vLnO
1EPDaLIbfCyA7oG0yeWxIMhSgb/j2n0Wab3xzIv1ASAwv5J6FZ5WK+fel7vpWX3CVF8ld3m8Hxzw
/itQJka99vdbhiocB4T+nHtHFXOi1aK52SEdvNt4jLA6KK4Prfnqi+pAoFYhm9bwHrLT4YcICNqU
U+LCkrSFs5mvVfbHTV4L+WbAiFxSgcNbIkF09FeoHPMbBzB07NznEi/8Ei8WrWxV6AQQ1GQZuHIl
VxVpVLRTCfcNfZEYboZnyJcGzMYUyV+uqRW3UN/42j1pmrSDMuuBJAEJaaKnDo+2CUC/MMj2mBng
TLOJHv+suMO3Q9vynFT/S4R5EJFx4LRi4KNdl3yleC4Gu3+f49EG9AxlP/NkJZZ4sxT39WXJcpp9
ktnWgsXFrcg9dTe55h2QLrnsyHi+qWnXH1cOZ3PaNhBbU1jAegNejSWJuqPiaY2a447OBG7KuurG
Y5tQoHXghaNXkACblQcZPQtBGVSGIpbjitv5Or6wk93pStrMeTlyB1b3wR/S4ziYBzf80rbxRxih
mMZ21VzaOC8EjrZsRZThGgbtX3RYNv3oX88GS8RDCGQ0ItwETx538q9DBtcz7ZWTPMmSP+x57Ji8
Oi1nsDNR3X+48ph3jGOAiORIHZNYwmKr/ccWj65Su+HgN54YW4jyBUZ3l6VwNDhWC+vvlR7pVGT6
BIzmME9/erDrAMSG/tQ4vWLoslXyWB5uIiSyCsp6UEqv/G4NVJL0JMu49AEb8btP8VcsyGYoRrzn
VXRkbSaOBkWrf90mjfH6AyhgEcE6oEtWmNMbP/gvhRg0qPJx6LeswyNTeI+hsH+zjplPJ6/pADVC
ddCG5jayFRvlg+EwnAGcL4tpm/9hWyncB1f5Ej6DsrYqivC2w8gCm1s9/6Lcjkog1Ju4Q0P+X6Ze
lvs1FGIR4HbsqxTENYsLWS/XPzHVZ1VggJBOTG+oL+sSqbn7V8VFv39daIXDKOtNzJRnWcIYW3gd
m6TjqroSuLR1Sk2wbuGxVij91BsyLHgrA7GVZOnEH3Sh4oT9LlzRkCvfYh0ZX8CFoI+L77iZpDPu
a/O2mbYRS8GCSIifbZhwTAYkdyTju8j3f+4TYSa7ZHS9SNBF3jWtk2V0arpOu5kLILpGNmVurjT2
rYrfEtax3qmHomkCNFdqYLtlFhFaW8l4tpNONqV5bR1PXJ7j+mebLAO1Z7RN0wi1dFwwR0orGLQC
HbiU7VdmEHQQCnlhr77yUPKxIKB8RMo9ioUL1+M3+hP16OoOWNEYkp+xbLzyQwEoyjwLteJ8J09z
oRd34fZLRRanPZ/RhWpz2UZ81USSek6WG0RPV6UTdQx7Bcw01GdHEXLA81Xtt/2kDLTJDbZoUYxo
Ft/nghhLbF9ll3MMsY+g3ppAtHCEa+KcbvX1RKNrNu3mLnqg26z301YHJTGhfDinsFq77P0djpvl
hYJJ6eIQUZieHhohyfwjN12I/ffpQuVHtoyaumtjNI56QqxneS2+v8jMC1Egrn5cgdfQcyMNxHVL
+rRW6onA//V8/OcvdAH54upq46qeP8kmUP57rr+HYlt2OyIpbgcuUYTDFSvD3i0kfMIMdaK8a/NT
8Tiurk+zPyOV8Iiidxgim6CYzeGPmd7Xs3i6WMSrlHCKwN7/y9KW3mwBlEQrBaUVpFxA8qMX4lQv
pZr3gPqjWfoosnPGpQm0EXnvJmcCaSQQis/A6LDX8KJhlt2bWdMgLB6JsVlvE+jAGrbb0x8lX2r9
dwX2RpI4bi6dCbH9ed0H5/lmVj4SFh/5TN3aNMcPSG5kzjlL6k6YE8dcS4dKTcBDSfHxO5K3el3w
mw9hyDzCyzwHnHzCkbT8AIHA6R2NZ4/wBZcRBiBXo0o6QM5ojVMIIOjVO6LlgoEt3DhJ84G0dag4
b6Mo83UbCDHxSfx/o1P6ReJ11CD78m/u0pmXxMz5AHKCguX92qkJbgoTNgYncHaVU/MKJAO+/vUZ
xcsWK9VIoTcW3bb39Cp1ZOQwFTtzLVSKJ4QcPIgRJ1gh1x4qt5bAAlyHsyM7MoTWqatZ/ARfpSxo
81d/kLV95EcwwdIFJ8owMvluDnSAhDaUMmqkRbq6ck1rMhg/SuUTUlumhsAUBohvKtB+SHlX96fA
sAbCRqM5wi6FQt0C1ZmH+S6wVqIY1Me3iXnWqzPNWbLTKfizKAEg6hSXcdYF1/WyACX4bE+uqOjQ
INSAYlejb2JTIVTnUSOMhuYmjxF5LulKxnGXf4i+a4ow8GkWFDaoDvBXalGVKpQhWqgAwWN52OqV
AdmCGFg5YGfFPKq0acueTa4i+UitCOuFAAqWz9v/1ZJ/piE7vjQPdzwE4tk05ayopTsz/MuvWOrP
jBkqcqfCm0lSO4/z0MijoIvAUmAwcQ0kYtP3ShS7G6NKR5RFREYCDZSs3yrI5l6XuqDrdpWQqbqO
vbHNJ0QAIIh+BIt0f9GMKqU+WrsvQuLnIlYPKDZ8SX5WDEb8AB5sqmcaBIljoDCbmcfm7fZPd65u
gGvAFQi/Yu6SVYFFnvauW6wnGl1Eww9usotYM6WsEcpNiHHhjM+JrKLiNqp+OWNw7G1ZRs0YY/Ru
eKoO22isvQsn0fAjeezf81R4VnBJJdMJhFdvFytIdVcDJ7tEaMe+dWr6jYhHClcVd65hy1f9lihc
0hywstPFrZO4zOVu89u6U/3Bvwaf2Z3mD8K+Bs7TPAA8zT31ruSbgsZcu1NY4lh2kHGUTwLgXnuV
so6V9N8VlF/xKpyBELV04yIsbD3jRZ9vAs7+Ljtd8ejDrCqesJimHQeLAOlqYSnmlhZIe5o9MbYR
qSn0CQMNBn5DLLn+js2b9W9ED/iu0dGfqK5a5vDCC2b0QAzuLNfSb+U/jWX2k07/jK4pOLHs4rIF
fmwdpIjAy+JDz4OdNKOypfp2bxPcwVNOcY7sAHSRUV28e3Cyp4VT8Pj9c3GQ1wIAsEKfFZW23joy
xUolvxLLxGFg4uxJDfBIjaVbF9RivExmZ8JECUUQ4+dutI9EBY5mAaHTGiP6w7csA5kCAazPIffp
74BCOTJobGdIQ7Zrn3qB8QhC/d2t8MKhVRDwUI3eN3VCZqfuA18jgbkK5bD89ab5OzywW76Mr+SV
w/CrptWwBihW9CTiwwdx9CiDaoW+xAExjDFVO7Z9ogtIuZofGBgpb9dBwqT44RtYYPpfjebHZx0k
EZY23A2w4V3FRJYOEDZGZFzoC4Bgw2j0A/dswKSyjPvKXt4IXmPNWQ2EHDDmwG7pcMIX/UNy7Sal
jxZUPpCRyO2LczmTQhDHsDdxJOAP5RtKooUa0tVmP0sFAYr1f8EN+i6MHh/isJGCYezkWEY0ln+r
LkQBgtzqtEgQZaZqjrmw+otFcCId/BZ3Ole4Q4d9WvPMITtTEE8Rqb5spLwo0QLIfsXYMVolJJFn
JGVTd32SykuUUf44ELpB+9jbuwDD6YTUz6GaTJLBkoPDFsmULw29AWYMgZlbUm0/CYVNBtUhiRpZ
AaTdqjGby2hpph8YCLRnIIKSsRZOgQqGIihW49LOtu2ZNeHYitPRgwdY+fNA17QnKaSQEGRsCjYc
xvrgTl07ccrzFKxiCTqIaf/kRysdXtvH5gQolzXu6nahKmdcvgtN8jlj+/wczUEZPn13YPJH5c55
X6dbAdbeWldW1gVUcUOtD5xwtWI/fb4pCWwVHwwLatUHMJs1xEB3cnGCBhPl7k6avpzpLgT6WNhR
bRuhRXRxXaRwOgD4wUOEc2ZAdtM6d+civcAcOY3aTG1mwYmiVeDfP+byB3rI5oyiesdwXliCL+Zx
4yaLpJ/O3RWTryv6ws15rZ0/b5uQIVTUZaGnRkcNjYW+t0V0oVd8sDgf5zR3LmNZQZASdpjqF1Bo
d+jpUEGul7T+lMc1vossTBTuoSxmilzWWidwOSLY6ziTcgjRyHzVlG6L+SyWhmLAgkYmetYNBDyR
ARS+U2qkko4RsQllcvCGzbaQMcCYvCB9U/O/8f0q8thKvrbuqnwBMpgPrsUHXdAckhLOhZwHcd4r
ECiXnN9qBTtE3MBuH9Vd/PeHHY6Y4xsD5HqTAbx4lmdSYmAesqQk51sc+CnGbBxNt+205QzyyQb7
SxO3HXCDLujs8qdnctkSQEFksMMELfxTlLeRd/He11UDCh8TbmTe6YrYGcsXM+pofXJxdejFNyTw
AO77dYqwSgZ7P0BuAE6CRyqD4fZsnlpWFTJYFQO8QtzPB29P4l+LvJbZjK2U/0amevkwF5pYXw/K
JMrp6VMfFoihDAz0Za5QCs1Mjm7+Y5pkfnNf6jUfelWPIu2lDgESg5D/BeP7MGnGJm9IcjEao+8j
d1C0OfcI97SAngP2g13AWp1MdBpBymiKKPaSE5HmZjpBkya7bKj1jfh410loO/OV/F2ZDRoZBVmb
ZDmFf4+kRT5pgo+s5RG/Div/AMLCQakrfesBqrGk+R/7V2nspeY2sHVKjRNzI37jCZi8PVWHpBFh
X771bINMf4NvasZDCGWlHGHeZXLIa86B5D7ZTIQfx+l0/zxtHnDA517NlXvfIoz3uSuDAcALEbXq
b1XwM6JPXc1cDkhOhEPU+vQwkiOZwKdDoZrMBBoY788SW5nGz4hFCxzICCfPqI3+sRSab4nldYkK
MoDOjVXrxnICqmrgAbMbqec3Zsi91kgVkp8u5bo1gyY7+DPZPYNV0K6CGHaUuB5B8VJDpoEN/PFd
nA2IvmXubTj/z2vCuXmNj7mYTbBgQzqqN8RmuOiEL0XGwXcKQGd+V23be8dQIIywRb1huOnQrk3W
Rgdbo+5ki3VKM4Tgm0fEdxDoSnv5+43Xk2MD/NGyZFuQE1C9nkgOGubbQa+wd4EwG4fCmqS3LLDv
PSfQGK1JHHbHriFyLEzaNpzyATR8AevpGQKy76AW+s2ztcvnig1ruzZAiRWqpDDJHM1OaAlXotdk
Y5BhEnuciF2EEWk+dkLTbK7UpOKOfvtzs9d/wDK6MOG/i3IvItS27oleglqCER8xNlUmuNSucBvi
p2qWjvhhz1/ZyJE+JO0goNcDZQj4ru0FbOyfydUhMXvFlx0j7VQT4bi7yzH4Btzd7JwlPnS7h1uV
7fhCQOK23VgmaoUple+RDVUlAj5CjpXmiI/L4b45/UjmsnzNpbjZZl/KKMS+DvpppmmVxAMhM1Zm
oj18AEZDsXVnGSASNLlv7vjDiMuGc8dXr9sb59T/n/lAV/hv0yQL/8nSADgfC/6cl4d0l17LZdYe
gNYFmM7rymFmfQNhxxzsgKfApKZ5r6O5Ov06jRXaFLbKUr7764/3GphBLKCWGxQYq2gKC9EXsFwa
qkIafX8KtEV2OYyxsj2RsQpDcdqG5C5tPJ5e4c1F6R56Vs36+ehcLfHij5+5eNJIIyUbj1S6dYrj
LdFylBxXPEr8R8WNj9oWoGxT+zz7KnkqQU4elXq5NUndL7As+jxYUEpNwIbymbn3cft9BNLhTh+W
qBNaMbj1cAQugHDzLsXUlsur9pgchdsdrCv0IPnu67ETO6e7mqMz5qllK5NnCJYmkaZJUX02Ir1D
5CuidItCi4K1mRifqFCQy/9uYt/+8S00GkGyE6LX24b/LYuD0iiaNCOyA269qg9Eh/CcoWTZuUSf
zB5mJUMgQ8/hM+Ub7dy8uIlyF8IiHKccWC4kUtsKT77OST27tS3TJ+km73GsPAPc2Zac0CP6bLKd
CCvxk5q71x8nm/NP2QnCOnyjgG8setG7ty/ruIOTApyfDi0seUFZDNMdzsZOtbtfz7vGvxXCyyIB
K/8znmCk6M4Fxpua3+iP0t4+oDO21rb0eUBug8tg0lcp3+wXUjO/wFOm+9VXT75zLF7HVPgvHa/X
uXdDGVYzrCpN9XZ7hwLAYuvlDznP9wTdR/Kabiuqr1ScbiZoz0GvD3GyPFiTIyXqLnrMC22preAj
1ddQo8lQa7qz11kcHM2vT+NcmteqqX9PbU8H/tAg4FMzgylVMyFryG+7JX6OqA9gHoNqFz450F2/
Aj6THSDepQwIoB+S4kqQRfLufZkkan79a7GVeSc0z5+NyjwonfFuI5bcGEpfJZab0vaguxVp8XFN
6wz+Dy2QIC6M9O/UzTACdeXB8bznl+zD/+T2HwmiC+QlPrxyprMYRHOe2hpBggWHmUHyvMRk36Ht
hvNyHDN8KrKs7UAuObEHQngMVwBpXF2qhVQvC3a+b7VCLgjF5ojbFtwqHY311XqI9P5C+9w8UxPt
pUdGrXbVAmvgxpBt1wpXrzhzxiJHWZtbueUeliXpm8VWhO988nIS94rckFR6guLH7gtR/p6JWJYY
QAaoivDbWDD2yfzw8hXRrW97xcCmZ5uVrS3vdbGYgcAl2CERle2foyNnZ7X4hI00fhNek+jeJsa0
M3SR8BFns3eN/ZzULY8sZQcOK1Mh79PTj0EufKcCrupIkH+BQB2qko60cO7C8PfgpAWA1u4wDuLA
oj36lzhLO2QUxNEMUxnidXQBpGpjv+p07IXwvGy3kRQhumvo7bWFGqCeu3v3vPs8qvE3F9usUg2+
M7IqbmEFquTQwS621mqlrJYi8qJJ6V93sgtDr7p0CvUHyvVTUe8N0lyjKOHK41HNnKmcbvZB0DJa
KWH4oAazmIYAM+sr/P4rVBjGpngzvIk+8hx5+TB/zct3gDxainhnACIpyreheOmIamppO/CDTrte
eib/GPIfRWjyXUGPQqP6B4uWhOya65FDzlVLp1gZSaqcqvgqT1qGum2bV6tLGUzXBWd/IaTohJs2
gclrf1Zr9PUvZktnsKeoGtgvMk4LX54rGPNe8MY6UdeNX/pPCb2Z1ALPKiCZEBuO0G5JvTsZ3DJq
NKwUqZ2p9mDMJRXPt30H7hWupLNoUfvFCuJuA8TrpKAI6o+AXvfzi7IGXUIanIAb+NvEb3jxqZqM
Cm4naHhPWGJwvqzwYYFx+0ffLev8GZRS4N4DR2sHaXUlWy8QMdeCfZex5JnamvizlGwNstpXRHyE
Mg1cz66Uz9VAmSK0Qf5g6CkIhhjZ4ZqE7evvuZqP0V7nclPMAVSpagwTskETkPxLNvaEn/+PJiK8
GkpaNbuo3u0lyCL70rhDqHKzAzB2+PYbr+qE2x1Ij9D2K579iTZk4rnBabHmWLeFn77iESx4jbJT
51d8ePivLLUqZAH/3kgw8cgmtq7nuvWuPMSm84D8xF0VSAKQNYsP6ZgJOgkHrtwXuHf3hkWXm7Pd
fnV4aGDHACZ/EoyBzEOUQ/ftqtlBKe/jV0Uc6J9vIE6/LCoxnPha5clkxHp+fFqoJj6yrNmxLT1E
lf4x25yCQaMY5JINrnPaTEK57+RA3RBkk8svETPRGNqsgCH1zg4Gi+JYqA+f728d9Lxc7FEKbwJM
V/kFcchZZGg1ctRVO4Ua+RegbdNvjvsx5+imQ62oxeHqmENNBcsJF12E521Q3/quSByLa2yWGL9m
E/cBEa2EbvQwoVPG1sChs5utZapMqVaAqIB2var9OKZGHUCnOJOfBGu+OjgEVIxUqASGe1ZYPpt+
AjKEI3kmrqVTBCq1QrWtzV/N//o0BigJnVdOQzzq4HfuEVwLvn+Hp8zBN/eUcK+Kzy/7F5qn/PTi
0iUOHd3CLn6ZlHOKSB9BJdnN6z5eqM8VV+a0TjgHMrQDkDINH0C/TnbvBBKo9bjuiZgirzJXQSyJ
3L9aSxBG8WR2fkPtiwdO+4UqwvVzl1sYSBgeutXK7/mGLybuvJb9GdLURMlELdOaVOsRQtusw5qE
l3GaA6n5LTOwNiJc+2i9tOcvJ6e+Jxd7wxEwye4rTCBZxM/Lnxg5R449FTkYXVN1yB/xzIawIpit
gMB/6TZ2Me9L5/fVu4Sd/4w1BIxE5fqMDkXYOFNcCgoqRo5WtqZko0TglIpNeo6jWFZTupDfQl8z
eKTJPICoogU7htMGEckO+a6oMjG0y9FF6P1VEB7Hl7HxU35qPWoUkRZPKKLXV81ubre9KMGxecXv
eSS8/3LAt3Ye55rHLGeeZ++itqciSURyfUml1XPexd8AP1CfUKg//7X31zWASmKMD8FfX1CHcUZD
TuMbMAeZJ6XthBG7f1nCCO/lB8MvRQbI78L9UiFCMremcXmHGNK+b0sGYObvaeTb+1xM69PILD5Y
8448fziMdgBLA0PLk0a4u7msmhJEb33zgvVbMe7g7LEEOmFjA4DDZb/LPf2ggGt1m5VBBTd1tABA
M7UxmqyqgqVQ2LLsOcGx1VNsu09LJQKVg0Ct+nvXWMudglWl0I+QDX7POtuPr8BQp4qmAlhMr2np
tQG+smIaYzD6IznMPmX2SD4RnK1cwDWQUBDHOiuqAWPlBvctNWxOBt5U5JDZvdSwvPSwemOroj8K
8BLitAcAGXaU6IDLGJnzlEtH86lJZsnMg+zBf11Go8howU7HwvOu4MVD3LK7xi9IchWUjSY2XJHP
MKJlUJ7wMRE5DfkzZSB2xj9a1qD6hS4AJXLfYQctIi0BFms3YJIcCfxaI7Pn25A41J7XzwqI+06s
4WzAGmjVCrOfTxzbSQepoqxVF++2EDdMwHWoSeaVMmijFg8Ueii4RaPGuGHvHxSMwx3YCL/zz+Uc
aLY1m5hchq3Uig/CVhz2eRm2so2YnBxekZvRKlXgti7svJfpnMUyF+uY3cSRnmzUZgYmSBQ2anmz
Hj34pJ59y0Y5TENMKp61yQ3g9j4PIgS6yXQv7TftMV7oCG9CMprfx5zWB4zxsiHnUoKr5h/Lc93e
ywyNJJk/XibVnl2lTi6k9Rq/oUN5/1zudXf/LoM+mAfOOvJm+4A3IRd1FTuWOXhBpHPAhnAOgC8d
DEwv88ZSuA8OujKemmxWsBsIDqAWilYXBccRexxi9mT5xmL7LuSGn37pNyktbkG+0mS2sSDjeqJ8
n+56TCkJ/kiEPakotW0rEi9o/FLTmVTRt1xOaI5GD+M/JbTId5Vo6K/Iqn2gA7s2XX99frm51upB
bshTN/fz3f36lWsjMGA5wUDBd2kRifa9lM9D97GTcNk4oJS9GEIKUlcaLpOYM93nTC2875yBkd3u
YbfmyzlZfj1C1jDyYnlqIq9a07Y54FSQIEJRBMipIAFjJnD0Ivb/X2xU8w9EAWyPWDkFB7InidIb
7upXjgnly8rsL5beQFvIkZI4r/OJqg+drfz1JQ9ERrp7UbWB8KiE9nEsMG2rqKwra4+2H2isGRCC
LLsRq32UQloeCBGDxBo0eUkL08V4bqcYVp5xAOJbHuQim41HaRCphYQXzhHAKGngvvbrqSAdJtwP
CRQdZshD6dUZPbVpPTwr0rcLGHkILWnIgvqMKBcwv00Qy3fXNK3n5TEWuQhja/LZr07cM4uWp0O+
Ftz75pc2nGpbnysdcfELvul0TRrIhIxkG/LH3iVt1Yvor4hvgasqTw+gTp6h6Ymz38BIWOTGUarw
JeBl/+6OHDfod68e0yNPI7Sn2YWz9cZGJt1VWeV+yZFfFn1MRI5qfk2AThraqP9LKeJX2G0XanBk
ZxRqOZ5iNGVGgJ8DJ24EE+rhnqOuJEHWG6dq0YX5SaSgNol1Jt9uV8uXB9sW5wxEbcJuWASYJbx6
mg/ReJiHtz6FAo1+A8isDJAqba6nup6ShEHk6R5Y1ntkmmBhHLsM3SMFvqN8Hznv2fX1BgCJlcDR
Sx1RPHkTPBRaCjqYhsIaxyqKgDMmfGkahJeGsUa5Y8G0ogMNvBG9Sw/TAJGXb7HNZXIvEPYsNYQl
190NvK8BpVl+himaSz7EQktb1uJUXkIIjGM4zIMEEZz3i5PeLKmbl+tK0U8/MffNIWL6/VEya6vP
SzF1Otq3tOcals2IzL1Idt/uBZGivJ35uXB1q8WwfSFLP1xOvjBxgaT71MTD1+MesvSPTBkuo8Ky
Fa85GR5Kj10Aihdznw36mSyeqRjvkXxTZDL0yB57pc8GIVbosPFc2n16uxq80lyK1e6r1xv8kc2u
Z4n3QVEDFeeNZjSYqMLIw+6vE/hQiTmsTOtHA9vvGDA+1HTOlMstuOa488Z2Lw++4yfXG4kAZX02
F9YpJwg5DKz1weV5gfP05NPCRwbM1cD8+SbQQP+LfEmrzl8CaCOSs8HyvyDqZuNE+tdC77gKnevy
4+yTPT5i6rpciE/UwSlI6YroODZN1mLqSx2UkwBhNY6RvWkJzaWGNclNb5mdW9WrIOOysCLky0FY
APgFuHysB2Lo5XiDCd2CXvQVnxAqBu1L3okF2TJUO77h37CZ8Guez/2TVYuPdo8td5Qz7SyzUoof
aJBsZTWgGAxDV5D1uRkIUCl7FE35wMa4+RTdHV8EceCgTc+DXpLBo/s9Ylfx/GxfFeC0MFdaoNpT
+/JoNu1f2WVbnfdAdOPTagGp6oJHlVVqcwIPxGDDrZ80R469njiq+Q7O4nEfaAN/klo9z5wHB71w
DJLNs4AB3l574hwCjK7Mzey8wDW7yAkvoLmwpTrR8AOYSvrWwzTsv2f4ztGCDbRnrZ9skwOA39XY
jcu+Wyjq/RugSn6iDl5UNjGCyvSFUaWM1/EtaepvogsmlkpZz2kdl3RfebRo4Ybk/1BLixp0mSRu
VRJKaiC9aIEyRsxgPx9iTfeDFvqaUd5L5dh2OKcCzg8hiCziUM+AdYRyOUSORQS9XYW65U665coZ
9wOPQNs3xuXsjSxqLokbZLhfJtybc305vWLafa06Vkamu/so9FBnwsLGBLYeYer73fC3AFXF43c6
wLAxbg2KofTb5dLWIZ/SvzUwW03GYH0LoCVR5GxlIxjuMOyjnAX543BuQWOGP3a6CzQTA5rb9A+U
p/CFBnHN8e5FyV4cN75wFO/x3qBVxTFeGbDoKe20aXD9D12/pRdEZAaA4Hp790dtnXY8NrCv39pO
enTc/myp0t8TKH5nz0Ibz/ATDxoWSHbBWp0CPozAsnyF5iunMHm8tnIeSYE/RmuKSlKE2fXoGoLy
3csv+lFo6aPb2+dF6DKl8Y88QCgWb9xFisZWxCBW83JNj19GcFLfSu4alrbFFWG4iz+P70qOZ+Wj
JbDzwCMu8G+QLXAonz6Fsn3CkpneRovqlRysJWgqP3nprtJvrhF8j45jWEJZGDLLBT1PljDz1Nza
T6To+RBBajRuBolXG6YKEtD+k/3i9nCPzFEAt2E6avQgrQHyZwIC6CivVRor4vqkXUSyhPfL5UJr
8zUl6k/i7tu62ChCigDVLbquQVupfEbtxNcvyfHeNxL5u3215MZgKcFbKAjQ9uqoIPr0bYl9hVa5
e1wcguPWLwWP9fhFsKHSOy+tCY5qpX1U1oCrJZDdv3c4ShebHUTxH1e8yx6Kl8iZ9EwGiVqW/f1B
HMC92kqJAy2oXaOBj3ubHUs8FBzZNg2jAK7o39bJrBSQ/jS8b1B7dI5H2Q+2i/ayOHt3V1Jhkx9H
CNtNx8ZK/VD3d6fPgL9Xl0JblqWNC6vP6wUCr5cK+/FEQo8lq1/VpYdGt0p57OEInTHNBzOq1I51
gm3rFMIlq4l7Xo/bhPfKkNN5h8gDzFd0bi7o2doL1v/dRfiSLrsqSwjbuaDHgJce25NOS+fe168t
myW3cA1V3BmwuBANRKuZ2kLAO3OFTeBYhORtzX1CMw0o5YZuVPECKj+YPGPWeVccyQ7hlGu/za2w
oXfolwEgCsfFCkZ+br+NaEt/ii7tb3D498qxucRZPBbkbQgDzGyoUY84XI7O3xsEyJ6Ts6r1HcK3
Sh8eIyMCnXdIFxliKGstuv4czSDYVc5GN5ztKipEgTv+s/xZXz9U2fCMgLExisuY+QCR5C48ZQ/I
iQ7s4VyftxtivRKvv4/RMmU6m3bxI1BuBOW4Xp60QzEEYIvIsElv5Mh1bT6EGbBsiJVJSU9SZX70
A8drTeSbSmZkcVqYnWtzLfoT2ErLFMUmxjrUx1qhFC3gQ6j0DUta1V0mSt4e1NZDZG7bYVUTGSxT
1K6gg/e9jnP6eG6CB3swwnRJ3uXnGomwKGZ5p5D4DfhMwTJHfI4DTSjMOUJ+YNwrSocPM7ofv0gg
YGyGvEvgK2Awt4YHHgSaHaJcy7ucsx9aG3J8yx50741k3+ixi93PmXlhTknJIZc9QROVN26BQR0D
hHNxTPJZX0o4jPEH3eugK5S52CjkuvPa8Z5qqSUkCvTpP79A1WnNyhpTRDEFC3z37OtTDN3OKj5P
C6I/SLpkvlI+Xr0iiP1tlaooErYRNrCnuqBqsq3wmHnl2yuMaKtDUAVofaEZ2M/a6cNtvEMAUOzY
ifTiHi4xfxzAh1zTrIM/+1QNQ5TSbaKjigEtqRu5kJfeRYt9CUQVE9w7OIkQiD/oJ857vYMlWM+0
WGiRYovUzHD+e42T9fK2Tee6EpoCt4mT6FSQKrcS3M1d3BrNmYsNj7kuFP2uvN++/7pgJmQPWUk4
AOE6Ru6b7abq09pqg+AfdLjaPlSlx9rY4TcLIMk3t6UGqIAlLa72XLTsD2ApNVJ//Qop16OKUJnI
43ZZb2CANqR7mWmZtZUqV3qRwGxesKLR4Kp+s0vbHzOmbhgf3mres5gpv4m/WgGTs1cgt27JIs1j
PNfBEYtdTLZuZiNVBUdBx8u9UQmEyoAAhKiB4a8VdsbgUN4/BTrChTSSqzwKSIs4SNdGivr5YEQH
5SC5sEkiRRh0Kf+XiFi25yyZ147BRd9x46YH8GAlEUb48ezkvAN2hWAGr2FmvV+FUSQzy6p5l9Qo
J98PKVP+3nst1HbzR1YoDNaBemBri4RtpTruzfaXE7flqJFhfeKnK2fcSsFLY8IcXszIZmRzin7B
ugH5RQUplTCyQ1NL5jZ2NnFm8WNAe8XMgTD/6m26rwvCfSckVqHyBXeriGzBiFBgO1t+K3bPo3Bf
XX3Myd4JgKZQtYTi0vJR8YQsWVjHQdZlX2iDNe5tIGjZW95MpNMkX/w56a3+NujZ6C2L+j//VUU6
a8IxMFZU5vx9EQ6eQuPQ/YdLbb1ONolE1G/6w/i77k+oWRUXy5J31pPWphL/zJWK8jyaVhu1g2sE
W3o/f0hRwStM5HmRqgvgfzSmotn7x8ZIRkqOi+UNArfx6idfTNzMwTrtRhUwe6KSfvTZ/SYEWOi/
yueXUBa/qnwuYC50w7K6279xZMFEyvWqtqCt6qTQtz21gjzhr6cPLXCUqpZWEgw6BAVJgIn3Wgln
QrWMD4QOsiMpoCLLU6qFhbq1S2CwA2IX7DYuDKCEKNLZ9HqOtS7Z7Ty/d/bRrQBjdYBfDl0NKBB0
Rf2MiWp/KduufPhhgWjZncBEVaG/vtRox9UUaws9hEGeEMpAWt09HNhqGuxBE4WXbjcVWdiLqY+g
/dtTmuM3KBCJNTQHr7krjjC1gePu8DLdYf2IxPtlbMqYDMqIylp9m3i42X56X/fgjIK2CVQaGTci
B7Dftnt9FiNAVly+lSi2HtXXvSqKrqLqHaKnl2CiMX4qprDnr33Ap4DvLwBAlXodb3WNi0zuvFwb
sQK0V0NlxyJwZycldeMj1y/hmPrbMcJEmxHqYlXh6rMaFz9mwSItuwZAab/r3IS0IBsW+4Dnt9Fi
W9MqemeN8Km2z5Jr6jyQheR0O+6D7ATE3cP/dJUw6gemZFex1LfMpEVjrWcII39MJXoXd5GvX+GO
j/NiOHYdIpuXWhW0Xa94wmj84j+pXw0QDcjSHExLJfqZ3/dElQ5PaxR13sPqMnHvVfkkqSwPRZna
OEPOu2JLDwlWOvNHxb92+P5pWl+dVDWJkyaD6Ap4htyUY0bGbm9hprhzc8jWpt8uCtel2SxKvG2y
GmKaUqe2v79Vpq3ovaHv4rXIcwRHUnaALMORUkkLRl0rpYYfwqQG7LPw3dkEHzc1qoOfb3/YsMGV
+zMs0o/vJeffJAjrdYCW8BZ5wiILa6m5/7If+O8sqMnQOwGR9e9nC7tAnkB0QKn/XbzPORuCuVUm
Fkw/DvNOysUI2SBD7XderFL37J8RkPL9yv8kgh68PdSxFMne4OwQpI3RMJLbZhCLC4Rrw8XtShXb
xAGD1Rse/foyGqJ8b7Qf0SG2LmbN/XV10jUBPXL5Jflh2l8DuGC89Rb12ICRoTbd+KuoKseHCF+V
B/6cOhQv2jbgV6YMeb0PMuAxLp1aCRlvVyyfWuvUFYAnCRrbCA7dCPx2JUl6PY+XU9d8OaCYqLNk
yA2KDbyzU/vn4GMup37HeK9TdYWfQkPfhPnkrsbYwg31T1k36rVsBvAPMZ5lyaNm4sOjwh94jyZ4
XLbYfjGiTtC7vOOms0/O9gUmhXPQ2clWVfjW7zTDWIc8kbRtEEBKcJCCINqtkIOIgQisppNe23za
4KKOq8RuJBieiuv/oSQch3KNGyoO8r48ltZiqPXv6P96WFBaQOqpPcoiFc5Dy4MwcXf0Cw5uderp
9sBtRjCL1AFZnCiv/ttyODlJ/nC0KywAfo4Qma8JTHXmsSu6+HexZ3vl7OyyMvRRKHpFg3RIiscd
0ETq9+CM05nxs2Y9P1SJ5dJ71nyk4lNR7o1o2zkVtKC/IIPyex/aIsmSNX9j9Dk5/RRbFMax5Gup
HsxfAi3BNuklB86LYSc5BYA/Trn8G5ta8sFWdVLIwkFdc3t9is6gCwL//yyFp+WLvgfrDkU3TQ1+
B1KUkCyTzTNrsbrKcvFizu7Sh07aI61x6Np4/xxiPhHcIDvZoxlh9p0qX2JMjOMK3eyN65NzBjzH
TvhMW495nKZXza2yNLHQiwck8x416QHW4tbR7eL+O4p128gzi/s5qIN65juUxsDmKK65vD5bqhuL
jSr03jhn5DogTShqoPV33zUWAso03DM8AyGU4x+LmDcF6tLft/7WElhvdKlBWoTmCubHrxbazCyn
2yhwHUaGoeq8dCCpYnEj8VMOcIOwWg9tyRJOHgees2R6n3vGgiM6U7g1dZS/lkdUni4C8swZ8UFa
pf03nx8+qCdif/mCePs9ntXjMV8SjFqjZh4jcLyBy3Lil8YYYY+aKu6lwh+wXozidHzXdmNGoX9g
q9gnCQkYER9ZFp8adann+i4083a0NtIyEOnzD/ts82B2J5uGEBYuZPD/PLbjLyQcJOAjJosD61NT
uQ8yWwqr9hhXxV4osMwVAFvObuHS8Mf6ccj3L3uQx5pBfJUXPQ1S9oq7z87ZROuxDOk1kh7TjgZ3
y+/4GVRo6gLjMKqopRGC5HdApfUSxlOiy+1egjPsomGG1rvGNS+utXFC59cdMOd+fG5yx2Dd9jww
nA3GfWEWx5o1Sb9c/aWX4zht6yJd6XZfuLkzxLFO1QHTjS4Cdxyj2jzq1kyxtL9uR/ch2dM7Z/Cv
TEm+wKfsWKAWWlXxQr6N3gGsPBYn9EicGHe5bQNnyvmRj85l0DdWVhRcIG44e0KJgFTgvILdaF21
G5PKuOhLhmYjEt+gjTZ03j1odqa3lAlCK00YfR3qZsHhAPWrF/slpkIqRv48YNNBtD7HkNHWM5X2
fipYG35wNp/pC4j3nHaMLw5ShR7vhXQ11CoC7aXfN241iK/5cPKNbbsSyZrOq+HDfDThRYNqonmK
wj7dvMRoogNavl06CgkPJ9239/YW0AklE/gS+z7vi6TBl/OksYrHaO2BBjgK/HVn6tpKhPflk7lB
T4DI/0R/mCTSiPw6gj5wHPtMQD8Ul31ru6Mciix9okL/x6xlWXBP+NPfcdbEMFjOvpizVzwlDaa7
HYCeRe9bKzsUgx46i1kK9gto2agWh1ewSUU8aXZRfpj1BZdnrd2dzc1j6i5zBjvj+ClwXF5koJVR
Y0h8eQuBtcvHXS0D5t5GKKaPtx6U87guAycsi6FIM/UBkINfeyAiF2TNw4kmJEKeDyyyIdgu8jeL
ksU5GYz+i3JitoM5YMKp3AjBYMzSrWEahksQLd0NFDAf/J2nPW1XHjD4V4ncik9R/tcCg3ELERod
1XXxHd6rG1iAgcCl9aQyuo6vlQ4b0ZE7NO/qQPApic9bXrvsvhiuCaQ5fZm9x0WY+A1ionbSJH98
6Pb+DXjkUFDSC5Tp02m3mb5HhrZSEMRrPChWy9BF/UR11nyQfg2jFiHusSUQ/z350o9UjVCnYbUB
Rw2aJXw78adOjRq7TJ8tPJqwq+e60xKdkR4ql8vXU1GlTqnt/tHvEeWc4LprDKZwEnVl/Z3jM2Kf
+FePCLsuP1a3ruJf48Gy8DkqeK0NI/mXeV6thGszBRJGr1s8ZblxsYeEEM/o62phqI4J/zsbXgG4
SN54bdTvqlUsyOPn4ljDeBYzsJIL6FErm+cMBax7Wvk8hb87AmCp6KheBX2vYcN8QvRHzL94lWtE
bnEsZlhVS291SQ8tR2QxA98ekzhkKt0p8vnRH9FVGbdfGVVG3W1gEaUwsacPBv8Gdq2qrHH9GoH4
D6EsAX6Ib4OgXoOsLbKJMviHYLtwpRloilDaalAszswQ2z8VzKfWkLaffr8gxO8bicCGxs/nMWFX
9aYFsWlBHv/qyqZtgCIUPZHfqAHB6Qtmf9QYvS9m3XfJQjSCM3q40CBttacOZV7lM0wZTaYGH8Iz
mE75u92ikaS+LXOXOojZTIMRaIv3AWTNM9sj/I6p1XpEw4R7CykM1QpwsC0mSfrl10xQyu6ZM2aI
juAanejiWja7aiIeWSpmrFa8Wz2p06G68m2fYqXI6RGYx+3eTrmCIZxhtHsyRhJDJ02FhDHfMNtd
hOA1h4PPFexmpy15PlhIHwPpBX0t8G+D8h8AiMi1g/U6Gno1SC0ZJmyyga3k4kcJqDM43DfpKP83
SQb6QIHiilhbcW5eQ2owAyPnPvqM2NbeSlDuX6ehS9eqIVnSjF+yxFAVG0d2NeECXWWITw/b6ggo
OyqahtDuroZpanNxafo/XSJ4l3NYnXofBObaTMREAy57NgjX28w29YQuTvfrIClTzCQDa0UX/u9f
Nj8ZLcHthZ9r4g/CA8LiCnzBkTQt36vTL6UuN/rY13RiKqC4BreE8R8Qt+GlCzLOh/g4L3TkLgS/
086ttMKGO84dvnkuwihL6x2hbYIkaMC3elbVI3+Oag7EqYd6dhFpC3+jmo878W5d8vGt2Xsj8NU1
C5PpDkje+0lj31ucCOhM0BaBxh5wEfmFGf1iiJCng8wHt+8POmSDAD7mC2GLm266HppvayHGweNm
Rq28uzAc3Z4kEJ/tPt9bvm8GeYdORzUAvfNlVSG//eLPjL3WBafqt7LBw6rCu3hcn8ziiub8SSBT
DRwISmqUlf+z0MF8ATT5C4F0Ev1tbo6tMJ/d2XYmRVJFSN4X4WcBixoR2Vdc4748M8z/Q2xjH2Zn
C3mcxxrPbR7RH6IJJDAmG0AtNOXFT9GYvldViXBTAMrahTimspmayXt262He2dgbXWxmmtnLV/WG
n7PmGrbXnhUiRcXDY4rmHf1+vQmJc/m8azFvyGVdMMYmoATJmSA7KuAgrbuFkO/2SBcerU2XL6OE
sBpw+1FuInBjRxvxYo53qA0UKTYdlKuaW/SqhgVoz+u5h+VSo/+I0BX8FfG0fZ8Gwh/7XWluOC9r
x8qagbL7Rm7ezCw2Ks9lyGweTyvu7pwGO6djxiYPMUvFgian6H54HQgJvMPoXROzakZBnjEyBLWM
z0YiOXmcLM28eWPdbqUvJIwtK83cHM5q0znefdCSlfxveWwLDMAIyN7VBKp8ImxgA/+EeA8jh+fn
6DTD98N55bsy2RSW+F+5uF3D3/z3uZ4FfQVFs+rOSZign8f7iSzRytbs2GD9q8M28Zag1va9hcGR
K6DmSyG0JY5qC0lfD2uLJPt1ziUOgPWKlAQyS5nwgDdETKHadced4rso0w3lYlZDLU5UhbkYJLJD
h0bdCimiAoaXPOA1ccgoZkvPD49BP3RHY8wDqlOBUHF8oVvShUWSQK3lonx5XDIn39feC+Ss5p4P
/MmwDCrIWnLaQAVYeE1IsMsowEM8WANY5YEyKD1tNZKkDHGYaq8RHk4NzC729D8FJKGmegoEbpWI
LkEc2VkxQX9lp8Ag53fqZ4DJJrY3YeCaVoMm8z7xWIgsihCnbsY193Vr7NCvB4fzjgkAEMB4pM2o
YB1L6EI/N+h/ja+Md5Nb6zddATdxAF/NiuvYBbV+k0Hp1EzxMlmT58a147DrdFkXeFpWA47hraXu
m5PGV+MvLPVqY19vrXS+lFgWy783cPqpZ1CnTnS5YdYKvguIfDl9D2Q5JYV//sL7vNF/SuOmwonY
IxijF7PdYNArowxkznas7yvfBbD6v0FyWcQKEo/a0eqGQFIyco4107/rnLoGph8M2YQSzM5zXBAO
Lp6Mlm6bURY+UHXBKj/c95AwXU7wvn72dLv2KN3r2nXOg/rxr9ecF6kRSDPn6Muy0R3l42FpP/wH
NQwepjGbgXkucHFg20IFV9Glbrpz8iJIPHg1yGfJ9Xy+PL8InlLB1RRTb3avP1D1T9Y+c8Zm1FCg
CTQE33SqH+3AsPlPCvjk6Z4NJCj6jq32XkZbcdRJLsWWlCPWXQ+3Icjfs2XYCs5T2cI+Mzjl2D34
STv0XEWpWI66ZWP9nFA8ZCDMssnmljY9ocpzXwr2FCmH6HF4ctiCZBltQlqq/FgIkXnV8ipptQ8z
N5BEDCbXf88RBBwhx3aM2aoPgIUvIgNkM0uxC39/cd6XhgZV/GweeCVaoHMzvFBGKmEGOaw+PH+P
y8uZw7BQiVv46C6bCb8xUQlXE81Y/o3VrAV3fsOx+qaICZG/icxMQraBH8lxHIrgrleiYTZ1UxtF
avFDIIUrMdPOzqECqhJQj/f3QVPppPUunJ/83A0TFhlD1idWL7x5Wl22h9gN2WraijFilQlB4Tfm
Pyjwrq/IIIirThwvMumn2zHf1X0wxpo3ebVo3+d3XDtyGDR5GYm72sShS8z5C6bN+SsyZgl9eN76
tF3bRcv1TQpKxYrHAMMFVUy4dFcYeUjFy58eaMc1+c+sG5G78B1VcaXltzH5mASAGJWTrPArEPhO
TcD/DiPRIWfmX6FVvtP/ggM08RSgvaGVqjm6AufjuXI5ky4Qem9cexjeldZIvXar2EKgOxap7EWB
BwPJc14lcGdC2vACk8Z9skO8BHNogoZ/7v9i68ab5y1XJj4V3dxbTQWRMOcpKHhaucBVh45Fzo03
xxrhM7G9+SQKTGaKlHxSgglNRZ1uieHpd2Nx+3otgyPqqlCQPuOhfMXQDHWSQO4ySkjX6Ke4sTIe
RL0FCNe6zsi1bGVUQn2I+Q4TzQV4Z0IVkR6/dZbSR8U3y3dPi+P9wpiQPam7FEMzB9rIZ91KLHc+
1HU2RfxRuScg/pEB7Hv2YIGsLVQTfqADvsWPPaD4YtsjwZDezPCU/165KGv0/9hHMREprX/a79/B
lA9vrsXt45GpB7+GdCacY95PWsQVKGTGFaQ4Sr/QgmQR4Zp0y4WIVHBgWTEzeOxk/lTYnyJlBzSA
E6EuSiDq6ui7GTRWKltynmPshHa3qHC/zUSTVoj9FjMo+6EWiYBJTjYGSqvqhRZZl9u8pCHWbpb+
j5ij/g8jRhAlbJYlZWrJbflw2BXZtM3RYAzroAljxODs664RAsEUA9RdaF3WbA7PYHvcsylQcnGA
CbPDsirIbJYRd8MjRXTj3glHqRQD5wFd4RkMFlO/pZjc7ktqM5ZWRW0GaOtqwylXa2ONY5zXTETN
NsQJhxkHTvCIah913MWJ4R/rBbd4RCn/w/Ff+NKY5oVx7nqmR4KnLhpWUwrGWX1EEjErGGa4Fl0m
iF0GmtKlx9kxd7O9hyeg/uRffNv6Zyi7r/y4fmnGpv81I6hmi7OaWsay8r9p0JXP5hONQOrxopDN
u1Dco+2AcJk4Q63z+JO9DZdehpl+UeBloonVKqRQ7fcNvdNLFRYVbdE4Ufh9LobPEqQgZyAP31JG
pElBfbANB1NzMN2wvSYQr3FL4blOTzwrLMyNckKG6G02F9/48pgRa2T/2HUXCTdhNua7EtlWcLsN
Ptj58vbplsABgSYhLu7a1PCioWTSKHLCpPEiklp5c3fV8DSqFzhXmDr/gNKp7/5lNVuc5YiW45vS
7RN5C8ziwgwZUqtaxnlzHSdzAEd8WZLbpwBXjN/Jv7cHcblgvIQAmjwR2NmJ49Paf8TzB/cMmKUE
m80U+NvxF9asB7xkXAXbQFZUsSPSvBTDKeDNKoT5G/CeT6chskehh/VpiX15gh/sMZsCdai7InXh
7aEOuhjxCVQB6q7L7wupnyaS0OgvYt9KG6nBuJ5lrjBNI7+NtP/KwGPtX6wOiqltiYSI7dNNh0yh
hqKycb/icDWszMQ7p150Kr+nSgK9hmz1h+SuvCrO4FyRr2c44WIwb4f+KDQa0D5l+nBaQY4G8ohk
MveRObpomY7olk7+Vn9CvEfKA616FYxFlOSSxGWeA4PJjyZWD+PH1n9gixtGzIyY4xvleGGIV4V4
29Le+BdO8wwqyZnwAaf1gxr0GyCr1TTBD8lk3dgZf2C45PHM4hjO9Cj5jxtGCXGbVYTbRn8Gli93
tG1LyxneCTC8j5k+idylj8u/goJygPnxoyAKh0rr8dsI/yw9vNTMv7EI0oBVm+Pz5wJH8EItRIej
unIAZIBfuTMAmqHmQyfyLUlTqMD54hp68uupUcJtnKY+NDjpPq8g5ntkFy6Ke7l+VNvKY2yIgp/9
Fs6jiRdYKa2JM26ypRtuu0XROSDGqJgW1C0fE/kgXTIdIgr1T1tzRABMtkjIg8WACFfhYTgRzIDH
H36DIp5z8QjjHrDlGbbvARGBhTujnCVCbNtN+P/0ty0oWBho0ObjrCRsct1btIPO2Z0BWbpBQiCM
jZbpj2tZ/2WlIjkjkpT3Dyg2CF3V820254AnWl469hDqGieCTUuhgwBUSAfBO2ggdGo33Up8XKZ0
VnPAFlCuH8hSZiMnG9gdPRYltna7YIRiGrpNsvptVYoHj0ck/LYQawX0auAwv4rZbOmLvSFhQtit
G+VSDRMwnHeaBFXVa/y/9CNSfPkfS0Y5nMex5Be4pKmVJYxB6M0SfJ8SQNlejmgln33Qi8iJYBQA
IdpibfLDXNnIRxxdJKwjy5WulaEF5yN7DaAKWXBAqwN7n4M9MsmJEiB7YqMa502ujF9cxAPvRIZW
R9jEQNkHQacxpxv5spCcP0EbZqpORXx+8991g301V9mAwatEi6EyCWcacyRof2pyCGukqXl+LZRE
z7JFbZtnD+xG7w0wEikE86u690I3fib7dVEyLCDcrMdNi7LBNfqaUU8gx74W/tPvJZbXXwXB+vzV
tO1/CSo9zejxWX6DQ/irKRIWGZEF+lwekRbQvRQ5xzPUSLYXEmG1vgy7TE7mXn9UKr2m8zb3PbAf
fzpByMImdzArNi29ppk6HTTyVwLx5q/F/r+VqlvkSVz8cSxNHu/Kf1FS3SM491uDaHuogXKYAw8m
m8U0gqdIY3nQt9Hyo75YmrRHvOwmHSTBQCVUPecS/1e5VJu1Xar+gQCjQ+YP4LISxaJQnw+bUTLC
DYP9bGpiOQOOV1S0xLi+IFv2cbCPP8Vvv2wRbIndcwk2cszTTZ/WZhq7K91OQtbsiNV5vamYEUlL
6fMVAmb4rZFJFwcoNSSt02Igkzz7W9Xob6CZsZs2zPliVuwiX1yGRv71arODf/DrzjTvoUxYzQUT
uJEmvl9HokxoqG3j8kqoWbgzvxbptkbqB/AB8mMn3LaPag1+NaA0D9ZZ7oXcg4yR8FtfL4D/Pxha
1B21bFaVELWU2SRL/KNSbedEjKhqGkHKUBn6MNeJTMXU0dQeErO/nPhNVM49yzf61D4Y4XpTwcjK
dLKK8cGwOkC0CSi6H16KseZN3TyeHjEf0Se89uetDwvjWZ+TA34SR/EdOQYAUGNAHAqG9BsJ8fU4
n/7CCefbdj8yWuSGYAT5oqEQPykmeCRYDaUJsKoHBg/JaK8t19mRBfu/6S77WfY2nF2NczlHUr+2
g+ngvhSsyk0HvA7EhdHk6f5xHP++ijeZX31qlkf40cNNy36iE7CIrS1hdnemzUljQRjVVtu7OOae
8ty7MBDh8QvXJF3LQiQSGS+2WYnZFXsgQR1Hksdxrf+zQA/ScDauIILkAmzxoc6JJB6ooLUMPJYI
Pl+oI80HNe5zqtLCFcRy3rFdvZvh+KrAUuKgjtUQyd8hB3TiM8Ftea0tVGMCKv/aojazJi5iIpz7
Rg2M8TpoCrjH9gay3juQY4xVGxGxCHgBMHZCFVepyvac5MNpjiQ+dUaGazUobewp4NUduUQOu3li
4+Z+rHIO19zk5ZO1QArAgWH2BSdx0uWxjoP7Cf+lpHUXH0WXlfE1nTCJKFxw4jwyLpSiGZ5EntFl
CTA2zJZu66o8Ud5UtwNLnM5YHNMX4wUaQhVOq98l927fYAaK7g8Ykp1a25yrWZQSfGYXVnzhgt50
UY8BsnAzSS9UyjrK171L7mDFbDlv1QFEqE9XmLqHtqOMYm8jFIL6HEt83IOGUVdgSLOZG6V+GI1E
yBam+UHdxdil7jJziuz7RfgbZ1X+q3NwhQmhU1hq2KKo14egTmeYqYE14ccJlyhzymqisA22g4rK
dbVDGc2cIN8osgSEt6g2Q54UDn6yW6Hp1m7S69GpaintYkN0GjUWdeU5C4uBOeamwnpbZlVyeWID
PyhC+3tJZi0+zu6ZnRe92ZnXw8SS6lh0kxYEwJXUt6h+v/ZtJwnhU/8tyhTnmeTeZFqeBd5FVwme
3gvrQEE794F4zXaQeZgyb0jQ/xyFuXqtDDlLilheQkRoPBeZ826MOk6Q/9nCIoKf3r6Xi8v6bht7
aihVTB3ZHKzgwUkt1x1lNxkXgayMr0Ncm5lH1p1MSfHSTtbswEIlGrA3WJvuhJ2DTcCZ7HWlT0IH
fkc1T28HpU4oJhROPuZhfPZtbAFzLokNJyg7msrxdSeJcJP9YTJGVU7xOA7O+JyFVfnz5j/IbwUF
HM7kTu25vLrnlvlcLSSmUSiQczKLaKJ0cc45ygBUYF6SDRMxHQdjjexZZXz4KzYyPGBzT3BX+5q+
RvbghyaE6fzVAWJPC7teBGY/tG1rVtVVo1F2h7zIXp129DCVCJJnrG4I1hZHlUQ9f0GCC0wePVB4
p+V3OAH6XgvcOKPRblHXj9/LWDjRdU4wAFizhN3EPwQ+U/R2c/5s7KnxfXsqosTPDt8wQf+ahmQr
9ULCRLWrECq7cCQk5Zk3fXSrEyeTqxKXE1p5Uh0+7V5PpKDIB+Qu8u1UWV76IAR+MWZttiUIu+Qo
xoBCh5jMgTxyX8r+yBZZkRCGTGMdODscLEa21URZ5GJQIjs4i8aX/HEZZm67egbqpG9BhYBAVyir
1FokrooOuGDEXMR6whasKgXXzTRVX7REDSmuGiHfMtJD5gYr0yjN7T4qfemfhZbMRHii/bVFIpdo
ewl+v/0RXRM2zXt7PrCQ0Dvz2zO+Vd2kwQUZMjknsUVf4mM83jyCVwMzVINSgq4RcW1Votc3a5Zs
+CRJwMQ3lLHvxXBNTp+HQKALZtPij0i8/1NbVnfgFfGbp97pUWOmyA9oZZhjqCmSHy11zLQZEbv0
DD8DJ0pFU2bIqmxGWuAbsf9dVMgP2213btfCcWj+R4FATm4O8XHKCRXF4Eo/9Ta5s5mUtAIy+hjC
ZVq7+ZDMYJGpRtggFgY7Anr9lME/29zGaG0L80KlVR/uQ1gOVUPLHBwAryOMAnjgtO5Q1s4jE7MY
Ei/OdcM47lutigW0pTWjHLuV8iSCXuDpXYYHrXeMvH+UZjdeJJaiPPRD+YabUSpDENQieioKnlXe
+JB1Joqgld6YmRDOenkltlecjYQkP8iM+zvpYxeiTPVHiCKMMDhQX3jgeVsrwmXy5lK/3OVlah7q
MPLvYOW0K/ev7B+J9k0uIenPgP7hPSrdulSC4LhjwwPuXHqd6SJ0heRg1Vr2wvFPAxuk+zAWNyjD
ljjrMfbpcEzO9bwXyf1IVwNbkNVb+S8eGOsl08/9uT9OAKn5mjbDRXWYqDPWnq3oicJNjwRkzeKk
ET5/hbXV0/r0v2kQK/BYMIzBJ5Tnkri+1Wzd7FpPb5Z67xlBkRicZl8ZynCz8/CwWIJ2SMzW3b4W
xEZ8+Jb4pSROxqRLrtu6u4Te5HirWC2FNCINi29tT1AT/Bdz8cANYKqDxKsMfcFdvIf2qrtXEdHU
FTfpAbNST463vzm+a7a0OfmOOJ+yCccfPIa9O5qC5i+RT4yBMqb7O60EL5+3QhGGcMjX92ZbveLV
Vyo3mHUr+jzwaS4r8vK90PbsecwR338agDgRwT4VZ2SnUG2CIlj+FrPLX14DSs1KYOYz9u9Yu0OA
8YwgUC0+V+0hNrPxMeDdUBI6q9udv0DO1GQ389vDKdbvfdMflvyxZoIbJTIsSinQfkdPTqegNG8O
cOX/2OZCrRCWSUyl+eTpAWurDqMS7jCylTUWdLb83ulg5G8o4ZzE+rFBBKpQ69BEqMNTCxNsBzoO
1iZEcWJAIbxiW7B2FEPvD2u6yTQtueiT1GGJb8JG9Y7I1SKCtaSUrAiYZPoHbN/LpE+2f/D89zvt
B6yw2Eu98IGbwJ7C7NFKb2M84kTFkPRMOyiOD4SnizEahVzF8jtXnRKuIfBfyIUBY1IsZDYYa70U
jsNw14KK8sx1XGG3sKlseZWFItsAgmA4izdyNqkfZ7XaI0v2dzorQo6l//ScALorIUG7BpZnsj+W
vcCmfLdbblgpOievoMvx1b/NZcHcziddG6M7srupVmegphUvxPj/zisogFW7uOFCYyXuKLrMTgFp
9jmrLMX8bIcShLPGeehLt9z68jL2HX1otVbPQGjy8DGRffy3gCO3Pli++dXyohh9ws44Ewg7rNfN
C2x/K8Ut4i20vheRvLsHDjs7AhX8yE16Pu/bRNYiQfjk8Z66wtdr2MpfI9NhDZ0wSTPc6MN4al+m
WKZDB/9VuqZ9PYTLSwXFCLPoedezdG1WTFoMMzFhWjxqPjn6R4pg0xFJJqWvkOfWJhvP36L66kmW
TW9HillE2jJIDFhMCb2n4oIMcl4YMfJ2UVroHGjHvZxuB3zkukGxl10xv/tgM+KBuXoOgcOcheht
PfIKZEgk/PygT+P7lMNDGlD6VeQF5cwZaMSDvoKAZIg87aq+pK8SG6wmYcCLWYBFyYlnf99RtgFw
YAO/WBzcxutYnG6n+ZGH/I7NTkjBLzik6I4byfcW5KIw5jF5oPgv+pD7qCM57TUeTvJ0Fer0oQsf
noOeZU+9XuxohVDpiLHmWTvvEAfkeT/O99t25Xkgp6qhKAc67rbFPN8i6Nhoh+2ZjV0LyIPQgIu4
H6hNXe9wfnJ0989LysXvEbnF7O+YyRQEEbJMGs5QDk+PUHZuS4Ph1VZn10jZ7O0JIV8GWzYIAEn3
VKgKFlSVxluS989fPjqwknVZOIOapY+c97Wdu5BhnqaNuw36x7ct9OnJ/QaWNh/k/j2PjVZsbiFY
LX+V/VpL00BTcdXdaI4ak5zNp8VeVzidFRM7kzRxdE778t7kNHkubICkhU9yr4RHzKmLoWqnzCFW
lBZoiY4dhG5G8DCkm7Q5RQepiSz0VwuVlNm49h2RH9HbtKq4Rw7uLCxA4ZhEo1jlD/vdY6MyOCsp
iTq4+5CnAJo8tP49+luTBt2MXcTJDFSZseTPfXWDh/JU/qkwiVCw85w13dGghVUhCNwOlnrb2zrS
brDN0wjdHkovDs0nSev/3kkUEhgjGuBhZlEi0RlCTFSRkz9ebrlm6qKQXagiJla3Uxa0AEacYJvK
Wxw1aDdtTDkPFKEbxi7UUiM+MQaVlFU5GDoKqo3tM6LNXLv/J/IR+M7rZaxFH8zyeYYgsMrPHRD3
9kWpc29E8FgU4YMAYYBnyf9ZBsFNbi87H4ka2KFoxuiZePsMDsB4JKg4YKVAHKCMm/FK2JK6CfVs
d3fVlVbRtZgyJfP/8DGxjOB1k93osandXKaQyC5ci2BnE2+HkwDXL/6sC6GASDc5r+6Oxwea2B1D
J8/g/PMbw+M5xkrbKoyi3ryD/0ihac+6LImpkiBa9g3GMWK7jTXQD2DptAkav2+wtgAUGMbuvvrn
cHZc68YhSQ+aNNP01ehT5AXUJVZmvXWIpAttsCsEsv2fOfYN587TwNcLshjaD9WI8i9gGM7HLhxg
OLrOXcQ8AJaaUTrdwXV77KEt/yFNPEEEEgzn5GssABLmX38PAoJ8jK+lFoCqhP7Ru8gaacEhBHL4
RHIAoQ8RoQDGdq0Eh1R7ERnQE9/6xAc+nNyTJ1DdoViKoEl3/PGlQ2xnaDnX7RZY4bv3bm8tMb4s
iUmYxfjXmcgt9CcUp/EDbXfoRnzcOXlkFDGQ0vCS9HCn3EwPAaR5yG8S52Ddx6m41wsPejGkuaa6
yxPOyxbF9D7qeMklYLN3XgI4W9SgJSHSOPijlHsFY1b706r9+otQ8zmOWxKYqYSdVrUHCTV0VCT1
9yXiMLQ84mzHpaHHa2jVdmENmKMcZXqX27F4yzZ85ruB50XoE9zTfDS7Ziyl98iiShlR2ngGazZN
WPEuTbr+sJyZZk//3SjbaXjWr1PqyqfkoXMmXm+oTMBhmlJt0HTWFF9nK+Un6YPSJinE/XrktBGs
zTYv87QFxJTZmM7BRzcYxnUMrI0Io+U1/GLoJEAfXoTCZdOF46GKuAweb937/MdFeSse5yjnug70
owBg6eUV7eXleN2inn1qYCNcJax88yybC1ONKR2KoA+RqVLRJ9E0C9FiyY69zLvQ+PVdof484lIS
n6h5lZHB6qauJnXtmlhk2MqEv9F/dB+8h1wrLn5FYs67coGWuKZth1rEWbH7s5tluyqJEZrZSoDG
1rDy5Ep2CaHqL32f8TudV003jvHhqZ0VZTCMK43E5a7O52HV0G4ZqqaVsu/Vi6waQCrWNlElD4Dy
X70c7ocycprFI1ea1rQlNaZw8D2vO/bgmymExRKjDIe6Ddg2zHC9NRLBID2ayEGZobZRCm3EsyMH
wDy0iXAAj88u2QrtTc48pLlr7laphVBZq9DAm0qoGQKjmK09AAz6kQFP7KJKGRcgZPw+TjThzUS8
buOPmVbq98nu6NUyP7CzF0oOmp/FUhj+t1teVbguOYSeEKQ7a30Ti+J+GIcKlmhh1NuHE3f9Q+mv
vw3M71W20m4aP/GP+Ch79mdLwRt9fqgIL3Gos3WpPKmlHG9Z1sAXblzrYRkqolLCfHlo1tDKRVgG
afkaq/OR4w9lfVjujwPBKbfDboM2WMQ9ZiKmxydFaxh1BB5OQITyL2xMjc/j0SbKh7MtOkVr3ouE
DSQyyfQN2RyCykTZHjS7JyNWYCc7Gk4elbjKkh4ScjW1YYIdf3qvefn7UfplqVr8miM1B892mmx0
wKZO4V0ZHLVnUXlt718r164jK80VugeOuIyP4Wvxlt3RAGdbLdVPDk1m4w5q8gZqMEuI6p3lx/KB
FQbUT8BQbLbv4nzka3op+weZYAJK3TTI274VB/gpvKyig/ltz7XzB4tFw7Pw2E+/00VHBhsErn6K
cNalgLiv38QjdYRyECPrx8fTzobWiWvwmFBxkskjRnFR4Mj1kTbSRcrkg8Ux5KftFiStRc2aM98i
e9rBXj00Bpf5N8p3kuRJKFNosjjNnoMdmbVCXdNvptTSvuvounPAY61Sxus3kMeCLYwfl9++7YGY
AW11PGh346DYY8lF5e/xyFSUkxS29uDWSf5Bxsl4Oniqi3lANpGf3EbwX1uCoOUKHe9nkB/vHLgm
x7RVUnv8+0DVJtWIZtDu3lCXeLeGHjhIvDtp2SLoXgNpKzFhw72Vsy6+78nBWIjQZeALnXZd9GUe
//eJd57HqB8xMQF3OylH7gDfjAUuVkkZVbb8Ma7uQAf2k1n/Lb1s15HlLYaP6G3QilUIzAB7NxYu
/ZmorUmMsYQVMpPwRWlMp2B4CXdQIp3pooa4jdjkupv0CKrN6qKwCW/KKl/8I3M17fY/lc2lw+mZ
rX87mhIuOStB7GdI9i0Zg3abscmtyaImHoVi69WudKNthunnf/v0Hrq8KvBxVhtZR7eX8UQkaL21
Ih1RJqKssGFXcTSEsDzPx4xxjUi66BTXBHExsekxJ2s6saJzIPwzv01jAvOVrvYx42wWix0anJER
/OXPWU19VAFsI/0bIomhuqvEaanv9GUCrPEq8QLeIyNsPfkWwFlG1Wee+6hilvDRvCM9t0E7TnbR
jXCq5eV+UgLNzyC2v0+lLUkf/dSz9is6mzFJSmntB8iyaK+AqlpbofMPEyS1a+BPGbNrWSdye5lJ
WzUDy7twMD9obmcC8EHItYbADdMHoemmITutkBvtZzwUtMH9V/23Wz9OV+oeYCa7He9USrmirmFo
R/o4YNQO37Wf7PzBKJkhgw5qzpGk2yLXSks886Mr8iHOId2vD0Cn1NRfz5Lm94fGm5o0X4/FzjZg
GjGTpjkOjCnJxwHHk3pvALCv+DP8R4oSSUIoc5ooJvLcTEJe43MC6lgpsKP9dLl38UKmEAj0Svqk
Ud2mP/Z57oTpStWY1xryO5LfFyO4Tt3gt2tzEoTOA1ABXFxqxTMU/kz/gVc19lxNHWtlIc3oSXZx
G9kFdolAlTUi0lgk/iiQEnLL1B5D6TiScXKt2XdCly4DJmNlikHLZRTLqGmEkNzDSgxomPaiS7//
DpilejRgpvskd8iELAcOkaQeoFc1G2E5IZUOXMNqlyVyqc8YYkKqrCCPsrXiV2fAuj9tDfzp/YGS
/C/zZveJWceZSSVrVxWSiHcNxhTSVWfQJ4NKSCKv1NRk2gb2LiP+CZrzXjT1WCUxQzkGyQyMBiyR
J1GKZKcBWsErveVOikKkvegrUBdvSpUHpOIqS9mywIzks9n8A4ehhrq663xS7lCNwRDT1r+TwZJ1
vSQz1riqlY+0T7ek2zEukTFwHDO9Nv2QBwf1p1wMk5Gxt5DKa+znNpdhGt3BQIIypY0V3wvgkxGq
jO38B2B2n1Vc9q8O3lUWxMbZoLjj0tXO6ICUZKcRb8kJ1plyzb9DE2VCKZQtQ2jHSjuGdvTERR9T
MJb2MGpfQYXBTvMJedNKIlR+vYthdn3iM9HloIKfgW9WyFJYoIsqyukKOExNKhwGv4eki8i1Gm+i
9menTYUFp8mRgJfPUx5ejeal+tTwVkcDwO4VDHrwj+6SpmYHGD+dWYWp+BV8omyMZJ2S4lLRi2ty
A7vOYxRybBCuXEtkHoVNyRlXssGKaQYHtUzHcgw+QfWHT09EtPZs2oxBVS9PZXVRCGJl3px20A3e
90SX4i4Pc0tIdX9ae1mQ5q7khxpvTRexd0uZ1btsw2DgALSEnj/3gXIpE4R9hQ/9okm97jkPo2DT
/IOpAbYKfw5+IB3JAtMDy28rsCYQafHnpBNywWQaNNXD3/df0d2+P+hYIoI+kNU3ASLnqDW1LDY6
ecQPx3FxD3NvX9Bf89fux4TD1mbXbE9LmNN3AuiptoLU150r1V11/4UbHShJfXIRxAI/yxj6JdS9
mQDPcDj6GwNcj2HDFN7PYSmWHywqIPquYFIcMP+5RkyKDXbAk68KWOKAkWh67tbKjoLBx0oPwWxg
v/+Suv7it/XrhzbC1Yd65pBAOieAsG1edFsl5Ov0oXq3JT9e18cSQrRiJ2fzjwCt6yVEq1rmHE10
Bp/yc1Cu6Xb6NCP3Pcjph+6SmlDlNmXdUNmCnwnx7x4IW7tcf6kg337TAErmx9wyEkZ5D6b+tzB7
aH79FqZzxwM6o60HCTWgmYx9hNW6isQatR/0PvGABqUU/kgalD8it0MD9j7lFfNeRcIKngJdhhRa
/G6JLebj6t8Ofo6lu3UpprxEE1ro1DwHebUXrTahgzz0NSA0YfzJ+X3duukIMWoZcIh4vxowa/4A
Wl67ENykJhhqVgmSytJp26CB2Wi9qqUVtjx+jTzIZlygzOPrdwuHNW1+unoN2FIc7xiSZJ5lrBL4
qCRXnAWEmKffhlpjF2O1sZlKz8jPTK7DfFGy8VEwlGPpwUzFe+3/+Z8zxbcC811fX3Wf5EeEeB3J
ccTEDvACGLpgXs+l3mIPexH5qQN9jzllSbju2KZRA5coa7Wiw44wM0ItQD2gN9PScEKpuK56E7mT
kd8d4sNVInFvL9oEvm2ra0R3592WspCKMcBx3KaiIBL63FmBM+BEhi0tL9+ExMn1d/jBUGEm8GQ4
uTIj2G9O+ymmiqjqRehlbimnFLj7mQio6e9dUdcKiov7YJxVJqJpcwPxx/gdsHSVBmNKR/S/Z9nc
Fi8riB3mhMuusvPy6+BBSzZb1JawTqiKGIoMqm06Nxt7a5yGSfLG9UUbTfcUOa3GYIFEkCS7w5Ih
J4CE2t00DxPSMzP2n/JJasdJxn2nHDYqO3nCQiWqsRhz+e4nekd+em+QuMt18BqSsx0Mq/bTaDnB
QJAHTXaPTdK4FTmaaJ/Ozb7sVrXACc8thEvDecGT1Nb9B6GOSULP+aXxvPnovSsyMBDcKsZlpRRx
lWcWoTSCKhGYojnP903OJKqnmGqHG8Osmm9e/9lbFltlIPZRD2jZryFE2AOz7KlY8Px41wP9eJsh
2cw1L36KLqXgj2kvtKrx+9uHB8BxgmR6Imhb9ICDFQFAIwMqt/+eqtmBoE/Ha1UVYR4L2XZktnjM
M2MM2sdos7erPXs0QUoKDolz7zDMfdR4hVpqaG9IwLnlF5cKdySC9QjA4PG8xF8pm/I5P5wgYG1c
7ceoSYhSmgLBRFaTCUpkKbGhOTXx/jqkvhdCEZSA/Em75lyGXMKVRoPogOtazJXNtlFYLgZwLfYf
FGnfEK2tHj7Uj2PhsZA+suN8tdCslVOgT08d4DGHeTQhUMLcVijnw8+gDpP8rp+mdivfE5S1kJFs
4K9dd5nOjXFNFbIQLYENomIG2MXdirrneds1QFPzzbwzSdMupZ0c0veTrcLNq9C1CtrW8FTeSolC
7IsuHaH/5KgxDypjIE0tSAIvEf46pg+fWohxmOZ3K+Lun6eHQggc9TlChz225ejk5a95VzEZdB3i
wvIWf1pFXXGWbMKCj2FEgijhN6sxo70eQtU5dUeIbn6OzypDNAFDZ3xTDak/pPehgaPxLDe7/pFH
ttiamKOeVbWegD0mfbxJA9bqFOtZyFP7FT5oN7N1C8jihQOHVBvnNI6r3SdU9nCVU6XJu6RJzD3h
7w+YW5gizmV/A483Cst6SF8GBAlxOIEPCE5AeieJRUgNvYP/BEcNy/lBkiuAUb/TBw0md1NXZkNn
qI4cuQiPnpFkRLZPPVnTOmNQf7wWaydXJGPlmjWqKT4iIIPwEfuRlp14I9ZnevoXzWEmS1vxR/AD
fNrd4I+PnekHNPDFz8EQn9yVOtJZlyhJyNENv98qjl8g3D5kPoK7zsAXBmdbMWq0S9bLzQC20cSR
ByKPfN0S7ZWg6tgRX0Y1HfyRL1QGx/eaIRrQoZKaar0bsICbPmeCgmm6/xrIcuX+GorGxPtITMjW
mbGp3ghk5RxxhF5ROyrIH1DKsb4StkoI6xEOrX22tw5Cug604pya8LIyNIO5P6wc9tfJpg6oxy1r
DMAsLEYRP54OpDVT9DNy94pkhu5W5PY6SE12w8ltJpCWjnnSUPtfFRH9Yww5tACYhSjGO27JpcK9
4C8+HNtZzBe8nfgOLaI1zXgCrT1OFfi74OWQX9WVQUh1lcE7IZJtg8WNJaGlbYE1cPT1/HfwjMhV
suLwVbq4tLdZjgsVkdIZb0lBTimckvVDVOvfCWiCWCus3av0xpT6oP/lyCPbMhZUlN72pFoGEkyW
7FB0twYhzqXOdNc5rNJLA7Gq5PVa4FEWwe/t7j1zaQlQguDCwf6l9ZQ7eP/0GdVSvxnXZOPnOQAa
3xUPocvy/oQXemnZ1yX/V2FV3vAWdlNhp5MpA4d7rE1MxHCD3Koa118SNaUgS4HtG70uM3Q3Tsnn
S1GzWi/7Rhyrzd+7DXeoH/qksyNmMLg0nFL3DpHbgtOfH5WoReuu2r7MOuVwZceaheaVRTH6w/CH
ADEnH9ydN+fINsPWuxHJEt+OE1Bw+XRnRD3lO8euRikIP8Ud2lTDdAe+/Sfi6Ddoxgp/nUY1dszF
Zz4x/4nTkIUkwR4WqB9/3h4obpWkYMOImJMunefX/I8wAyxA5MnKb2GwcsK65sgAS4AomSVitrcB
kBrS8ZUyWD1F0fxL5RI6PsFpbn5A4zkgEiBLYDYEdD2Radq5z3Y8xjnDqBlrld87+SqAoFP22Aku
hGgmxnb4JZwrF/MktQ6PnJ1TRcO3G8GWB3n4n1Mh/+CI42S39hzBHCVeIu3M8kZlVRzwMSrhbvUv
3EeboYephsTHAZbp0M3Pg5pwuC+kSo0Jl4bWipQXjxiMJAe6AQfGU4fJGVM7qQ5X3+jIm+36tyQm
EVByPXiRVNEPOI5ghrqf9aQEyO8GuVLEaE9NAqfRvTST5tnZKiluQ4T95BFD66sTB+6YaOGGRadN
z7L5leXkPL2V3+7fKKIdEbgBUQ3v23RFLeD6x0OZHiryfOQtnAV/2v6SoI+MPiXBSEPkAQjkVJ3p
xCYBnZbskbctls6oI+gM+0ROFvkk9GoC8Y9+v4lem3NRINogRO0w9AiXbzIe8esu5GdudXBtNzlL
VdEa/HxRULALHyRft9XH5P7w0Anmb1xoNZ70WMKaE/oDiJKisU0YKbFvwqxCqT24B9x94QVKQXH6
D1KzVIHhVnQLqpiBeK8soyMakQ6Ly3l0MeEr/J8lvHgMXTgD3d9/qLZUmmJToAGNKMgPlPxKXJYJ
O/lFERH8S/1hl/phrgmsm1sbu4hqOmsbPe0niNewWY3LM+W5UDDEzWWYrlURi38zNX/auEDYvV4F
B0knwsn7h3DXgeRH2RdtpzVXyh7AqlqyojeMZAaZd0lNYQdbyPeO2MOE7yO2jyWi+3n5d4d3P6vj
R/Kfsn14Pcv3wE4L1hr1UaJtMR/lUc9T9p9UOqkDeXwiG09zXErN34nxy+ftX05lBD4SVFvGuSme
dew/oWtG1UdH9Hf06ANkNQhXtxW6A4Gcdl6Ja6Xfd2QvuVqa7UZo6Ysyj/IaCyFexXKYNgEl0+CA
b5wUWlGsVh2sV7uPjl38ds8/ccJsQebvU2Z3tkl8/S4mE9Qm/5W83zof8xEPgzuspU+KswMeTTtW
DT6K6VKbONgQ4lcI6wSKkMdGnxRG2MXWKH8GvnNFOV+6a0BTX2CQ29spqw9mcrtNn/TM3HwZ/4gX
Y15Z56YNwFQ0kDVvm2laDDLKu4k3NPbDj1416wCYWdapo7f0I8BbqiKn5AwpjWTEW8V8lXSr0l9M
+wc2VfXy0R/LxefPcKGsFQzDNHvfEvoWjYiSiEssj1rRAPQq17ob5l6COEj33THfWDy0gtEgO8yC
7tvrlmLwvrXKjItxjfdibJjS/vHRfNIyz1avULJen86WbngO2DFuh0SHvN3R5fYwVsEr1Am8vf3f
waY/8cFww7tuWCMMkjuVb7EhEHSu5EkacMFegR8DTMg6mBKnrwTFLvt10ctNk4bcCtgcvE6CTXsJ
ef1tBGX+1n0+KYlwERJnZT7zlIvqD+a+Gsup3br/s+dI8/xJV+OO7XxtSu7FoFAd8c5nZ/sZJ9/E
TZMkG8+tQUZesbEcw4na8IRbPpEeWgqF4Zu+fALeDGDdEtGj4Z7yFfPh48CXVUx3fxY3DAzyBXfZ
DRIDqTj+yUJH+yQoo4eV8LFiNISQmu4y0lyUCu79d4RfVzKncJs/gBNHM1D7VaTX4iOAttUkuIha
5y2vu0kgRZbfCGVF2b0xvMnqQu6XE1F2T3HrsE2cMIgg0rHgRJMkXTVIBDU+N/8oJOUgAnuq/Qi+
Jpn20ucUcswNNYD15oPm3Z4GbMm47iEWXO48ohYtmj11ZqjgBJ0/PlUvkmC2uUABeMsUAhKFgT45
axLiMQjw6cWkHwYSRuQATeh2BSxOKKpznIep2mtVTZiPt1caYOXS6XuQOtLMRf05Cdbbr8/ymaID
qOuoVYlUXY+vhpJz0qeXH71kjva1kELB9b/BQePOq7uOuQ9okcM7fR1Bfd8aWUmeCxw1Qhud1Y/B
yzCTzxWqAldl1UlEHL8PancWekkdfQWuADL9DPgtOl2YjK25nSqR8qxGWZK31lnltLbid61PRQKr
1xli1PRxnr+IT9JOST/3J6J4vOeWz7dmyOThphGwbuilAlaPPU2p3+8eL5FYm6GTUUC31hNT6lJB
0yDZXiSig1JkrCgsuz7d8pKdEwIgqcK0Strm+TPzX2KGJLXinqrhk4uJsxvoQtytpV0jWQ+mMnpK
646qbDuw3i/cHDiyfmnBAiJNj0cj7ofIUQSYoxBfGUBzycp8N2j0eagFay6QTGCuuVBE/jYU0d8H
qInPT6BtwxmmdNVsnrvzE1UTReE6aTkiQXzdusFkE7Tc6v9PgEsxCQMM9f0VY5akx+Wrf0aulgPI
KbH99yIknZ3Hr0nFoGpTcMRVfkAzzY0GtCHR/GcbycWgtjab9rQKSJG9Bko4edcNepO6zdNZhmhN
xjkBC7THZk4usRTcRXhloz48i4PPmifXd5D1LoVtP6f+ar71tUR2cU/4NmhuUZSzvcttmNYhC2yO
X6PAjYIC4/SwirJuQOyUSopXrhcmXKpTFYuAPqHaOa7OEVNtC2Q+MEDLE6C4xjSdqziO7uQviSTg
gnYClRHVAgGtrdDbDfi5rLEoaovVTKOYairkt5f7W2MFcYdK0KzGq2uiyG0wTND792axdTAFtojJ
DIvHDXmo4kAt0POcs1RyxvU74DxZ6WwsQAmUYwkP9jBfxSAcoX4oEvJoHBc54NbDVa4Fxvysm2Oa
pRitKEwaevK71a5M4Sk3Kc8STO0LhVsZvGoFZHyKgkWyK3RYOsLG1YNvfxSMgu1XJekWrVA9Z6XJ
ogVK/+1us/dpnaytIamwIr5JTHDCJmax8CeZrs2qe30rTdMjlt5bxrbSF9Hfx1nBPV/56i5pFQZg
iOX7cVKu5snPRzXiMdCcFok/xSK0fG8GkmUjXatwOaNj9xUPOI7WQFHPtF+b2kAtjJhczN8NHv6M
P7U7mL6aePzyukqAx2ff18ki6QUM9FVZgjjkT+qOYHFfIXDm52+J6iUZr7ljCLHgx9L09DRtgw9I
AiUk+icSu5XxxoweWY5f8zf9xA3sJeznf7HjweymfsCAeJOG8Ct14/e4vM0m0TjJbRex2ZoIzcNH
tXC0IToVNdK/jOVJMo4B3paDr6fP18airC2Hr41zI7est0mp5CdsoueQA5XVoBXW0Tr0WtKn4+HD
yk6llvJ6e8RWEu1vUMW6xhna+AFoBVT7ZEWSsoDLBLA5GK5frZP+XxS067094G4FNLf9BJTci+PE
vQWRzokavpbzKCok3qR8ZfwLrJGPEDIFnu7wrHLQ524GWeLjnl8L0y6raDep1grXWABTCSi7LeIh
KU9ocUeDux2I3Y54Jb7neqXC605pZRYreNnjmjFaweM8SkJk6c/9hdGoJV0n1OF9AXqg1cnmuGKX
y1ib8H/L7q9+OCHG44bG36kxbCujglc/vTS0d296pkRc1fjxk6pLMMSTVG5WbKRXE96OI+tRhWtn
Y2H46bxuFLlvaYUnKzA/j7hLdr20ym2Xey/Yv7oA1rTCHsKEE3z9XlP71X/8LC/sao2LnbZ7HSgz
XnwCOCKilIG1BsW4qC0ZiEvetByF1abFU2W1x6QMA6/CoaOFZzZg3CRAICHJ9Wrj7n2QcdlynxpQ
aqfBiDKr55l4ySziujcjJ/r4+5KPoMHecCcWemc7rZx9JiWP8/QJ8AodZJUcOkHiDeREq1PmW30t
FhyNVt4fCmXOo8TD818LMv9DToZcLOmmN8Ciia5Iz8CUBZ+9l/3gHZ4ZekiM08A8hThFHNZ0ENFe
x7wWVnzvXKdUxZYYoZf/DNfrcnD0I7r7SSh343Rb9HfFpNSUHVkPjj+mmHKqIIRCK3m8s52MDbEz
FEMd2Lmc/uwPuJQp5Q8rZfOL9w+AXPsFQeQcoCM/1kI8kQqGkLXNmlrc1xO8I+MwNLaXrPaX5yoO
zCGDDDYleopQtOpwaknyg+LqZ8wyVZPEoYAxaJbbSVOn+My+sHzRTMyCBtx7Gb6yRTzNmUxedBO0
Nc/EljCK23BfV6NzJMp2ZWhn3JvOWXhVTqfjwrCNV9x4OK0PyppfLM23BJenZqrQ7qlT2ZQN8Tfo
4/9WLxdXnFCqnQZsAYIIxgsBKsz3XE6PQQQmJg/bNu6V/5HnSiTLM9BJCPPstVSriY3Ddt6PpL+4
JSEHSIpIK7ENMl2e1DZxBSHNotTnmMq2Qf4i47YcbT7FZ4HrSy3+y5PpGsC9uS2zeNqpCVYZqOPa
IuIMjhFFNktwG0WdJmfhd1KDuaUdMbCva0YXcpQkgQhgRtfHRDGh4PCQzT7SdWFiKeBRkGP5eZC+
qMslQmlxEjrflS6N6T/7w0PdSR0edF6ARskggCwOkWa+/ZLazyBQqe4IVFDi0ab6MyBYUtBdTi9G
B76/YkQ9KhI7d9zbCa91Cvky6OJm6tLNvzVO1jE0aIngeSSfNdhmV0Q+/qIAFkzSWUYTC6hCGVRk
GAOs3hBja4Bvz0i/RHRXvM1OCf4Uiiw60FVVCRhk89JD5CiR9f70MBJrgsOCs8qfSu7GGhwJRiNF
kAQ/rku1bcC2gh33MAkIeZ+yoiiCkf05/sh1sG0GtIycZtvM1AuigUXuGU+6i9qpaJClBWSQG6Rt
4A4qoFKp8U1o4QTEK7/Zz64u2zVhY1n51DlwxgOH20GnyB54WM2PNK9ZgjA4Unt38RXowYpHufEr
HwfD1pIPge5bu64VsLh6Or8iI7ZNj4TWqysVhOLRU/Rcs1nUFcg6xB5w7TFwoCN7ikVV9L4Ap/Nm
Qfi/p1u9bDTIvGar3LqfSZU71/eZfwoZyyQJi5AAB7C8WpSXa8B1XmesFy/11kvMlZKvh7aDqS0N
TTqyt6rfO4h/KwhXPgnTkAreb9ZpEgbncP+j1hGCsmPz70Ir+lGa3L8yeprOAbz514tstXGG20Ha
bP006Ca8bInj0139mquQgrDpy0htrC/CMVweOb6CVcz5jhkWU7J8sX5lPi5XuHDV53Sv22noTsma
//3TpPjOrY/6VV5rIztL0c9eSxicbbPmK1CAKt5AYWvTYPStaT8m4J7JQpWWc8Yu1QB5NtAghB7N
luSz5EpMl2j/qT2F1HU+yko1zkl5GDugHfdGj5FMq9ae7N6N6KXhDCfrk3z1XJa3disUFSl3vr4S
h8/4wVyExr1i08Lgy32HWCozXUwhhMHTYWYCXk6sV5xLnlgoA0o7YmBWvj+yvgl55enXzl6cke38
Py70CpVktitZJpnMV/ZEixM3cxhhfYg+V/lcI55xCTusZHAbKiQ/XytpuDI9Xi1RvfP2XjXRK6CN
4jm691nvBumrRYTlf2gqWmsL7whsf1hsLvQQc2Q/r0Y/MRASAtvCSr3GhEZv2oCczjTCcP3EP/gS
lSaaacELH7uL/OgzGYF/BVAUGAgpY8q63RNt95exLoBvc3LcCMJLvzOZAPaHCGBPvpvH8xxCQf7a
kXfRvjJi3JpvoPYq0Mdr9Tp1IwGRHjz/lHgD9gFthcNIxlTmkugbLEUqSTyNMZC5AgxDCF0+95h3
GILmgrh7rQAmeLIuwdpp0VvWQaNwpQM8gNPN99eK8kq333BqG41eEvdv8bQKRj9UhQUsIzaykxK0
r67+LktPZ4IVHiADqn5KMwoMtWCW0hwjwv8D5wAsTWpEGamkJDAaCaAdJK4lu3p6VuO9qi5h6+l5
oNVJqm35VrGobU10SXc2yo2entw2IkDzIcAmgKiLmC+XIayjAsQ8UqGKq29dgZcHxL6Qej5uGFuU
XOwleZAsBsDImr0gFwUYRr6wMvUiXPod9OjMuClSSyq1B5sH+TqX0YnBMbO7XZaK/XGNQ+sDi+sV
Fs2amL4h6FK9H9fdUFeTk9Qxh+/BS7vYPqL9Ya7BvhjrIHX9ErKi0umNBBK+LSrhy8HiPVOcHjSh
Nm5BxlGCpi3bQ9oaioVMN5peRn9WJ8jBBZFKYDrsn5LhVshVPIpGZAJhJh9IBB0LzRghoybJxn87
0lPI/adnlx9veD98y78NoWmaIyz0hNBSBkNdclAhDs2qzGan1CUUqrHdJHe0+t75ALAhbuYCrwrk
RJm+0yUz5+d24YuzEqRQ9ySW1v++B9d5Z8/IN0JcRPDoOgyt1nsitJrZnRQq7ovnXwMyYPEuZm3k
A4I0KKVCBJxmqmdCUeRq7LpDsQ6BxohYJ2Oyqw0l6j2nPIs0/AJWPJFen0Aavf82HU5AJPY017JK
WIYizLP2lOOSisZ+CBajUdaVjpu9fdayOJQUCxaO67al4b+SvIsW/YZg+wdGl4uGQcwIQlRiPCwu
qVgy0t9LtehY78KCmqaKd6PGZLeSbVD1j0cZ6DJ1ezi6Nm6UNcZfHAaT6/yYyAEYy5XClVCYNN38
MaucwBLTkrrVf5ROBVcw08OaDS16dyvPPltDmYY51VDofxvDMhlW0yHFsEz690M52TMEZc3toE+r
o2/rZNO8GiGwSLU1eefK4xajz0tnVD1MylUuMvJ+LS8hXgN9MhBl/NA2H6+4NQazEMRKA7c71vz8
h3Y0wROJ7Gp32c4oJk/l4UQVwFT09DDXYwmdiq06GundEnfwvloruhsts8QmLGVYfittUQgB38wO
BLrqQ/f9MLp0UQOMiNRslZn6/GSlA3PO/GK1fppQyNvt4/26XbRW9vszydpKoOvm0P+ce9k+NcIH
WwI840D7hWd2dLpppfewYFWtQznkdcYYdz9cbiXTE+javU+ReM8vTLXwtbY74vgXqhbP/YTpPSgC
GEG0LdTbJWdt0eVX/zT3oHh0DQ1v9ONEOIxqFeksWPm7jZHYvLHvyoc/fcrBLKMzscNWx16ReEPu
B8JOoDW+5xamX1qHqsLsoQ+S/k+N84UrDPmUMRapfCXfS4/y6E3zudjUYGIViPbmUw8AfzpO7JKz
jyWbtT2rFieCPQeuS8z1xR3HyKNC5nL9vwa+lOunoEXxA0SesHdM/9VXLsBjPCOg+zvd0Vf294oM
nPjJy3J8/Ud9JXR/dHx2kh1GEDOqoXrmnQo2snS56tt7sVZquM/X6OKMN92JuWzmODglx/7FAd+G
ZmbuQFWoWoMv/VOWvUr2egxwgKwkb8Hw0AraRoEFrA3SpzsvmQoaEuhwpikziciDMJ0SNl9PMF/O
GF9r/fehqWVZijHVmgVZSnUY7IhHHCyKb+iPcYJvFW6eRk+82BFPTP6oJcJh7eBYURp6TdEc9CL0
yxMhwuB+CRFSRT74yezzAyAG7DaXFuTqf1MpWW40nzOoQvrNZpznYcFE2g3HFOiOm3Q7mtveSRWf
aeE6WjAnfWgL83BjKPEvqcmRhuVm5qHsPYigLAANf0jgmUq8q4+RYPwSDKKipRhN/lFqJy0HJ0Rg
02A1ympW56liVvT/8cakAXvmI5BQLX6zE63SkV3l9i3w11on2fARr2Atu3IW0ZtqTzX97+Wns1Dp
zTVQe+7sjDnKK2qr//QvrRFuUkjPBx0dmJF3huwTguGGQ/ceS6ZPts5vZgBTd9iWePTlRIoTa1xr
lsBMlLCn2BDVVOm0o1MQVdrkZ0TsxhQbiOXVJw6JP9bq3gNbuyi/1Ulcpl+V/Z2b96sevOp+SfUg
FgT+FUQ+8eSmcMkjQiguFy9OcTy+g+wqbCOafVwo4AqmclHDlh42AmUk3ao/pdgDJMXsGBZXg4p1
V2r+v0IjOjugOWGNgpGtMhhQEyxh4couA6/bddXHDRtEr3TP5i14dbm94LKEhXmyM9emHuf9lDOt
FXbLVoJnMF4aWzy3YNNCJ5eS2s57M2XUcy2KlUoQZfVsAoWhDMv5iwz1U+Ln8ol0ZwjX2vkpA8Em
RsA5gIuHsb5GYmDa0xckDPXhminQJUC363pBOAaAaiGHTg9FwRaklD9HoSSUTtsmuaq+s6jyH8t3
0d/A3w3IIv4hm7fl1ZlEnrJW43G2hoLrjknKmG7NsgUw/+5wU5vRYba6CmuqWkK2VXO9YiUeRj4L
byOV1O/8b640MhjPmxZhVjEEIjVlKtBMdmsQ0ArcG4t5jc+SKl5swtZ2cXepefo3A8++KnIBHtEF
8TfUYcAMdhddA0TKSfbKKG96T8yK7BiBX/WeInUYHxX315tPyzqGd3fn/I9gPhVnJTqjTkxp/XhT
tbvxSo0318iTJ6NqnFIz12uwi/bo7pPplHo5Dgtabh/m3myrogGUqs9NqRu0LvuFRvz94BO2eKCj
Vp3Ov8zSissU7vkzLPNEuLckThZm72rJ3HJ5hMX+GMp664phnTJ/I//RIcdMzB/N6tcgb8op10y4
5W/y1swDIx25KH5UapPMCUJmi66UxoCObNzaDCVsCEDkFV0ShEI+X94T+TPjU52TEPeMBfVlKAAJ
2pgPCICte4ujsxKHShjRRI4xOuKg+uOd5wSdHRQXdrTRdjiS/KoLXTJJruQoIOTm9BOvpaSf3l1+
DtjbB/tmiQUz5J8N5dqMsY92yUUgpR21kdWKdyrTgIa2ig5L+kOjXg8zeDyxc6QJ36gUG4yx+pEU
oMd+XzbPX4us6SOqs87PhyJnN2BXE1qAJxEeQL48czHbw/SE2vHJeYwV3JNMxkXO/G0O/KG6tGUw
z5WpQXJPmsZakQkGiCDfzQQyoBl6Tl8r4A78g2wwwx6YJQT+qSwkeC0Fc+/prMkHmTzibvvlNbHF
qLgHkqhDwz0U+YkIbsK2qJSF069TkASCrpDONOZxqCqFkVfaLVx9zRE8jEbi3Aco3G789YiNXXA2
WdmNLudsL9g/M1xQx/eEJKjK1oIR7J2c6h6Y8IGuj/BnOJgiAKQSjLo8I4yC1lB3TiYLD8JooQKX
dYtsTLHNvouHkgVhIZst5WTydyahGPOMKVWw3pTmSbXGLy3WxmAokyMJpkh2YOeaE1mN+D7PONpn
EjjKth1EJ1qGlRsV50VDqrNXTGjVeqWVH7XSQMm0/Ef3zvHWUyvOYkt3qch17TlpZfGkuNld6uPs
Wa6wM6YpiVc2v1Pu+8QpqJhQaiZPw3rXtND9mgz5TYT/80hxOy48k4bcYCom4KUQbegiNC2L7in2
zoNw5Q21RM/Fn2tQ+VItU2IdRnDWLN5ztLll0v6KbeNMED+nqyX9KjykTTm7iOBrNuePdVXlQHES
md4WQtva74qwTphJvHw5AUS8xtTdqkSp6Xds6ZnIDZB+IwcNN5W3P/toSlXcgBkcMf92Hyh6hI8V
9an09+e5Fb7q6kAE89yQXt/mvMSDhlKStFMNwkKtRvq0Soj0JOXjSQicE+6iazdknFsg5WVjBcEA
ZdqacgHwm1pz8qL3GS7tEyY8UNfIyLXBt4zrfsHP0bvPp8tvlRh8K7HnG0uyIt7NX02xESwTFFuG
5BxSmCl06e6B3YGTDM/+voJJJWuKwJJ/T+inAcCrAkBokMB8gL1Q1uwIPaqi/AmBZue2/7WnftwA
gK4kPOhyQdi/RZ/h3MiWS/6hoHvW2iUz47Qu7FrApqO7K4GWTGYAgYHJOoOGsb+QGDPC5XsfRWTx
e5aVBXT90gRgKHWLO0GH9coq4qUeqULJorVny16oyFRApjtDQPdI+PWvrtN65qnOFYbRVYNqdYiZ
jKmSztaphI5mcK5xP+926Zzq5SBPpSyAtouRkM62u9isNbX30gtin316X5vc+TvIOiwlNO9Z/KM9
8H711D2klOTFN1nFNaVC4Nz20XVi/3cNPDZqym/We1ZwuM36zuH06Ht+VhU003xCCF6k38KM93Eo
0cRhqKyJk1SFlYEy8TWZIha5cbJlxnOyh9H1a5my+vyUJqavzuFsW4dbtbFOM08QLLC4CRFGxam2
+PLq6DLnte8cn1ulhA9xmea3S5LkBU+NilL189w735BFdXb3UXvBjY/up+hJBv6aIhZ5N3jgydqz
WKI6GZehT3s1zQsgEzKVkaCPrc0tM3nqloBaIs8gFjqybWYfn/u3ItqLD+qWnL4U3Ja/xINh1f4R
Ci+VwD9SA+ZVBr95PP4ruD59mkNyUVxlg9hRdbiewO+CbVd30hUj6x/cQqClGTcJxwmUgC1P+8/b
n2d2Dx+S61u4FEfaAq0wQ/WC+N6ZjlH/takYq8u+NtbW0LatevQjLlGxC4F8H8ruqRbLLqdPUjmj
BNbHNa16+maiPBTzlTX3qw7OMKXOsNIFAkMncJ9rEhwmTUM+1dGD7Z3iKDUxajjPwTzd4Fow/7o3
MexgfZqkpSvjvw8SH7Y/nIoBn+PXKDj6pgp5ZgdyE/mtntHz8MeTh8vdgz933fS7XnY8xl2rh/Rl
jpiVA+pxVlq35inmKZNiZz3Fk2fd6i0ma1hrOB47jOQyNAIeH+gWor3iiaUusIJoINoF419eqqrf
l9W+4dokKOR7Q5oZ5gi0CYV7g0ErXDzZR8e9CXHnlSBrydil0we9L7t4uZT7IFh4Ve2kuYixwiaW
ChtX53QIV3RHCap9fAflW6zJlhFlv4HJWQ1duAqWkx+AgpYq6zP0+lbAq72lXR7uPHlOSI5Nc509
jJkZLabzDRZ4ZBCc+NhdR4VIaKRWDV60PW7UjusTSSc5wnEZp2xKEDn3FTUMU+KW5CMWm7fTopSu
8gDibKQSfvuYSN4Ogj/AD/3k6GOBRy6o3AFapf5ylQ5YO7zvgKO32W7uf11bkFaz1x15LciHNXk9
eV3ftxYt4ikRZDHgl9LKgPU23RjLIQIj/8l0p1RIn/cjYiFSz4V/0wtWZqmFw/2SMQtwWl6uNlgg
QcrVmG6k+m7VV49sdWU+DirkzVtWGKhOFqRtZlqS3yQlO5oY4c8qdcCGOKqJfkawtPH6TfmSbjHb
vxQeNQUvPDRSPUEwnPO9ZpG8m2Gmh0vWekdJbF4gIQaQ0GYcwMXE1igJAKS83n5kMWRCaqEgaqDD
kvTdALpnW2HXDWg+9JYTIH5aDs7m1tpcpFtOGQhhyQFdJejAoIrhzljOLtGBaYG0ctzz6BVxDa2Y
CqMpV84CSwMcaTs/X/BWbObRPBWJ37WCyzZuM3IVwo1I6hGWWsJhPc0Thlsi8rSIcUtncVRFLevt
H0NYCd+t3fyfAor1/1Y7ELkcjoZapPsy8NRNkHAAT5aNItRMHhbsi+Fbxlb2aNxT5WemudhUuIXJ
bXAxnH+TBuUOAFwxPfTJqo8+aCHVaNwVhwG9jGkcY1cm0ui3+kP1KY+a9Y6jZ8cGBPKV31UTpTVm
QUeZKfcBkKbzFYxK8Jo/8q8BHIlo9/GdO4EWQfEHrPIcPJflpwWG4ZmHUFZTGerilf3opFdH6rOS
BkXvQA7GFI744paybTPLzngXPI8u0z9gbFBuW6HGOU0XeNaGCS7qAgM3wyD05cUXoZUghffMGx8i
4nnvAQKloRs/VUkinW/MoMOaChKLCZZnvbkuA9JJG3XLos8bvOTzVYjgpdhshLuZzzciWpGEodf2
xguFr5OklmQLScIYDwUP/Fvwn+p9tYtLopN9TtxzIydN2seXzgr1dVFIlWmKwenlQ9iGaDWnI3uV
f3nCRTB+qWhQ89uhYRExUlWkiJmi4ayRieRHMrlIhp29tdO4vvnUcI4o9c2UnGwHp6ROVJwqrsmg
mvKACmfVn354yXiQDUiiAiJOowPRZuX8/szaeN+kdO9Ajg/MpAQrLns/+9W1laViukhLqji6hwUc
+LHOwb/ldxJJV+L37kpXCAkS5NaAiPh48sr8iZG1oPK0Cpcfs3aK3X1YAwDpQ0x3STRe1TpOJ7Za
ObZnWbD4uSgcL8VDc2qX3TgL7QXWw/w83wzK+8Bt/ZYIDBt32iKGyGUMKArwUu1QjwpOyf0XHTeK
P70EdLQmrkUrYzHAMTx9K0LxBnJDA8o0VOqQJTMcqLg7pYjnI4hA3jVR+bySB/ao+5UU9okQCi/I
QvQ0QB7JP2pNRGQ+nbL4cBXv9hfEovxiCib8XhTsDL+qn1J8802NrZAM5wTL6NeFrKyvSFWyMbHv
LEM0Z8g0D1tfmZSoRn5PBNfSMj3jYgbg3s4rg6G2XOoPkNYfNSJlAd6Gls8StT1qpHgvykAoUtuD
hRH3Z6YU7YOwzZXBJ/u6BGoxhXK1PPirzoHFPBzxKBnhbqZrBcYymubjXVKkZuQXASTanFK/BHvv
P/ERqxbrkGijquwbotCkm9orUDcVpnkVJYYXOLG8FiUAZ2AEiA1SqA07nHhCNLD+QA71BpYhpnYl
qnr/uEJoc9dE+aoXnVN4OCHGmhy0HsoPGE9pgzEYk5ZrSCsfsN0rilQcUic/dUjnd+PQ5G7Yhxq3
YypDOsqddI4coR5yrio/gbGq+6HyQfdOgyc9QeYIkyQfh6SWJSTSMQXQItJ2Odbe0i62i/dgGNcI
tABAhV3PgM1T6da++A4YAaxlT5I874dElP2q1AxyE7Cdx2uOW3CKGWa69R8tbd2tQoHjKTBZFBpb
K/p2xiuXNYujF9SXwMSKfCLSKrgWFHFGvudsLq1SW3s18nz+tVdgVf+TYC73sS3LIn0S0RxEgo0L
xmUMTKPijuxzrFoZ/zuVuKu8uzumn7ZsfabS45RxdKAC4Ynpf9zCeGylCQUubrxi3EN/Y4irr1bF
VUo6mPljqoqEX3WQgJo0jWTNQk1t95CR0vL84/hqTw8BpACJUfF4/r26017EsImTpSy/RTv2uTjM
zVJ8f/hYsDw+GiYroUTHe28Nfgb/TC8dkXzl5ty0WTXUQgwlXnozjBtQZgsliQOq3MJA6ybUPyuV
X0mP9ohYxAaD/4sCvoxmTYP/h5N+tGhd1o+8IsZYX+++1KxXyXJdnBns5HWjmOKqGlZIMWN/7Gy5
MvXhS5zJmElW0LVP8iTenzL5cMZ1ULSETyvI8aLZmv4kKbRhiGoxgISwpD7H9z6HUggLFcGcy7qR
tunJjtMAAoc/CHlDsxhpsaFyJG4lP7JeRAjz8A3KC7MNifIZ+ZdU+nlQLj7egMWF3rK+42q5P/O+
z5ek+gwjajfyca2MRUI4enrUoxZOJwOIiR+cnYL+cjt0cswKfQbl41Unt3d3HfHP+eZ95lv+jvmW
ZsdPsti/pCwGlLT9PTzlcBVkdElxhbSb5Id31mXfpIrWs/McHOw1ZrsgXnXn1Llg82Z9pA6JQviz
tNvsWT5fs1Oa4IaHhUMUgUMTqzIIvzaOWn1bQlHMQriSfXsrfLC2eaKcyc0OzTnC2iVqumpY+Rpw
7uVWDoDUvYwaE6igg+xE4anhAUSVjyaIIQd1KTOOUoJ1Zgwh5431WjPrvrCQRfmvQ2rlR5L3+u5Z
MKe8gfWOz2Ht3xcBdEx4v537y0sjTCFSQXc/brkj+BnqZxKUy7TnejoVDYr4/POuH1Gf7bNLxk78
CKmuINCeKhqrQtfi+KYNd/+fzgkACnnfbWnsiOxRmBc2d0uNaCwYNBuv1W7aY0uG3zRstoFc3O/G
uD/64A1eU/jrDHNa1W7J7e6rkmyP4M8icaxRrxvVyBafcDUuXKkpez1cWZilF+dyHtdFwhUsX9ap
nbnxtyeKtTvE2VbkADAykMLZLIvfzdOC2qNmjmVs+mGFlxhyPbR+YzzXGoV+8UNuzlI1y4gSkdWt
mzi4OwhI2dudD1/7xf4PpsX/xkc5tcrdTDQZwlUQON6J4kQmoR3lQX6Y6FqgWk2+IBWIkybQrZC/
SN/ub1OBaMDbF5eWyLXEY1L1p2geCfL1xWzRCt/oChk89WSUyyYwB+kx+gzy5BCujuIqUgpjg7a2
kOITr5Kn2g0xYh+m6wOflmU+yFB9ohq2JXriDOU9NDhTzqFQEBCN8fSTLr5EfGGzYO42wOjrzDXf
NanjL8F5p/s3J+gO2jf3dqWc6d/OAvCHMOkIggEq7IEcW0/FJpu6ATo/c3nCi4J9OARf/+gtCbgi
VbYysd4U1sDDotkZRWgKdvDlDmbZLCM0zKzoNAm7+G9+B1xxxNMmHxh1X4vnSdE8JvrVMavhYpJo
FS28sc9WHFTtGgr50aGs3Rq/4F04aIPzF9ypQi8dovaifUBUIV+buJTfqILHE5AUje5h8mEY3erd
lrPu7ftLfgx1sc6OSzkHIU4XrOiV1d2lhj62d+J5t8Jp5oEw3YooBI+DfTraXEHSz3Yzwn5d9piR
1ahwtJsnmNgDYtUG0lC5dLWFMW/9CiUShNsm8x3YmE4XUR8Szd8Kz+xfQptj6Ehmv6PuedivLvy4
SDXu5EfEooPxlVu8ztNxHMzfVj8CQhyFkBN4O+KEhQZ/Pm3jGrCp7P+U+fRfyibow9l1n1fxvyce
kl9OQ3kJEoFot5UfxNJGI7lY5/sf2jdkt7G8gtRkFLbDahs/7i1uFhbYysHRwOaomo1bDhazokaK
b0QfDWVCqSW7SNkAdI+3vVXqhM9nvxBgZYuY1ia+r8RVXkHbJadioUy01PWKoUCu+IK9ohnhLX7o
xZ1nIhm+4QLoTRix0O1KYiXGIbFI5g5anauec6/JkyRHAXn+fHp6LlcF5lv8HFbN4+DdkAfNTE/8
EzP4VGBvwxwvi0oBKwB+tebIivNb21Iwqw6JiwCVUIvsvm36U9wfT9CgwosJCXZt8VDgcoPyrjvH
c910bKu32BTmnOZ+9S9/UUexw7S0fcvoku8QHURySEGUhSIRF6sgA/ZbAb0gd0wRYc5MIXa5kH+c
8/RmE477XrRMG9lT5on7Qd6m6OPi6gDl2Bdj3ZvIc32voKPofDaGd9KxZ+Z1ekIqAx9gS4Tm9w5x
Uf859MCdBR61tqEcAEowWuM2GI+GvJl87XwKdGNKIDnr85QLwxmWBZfUhvuH6POGlWyjpyQZ2sBK
lIBVMLUYngtb6MHkJ9O3dEoB1bi2EdBB13TvF98pGLKd7YsLo+Jsly5CZq1n05jlVZ8c0jbx7O9E
quOESlbi0sbsPwulX+hsPYpMgDbQwMTRp2rLzVBJGMcdShADx9qqHNiK5pGfY2UfZfoeMNo0EtzG
VlSJdLlNLZk6wTzTuvxn8ibGUxDpe3l44REc6aIw5E0PEkULr28l+fBOCM3f9PW0N2eNv4Ufljhu
2MM4vBXh0340LjLlA97Ch3Zva0UlHy622OZAU9ADFKe2dewBlVXRnuZZ2/CmQrpg4l3U3pqy4ivS
hCdg+eGCu4lDnlmyaIgciupqiMzIwHl3BVzBrInxiYno4/PKZyhEyqN0ed9f8ZThvzbOure6xlFE
yluTPl+mSuWIbdIOBudJQDNKhTBRtUI8RqfZQkw2oBkxejubqzX3mU96EaHAomtdsXF5rcmgVtk7
SprSdh7S591wgO3dujzAIqtvDpD2IP4126gZGjjsFMJx9a3gORVWK5gsCPQCOi81+W3uTv0O2aY0
UjY1g1uO4p2vDcrTYWIFeCg7OLT96CIjcEyKeIElq4bn4vrp+R22u4iNeh6oRKrrIUPc7XHlyntX
TBDZzZ85R+/M0cPHcDNfI7hKAKTTqoJe3ZOWeKUnJhXeRC9KzqJ/MLSzRNbaPsZ6ioUa/uJ3HzTe
T7kXrUUGWqK2n+N5SQ7R8WIMHAOmlcSMKWG/Du5ggnbreAOyY7WP0+Lrjb+Nluhs9yj9cSN57byr
bQ2doN4TdtpKwkp8Gloq9t4x+gmZaEpYowX1YY2fcDJSiF2vRT9eoERp8WqaxREX0/0UZVuiXZyo
UfFjIqmuQVGImPKlLiQ7YxSZfVBiQkEwoD0GM2itGEYqEbAOP3VnOz1CpyUNBZd0oj30yFISNDpK
nGfrTxJUIt7/WInU18+fskJdzlxvZCko4T8BJ4z7AAuzgI75TCOUHj3Wf7uu8wpVpMLbCSo5R6l/
KThQ3oipWR+00gFAM/JNZ7aV8fSPaPUvFPr1EhuHfsjWSrR1UeXTJ6Xo7GH54/TSbbGa8wCLPYWd
VwZJzPWlAthA9Wj5c+UHFUat3LpuxKVR9RX5xp0C5RGw/eL15x1QjdUkXmIsztrMyGFGyNB9XXZP
XlPyrLjjiikCdK4i1Gv0xKwtqwUw+wWvFHogvrhEZBRWm4Pl/x1s1cA9Ft/e7NkMXV29d9DO/4yF
W2NGNzD/a6yQUh6yKfJyvc4rPWCXMfZig8plSVWt/fWPPZAK1ZkXwyDR2kVUIV0+yD9opdqhydGH
zlgsM/QSKBSMI/0R9e3cRl3Gj4CysIbZnmmHCJcLCVfklXf93rNxTM0u/OnaAI9G19M/t3Lp1E8e
JDp5xMO+eGi7MiCpk6P0QpTz7WYL2MSBzt8jphmbQIoE4oYZi7239BsEoGn1TZCvW/dz07coMNYj
Ut4kq2VyMWfsljTTOMvEAMsbwOTXuuV/i6R9Ub8IDjNb6j/cOHeNUoca+nbBX18woYYvjZWLTcHI
/ejh/0/Iq95eQNbWEtlSD9fyMfJg03GIg5tL2Kt/iGRvtt58cpjyodYvNERqSH6DEsoQ9pS3kI1Z
zhSmmK4/VUpEB0VFf9resbXLNgqxNZ1k6BlLMAjemrpU3PKker4JIsOYTsQZcFlTeodNc0e6/zT/
lT6ZkEc5u1rPvD4dOG1ZipK0qQy5sqQ0ZdyaHSIGRnLPEJvM+qLJ6JI1UWBvHcuQoUOf0+Yg6yF8
HOL9uR16i2pITnSh4h/Gpq/yM+2+Ge/N3tl/AfDxtbrKKAxfNBWGj9+EFMwO62IrhoClZY8qChTO
/qeqiUb4QaKLkwA/2UTekfnbhjzcdW1N61UrDqLflprsPPbyhU7/DagBmTrYQZ/78NbVyisEEq/7
20ginC26Kk8Zq2PZ/sP2Fg77MWlaISTxPAojaaFia+QfJx36BirlgtTh/XdkigbvRodrbb7WCiZv
396UNeozFlshx1Otb0+Vxf3efqbAshgF0kdbBHIsEwIvzpOKgxGx+/+flzr6+nBhYfcuRcJ+74me
i04eKgI/HveM4gyv0Jb2OnuJbyNrufamcH+A0AjP/NlOnkhiyXN889JfbIOCOxdLV6AeTlfp5vV5
jdZMRNWWxt6BtrM4CrGPWma5TzzH4tNEaMqmr1BzheACkmu6IdjxAccJzKKfx7i/BM20Cws4ILFg
rFFJm6gRW2iyRX143CT7Xv+hXKy4i0H8yRIwkUEQUMhZqFmhwj4XKLwwpeHDRb/7GEBy1ux5P5xx
EQqrRQ8rBmuDu/ad2O4ivcfXTTJxs+HZ3/nULBV3MF9O/fRFLgUC6JxNMxBWx+R5tvgAzM2OBwMC
fmTbrJsW6PGT/sI5w7+iv117fUw4dWeqOLH/MfIb05HCmb0H8GoTw6zjVnlLv3+d0K+Jf1atRNrv
+Jl4PUQrR0eNHLDKdLKBWMpFaduWGu+NrRPh6cmCq2wf0yWBZiohkNVl9qoGOqlNzG1Lea9+R7OR
1vBNvS5SE6Xvcq9afFMANjjmj731gKXcyntzQMPIr01nIZYSpWqc1myYTGZKdrdiQL0FR5ToG11J
ELGDEp275GMwip5CPlQaFasMgLFF8T2Bq1OKujzCyM/jCHxOeml62m5vUL7aVwnQchEQKuCfj4mC
RW7IqVLZcQHbEVG670x/AQn9RreVtT3PlmvNsK+sHa54IeRvxt069jy03STkyc280QAsaQhnVt3I
9OCipxhXB1m1x9C7vS9TIjvlLsBytjByb5JfuvfLePyAmuoWD+A+CDHpxpt9GCb7HWIdPley7eKR
VZDsCB8bvMFUic9Ii+lGCSnGWrFywOmJMmL2H1dcG6fg6ToD8ibViK79aWn6tL7TgzgZOA545EV+
5H6h0UexDcDX/iLgPDnmip67/D5xAqFivtbmYXSbC8bczaqMr2xJ9V949cwA0EOtr7K6IeS0MsbF
Sj3SEh0JTZXRp+/AdX7hFEPqUtj9WbFImDB+8KJD7GaLYxab0DnSoJuoDpcx89tqqZDoZpHvKO31
SuCeLUmd9JNLRy3wy1kgtOivD6BSlG9xZnjeeKV5og4aQYShaS0BviM2xvR0TRGeieqz/RlKGrRC
J3+C0KYymBAUXvL8TVPd3WQoPcanToUR/PtaRAxJ8WigaA2zRrSPFyK8YIfhVqI3vojTFxJj2OlS
3zx7WVjkvoyZUmz2DZPw4IuvtP3DjxQUc1k8ty2gGOrZxZJ/lgodnEqKSWu07yLeKnbv1MXjZWXr
DWt/b+xQBKSdx26ulSG80wLwlS8i/BMf2k0Z8Gj4L/Whs/Wn+zqdQHXrPQuNSiJ495gXFj6/J619
Ad5RWRk45lFWxqHUWC8j3vkigHbYUJRkJItbsr+uBA0+mAbLp3fTopLjv5ejb5xpP7b+t0CBvAGz
T1BwNw/LhqM3+/ZhFl0lM5YFa6W62OdUlKcR1pPcSwGWoZJnWxQFXkLVXZHIjT5FIXv6HeNF8oZZ
wqn2GfAyBQtwddB0y4+EOHbA3ZQuE6kt2SQ3bn6JGeWfisFyd/vHEy9+SM5qUt7FNUZzXxXWHXuX
1elYDPKVuVwAYTFqIZcxcDGJw9w9vasNL1xKi4FVJ48CDRChfwkYtljz76exg593bTJoVPA8npYQ
K0kuNmpYtC6V6hJ4M98lsjN8srPuubEs16395zLLxbMWoGuYpDV0iYIYL9/KRGYIobBu3+5x96in
OijQrvWytNquIXbDDjieABtSWMCCYtOMFE3wo4z2cPaEAag1KnUmdAkd3Uwr4D2VUkhofYNKx3j6
rjMR22iqMtLupFj0k3j2gPJFUVyUeVYfsKXu2JCV0Mg9z+j/HjH0P99qytPc+eHLVIyg6F/vORNB
9VrKJ2o1clOERjz37o49Jr3N3qFQIKYZjjZkwGkmNdU0AJKsJptRhNscVN9v2PmlImw3kgFZ4VoU
f4tAwYa1CEHq2wzrtEMwoBsDXJNGCydV36v9BSo+jlBCtY9fH3GgUwWEvytGnfZ5cYxioYaYnXgV
G6V3Jaz8+USlABSp4p4f0mFax5wX4MU3Ww/2tyULlBIg7UjBpFKuDcTBxDdvih0JcP8sR/Tow43h
0qxaj6abnGdPF81F1UUraA4iTOMoYU4xmIehHXMTx2oVldRyskp0wXRRcPS6e1LDrI4/WDN2+wqu
KJqbrg1yCiOqIp6WXusUQ2EkVP9VqGOw95sinaVO/rn+2G9zzBVaVTjG78P8C45kyJ3s1Sp8p9wZ
NOicN6WvmJ7xlvuLcmgrCVFIZLQCESLolVpj4hwt0dvmuR+J/R5ZV/7yYE21ZjXFQnAL9/FpCjoH
HPt2DWqmh0uMeH8AJXcrU77GKchCZ/tw3ZFo+xFtTfIuLkWBLgxVpsLc4U+uo3l1QQpk8zLubdd6
sWqPvwED4g7z9LzujPzFYxdYEEm16c4seFnKpK3LfCmrMr9Of+8fxzhbjShxS6TYJ6ajRGa4sKIg
O9MTr8JUX+vu3UhRrwgJdGVX9KWIa2hSr8ptTgCxjdYMvEsRyy3DMBIboF/vtY00lz5QL3u8CJzB
XQbIFpIJBnLUgSwSdbqLqvxAFzkI+ZlJdtNw2vL1GFMm5619WtP3c2pXz9VNduguLBrzA0xyiiOG
qePEIgKcMk9w2KV/vkap0LV0ECVqOwzg238aHgRfdsf9se6jqMOcu1o1r5ChLd8rxsVRqcNN9/FU
N/+VM85C+I7AzZsNTcZxtAZZJadlQFPgWlhhYCGaN02l41bkuBqZOZL1H4kSu6i29i7xvL7FdD1g
LPxfQ5hvdoRlYUbu89GGU1HPVkHsy0m21qDb3vKOIL0l1Qwd6ppR4xWgD8TSXQ8rhxorIJPAV/Zj
xPsq6lsf4TpNKqpaLnxoKio06l9watbOYPkeMgT4v8FEjww8bhviUHXGAHIdKQ8Ij7N644aQpxII
A8KkbU+Lq8k3zpY4aNNKOMT9rcmPWgo3c402JhDzPAtJd8vPRijeUGB/ow2/RgOCZC1w4ixy11os
u/dbGnCeYvKGd9l388VX79lp5eg2Kvfg7/XFPgTXxWqLfMyfiQbA7V6P8oOAqz7jjjH7EvLvdajv
qstD8AePQeAPLwaFmgOpPbJGpM/OBK8KPAJ0HzMYXAPLmLU2S/oxeRCshtzX3ynCBvGesI9JUSHj
iJh2Z2jHYCgbBcRkY1qWZBdeZQ/WlyD5Y4VEtJEbf4YmrqqZtNC/M9Pyet5CYXSunz0g8qrIa9sv
/WYFbt1pD+HHjNmUGc0unwKmj/DAfkzCwCi8P3WEJ3bNcslUDL2zT06e64kGWzTkQqQrzHL1GZVh
qGYI5kCQrIxKih1IeWMBoke2ONzh5lfHmLOa/dwXTyB5NAPEUKohCZjIbO6pyjLp5hlXE5ShW/Mu
8onEMuHZtA/wA38dNfn1U/dqCsbhQfm7eeDKsZqPRs/IJ0MKowxWxtLOmtUrapKeyBMjD0xcqyYU
7htNIWy6sNz5eOGSG7pP0xG59RR15TMitFuU8qjs87Euq9y5uTqHPRfvBFrJRfh5Ez5v1CuzHraw
mhRqONLwBkbFPdOixo6FBSfPmJxZZNdyC7zWc+swCR450Rcru2+gWYS70mw6pHUnmOI1oVBkR0Vd
cEp5OOXRDVJ/uyGtkRZeF/C4xc68MmcTE5n+aCuLEtqQoQ2FOasHFDqVqV4++cE6bDxh/XnRt1ow
RIrLUtfsRXLZk69QCXBqtlwDzNTi0F153ojMNyUhSc826Gi9pNgGe7WXg5ejatxPwQDCQ8O3qdiW
bIMqwltLtjp2zkWFA/6/9Y2D6ryOuLySJEUcVWgGKo7iNuMrA1a7ImXB/bpPxZq4SqfSq8qM/Ioa
dTjgJ4mubweQiWcQWyUmBwJU37q5eyzJFLntUEBI2C4StUoNhnizFDyLAyKXyax2iTG69UDIAnzG
YPg0cks/0rts/e/1FyzR0g0Vy2WsNs6NGy31c0bC942snd7tUEVykULto4UCCNC1nEe+qgHrkDuz
NoPc2bNcHXx4Y50d/4EV7o5k56XDRe25P9wJUxoPrIkcLE/SE3AtQdI4oxyXwmZm9HI4Sg21/wz+
7trcqaDdLyxiAFBrmycwAjj1WxOsOUhTc/qX/xKG4ZgjW9wGgXiKgxyH11GS6TI+tpVCLQNffkmB
DfmlCOdsifW2f21Hx7VCil58oZxGCe22zxGpJ7P/c6hr60o5latBUw3VLQ/6ywNbKp13frTQs/WJ
rvUbPcW4iDgYr4Jd6c8VmPOG3nAPeXE0ulHOhIsslBeyg2EnFJceKINFbk3rLvMEH2s4HmPvFa0X
PjV14W9WmdYah9mNvlHlVw+K4Mxqqau2c15yZlLmXsVXW2IeRlWZSVBKFlo3w2JvZccn4bhp7Ran
lDT3UhNa4vxCybpBkSXVav3chBX8mbGT7g+k3pfGwuQFGthqoRaNkk+68QwiZkhdSXZTsEBpR5Wd
x8VNuWPXd+MWMVmVVemWCgjyPkcI7rgBXKO8cqCHYEFGc8TLcsiYiuBZ+YbPNgE7aDAJvSddtZBy
LyAi5msOCClrCWaSWsopRIBxMMs835jB86tlOeek4frAEAWG0cpaTnR1YT8XEZq5qbxkK3k8t8+U
4CdAZotMMkTn1v6R74x3UzA3oB8Vv0dr38lnUSNG+AN8p2WpfprrjGArv461gixALrBvS+PaV/Oy
/DmHSuPJSCo5H7XnyXRTagUfNH3IXbaQGZR/h0x6XIEEB/wtvfSDs9K9de/n+TQ9Iuchp67JFXB8
UWGI2iZVaclBUoQJ5PKbwvErCLZwhBZka9P4R4cLyOSwqYjS6tFTV7bgppQ4S9yavotf8yIECo7Q
0lhTl3v0tlzFbpWMskPMiRkzJmfILHM0JuQ5Jnlh2c96m9i00oe9SBdmnHy4t+/ChPoKW9Pspe84
cPHhWM87nLUf0TrYMfxl6IiPTHHZpnJgdeXqnVwQkLvc/kaxWXCVReLXnqjUfqSKJ8JVL5+KcD++
Q4KH2FK8L8d3IFq+e5Je32kdizkzmtSXWgAlQWzm1HG7cw0CzULhg6LcJt5Y/lqr41B0LiQqJBKM
LIECbYxJI5S5A5ei+B2HixvS/fnLhb2+gapmRu7TwPS3/d4tdGyaiCeBCmbKGJs8SZvF3cBa82hM
7yABDIj+l/qdWj/vmJ9qH6OUTKORnYRVeQxp/3VVEL5TV5dkp+sl1lCQhVWNv2fvN1Ifpg1caXK5
uJaKxSNeI3TnxAv5IUdGd13qR1BhuyCHRbTp6WAfIrTn9MUUddnMPIbh8fAdhkyF+eOeVItYIF6Z
xzLafyrkal8YsdRhE5GqTyDevlncqqcpf/SL6K2cHx2gdyus/ck2liRV9ZVcOBQRy53Zn49LFMbg
M0m9qAMfunFdN7NWmiRC4EJpSBpcJrQ+q2Rg2pCP4xhaQ+kklMPZt6wxFRHR8gXqbA3kANY6cg9U
bmOma33qCgcBuuhNEBt/bCzEw4sJqJgo6JGlT7Vrr1wdebXI20dxLm0RjHkn1N0W1ZG3+abuxVcG
31T86khs0vsl2GNhC/wNdJoQ8DVahMhmag0mzKY4Wh0icfXTi8VJctZ3ajnJB54M3P3fT+4aMXqa
EaAPK9nOPDVOAnAdlk6FybGAjPPBPuwIvtWeRBR96+a8nticu7mRvwloDwdL9zrzv711ecT1TasH
I4qTTALZWV/hNSpiwEOMhJvW0uArfvs2OUfm4YDA8L5u1kGbAS8bTYU1rFeSWQXhEJULLvS+l5WR
sPEm51DHW9upg5SQsufsI6Nb8PmLycHx2W7YhydAx+OSKJk8wnZRSU1VTGlOiFTGHZoiDfi/YK/l
eTQleHa5HsWPhNHgsFFSPnpD8nIMvAf4fX9+wtrTW9SjT3ehd2hO4g/TRGutKjChCVWVV1S/Bf+k
LLi86546p6aSVw9a/SEnnp+19y2rCh926w2FugO64Ru9CucSX+JQ8Htt8/NMcoMrooi+b7WKzQKN
3QI29AmLHHK6Denks85HTRgNczp85xHjjguQX2F2au4PaagQ8QHJzcApMt3PLW5RLoLXq2rsNRcY
cVaA8VIbZ9dJ/h4sMm5we10Jv+cHqeY180hgM1ysPizfLo7UPyrszSOVVr6Rsw0Jzu/JJNEotrFF
OTu6uZIN7TqmGYQ/hOwGSOD91+5MSg2uVClsQUpKrUwCT6EPM4lfjZc8+qJj9np82WFchJjCZWD5
N1XCA7bX0hR0vFGAkGeXBWAt9dwHa4d+s62GNx4ygRTWhSIa9CTspoTmq7DICgscjuQFZi7vI+dK
2gKaTdtwLSYKpadOI7UCVSDt/zB/lFVKB828HnKRZ6M5Dnpyk44p8OLQmdnRMpt+s6zp+jc8wIql
jLJqXkdp+vlHQFxO937ZopEUeasqMXlMryAxR5Kd1VBweD5Q+NWT+/oRGeaZiqwgTVg4HYP7DZXO
7k45aEjPY5eFnj7HlBXOk6OpTONSkQG+Nyv/jw18XsykuEN2xQmBTY22Q8L8lZz2NDB5t9eIHBaY
cOLshj8e7+LQYG+wHNfZtXyCZQwsA1oTCBC5kMxA1shosa/nS4+niEO21nBfTIAzyhX0YkglGpTT
3yUyG6uwoL4EmRk0gMVzoBAA6Je58zz3HoOn1LJUHMuJzA1VQIQNVBa5TnmF9IVuo4Oh1HCLu4cJ
bB53a/CMB2i7FYmUKB8SOl2o8aSjTwEq2Agt/5uxJd3fBsXvphDFTOuHgaKTMhhEJBH9ZXyVkYOL
kIyTkWLkrDHqeWpiR3EDZ8WrPOIpvy1lndhRrh+7Mj9wudHlN4fGN1tQGOYt33ERzb7YxQy4wj7/
Udwa3pxf0NYy6kHND+ua4hbEXRRcyDQ2NvNhdTmORe1ee2ByVe7f/6ffGX/h00u9sJ10vW+famhp
8agDjd1RW6NPck68G3uDu/bIIRnjCdwi7btaWkhjAkungazDRVCBIJpaZQTBS5MizOmSewPguf8E
XwsbK9Fpv7icCFRWKmVPmYnZ7Po7I0HuDHcikRCsn7S5Sl1xcYNsJwHRnq1bjDdkgl5bcsW0iDjV
8TBequiCdS368ZiUdWTtJ7VM2YE+QUzG/ciVcFv8UsI9dXaI157YXmOWG+4naR/bIj3J8Odpu583
FvwFWKWjPfYcpoxVpcAwiEpCQBa4r0yjT+05DRmHPySW5hI2XMntNNg07yONEgUCysPSUTv81vuU
PpgneESp0gZZrLYraY6CIFj1igddxKKlL9PO/dOLc26shj7fFfYG3TjPX4LeAJP15/x30J+hDqkp
97A8maoVu+cD5LVR5SyumSyHubQmWOAp6Z+TvDH6fAPntJddn5pjS4JbT0/uPle0A7Hca9TSPzaQ
hr11WaqR7dsA/Ucr7ejiZ6Me5BXGYpNEaszfJqiu2MRJ6JOV1Q3R8dZbxpvHKhJunEiMfDhAOBPj
zfEM/WynR7WBunYhBHoBGIVLgGoNg9tV5EszK6pw8mHYaz931XGEsVdW4RvAXV8UVaT154LsNFtM
vRiv+dIl2DBHK9WbZ/zLTYhTJYWkB8vHj4kOIItQqfCOGmono70M15VKwZbdslsANQKt3BRpND5J
al8hUGQKw47ocf8EwJZjEqJCRkVJ/MmHHKvBaBQWkdxD/oXrUrm50deWQat3iQSftTv6RWeW2RfK
BjKmlslS2RHsoxj7QxbIS+tEVeg2jrfP/CnITGZhOQ3PN+SB1KH+jgffb0OpPGu+hYD7nDyYfBD3
OIgZ+d9uxk5GR0lNr7Nwa1TJnETRt4XRnKpwWxBjJbQsRzI6V+5pvKxyM00+DJWYhIUJYRXDn2x6
snSeb1ZVjmH9GXamI777n7raS56L7AHs6QAkr1ndpcgXYf2f/xm9RhiGwuIrjneVlMXoiL3kvX2X
VnRccdxeL/BAs5U5Kv0sG8ek6H9t/Kz6y1Ab3fUeTogF5ObBmiEUacyRFHH5je5iZaBSK8DLDEoH
wCDVcIrWOkPz5JY8KLN/FOiHsDhQZaFRbIlBSIQulc8BrJFTV+Px6fNZjIXP2le/ZVMNZl+po4zg
/dipF+R8anAUMghra7YKnogsSc7Rh6GdolbiekgBM2DdEb5X6/EpZR+5/vmK/7sLHXCteRF+3cjG
W00BDhOmiH3Y1C3JSjr3iKfOeuyppAjdfDjfFYzvvua1tgVcd4euE8hB0OQYbOEnJdrtA1ZeWito
Duwz/pO01hRBWxu6Nv1C9S9GOOeA+mFa/IwF2Iu/IUf2p8fdv1HMHoKyw7UoTg+5G0aKowXzFG/N
BNR357+Dn4f4wiAxxfa7gSBxPt4pCmv3BCKJFynrPanJUG8EnUaHVzp0EKRJMQ+uwgt8qYoiwhO1
MtMS1yJkkKcvVkt69fNYeYKDqx/3VAZuyA/D7BpnaAgNM8DRfRYRDo+XovUyzyIhZlpjscieFI5r
0gfnQnVOk3ZQm0Nl35HwpsbB2Ec7qgOVke2+JEerDc6VzkLzoJy5IMcRlUwOxYROyxD8HV4rrUif
XJoCK3yvb3st1r7aGyiPsMgq6WVorYslnXCELAW6IpcMn2ixAoJs79/68vkTpnZnaKWPjnti/c7p
Z5IDkULje6FRQBZFE/67euwCdrJjJrcb6oOuokKndv7FzNXpWJYNGIt6tWdYGB/Ea6DhHBs8/FaH
cnoxz7H+gaARZa2PiF/GCvpVBRLqJXdQuhGyOBBp+Mm3zmnJF1EEVua+AJFm2GjH++0a/ggMceuK
A8X/OqygdUH+W+yiph+fHHSJGmniY2xbOkGpYIFE5HwChOSxdlV1xH49Tqz4j+HBvaanl4wShHZ8
mBibQ1L1BxjOO0R4BVsN5Um8cLZfTzl4ZSeB7iC/uUkZl49f64cpCLrQEHaFztrPRsGCu2vkevcQ
6Q+Sfs1lXKCBZVYY5ZtQFpj3Xhhys2UiFnN6g1GaqdJTIKrQ1n11zIrBN9LChVCQv8axEFUU0qYS
qBx4WHoi7+Lkx2Ub5rjYbM0e80Wogcw31QW6xX655268SnZ5vzIL6p7Zt6E9jYgznCDYG8nucF5c
8Lv8+Jz5TZLjCufM49R1u9/yAFB/tzzGbI1f39khKH9XLI75U1tEjQ2+cel/xhBtdiW5GHjAliAv
03gibNkA2LlFzUbZE6QCMg+EwscJJRUrJY1MIibd9qq6DRjWxdiea5lN+CmGTBpnJuVTuQcVYtWt
lL1ncy6fV8Tnh7EZU857nB5denSCHQvzPTueGCp1WKRu9SbC+aH1glHNVuSG4NKiReFp6W8BUApM
rssvG2ckqjZ58S4aYubd7BePAFu/YdPi/zO3GJZmlARBfQHOhjSfSrVh8XLpKMKApqjjvSuPEUud
0Ca5m6JpZLrTGi+8s8vDIDz0di0HnM7g0Czdaxf1Odn+FdROy8FNy72Hv3Bvz4ofVCncXXWcF+Ya
R2JZZvGxVk0oiveuiw6zODhEgV8BRlDWdLnsz1VnHqx0MegfLEtj5Ahpy3pMgRjDkiqVvcK/Yy1h
mHqICnfDDTwHUIBE8xjm3xPn0Jh/6cId4Bxu3a6LPt+BfpOJ7uYqFRWml1kebaEaUFdy72Z7Ct9b
2o7emV/3oogoocjDDp8GZ7ffbVKU0orC/w0qjdAeUySLPOw/JjbwXD8V4rRWC9IqGAGYFHHwfH4a
xRWKmjfDQob3bqwMhA6lTFDaodsUiErtCMWhi43P87UiaaRpedGVOa8vKJ8SGID/GB92tTHEK71s
78j05B3+VWkG8ZaaEO8cKvUzlz45EWkeuWeUvsbgouJVmuiPtzW36vaSG1XkeTYqGKW1WXnynUJm
gB7O8FWStx3MxOJgqOvqXsYFjlNRPqCBcpUkPBHc0kb5k63r3cm86hok6AtK5cLscsEd73MBxY7f
usALr2P9CcgFp9CLgbXvuivnlWtQu8D0l8hjxXAYwI5LcrDhqEeDxmDL0+PgSggSsAGYm2B/ys58
ss67eO0AA3fOOPfDVZqovGoM4Lt5NirxZjT2T5345zcYbnX7QxumwzNjO6y4XA2YSJnZ/sj3wIlT
LjYXA5Q/37d717AWUuLbjbtfzVTe+t3ONjy0G887L/aq8QmPJrdvvash/9EIn/PmnmAN6GQEJZRR
1PJrGs0XrvzaaNZYnt/222WeVmK7Y4ZQTpJYAhdncjZWSt0e8U8cdUyYYlrM07VF4EzTNwAQ7B5e
LC//uZxfNHpTihHTANyi5yTkA4/Uv+q0/qcJo2HOau/dk0k2TXR1t/lJxLhP8mtB9RS2F4u6mVPT
zkypFV+t5oPahq6k5CTTAj2uuo1aAwmeKfF7lw4GQfmKoEcLbErUmUXvPwZkWGnX05j+wSVu5dGF
NADwIHBk9Ci8dlACslbEWbhdlVPuh4itIkkhC+g6El+0K/d9qXTyMbOgclshuZ5PlmdGvb5ZaRPy
9w1cbA+MsE1HX9C4uMPaB6wG0JBO69BKOWjVsjlpmiNj7Cyk3Drf82epMpnbpYN+QvwylS2hjHfS
I8lJsC0pAnplfdRnkaeVw5HPZTkBpOYvkQO1wxupqe7SX3AZqYEvMrtRJ2QlTYeoEnzMcQZgUewJ
9Uf5Uc3PWOlv/VXICyxo2Rd9IuXZlufYwEExmEcO48aGAtwopV70aQqPSZZlHX69+lSE6RE8sGZT
ERVq1YFPcrD1I4xS6RQwy+94YI6QpYInfsCdD87fekWwHnd31DAslnLHnAAuB9k1lbUqqRWFw+qz
5bWV5c8Q8injPXkSQHwG6Bk0FPCvy8Yr63woovGGIvtI+hBNwBEdjzZXVYLcrk9bbY/tnH/qEIm2
6uBqG6NjnNbxfXc5ER4rqv06tNXBuRZGgGzyfMUk8whlyp2130GBgJny6i5+88i9JXTuevB1mhba
+yVLybTRcPWZhnzLz8YObTMVaYZcWvdiFef882Jsou0O+7XY02Ami6yqAywRQdzQhPlnUWNORUsk
HR8UBzVFAExUizRWJhEQds1N40ETbBrT6ShyvX/rbqByF1++gTdkfZ0EbTEWkC3MTK0brmKKoCfy
N1J2SHbJua0tU0ob57oqOvzK4o6D1yocInLL5oziRuYsjL2hEluTzgfRvY7KyHpx+3XlxguC0hdB
27P9/hbBf5BcBQYO5HP57DzjF+e7BO4+QiT4auS2H6YifwA8JXy+inqxdn0lSV/yQwwTPjQOPUOf
pVY1IjifM+KMKdDk51Ww0j1YA748MdN+Yk5+agjS1dZIt6oubEzcSkcJGre6UOTdpEmswj0FDh2p
NpIv7zYZ3MGXH/u9HUtHggqLIdiHPKiSwMaUshIXl2l/KC3uN8CMMdMIB80N1CyinbaMcNuviQWY
acZ+7NH+ObzvJpIP7SqDxk0/TiiKQG0OlMrQQvBZKVngzLa9nlNputJ5uiPbFEYR+NPQ/CyXoSLQ
ILCOPszd19bDsbh4RZnZL5MS8yPvDdQQRv5LOhV86PNSU+OBdchqmFbsAKb4WYxu0wrhX35SAYWb
3vG6/Ia1ZdG9UhTDt1py47/YBze5uE64eTL8nlYoMLwNMb0NRVsg/sKQatHc93CqMg9M5HSiecQn
9wEByc9Vao1OgUndeJB4W7haMUvY7TOIHa7GU0B2aVlgSOfS1YPsbHZQwND/nHH7FoyFFkayfGW1
h5HUuJ0uvY+01HACYhZzCDQxkzcXsOrYu1yhf2/xrjjvA5ITHWckp+5hUSHFhgMqHRFBMuIZI3rg
CL+lLUSMvRG+4SbszVCIjjLEfk7DLx3iZuGR4Yex/8TAEwJr1i12m2znuYas21wmDg/9HyKPDCmf
VpNeJ2ExFfiGkPXpy1pIfWQhjBmQgiZUFOKjHxj427aKuCqdi5dYN32waNCEVYWrF9JBqgBW4h3z
ZCixyFYaqCxGd1usiqXeCd+HqGxxBAjZVVEpMi7rkmjbkl9aqh4n2Od7x0kTtpwYfHJY3hovxnUC
j10k4JmsuPPV17TgxNlzQEy3I8cp51S6v0AIUke+U/02g42L1a4GmWjrqCWHGpcsH2wf/InUfuC0
iq0zVIUjjpB4AqZgTKhMO4aKxpc4dDqjo04CqknYfv8bm0PzuISszqDjGan9GxICvs5+G89pIlIm
LxIoD6DsstGn86OwqudRRDTB/K8KDaa0P88AB4rmQ4A+Mb8+ddCoRmf8a691jNbD0UOAYxE7bXkM
QxT5TuyuCLUEpxqZYMm9MPmnaggpxMIMdZhrE9DdQqqfxJZGnlmYa1pC7RxWPCn0ueMsjp6d/4jZ
SGHnCvw9+BeGB6dHDzjHM2J1NYTSTwHWjia4AOn3VyA5QXVHzOIB94x+XmPX2StfxLRDlBSygvy1
DDe5iUIM5snclW5VB6PBlL0STygQl+/ZFVM4PMfubdBVa2NL/EWEawHu6mlwOQ8PhpAi9Hz16Ah9
yQJtYlP/f3YH3mbuJASFWABpol0NjLi2PFgV2xyV62VAFZvPNVLXyWSycyOiAFRogO+FMUmUm/eR
S6I5M42l3MXLytmPRRQ/N2wbXZuC9ebwlRa0kh76sVVVmmwtkSgHNZVJp0UB+/y7NsBzImTq26gr
pE3E3Q6PM1GEFcZYp7cLIpXJ5gEkGEw0Jwx2VF50b5qicD7iugzShWjoJg4Wwe/gX6IAhCHrcNHO
3VvPokdUg6esykxegZUy2dm8IoLMy+jceRXt7K8PA/EQaBb9ta/ISipPxJTL0qFLVLj/4sejrOMG
mNWY5cYSQlTfQ8zVYXzIHg0fOyJ/7Ugux178UpZJV4/oGuA8CLaXMZWxC8+nSch29m+wkx6rv/k3
t4DdfstZUDPJI03X1sVB5X2uli5gOdgZ9IWz53OCTxMQuYSvMxC96kQw9TXcUzehk8bt7eiCqwXF
0gfv91JGvdCzO2WDS5TR6uTNZb/JYs/LfTZa9bCLoiIOm4s0Rpg5ewHMAcjto6LQ/I4jTESHEPoB
+lEx+aKX7gXuUJWMms9b5bhFuQ4C9VjQl03f2XWWEDczhCOqN5oCB0trOpVy5WNoCs4lfk32g8By
CWJVRp1sO4LGM6xAh/IUYMnWZv7nl7+Hi6GULBFe44toGf497noaIW+XvtAhzmmpMpOiLkpQuWLB
Enk48wxFK5p1L1ZJ/UoWkXbGK3RyEs9QsegZlCd0S3bb9TMdB96mBqD0RM/oQGKCrLQ6Px9BZ63W
WMdXL/W6NiGju5SrBjDRRYPvFSp9QXQ20TCxA314C2j2zfCrdHnX5hr2sieFh/Fb951kKgoLx4Lz
/Yp/nyuMloKsdzyO/LofQLzcAasdHjOYd1eMP/7LDhoktTrhQwgY0Aqg+HduuYCNYtg85niaqDSt
AR/wzz9oVZFaV13X8cuH/F7PUypLoEPR8RjkhbnR4c5+SRfz6ooRnZdDRbWWeGpR1AD4baZFxkhg
KmcYUhuDX5p8KMsQjQOQV0WfGlk0Konl4UHzssA/FbMDxtBLYtWyHuCJHQ2SnSjXxmlWdQ5IoiYK
3K0jpgHQbpqGHiyY/Bsm46vjVmdCpC+MwWHj+0nDBALEeK9dkHCbv/AvqyES+YVdzuOB8/HjkLzJ
cYvuRXP29qNr4SpcL0CErnVoO9B6ZnqDF1yewEQlaObHZcf2yx+9dkZDsIMPke7Yoc1lTZk//TJ/
cEDpLEKPpHQ3cNhl9N98zVWzaN0zp2mrv7oZXFT5URaUso0Q/Ov4pr68UEf9CPH2EA7QIM7Nd6HD
8kg4mZ2ZSpTs9MHNoT1cCjXf+8ytspyML3woBBj39lYXP2b9LooBB/PWhcAg8I8xi1bNJriIx01c
mwiSlMivw3xxD224ZX0IAWKNipF9lfMZHJW/kLT9/p7S9Z8f8HS21ipvz5I7pAPyt6DJeOBM0EoW
1+u12h9QY7Cs07WAFOhgX2WmONvdK/Czx3GM2CF58mdVqs/+FUUXoWzK/Ar5lb90Izw8JqGgG7OI
EvbiNLllusHMjpGR3ppooZwDI5P8rEFcQv5OMMvgY+Kpj1ynMK+r3i1Q3Cz6fmLlTRUNNZ1HAg9X
sygA0AZuc+Pv3f5EURFibuR3+lZh+Fak5qIewpglrStXXDpYCkCRQAKpYengMnVdr7CCEd8p4XFf
lo4XdfAFXs6vswhZA8JBgvuPX/+gsLYXIHcbqDy3tedTxDZYJJv1tCO+hGsB9sS7bsO5csMCbduo
jYhenovrlfaNoZaI7BIuN1NooR/AC5GDGyG6qggVA9hYDT+msg2xncN37CTlTc8nQGyZjORw8a0w
+/qzNHJrM+ThkilFmUUOuaMIGkx6PE5MAQnGK1MY/fN/LyNfVI4Kt1l0VutGX3hJ+Lf5h/gL59Fh
wSHW5sgylZH487N8U66HEm7DVOHr7RUve2+fOnsVKhLjk1rH+ZWEBbTa5W3+dI43yupJrqNJoB99
Uj+NSCllQfhM9NoX8LIKVTswS9NvBPpmFsRAGjZU4OHZ5BHStMQTG1gKPzFmuZTphdaUoCTD5NfU
UozhYjSiD/Kbp/UrfnEAq873/C1LNgAJftUswKLo73b7ZTHkGdWbhyujLuqx5Ea9mh3cUC1O1pd3
qh2uyZopLUnPsjZndW4xQkEsfTEnEgh0PlkaHd/YfjfWCP9tZQF+5lv6JQpVnsHNoHSh2hMG0s6k
YbnYFlm6TG9E6uRoqnQRJUCFeRb543ILDSGM91oZ/qPTNo9e+QxD7tl+W8QwCJBoVNrXqeG3qewj
Sy5ZzW8wB+380vIBrjlr1aKj4lbxoWUjiTTZsXMIiDv0nSDT60PVIhiBDgADr1Smym4wOzyjkbYi
5bBK8zm1gj6BjatfoRyAsXmM13N2TJ7A9lUUE9REh+WmjziMMlW3/yVCXZHyUwOrEGqHFid2fMgy
Zy7638dNxqW5cyCKioc2KpObpov9IRZ2SkEbOx461m7s5T+uXEQDeHLUquZUC8Zuq8oTuf81yUoU
ieUkf81cL0lFAprzkKOFz7Lic8Q2B7tiAnGHuD+3dzmwctByPvqAj0W4494geIMhopdacyQ8sL8O
Uur8M4jLPeiz51cg5mq0wli8rhn+R2ppIL/Njfv+3OhSnOl0Uvo4E7pHpM6eMwVji50MZRyaDOYG
IbZBbLOl5/BItxiIPh+Pc+QQePLstbLLShcJ9zwFT+sQCHkp3tJCBcV3GCV4avNMKG3TEj2/qv1P
ZJFnWihUBkYRjBbv196hVI/YN9731YnvayZOvR/YTtXSdYY4Rg5WnSeIqxZ1QyEfilDq4qGwKZAe
JY8Mw9YHhJeZohGFQSaIUs6zP6Q/EE3HER8kPALguj+xtcNCMdFAflEbJxlJcRGVK3p1CuDieDMC
jHbdv0/x3GpruqMHZP5cESA9GS2HjbFur4xzoBTH/DwHcuzh4whOYAsY4IdoU6lUOAvF8/Y3yqQb
HVPLhauohHmrUG/tiJyPAuEwdUeI8Lv9Oo7XfU/XIgd3Wn2DcpE1Cn24lK6b7/azT23iF3QId07j
eCUrlvNXSmDlImzA97oogcUhxShkQASYFff1030rZ9t8nZ99SnNXY/WP3K3MJYshY8wNATpCgkgr
Oa1/QMIYfSfQn84NCth5FHdHQN6wPXBdCN6r7vFtwwt1+uL486rKfjRP97VbCman7zXmIsyJTODp
3puvvfnchPyixPrA8zj0sJ5tIG4Kl5UEnHkSloI/1e6yBlBaoQ0/omNN4yE9kwZmEqFyIoK6kZNw
Rpog4TQEUkUAKQAUme0EBx5PtkpkJqqY002SXow52JDvNeukWyi/52lKRJWK+HoX+Y6wxvizNsdg
HLxtUrhXj6G/glKtr0i01zmTFQqoIwhNMNJ9tDK7Jo6Pom2rI41qT19Ph8Z3/Jkv9uJVf0RVxcri
0yPE/Op2M65QIcKxBUinsxn3uf7vA1tLP9RM4dfdldw6mNLp5y2lSWkxJ8myneWvimTYHgs1+Lhz
VtzVXIPKzBIkOxw0IgkshlFAYHZX8QZyC2KGTtQhBr+xuNOE7qv6IgUjLpm7rK/d7jvR/0fbvPTa
nmicujFMQIXPVRF6CGHXpr0tLgosQKEef+5gvWjvT8/X6xTJfueapU4ya9sptuQDogO3DPivWXRp
iZhZgVCzUEIs9pvBxiLGJX3yBVuN1o7FWSxohI7A88tKTrDB/xW7rden8ZZ3g/pPOuzS9c0QzpGq
oL+Izdje8RmI3iPjFM7Htt8d7jRj+y9AVuJoRqQQFRWemsT6ZrUkKVa52BWctqFcsULBUeXZ653Z
hezMLw29mS/kMjMF/gISQ/VJAax63sc3jaKJLqe7nT4akmLXaE4bbylVHTzTu4j8e8Ho32J2GNcZ
0lXViTZutQNabKfZ7hUvzjqT0tITDRyA5GQ0LwV8tRLuaaLvDXNdIAonHW0R/1QyS/LC2A0IOlUO
X3zlgbQH1kgtmy1GBbLjepC/pO2bBvzhhvQe89HBGtlqviwCJc7uglclfr7m3EIVmq+rac8PTqUV
SsVJw9B2olSMRywMf2Rh7AltWLGrrzTWlZvQovuj8Y9Xw30H/5k5qzRyLGODCAVKFTQxIoFhesM1
U+QMo1E3SMV7fUUI/3xHYNhutL3jFgzSsrOLd30k91cNNiynkCIxrGDIhzkue0VOj1xF64SW21GP
4Ma2FkPr4VsIiC57sEUOFbJlSgQV2c1pwxb9v2ckOF5x1Wug1i+oZWEbC23/JiF1q9BxSNmQUtk7
q4h+s+fnI3SH935gcHQ03QtfIkn/ANzqhO9ViQqoQ+K21IKwctV845WGUoL+xMLiN+OvkElQOpFK
BdqBzqBO+0lr0alzoW6vUY5fcZK57YjM2FkRw3BRRJ78+yeVTLvUxkEF7P7YVfcvIMFoXnlvuteP
k0Zx/VinDXlgSf/X74uYFU7R2kCenOGXLFEVsEKyoQLKhBB3SFVk2GGt3B/MVoy/PCZaj+mtxPBM
UIYbjg7SvI/cfXODbEB4gTHI/9FgXTozgs9sDUZC9zT555Va06UQR4xBEwHTpn8HzyLEQUcvk2gz
KtSHFV/KUXwVJILbskiAlDheFbUzGKUZ+de6904fx0tZ2VEUwvCJDQI4e1HVzFuoKX/nlHdfP5bl
eJK3RO1pISlRYjEN6NAn8BhCwtgRq9y48m6hSlBgIVKBVUqpPvoIUi/EVjdBLNl3keheQarEbtyD
Ry63A/L46vUaQ+YKEhTQO/2qnpHDMYGY+MmR+QuE6dglYZ7TBYhQOsPQet5dsstRcbuE1YxdhCxe
havPXTnjuyxiq6ZSh/5Rt3aZjUBF12a5JW3MnIkbdb9wohccOL+XCXCbv/kr/JY5n7OQwTWSBFDx
Qjt/VlCU6Ncd1EhI+gQ+BPYpEy/Cu+ZbyMrW6DzT8T2IUh+KfSIzlNCBvVlkusDG3C241xBQ4/xj
+L70eL0tpx9XX7fwwdBO9oxcLZriN68VLyejdxao6kjJ/iH19QPCr5c96rpePcZc8QR4RRvwcQiZ
8xLBojbUbPD8Y2hmWg2mY3x9sDCaerjjT3Fek9B928CHzsN4ayp0E7+JYF+dEazDfVFYKQKUxEVm
AoZlCCtRqZgXN/BNf4v8Of0VF1G2jCryVq3guvBk1w7tZjQpgVXyJiKMQn3x4YkIED1stbeQK9vJ
EfO5JapLoCe3jFDPG7+LCgJ8jCrWhnBWOLBGLec63nF4/KX4K4PISd/UYDhbdIN9Op4rsiMYka/n
+XUdE35Y8DzOIYqIS1y5fXZW9fi8XdA7cM7ldtg7hUDehpu7d10KnUGNNtmj/Rd2tfhLiTKCfZ6Q
xbacHVnOuPDtK2lBw7jXtOQXYeDzIi2bPubONboORySzu4nHJSQXALkIx/zDhvshyrC68yiyvw93
DVGzoODCiR8jTi7IanrnvPERP2C6Q5FVC4p0mCJ/hd5bOmgIp1+7zeNljAGcsJs5YE8vw9M86Shf
7NkhXLmHZEbSA0qy3MBNbakUb+RilQFKYbQTz1CdrE3i74IlA0cWGWIAqO/jlEMBBewirKzsEyY8
zvnYB1tYjc8EjgC+XGk8DdfhPOjNDx7B4ftnIed3qeuiBmoapZ3RieX1N+KQUg9FF4PXV+plJ0NT
jpXPKoCJJEcSyqk2GpqEadEvQKGzo3RT2J3uuKkZb7rjzApTJpbZDoPrDiTlBqLfuDiZem1goeg7
JL3E+IlHj9YqOV86c9joXhjbMuHBLcKt526iVda/eXvlPvMpzwz3y4EMDS9qUrnhi2IQE1O9NHtm
40P/K37P3Z96YS8cGEZaxlXEWWFw9Kq9vP9fxaDyRlDv10joB0kmHf46Uz805I36uxU8vb6fa6iO
jYbb5rc6lLX+iszo+e9OehQ3D6nzdY5Qx/LLlyXsifWcM1NdBb+Pjzo7g0qZBCNg4Srqze4tExio
mcbDvDalH9ktS08xCZzWzuUd0iLa9FoFJTK4mESXSIOAaN85M5DGl3pqincdXX+u83tMAn3xZVQ2
jLQniW3QIgwqMXC2thiWuSLioZxqEa1MP2/WfLjHbDu4kSs/UmtpeQBBwqzeJB5b2fQY1JlKmXJZ
8wFg36tvrvJQBOu0wQLCaqUyouX9xrFdDTaoYfJQAef+tMcc8tVGgAekRlQDnuvuqozPZHgXDr9s
JfAxiEgQkvJxNCxCqfHljbgmZgOVCcyv5ZUGsxzp34uVcSl/WImwANlXTLz7KG2WpifkFwouxnq9
uGcK7DGd1g1KRnouLZR3l2wbG7IxFO9vlhYZUPF8URbT9ZKSTgO7NPvH/Mn9jMHAs1tcOueEoJxw
YyQ7ZyPC7IdfdCQAEUf12KZ+/aVYngnsTtF6529GIgJcbRG7hs6oQfxA2pfyqcqqscsV7XCY+vuf
QK79unfELb2CWgsY2vAwZ1+FOShnabOBt04lTon6ppN0NyWQY1pZtp27m/t01j6XK6fIYqFXi0Yk
tRuyjZBvsi1hcj5woADipa5Z07fuqDPK//JSP2EoUIdY8Jug1R2heym0CZ6bjr3QzTy79ykWhP7H
9ogiYsGl/dcz/cotqligBN2nUDPUbZrsO0xmfK3fJ3XBBWGJ5kVBsNDnsXqzlRDE5upDzWewKMMd
elhxbGeQ3Y55P++pP5ueuQcU2LeEwCfKO25UwaW3+A09RAm97xt0teWhczGOqhcPrNFisXU8h45q
bgshE3PjqF/caFvKHYdHBpvJwneqx72qFzNX/Wtc3G4bFQPcAGCuMfPnHzwh2rGp05cUZM5XOz1F
H8SI8bUKLZZboukGI2JGzlDsywVpBczWXRTDNnYZmiiKscAba6SFUQ2BZj/SkGoiDTxp4urbP/0p
NY1mv/PZh4uM2fZx9Hvir33tXSHj7HYB6D3p9ulNEeUC2BGdosvL9Xg2NGaOWoPQJZymxd6re/bN
AG88YExsUrvLX12rCBEqqrBlqSrCZOsGdOJ1tlUsmSvNmqvAgPScB2OWBcGX1xSgxdKlz2tezxBB
4irfJQNOfRHohYOV3ta/AbK4VuHhG8Rd8yFu9Y4yz4IsRUBzDgwRwO5PQGor6gXQ8Jj3pvKT3goS
iBLAqwo8ziKjETvDceqOqGiS6PFRoXulozUP5/OMAe9yCm6k4DWdxuiJ/3gsCYomoqMAs3Mycjl6
Mg5x3WPJHd9iqJIL3q33lf2O19JMzFT8CXrglVrUHVQ1BtgskzlnKH7cYW1qY1xe9I0S93O+hX+a
VLwbSx6jYl7NrO9ERld1t+LlmArfzY0dWmVKIoQiJAwcFdyJvf2DStkFLIc+oOpqp+kUt6qd0v1m
xeKDBRCEyvASA1NsLykSV32M2Htj7HibafJ9muo5dD0d3cB9IHlRKv39HFu9nGTnGX2MHGBG/oUI
815UTU8PiJ3OplvUsjfAmsEuOgrG913yHw+aM6KSG0jilYOkxvegu8KdxDRpm1uQFSrHruDEE/+l
1GT8zcIE5qJvYvY1xSk/xn2RUEOikQluU0lriY2xVZYwnbIzl9gFy9/c9Q/naIWFo13IdznwbiJf
FLC+iH8x350AnffAgKFUqMEJ6aAh5C2i1bkT7C2c28YqJtg6Fztf5TeFz+x71pPru7MOwVJDxqYl
/r21VrXDa7cssp6LwbIPZnDE7BuE0clZHkEeOjr7OxKc/SGxBdYT3Xq7yHbvo8NkPCUGpapfjrK1
sRRgryBjrAMzJYxlHTjBrnKAEV2rKZ+/SFlL7nUnr48/pji4h6hSoN6cxMLg7+5aZzX6fm39ZkUZ
laUlw5NwAmhZgnpoxRhsvbfh+ZbwFNtgWJAr6iRUea9AhHZPKCkxkkXt8ZtQKptJl288ZdrmmGL2
qwP04HCnPK/9B5TDqMI8HAWHRDUP3GfERYMdUYnIx+n/VtzYUepba8fNnmUGUuQop6EawBh+M/Bl
9oyFl6aINhsTUjGXrHLYbYS6+3RSd6lTdb7o0W0rqoIWocHYhYPHL5cRrx+ghILJSlipgWJ7QTIZ
eNVeX4gBtIdf1NyjDvrzU/MYDNqZMCp1eFeIQLT8pdwjwBBa8N8L8JPSFMVEqsdjtFwgWzhaARyk
/CtJYA/NkFljqwd+E9l2wOUkIZabWnTquRhkXMxPaF3pT5OaGt+mgQ9DeQynWTkddN09nTRfL5CS
MHGY1dgbEY0X+He8lfFlVLFJp+o0yOVl50+nZ4Pq/v7m2PBc5dQciSlBLVkhCDCN6u1jQcn2QtKX
khvR2DMpj37MwQnDoVS5alpwQqrS0nDqe/UBlRjTgVRLs0pgVw7QzbHlTO/R/TSNkx+oCRQ2/s/t
TN8bzb4lNVa3h20pZUFd4PWWh/kux+RRoxr/kzhkHyj4WvQ1EOOP6/KTwvIqaswKnogoDPzq7uJB
Yacjh9b7EuWIqeKcjE/bphDaa0mcqvmFp2V64cEBH6UdXZRbVz1Jn7rqylPb9ZA0zDEpfP9iaCMT
/8kuKYptX1b8R8CBINeFghNhgxyMILE7b3qvjM9b+YiVycw6J2tOPqYWnXNqQMT9WZqq5fT5UGpB
ZyznAKBeuWq5o++moB/EvpyK6fvIvaFLe/Dpm9Ag97m5zhgOCSa573OuemZULKCixnkrlWKdR1t9
S+0hayEC++79NVbsTKTNBUCVkyQfJ76g1Mdmj4tejjEtzWAzLDb8d3b/cfuFrdvL268uDU7aIc9q
T+uQGQ0dlakrnR/WSLueqIhnVPDGK2dB6WgfDNSiyQzV0q2SAckijf2FmKdqxNheTyF0K5qReV/K
P+2xOlKBp21iHX3BnK38zaUQ4Zmjv5Zb8u33Dt1dXm4L+UdMprJS5/Zcvwd89X5pL1d1A2sfYDfL
kSkHPptuvGMhTYMeycXYuo8ezbNpvzHvpMHmQiVcJ1PY7ybR6qApHYyGXZM4pjqa1QNMji1F/ZxS
9t/p26RX1lF+VKFgPuJgWWj4pXWJbv+Ib3KxeDom746j3SX7jnSlwGuOZhjf2Ql9xKAC3C5cEpVE
7+6d17UZV45lkfiz88MmLhd7CGRb+FZGrNJPnj7mTro8v5aXDk9OpBcXbiylDWneoyoA7Imtna7h
gyvK4BRF+eI0imOE5wIqlf6yuI2p52U/cudqrDSyLiJnUKkN6SukwqlvzZSyS8+pk3KMJMC8afgU
dqOM/adMpFEJhbhHAz3x0rmko/ZDynvhJrswq/fK2D7iChaNHgGyYTgxQNthguV9hEtPB10NwnHp
ZmML0IdTtsKsQhdlGDn1NT7DzZKHoEObr4erHhPqMHIxkonFLteEx7Er/silJrZZhnM1QSMa3heh
/GVhEdZaS+TQT2C+LNYDVEwrmfoKmxgrBvQnqlrDwobGmuQ4ZXLsfbEnaH0KqrRLSxxd4QTjNMVl
FaP4nloRNQZuPpjwDwzcWsxa83zFvledWTo2IBDNSicGbzdAFZvD/1diBP/QtKVQxjWZV7IrHTT7
uwIDFmx79kGI2tlapUmiRbuMxbLE7PJxii73rhaK+RgpBuBcH4t/uTf81R3qIFXjOmKewqbBAeku
diHJ3tfaxLHh+UeT/WypiEWMM7oWOpstwJddCDsjArUX4PXuj5npkkWduQ/i+NFusF5iR7LOki5U
bP8y3GbxXxjbdiTIzA6qG/SJHQ71bB1TzZYH7xtvdwElj/FaXVT64fKUtOP9FEBbwM7h0j1OXO1a
Ga2qI8QeFYramMYNqHiWXCxV8eJqN3CcjkSSe6QlihOYzHWhhK1DK8JsDpkuZFGtDTrW4IsvPrMA
cc4jF2i436BtS7XFoH0bThCsL9djijc58F5jss8L3dUQht6LgnaumuhG+c8b3aia4HNeqRGHmjy6
geEYFxvRc3KUcPSBH3Qoh6UfhT8iTdUYh+gpXL4cYlLyJkGUfIVafYvWwuQYxr4pbawEgKfWR0xD
ydAzMvtwV5WJbXFZbKhFtuS/aBNl4jZOxXw6zk9Qsp2iZjA3WAW0oaUEVM/G6P/f6G7gLNmgHTTd
N3JuQW1lPV7hqO2vAtI0Go5Q0LTk7OloTeTjaGzjdXQnKFgBUGB0Amgp+Oj+Z2E4jVaCeyXpIXk7
6qoNEaWUgJViP8Z1DnRFLZxw11Rf/wEYlZQ3NQe4+JKCqS1fUo7sqVAhJ5cKVsfInFLj+SSJHH6Z
zeYQaxP78o9ym0YtELBynDXboAIjhpIwrfwnJk9wCb3MDQQBW/D36nR3Z+9dyM/1rj4yiWHTmDHO
PuzeVzrL2LdPDc5TtElfiMVyhUU406tmSZDgz2DgwmrPlSsDMpaJKMWPEpVCIe+yhZS6MF1ctXl1
zYEmAYFbF61O04Igq7sIQa4eE5bwBl4iitBdxnYL0yWhHNtSsmg/W1lCtClHSoz3v8cgQM9nm9BU
nWJQOvKZ9adF5cUfkg8sLgpwgh2PZOugm4IXuCCitHP6/R0lyBm1EbGd8jeJUFxCw0yxyoiCQ99H
RJDGYhxo62WQOi5/ncdgerBLXkY3L1BJkQc+nZgwvXJ2QOBX7azmdKyOGvlcJMQy89/Y+UN5MLnj
LIE9dwE83gbnyKf/JDDWSh9jTUzlvT4cQI7gTwiBrBddysKw01WCStO+gss0ci1cz501tTAub9gV
38jYzQAOHDDJ6k2wS3Kf6WHuPMJJ7sImwzE51qikYKJI4x4WYb/7o9g45LDs4ze5UgMqf0EQ2QyG
j4pwLklTz5vq+Qz2YjHnki2rU29Gr0+KO1BasIMCDF4gspjPyW3hx8gnSuoHZ/7j1IjSxAzy5bZk
z1r4EVCq5MaKHmcxjceOa2PT91RlvE/N6JTne84GyDh0+F6xPCkwW0WvVjyBWy9rCkDlJUpiQXyx
Fjx98WEucamAPPvKDeGmNmUcrzWHosawjKvOmqhxBZu3RkoBf4w2iu9V0XUT28xnE7sCewWSpIes
KHwl21gXecbGfEA1SuzFkr+rbA8XxB8I4i8/S9hl9n2RYbsgaUfwaSa1l3vL9dr10TirwJNCPtsW
dWid6AbxWfWi9cKAcsrNJIkCBI08Uo1ytNx02bAAZv+hkwHiAXj3uJHWr7zILdVmLGIGB1VVTszo
SZxD3RWGY2XWdzdNbyXKd0tYk9lV3R3Ndy/COL+aOElo+xvWqp0eAg053gUY5YDr66BrJUREOgSu
eSspbZsWOXttG8kT7CI23W0rL8vcgmxdX6NEHaRTaZgFY9D+2IMHZ12rXQcLQWmtAwT98pb0IcxP
mpkJpLKOWDeaxaOxhPYpWJof5hsbpQDTb0VnGlwrdMLltiSX1negDV+yJQ2i3C3rioE+MzBzypvm
ZwOZoxgnlV20BbyvfnSMZnbXYHzVdWSoWT+oOj2H8/ziRo1F79RXK/ntp/cXM4zwYXRuCsw49XOX
C6AmAJccgKewADyOZvEMA6YIAXG0CjnB9JGN1ePetxJ9IqWibz794A4Pl3CFUw7B/v6f2iLeQyv9
SLIEocetPiY4ykkgXfCwvaL7tJ1SzLwGMD4j3Rvni27m+AxoQo9M6U8p+2DwGFlv0qOdfRqs7tIm
2pXsch9Yw6cXZ/FtGi3tyB+mmQ7bDggGbhG58QsSoOYbN0o/WtLi5isoYOJwMZNm6f8Ks8a1SKMP
aBtLAu9dYVkazuR2fyyEipz7BC/ckNYgytkSA49n4qvuZZDGoaM2xu4CRbayBvvYeik8udQDTDEf
6ADvTk5l2KRTIjlHVG20nOMvEmg7+hiaYcRhQqqPDyCwKj40qTgmparz59sQVSAkUwc5OPhUfjbo
xAvTgSvkECBiakm6tBl7WJ2SsrP/grFbdcm6UctTsWaZhl7TmwQpPmgx4QCbgoUxjsY0CDqSNGvN
GXv+OQj3OQklS5g4NOtKapEAqEKVk6OBlid2XYcijWw8DiOXocRB4yEoquPnmip+GRw1U+corfiv
U1JUdnDf+6KMfQN2aouytGePg8JcQlSkmbdocVGbCTU4DNZHktkHRDFk12bV4U9Q3XmyMcZfxURX
J0AbInXN9pyeDtZCvqBYARMAExM/eczOAPW0mC7SOJbGfmGXhsOm5uqLr2EE8kmAH1unHdjD5eOe
LomrbZy17Dw6eoALM4iLh7dBww9JbfeG7X38minJMLHVLw3vG6G26PFhanpxadlRmzupjUxvsZIU
w4EZHELeS0oADKdKxvdkQKdWvtGorp3Wx+oPkasNJ+J/PJ2vBB2XJNmbl12KHuoSMhZqRkyWnAdC
zBxjmrB0eHfpF0A8zrWv1BxEYVDQsYHNCcjlr1at6JGEahyaA20k9bV8WLI3p8z7DyuLvTTbsHJ8
mGsZRwNAMqU8Ln7OnsEetVpg3wUM7MYm+4wiqywwc+EujXnxhQWm1P7S899AyICA+FRhl0Q16iJL
hVO/H6OeF1J1ffJOFMMN0d3+Sa9IkR16N5yYhDdtbkzpMYBJUNoq4ysJDwvJOyjS9pNiIVnG/1go
yeAR2Qs2D6qbSbXKUOGT8wrebUaxTLPiYfXmmofrRvtLrxSUn7IyZh737KVJZ4ZebKVuKA67hWtl
sAzAVgatz6C8FGqcUKwWq8ujNGxI6dHCPgli5QLsY/CXhH6fOJQxQ/Si/wJgJi78/c2AO/lmvfsh
iOM795j2xlTnEaFk0w0wVrhyznReqlh7hcghd8/SnEWpwfuA6KKMe9a1WB66SGidIyR/CvUz+F/G
q953OtcLESir80n+KQFc0snkoEsjrYXtBd5tK33cZ/TUXVVs92Ai5mseO5beUj7AAjySx4n9P4oQ
qx19TLquuV/8U6Qi8NiK2AUlVmYxcZvHkwV3srefDQx9naQhj0+IW1A9lJtDrdtLRwKp50pkKcXC
KrlJrS3tjG8sjr+2rwb4mmGdbUV1Z5RC1mVCpkTHTSnaxC7R+xB3r54J/gBswvhvqxn6n+MO5yib
AG98iXY+rxKeSnpu7hYv9Qt86wdrLY9w23VfoSG1OeMOtzwN1/0/TydqkxJ3Bc2w6uyOoPNDlYIj
vm8fvQLN6dvC1A+6B+x+p+bFC5xilZah1WoQPOBA4WVu3PaEgxe7TuungJiBSef6mkn7Spw2NSlP
ki7XyndvEQi11JLuxT8UWsR9mXWjq84p6JmlZne1YboqSyQoc4G5hjgtY+k1foD6rhbLE1CqHu/F
KChdEdI4jmDOraymWpRmUhfePtPunLi+6obRgWMmLmy2h+n72f4xCxYhqsrLOaEAn+aXXkHwOwS0
d4MrXJeQtRFxNzs6R/U2hYA6RPCnrnvZEemokbBwSHnj0eGhJqf1Fz4krGfYzPUMiRdy3fHqkPdW
FpSLdSinWdR1JnM5FaFkaZA3r99TFAK0cpaFet4oGdK+YxuKT64rB8rAnQGiyDXmWdAJuNiGoFVU
i+AeiwAHHKs/bYsISUPBH9Kex8wFxCn51cu41Y+SPxy7He9VzYhXhCrfKs9Z24Ex+DTdnb1nTTm3
u499E0J9CttTvSPm77E778b20kVxl37t3dcgdVB5AWvUNov8/qeJ3qVqp30bgCNShC1CU93+yJrW
mwiPWIX5puUuotb2qFXAQVY5Jlc4pEZUQDzsj34wynO8OSRpsxRRQScnOKEflvQK3ss+wRA4dCk+
b+NpaHfJP7fot0oqbHrm8hhwXE9dZbNYttBc0CfvB4H+RdSb/noHQc3x75Va7ECudlf8KResPNTT
CP56L5XyUoMapZvppXK2HyUniR6YxUo99GhE3/R+cdXm6kdBpvYp92iDlBIfmRXNrytN+zxjz7ji
VeJS8oz0N1XyttCy6K4/uPP3fSR2MqHbDjzQmhjFJEzNgZiGf7vfbPoWio9/QUOrqkRUj3h3Gkj6
XONpd/CKNB7iOhZ2kUVP2dA5EQuK7eDHpwzigG8WT+WC7UJEYnBJj675lhUjDCeXZIR0dJBmSZ3j
efoA5PlUNT29DrnbP8OaXu1EZccuIaSH4Pkh0UAbFIp3iGqlZyWqfxZ1Yh2j9RSaOkh2JJEymTHO
bPkFB7/tbO2YhP/TlloZ8DScR95ykvtO65IlmRVBLWDT2dGcvXQzqy3eSGXKzUr/NtHJJjV28Y5D
+JzdF9kVk1vw8Gh+fbrTgDmDamv/smmV7YKuh2IJIm9qFALV0lrCaXqcVcLObdJIIDrhtOnEBQox
OUBrC/QrzWstBVMvUtLsSY8PD4fkOAFa1oA0Uht2fzVfy4xLlq/C0TbnuIt0ppetcsQiVrK9nDho
wLmkFA0L/4CTsbz80uOEP59PZeyaZjtRN+gwQsMaWYkYn0+77e5N+ITY4tRWnYnRBOMJQK9WN57a
WuMN2OyOx0urwQRqfcltRoTYok+e3OEtlqgKgCoy4w9M7VqaLJHdBnCXm8cmWzq3YFEzFVCAYRvg
u+rJ1wRRYukM+fGo47u41OZx75VtFUyrRadBRz1q35x7ScwGMofBEyLZqOKxzj/OTHzlNaKrRvLI
B6wE3NuK5Ze5cuyq3VjhBY8YBUzkWcv2N0YgddF4+f4bEp4pqQo3MDqWjY9unq9pgL21Tif8l/Mk
iNY83ZfQaIDTfmyJ6zkSG3vTFbqdSzrbHZp81cngkkrOZCJagKasanAco9sMR7HSF1HBy6VH/3JP
VsqukugyiH6fbSqQePHwkgxCL+hX7OAj8m9e4neufGnVNc6RmOJOZxElk3+X9VBpCdgahJl0Xiy0
OTromA4Y/2ms9+j9xrJ+mlNOq/qlNB5LalYQH/u0R9zrhRQXfpRvtvH6NlAAabulIpAD869rmLnr
7El5xpm8QpTbIACkxYnem4BCyzx5XYMgS8ltpzF06LDDFV0mJfPqTv3ISu/DZJmD17Uoomw7JepA
OX6FMbQd+TBf772vzcZyLkZV/ro8un9Du/esaNI3vTgaEeBmJZMqoRE+wCUZbOXPjTKqxa7gSnf2
oIm84nt3c5Gv13UA0Ttz3mtt14/5SYr/aQzxhEpL2fp+oLGZ0Kiojh2Prqi8ZNJQFkcEzH/6/Oxp
qTNWqTGFbzYo24HeUCm4rY1oWuo8QtL3d2RftNOPX5tPhUIiZ/Ye32QbygghojK/zopKo1uexIvU
WEOiz/IxO+mw6hJTCKQvFuvzlXIHRgFZEdYJD8OdZsuxQX1gS+3lqTKwomI+NLi2KbWm09g8OHTg
vdkrbZKclxxZG0zcTkTH8Ut1eA04B++sQRmRmcQ/CLXPS56f8MFen0QfiyR/wk31D8EQmucBJ+XK
5Z+yWi09Wra8DgOVHJ/0AIv/EG4TKxyU1rm8xkXkMyIeSFSUzOouS8xYfsoq2r02p3DYE8EnmIcH
NAP2nm2bzHFzpfiOsJxIwojDrDe4rEi9j38aL09IStRDVE8xo0MCdnx1kLPN20XRPrLM/OxQMp0G
8Di7ir4whqFkbHjKCt7a6JYeiFdmz/MpEAlQ3VKMm3IUdkSJ3CLLFofxcH5+INvwrwp/uk/hui8q
IiNmy8ueSXSiKUgLthOPhhw8KPw5MZhXz/2y5pa3oGk2hFQHaU2bAxZ7pIluzrGNQHGd6m+G7E8v
H6QbxdVrphY0Zl1JRa4eFTw54xvNfqBVUdNLApGnryR3tfySoEiqiWEOtehSiX3VrFEr8duMJ73F
qIViHZh0Fj9N2CnsS7AjZkl56++myMtXOfq68RqGkDxf6UVS2l1e2uZW0p3RUq7Ift8nO066qhfj
gMxbOuj7Ve8Sxo29lPISX5CpGsxx7bcONOf0KNh8U8dBou0Ka1uvhujNkdhWVbhbK5Vf7H8TwktD
ARq3enTypG/NABU+GVSIWI8hiOybjjr0V3rctegtoBG+sJtkLai+IRDhDnBxPmR8KzB4QvyLd2vk
1smaKlrzUilSWVvVdUpFM/f81wmtHbj5ZSEQ8ZoxA/47Xk0++SDNc9LVN0PUMa3CvtSmOEUskr21
DQg+HqSDjGdXuiHs2Zi3dS5o5EFORUH+EwTQoXxTRF29FxLvEfvfJDDQOE469Fm9CdufhgJ7oOTl
BZvhC4xxVanZvcEDUO7gHedik4JliYMlbqyXaUW+VaxWSBEYjVN6KrKENmwr/LSm9URW16BPOAcp
D4vRCEHf4uWxDMSG/z1BX2JOK6Ba1dSwdvgd6eLetKRmiYp1kSP/ZksgKr5UpOjs//2Y8OcVeG0v
Ve+PBj6WvdqTqyMnCiFp99aZhWhs3ROvYN4XY6VXl16uuenK37yRYWZvrcfry81nMo91GNl0frPt
UJXkrs7GsgWns5fTeIrvkNIZOKhj+UL0gfaoL32ADbutlomH6fojs39Ml9WBDYG2fSQa2blEU4ZO
TR3juCSwWoIdPEwQ+MVEV+JHpGAMim4GZXLc4b6uh0Cu3Du1lHb46YQsMmAfjQdj9BjExdWKXKiK
2mVEe0GtxYoT4djp4RFFwPJhXGNXrs2bfOELNWeeAWa4wY7daxxlk1bzJ13YKyS4ntrNvkrNT4hW
EZtqenzLsKrAJg/54xiXZjz2chXORkPK9jBGp6O/D8LK+Uk/WjhdN3YR8s/HlKPC8k9Q981CBffA
Z7DfW7x/8p+c1rjnbNEOus3YPk3HxFqj3BJnYUVF0rnpcAJP834n0LETxKE9PMGQCq0jIg7oJsGY
t/XTveXwW3T3I9go2piAKsedaJGWTWpRXeVuwUQsnvJc3qnKxbiMsr1YsQ3fwe50B/QWgR7yC7wR
7MsAddjmFg4JHEs3eOdDHwHUrgbyftP6EkSCHfZNCDwjIdJMA6u2cOpvWUTUKI8FqKoMD5laqD5n
y79ftQ2ExDARexky04lmyqlEb8va6KcPFQiL8Mi2a6FlUcJzv2SZUKxmkDWQkOkVH5vLLmQNmwT1
gs9nW1NooVrD7DpWtpfYZ7kWwh4ONqs03QO2SL5A+go6IUNGC1uVgaDm+TqFOJbjJ3obxASFJOtS
AJGrEonyeS8yDEaKy2reUyuk6ptNXMiQX8rmxcPqDoJ9TYx2GJFv1FhJoQr6t7AbC05tKUMxGg1G
e09Mn4B9PWaVkpj16nHaaHOtfZBfhwkqZDYqWMJ7rtieol2jC4/PV9GEDIYxn0gw73kg7JbL3DxJ
B6Px1owesEWy83phn+epwScsA8U2rZ70F0PzMVGaeSMpPXSdYXH6yD9M002Pqop7tYDxpwsCxKcv
yZ69mQaVVGKi5cIbDj4hbR4wAvcRdIhsdX4l/HHWcl3g095IPfGqzrq26X1g2ERfjm344e73xK7v
pY+vMd+7PIV/0MPPTgKhqrBiXcKh1QmuNHHtGkf7zBTJO49ydMXsbE3ThQ4dhi2RlqBJGYlMjMmE
8Ae40ePu7X+pZ83Be0ghoYFMaoRBcykEQRZKVSaijzWf5g6PK3p+shvpImY102IBSOOjSK+JJahb
3nDhkemnXBLkLaaq6kPrWqIlrhL+YcPCrglgV8//abtDWxHXGRoswaLyPc/g6MFsTSSxT3LVcCrB
e+EWgDgvq3MT5a9iSCooA7E2yMrovD54xtm6hELlUmZ8zzGDYcnJoY+8RvX/VHZPJKIyCXKjhUj7
qU5F5orhQEt/5TMIQG1cNM1a7K5TJXqtnOxhOsgu1/lE2PwhIgP3CCcw3AriNtyAax+Fe0LIe0gQ
HeWAn2rVIEbQrCy3wXMPTdxM6GdzNCbTmJvdoxaVT+cnexLNbGl64k80PQX7rbiwgf2UiSMaiogJ
P4meK79IZGxoHmsc3CmMssuV9cFbeeAJhlk4DlnIj3A7guuKfg7DWOXsdvijnta2HquD3DQxY+tk
4zJRTrOxkiL63kmhAwK2gi34nmUgg/NghD4S9phtRcRdLWiOuTxMQzqh4h9VnEIofsgghvg21kwF
+sfgylFN/qDrmbv3XybctW88poQiAXNAK+SnQ1HcQGB6zK88w6ccxdDUPlOb2MhF2TsLmd7fMfDF
4c3Sbx5BB1JuLOxckCFw3hRvEsEu7EQ32Xm3cjywR2D++M/flC6DfEA8jopwUJ+p8tIVDcc4ITbl
HtKCaiMmz5Bx+X4e8qtslD6mDwfopxJOTMaJRVvXNau4IyYGttQZ8xfcMGJghXD7V5ccFqi1i8yW
tG8mdCfw6jhiBpSTe70+J6uTEsD/62FP0Amb82ycLUtTI5GU/m61vMGkPBheyRsf/GmxzhYaUmub
CH01dBTl4MfyYZWWsz7odKIegBreB2TEFg5uRuYcnrShIfObjm2x1qDjJ0WbU+xY8/lOxj6vb7tz
5YpQ10i5RnHdpKLRQeULqkPnv1xcQaIosSSBMfWX5ElaK870kuoeWYi+EK1006M3IvgF4oVx8JMm
90RGbzEzDFPfTJ/wmlm8IZLTppQSccHDZ+oSL6Ev1FDNVjVzjg6f7Ik6cZqMMZzG3jCDmHwn+6RS
sSXyv8U7+Yph2qadBW6gVb54BccUtmVeB3Hv40Q819KOLXietOlwo8NBkYn/lJnZ4BX8fR0Kjn/P
vclQxMIBoM6NZFkYMYuCHcNcfCa+a2DTdFv57BiQQVgVeMaVVZ1WMNANSmnM6siqnBUImHp4Cc7J
OqsvcVpDPxPRQR3KKiM35IqMcjUzJMFb43QlKkDoqNB7noDBPIHqeBS5TeY6JtUbF7kU0E2SqHTp
WxNaNGzSZBoblNXRSMyhYEsIAILE+g0+zqBoiBOEKhAEbdbylCNQCtOGlJQrxXrXPHUoTJ0VCrMv
E4TL/mZX9/ohv6ZHcuDl7oV0Qubu86VyKxujcxwTXVVYYtGmN+FbSROQ8+FygUF1u4WaZ1Ic+NEK
csEgJPwzmXX9ex8G/YxFzqw2WJUTieUhimdwyvlze/Xt7rdSoy12Hyp5RLAtNR3qkzc58Fzw4S7S
1RaJpdUcnG4Ux+MqOHTy1DAwzWAnaHqg1RqCrhY9SECGpnIc24uZmnve7a8rkS5VlOKWRmYnSJGh
BqqLBubkQYppJmtoufoQwR7XErjeZyWyVPbAzgtCM0DfXmTkV8XbNpOdEvCd/Zt57rVkZ3/+dboX
fgTiLV22ekIueqwUlMTlfOMP80EHOdPJTmP6VEapeyB2FJGSaw3JP0CqASX/12paYg9p/P3yHjwC
mpnqpjqsA788AZfKWtJoOrE2atkjnq+qQDjXTytOCV1HN+egE9cpkHfKZ5IvH0Liev7jc7Cm1sUn
IvPoM75vgy5S7cLcVyd1LdAiM6nuClhARNpBNqY/PZzT5lrUZEHjxss36M5NGGYNvzrR0xrtkqx6
5Yemf6eHDZtXocIcgf9bcOftf6OTnYOVmXqy6E8btv5S3AYqPtLzEsYL5T78Kz0JTgDVc//V16of
oAVm23pJY0DIa0rdCeVAKpAHWT83lR7SYWFih9GC5haMGbz9fidsygu3lofGCkJYvFTMFF65J0QD
noYcauceTHP1wSsZkgqO6FZ7vcBN8kijMh2H8cMzY4EQ4luktGkhRynikuP0mzjY/XFSB9842VSg
WpnlLKwheGBu5gJHWK5YlzGDJWv37HptD324ZPCXCaaaY7IhWz1J5bHvRPD264zmZYGNbweMEBDN
3C1zF/7D7b4A4wweIfCOc8DtWNdLBtG2FzTJX6pjK6BoZFcITR8lsYzzLWJZuLsvGKmeZiZ+pdJe
tXLR2N12QwUr7m1EULhMlXFGqjV4mZA/9uuE3x6LN8XSzW3F94YoEBCdVeuJ8xnTRK3A7zmVM6Gd
myqFGn/ha3T9th1ohO0sPR+yTRzqdc1xrT9wUKwcrqdASA0H2AB0eP2sfl3c8+rRuLuHE942Tu00
buzdM4ZC2DiEoXbGHJ3H2GytH2mOPLfRxSC4MnKLbm19JapG8UzznVirT5NiWxJtbqYCorhKEnpP
m2UF7F6aYAl9hrEvFYX8aP7+iDYfqU1sOnff4wS2Qt3BCBUkz4nypOeC2sYeVyDZOJAGdM4sI4xI
v98p5Co3lmXYJENDZvQTnT0sTmbWOL7s4oy1zh5jKq2oy8b5NCJfKpjoTgtAyF2DoND79aogpj3S
OtqlPKMcEjPJnlvnDa9yhPuJJnKcopRw01iq8gEydqymEcY8XTW/yLXgAIY82u5tjBgvp+zcJQIj
EZ5UsdcIVEmoXKovveYuUbvHWNwwMoxgWZCBzEi1kfVQDWF0HmVaOxUeO9e6SSssmYqX34BtKLhK
915Oh6I7GXMUBZYXb7XNrU2vXy7ulUyw1GzMjXsqIJ3jkLrmikP77k6w6s/uqbnEejJKIGzUaLo1
CGtJrXGZR4J6t1AyGf2EBLsiyNQPMIuUcUHH7BLOYyIAW8e+FK/BmHQDCJN5zOTFjcxpYPPcwyWT
oH7lPWi8OpolBYZ7yjbZPwqr8L0oWIRWjDUUAaMoGYPyB/aXAMqaYVfJFNaHeEfbB4st6mryKdTy
T2bXFmQGXRFElKN84ALm4Ix9n4tRqqCMvRGS9ZrddnlTtEJfyZEK4Jb5DprlOdclceDmuJj2c3uA
s71j1yuWpeVsK6rAiHwVZF7ZsxkA1y4MMc5kzalmtUqppH+KyNo9uXFM/XSX0GiLGgPO0NVFI77W
gr6P64ApjXgZFueMXLXkUYy7/Vxd4V+f9X2+bZIR83y2QzqhkataM5e7QI4U8D8eW+2etWTCsE36
CHe7GbYuHTthc9FRsB1Rz2fbttf856UsYBGf+9E661bc4PtYTlepVrPypdDUOajiYvdjBJhL764C
1QEhAHNU3zsslgbbwe0prxhTJh0oAn0yFfcPu/V9qSVpejShgmEl2Z1beQzAl10UfDQ8ZqG9Lq+X
8tYwMzADi07wWTeqnZEWU6RSbGJm5/NXSmOrnRYPpU6JApDjslExV1XC/KhuWN0bBnHgQFmLWmea
1ECQyENAawZPA0liCCY1vG1eGNVEZazytbz83/6UNefPhgPujXw/mUQaj+M5cNnMDHEyu0qiKr0J
Bnqi/VGBu2iVnE/1zUqpW+bZiuweZZDna1mR6RsSREVTGt6ZWO1Hv16rgr1dHaTRQg4yCP4FS27O
dPeKeQf6VxfIK4I28N8mBv5RaEYnhf2a6BaBox4jizosEvldPs9A4uifoKSxRI8OpwX5pKI7JST/
jH3rBS/8FapeRgAOTFzc3HSJ4FQMT4QhB2esZU1DJY/JTVscwfHuF+7Ma4MzHdO09pnWXsTyJkf3
xTvTSvPJxZf/ItMaikaeYv0ASCV3agGkD1D6zwQ2PDb2N4vv+0R9X19zMZfAMUhzdI+Shh2Ymyc3
m8EDtvdGbLjqFgLcfVFkwQkIhMb1H8v8Icdmp4N/RidhrcpsXzXPzyD/F8aCBZnSVbi6CCIEdJjL
ZLNaNoj2jwEbkjy1WzRrh0Skiu3NYSA+uwtyn7UBa4VYNvpyKv4fXttp1PBVdsscc/QXipmrDLzH
GzcSj7qQHh2gxOCYucALQ2fpzeGg1zpAxZDW5anXOuDMx8RhJmPuntFveBNg8ZlsUuJoCZ6mMu5+
rnfX2EiM3rxmAKQyWuRyYELuBAZNxAdx+012UqWJQZXRVLInGSItGgsbax1t3ItHqvvmiYy8irlE
Dt7l3yLEhz91T7RjkPcRKlZtdlrYzbheM/Pc2Rk0ukUajZV+Ud4n8c02gKa/xjR0ou3OUQfdTlfg
Q9QfOszu1n1CjQE/9gjr7d2+27B9Ywv33oh5ERYQDGeK/k695SpHHokB6t94ch0yiHMVNDMGY+w+
uaJsBoke1PU63bbUgLyYUVpCIJdjyft6gK3ARdxwNfwCdQGhYfEza/28lwxTxc8GiN6UW+R8fIuS
6H9yZG0QkEqusU28ZlcWeFsF7VZ85P67Xy3UesCKAvxxopIqcYxUvcdNs7Zd0AJdlCUayTu7rDY8
ms3RRK4qrpnuvhH7AX6n4tmmVyQqx2R4kAx2ZU0cWOn/Ef4VzRZrjPdIcx7CdLqY0tFqTvdAkAP2
e6NRdrJ8ZbyBuAqhX+0rVhKkMNlW5i7Jmu7JiY50V/hXBwyg9EFkkc80WM84Dx/snRYowdYVT6sE
soxdYJ71ehRp67hwGr++qi25IVpajKK7MRsZm1u5VgetUf0a110Bpru2azX5LGoXReObyaYeEpK6
w4nmrxU8zCyJknYtKqbLBOI+FWQmYbS26PRsAm+tg03KdYU7oDSsLealUyOXO9P8RRXluR5Sv6ks
Qhh6xEX7B9+nSicE571WgqT9CLL3iomcVfYonc7cT/xWe+xi8hmdzyTWFf2hneAjbQvb3tOFe29x
7EV0roDphZ58PwgT1MS+f18PA+OXyORTUZ1QytBSvqybDiQTUxh2uhoFcqcId1bRoA0JBQclY9MO
gZxPK+L1i2mCjrLjNb5dnwWdceKwXwbR1zbcJfmer+7+nuQ5L9TfEaVBTVNfsVmKCupa39qBk9ZL
Sm1yGYo3e+LQtAEYIn17Dera4yUuhI/7c6has143FQPg7lnxnuUwB2A6KZ2SkF6HouEqAqN/hUtV
JNCcf+KjwQb1OmTF1NwDN7ZwT3EyfW9J3v2ZoLFqKG9907aG9bfQosPBtTXAMfG8ehSEbVDuVrXp
yOdY41dHcIyFBwYgPGSp31PazJVykDvpZq2WR6gM3Dhd3QaXBOibJe12KwLSzjcRfaqmZxTQygcv
gWnkffSJAc+KU7zAJjBQOX4ImUTBVClovb7BUXceBC92myYM1b9oWSOsA7VGkxGRx3Q+I8P+gonD
nXNJ+/Im1Tkz8xssFnBG9tscaWS7stlL/tnR1MgJ43ZYoQXuuJCKcyBdpPirJHH7n1PIyLhNIuOs
kdREt5CoycDyiG822Z/kaDVg9DK3PtvfpvlDTwKQgm2hC+WI4M79itpDo11aqFiYuEaIdiNMv8cs
f6FsV/uAuWDd4FpuyWnQQmYGSUuH9zo0GBPspi8cbce/cndRTVwTuzl/CjpoN1WIENL7FUiiSIlj
hfWVSM1HdimXfmHA6GjnE+1SfUSFMDwS/utQAVxR7EjuR1abcrMY33Y4IBBA78rtzdc6SPmMNW0Q
fv6C9kkozgffRZFl5d7ixR0rRAwz72oeNhNUiPSV82LZcF2sk1OZSjl9nO8TYPFpCrPYEyZyXG4k
2Ohae9+3RypdaBg6dFj3AviF00DW8zF3KyjMUOYeRJamgQU6ezEJUVuSFsTKOo4OFfpeepRbatAF
EEY2GuqpbNrf/7t5JjN8/JLSuQiPaGq6TlSYkp0R/uICDpK/+Q3ra3gPG9iFDzvDP/v6JwVjjB0H
qqVUqZFMgFzuiZncS8+JSFutJYc6zrEshdmvx2NJSTG6j90XNny1kEfYZxGoJ2OOrC6sHuz47ieX
eiwJSdFdqmY4UEaqtBYjntmtaN1jTfXebBL+hyNX/wUHjlqL9XMj8Amv3VH47DTI7GQuIkTEaBYK
BraQ2L29uxuWd3Yj8U0ZRMwvA93tz2STOKO2YDYMhwPeMrIcO4ve2I3s7W0R/EP8Xt/fzUxqtm0h
vpFliCfDJCBS7QXIXvMvEPk/YHxm7ESJrrv+lfMbyl2RL2QkM42KSBrcnOIojCetb1P/54sm7Q6q
dKnoRKcInJJ852KMM8NglEqtx2G4VYPj1hb+MdCeHRfmLSGAuht8w76swHIgYy/Zi/94tI9XLSka
Mkc/OOIJeSOwZxRv+Mk6k22VYbYMUpO231NVZqeWBy4Mcwx1bGvgv5VTMt0j9U/7E4qLp+fwq0+P
1sNuzNS2q5OzQDxz70BVoACS51HMoto3najKGmYFu7YI5SipVFUqyjLCfutrX55j91W6u+3K60ne
qBw8aenKx37G1kKYClxONx4IJEs07fb8WAv5laU8AJPc9xjsorDrD6K9JBb1FskOV4DlxwsDYDRl
VnPHk5MXWnOofmIqs6hGe0sF7w+4HeMJ+qRJPYKgaZJW4esj8g6S0YUAVDSJv5I589pcp9W5HB4c
17KrvfEBxWxpc8erjte1W7nEXEo0fQVAy8YonrlYC0z3Gag/Z0yxsX16B3o6IOz/8RZVMUouUukj
NCagshJw8H/ZgK59pVg9ber1GQTaTU55Shm+quvC4YTm+b8AykN8m0XYnXLZdYHCAu6CD4eD7Ocl
dtxsUg/qFHM3iWKCtDyvIJSvxnDF7nf367EbKPlWY8CFsB0j+pXPMy/JqgbNIShBHkEZRgsMyoPo
qT0BNeArnRQL4rsqdvf6gmJV0pRsmZx/FVF93aNM80rKh7J+sf89m+ZSbH4Ai/smaMkgIh+EZQrI
Q7JFXD7hMHnWAc58UHacUhezM+6lDiDCIWNViJ2GfmsmeM5Kd6IiOP27ZwTmBr98rz9IQJuCdwui
/eiKGj+wW8XDoyYRQ7uUDx/42pCOfeLNtM7d08bmVo8UqUzQdFXnzzbeDbrQK1NDyg88iTt1w8uR
jsAbE6is4oL8XSxTXcJtd0B28UgWnC2Hp3OOQADQb3KhA5XY7C9FqeNt3smFKrrbSSo0l3ukDi+g
Cqp5lNQ5j1+L4ucRsZlziriRkQFrFie0H1Hair6N2hB+0sq2hhpcZBL0zxLZOWyAyHogAdhc/DV0
8T8F8GS/MK42vw0E+c3Hi02Rd7hetskzdvostDmPvlNVkZ6C7NmSK0z0yM2hX5xNT+3ySwL/aNgh
UGR7nkqQgl4g/8X9lICX2woSIvH0a7UIQT6Bu5ifZXPyFNdWNuIl75PGufECPUBdGrTRmXbdkJ7o
8+Lqd5ovKUovyeqIJxWTsxtm9Fd26D1B40bupwJmx0iSZIuLXO3d4EG9zaj/pWDGjFEGnSTwVc/v
NscM4Ykae4BYw0Suslmy1Wgg9vt5SY7lCeL9O+zgs3EubF/3Fx2VSKeiqQPIApZqkVb2QiOs8kCb
PUpcuth4cuBkOuEEv5hc4StMYRxuL1tZ0E4uIQXaG8Q2pF5zqGCjCkYXYK6slraYGLEoZa/xZ5a3
7pJPV0HABwA9Ln/Fy4ODsGZ98M0cfAAvoAu7h+gCErnEZdttQjzqkeqgWGD3YjdT3DxP72jIpuNb
dsjiZPd843h+7c8hmHaV7ZRJg8PS+qbhraba4UOTPbdtPESquXtggaqkR0k0+FwTpNheN+o3ehw4
HAdKdqs73/JWsa2kM7HIS1igFx9PqwHD0BnSdU2iqVIXfQTpnumdrEDtjaNVguhxf4v+dogtYQWk
Kn5WDA5YRh2VprsfYmvw4HpdoHcqodo4jSrONKFW+G0vX9vfniy/TMzLY15SKsfNLH1DbXw5kUiJ
RjEMT0ifZ4hjAA8AqQeS/xWpoxRKT8zX7J6AlMK8Da9rDjIOIBBpktdSLzbkoF3lP932Uu+qGl5R
/kocc9dcQGGgHPyDReBNeRI06WZy/KRtn7A58SQtadf8d3yqyH2ciymHpYKoRo8t/jOE8ai6tVRi
vCT7xXjvncI/4PEhVzZfUUGMnJsMg0g2Pb0gfCStJaXKhdyOonls3uMotLw4ObcBA/ckaPC1rL7p
qBE4T7gx8pJ/hfjlDp4AAwQe3QadtoCT6DPNiYY4L8cAV8NHIgo+De2qenKyy9qOdb/lQUk6d7Ti
dd+/QlbNf+C9QwC41DlYkriMhS8rDkw+3lZaE20diU5NOumEEs6Xsrqz/g9xoJ9dkGV/XDgPNEQc
cxfzXn75uFP5xdDzLnJCgkXkny/5GeWf51AQD3CfFErnYpxHPvF9GOKYiI7YqJAGBnbYWleUsI0/
r/c/wVJPbOHe+M/jzlFqfHAbrIHi7cvxHKdwsLY9F0VIEtousRSflX/wcrxbFcXtMEXQ245FGoj4
HuUxpdM6Bx/ngbKFl1KLMXTiNy/AJMYJ7P5cUi9L3e7E873V3RovWxI+cTEFUdUxfVzxMgX1w+ym
IQjgHVxigc02M/6+WDR1fTeDAAOgUpyq92pWzKcy+36Mtygg/7o9CU6m7glk27nfdmNHui8vzxgu
P13i+cAkFPLeRBKIJxhPZDmyZMRby8nhhS0JulXZEu0ufTR6KhwfROa5JKsFeYvYXhrARWPBBlO+
FZ7t+Wmq9bp2R5+bfHrk8ZrbnOLEPZT3eJMsrB/jGSNh2D1KOdZ6jUVUj/64EFSzelAl3aGdFNgo
mEb+LVjuZEn+qTOhN9qyWWk/gMvG+C7igfsbgXUbxnUAfU+vjn4KRdltMIN9d+ksC5Ty43+uHQH0
A3Jhk6/GX0GvaU3kpCO4B3z6FHdkvq7UEcTANT8bNCNUW2NQaDzwY2xCWjj7wS3AnO4Ca4fKrP7c
RUAvHZLrYmqMEB9Av/wBmaknTyf8+a+TyXIxiPsj+f3wB4VVbChGzACUPoVl+jxlVh+rOh7/OPGh
7Ai97nz/qP946c3bQjVzx+KS/EnhVCmg8juVcU2KwKw+bb/zfu4eU4vR4BPfYOZkKksvTyK9bRfP
D65QoWn8y4b6VWen5Wav1kyzBUMCZrKjVDbsNGmy6BcjiPT4mtQPKh51R/C+q8AQAeVzHcyEXQkG
ROEyEDhGeM16Px5YdPkOAUxnsgfPbTeIveKUG7mdFPhcpL9C+87wlr1wBolaOPkVNwqiTfdTjYDW
z9UZCn34W4uRFuCdMBA4yd4SeruAOalsqJMRr02G3YbeyIA98FUDc6z2FQQgCNxfQsaoM4Cm/uOV
xwfhDwVSdLvUPY7GNJ2fh1hcACp/TaSbi/yEOJGzkZjpLEtVtcs/tEDkoO0fDrwbY2YF7Aohk6CK
WZfZgeuynbv/Im1qy5n94WLjHVgM/drO+Mhig47gzUzs7du9g0K8pWyrNXRHmqcbb2nIoCwGoI4P
df6k/40oEGiv593kQRaBLY+y0B4lxRYa545BQOkdyQSrUxjDLvx72guVB/UjAFDYFczJw1HVCjQN
XiKrFhD8KnTBnAEd5P3EmT03+E2xD8kZFrQJNXQkKKo1MDC2DlbQO0P7u5Pa13W0WpNHBz/QIzkA
RZAVG+G58jNyM80FD1m+wEP/12IlSdmzH9ud8lx0mGs5GzzQvgwKwbSrq/4DaUpdmU184CAxsOcB
XX5uEW2De+4sJtXsdmJXg7qmWPQdNy5q4ojgRf+G+wTR2JfecBOU8qhxsAbmFb8WjQaC7tp+XOGx
s2wLaSmAoXOAST9PNVrb4CmBj8uAFBBpZgdG602+kkjQlvoom7tgE422ODFKloJbt/V6sUC+FUkp
GfCQbGjqbzPF4MjJLVpXVefAjvU3ytOlamVCpobkbfqpz/YPScd27bVQxU4I68m+BBmEnskf5NRb
Jbdk+6zbvhDbK95N3oZF4lFOMD5PxVvAG2NXKQQCGUtIHMUK83YUB7TjGyOMCrkUSS06wsPqAEgu
yamNtH7wHrnsmbx5ifOcM0+/VbeH2CtpphyPN0YzFnVJZSKmLbLJPj7o2p94inlftKrfPiQl9767
mtStE8UYKCtwVNusYOIALPPHLgg23YAVf5qqcbWZ5iplf43AHW8xGiN5Zwf9H4sJfRyZ8kDwRssC
F1zfKuczIbolH+B3D2HS9q9FdmHXpleBwUgUJLcIZUsgpBdPXZq8TIW3lWmU6cRfpTlxT6anKzzx
jWzuQqEUe2z1utmJXQ71nnHF2VaQj7F5TImEH1jnZ58yaiNTvx3vlnOKoIYswKZQTm82LXkqlsFC
T+ljFL6pKSU6Qc64OUaEnHzumtwEFlxMOjTeIvNA8P/3hJhqcRW+YC8aiE8RgvYPlH4byYG5rc3E
iaVUwLrjsg/rTbgoe+vUcD0aDTBU/VDTDJomVRTh6OYPhcoaAT8jZhxjJKAflkc/mNX0uMWV+chR
fQ4Dqr3EjUPFpcZu5eSApOPRY+2W1q3dKSgtCSypOYZEEFAzEhvRGPr1ua707KDg8bwqjeyYRJSK
5yOlrwkIAUzCadoZN87J1/hH6OTftzAhFtqwGfNNgcsva7bAAaNgtMfBQfcLzVhilUgS3qu7UbHg
HpJTMVfyLvDV8CvAfDoouiEcmlqYJ7xWdVF/gnaxRgm8zDX5jpTsa+gpoUPk4FnDatEhi42+lK6a
Z6lK3hfApfu7MzLtXwCJK+jcWohc0XyHf1VjWCaoOh+fQUSS+ahMY4uZvlnBK1QaI8Zd4Hv9U+rm
Wy8o/0z1e16XE1/b3NkcwZdspRkYDzcoUL8ins6BIGN5oI5zAlshP0nIXTZoVXlL3o/90saYQVUo
5FBftwYxhhdN5eChyNncZrpEctcUa9xQPItMwHG0evEUEa/yewLdyj95LgQlvqSLsiHzYizUltQD
XhxS6/o6JtiAv2VrYbK5ol/4J3e+dfGSCWn7BocQPkPq8zd9rVm4IbUjlZO067rFojNpoy8BANVZ
ANMvOnG0iXlEEoIKB7l08Vqq8ISdMOEk57ua26Y+BtLR24KwrK8+ALgYMUaOrqZjAJSgJ0nZCpab
0pE99bqR6cihLJeDfw+LxWLoIqqcTeDEgdi2MmHr3BWG+fngSFCLGs7pbCmNdffQgsYhzIzp22RW
F8v1BaNIjtcgueHomR5cePvriCSLxf9k/pOl0QmnjMIXJdPfaDY5Vj1OASFukdx31jXfml8a5jKX
2IuKTRHFq2MQqACBZQAGhOmKCbiMEj9kTmWNg2vYS5b6nr5HzqT2HGewRFXzcwFWIQuKIJaGRKRo
Nk7MTJirl/2YW6lI2SnaTWa0a1nsHfogjOxTTLqe8ECDmD4WWME2SOZ23fx7Tnf7R+kEmc74RZ1U
nhz2HZxsJFwb8PqKDkP+SwE81/f6NQOytRPxpDjnde3qQ/gBM3jeE6I0XmR9D+HBcrdvREoDxqSn
m/9052IJh2ulbnS0ZITSBxsLeuA5ctiB98y7d4L61Ds59DZX/ukLq03A8tlGRSw0o+LlYd0JdBB5
Y1YyK8DguZptOsqQw9DLSJC5KwoDQAjf+FBYphDgQE8Clvez/KiO0Mz1AdgmQBI426QyUlzXsChq
MtzgaIHw3fY0omaVUMbO5TKKjtxbjyfm8nw7gWd/QMoVW1wL37ucGzKkmChsTJ86uA3TGtklMjGc
TuFTO8yVTaIRdpWU95QyTZgKlnMZeyYZmq3oFzkWDokJTBQQd6plzqeneEhkaoIyVvsPrSQKD5xA
WV6yPmjDcTbkyuRYNvn3nnEbOokUlM0Z9vl9oV5v/uhueKrc3Z0Oebe+tJN8v8rs+Wg3xabaengH
R8S1deMiQ1VkeMmWO9L+HOoYZXVkXBmwk88RPDEQsUDVX7yuViM3mL9I+cikG4fHKrOHHs0yAYyY
AIwRTGYcCZiVWoMqanp8aXCbZs8ojzyfQ8m8vgr8aQPqFL6m6aDgKSoxqqAJcIlEn8sWiEYeyDrs
+aDkxSFkZn8O828n10TCg/PgwdzfFcIuKdnc8CFO3LyiDwL4jOVLuVWrXDTO25x8XcuX8oruqxHu
LbIRSZzmNu9XPuhsi3D61re8fwQtIaq3B/vT4UpnFXUyAKn+6nzWbXJ9eHmzQORJ10MpeFHTwPRw
1GS9JfGXtTC2FH0y2akvf0CqwkyofwQyaJIOLAR36phUEtdWQAYhvc4cNzZbTxEkcA7nKFky8Npl
UQyauHihpGCraEGUZQgui4o6iSO5c+wURgGbWR6LXQEYfmrClh9P9Mdb/75WfLmpnaD1YAkEF77N
rx0LysXqqBDOao2OFIhe58wchOCw59ZERlPerIKl6S2ADB2LsfRrWF/7PkPsQTzgJCo+KbLjG8gZ
zI/KXbR4amTuMcW+fMGVgNsmIHpfHtFwun5sLC1m8iRBHP48QNG4hg/5Ps2KfpJ7GLvZXwaCPG4B
tpUv30vzeZq/jrwO1FRlzFvEWa6ER279dlYNMCo6kNuF2NH7c6taafasF52SAypq47RjegtKTCSB
1fS9LBujUswU8fOg3ZMTydl8diXyFvCUwjFogbGa0FsefKa1uM29Z8UTMuYrGr47gdJRkLkz3LMj
Wqijnhf3iYi062uxSAE9loVkdr6jz58TJtTuyEmSOQ3H2KW8Wn+fshn9JMDqEtu/UDt+cHveA0PE
LFwqQiAcvczF72tHo5GfeLgBfL3CfmMEkYsyhSixKoUBtjPR+5/khXoqSs3oyGp85LdVOGpfrfC8
7HmIYDJ5rrs5uLaOaHkaLtYRB+mvzNC6GL70GsjU521qBxsAVGgbyiE/S/NsJMO5ZT8kVAPnKePj
3GL0SeoTyKy9/0N3bUKWXiVS63Rjvwob9iT7Jl5ng5jSXuYUNUVYg1W0QAreuuVp5BmjJvTJZjWS
89BXgWBIT/Rl9f4if2+zvDcU2UGKzq8vtOfsIkhZaXrxNbjHFwTd1cWgSIxaOdKanLnbz9wDwQza
AfHwL3DqEOEAw4gq0NZqM1BtWB20x0qI6jjAOyjLbexNT2tDCAj5Q/AIwGhBJ+MNE/E/fkbDgNGr
2mK5bcqnN5m61Fo6mHl/BzmFVcz1+3X5iiGuEiKKxostdmDhe+2eiVjFuVdWuJTMeTV5UfuU6Wqn
et+pdONA8EOPNedJx7GdxxXcIgQWOJVUCI6tv24xd9Fgia814bugHJDclZF8iB37x0ff2NTiNdTe
UxM2RNBA+215QKlfBVsBriImkZRf3z7LZ/jfHnezoEa2Nbc6I7Elush07Zv44TmShJ+PlGNnKV2h
rmuoGvfKxlujG++mrq8RyTtqclFDf7QDsmXX7FZ4TL1AKDxLd2uylHvxjQqh9KQeVJ/BlpGxgj1a
6LnDD6ij5PYHVBev8ZJr+YBLBlhcpiWMFxKo2VixDrls294J1Feqk/FuN4EkFdQ3zFJPTVz1u9TE
hrseGEhdqGl/ak2/BDvo2YFtjyuRJoABwhJqD85QMjurXd6dS6/3GJvOEz2whTAupCb/KB/OWy5e
KNfD25+c8CuFNtnniiTK0Kk01sLd1MkUyppL6FwrBi+qkdzEop8ZGL7wcCbrmEEfEubrB7XM4hHD
PaICjAOCMxebFaBYXO+6Zp7LbqACUYpMIUhbbV9akTEOeIQE/WbE6XdLwPHh1r+f5NKZJlwK3tGK
Ogih4/crX4eGMOPYLGEP1tezY8wJ6r4UUjXLPlLBNhWGhXS6T748wYcuiJJpesSESHB4xGMB1yIY
f/5DmE9aCqpRvsI2Jk/GZn9HSGkuY7FT7Vng+ZbVt5+3G7xLDEZKKa6H8i5aGgKI5pzo20uaczyZ
mBN6t1EgYWpNOC9VjQsXgugUVbP5MYs9jA4z8V9UQ4c6dTDBidEQVAsjnaS9DDDPRyqoC28YEbOi
gqbgSdbjnpskCqJUkAAKcGZ9x8XKON28WAQLldyHju8c9iKGUcfGcMv55fwwo++QJ1pCugKcDeuv
5utTLnTsbeMab9eefUFeSkUUXZQr0jXMUZH05uYEolr6V7IngUEmm+natMkI90l/tCqBS0fde5Bj
2ObTGQwiZI3QF10zaVRaNENtnPN4/RqsqNTWi/W2y744okv6PPNlxZTOJgp11Xr0OyXGkbo1DJZj
5sXQxz+uPmvcrqqORG5wsz21aJhgyY3h+VtAeey5T5v/hOl8JXh0IxZwfUuuLTvjUnxRqPYA7ShE
ngtSKbwDQgvhCu5ze4j0TJmx34gm+4fd/bDnyYQ4ZFswi4HyoVbGTEslf0Dm8/x+nn1GMhfcJ655
jxLHP9DEgoTG2VkBf94acEIXC4VKQo4e7nH8HCDl02nR1x9k6j1IHjHrWV18MBoqrsGBSgWPBet/
/GRT5bqC84hxP6vew4LoqPx+HlE0sq9Il9ozhb7JtJkmeEuEtZtYJdjxBOF6R/k2h9/5d2PxgSPO
CmTUaM7RmEqDrpzLW2XesfP+gK3Uu+3ylZoIn/1vzNTplKJemAcTUcoj8/7eLmS13HRCWeEXs/K1
6/PgZaUM4OTfM753WiTDYiltmnrAsOh5mMXZM8Mp0rlx+k0IGKN6hgwv/2fTUCEVUDqdr6qC/2Zz
iDcATOYpHxAfvkmUz3uiXucyeBrBXr1HGLhjx3ya0oAut01kH6xWd2jKVxFxb0TuIknHvCUqZREd
pgVEhnakhkQBMs14eWPvG2JnEgGL0LINxunx9RdGH+XrWDoDb4sNIFvd/qFmsHMyvQJ9oHh7B5ZW
6EBglOhu6TTD0p+8hEN0SN4Hh73Z7UR/usJiRliD+jVI2vxeBGmdAQ2bkR0aJiyo/cncBjxqoHJD
fTP04S9xACO9P8ckzF9vZ3GPv98YhtGNMMjFq1P61/NOTs5UDiVn/NH1Q5CXm4YjXEomIw34REih
O1K75x5RbmJu1rMnIZ6gbvVh94ufutEFqldwEQ0QBnSHu4//3VuuCXCWZ716LmvGFeSYwXpxj9xK
iDMSj8PJcdlN1PUtwZywns/WyLNhsatjiokQawEG4vCqDu86irDICW68pBdc+8B1rX6AA0Jx7i11
MHAT4Hx3+wYV3siGVn3R0UEwtBT9ZElLZmfR14AofmpMYJU2b1h1RPcEbenVz1UySYxhhwZIjuxS
ab9gG52+3vD6SLpjJlNc18180sX0GXyKOvgx8EJLeuIdqm9aUIvYDK8JQKCQvaEJNO1UIdf1sYDl
TuyrWfwafMwir56DuYMyU3QkKAczcq30BOJ9q6F+4GKiPUaEGJN+yq25WJKZRghxnvgspMJExK0A
f5j2cX6vQBQLWWyle5jkH7yHtQMmk/TkqZ6npzysriOsgr6wkjK39oaH+zLJG2nvgMpOsZWwtKVz
CAySM7+/KmBhFMDmHKT4OkhYQUKxkh2eCBNx+dPfiUq1/7BrIryaATRs4WFdEdHKthqsj7iVY9zw
akKZ4uWk3XbatpJEcMoLDyowb/LTepHF5pOtc9pRSEFtRJ2Nk14vpyOiCDqsh9UdXueIq6DoI3i9
Yq/pQLP5w2vU8XM7cGodFMfTC8NdYfBRszXBm73AV+qZKMlbfJdvK8MpVsT30NWAVbhrnGm+nG3a
Dmny6U71z89iSvWiscHbOeGFEB3oAF4MbqgybLDY8LibVrpz/oy3QSRKkzKsZJbOaidhNmveZFRy
4yoSw/mKoPXYTNh5uYrBny47Om/+gKKUPcPIBbg6BG6L/C9fbI9+fzvaXow9FwfE12qJraaq2ARP
bWLAjRNwSjPLYypZJbs4VgeJ2gCT6wfb5viD0jc9iJhuh1/UE74cywUS28DUK89ZN1gxydb1EslI
/0okY5govhMlC03zuexnd0alSBBg3FKje/ONNk+zWeasn4M1O/Rd8qrMHGOWBiVX+P5yHaKEZNVq
P2oQrXZ+c0o471m5bOjQWWTyLldQJDgPCtisqI6e+srnIdP11y9yBOqi/Iy3nBM9hXyJUj5pa5Js
GTFURu7+cu5mvXnJEelz1rL9hvj7pH53gBl9tjByZqqaWiJyMjLv7uX5VM8rhuJz68V98rMIsR/D
PDzEV7LUhaKeW44wfMkvGZXA1Rb+4kp7KmG/FxwsKwLa3I7FwZZFiYY4Y+8TvnQkMFFIcX4BrduL
qrVsFUKyHIwm7Fo/Nr6rOx5Sx5YyYQMsuOhQlsNdvsAm0f9o9SM/UEr57NMLHL3dTLB1UWUOA5jy
f0bLjMcHfM2dL6QN9c5jCslTxwWW4f9Swz4ryxKR4Eys23+1wzjfBbSg5DWWGdEQ3cRriYra5HJk
T1CHr46anbdHOpdXcgtKGLNY8KyAT7DR6GACm0B1LENJTOMDrAeB2DzdJKWZo1cze7bGBB3/idK3
POhdhpKp+xgGThrtGN5g13KMn5FHmuRQGVbL46DoLzEAL0qkFIFJD7sTG4kGNUtBTtw5X2iKGCa5
R0OuAaD22tp9LGnLqDH7A2KZ11MU2fbnko/I2DEqnoZqNMs99xWhvZWNoLirgl7OEtWkH3wNcKRe
pynEOJyu8fE1GDHwcXxxw1m7vqpoT9qOktcbfdqccetzEgUmtOLcjtxD1TKkBLqT7ploNGXUJjlQ
5ekU6yreeLgg+4wHVwIQQ/ZCS6JaB/2PXHJOmfav3RIwosZrXmiLJfK9EG309kj6FlzhxOJLAHrk
KLgaRgIV3fRqaS1n0AvmtNRBEx6pORE1Qc/YsU9bxJvroDJIIILQ5H7XnBQRNCxT1RCzbAl7Bg9D
IHiUMeRO6JT60tI9JPGDRHobADQQ3x3T28S7nTV0k0Ta5FUxenvvNq9X7iSw0JgTxWVqWJ4NM2NC
emwuFx5b9dbaT+RclXAwU5yTWo07XWYDugDhLGkA+i9UgQmQYH44T50W0dpeGP8P37osfdJmrmYH
q4UEEmxNFN8MQpPUHLURTFR+/MGmBixGfVat9leD2aeBUGAJReetnrHToRJJwYbz5PvxXOXcRr7u
tAbNOVGdu73839M2Enf32sRj/KHYMJVC4Ggq1BvXwMFpvTBlXqJQP46GBN1AwpdHazVx6uyWjpkH
Yq/Y0bOa1l28ODBrxWj5Ncy2AG2EcesoUeXDSk1PQyoYv/KSks58RgZU3MGuSxe2kNZAuZfFyJWG
1iMwE18+ZR67L4jlblFVrDppYPsP7RqUov01ypGrbIj1VvAv0/kA2GxOh5T+vyiwOz2//ZU9Athz
kZe0Xj52JfUTc5GIOgJR8cMu0vva5HjHiyzeLtxMBgTVT9sPaj8D2Srz/lkn1UWahvpBP94hNDyK
6jqD9AoOb8OpKbSqScFE/RHA0X1o9k2uXUiwNgXFxtJaxcIe1UC+vpZoHJrrif0K7TiSjxF6Rj1g
v7gnRa5L7l3QxysUuoEwCA+4PNhsG+qcOUtsabd9FzdvZwFz3761Ns7+R77nBQfgKi+CzEW1EoKu
hfyyP2BkATJyVhnoN3Xot654EfWbn02yqzgpncW66KMAr29euwh7BOjR7B5LmgM5knjSqpbJ9Vmx
a+VU0tFbleyH9MTpt1D88l4HBhpsXmonJvXu/XPxi2f7zleuGjqkRrVJPshlrlhkVwnZb9RWZo2F
xuDp0c4aHlIRYyD9tc/r//9X5pzTA6BFRm/nkZxhfeyyDkfAjp8WIdePxudEGSL7G4x2rRz8SlYN
SLAqJEuXNx40v7cuNqoje9VswP/2rep7kS6/TRPzoQD5ogOi4MN0wbbeGna21n26NC0hAVZ2GyGO
pCcUZbEfD8ojrAaiu7b2KfVYlMvTcZmKQUH5g4GHKIE0ms6LG5ssHrg0r5ms0qifQEX51lKHKQmW
7fJvfrdoRvbzwvM5BnVnyFAWmBE2+yavIwhz0ojlN3SFE7Ynz/uoMTzaeUjnJxbhGcO0KSxbtQ22
aHWopK5tOR/ItTUg/Ei80/HfSl9hsk6oZXOBP5kokiDMCDidrhE5cY7N0x/SGNimmgi3tkLOY3oL
mbrMxxhKgyHcMup54maRAcDyrFlkbLU6AOSi+Ra5/48a0HtICRQxv99Y5WTomapTYFzzD0gNYmwx
A6nw+7DWB5eukosF85j4MU2AIdzkcqs5c1q4NG+Z6Cizd2X+rLFOz+5p8PzHAUsiLHYYH/5jxsrF
Hx0MGJUjq6cL6Zgvk4guoCArj6TCKKku7C5JOZO5GeUSP/gK5rmq3v8cPTgrhnJ2naX4aXcErRNh
NCx4YjaRYgRXkc8DkbP+pHeaEtAZV+0pmdKPcsWATDKvUCtRmzxQDPc725s5pn7WYyMeXzc/NDBq
X7o67GnrdzsfvqFeWJvD0i/XhebdN6b0QsZAyLwGJqjkd5Ai/UW8rp5C2IAQEkj/n7n48pavJ68F
DT7++p0a4XSVUquCldQiLlgPL/6MOY/QTQZikJSFaz63Xj8hBHqjJwFubREVvBKbzjG+5AXufp48
NogUao3n5juZSn0BFNnPJD4xQEE+Cv6yIBGOLHMvVqyJLgUUNBKgQX0wEwZfWaE5+AqLljkQfBFG
9BpsmVq7+JG130L4Im5eSIbtjtqUar0cIvHciJFdPw+oLIS55i3uSBX7pX/3exqDh5Kds8idCF8m
0ulfykrRKqEeI5IQC5B0GCEgsQdwio4tm0OEwIxeWY655eILh7wYDyLrNO7PBZ8CBHUsIvA+o70X
KbPMg0dx8cClGQ3HOV4m67G+jcuxK2LjN0rbbPzOIWnytOrVGLd4x4BkfSj/iyI0ZBw+T6YSoXIc
f/X99h3oNJl803yjzA7WR7ufez0OZdyrITSAZM7VnVcf2x6zQxVAw0ENp5vAy5suYxzzEo2v9rbg
eTzx6Oo5XmwU9uWDPoCKqEK+CdoOQZqdeU166AfotJDyPxll5CNzwuq2AbX/dGvV4Gzd/2rAYj3N
pxdqrDEnFOocyGzuTm40D09Mhhy39vFGyX7OtnPQz/QbJUuM3vTtefBN3JcKI+jNKCHRo2PbTelk
jrjZNZ7EQz7H/McqZw/VewzNq/6TqSaLgStGSLpsuxJxDPJXkYDVqzuGHPSVMpsDyW84nqwwTYBB
bZLVyzf1bTZcGhLNnogn8fP6UKErkY4QFCxNuKrylV1K7LtkBZZoYLUGNk1uBu/VD9oo36roUobs
DUQA4WQkPuVgn3WvEsaMPpnt88Dm4+/vWKO4NBMSMaEk9At5FZ54nDo1ibcgxhB3CUEec7IX6/bh
00xoLtKATWh5tL/u/jUSa+DcitYVRB7NYv4reUwaDM28W9BsjSCjilqtJHkvyLbWXAs+0b6LH9rO
5EEaISx2n1TW79iA2psRn6GOsAzZHyCIDXhdcYwhkz3m29YwVnkiz2i5c4CgdFiJYcYvdN3MyqID
0WPcdK42WHptjpAaH8dGvnkzFJRFvCUCxPc0PttfGJMuduaP7kZYGRVceCeA2uysPjQ1cC96DTyU
a9bTyLCz1scWjzM9t7SZcn++/0efYI3XqmUoDpii84et8xePu920WpZJ8JSqc5s5nukwIXPNsgj0
FgG+k6JAa4OKZOD6RuKQnlf48ne9uKpULFfco6C7dLVAu0fvAXOHbOnjGwzJrx5w8IIQynWsDTmb
h3F+ESA5lu75GqQ3FHUDycWsRVRIkrAfA60iVgCXoErUi/5WEnlvZOiBxUr8TjBJDKpu4Jl4Tkm8
f/jshkAbq8dnElVfL8K8VyF/jHArVP2s7X2Z3MQq9FU8CZqoixXi/Si3vwefT/ovzEMiN7nApM19
Pl0W419Y5kXijyK+TmavCqwhljXHleZWL3i/7Q38LrUZhVqnpdO75H1RVGCoEO7vEPbf5M7I4IV8
HaiJOeZ5jxWihDX9MW5Mzy34NwkexjX7bxgwe4BvG5NCHmHqA0JcFUV8ivb57QAIUNsv0WCQPin0
L6foQtUfDUJ8zbwMSxTOavfqhpl+bLxkhBCOp7hvoeV0/PJYHZDaHmoENqydllM93tRPnNLho5MJ
SRtr5Vld6RJQNR4o+Njb6STaVofev51u0P/lfkl5t+IH+PvB2s+C1eRzDseZbOtDCGIk5eMkhHZV
J9InlIfiVcyWrXqgRl2mYAErCAJz8X0byivZWwjXd/2zePQ1/QJyts4eB8D5JLm2qi9PSbTMaDHs
y9tso2rdkAB92RiNqMx8ew8yCyo1xF5uiKarTxL110/foyrIzrvPs8DjZoG/jMrMoYpUZwBemf31
KAezT3+GGB7MLSGKiw2bH6dihL+wg6T5L//mDQ+McPHPf+oEpR1w/nt4ZSWH5vFLe94ggcAimEGQ
VkViRixogojS2jYwY411Cc60kZTqaXSYPZ26o6lnRTBKIPhmAqjhmk8SDq2n4OI8f5PC/D4Jdzk3
+/ASuk70vrXoyPUTIFwbuikoFMdmth8VwqQ/33WsX23KOSaToOc1eg2QKLV6ccCAso0twHsAB4Sx
DM19E0ffzButAwdhWp1PbbbIYpuFIMWVs2N71lghBZv+Mvf4KlUF5IZelT27hZsZljtr65zZTyy9
LuhZq+fJCQ3WDgCqcsvtfSlJz2yhxDjT6eOZTQHxrKEC+gYkz2SoqjmB/kz/1W+lE+uOzoMq/6u8
YCCXhJDDoWZNJMV5NNg2+AXedgXaN6YiEJKfFiS4IcRs0fP/a2jhthK5jKG6KNsceB3+QgWrtWJH
vZ7C9juLGluemctlEjZWW43Z7hc0tbtQWubHh8mPrr/Y1BdxgQ4SQ8Wu8pnjST7W3QDDuCjr6zDQ
J1BBEycjCheSBI2CS4LMbhRST7WlrBDXFlVQFICV0VgksinxoTeLEFGwWFTPWYRasY4VqhDyLBLN
xJylLozTw/fPBreznbd7NC6E/JEz5IFD5BElT+jH2gJVJ+KDlHhr+63fNf6IFBuVr2GJlW3qooQ4
h53PPIxIu/eEXNZ5/i0uue8idh7AlMpZeWdVLErQ+cOre/nRVgwiLFl8jFYVT/pfvGUYFSa4gvyB
0UQ1pTm9LnuUXuPfdFhT+SidpEcUCvKBp+xI++Ecwch6zcGyASN2Zrsdat8Oaah3Iv61p8p8hGI6
os9uuAU9J2Q0YxjEAXGSxyv0aIvmaxluFR++8ecHQy6JmkrnARf0gp/hC/3vMWhQIDIrlNXuQSIn
0kG7cfF4Yn1JmZqT8P2OY34yxrjdw/7vthHVGW1/edEdyxv894ST+tn+UbuBFF8jJeskf8Yjq4R6
hQsgxLPpgRZN2g2Fl4xuepI5FfHsZktp4FU43P5vi2fh1iwICORnyhXkOxboupD6wwAEngEf6aip
ut9/0d8jf9LEKpm0vsk1dLV9rK/RdRxQqDpulZJC34HwJVhvzCdHC633vhtNthaXXEWxmoaU4y5v
JaDt7wMMxn7qm1Pu477VtGi6sZJoHv/Rr/K3SAaP3lR/Fiy5fAqxqO9yki9cnjywFOSXflx1UYXg
Dky50F38Q1IL4hzl6qS6CZ4IiPyCp1WqgLVZipYcd40HT9owhG2TaBVfDMAXZoUbY9645Ki5kJ/x
Cd7Gwsr7jD1hWZCuif2MMiZExS29zLOU58xfYE2jxcx27dBQmmW7hd4ta6IYnoWTPC4gjuesDjMS
4RyzwhSBZaUjo/q8RWi90nB6B4LpJvahx/8ZbgkDcGcTtDUBPB/Yh49Cxe3xwl8ESpYevX35UmGT
CIEtvbztVkyZWd3QRpe4OXnSob50B93FpIVYK4cZa/xfCN4tnqUK+0EQzICuHY6o11/sH/fMFqla
huSLXVwE/kXZg9blri3d06zNY/sqFlbimWT9UbQSPYfsLoVz2A16dxF2fY3q2CkK6/wZw8jYXL+i
pjIo8RTbZ6bsS+GlMT8TODUsxJEpoNQWvlaK56bIBnBaWpT4c4CKTPBMI2jOrMGxa/xe66yM4Xso
mpL5BHPLFtgWlVXtKNnYnEa87djggIJQH3ra61kKuFkW5tvU/48uVxED6CTWjdstvB5hCBjFRo56
lFBC8v6NskoHp//9FtC4lVDGlyMhuG5Dlrfut+3qXJq+YrgKKgysqE8BLsg47ZVFpQKy38klsGzb
KBXgcHiuSshw+vYigJP8Xfjzt/w2nNf6AHo08TGy4cyR1shCxA7JSfNV1H1MvOtLVsFc9M0riNp9
Y54xeG7GQ45WptQWVfQPmPIXKpSWveV0SdXdubO1QN8oLvl3u+RkR5uY/RuwWy5l3EGLxYriDJR8
Uvtqsi5M6SS1uf2vw2AcfM1Xy0WDIEcS32sWW7SKcAOG+2m+f/9BoDeBnJx/8ysOTMMK51ea733J
At4pXmgXet+GXyTeGOb1VTjkC781kq84L5MiS85MTToJO6fZsMOdnxX7ziiX+TcMh/kCACSW0HCc
gnx4ocQWCmj+1qyyW/S5WjXMQLcx4t/URuBYUiW9ejgyuyqDp9q/xThlXu/dos3ryjY/6zNmJVxp
8T0MALNoJWtJG126uEreXQOh6e/n4JwTO/q0ZF4zUDs7PNZloKcKCexc/NKhuSMaLSRSiouIoHPK
40zzd21ZGvtTMKTHKxdXWDAiSMpqPeL6euM/0HljWSechX2kmO3ssWubNSagQbLR5wtqCfAOYkrp
087f4lfhQH17jWxbP22RquUB4Kif4xHzXBx3sYg9ol9W/SLWg2N1Kz5cFYEBSVwd05IEryx2477E
68IDCeabytyrd1bNKzpy6V1nJKP2W6Ix+LvHIwPPGw7+m+59+7bcaIWPENEJWkrW6SvAByU8YEWD
bca8jBT9NGsZFkXp5q3FoRpmcmuJDpJNAOjpO5BhMNLUNWZAdEDPhFie29dgOqtmyL5OD3RBmGnB
QwaeADO207AKag1CoGlEsGLzrYvTtw03COcblTcsGv+1d0SEPoJFw+8WVnyUwGbt7Z0PCu81iQfK
cZkNlrUQjM1rUepesBhZO0twXhdkcRsuZfJiwnhapSi2yF5HuKFOrm7BuHtdfeN4Ec8d2s6AJQZL
ivkcNNymsbUa4/TRXPlSuH3g0Gf/7R+DzYGSp8t6YnFEA0pRin7o7u985wqds7/MlOL4+GP4mRFi
4uDjXGq1SMN8bhopCnOROige0ckDiCH1LmNzWA4b5kc2DQImVMj4fFOc2lMtXeCt7EAODsKIVTy9
aPrK1f4YZZYYax6YhXy8ywUX1EwG7qtd6XVC3wc2hgcfXhq/IqQ/ZXtVGuh9IBRR3nvecXwNvPt0
MJZXSOReHcNbHFY2Y2+9Ce2sefM8TKCR2nE8oHYqVUNPRGXeCE0DKKHIHNSNvFVIE4CBASEFkzEA
aTg6GY1juf/Lqsdb0z+I+q+Y+7mKtBRGZnJR5/yWxfHOItU54tsHaiW/8mP2a77xERtC9E+7a3Pr
9TKYlYoT/ei2jG/WKc3ey79BMqJj/6tTSSu4ENavafY+EIZOOYF7+7bUWt+DTLSId70cpQQ2qb4i
9bFVojYDszi0XKclPd/+pm4O+DpdEv2ZSiW+pTuClSvoKiVs4X9lRucXZPAE57cYs7pHgG+NHOnr
xVqGax/bBdPIRX2EDiwKQ89MJb7ZygI9kdaasZZmGhLnf8zj0C3JzPErgujLZkOLO189x1fn+VvU
GqSaeikAMsq9zhRVW/B8RUwIDWruqcJtDUqdqqkgyEAa6V4kqo6bvVQ5DsshK0idCD2UyKiDmcie
eZATIl0w0Bro3cmdjGQ6zPteiR9O6C0q0pgjY/1qmP+GJompE88zbuWtmoSWACCaq14WD6okAOxf
rtzWg3n7LMS9UWwW36MM8UPMUPyi8b7igcoSMNBCkfyNwgEUjIEtoFJBcBRlpGmmPQCouMoANvkg
L6DYKgc61gNM5zAF+eZQx3kZj+3c+4yJHnH2YNRlI36bC3M3CUsyIHPohU3DiMnZw906zaXFx8MC
eUTEcRSfF9muA20tXv/ZmGr0ah07r4g+t4joQ3ypsJxkqqsH5pCVh4zywcaKb+1ca0jVGyRKXTdY
u44++mQwB6hJxim9UeeANJ4J2Pqn0eV/S2o2xzvFIEsZAsleujZ1+m5lflnOpl4UqNdjPZf09qta
8pENJ0KpIP2DXscAz7p6MLHXgpXdD6XJT3g2DIObrQwdZITJXQ3GnA6uC7Xx67G3RYwin33gd5BP
hueaHOFFYxjTNO4V/Od0y651wpdorq304PZsUcJdYLKyh5Oj/EBMxpP2ZKA7yzv1GtETKj3oYH4y
IgCe3fXKXpSUPuRWiIvRo+/Itqmo1rzQlwF4hb2tXy/qkwNqpgh3Ze4l6Aasr0ZbsI9tvSUBJh7c
g+QlCVpreIhsBk4WL+k1KrNXTJDlnilzxSMJizeLGPOTX9uQNtwF29O4d7lhN/oMXQgPfFl9m7q3
fQ/ZCHQv29u62rXp9FQphcI7JbnhnPh+bUfg1eP4MyBkYEwGDP0Vyd6PvyExK/X0zFnALYzQGvKi
LI/jPseKl2kV7Zw2i8lJrIurgSdmhqDLv5HfYEGonfi2Ih90jczTx9iF1cf7Aeo7I0TPJbZjzpqk
46mMBwu1dlDAmx4NO2Be5V9DvNGatAGfe2Qm84qj9l0Rp/1oWDAzKOft6+19q8pIFO58tZGKuLYd
tbV7NsEbqSfa2innk5aw9xnpnBm+5Z7v78FinHRkwIEvxkeGK/Oemu4dxl2f6fBZXZ3Bl91LFbmf
2jVUCSFheuJtbXKx46yS+6DKWRpHdrp4IbSpw9S8U6MDfLTwVFfcP4xdrxs8XwvnauMt/yq1hndR
5xp/9A0h8S8NNaCfIhAFU51cmCtkTpRjgnhBsDygP2jKqhGQPei9SCBQgeZkQXELwsMY4zTonfTx
AmSGdeOiAP8iZjoxif+3KTRd8N+UKRkYvyrFVzouj5tj91NykN8CEO6BDIX/aa/3hyG9BsqUPh97
BRX6Fj+5ski4s/RSle7+FIxNnnE2QCufVsUIZcssFH5d1cTKCyJevfxczx7zyijyEcmnUABImWXE
q3ZA2wdeJWMhrPwmWhoUZspvGti5imrnmsDwrKRIU4XK0ZY0BFk8x76ClBo1byn/TM+cC12MEtgR
D+Llhws2cDkUR2beo1wpBWjs2t7Kbj2hq0paLYlY0uJEOAF3neFqV6z9N3/mr2Hs7W9UYXmW7qIA
c+OBnhZhV3uJRC677NOM+5/PpdrdvEjh080qgYwwzNfAtPibbUcTVqOsibiZ5l0Be1tMGZOIvWGd
GTFCQFDR7s2NFN62sBh0mFxMjOSfzoAodZapKp/VDD/FHy4IJ2Uy6pQyxustd44eoCFpBZAqM5jF
EigM8ASefEAttUIIo0XGWUTLk4W9LCfBrh/lkM5d8RP23DBLrTZODiUGbpRhubxX8znK5ri7Ku/E
FWctRoezdfnztZ/rYP/DVy9Uqs+gL5qOdt2RF3lPNYx6PZeh1Owqw7/RPEmNkmGhj2wM8vSsxut9
LW5eHUH8eg0B1vYg7IdK93ScGWX5W+88J1HnV3aEdXXukrFv8u6ZByQ5sXLQxkIgchQUtMWZDJLA
GmXDNba7ncbbIaAjpBbpXLXzEyvaJ6ByHKKzFmCmEHoa02meJlQktnHi76tgX7iY8CKjj4owiF4W
eO6poNvbd21GPkY27fgkVE1VKL0Hd5EfwUjbQURIMuuKy07X6oyIESCe+1nlxnCGOF6Pq6GENQHA
Z0ZctQ5qxjlh/q0NrlHT6O/VtgcVbk+qlaupHz+pWcLruN4ly0s8fWyA0k+CbNkQG6h7LKSuM/Nb
Cj9ifwSBpnHXP3jsYZOo1x4cdyrawbXrzw5yW5K+n2wtHxq/j5L5q1UT5hH0k0qa4+dhMak1xbg2
gHukmOTo/eJhmU5YQTxNYd3RTON9HFGnfMoPCtZSaIuU0mZmDlbvUGyGvkkjoXTaUB3V6NEXPrQX
Vkh+BJWR6YZoE9zTuAk+kfpk1/vKEBEu7gwF/XLlVmdwpYYdU4o9QK06c7h14Rqf74SpBSK+iyUz
m2msJmaxTmWMDq2xto5GE/tjA6ojG9OiXOdJMRDWK/wUo/jkD1IiSCGL+ZQTuOIdravSoEDAaNap
E6BEQ4s9Lv/Jcg5OU+AkkxPCjcjNHUPNcvq+SdpONqMwoDz3s3/m90QwQqjiHL6plmkiboYsCtcw
RE8LsBFtsTuI5oHdgF5hQBpQACiPBysGa7MyvlaJYNgK+d0dwPofEDMI/MGMoZsyxWEpJpT8Fn98
xhvvq7iO7sk8iQEWPt8V2vBF2qrmeUFHAV7CfgsH5dK/X7cRXbg82SWCejBJo2agdhrDLJRXwaE/
Ol5KzjEkQDqylF1zi2XHES4KC94Rryo2dy19bmAS5uaWGTBxN/aD38luv3sjKhI3Ka1bHZLVvmfX
mIRAnPA3MsqWbBh0OZiUbAowvsQBLDALybQt9i+kgVVDwScQPNqVTl1w1KBluuqhKTSigiErV+A9
Luzz6XdX8U8jIxF4zEswVz/pKBjkqYidrroXoR3NXBp/80PO2VYrulSBsm6M3mimW3tiYoob2+pZ
nUDtE03mRTmLkdH+EAMqzvOVaO0GnISP0O35ktZrvAK0KofG4tmDO0tUI3xh98bFoIjourFeIIHH
ENT1mM31QHDlOMFIC0iFMaM2ucQP5cRtxESR9Wy+4WTyPxtB1/BrshY+eqrRw3DBZMxS4iqqtIV1
7IGwCR/uGShhg8VLRI2wBbBhZCJYx/CaIezxdubOoT24u1xUEQPY0MA/WMVFEyee8WJ/T3jg2Wkr
AP0Yc7P9Da/Y+OffX+vt9SL9fEXSEfn4ROAGOKgC8EBKUeoEOtwEctnpi6vB4jyGzq4gWV06lWE0
Q3jHC6eMk+XovJA3Wx8+SYlILOzVkpit39hF91YHNvB6tDxV+o8WrQPdCtGt4yGDQJS2xkmepmtX
ne7f/iM/N7Xi7lGZFNJzwcBx0YWM24L5bcIXLf0ENsvjpqeGEushu+FztULY/J8zXsADX2EuLAzD
0yXwJOvfUXtHoTFeIGAVmZl7Jcq1gYtSNOQu8BnWUYHC5nzg9UUyDK34XRzXB/yccGN/onvVyOSZ
3BYzf7Wruu6c4vPaXyp989l39UYskMF6P0lI04mSwqALZm3qyed9POoxWmvUcQqckDvS9o/WO4MN
VjvKpMKGRGfPyrLl9EBhI4MNFjMKP18ALXHxU+FUGFbmwN1DLGYRP+npobk32zdEqc+HJvz9TgRb
n/NBns3NQQwLHsyTMtr/y73Y9duPhhPEebRgRBOL6cNqkLWR1POZYQkHoh4HCbu9AKPxC19lrJxC
JAtEIDjvU9XbDCOFK9ZHs51VTo59p5iIDD5hPnSfU8XIqN5iE51ivKHD0yiXIufYUv4qvQXPXhU6
2FjD5+7RR9yMs1IEP8ebCZsL2IY2fT1neqA9NZQPUDDYkvyM4yO1/5Pi7+Kp7sAtXmB7TPPxdZ6a
e6jI5pmDaRnV63HNX2KBYR8cZrbrUU2FD4jBxKbwc5S2TDw4yf1hb+DgrxhE+KrE/kCEJ0ubDqjs
R0cUu/F5GS1sWMzmlvaawBUifUQrd3wFx3gn1/2u46ylK+8nGkFFXpCp20X3DKpBqeB9wMteCgBy
a5MCrY33vlk6rkcSW0Hyt5kXCaEfkcQQTtEv3xPwqOJL1NC+QB+gt2ppcZVhRAt5sbK0rh53Y0K/
3eqQoYqU9vtWbc+ctdC/a51wpK9ZmS3U1+ICSpmROGHlSYt26UBmvCzJsjfxHkVoP5efCJF2CQy2
0lFI23CTOQXlUN1iAJPazO0w3w+vu61iXO9HUW3INDx3w0Hdm1vGiawBgrvMVVXhvqKDbzDUXcyN
4SGfdKYnCBAEwSQw7a6OaC0q1Tk/+F71T3fBIBJPcTkQZYJBP30Z3DJPOL9eTustoFOy4O44sCKX
yr+umY8yfcy9gmslPMoRfL0RHfq7Fo0+mLg/CnL+mY6wnmhRJDB50dcNwO/YuVVPRahuEK12yBIG
8IdPBBeYjJLi8w8drltd8y0cbRGoD1VV/2OQunRytsUKnVo+WIvttVJTgciC+IKM7WZCkDzrPNvS
W3Tur5YL5s6kYc4pub0Vfa2Obzi06UC2E4yhNfTxpFb4uA5ZfBpRH6ibt5jB+yrG8cMxh1KN+fy9
Ce110E3vp4uC1jxMI6e1Dmu2/OLiGgCUODnSionRWNjtdxljjB1gTQs3N4ROqp/Se/hozY344Rct
eztbIluo+nQlogaTj/uldXP1PN7QuzJtImoOiaHuGjQODTL9H4MWBY/aLEAx0gDOXdKDEoblvb9X
O/W6yNuoVzAGGkzO5mvu97VGMqCZ/dFcqoRzgs23HNtUNF5BwJpXHL+Qqm4TPJwPzM8ncHgDIPUe
XEF72k3ka7tj0C48sifEOJWphKrBg3b/qanoTI37lNmWyeSDxMGZjJqYWLp1M0BGpMg4s4Cadsc1
pdq+Rna5eNICpuw8zrwaxJl8yHBzzUGh9czwiIL54OUYsLlGno2b5FY4DrUP5OXl140lrzm+HBo2
MpXFc/Bfc7rXWxS+p3IKy0puhnYl69qYVLFXThWM9zPBUbtWj4Aea0BstcWaOCGpYFSz+KqfBqj/
fYDMa93X/PBVwh0gb5K8QWdHZefz450kUoeSkiFkI1GsluA20mY5wfQVPTIYN4tT3smaP9J33uGD
eIlZqU1L8kDNekZMhCl32ZUMNU63Ah+KeXY70KgOeFGo3ojcEUPB05O8PSyvYpN5DuAb25cAI6gF
tTwH4IYqUxz7G5It36QA9Z/A4fIz8DniR2EaqY0CLc/pUaGLQpsCvj80Z8dLTejseNp2+CuVTaDc
so1YE+9yCCenZBzp4l/mn5UxlV/gm5Ks9HiPiWj6PlLyxI9JNKz0qcfH2dakU1PdIJJkRoq3IxRe
cnJjXjHsb1FDnxwV4u4K9uSL+QLlfX0uL/m3/aLZlckFN8SVUlApIUZozDrmpWsCqX2Z4lsk83Lp
vhCi3ttLm75vnarSHAUrfU0KeIjyBKXJV/B15Y6yhVLbL5RGe8dBSjVEJWkGCXLHA7sdLw/4LpYV
Y1Vg6VbwbnjVgNTR+alfqrV9fJD9r87+kLlGgbiZQSw6wgnj/Ykvpaxz31EXSivDnOD8wgtmZY0W
OAwUgQ+XCurYioqIqIka86kyIR03eQNX//QkWBbRWT3wBSxTpW1X3px7ga92LebQ+Hsjik1tKU0A
EkzZgJz5yWK/3LqPt979qkR90+RnMUYRQGU818rUcGs/u9DgZ5rgoLM9jBBplSrtEkHMOjP2sVMN
3/Np3ucX9x0dQTZz2XRFCv1zBZGrJmPPT2Bb/top9Lx+6WJzLifx1+qqDTdqfUusWwwWxeXFlhWn
0X2vBQGUtmbYiAaVlqtApP7g0WQNvZ+p7+OE1b3wiwiw2lwgqtL1Sqs8P2jV+LHu9/JP2L631/gQ
IgYi+1nVVkAk/rL8ZTPZx1jn0GPAjwvPi6vIzrEwWqvY7YgohKP/+1lADcpOdWbCkCgZUiPqYj7G
S/0xE1GTwqGkrxg9wEXdfCt+OPqG4rOSGMbN0uafXR66ErChUwZNquvaST/J+0IF5nFny+fqvYsV
4nqjJF3dpT00YEeFwNf2x9HHXamTUSsZLYN0+v3k6C6VUcoMGJFD1unsaNUSAC8irM2pmzw3teFM
xDYo0OBS9Vhqx6QUzXOyopotcvqgeSZ7BqluEZDZ2Z7dGGQ05UUMnmMGxqAMGk5jrlFFxmbHQgeK
Y9Ceaxt+JcoC7nmaAN2DqwlE0Sw7wJ3CyOfGFnLv0zcejWeiLNeHgO4if5vLU7rPVm3o3fke39qo
j//xFXuyrkyOjLYagJ4qDGrYfsiGJn0FvKBqpT/T95lHv5pNEtji0xr8Gfs/kGkNsYfdTXrA6sSq
EpBROqLrMzUtlchSMr1f6F0v0td6TOv0T06ncSK1PB+uNKbmGm0YeC3yW2/0sKJN+g/70ZOsjcBa
ZR9vQjPTNcmq5okUUp82WUOxaJXBHBtCV+NqIIv1D/ojjm0QQnpSc1yWleVyDLzjIx6FTUKdOsNY
gkZde6vFt8psaQVhzGpUMfPGIcUVcqsuaD8q2CcgBJdj1X/9bqZ12y94jxxepLVAzoTxi2GJN0qv
ipNEIFGGBXiHvOke2VJzryMbUmCx+dYB3EIkHWvj5DSgHIwriw2XdLLrPi5A60rJ88MHL57GpM46
GeWjYLso17KlDplFiENFiNmDSccg8hpndXXKsp6u6dm4x8/y9ve5WDidYa5OmEWDLrN0LHJE2Rcg
qjPY2sngqqGFm5HsetX84ApX9BZwK8LpEreP3+dTYGhYJy90uDD5dX2xCwNc6ZCFJhTJtpYOJdkX
uK6YAk9lQpg3O098RoSBXuyj8d4soIPbX8MAyQr0yrQNTIWYSzqxvLEg5JLyDq2ukW0tYYcB6UHI
GwY3jUkS9g4yMCSsO56dxcqc2hH1CzuIAFAV+i97wa9C+bKggu/pSzcHSWVITEAzCnqKXtiDXSI5
5gqNtW82SB3MiIn/m8Nq52P/QfN5bfy9d4GIfuSnfkpO7KII/DNHX8MB+PErGsqwzIfHksGwcq2T
zIU0RzrK+dAirrtmllpCkpVC18AMQFvWG1yNe2gJTDu8GKrdCRPt4YG6W/2R2PacTm61kEAWqGvx
6iQab0x3Y22rJWeW7xN9vlWHfxpK1BgJ+lpipBNamHENgOXEO6JukIkQzHPHr3YDNzyiDoLUo+Rp
uGBFaXKcqzYBFWhRQbyH3Dv46Ipoq5UkDjF1cj+poiYAmTL6IUxGzqMZ5MXT101n6hm0LrlZF7YJ
3SV4eVms91FDSRUmQEElfMoPf9T7zYQpS1gD00/ru9zq3pxMLY3fEPMdv2AK36OkuLiyU/ctDaNe
4+VbV9irfX5rbBe/y2wahK6QQz3DBBmc7490eNKiR7M8xG1+PIzjdzZT3DuHTmnq7okr7uSJPPtO
agoWOiu4Bz8qh6E5gqy2+g3t/2hBvjiIHciQgsCbwFJP8adLnRSLObxeGpQFfYMVDUGI28KUQ+i/
pm1W5XoXPxdhzZ2OYXK23T4lKupvN0RXNBMK/+AZ7CryE4fd2YbCLH/Abb/BQgb6AGID2DwWKkci
NDnRYs1zrwZ6d4ch2SSqvjQQCfDGvnhBUoULYpiPeTCDs/ijMm0dVDHGSKgFgNSRBdLOedcUvFf9
k1AldxAu+/3h1XyjGCQXkBh62lLB0GeptcN6tfK+OMt5QS9F1mqiziYkeG0RIFVZW/1cTxwUtou3
stI/GTCabQwfW4+arnpcHBYSh5ZBZo6Dgq7V+MZqI9/UeOSS1CK6pczvESfXoRVhrbeLOB+gcbK/
4ap1sb8Qr/0Vt/OyoVkQbQI1CAVsW7eHf2LyNNrAC6cN9b6MjtD4kWdO0r9ZZ9WNqnclk8SGdmlV
tYWRGVlcdnCth+7igdxPCWPdvDkug2Xhu9qsRj+Iua2Y0j6vUlXElb2GCCnQv4YR7lNrpWYvE/rG
bj8ElnpO/02btIbqrRHFrxWpNqZm2I1hXw46CvAxF04NwsXci64qdns14CFRpsem8eFdMwIGUwsj
DzSmspVjIiKZ4d9R2hhJUoiNWl/bK3Y2X+oLEFNee8jZDV3ywiSvptt8MtVMmIXnryL97xdy6Hr0
TBHk9gZo36UiyB1MyjN6azjMecU4JQPzR7ZewgtA52QWtKLYJ3koFH5yw/k8Vo2SzuT1jHpQsVkn
5vwBDGvcWYUlLlI1PRmeoRCx9MDmrE4fnSiXOkDu36aqvMulB9GdeLcAcqkWVctftK2vnJz5EM2Z
3g04EM3VCxGJb5KN8OeRKOGHNW4CTHgeW5CHO8vGvUJ6Eq9eAKYVyr/cbLsjba+Kk5bXK3wUqYZa
TB1XyDHuGt07qJ8TrUgIb19wXLhzA9egybmd6DtJacVpxbSvSWFE+WuQixeP3AHgfKIdtG6Yw3MZ
FYfRo2MxvEdtk+x7zHwrlA+HVttYrQPGMx/H0WSuHY1xqnugLN3SiH/d2YxHkN/nI2v/6xxWbb3J
B4Kd5oVuKDzGEKucXr6COroXzrm3G16sAC+O9UMV3L9rdoarPlPaFNY0lg7+lhvEMiRV+PEnN08Q
NIikrrTAu1ShOK9x5kJw6wJC80Wj4dx/tX7de0ROgDem+g6Ch9i5+FqDv0nczif7EfN1dF9euQhW
mkSobqsA6wFCkfCzo5sX6emBMUihQ4ATUm2C7wV1i/zctdryMsow38OyN9npg+IPHEUN2sUKYlwz
SLQM18nLZCzx+eWC4I6o2N5z5PPtyloUOmDmXjwsL1Z21Hdh8yrIV1YycaK7KHLg2Dm41IC3IDPr
7q4Wz1M4U04qThxVt8mtwLx2UeCCUwRNeer/x4ofhIBxN+7klXTei71u6gLsjIyGgFYP0o+LfeVd
0sbT3QaZIZlcGj8IY/8QsPCqkhEayY10TYluAYD8OzBJTvFt9BEJo8iBCQN1uafqWXa1JSajrNaT
Hlpgc4v69cV8AmseQvTRp3oaXqa4mZgAyGTDW8itID+sNMmBCTQD1XxnmZXACtIeJjOuWc3JcnLR
y7NYYLzzsVVNeZGBtx2dX2HSndmrnzIAVKWtVOZ3ZcwiVk5AGqCC1Z5HQ/P2wzP4nYBVbWxmTQa1
pnvMXVMLAa5AszHQNkNU6To1G34x0GKLhnQlpqDG/IQmBaQt0uFfMd3tM6MfT/65TlJIcA3Khq7O
jjOWIIuFl2yGhydwjaOiMsAiUxWfV5gZXE1WbwuqlPFWML3sxeogKgI1TxoKN/xOK1Aj2QzzOWJy
15SnxL09q5lsDe+mN+dQDjuE4AFpfuSo/Lq4CcO8VfrYgQa1Jd1AwkUp9O1DBevYnmutU7geSHiH
ynwgywAC56GLOdDNLfRj7QuyL53RRiK31A1p96CTUtSqe9T0jAbCkSO3y325YcAKKDuzejy4bygV
Nbj3fbIOS0e3X/rcmEuGEYT3KgoJEHVJqVhswfugi0y5blGhzoKqnuzsSAPY9+/GwQQ4EGRk1iLL
k6SVTJbUdhzjEurS61nWaOZPav3ym55A5N05aEyfO7SRzCsxZ+JajEXXLOEd3EyvPRWKas491GhJ
MU0DC7Qwy4q34DJuwonjQMlwfLYTleWI0YsrkHrxjrVBwG9MJ0TwFW5EjiG/J2hotqrMZKNWPq1N
UxKhnGEIZgSHq7Mt7p+tgealcjVaPrfdnTP4rNlm2dKDfLAGU2mQe41NfG3jvPF3zB3HYyiC5uMz
PTVugy6G5UZq8vbYhsvMcEelREfpxCJy/JPxgYmkJDLR/7c7O3fs7NENW8t33lj9UHTSXjWxRNT/
WmzwmKdyzLcf4Hlgetq+ySLkq1j2MQpOwSYw3Gr+r6Qhc0laaNfzg+fW/O4/Myryp6gT5ld/jHD7
B7xio++a7gpYnBY08IHtGWT/jbA4hEXff31Hb/5jYMR5ZJDlrzlssknCNI/LO6inhGxUJ8Hd+eu0
jv60YlYZdd0BHye10dQx6gCSJOtoGqTKxK/bA3k3zQOMifN9b6fAzS6Lj6DQDMU7jsupC4gx3UDC
8hplEf79XViW7z/T6B1r3CjI0fyVrp8cZaXliDLXJokMJ5cC1Jihx73uXSdOd/k72LE1S2I2kYps
Q0t1W4k4KcSS6U6uudsJx+KmyYb3DWtJ00HIKPcpOja1UP4FVW0P9juvuqbx77J2q2cWRGYO0/EH
5EVb1TYp7Q83FaOaL77LvS9FZ3ojYyZiRpqtuE48QuSbOTBytA5ZvrmKOwV21qcvf9vDnaci6OHM
vPeIBOZm3JsrIXmIT7boUJrxSiHcwx8WIrd+U+ZLRdbMseZddw6QCBh/l4IMsOdOH2b1ycZyT2ug
gP2On+Kag6GLHb37LKeDwsjIgrDvGlJx9lSYHNgJrFFXJPDVNOAT0SWd66qp9VFaolRZhm742gAC
T2JizWdhsFU6phnWX7p1vKDmBJuBoLcHpvbkFg8oMxuZsNHqOubHlvDx6bqwIUf7YANjmkhwU/vM
KsMIkjkoJnm5CFSdzknGsuM07bjY/OxB9RmlTDUVXtpeNQAas3FNNQ2owLIbEOGxySUlKfyaTeZw
8ziJMkyK6LKXqPO6DCwew0zjRSWDy5XBG0p3xZ/qz6NhH5RXuKmeZDmRpgNKbp/Kj0uN4Ylv0JPd
8QawU/OiUavWh7l5WQw6DHRkab0xm/fhqLTmkqN0aqs/gFs1KqTnYcNDtBgAxzKSNrEia6w6PfOH
uu9gy6HgcToYxd9JOpGD7GxIyY0AogtT9Epc4FfDuR6WT//7l2ZFYVM8R1aXEUr6uztbxZx0tZJ0
3EWpOcZ4EfS5ZKAWw9Ukjx/y7EYZf0M8HOt9/ZVN/ImF71KF4cxBmj6olsPg1Wfj+xzTnLA0BkDT
2tf4RMEOVAWjOLorp6op+VlJC9IiFWQlvi5npgOspPKaZB/epCsbPtnaeUlUQskkKzyGsT6sCndq
sJ8Og12kPLJ1bpniXRaBhhJR6rDamJD+gvRXj+xb2e4TODXC9FycP2fWAbHqF/2lr1T16UuOzu6f
YLRweRfq9ScQX35XiUaAi3JLio7iwJVh1zjNOrh1Ka9jA9LZLhTb+SY1MyfMame7fLiinKT0ihsg
VLK8ogjHhrz/q9QSHKnrmNcoDtT4tZauPxIYlpyMoMzclL+O2UlTTbZBZoENEgh0Lq/Rc8Caonb8
F4gtW3Axlng1FYV2PPkLXj07/onU9IGsladyPu1oPCCfVzWSr0CNgn56oVZjPfnAFh0RKixHpzxH
s76hTtOTYxFde0W2NWiXmob/AR9uxqAviCxAW7dLuX1CiAfrana7pm+HtvIBk1TDIVL6kWEwqbiq
hxLceXLxIxWdrtlKiq98NiF53E5s7Sw4QNlTcSX87ZgZ7uvCW5pHdRfStOay5rp4K4L1MOp3+v/t
J9RnqNXt1D+Jv6sQvbvvXNCY5C2jb+Ge24lUVeIKYwVUwRwLTYHI13SeKvtpXDbkiV0936IHzX2r
0QYxuPtiU53T2WXF/xFXXuogN1XhaXFuuO5w9bQ7rIEbTJoc0n4fRV32MbV2doKgkkq4iTUC/okU
z6wRzHfvzf7LDYmvEA/irUGmcbkQ0ZKajeEFRS8ebrxm/KbJkkatQDNWLah8HzbHCFQP1MsxNHTv
Jo5EVwFbAxZSOhpMmi0qL14NwI9AhtYSgCBEk8BjDbeLqTbibj51v0jRs+mKdoJ/pQ/VOI95brBI
qgycZXImTbWP3hcnnfmkFp6EleZiNtnZg/WvRdxY1ZRr1TpPPrM8EDS8hc5TxXovJTekphjdZoFH
2MvowLSZFTBsi6VNbJdi74fvIaqLDAUZxMPuiEU34ps7/4/i11ciXsoUoawjXscGaWtnKmn7qsSA
AhNtAJrODVkIzWwwQ5E5hTJh6aB/kiQO+NN+eDESHBFZTYoV7TNMjLxavGT8sugMSxLIcjf1QCQB
8J5YRT1YTiHFyC/0R+vyOL+FQs0hv9ZZfDUV+EQDffVg2VsPJ/etDDMBYuQ97NcvvAc3cS/KMZRc
7IKoMGPUfD7NYMchZkqRBfY9+/A3I4COdUZSb0NTB+zWzGwt9xdJM4/zr/Ec6AcsVLyITs8YXZJ3
bVsuG1D1tl/a6USU+BDcp1Dp76xpOloeL64a4+ntjUTR3m1nRAMsw9jIu914I3VzcOtEoKRNcVC7
JjT7A7lvhbjVxQZu+URuiBM9px1EfzpPC4vcALf/E7+ljrGL4kW1ks76qWjAusvaJ5J/zOeasKjW
qE1moJ94tUF7fVKUhJLKYMgvMO0ueqAwgEM1WnH8Y40ifKaKcYT180Tp7acSoF4tHw2zhtHRmFP1
5lWGI0L+D6LwVq+lAWxtXsIakifF03tXqSQox0xhqS7F/LPHKhasp+ZQbWDUbRXG6gdLH2R5gTws
/AvpgC3urT5l3ZoZyIPCK6GLf7fpyxZIvvPxtLFXUOueMQ+uLR2O7feTEaVWub87GcdAbAGFTPST
qFGN59kLjeQCxCAWqsAX742JgspgrNX5+Mh75mQQBziUXDfSI/wMW2xdIU6MNO3gRIkDvuX11ZI7
B8lbvW3q2YMQWPLi6bk2zYdhV/1SAswhd8WI7xk8i4za6gCLMdYhSKzyeROTom3Pk2Osj6jcc1py
J0YgNMwnKZng58rDZQ7T3yQpJZSd/tOLAyK3GdQeFx/VdJuogzkCHHyVbubjk/0kAUIR25w7gkMh
2etwXu9mrKo8xoppb1LDlCXuBcS/f2KU8Bn162eeFwPQ+NadIwI/QzqZ7yiBkiV7gT1ks1fFa1zo
GAGPeSv2LbRQxrB3vF4b34fPJEJ1OY1AUIgMnp1gBNs9YwKCsZYZL9OLT6Tc6RxURwvH32IDqK3/
/BKZPQAAWf2dAxIZpfnOO5WBlXYHGv+mD9+quybRdish6f/io0NzIQo9wZkf4iaHx2vUKholOd1l
QZ+nXTXPepagcQojkiAFMwjA3zrN+LVCH6fdzwE2qulzR6J8CaaPQ6ki/+h7BtPSg66wxOzcn+cG
G2xHiWv1GmGNM0O9L+od0BRNpXl2koHdSThX3FzlYk507etW2LeQZ+XTog5NMAoHHDU1nJew2dGI
fUScVhM8y02QaRmq5VKF3mAYbDRQUT7BvYSy8dPDoGK3ZuyzYoOBBpgoAeiy8f6tdbghr4EzmiBB
SertolnIo1gACxRQ1iYdoF8IyqsqMWc31HEONl3ZHYDvF0PJALLT+fXUHR8aECQn6ql73AT3asMv
5bhRqQ4LQmsN/h38BynQihNq42YyhW3FLe9vq3n7LNUVtfmybto+lp/gVuQ7SAWdEUj8HynAiqGk
9dZKJ4AcyYjO8/bFtLzzZ4fLlFbowZhC4v2QQ2mN/rmwxarFJt6oRz0kxJEt51wXdemlDN63NZOb
NTziIpjq/bTWSRjHA2sO/diGtwW6XMylHykwBQJDOvgSWsRlxs6SOLdoiZwAEpufDogEX71e6lj3
x19vwV6jGLYXH2rKe8MAhjF4P4BLCgxgHw9sUGl0BtSfSk1RbFf5c7PAOuUjvC8B55M4nBpzlQnl
mXPbkxachB2vDilOiSkQiFKPRbAVeaHAnV0dgg+ZZmLRgPvIfCq0kdNvelcDQUvET0AivwIGzibr
Hi7OGntfctzgd5X+99nMnd2mTRQNr7w+4WCEabCXc9+c0XXARePY2TpiVH+OlNxd1u3NPUXjVdEY
8JFjZOoEExFH1EecsLHBZWusOQOSwwLqQFfQ3ZaDcfgM5Auo2gOhyLu3COdX4FsPD9JxOae7T1P1
3PXWqTVxWUD1peagRAtNdssEQsoESb7yb+OGJoGFS+3rW05SxqGJ3L7DB79sECxcHoEGp/bITSuU
E2rXZTl+QlfIEYxpowd/LGBgFVMsm3j+aZXmXW59PGk1EBI7lYqxgOmTyCj84MW93MJ9iYldblgn
G4a7fPnjoegd6NxnboWvQpyFD8TkK9hTh1wb0tP2AHV5fw2B82PRNbZRi9UQxsyqfK1x9vKdQ2GS
WyZq9uZ7aAgjESlWIdEm+GWG6JdyuJxA//uTA1ibKgO+A0+bBlT+6zKQ2UbRPMaw6J+VntJDcDzd
TjJkQV4en/Yc80+JdqsMzxZNqMiyVyBcJARCUi2bn/c9TzwmAP/NIG+F1/J6tHCTJPVS3iD+NRFS
6OYR3r33ZHbYDymEjrMJIFCRa8Lj2QVhLApNJMw9WgRxgWO41pkN8oaxftb4DwgUhZ6C9Obbi3ts
CF7UDmTCWHPpzy4Lh+0t/lBqqmr1AqtDevaW9Dh6X8V+FBEprAYmYHZbPJxIcOGIw1+cRjyysp0D
4cjxrxuy/WaNSB3eE6UGybh5joUWMSWe1gaVfc6HQCqtVIFG2cwSYZefgXqkEBFyTIF0Uc032W7/
FbjzRGZhRVmNko8QKp6vv4RzXzZ9fc7Adsfo8MV6aE6OqZ8m7S9f0RQh35zb6sBbYdOSuvdgN0ok
OkYPAt4UOhrnG5XdgsM7eIMZJd4xKNdCBPnKipM+L7jdmsVS9JxDjOcRiDNt05krRYfROWjhp6mC
UMyJW5vlDjB8oszNmmPfJOIdwOkLot6e4oKO5FM5HJROfwVgUFfZFPIuAfAJstCqNHPTkkEf8ehL
q4EFZtiV2YI7ga0PkDf8980hfVRSITyreWUEphyBFamxJrFDUykMjwzoPpwm4LTtcjgRtKIDd9gn
m5a7ZfavIIAm/Fe0wx/0EMSK+2KKW36vTVdAmLgOyrkqigoFivv9z4OiefZWfwK6iPOK6dyTLkCb
cgqkh6vQhDG02DV2SXzDID4Y5+NhJwxNgU1Vd26heAdzbEFQZ8s60P+iAB/SZSEyJ8dmEvcnb5Mo
QAjhATD8ZY+OJEyX6Z0AKnETZfzjTaM4rZ4xANydJE+1dSIvF4R5WihZTuVF4LkB+RngDev66O9T
AHoHnTUiRC/x6eyXx07VJfveGnLoIL6ZcHNUtI+s54R+BUgaKFIv1VDl3HsQlcAw1DiPGrVpiT32
i/hEh6PBPYGhMdPGof1dw/wwa70fhe24BIuPsI6FV2ZlZtpfDRiAVDbuZTho5Awb+FLQZWhAtlGr
Cqm63mQqIwRTHJeLKl0GFSkb7wkPz2mfNIVvRxFwQGWpg7Wdhr8SajYBvy1gCQYa1KrBbhvX6xZz
CoHBNRoES+M0pp66KNbGPh6Y1NDsb5yNL1l0YY83D9W9WBJ4jI5kvoC10Z+CIxvenfxsZ1LVYzL2
+vk6/SIDzXQtd8IrMJkg+2Be51kMguMRumm8BaOX4q5vwObWFkyEs52lE0uaPXVIkODTmWA7rbnE
3Hi7JcHffbf+aSK10/jf8cjBbrh0nmrtSuTW6KwyLPafc5+xoKWhSFYJYIqQf00RlOkFnkix5Qzq
l/kVBFy60rp2kUTYske0NCImSCsuIqbYPJy46fJFnUesBvDM+o2oIiS3AByCSPUDy14kdmQcd7/r
P5TB14WHKRUK/VtIm/UemZvkDZRUH5IAOp547kDt3q7eKkY6d0+y0GJprvr/jtCZbLEjQgneJr+D
YOFdb8nm+wXpPptBGD7mfQMNMMEQyWoIUMFprZ6PFyatZIv/zHfMCVshCwhdfu3pg5FABg9StQ1p
fb0aK2YqINLDc8FWzRELjZKt84d1Pv3ThSAj66xaKoQ+o0eEtmh2XHiWIo1IYnrOmGtpWztk3gIK
WfTPkACgE2sljZYE1gJl2NPIn7n3S0FFV1g74a0UkzlFRu/7YI3LOlvhteDs9EtRSWDuOCYDRyLo
6fF6o//A6MmQz3QnCDFMv7YQD8kAVxxngZ3pnqRn7x3R7B+0FdPWp1CFKSG+4/1RqMMmOhnq8Bm3
dYpggXWHhPfNiGZ3nobAzTn8+mMX03JuHNj/K/3WLwNLfCqC43OXNOzRfK9xv5vXznZkysTYKRcM
jcZ3OeuIPNoENkKAxBSyKXitGHYyKNh6BlTZPeSVCAEw9eVomfC5sUHboz7xoE+hbhKX4b0twunw
lhdtGRqdXVFZ7ztbhzChqnwW3BJ18kucXWqKdRnfF3biRsCEzT/yEMxfHwiyR7O6rY2pZvAGoXyH
KQwFdHXFflq1LLwZ0eHvQsH85uHq3vgdrtd68dMG9HRgXuxX4q1jQfZDgKCKXzMMQvZQnvPaGAf4
Jfmp1hlynCJwhFQpzZ2e+E8eiGpKVtO9GwUoeBYlHYG+sVnBhtUPVnGePvARSWFAbX3ZcOghzsYu
c5LPYRthKMhI/YAyolMAoxKuTOF3b7LLBjUfkoZafmMOLAoUcSh8QI78O7MsR6HJO3SkoupPl0Yv
2t80ruylEtJ312eQSu/AEfNKVMo4yG+4WAHapZ0TZQAraxZY47XJYTmmJHNNE4nS5HK9ovIv/NEG
6LahszF1AEsmteN3Lg+mnGnVo7xDGq4tapSvWJDDP1xcuGmT2n6Vn4n/4IpsdusCm3Y3ivs7Qd1N
me4k/9wDk5F+uWVItQ8BWTbDeT7nCjqoXHWRKWD9uN3o43FL4G9So90IgCx3t67DRYFHK8hYDnF7
VoRwkCbDVVgqopfpIjEJvJpHqIuSc/vDyiUahmgBw6FPjZy2nDOBUdaj9kSMgMRSObUeVNLsBcV5
BGpNUdAmsyFV6KhTf1hckHT3q4xP/De7lljylKDw1T4ZzmILtkCffjqjFE/do+iD9elq9e1gLpS9
xobDVTvgXFwrbgsVZT4ikMH5gJWO3ywbyKOeZqPUubnv++357ZSv8tGI9fAQOtST2uMSo0H2MAZv
WV4XZprKxi7iyc9nljdFYmae+xu/IjhyWggcm1NTPaUSch9PEO+AdLUP+bUtaA13BAWHXegQ6Q4E
vVyhdcftPGdla77VONdF6ChfAK1Iuxxf0EzOJp5yV6BneQ3jJTF+Yr38vcK1Ho7EX9K/OF6snjd7
/RUeyRI8ujPFnVrZiwhoAbGiEd/B3W2hFFWZi8UHBZR3JUrKdWq9Nwf9tAG4luXnbf7eWKjeBBgT
0QvppIJZgsAec4D1vrEWW6JZ2BCmk9BvIdTgZMvsdnlPVjA6zFF8gZ+LYNdm7Cd58fG0Aa6ZnWex
XK5LhDmjSZWJzFlcrUWEgl94ZnlOtRTRVytV8t3Cj/BMu2IKOwblm/dv6bmbsGHRhDed7y2Mfu71
dMyn1dWQ2sJ4osYbfWdV+p4NoLryKY6h8K9ggz5/WfGcahCV7PpodSE1vdbxImIi1uSZEwYuoEoJ
stBii3hiX6wgaB0LI0GcnW6t8YPi4KQFht6p+r/6QyMbEnIimfc/A0kP+Olv/VN9h/05EoMEYXAE
dSUIasIllXuIjVKNl5LfGgl924Hhb+fYAvf2ykjT9h7nenWwT2Qvzxqt/lVm0h0W5SGi4jCsrhaX
fh8OFU6/E5OGWrRIQWoAiUqwPrPF69TDF4QxwXDdTPRbQ6Ep2I5ukefogwh6QuGPG1pSqFFo9Ml/
OwYUJCbIcNgFO/HfcbxnnDdVV4pM6w1+t8yxmfLJiKZhjgp2MOoUSaBto1+1zno5lGOlFWeVtYDr
ZlTb3CUKLMQzFf0OUkSXhnRFt90RZc5pQcixaVeHFrxw6wg2cUfNLy/TqBdViJzdkgWBgLoKuO3n
MsoL39iO85a3E/C0lhDNnhCzi2vOLCYkEtG6Jj4sMkK2EQ7xvY4hAX3WEIh7fPaQN+mUVPuvzjLl
LWkVZiqoXXtMZ++jUpHn+F9e3OVKnZJfoiTmzhYWfUfpEzUsX27nGRbrnqQFhh2+rx3p+CMZGGQL
TnQQe1YefmxOcgfkiNAlVsN9VCa1B77xQ2luVyfFKgzXg6o6f8JjJJCfP7rZejDjuymlGx5Z5cOG
bsTVtgkR7/abcjroWME1Oxg5s2VrIf5w1oTGqNv364XIX2VCD6gaV9luv5vFQQVfxnzIXB2yqCTt
4yTG7cnoUBJsun2jvnd0Ba13fLmRLJyh8Hbl+mzZv3aQWQXrF0YQowJ0hoOX+W4lMvEAWm5TcjT+
fHLom8qYiKdynsh7JFZouWgVLxpL1VOLng5i3cJxOblYA405qXF/S6ESp9jR/BvUeEiLFJUUGsD/
K0wdtDyG9thDi0ly8bl+wmcbuS3kRVnT+IQuyDyMY85fG8DxnGMriVcqZCaz86UM5rhEcL+MmY4C
tisX+EvYF7l4LoyL6yohB2Tj+IUuavGkVDoq+WF2CAqiT/22No6+8CKj02iTDljZf/hMJ5eha/h7
5tvc1ujjisO9YtF8xLEpMj9Hsehs9ty3DmRdYyf4EaTGJXkbxMLGqp/Hwv96uSdyA73Blm120h8G
AVNC304Nu4/mbyxrgdl5+KCjWZDzc/4mjN7dSKjAuhlN+tDSA4eQhsCIE3SCNbhYnlLSHHy6tXoc
DZY4ldvMfwq8xMr2RvrfuITuJcx1WmVOmCvnRU+AFnumW0X06WZ9Buoo77V4z97rUcxdzZg1MH1p
VTriZuj3hLmjzA73bP1+ICWYvm5roV33GHVGAawSuPbss0JpExrdNYsc19Mvl9aRn82A8uneI0s4
5bF620mSeX6cORTFKLzzupw8r5LAtv3aSnd8YQiVI/0nrWx7SobQH1VBvnhVM0ECXBPncb7Ozs+t
b1LdgE/dHf+uIRI6RsHt6pfm/Q/AcFTF1qCiq66mOZWZ8ki+BvR8AZPgQZJllIVGpJPzf7MSgaFQ
wdm7+r7W2r8sy9S60ALh9oTHR8SEZhMug4YsiFCXFZ9BJIpC29hWRIGaRJ2CdrTl0Iv0obNJxIFH
JLJTEowfN9yZ0DvGSZvnx17fWEdB2QGBh9V85GoEsqweLw/wMgmZ3xGvjw8nP4xVvVdPdqw4kja6
Oc43dqTtpFrWqRU072X1vphfs51VRqo9hIMfnFEmaDgbDSQ255B452u/KhtHQ4MsRlDite7+An9S
ZwtHrgNPyCCDZ6FNYVVzwycWfnD8GbODhNfwArh1yf4Ww4YhQHdQUZGO9j1wmID0uQ48WgDhMV8Q
ku02L88XLcsxhwrc4n4l3IdX7mGzDfiE8qsrsTJozezJCbgJTANPvy0R1Dr/3DitdCudhLMr8wDH
tsJM2vu2zncPqYWCMoZ4IZ8dVTBkKnC/4uJMWlWPYSTs6UXSLgLTvzDQnK0JAkq8A3peF15Ngb89
hXz9gtdl9uEgKVrK9BmSlsC6lGYJrv+7mM8aQRP3WKvZgmCiABNaOXI0hsEpGhIixYytllKCq9+B
S+OolW6ufOQohGVVxgFJuRMGN9maqVCTn6vHa+bZ8ls31DzWU3XbZp2vtljIR4lfiwIKt4X8bxRs
UhAMrN+BCkhyyjiKvXn96D6rSZTnXgEp7d1f6l0X13gRFZ35cn3mthwdcZq8WIW7w6Sx2zRtwRrt
l4fQqREy6i3ZNc1Yj4IjseniRspyqaq/neSwYpxsm7koLsHL5hsfpnIpyKjXXyuUf07O2Dh9l8eV
ImPGrPgeNC12PoUxAjzZRcvjHBpfdTVqYPeqNCzk7FdwNEU7r99+F4ZxV18RO9Oymz8Cgfz+dcwR
Xpf95AWWmvtG40gljXb0dwJMyojUKDqWbWQsvOKAXM/gwqTxq8V1XhpldHNy3VCM5XNgn1CA7N+k
9jOxS542/ULvqfAG66jBhYaaXsHHX2YWnfQcSd2RQUOQfoq9jwdi0o4ulVxHgtuYjr3nDCQ3yu6H
UmpQxt21r+wBBK+kv1wsydTQEdq8o0mlKutb8TTMVC0ibR//7OSAQNJ/3Hrgw9sfwLPab5dYrKMB
yd8D1KTQcuxepJWXS+sjY/XChjODVxQW81xcLTWh/i1/u7ijC3v4VhwtKqkWBeZqsamjIPy1nQkL
5bSNO0jPgzE8eQbcfjNsHhkkTneWQKQkJCOwvmHpQlmkE6U8x2GnXc7q+929Vt3ltRLH4KWW+Z8d
k4dCAoyMHpWg1JcDyv16LOkvJW/kYzSvNngyvS4mZfEyxG/3O7+8sFvYx64wE/C+ptvJTDuredbf
dm3Zygd4uiI+JNA1qIlsL3TxmtF8gWd5cyoq9JAOvEdKEIKe7j6PBZWJI/VUnND+dtNlZwGytTSD
ei3QU3VF34NJKBR/2OADn53b0daz2J8EyqunLCKWl46TOiuxBXIrs6XQtARPKoEKVb4jwWTF647I
LD7UZgLMT1IXJildoL4/G1Mt22XgfTAw5WpKUFdxPg7MqdHN6hrL9H0eBtE15iQ7fR7ql1anS+SM
Ba2k0b5PedM1q0tKhu/LMko7ZOV+2DYAprHRUs0RzaGzKhH69LJ8aM4Gu3UqA4J85R2NLZ5hPJ/x
ojlaBpf9xSG02buIVDqcwyIzTtfcghBKENbfiZ4FSMHlPRlpyKto8n5J4b9q9anRF4lJKSI+muh1
tXidCROVL27S25QBuek+IDYyO7I5agsSCxUeNO5I+gV00cNAHerZ2hTHHPnz4WBRSHfFAPNeoQlT
QPk08ZkR1/qOIAEVFU5kH9hZyDhLxdp4F/8ZFmlQSWQnnUM69RhhH0LBVQXPEVg0LmxDb46pvABZ
beJkVzW9xivTX2HkBHcjSnrJyCgvRZYsg0q9BKza/XwaLEvNnuc5tMqqdz0Jq9ZMKWBztlpn71En
ZoOeYb/Y5YMAfvP37YM4Y3Pfm14L1hcBQ36sQ1B8YRid84N9zU1g7qUtuG3naeu+l3GN8p8pKcya
L/Px29r2zAw8FljW+aSWA2J4me07z0jdPTyxfVDq2Yomge2IFK1+XeBsF5hKoy6TimVOzOMNyIx8
dfphFIULcKo8eBCVLkg5GmrUAV5qSgUKjCVxQ51zfYoaTIIHdr6JDHvzoFs17MyBaBptiZJ0DUSS
my7CmNdC7uBf3TDyNFhJ1ZIhGsibvZ9s5riUtsqsxtRoHME3HsTHNkU8kaVXIyQeXkFGBrGhIhz4
iD86W6Q1TLNZ/TGh9yRsT/wH8Lqo89ob3l9X8/kFWfPyr/OwdiKPsn2nScvqJ1/DyoGkulRFdLYq
/gGsrvhrS8U09/9dOSY78cZO/W2WWqUL58kY1izgh30AXJxJG/iXJYoPuvgT8WWiA9W3tnuf+5SC
ySt8HRs7LCLH/fPuqJSCIwtikOG/l4C8XyWGFoE/+SGMLNYULY9UkSVXLMQBTTkchlCfg6mMrvhX
SY3kabP3wbbrsupS9HqgGjlQewwWY6zsPhC1qQimTn8imixKJDeZFM27O7Nag5iEsKiZm/n4LBlk
9yVjW9zUf6Vc7uyajnNCO2/mJROXJmsiKzp3HUHc6tzMeOlAQF3y4acGeZ/fr2gU5L70mGda8O0h
AI8K/1A+pdglzOp0yk4JytY65/VtpvQseAACo+B9bGYVsEtCT45NMwc2naeDoxYnwpnfcxrFi4n/
P6rIxSQMkatWFd7xjrHBnietoAJCAJFcT2IMQGzmghUpKutjIFdosafXUkby6MoholoNS6z15lke
LJC9W4O7lk+gzeb2xcpoaFSXP4pyh/Hkm4WGNtOdkDwjaaUH+bZs3eIOxqdmqY6+LtwgIsJj+oXE
FtKMapMtSfGa/0DUdDD18OMkLkx1ASJWDNLZ6FLelKuGDpmSOFxEMcnhCA1VGRneJpZbzTvEsZbT
2aYPX749xhGDoa3EtkFlZSsasShUoOVVp4ejZEmdA01Duy9/QFex9EMm3HpnYpakcVwn4c4v4IS3
Rzkx9KWr8H2TFLDqi9pWkAhmp1oIwU/XakQqPqRN6vnwVumSsOh7mqdQNogp2n50d5guxabXhj5j
TxZzWzfWlT9rxOODMmNvEo8pncmMVtXwVwpx9MGhgcy3mIBwpw6s64qqrcSPnOHSyfHyE86SiYqK
NOqEawcPIblvktuwJ02DzZb5vyJCI+jCulbytb0jf+wLegpZIfDNY/fVVUb9yUV1wI0i8T7OUjz7
eZZ57dhAyY+2vo7ux5PeI+vj7+mcOaUVQqI9GYnoA1nzNBj2aSy0mjbX4TtbVjlUD9NTpVH/uwhZ
VaBXSAUIRA6c4PduUTkQWTzzqHO9Jc733X5m8Uzwuqs0GrOMfuKuVc21GDQ3S/QlF7Elyw0ke61u
apxH6p/p4RakUHSM9ZFR5AFUSpj6gqpYYwgXmdvRv5riJ+Lb32fuYmnMhV4jZ2U5AZxVnxZMy1R9
fMjnB/javF7rDHQCd/bA3FPam667zCA/XeAN5SMTV04P6frRPNTdtfVC2ksbTWKwJcFHB2EH/8Zt
xpuQczUd/2A9YDYMwFpSkpPsw8bhZqttjtzZV0j858M01fxdJVglmjDBCWH4+LivG3O/eWQSIVm6
SqKWDsQGn6QsnQI7a3sViAPgtIqxNXouLH3eJsGSWN6Cz1DGWyeFbMYszXxEZHIDQGNHfeJwC/KH
zW8gP7RjnLPuF0prhYErK03YSx/8SkU0l2ytOSgfBf6fGRiWEccETdkoAJkpK2Zs0sLYvCjwhruk
OI3HllNqvHRGOwtwAI/bgiHQC16UnDWYfL8lyIQjUURmoLwZnCu70qhy/17EXu9ac2BOTNG95yst
DXwqG9EpJ2XRek19mVKMDmmBTyA5iMSKhvFVhxnTwSrUDmQvCqr1qcNZAE/KjqxIvzmgjm4xXVkf
eI/qDKXsQNr+EcAcUEkz4alSsV6cItfhGFHpklY8jNS6V6wEkbvgQufMkdTD4Lbb6DmtJFUQp7b4
XStfffeAWySm2GlN6NAW2U4SH7ZO2UzJK2F2NMDHI8lFRcbSGZPGD10FOqR7MqqqTqosauzMjAg/
WGudt4lttDXnYsA/I+rgXvJ1p27xDc57CYZZOYjPQmNRMSJHkUm+kANPZHKmuK+cwZEoxN7r48Z0
LnFjb01UzdMZvdHyf0zvTNPeUZGnlXjaoO78COxpj1R7j3LQx3YtcWblaWYAg+qVxqxKbJhoCZar
yei9OXnXhLvtdXpkVKAc6Hxf6Zm/Z24imJNi33ydo6p+OdzazDbjDxRS9VUTy4xXZp+WvjF/wpJG
w8uX0NF+NMq1ApbmZzOTmyFnTxY0hNC7uRqgiQ1LNEd+B4azZwiwU5pUiT1y0wcAQoQQLlcMwTdk
FFSJ9YAbDu96dnZ9wvDJwruIAKTy/ToGV/JvuaGt17jwbuC9eGDDllaVbAmaDcywNIplhy1j80Hh
cT+qsLM+HqA4GD3275hU/F0+3s2yMOaLViII2Nswp4iaIO5Wj//+C+YLJAXRJ/W2DrGCC2PdygTv
8xgImY9UhGPp56qPi115IxRddgKnzcPdD+G4jgVejg+rj3K5YTNm0Ucm2T3MGm5G21wCpl8c3XAF
mpkq1ckdCFkq6BGVGrCxG5YlXv9ZI4kJRv6y99JGl7ovUmfkb3c4Q3ZAAxbpHQTDuRdhfbfwXnf1
DNXeVLHrFiyRJ8qhTOI87LMucWvWxAqpRObPS0P/6uvBzaq64TnSKMTlRIsuNOFloCj1uNdMmx9x
S6GhXXgfUS53MmpyRW1yLhDnQlH/ZRqEK4W9RJ+X0KDVWWnEOigu6H9E8/1bKJDMspOzaCaCP0rw
7gfrW0rgAf3IksI980XSIvTHtFLXJxIqJ3O9lJCTNPvc9HcbADpbvXahiQBXicT0qrwPMnugMjtC
DCoLwiETddLzaUV58fsNc5DicQfsxwTPHQfwALFFfcxr/FxFy7hKwKca4Ifzb/INEabel7kaGkvM
R22uLLP8e0cdUAkMDPuspoXF5EhupiA6iSP5ob1TXyBymhF4XqEMdm3byeFLSf5ANUNKLSgva9O/
CgRXzG42qRM6AmuEkPyzbXEtSnvoi1oP5bX4BugfNqsosyQpNToFNqtQHdTAfzsQNDW5zMnLe1dC
t0k8bNafZLnoLESUPXsrHUoYTOWtkVTHvNDP8NmSXkOhFl2ZCiuWe0aOshVf6yZmQ5xaftI0d4D7
SaK/c5SrrAYUtPP1QJELVSiEP6u7cfGxgdDrIw+zh03fSssEnR26Q5TeAGrus1I9bhJFDtEcASpp
F8Od4F6g1Q9QIaLdzbAwbanQMd9YKwHsYOdHRQ4NslY8SSye0oDBPHB/K9SLuHPzTXOwjH1t0vN6
n23bD28vk7zr1cvgSW3iB2UJU3L/h8lVnelV+9dvUOrNY8lptOBKesszbX3i5Hd02Vv11imSnwU1
TqGsTUGoVGf8ax+RfT23TxjgecrLQakMoXBHhHAVziEs5JPu96UVkt+yo3/67FuzCiuqmhZ9fxbx
jIPh2R80hATIAQ+3sTDHjeiOV0yScycs7nG41dge6gdIrbscoUfZz67oPEjEU6TroovnYDkEKs8g
ONqJIQSTdikbir/jZCIym52SRwhl7EdPGUFxSsu+x1t+SCy+mHX7F6onIWlJi14hUWMILsnpbCy4
Fpav3uLIJalvWdAyo5PEQ2paADBh/WRaclgYi9ZBAl5etqEbZe2SyuduRAnGZZoVN4EqorYomCYj
osp60YObUjbHC245okNH57WPKskabgyKhjy9LTqwbgMxkPxue/9VthteEzgVOMqm78bBD8TF0Ds4
db52NFJJdMJpSqDPLbqpf886HDenOaRgzQYSn6YiP03Q3RFfWXRiWBOO8ob8ZCqKXaAeGwnSyhRH
zAr2Q7tpuVNDskpX1+QZ0YDIG42ZGqsNcAwnH66cdUzI+Qnm7D6AlbnVjEau7W5SSbaG0mwtLgQC
8tCui9dvu1cGUwLHsaetNuE96wxW5dJGkH8ydLbLNTF+VJfAL+iAVkclrPBVHn6XFTdAiqo1Xq2o
syXZ1L7mv4MlQMdFcbTn8907oqpOwEF2pD72KJnCGxjnCZsmNIPwG9zyBFokPgQYFdVzi3vRgnwi
O3oCmUyOTxANs7t637hKocTu8i5UUlKLbrL08Wwp46L2MyM38LQGwiJu3QfMUa/D8CaTL4Z1rQLv
IRLCSB55HGELGiQdy/P5wVuNvOqcI6gf2BJX4jz+Ns/NHcJdrL0NhT12qiOlllhXVT51bvKsWcn/
pxhirWRPebOa9TNXRl35POZjCHeSfL262g3TfentqTKxWUUlaetyyOamZFhKBNLROLWaQ6B7mS6J
jcQ0qBTrK2qE6Qu6Q5sen3kEjstch+fVcJyPkFdI8JkdXe3K1RuUq1utoiETuePtN8M4aZuHA6Z4
2pvcl2jq9fsRnBg0imz0i105ShQGUfqoTwK2IRoUxLDdLrn3TVlbSr0uF9iv7XtToIs2sMNwLCqH
KsiZCiG4x9oQdD7uU08OZf14TAnqQXybHUWu5n/TIMk/A6jfEMxH6j9sTOMVzFOnJp7juhutbJF1
J8Ds2ErpVcOhm2Vvf+wOpMLsdB81GaC//d866vlvkgZX/ZuQ9vawh1uWa1T96OMlTym7y5w9I0Rc
Fy7APOzDtoEPALllP9FzELbc+o3rNye3wXdfKsmQaEkrwU2FKsB+r5zVqFl1KcWv15ZDQR/OK6tQ
7l9Dn1ksxRHSMpaXWbHT4yY2tYiUnrh0TA7e80rSI0817135GYuvTBM2hKWj8mkaSTLbLWmM9wT2
jvtRhnNE04yx9nGsnfgDOpxy7E7nx6KhkU5mk2DwJPqUx52eoPoSjrqdV3kvxm3n9MHqKKthAC/s
0RHg0xKv5ofD+cCq+k8A0krrLcnFrPcDn8nlAIt+SAc9Wb5w9OLe/gFt1xn2sjh9b8oEEVUA2La6
SxKIiH95cOb3OkvC008EAl0bGMpesNRkJicqo2LkyUNrM40b2Hn0B84KXrcU+cgeTsUEHNBj0CGR
aOlQ8O4XRYADH46ftAYNng0k8+PZL4JZYncwjpH9ITTrm/0dx/fzutkz6ngratyU44yUNtVolWfa
cLw4GoVgdlbkDhUXedIDhYur2p+ZdkXNFlg77jzo9aCsxaW5AuuBwONb+Oqqwf0b2++jXQ1E6ZeF
e/1WYXUScpBdul6F6xGSaemcYd8d5tP2hzM+7TZmz7MQaNLZLiuElqPtC3jPJE23Gw8LV8odwWbp
cABBcyUHgUVYsJoEXbCTzUbG6XnYcSwiwkHB7Ym/3VF+IiTupg57wDZ+rGhItd2daN89XAPzurl+
jVZRS29K1Kpwe8B1PPQ3CDX94KX7JQjSzlFc5gD7KhgyUkK5IA+jgn/GBDQ/F/UEPAA+lpXLP5sV
MZQqnUVrGjxHnInhavvwS6X3QHV1RF+kBrcK37cWzbl6VV96aweCYTmZ+/Wj43c1An5QpDhm1L8r
IL/iGiaKpgrGIVXW05YGkDnXvO3w5jsr5pZzlDdaObHivFSPMfEpxgMy+HPwMMdrHjVqs9AX7odw
dfKlZDTmYUxRgBnZLfMHLV6I5dqGWx9/ilDHnFCS0QAHhsCxsy3RsEyfB7J2ehnTg+nJt2qHlhkb
SwYIgED7ocjnQIyc7JMgg9Ck9EWHt3/smahiwromAVpVZfUF7+VRMpZsM2sYAAIWkUIePSgT7De2
7iV3kSmDDasGfzYNUQJ0orpX00oOsE+kprCDbJuWNibgC7TWV4lrYdeiM+gpQWtkcZmjTI/qWHMN
hdb46lAz3aVgC/IKaP2Q6iLOpCVgWGvnWHtft9l6du7Nn0QIhWueOPjJByDmZ4NYWpfnn0Pa04Vl
ozkHWgQLwon90GSqZfcdMFdo3A9ZdKjWWt7SECQAzpJAvfKWIntK0CdtHogigD7nIpad8IsGc73c
wPT3AdK+Asgd3ODtn6aliZRTr0+rXvbTG8YBXkBcBVPKRoPmsSbRtkJ7FfyMTWTjCZ+e8ffLq1EP
Q/1/NLo3k+A3tLkwd9H0U405lEfne3d0Izjexk3FsWQ7SnH1zgHszqYlmu4d9i4d3yjs0P/Lec/R
/C7KWXDikuAARfpBuGES0MoUEWPpGNX5bOwwLQFnTvLX6Ai6gIMT7xSWhXYd1ijmQmeGaZDkw/O6
dIymqwCBIh5PGiHk1xfcTo+dXYAdRtDmvIk0hsEv3v6borDUstKQ48JqhuyYqG1SQesbjXNaaZif
oriCtf3JildAFZWRp5aBgbA/bnGZ8yCg0z/VATbKVeb6YWEtSOX5/2/JpVnoLj16hi08YaKcxCV2
Ppr14RhbSXV4L4WqjeWLKaL36AIL6K7nfnD1WQgHnmAS3h7Kx8HJMtuHg925qIays0eHlKJ3y/Xw
/XHE61uRjN/3g+HJXk0ajDQZok37MMfKcY0Wv0AWyq9E25zkgxoCJiiU+lUF3W3O+QEW9EaQQ8dL
JaK5UHqaJFCfR/IXUJr8mWq8pktfiEwH4Zy2Y2VPsUALK3Kn8FCfRAHiT3TLLs0bGO3Gtk/3skg4
no4SnJ1Xx/tYl6RVYLSx/XNfMfW0qMqh2WsAkkQdTrESoQXojkTBEN01BOk8NBgtigy14vIM9IpK
kb/M7MeUcwbDEk8w15YV6dvdxDXObzqeiQEG2Q1eyYjjvYsZbXyxxUJwIsT3c84Jsg4tAFS0Pe1N
JiKZbMxl3tAetu5eb6QriNYSW6VQOHhnwjELIP3VGXGYQbqJ58NPiU8KPs4zf4V2VRKd3p5pGFUW
A+zqAH+HZfnO8lcKyIxLSH9iBkdYSlwQhlgxBogpywNb5YSp23modgIoi+Ec40QXjWvg7hjUgwgV
E00dIvRIJ2ZpXTRo9N4vn2c5j449QnY1Nva9V4IZLHnyNUCPmYR5/zK64OePKmdC4E+j4fWYGP9M
eRPrbW/n0JKrW5d32MEdxYP7JZFkqSjLcotO0mcwlHT/RKh+8Ckw8vZH5Pm4KaPDKF2VJ8xbmTAD
6raVCNaAk0E3/IcSTqVbk+1rUoz0BH6MD38UbjDXuyjb5zbPhRB/I8bvO/Oy1wc/y5HtlLgle5/o
yd8Qo9KGROH0eMqaYtP8gJiP8idwgT0A+MQAIFyEkd6DQNSMH8O6qdoyxoVmQNjk1aluEig3gTw7
F/BS6bhzmyOPKsyn2H0v8BKiQ+DL3+f8uW0ZnLMWVVu+na6QPPkSKeM+nw2d7Y9ZKsncMQtq4go4
/x/bwZPw72LlOIvJVaUvFyDuACpcdLrM3APtsI2jEu1sNoYewQ1qDUt2sd7wmoTolXDsA3XxtFhF
ZXn5JSEjCSSOKygCOapti1SehLS0UHJ4ySFtNSz+uVjoZ7bmG5gZ+9usr5tcsW+fii2ikbm+qnho
00/PaQ78TTNgKKdBELM4xIOe9oljVVbTw8gR4XOtuWdrNBa6rRTH7k1oDjN5CQ7UZNdL5sU5Lx8K
5KyKbtIpNoKyAv3+xqc4ahJNVOrnAQ7ODead3rhy3w4d/+x8k5gND9N37Elm8kJgibmb2dStUQR8
XgPbGvvZJUALLP5bYfQGjujWht6P7jLAjqbCmkOgJbJ0z9LyrJZ2eGkv/8IPpTJL4cXCNuM3M7jg
aIguTDSJDz+vIAAPiDd+4MAc5AkmTCUW4hgMxKx4leV95nwtUoM6w5qq3SmyLY3gsVi7fhgbJJ+R
seP2s0ylM8WQkwL5DcyJLq81TKtHl7xr5doSkWzS91wt5myIh58aX9K+j1zWyAgMc33fEXkbwx3C
HJaJL43CL64/piI3RdyxGphksxMrx6dBhuG8UjGmKI79vtd5zoTgXC982sFGK2PgA874nVkzn+ei
rT2cDLnHWvLtgT47HLuuzJdOZ3TUhm29CAkM5zdSMYpAtgKswkELlTHMj/DshIvf6IpDsAJBGrD3
VWq8BOWEP6/1ftOXu6gT8HlynKwrNQ9wNKZ1Y4hZBJMKZpWumSruVI4sfPOgGYFuPbrG0F4umiyy
b/qMVtqtygneAnrJj9LpvtB3L21ELZvpdanxGj0ZEEWayTaJdOaC1sn+iHKFVsMkxiU4cGx8s88k
a8aTKseo/1my+7e4vLiCTUReFLUqdnGsKsnkPlsG2VFonSRBup4L4gCItgXyfxmSPSfb/aK2/a4E
n8qOVGFwIOXK8M1fdKCIFk+gO2ZdYsT7eLgQ0+oE+AKReI3zciq9GFFgqx6kLcHx8r7L8LlBG+YL
g3oBDsdMfUMVWYGIpt+g66I5bZgjxV/pNMkF+a50nn4cmZcOcvapqtiT8V0opJVockw+NRP6ereY
1Qd0Mv+AknPwQjk3wxDpVlp6h5vHfTDoOkSv3RK1IBXYyRlfeM3hISj5zXZy5U0SiKS7uLQREmyD
/tFyHbW9sekEp7TOyzYNS2nrFnOyUTtwqIUR2Sy9o/tcxUvKoZxGcosrziI1CGhFJ1Mx00RgbgWz
oGZGPmCIez0VDh2oMqZE0PnIgtkaULR4GgFm/AJ7x+rrDJ9jygnHm7Uf8jBjiuQW94x70tJgimHn
+MSIIq28h+c8IyfwNzhtUYJ63puYlkUWQzzCtMTV8fJs0Ig1h7zrrzXSzx07zL/0+Sk73AqFJxMu
A3h3I1NMc7CuizwJ8+fUbx6uohPfbKU4N2VLDOVVMOHEHE5YIUht1RkmMsFghjqi0/ESsbb1jl42
2h9cB5vt7RCHb3o298YcIZya6ej5VZrRuxIYNHcMN7b/j08tzxovqnTQfHa9W0iL4ODBHK63I9i5
/QU2PrTZUgtGINDdh9IaCkJaIgXNE9pvAFpbT4DANOmR9iq7nN2YbnUDObIMJbYpLF8KnJf0ZK9Y
9We68W7RYqWqEOSxiB2blSNturIH3UDSRXsQU3QsxVkFkIoIrjqnpDwTFSqHckMrfs1JqDvsBQEf
IOV1TQ6VO+Z3zvqOhZzktbszbXwNj8kxGaUtjRgss1qA89Aqq5pgkG1Gbgc7nMt5AAIDm324AaOR
YmHnxoj9WiVv4TfXXnfAcfU3Trshm4sgIs+a3tpKOOydEeJbq8OGofkQ8LypE7v/5dFA5kuS2aju
3OYEWdppV2O4af4IileqmX8WTSxjWISjUyl64F0Rg/ByRkx6b4AvI7bb2N295xk+qqXIjCKPGuPs
8Ij9goErmP3mTV+EEX4KqlfgTfG9nwnBMJjcgBVYgbERfnPaD/BA3Y3VAkjrbHN3LMUhv+1Lpf+W
44jAo7JdyT9eF7hkzlaQrKEiJwplIKPSqTcZSFPAOYxy7+kyaXU82xAzpxAgHNJHdBeHrs0jwMmY
B76OgXJgxkZSZuplUJQDyZGa80tEmMBd49PbxCdmmSfkYDaT1phoOMuR+zxW3G84CAkpXEJCqSNF
UvYtm/WPD+rbGPxKdwulc/1u0Is568L8DVtSDDAcwfqlQ4g/z3D4cWU5BMLFnl6j5gSL7VfjdsyB
ePcrSdEDJppLmB4UwGIi0Yj6QEh+DlMKvhVF5IPbQzBpz/4K4Xo5lBTwwHns0E4Nr2Eq3mpI7M+i
tc10GEJbj5eX3s8KoVdEwwW3hPKv+oKpswBbyirPNN21p0omBraNctHJcZ92IZ9SIWs4JzxECopj
8jeqsMPJxnS+A9stxanhfoTHj4MXTtIVBexBO/CYcuoedGM912/g+In/PfN7nRl0aQYSzjGA4Z3Z
YY/BZtifz1vtIgbl43JlO0iaU9GKBioGCHdWWBaJk9DDebJNMzcAkfLQxyhXG23mqmTgSFrSiv93
YdDCZjknqLOn7cpAUDjEsl15r2QGa2d7mzB06x143bo2nKodmxD+kDDfOtbBkW5y5ntFM6BUH9yy
0MBJ/PGEkRmtkjg0I7UBOueu1WjgyjM0qDaAe2+gNkxVv6HNQZPPwwF8i9m5ZeIPnk2i8o3muXBM
IQD1tL7A9i2l4nFRaUshWuYrTF74uFJ0uji8dHd1D7GsxAZZV9fjZRgtL2BnKKYKmpTR1bkGCAsw
8n/Vt3fvcoEpqqvoH4lcgGrF+aFhhaaamAqAAAzulCeEOxDaU6mGhX+m6JgSMpoJDoeKxGMTQ5R0
OMOLQwdD7HmQHs7d6v0qtsrMnjVpxT93v8ihkBhwZkMSyH7LiLDnRXt8xiv8EvLwRnkJUWWihCIo
U9Q87Dcexs7NrfB5gX6/8beKjtpMpLe6w3NiqqSeqxlm9kizcWNKrCyg93FCPUZm/OGmVpCfuiW+
J/NGgZQ+uwXLFxg1rDdt2sCtts/cgoUleTeKZQ+qGCqiIMlviREjpjEvWA8cc3MaizDUAyoNNm89
aIPP8U3Z9+Fmdd19sJcuknbQBZ+YTXQaWnLSINXz/Ff7lM3WkEfAKlKD9nCvylnrqPAT2AqWBQZV
z6hBCXLOSpWY+eDHHy36ZKxeY5oif1PwFgOu8qxnsjl3BFQYL/lENpkhVOVFWrOpmhEGZ3qqhCP5
7RSn3lv7dYe+spSQ/PcbxdQtmQlhVHlBKvqgMmjg53hpROFds/KaGjSRKhQC07i5aEN9pb/Q+LHN
FTZwgI6XbZuBsJ8DLL6ZJltUihAIDlRc4jnJvvdM7wNrHHN0KSvfG+iJDWkGXWOrEO+VC7hqiiYK
mxsc04dM0AY2aUK+fwdztSKvb8wYvGNRStkGpAO7fwl8WgbHgFKwlpSfsE2ALaILhPTKRv5cVMMx
J2YmTQgvRocCH7LrJfT/U0DSZ1rmR9/HWvYTLP/hngOwyuoLmoh2YPurBTMDuY1NAP0ciMYjB0CZ
frlDWmejesCAV9gKtsjLE1A1VevdyNu2KUQbJmp6ZH+gSvPkFx2BlBGezbiNaV0hzP8eB+Vp4kbE
gOObyFy3cUk8oAlATKL+AEP9nzpIwQbuTr2zYD/Z+Z8/MNxafQOsbK0DW0Ikt6YBzU/6ff28NHPh
YSI+bjvE8i/ST5L2dgSIeDc+SVFpXuf3XZbQIqEAfC1J0yKE9dCW+Nsxt4aaBlUqiKzAfELCTYIc
ZOxe9BMFSEamU6vi9orve+2Y1Hh/o4k3suCpPwC55srNlgs3VtyqrGZvwUcsRLavaKNQhHbpYDqH
5jugt5XJvVdV2SwLHOVcjLODSIkume1vm/TA4TjFW4uddHQm94u/wcfn5Ji7jfOY7GYGEmQDhr68
Neipb5dLShnPidnbYJ+oeO5z0je9h4j8MY3mSdxmyE0oxsJdonscx3IDNHvBp6LUOHwuK7SZIRFy
5r9hB77sMNJGN8Tyu8bEEKNSxTaw+I5JOmHI6GCeXEqA3ohdGqR95kTyXEMLsciSOm/X3KD6Cyqp
EqAR2E6Mn8SldyYIhpHjcwFx0+wEQOyqKGl8VGUtVUvhVT8s62FiSpIzDDLlnD5Eq5ASRbW96aAb
xjU6GUfTD51Ryne4YLriIOzHyFbtGZCclkAAe/9uQYOKmuclR0CUL9H0foXuNI/J9ZpYpSpVKglz
ZspAkvjZkl5UTg/8BXSqy7GqW9NaxlJk9VaepRoyMnIAkhiVF5FTzIgqoUCxoOzSW9Kwxe04iOg3
YxmID4tliYuF/8MxdATBUqC3w8si5GmQ8xTlIVpEAjare3DkOFvJVQEY9umdp4yH7l16nxVHCKlx
xNem7FLDimjQWAD+NBbHbnvgoXA/WqxQ3CCc38mbnNLef2ttFV8s5P4L1WFzQxXuem/I7Z2XT/MZ
xJs9YrlGc/pXBZ72+fm6cQQtwF4J/eghzUX1qz6SKmpCXsgq8ETgssdGR22LSA9C+H/AdXBgJN5V
1HGG8F7TiPekU3m6RqceEkGN3ZtczsgnkQLQ9DMswQGWJ5xoCZEyHmqYkhOphpEGBb/szAMv1gYk
Leuqg/dfj7mQuFQp6B45p14Uh46XckY3DQRkoLbZE8Qu33QxXo0MehyExHy1V6e0gV93pm9AWzbf
LIhPl4u1SjfKLOJzR1KbeF988CAOFygGegr7TDkCO5M3RusEYBFUyd57az3TxEdzUq1EDihxL5jn
9gP1+15kMTLwo+SDQl7fT9sXedGk5tZi1wPT8WyJq1wn9y72QVcigLsnGP2m5Eca9nCG9oMUQqlJ
OAK5lAk/zVR2YrzA9AS/kEb10DU/wL1BHtSZNMuf5XQvGnR1LLBuI+GVEqVORLhp9VbXgtoHSSCL
kvTi814T+k/B64BuItTKqfHpWu2B7dyWZIhRxZwTfdhjJ7El7JktQpyfoeQ7mIpA3BAnEvzGnKI3
f8+N2xYTvmpdWgZgvLGxIISbUknQ07FTfFS43pRRgGKLyMNKpTk9/uvGjBb6+J9wjEjbZT+CJmts
ygQyPHB6pIkNIVns0kDd+ddB3RrjiUIMCiPgq43QdLnMKqO5YuPlG6+7yv5FOoADSnXhejjZpeN2
wsNj+dDOg+8AxwIadBlRrboOQO6yXDFgrAGDSXWaZJEMij7i4ILFsE1CiSLWQETFkX2uuHNnN45U
7qcl+Dv/Xk3JyhUF2yiql2EqT2cC9xr5sH6CJ5r4Ad+kJsWaZxr+LLPJEz6jrTntn+XvkEpNSxFy
cVyQklY4OSon/1s3KZudntktmeouvAckvOGjADZrLoTuHNzA3jFX8F1ctGMISmsWF5YrKa4TVRK2
clZrk/ecoONtgy9eHLhQZr4i8crQAayuHT5GrYkifq3Lm3IFC/hMcjpOFnlCXv4fHxgYuIIxbtJ8
JjzDoirPpfbstzW9nurR45VwxXBglscwC3wAuA/YMAR9jMfV33PF1Cl49Xr2SkQvKcAIXKuVPfkZ
ex/sXMUHjarNjaxdnkX6H4crolnQXkx6DNIkCyz8dZj61wnNC6QpDRmMuLR4ZO4ty0DL9HKqtTTF
6jPi9nvJ1qV+ZrheJYMSWD4DtuJ3cQWcJCD1lgDLybYPLT5tLcxxTP90AP/28KD/qd9yw6XXzyLX
dALOdr1Px1SHYSAMp5Iz7sLsGwhvo/B9MDqZhWDOrA/YLCkhCUWVezJ6qssk0NMxH7bT5mc/YtBu
m7iysxwOIJRgQvabHCRpp/OXV3KGc5NIInlJDmqhTm6Om2ubZXEG+S8inXzidf23B4RTO3O2Hc6S
9smY3/ayyeyBQ9QgcOzJR3nx39841ZskDBfOCMzrUfWF5h0C1uEwfNPxFWnrc8XOKCpxtBIUjTsv
Gi2UTVjT/R5BJxRFH7mEi7G9IMwwyRrgimnPFayQPUO0TpSENnVm4cDBi0gkHc8Q8j3QdSNehc0l
hGww7wRovxZF2Jw6aQq01QJkxpkiZNiuUqvgMDXXPgTiSUFYpM9uRi25D4tNF6BKrwgpv4Jd3PAg
8YXcB18tlnxpWNMDqX6R6qv6I4SgK19wbTrRLccS5SFuu7D94AEdZ0IXEOT3ffqjNqYpV5J4iDJv
t62AJjPJdBHqSZHSmRSDIHivs/BXgdjbKeB4reLvr9nBqn7R4/N9anI1OMpAiYhK5A/2n8CBvt64
ynvcmg/RH+a2z+7HwokJxKmNKkkRFGE+0vGPRlw/jmfHPIFVhnbgWuMjpCr8inKEjxHA66HDB8gA
pvFLJN75ZsffmDUEzARF2iNVRWW9OmwuqoZWDORM61l9ZGFFlkpaeMgsQfOGULuipHdNP0Rdlqvc
YG9elvfAEz+dQ/ys/vWRUoNLZINvF2uiTfmaAOzHXE3V5IzLoI8G+XgY2oPXhSC8MG4jDUooqjvi
TfbE5K/0o1nJYfFT9uTNcg6xJ+JWVzr01AuWzIl6yCWLbK3v80HxRxTS5Wa0fbdOF2i/MT8HaF0V
RPfgX11alDMSA+MflO+15qmSjmpGb5ow0SjCTwIXt91oOvhW5vDHPX6s3vt5RWChlYuUFDSeqtqE
abkgd0wgxfOwZmprYi0VQDnfac0KVuERfAUzI7Kjw03EoW/MQVGpXupuJQNhtDcH7ZqZ9jHuE+RT
vpy/xepxH+oDPujmSfZDFRl84nVyKfCv/OS6vghbRV7xw1UlDqQa8870NGYPvhIuPh8K6ECqZVyk
DxHuWMyAeCGUu6nRijAwJimRkQ/N+LUlYwvBMYEhEGdJHybB8L3nKFsp4nAX0gyiUWbo8OxAJqOL
zF/PbS4jFGR90y9Kx2HAdQEQB3Rx79dxk/2JHg7E+uT2Vv6OUOkbcS1ZoYYInUZMGcbNkZt5eGwI
Uoz9toLv7PEG52KeP0C1h2a9+AxcZTlMrHyGT41w8V+sk75LUTtgjpn6EaGUsJu23m4nfdLA+kx2
wLc0GB4vFUD+lVM3gYUJLxB5TbLLmTRFQS1uWNvCShOHcHelcUEcWh+wwzjt5z9OtKVL7zhsd3Tf
7s5pwFT2VSiJd6j7tpUsZZXLAOtwdoocHIuvFpbh9vHjnlKMLc/52iHMjFBabJzZxWEw6pzRFHo9
JtS0ruGnUEa1eXsH078qw9gxrf0fTATPAXoSLxnNRTo5XRHBR/zctGgs542w7lYgnZ4dgtn/qok7
k0mUyT72/8O2EJiEECoxfILF6HkyInczCuia5Q3BiPbXmjBrj5bM4MWVpQtxmIs3HwTvUr6U/Hi+
IgOqO0/5OlLuZbSCqPUNJYRaeOUdqU7XQtX4FLLT1LP1zsH0meqwRsVPmd36z1NqfZ8BZcgxCRZH
3mgBxrhpMoS6J4bhqofL5tqs0G8h4mZapp+hvDelCPqhQL+5hnXQ8KUN2qAeBcRRc+7FGt2hpYrN
SqU2dGb7XArFniwFV8Q2ovzu1EBHoLjXqzbV6uYSeOhL1+Th/HWc3orFaLMRW2IMrCjHmOXqCfTx
OgEez3u4D2aIQUm1wLrFsAZndUqpM35pe98+e82vMbz4gBKAbm4f9yfFu+U8pnF60qQxicJ9Xf84
KphNjmM64XAScWtXZ9lMhTSieuy0wQmnZV0tCWh3pkUJGnzvfIFaW8mEd8f7eAIeSaIZ2DhtI4u0
JTPwW4xFtnUkX+nzzGm44x/NPaB2/Lfr3voQdqtLYbpHEwgEaZl7EzFqrM4BxxTkwG+c2Xg8OqhJ
6z3ZlMVvpGJYQUypkKpDxYGdlDFWCSTolxH1XAJM88maqdsXg3CzqFmqEgWkocH1Py8PQCfOnehq
iMCWGh3iz4Fx19ikhZOkUopVwxUY+1jLKu044kP1yr1m8slWsIennC0lLx0/mgp0YEtmz+rCyUD/
B+r4MJ38su+G26FoglGA/tgw6hYKoKW4XzjupPR3Pl904YK6WHWYyrhjAeHrOS1xnEDLaiQB7umY
0VVz0h1K8X0twRIslsQDt5SS7cMUyd94CDy2LatweOUK2BZOC4IfN4bZpE+cybLNE4GPrl2kutDj
Q4S2OZABTq9TprBOyBN4CqeEzzM2y8T64DVv2mJyPApHMGQYx3ny0udN1WfjimAy9D/zz+0XaVaQ
telP54e63xp3DoqU4JE7PgXIdKg5G6XLuA076nGG0Sfp+zLuOCN8l8jG65CBOkkxQn/gh3zDnpYJ
n5QouIExYHXwJxpdDM4G4HS7+h/IVla00v93JOplLX2OTQXg0p8QZCLOOZANAeyX/zC9folGF3/K
K65Xy3GIboRC3fBTuskX3rqaEFILjpFWKQs7E2ssK1oE+uvlfvzLDnh+szYILSnP5jL27RCA7uY2
ZYlUq0HAfawySZmy/n9fSI4xGBWCOCIkoiOq4sz2Bl02zwiALUidflTwOCsuE6uixLnhti4kayhG
wySX4sbMcxwcmHdjYFHF2vpuLDPKBYoQo9uuF4Oxs96Api9nRO+0lcOLdzieoqwc5Pmf1mwSQgZW
K9DChrprqYClQ7J3lOXjiPW5vY0hi5SZpKtBydUtIs3ZRhCmluEHrX4aGwVzMWsqHELOLy3ohs+y
66BKOg82DYZjLduo3qNuLVj5LdN2WxO21hP++/hJ5/vyLueI//8XlCe4Uc4PoDVw6pFrrt/hY10a
9TzelmUGk5WXD1t17p0/bxoBOPYSube2G6/I/b/fk82ydos8KwnwBJY+jT7KGL9bB5VtWLKQBVdi
SjfQrxKZE3iik6lZ38a/WSywRTIVl2JLMfynhyXR61+htknEUv7HKM+xmWmL0cVj73+yHcjc1ZmR
Mp+Q2Ly7wv8f5e9tct4XjujaaW96EjGYf1FZrYCaGSK6mKWC2bqOpLKaSKDvypGlyXmfUBt3/cg3
qCfojD6j1JzrAKJTgq+wfiuAP6dxrZ9dd/IAAgmo+ojdc+IWy93xHIVvO2v3xtJNYHpoosxjZUjI
yuYRk6LHZpx9wJOPGwWWih1DhLQZ+22AoLED7MROM/Y/7Ytd9R6V2Irmy1eICRpi7XHMlWqruGTX
SbAHBWK/wYl6BvqCPEEos9a5qxjuu69ZRQwP4SkyKSHdZs1lWQ4FCpw4BdaCg6TpKVkH0F8VK58D
3vaOf3PAkhTt/qMBCCMImXNx0djtlnByuzYHESnwbcrkYxhrjcLg04E2nyY+hQ60ypNnxMEIN55I
swaCjls1zi1cQcQ/ZX3XJUhsrIBVUM+xN6Zimh2aNvweTXzpE5mkA8+dwuOdj5qWBOUK5fcoR3S3
3M+IWdyndVn87u4tRzlWYuYB/82sZHsroVj03kjxQUQXqIiocM7efB9AUqQQbm1+u+SIJvCvcJTR
nOais/3QGhv6CAZFK7YCizOxCRy2QHjHGyDzVDJ7OOK3q4bkYc4TZzd0US8XyOkmoupk4yNOtVE4
eAqoA3zB2w6+cCkfjTILFztqwpq8vqQxWqQr8WBMnjnBRSNCrty6KXTaANgneuWLuIyVF+69FcEQ
8PsS2WnBawj0W+NNEcywFy9QXYmv3X9Hbuby+jwa5Dxj3ks6+1uALthSHgVbSqJHayi6b0PSnHHu
De+vRj8MmD0yebRQHwbralufU58tFK9vKyZDTekRNFErfNgIpNNaTlyOKCspKrk9uAFOOCXNW6TH
q+xI+SexjrX4tkbLHRLlVhQvNm/illRmz3X/AmANZ9tq3soLyY9ts+hhrRfKhIArRVw03+6ZRIjr
q7izKVKB4eXSfUqjWePQDHioW9/UBtiUdCyChTFc9j0QFgoI2TN2ajBeUliCsfmA/PdtiCJMW0vm
mze2nl4Fp7HOZD3kBkM6W48cXvQWjaU5M7xOJ2AgVR8CgC/ktbLL8rfDfFhuwdzSeolbuGFVjSOK
DxzplGwsq3KUn/zSiMoKiExCsV0bm0ZkbGBOq4pDPg/teB1NDWy2h7329aorrbtfVUcq+At+FgsR
+P4e746p3sKkQTJfXDjlwJALCaD/cHH0hrzOdbnH4kbHsntOBMRpCrra+rHVMttRP9NEeMwx271H
fGwOFL5+DNIu/dxTS5VK4Z8DZLr8zAGA46xVSu9OHcNt+PKQ6/xmPrwwsiff6u+bVd5UAsEXBN0O
tmQ+TMmy6xeFVG9S1zIXGgTuIACZNoVgRbI1uQH4C6nErVU0RNsDnvHJ4tr6Ecw2YBJn1BrB9x9v
tSGkWZbuDKUl/+FUyqJUdJttXtNUH+XJZPRD4mv1XK1lcf8OcVhAkDUl393mZdI/OVoYBiEpju6h
RJ2lPNiyI7SyrKIGNJD/fVjaHv43bt8IvxMQwJJdPjxwqizDNZqUuThpHn/gGXg2YuVFI1XInh/L
0tZFWmF0dc8GhTyOVNC4+z0p+OaGewLJaWJw6rvG7EFw6wGGCm6nl+T3oCA4qFRlIFeZXe060ctc
doT8ZVi5KwJ6/ER8lj4NlvCbFvqnZJB+/zwcNXWjdzygYv3qkviUSsjS0duknROknskopHgr/wlV
UfcE+hkiNIKcVWGg4RnCLdrTYTUQqZSE9kfwVN1YNqrxQwOe7xXkNYI2AjJaXN7+GWplWi6RAORY
1DeeX/VC9ndbyDnvrfwz+QxZuc92sIZni6q57Ey6r9MLyFiFckitp150drfw8XZ/1OZXOLBK+T7H
hiY9twucUwZr4pFIzOcbYjPtwf8GagMLGoRv76Mql2ESrtborxS4DYJm2+8RteSuUfKqrRQ+vT9m
sQW6TruIIfRIqIx0a2Rd7HJvvXn1zXunER7Heyfi5IIrk6V6kM8LrJW1c/p9r4o+n15pGZI/2TtX
rFT5ifdMPncAzCSKxtilA4xSii8Xq2Hp/G5nP5FyMF5TcESEIz4yU1G2OJTwxmIChjWSse60LW4T
kUgH6WuamiL/JwGikBlqCyQw8dOuxNxRT/O/az+4N2E/ai3vFTU31WEE+Y3V59LH2QXvKabi32fW
ESdc/7lRhJ/roBP5qLzz6k1Sc76Pd8AZKBUzkQCfGeZcKrsvEyAL0k2Xy2uRN7gqL/XHd2q/qx3S
JGlbOAL64sUzBfF+CS0HIKkSIuqlmwzrhs/IaGY4zoy0jrBic6dvYGx/3NynSH01JtdfR4LwWsWW
4rqPsBlfYQ2uzgjjboFas+0blW7QB5pPFVCvHHCzawMaNu24qlqvxAqq4xKJT1CjOjJtpv+f+1yq
mED89PJM9TmNh/38KbXbBYTW+5/TYv50722GqPA8cJhjLcNYxxEK319tifI6NxAlJy6CV+uFpXsX
J55KoaFKzHuXdzt5LD5xvsZiloji7hRLSVsOwZi35rlDGPNgPa94xeDZ6S1wyrUBe1KfClhUWs6j
2D2AfEq0rpf6ywMAA2lyCzDaIaWvvXVK4d6zvPPvn5eZRSjUC4Z8zC6sqD6vQ4eGeYWNaMviDY/U
nqQxPL+cgiPUPMC+0cR4TdII8yOVe3tMy+PhKWBQFjJnxRdI73tYTvcMK7AMOu6bfuq2JtVoJxee
XZwk+kUHVol/VmCETARXPJpFctmsTkkSdqvXvZL8Oqo35uzCWTCkk12yhhm8er6PputuFMu+qIgd
g3nd2StKu9vQJ2rDqNef8RCoSN+4ITqNnZ2frQTnxMicHuELLfJj4nNIkBMSxXj2nUMqM+bmiN4X
0G5mz3UD4QnWYj4xucMSSzappvjVHqOfLkoCONo7DYKNl4ThLPSsdruzRY1ReTiNc2zcqrR1l2pu
k9R/xpshB6nYPz2Nn+MXZP0YN29e++J2LVdHMuaj3dt67Fp9AtyQgu8bMHagFG5igJwZfevp7wQD
04MFFwsu2hxO156aI47fv+Dee46I3QRL4qKd1Fyo+mLT9BW8nw1E0JxQWDq9E7pk87w07UteNH9K
7zkGHa2Zdn+0dXOB2iLarPXTjqQzOP9YykOq9s3nU2Hq4CPPWyU4r2H6WIRp6FiWi485vcakkISv
5PiLvRv9NbAtnCaVpJiLFKBQBKHxjzlR6vB6Q4Lh2fCA2CHuupSu4FA4WbvAIpdnfRaYrRnDI1WF
JRgNa8uMwwFZzFTQgaSfONnquqYxFXxqm2zM5HkK1hO2WilwiqaHz9oIdwYWW0uHEd/d4VxlCNB5
6WsuRjIYf68IP8Dj+AXap/gl3ZBjkD61uGMGG5oUVet/uNP+FtxeTy+yFH7NqEzWmYM8mmVwfYkd
AnH5XXA8gbsvqko3nCtOaqzgbZ2P9YNIsi1Zi7OLKGBkBCe+IN6Tas7xFgu/65PtVkTUSoND7iNI
zRtMgc/+9PNVfIVWJ3DMSUIOJxnU4w73vLTm6Ka7H4ac0G/5F9kYWnciu9gPRx1RzvvICrw54zpL
xWeyQD6UgyAVhDxqCS1zuuGY4lM/3MKgTqClVjw6gIO3jHgAXddrvVJ12kCkqVf3XE4ihw4BDeQ9
xymkh3yBk0roK1cJ+jD7p+7Ujrj2yHZcKXD0XrBsCg6oV8u/jbrxmrVdr2WG3oe3G/yn+JED8X+x
LYKJmVmIWO//iyz4pb1lqTIIN7/SZ5yKy+1OKKCPCPeD0QtxK7E3N2crBjYg82jWPr+liz4AVCsg
WXXAg1fKXxKf6hT2u9M4dYHekKhUhHwyKcHh4CfReQjVEK7EbB77bTEAdOTRycWCtT3imbgJvLTi
G0KCXrDd0/C+ELb0+MOYD4ZoijerfMJkNhUjgVvAwajbSRvx/ozgJlqAUJro1oQSxS1ooDMi7t6c
5btHsGTfgeKn9ZvOZC3mD87HviJ17sdrAKEGg5HbEsFkYZQDacNSsDXjiHnNhxa75ff07dK+hXd0
2E1of0aiaDoaqjtk5v2WsbQdEQtluNBpC1OYelwgTGayxo49Nt3onzG7mwMw5WDYAJYMtLrKZyZ+
FeC6ZweaMCWIILurBEfZis1P3/QnCciG5QeGdasrPy0AQ0mGE7A0lM6mS+bqyVEgkWkwjNaN6ned
qahda2PaAHskj93TXROohy2u9l+pYdUEIAXSv39/Dd1/lsUUhtgQUs2dcjAN0BeU4hkWjtTcT32V
/h+oSiDYpiqryG6+nruiWKWS91mirnCadjdAHpNQGV6OIFfeZXR0PiyZ3YAGXSnGmswieiAXypj2
x6grEvjq8CqS0qCXuewqVDwQPWxCsQyfh2stcqFHdEG9j2WJrpfxGA4HXF8MpYSiEScE6OujAMCg
JgbdZ6GwqKc2MUQt9/Q1qrrJWu81+pWDtuo0xos2SWCUhEEJs4yRikjdxesXYCPtfeyQhoMvUuHk
MEclEBKuIQBoRZSq4pkfFVq/Sbqz3Ly15IxQtqZVgIAae/d3Yu53cZF7xU1zYGi/XjuMyqR6V/xX
WWeZtnCCAGEEJ/UD98gudKOh2XA7eKWOs7xp7p/BVti6SUy6gC1kR4HxvzjiMer0lAmp5eMkytNI
KvD0RO2Xjy5sCY15PlihFKWwLEZWuKi5S6V+UiG/rZDeyt3PmUgzp0jcrFxIukP2xBto/ZApG9dG
WXOhemkpYTN/4V27CZ/CUpeYIfPqWZhEwOmbQ6Rg0mgV/5ZEjjOXXKNK709ZBi+NQ7F7poeZhFAc
VJFtvvuw4qLH5SNBOX3ogaxoWllRk0/s7a9Z8xX5OLOyjPOw3DO5LI/PE3SmFZIphfttxfibD2qh
6OsYocFiRpZtEV84R9u1C2kizhCPZWkBeuL5/8+agMjLapih50AUMODW/vB0IH2UJNq5+IT7BHtp
Zmstex8Iw2Tq323W4SgQsrlOzaYvHg87fDyy7VG7RHggcsH/zrb2xkvI7vVJqE6Zz3UUL/oYAl2T
osOEiubGR0MAU6cif0leliAGhP2cXffpG9+qE/x/VJmrPmqIjZBvQylXgs+lbSOWUD3Xb9yuy7qk
wc6v/2JcFr2hvkHyc4E6xbDBUegOqTtZpMyvYRm3aFnDYhQ8W3IElGCCOYEelkb67EN6VRR/hHkH
to9V5h5BjBMJUZnBEClPj2NmT88XRoTbooR7V9oFYqPk0FxPg8pM+BgWAQ8g1XBlRBWjeKTfpPNn
dGyI51J3W3Es/HLY2D1QL1DlXS91QdqhUDK1AXE+26E+CJ8cAYZV333LHxgmQJ+XuT/IYLbh0rJB
i8Kd7/bvDM43mhoWJ7mQbX0VO75pnp0TcLm8IF9NfA2yFUSHgOqdTZ2YHLsUvhAxBlY432hD5Y5n
/pcUhd2OcUEWas/gNfRggdz6QmYNGHp6/P1QEdarKJi1Q2zT0mmISmeOAFwo66iEZGFqS047R62g
B+PVf3xxpnyk7HmXvTob1RTGB98BeNk9sX+SUS8/N+/qAerR5ox2LtAE8R1JdVx4g7jwfmEXOuGL
HdT3AYxLCd4P5rCKVTlpETHcYvmp5evOON35W1ZUsEHTG90SKX0qnGeIIqSxbEgXJdyS74rnX9qS
uPA3jB19z5uNJm50ewaULotVBL7CrXsDvylHNYDTKCve8KXENZ6VqP7OgZq7fGy7V0uoVa1GoXMg
c+WdRDHME+uAbuZOiytbsKM+yyzsX4mqtebWf2Hw37Etd6pcJELLpB/KwtSSarjIqanDBRQ657ns
KoghK6FstnpIcSrvR9TZOdqIXW63RrweELLV/YD/dfoJtZMOrru1XA5JYnp8EC0iMWIReOasjGum
u0yBzm0mdju3wETjg7C+Qqug5A3dLRLPAjpPU71uiKImsQm0SUoMVp0N9g3bKsjlsSr1Cdc6Nk5Y
jMi9UcWHfn7OtY721nZIw6YBre1/IwgPPS5oeT7AGfG5fXB3+ywX0986uE9uSjgDqCbIFGg4wq2E
cWusv4xFoT4tIkAa7G3EirIakCvPy8vYQ0QwAIZLuX5WbtxG74k8IC2zAIDtVYKEGBGC559OUnQa
W0I41POB7I7pCYNxDvCpFIdVr11aPVVn4vICAvkm5uIflTSnVlrBB+v8nVR9QKUxoCqfubbwAeUa
29YASx+AdMzzSBReBc3gQzKbU+enPhGWPJ0CUCNYAzf2mNckmm8BvEEt2shm2ZQUk2KdOvSrZ8OP
XKt2L8SEdaQlO9ez7m9bATJjdDv6VZeW37UW5OVKlqwjY/odpL7g4LDXT730wEZI9VVkZcWSXsxr
xxGjG7KmljFPk7MEo40WZgHvW69m4t7wIQZT+ntyISW0HhK769wRXfP49cWI9G+rxxq6s5bZ4L/I
SGqpEoVmPaRrq+cru0vhYepiDUUXAuwfXhgD6AfPx0qfu1VBEW+6SwLpbxCikiODZrjX+fyVf903
9bW/cM6lD/ZebowtNiv009hy4+Pwdo0dJ69vUlEA8hUqHxVko3+l9Fw8LZOYM9gpTiJpOWYkAWa7
lr7hUExndZOgZFQOspz5YL3i9OdlvRkeoJHCmPaCNJgKHvV90PfQEeuEwNcELwpWBH+puq+9D6Vk
D4ZqeiybEfDwdJ4mC/MsbsXCgTqLyNATNBWG45HW3iAGVApisrf8Lnhl88jyuOJT+s7Y1+ow3URp
BUselcq5n1lhygTlZiDccl66zgQCT8Etevx4C9fZSJgapukAl7ibse8jcVJs27YD5GeyTn/GIxy7
jPAk7AaUm5V3/C7op57ORcnF0TC0QYNUl4lQHX1t4N5rh3wfXLvjzif7J2UOzLc+UUHZOhGcHMoN
58gZZ7Hr8Q0D0pns3HSA3FAy6HpBKkPI796BIapT9RF1MwLOUSA/hYZoE48ePBMPGlH9nrvYomHz
y20+uvmaHNGQn/Ck5RkORaHtuQp+jXfbtkT+JUOnXNbwyNqXCVmbrYIvwOFHSsCNl3cZUi/+rBPy
oGFPZTT+MYnwLBqw9cUAouOlmJRxNvGC7w+7PfGCWKu11k0Uy+JiuLYVrK9COwgyLtNyxVQ50ZQM
uE8iR/2mq+5J1olPKryqbMxr9Ww1u9PKthqTSAuf7RHn0bUwn6e2gkT+SP6txZXj2gP0qDYyTmDH
M8fstGL/0+EkLTZXVkj7I6S3ZKvnEsOihm/NopGtStnVx9rGh0+J5fUrQNpLbBieqMkB+uSxuU7S
LUXIOk677fH1NySRVAeL6NSHhjhaJgQbgBhtxBZfbdU2QOZKaIsmSpurZGyC7//CNLH1AWQMBm9H
CaFD/npydIj+iTq81k1/JpzotC/jO1SI8rbcDEPkuuqa//g+VxtZ2Deddx6hGV7pyKq11fBGZsWO
yde66CYSGKr9Xj8sSdjsPGLntF4CD64cwPp8isPRMqK8naAZE2Icx2F//cbIVqIgHmvj7K8uX+7B
KmPX+BHByzWQ1DdLBxrOtOmt6gt2v4UsOPdiKhBWKz9uQTAyknIGYyWIZVzy0UDzVZcdFTNw3Dx/
D1YG8TLQC7b7poUPBx35I9zAOYrDIb1nc0ujfKRWKZBgUWkTOBbkY1JMjzFoLoACY+2h2k0+P7aA
/my3SSU6MeqiPrJ/2kK9bFbACveMPMiJh+1LMngEDhHwGHbbuUxlaeEpuwyTz/6BuWScKfxjFxVn
kQP4X12wEW/dKa/NVeY5Tp09dSVS7HFOMoNt++C9lov+IjNToChozwUe7TZeAk3n49Cn/RLhZQ16
PG/X48shfNv2gvFxuzZQAWDjdwAMGWquzUvu2RXXyIcavDSmbWCCgUL8KGvpUqoNses//HAFGlqL
GqROcVRBENVUVOFRCz1Uafayqd0NLPZex8HxyXRpI6o1SyvhBVAD8XX4OzWZ4nWaL/z9hy1NWeld
kHmmJDX13CePazPiDdvzIenGGr3/rk88wQfD5NVqAIzrR88FDixkObpI8WqeEcZWOqyB79W5q86s
lSv1pbYvUAYmcaUKtoJAS9+ql03yr7D5+XYq/Rd2L/ymdY9zXrYwu0+LpZtEKEpTjxCFCfRxT5ik
HJ/j1Te63VUBCyWYP5pRpmpyzUVqJwMfbEII9u94xwR0qBpSUwc/m6sQM+GuiErkr+u6Y0PIuVFB
8WDe4D3cy4MQEmINTp7NvvqMoFVMrTgAfPLB7fReaQom+dF/yUF5QnHhCzzGRbqVzsoyV2yYalrR
aBS1OvmF8CrJ1j5cGtFSt0VW77eb/ikD0JlJREeV/2o6+wo0ug9cawRD58doQQUHXQM6TYvHEZZW
/NmYqlUYmd9AmZYOWDfnuOYgENCP/URV5GedpKB+ocMrWHGGJx6lvU/a/YyCQ1s8g7cpqG2UoHS4
WyigKIdRK58MKTqgTWbaC7vq8/gQ09Vt5/aBSX8aayVZkVSYNUZYBUZiDr/MMnqBcYKKTW2n/OGR
Bb12IMVVPiJHo4AJwB+BFL7AwCCMg4GZInWbml5ecQ8bmw1XeObbk3aIcma85vzYMsd33DWqcy7P
LGQQ9v7i93X6sT0RreL7RZ6tATRgrM487YSQQ6WndQbCrf+mAnLDlnMyoInB+ZqXv5FNfjmjmQcF
Meof43UMV4ETJH/qo0CTcu25RnnTH/FgcJVyqh+tRlTbwVmqalvtUqLdQb9Uhpn7/Vy+J2AJeKOy
fpgo7H4GStFKywyGxT701Htzi+jrGT5Remf9h3zFbIWmInPON7ua6zUxkESJ3FjzlnJ9JOqsf1jr
czGn/+XN+c9WS80mfTYCqVHzwV50ZVdxL/CydKy+wV+Z6xuGubdmhzDYbv+WNl1xx5Em933/aRe0
ju5ATz6mIyL0yBHCJ3qLX7y+ArmdNsRivy5hkqCG2D2hzeaGm+0RHYbpW3mmfCsxvZK9/namDCIX
Xd+Fw4qGfga+JJQ+/oGWLq80vAv0Y6XDNc0TGHU8v/LVMjRSJEAGyo/c+I5UZohZH+LOy2l4VeGG
fG7f8z9C9TW9rd8FYv03CjatyeZ/yQm7V4lVAuvjFzbLdi7w2UcWN1eMK4DKI7Nzoxdz6hgeJNe3
etnyA8X+VAiPxN+NMFZq80FUMn+adUw3ZdH8yTH6hvgvAE2sDkTfdaJ9gA0H8ukqleigBYaNAEuL
uvUAwFNfOqiRa7wTN6OkqwbprpiuFbLKVErlY1w3zb8QJVZi/W7A135r4rkW76m8CzWFX+4RsDh8
33zQ4i5BJCY5lwbqszN1xSJiIBUrCC7aNIU9DOArGvrX18TgowW8vZ9E0XmysdSh9R7vfmDNqF2z
6Y1aWooTAYv5wWEhYdV6wVOv5d+keEAv3xU5k8dLmoYMfmTMV6j2KUY/gFjobN7LjLbxWUFU9Rg4
+AQDQyCalnA7UgSZ3sha18xTWaZ51sVTncfVORkz/inDACJWWr8G32bJ5ZypXPzpsbv0gXClzvbc
5NpdiPJz6e3H3G71Ygo4uvblAPOlLTNTldX+MCxjiM8r6Hbj3KeNGv15bpcgI5LBFutHJAm0RaJw
8oNLV9lbAikJ8AwA/D86mw9Fz2cvIUdzINvc1P5Ryut1fEH3g0q4fnndl0Mn3uPZ5nm1ySmVH7SN
vkKeK9VnF7TNr2G53RuUyLVsEQe1N2hOvjQ6z/7D8r2E8rLwt1wMrbrbtjMf3rEdp81iyXubZ0ju
8eG8fx+krWWY5DRnTNt0BO2TvyX9WRtId8UyakJJ9qoKIJgf7KSFLyQNVpjgWmbZyg3DqFpdKGpI
pX9K2tFMYOPzUS2OF4izZa5gfUoV51DObEEtSryCbY6aM2k6EAuUK2cFxcg3CDLTxsRPwNvmpKd2
HkJ3WQ8feLwHISp7FG+RoIPhuJcxRyWjTM2Fpzs4Ly+NgH8rEDMIa1DUE656LGwXIXRw5SnfD7AG
JsYEMs1QQap153OlWhamYUsuovDaC5GOymZ1O4BGqdu6jsJ2txmtcrn2wAf+3MQV4UNYAAyVSRD6
mpzqsx25unWIchCPj/x/akIIcjbcCr0cu4EqYYSr16gZ+gH658lAViY5geiCOPhyEcIqggG26Odm
8w0bv+MYhVWGn1VHOPzVPV/Eeb7mkqwC9LWzzn8j6QUQLrNuGYSHJ6c+vC34WeTA4j2V9zaqv0Z2
74FTg7OeXSDkAF43AAQ8o6yI1JVCThYzH5xq6gjTdjOf2Dy9Gv2/04QkUX67ux25IGvz+8ZOYqUC
eEcs95yJEetdZkiWy5dR5inZ2LEGUYy4vd04quYedwzokZJLxa2GGXRIxTK2cQAywnwNGZOPwVjH
dpXfNL3nPicwAerz5UQEsg7j9vz7YC1ko5T7BZslZEhMYZiP1xObaPDNTcoMc66i5g4rhIWbAa4X
wq624rh5kR2ddxNZz9Jy8B6DS7fbi5elQZMLcxUbHn4vgWiBt3NPjyjoEWAptBzi8Toev1TC3VQR
wz+b+bMoFfqMBXlkZ2Zm/EdH7N6BAGsyg6I+HC87IiXSFoCCst3d6vXPa4kvsMxDvI8DHyYyvkZM
LXxL90jpNCDFvybYnBwrJNi7g2dY7LWpXUSitReXa/TihRRs/M7EP6bWsSNgEhaDc5mFLKojmbLh
0T1C5yt3KwSKuZ1gg5OxOuu4fveVIvZwIzsJGbVQhK4h2gf3PA0RZHMt+ZBwYjSYVyEQejI8gcNF
ggYnYV/yTsurLKpf1FLIKgIP3Wk4glnWCn7kAEOuioGw6Gs403FnsQHI4CnpLIRjk9JBqnatXvy+
lrlQFGhcobGCWh2h1OIJs0c2iEJ/qTdJGXF6JHuY3e6IN8iabf1R4J1nwpwzNFm27J5mYa8U/DQB
m1jD22Cyfxq+ZqIioogqC/ZAGXOWVCRTN4OBX/Ws9AlndGcWCZJozo1PT91VhOy9zMz78cLi0mkl
k2wOjkbSQWkgvT8C8X3xvrEEzbgGN6eDRMCdTsZiZYV/1kS4xoj05uFRzYyCi+WS48bb4vyntoa5
of9pI3eP9Z7kR1RirN2O9BWPMce2cn9+8tNFBgs18T+zOsmIM/SQTRHkcrIVoa8VFuocUAedHUcv
RjN+6xkY7C82oz0eFjGjHjNBwV7T+jeM4nFSkqwO7wZkgpWc8WtDrA+3cOG+igeMMsNf6n1MkaSu
O9k2FmkcQ16XOrQizN6dnTEsKAS4eV82kQduC3X9PyqLB8ykgPckQPY/+/5GOE+pw5iYNWPalfEC
7x2xzXWLzBFi76HG+M4FOokP32chDR9D3PahhXjnzAXgphTJvAL2AG+L2/yYolTE/SLkGclQPRCM
/Y5vPJeaxRmQEOTtPaCqT2NTEVdOre/TXyWdLf8FlTeB0OnKkihvRYW9xw4jyBIhsO4r58W6B/nq
nwNrAY76wdTbrvnBBEV0TonbU56uBuMzDttJHpOtN1csi+AZWWZybzZzMrQnGeppaa+6sBtsWmLs
onOgAjCrdwUbjCNsokv7AwMiBo0RsFTEfzEh3xNaOxOswxQYg4+avBG0lFRykZWrdS1YM4qDr5xU
q2WqHMXV6FL6vUKE/KZX2SUvYzi+CyYPVMucHyBUPcWU8K5jVqubSYMV0kQVIVAsdeo+Nm+RnjD8
xx8SUOlryCzICtb8na1RF+J8n1O2nUD/rC2wpknKBJTURtKGYwXDAQNT3jWtw/aK2w7uBVGw/Pul
dztQ0t8fzJ3/2GICxipP4sFIdfXbI1Exu/tp4JMzYoSah4MsdfY303MHDpJTOka26KzSLRgAUP9x
BBDHEV9oI0gsFzPei8pVM0Brt5KyhrN+jzrjelFGmtgdpHLGRWn2vQqOo8Pn2G0dZYf0m/rdLTDe
e+1PB2oogJBpKszIvKoGipAO42FTi7OhwtHTqrWx4ynzP04f3xEEzr/0ScSByGgSCzpBt4x1heBC
QiIe2Ci4YX8n6R2URDO2E3r0AoyKz3QJWL4GCc9MLr8Psp78u5RIA7i7KpbAKeswTrxzjXBLqPio
HyQ1bGJAsqLEbhJYbxZ/foGGTg9sROzEKj601yoWkNIl5q+F41Zz0oL+Ql4sOXPrbbtl+dZ055A2
ajp+bcUs/18WfaSC3+GCZb8a7COlTJdhT+FaCVWXU2og8FT2wFN5WYRJQiG5BLT6M41JB1zfn8WH
NTzUaQMNRNoccnvK1G6vkD/65/kCwAgUB1W8fyajYTqTXdHiUeEYBZNqm1cx227B+t1bTx/gn+Py
mRFGrQW05PD4Nq+ha/qAZN9F5IxP22gUsfqWDH/ddsp36Bib/S1r75TrNDK3S21P19IAtfqCaHSj
KXk7yWbCrnGKMB8ZgHgBwH1WnmlDmB2Tz5EhGgpj6Jwj+YFiuXG8RBz34dSGxI540/Wro6Trj0fl
XD0ctO0JJ9oXZre1E7O7IteNzIDCMaAdpT2Mr0z0i51Oywgo5LWq+ONlUvrENwJUCzF/sz/GZh02
0B4QioXNh/EPk1e9IRPW1epgtzTV/U5393Wcv0oJtsRji2uRl6tLM9PC499bFnrAufv0M+uO6qPk
Rc2NuKd7Eu7kh+gaxAB5qb53/r+mcFfDUf1EcpSvM/CSLCpz1p0C6evbc/il2pNlVRwm2dqUuCsw
//jVeFWcNw9iGABl57IJKjGkKT2As81C8lQkZg6ERgB0UDXsd2M4HYQIVYDNuHdaWTswzaQWRy9N
+WxoCbxhPDjY7WQnr5e3FZ5K/bx3QtZxEVnlc39Lw7sT5VgjDkE4nMwcusUvU8t7gMb/el0MmHzJ
FH2rcFTpN2rhAxKJ0/vATTBMzxlh+SqzLN99J6YxfMdKyR3yD7HR4LVRUzvNjveYcDhCcX7pmAl5
h+DpXri09pWXae801Mr5fnqqaNMXQifTjyOYf9XWDiJmzcB6KFnQTPQ7vmtiuKVqhaqFUO+ZKcw5
K1HSsIYbHS1pQv6XIfAVq+cAoy/qbCwUoDJG31eI6vmfg+8U0ZzWrKE05/pXZR1n34pqBukwdsLm
m0AVhLcnaDdLcEsEZv7EKjHhRjhsg6xdgtcUt5uElU97z0IAhRn6h/hi7+t7hP2K+3TM7xGqhpRO
VIMoSrZNpFO0x3Phx4PJBQYzN8y1oaQPTM4RD9gmM69exYAZMrK/Nq2DmenVZYYju/5JYuSlNw7w
0BywwrbJbw6L0jYPem7EVqkeMKlQhfRdUyh4SU7+h8ml9BCJaq3T37nY1Lbz2M85ht50zcGviBSp
sfauBQKWWnlTqfvd7SNRSWOc9IFlq5f8/k3XLekq83KBo6Mz/0hsi2fMJBJBoNNK25Z+tmaOZMOJ
u3fc1mgqXn9a0e/vI3a2EhlwbLtW/knh2hSOdBfL3QWbLOr3Wu6hkRonHy21L7SrjwMCn3aT3aKs
8aht5hGmjj07cyl4xSQJli8yaVDmxAvgamhpwQ1ChdlDZJlOq5rDZ7PMLBXQ+CAxp1EkjxMZw/3t
+iWwU5MRzH7wG1O/TpdApr4hv60DxLr+aN/BAYWPyKg8L4I4h0CrZV+ybixw9WP9kLRYJ3bLndBA
6NOJtSKa4KNOgJNFHkPeeT1oJM3Q8dGrR+hFT6kvM3jUYo2vuNIlYxLpaPB6Y2/y/HcCFmNdWe8D
gKgnXVVwF/dVADwnjfFHyG+5a+t16fm/swptFakWfw8O+ZAkvz1iSqiY4it0FANAt3vwO/RQoKkj
fErmwi83OGTVAsTpFCtYQNvEQWJwk0T7o26WsqHypAcVfMU+dKytEgjEdRv5BtNiLc6Qs5TRjj/z
zAG/iERPLsVoaDgkvQT60unLtMOhfT5p/Grq1PxX0fBzvkkd9YKb5elOME9U2UQ1U/oddVI2SkQW
/YDV/8z8fb5J3YUlNSbF2TK1Krtr0LWBKagDQrP/AtMbYVxsuMN2SRJMcfgvUgLoxKD+10bN9+23
eDW0Xg00K/aJBgUfeTlNvihx4kQA997pBCICxNYI4tYMjPWGm1YRv/q8k2YPA5hiLTXs22/QiLTn
D4aZLJ9lAMD4Liah4xImYe0PAfkbY5RirwUTYoru2ouD67CXibjoHO7mbkHCBedsTDWMOZiH7WWs
xMqfMBtll3h8cf1kSMckwvC1viK2Z/p4xzFkEkiEaADWT/KlzjMAl2SW/npUn0ta3XzWfsmvQDBP
wAbADOdv8nynkTI/BaYkqP8CnkMqu8ve8HqIfM1lbu7Qw+/JMwof4XRJwGrI+lvqtyznp1V4VaCR
ci5ykygPStXDY4NpGu5Y8SNYn7+7HZKiTLx5R+MelF3yvWoIQU86S2GsDkndibAdwykCqivkskdp
B9tcFjG4QEhw3EH+cNKhRKptVQObdEIjtoSdV7PI5p72LcTT8/rIS3BRXVjvTomLLsVnfc5wTCr1
kiN+x6BPqLGdqpJEvTMyV8wU7lK1JP2EDLRcZ58nK31Yv+MIlGijs8F32Sap59anvNpjb2kDBHNS
ndQO1CtG+RQ5uFA2ESXo+mSSlwnuWJMsZFdd0ECEj9jhvPh4BfGXPeoj8598Z2bIlM6E5rbl6QpY
uZQyCklomsyz6JoTi3nxsMKIB1GZToJ4weRh4VKzN1KERX4E1olP4u3GD7Yq+lJwh8C9ymsRyKS6
vobj2//2/hnKGTq/xdYo7XQBZ5BqWdtsUB5vJ4NmAZhfUe092/l7YfxKW+Ys5ZqNiPY4X1f/dUG9
SrG0UVhB/sf/gBxN+jdb4y0LJcprqeSOTdrvLhahPg5IrSkRJCd7RSb6AsRqXDrkxmRQcpzb73bB
+WeKXnCXZSUgqbivTlLWcgijn5aqsa9+mW5uiJxpEFv12C6HxMPPkxL3BI4wlfruiH94HsRikJ0V
jqvELT5revJl4di3Hrd81Xmumo9EVe69vTsS02dRyvxrN7chDxoRNBFfn66C8s9UVxwonEcEol2C
89Vp81Szthv53oyBnZ4c5H9vKqwks7WqaMh/v5bxHyvSi9vIlPbxTIaKto901nGg0H8WxVlOwzFu
etavCeTYU5Wdx08Kbxg00U+unNUOGKLGiofysAO3zs5fIn+OEEuIXz3zMST7Hy3lC3k3H4J4glxT
LG+11JnyZRUQKiqvAI7RoLcNWzUbib0wB8JWk6TLnic7xlz1lgw1Wl0DXD8icPkd/DQRfSkSF/uH
aTYtefEylQHFRUOhJMlXK7caFC1mbrBcbwVNsE3Byu2eKC7VzFM5QvBoGWEE69kRWjlpNAV2mvYv
KmgqMRpqM2VSiKGGBTZHDWa5Bv53eJDaSs2u3dSyDoLgN3Awk3gZIEXHIVi4ANyT6gryNZmgM3ks
6V7aY7cl/hK5PwuIcJju1aC6Fdt8xNq32vVKur0jsiOq+MNTyzwIDzOENd3XcmZW0NmvABeM92t3
PucVSwH79TYkcVCQgIxWaLNdBk6FodCLDpLiv/MFKkQdQgQS2s21+gXX6oRMQfitVUaivGhm0JsP
uTRNoI2HjRlfEn4LPiN7LAeJ4jHg6c2Fc3KXcguahrNvsP9OihBvNcuMBOJ4bRM83SY5ohkYAHKO
dtgYLuyYw9kFId3Tq+7nm/MUzictw6bmjesPneusp0El60xiHma0sqHaXjxQpqU5PfukSxCg4czn
IK2QYZ+zeHnZXQV2q+smx0rNDq4pe60kmfYHo0fAlIUrxAvlc1DyqxW3SlX6E+x0e5edYVY2M4Wc
P/RJuTSTl3IFKPuTvX40VyMQGHX0r7AOQKhWaPuu/sELOini/LI18gHzJqHIqvsj60v7ye0yC+Ll
eW0iVoshSaSrpjMpxiF24cSefbSr5uH+qOzC/NTXt4a+LIidrmtslg3j/0jDAak2YmP1a6kUvHl4
bk+8d224Xbh1LbtB0NORuo+BXhpU1OHnDxwXXsTVMMRqxxFYjYz6MbViZS5ZQm71mo75HtcMGH+u
g0XHV4kfUcQI2JDA+8zw7hnuZJNWRF31uwqTpTBg3wro9jCkJSkUTUDc1A/z9dlbrHpeEA+zWOPx
ztrFpgxUjagYkCNZEGioqrh/WF7apgAKrw+NvOG7vG+35H29OJKX163mCWg8GRrHx/Om0pMK4aWs
sIezgcpjdqqiPDK9pKkjnRPEjqhLrmNGAubZpytr7aQMZzBdT4Zhr10KDwl6EmU0rhnoNScQwtAl
e3cyBVEzFddlW3oiuIR2UgIn4Dw361T5NLriR6g2zOTEYn2BVViqSyMZRmrgYEMfiEhsTb0SHxLb
v4mqrOQ55YjSsgMzYQGt/YZn4Ybh/rJGP9nWB81ytWhqQj0KmdI9WObvuCIvyqUN2IDwHTOcbqeA
/PoBCxpPLJagb6e81b1mSCKK1nEv9ls6kyDTiNwuxFR4Jjy3TaN/flee0nelsQOQE0XU/7NAd5LP
tI6JqKGnZq8l7rv0bVpmZBawgwoLCG4Gs/OUK2YTKBurpn8JdjfBdw1NzNPPBMV0KXq7ve5ghYlG
T9ntUm7cjaELTky7SmesiV/8njuumZSYmcdldF73XYqxBUtkXrr43C5K+z97sNBs9RtkoO2NGvmA
0hgzkCwRvjqIaEhLHUbILzkxodunj3YoTsXyk1cV8FNw3ejQkWu0SaCd7yUE+P+lxgyxx7p/A1q4
JivXtuQz4rQAwHHFJ5NMG0qpU7lOMATzCxLL+BHsLRNKN+66WqtCn1OqHw9CIF9N0Avsu3EMrTs+
qvvCMSxVg4IsPluJh7WbwbPK3N0QP3C8AGniUYKGGf9wc3mk8JVitudNSjlhyY2H6/H7SAinaTsa
juh0TM5lSb6PlMniistmJ5ojgtZeSz+Ci7hgaF5rYjtSq0BflGZlowt2FsOjWGioe4n57HeXQEUs
jeIwf8yOzqlt+UjTsAcGbbKtZh1KMQnVgZqDh5/JLHu+oHjx7Sf2GZ/rxkmD5ZxQZXafpt4E7yjw
E9fT+jpjq1pGK7rvgqIvewKXJlBnBXYSdeDxs37S/jKDd81R9j3R7Nbp2f/2AYrrGztDMOqIh5Z/
qQX5cxmbYT6jtr9V4kuZbiOfNC88VBwczn1IVAqd+iveyfQShDF6NDSq2TX5QMthhDLNK52xUwV2
DmBhH993r21S0o0txK6YfKmxLM9FMGKCOpY6ZvNw6NzuFbDK/rWVM7e0ppxT66Dr6sZ0D4dbFKJD
leaPim2bRBUZiGojml3YFjkBgDFVBYqW97JIbNjByT09I0iK8gNp+xLi0JJkg4I6n544Uzl/euqZ
u7bXSgwYEil7HCRsQJt2eyZtYVwo8tJgKdpmH9bKh5vYR2n9AiADqHsTPj+XetzgmZSd5jpl0Y5q
geO3pd26lX3CC4zLbQ8VugNHjNyrU5j13FG5Yi1xFtDYjfS0KiIPcDlb5w7QIQL1ciBFUrvoSmCc
t7dZo6istMbuJsVsgLc7FBkYrvYugG1kCRKx2NPDbzb0KA4myQB7qrBe+QE7mdL4N9+1CJpX56Da
b8rF/5pPoCY+r/2USwKIeqLwf3QSdmnad8BsMBfeZmeeia/nLxzt/HKOQq0gq1VxU7Fwh229R2p6
wYnJuGIb9L2EcnxjzIXd2alIlChte1CWfOtujfDTfLHmk4bBd5MsUDyoMBG79DdchKOxKcZwYoRV
cG+2oodUFsZeu7GDcymd+pNZEo/snENGzt5YpEkhvRg8oCapknCOICOwAA5DVP29UT9vOMnJSHYP
1KCjhxJqE0HlWo2gVeizN1w5mKgun4ACRTO9wwH10jMwLJ73OzGifHK5qMkS7TRJHbpvnHjjF5f6
gclEmGMRHpR40TQNQihEjgt2tJ/SvjqcPJqRknafy1ubEu8PdfyCl3OgkV2pzZ7x5F1TUTy8gLSx
DhuWqRvhNKTPrOEWaVjKJfLV8Yel0FWU1JYbylViD20qAaTGkEJHPu2cBJnmDCGBKBHcFcReKMfX
S2tTL10+uaz9SzOi68SCFSUQhIGoXH6RHusvpfr83VWYdwJNpW6eoiypk5XEz9MEjr3080+v+oS3
yOIu3V2kBq8noE0kpjCmJcBOBGYZ80CAO/5NelhbSzhmK7T3fGeTEE+RizK6l+nDtejOzV6PJCZd
G6G4WanKs57iDIl9EXXKI6fzAbIS0xOe5tHzfUHmybjN38HjRTMvSiSF+yS8aNjAGOSQMikdYcap
wSWc13FJ53N4zT1dUoTb9ESzQXcIAylQ2uPxG77qrhAubzChV+9+6Z3ODy5F4CxJgJ7aWZSxhOkL
6UfAHZbYbDwwR6emf92q0tKYq6doa6eRYAsFvhgkgZlJeLX9cTdDH8gugyb6lez4xioluPriHAZr
KRqwK2tId0Z+EHzTcIpbD3/r/xLXI7S1F+p7/F714/iR0+ltBkR3h0lmxBzNsIqebiYx+71V0oG8
gLhrmxRxnkNW/r/OPZXfDDP841/HpEyDdD+Rw8LltkxuVBhk+KZnSsIuhxjU+W4FAZ0kPG0W2gdE
jX/fVc26FCpd3p/bMxOkfxOpBNEscJ/i21ZCfRC03xIvPkVmvNm2mECq4wIsjxVt0Q4elaXck3au
KIIABGDYFaVXNw5vjeJzi0MZCNXL0cwzMjdbKxUxemPPchChfMEFtOAUgrRV/9FDllRbZCHFvFvw
A3Lnp06lEq+mqchJHFf7yp6QQLp5+HD97MhOzM361H4t4XYnj/jnMa/vAHiemIH8VP6SZswoAvhm
xmGlpgD8lzZSuyKDf/ktiEweKgJX2O8q5tZG6V87U/ni/vKYfOZYNuNY/CLX2t0i28yZNczvaXta
FlYCIfs5jreKrL1GeS1UHsNQXXYlZeXRCXUNxowY77xKRJZBigEXYNcQBfaf+4+loLnw8krdfshc
Xi/JrRBieL2LlhadxJNDeggwadQhYYAk6dEWrMp1/fDqnpYTod7u8ktsDjPNNyRipcdpkZmPst4y
SCV0+dnVEP5GF9sxU8yT++G1EAhOrpCYJk2RchdIWifjrnivfv0a3yIf6/JPyDeHN4TE6m6fd8t5
Tzn+a9paOYkBk2pgZnKSMyChSQLxP6WM0bxcLmgG8PsUuAsYkqXwWsdawAJib7xEs677OQRRga9T
LJiOLpxn54lQFbfPLSZtJl1o6kB+SAQZILNOO5W9qz8E6c3aN23my915PDtkz3UBpE5fiyABt1pE
7GYB4gQEcXJp1UoYNxU8ufkVVFG3V2HR/vUsMGCo0AQDeyr+Bu9+iDy9c654KnkSzyBTHB+aZbID
/vsVjfFvxbWGMIn5063YRs+Lr8kOGdKwXoW85RgSnw7tibiwrb4HvrB0J10OuXJ7zURgYZZ7L2Ah
+C1pVxYNPaiDSWIq/zZk5TfYOpMyQwT9krAn0TBAHI2wxKqeRBU3FN4BV30UzcnxTwhgtIcBxvFc
A1P3iLXdWbbIvuLkoeb/5FV4bqD9jkQk4fPLXif3reCOuEqr5agHlZg/JQ3OupyGAT6zuwpghKyl
KEJvwlA4nY7gG2Vw3tspss1MWFwCENaYsZApb07Q8QwwnCgxtA1V3FW1fOTAcCXSKAqtHulOToFV
4yYMkxvAbgPrG2dMDll+Td8RxD4MXAXKv/cmG7DOVyFkaF4b7EdFkpyEqkF9SxbmwgWl5JlnqW0k
61VDQGABK+YF3zs/qLtgca6B6YTNnGM9f9WnDOjNuEAtS6T2tWiY8ia5Oj7vzbuYAMf8HxjPWOqj
xz4oNdMx3hRt5ognQznOP42Dr0wCdT9/kkmymIApJNdz/aA6RsrYDbOmg3813X5qAVF4tXSgZHvg
5q/ic7J4jEsKW1spqgA2riI7KvR82XvOXQ3ks05B+WSZrZYQ+3759D6G+UEveJwKE8opAyVE6bCW
9KAg5a/Qsspp6w6QdxBYLUxCMQGrsiRKCJ+gfSPWfi2Gh189bq/F4xBZfbV/T2JXn7Dy1VqdaA/S
fAjHcggxqZsd6w0xsF5Fsrzu04Drsw1K7rmwESl7xwrprvoAioQskNSnn5lbsOVAfntsYIgK+I5g
wwjl+/GtNaHIriUhAkHuTOYVq0ppXieNtczKWhoHZeR4eW1B/DXf7/kEWPK8KJPNvcEr9bsTOXRt
dGOBj1idW1GljyeyAaEh0RfenuHfnEJY/C9QLdtlvad83b/KCqU4INm1npsCHT6jI+j0Xs6ILhD7
dDAdhVigsRxTh6reOt5k63/+qEgDTOyFcGwT22xw9ThT2E40hRslKAHxpYByd9xbqIr2afKt9uj0
A2n7paQY+4AYa9LVPrJEMwLJOJrpnqL3bhsMeS0oiMe+l6zeMcot49nPA2P38NaHx6MfJ8iauIWg
hejYiG+rNhj0H90dnQF/KFeyxh595YjphPyplWyEl9PlPQnSq7UFllwV/7zBPIutSr+NC/Y/I/yE
08Z6YxU5SLK3r2l8h0P3Lw2M7elS0Gp/UhKi4BmKZDGt1jhMwJiYMnAS2Fo74UwOkU4AIPUo1kBu
NcUPyEQ2A1XyRpdDbZ4yRTX5WhJRAc6vxl/kGwGYA1hdZfnbt85P19CVU6jVApMOP/OGhWnuDR7r
fTAveceweIqUkq1OBSNuCXGpZ8CaaMmv3oRBtYaPVeple4cUoOuxC0GHG0aPn+Rh7BNIj5cbtGEL
ccgTVP3jhp6dzMZmu9DC86OMka7BIs7OQ8CRBr8aWYwImnosf+Kq/dVjWVX/YTogvWDF2vR6ffQh
B67HfQ9MbIpq7WHQqvzyEjuntRVW3Xzi7mFfm00CyWTmAxybG/hW+KgUEp3GCE7AEQilAFtg4vVV
LbrxzF/b3VWzFnxCbyqOrkyj2DXwt+37PWF1b910TszJ9DhwPbsg4hUo0lQvzY9N/0rXxgoGE47S
Xowpz6iyfFd3kjNEqz9ksVxM1uKt9ICdZorJiFdj00g7ScpfJJmYKE/kPt/GoCMmDJib1HfMvDS2
8/u/kEHMHYnDK+sZtukUb25AQ6pmOanRAWbn0+/CYde8WWSkQHPnSIXrTFOj662qOGD/tnZPt3Qh
AE8SY7pM9wVUAtMKBAXS4rtJNIqmHrZ88o93MYkoGcic2VR1tCuYltuMD8BcEwdmUcV0htB/yJnV
xa4VgUh+hdgSVMtjxRxuv4oHeqc95E1qNNao2By51OAY9ceeflT9c+uF1DQ6GEnL/MvRpF8DbCsA
pYNDobgqAbh/IWoFnT3PbUy8K+qNM5GApu+LSO03XlufEGDC5cE7EpgvKinMLlR1jXZNQXUOJd9G
0x3drJXR6byM43vFJjJ7RTZi2fB0/e9qyAd38sjQa3dmeUMXOeCf/ybPJqSDS5qbHsY2+WgBOKYM
uQaJN/eKrRUR3kqVmDUXou+4qmsOXJL6USwUaNKaKQQJz72xMRhLsK6VpsJDpvKxNSOGQ+d+K/7g
8lBc6ouPm2/Ge7a0HRbz33EHe0V8Pd2qNSUYvgjZV8j0PYlRN6UbED1XyIaXi4HsZs8K6l7emFFO
uAFmyRFI2P6rqmrOyLRzyDaWabZfA8+OjAKwWDb6FL/Mt2ByESZw4Pa/TJTBEyBjh7BB+w6t3Jqa
5S1gpY/veaU5LwiHmT4Su30SwFFwgSoTTCespgNS030RRhlcJel7HHtvXWLvk4mMle6tWvnu7gQP
FOVYJxRmGwfaLyhnZG65D/0ks0lGLW7Tw5wK6VP+2AiN6ckyM7x8wVJpAVNev6MaMCy8nEd8sV/o
oY85DgJ7VcAn2scqF/GrB29Fn/WwgdZ37h8nt2/nlyn2gVuHq54CBlSdF8hPD4C199Lee7rXQZXH
/5ugPLiOH7p7usW0Kfk9jIUwEftLJyusDIyFgH55qDtiu1V8UXcDB5u1Qk/Q7MXho6SONMh0TR7a
E72L8WwW/IXq8Av865lVfArvh6kw+jJb+O1gsrK7Z4P91qv9V90hOyiAQh2gdpcPLvTRbgxMdaRl
U+8erF0y42skBjy22QRorsQD3JhUnad9xULtIIulen92/ldHNlVR26QtIJMDaBuh1PKm4BIo5JjH
5S2oxdCNrUxW39q2lHWDd2Eb1iiJ6ERutay/0aunjXUtZHmGR9dlLPwqGnlO3MEb2WeqP9QQQRg9
/yD+2/oQ7DiIMjrhgEhVEsvqYx0OBAVU2L7ChGLVsLxq/6OjwWHdxB4X+X2CLDMLiwy0qPIvLW+b
W3yBXyQ8kMZg4YBHNhwW0qhjFCwfghgYa1Pg3WxrwDcQ2TEz2IN16cd2SbXF2Ti6sGjT6m2M5fWY
FnmbvjNrkbz9EgPugw5ilAqhoLqiEp4uErvQu5sD5MNnM2Neb8x3liZKfrqL7G8SEYWx4w6ZnjgA
e+kOVMl5Eff+iXd5Wglic9vwwhrfPZF0scnUgtAo1BUhygpc4q06OQrU54oa7E1cxIdAUp68OyiV
3V4yRy7Z9LpZZa9hE+FndBL9hekSTNalWUzcMJQPBCHo6t/wLk5I8O+b8ZJbBhMBLNSzm/Ixql+R
1kft2MxcObYvOw6oBwKBPTuDpDAH3m9U1c4dV3rSvZpstLoxGorv/zhLocb2X6u3P6lcSxU0O+Bt
gR5OE9/7kzR1eR0mx1b9W8/XXgtv0K3nuD+ll6V5fynIL+fKKsPM1WfRI2KMxwz6v4d8UeRB2B9p
QeGrnIn985b2l8kR62CUMPEO//5yGRPuPRiZ5HdHHTLZcDAuhOdaIVqOgmjg5kaHP6haHxkcyYZQ
kNncgYazamFAwpnCBtfawvXVGunM44HiEDZa2BT4cD6on434RiEE6pWvKYSLX6uOD6jrW9Rb9Q7k
4/7sQ80Z+8xAiO73709kFBW9/awGzyqL2WGCzouvsOvrte320KVeXkjxt3ip/116F8scgvLn1kzt
cw2YqvMEpuEOnTeJ5k0YfCU7xIaXI9ZU2D5hT3ZoNQvn68BxlO72QrSLvOiJG5zUaJbosGZzkPAs
YAdbBFOFpeCdhgytsKcDn6YQtiMsb42jD+qEHthdHGeSBwJ6ozIhujJ7kPQwyVlrGEjIvcAuGVGW
tE3N3pfrteHl7grF7Nqk9Hc9XgYCx1W7X5V4hGKmL2Ok7JxQuEvUuFlXF2fPg7LrOZherPm8JRsO
TwQVgPVByBoPbZdsic/as2eJ6EtMZh+zSocATFYY7/smD5zkuk1iyWMBkePEL3m1i2V7QAlnndmC
+M8R88/CGYAPNaPJYUa2JU1n2ByaBKaPXCYzfrFKXPVgFIG9sQg/sFWsG7Q6NZajrYUYbmtS7mPI
o+E5jsJ6Er+NgbLEkrr52kih6SpecOpK9TlMDQlH5CWbTcxk2DFiNpFA4936Uak4IDklvYLqQHYy
+FTzHAawkvaxRiPS/YLiO4rjqC0b2h+h3npEIBcalgwtk4FBb94nPtNGQLlpro9cD57x8L4io57q
9GEPJ7vXs00drz2s4XsSTwF6Nb15/uSSHa4tZRngZqfpB06/DoyjmnfF7E9Eo8jt4f6Cf3qXxAIH
OkLPlymLXDS1mJhq5vZHp2cTaSKRS8VRBXyi+nZzfqXkbyVBpsl95TQx99bFXM5T2L5gbPQorwya
LoPToDdqr9GVBYfxvOYNUF6wKO3vFedyDgFoZ2KEppM9VCjmJw1Q2GFfdMECnLPW+PK+8vubPDO+
dORuC+/G1/V3qYMmjrzfGs0ID8W6dziqj9ENlIW8asFSErmpQfGA8dnUxLuU9rC6gLiiOlxPEgwu
U8X76axtjh1+cj8uiAU+oTQLMP+NPmW6j1Ch6XsUlLwG2JOGV99sYqJG5GLb2sstWnivApjOEpxL
urvH5h+kHbcx7zYSsF9L1ILCBGJBmuJttoNRdHo0P6bWBgDE/KwTh7gdyZxT8mX/Kr4/JTDvSGm4
jTkttABwqfpLH1ioJXrR0C0cZpq9EtU3lIEKXjFKuDWlrdMAkaqLOQ0aImd0CzAd/CGCmYYv51Sh
e/vOgkfyUDIAzlEK9niLO+aVBpY6HZFm128I3bI3m/1w3e+/z+vN+x72Lg2LI/Qhc7WByZZTS108
6E4/DfrAvfkGszJ0LjEO25MDEputf/TEVN1a8RFpTU0GGsZtv8GRfEHUQuqY1MrUDyrlRuQqa6+D
5c8yeKHfuuOCFHeEtECfjAQGJVT30V0YF+ZMHLZSMq0j72HxMeA/ILt7NpOa/vJA7g5CXgHRb83T
A6m86KVOxA9a7Q9zaeh/qxiafw2LWYADd9XjfsxgzkD/ahoeuEnfYJqL2bT1WI+A6nMMVQqdjyer
F9vpKHHUMVvQCqZpn075kmTEY3F8k60U84czZCS5B7C4AhFm6rggD73C69HFHnNW1i9hzn5S/Tx7
gEEy82t0O45dJiqJt9yfPbzzhxRYs1tSRL74TSEphIdw9W22HiHiKWJiunc0zb79SBW9/Q0/tcr5
abdDXSWUFBA3N9FdRTvRqN8F5OeBDcoYN2jQ/2pC+5v4LCPnOhB5ILOtEWDlJcFIRFUSiYf5nfl2
WQLYOkRsEvFMlxcM/j4hZ5yixDiUATAkpGQWY6NR0IzJB6i1GVqR5ow39vrg2hRlWnO0hwW1NYZ8
Kdvb0VGsQFlGSN2vel1NzTBw6ULVvZD83PmZ9unx30/aaF6duAthCOblRwGUIrzKDY6RgbKozSl1
99+zpufesMaVcsG7Y8rsOF/wRGThCz8YqRNyP0x9sohD1vgJo6cDWkiVT8YyupRTa9sphFXcWAiE
Ah2cK2lnT8RKrzO25owtMFK1KKa1oBJIOPesttkFGKtlNWjSh1krHzSZYA3J17APZpnRMPelgB83
WA3i/FjLnpvwcFTZaoLv0Dc1uHPawQ23mavPY6AuQxqI5jAfAusolthAems+nXfjCIZc8hKbVxcI
P9x3ybouazsq1R2hABIhcfSPqTD0mKEldf3LKBOGAS6Lv2yHjtiDdKGQoDK7hA1qwybsfMiJZeaX
pe5ahQRfhuJ/Napn6Pqex5Fo20P9R0nDNa/ONrnwAAdy0+6f+VeunZtG716MCqWzrBbcKW1hkf3I
P55zSzBSAu9drBPOa+cfkTY2VtqP3F7NhkPmxQCT5YnRxTSkk1aGzgBBVWvHMtyqsI6+4vZXwV19
rJ0gudOAk4hr0fQA5ycMwenbbqDtxWuc0092OniCJqhlUI8MElsTv7/LleuMKIG1YUlxpB5YK3fP
Bx34BZG9tic3M/cgJ1m5r+dgRxaTLzc/vZHb7uBLz1i1Pl1zo5CWk0eT3i0J9xI+1v2q2nMTCFIs
YH5F74XBXzGyhifaUhw9EA963n1wGlTD/dHoIyh0v8Ll7++27xMVTKm3K3GrtSoaFqx9PHGyxD8Z
edJxmoSbEN0KRxXqGzTN+AKhgLRCNbG6ST4WOS9AWrIlJnYhtE+bhoQX33SkdyYP3DamGVGmSdxJ
NceaJ0JNLdyMEUgOZOEHXUr2LPHl2cNePXCd0BgpHwskkGBbc1K/kyXLFk6cF82FFfmFcIg6Ko1/
p2NXBzwYPSfUj6RLLNjeXS6RBCKVQnOYm/s8RKANHUzYi7dWMXKoWS9cs7ew3SJmLfjfNjzqp1MZ
Ibv9nh6GyhENdqQjdgN2a83dxkY2vWdPF+vD6yFv2FbiSqpX73WWIbjeY20FOAA+4P92r/mZ5qlq
ErLVlldevebmjtUX5yE18xWdu8yvpH05ZXgG0uAnPWThet8PZfE+B4bnF4GnQkg7Zse3674Hb9cZ
vpdL0c+JZCIgjboMAvttqLPyATaVsVMG8BdzO936oTfK675gsLYmorUcREKeZmxBx1EyzFaW0YCk
QDFxJZ1RkagY6BpF7n3PBsBC71hIYgl+6p1BOWkj4yaIvktSSj+JVjnocVi9NlNHWWk+6RqNlxOU
WDqJWaBxh7D8fa5XpRjh7MP7V5r5GeBbeWS57iNWMI2R2TxPRO+WUCEI32J1EGRz+cy3lNwUkFCc
pV5zkxt44qWfGgaJJ6q6xbSKGk4ihwre2EL4lhzoN6Hot2n5r92CFhFkRCeBhFqHYW+IDcFjjzsp
WC2B62vpnvmjIeRfxHOahSnnQ3nbEisUjsJ1CkXj9PYF8+zGnQ9ItuOMTi7cSxaoiKj5OODn9qHZ
yVUaQu4li5nCgL6lNsRCZNKMoH4i8qfHsYcD1QRim0YybmrPVnNaDfpSWSHxXmRmrNfuIBdHVJCc
tPkUYj62XRp7EpD409I2ytY77I61AN0O40ECB6MTHn4nHRvvFqBJwkfOvXuGyd2C0bRUa6M9MztW
Jqdn6f0goL0mXdg7WwZzzF3VF9I5b9my8ZWXrYN+f8DothYF3vXvfOKxjYIb8QkSPUS63EOLXmtc
aHAZMPqq6vApHxSC03vau/6RobWjbLxkSTVtL3sFrekShMpQh+r2CVL/2xrD3Zpyv/jSdnX1jJFd
7spdYVxrDfW2dBCBtUyWusF/OnixXH/imvnKFq6zJldQmYSMtOQMVie5Vl9hNG6x2YasE1Mrn7ak
Z5nYWJmRoEuW5vWiGSSHt+h9vLpJWV9YuwkcFHDC0lH2nSdT8ru+pCwMHs2buIfHJcZqA8g9OZIB
+RJOf4NqMONkYh40uSn4F2dnNFJ8kFa9pjvIYSurGDhXdjbjjqktno/Zqaa/bMuN+lh31B6XejGW
ZrQ6DWI4nFbDbjkTfZDsSOpaX/YE1f6W3MUh7XKJn8Jd9axtsCd0KUgnHqqiYWTbjG9/VJaEpVgi
AU+3zPoo7WdZgD3OBdJW7jo0tDiyu31c9xCMU3V0By39SVWBMpDAJ2Ap/lh/uzJ/PzeF4Qs863S3
xgMKSCUleNMeLbOGCPTeitYpbXM9NSXmhydM6MtJlybRM57Lg9loi0PYhPdhDGm8DQS2au95THIl
SWn3kdJyawKtyWcZTWY4a18nya8R0pHu60W5aUDAKC0xhlOBjErWVNK65/xN7+wREFBs1csaMIL6
9VcpOIPVYcmKDsS9l1D60OdMiq1fGBsRz+pGmHIh+xQ+D0Q1cU6kmvESUNgtr+d2bJ/t2+pASzIg
COreetAhj7iaY2G1OWnGxvAzjb7qjdjX9qiAdIFrRUsvtfiMpERdhZYRh+NYgv7Sm2s8huBSXSdZ
pmD/fOuJaqeXUsUmXi/O8ohtbpcdS60yylOx6rjMzdZ8LeYr8/uqEORWKEnHgUqSchqOHiONijOL
lggLiCcKzfP12IR0BsszJJgRRGb9XvgETiuVW6xlgd+SxZ4UYro5V5vgQ1UAzIIdzOkBXK1CGpAp
ajTivEc/yo3VaYmqG0JHjiH8gS+uFQ9a0PbkfnZDIcovEz+fhsWhLHR8BV4/HhQZfqxsjUMrjAUj
U41ArBAt3hGk8XeQTbLljxF7TIAQM4SAwc+LPIY1JwCaBMe/HnIUl75cBYLh4q7MkkXg0zPUxeMY
4aZQcY9kTSwLb5QXtvMhP1UQ/A8AbG0ZexDTYMPltRt6Oe0J3C1J0MSl7h/YbDLxBLjbNXRJW5hn
DEXG5gGbFs1SKppEzNOqybed4izq8n95Zgbj8OXAhZRSMTkaSeMD+nDRO7YWAlBS69yQx98XmIUY
/RWv/KJv8WtN5WyunFdGZV+CWgakmOHoCHV2z79W/7p27dBXs/TC7MeStgsJTpelh5KyCKD4yDDT
rqveJG2uIuufr5jHlNae1UEmyMVHWH9XVXOFjITLTOiyD7AOiOIAUOrldI46wWvU5ghG2QEXyno4
Rqrdp9KqkjwyUDHUPHH1igm/6dwkfWCGoec0+VUsUx3O4MOEWAS1J7+IkPp828E2h15u/Qlx1Yw2
ISty/X1pn4lqYYDvvZoiuzdYsC2nWTyD/eOr8kgrzh2iYGuuxC0MXZC6YOQmpht9muOJXxElDCp4
muAW6mjDR2aNzV6lEDv/OyzMuGN9Qsj0gFVaNnjOOuQ45MDKJeIl2uNLC+7OjSmpHzoBV6GL4x1H
fU1Ue9KlwYzCYnrwL1rmqNm6hZVpLgrQ9kduDqlammt0aSt9yjWOYN3yXszAQ7wpLLr00gnkwu12
BOAFBSZB/J9CqSfWEkE25E6OHuvOAndXuykxTEvlt4N44pnItEZTbpYA7lHxfqCynXm4pkV+wdD7
US0a1jchxsFwOg/3RI5/k2FZmWgjr+3OTrjy5dhZNig04s7PrcMtc+dHPirIa/VadeczQV1TIenb
zjgUckXk5ED5qby/ScKMM8W8ouKxuXBl5K4g8HHGia2g9W7dJJkhwqxk22Ls4fpPDY9gz5K7+26u
paMyQ3Xi0NLQ8KjpgmdIiJFUux1sn3oPteIbtkJTMyZDjco6dpJNwry+vWvp9c83H4gCSg+nRTje
pMfzpHX5tyx6yKHgDHcIOzPzQO7ehk/y3d4UF7XsbeQy6hmJFKtb+ZLVweSAcZE4EgY1aqO2cQUv
VP7wOg+y4HNOGgdp6AePR9aUTRyJYp94XW95mh1VuT31VUQ8YrzKi+9A4GbgL4dWqrE9nJRFk7tP
xzLS2RvqtkJlqYai4wGRPbc4qiiE8C7REv8M8BtIDcclW3wDGzI0V8TcvoxEEZ1Pr9l/F6PQ8KUt
jYIasxGedKpanJix1GnWmjM2CtmKyDEvKEJdykhIMmIb3KyuhT+fbxJGpXrxONXRlKXF+UuVMGyQ
jyYTGpj8u0DSCpmFw2hYP6ze33u6MTk18MHjQ4xzld5XHGMBeppVo+w6lxzYj+FVIZKDGVAKxZrt
2lCsK9OiX7LmzAFd6Yww05cFvzEboNlq+aYIZFpLyfpSq/caQBm50ubNpkbXAMqew8VBEkg1pJXC
Q8gARehG6sYHK3aDhFOxX96TYyqTWMHv+RhFvpBBaDuzvG5qlaTg/3LUVBHI4z0pb3jDi5g8M0QE
fQyNIaW+MiFNf3wiowPVmKIl3zpsxgprbfFfHqrUgERQ//gAlW94ys2xwsStwqGTHep4WAmgAnQi
3biQSIsEAkiwUpUGIeO9tuZSARs2wNVhiZKojx10KwMeGKCWAb3ygUvjhcWkpdQU1YdqNkqAJx8L
/GO7jcbascy7q2H3WTW+SBaQNnU0TJETnrLEoxcrgusI/AECvB2K1pWYb8BRdxSRbtXGM3mFhROw
zlWo2LQdumn/CLpp9F+GOyY7p+UJZ92QnG0O7/j+TSin+5XFA8HNRE97e2JZJw5ZzBsHEmAmWRH5
EdAwkoClufl6eBw/560+nLy810ubt9eXMeYJb35OJ+7X8xFAwl398dckWq79KON1GQp7+7P84ylu
7GRq/m8/tO4/jG8KR0b2B9SvSl8fqnS/wvdrf46TS2RRgQ2+FBtOOyP3ikYzrXFg542lRsE/R9VH
VEs8cSl2HgDY7FbURxlUmtQ0RGx/Qawa3PoazEAwT08H6efOz04RbBd5Wuno0Q2rsEp9aGEcrqnj
kM827m2cZdj3r8F49NsnJd1Fbd4tWrXC+IebUq7rtHJXsC5EP1Wy6CI4DR6u1NKnXbV543m27i6A
FtLbuKH0xvyq3HWB2pUwxOeOMgNu3f+/fdxVTBV7hVIAO+/Nw7qMenB/wdyEblRq6ZO9GPf7ZL2J
oo/Ue8+CFfQExzYW+zSnUb+qSkm+zrVLcceoXLQFMvVkVAhYromBH8Le/XTsIHSEgvNEPAtoSkjC
HngTWV7A46R1lGprqs6CGxh3cFGqCJE+k8IkXL9sQPyPn2DZV5ZEbqKPOsHSUYNTVy6ec9UeBst/
texCFyh3zXyAhNKxZY4F/baz75U9t8FJsmokltLbtKjrFo55ftZWcdbRKPTMv1dgMTQ9fizyph9J
3M6FTiI3Vib7j42zyXXLPgtmepizFR6y+55T08aU83WObtdl8WLctCN8Y15m7TLvxiaWZLofTnVo
nDfHUFBq7RUj+NVLzWvf/UCvgqeX+gGV9NQ7DTCOKk9huGmirRXZDmvCKDIc8EiSjILyLhyuUKAi
EFiSHWot+dlDIC/0ElQ9wsLejTmifQpf61zo6f2R11axlmcZs8Mf+CCMlj0TOTDa7Rix7yaxdY7N
5/w0Vuz2c2I2xjeWaYvQobzkQFUONuoyhItdK64IbI5WfVfYAw9MmPp9/mOya6hmE7GyTf5gQgKR
j8Xf2/Rw0OM2SK7BywjONnDeyf78Eu5pdpNzzDXp33BVDs9lpNfXE6R8BDCgzkTq+AJoZm5vI6wC
GYrgNM74Ad3/Tw2T5ioo/ynJfNYC7PbAGSPgNt9kUXj1XS/fL/KvAAocfCsYX+W6smSBm8E/XpKj
kFwp2VxADf6ilA4MjS5sqBpFKFik4bKOOKhe+4gnNlIPcndIIDmwiBk9n85ErEfGpvbseJETPSoa
Xgs5OEyzkL+wpuYbOO135PSWXovQhvvpo+Su89vP3E0hSB2Qtl+/gmhvKi375HPMaGcnC0eC60Hc
I8vc1n61MrlQVcjAeOXQXaJuGEIRKFbdWTU7vEVgIoYQ2iKpZsB+sB1KevK7KY/hcAk/J8VbmnT4
V1XIK8AWZEsK57BnxXT9dtJcFo02zE9ofi6MRE7paZfyyNra/6ktRXm9ifTKz+dsK3MCNwsuPGSA
gs01IYjK1NBWci2a12v6dmbkwdaskNBnFb0i2PBf/A+pNN8iRmpAYtZHC+M60RKwZ4dnTEimX4XV
0rfa70/2jNDgAZ3ckmF4blxF4sOfH+8idFMd6SqrsA+MxeafM3pOBzTHTxj5tqV90SAP7env/V36
3cMwzx5MASLWCJH+a7ru7e1SXACAXcxM0mNqchVjuRcKhUtlR+x4OHGV4dDUd1KRr6KoQc2yPFFs
ALveN7zkAhlTu9TQEWtCpLKAmU82iL1U1nroG191l5qQH2l7db7OScgwkiz1jwKtai26SFzlie8N
MVi8ZGzZqJWknTxFr2OoGlhuV3Rn46YntQ5xZ0S+cXajO75GAeVZC3/KRDpPsai3Gs8ZBeCAJ9YO
Me24yDh+fdaQjfI6BZtiY/znO5r6fdc7EcPwZYjfWLWIOkeYBEooQ9qjjURx6Y9XybyWe60nR4o6
X84jKs74Pq8JOYSd8N44wMOucaSbotE9z2TK70bUHsRfhMyic74Rkqw7WD4AFTHa2NeFUoHTwCxk
z+M1jwz4Zq5R119ZLO25yJ2UEnXDk19MZPw89X0X4tVh2PgfJqudUP/5kNlwrMkIIQfnxh29U+Hk
RLKwWhcKPRtIcR1CokHoXfPufXlM0qB4cGFeO4uD1yS+BWWalRnjQ4lanL0lC7Yz68y0JkZjuxiY
Mi0auzX7liq5wL7CeJ9n6NAsQyqc6pnVpZ7GSEXtu7C+UQPDdJkv4IeAxqknSylgCChZkrVoIWcv
/xVTbDwNh/EpiLwROBeQEPNqBBe6jf9yUXy7YYEfR7SFeSDhit+x3gaiLxabH9kkhaNYR8arXWQ0
SZjwANc/Akt0ZlGUgVUZRVa1mWiDUUvc396UnMp/O+BsOz4lKCy9PSMDgZg3EzVjykjiRV52UwRG
KDEFwQelulaUp2iqMz88Nq0R7K9FtKvfDyt9vFK3LPEI3nKn171ReLU7UXWxvQNZ/LIlaC5kXUqp
/wbMNLcAx3jXriyYB4kxyc4M9D0Os0wFGg2j4fq48KDxwwb18q494SKfYyuDY/51/G9KukNiPa0Z
ze9Z2Mj694BAWzCJXCGppv1oK6hG0WynuQG8Fsbe4NXx+9+f2nkgr0DuDx7duYPsQ2fdByr8mEwS
UPetivUKYcjwaqB6RSrfO54QDsLyvzHxrs5FMnSNJEhM1bKJLnQ9l/thz3OjIytDEa5VLFvcWaCo
r1KwJk9Bop2ONrMx7XGL4E0Ont/UZe01JvFiwv6lPaC9qfMj4/xuHZHNTooXfbQsLMaYUL2GNkBH
FPKUe3WGwv4mlgFXURMZI0sMidpGhiLl1c80YKbjowyvl6fiVzKr4OgkajVUZwx8kN9bWfXiT3py
LuTepPvXTdxLgK996cM64X7JMrysVogYQ+Y9jhERTpSsYACxD6KMocnGbuJNCjr7/Xs6tYe04dTZ
r31HxeQ8kfGHLJbg1o0ONMeFeXb8cEDlFkzXW/FX/TtAJwGKQDiclkL6ZW6aSgJ0dFy/NqAKmK6x
tPWjHiVC/reH4tuYQX1/YfS+5DamWuGeRtOBVSmRUQN53n7LmdaewncUv/4Bz47tYneya9PInOxS
UWJZiG70Roequl+wAJR6Mbth/UJeexcyWQYL2z41qOG1r0W92eksKhD+m28m4X2bVib4/dLQOpXF
Xh47EYQfzoAyZA/DNjLaPm7Kg1JRsEEwfRBHkNUIH42amjJpeWlY609eM4TEx7J0v+j5zkxpMNRO
s6vK39ZlgpuENYAWeeM8+NbEvNbuPwNTFRAU6q9etwmB7mK9BqQA4QtwYuAmMtYT/iL1XdfsX812
Wgt2z8ofujJ8Ef8mLN3AiJP30AOD12sYdouQKJYZ1JwxPWJRHA46hdDUubVQUlhqTA/ng1ahuAe9
zCxZdOBee8zyxXvGZO/Hv5yDd5gWVOc+CnX8ruqdV5OEZ4NocygoGYQhx6jW9SpgibpMO48+GoCu
FyOeO2nPbp5omCs7siS+sUeDwTM/zyeD9w97LUS719xPZE9b/SmxvoLAW+gzH1ZiRux7syMT7zAH
TjS9PrcjJf+4LbupSXw/1w3i5eRTIprzR9YTy+vo5PBjtTWI4MPlz3LKKoePycI36SVNKMmmKCcE
aiJBXph3xjqTZdjKPXKh+puI9loC/JDu1GqoX3uVCahn7yfvrNfzWBZKCYykKxLfO60vrelO9Lfj
jb8njrWQQag9y60dFrF2C5lN+hr0AuCGMGcZsaKu5PP7FpO88Si/cp9fQPqwdOJSU+WAlKDn3QEH
E2hHTu5X7t5bTDHLE6VNRKObb7AJs2cdhDTBpOO59xj5htsVw+9O1j+gIYoHQ1Wm+5FZHR530xyT
Gm82E6G54IZwC3yDYhz0RbPa8SmF/ag36zjSVllfq23mguX/kvzWgOAhK2Wscfhk78AtjWBzdQoT
nBc2ItZGUS9c9PJsaLmYj7YNqoojvxT0+/I/6xz89gOYspUPM1u6oMyiUEGQyKmjfLpRVogUH/Xb
rMl9b8eMAYOIozQs0gqtXCOAbJPNtNnmBRelPcDsCRbocdeHjn5lwwzUN3nT1soDBQmZBAkgbSYE
LuA8nrPQB0anyV9Ip6qP4H/IVsZjEUd7e0us1dgWV9GxXsc4CkORZ9F31FyGi13y2RHCLDqzE0D+
tIb8d3x5/vYtqidToLhsWwRGpRTQq4Jc1eFgJGuHFBua8QYGx5DtaKZ6AHVlyuv2CNrJyPEZpmMs
HvWrid3Zebnod2KmooK5+pq28lgZru7dNMHo/aqSrsbkf5R+NX/1dMPncf4k3kb4PLR0ZaW/exhL
F8OTMFjSxcC62UeY21AxYx3fU7LLTpu8Fuc0LI/kF8XQVVRBRg5ugQfKDR6GUVKpdVG7RcLgwC0p
fqOKfpYbnb6oMuqtrOCoEcN20LUB8e2C3zzfI0M8jr77tEdByfMleqYiUfpcBLUAEEZQy5QZFeVr
PM3MyXcNPKJw7JRwaF3xNwVfJ4fSoAnXFPurKKctpu+HCOkqtEhYpsKDQpWX6rEbdnOGbTRJzqhE
iE7qV3YdPU3nqDSoVLVtlUm/lhtRtk6wfHZXSP3RIJNk5ZKJeqdur7pLhXMLLAB5RVkLKMm12Azd
zD/1m1j2nXkwH30zXDhZzUmduTI05KpzVjY5F9xKH0m1kwPI9heWsI3Qk63uTEI8Aybx2wt2k8za
YVepNFjoEAMfI7Cfz1lH6RYyywcp4ihsAQa3bsDuEJMxepEu8hNOLu2DRjDMj2lXLTUMEAdr2l15
mXVr3qiLPVumHKYDXst6ljLgOTxhlleJSIse8BkEJ0m+d4R3qmcuawn6vRboA79fIUS9S0AjhBwE
FG71F/SKk0ck1MFPnTw0QfCkIiZL/pkPluWdiieGkxpVq6eZFtcCVKo8E+/M6QVX57Lon1FIB+YQ
JJMGPCKnhyvkDTm5tdqdm6C/5RRyL74EdV24mDiNzXyfQXOFzCfDSUBpa2m1nQWwzvGeEA7SxOmD
AytTrV0AV/BOUIP39FHL9H0nXQfiPCb8fXg68Zcuny+o1zgW8f/Hh6vA2OxyRDRc1TrKGWPg2LWh
oDe+neaWWAZyApMWEkZjvNY5MYyDNL5W/n02VxOUkzqQkYDzdSAQrflcQ+WCSqIf/O8KY9x7TcO+
3zSR3DxWoTAQWg2/ASpX38erMVAkBOXrjX/BwlMkWRKzd/aBQzOaoZHXta6RxKpvDsZvCR//Bsy3
JmU53KA1rl3jRVFVAZRY86FOlBYkFAB5E6ZrVj2FV7+MC3aca+EODNwpQABrB97JIyokmA17u8k9
YSVd+SJy+8wWNh6akphTojLq+cGqV8SUyXEs7M0c6Iy8LK+hu8kb1o3eeMOkidxM5qnBhNwqwFXj
v+Jmk2jhR6Wrn1Vj8S0vKlCoeToqESUvEXRWW0TDEqX9HCUGxE97byvs5clJI1E6ZQx2LhlU4ZO+
9cmtsRIFP3nNPbCYqyke6VKH18MO3/vhdVjUtKvhW+voe1nlHYSpPW26vPwyDQthkSU/72YcIciw
JqnNbQBx/m9Nle8muwuBBWys3qajs8J/U/zB6NMT5/5Tjkw2cLZ5a4HQmyewpDVkFU7peiDr+U/y
6hHAZeJVYU1yhOe2gJ5UQhfbF9hlt4zJnT9zTQjZgpaLacluDZv6B0g8EAtWBlFroVqlWIXDtxcb
w3mDOCcCooKOwr5hXaem28eanxSc5e8n216BcOQC3pWf6nlAKKh1ElatCva16nX1yrL5xOjvFSWq
1cCx+oBxXjjCUeRPmt5KwpgkNbnP+uQH91zmxzAoYt+Wq3yZrWXlaOgzaFclm4tf7VIV67Qr1MmD
YRNQ+y/dJaoRkMD5vQUPWNXhZk1XQhSu1wecuO1lUavMNyR8K1yBp6r7r2dTcw9mfKqz7xeFJwyh
Eg+ckaAsJHKHoi4wrqaDQAvAZIOjFRqnB0Qd/Rt1eJnY9eh9pIn25i/q0EfM97DxJd6KndxdNyFM
bqrgieLZch1k+ZQ1VtOnh0Uo0OKlG8M0TBSbwtQJb7Ji7Kvy9etUCwKBrIYpkRkIaJE/zR2kx2Fa
zxgUtYmCdcibe3gNJ+82TIGxEAO/OBNGYsgpRvGfEZYmhhTZdLzhbw0xXHxZaZ13LwVC/qxEKtTs
ukcE7+r/heCmZ3q/KVcpsXUFBfuf77HaNsdRSGPG2BaOoVpJcqvZdWT0P17jKKJ5uPAFllZWQtkw
b2VYQ5j3NCzhZUsJWGx1FWmd7FjmqzMSy1GRqJYIZQFImEwXKK0sSAXU+7hQUfRp0GHcryeBosGA
eSYOpzGU07s8DIf3HO/AKEsFYT8AzAGHzLDf1BcM9XfdE7E0Q+Uff9DpCfFHVLBmIM02qyJzF7Lt
7/fWJAQe758ywbaEE4FrX2bFlR0ez4Xjf1eGBluj9KZid0JDvvqQZz5jGIDNna2aLiha6V9CbSCi
6KmUv9saJEMl6OWugao0kjhluKThZ06BLh3PWzlE0jicL4qDB2LgYcyyljPb87noHC3uQaAA8HxQ
FvlIDIR8KBwVeT7RuVdno9IWvsjO8xOichzD0KZN4u75Xs0n15saRHA+B27lG+NZZK2Y1pRnwa6f
BrrDY/QW+M6XUzZ12kdFzLZpWnLxXjv45uWP4wX1ZarPaOylrYwCR5Kvm+e+RkX3qkY192TP/EEn
DFfjz2ll2B3J+qpQ+oVcemQPDbXAHbMtzROes7wyzOc388jMW7b//qFZDOKFQxnJxysKzZXLgow+
x9iK81I5Iw7RP8+ZV819XjrzukO4Lqf7SU37QbMA3YpPEc3Mt4UtTUPxAl7GaNzJC8fteUdziA+t
4384fjPdMfPohRdQP60NZDG7oA+VtxldxwahJ+BC8Wy9LJ/o6xnD6V9VaQFVJFnJefP1wjFOyS6n
HNYlUF1XoWELz81c5gsuKfIUU9eVLoSm7m+B9auqPEIa5nHEqH7IJVEffCbOnfrOE/kCuol8nUM3
66piEBwv8MiVfyXk8Ik31GeOfWH5/2z+nQKnHtta74eLzVuJjTB/xziU8sOFVe8wSxzQEmtMLcTM
WCOlrnzvb7QC1qKs+yBLqt6Oa5xTj0kDD/PTpIsgoZHkfHLgmo15wP5VNVgo6y9LeT3PwfANKk2y
w1bchZ3HOsTa26Y+7FWBO5pQq586s6J+Qj2epr9Szg8uGSVF6Z6i07xz0AxbisaNSYMI6TxGnqqk
hf0H6ZVOuG1Tg1Xa7v1IL7QybhO1VhmUKPUeyMrPN2ve/BDzGuYJlEYZQ9y2JwrNqbZ4e848K1b0
2vCS3NLqQekclkoAVTH4EEEJCbL5jPpdxcfR6Kr7gIJ0A1yrmYOA8RlfKMe+bRvemEmLfkyBur5K
Kr2iJy1TTeBtDG1QalBiggJeKn5UdC4Lzd+9EWAzOm1IgtSWVtw37AitWA14fvgflqKCFb1lgD7e
vzK14wcZygjuSR/QjJNtHZqkwlZxcOzYMe8Fhm8wcxYIWBDkkr8OESU+8sHZPPqYaqzb0GfnbefM
oXiCjbefUebSQ4kt0Onq/91kPbhsFee1J0EFjUiV4nkCkDHGJbCJN3k/PZ4HCJHqRYJr0OYgyo3J
g3r/RG1ndYCqMA+81byyzS76EhNb+nNo6PcvkH+85E3UWxIPr5E9f/nnsL/nvG5W18cr899ZmZef
zgK7nsJfetfB22WjFE8TWjkvE4qA9gwOo/LWaY/uVRHkNLxYhSToL56QKwyz31MggQp+IXOu4jQS
o5xzqyB6rCScbqIeA1ZGiuvinHXExMCOJK6zj7y+Sx6o01QiEp9V4syE2N6RuOY7t3bwVcb5xsTw
RLz+8B+XFz+4CHceqgHgMXQaF7+zgVV/w1TvNM1p5+mKeh4BgXoO6ub4Y4rB36y28M8EOdXcCXV6
yLrsQhrqpMPu2Mot59EMKtjA66TjeEqSXS9aO9KvsmNUUajoLHInp/vw/bBJTqnOkHPCVFf5k/LW
yvivm5X4Xly5ZxIkSW7LCN3ImWHcPJbWRGwBBiLiRck7k+49LPZTExjdrzw1Cg+6p8qO2W0zjW5n
FU/S1Fgl0CQWxqLImwwvN4W1wYPV2QuAWt3btfouT8WFEzMaB87NJJJimI4aENC6crmTNAA1ZfZj
Q19DWpdZontGEnwNNQ0J/OdJlNTULD6STx29ELjNL7NU8zz0KqTGdgKqpbNnWe+g/IXbjGtnhMek
J/VD4qqfTd9/m85GWueW9CJzSX6kP1b0EDZ6knfmm8jPrUBnVkmQKfYKAvwGeeCjvYbI8Vnlb+om
SSjonotMudjCFiUl+RPBOmkmhsFFr1nqXDflse2jPZ6UKV8sr9klcFqPHoPqiPjvCd6sXnQK6aFA
W6P1QMJzuUtTWIkX4V6ivyMNg2R6QPGejlFKW9MDlQ/oJtDtMvlorYaONYf8zhJwnUYX8KJZCjy7
uZuapKnH0jSFGhWe12RmgPmZT25p44oSVRGeY2TvZKAG8FiktnRLaGyYeBCwPHNqFCT8x9+Jx1pk
hrTWRmOz1iOUg5t58e51/UP8Wfwtsr9f+jLZqux5wfzJwUK7DE32ytHz/it4oUAe4S88frAZKtt8
sB/ay1aKlsMkVUpow9So5L4rG5Ei+wud1YNEudU4qy32F2VnJwUm/uxpqet+5IJtdhjN8iskB+r7
exqzlznhf+gXebGW/QJDtRLMCXIHPdMvOzhfIn2TJB5p14gTFnTyV51LfrCmMhwNZ3AfEFHJ8N0e
+Z+t/wH0bJDsAORxmnXFvlRgb9lfXgwiCGgw78wcRI8w9XXd+jREuAqCY8PHvuP91d0mXVnZHGVO
96rlQPFzTmLi9gO8tJGgrc/qSj44PDtUbB1NyO1B9X9k0gmo4p5DG12RpienJOsnvmjglPA4tEow
+JJbr2ZG3y0zMpyzul83A83WT9So4O4cKNI0fkaX6SyPSXq+aTHxdXZfHoJVcty1/A1FHFDfsx1r
q2kgMpt3m5/nJRlNsn5a3ALxp5qLfjObQhf3bVUwHnEn7dNw5uFLXcZ/T1LjJDaOj6GKNgvuFicr
D5b6UgGl0O3+CMSoZYYTogE9LyRW9LfCdaUUt3ub+ry5IDTP5fdFArL6O+uvZThtKjQp2g5fIEDA
wnEWmI0M1ggr05DLsTNzQlvPVSLl0HdYeN20c5aVyos9htv3HZvtsOKRuyJzCIKu6a9II0wQ3RR2
mzINXRiAUBmc6J9mAhvoNf7CbEb15ThrpTjpEhlBm97g1aHVx/+1F/tnz8QkPdMXrf39X333Dl46
LYrTJBnv/kUOpF5eiKulVRewBcGakU+YWcVyc3T4Mx3RiWh4ntOh/MVlHBgC9TraHiFBDK76D+Bf
MaDFtTUJn13XpISDUZhIYAoddGFlpqhAnNQ4uPoA7IlHkPFqf+cmKgf7vKJaUc5a/sYx/oJ7sHeZ
75Wu+QMwnYFcnXnNaYXMuSM6xAuG4dFBFtjmO44prN6Vm62+7sgerXI/SczsG+mxdl1KNxiE4S7e
4Oj2cNTA/LpMCDQ1OuzhKrtB9ZmuAQkntQpFyVB8DXdfNaCosW6RGoistOYDAzlU90a4Pa8RpGlN
D5xJ2a6IEM/Tys08iCMbHnoRpOpuujcvyG6LzUpYoU35lIRgngEZQAwU7sdiuS67CE6Dxdzy30eA
fqPFvPyOMQyAqrpTsv6ZMJ5GSbj00o81MwLikxKW1sTqE43SBZ34t7bm+o6Cb4rzuNYWbNiF9VIm
dr1mzohWXxk+uGbXbcEdea5NhEg0+hqYV3utZyIdrv2KWxKoKLY/JEY2x4q8NT5moaLQ92GWrB2h
RojU53ZnEFipUVSdlOn1izsjXA8sylq8JZ3VqK/4AwcBAPSlyKQ6rb6tukqXS7HzXFbfkog6dv+j
3XI3BVYI71wArREaYmkFKC9YD6+rWE9A5B4jdCMwhiOQ8906NmL9JqcVX8MFlMhk+g54qAb+TKlX
n/rD7C/aErthlkhu0LXKWblc5QCVGPh3r+qE2j+h+eLV2I9/qb7cROrdlXKc9ryJH9MN/goGw9AJ
ldZLJ841fPBzhkFpNBS5pUCOM873dbFXCVl4FtOFOcKtoSl0siBOI9/0VHlCRS1AapwdCcI8YX73
7ErOhGLbGYyREJ7vwvRAq4cdxS8lRPfxG79TlC1LKWnuD1Wl18zKOztqhsJNB0hpoS6+wMrVYljp
J8iitXoYG3FUNBg3Z/LgyWS5gWgjoV+L8KWa9BSXroPPOd/JVZaU+S0dADZVv+WXkQW2E5IfFzmX
PG/njeN3fKyB4IGioMf++E7FgdskGxSmctiKY6KDkmgYnMsHTxyaLlWXc2T3xYy7mx3VNd1AcnpE
nf9BSBukCsS4iYDEX3FlaoMYlnDBDjosf8KJKtBtrXhHwhf21cXZ/zjeNyJMiHGlRUYMLqMvXgQT
OqyfoqF9ObxcIWZO2l1IMzVBKMa1HKkugD+J7HS7+aa9c/feYxWbpb/Hqy8QVbX4SM5kc7qN7fMF
arykrJar8Qs4hH1M2LK7looJzFMPBFTI5dsnzfYZoNcvVLtZ6y4fJ/uk0LtwgRyEKR+HZ9HGmkS7
2qF4RFGsy+r27Dn9O9T70bDdPJzWXd6x8tsf+ts+IX7wFWa1IajaXBJxCcY3WAVGLA8jc4I8YhdT
Q5X5Evlb135rXz9ERBlgIroxfhpxCMuM1jj3KD1BLNNNn5yd4RBqE+c8NAUvz1m5AWxirVvoKKUy
YvdUCZc/Y9QUxoLhvO5WCovVDlATuBlJUlUoVGU/sArys80aSiHLCamWN85b+ABTSCbrr285TYch
zlvltvGWmse9m+baC4SfoUP+Be4s/bKyHQ6WRjV4B4yf7PRMvQ9eB05SdDwo4rKpimct/0KG+NfO
dol4levKliRKlXPoP8FQyHKKAM+tRSvfxCxgM5V2t55f8IJPFsAGsjuq+MSYNq+9bCGLyxWeCU6I
z2Ji12eX/qzEAjJQNND2kvZAakMYKKwF9K9ER63OPwf5Lfwh7dXZfYVe+NFdLCx8LZyBv31/TI9B
PetbF1wKCPmT5s5Pyrkjin6fNLMoKt52Mtip6T4831rCEirA6YLMkpyCpgwZDko9Hfw9redAjgAE
QmMsOchaMgo3fDEAf4NlcFHE3TvEuCChQjXbwJs2BgoFDf5nCOPkwwe8snXFpwYATciSE2xmgIYT
uNdEUgMxb4QNOdtvKZeZf2Wb7m7zdav7/ZvtZLJoZdfIpFc3K1X2JaPyHCH7PH3etJQA4NlGn/ph
J0MdaqEKKdieKBj3Hz8TQWCcqR64hYkPauVAPt6hVrVQxBKBpFd8j6wps0pvvdZPIhnv3KbFcr2d
hp38Eb1t4TV/20UtGwrE827nigz42NdTdQHrJ9nxF/Kr8u24/kUdkTYgFY9Kb4IXDqguuNqOHzbv
+lrZbrPK2HJt8QPv5UTti6BjN8ZuV9Kc0deUO7JxA+hzLibvP9/2AC2hy/qJ4inzS8lYFJU79Z5X
BvqN0o2ZrqqJOe5YKMbWGRiEBlGPCjD6SrhadoFR2d52/RSwFQd6yT+T5+kpuXphP2qGIMSp0Nz1
i0r+4cblxRgSqN6k3Ihe8oZDGje5jfh47O1t2S1JkEdNQbcYOUsJZQoPFHh4VCbksXDI2IL/oCtt
3+bXrN91tz/TeP1PPnNOCJvhuDFNvzPkNpavI3hHa6M1NEcr1dLGCAzG/sdN9brm4oJexaUyAbCK
5yZNkS9LcqVyuubf49CgiFUCMHpyaH+B1dnTVXCtTnjUAZxj4fK95ksra2JqV8pDEJhuaQr3iNxK
Wc9VpuRhw0X4Acxqk0eqpPjKSs9q+rynlq+GOYrBT6Sp9D1iqzLk4cZzLeIGsN6gI9jam+bgjEZ7
H43vSsb6rRT0Ha+EjC5w1BXa+9DAJn5QfnrQhqVqqPjGEfzIRZKA4hXb42Aq/64A7ecjk2TV3Spr
eWdPDySNo6ypk1LNBTNOY3HHbw3/bsNgsq0BfeeYwtb6C8iZjhay3uHj+DHLrFZbro9awE4nDCLA
Ldkzk2Hyl2AviLqzvqFUDO+53Ao3xak2Y13q2DVbr9WlWmm3BG5O4eoSLN33+OlUdAANftDm6k0S
2KDySN4YP7IHgfkle1Zcyl0C4ZYwBfCY59gWCjJgWvDZd097Ptc57kcrLrSmn8g6dbjd2tMIkuFp
55yws2N0562X9h51F1/deUcvKdfGUvJeCzyowjs0ilKtu6Tp3EtpZPjeFJqPA7oiHe52mox8cNUx
4E7PGvXoprCBhKk2Xx6ZnZMI41DR9AvxWpV1LrkO2eSpK1cOHdrwVpPcPMZb+VVDeKAnOCVCmdgi
wNmt7DfleW4qXLg1gtFWnafPISxrImcsHj4rwe2S/ZkyAc49tjkFecO70VjF/UbdKOL6dMer+Weq
V5KSQz4BdA1UD4B/SIMwZdpC6+Kf2MH8d+Xkqsl/7UfIQTUabx02Ofb0LBG5qhj5W3j2az7QeXfk
osmqHWq5+D2AOuur5MeWoP+MU8mVMSth5r4SKEMTvnI6xIkf6UP3TvMXZIqvpf1cjElEeGQyYTv3
Puajqpk5RVf1RwsTfi0O+m1lzyToG4Nt4HZob/CeqlmHwOqssc8NX03GK5ltmscGP2y+QCwzjTCz
wXanfjlmRQwvnJ1628fmpFoUnJfa8HoNvcpzuDYUq5bPpiFK7q1Auww+O9HyPHYaKBajsYwWpEFs
R5SflBWnpiiFAiaf5gOd+1ohdka7JVNih4VnKIcsODA27JCoKUDUyY5eLxItETNARF2TvoK+G1lm
LukmPE3gYTIFjvUH8AcUPT7ziieraajRFj4FFMR2jdCvmyZHAfSUd7mVvMd7OWtinAIEiN4i8jYw
hzww4dQ+M0eEn02XxFRkHRKJ4ddaKLS1dmRcTLR6YHaB5BB2C6Jejqnu0AR6Rw0fhQUd5QiGIDtD
WVANGSzdyTWiYnfPHgWEa1Io6kOmdzthp/OgHcZTKdLgqjG6GVgbhVF3Z1RF+VYxyA9uvoTnRTma
KWr9Man5oaccgYU5vxW4MsHJ5Bxeina60xCN1gECnxMG+TCxUI/Q4byKBpv7S7GP4EFXDptjq75V
K/h5Hn4/rGdeCnGFqZHYrEmJAgFE884kp3q/mNgYrh3nfgIMo1QfuM24P476cBNSh0hHGkL6ZCfu
2H36A98QFDHP2NXQpDNlYZmZ2hejrB/EVLvfa9QgYo/V0E4NHXvgO4itniFJeCsbgcpxLgeyaGj0
qf3ZpApgqSaiJUqv3WKpqQjnZ3QB7+Y+YBY+CZ7tNLyBVSVc35DB98fzW0hmKyV8peTnM2V/spas
PiKSTNR5sWr4NcnEKZ3ZZuiwvGUcF+0wxkf0wY5H+3Mu6z+BatZoYd9YFeJ/CXSon8T7jILhggcH
zBAMQOYOu2F3MtGEgFCp9Mmw796u2n8jxVsUI5FZ3AXNsV7IRgywPvWh5trL4uw8UnbFaM9DkANO
YrkYW0DKrrBpKMAwsYk2UE1ljxtzYU7ll1T4ubTSrKX3gpmbC71wpDbwOfGGulQrLb7V9RUXPQs6
H8VX7t2FT2Oz+GXCliNSwsWSYd3+lDNW2iJQTc/nzEFv8RV4MPFhVV1r9PiQl3YePtH7JDsQv8a0
Kc1UbBTHyAdxymCMqQWgb1uYupwy24213BCQvvOnS8iutDFVG/kEjnz41dAgemgDjLOLnLWZDU0I
Qjcyg7oh9YSlTOyJ8QOKh4/IdJcR3UudgIUaJBUvKsCFMcV8+R2weSzO6yDMR+Uw4z66IcYEB56F
PIOsPRHPW5D5muCxrK2F/fvB+mYRvIi7qXyIf9154XJcg7kF5Pkt1v/JaGeWE3QrDdQJqKVRYUDe
kVS7oJjwfjp0e4DVns9bKoTWq3Ztmgfa34cVVsGGquQe0WyEx+3xyfGoNdh9Vx8ZcPOm7wCnBOXL
zg2qMq61bkcv3cuoCXfTYP2LDdoK/SBJVH8yBQ5EHxHZ0jP2mQA7llo4GBehcpdX/EbBuhEXk0uA
NPrb0QUC7XXuDJ2vutn1OhLVogytZX/CRjq7X8qqNBxiD+M0mAOHb+YZToek+WqRgStYUtTp9kVE
YjTMTebxFglz3aPP0qaFgjfHii0+zj+LqC35VmbW3R6RrPIM2DHHVKKkhJNUQiXeWAOtkHEQaTCd
j7K78vex/jnefhnRJXl82plYh2tJTU2t9EZvXhSbAXHmBPLI+MLaqkdxFCenp6PxiJrxiMd3ETD3
pCNodRW2JImYb97fKeAYKyIeO5U2pRsJNVg8pozBaUZzuNSGbAnKya40S4a+KGWFBnN35zzbPpq5
rPogwauEeSkUBP6DU5CtABswikBC/SsAg1ztBVN81h1kuBj8g8BShrMkqxI8Bkw3rVTI+QDpSjcK
DbjxgNR3DQ0/pQv9Q22bBhGWJlOu2GigEH/hNS1XyRfK7jriyhQXNSmDEkJqJqsJznYyEZ5ED3a/
C6tXwZXOGBo8+mSrbP9RhrbDwLubCrl3AF/lz5sAhv6hi2EWs8fvCv7c3zA+sWX8V2tOx39mio9D
qViTKZ8mlcWRk5nGSi8uGozOtyecUl4CR+cPUs1dY2buydyOmalz52jA/AMIL3u54dZQGXYIWEQe
GRDsxld+CwcXsEBh/4AJM7tdE6I4sMwSWFhdGYfEAR9FIeznCt1ZA97ayMvRLGlFaFt/sZZmFQxn
MVAvRPhEEACF8rtM486mmyZtuHlZm6nF5CUmguquvhKb3JODMuIFapansacv5WcOD3lw4W+HesLO
gTIjELfd/+N6g0Z3YRw/RST4x9yWalrDs9E2TTVn8Ooc3pCIA2Pk2hH/ayPZ4cGDZWszclEKBv/l
WhXN7K332CvP4RPo5TVkEg03M5rnfPV1SUgwNLplxniaKbQ+VVqawdt4VSujokYfp0z92g7rBVDY
nsfexdM2AK8Rm9lfxsDgw11rQR9R8WygS0johY1ddWK68s19hkLKRpbXhujVT+xo9XiGZPHXV5ch
N7uHykwxQzOiYBHKzZlayTf+dA4aJ4VvA7k4iivh+iKiWlIKscWPCblF+yvDn5HxkCbXgaozjotL
k2Y/hxQCI7u51plnwFfQWzs/7EO0VGMu1JYFvWm79YqNyzchI+0fgUxdFo5C7nu3EDweECT/QLWy
8cIWOyquo8bvDku7/e6WWA+61zMWaZik1k6NHSvVx2/uq3iXFCWx40HnmyDTOJI+bNHt4sOsyCia
DtircECcLt9EWCH2ngV/oTIwOSTjKmr4guri5f/QhYRhwMdKlAsOVKLf0TFiFje7/2+pHQJ0V1Sb
QJHVQ1c2VyY42123pmtnAt19wiJprTjFRYQ2B4PoavXnOA5P7QTUyyDF8Zm7v2J/dnsyjjSaO92m
yQ1bRrTg8CFTtpvtPuNKrjazfyYhQoh2ry9pPq+nlftV5VNj04uxYJtLLehL0Vh138xrgy+iH/rL
rmuMCk7+e4doB2wQjgFTIwRI7tyLlWblFpNZMh+4qqRWrEIVTLSFN/jjzf++Oj0Mw//ujjd1tMkM
MMdipsJrTrekZ5PLZ07jYanpeiNxkwf+vJ9NRqPwNqmp8/Itc1gu0cSXyUgwFhBN0+tPDvO6pCo+
6SmZqNYzJl6+gepB7nhCzfj68CT9YCFnj0kC+oPu/82jBrZRNfHdgWwPsqGMWx4YfJ239Zz3Ix5m
2ROJSgSwo/EJkfXGiAhdHJL9p53LuTOUk26TT2adFYTwkPdZ9OxPuvJg6vQlO83AlC14VJxVxjBb
QEers+n/RwHN/c3semIHtjGrQGK886bfhNMr/gmBn7sS9f7ferNfG/Y/tj9nPgBZav/wVxci2QtP
+2IWIGKD70D9l22uf10eq7HaaM1C/JmwTEXCb7As/NEZVmtX7P3wzmm4x04dEB8MsxmJa6H4ZDSK
lhdrP+jyeQHYtRyRbWoVCO1WT4Q5LWhBmochcXyTkd9SChKlUmuaR/R1Hzfrd9zrf3KzWA68qMAF
QIw24YTUxiY+W7r4MYlbKKLsgPF7rIMP7/dOTrYZ40Oh+V0vo7t9naXQ4D0Himf1Kk2eyWvQw+jF
zZOnkLnC+2qzWWJWLrlfgx73+/Vb/HDSO3BTei0IkJ7i3odjKqq9GhqK9oCdmXjUZjNkMtkDJDFP
X34aeSHhuPOSomY0TgzgzpTFUva6MzscfeI1nDk3y97gUsT0LGM+qXhW++9H0+0SAVpEa5fs6jSt
jp+9qvu1FKQ5n2pAOrvDUdak+m5pfKyhtPFIbvp8miNgs5aFK5vx0Zaaw9ADR0uGBRmb/AlHo+hK
UW7OyXvscPWuzbO4jX21QHCshnMzwkiZaUOzeXMdFsTl7EsgXoTXwmX9eUL0Pj/keczQdin5gmw3
SMOEqOKLt9+q1CwhhJOnZN3b2RgXUTsfwHIsQcMX9GaHoGPyMMkmnfuPX8x0GR1E1QCwj3re1jwq
b/58sX1KuJSkubQAaWhpTkO7Zyf4rlggrO7ytF1oBDdDwPXebNAbUxwBLAsAsu5iGRmkeFA1Gk+x
Y5uQZyVeP/D7Y/4wrO/0KKlu+yKvqetFTCNVTdontf0C8fdojKCXBseoqybJa0dAlWdISJtSl5io
edIKOb3xUY26abI9MFOzVn98zOnVohqvtsLs5/D4dVKJa57duigT7Q+DkDo7n6142y+m+EUsE1Qk
z4HUJBCwRpVhHTz55I5yT1M5S/3ETHCTLNjFw7Ci1bspaLO7fDHE1uz3F/e4ioiBpeFqAgecJ1gY
iUSLnJL21soAfLz4Mo74zboEweJr68DFUzt+I1N3BV7OH8zaiILd7qWGs+zr6zkQkjDZ3N/HaN7Z
2JyvIcdpYHA8TGCPFOmrZL9SEOAhagiUkJpLYWlvnoyORYIx6vzW6nrzckmAh3L14pB8NRObOZhI
CoiFLesWCCLxocH0j5zd2wUPPlKyOliKfBnebkIfvhL96t/6KbM3hJB4hhPC7stDtOamHwKYsf9O
5Zv26AjynlBpL5IYjN5ZOo6NjWx6KxeRxpsBDsuWrdxwmAF5TJmgsYHW+rl+hCtGMY0s0yGOtHvg
7xnwiKXY3USrCNawazbTAB4ONK5KxF6xy6M9Ch34elov4JHxO8/F1as5cR1NYEdqgMk0t/yGxqnx
vTmjBS6sARNHSuUb3y3KeB74ehSrt9MQoMIzmPj3Gh7rMXvE9NbraZMQNmkyMwrYigJY/sr6dv7I
05WG+no1lnlrXsbQPbLVpwxVlLRlB0OPc0QJOoe1EKFQ7em+SAPgYStJVJ4KcsXoOvh51TlLOiJ9
YLMlBYB8Iodky5YjlGmquN9xIyD5F1nV76Zu2SCglP44NwB3/x3OzrrCkHzDVmL8hv/XxtFk8u0s
XS6ZIyVz9HSptkQeDfkWG2u7vB5jBjV8c0IjGDcgdU1UBGyjAhjJaQh8GVkZQiXU+0dV0fah+xNF
Ll0VBZb6rLdtpV1Zm9H52OpArSIiRio1AsCDaq0q6u1vaHip/KRY659muq8dGCnZyCXmzImC17u7
RzuulatQPkNwXIVLvX64DaJBLHYAiKor5NYoYFrJy2jl+rRxltEZn4ATQrCkDPGHMk7LDUX4xAw6
60J/7dUbSPezDgK7J+NERPG8K73DIyS82bAE8nfe/Ntby+mPi/MvGdALDG0tRSOVmbfA4KBQgfkJ
fOhr5Tprei/6ikBKPxmKercVJBXZSEInNAWvEyORY3YyrxdB/zT046jK6PBBa6xyyL0R7lUerSHX
JWTvxCAgeSS3lnWBPCNTUWlI7c7Cugvo016UMES3wZIMsGq7MxwSJ223YV2N/buYjTSC0IvSjLnu
UVvkwZ11VSTXTCGldlA/5utR56aLmY+cR3L0gLFcRCUMONJ22plhl+S09tkLKnQx1NyPiWTB4VvC
fJ110aJKmDH6Ujk9tll26HPArglN22i0yo/JAtBw0Dg4RYSTz54COX9SK+qTF5JWUhaAhHz1Mj/D
F69jA+db0mnPozd7TpVpTcCyjiMt6tSTL8VpWpcxbxO6qzFJ50IHsfM0i95MDN+NAIzY9dOOR3FP
zZ2LxZycT6a6Z7naLv0Lbv155KOiTABZsakKVBS5tjaGePmtl/yo/vvLBTtS6MVOdsZw9PnTy8Va
QYPiZBiJNgk3rov8carjQCfYBcrRn8j76MA6zXyQClIj5j0j0yoVhMxdpMiJGaI9szfYx10kSSBW
cBJZMNez1iIzwxBwSgDuM2gwwrU4A5bZHMztu3fCOVP40sSHk5DFdXyMDwcReNuZ++xb/F+lPwES
Foe1gZX8SiNDNkiGdjBbhRR7ezgpra2l/tD2DnbSf2G5cReswyLspAASq8vqxWmyqn2H53Ixud55
RfX7N6lr3V5qov2ltPugoEAYOjnBFtuOGRQTgbDk99RkoBWI7jff6CrqLy8+WdPWTl0y4cXTTzWc
ccG5+hLYjR3IaOLMsLbiPnkO2WeBMcWS1eTnQLnVosnjBiicc3tsyQSo4bys3otOUxXzB7fCRco4
76sYx2Ml9JghV3UfUC5UhJB1G8NKwDZ/0RqfYh17AL3SxuUB4s01bTvjOuRWdXpSBqh1j7d48qpL
0mASW6wWaJnBJB1PgUXoJUXkY5W8o/tcKxGGSmZbrz6keuuq2qMOmrxFw0irWfp/ZaByT5nIstHF
zeuRbpYFLV0fHydUiymZMTVNkhicr0weGtiOl9jY/bu3RqOSwsn4CPiAP7TPGyDnjsTuZZ66RBS/
F9c6RTLnDIv2mpw1cUL9InujRL+wUXRB+kcPQBiNu76x/VFK1lv9L4L+2OptW0XeilKmEOWy+YV2
9nIRbzP5xaDOrfTTE0EPnsEBflDBhwGnJNeXxBZoBQN5Hcs4vdfVyFyGsdULcwz8nq4Ld3jnNJ8Q
7CpvVBjNnsRVR9lEsw1LOOsPuUIctgwrd+DL8Kzjx1f3xqTWMZL/3BNLvHYMDJjsE9M0VJUNXYvQ
9LROunnKl58cwli2OwBJcUTWgxOaQqAoUR7IeLYfK2dZPzoM587glMqI4OvhLLAq0zJ/9RsFjiYK
eqQQBzKHOffwDOCYrG+psEPyti8mP85EYJJuPFNen7MF9TVbkKv0Pi0Tna5MGIP3yIXTUilECusp
UtdHbyF0pnGolNMdMQHJE7JJSJ0QKLXyEwpiscOIESza3OaUthvU+sFsFJwKqGEC3O/OcXt1QgDu
Q19E3PV9CODNgDuDWQYHyK6cpxchiSu/yKOTxeN0Y4lXCVoBPuEpqAGc1bnLX9WCo1NtTf231JW+
l4EiwB9+ZWzuttElmkVgSUBOXhzdCrCCkbtLJOnddky29W0/sjiJzd/sy8+KTZyu442g7j8oAL3+
RZdHpd9Z3O1gvjQsm/8O/2+xEDoO0JfROy6TtNP+Ug6i/opXcme4LtJ+9DoPPye1li+4clke57a1
hIuR7lMbzzhIYN7RAx2FpTcGStCJFhIsDRfWyciMNcDsOwEEiuB/DoH5cEwX7o8+eQBEumaMVfu4
yqf3/B8yHY/RNDVXB5FKYUmOycyk9GApj/88vWoQBbUU7CG0yZ2y+BVFznQRxQUiYBMg2bJqAk5N
Ip9dICPCHz4rrFSQ7pJfXkT8py3/rdd78EXk1hbl6GvFwglSb8WVAnH/yhUtkCks2eU5JQUQdCYb
AjrRbvQeaJjuoeHeRbK6qa/NEkONMPpEk80i0p4s5SunL40H7KVVICs7KEoQ1a8pTSelzOTf4Ben
t49vZhC6OtfEtx5QFzAGCcFsZSozRK/Qg39nwl2WLCXIMYNH4meP4tzU1V3XLAxwPm/AQWLYCdtc
qbK/sB7ylP93FcbFilOTLSfW6dgABWORP6Wj+gTC7bnANR2LBRBQOtL8P1HCwJ92G0a4hcRbT7CZ
8G3V99tnKmBjH3n63W/GNZ5X3OxvDruPeskiApYzZIEsxU+qZjZ4gD/j2S1jSx+zwQOyDyJON+8O
X9xllS2Hc9KDz8awaIKw8bcGUd2OVZS70I99V8gvdchUeO3wUTRwKTqthVyG9CrfQnqqmIH0biia
tLom/1ci2ybMnOmEZgoHIb5cd/cTYUeCLCU9Jeqn27IHCIJy+EcPymgJbJqoosxLNYBUhuaQ++qy
ahY2WGnAbr+579pQCygYBHVw62VE3GKPD1C32kZmtE9Vq/GgVnCTrIbvWKLyviGtPl/SZWVpIhRc
6gaf9YSfRMWbAPzJUL8SA4T7pALkHUzru/MaPgVQfb5owzhY3mdtVWvexDmNyfm1cS1CZhtg1v3o
fiDbYLsbV9rcMIHqIedm7h8Atc+x+42ARq2n7Px010NZIPhDooQpgwS8b1ZebszRHu6OLUJr5OUr
CoIyZPAi+pRE29ixfC/kTWaxeOJ2Me46cRDEV58oLs49tIo+3dk1R3N70kKewQhlbZvz6nTVWcwp
AT6J9WymV2D4tVY/wDBjX/PKdMm5UJLKUrQEhF7dEwi4/8wX3Zf66jSrK2hFnbkq+rVcslHsCE7/
k6MDLXUnyxtEi0HWdnlCZYpGqBp6AArijXpfptVdzqXsfB9Sf8SYg1+4VTfJlOncMSBM/NCXE7FE
4DqdBs7SvdhwMzXWOvGLnHz6DAjzRgac+RyY6EnlPtHv53FB8wjQDpxxWbRKm+/8MaqdBB/mUAxD
EK+dThlUFEXSyQkMKmcCw4IVAqx67XReFPYCNr12HiX9LRcL/dUT+JVy9TmvSXF8vYAj6MlWGD0O
D9+bOoIPcq2wRKszatHXclaZdp3/JhbPUww6ntC5hl+9DbcurwkeiHEzWkGb67ipYEPLDDBZrlWc
unCqojrzmn53kG5oJADcWF0zBbA3R7QzWaqr6gQanIqayCM5h92KbOj5yOC/Xf1M1bmAhVd9hURQ
kobPXcxKO0X0WAoNBUl+zTCMW72lqi28zqOBTXVrs4t2sVVQ4rsso8fZnxpY5YBZVADwskdTdNgL
tQLcNY3CTt3RnaSeODAwosId9PdjtGW2A0rKoXVnzQbq0zXdnbu/CAQkI/+aS0A7t8fZJ0GOkXVM
MGnXs6JbRKMY+bidebeWnK4VkzrJCYkLwa098SS7LuOXKclfxN0wcwcUSVhKyGqvVAdWhynqioS1
LvrqsEydCcFggYwkkIzrLrcDTqb8ha/Xp6/5QibdynfvJMEGx+N9nQsvhZR0Z7bxWFAHnKrU2tj6
AFSfP2ugA5iQIEvrfmibhTRYIV4CtN66b69kovlHU1XBal9ju19B3lreZprF11vdjvlzXMlkRyLi
qX3yu7ZMxElsMDFBLFzec+lLQjJ/zSPMjjrI/NsPFEJCPNNkoaOKLclyseT9pxEeRFo3BPZ7VPh0
/dkubAnHSU6PmO/dsWPrzJpgVy16VdCUzcloD1wTw5l+0sXmlfe/f1tIi/sDDK8A97rHcM163Cyi
f63FCVoySQAjGqwyhsGwubr/aD0E0rvVPCs5DNx5vTepmkeFgvTtu2l5eepPyvhKW1+612MPbt8J
0TCY5GbesgDGouAkcCzYCKB9hHNp9tH1ESUQXaKiA8prrfAgAxqDvQQKN+cRvGzyi7wamJj68/m1
Ie5KQr6t+ElJsTZwupUr6Et0rO6Uz70lpDvYM5YJCrwVpCsWm/1BbodId2J+r4gz4WamdBbcI44Y
qadv2DCe9N4G0zzoKrJqocUf65bDxpZBYSOQ0YhFJozkDSBSqfLLpMcltVyA7OH9oYGB7gFfxicL
PVYBkoQbm48kETE1Bk96USmlYETwRLuQepfYx6/pWhDqjvAmm2d7UDOQxEax0/CftSA/k/eblerM
qn94TkPfPLNofMZdNYR6a1Cu5QeAwwERi1HwNEPAlX1/FH/PCRAq1aPT0t79zj1DKnl/7v0uWRM8
KHlo7CU18LFaw5HP/sQMRxVua/TepkCr22vd0PjW4jsw6JetabxNpUjP5koM4KFTgxnSUpXSkf8D
EZeTWHS6qG8enx0o8Zis4Od0AFiZuu5YIwBh20kOftcrWzvRlGLSEina5LHBubMn/7r5+FKDeNxs
1K8PIFviUbeBpKc+w3+RqIVjJdzvssitslNlPZ+ZvmuLn3MHDXPP6uk6cXbe9+piiP/7bicFhnQb
0KBr0eNjMbx2Y7PvNV0SchJSwy77nlJblHam4b2yj15UCvwd7hYxKnQC/K5GMexGfIA+9n4iTX4m
4IRTHS98OyBVGhO8iYzu9Rtx6cJ6Ugc/xrcgEZHwep3BBr6xjiOYs9VBAz+Rhvhke0Wa8fLoSl1X
ibnr00Z1BpyytcltXWe/LWBcDJL4uQ16ILhFmvlHfExWHzyd/kCefdcHBLe/czlwgd4poK6ak2cO
jGAIPco7pHeRkMUxRgH5qawX447x0ivD9XiwU3aZuXysRnKCkDD30L0kzdVy1YhxXLLk89bUiIkW
6mSuVmX0sn7me4yBgoSimpCStq5Z7/jX3xSxOGdqhR03mTiB3XWum1Vo8txgfHYy0PfLVq3zLCpk
/KoaPa3Wl9zL0y2XBRg7Z27ANGawUVUmzC0KGv9wAAbFKgvhBTl8mFKO6D7mDAcUF3n7rbaKc2Y7
svcPXO724GExpVftiaXBOgqQKdh4T+VrqMCIClyrkQHbHBETYUdGDqnmdh/vYO9tSbBXpSUgdarM
l7blEJ4Arq6Rgjzo6h5CyIWSRwdvKpXkCSxaysEpBr7G+k8hYRb0XfdGqC1ZY7UIBWeflVoLhb66
DcgZGrGajEZzULlQVKSV7iVotIvM3EzdE4yKTOu0NPAgrM7QSMolJw97H0ZPpPGpBAyLSPfuSWwu
HVtV0/3b2VUynSb01KcmSvurTjBSSHyRwpJFOSbGTqz4EcRlI6U3ccJXAK8IYzvFkg6Jxg8/O4QF
jbE3ZWd46PdLAN5oTHFqnuhmDMoo2wylEAtxzZnTNc09/9wZZWSX0QLcS5k0jcGru/S3JYUP0YYB
qRItR0WrJVo+eJUUPsPYX1fXYegGxT/zf35pbnoGT3+DeoIPNUJUJKiEfCYfoXHHPlw77vqp5Ddx
G878KxQ7vjYPBtIAKMyG2P16zVDO36mVhoPMZ06eMO0y3efe6scSMkSeAD4oDVnn26VZ7NX6CVNZ
aB+VgvDgMq4LCnoQqO/p+hRMXZWH9bwsqtlaNTMxp0+0AxJFsWH0IBfT3hsNIE0zovgIkLlSNftC
2mpPO4KsGklk2pQGYK11wFvsNJbgBGc6muZ69uMLSYbYWBf1G3AocrVWBdDT4ioW6DmMpY41L8lH
PKbbWW8+kq+ZHJWTztDyzLMtpqtqGycaNtlmGZPgIDgURUCEnRBaqsHghetKAOE62+Dg4q/MuwVY
6ObutgmIUIkPVI/UfnBNVdcSyE0GbYXjJZLVygQpJ4vJ8SPu8Z6VoIJXrN+mgulX1Refl4cZsEnu
OEOuzi7VbYj1GU8yZIv9HTfE/bBCMr6P9wyl53wPRITWnC5YLCxnQPMkvWhHf8onWJPqrgPLKcyy
sTPlcqbm/4rGDgq8VMiOI2SE2Bi98HIMIl0wWnt4gvDwStVqmwkSJMGI47774DoYu4kz31LDR+Ud
hEviyDcA9WxNRvU8DPCKMwibpHWnSUw5XFMUHxkluUQ/81AeRf5nVtFWn65Ds4+yuNl71rAOmd0P
ybQcKW6ndOsAnjSvT2aZJbqEEh0lBBLd+WXHNatac5yUzxVG02CrmYcVH16jvQM3OX0psxjiEyeU
z2NJ0vy0cQVQ51WNQVnbJhwzBxbZDTvxnZjwtdWq1gZvJcks2L4KILxx/Tb97wqga1n8XE9HlhBV
11dJNzoWgUgujqJNTPP/Utwx9ZsWzmmZWHKBehFD0vrG0pfrlxLEaLCVhtfFTj+LzkqsGvD38a2z
dfBzaAiTJdycnYX6ggVQ+b4aDcIkgN+dprpP7IUzCgwz7CPWC59MXti7Dj1xmfJtl/khC9sTD+Pj
JLm96L7iOdezW3io8PnRTOMnvqgld4CQYtslm7l//IMhz/Zo6ySuj8K7HOBmYa3n4vcXSemGFg5/
NQXgsN7090OQbPTUvMAHsMB4M2s+Y+HMCgrsKxB+S4RyHZk4RyG1xxF8obt1rmbHMBV+M89KOIqJ
uy2STFUsvDBwPBCwIVoNgKeC+z30z0LcjTZTZsPU/xKxEJeuqk1bJBSBk2IPh2f6Z7EEiBuE2Sm+
NMNcfdvGCkZAILJpVe1wbrlbqrQcJBdCrvIAQW1WmC8jKLoAsEkPBkFYe7747LYMXEeh0xiuodIr
Gk+VJ+QNU7Pp873XdIk3DHL2wP1bVib6BvVKiudyrA3l1Mf6N30qs3vCRzmvfbDrOLsISBTAJpBX
tIp+W8jbUWcFJnPqgbJ99cMZ5HIIfxC5K4dcvGLLCQQgGj4qfVxhScML1hcl+H7cPZwk0aP1f10n
lFGbpRZY6AwdpaTzkI6e9G9iwUrrqboxIJt81BTv6QKHQ1D/9wskH0hFzCNK4+F8T4bTN+dm3x8B
DqMM6zUTcRdli93hdUrvOsIkxaCrzlyuU5rGZMcWoxHx6VLE1zmIUUpZK4yepY0g0AMAfZ4uf+Rn
3gWQXQ/wzorCD9gNSEryf6L4ZgCFooCAqj4epQqIFDTpZ7DLtjR7mvsZw/XiSlIoQcrCH52T1LR1
joNJN/fAfclJ91Io8cAcIMK7wCZJbSPBYK7B/PLxN9pvwFV3tdCoL7vuS8gaOmY8310nuNj81Eyo
nr3DhNM2Fx37bo/4zq6xJy4AmDuxKD4XXjf3qU+zp7SJhYvjDihrUmQPw32N6kFmLdtjqqURRSyp
yfykLB/QnqVq1oI5qf/3Nj3l10DGzEfduo5uiu3U+F8GdoJKR+YvFTdcC5svaHIbGq7AwRvLfP6Z
bMcWVCAqubpQw5VO5O9yOnFjrQvgJn+sS0uyI0sw4vs4kT/Xa6KWQMdf6bHZ7t300jtmYhwY3XDf
PO2T+oXWDQijsPo18b0ubkv8WZCCRPXa2rSDqw1bENbu+mBypdRc3bXnyayVivFzm/P/sfK33jkt
82AcnXYGN4T4x9MSk9QccHcm9lSIzfNqxIeRiWJ6uK2E9B/LMJk3AC1P5v1GM7WUCz3tOp3VR2GR
co3dk8IRRJxGGmyqhPYqIp9wzkvhkYRzlGpuZwhg/TRm9zH/a1w0mHkQ99RnJ7r4s3nQLf6yEXm5
HUxkz+1y0vnEDTwtUarKYVPuv/tOjMw6axCgabDF6oUakl/thmzkpK5aNaL2UKYowc9VTmmmAzDP
TpN5tA1hhoUpIRyqXcXvvYOZSmk1wSeaDg20ZTf1UEkkiNcCWjKIxd99URoAEzOg9fAWfffww9jW
/F2iIqouPbIhxAngAA6xNQGoXUBdMmmCmojkXGqlSD/T0qLdyoekfUbxWq7fU59qCCCJaAftcfQS
2/+KhbSY7XFNjJ7Ijvf+yLjA0/1+wQZg8h71sP0N780A91cf99BFzJaUcWkkDOxUfR/MtFVOo0VC
66Gjbn1uiTGk6JcUs25zSyTgBEF5sY+f131Z750/FJTBNEwYzQ24fR2VTt1xG+MPcJV+GIhSbN4u
KuaZ0mdpUdOC8ce1dr0FO2mDtnqEDDtJ7EWQH7VZKJBacP0lOUw/EHR88LbQ+x7bnexyU4mEZQVW
jmyxvVOV9wHaEqORnyoNuXJouCvJ3JUU+Vu2urXXh7ynhEWuxRLJ7rz2avsgMhhvsDXNpIJKevQt
UC6l28nb8LFi+cAkppjuBBzH741mwCvnzb0XL/zbqVEJ/USLTH7b4Vkmgd3sPwZGmflekfdzNLd7
cJ3R3I5u2eDBHOcw6W2mJ7MFBOnr+wPUXOLjXz8paO8uprd/StDzhXwbSKFMHjdHNxSbMABvQrjs
jIWhwQVYj+9IAQ/Zqk+kFHB1vLHHPmBbZ3zJnJO11tI86ZSI4FptUlv2vkeqDWFdXdlfDvXe7G4W
3s6Gtb7eydG3xgPyyyf6mazyxLzcZO+OVQvouJTxtVwyzKYOUxqnVDpfkcrGYzHQgIni3VnXOM3q
taRSoIe2MeK7S2b8bGYLZ7ZoKH0YYLVhLjSCdvtX9Kd0nxpOVyiZg6qbo84mN/UdwF9KTyFQlMhQ
9iu+TmF8JXmImCd2R4kVcb+UDtJ40ccQ6ghfLNepKF59nmRTrsbd1mcJk4aUmfAmdtGtezM95Imw
nf0ofUKQOwA9H9VT5ahxViOIfh5SSUcaPYm9+XR5aANu/Fxx4JngvF7YEPKZOu7YyjUGT/yekVH+
crIyWlr4jCQ2O557MvKfseArlIUNXacyRpyXreJUvfPrPrP6zBhSsX6KjJS3N5tJSH2SuLqA9rHq
Tp7DJsTLU823x+GwWmPoWGCWg2X4p94YCpzIC+xwjcCRrUfdqbhU1RNUlB+IIYpfOGR6FvTBn8h+
qmDEp1DsJZJMbyiKBw9MioscH/5Gm0OVOpiYpG/ruRTxS0zL81UfKUy9IT9RQCpCpGbLH6YnpcHs
qCA32bGZQ5pmbGNBGefTHCrh/NAr5DjaI/Asc4CNib4hWX1a7AT1zY0r+wBnaDE8402s0JJ/YCH7
nVuhSqfQplRHH4ohQ6WBlt6iRgyJVBnYgawNqbKdWv5xZsNfQQXT840w5rt+kvQNxPUc2MP/0MY0
oc6jum1lQMtRxR3NJVfz/DbfloA9N+eVYywERTAEWur4HnT9OBoBCUwDcxts81V6p1SPoPRWjOvi
4smtRvC2PyYevpnl7djApLYDImm9Sgy96hOS9ImLvCtluAd56zGUzeNH7cC5lryYN9aHpOvHch+r
D3kG+YktexRIwXhxsoTLEKFd4wbAd8sY/CCo5D/3ACDHAebrYFJ0szNfXWQvlOfxXQwTWVoCVHmi
uLk/XN3642fdPHvs8nC7GRP2VUBvjHM2oanR5rI/L1GwOnG5mceMcIJipUC1LXUE1a4wljTZ9Tib
w+5hKwCD7X/sqJV6g5t+Ct75lGlGUmZ5q7/EcGt1b979RutkUkFAAqqqXrkSKaEVstg8zGQvPQMj
+pQ9tFYx41rFd1Pfq5FCDbE9yZBhG3Fp2tkp5XyMSj2Iz9xV31256+BCoHidytmljT0iQgF5c/2S
T0uv6F119WvRJaU+PXrbIR2Jvb/3xrtv+v0ESm8Mm7QMwQtgz3CCOAjoXvJm4/fvFluNpyvdzfvE
7WEH8ZIQL5s+SUjTD2k/5UnTi63iJAJxIUOPSm6uzg/0WVmZ422wCYu5TkI+NgyDPWDmbxkDQnn5
CDyAfQJuuq7VySbnWiKb9CE9JzbpVcn1aTBjH1DN3PbbHVh0lwZEHDrOkuaT9dmGx/XsICKzl0R3
tmR29uyNo4l+mD/dXLyavQyHup8haGOnDybq8eGxecy18XhCk0A+7nZXQIn0DmVRR3qsWzSgQ2Vh
Cev1PHGOeS0mp231EHPg0971Xklek3zx1f4gt6BpqE6JGBXyxWgXNw/eTrgbn7OaNGc+CASB9bRO
4aC8CdeEbjJ5yt9ZZqu6fX+zsfBfcv+lapgiIezWDaSdUFr71rEEwIoLdHk/ef7CmmhU5xj4BOGy
VDkTKMAJy+DhL10zKQSDLIyxMEKe0eGiKFrWRRelfKmE8Ge1PcswdU6rphFBuUdOHaJjwl0FwBN9
gtJtXU+58FZjtCEa2bHw0DAj0LPJwD2vvmAdPUbsjLQ8ZDi/8MmSYz8aNXaDXLHDUq8Vob8650vb
o6VaJdb8FWSMac7wgN9r4CLflvh/epBylS20ppaaDLGG316u1hI1GKqwP2KCOOFimETi2BycL7YJ
ZfpNvUDhL/75waWRMbOofdI7oKclh3T68ojUY4F5A7i9imK44AkcEV4TuxAkhEZ8dXHoAOE9PU61
f9RLvupkFFxg+hXsQkJxrwk89bXP0uJL77NzOpz7PYQ7zhUA4WHEGs2bAsDS2OE+X2upsylvaUEf
Di+fk5Ux47QX0U3gq6cLBtSwQq7R5fv+oXfg/A88En3RXbIHt0VMnz9ewfmGEWv6bMUxdNCnVbwj
PqhFuU1Mw3hmGchgzbfMPWmzpvaU2YVE2MhcSELMsUYFBm3Bxu2YaUj4AMCtij48AjKfSwnqGSgk
3Kmj4Vr4LCd0ziCtv4UW/U72lnsGkzP8zG6WxMRrjvNN5PsyKtGCtdnT9Y4vU53KAvFZV+El+D00
3LBcUXW6p3urezdo0jHo6mfKdPcoX0+Nxgmo19vHR8YryJZs5ofP83w4YolDr6jrroW554jgMFDq
XddDfyqXNmAI72/S9iYwejUsLuQ/bh9oWpKLxPbho1RI06DQ0EaE7a0uaeNwAG6+ReqyXT6Wi2tr
zDoMpoRk6I2t7g9nCxA7g4axlj23dJILONShhb1DBznxhGKl7KFdLeu8W5vcp/PrtXoRNT43KU1g
gM2Btxh6H9Zc5jGMFx3diEt3EPEYYPupr0SGM2Dn2ZA078PjG3qFogxOg0qru3IXooi5RJPIzNxU
8dLcSB8Di1D/Pj8bKq1AMjoaIgpfSRj6hxOz27QvsRn449+zzhMXP5tIScTnpIXwLlkWJSsU7IQY
W36IJn+aSfBuzMeggh40AxiO5s1hp53rQkSoqdotCMju1up+DhTBObiZUbTAHU5HQKN4Uj2ClB3P
BaGP8U3+z6ROO8traLkEIm8RMaGMetGXZAPlFH8khbvTf64cPss1RWwBHA/TuS63QQyqq1Wt/4ts
yT49P+dYGS+z2fAfQCVATdVIocI2kd5ZAJBIEu/4hP3OWoGbcv+MtISSNK5LJgI79mFu26/gJZ8c
45IJW+rbJb+pwJJiblgnqaAnja+ddjf1D+s5gKxNxaGUTgXvMFBj7mv4flFylc+fFASHKP80QJYw
HUSIrfhAqsCbM/KRaFEkPQSJMRD2m3Thz42Iq85E+FnnYOlBMt4xKIgnNtZrP3oYj8+pbxgOan2O
AwOQewayBi+5FGDFaTZWyba+TscSErXZINJ42NswPo/J6F7jMyCu58TFtNgzUSRx7puMMzdewuZ/
E8DYMGtCJl4lxqQCKQ72uKSwO4eqajQFxsMEZ7gqlmKtsy6yDfjVbHihii+1078ubNCCJYTn6DOC
cqQtEvVFwQ0m1kB11Les2BfBI/keO6lN7LE6xvtE9XBNYYwr3sZcasb/ZHjgZ6Ag5Owr0/bf1of2
vLuPhv/mJ67my5kUyj4tTqO73wdiATu6nlQnd4rzkAYg3joNOEllIZsDFsBbgGPTNVLZqw/UIY0t
S0ACHuSYutaxaMsvFn/qnCy/bv3D6qcpxle6czrBGYhR/j613NAZfJJlrk86fnY/k2r0QdvK3fVW
7mnST7rRjH9hi2nk4SKIK61Nt8eC+7dqIRsV6xybUtn/jER+Qi685Dc7v1DDsX79GDsUP9XXculp
f9+YqmyHD8x2sIMohFK4WXi7yXlT8/a2ryf12RMGOGqOcusEJOb2zgZ72z0Iw+oHp+AYbyqOBO8t
sIOdMDivZmag9s9e9jgJiFETwT/TuDZd5r2LnHMInfGIgM64afOJNlwqmZ0m2TEKRrodyLs/uIn7
US2ondbFTk4raZNY1rK8rNpA14g4BESht8VWt4OwDBs1A487YLH9Lxex8CLZkM8Jx0VV6q94thZS
u4EZvMFI4lEcfrynCI0JOEFYXTVS8ORQllnHH8JF+o8bgZpr2Z4a06ThEw3T1xUEHp//DGEexzT9
WdgZu+5SjHuSRr4l/1YhskPtp76Cug0XDiOHAyiG1Dywh0xruXS9bWSSWSn6xMZTGEKnAg5+8O9t
kCWwV/895gD4D8aCenvpZGyY78fiqivlgEY65JYfTTXnVbcbapqMLhTV80KQ1CIROJzvUUqvc6Hv
Y5znWQhj6w8zHQ+avvXaMG8snyH+dIGrrBje/OLTv3h5YnbsacH0TJ2zbUxH7Lt1CxRjQYl832RM
fbpImO14r8RbkIfXMktjrmJLUZoZpbGS/5rVEdZqbqa5s1GyE+Eve90aYAZ82lVgl1dgC8KT5U2r
7rrBIU3YqJScQAAvf8bhWGCk7LvpTFv+VLA0M2E0XJejJT4q1fboVdM/Htkgkug4L4U4zwVNJfz3
LgM8G7eLMIhWCW312JAUPG4m1Ap1g1k19HkLoxNON4wfsxXqpEjIfmJFjiZ8C7c4ov3LvxTjHq7U
NX00egd5s9F2Gh5i63/dPXOkadV51qVcQFUK2+ddO90kkpslfI3H734VT50SV5essMMH50grd8pT
4+b2y7B2kVR0bNmT69Db8TtS8WszM4FaMhE/CWWh4nbdkdX/sXfUxP013vLajfGozWXenqsRl47i
/qF6asq80q/fKUu1dVG0rVLrUuBQ+y1PX+lOONfik8nC7gsT0ZC6UccdX/XXygHEsZiUKqqwZM6X
8gaegoGO0Bc+WACELT2RWxtaV0DUZfUzbX6FEQd5jo8397pB0JdmxWC2GFvkgYoTRJl38MbYDDXZ
pscTkv8ic99/ACzQmED9abZgLcwDvw0LW9YL2Krp7TMGimIbUe5Qrqzx0RHRNG0aUDVfF5ajfAEO
616R6VbKJXNktmyr4MAlk4NTnmkTMwe2jcve6/eKfm0A7d35qXPZTSgmSPrIoLN3+D7zdRBvSuA6
Rp1q1WgysTiSPILDyHUwUyjPEXR6K8Y+RNTIgTDFtBUDDP5r2wYkwRAxQYHnpRKcsBkJykIkHa7h
5IELEZmob3eElbHSqoA8B0RVOQde0R31i6EkZH6+de8njN2jaqZlHBhCkLPDqccuDGtAeQrZ/yl6
VzGvINWWtBNLHVRNhmY6jfQDoc0ynQz+JGts6fphGCGILthLOElzN4L5Mow0oH2g+ik+F0UgBUq9
Rgf3ksPSlxTXGeegdnSDUmYoLwumHgf5KgunyApM+MPp0cy5aJXHW6eK/r7U7IW8mYujw0e2+xzW
IF4Jlfyf4bq/lTKFtvHdkXg4kgY8GDt72YZKSWb6K8639rxdK8QxmwI4weg7cv5H2jB2McB7zhxS
ZZPlgrpcGy8+xQ5aKonOZtPJ3h3a93jkLJ35fS3nnLAaK+Ylp2de4vSc7k9i/Dd5LE7JDe5XeAvy
y0Odsg2et/oIRwzXSNOl6dkXASHF5A54HYrfUFdZDzBZSwJzeI/JTYiUUVMKMHw2t42pfUfb4bvE
dNe6vVV5NjRFSIC6WeRHM7pNEzYc/xaR83UTDdrvhNl6nRlG4QDX2VEmB0mbZwUFkGmGQVjmpqUU
uTCxJTV/n+py2CZAz1NR/7J3go4pjg6LbY2ggLaCvF/axvx+yzDYoh7QeVcPCz8hLJwvTT8TgSE+
hLtp4XuxcQ7vcr9s1MEYLwbm/zqBgfJdVnVCUMLXyf4M+zNDwbXqos9Nbt8yhMkG1xsuVe3LS5vO
Y1BHA3es5DVcn6wHrH5/kHppHc9Xyzkm59cTqkFghROQsuAp0PsN78QeZhBMfTkGOHF8H+65CKKQ
pVgGl8cYQeb5qwDl2jtUdVwl467fA6a/0tgMid80a8H5LzBgzyY7HQ/uzze8a6AwCc6916O/Lsie
vOgl38n4OSEH3GgzQW+rDYQkDrIFr+SRIBNGFBWspQ9pwfaMJzb7FzLYXEnq5/20g87b5DTlCToQ
fYjxX0JytsQ6pCj5o9qDhxG2qLAzfBDt0Waz2sPrW33dvX3r7pgA+qYdBJ1tG0YFszNhSIZnQlHB
iSiOHgYflddvxFAD8odcIehqP+jTHffQJ0cD5HuhKgVq3qnAcckztjDIm3BCsZalWOEjLXbzmeq6
V9xeLS1nyNnfV0EAuhEcBe57pqCROebfV+Iit9qtD0tuv8S5+y36RAVF289bGXlQI1xmcYLvVbJZ
3lGrwnl22BFUFWR7nBA+v3sioTQpQ3CQ2Ze99pOA75fE4iTT1j0WedUBy3SobnuBvCNQ2hHBnrFo
c9r5NlCZuF1MCZn7nGwlpk8URuKeC41bHUMBRM3NTs4UFlJByfrdsItMIem+eIjFx/3wEZN/j4S/
HmMPWJPxmQaYnOM2O6WF2955Gk6xpD3U/Nh0IK6Lm9ejCOHTVf2Rcsy8w/oZJBd9zWAeqM0db6nx
ANQGg39nHjs4ECAB4rTnv/4723OSwpGMkInvtUqP1EVyqo3fvWI8+MKOtQ2g6einoqEkSbFuiTpy
EtncHnCdudyjowrveGrV9fT+avnGatzOYOS1tLbHpoIZlDSSETvbAohfXOC2DxI0WKDk5xH7w6K+
cUPPx0HV7Sd2VnqpJo4XQGkB3Lp+knGwccwKMaYeY1D4nkwW49IorpQwl7oB022AdxBs9UWbY6am
TF2ytFaLMj9YkI65OxoONKe1QMIBKXXPqlH/9UiHvpMsY8Q5VKZFFdeFbty7UrmAd0DHZV5vAcxd
AA/ghsTctn1QvP0MvuUO3xAV8ekh6IngdJYKPmjG1HyD1RNcVBbJIQBBX3dSDHPgaj5cE3DPKmcS
4ivkgrjQ7haY0Bhf+/U57VVWT+6qfNBKyinRCl+hxqayDnk7sUC5dZjhsp5jk03MM0NPgWdoBNUo
+LUad54B6GeuWsbG1JLkoBTQ9xfD4UqfCveSge9N9fwCqYApmCUNNrsuZaJn0qFFtTP/04q/7m4M
CzK4IBX8T6IiuhiYdZlOUS2ukm/VbjgqimtXIpkSxitzUcRYZwAcNmIc2BvBWfY96JY1YgRh2vDX
P6BL9+C07pF6jW2vb/ypjXAfDjVAydclCJP9DQ/aUtAnYIZCAXpTBCXH16z3c6JceGYRlOxptNAR
kkL05hoILXLBMYb2Eq3lt8xUYBus5uKn2q/YZe1il6fMiVhMfvW6rJ7ga3MgsaqDcsWzAEy7zwIm
2/13677O80u9gA+1wqnL1FZBmCU/XOH9hPp9H0lHd3rQGzy5csWP99Xor4RQUOWsdifLu9FYWflZ
FdWM5z0/D10mhmXHlQJXFp7mRUIk16hMkoUh7mIyHprXkj+CnI+GLDZAAQ1B+VSlivo2N+D89eSs
dqEN0KWW+x/JFtXPun4GfYUYyE0qJo/gb9f3eJP249kWm8jrNa/qIF0nUkeA9AHe9w34EH5SyHN8
/iXSS+A4SFfzxdp0msHGh2/JZNIdOzJebm8LxuDHv2edBFw/vFSpdKE5pPjZxCo4E6cGJ1tGTOR8
PSqUy5AHyzWl1FZAuhKnv7aRnCevBNR1xfj2lBA/F4mmt+MD17wZ7HKO4bcYLnyWSaXDex6nX4OK
xri89QVGmwVobzxSLtv83K+2gb51lVGhuqg7NDEvpgrO/jX7k3i+H0heee1i4Bb7rb/nKN2drggn
WA0pF4aN3Pmqyg65Er5VUonw/DcJstUuUvT1uI89vXbrssiue3bzxMiiPgX56UUGQt0jjlzGHtij
1ijUD5u/9iVizc+sI4SnOKrhjIPmueBcBV99wJsFXgF+crgx6ZBlRI+rp9uG1UxKMAUl7zXjmZiT
Jc1eQHEnzM2EYHpgr+Ke0LjMJ/jBrAcgvOMHa8F4WZErSw6JCwJhoSzdZr4jErlVm/UyAatPfXyk
Em51jUnVz+S65WmatgwXHo6+wJt22ak8rLzYIMQZqe57oxODPZp8KTdrQR1o0PLmAcizlmmRhGYI
7b6XQVfM8LoEtyFd35ZfnVG4OVQ28UXCqRhr6YSKa7PH03Xghug3bZgaTtqXCv9sZxFWX8AKKdJH
5tongt2is6wHYMObLAhcM6BmoxCsOcO4Wp73EI/CEngsi+cXsWAubdZWNrE3C86YONjBr1VOuY9S
ctHMLL7fXbRJppm/Kw6g7vlSJCTDLY7roSqU39HDgd/jgFjUeMaIkDtOzLma4dNJ8/IrwG/MaHLZ
QRo/1LEF4CfWq0CeKiOFVk6O3zHrVjdsUjlYR8ZskP4vLxbzt+RQw4RVPjhmoHQS9JydmIZ06vQu
YBqWjiEGIpU4UsAyM3EEF9qMiz3cqYv5XNcgUgNHQR+hqSxeraNVyjF4whOusRMBKIg23gFTdNsa
Q9gmQHpr/yohFkQ0UW8KFPym5wmEA71jbh3K3P4oE66Jsxb8UtjWVx8rEdSZc38h2prG7l7dofGb
VDFMBTYIB52GAYIIHONH5htyPk232T/r1F+PIDCWOga3AmSARXF/DYWRJJRkco4UcoucJ5NX35hR
xZ2SE9mhdXyiIMZkWlvV7Fp1SByKFOKriKyfv6E/LdFEQLzXvjoWoer0jB1kwqegSpU0PNIW5fv8
jG3rnCQCh/rzoRb3xR5McxnhvExhDoKsMT8BbdAJWGNWvKSby1H40jR9RiNE8DFJzQ4GMZIWwJ3T
xRe2C7Wk1UmfPbZ7L5GE5/h2PsiurRBr7FHD/2405jTT2hR1IUr6zXyRvTIgaBVRT+lpkaLQh2pl
CqpYANISZ9tTDI/5zJ6GJ9tL781YGCjxus3NE5jaZxrqyf/CyP9oyX0u3Mvye5zETKdoKpVSkqma
BPGD690YH82D1qMFFR8e6RdcaM9O0CcbtBAHgyQlwvxDZfI3GBgsZJPrb7YpWvee2rmWwt2HN8Bj
Hn7BHM4b7upEqO7wZzCv+c7cDnUCGVzZ/K9BhR9b6+AurhIAlcdeb+u3UY+RUUyB4jzxYvCmyigo
y8Ib7HbCenfdQAYK6Mk65gl1EZhjOz7HIj7L7PpECHKUPeK0HjWyUkkojaesCXl93SVM79RL0kwe
0Fy4XiqFVErDAY0ucaUfFYEI9rTedB6/S1nFTzPe5JDk8hJUFWvrKpGoNsmD0VjHQ5whneTTOEkG
ieHJ4lsHzatveKKaMpkgFgkpdBB1tfpdcttNDuL0Ef3WWahYzlmQ1gCnlzfAalJggMUgIzea8soG
UITmMmJVPrk2uDKSYE5B4y/Zi/yY2loRgyvlFK7Syb8Uzt57aJK5C0jpO+J0OM/Lk42NvjjMuPUc
PyOW9gSMeOzKR9ZSwjeaZZ3cFyLrPN8tIcVywdwwNHDlNdo8Yb21JzMapVicboJ0A0D1J3WJskJT
F4FZyizTAX5r7lD/9+5VwzKmsNzmPqdK/aTUnqkC7WcpmCYq8+tna4eEOaY5fu/wU4Km62PAPM+V
uT8s9KXj//XZ2UGqt/kZzBnVE1N1xD2Y0o0TR9BfOSZfbaUUmtIzc8QgNkGuAHoYdHmlhF6kYwoH
zIeSv8c8ME8vjxK7QDS8QYg90oG0RdkRg3w8BlSmygEgft1YQiJX+t32aFrXKg+aQ7jRhHUcmlTA
i4DmEyDh09rO7qcyYLepfIn4iPCtuRDcmVDzCzIbQNrcPa4Wfynnety9hOPaxwvr+iWyECqXNKNJ
S1bMWIg5Y1uGzcbYZK2ChuPPxQMolFUcpXNkFsI0MuSy/TpO4rWpnAoZjj13UIpBMHWoGSn23UCA
cpgnHdIC+8syySnSb3OfAOL/HAyEmSHZz9OrfsZ49/2Q2ffVSJUPAp8o7WGph2VZikmoCoKtkUQe
/gooebja2E5RifABY5WKbkwIVwpt0O/YXfV1k1D0MYHEo7EKQccnJjhyZk/JUTHmW031p16ngbUH
fnlkNHls9ZTXWGRELWwnGCkP21I/9DNoGfw4JV8XDXlNtXoLbvRypOlu/LJh8coi3Mv1PmK0JmS6
O2ybFI/nAUtw3H52JGTFe0oXAg3G2OqfTsct+lZkFEiF3QhmH4s8jruJdwe7Ocy4tvMT8JPDZ9+d
/IfSPeszy0CEDWrtT+j2x1F0GmWIGAD6uPnJKTyMBxo7Q+MUbTf5CxhxGiSiV9eEFBEx/JLk6D2q
Eqmdne1t/043/11dERnIMeGUJHMcUVwvdWVeZezOs84t7RZfiECXRwv1NbtGM5k21YkjsCcdLTGV
CeI0jL0/7HU9LlUIpMHy41aM9dEmFpHHFaQtsamYT5mYouy1q/Uh4n3I+sfU0YXDbgqSUkUHhSxu
KzsI//gYw8/zrvAtZEffoA4sfwGeSfPQUJwBeslm2aqLo8QMloQ5wL88CxfbOxA274yDunr5lBfT
aKqiWCy2aeREhVm8kq/w4XyORatsb/GL5eB/pDOIUMRVxsrEGbm30skIntymGftSdzbXC5FvdPYM
6GqnABYioG8XjJbeCXumENxP2L/uLDGW5stdGBFRG0XwO/9hlkFS5LM9LQFXjq/Z0pBtYXIaJu3s
xjqiVUykLU9etfUaRAH1IWWXFBOeSL1pzSfwzTgD3Ome3HnZFPpt1E9TvS3Dpj7UVrATECV8/Bnw
Uzj3BIOPwmdJo1FtSci8QADIQluRscoHlkUW++lLCU9BIlHr7I6TaIjJrhdHmd89TnFzqghtNL+b
HqgMcZWnsnISZKLTRKyNcSZUrVPOllhWXHZFHlOPUKs7qWFBdXV/vHL6V9OWZmZkltDai/NzmXYY
d5pgonTCZIFOqeUuoK7EHegjwQ07Omyq1U28Ctai7chfS3oKiTNTnVjf01S9U4QrIMqOjOXCmvaC
wF5RLYarkOKPB2KvbJMlPC0P253PYIycroi3BTGRJ5GdN6eqb5rVkbGTCF06ZV9JJ3gR+vknT4U/
ikpqkHoL12pqTn8iH3JKrZulGqfaS4/IGMRQXkpxHh6LTWe997X/pXTIw382Le//k+chtWAR//UR
iie8eepEw+dOirYuUCJ6RA+JaGhZVmHcWs6pwh7mG5LL5lSMHqXDj0FV2x53EhqsQjEWqZCrpM1R
qb/sLjWWyH5DzAruc/gcUXLt9IPN59aRq0FcPtnKaC3hUq5fuzUJySsb/Otlgf/A8uueAUJX2nh8
kXro4vlqmO7ir7fzPh6/Xbb6yAIwZOsU+z5xkuyiyzJbYJJKyWf4UEAkIBsUIW51g1f+v4hJr9QL
aiWHUnnffxFGmMWNsUrPmSENTFeQYjy1XRcTPn8Cqsi8AMovjX2ke/CVN8TUlzbzUuzMtxjddgaw
3VVvCptvOJVuTBVgd5uFVCVm7glQ3TtHblVTmsShl8OY5/tr8u65NWOpU/0u0SxAnNL3exxogF3T
39UlpQm/8WR6yt1bTJtY3yR5SCbKNlY3QVLs0pRW4HjHzf5b+pHjQZ1MxI7ZvTGjR+RdM26UxFqd
UdeFuAi0aFDBu2PiAGO119urWKkMrEHrC3Gq0lntkzt3Q047KjxLNhbhHwstb7uLnCMiwjiWgG1J
joiq8URi6I9dyoZnYxm9VTT07jfqDyRGEp6Lq9PzuCgjKTdXvwwqxtg9t4bNj1P0RT7wpO5kTEj1
mZcjscGt4ZBjGRdJV9M5vxcBkyDOfGzzX/mlIKohQErov43Bl2IhZ6aMqwqs3678FjIKPJBDiLcE
xqJ2UT4Ojd96g3e/jagO85LlaV/xe/zZTm+fM+w3Z69bX1AhegdFW79uKHjfiRW6qAdAcHKCd6hC
vbegNoTfpoi6WqxosxcUP+eL5gDHbbIOU8GL5kMxD7wHlXy2MU06WyZf2x5f+Z6uIl3Tq1kWiFm2
AWgtRMz0UXsiC1ROlIMdUGQ2JqpvBvi4qKnMQmUQppfZmuhQdZNBsQg/B+1tYqPQBKPFK/tjBmwH
QrgwrgPVKoBss12868iQZ4TmshCYKJ8HFQKZw3II0k6xgLcsmJLjafcaXYpgdGX7cRc+vKhi6JzJ
hyaQFoNMnAQZwEhcFipm0yP1WGPtuh9s8vUQNkYcneshiDDvpesMQUcPrqtBVRPJldRShWqxDPjm
p++B+M8vkC1jv1xgnF+PQfjb8yuHZcBb2+x5nstBu5pCmSGMknRJWLgyoGduwNTaXyjJ5gcnEQc3
/mo3ihozASCnI0ThdyfItTejCALnqSuVJta98Z8YIYY0/GTT/HVQDMigEYNBCRLbCDF9yRfyBeXc
YvdJnYtP+7J5obvEonvp4EUr5DRlf2/tbdOrgtIf+vSGcDvMusJ33qKr2BeGnsilkEaH2jPpv+Pr
2FzuOqSqDLcwJQISD2pak9Zj33kGA+O4OCXtnLXqtqw3L1bWI87yjcw27WzsC4+gVkAKKO5sh2HM
2xp+E8XX2LiprCXcHm92bQ/M31UZS9JEOtV2W2xT6gP+zfZa+u7aX9yFAmMJGSERlNpzPlwlK2GO
JaamsDk2OuQEY9iAI0xWGj+qMhE6tWyeokKMgSmbSGfJr1H92VTwzOcfyBLAi3UqbUL89OmwwrTN
zQIJ+gulSoMx7mvl1nyGU2Gdvl+rTULqaYuMmh8A9aVZfuN6ogyMW81fXdLcs4w6PPH2G+hRrxlZ
BITM+lv9ONKr9sVLBJLRp/nSMx1C/X55LzGB6p3GG2SIC4W2bDp4u0dHFK3dUfhniueiQ0B5rjCm
z+r1LNpXz3oweIPKTvwOIJ2hGONR6tX6SH1XeaavHJWIs7ewD0lmQPFDHkRZPsVbbbRoWtEWECkK
2g6rFdAtsY05TkRTSH8OoeILccHS4ovFgGcg19fnHVW+sEPfLRb+DiwP+O4gD/qgqw7C3AeBEpsw
q1Wv+k4o4qYKEs2dpjz1HS8KthxchkscnRFWwO4cknKWYI2FogXBT84QJeSnHDPF6Gi2I+9hU8C/
FllPWTppOlem2Zh/R/UnNCZP3D+mf++I+wtnwsApvSb5OoPytkguIuArFBcK6SodTHFQQ3RrJIN0
ojhfIe8dAHOMmwpecIr7+k/jjU+FBSL7qJ+OP6PNlLnZMH/vO/1gtM7uZGYDz0wcfeufYqmEj7ie
6I5S43nUO0T19ZuXqUZJ7ABeGR8IVGoqF2ZDU8+uaV90GTCV9WHh1798Ia5li0anULgvBcwH+Azm
Y92Jkx/qmY0yVvB5zj7m34Y+1Db++sAHO0ZG0F7kuHD479ubTTeqDEfu8XTN/WVnn+aNQn3cHXHy
WzhczcSDDrF1N9TvVF7eQ0x+iiGGSyIdtubI9kFMqXNZQvTqaunUbOTb1kf6qDCU2Ebx80AriKxp
XYvByKSBLM1fdAf9DdAs9sOQTVj2vEDUvWc0ZIJxuDS/+LYXy1tnwINaJUsPn3om6ond+O+13vOy
Y9crii+mr48upqFa28vbmbw4Vkn7H190ZtIU0canWiUrUIfkR1QfUWfkclTRqly+ePP2i3wE883G
RAUspA/zHEhwCcEeVg2C/Jcg0q1DtYPTcLGaEo7r7JjmSfYFGDUBKkghslOxDcDQYtYvMalpOJP4
EvezdYlEi2q4dg6mbgDs3hEMXwuqT4duppfr+TFuivdZbRq3p2c7bVewKCTeOm8DJ7Cr4UehkEC3
Q7VdbPNLCFp0OaPuFA2O/7PsGDwKuTMtrRZ8gtTrRrJ/olMTBdaJJxaZeArjNV+TOiGXQSL7A3Yy
sm0+ozBdfTmgwK7U4Gd6aHXvPlUxhwsUt1voamFfmAdA/I64BWXKul4IHtLxCzbnNwk+ActQ+Ezt
vvrLqH3uE9ZVpV5Rt1kIyRqeX1wzun/74bVepU+LuAhw2uTJSV8FK4HgdlAcqTB58fBh8UoAxMsG
Y90iR2kq1nl6ngqp1F6sL8fHlY8Vz50JV7n4qB2n0FdQG3kkNsMU2WqGln3ZvZRNWE4NEE4MOcu6
PltAurkLzHtb2xZrvc8m6ayHuMm4Kq8i6DNeGjkX0MaXeJWWrFPld3Liz3VR5X3tHgE1hRn92W8l
A+dOCb95uzk4jhpqO+3sxCxZgWDe4KVYgcvZxvp9GRhoVCg74wpucDb89McsE2jF3cD+8e3Yqcm4
VfnWMuxWz1E4J4V1i8YQj1IhmULthaniLbs7c9uJ7AGhWlGVK2IG+UA4r3lWUEvn11jEKl1Ecfwo
WEWpldi55tNbfoN+DqBAdc8jr7hvrnfjAt0xqj+LyR10peaeYncWYABCG2y/Zq/RNkHV1DIXszZY
+F7Pj48nCkA6IQam+x00EyUmXJp+1bnP2npcMEx85fNi1U0zlaaESJ2jJuzpYtRN037jO0HJsySc
v8NlA7k0NeSd6j2cJolO0Hk3euOQSTl4xAXy7EzMVCw9T0EanLhDaj5CHReElpgu6epeuGT6K9sj
X37pL7lqrWBMAFgRp6C62aadvH9eanTMtZWwcIIPx0LuQdibl64no5dRIr10Jtk0+fl6lki9X9aH
8Vr9AkJ4dX8MJanctEUr3FC/jRDWqcZaeRA2VtGQIqT852UphGWbLvDpbLklIMKRPETw63CYZjtP
01iI4IAUWs6NEtUuzQfUZnOhqtOpRFEd/dMw2WHgbdoeZ9IU/nQLZwesh7DeDXKMO/dRJ/B8zHsb
3rVmuhskg4W8Z411sIZTEMRP95oNJBaFHDbyCUXSWXD/AIeiFqDlUEpobOrinOqXeJ9po9oyMh72
Kw9fARwr9JKUFDY504pN/guojWuLU3F48h93WbUv1J7Oh2LbQV7ifAAOK91yCFJmsgpyAKVq5EtS
xC+ENg1d+TT8DDdPR1e6MuEmZvXHMgFeMeL8LMyo70IkaXaX2uv/Aee0i/CHPvTO7pwvnc6ExD9y
UmoX5YXehx+JoJfO0T5B0ODE4rOafHgUgPfPVOLwAp5xKapEECibSBDYrK1RixHy8Fzt+Ug2aMec
vEwsk+RrC5bDZcURHjctR8EshBPx/TIkchZ9QyVc4KJp+OTIZTpWLpFk9BULb6MAbgU2pX6Qf2/w
1PiAVH3x5G8bCgb4JNC7MqSXIhFW0MM+t82Q/hTvcPaHO0I0Ey5F0S27SuQjx81IsB150qk3TenQ
XPQFm64qFbttNECvuwP1F32YfziQFN9XTMtj5Oxd78MC+6/fFHPWv25xNsorZHw5hdUELlBG2Mgd
4FpUB24XE5pRVVsWLZfCGZVBjoSBkbC8N1BJD06btwi3JTwwQcB9Pnm0HGa7DBoXhMbh7pbeyWBs
cKQ7KQr1C9N17Pa/D+LGsim6NPFpQt60ZQgi6nZkDmlD32ja+v0PHwSOqPmX98iqrvC5WfaBl8DE
HkXXvLdHTpE3QhqAT+x9x8ewhbAs1l2hoY0QTpt75B4doouM9Kf98Bv+HBIHkoZcx9vw9tYBYfEt
A5ayTfHM+XkOvHIsu/CE9f8uLwzPD91Zj0dqNR0wLKCGB7QVidhw3nrWfCMQrGxhwnXltzJ9MYsj
9GoZIkHkpomyH7NJUlMTcPzuYD+7dDWMjZGzcFh/RYEtbRRvURQXSueRO4OIVpnC/QneXIscl4sj
KHcBX2hnxusZjOxYLb9z7X8XmG/xz4sZCOB/khIFWqmh7yxfRsh5WpjIfUEi8mtLyXACdjLqoQTs
FgZ2y6Dy4X3Ev01JBTcoSHcLud3Dw+44K5Cu9UxFxYJJOf/ITYf7Un7KyuhP4y0lFaG65cK0hxEy
yuk0/QvAH4TEnTZCAaaXq+07bmN1S3gttesAWsPFwUElVsxp9UOnvIQuUVHCAcinYihzHQsgm/5G
d7YCVuWe4/xl48oAVKq7sRbbjpno4x5iPvtjwmx80jsiVeqf+k+po0l9ddB7NB1aWYPrhcw2EtZG
tbZ5Hj6inoeLwzZlQUdMYrCxfXsuWe/iCNnAn9xUvfUtE7S6NRB1xo5EV6zxQs3TzWPuLu4nKVxf
sKM2Y+DDQpggXWWlDEd7T2hikMdAd0HeOAGf3F9HZXc4aAhy2pP8hebe2/gvM/E9LJ7nCOjuZIzz
VQkjN/h2CNBt4bYo1lwApllx4vaQ+ajU6JoaxdTF0e75ON6T9ghWvVAo6z2JuHnIVJmLiV4Jw3PG
rzY36zwIEwUPWYbZnqcLB8yrINGvd8t8yn+OO85EIw04MzSMsi4IQFMNDZS4pm5pMB7HLBoPW2Jx
Q1O/YokOT9Ucf8CIt/AlwcgDFU+FFosPiQvIq3pdel/cPh6CnytN3KBCHI5kWjgLfdI4nJoSuyGt
dv7+2hLbRWlD7zKLyh/YuZHnE8B6HapFt/QGJ4D9oq1TspIeRAMFpaTwiug3rXQA4X4fd6EKggK2
Nu0suhUQ41sagYrMlcW45ijOoweMSYZNKwvCQRTLPV5jM9uvaaclTBkpU7b42KEzpHW9JAWO6OXl
nuFLSdD2pVDn7d7WwWfqw1VI3G2URM7m9jOxunXADlhlh8u3RymuVUcAr9kwxaBNOdtri/bdfLrl
QyUeqiUUv2gFbB6c//iYO4IdPhq/pHUy6MWJQozTVVuT23RxtpqWs8O+6rkKHoQ5j5WsIUkwShcD
U/LdMWPC+EJfI1busGLjEi8Dg2IanXJNGCuixT9byM8kCV/4rr42C2jNvEClAxW1/EP5PFfYJSBl
r6LIIU8UlrMcelBNaCU2blnWtBZSscxb1GnDKgUQwCQqWtZEzuOYA/r0vjtSLFs6Bg1EbmSA1gof
+jsz2pIDaYYqfXscZSA0iJt8iR2nGqJlLfeJjQqqmaeDbcPT7z2C9O/YjCTjzTImjaeNuAq+nI0Q
CVuDt9/mfJW4psima9DYasN1vUAkDY0OutZa+ILAkwHIcDnKaPfSkgDRHRBrPLBT6mgzERDZIdtj
iIMNm3M5w5rr++QOcaDzwkrMsIlouROOYJ2g/LqS7yqZvmK0bngvD6p4f9foJ8wb6EL6dXenUM7j
IbfDXr2lSU1owimB2Ct0/M1KmxoyJ2LlnkhBsUn9xNP+7mdDS0sG29dgxb7MVGq5H0DXwyyK0lvn
+mRXmdH69WZJkI1g+hhGqT2bNUnlBELAsnuuX93p2rl4uYbf+mr/KLqpt0SY0CNPErbwATgtYYtY
hwBeJl/Q4QJZ55tP864MSXp5yyovQWD6FSFAnukdwAXM/VhYNCFK28U5rYZg+bFAnXaOz8/0YWvW
4BSMzktlPPmaISpn+w6/EzcXI6eTTbOQffZxvkWpa1yYtVFDQu5KyRmQa1VucRh09PYyVqXD8dUK
B+J6NxDivqAhl6nI5KO1FazAkpS1OofVeu4CvlsJlwbm6ZM2ZdFQxtJLataNuEFAiJt8D4zFGfMJ
f/eVk8W4eXowbf2ovBQ1B+Ntsyj2dqd2rQJ3zTuai1RxKTTitl6h8EtK8dBn74F5vEEKIRZrg9W3
KqUdcH/aApNK7J8+PhbPMbVL5baByl+gMqGyyOyapkdPDb7+kts8IQSkpfntFFZHYywhvQm1X+SR
7uOaOa4Ojx9dvoIO17Clao7XEk7jkyszFdK21oZW8AHpIHpU1k5x0VwKjRJm+8lq1u8tBX73O07V
ENzieAb2K07MDWTH90EkTiDn/VLz4d20DsEKMx0Tv96zeZgusEkkpqUILdfcjBybd+xqClSWk+M/
N9PXHp2ZdYV51CjLqX9u6XZKOoAMBf+te25mb47W4bPfr9Z6RsNZl7nRBW7HY6qDaKX0F/lSpOor
/Va+Daiuk14O33s5dhLWz1940c0tRCxGJcT+/1bCC2TJT54S7wXiwof4DayhjmRFhAOsfhGuECAR
eQsQVxE/R1U9k/ieuaqlqx6K4OKpKQDHYzA2SlgKiFNL+W3+/9EQRTYR80bo6oLd5sJFgjPYylsu
p07vtLUAARevjSwy0NknDOdklkilG3aebAvuYu2+F239Dn3sS1nCQa+tz4UWIjvTTCVO8a9DrwW5
iHxerdxF2JO9vYTBVcUxQ6cunXx9wA1N4wIPgolbRsrovbY5AcDsk9fFdnORJccpUivXzuqCwZRz
0kUTRhGZtYiTWiCLPcaMgqMr6RMquU4ERDIxv7uiWC2KwiQjwyicf0pFIYuHfGVasIyzAQpEzClm
7rG0XuyjAPcmPX8U7MZNi8C/PgTtPbVVkrsbyt3UuOBbCpgQzJvPiu/8A62rUJ/HFprTK/CUyxvR
G5516wzpc2ByVWkMkMKLOmSrlnmBD54VSLrU+0Qhg8Z4ytSapFVtB0E/35T3ysy2QPzDm/IRjxjS
nZfC3AqCfmVMGQZj9bQARgWyj3RuszMb90EJApwI50QgbsmLtxx4q5sKrb+2f2T8VlGe9xRjgQWG
93EalKWZ8GjYQz92PZHkhvDwEfcakxd/FYHnn92Ic02+i6DHC6kF1/U1QD1UrhtOEgAsSUi4+DYp
rr10j1DUHry8iZZIeaHffYloa6IiJjtPPkHFkU2paCzBYC3TAB9tFiiRSko69Mq9z+OEtLOEtPMp
vUTi0dukv1jwLQEgHw4FidrDj8eMDe8lHUHVlge9oc4H56+1dIuSNE27k/vZbO0hH3bzjouVn09r
r7x0k8tn5ggsTd21IBMyMI/6RVPZdxOEuuwa3oat5p8520zwIlzCG5zG8xi4FKGhpkLooktCjavu
KhBtDS5z4/oQk+0BZHuXDPJTHVpLsFIbuIJfuo3XZBWR2gPexdKppSagDTw+ru4To2Yw8PQFutZ8
DfNhMj64265i+Mo8KxuvBEEyN4FPFkv+qzFAS7waH8AQJ2dMpQHtGwX5n4e92Rht+gSc8BAeoSUK
VY222ofv//XUg1bBY6cTjwwmVkfMfbMW3CJpwHDTs3EDooPCMgwZKn6ZcUEFpKUXO0WI8iP1Tpj/
kxq7RA13EBsju0Hlpc18CgozcEazrlOx01ip91b/FcKsBkJ2ogAk7fX55brMGjBcItSV8xiWsnit
Its2QRk4PTYcsBiIKlHlkpRykuwS6r2Vl2LNt28StbpSB2+4g11dFLaxyg28WIimH8PePr48CiDe
HREKvgViOiVa6L2ynjoqj2mBAwdmzlCF2123gpXpNZ3vZOXQTaHUXxayEoS8QdrpEusnsye8H37Y
Cofw174LyrnTjvzLhKZQt5Uxd0N4slKyqYPAC9sVL3PvaMHyICCgLdBkP3myCvx9gdvvyeaDHVI5
BQ8NlMd6EW979A4UkBCi15aQKm9gBBZiUnughLt8z17xoY71LXP8BU00o1O0dNp6BOz9Wo3VLh4+
tM6wp9XajR6vWvOkbySPZNPHOVHSqgbpu5UBGF/wMm4ekhtsOQlYxX4FkBvwsmb5FOc2889xuEEY
GABbqyschLmAaIMyNVFB5eguuY8UUN4JjKO9LfPlvsDMeMbzpCCkEm56mTziOPAj+slRYS3jnXcp
+IxzV5lhqvGQBBXA4gi4Vs9ov4ZFuQXGSn2TvyH/xY+kcxnQ45ni/kLLS6aWza2WocG6x2WHN/6M
uG3TQKRUw+8lG+zTlmRNwJaHVC5HALc9JPhe/lpJ3mZ4UOhnCZ7/5+uhIXGGURujEmOZFdmPwBgP
BqbAMpshCdwb+J4ug4XjkwoJbxaVcJ4+mjo8An3NCoKwZ2tPTz5NRr3Knhn3/lXOMsSqhynQw0mp
9ar3TsdBIPPqBhqLeXhFtlmiCzyNuSOEnEEF29+iRZrKL7G3XTUd4+UMjcF62QtQJTGq1JekHdty
/WfcXw1jbvnUT+oezves6QxFc1svNjWZlx7AQNius+zsZ2CarmE/AOCEutsA2zLflEzp4PXkmY2s
/qfx6TKUyzUFH54LpHOMf10F8Mt2YJ1rfzImsVLxL/CJvOzoa4VVjclfyxyN4XgNzzJECOTdP1WT
QxgSNqZOqWxVguRjsjLhApDCbCrKlqbFndxxIlLlhEvyXm6QQpadlTS/GB2klpoUZtsYDLpiT2sE
vE4DJlXOYbU7UV05BsSM+jBJjOxwrIAl4jp1Usl2t8wrS4No/mQ2jB8DPpyRe77C8rqOwigpVOvj
3PZcJPmoYURCA51PgHY5s89GlBaa9CZrseTpq2Zna7w4J8dgvQBGHwqLEv4LaTwVzFeMi9Kj74td
lyCjBx0lB58PpIbheKlMU4c6ai2TPoe/aDvDp59rnwmRNCmeuYYBQr35aayr6rpASa+VzsRtYMJd
P2YjIuKtY9kTh5HhPLIweYMvgBgsXaGE5IsPStdCPY6wEVNeeQpgcXryCTIZjrksRa6yPrbwfLVW
ZBnkndrCVEI2R8vwWxqxnteOra5JFT6WCpeidWvrUufhD00kku0lFukAdrMEgYvH9HJQyI1z+RQ+
BlwUfsi2DDUOtH7+rI4UTjOWh+sfs0GCa52aPY+r4Abq/ge4YiDVUwKr85WM24mNAD8zxCZukccd
SlcFXAq8OQkrSr7ICXSZttjia+f61nOGziUsqFoRVmZtnNAT/GF4w9Q6b9iFIH8RyxfnDhrub1DG
yXjQFOoop29HQ/krixgiz+ORMLfDGEfPv8eUMhK76Q+xWSMrl1Vt2U7PBxjVSx7yAZsIl6eRvtJy
bzELWxQutT5rL/4vHhvElrHldjX78pEhTRL8NpdC6h3AqK08U19SBmq9aL8W3MXKkeydDKhsIdTu
SWF2adFb14JcLz6rCPmfd6WR777m1YzwofU9JiaTWIa8HLKVAg0W8PUcSoqoosordepvnejx/+Qv
+HWX53sWarzTPHgII9oS9ujhhNECB7+rOdtKqfm18BL55BzsXbz3YThMfSTpgs/RA5kpp67EdVRR
VId5qntSBRDE+io23yQsWEfCSXIq5/OqQOTgOdAZa1tt3+kfQPKF7wDh9djrNOmt3CEFIvfuy2B+
FPOYQuaQasFCH1yG2tjqXfP/eQiJK2f/fbPUND3IUVGVtMajTD+1ocE/9DaqVAPK8+6wxdK9AOez
aymkRFedGQ6yoKsmu8sMyNfwBbaVSnQbES9gsVDIQyi7oU8PLrYsdH11MHvcd6/qH8m8BWPjxzJU
XsVjtM5XA6Uh8DnhAWDVK387UNGVtcwbFIw6eRWV6uS5ebDcDN/uL1A2XZQVPb+EICr3aZ4/Kp1Q
f1RmcvDo3BBQAvqjC9i9GKJJ2/ZwpGuyUBI9DMDO05bW50YxZFN4cSMqCSK6/gdRdIyzsw6cE8CW
4XJwqpleKsoB9zHkQ8MYNBeTA/FPVNL9yJHSjnrHGUFYnBAO1adey8XbtSffm4Gl0WCl9UULHVyW
5NHDNSlDEnSfgLxprfQ1dm/5AJY6jECJj6ysRsxFXcrQTK8gQ/Pi2bL+ZolEw0lErkWfV9Xvzbhl
L1yG95vd7g0a5KRv4yh67gtJPk2BajShtpyU0uzSOrvvgI+w6WA6JZh1Ijdy/JBFALq1ky0io4xV
a3Inh1XvM7VEyxh0ruQwQspf+LBmGE8Q7fUsgOZklrg7ISMfz4tXgPgFEUT+G+dSFQ3oG+0PMzcM
Q1zkrG6UtKTP7POERFMTg5cLpU5mEbh6i1S4PC0aUlpqxqSGTT3GykSbmUVZEynCu5RE5T0bmTE/
EO36YWKLiPFERIuJZh8/vW4HME47vfgViwTVREmd9V+qBmYojPE10yzm0wUY+zH/7nY7rFIBNyGd
E8p1fVZX5r0TAFNjkCR92SOSRZIcLB8iE15abbl1C7v8DNcNlAo7ZsZ74rOYgMh56OoLRvThQtsG
O4XhPpQeDgept0IsR6bdwsr+sflaAH6anpiemh3g+ix5eFZA+GVXolb3Oov04z+OGg48XhHrF9Ha
7kyi5jXlpL9Io8CxOIR4YU5NAiKBHWzVMjPcg+4VXaE1U1CDfTMgNDPHnp+mqDavWF5VABlnS0q9
ugsCjxam04AYXvrbDJDhxs87HyLCpLeSUBDTzoqeUukOEc5Hpn1mCzHCHPrDm9u1O32H4ntkOAZo
h9VjvyCztFdmtsKI+HONP1lgWgPqS/KIa0oDMdTnw5Tu9B7VcSFpQDrdgNfi+xPBNE3O2EsbBTxS
SPlIlERpvXN7FaVwCEd1+sHjjQpfSrSZjE4sGJQA0NSn4aMRL/slriav8e+xFHKChA2LxMWwiYl2
nzkQEtxuCc2lIFyhTG+jO/Uc4fsZZR0yJ347AwDZx7mQmLT6OPeKMaXOpRvFwiNcwR/mPbZK/LxS
qtEb/MuOUppikXtcjj2ugpdC4LoEEOoDddXpKMyD6H03y1VgPQDQBFO1/1EoDYPJQEXUttEXYZ+l
TMutgO5R+tWm09lTCiD1leBVPq5BwnwMsjUjFb+HdmcVW6Hfh4Wwqzt2WSDgYaT7SZPehGSxQj7v
BF/P1cRbufBIHN2RxCKdT1MacySEP+fDDvGXnQ6SgzX+Fp3v5pSxYULz95QMa6+c0TH1fpqlISiG
UtHVW29DpM3mqvg0pe5JJv4hmmLbqXR2+YI89yxHoe7ecli334HX7YCaH3HWmPycbvTx0ivNtedb
foxaBGAWKgFwIJ0yHPqDd6DpGZPXEmmER4xYVLRQ9pIui0Oh5StRgmW95imzXqDb31tDDFZ+SRMn
yAqeDvDs2yXFXzX11zvxrSeO9feYIVbwLJgIpKnIyMqF7gdBcYY7QyP2uJlAXe2BWfb3CNdFwuGk
fUyNUdCV/fsroRZEj6NZn2I2yAcBKxD90/RmyzxTxngqtWpcRoHDt+kUtAFPmawEL3VtCXXy5Gan
NDnZbd6kvkMtb9F6JOq6obP/F5/A9Ori3AonjaULVHrZJTSarK2DNJuF9fDCmclC/7ri0vkFWTrS
axr8W6vdFZfh0yLgghLsdBTTyKL0l70oFhglosvsnacvGRBIcEsZGeq6G7TEZBpsLaGXEP4FAM8v
hZD+cVYConturkl5Dl6tgj6RgYK0A7OjHKLnbtlKqNCSP1JRexCNSGwaWHczD/Uxp6zsCW4LT1oG
fEcKWEZY93b2UNrmiQQBd9k8PsTTNCZp8/aoUTXIjhvqKWC6xEwH3/33DDvj9EOeuhzNFFUQIivC
08n2YEWwXdM+qjtZFHUatyiSAkg5P3ST3c4yeEn0GbjUvAmgIpy/WfsVqDjSqRhCyRI2/T2jrs3I
EnFJGuijmikvXrEx/fmRPQxoCzGf7H/+3BwHjvMTlO3f/iq4GoA+EXSUCTFaHDRATH9NgrDFwNM3
QFj8NaIZMkRjllSGnnC6bxM47JI820yjq9ERgR/6cu1KNZYz1j//STqKveY3xkbRY0nAXocI8C5H
dF1IuP+VzHOiGworhHzyjGXMzpUj5i5ag7+1Tw9iFze7Y+O+OG6iZJsLYluUtFqENs0PH0yfc3YV
L4ThML/QQbc60/pA8q58FtTvfWcTuxLSTXy+IpcgkjY1M84kfi8X1hIoIZd4rkoLWiwo5T56YDcV
PY+s0ZXFnth7zOyrTZmT+ZerPnBOhJac83UbLGqYIYtMlD+J2GZe2jcua/T4FhQg3L4ISgpPYXhw
cEoNhSdfkZaDAGevl2/QanDutNdCLzmrugxQiN+DY4mu4U5D1QKDzzTR//laYH4tqMVcdIrgqx77
ns8+qFSBAq6qqTUr/i7aC2j4HDsYOMfklAf5FL7lCQneHpwSjNwZ5h+NyXiCvZrySB6d7JmK2Yqb
IH0jpDJF2zwy7AbQScoclfPNeoUkmbAXAxSpa5MM+VH6KUTUm6oKM0OgEFYWTaKKcDOXxf0gZZPM
c2SpIEW3C5vg5mRK4rcWArbWtaN5I+SDssbNz4SnTepXMZi7cXzbkeKRCo400T6G8p4COAXfzI+l
cnmA9yV3CAXJ3BJsvhsRAlDwhvxRPSpQqb+8w+fxp+JrWPYnN9RXGmLcQzOSsFfBpVVKPseFY6mv
KX3aOGUpdpZXo/1WtEWxzzH4GktrntHSC7EJfyYcOmFSS6FIuUue3GfO+xUEhHxvEnCUL0ITdBZj
mwz40ywqtU0454l4hKdonCwwlzXGem8qEFiMdiu/vYyn9cyN7101Cf76tupgQrbWTqqGFWEusawq
EqdIYuBHr39v+knGMuGpqSelqyYhyCAlylP2TG5iWp5OiDEil2OV5xCx2kfgwMx7+j47RQnPo1VL
KR5xgXYYRTmCIsuFZb0mRADXUJR0e0p1b5TdKacGr8KnPyQWX+BYY2K9eEFkk9IzmHwF8HN1msR2
LPxhufam/Vmu1E/Rbeia76PNqWAV8vO9heKvodnG/pXVOR8Ph8h9VOQq/R2UNh6Ft2emvcUl9vGh
47lhjlBqMDl3aGZjFGn0NXbPjMbcPwBUcRkuJ98VbgChtbdl7CbBKzBOAXYRvd47QOnLPRonVu1X
BBg8rLf+rH9Ru3Wg0t6A2H/U61B9lg/oV04NCvnEgNjG268UMw/sBSTBGh/lH/Zo5LoFd4QIY6xs
9/ueoPL4ESnLY7mlhIDyRNdrw8jztbDKHbHvWq+7CBHHDsHHeKDY/YFFEVicgmadMRPT3hcSll4L
acwx+UtjJirZT6O/0GlnR2gfHW74U3g5qkV1fyza2PJUlanUqR3YnBqGR8n8pvQLdSb0QC9C/PMw
lgBkNyqmSfSMRCYSU0fRjc3OgpCqvTgNFkPvzI0fzWSwBqMQ3D9XXqGPzhgtrziW5ZJ57PLAVVU9
x9kJ37q8pln7rlfJZIoU2DREHzaltduM8P2I8hB5fur9SueuHTRZQJCG3LHVA4S+BZC6yQjvJtk7
YRZEEAqVbzPqoTBcaoq1FnF1RP0jExJ4Ldgd3h4s+uuwUzzw/gvDZmNfrrb2/iYxVpTkVGwlXdzo
nGE7xaoBXQxt3mVmDqj+YOmOYZU6601IqcWMv/UOT5FT3Xifk41ncHXXIwyRV4EjbwEXq/BWfHXE
DYhcxhsXMBrxdO8l1mR3rXtqz/A1mlV1JHhBR9WmUn7i9gKaFce+Eog+xkQjPCNJPc90wBn3YOPO
sh1RLVYO0Nje9Yjj6ve3539I6xcd6QR+j7TgI1DWjt7tOaSHaWbMrXkJK1icCD6F0euwf/YRjuGM
KFQkm/xz1CTvbtq+fipTqgRr6wP8VydjdII3ha7AWyiNhy0cGbM/GGg4PAjdokL5uoJ8zWR9KFRz
YObDseTNpHs3SPhiZ3b7HDS1K/OemuI2yE2FKhdQqeP8pWalkIQNE9ZPuM4N9b1pALOmUtWcq8Tl
4rf72/1iNMbg+jWYMqzhG/c/2+R8dCmZTNFQ3wNs/9JRxooE3zFVP6ptdQEgQqWiDAEAxHVFfyPe
xNF+SSXtNsWaGq5dhfmvXD3MkOavCJpZa3zU3U2Fd1niYVjevYJqYPtgGUktJlsUu+N2RstWEY8V
DLix9Q/yFqry3g8S0YUNQl0NkAiUENmnz5tI6o9ubiFq6S+7spmO9/+kYZgQrOybviJMkjhzXy5c
ZGixcg5beaUWOOO8Dyo861n0ZOJiJjdY0kQfuSxN/j0Xk7RTAwvhU7wGWiVWG4QGTHzS1W50XzvP
suEcdU6lTulPFqTUGBZhOIjWhx3wh/gaIqfHvCSqrCVddNi31tQlaAf0DNFZs6t7ymkpVVFqmYVN
8wQHbnab2zodY5RvxfI+k80kM7JfrTGXpLYZahFSU1YHVDmqvpM2lUmhWNoZJn6tXqIrlpeQvmdY
OosO+vK3TC0Hlh6qEkrMB04Bl8D5h2uItVh+908UIIr/DivxdxtOEL66Mh64iui2godR5BAELI80
C05diTHKeJJ+Mq1WOooq8xjyf02iQhMUKxQV9megA97JskchHJdY/muXkHhpIVvsLSrygu3qB2w1
4CXmO573KAratXl1nEY2srWCnWKziT2dKQeTMrUkEby4VU4AhfW78FVSh4I4q/+CiaJChC40pbFl
YMXAgqTgQHiXkCymER824PunQjw6qZxfkKocozSFg/kpCArpgqZ1RA46EEjkNXExr3cYdJad6Xhc
PZXzu9D7wAVZOG31PFGI9jIHoa4mVa/nBobT6SysXcNJSEGvBhm4zgJfoawKk1BDj/cHljuruui3
w/VTL3cZcO7q+lmTCejIHYFDzYwgn5HL0o6ZZ7pUL8EWSK025Kski5PExkGQkSX76NIBu6Jt9D/k
EmwrAQ4/kaPNZs8DW3AwUU3ukY124eHQF0vP1wn3jtpdkmQFhZZ5ePcQpRkKZqiaATKx+Z0IzfeM
oY859frvNf60eTg1xuepyhxL6VOPOMn/asnhSbU/U13vKHqyV499uD7M/AwPE7aBtvctkRY9gBNh
9Pt4QkJQtInpmxOajGBFwx1vWjcZXAPuZDCc1vraP9dQJOX8fEIYtW8YM1BDF9NHwF0dgAvKFx6c
wTT9AKip3aFzSqzuWFvmWIFPMVpzz3nepHkgbjFQk/E5UdXMRC156oCcWkgB51oByUtICSblJO+D
XuDpUFvdtIABZ1z9AkS/3rqU5nyuHc/aRSqjVjzb+dHrwPEJdLD9OjArmm7ABf1EItYZDlGCyEyN
zllhbIR/qoy6KMDXPauu56bqs853bEEhs0p/OnLfVKG/E88doUW3m5LmgQaSlzJ+A17OkjoEvy+7
bflIt90lW5tPWFmeKI0H5YyeAGQq5hjv1TbMNLikeMiI8sP8hpXr0oIPLOam94mLDzG89GrLVHGk
OR2lXUbOLPwvPVXlM1ewNQEE++RMhJFblq3dekyiaqlGT1oYKJEzlVNkaybUsF3K3fCqBrqDqFbX
n+eu4mxvOlpusc5YzN3MRu+/e7kJK7Vyxxile0PxpxNVmZoDPHcoD7gxJtKWk21vXnIhYZiAAUkL
evA8zZ9LpyZeOZ4FJ8AL1YmZFLak00Z5X0WUW2WFf7fN5mxponMN4KXLpMOFNzSGUtlcY9PrscyW
/ViCpTTdRymcciREee4VjVjdxRenPLWji9dKqf4VQ4jy/2tmYYxhYeQSbMnS53YivHgClk5/tAjV
UUJ+Em/+myYUK32wtNO0LEDAbMOrpLz6ZVTSKsO5Bcd22DHHCPX3IoLAdcx3EfvEQBy2Cw4DA+0V
zFBUiMBIOKpvOGo+tNljPjoBjT5Nh646S/5yiW9toUa8i0IUbk5tDqxxEp3mHRBBHzbjbs4twDK7
73JJMdI9l9WfsIcxsDphPZ1CIahHoCiqW7w3qoN6KP2OgfrHnOfX8KDxTnBNmdcRuVpnRU+sQpJz
DfynIuB+8WCflJOtLIFoI+k4tsiHMOSukcqWgwpi6AbDhhSqN3oyO/E/eBW+JdFJZ3pJhmCPxXs7
zKJxKgR3EjHa+YffoPP5vwnUcYOQ0OcwdhDwC5VF49gA6bnxGHzlUbFq2As5DrcqC6J/tdNX3gO1
mrJcR9hLghlIB9kMiK0RvtyANKKbeDqogYc1+rtwKe5u9GJcdGIhhiG5jv3XEW7KlGZS6kocwkD7
9PDb3wfTQd45pOAN9tQ+4e5jxAb2RDTx9+K+t1V1n1FPzOA7Jown/xLRoztKdia34Y/PYziQ5gsD
568xvnuJ7nFvh+8E61U17NO2eY6Fyo1Tlu4VtrMp4iRGRwBWb9LZ7Tt7G2DidIXPF6mdOC9lXnSK
Am0QGhuSTuz1P+zX1mO7RclLE7Sm45kNN50s9w23tbfIb4Y6Vs/+kdF2xDWcM9fQMQXpygvDTEkH
XmiHNFwnV7lCYHdRt4TShpxiMHbmaZbygk5HiJVhmSO4Nuso+1h+NHo3TLPk/hWPR4rCzrBOrcRQ
6fBs/Gnclhu9+EDvSI5F8edSVjeckrhycMAzCOgsNWhuttFnpn4CZQs+ttWExkJDG0Zq6T6hRAOD
lZoFZnu+EYBcVQhENRi2FwWU+yYRDFDhiv4eBqdksIVdKIWkegvY8eFXwchxLDpwdEIkcPmxtGeY
PyIrtjGuyG1/GInOMc0Q8OtSW9obySNuPFCPBWwNzOGedIufeHqQmpYF8J+j22YbDcDXRU11CoNN
rMfGsaVBIao61txuR7BDIi1e0wEAhiKhLDeqPoU7vsIp7yvv2yULhWmLHYfBvc3Yi22Ql/P+Ma6N
rF17dlzMnC1XROk7I2V5yUDm01Zqk6M+3G3l8RCEiPfAk8LN2G4vxXzJFa4BiscQwEpoPpNHx6Wi
R4R3D3Zz307z73NEaRI/2reRUQvW70OXAL3/nU4k0HPBB4wsWMpY81dfqb6D5XCYHrCO+kUg5uKx
09vhjhp3M+ZwLHV9csg2QlEUgCL9q+fHeOk6grNcdfquoHzP+zKhMsll+NRLIO3aOhuw0jjPkfAK
ZPWV/pcP3PPbm77CClLVk/bErEMJBR5DLqaCz9GDKEiJnA++RzLqmwMFA4cpS4h6j/za+rW1ZOWi
Ls0yPAzEYr5khBRGnImHjtByKKasFkC+Y7tFk+qtcC4zIfvcLudZeNrSAN91R6aRxraltK1YUAlc
gt9fpnGkfyZ+m0SKCteG7FdgTuOM++TRBOh9IL8t6CpXAi3GmEB5XR6B2/Insuzg4/MHGM56sKIU
TSqFI/4kipbEvoQXwHjBKv9w6WeFgZonmoATsgJD7Y8IMFzt5kxWk7/qeOepnQ4Owe9abdAb/1Nj
yfvhS2iW4hYTpC7zVWcxZrbPYOl8CUjNHDOaYyetKdsYMKqbimGeMt9KD/g1RYsjY5GcJItDThDJ
iPvFKJ42jI0AoiLx9rB3BN08W8GT9gUjO1d3CZq2GfCdakeKLvEYSavcQbLHU2bliz6PIBpPa+1+
umwG0Tl2kX9+aoTODiyG6qqIxkknkL9lHPiRLMaCYKdVOkgK7jak6JacdcVxRuelxywwv26WtO6C
Kuf6LAH8vtXRd15Bff+IR8slwPT7YkYtjhXMmaMxMYxo/7enTehuhzXefJuY2x3fCmh7ivIH+stK
H7jDuddQ439rn2KvP2J3WyFW2NZgaGCsHVW0mklL9G+VTXCNleg+9mriKY8GyJj28ytEg2uz4YYZ
CzEuTFHpSHqdHAUxK82HkoBxBLXicOhUXfQaK/rYRg7pbuxO4XQUyfFkeortfuZ0KYPbmg0e4AF4
nyxNnPDhsHpk7BldRBBrpW3p+4b8V0aUgPDNtOsgorDQedJDuo7rCw0pxf+QL2cHROja2vc5iCdh
mn7Yklxx8RMp/sTGdDslAO5cXZmayAPh1pQdq/X/XQge3hNo5Frfr8XdYDAVaSy/ReqBAn2I85gk
rzxoumMwuVowvmbF39cFeAxF+ke+w8+WHm+XBOkgDjwtKVJbrohLzOmkBZl2vHYilBwLmCFAqw/t
vvcExNLgU6Y5INjQsBvfOenLtyhixYlMCrvS2D5DNNLZOY2qtQlPQLwc4947IUy9OYc+SgWePXuu
/437ZZkuzPY4cUkwWnWvKBeih4+z+0y525mF2yp0/gC519W1Ye42hSBAS/SMWNChpHXC3XM17mXj
Sa0bSCK+jP5KJHUgfJzi3aM/vkhCVpQH0agYBbyOxRAVHHmz6BR4MDaq2mM+Po7oGT6+KsJLBIS0
OkUA/JGB4WaVJuEMxZOp8MYh95kMnA7rrRfSpItrBmiVMC/vcqVorDXGwfNiZAGIWiwJBRBXHf3t
zR7v6x4sp1St358o0ndt+QL/UsPcgct1YCoNGqwZqZay0Q/LlVjOk9WH2HvD9L6RtyDGDhxOwggY
Tqi0XMm1YXQ6XCu+k//3TfozVlB2EczNEDIZnTaQcp7yPNaye3qZX+26pfPEHxCtfEJBi5lraAII
ow9EO7kdgR2mCSPJfwRKEuiM7A8W4YB//9C6M+mEycOFlHITCmp1N5CiAYE+utROR7Bs8onkyrUe
iaEpyCMf5aDBLkZJhavS3P+ywMiGYGWsaRMVTKgO6Ja5XMkwsFIxd2F+PCanvoMrJhlQsN7aT6KL
Dwv4nbSI2Bu8t4Zy8M2fIaiCeXlGTcmeWWBNo66ZpXTPLyivGTp/fWtJc6w6x3QfFXa3HOJJ4npW
qlweh/NfCz5wCpGNzwifEl6AMDX350CxS9FMztMvsy61cMM4Qt3Fdz1vFlVO2/V/p+c482AqofzV
PODeOzLrZFnOTLmLKARfqOQ75NJxN21r2gVlD0CSw8qX2jI3/jMER/F98nCWE5hMxXIB8J4i7orW
g2Q8i4CGdt2+yQ65N7NlLbaLP7T4KKnVNaBEvNk/ggYngQgkgCu2nqAXF6PjvYvIsYiefccAuz/o
L5uz5ZLvWcw/AcivZCgwVBI8XxqrONy0xG7dgmdVGXlsqUmJLltdSbA+cJFjHDjcIqYmdGb2CZ3w
+zWLp+puUrPwHg4I5qwJVWfMMcctOyl/qpT1AbuRrCr1y3j6qH7VDDzHJKuIC1wfxrK5d+8Ti8X/
6s9zJGHsMnjP9NchU/wEJAa5/JGzs+MU3/7WOTYhQ9XX/2yGW6ZhCP4YNErKEkvZ4uvz2vjXaQbf
cWEtPQAOzuUyr6rwopO2Qwenfel1T5VyIQ0dJrk3OPIH91IBlHUKReNYLYxZI2F5fBl+AkbNvDJf
9fcdKvfMzNVq2c73X0v/oavCNJcs5tL7c1ajSRVhvg76zAx8bBLfID2SZOrLXVHYT1toQJt40aI6
+pgqP5yVRHU8yKG1Uuxirpl6exqbzxA2wn3uCb5fRyqUxJxycflJumRNbdTxEEnWkSKOlKSli5ma
1vh/7m79lAi0VmiGwJyIkR8K4nV2mAO4oUfQQThPMdtxRmP7x6cC3KvLgSxCXgfHwyGs8NgmXu6d
cj1/dpj0XzLo7bBBE2a+m0opRqImyrK4JBQQiPjUyv4K5Ir9mRZA0wD9qQYSyzBhsRbFbL0HVPfJ
lu8uUudCNO2JGkllHeSYBMnVuvTVDszWbkkpBXMxzHdzsMKicNld6/csBc1G9cujUlmTndCDfdVk
BjEdfRse5NHQOVp0/BUlTzCvnZye109jHFew0KIfl37LSqmfqB8x1oRfnc1E5W9oiEH0LEzeEP/d
gPa7iDyxyweK2WXWuqqk+fDyj78D8xMYVyXgCYW672Lk9BKMt6X7OTdj8eJ3ygL8N1Uxw37SY1ns
vMBi3LJaY2/E8McrTgmyRAQbcdROH7Y+zwW4LnILx5yPVB/pUJl0hj3RsgIVJjH1V+YHsoz22Mjr
IRy9OH1f1hgMKL9kexsTJk3J8upHOjrUeMRhHzb/6JTqdM7PiIpx0ZTSHDiUdWT4IaYlSoZTxV2r
6BopCbmsUKZkcWodPQiHpaOIKq3+XTRAizc7hOv9SuWHi5CHvDo+3ZVPRgAxDAaLf/ZmfksbiBD1
JuqwAwBcTz7O4s9sx4NJyZ/ND4FGGtd1gBQirvyhi/d/XpWvD+Vccew/61Jc59MKGSrhUc3rHAF0
/1OyApt2oRjEaehFCUGZ27RAMSeEtQk4wJbThCeTZscELXnibZrhuwOy11BflU1gQZbjPz8fZ6qn
b13UuYOn2CDmtX9ZRu+cRa1eRC0yTbYdnNhpSsj6JDCSJHgHlXivnLXmj7ei8G5wMgL8Ot56THx8
y/5NcgpgYut1PGvEGaBZoxlTTFDg0n7lpe0T37t6K1+cTRdaow0N+z77jzeG7X1NF1bVr0u9Wa1d
pxROOByQw8xapxNqweMAVclSgtDaCQ5IJtpNQaQUncxwRQ9xMiD7oBjr+ii6CnPmoqyVsTChVskB
1rQpi2e5myZwkrFuZRycB23ZaGtEm8MwK/89EdevBNaYgfbIoCPMXB3WmWCqBRXGGgNa8MeQ7uyk
uGsoVh4Ply/76dUeHSQxzFn58SOzdL/2hslrQ+DioZVIlhSh8oqv1Y0xsNVadDljgpLGzWiIcB2y
+z475LQ9IfEXZyeJ0UaprRgFXqs71811hJK+g+eOcEJeqcyaLfdcQWCIofPwQKfAmQ5T9InwEsK9
h58is4FBpMaGv+uJMH+s7zUE0j972yPBs5vOCF6MfApp4BpNMyG0mjOoUdueaqu5tmaL/Aes72zT
umqMa8zPek7ZCYL0mPBo2X0/PZ/2pma3/AvqsLM5wcUOE6cLmJoZm9eSDT6f/oY7uN5Oj3QLJ0w3
mSb61/i3ga4IxGkC9zbUQbIUt4UD4l1wPvMy785oNLIEudPL6cJPXgWaOXePPWVeU47M7/oIskRV
VIu5RU2meZDNy8KuYp2tp+la9Urkg47mAzr40gBZ9++2FFaRJgO+2JhbCkU/LSd57LV6C0GqS+f4
F0dMQMJ8rkh/akXYc68vYPmz4sI0fexwH3nR+HF2EycBEXRvj9gDD8XqTTDDKFsz3++qU83RSOYZ
pO0yvkN6FoOa2l6N8on+xBXeuPFXxiY5Qkpy2zFXXRUjCB/aU8a2YUe38GNxv9BJ/ZpfLGDMlYiU
g1jmAqHC0/huQ7ewpoDd53EiNMH6UU8Vi036/armU42x3EmkfhlhSHRN7wDM9xUlkibsm9s2PoOp
b8zQIR5xMNkvzdh1CSBlFLhm+snf5YFYPn9rowCLYxgIp9AnkQCDlrYjaNAvzByIYL2hzfXRe08n
NyQJ4wqkVCZewK9m/MhznWrihbczOAM98Paoasf+YTLU9LqUUo/rJEbbjGNenfspg4SRYsfkFy8R
3g7SffdMJtdu/yL2UjCNBFEvB+6cvWh89i95FkjbSR8tKdy9yPdjSqb/3iz2YMnDV3AjkOCucGzy
6UE8x3npWRgS3kGmYw5BUBpyXxbS17daKg4nSFMq0Lxdrz1wcwkCUP7W2Ie6D9P1SeO7YiCUoY0B
9UjQAkzgGDkIhcjcXlrV1dnZlWc0yuSAJHaQVhNejKqyxHVyw1LN16eEbcOYfHHlgV8OSurpXmFb
e7Zfb5mv837gy8sVY4zdrlakHnVPXVh7FHSjlkHwbq4dn4D5jjNUKKSEjn8umJrvrpu/0t3qLqFR
egJ5iWDYiE0aIGCilGB7W03pdCQtZ+ClMx66HKhACrBUHfQaT2Xjz9xrgxxa80vvtjWGRkkrryz6
PM2K4RBFL9V1q5/6d5HPDcBMkESkS7xa/jFhTbl5kKcGvPw+4bnZGvZmvRsSBp+TJrTl/ah7wAXL
jGApmA4CFynOM0IfiTyrqDZE/9WRgM21JV1pVzX+RHTaVgEF2xYrrKUmPQr4nGvxOL5a6HjaIcnx
TgXNLocYgzPzLgvcF5BIfSIwDEEyHCIAEcDh/94NNZJ60aOrfchT6WdBGnd6g55OVE3lGiueMQOh
KR40YpHZMaKIoi/wbMx/uepqbyFhEFHPevQ8DPEO+0S0Dlux6zLZLzI1Fa2ngPalENIiZ6jvxDZM
AYXjTwJpCoUrsT7wgDsg2kvNKcG5VXfQZmjEU8m0M3p/DeUa6IlPbfwpUhyMTc32B7zs+UjgbK3E
gVw2fD177NBeFm+REMHBZfGCkAYDmvdtMG+SQY0Ggh+/T/Wuf2jiO/crl0qXDpKIw/MB7FHPN8Ez
D496BPFH95BrcP/gysMS3s+K6hi4LFYPcpX6iCYpn4ea3EpJiMiOoMEYwtZGljWa/tIFnGxzJIgg
tRCz60AEndGPChJcQaxNWFEw3igCvb3WLzpdyDOlIRYj9A8SvLStjax/+5NzRAzNMYphBU4sbTfy
0lWaPZ+9fj2FE63t+VKBKnqjPdcfeg7m6ESa3Uk53i9oFlzp9VBWczsJVfOzN5jEBXbbi2Dr3MD+
n+RqEdxPymlYGAcYcZn2TXutNETxdNAM1oMXLYI/H+ZSHddeepgOjUW4SKlhHLZi0QEa4sXVPJxw
wUBb7k46qQJExkRCmdkLmGGaephLV3Mce6aMFkEuzPl7J8RgdiUaJcm5HuNhYIES2vALJag3aAt9
H5C8mDYyLYBJIT/Tw8JNbxqIG0L0Bhr17/ppQ1Y6IufrxkI6DKfDkFdEpi8IKYSHQnMxVdm8Apim
8Er1nZ6wiN6dL/AsIyp151PUpHI/vkDTXZrcdPth36xzmYBz149SjT5SEN1v8I0uaH7HRQtfEXXg
V1V9zX8/VvrwdkLqOYX3ceQCHke/MTsJamRlZgHr2mJIoCvFoO01o/1j8REUKG1tgiVbZWO5dt6u
iBmhQkrhfDScxUj/mM2x1Daiwphi1+PzVB9/3AhzqUPDNTSdntvDTzT5T29F9Tw/YjViKSNzHiOQ
CQ0Pq5bFVH402deox7VFIYFS4KU83RtNFGS071jlwary5wiDGwnYfOh7S6CNS4oUfVobhsTVmLWF
gIWyg/foBUU0m/GINNXnO3WVB+rJzDlNdYcLmNZYFrTo+TpNC7eudeOueS2A1Lv3Rysmox7F/8fr
UqGAgRSxrx4l1/Jc16dAbGZeUP6Usnf30c9kO8cpcJazFJal+7UEkbDaHvAlvWwcjXLAlZqW2Jh3
ZJgGPDN8gTdtgjQfs3RMScxUEXnB0wWIV7UYAdJCwMZdU6PXo1bF6E58g5Da4G0+OGjx4A5Ac5vJ
W1VJPZ+tVts+gQUN2sC3ZjUBqzg2zWPv2ik+uYGSUjGyiTqDysoXowPZps0deaybm8kT3hqjarMt
3LVw++LHMTNtkfHeW14ZvkPypA4GQakK9cELQ4sUect7XGFjKyV3/Hb/UVK4LdsguvvU37lNB8hR
QGZw04+zR/QYRUIo5uk14IwtfMs0j9fWMjyAX5t5dLk8rUK/2U5yVBQqoC94QYqc+u5KaVPlDwfC
h0SJH2Xe5/eLFQHk53S6XVQ41oACZIOr+vuOt55T8pBWnrOSENOc2znA6p5b7IeQfW+YyEmXbg71
ZCZVIae4M+vPT70HuSljZuuL8pV+Ae+urnjtnuEH0cSxs4xODB+EymfZajZg9h3R2BC+yiXPxTju
N5V5LSSRALS9HrK/Ss6ymiTBLJPNkzYiLYaPTGIUxhBYgYcei2lTXdZrbUFs1+NCSGUGYZsYlzcc
5W45TjMhUrUbdymvQMh/k1B7b938nlZ6SueUcTE7FPrGSGZVRsHhjqZiE28JC8yRU9n+ydBhLTWc
+PNC0n0AANAfuJZGXLpRRXCr3erNxClJbtTl40WH5MIPV2nmbcWsr55ZGgGzmpcKcCUJwTc04Itq
QBktTU6+nApgB+QhYzC/LXjasn9Iv0ht0+m13ppuZ4Ex5WfljoiVVYB4sZst9oUiYqS3/Wib2c80
9cUTrCeO7xtY0R1/Kn99pMUX4p7Q58NNDmAjCfYtU3VjUrj7+LbuNb6JadY2LAV6+zXKhCGGvcQ4
UUBjch6dBsg1QFmY+Yu9OpTb4i8JF3G4oKG3SojvCk1cMHiEpEjqXyiJx0FKobMdPTojpofq+Wh3
P4HSvu7PCilfQyxSPwu71jFY1nTN+nlB+lYLxPWK0CP6cz9iMiIl3xky8EAseSIYJXoolqqFzkpU
YCPEAUSf5Q0ywXk7LI/rDJ3pKCJq5kGEbeWzFlcAjxK3ha06x1MNq/x/f+2oXpMEbdszxQYP2HRQ
iUt88GjxyQL9XfY92o8qtyICrvUKo4d68F9/qS+DSE2YpBZ1pIYfiR7dou8EZUi4+Qqe+Ew5b/h/
ETIKIJZKZF4a8QS7N476iyBnF/9NSgS0WGy1MC08xfVBbNPL0j3+CFJhccE97lfBgRcrduk7rqY9
NEtM/wTAcxIEdP9BoKcAYT1uYRC1Wh0289RB9Wt3kdTCe8VXmlo7PuFPISX39S/9N+QdRwjElvuE
m8e2DOO5R/2lNlglbZJ/Sl2TMMe1QU1o++6+aTuwaWgzf9/77nopbAQ+uLIOs1IcGKn14WSnkYZn
7/VPQiJGfJlj6Iz2heofNFofNNCOSgyH6SXkooQuKKNi5rLV4XhLtAxczkuNFnja91qVK5YlCvbE
4xldJVQiso0SrXs6dDIKQGn2rjFUGMdiubXjZTVYQ1G5a3jOT7q5ql6fi7erO1wDT+S4n9HtUw99
nw1StgXiZ5Jb0kCrls5QwM1Pnuo4wrhTS64ayWl6iTpEkIoIkR1A2BY44cOlILw8UoHaxniCY4/u
4+BtcL1xZMKaZeVZPAIKKoE8NyF8wWLXGNiAhXxNjpAhHOtcr9Msk+zul016p0mSG3xCzk6wcQ/M
itu7UaP6I4l4D4BCvax951UgmJDtVcoHGmZICxFaKzYMoc72NC+8ZIXBg80es7J0bgZ7+AEQamKi
861QRNEmvqbQiqAHXgxYe2AOcdorUEMCMn8WdtWql5JOId2bwvDipqg8IUgwsM90wm/evGAjzdCI
+ccdMz4kp35UByrIKWxyXhQLlef539VT0oxzZhl19jo/GjKj9YABJSIku/EptU+WTrySgZzi4ugt
ig9YOFD3ieZxIp5mO3avjq4i3/nUbqGqYAzwJOJosb3BNM2uYtPlgIbn7j6Hk1TFP0xk1RPzfHXk
JvNjV+4eH/3YoBMHAt0PNgn+yGkK5tQNhYL/jVUKpAIK8alXzriteljCcVLPATbhqpqYqsLkUUu2
MYbG4DrTIW7osazgux2PuO87jgQbU1cTsFunpAw9nlePA/tWY22Y/Gab9owIKh/dDwzO42dXKkrU
P6+NVvCqTTjh8PL6SKOZVClVsYyfs90GeA43csLWVNl47QcxMiXaNp1rZSRDkjDn+CJJuTcq/zjh
GJgnkG9rL5OKckiEPCm/HbuubGO38rLQOIvdxVH+RpssiVG8foTNjKnrhu6fa5MBIKE8Rwkns6P3
jBAuIaEhvkFVw2kKMaJw0l4TBWaqHPiRQsL1EWUgK5A8R7Nr3969pxfa+wPjZ8IsfpAUJejpb5nz
GUtJyd/tFFze+Tm9xzJxHtp9JZas6DhWteEHyz2QxukVXhA75mfBowypm3hzvFuRQboJkJiP/yMw
cYRVjj2zMhV/tOENBfIppAAxRBiTBlFv6WAoC1tWUJSqVmKa+8UHRAKsDRVU8ReUQ9MfLxDnoooJ
7OBmamst+rBrevXhS8jIItX8A7Vc4lv1p23UdwBl2dgduvYmKjL+38ijv1ThKdR65Uv3bgYtUNAO
qjLh6YZXbiMR6r6YQ+HpsvZ9taGU30mQ8dMpc4LRmK8pWART30J2TJ0yWn7ObDtdWmwZ7GktEDBm
NDtaQ7tpGaBim87j5iPOJVtIa1ofkCxtyULIrwPYtoE2uEbCm4BZfiCUXGTcuGvsYufQkmmzoCSs
lSLH+4uqWdZpxs1F3/TnOydFjguhUkppI4iG6GolekMcm4pafVKDfkldgGzJ3pRvAmw3x7q+PM3R
tvNlUCLVZiP/JDTY07wX1PJDl7oDhH1Um+LPG7jDuRvwjQEinUWfGSWxvgUmdz+8ijHtywOWV7/L
Rj1bCnEt8oNHEEm9ajgQFAqO5RgRN7GmCS3KsbHBT0BO1jlp7dJzscoHpZv7Wl1qbMR9zA7WDrkq
ftWwjUxlfiBCaWvmJokuusYW+2xGbbYaEd2NyCJBZYryENUU/X+OJDbcA7Rm7AGAW3TSmblrszeQ
HGaUA2hW7ddaIDyozxK1IxlC3ZdP25T3Yg1ZjfGIN76IVHmuxRPaJloi11TyVRmHkw7fqhdLEiHK
1aHZw+YxTbbhOfmstbOrU+aFuju186VGeY/kmO/4fgs6gFeqCS0kelpyGjS/pfwEC08geaDsR1Iy
dnzC+811gPE9bnhIOWfs/2H3zspiqNl+OA9wbMre5fAsEGWgu6eASxnbjRX1epnaMMgeFdNMW+fZ
rF+5YWMXbCV9Pzb1KU6KCvPeC3eHLI3Cd83eN5sQrDluhjDw1d71G9v1XmZd/4vvG0hUjleyrJyC
XFEgMrogfx7qpQG26IjEns47JLi4WJRx5YkFRCMxKLSI13CrEXq+cMJ6RIsBth/mIGwG8TGD5Vyt
FuNUJhApimZ/p+RKBWmsEi5RdjGXtMct5RAe6z0Q7PZo0ebCfGtDZtnw6lS/sSEjZUOsasmC+U3d
0OBx639tbWQQGf/8udoETZ1ZnnjYxbxJTf4AtC/f7IzEpyK+jifhpPSjq9XVviCP6pm2Y/GXJ0qc
V7a9EMl8lXxvHYiTnmfJxAoO70oL1YM/SrBV0rjS5oY+z99mm2u2Jf5WwQrO+6uYV4QqpEh7RtOM
ITPsyR74BSINbXBPTUtbg+NISnAHw3qB2TXTLIRwJzQu8Ui50RXDhlbcjsNwe/W5TnvZ9h0KhQQu
Vmt0NOSdLZ2zQoM0VLGGG5nXHTN0OeuedXzIgWmAwNC7Ueoycoh+y5++Kw066YlPsgLBAsEVXwbw
O4VxuUx3qPRLqqfv4J/z3pDc3WLIWrTVO81p5uXeAAp8Tdt3HUt6ITyI5hRHOsLERkeHHG1V9tKS
87PH/ein3Pu5PshMzQIrUth+S6bNj8MjNrJ5htNspeJIvpo8RT++6Wd6WYDNYnIZifQaBYtCNyEk
H3RcJLvERMlhkZhb9Gyr1q+Jde5wKO58rxKGcydVaYhrqLbvREGzO62z+nDqkgsYihclWijluaY6
tqLK4GlKbRzzzQtFcaq6bGXpqdP2Yri9guI005PCfkauswgAvPldBdk5wb1OPW6cyJ4poBh6EzJ2
OPXiPs+xL0xxl+wlPx79Xh6GfSjlkQ/XzK/t1hj7p0GsRhOxpHYThJHpIePrqSO5axQ3UaGXJ+S2
bv09jsktQHuj8HR0eNgRP94mUZygYBBDgnfzo01pIUmPZ4gcYtptzTx3PCht/Ry+WRDVIziJSrAF
QUplDby7Nl/+xo0erXlVb2Oye5Gv8LeyB8UdL2szLPcYBwWjFxAUABpdqs/Lfwr8QCnH/61ZltUE
dAlWUQ0IwMcoQ4iQQMfsuOEH7nhtj+juGCYkZbg103JVezx/UPQKgSunAor4e83kOb2eIhJgdn21
09NzxdsT33VNclmqyr/y92PE6JYdRSr1mTBuc2iFTm20r2PXi4YZWcpB+Gcs6Hazh5mTsgSvrALd
9ZTT2g73g3Qei+/9vuHrFGdGez2J+4IZWiemnnj9RE8QA6/5IowJsCaHsln/BmuJ0osBOx2FXDgb
5PYKkU6ziOCWGIffkWj6sYlhxs7jPU6hZZ0VQUbQsGmDqA0Slr08IDWKR23Y4z4eCbVqnqogvV12
MGJDXhJvAjKJ32tC/RSlapDxFBUG8W9U8RrH5+Yvc8nCNtA3s2H8IGXEZRrNa56XYo1HrgFKe0Xp
KvTiXaSa1uZ/YW/DfWeVg8tLxlRfW34D01pLdiKVlU0ZxP7bqJG/micCua1ICnZMDHOLU/rpLgit
LRPvB7k/FhkFleVf1eVdoUfPbHZzLhNKPRbHaL+FdQl2zBmup2dHN0K/fDYCk+j1E2G5dfCvc8oi
zPcLUE7qxTNq9OAatdE88T6RMVI78h1Rde2z4SVJvEGQ3oPDZ4VTW90YaLG4Zk7i/az9JLbiWYdt
ggCAq2VsGjqkZxQ9TENWVNfhMSPvQ2eETtNlPRxP2AVlspvtQy67hIiTwlSkn2GgvgjmclKEdCzl
0m5v3NE1hqOxEqPTZ04+EBEkVD4R5FuGISEbOD1k48MWmGMnkWiaZXg0mKd4ziUSUv60m/AIzrLd
KTLtunM09nCTbRmWPrGf8u3PPJHMj2nfv6GaDwG02aSxBKwB2QndsZFALX3uhCLUYWSuyhA1JIhK
l1Rxh45ZFl/arLQp45X3joa5weqFiX53RdCZaapL7tNhCh59U3fbh9DAEICjiFSWA/8QipxW15lg
4oJZfNKDDUIHIcby9y17prdrQM+POCj/lmbaxwMxkjLsFObgby459oub9gg1PkAAzapP/ISE5p63
MzXVbqJaq8fYE1Fuf1mHAwxXGbrI7SF2xDNd7L3fyQlX8LuShzrXZ9QrmwpHSKl6frWa3q63dVV2
/p1NlM9hrb4rukx57jjMQcuAcLzdE3VSIMlzdCbJQFQopuBJ6B8JFWuCdys6X9nWzr5gMSebZ758
ONaCp2XPXiZ+3Z2v4o/XQXbWjhFFiHy+HIiNJLnHEEDBQrpexnDJxeIq2PUXOocxnF0PpHXQyLDX
MjoM3+V89FYpVM0IY2yRnEP0KOkJgDkMEtuKc+MrGeZOrO9P6pkPhUbi5+lsVeY0zvNI0GEVOaT2
gYB8n58W0GFlapzoBYj25Y+qhYlgyMb6/nEfxqa8FS/LsU5CjvYEY1FuD5IeeQHWg9SjnoX4PXdX
/VGxMfM/OHNiOrj9TdN5zVjHD4I7j77m9ewaFhOR+do43qQw/rc/ZWGWIMo6z93+rZLOa88ssu0W
QKQcZHBAus53ed9u0jTfLavvhlYfLt4aSnHDD7YvWtzkkeob7GhgVxXrtzV2JcSrc+s+NPevXIIo
CDqn+o6NvSKf47mpofHP64KoRyAowRhiiKOtQ9HhS8Rtp+yv2G3Jum2zKrEi56+TaIeUUUim1z3H
XcQ0G8yCl7oAIJ8nBXzeEW4B9j52NqOQ47D4Bc32uwUBGn5zp/fhbu7mK7uIRSlExont9bwtAyRU
aq9p/ypUEtLlOjjfAb/pKTxaxFzFTD2d3/1u0hY8NFi9BeXFLhiDsRLe7mrebtkPeOpGPxNKncQQ
C2JE+0FsXFrB5NkvBD7QHPJG5JQycKxi9vBL9yZFv3Rg/pS7BC1I1iZZ59SYcOXdM0AW4k9wxArl
ITJOPffIxj5cbyKmYaOzyuUchAIkzrQy6Jf6IEJnYghzX6XYM2Ngrqdj4MdiRZCvfOzOO6FA65st
pLIzWlkcrXcKyclzcsdV1JA7bBYta5WEM/MsVZJwBjdcJGj0QTpnjkGWhXsGlBFj6oeo86DE9f6I
mGeTzoxCy3C39HPiij7iOWqNVTsVMxaeKWIfqvPWikj3uGvJFcRuC5E/kf7rQPxwQdwV+kjGeYsw
rDjzd2gLCqdTWzv5fRsht07tJngoAkDZZoONwAiSBXpe1BgNNEjsrnDujZtxVumQU0b+odWHIwYQ
AEdjr99Uri1sYeSzd1mJcWFdRMxWiNyB1LB5ZFE+pddKTqqWqeCocAFaIor7ztHXYwl7iEnHCW3c
U8K/h0AVMhicvJAQdlFIO4av+DBbcdPiwx7bMizK7HDGQHLudBeB3IA+CAeUJtFvK9PChvOKqbz1
zA3g7I0kH3KKUoXWx6oxgYLVJ2PWshwFTgK7vkQLkrDb77WVaPK+1bEtVmkhSawFHCIrLOYv2kyc
bKs3Y3B1pJHILct2PUIeeDaqcinptdxVKIkr1J7TQ8EaI3Egv0QCe5/gOIHAboVLUPwvoJZMGX3D
vXiTNit5aLcu1Z8QvvidgS0oeFsXbnzpJ3KnL/Fev1vpw3hwQA9vpsZP1Z+skv6h6ks803Ifm5p4
BHEEb5NerHVeSVMwGyjrAwiHMYaGWxSP8Z45nkyY4hG8dx7XBUybFSFWn4Wq3A1fXbYP73hxHWwE
ONxCbq/CoQIUqaIcoPE48NU27oGf3PIqDAsOges1IazcxsgiDh88EE4M0nis5aYXE10UTpfKfJTd
TxqfnATcmJHxLsFITg/gSzuTzNF3cE8tUi2xiDgoxs361kZby5wzBIszEO5kk9Lo2xgpIrwhNz7+
ncm80RViYccVf3SYZAyvNSAdRsPxOlyjstN84ftdK7PHu9kcRptbqZNZXggBFStYz2ojRy0NDksz
7fuwWmmx10tTXq3gv14n1AO2YOzLqo1tcT0KDTi94JxqATQa4//O6RwQsBbNoDnysxe/8mBxt8HR
eokdQ8dkTkUuKBSG8gx+GuJciazBoXeE8cGeHwrlUynnCjZ20V94ngPb67lM/Fht/FBjsUhnL16T
jtdMk/QYd3ES5VzKx77+d1qqRTYxHUJQPfcpcKT0Psx53iLyx1DdwlVBeaSTpv9SbcjZOiSXF9LK
CBmX2SyK4u9MfE0Z+jGamRaTY7CrFp3MgixYBbLi/5/0Adb/v4n7r/jgij3vMQgTR6ryayKMgFu/
MSu7spHLOVj4Qt6nPeT8g5l3+xl/1+PCankXeNdF12IzhgSn8uErb5eYQaJSiCEK2IlHYVJfQvcx
xehV1hwdMnbqIHKrSvVh0JelhnsMl1IcsoQfAXBXGl07kv+6ztEWhO0KyQjU82HUNV7PX3TbYhbO
tCAZvNScw28LdZzVwR04nLTFBQe546Dz7DQa9bnmEcjb3Vz0NehpibcHBpyhM5ZF1EGPpCgpQPoP
AiYYOxkjz+Ix+EFIzYKdaC/jwpC+hZsLQ1XWpz2SYrnzBpaRKS5ACphh7GNVPk2bM9iEe6pZMOYb
RuhVQFjYifJcXh+z4svxJdM9Ev4CjtV7nZ5tPUy1BKWE4LdxkJymaOkUUclgndaVkxhXkMSNLjuS
FJvxdsItkLK81E3Fp5rhnVqmESMss6zGe04l2GpOZL/+/6zRK0iNspgeOYTAhYcWei09/WP6wDOw
oJiddkk7+8wF+6vLMm+jdM5BCOudGi5C3gXshcHSiJdEhCnp0s9vG9xylgG5bO0GZmG5ej1mC/vu
hVfunA1n0C6/qE2mKg/F/TpitsJmp/SmiuQJGKcmnp1sj/WHRXL2Kso1NB9y093pm8semSjEMbfT
AIV89lzLF8XdqiFi7VrK+CUr3ceskOD++VzgbEjlSwRgEJVylHUg88F2ws0i8clObVLNqfnnUECK
ZLPy1VK61fAQGOXVCLJqJniK8bF7UElC9t0VfxS/RYIkCRyiFIbDMBrePqQKWITyhRTIBJxgrPib
B3MaaEvT+lb51MveUEGOqiuWE+Ab4IZT1saXvRrog8VPAEe0MBu7+SrQKxzUqOKc/ktdk+ORm3h9
SHwcdILudaOkWslllWuThDtTvLTayKoYGjiOd3xe/6+wvut4/uco8MNV6arPAEjjMw/2hYXkave6
3pQuc+/4AlFlFNEM+BxmFSIbz7FAilu1oMQLfv8Iblqyu2kyNtDSfCuuLtrHKKP5c/iBugTRJa6k
3o8zPFWGPem0uEKgK+yhwpW9615+IliOXPAnOLaF0U3C7uqqPLwxJfxZfSlNq3QjwZe/xodb8diP
FpMCt8kmRpSFa26Ji9fO4RY1ebfgrVpKSm68GDgP+w1EWYgujn4HncyGRDU1d0iGfNsyOkDfm5OJ
VD1+Pdt/WiKoGJL5jyP1gDZnISZZM6pNkKBul0gTTBNhfvE1TnGxlVDuN8GaldNsUYCl5HZG4sDZ
87z7Gg/4+vnZOL9oqTNcjODkMkwfhi1YZva87KLSieARLpF0k4QksWKvv+mQfMDBLrh/WoBc1Nxz
q6ohOergMWjh91pdZbbhy4d2+9wQ6q2oTtQXYWy5ATs22nfOpyeAz0pI2pf6uEku0RFUX2YQc895
dDB93HygLm2OjcluQ9HrkewmZ/A37zDOYSi7nCUVxZCxTYElX0mqRDdLBb5Rui+7bIDDyQj7Jing
eKKaOKzh855scVExnnxdhLpWyaajNuFUb5MyUa0fWZ0y2YYbRibRPRXe4NXqGaJ1Y1z6p/vpRqHb
pSLljnRX0as1h3HjNLf1drBnuHqAE+Dp4gmrMM0V2wytzPaa7H/KPA/FI29hIH4PXyxPDiIpR2gO
JFmpsFqmeXnKl5+Kqh9OozjAb9OLAGNISpU2YbTkOr5AKjLySwBu1Er8sviOJ+2G8cSqTmxDAgWO
FMufaQpoRpmIZwRG7IDrNad4kFx+oFyDz+S0YBQ64Dh7TeQuVIDpBzlc9odrkNqxdpsctYpapuZB
0Mzif20yv25+jeEkwYBYll5d7CqlTkpmlObCESjdHmCaUBT9KZKEYLol2KhwF7+RBppJWLAhNW2Q
eHDVlazH5J0mdVaTUtqWPKOlmovKp3GYXpwmjMY/oKIZ3IrDI+mPMO63lu3NBPGs8JOCOmLMy+bO
4G3Cy8teFX70+3lp860C6pLOU048M6R3uxBR0OzPwrXSyq1ZGo/R30MVDX4eP3AAqZ1aEFFsceyi
cidwGyBpmKJqlnRmpQOPLfLm7CxrCsfMOpbuaM61baTn0Xap8IcVJIh/cUOvLCgsp++Psx5yDnjn
u2ECjJK/Wo0KLSS4OQJEPsm7vsNdz6KTlQGSQFrsOVr7DxvzwtgqwgXv3tem8Ml3A19ykm+OHMEg
u59jzKKKFGGmRMzU22VnZLZSGqLoSGCPM47Y61j7IWq2jsVi4u8VmnhahrVkj8Ml0LoNuNjZJerR
2O/h4hRpVqbPUV4Dq1zaUcVGzqzesQ6zpoEbGTs1SqYTaLgbDmBYv4c9OA6N+mNzMEg5mkDMM+dV
ZnLasfZ12wd9epTbZp+4FtmgQRttX54bC74kCo0vDpMcuBbX9QPiDotWHhmb9jAl2mJMEVR603GV
ybLF3e9+8BiRIVfhwCGvLcEvc6vDykNqvJw1lgGoJt0lpsrzR+1lZVesWbh71z6YXrJQPIbNZyau
EHL6YDFXs8sdTPxmuK3wJE7zuxeBeZoGkP4vvCvhPIQ3ZTMtBWhEB9iXn1w0lsHfQ/wkYjawqW7S
lyeR7hEiObiD12H4hzFwdCk+8CbvPtsXr7QNm6tRKo6fZt9/VD6XtzTLb3sNQ+ROyOojFcN7wbCx
FFlCr9+qAmM86ofACbAPMBlhbwi+L8xEGk4zL39SUfvlo9JmEwXJdfLcpErkUI6gZTUQHzsN/2rT
3r+38GHfxQrIynWVngJKO0boGLO9HuJtlVyUGLX/YSkFO//h024FUfrihqaweM0+viFnnZ27x1Bv
x+aScRsLhabVilM6ILSEiV8/ncpeE4ji9We0VlKJ1GpR9zqSgBJuCW6loZy3nYimAhmWAH9VHnhL
/uBXyZrNXJcBoU9YHMLtVaqlj64sYpgw2+FuxdjOs9HBcmDxQaUMxb4EhOXZlDSFP6affQztNwJS
zID0HB+m7cmHoIcgIHLYn3DieanHA3k1G4IzBMAozWMvqtE+tOvb/vwPK6jWR8Dlc6Q/VEPSlq61
AOT+tu5WJO3E0/wopjjLWBd9aRQHECwD2mXS+plUHc0daOXHIk8F8um0ErWFtWm/5lpfB03x7fng
dkQcLaOmTaewgQLMPClPDZod9j9J5ir9jn4pj99xlIBTEXQ3dJUuooxiEbUhPgD/NWIKIou8KqEY
zYUoWuCmh4WSMvu4tOm+WqD34oeLUPwggPmDEVLjTk6qwfo7LKs/MpSFU8JppjNTZYl8ctw/719w
7kJ9q5E6m9yex9klBkb0ato9lkj/lyVQB287oCtebbE2qu0o8TfyyVf41nbQofs2XAgYxnJFoI62
oUkZbokLMqnL528mm/NIx+CWJqbA8cvLgLA/74ViryeTtAYZRCTzqyvL6HBNpVWCX5/lfsvCImn1
MwDqqqcNC6qbzA6NdZ4Rzo2JxFT2OSb1Vu0OYHQgeGwNtHWm2HxbwFJbaobxAFeYM6buUIB9YCU2
6Ki/N/45gYKukaOz8z+7i+aPMuqk7O4Qp3aXEQlAuo+dQTK9GsqYrLp8Elul/sa07g9haOytMlrl
TU+whSd0bugDiydM67qMu4JsilulmthSoqHp2MPTBCHNWuM6NB11a7bAdaKvCnMU0HBmupqm3FN0
XHkJlK+EL+e9qawq04sE07r05imUcUbCNdks7SgQ1rBdgTzf2shcJIRQ/EKA7K06673rYh35uXvr
4OUqzrko5kZR57bw4iJibAnLYhq5fITSRFHua1oIPx1wKPTNlcuz4U4puYkBBaehPgzieBJBAU+i
XPmhBwzGBZ8/FNA8cblaeiNOZq2FYudKTr1mSP9EHI+kdA7okrY7L3HV2/1jKvpYFDVmwiKoCJAr
307IE0aX37jocAtLcjMIc43cNYReoAHAbhPj8jvPw8zt98v86eVkVXzKtOL8DoQ13QQ9fDTAYdg4
FHMm4VAIVZ6gt5iHEI0LhtueAnYoiq5O5WwBHp5b2HcKUpHYZvqZTDGkn5atGm2vu5O5SdyR8QS4
sS33TnJP+5qZGhfgwUBIzxAL6qjXlJUYbeQJ+YTWluwjZjw7gZZ0Pm1CZ1IwHbRUFE9K3hS6BAVo
4BaB+4oPYAZp71cklS3Q+HAwniwa8uYnHa8v0MPS+kwM3Pq1dY8uGXSvQ7ltx+Ft/ZXO1IVityDe
+4Yjv16l86w4cZxr2Xv+pVM2pA9Rw1kpFsp0fF0AScnkFG9Ly2GZrTsQyDeU6G9dTH9RqMmrmQjN
kHB3t0ys87NqFxQ5P5/E0hNdAB+CdYxUE6Rx0IQsbNM/BAXpKnZNLScKghTrOj5QhER3FCVfWPHU
rCCXUiYttNLVqk8ASqRKzNvkmFquvqpJygRYHCX2eL7ReJJ5Rvmyc7jVi6FtVkioI6PYAJxTGwLL
S8XfCntJwFvvgThaTmK1Hk9V9eJOHHcLzhW0z9B4qZKXxZyTydj3ci2O6mMGsjtgokf8Z2L4Rrsl
Z0FbSV7MFtWeuglR8CXkGN/VWZMNjuNDRaknXSKKh2juXiAv4WQg0ijGCQH3zdiqIYQPXEaTJNJL
aHWWP3RiOpNhGdzj8X2SYWRNvht7Q8QnPO8avg16LESSnogDb99azpGCbA2d5QZRP6m9SdbMyrbZ
HyZzV8J9qJRsMUOhIJXjqvZMdm4sDn7KRbAl/7UJ+CvTgl8Od3KYGotJYT5f92aZNvxrqAFr9mqq
qcKZimiiXXdAb/MF307bcf3YVUWanCuVlsHQlYI33NK4hfLKBz4WUo7qpFrCG/DlSnbM1Ic9iSSQ
5LIsbpn6NpuHDYbU6Oa8nLgzedH7DP9+NrYbu79yv6DZH2RDZvzRwrcW0rCY6VnvvCMZqjZlMcwz
b7MbtgK/nrG9LRsDJLpF1d94F28WbOv8pzJKgQyH52+Y837ICEqWX2x5+8uPbEKtezH4K+PqlGAy
Val1Qt//a8LftXcj+zf/i7O2DoD3GnkVAITXuqg3Lb4cv5//td4bumhD5m3BRIX/Oqns5C59xRqc
jIXXt58d7h48w5IWgYHQzSWwBG2kFNCQtrEt2E9tMdqlwoNEoc7q47HH698a8e0tujSfx0rMIRUa
2KFdrNKH6QO18OqVLODE4CikWj7tfZCtR+mgdh68AX6f/UBpnkzpVizPJzfh43G7I32BQd0AznEs
5znxn8Dud8EprQTEALFSj0/okeHa5HftogvNC2SgO1808+nEb6jFc2AelcZcM+/L87uJX6B+osL2
lJzl6vWWzPsoMcOc99jBZeWw9QnfY1d0SBkUzQqJ/uDVePR+byUSzYGdscLjXMGkUmtzwQTbTZTM
tirPmbE+IQ+LCfVH7dLdTz1WgeoiYXN8aNvZsYOSDAtvRhGubSbXXpaFLZJrTfVnUVEfOr6HSywM
4smR2F5OQTrraVsDKOfuoQoUc0Tb/aV+/eQIRasRzOhqVWAoVXWc6WcqHlRUTmldlBpM3g6SrJ2i
H+og4HRWMEMTBZeEL8yZ1UOM1YEmRdfjjU7f+Rd5lyv9I2IVuHktiRFbzV9SMEaF7RDQCrZqKvfX
xR7OuzxfNSt95YmVNMOtlpfbaT5eAPG6qV1d6ygseKQR8x++R8tKxtJdtPP2wVaE8NMOqKpHMs7u
hFsHTYXesMARgqd86VMVsVgbWSaTIzn03hDuXVuLXXTfGF7+wyrv2K5ynOudUVHPoObKysHFEQ/K
OAyx5cIY6wk4FLVaO2ISDlOBuWlUuNqyU9T9fB4vzJ28Xvtu6IyOCQyBp17vFEbNLQ7rinSl80gP
avck0RP8VwLn39Ef9twfFyhSvxEINBS7bSuVQQ29R84/UwtNpSsnxLLVx1UUiMUWmjmPD6i9Cfck
Ocs4IRhm2PmOfpypX7GNUgVDsBewA2eZeGx8ejVBCsaX9MIxdlyelgz6gNfJiUj+OoB2t5ntEAio
G8XA8/XUN9b+Jct0y5kJVBKBdc/VQoEH/jWTLP1YiJsEZLcF9b5VeRkvZeNuA456eBFhsMeDZJ5x
Gk1fFvTl0/E7OiNumEYlAQO6prc0EuspSJHUa47FabSx5ImQcHJidbdrYeqTFLEGdeOAcYGAIVVW
ToOzoIyQxYqTq+e9uQ1H3JOI3A2e3dtUqqI/HyFXvsx629sVYEe8srL6U7UBDclcKZrTTVbICUPa
UtGC0ISLK4NrCJFKitEekc+m+dA+fFwB8/7G5nJE97PjH4Jbj4W0mc+yRjoQs5rxvQC3zQsg0tsg
CozNwpP75+K2uAA8Yz7lZRJwHA3F07JTKG59SzPSEMoNEpHCT55yEGgvdEuclSXiMi/s9sJ70BLY
86unDsImg7heJMWX0FexoNZTCp08OoD7a12Jib4cVhzUV2ui/oOgrINqvyzwLljeUS3US5xctLXt
WyW4GLFUMelBpRaKfYZ5tMqN7QhInva86jazdiuLB2sxq6HLTHJCHwi6RnRdE8pD3OzKAWNJWZiP
QwXFuamsHdgOBJBP3RrIev2cibtce4vfsbxFSIe6r0RMdDoEkSsasxYhMrF6sfTsHDz267gwKMvo
6oM3KEixqd5dt/sGnnzl1rVUWqI8DmJRYEx83uIYZny4R4cEyURfAcLVZmilZD5DzHHl1qkuGm7t
mW+ODaTU+T0P+KUVOV15iXn4Xuevl9Nk7uerMNALdZAgZkPQWldCGccO2E+CAoln/tSPCmObW8pG
QvHQvlfE9fR6HPEM4oT7ljmyaqzakQ1sNaHhgkjfIAx968uug/8JHjIfAO7RNiSB3SfZ41B/P/4N
kF3byiMmNt98h3zRI2ByRpVHSIb3sHDsRy+yqQNeHZfdRZ/ltjycoSAKTY/oFFHC/nXiPCtCKtzm
+sImeNxHZn01N52fBeSvxYJ+szcLs3r4Vt16Wnq8tiWmqWiTHep7BC2V0oyNhpPQpfUeJltQOpZV
StvR0Dz4Xi/hmK4WzX1hwklVJ4FMdapDG0dpzGtCbBJ05PLYG9QeyYvP6yMmS8xRq1G1sol0r7iI
ael6wJGrqk+AMtuMp6DcAJXp+0td711q3kurGM0YQw0P6uAUOX32NcS0Ltipx4gt/3POshgtDbka
N9iuV3AdpAVsbj8+yo10LqPXsaSRfdGBURjLoFrIdat71GdmJdIlGrGbgjnM//auuHlNuC2KjQey
nXdc3dMZmltN1at8fDP2X7ZZOpX2fZMqNDygliYPg53aSSErD58xuzfBpHKMEeqUMmJCXrerkiPe
ZdOPrvrZ9EuGS8J2RhRAB0ZaQib3dCgk+0EidInRnlnODoS0MyJ79ClC4qkvBrwnc2lRbznho7tX
ya64R3pD3FB6pZMA+SYJaW3MKEbmD1yoK7nrEcBk69MPy2nipC0gIxTCl5S1Z88RiNlogcphFjl+
/k9EYCTKzn4/JeH0YY/2d575vf2e0XwkqSUjs/VUJKpsZnqlZg869HxkqBRhXQea2c18J0rg38XP
gGFZHhKg+vZ6cHOs58qWrfFHBfxUhOrJYe9+HN8c7hiHv5sr19WZlqZuq4CJdqYL+5B4vF3+yDY4
2JLtVIH9r1ihwe6gH6TSZTK6ZJ2g7X4NiFBBixbenvZVZVaRPgiybD1ZM1clK5twKH8a+Dnb7AFo
PhOA51s12MabqVoPETvyiPg9yVTFPJjSVNdIjAWbgO6oO/Yi4ProCn2tmcnDHtbTja7Zq470A0xv
oe3HIaUXzA4FkJ43vS9CoW0cytqRG3OGuQrHkl+0YDtnvYrYF+LN8KT7eVEpujbfc1bZh1CSk9Ph
WQMice6dt6BNn18IPQ3eJCGqfp0ot5gdr+jbIq04Dwg2j8bzpr2LlIH0xYWAQE/84M7oP3KFRbS0
ZxWEb4xB/ppoQeX+LWc4kKZBb8Sm/8ARrtEPTDyIH7OunJ6qR47CV4tqiARU8PBgFJHE4PwUP2U1
OQiYdde06DdPuyup/DaHNnX4nziuzcJQKdCK3E+D6A9xSDVNUKV2GPptcufU/lZRCVFLyUo36R17
vQmtvyjGFa5uECq8tj+AArMvpuc4nJEunutAk+IAqvSRf3yx5F0Zxc1gr4r4esZ1YKadZWWilrmq
b9MP2xy2Qun0VVMYp2GMwjFsEHk4sfYn61GOeZobcz0zvknQWrUsCWgt1mEIuz4Ob5ILY4975CB3
IBxBV/6CPIwdeOSS+dwPmmoCt2dzBzaj5/WzP1cV4GhifyhYh5DYVHm04RKYpSYZ+pjJkd6W26rj
WD4g/hBU73LHeoFfl73jdpbfx9caVWjC8B0qPFgh67YB3zHg7lzrXaiQdAMxx+pgxsTZT5x07X/P
Vv0O+rNLkF76ck4OWl4RiyO1m5xlnHqWHRIqn8+hPaLJ7GZsY6dWBR6CzxqWBMj9Rb6jmsjfv/4C
Erq+zjoVG2ql3BZ9gyygHJOwSkHR90Nb2WV4SVJ1z6cHtHSQDwSAVava97Fuy9yVwacvMDnA+Au+
RL1PVvFB2dgyEP/5j2K2LkgZrrufMQGE/avHFQp2r86SmNTtGK5t7sMrXeAgFJefJfTuXh1hu3f0
aVier7cwom6sOI+H1RWNKUjJ31kkElvrvtS1L6v1vJ0OeVDwP7E3lmCT0AqYMrAHr+MKsnwN4R7F
m1esMi/W/ihHHCtusL47QOi+UrUw1Ev8wo1PJFOWY+sfRS4pT5BKHu8IDSWL7VgQ8bUKLv1JpNce
cbGkJJsXnQE0T1htPFXYcnu1LRFWdIvSEvOgS2Za9Q21HKFpYBmMY/5OGp7QTB1F8IVQhckdrt/S
2qZAed0C8U/cMPbTdzDx89WX6CGtSkMNwogOZbSLhcJpxidjIm2MSAz8nSeQPBTNBFhE6pfLlKEY
J2at7Q8cTODeB1+AO0isr7fG5lOdWHZxH63bgyrBry1WqInIy9vFoKfQUFYBmyDspJbmH1L9DYYC
rhD7nOdzm2Sv4BB2Zn46gnHEEt3iLhLVMfUz6ajWh572XidjCov7hW0rbbzzMTfC4KEcBsmpgdLL
HB/7fi4wOAADRk2WPZIrCEuF5UZmsL+dsXWhanJhvwOZ7Dvpy4HRHCqTJm9GBnW/e1s/MfjlN3P4
TCzG1vhE/gwbWbU3Fb3wfa7otJvkQENXCmMDvsFE3FeOisMcpOcXMAxs7vt8U5ngWWoCZgUj3LCt
uYzvxrrbN4PNJ492ClY8ZQFiM9RR6keHkPTl0c/pqkw/7JSwTbExNO3Q74iU5eI8D0ncZNCEHvNJ
CqoKP3zhsqAjGxy9WnqgvkLjW7VAPBAc4XvbvvpCik6oodOLCzXqBOJfv9aIdf6a0O8Q3gc1hogC
9xhXPfdstkZFUtMWOIAHS0d3J3HFHP0BjYk8fB22bJyRqL0eg8NbOmwjSvNdOV+9OJv90AxjEU4d
aG5zpDBC9DIgI+s6nnMaVFhMASYGy194/NK6WOJNCCzOf/NPv2OXTfkn7PHvdw4Xnr5y7B1iKFWb
MjMRT/tB8iV4kT/dPGkTW+gQ6mbRCh8AG55E34R7llAc4kh6D8QMsYgYgGhZngVP6v/1/uuzQB3r
LBTvD1dTwPAGjtnFbQKflZO4ZVIHsuHag//DqlcMutfkpI/55qnBAZW7cXmfbgYSJHqIjYK5ecdT
STKvbMyZX3Q61/Hsap+XXI+k88HtTXQj67vpwqFbVNiPkZVm0ep1anGqYWGHXaxSFBM5mdnrrRRK
TO3lE4uc7hyBWftpI/2zixxPIhxA3navph/fmclDevLCRxxjdGuKpz+dOKQzW8iMLv13tPi/ciuL
JDvT4x4in/3ovncINNNAPNi51TU/dSn17UNVO0nvEXCgvN5G5pL8rPnRN6O5r9uI/fSxdVk82dvv
RrvU7YWWnei1yDx8Yw0zL0gxBFKCEKv1lGz4Ul1ara5bm7zpqfWim668KJIOTHMCr/I+Xlud/F9c
bb5181IxRo8J/Fj1WEMwEMGZippeYGgW9vwYuIex8Xy5x12Q9ELQ7ysIhkMQBk0FUsEzkVYVVsbz
WP/bk3+icuKasp1upFzzS1OLkE4oZBECmTIJokBj6mLIpXu+oYb+4t+oIljQqznIxbdGtjrLHLDm
8Boyy7t2623KsRf2m8TBHyV112mNg5piNDkdC8jm+0dGMD1R/3HWP2/RPm+RjBoaGKUIiNB5zPsG
V/UavY/mbBfX3EPxL4aDTWy69WSheUu1OPZHFhaAMVtyHFh+w1iQN1Y7lMrLFRaAyLhlHMIRjdyn
9GCbxaF6OXp0opj6RZf9NZKbpzFzhFAoW2RoD09bLl+X+uxftKrMc+7GWOcp8pAM/9uje0dZEKuq
qMklMrN63rUaix7XUWaR6+06qirpOSeuDzPlS8uc6uPI0vWNaFMo5hqV0CX1w3ZHbUhzav0GLcRI
VvGLmnkakXQHOpnnqvlAYzY7g5Wp1FvJuEYLLE3ZK4rmmALdxG89ocWqvzpM2DQSVOf5F9p/vnvd
YcWTx9lcJvSZf/xQs7CCdNnMwWoirgvvPljZZeyzwdG/a3vW41yb5QenAB2wotkk1hbvHS/3icnJ
CKppHnlBYV2JzwyhfmenELdcQ1MPnG96ieaHYtcnpkKBQwQQUd+EboB66AYLM7tzN/997nMO8cDS
6KmUq+q4OjAfQb8fE43NFXAzY6v3vSqkK+CIf3IKHqFz3NstWCO2tTbe1KRrGUccWuOto/B3G4lh
2ADGncWlDsHaGszsqMJDC4MSlrYU4uK1Xwt9X/S3L9rynTssJdSyk7iInx68P3wVyJ/DjnEn6wYy
2eamZypGJPdmjx2Ccfa4sN/1zjg8+U9iH/j7EPc20F82/NNEslQKqUp3SieFozZeHPZjOQW+9cox
zBFpRFbiBwlEYqtASGEDegELo2VzVqEfE6o2DjiXp6VYFZxjOzhUNKPes4fW2+xzesqFPHLfnhB2
N2JqSYRWrxN29eXLMOYiMbif5bESq4jxXlIXNeJnIGJgYWP41GajhNkpcKEZOi/pdKgOIJvYueMW
Ib3A3kgxvbrRwbFzrG1r23ZPJqhKNlI1SDLlT+Q7XVCTGmkr9ebEOr7j2q6c9qVBhhVIZY8/VaXr
RDy00W4vK8qmqLrpH1juPxLzNVb3oHQK15jmhx/+Hn6JTEiKiUPYswRSv1CdmrD2P93syV1hOgS8
0Eplhib/Gkg1ALBZEV+5glgOzha6tRjBFssavDof28w7U2F6DB6NoCJkW4I9aObUAsRMwjBNXxGO
Dv7Uho+ca6DUh/s96nvOP2QL6E6BXve+vZNH7Dra/4r3LOByfr6TfStX6f46dWgGEVSVyyFiSOxs
kvNvdTp1E8DaO7a9odukMxxzqEongrxPyIG9PBVbEe7XXebioVtZ4Fai5BLAVDQyM8tKiZqtd1pZ
jO3evk1SuxVrN3cS1/+4lSfJdMrkCljvScqXQfOHyTdYW2vFLBIuKV7wiXrFp8gRBKhLOMTvkkAU
578K+GuW8rbuT2tJBLw7OCpQLnDbt7dRBWDY35d0ZlcD1WXirqX22jBAf+Vr14yNQobnE4Ql3fyK
ENtFpcGai6x8ZpiXA0F6YDkiMEynGMg/TXkRK06LVuTrQFxfZlyf/J6jyzTf72hSNcSWL/3DqJFM
upJj79ehlRoEgT+C/mffAxfwUQkvKB2+15zlfePWq5liECXhRFs1rAitcNVlPHlJl5WnynSGj+vT
CisUK3Jv4al0sMLmrkUiHTjEn5ufNup6jQjR1g0n6yW8kzIDfJ5l+ymSnAD71Ez0oBXLBpQMYXTq
cYsfR3oxwRnVASP6k9t488fNHwC3KRuwBDgtwWys8X70jppL2F9XPg/dJYBxaCUK07tNXETeJRah
PfbScsp4Mv1uYwQVwLbK1Jn61iK1YBomp6HfHDKAZ9cj/MJrPfPDVsuJHNtvg+FYgZgm0l+HzwsM
87Bjrwekc+OBA97qX9kd4gLDaIGwL4Mi/kPtRaceaUDs5ULP83Dd0iOWS5e+xzwbEPlNouHhF0P8
2Z5vE5WJO/wODP77rESLFlbWhfejxDE+DF5ScSKZECl09MVmwJyTnexYrMXjrhcpPAkjTviXHkzN
oLUowghLYAP9qe9OYXH7VP5zPENOCdytTHpJnsyodFxB3QkVb3HwLyG7vGzfSfJYvqWNSNycCDZs
dQfjCDJnVVrt/vhoyeBS85Pp3WCQM5vNe0hFRZFrSzRS1lCzE3yd38Cp99g/TRyNVA8xMU8tY+kh
HJlsXKwegkM3UgwRrLvx5wYwOGPY/r0HjQpQfuHy6kmT+trrXtZ2jo3LWet+CIYp9/aN5JAGaKan
uVEYALZ7P/ZItjjFOBiPqLgX0nBrf1LzJWtEnPMOfw6DhRxQTKxE7S/DIf0ybHJdwQDFX8IlVyUm
nuoTPMj/zr76wH2HnTRfWBL4KmutRFd0Qt1sUdA7aj2yoWHACL1ViFJk4xJRKOV/mkBIBZSiWRdJ
ExxUkz9vWKV+8596rmvt42EQvjWsaQtHTJuouE1A9B69kAq/xammtT0Au3DZ9gcUWIZQM6DuSHdE
SYQv/2FQky+EneYxPWPrmwYAt73OS2XARsRtKsabXFLYGT8hxBO/zsSpIQ394G4F4ejlckhbsDyU
1bWMf/69YFzXDnEgw08mF56vnDYnXpiHUsBrVM3IaSgWNjBP1K5KDstlPHtpCBYAV0UwFeOrf6Ht
/yS88/+qG3/pB4kZBp4MozjOFw87U3TX1T7DS4/CyXw8zNPAle2J2dczkHoJNNufokU3OwWT/HUj
EzZUcmH1qhxXveLXhcEo76JZ9AUeqtT0ArgkFG+k/dx7tfmTkz/DRWoJg3Fky/xVW8R8c0dq7aqe
Y31DC6uFWb9fDKGHmPdApUtUbl90YFxKdEmEIkaI9XLk8PU5wtas3IKMlovue8Ydbk9Gsp6lNv51
rcOZdm92VRIric3z45ayy4D4kj+Ba7f+lA+5W4XLkvqUNGh7T1RZvpZhW++csQArOX+ZM8IqD8nA
/GCvIdrtHFoTCAppGtgPP8if0wo2UiIbyNiEzSn+0UMdkMrJt5cf12Pt1tj17Dvj2xfZA5c4S7dw
IXS9lMANiMTN7QwJp0X9H9f6hNQI+2xS0J+WJWZzGS12dRXsvMtmYJtbhXy3+CvX8/GC0n6K5O4P
9Tq/VoYSGWFuTfAiswxwN5SRNxDe7hVProxjtixR5vC3wCjHK1fDtQHkX0LQlxwDrPpojIdNoSGO
hHEK3LYOhpCXxC/O5RX7CyHg2zqqpkpVompzVTU/NO3hKCmuXGb4SpfK3Dco8+jzZdCJOpBO7qma
Avo4pGU5kDd48hNGsfEwaLr+XSt6SbzhvKjtGbFiYf6BTSzPUnT/Ckt4Yv8K0X4buUsvlQYLpcGh
CTCxqYJeRlCpHKeBXUH0RL/9lQx7kW/n4lZJke8y5IXF6968EISLDgY4rd+jtcIxHby+NKNV9P3Y
o/uAvCkdAP6sStgb9675QOAGI3I6jNH4nl6t8cFVG28u/LpPFwmwq9rE70bbnSNMU8ivJhiNoQbA
PwdJk9k6RVg9xjgokLbK5KMhcaam17BkEoLjZn6jkhZhuKu5/tBl0RIWuoL7EX4jBmfmHoSqhIir
uzcRqZtwfYwtyYdLh6Tlh/zbqkplAxiY8tvs/W+3MkYGvSk92aAS4MIqTArQ5gvrcvwfhsNSG+TM
Kb0aQq6z3TNN6xO+Eplh0FSIUR9C6iat8uUY1lBm8KkVDDBpmWcRIv1ujW3kKMFZ0/4ib5aIa7k0
NO32oJKzRJ2cVA4Bcu8atyFbA3wNCKoSffWSVUD9m1RsC9ttneynvCb90jbgwm/ACzljTNKR0gX0
LYJOqK2QuTAcSGhMlqQNZVaHeZUP1BxyaNyn1f422AYevJ1b1Kflu4YmcQJKLJFYjSHTgSekPz2K
XC1gK3t5WvZ1oTsSAn2MPg0P9IlM7WpY1Arkkm8Hk5ntLE3hspz3vUUWsk0g2G/2AMCkZLKKt2NK
NQTdqJMI2XvKUtU3fPGRDYZGE0yxCbbx741U7crFkd4xhj68DLxiFgYuWKgCSzx1bBdIbFXJ3pRJ
GUlLt6m87kwt6F2a9j/kZxyOb88G9VPk2EFMmtqHt03TN1v3mv8FOZhaCaAugO+YhZKtc/eoGmIi
gS9/ICCYKZ1KR3/NEGUV+tc3WBskk9RZHYfLBFIuME4UOteDS8hMZOWstOXsG5l/W7u/81PuHJKR
F0qfATAoc7D+vfAn0EIwi+RSbZG33arZ5KlowQs8X079UH4MrEUjjK8aQ3+ri2/9rFK5S1afgJeZ
j0jqavxhWjBzy6KCz25wte58n9gdPbAz6mKuGmeSCz1JUSC6qM7vvkwL0zFIczR1lVNvMomJrRa+
aWuYm9S3aN9TH4KZM7XI7lepCdQ3yGbRqLYORJ/am7zVh9orXWJHNpm9aqH7a1uMpJ9esL5T1Q8N
dqzhyZFvhOxaiHgxeh+pQY7mNFr7wD9Is6rO5e8ZQ6fRrrwhKADpJvlz15mZknQWW+PoOzxj0VCY
U0r6QR8VWBd1sii/0hibZ/qM3we0ZXQOKsEzAzEJ1MkTHH2HZ6VVl/fAKIgQMCHBY5OAvRwHJtQY
k1FeL24fKEdc+HZsO22EB3GmCPhfH5XJMauHlR1dTClARxMaoEpcW8WMhc1VQjKQ3DrfkkvPgrGb
warZ2XA1TFbpt0RwfS/RgEW4mwRStym73Pz57cr0dCBqdPWgVEuap81LtTF6ZRF5cpZ4LLu3QvFo
UELVSGG97ohFNaG0u6VQKs4RPefqog9ShExHwZx6pf+nGwjV6j8+SYdhmxKFv5kLsuUPb376Y81O
VzY0XREwKFnX/fmRM6CTyqRzIDDCzD+1ZHde/Tp9lLw6Xvo4SJFbrwgTMtUGZSfqk0bPfwFfPLKa
rSp7gShS9n0pPk9b1Z6PPsIkcQmJxvQSUerPxMpSW3GK7WLAVkxQUck7r394atVYO7n/o3V96tQI
EpiMJLrxDzHYZsn7kVpr3iiKrhu1BRMFNb/RiUinNcEdpfxSTSElocrWq44GFfD8wBwjf7NLJSxk
luLD7eDLLZ3iYjppSLyQ0D3hJYdYWiC9/x7r49XitKm4zr8ceIWltoDNQTvrWLzu7ZnfAn0LHAbr
WSGg+Eqhboww+oMpTfWCKzod+mR6gXxGfAHcnRp/VDc9sB4THngjMPJFOvfjmJZjDGIvk6HD4Yun
dZKXHNbjbmFC4vBeo/YosPLXsc3JTB0jKsESmJabtUdfi4zfa+8Xy8wMmCBOvo+oEnrY6TO9jYWd
M7YZwnJ7IwA0QeWijgY1dCimVOnakWnSuJsvaQsi/eTnanM8CNP9uPfW/xnCxcq/A9yOqLAzNzLB
ZpTKeWD58fFvMSCZyT4BcU7m4SwIF7DErlqsLmyzMo2iGddpQE2Vuex0VfOKex05BVDWdqhFbPYR
7hCvEoP52JJyydKEM/i4K4ptGnMzzcBXfTPXpJaw3kSuiVeTou7Euh8jVPoRzLCGc8a1wS6J8RH0
rnySDEy5249oQQ9ZPG4CyZWLyUDv+oHhR+fo6xWU1ocdkGHqXHXMtQ0y0/5qTCuhrvzWYLBY5tox
EKRE/1unWwwJtGKkpZgQNkkALjaLzXwLYKPMlAzKV2FzGtuzljkThs+zvWcwhJNyNuBMfGpA25xA
8iOIaMjZvtl6YxxtmQzyWGio58YJ6EFc56tccZ1lq+gBZiYA1IpDPyRk5pr8G+ZeWRn8fsccSqIN
0wkvgpQ1VNEIelT5mDMxqun8XbCLE4N4CLT6jkYKvVCO7BIq3qe4IaoQHYr1AMHIXzNgji5QT+lT
dbLjuzdNgqHXyZzsLEEKg70qcNcYvBaYxT4tw1PjO4/+wv2qYGiKGaungppkVxaecJQfOhbCqThC
hsdtV3PHEPRR/JDMjkVrIXI80J0cKiH2+VP63Dk5EsNx8KOfeiAWsrlnoxHmPZAUK7rXNOM+8pen
D0s66HlxBI+qVpokKIwnqGTIyywTYnARreHvbct0VyNwj+Ixp9M5u+jZWQcbCsjxR439l6A84jB0
JWete3ak4Vu5UT4DzDBG4xWfxooFtinhIKM101+qhF0yjqhizj5zWYRcsA6j0lrNj5pQveqEjU/F
CfCwGhPD90uoyeAVUIlk+qHUyifwIjBkw7ik6WlBi5hYFxIOWaMIkwK1rWtnKFldmLzSTXKhZWhH
O5olWB3sgUO7AUp0Hkn9q4EddWSyWgEIZOP/Cnq0yzxW/X9pfnpxyM+qpNbecgJE6MYs282G2xOH
PvE2+etvF7C2luwaNEUp+uoxylZCFq1XNPqrTfW2AzTaNsnOQYHQcuZMb6auBbKa1B6knmOCkeRR
7Ek2TK/XDzrEVahXA4YDvxY9zj6dUQAeatHHLATod1eC33RZGqX1j7fgJAWtQrrLaYygubKY5Oec
DFn5Lde1aH/TQOz8rzyxMsuadV6t9VCXO5k9h8cmL5DUh58Wsvcc8BVVe1F9E7FJeDy2byj3hlDF
Kg2WbIYDfiEw0vI6qu+m2+1crBnLViEKj0Fun17gIM2aQKPE1EPfQAG4xXR9ESDAgi7uR9mhTu31
FpTztWCcKxSj1khheSfRTGIvN05obpLFWjio1VDIGSbUaIgEfo7tVvbOZyqrF/ziSl626ITsYejl
WLNVj47MuqevMYbiKQEjXjhAk1DvXV938Fz35oakZFHweJMc1GKRWQ90+NLEziZ0iNAwa75IGDmx
Zw0FcudsRG8NJTVEt96jbbl1MJBmg5Hp2jlSU3+XCg48J84yjr0KU/aM3hygdPVPkQuyVAyIkyLx
tEtg9CogbZVKVQbtq3cPDpMLyHgA0eMvO+mizE3HA40KHE6v0JHrY0PkE+Q9gVSbYGMbMPQ9q6eO
hRyWFRRPQjxnra1MJSGnPmWD2pnej6RMrf19JJbtJLhp+KEXUq8IG8KGs37wbYcHCsYlf0PPL7ER
RX25/6tNmsI9Rlb2jTmO9lG7WeFWCT/mgvTDIWP7EClzIY2DFzRBa+0+Tg/smPPzFXrVgfSWvwHT
E9DRbxndUfB9GCgDdWV7WqTm8hYVm89xsOy9PriItkwV0oVmYUP2R8pMDKaHzc1bBthQgamKsy4d
madS2y1/lnPzXqtVUaQC5BdSGR+cNLHJJl+HSN3dDkdHkmUOhH65Ye3boLtL19QLpgkOQqrteFNZ
i5JedC0KLaQCKR02ZWBgvmge8iJ9lRcbvbBq+C0g5kEf27E/hLkcMUuujrGqmQRhtO8kiKJiDggR
lB0ifhPSRCrQRtzejE22ilbyV/l3Fj9hoYdsNjnkXU7HHr1mnU5UcNyPRJCuKn7fgD52KnUD3RNZ
plNtwif1V/I8mnOZ1pm9hZkaVYWTM4vkfYEid5AzwKfR9TsOOUgI2rk+WoNP+QIdD9A7HQ5lHYSb
7VqtLsCMZtdxioDBLU6pXgeL2dS4OxSX5nBaKI2URO3gZJ4oK7b9UcaNELPaqDTB8lyH7vEtJAaD
5Rah9op/WdNh6ehW+nK1ly6cZ6L6cLnoio3DmPMBJfZpeCxhqpSo9X+rM5LcUInXRKcuKhzY39c2
8ljN7bSJrhDM1kNHxvke4X4YWx10a5bcfeiDi5tc1ttcfn04FfNiBFW3ALfO1rpIEQ9EJSk3bk8e
WM/pFJAQeQHZDK579QVhVFmTS8fYZSIqI4SxBwTVnq/6hPjE64Fa22QfefTg92aQn5X3mWMXxCF2
Z8T2cp71fxzyxqOZIlYslT4JbmAJ2N/vyMZkhmaxv97u0yCJ441jr6FJl3BikVh2IbuWmeqW5CnQ
UBvSeSzVyGi7a8H0PXsdHVE1awGawrOa5Cl4vhTJLlMv071CYUfgrFOyTXYh3DCYGmuk8Ol/PBFI
KHGLW+3sXhfDFhmnwlzriqjfR9D2fSsxWGa3obEMnpf324ATasFxKf//aZVvqO7JMS1OPBX3GCik
Z2wShIfq6ZtdKTkHBBVnlmeE+hCvIMJ5QOrQanYbzj/ZrcSljPtkW4UEAoMIDyCd7qvGB/6O7vm7
0tlSQQCr6vJdukmOfqSZHDStMOtE7sUT8ROZeLM5TK6UnAONfF5IGHBw+4LhuWhdJj8xFC0dgFQN
/G4DA3NQOzk5+KRaehRziSUA5CK2bNWt5HrBJJCHZUQdj08DrjTMC6u6skMGVnd/kLRy0iri33vF
k8henJMyWP97bD520sV/ZadXn8jDJOUSd8yoT6KhHQqVbrHGfsI+XoStyqOfc2cIy23aJir/br+T
LeXXbZXTDDcg8HRFyelO1dwHMfswfVNrR8niV8N0n7r3zVILVuXshAhgP7G6++luZ8DOPytcDcMn
iB4iW1nad7EBet/Umb3JMrlI+zc/IJaG6uoEygD+ABXi8EBKyw5xpCCj4eFhovj9SQsZk47zTAyl
q+GrDDejW+laxdd2ilYEK7StO7LJDohIlptpUM29tafa0RO7l2hS42EF9Y9N1Rbxb5Dvm8egkDTi
cLR5pwMxmUyTKc8je/tMMp135P9km3ZZOH5C8nmBjn1kshVooSjqzD30b561adykUt65mzDwuw1a
Tz6bJ/SXcxWPUt1ua1JwNLaKqVKHsd5Kk8romgQD5GYTjipOSrpWH83MxmBX+O6bzBLMj4+VOSh2
UeaHbuYD6Uj95hw7waGJXVxD36T7yZEG95af9HNU/mKXXgxTc1lw23gg+/wgRyAIKaLwd6FhpIrU
z8CSqSOdqEEQ2q06GidPrGMugLA23pD8ySXAadKJkHRiJ2pzBbjiufQN4am83t+wM4zlmLfSK0Ib
OqiD4iwNL8wk1MKNOL1d2xiLhGgf7eVzwaq1wu6E4ctxqKgyBVkVllGeIwgVQTU/iXetIabkWtZA
YLorUIpxhj1SXqFxBJLgfR3o6DhgQ8wncbedP0lZtr0ow5eY9qqahrNrSUgMWieCPM8zfzYTPcpV
6oSGuo+LDLay+7OZidm031SZ0RKczxTHhkYBtTlLIaD3pIYO1q6uB6NssyXb7BmKqUD8UJx/asHE
Osad6EEm3N3iWcMBvuzs2fV4L2IR9VfdnJRmbdaOn93MDSOH6VTAzdedPFznCV3uy3Hlu0cnLNIe
VFUUw7RowSZcFhV0PyKYnv3fPQdd+77puoMDRQ0lHLWeskEke9k9e5rH+s3/XI3etFbfyd+d2SjE
NM9TS+ectdu401qbT/kkSjiqIMlgDOBFKkyzbvODbUdf4WBzDh2E3lrKpj0KX6w2s3MbAnqK18Ay
8XEaUjm3bK7V4RjYYkuRng3q9hnvHanwnOD8adi2uRadcgudeGkgY7gdjEUfyz52k8ZoMpJH4cYx
xJ45Hn95pDOun8D5oEDXPzGjo1Rb51k0udhvx0THPFPVHcsTB/YaYNxonde81yFmMiCJNnX7V9FW
nIilKsTvcm0nBc1hCKA/YfYGim6jQ8/QHpwvUF3pOIHcSgoLNiKB4+MwmSny02AsQyBgK60IJzHO
QS7pal1pQ2IHBM7VGDSFD4tWBSv/Q0sm9nWt/wxE7IPnsmGpPpYmnKYcU6ezcuSsACls9HMDmJ8/
bGXllWH9DnQJvMTZPsj/sUaQ6bSuabYz6FMTx80QhGgnriFrGDHzAmj1+qGlUjVGnBlaamIxXsT2
WLiparGnJUmNQVvXB6+ihTzua8CQxhSfeuJva5d1UujbAQNzmPdNCj6b0HpatUG+sFCwy4qtQ4Uw
sQSFaBRVNz9YmhbWZcHSBpfeAkw4UvrCwwk/wQQ5WnG4uilA5XmPMxbyXK4Dklmw8zywqhNDXEMN
xP4KjrbRsub1OJN9RQkZrHKnvqfRjYijtOZ4Ao89Uw18npFCqNZEGFZ3uscCxhT4xQunl+D4VYdc
eikrNZHHJWbgPqqs/bArPvK74ivamcYP9UQxt7dHfXMQ9ZgTeUKv+jXPdMIfFCYrXltV2wtLDpzr
7jJ7CvNdpdwMicLkeSwoS3kh4dPyrAQNWxPWloHF4dYE/nBKu7xDLn+1y9f32cCLkjUkXmgo7Skr
zamKLJnbWqiGpo4hq3YtmVCxtUzGQGdCX3/A4qPA30ZzraPDRRgFbpe5rh3Ikax3dVwnQfY24Wo6
7YePLNFbJuN4xiyHpm5UXlorSxdfdQhvuDW3KD62yHFXDbkB7XRwMG2t1Urr8ncePmla64WBtl7b
jmUSkLi4glC3bXx8z0deiAKEU5+D1HyymOETMqy+jCbnP3AktjGkc8fPr9Rp9B7NnofOJqF4IO0t
+irA8nXhNs0z4VtK9TT8i5sKH+cK95mnHZaaagqOCg4IrauP4acYk+KcPsM2E+PNf951clxjsmFx
FUzSJmOtNQNn5fxIliJTYu8sUYOs5J+irGJq6Ujp8HI6FZZnCsFYP8gpZhiaogG4dUmsGlFMv9im
exwL5yUOgFTw0ZloKRk0Wjs3Gb9HTfiJ8XWyavYyAZhBUJtML6J5TdOxdpg9ULMLlKpWjySu8IeX
o8wqvc5P66r4fkC4ZuTzCMX1f0F1GUd8y13eUjXjjb3enwR6yLXiZNMZjJkaNTQsi2XHe6yfNPIJ
PmNXbS6m4s/xvJ0rPQBCdVNLmupUP2jOmvSkw8AcU0CNUYNO0QjnFKUG2gqv/2o3m0Ukwim9RQos
gihLSBZls1NlwdXJovYdR+1yWeWAVj6zJ0YGwpfVSxxppQsvXSfNeqgkdnkk8XmES1zATS/BrRrP
iN1/4oehnguiAC6MkfRiPhxDbgmHeQcj7Z+bjEsVdjJss7yQ2wacYekzSMm/4m3bGmk42CRmGpzT
gmc3r5C6UHO1QKQ5XPu8swoCRRdQzBB7p5sGsDhP3AStDqQ/vFaHz/lKek6qnAgYSM4/2ev/CHO9
21pUgGJnKiRR4JZknXLnMaA7B4XaIoqm3tkTWUV+31Kha7T4Qi6YONB2bkIblzU3+B5bpc7qZspz
zQNTq3LTTeRY3B4lmWR4bKakKgxueSCJWMxthitURffe7lJETHOimEYrZjBPdIq++w5zIrOv8OtF
xAPuOuw8s5nd+hgGgeuyFDbrxqWEJQHL197ROY8ym/AL2PUr3BQYR7D1ft4EKHkQIoG5wi9VMHe4
TsxvPWGYCICMwL66p+/bgTTSFIPa8GT67uePFSERXRVnbAJfcfT9aQyMMDC+4Vv3aogxT0MwV0A1
/XQ4GOZlUe5gSSespCq+C94Jx97pw5jHEvozVwbBkDy32Pk/dn27GLeG12TweaarioWxYoxvUd/s
qiZukSaqSzWCDde5xtbARDBXKO53lM9YMJc4NK0qCtSvB6sVL9xUSQh7fY8AW8Q1D0DUuTVmjwTC
I/3hnOF01og9eiKbcC7ZBhQ0OCPWrQV45JYccBLu/qOZx56uZf7dvWbEdTOWcdWcAa8MFftPghT6
vUgaRTY9lUjaUBuMNNJHxxTMkTewLDqwz6CzLQ4jWgMpF4UnnAp4Lb6XJn6mEn5leXKU7Ap/nj/2
I2GUzALjhAWOpLRRhLopGXGB1mTNT0yXDD2jEWwNKitJWQkAivTvhpUf6+cUwYXvDZtnIIowyxpW
D+MWv7b5TDmFjfjxcw2LXZvl4KQZ+YaoKAR8eME+uG7lYM/qhkx42azcSOcgSG1zdTAV6AJMp+LS
4qUSPjXq6xqFm70xOHoTEknxNj0xzI2VoTluLqxbEz+VsAiICwnhjWbcP8qBXfSlYhOfjQu0SfWV
FRzGQRGreBfLqKNhOE9QRhrS8GRev8+m3zXlspw//tNqBzFiQlRJKrFQd25aVI8b76XlzWxJ+I9k
qT3wBpyo6xJmVtDbFahBlURitMlbqmgRGXB82QkZByFhS8YILoAMA52J8Qhdt8l5FvMC5jsUF8kf
0lfe2F+muHmcDkLnFtwTqaKFv2fommvFIZmdcJMs+K5dmae3htHIB7qKVKuaMC62z01E52IhDl9+
KZBJEVRfDubVyQiuTy0AVX8VWgVbqldeI26siSIfYuHPurZZ3JHeJxG6K/vdrPP6Om2pKyueF1km
rJx0rrWys5APYcD/habpIlV+YHpsXtH1VmlXdn0ctS0127gZPUD/5PAw0gTTOXkVd7pUHq7NAxUD
n1CDtu3B/bJU7rzPKaYfrFeG9mhy+RaFO6uk+PcG6b08zKPmHCWdYki26OWoXCemWRTxCGzGxqXS
IKIQLPmJSDp8ExXMrk3kwGhun/hpyMlTGT1st+bAYyfwfpYZ2yrYggYEWMoBP4UOFpyR8SWsmhtA
xmso3w+0ITzH1bvLZU/FboF2VDZfju9tvft6kJRVDd8zYZ7IdbHWxQBEoOp3Hl3euFCcxmBXncyd
hmAs0gpNIOoja+MpEA7vVgNllqJiM6jyREFArLKDlmG8/k8gfuj0XJxOWwwlDz0H7z10KvN4b8NM
bS/QVAItvThGZNnD+FAPPZygtoOQrfeBoEoQjQjEVCmVqZkjkXNWrGOBRt8HXK3tVC7Tmg0P7sn1
yKB28ixNYp1AhNoRvwET1whAFO6nLX88HGOnahmcQIf4BJUs5iuPlivAFAVpXIZlt9Uq5O7PwY79
ZGRAsfqujEp2g5iHbJaWHDwah01EjeNiDb1PelHdJPXdKahqr95ylwMiVC5Bor9HMgqYxB/1kH1+
vLY0oT6s6sbrecFnzD/xbfRxo+MSkaLztw0hV2tkHSfHwv5R1dU/jOQ+Z5IU58yxmcAdc5x2vh38
KpU+FjSqP0oRrtsnY5ThR0s6815B9/qsCE9LctdoYPq9RnYZgpKPnIi8q/XhTG+TFmW6gq8AWUil
6fGlkgeXrfbQ/zNcULNOMKrKkbd2DbgaxDSwpEDXh6KWSmwBG4FQr7MBybjOpJQS9hIXDMAo96MO
RxfJxrhY0Fq5U6WVAvr9mH8LmYrAQuoq9KKeJ2sXBiXqOCcZqWjR9NLHgjS50pjElseqHy0lhn0B
ICScTXAPlQZt5tQR8NBbwIGZXxLX1D2jvwzGkg93yAppDhNwJDL4lbmvQQzq81UtFtpEFCi6nwsP
XSC6wU2T/GnYLX+ECWM32b0kUvBFz1ryO36zmKjVyfWZ0W2VUK7lH7QD916u7RChSZu+7oKpPWrq
i2xAqXNcWlNR7cwAMcrW+Ixv0mbTZPuiL1OOhlzf4gzC++aeCFn64YlLUa7goTurB3WTh4+bZXug
WW5nSKp/iIaYVBxay4mYEQWojsyB/UTxzbxeEvKOPQjZOj9HbBLV55giTRqmXR+2VQesNBBa2rat
TUA2pSCTkatTzSYbHif8n08c+KWO9X6GStw7aYKxbvNd/PbOTkQN9rBd2ThYzHdqqf/5szu/NbX1
OFuSe82FqsBTBXQAwpMvY1jBKZS7OOy6nOLYIIROdK1WgkB/QOwpsAC0KUceCTOAxggxQbKQy/r+
MYPtn4dT8DLVO3vjvBsTGzpIg/Z7xmYvfYlphvufRD8LO/P9sAqgNXxvHzj3mb4uECgWcfknfp3q
GqiRa9xRfSGU1a4AcHxJclMTFtWSLHlkzfIb/Z/K7qhR7yz0nWEDyHq11ZIsuGN2DNEiVAMbnRBQ
9glvHiko5djJGty8j9pN00BjyqH0aMqrPOyWQk7mtK6XLl2ehdMjOo9g1AKAq5AS7exuRn1cMR4X
491KOoXvNFD5euCOAOeszgIuWuzfEcxLKKqNkywS9hoeL/IBH67b04BZGlK2fwwIwIzWsGtg6tMa
vU8ChRv3yJSRcJAlxo8xi9CtXLZwzgbaPpf5JOvfCpOPFrGjs/+cMCqf9ZlScuaobpwws87rTVVO
PkzlIpJBEWxme4HWS0xaA3b1ka0VL3D0iMroXPgFkRDksHSncj29wiustV297MAriHyK6oL7SsPx
9SxFmoYu/1kAvZX81KCPbeAA/sa7RLAl0Ul0N+2tv7hLea+tEs11XQbuUkdujvyDtSeMMHA6J+6L
0wv5JxKF+EJKnNODQtTSDcKFIeVz3SuFX4itQ93JykWON4tIs6DNiS2/SFcIqGaAWCuOHXWkKO08
+G9ft8HgkDsz/EX9LZqfXJKLtfMlRHUZuO2hhUNsgXZlXhciBWg7uRgIOHQ/dqT6xfbzZDOuo8xc
sB7j/FdrpdMWsUR7YT8zmUVlDDVfG3Zb/i4phkwEAi0zFlbkUi/nZIMZc920bdghn+sntUJTH697
nXcGdECX43vDSk+M1+OYKnbRHSVRywjwLEjzVy7kb766Cb+1qRQZDZ/dHEiOCczqAzG9d0DoNbrh
6IuXPkyG/y7dWyUSehYj12QYIQjDORI6Mmp3ZSO9wo4mroHEUNuM/2kHJOq91+ivEQA6iRo2oc9G
Jt3e8pysFcudvAs53UMf+ytvjJMY6JDpKqyn3MgHAhKJw8sDxhAOtW+tmC7yK6qKU3o3g6ktZdad
9ceduYzLjx7u46SAs6m0TWqfhaN1dHX1C0G7M+6jtIixk32TbBI6UlM+NGpI/Xjvunjcwj58BmjN
f/0ZU7Ra1itFn7pGyi134YWSHo2nXfGWK0Zhd3G9/ES8Ui1rugmjYy3MjMIL14BqS194VdUYaWOk
0sTVeg7V0WJGC9Io5dbKF7WL9F5Bznrwenrcn3CvCj/SEr052O0vG9PUUtVXKEjqyQVtPbXh6aUh
JDTSJNBjTP9dl3h/JnZSVA1lX/CkgUlv5USqevK2KlHrmuz/XMA/TjYOKwOw40ybQnamJH3OveX1
duq9TaXNVDZW1ClkHkV+Ep5EsLL1eUlwMCy4qcqr4K9I5nz4AXedvCfCJgqJIDwH2720S5ax79Z7
a0UqMqaOlj+TRGiX/LUOjn4zd9bouuEteBzQrvs02UxOe3fNW0+j2NqarQZC+0tYR/561hOE+tZb
VUMqLB584ECVlewGHHaoQmtq8WfHRTuzT+92Clfp4xPjoOlRRyAho8BRCWX1fcrbA3yt8TfQ+WuQ
Z5Vicv+GVj0ktPOLz6Y3ExG0PjQSLQOMnAxBp1QYGWYLMgxvPhe7IGadk+CTlvDQ76OagXmKD2lS
yjcoFTgQkhTN8OR87kGEbdY+/fyJsZovHFgNJ47Od9x0eYfR4YlqOC+0LXpixTueXaWgjGV/Kk2F
+aT0pyhkogj05Fe3W8FMAhDJ6bi9ncSKnXtk1PO+TLMnw1ruuyH0nd7lB5ccPyJ8Cp4TLWQJhT+O
ym7hZ9PvTRhzjOQ64r8oztWLcYVpKlshcttwtDG0XwHlQXFnYzkNJMVGGFakCnv5eVZ67jJfTVeH
F0LVeETtoA/OaOoi8/QDzi9qyJPk5hC02IUyvlgpRSt0YgR7jeE22Xi0sG/O36sJPoqutHHmQ/BO
KCeCO1+YZYQCnQLDvUYRReh8Y9kRhNrYxqlr7pWe/0cJIg4RnswdNwq74MZjTB1tuHw3AoGC+qVj
85VYjWkVpWjCAINBXy4iSZYMsEi4d6/ozduxp8DolHcqKLqpTErkUxZSPQ9X8KTJhzwi0JI6yKCj
UVKB0TVmxAD+Y2xOMTZ1SqP22QK3sNx9KMUZm2NBUREgoug53LKb9Zw9jzZcG8/xpr4v+nS8dpwA
9Pku6BzlfGS9B7l3y+i/zAI6mb7KHLjQaX6/dtveHnew5LBAMgpP0Aw9FmhgTroYW7sxj3JB9QTH
YvYdIBL/ZhJf4ZoUHtkNL5AdQeQtjfEkJ2nH0Bcnom7CXmbKEOnmWyu9FyfUGv3HsIBs3jtaNOE9
QG3goUKVDzJt6dgvu/3EZGhgU+5iFMXGJ900NO7vl7XBl6ylB+09CSnmJ++ZDWlC4YSvw5hzXnxe
CbIXqZHSB77uvJszM/9KXbO5McDsh5U5s/+g5JSBLZy8vgmaJ6UN7ydQvuuI7/qX2AztXp7FAbVh
LygW4Ga6ZIrjn9bZX5hqSLLqs+YiwP1BwCMGYqatQcuDLuhzHDOgk9ODhyDc7zFk6UlJASVT6eB/
XAEWh2IAhp6RCv6ANtMLFUpaG07YUdSsR+JotNYrRRGBQztYLhskd9Tod6FCAj5tq4vzkR70FDrX
wyZYOW3BxdaRkTtJu5MwKrH/rNQlawlnNRFFsVwlwm1evb8n9JL7uqEMg+KQ8deZFv2e5y4fmqan
FXM7fc36eH6CClVootGIiAuBtWjbECFX2OJNXS36owyXFOaSSI+OtW3wjoPKVJKJluZSgJW2q3uO
EPqoLxt+GEXLMzFWiUyuunCv3GUgCdKbh7rzzVEiYwt5JrB5H+pmBDeOxyKCa19u9UBC95w6kEaD
I8LPp2OKG92sA/tshsswcjkQcl5yJMf42Amzo7Kip57+lwiMJG9KSv+Yqv315Or3HCJ9NrSLHHan
hcKscgTduTwnJXe7ERe6+SKr652RH+eUgqiheanwrv2VXOTwsMSLlJGAdHCPCUd7VZVLpKWjhl0T
9zy675LgMgEbRWkKbierpV2QeB2T6Y6DqV99ipFVDJfX5/oqg3ycVLsQklzD26Ckxyv5LnNi228q
AqZJCycq5eryRRB5aiT79TUBiVNQg3prV2YuKjZ4OOjEX+XhyP9DYgS0J+rKHVNKmOVh3kgDptRq
l3qv+ro9Uuo6Rienq2U/LTfFK1yxVthXtXcUOw9Q7JA7Gvm4ggx5HgDqgoo/elTGArN4PgtGZ15Z
z0SQ4ayybJ7qn8IRtD1C1ahDqgO7PDieK+g79Co2hBiA7232K1zpRrTUwm4k10zzwWP0xrLfSTEW
cVmVJ6ZqQ1fzL3eC8Gu8SSP3hyKKcFzw3ART7m6sRyWgy7fXzh1FdZ1nyRhP52ES2uGl/xexVQkb
BV51nesT8xZyYDKxtw7TWe0EsDT4IFA/VxHMNp24EoyZ1ekQF1Ffe9SFHd/Q/je1P40hT+vwfW80
fMjQI4R9S2G17+EMRJpYAICd7XyjAADmYI+ivAwFb1Jh58FjM799rDX9VMc2Mz+9RVb9ICKilAY4
qYRomynavooe5DjBqPaUyLMbOXWbGdWZUEy61Kc+eEZnyLMKShBhdzzeGKIAbh3r89O0J+LTri6Q
QABE5DhX+YRnq0YYLV6TmE0fz9DCIJ62MJRRht1WG+Cp/E6pTJlpjK/VUF0JkfUVfLroaeUsdDrP
3HIlJxPKnTqL+iuZGuKfOC296DUvgYbgVUQyp0qt65KAt65B8743BjGEwtL5epb2FvybJoejuep6
srjXNzoJjJzOxXNmOeauMv6ziLKcb7ghTDn7muiRBeq0JmGVVdT66jXt8S3CQhKGSqp7abEy4P0W
QJ03YRMg8XP7PCtiH30sCeCBJ7uclxrfW+VXSZdvj4iC25xs9WEc3zVYBn3PsjIDbbpK8GMKGM7f
x1loXS6o7vN/IFQUEXW4Dj917fT+n16v5auB6IgbiMIxXI2n7iAQiOvya0BaoqWtVrnFWt2um3Dp
jrdLTXt6h4QYAkh90ewsisHfUYb9CIAnRQLRsQqF7RKWWqxG3x8h/M9MvLb3PY7jA7axeogENLRd
BXGiI7PvnsCoyGMiKgPoGLBCfGkNSEG/BxrRTIBtyEf3iwhivE3rDTP5vlz1E+GyB/xvJe0A3+bJ
e2+2XHyhC6uYYaumVIei+YmY/PTPRw9SeRYTZRwA+1KGU5vgFgP/b26akCgMxchFAGbjpBdFi/kN
/tbde+IgVb2IBTvR9ooa7un6fzF2Y7/uU1WkYUdGi9hA9cBfkTFyJo+3tP4E7akvAWICF6Ss9inM
cw7eqhvs5HOq7eBMztBMySy9RTsJ6hUJPN2/yqRP+u2FihlkHXj9HbgczoYtdLB8rCCVyCK+/hj7
j63QmDMqn4wzGD7hH1rnBnDprQumgSAZLV6fC9LjqO3IsZaBabJmo5fBz2rL5Kab69VlBethyxl1
5/otqZzT84urgdMf77TccjrFIjX81WIO1IzdaKAvHV2rB/RufcbnJ+COCfO0GNKF3t5NIrCJigXG
0NfSN66SzJrIh4GnmtUO22oKjgeoLh49ETzy3jWPTgTdH+PhlC9YL/0bgyLlhkfbp7j7f+2jvfP4
9beIm31e+J/CQC0fUHOwMXjDqkJ8JrnvnbHFez3JNSzFxm+3n0ut/Jr4WAxFIHrDdU6vmAGy7HDG
LIw97s47WeDDCcfeDDSXAjNUb8gk7GxFJqyu/2SxK7Nmep6KjqJ9/F5LYwNdFt/neoE4LB4XxQ/2
MHCjOQZl2S8yh4HlDME+50Gu28vGQoKhb9j4g9bYu+uPq9FeA0LNFXsFWX1JheCAYG5WXoBHEMBs
fgvINvP9eEty4F77Dwlx7ESVkBZUvb/TyaNr+9WugolYm5PCqTuVPbvt6chjIypeLd+8FHSbQAQI
BEwtW91lrZNgIUBJKLInCvA8HcifjWq7itdXxoyUKc2IUi0ZJ+hKoSjaa0WZnGNcJA80mYnplS9A
BFNnhNPGadp7F6M8r88Du9NLz6UbmGKmiwZcZN856oFXeL4Z7zh31b9i2p+7PjNj6Uketouz30eT
FD7Cih3kzTX7tyrEJ3b4HiQNjsa3RlRDgAPgy4u0UB+h3B2H/5IloXf2ofH+Audfy97KU+8ZiX/X
knBDN7Uv7GNZN3SiZTQvynj+BuyBo5AqkI3+C5GIkTdxD91ExmTQ/5OgcZUYgpK2fRHm8lYwB6Yc
gNpAirMRiMtxOn6iA/pfVbaVIjv8C34SWiKEeLVoBU7sG3BfwGrPLlR95CFLg5FIEhLMMS7JB8fE
zqPKKWIcnKZinDdU7C/J4ymCRqPWof/rqeyhyq5UlUDdzdjXwBDaVXs9hm7HP84wHr88XCgl1Ilf
rbt/752bMZpR6vfq7vyfzpfTxP/cMzY97yXYBDHIWrRkCv7SmOOf97CjswYoDrU8UFyJwztoczUC
0Mr9YO8TAHelYegHX+Mole7h3OQEgdekRqL9adDbIXi/r61yFKLZ/F6rblSMPTXF+LoomRVoR/KJ
gmVTppXxB1WoKVfV5PW0oBgyoF8n0tRnbmqX2sZTfkbMVHHK8Sq21mm9F2JUrMs0OwpK21MNpCRN
JA1o09T/mJNt6+Ab2dcsSTO5gtAyUq2wP7RAj5kw0xWN7vT6yfR5/z+8ES8TfUQ5ko7jDns8UBEX
hMwuyt67dSs0zIEasvZCj5Rwd5xkefhb0OCPrNCr3X81nWC3vnJQ0mma6C1rTRyODYiV88n7W3iW
hHkHWfB3UaZF0rSlWl2b03q7rciSeIVQPXwQ8SUBqlQnFwtVie0NIUgHmmdkYO01TTi+ei8JnDjO
OMrlFpWeo6v6bGg4BaxAGN9eW3J/scrvmlqbnhhvnyGH741nombGO3WrL/Xs77u8xKRIA6z4ej7g
d6y6B4k3xG0XDksyoGZM8g/hAeAUi0I0bl1DhSLAg47Rj6GQjzcEabUTPcdIQ4y7w4MqNE12a6Zn
o3e5sWuWDOKEAG3TM7ine+blX/Kn3lnODkPxBLO1uuKtZR9kKndiJteRLq0EXTJBRSJE3wkJGcR6
Mpm+08ad8rZ7akFFvPngrLQnH3qwP/OP9GWs7TjhK1erI7+Lt+x3Yi8zg5aBO/F2CD0Hbf3IzTOh
Q9gDx993OySyg5dYSZz+Hcvfpmw3aZIRYnltmwnVb87y3s+3O0R0rvCBpkT65DyONdKLvdkChz/9
AUeDiXFc4CCklJIW6pm7Hks79HtG88qWWlCr7YS3oX+iSMZKgysEpiNsC+i2tJOkZQvp4qbRtqTG
EHN0SxMka7B9mHTuAeombDHIK1lmbwfwHfJIfiNFVzVTBs4jfcPY+gn/OPypeFYQLfcPb7fdSOu+
S2TRrYVJrU14Ga/flJtYFrXBHk11b5o1zXHk8lUv5vJsNyxDoM/B+rjpS7gRhsnEj/R85cjJGcki
Q7V61P+Rz6W5aF/Dtv8PwVquqgRl4W/90+Ye2ap0ojOywzim6aUTQvf2+MaZ744iwUyz2EmM8PL9
oqmEJ6DYLHWUHbagKlLn29D+GbOPJ641kfTJIp2UI4mRbKA7pjj9mivPHNQy6SRZjBhAxvJ+5u5N
RdWRM6TZSG1CHcG9usFsN3jBoI846pAsisytixcV5/YNnodU8AH4JZw/BJP7dey49UDzd3vC37RD
Zmecdxqk5RlzkGd2VY4gxa4hKVwy2OkzJX4CnEvmAkMXjIzJMg2gcWJnjNkkz8+mSKqioru8vb/3
oPSmvSibd8WwQncce/yMr1nXjb7sWnls1yiMFmRr/NQoD7laBGPckmDbEjAMcMYZtCb5h+xgckc9
8ebLg2Fb/z2Rp4dlWGIU6FumtT9ojPHVcp90F2/pPKlmNlV/CxOgnb+ZDhoQStLS6krwtAE6GMea
7z0rtKVu2zldMUAZUZNUGMgQaz0krwORG1HxJV7xi/XWpZ8dIElGyYEaOhZRVYuqY5HH6eKQunAq
kcPffg2xTDVJCQcnLeVnmnxXgB0KzhTkLtrY8iCqPUcXXhiw7PHUWjmRyZif6rRcdOv1rZS/63JD
FNzU647ZTnA7u4M5thWLs+TWribVdU3AzlLX2hoo6px2RYd7Y8D4jIp4RzBxtBAehcefBAYjmfr9
tK3jfhY6X461HORjWYKXuCVt9aOtClkXMdf/Cu0a4clTV9DngdO5HzTqFsRDI84uZjx6sSLVu68D
yeJEOOauoP3HPTxyAcr5kgidbC/RdiuA2i+j9b1X5nLG26p9pqQlQVkwUoiNSWimbl8CJfiiizqJ
8DqESd5QRT2LT9ND3CSJdBG+ONfQDjPL1dvWBeBERlESfYWCE+pO+VhvCNYZJWsy0jRZa4iu8STl
R1PRMsfQfOlsG6vKrfXk2a+gFQDs1eRhgZ6BwaQ5FetQ2TdpNiTMuaWWBu9uqLKZUQyziU035dT2
dHkaHEzOBuicwwuNME7nh/IEOVMfNV5wkWKLlaPFvCOVANn37bRB19KRxyfmSB+fS4KC31cJlZlN
Vcnb8EaTmIRfJ4fI7vFlWakVsJ+V5KwDPNLEf1xCEiglw094UWNK890Dzv9hLY1qyVaoB+FP/0JX
kPsd9+r7cfp2WVEf/DSOVNAs1DZrDuRY1hCckxG8hP4TtUbt8zH8qUeKDXV6Zf+49l0uonC0VYPb
qZGf7kMug1lhY8A8OFx0igeI8UBbttVOiZENbNyy9WbY5Qfs2eHASVvcNA6/kJUvnFlbastsRxz9
y5VwSXZ9N9m+e2f387cmDfgvGCSgj3ZQOy4H6z0/OQ2PWDezvkPi33a09ODDxfzrLDX2qNYM2gYx
MBkr7yceRrZN3gz0HL2YwuxS2+lfCTBvPxXIq6UX29RLMWJzhSx2VQtRNw3QHGbE9XWOhneWquOI
cqlnVgKhsVZEjFSyGjK36+XaPLKZW1M5oaGJ74N3xLp8HpHnnJLmU38pn8Z9zGz6pe8nQqxOr/hC
5ExNr/yBqGTwrETjZSIBW0n8uAx4lLAnQUXj50rqlirjj9meTu0ym4FgpwF8I/mXtkk7ARXFd3ru
p0XYRjZSC2ChaUC5dlwW5LtI5/eGl9f/1sy5zmfirNBE193dcxDiVVRMUpkldzKm9J+H3FvJhcDI
orAc7gyWHSbNtXrZd4FUrMOGIdl0XZtzx6DayTwidO9QqNV4Qy/aEeejR0Z9g0Unjt0uXkkVtmhb
8i3Uk1tFoauq107S5IOlOAex0ciQMibzpewfQ6YA6WZV5GjGCAHiIvctg1tnfKlHwYNCFpY4WSn+
5g6tD524qt5QtSn5vp/bUzFb/hqQTNXHgqOl3omLW2kiHDSZUh4sys2xt3ER87i8iUFiqx2ATJhn
WEV4+YYhTRUcYP/9MS4mQi5Y/WC1GkSWRSLesllqpvhv0CBfYVjL6ZPIgeWynh1nOYLdjNRwQ+E4
cC6eYJo6TEgglONfvnvOvG9N1i8xO4qwoMQ9H4jCZz6drrvxsXO/+6oaDG+pLz8/WhUWS81fKCEO
+o5wufJ7k2xE5I0AsdJq+gfDQtpaompMod/yMhJJCbpHlWprZrWz0eL8aaLhqJVCrFHZaOj+QurI
+/9BR8lMhLKfdqrbwKilEpz8mSokJ+NSmOXFCnkU40R/TJ4mIaCxn1WOm8i36ZH4uwFAj7hnQPw+
ZzcUeim5D7r2Q3yMcsQHlKrATpAyDIfa/oZG74rcINvBsU/f6oDpiKxGNtDA9xb5F1TFkvB241Uo
eFRYSJ0qEN9Rw6bvLYMgTCSELMb7hvBRssq8VoeISgD3y1zxWEzhlHP7Dd3+2es5cSAPe6qqFC+O
tJNL+aQQ85+hNJ86zFrhC2kj2MGUThQUKR5Sczril3M4LDBh2T96fe5nt32f3rpigabP2Tvh/po/
jJ59iD9nJ5UtnC2ED/R/qE9y+KvouPGBvkvK2IGAktFPXOked2nYzQEQ+kCpkIbeTProbgIZLf21
wqHe9CHrYspJjF9iwb/SMxNzq7kBtSMl1OYu9T2wL7SuSEFMb3VXpU3wRnKrUjvjccq2GFGHx0yd
ArKsPWg3TLnORmKXKfnkkBY8aHqx6nBHJ0v6xaUEePPe1Gs184ZpZrPbAqJYhxzclPxgFRLXFZmF
x4RdyP4bjI0OmEA5LwLACwZUmMEMlZG3cpHG8kvLB31O6ybhKEHAenhqI8lRTPVfqVnJq6qpan8p
Bmd9G5x5awmHzASmZYh8xAU8oCAIFq5GtowAiplOZPHq2w2hS+dwqgGTDOQoOXLHxBasjIxNKfyQ
kssIpofCIUd3PDB6K3ZWD50F1UdHP8UH6XCPjhbVwZGS4zxZ3+BpMDZBffFMJvvd3FLyKzQEe202
5YDk8sqXO7k1bv23q5UCWkN1wp/regV2u4iHxZkOwDeNXRkqkVNmvnYIdD4U0tRbY36l75HeHOjT
xLAb1ELh5hprK0TlFUuYMexu8xS43datOMB4KHazohOS6fj47yrTuCN80OWI5sW5K6sh7RZC/YNC
q9xlNA0nopWNZgSgBKLzzFaEAlOk8E6dXG5MTjDD4bSr3eikS6lV3WsOykFFhudIGGTvyLmakpdo
GB9yz0Yp5y76tM9o3zPKZ5mZ22z88IyhxQYv85TNP5dNh0a9brlRRmjnOlw2X2djb/HPewTUNQid
7gaMHjZdiOqWgZA2uZUgbtSGMFCRYHralPjBOYn+zIQwWmxCeNdoqGyb7EWqj72c97LaYWUG8JeN
vRyVx/yAOl1otXmsB/GnI5woYWLJI6YXVRdLhROKBHY4nnaA7Oeos2O9Xi2zHAtNvzKjEDc/8szC
FvZ9utz5TAzWti712K4YXxo02tsxfmRdiu3OHPTYUx6+HUCc4DoHJ2AoPXawT4n1oyzr8fXcfCa8
RtYMheTu81GJH/6opxKOqSHHQyUTAVjRnL/OKv0C8pyVO4Ti2pZHEZDuuCHxd39YLYfQ72dVidEg
vyXMOxKWRqsp3eFV5mFGQm0Pkt/gPZsEPVLzdqA6D77Gt14/1AK1rEH/anoTsQx+Tp5xeGHfD3wU
/LbIdr7gaalh3HIqCEdLoXj+bfREEwAPG54ngVzLwkqQpnyzwXkgCFtdiLhrkzGWdCOcSJ6dKXKs
YLrD35/UPorDLOT2kMtp2vlejn8gSWOrdVKfO8BZ21SPC8T6zsfdNElUffn7m9xQlTFG7sLKZu5I
We+BPADVnFMWbEsdCj9zxAlcIjcmeWwDIpvrDSQNeVpZi3Jk47RjlHej5R6dEiCwu8TPpv4O32/V
b6cTfmSI9IvxivxWS3BHtnDOk4XD06l6HE5hFBHo+DT0oIV+gmpPqOQwstCQFDH0QXeGvZ9wj/bz
TVJb+vrdG1FY+cqJH+YPxOuWGCMe400XrnrfoIfiKIV7GQAPT6/YehUjRPc7QytCLSj4HOc+1pag
geR8S4bWmybWngDS9nid4+Ongum2kr6HC9K7Po2dyHPRY+6qEi/UtIUCm4ui0bwcBMHrWN6ejQAJ
vmqqCyOdaol8avsAjfZo4mwLDWrx0MfQhTFyuvybVXqq0z7/sxUcNqIs9eHguNz4aGSr2S7PXrhB
niRq7nNy+u9rURMjeN2WCmTvmes/NuejSARNw2ikRnd85FJgszfLowtoDp4Ecxk2dwYv3Q/98i7b
s9R7gQH5PwgFW78qhPQrePKGmczhtb5gkTAM3R67Y8daQl8lhRrRSLUtJYan1pY8O3GQDdSCCckm
q6aJVDRgVdo1g3PNevR6dU0poImX02JpALzbkA19e0wrC8saxuaiYDLHWHQPIjVw5O2UuIwhtJLK
38hVz5YUCQkwOxX1yPdeoMbRPbHm+qnYKOg6/92Vt2/7GaIn6dN0ptGo2isKi3K+6geGc2XUe8dy
Lx3cmKsUFdDXT9ndZofJUepstzRiiYaJ+yiaZrVrcb/pyDNJkeInzMkMh0GfHqLjiCthxl2yPDl7
8kWR0spQN8f1auWjIAdfqS5Iwc8cZ5h8SFiJ1K4RY9qbsxJ3rF/5Eshp34KrI9EXJXeRozoCtQzW
LmRUFwmA1ksNwaoI4EwquLwju1hhu9yqe/gFf2qskljvVpaFtdGGWDNsDns+LhMkAQzgZV5c5xOP
haxlIUv/DFukwDKCGR0WndHBHkVnB6Riw0Fa4bkOoCmXY32TDU9Xg5RPhqP4DRaQDc7cXn7v3EyB
hJlB6KK+jvn4qHa55Ocd9DCUwuG1fLZS/UZf7eKhyxt6z4ODMbjvx+gJzX06H4fgAchRH1V7zq7G
EYcjJqfS+tcUNr6AeTKoBWgoq2J41fB6im9sH77eOnRCL7D8OWqbOJXEhpyOrtDwDq88WSDdnvJr
SI5YtNpbaWnc/ajCXLtiCg7NmB0o5rIEAx+h0BEm+ecsrqzrjlb+xnhuGSvNOnw8CiaD5T0sxJBl
M0XNBfE1aFjs2uauSxdurpR2SpNHSw51Ozw+/dh3NhvtSxFNC9H9dpjSHf4zihRXlevpzdwMx1Tr
MdY/mY8yvHphPHaBYQaSHvWxEdYfK/N2pEjYszIXiU06CXCe/0XNEPObTRMrNnVV+9TsHrCen4z1
0tAYiLcC45M/+WD3f0e8C96i9aYqFIudjsfwEFa4uZWnj2m5dqAwY7gCoGoHqM6Jvcz0pQ0lC5Iv
W7GsWyI2CBfrCaCQYF7jN0xIwuKDF8qdqrfv9X8DiknuqRwuJmeDklQklb6qWe6IqClIxEj5G5QQ
Z76Hbv40Oto7i/i84J7Hf+HkfNzREa8JVEFmOUFZ2wkriw8lV7bo/IUwVTkpZwLD4iP/JJnF+Tcv
KcGMPFdgpmDiYu9FfZeSIF2Q08ygs6H4+XShtJ13qy1XRZGtUhSrhjVZuke2jeDKG49v+d2o+o4d
ZKUjwakw4tENSieqG/vH6It0SQ5c/8E1kvlqq534CpZlG7GrxjZxfclapACn39ZVrLz1EUQtgulK
l4gj6AGqLVXW5aT01W15JiKtCHR1gYuaemtiByY3NULFyodM7UFO+eoBX+AOLKXU59js3S6eBE5c
0cANpo29RDd/ZeK+9dTKW8KZ05CRwmO81q/V7xQwWlXcE8yBi71Aty13TQiuNOVOLhITp4mkZkON
yTfTilcUJKVKJY7bLjLg9v76YgZjXkjZvHjtuQxN5Qw7nolJb1WfbwSsbRuiVKNGFikH67+g5y08
4ZRfSZeZdJjRGG3QiFH1G3IjUsdtRcLLF4JltaV74tbq4TRa9DH6ERYNQCxnXg8AVWC53dMDu/JD
tSdzJNzG56+JArZaJ/R/SnJzyWVf0JGnXlefMypvg8ShGJKxkAPJnrmf1mOc2BDDPMt6HOt7jUy9
RoxrvGWQfUOTF49Vir1/ey0/fPosrvHpNcvNfRlvEoeg4eULxvh/+zb0sXEgbIguI5fcq6qGA1kW
qAhPQ372Pz6XhesCVT1i9bJuOGETGV6kkFZ2BXy6u2Jamh6ORH14QTZI+74yPKkqy9QRrZIzMlQI
M9uoy1HAO21IOWAnEZbYRA2bujQ2E2FctsV1BWkTxvWGx5oy2qMC/xjpI9wb0tmCo8YPN4jyXHl6
c4DYXm8eIiVwC0K42jteN58mxPIV01Q2Z3gyzH3mY+YF7xPljN+8zf4l/VMGDcwneKFPxDGbQ3o3
OshiZlpqtdYceNI7h0lICovPP1AcnwWa8BV2B5nuNjvWnfvT+//5jS5RN8nlEEAseLlb5ssvLmSO
Fuch4i4Fetl887tLmX3z7JkwWiI2hRy/9JtIBq4DtiBGJgfgEE193s8LptrgO4H7AWiD7msNDm7q
ohjfARIaYPcMuqWV8HTHtOArQtjJG2UI6dhde8vSZ/sB6Hh748uH5D4cchiK+WGdibZ+Kzzx/oQZ
6F/dRwnQjZl17VeU8hzLiohZMuaxKXnpWLRga9SiX5xcxCBV2B0SUiyiLzLdtOCvyttwQ0ShbWA/
6MuLeIRVJvQCwtjSYCTjRQUzYBVX2ex6o60dih92A9AzwBuFHXoGaeSfD3MkjUzbOo5CBONVHQU6
HGapFKy88hK2pMQd9icbsyMkD+++dg09Jg6oKcJZji2/UohgOZSgfMFYE1CrkXFFP1pVuVZsGZSy
ShxD6Qtpo0BlYiS5f84oaYRCh71USqi705sG/CpUCpyf1rQ39I4EQgRw342RGBmmCHwKG8bw9iVf
z0IKxo0n2UeXzecZPfS8YWkEz3iSFcMK61V9b9Vzd+XdkQZRdyosnUl/OZJuppU3zRaOMx2UciqT
PYhf46MfT2mjg5SO5zS1ga4dFgRcdjc60DJQI/0dOvl2Rf2STcV516Hxg0Cz9f6o421kHD1XUCTV
HoTas+ZjZ3v4Iqhys8RLE1udY7lG8UE5waIM/NkPM15neL62Nwn4AeUBNrftBe86QFZJZATooQhl
Q1ZFDAP9J8HWQqnZBfFI+V6ooJtdq2T4c5IZXMnmyeSqeLTVa5KV2QMCEuW7Rfv1xT1cQprLjYWo
4DiIEI95svWVpi/XwvshPcPMWDSnSj7qezH0Sut2yZdjys6DBKVwD3Kv0lW77WvTdRo7rzxMQUZl
JVxpqtozYloaoMieVHKg6eNVGaguHWGzBVSEAN/OXqVIt0oCmCISq0tXeW7fRctu0wyMF+Oorj/x
v0pbWi72JvxULqClWnHoIvQYugEr8NyaEuhF0FAwYQVKrVganFMDHgW4nRB4cgVK9hiLbO71BvQn
s0HVcb2elmnG/6Q7WUVlN13/d2/kD1GuHPGW+LhoVmIc+62bojqZy3XAjjDXOsEGjtToxzIGl26/
Cgr4mIq98CCd9m48K2/xw52ofyEm0l1rtSW+EMUq7MeGtQZeFXSplOvOj07xBHBCJhHS2cHwp7C7
I9FHQ48uLKHHir4RsRo/YM+vTj9XfpGf1n46MAR+Vk41J+YhhOhBF6H8PJKdzy7ypDQ905lyKIqq
GxQLxnaIlp+wOupXfY4FbD0SJQ+ak1zkb4AypWxSumDZ5auXeXPcc9sw30+/77kVi8g91wmLrFxk
uXGNufAy/Jt81MCTo2m50DVLhM5PufZNYIXSHPMdeZ0wlFDmxsYU6f88QE0LO2sKVoAIEXG6ou/Y
swwzIK201+WIZBW0XotXa/cZlJPd0b5RoVXYHg2lu70efMObZGlkz3XB1Qw9Wgx76UN8KQt6NEv0
6PovLXUpQSG3elht/YYIQ5P1UY1HuQecuS9ueG/i2wpGMXVuqN2KULpRiJU6kJljqdVJTGak8qCV
eKojBbdK8pfv+h+FCQPieOg9lam1hNFb2KYyIOPsIxk9CdtMYt/t5pWyHCMxc57fY0c8cI3gV5Mt
808ALcXhOkaf1TG0+eEcIT3CtZ74vuQ9SdWJyjDMD9rgjbDaS4BrfmKCcAyoUhRoCreNUtJC4/wL
JjTJ+HxPWqj+x6bdF+mMf9F/lgdvQUn6d7rZF6bwAo7ivetDaommDdgJ5ViAoa8e4Ri0pN1zcz06
4m7/8Aa5rN8jNTaqZI0g1RZpGD/T+ApTsbD9tIkpti8u+RNw5WgdCMHkE8xLdwOFNUGADw60Ov+8
JqiigCEspfZCSzNOhrgyNzlTPk0kjq2hdEOI6L9yL+cXisDb0uSu1e7w17DMj9RbEziUQG0BibEx
9fVxDzT+qryrs7pLfEjInLzP2blN3bYNDNeWjd5xU7ZkfTYq/UoYKLV1S5qhbMkQW6Z1mWTqMoBl
R/JEw3YdZu5OdKKO+g8B6nwCXXMmLUVjQeSHs3g0xPdlqEiF4e0DvFDkuv6r07jRG6LgnM5XeY7w
+mEOuBXHtBE9ORWCv9JTVW5pEfcj+KxRrdy2wnLQAI9XwdsCRPWJ1V4YcIcEDXEVJ9iRRwnqs5DN
6Q2/1cSaXF3fLyFI26rv36DWlvWbrLgiQShnCH7bqJliz3TvGAsv6uluxauV+biiwVR9YwdNxR8k
xDulMaGfOAcMbcieo+MhMlzw7T22TLXVVK4fpFEVUqjRjIIgye6ym/YjFKalLUIitt8IQsiksce9
pZTjxU7bPe8149VS9GcLHBQmu6TDlR1xPDElFE7Yma/Q0MrR9ahWMxLqLT20jCfYjs4CF5s9mPNa
shk1vowqnfkeBvjx9keBSsZkzYQ6TuokgBwn9gCgA3VO3qIU5SXrliU7JWvw2QJ0l8trkCV/91yE
6sDfe8b9NchpenpV4hpx5GImyhBkDdktse8Y0nAd93g596U2yL7pHyhP9Nwrx8rFqausSxBrdR6I
2Ke65pW2U75A5Iqwqd/7/BYJ0JNU0ryCc8K4T7UUd4a1v6CuhWUOeYEtQofwx4IHt2Myts9oUi2k
JAdMTP2ufj2PEShiJxpNGecORob1xuxPTfMxpfzkY8fU2Bs3sA12tMOE2x0q36XYj8Tp9sgt3MpU
wV2l67SwckNPH3O81AAoiM0D7Ki+hUMTUWkv1mJ2bS+YWjFTdHdvmEBoV/Rwzvc7v+VruQ0wzNro
Dy0h+Vwe7091v+OXX7IfcRMuKnKsOdTTF2nELlE1Dk+gfcpHCVMxjzTfB3DGe9tKpezCpumwEqpO
Q6EBBS2LPBEkB1D+1cCshErVpvFOhQE53cSQsr40fHYiyKbJJcO2oG6zzLMutLiYBg7zOrUcSt9y
b3Ik/9cCx9vfENeJY6z84z7orMoNTJNV7VIDfGXQB16d0t7YDAggjJrqh0aXZVy37OpOolpKaGRf
oYj+j2nZF7YwZZpAvH/anh5eYKJ3E4+kJ6Pvb7Tu3peK6/lOJVdqqnWrC6I86qQL/uTEQ40dZT9g
0EGn7uzSSZZjhQ8hD04Llr/N/MbsOZ5o9Cq8FQ7j5fwWLLF39HVgE43DoJWNaLiQCDbPeyQ9bZg/
b4oL9cCY6GE//2+lk7sM0WCKaAL+M3KAaMESC/Hn0wFS0pO1a3LUJq1aw+bZbQk3FRlMH4hxFTd+
62WIs6Y/mARswxl1tkZYWZzoJt2q9/doNp28cy2/dVtx5iLTXvUTjf1fnDdKzix+Aq+tap6Rm2Fu
f0iTXo26KNwUrT/doV2choMo5S3lACPUqeNjJo2N8tUhwC//bmXAaWsh3iexssNWWGjfiraTCy4E
3SqfKv/NbCSnGZWktnWKSOiAbPT0L74Rk9tLlmIFGfwtnzysHk0uGuCsPPQRwxgTP6F/SuyrBYFX
hOjp/h9AUnx3FrUTXlNCIkonrInqGf9vcaxLn+b79w2yCEHljY3z8HxyXHVJO9jzGGMw6pn0GAkE
nfgUym22p9aiwndqlXQyCBDwGGLZltxvYne+pk7PAGuECYAKbiYormrq1tzAI6x5/HJ+ucX54cl+
sNptkjQcVkkpmSdNjwz2TmbQE/B/BNWrCcu4hBNPjbKiNFGXBmmw/VQg0FZr/zmZSJsJb/7oqdOl
RXCjneAz8qt5mo340bY/zyuoU2685zqq1khZSgB3OeFrvurfRXckOE3BHdbcCSIJKWh8VdON/prT
wu9jbs1Dzujk8jKtfhLL01cfkO3dwuCibAU33f1Jub2+2tJ1Me90nUyCyWPkk8XZoBsnUxsouvGh
vGhT6fKTCH5uyAwDw8o2H+INtF+YQMVcCUvgQ+wLN2/UXkGtbUsHPQ2wMEtOhy1nCkz1sYEYnmqE
uGFYsIJv4cium+uFbbZ0JqS+6ga/jShdpen5s18VseV91QNiZE+enCpUDkHg8ZEx014RHZ8LyoUC
awPDtQOVtkJ1uROVP928Hf7euHoRBwUiRxzvg+hum/l9lUjGzKqyXmgfvQm2gUPsNqw//3o4cjti
2IlA0x7ulUE5f43bmfiXqfd3x0uhSY/xNFxes5VePgf7iRKTa2cUf0CTAPoHzbuLGpFoPHbO8HOU
u8iWD6QHYbyicgbQD3W5Wak/wPIsKzWmgfLezUAgAKLTXuB6OgZIvMePXGaV8ARxGjmwFY0YJJL4
WG8Bw/lgHrNDz5EX6WlaY06v+Xkw3zsW1HqML6g1L7t7zimK/EjWU9OSWHeHjsaIm9b6ZFRqBqgG
2yfTxOiKJnDm58USOCZo5j+21YSYSdus30Fc7VXGsh3ZkIGNa9Ma94itaWfWGSzM2Gv9NKezkCD+
R/0bQsmCbah9EpcWwzP2QM97+dmu2o5SuTgZ5lx+x8csBH/LP46qToZQr5sV3hbWMiDHs3S5B38j
0EX6u482thSbN0EmZBMD7N24EswJ+dkbqadv2/7WjG+5J3otl4eR1+z3++FqNE1KWbb2Yalve3/M
q0t9CKChg1NR0ZEUKykDbD3fzi0bf3DlHJ7l+QIWqsgDYDTwS8PR2kznR6dD5mNTpOBWqphkr/Fn
IQk7XUqFEJwFb0Z3ESHYPF+g2W/HaONYWaMSky3T9B7KRXjaNT8FXPU9mXNUBVaS6MWSHxS9Jft4
DK0hY46gM9HZJXVOcCmXdjuYV1xrGFOzFxGOZ+YXyr9/2Lcsy3WQ2iXpkgRCcdWRLANnroVxOg34
F+c0WdVH/D3W2jTxl0Tx/g58hWpCAQRR4We/z1NIo+KOVPJ5a6d1g+8hjX72r+aJcLjw+02RHHzK
sudqGNzIvCUxm1gRMZVZ6Al17JMVhHWaKH8xdkHBGRydO0CzUSj+6uf3+/fCZacjakTLSln/f4f3
IaB39gie7BTfFGCIyDEcn02xvafX3/Hk5i4EUBR5jMBakx9wnrpVTaFsoWB7ogGz+8MtqzYLoOr7
UpvZvjx8Eza2nFtVKaq/fYPKAc0Vg8sE3UVhVWuI/PLiR0NqRHcuw3rmsV4iRUxZ2HUjgAzRflD1
omNveyzlvQqXR+m8HSXTrDBC/EwAMnGdmTEu58oosM7QXrMQUsD0LaDy1a4dVMCXBzwcNDCYLIC3
XAsHaYpU/vZbe0LHCErwL2+9rjU667JMoE99wpqW0jy8UjNxJDIG9/NeBGEMVEIrsynS+Sc/YiAX
qmi+vu4zty6xIdoObRRBJLXEbt3Cs8aWTCGiqjx3zCCcJzrm2/iZg7XOyFfXo4sIC4Kr17zbWIPl
009kqyTslWlD5IoLtmwc5VpXC6VqjgdxYYVnGfPgPasOtbGxYIEznvy2LiMC9soRyP/JalBdS55u
H+ii3sX8PpxyT4KbzJjLAEt3hieJzDJz45mwDs0zmipO3tz4ouruIl8uIFT3QmF2s3cbRK0m/aqA
6JasK8sahKtZksd/qKc8ZqOPtv+ZpWK07orulpbKrpIy8BUZUP7VngfL1uYHT5Vmadf9dq1CVrra
YgtkHTBDbwVAnND0sps0K6Wwu6l0G3PI/1PBwKeSbXmVtmCvaGbnZ5eLPAKi2mUHp7P71vDGCRhC
XOOdCmg5BsjSeaTeuLz0bNZqauhFkO5iIQeqgyuxPxdtJ0+MXEuW0xlXdg5rfuSu/BzMsnueTaEY
25YQp7SLcJsfUIapcdtG0nH2pjAKiFOpcHenH8k06ZkCVW7Sl+vSxUTGR5GgL4DX4TG7b3Pd8qOQ
Mi6Fvlh0PYhETKYDkegoSZLXlQy9Jf2cJzSLy6ytgDbMgB+aJy0XZXPXS7DGvLF9cGIm01ITuNaf
4ki2whK7+tEnX+Au+p6cBzxZuqLyCbzt96qRqurzy+gzBmY+ZtR1a7igNxgkcEkNPGe2iE0dJqNy
4daXDdolXUipnvNpF66Dk+E8yV4fNfU+zwneLDE4tMOpkZTNwHLoCUOz8Cd/z4JdHbbkSA4SVrYO
PMhCiaG1EY1UkRlz1c7fCkEh4VlvCdit6qDejNqNFEDUImzZne2A26JTtoJ0bc61ILXD+iVze7K+
a/KOvPZ1wPJ9kWaVcnZGEnNZZVSBfDNwXrtiysnUa0QUFmest1Mn13eIr9lb2fIU1ccWUSIOe2Iw
9Yu3Ihio8vpbmcHY3kzj/GSRsHMZZkqW5CYFELkKZdc/UFzoBeAohx5evOFakBHmYFyM62P1HVd4
qkUf5p8sfJ/iYWWJ8+BwhL4G7Ub1Ic3N+XtVpSfFazaIdYssvACt/d7ioS89b9LFhfpqK1qhpGDV
uCyF/ri2WQhMN7FkSFz+QdDP9YfBMmkX3fXG5hjrdEUD10InxiKAvvHXQTSboZtRo0gcw1p+d4eP
uWjwJGLjF8pvz6Td1OlzfHGGH8CeDwPtxwytXEOtJjZgPXZTciRRn1xNqOcQzjJq/tLM17Kfeqka
uZBjWAVMZ5SKHMpKRFmKuir1T8X9NCcNAW1SQz+aX904MOyTaz2cfDhqSvOFIumCZi62YVTWC9Mw
+j3EjBUPZLaC6uMflWIDtYV3yhqufTMYVhPj6WDZrOULj/Szhfr3Qfcwc6gpkkqKJJ9b+OU4s6DT
UAEXrVyuUZ0PvRGAnp/5r2LEX+YNOm2dfFXyXOxjtoUkwjKY4+cJJtnqzGVdGwzP12jTziXPhSeM
OAfAq4FRbh8Uuq/b7t3mylBHZ4WOapsfFgvBMDeowAUcRsmIpd7tyhQJ2AMUtbGT6+vTWiPW/a9r
v4ucdDI3GWHTT1h0XziJTUsJ71SYjDZmNNusRo7I51Xi26KDFt0WEEHE90PUHWLFez34DzzERd6u
7r5sJNmdef0ZwenuJFS0YTTCREgTyz7iv9+6+IPhhJm7gfbjFA1WWDjzNG+nd9TvCK9rCuRGJQwi
UxaZB28qyDsVTkwqRYtlJKRL/1Ouj5UPTmdJOyOQ14Hr5gKO5XhSS7dQmuY928UTyI2ZnkZkxrSy
5Jo+RyNxVFd1bPfaAhLYqFGnz4lVE0O23lZYmkEjMMWa7GU8w1glAexrHbcSwLEk8f0fe8HLiybP
LOYqphtybB5+x2p4YfHMz6r7r4nz3yPP64MR9byMBXfSU/0OsG24eZPeoNncPXSKFIRKhIAuSAWY
Z3NJUJUVwg8ed79w2C1kb8D4JneMfTSJ/rW7arp0rhC1AiPSTzEUr2GWmw4AhwjAf60+Jh8Pzq09
+VkNpMyGLSY9SILZUAuLNFyJ3tKNPDEUM0IJY2xPQ7WWvAqEz4PWWH/ehDUi5Qo1w1eNQqDQ4N3E
eK+LF90iJTyuLqQU7Hw+RKuRMTS1VinPr1krM4sAKLetI6eV8I2/iwj5HgMmWzqgwaFeMmsQmWCP
+2UIhZIRj9TsLO0Ap1l5rmNAHc4XJoB570dnlNX+sLDz/JO8p2/Ap62tYTZlT6DAHw4sg2jVCz4C
mKQB34GylD4JlXTW54NnUytFOzj1YtXDnGqFrSfZ1XFB3XCsQWJUX+Ov/MtcEzjBQ5EsPHFHyIvR
NUiOfGN6j643VZnHL1AhHrAOI78pmZRcweD3iNQO4dFqIFjZlkgRIICG5Nt7TpdlJD11Lg60dx+/
W/8wNy1DKDca/FSUEPPBy4TJEfT5h8IcdAL2VCCl8tSnIutGIUcuq5T/RUZ4ZwSNnzy/ZfHRzANc
3v93kiWxmKdTkM0CMyQI7tD8DBSu7lG34l7wBnJG4Y6bGpKW3Th87BEWAbLlI6y1DhgpBSE94CUs
RuZB3RvS8pwyKnXaOJV+9FY1ddlzQT2uwKVCRLU2MnRypx5ZaMKvclXTkVQ+gzVug/i9918CGosW
8fihwlNfVeTQAIUPXuliLY+f4/1MWCegw21WgYDBEJrjIQVWEsw1m2B6U/5HPXpULi9LA+cFr1vD
sFHaYbJbrudQ5GgCFwEjcpIfIwuAxj/hradOwyQEhwk9ilPpp9fFbAvCujZ2EmIcLsqmI5fO7xab
rrICepAmTUmyv0VLwfYfQnEVnAA+XB0uicohEEQfQ2gFz48rTBg74+LtA0Gn0gfr+EocBd5mKFi9
7h8x10YONOZOlh8hzJslAp2Oeb0I6vPOay/zH90mGTtn8tgAWz7/dm5oOFZiuEB8cUnytpbGJ7md
rJNBkZHOV/0ninlandM6kciOR4hItJzWu1DGvbXKMgzGJmxGh6sMdcF4EKI42L23L4lawcynE1uq
DGjc9aiO8t1AKqpXxTmE2xYdfdjjXr5c5HxvYVbfSN9BPmiKa5LJEeVB3el3j+y3wlZ0NaaxcSw1
LnIopOiZ7rHlq3suxykdElSgakQ1mknH2XGGaRr/EELNORBhF6O1kL9l8Xg9qIPxhjOZxPj+pr3u
U99JRnHHDnt2A05z7Af8KADFiEPZnRSrQhtwbcC0qgFDcxkuS8rtwjeBUUYnYyV1gFuWVnuhSgfU
+S9h5xPGT1CovcpKMAFNpwRH/gV/MnheM2Q//jPCFmGgbETlQaHW8dz3yUmNDjVFjMr74Zh+qvrB
2dSBMAnUxS9dYQFtcNvyyHin57lN6tjYmE2uHh5Jv4YkFT15igwanuQOGLwjKSboO6rOXRRBGn9s
v8W7m/d5F/Oz6aBEoNETOaDEP/PREQcQLTY7Mg/j8RWUBmv93D/g75trmREkLZfo7uuccQ8z9T1n
j1imXJyViQ1gccuOylLfb02vKT948hqhy826poV7cNOJ80oiCcKkL8Ai6xSNipvI08bIgc1uiwVf
l71fFjKZLbmG6kL5lWv47xU54jqjPlTYgFh2lnxwqgXq8N0vy61NUXfDBudICDrI6nfdrOeiZGZ8
xayWUc3UAbvB8O/KGT+5vAN9Ny7Yx0Fwu9iQ2P6OFZ1PaG5TvtvqLxu9yy3TYniknQltRCqmGin/
JCz/iD7KiBCjm3tkVduTZ8n7RgJl9tbpKyFdICz5xCliU3XDMMOD69nZyRsT3E0+EzjIeu9U3Dym
8dW/nipiBPos+kKjemWH2ktaiXu3xJpIP3f7ukyE/Ojl0vgZTxxxa/6BFoWitBW+XtalU+yyUzs3
KXJ8Gt2953sjAjFqYTZOmjDLOYSxgdL7ioBhWhdZezG0NMVkklKzTsfmRnDdWNXzVxdvcUnnvUIJ
LJuUB99PVf+gMcbBlrlh60p+KXVhLZ+3MVdTYT8qFV955Oo90pwJs5UtdLsp9oaemrHvuWrxibn8
J5IfVRRTi4q72j5m9oBCymyZ19YSRxC2OstTDUlQ7bIFHI6dnQwQ6RLvkwR73yILB43vd4lr42eW
bYOSRIn0vFI2l0HPxjZJo3WKty0if/lYmnSbnSligYRTE1CReuyCi/oD9F97txE61NKXONO4ruZQ
VcUeEEEm2nH8OoHKtvMAi30yuzwGnzpGhSwien/yyx2O3ZG7D0u0N7M+77GiJt5aLfl47K8eGa1n
3Ip0dDFY1g7aQhgF6g0yvJPrMOoBG2v/me2FjNp1MHOxI8JSKJEqgGwxJjuVOY1ER9b7i64OzUbO
ueNVeLpVAXLKSFmDFXj9e+OLSG0Ski1ka75sr37faLqXQPsdzyLjpcV4YMaiQnXBsBsjpMmPPbm6
jGnvGf1q3GhS9SgyzbaT6LcHAwwPe+G7+FEB042LJgbfv04CBfqSOx5azylNfJF71e0yF0JMUbu/
7xD3nkbOsM6I3xOEYiie2lSHEJEtNwrs+M6RjOpEjLDS/t6RrJiN1ZW7omvDvEgK6snSmpcDaYuy
a89aOeP2Gv+zPNqRkjHYsFQwyqiHsFrwYSQHjxr5hzCnJwpN1UWCTsvZsRLjuDfcgbsUDrxI1CWE
65ww7kiQvoKEgijEn140q78s+T+5TauGA1+N/E+Nb4AEQOIFq+Es4TeDhV0nHivGnmsT7FrZtYqB
U9N9IgXqQp5ElC55YjikfhT6fEB1J95T+yoWCz8U1+Qx4tm+s0tq9FzLQBL/cqUxTFT7x5eqWuRF
FlyAiCx08mONMPhvlA74pl6R+gJhF+D7YCdoy8lu8r4ZpWNiUNSLf4IJRb16VLUvpMzZCUJSlt1T
vlxj9ZS444FHso3/QlwfU/ZGzxDi4AAIuI/F7/4pUuK7blOf/FnHVoRm/HM/nxzoFHMmeRZD+lU/
FGJ2KuO3xTXPP1vAoVxzQ8lrPAYfxdaCVqy2b1dAOgONb8XqtSW75tMdkCQtgojZ3yR7Z0u3uvIO
+OXHThanyAyNIw9MLGVhKhe0y7gGJ+8rdirdptv3mStm1mkKl40fqweT7p/pv3chgmZJhnfF13Wi
FQaNgDYb2nih60fuzdXQIUdZ08n56jdv/VPf3KyCHfF4Lr0nWgZNc+DBvRJzEdlE23aEZos7kool
bAfRqjxYwDg2FlFfnRFLjUD26BowlB9/Um3TzAvgsbJdtBqlp7niTeTP/9MdACzbsohMRfLfJUoi
0Xn/n4OysTFqViB+j3+hbH9p6MlucrtmPijMLjPHDjFeQ1dsKi/r/V8ohdXHIzp/jgxQY9A7xgKo
CGRjQAvywpjDbZYNSGCddyJuundO6ILZYmVJGhZOrbphONOcH5i5aFTh1abjlG5pxXbptjmqntdU
MLVhbjylc8DnP/UXE29FtOMK8W5B2UKT112EfQn8h66flXp/ZA39VsTbrzFi5gv2x/yYkqY/YzrL
hvywvWfvSplS0Lbxcs6NeEZKJq7RC8PNyrOoW/yj4aDNTeiuGtwtR3pQYYB8tGmqdx1EzeLzJHOL
iQi98khMe6noaFa/TY+hdX0suuNOiyS1hjEmf/FP/qG6IVr9iMeV3992V4nq34+A5UtwTeVRf4JG
5eW/RDBbJ16RQICT0A81b5fJqCcXrUeJViIukBhgyIrqZYE82xWPZKVg+rL3GYXvcdCPVISQrYha
2rxt1pwVXU/PJ+1/f0V/R7NWfZXj6HROmd13gZUEqGQ9J8xIjNVnStT2DGih9aI0Q0gEvaVrMXQw
fuQT8oenTkQlReQE5yfLM9vqoUzhmkzOHChwlM/UGDMRmUkdXz7U5wbDgYu4LoZGAE40o1W8Kl/O
WRV8WZ+cb+la7UPB5L2nMMBa3+Y9gmhaNcJLqDCvHYFdaewoz0nMAeMfoNI/x2W+4zdBfrfy28Xs
fJjmNo+7UCUpx/xzLhZUID3F+QDd7QXlm6OFGaIlJmkmCEFOUkJPTv63VkPuDP3QQnnfMu/zcAaN
ZDf866TdjQTQCuyfjTob5q1oOJg+o374ZxJFcN1PnbdwO/ZVqMCKelV6Hj7Ed753bJOW9YWFnlI6
JrUN70uwGvycZUSYvFRBfxyPkvBp+fh0rQ1rCszhbjRSedRJ/H6I9C+B/swTGWcnYFRJiPmlqN7q
y5JFCDgqV+GZqzGsRUxioR68807bp0GklU5KsJaGFJWE8K3tjRfZEx1i9IoK817627y/8rHz9+SA
jg+H6PF1fdujEADWMp5h28Lvh0HCeoFFqwmnPZGp4/tZGOItOJ3iw+1L3Rf5HUaYLva7k+WkMDVO
9DeUJBGjfoEBa1K1RnPKVNctnshvTLmwBYA2OLI0KJ8bMen5s83jC5cmNLK7ovtz79EpfJwZ+p4/
T3rXbCTBValc8eWMzZRp2hn84hQamzHRGli3AxbIFbCpqgDmcmm0Dl6aR+gt15a5TytGPZFmW7RZ
VU1iYtuCKGWfYYOpccOjSxPLAw8m6TFwilx+6TTosTBVBZcJJYDMD7YDhzEtSWSGXppZFSOCyvPX
io/mmr7VMt+ybwJdWb3GN3WCbJXQVIiWHSfROXCWfX08XaghVj7MUGjOv5Jl2mZaZOuypb204qOw
Y8rQ1CYkTtAo+xEaQiDoztQ6btiPbsUhDLDLrUIaKW+3gja+Ta9GRop0cpLCQjOXvb18leQTyldb
j5MgGxXRvrJlC2mkTaAAzivLuU/loAH6Qda6iEzb6sH1KrsCCQRkb+Nzl5IvQ7RFNgLlq6DRaPWA
rlT3lirepFg2rgJSpJpdTBfBOtMzTAHI6GPm7RUNxMQF7SnOxBkT5yrUgwU6pq+Ms3jY5gJBIOQU
PlLIUTRm76jsOcO32dd8vXTQfAyy0JEnpmg8udjW0+39xfYrlMOGD/hYxSpRGg8XeoLlxKWPxz2e
/NW3FCB2bXCZuUBTkRFjw7KqQ0eEX8IEIkSOezcgZten5rsg2GGPYR8dcCsDts0WaiBW8aBnuvCX
OgxyU3mLOD7URhIh32UT8+TOptBzFTYKTZnOdrG3QyktmVz27gg0nqD6aYv7zPo0SbCLundqQq2B
6qOGWXNmCvHOicqEPlqs3gPym9ctZ1xddiKp5fHZ7Wpe2hnZ7MXLiVNg1HtqUN5O9764+4Es1z+j
a9KSZKbvn7QEDs9r9R5HQ/1u0xgUjxUFEX9CW6+uSbUkYrc2VfU6C4gQSmxhM/AnHjhncSOv89FD
ZJo3fwKG//VDLVTk4sKzS/DVoXnG6TrlUXF7c2NyjcJ3C3PKFlN9I/NOCMqtapAMaUCEXW0xIYXr
LKYRMwDMpm+tE/w8dYw4oWQo/hFRHdok0YuwPFl2cOdhKI3mYI3mDwnAPUHLX6B271sFuvxoEvDL
ZRjQfu3HZEd2Kkk179ean2tdTCKwQRQ01ZR91ym3Bi5AhsdMzT/yBvLmm6YcUZip65x3MPs3eNdw
IRlPBahDkn+vOK0kpyidRx5uw3FgXIP8vudIaIF8zJJ/IjsgqpVJ8nI+wtIE6nZNtmlda/8Ar13H
5ihiT2BimeA1YwQQWXoKuPasPyvEFZMs5Uw08YmeV6sErLxp+mrqvhAHCx+WX92T8K/M0blYPPoG
+WPcBfIMzqJNECmaXR/PQlV2EJzYPINjqkuQ/mKFC+JJaIOECz8WqJh/nz/BOH9wW8ZRE1qPtgGa
dBZjTGhdDN4s7TVEqTGuwPQtBANP38opW2yj1pCcwRF3px32ws6axzJbXROX5/SK8e4WSzOg2ouC
pK8KMzWn/56iy+pVekihs3hGaOpMnfxtqWcdbTXN5hyl+zuABD3bPhoyA5kEtS493ZQjc02YlNK7
POt9F6KnqC9/CK7pQH2himYQ+4f7AmeMGCArYAU6yKvsy3JBTLMkkQrJn6d9DsAeh5Ge4khIqU94
Or4PlL87aN19/0Ey3TAro0j7AdzS+rEqm5YxUTFrDk/wUKeBXCyhkmpS2zQ8Z0704ro7eddKa6rA
0TuvvLDveNW9hPH8f3DecDFFQbNwCmB5NPFz+E2Hwh7n3uH1H0e+hqZc5/D1sOZBcJTEPIlAoKQK
D4UGrBGZw8pG47lv4JBekMDSITZ9ij3pnqBQBehU5GTvKohJlj6y5/TDaI9jSiIj55r8n1qeXhx4
X4x3zmN8oq5t8DzmkbF84bXuvAzJmL8c3qPsLa1skj4QmoF1jVIG39gM6QS4CR0gKfQIHs8WuwzA
P8AUH+6APDDk+H0G1MA5oWAnzmP/gnKH3hIilMb6sH7iZSZmKrb+TeBYd7ciOmWznEFrWe3ctSJ2
UYNQFPqkFkLS78MDgXiZWuJvfOJNcXk/VOxGSqlWNhI5NCy2/h8hqNcNY8C1aFg9zfeQpsAU2w90
VBWmZXdwPx0yPiY96uV0Xb8WnRfqArl9R5k+0bzIt1k+yYohWCqmC/+D8l04F9kelzwTQOL4Wb3/
R6wW8s69MW0xwkK2SC1fnMmUNqnqFC71kbrWwSMqNJ0gr2KLL+1Oysrl0CMRU8ecjBOp3XBtxjWW
Kd5Rs5czVQAt2ms4FipXAXR+uzKD+qqVRFj08k/ze+9c4qUuS0GolM8s4swqexpFOsHvcfw0+K4Y
C0ND9tJL7EE55Y37C3oqPN5ZDQJAro+Z0BTrMDMnwzggcakHO+xaFKwvdV55JdIvfbvdQ0uBbcBI
mYMEYbkFG09Bxgmu9Wl/7ji9vTXTAHdSYKm+oYDYzywg+O2EZ7JY7/OYaZpmgqip2VpC7K2derXF
o//RBGRcquM2ROHO/0WdwCMwLELmL6OO5HfzO2LfS6/jwVsrJLR3hOIiNH1K9y8prXcH09T7B2Bg
0X4P5wV6PPid4hAfEPxPzEsW4PN2gVqj7dWQYTJ11zVJGi+jwErXeZo/Xs5xv9AS3pl14JmUdX43
FK2ej21F7fkZWMqXN+B8mv2DrltE75hEmQxwJpGZdXOVFUGu82iy3E0qFEG/atcaq+SAh2rURFlF
SlrPopBdUo1+9yeSsP+gD5ecHbyMKTBNVoEf+2UZ80MiNFrPvULoOKtrdn3+DeS3nz7I+EjPGNdm
AxuS+2xxW8ECE2JkA6acjMO2gIQxO6zDZatU5ON1guUfTaGsLGw4AQugpXSjghTcvmYmC4s6sejd
GDhhGQ2YT/gH1ecA6s79lPwTOshiboVzR93v4ugtFNBL9XdGimIWo24/OlXzd2c/k94IpydnI5ph
NNu4nCOHRvT5TloU9L0kjSP7AmjfH7Yuqg2n88Zf9qWcWTnNHGYjNwGIqlCaQrmKVyBO9qw/HbuG
bJeJxEW7KgjXccKCPxnPKlG7of4ebao8DC/jbp1fxVt6QY+G+BL6Ukh75eDiaXU/USEqhWRc6oU6
+PDto4K9g81Pps+J308my9IxacDzct4pRQ+zGxjNRISOR8pQF8ZdOkvCDo3EdFQXI2RKtSDBJXAx
xmtGcycKayeEOu7io1AJtLi0mwNMID0nDcaA3nC44S3OPmeE210rDMi4kkOTA3hMabMqNs0yAp1C
FOqJE5t86ks2yIbigug8vvHnBkMYSvQTPjhlQEpi4FaJpZ/Tt5MYAjmCFtgfGM1qKVLsLQb6x8/g
wMvxWTJkLhxOw6UJQOGGZH0ODx37Wk8vAJklNl0f71aQCDcSaAeynSP15yPTejHygbm3Nt/qURq5
p3uDCu1ud+xu/cZIe1c07wKwUMnA5XMHDE597LT6dX+O1Tc9nJryz+3ryMtr9EdkGNvaIyH35uo4
zM341VOttOnsW2UhBDpN5qjIFcyQtzIIjcO4p+LVzG+hkO9DFGF9QJYDBTBOY8xqpnynahmejN8f
rU2HLg/jStFMz7duZokscRp5wrpLI87YDvMZmlIttgPUSIBczXcdpoevNSTk9Jn5LOv3rueM/fEM
VD1pybQxT+qm/HNH+nsqROkhWu5R0TqeFGrMCbIg/du6Bt7AJlC9018HX9IcFYpezPdq4MzURpl4
lZzdL0qngWyOP9wYo1YeEDFpaX6DVDHq8eN62Nnwn34JNRDChU8xzUC75gw3+2AkOub70Hv00/Zx
r+U4OENsACnA6KGAm1MPVE68di1uq3BU9glI9r2l9CytJn7TUzdHF2Uz9Q/bg0N67XaWyyJGhi2r
MVr6MCYnxtUVrnsgSyhZbK8wVtH3b+sEygmzmr80XTo3RQ7wTeYTeePbNnats7VMKJIepKdy0hgF
wj4yrtIJg9CNuUTvJPMDXC4qBF6uzhUMbCbuJxj2/LIe0dvx+wnkE7mZpimPdLNtf0mGUDW/1Nea
98skjgq8IwBwyZN692qa3lp65tB+T/Wh0X/jO5IdjwUIXwrDQ/Z41HpRUHKsLIIdyeP8J+Qn3opb
r47s/t1COH9e42/FbiliMicaVHfopqXSaNExLcbrvhbS9+/A5RygcbhPNODPgizKPdgpOqVg9QAo
jkrQqJ+eSVQOKHhVgVJ65Gh+ilUwB4v/JgM/cuzdzEeq+J2AedPyW8N83ttj88xmVlE11V61xMxJ
C159BE9Lpl/9fD1fbtrBKtR+SaoTVvd432k56Oj/fTnu48a4vteD0TbTKQyPdyjenMuCZM/gqo0K
2QgCISCgnoRLvKuA/Y68QrIOxHi/afbteskXtiyZhqLRhrCrFylN+DYwOZ6vnuF7ZK4FHPhMMI9t
NILKpVWDdJUNLfFJXq1m6JcjPuzgIkDZaSjlvEey0VrrYB/k+sR6/dSR9r0fzdZFOgqOks5kACgI
2hqYW9Y/QeO2eLltTcNs1W8uW8Qq+Azkh1hf7Tcm/Q54p7CAoxFgRZOavnRxK9PP51aSZ4bkOvmq
/ed3n9WyJLXw8hItnZF5Vi17TCbMil2AyHLn7yJb0g0Ln4KWfwEnFGv+t8MFHhD6kAq6lg5iQgMu
2HpeGf/KDHo5yntpSHdphhotIFruv6w3oc1wp5OVwpjjdEaJ4pbNKRCrQnP++/6xW5d5t85dJiBh
4yGTCQz+qMfnoRV4YpVQ5Mi2HdRL09QJqv1Jz708P6dLlDEjufvrbcLgSiH/ucLIIcVWzrS1XQMm
rE6JWOO1AZuIRylvPadQa5t3d6Huz2Eq/VSCL0rkLjSCDgqcHNdK4sUfD7cv/oEsIBrrT1C19jOC
1d4fykZMVFQVU1fxMxnQLfYNYTbVHH/JuP0gwWM938TKETROpCpdjtBMe1Z7rFqMDh/p4nqqjLwW
IY8366iLkxpckwPGpGZPx2kJDFeYX+Y3kdjadRpcthrfvr6Fs0z2YCCffOieMXZaw2xP3yLCdOBL
qmXVX18EuSs/zwLwE3elUwkRwfJRr2Cbnuu/ovHlZVI0ano+q4XMEqHvlWHZBtvXD7zw+bSFE7VJ
f7YqAnrmWb3YvxRPpyK45edKPXL18ttGn+BY0FQ06wbnLPBaZCyA4lwbMCr49/YYL6OR0K+Wag9c
NhT7HSn+iERMKX9v9kIKKMpbPlB7B0929VYGAhljW0fdL6p8cHIIcP0vwQwnEZVsXVLeFoWHljU3
/p2EiuQSuPfPnbsncE+haywyk9GsrGWcWCpbWYxoSloMj4Pz3LxSXoHRuhNGk0s8hc9Q8VTSz2nU
6cJjxoX/6ZoWZWyBOUPNgb5PAC0IfwuzHrm0eh6R0Wrj8YNX/hk739mdOm9IPYgo/g/l4+Pst+N2
ej9MxYJ5QJZmy4ZObtFxxIcCHC2XFPShFalrtSRmbVGh4i0yXj0j24+LulqoUV56pkD5dmpsTyTS
wqk8sNYMcRe1y3UVo88Sm+8nuSWoSjAsEJkcwBawu1pseO+73/Dl06PIX5M1ffed21z/oVbMY6CR
L7VScQlzlPFYPXq6Kc+YBtRPfekM1k90cHUop9HecBcTaGvTicWevZBtoDMdp/B3S3d6GccVqeW4
wr2mffPLZqnF6mRWWc9YOvsRHNXujXP7PO8azM70LnQ90MmKYSYNXlhR+KJDyXTm7M3PFZFXFtt8
4oykKQzfLQ7L6zgkpv4N1yRHGPJjdMkPaUNEuHpN2e0HcDzv302sxaPG6NdtV41D23sX4YpVhJ4/
SDES51n1NVhZaOeGEEYlpBiHfNNVP2MaGOLPF5B5hmczHEABPr6fMehDtJKi9avvARQVDPSfqAA8
fBMPFUyZys27JSqLFWc2ylwy/ijsakKWY1I0vlL5r9aDVl4K9ZNWeBK9g7s8Y/oLKr3PQv/bDc4R
vRrWrq5YdyeGIUDlzrgcWGc3JeNmqMeoZk3CXjHIFg0HR1PrfFexYnZ8jrBwPdPGY4oeofdiF0Kd
XQRfN5Qn57dh+KrQ7ZJaQhvDZz5xyo1it/FLgMZAcwiCr6D/gQZXgSw13nrsth2yi+aSmWvzuCRo
VSmOKntNcA3wtGbR7cv3WOFAPeQr2jNC2X5a3Uy4WCns5xzkH9ClkZDW8PD6T1MDweocKMOH8OA6
+BsPrLg311H/F20AM0Q4IbXOZWU3uW/EM2cgWKtBBH03IBTjfzbI3/Zj+yOxXdGi+9Kx4E5kV3Pl
2CvmwlJ8O7HhhFSFIPnXN1MGLb7blgE+rNjM6gSJ3efSR1VNbt8cuo0gkqSg7qTqZz49Hknsg9u9
dsyLAOZG2/YJrxFqAy5jLnjF8XbP2RHtUW4l931oSJpxKZN+B+Kugl6W7mnCabnEjeAfvMG3AXQd
5Wg/6WLVE8Ck6hWz37PqTQlTPfaq2ggqsLbDvN/DF8oaIeUqYHRtE2faocFTtsggpSc7C7u3zZlH
2F2NtonkAWf2B8hYhsYSHIZVIMMjoJ15FnumDrkR41L+z7SgET2vnyx2WEpx4OfMDoQc75/8Q5JA
FcEKKTmJNgABa1jN2cYJqX/XMeJrMYc9Va0nPg21Wm0s67ABhh8u+PWQtwI+tsIp6dn1VVZVnJZe
SrEKhyPWYiT+mJE2eQUR5d9+FaGMJ9mCjg2TO8bscTbpr1H3uKWiw+v1GiM0WpiYyUOhwd0Ko3K0
GSbDGfbibhbI7AIP+jKM6ulNpvW831jvRyTuhdoHtk9nAKcYQtVxb34dRRxbqcOy8tn203CjpEuK
+SmFyUgEYXwA0mPw64UWnPTJlcDaHFzfbHj/iiMSv1avt64R71tDfcDWj+yvVlJDYzcSUHwOJI0r
r4ryCkTWA5SgbviwBy/cAzBIFGXSJ+BMy3JU+tXzaiquh72Njz/hgPVCphf25qgEaYXGvNB54Jev
AmiERinaRH9+zMNPYZdWLqVHbX2pTeqWit9fQMO83nnQ26u5EpgcLwou4rPSwWFSf6mJb66ZIWeP
2N0IWpudeouLV6dVoFIgocjAVdEwqRA9HFbREn/1AcdF790VkxbWwTF79FJNQ3fCdBdpuUqA5xwy
brm7vuO8njbnTUhNLFOlVuvXoIVjVjiRgJGmvTp9gHJ9gZYOyzaG2K7onE6sNbnm+S4v5uAcBDvt
iRVgCPcdgIWh40kVrhfwxUMo25EcCmUHaQ1aEVqq+JJLM9JNW5JK+1C3GKIjA6IjH6quwIdRPdr9
EL48kAKLoouUvsHkQeTsDktIkceDw9sKcE81x13rF44yD8FhhTC6TEYLtJDtmJBaYze+XnQucV84
gb2mhIS+bwxGCMVbvzXFzc64AedDnQI0fBurFelQyllRpRPdE9iBSvPbvAqmEasyWWbYA6d1nott
U/6RMJ7EH2SznrpwHctSIS0TZWu5Gwm3bM6xr3mlrp1dcfgc1UCUHu+gZEqvnppSvUU4galnkU4u
waKX2VTgmsU0BRdGm9nrLabie5M7MCGfiE+r5l05kWTfh0dv1jls7D2T8O1K/ZHBthDPdJTjPiR4
aZZwjFkDcFySweWlnlHngfMruTvxlQt9Zo3EFWA8jpU/Nhr5X5hxPsqMEXba1EzsQPSXHiJ43StO
0wWyXV2RjFBQHn6IVND6j4wmpDi1DRoJSyv4LbDQ4mRtD8i0N9DOOW5Y5Niso1vsL1fOzrSMKU3Z
ruegGHOptJBBhgHpHkTKkfMghtzBZtlfIcLHbrzZqOh70lA5RDVKry0XTr8Aispy8UxdHijoNAl/
Iy2IHmT6mtIFSi7JIBszEcVV/yyrPMpd8kzj1WmgK1yl8eiCGEdiv2nIoIqK1bwGI6CE3LUO9Jb6
5DYxlonpD7MQKzekEc8Yqfw7qsbiikFOuSioTK33Xzv8emiAyvsad3XQZM/LUo9oR1QC8yRLRJdh
sFbwmA9SZ4QHFcGkNBkB96XzbgvaEHHkFpu/L1oWFmsgvQgCLGc+3TZoOvq2iDdzd4G4zZ/Zpcpb
1sbdeoZY64ExheBa/wh0psdPooi35f2zrme0DrJLyMkHRf9L3RA82SNY6WVabpYlBIeUcF3XTKmS
KHWl3wQkHrBBFNDCJJPx9ubt2kTJ9MhCK6tXg3aLD7OujrIWT7fqg3bHLQcD6uHwwfi+fwwH5S3G
k8HQ0wxxqtOtcNEaLlbh+Gh7Wu1uE9Gof8Sprw9afKx4JIR8wbv09qh5BDX4FZuZkWhrTmAmNQ0R
kQUkD1GKo2wXYDUxcD5rhtUZlqRv7tQx1/Hh1WLdafCBzXgg0Pc0t6fwmDJBCg0b5F3akSc3VMyE
uY7LysGcKURzpy9kQIcUAI405TJYDOZBqG7Lo4Z9Spa5+4hr2cA2wYgMmjYtNJ9FMGdjlqART3OJ
q4UgPtIZCrjMbbcnMfvmRkcCGT2PU1Hg3gopIIkAams+UwKgTQ0qFplaWI/+CSZ0Yfowc4wj7qs6
Y6ACX9R2foWbVhQvLaGX/MH+ZwI4nWM6qWvmS74W9z8j0X2V3BLfIjmM52AwfhBxzt++L6YL542t
bDbX9ZPRCKI3N7xVISIhXIeQTGBBXnoQafbl02MnYL7mvkkH8aU8ITKdfs3+K+9PWfKF/71W2rU8
f/GXnZZl6+nJp/MJ5qgdDSUeX+OeLoRfpgrMs3ExSKDoKWToW/dc964s9Vl1ep/MagT98rEdN1+z
D/SacNxbu3SKAAivBDkwM0japPM4wcwkZHTrjBqhgXG5puEUwudO54i6tmEmipyMJG4rtkhRvQAg
heUYetkbVHCOWFd+N/nWnpnodLEkwLaza9Ykzp0ZzdENsRToNf0KlA1lCVj4rjqUFdF8tD+GyPGe
9BF8GO+Q/Gw2UGIYGP6t1nc++b4cUbyhWkIdj7Xxsg3912vfXXKyWcYykg5XMNs0zvlNgg90etOr
K5mWyPtd7LFl/FaOTsPmjZoGmo2GZnAFrn+SYwELh25ALyFvYJxAkteufizsI8EsDgl/HMJYwdoW
B1xsZE9CQcrAV8FCrR+K2J616Gd1Vm4Nl2c8l9+DqnvblQD88yJnd1XoHtBapxuho++zbSOMNMb2
OGjAIQvuL1l+r9Rh8OcJCh6qrbTm/qHxRKDbGBgRux0R4PAJzIbt0LzUGhRCY5fF8nGjNnnU1cux
i0a4vMyIk7Y8QN4HfA81aGHhDFJDwiVwLCmvBCuVPpAjNhfIz/xTLj67NqOwKeZS8Jq9OoyH5RaU
ZvKezeCtKqy6ew181/DFJNFsj5pHcgW2F5eAmMT3ng2YDdsj21w7mReQtrVtP1Z+OC6aBB3/9BeJ
e5+zxwe4NiJpw2E0YDgVaPnYSAv14ClaQgxmSU1iWeM7xC0Tnr0vGaoQ+hNtTEh1guh6zLyye3Cn
ak2iyHOhoasAD4i2mJZPxliw3TAz5ce6glnM7znDLH5nHGy283yxm++V8XIBIgu/Y6n/yg4BEEAr
YfEByuk4xlywElMB2xIG0KODsTZ9/vqZqKyIWdNS78DpLbRjXVOL40l2Y/GeIPLfDnYjo5KUh++T
gXwmma5dXYEbggIfX7q3G1sShiG+bLr/TutNKMaCN8JYKJTXisRJrEhuAz8yZWf6YLA8hvr27qll
+DZWXYHaMqyJ8b9awXdnRz+eKr0M05BomylW2RJwl/uduKQNVa9gLhJtmmwtINRRKbr7h5zXhXsD
y4kafDjWesiXtzZVnc9QYO37NOv5UzmNAR4SX7DgC2+IHG43YQMGX3rDa3mXCxN+5hWszxCY+vvZ
86DVW43D8MxDQLBIGVFJfC3tzbvHoYdEOlI18HYSOcILB0GTISe7EWyKf0/R6Ag+pi4s9pag0L4d
cEmAbiRJIq5XAnlcN280yM0lPBoIa8wtPHLKRCOw5+8QZaDiQAEnO6QSf4HI4xCMUJ33ZPUnnAHg
vXr693Mec4XUjWyFYXoR2zRSG0DL7jmBGhRdvlU3bT+vDfIdXEnYn7VqsQKvbV37GbO6dWyJYXBy
td0rKQUuuANP8v0o/AGMSlXdFOVMEufxgqFlCkuawNkp2AvumBZVSqDlSTzyeeh3lj09R3G6lJdQ
kv4U1NnoCdZCkVPPBexccKsJgHKK0N8qjNVJFJ44S+psU8dnMn8EDWydhHrjTi7N+GTBVJyAbmhU
7816SxQIHFb2ASsum5KKX3ejBpBqR6Jcy7XqI6HMtLPzdawzkDFUSUWCmZ3Qd4RLcyfba90B2bs1
sE3x0nt2+g85owotyR2Uz5ntfPCrLluijHXYeycct0gm0sR+xQp8g3WdEYqQpTz+oYAbYQbtNnwP
R7SPHoM7mZ1QQCkW5p+MV2NIdku6i35VZHrbIXstH2npxo4IlmbfSVJsx1ApOP2o4PjBqN8Awcwu
EnUbm3g0KAW5pDWNqktoQLRPfBzb85ViYL1MBwSUXHazr4Qh/wCKM9mnqtRDDfzJ0jRSuPJjkV/3
ARWBUZFMGYpazzBNUbbYDyRftcX+8b678tM9T/C/rbuKLRjwmIKf16kHoULce2el3cKvl8d7SlYT
UOPETeA+ax84tSLzNin84YFIOAH3ke3jTg1LqqEFmaL0SgSyhkXIzsazVyAz3vTzF6UpQ6I6oXYd
+HJnuqrRW4Q7ZB0++vGvTqCiqkZcesHYBMP/Gnk4F8OIoILtAJfN/Ai6yOkvcbyKLLOIm5X4or3s
Zof9zYUBU+rqbL/pikXqGkTa1pRBiBQ0ysxqGNcmtMjaAbrsNtV7mdkjFrbYh0gFC14iyQptoHUG
RFnsSDhEEIf2BWpl22iN/P0Za17dQ9TXqS2RV8rGnQhg3SHufymI66z0OZAiUUyc5ic05rrrQVht
Rp1QOEw0/y8xD9T+OxHWhypc4IPn5PdNHFVVrliMhN/cCTDTJJyxXnYWAC3vFArdDfzgShYdbUqq
xWrbgloQcU255nzF86F8zd43eheoCHPRLVcTcTcUGvL+30dDwBRItkpWdVJe8KPWtBjwddZ1DJPT
4/O3BLfAPWf6MnU2WO5jpM+/eLbx43/RBCuxw7GdlmAMchQQWUHSk0EEfObxfylO4wXpSDdp3w48
8XF2AmxlOA9IO2QdFvD+5Ejtr6a7OdiMw38+VXzgnFKBM2rM3zu270+Yf89ypssaihMU/a88Nwa7
sU+lzO7WBgUuXSXkZ8EB+mTpHQohaWUf1fICsYmt/JOVeo+DWf9JPa0/aR9xDTRhYCkTdvvJFYiR
mY7s2BXJDcfY0gL2NH5VKVkfQXe3/tJnJOY3t1A7xc1YVcLhMiRmoZiXQAS65PMHihJCxa6WLxTa
8laar3W68KZQuu0s1Yw6J/cimjCYJN5AjDkz1rHqTao91h6YxQ35hC+BEJGhwqLL10meqJ+gVw2U
o2dhCjQ3ysH4adww4EUVghTtTNhhuWvT5JDxHdbe/71DJxPQJ07OSsFXUrCFn3GuzM5Rxsnfz5qf
6GmhS3MiGexQDyQ3XNqhqroknolw9Fi3p0Xb/CGXABv1bf4VLDQvVGMoz+SfIMj9O7NN4T17Lrzb
uxWUPw9OYIcwPede+Kbo0VIKuT4mGb0L1sDyDYFgE1CheDOYekCq1FrieFRi4+97j+x10bkxzjhx
hzTN4XZkguUPjCV9zKgFbl3nCSVh1O9ssQRcbLGpYBlfaZ2lLuJpNOSLgXM/5Pts5EBvlRlY0j0j
Sc16HQf6WNUXI3m19/yRFO3nDXclbAmq6Gq2rWECrZHmMjtV1+xnoxbyC37tiQrOxWVR+vCps5g3
724lnuDU2bM4eOeRGcPcg2SnyF5zHGKK0EgbJE6+BtPTUlTNmNpzpYPPIycXS+XhBd9cyL9JnL39
7lOzhnctp5/voYapWEZm5//jVKQ8dtOAsIeY2OqlNiK5pB7sRubq2U4Fov5nzVSKFlQhVMBzIS0P
tBqJCe7P5PC9Mn3jkRRp8SQiUGaWlfzJAbZY4PI6SWaT1sEQv2rHpiIBOVFKNBvwuy+1jJqpjbFm
H52HWPF7EDoMmXAAVG1XTC6UCmJhB/fo79Ih864A69bCw9hHOvC8rIcPHbn94VrPj46zjkbfKafs
fJjVrzQHuZ3QECdWbCCCnVTMeIDMWDEf8EcCUa652X+uPACLYO8yF+gSxThgqFDraEvisgTFR7Um
9BR7LNp1BWgzFbClpjPoWkz6GmSS9+2NERXxAE0wVaKEFADzod+xrq1H2v4g9BUMmXlPPg2Bb7xS
k7Y+7jZSz9yEClAEBO5nZ8CRy18l0paxDwiksW3/+WOVgWNmwJk8ouN+0SwiL/1Z+SXtxrFSoawH
+AE9N5xfXOeF2UXe5Fp/yIQe2+OE/UGAGmR6ZLiaE4RKsOCoeBtGMs0KFCD+Ye1qNFwXvsH/TRAs
Q5ZSRlCIh0oYod8njsAKt+JbZE6fywM/vOGxnFCUq4gCWALF1N9xsqUgs0PJvgILcR+A8uALJJOh
wnGJKPkRS8Svt8bDR9zTGTiEMQFNCmX5MJGAj+vmRC7dzR4p1axkPRuQVLOIHWQBgjxpgEHuZJQ6
ucvLP9Qxx6NORzT7ktTKorEvAwasMgOnP42IN7Anjdwn+XucY2WbD1E37DyJ8GBUnXweiRN2Q410
f1HZIuzMJPwLsku6juz7rJIpfw3DhFSKuf/t/8KFVqBkqVWUnKZLmHfMexfS46C9yhbNHyp3r9qD
5Vn6gGnajqYA+rBsKwK5on6znk3kaBy/QhzAXu7F+0NiarWBqrUJSBc+csCmwe9pq0QP4el/bmQW
o0XVUuqpdN5xfAeTbcLZIi9yoMOyiv8ey85mp2YF0F7HG464q7Rw6dssS1v+EEN+vOD6yw83uyWr
Z45FWOJmwO6HZ7tXed31ea7TF1GcEqDMkwPTIFj7yhqzK16bgbBVGdRw8Q6lxLRToqM/csnhP/ys
zZbehrrEw7AOTThkv/qgr87m1BlN5TW89UHpmncrhySY68xJK17+WI9kjNap4885nrdIpGIHk2B2
KoHA0oZ+ahha4uPyt7d18AcLqHvofea14MEg2ejqXe8skSt2FTXoVwXeql57PE4Rjz1iI2ceveIi
kR00ge0lDs8M/gE2Mvnwa/VmtvoCJzKpUxZlEkoBPbIItJd9V5i2ulu3GbFyH+dZ/zGQvxg0BYor
4YJH9/j2VfyUv2EiQGLSaAMDnmgA+3mLudWIWVTgPNh4F3nCu8gWnyRcGPcGbO9saij6lEh4saYv
H8CZGXtZqpP1AZZh/2ij0tpQkwRstm+T8conOQ8NDmTmgVs0LcJ8YTP+tI8yZu6Ypkl9h/fypIA3
eoDYXAp0HrBp5i1eVjaHM+Rj1lPBxVAT/hRu/xL5iSMTSO7AYVwdbrJ3pVsp8qmzKa09P07k6/Qw
J/o8fOr8RjhbftIO1uU/KfHrR3haacIvomltG/+M8tLDSiNIAEgak81tKdLLhfWTc1ObuUE7AKau
CeaopISjdUl9AgILCihqX/TI5D2gWh8lsC953VaXfrBRCA8eYQyOAiRJZ3FujDSP84GegtLu+QE+
Dd/Kc1lDUujUD+Qkls9mDJy0GsL+6V/SdLNuSWGuZbadcPbmYyGpakogjzxqyKxj6qQSuxeVdhEM
4m5uI0bmpUvI2euvmDZ0Ai2CNjHZtUZPvg0HObvRt+dXYsWqvEpJP1VDpaKfirzgDxFpkFoOvtz7
Dz5ew9fyk6ol8g2RkIlElMsozU+cQOuy5XAzmxtF8g0RJOUFGr4oIpgwfIxz45VSHHEejEOI7Gek
PNZfmg3HKsW+bu72jrexxHIPDG1ARCAiQbaWP2H2JwnwAiLxDqll2ecfrxdYS0nTZRBKGb0xFShK
LF6W+KnkFKtql0Jg57WDsgxClmWU0mzuK+gnz7bKkuFr/QdrNLBiSVq5boZXkcK5bV4e6zEzFuRN
IpE2mL/dQw2dvOcOhxHLDmLKQ/wkazq82A4rXOQcf+XTHHnM5+YsHVGzdP7n9bxbD8w3d6c0X7GI
r5SljgtBkEiRUsT2KdTycMcfG0jdeZX2IZ2eAL+wi83iDm1fkQxK5+nP/NQnaY+T3kXzvR8ojiTH
IT8vbBnx9PtSY7nOLkxswXIHWrLP7cAkSOlyVuKN6YQWXaPBlJ7I/XyEFX1DE2js0AUm6sa6kMAo
tyPEgCdrSb4H4vbQYCB7ruWskYwIMAle6v40zxaptTVTJ/D55P1PJ+H7ySfS4Z8S4fI6Q2kuqrgu
lVG3+2PfiHa2QQ9VRxtt1gQV4VlN8mil3f1gWcX9ojhtaNPtib/7KmVG4iYbTdFPa3/rFzjpjrkf
glYz+cdqgvYadgPfXE2120jMReKsxtLHyVV/TINOLTfS4QIeVMeAEGlSREk3+abCRdWssjeruo8j
gG/VEjwSHZb6lH3WtQVrYn3F5icRrDGnE+VZ3euWCz1/cwoukoNGZm1FFjoZU+BWf166eY62GPax
bcqc2FLOK2RD6Rwqqb9N3quYG87lpQ9CZnRrN8nSSg42c8pZhGwaUdnLhwWwUZjInBfhwOpocwU9
90mHos4jccpJQLCkJsCToSskCC0esasnlwKDZblij/BeZrwIkgfRfO6H+QfX/g/K+F0hHOzKrQYH
ifXULH1jtjSSfQMMnMBugRJdJ8pqqnVlPtKYhf8uI7XWjJ6bl9Po6sXGsLTlP1G4NAzspFFOBXIb
6IwfwT9QZiSEFuXYDgZh5e9j9iPGii1dQxgUFiET4lueExmmessI+cKdwPgTZCDD9d0OWotGttKT
HUGRhyB4X9sD2jge8xoyhYpjwiQkcXzEvAoHlCWw92avMT7Y9UZ6Ppk0bmnYMh3raQundg6cVFAl
60HgYngws9XLARmw+pkDclWpWzxiThySGuwKUvtXBkf/+BYw3TdrI2S7BvHbzgkCTe64EcmYUGAj
SR4ZTmk5zyhHeC9QeYP38dUnoHQBZjYsAB4xZeamriJRkiSYHo23S9KtgzhhOIIgHVuBic9Zfoos
k4CtNJrNFhDxRo3aHuBNeVfawtkTD04802Nol+Lx/cUskvxE1mk25c/AtrJEfyDnVXNbYqpQJS/U
C/6/asLHHrD2L4H8Jl/lIxFKPtdgnDZJfGtUX3bF2MGAgomTGGVaNnbMF8WliHluc9FHaPMl+7mG
i85Zlkr6f0Bv4r0Uf9drJ9v/ou1MLXKpXEepf/reLCKYOWNl3yem8vezNflLgY+l1oaDm6bMAW9W
Z3UmCPHaNsLjID0eQRw6scpJvLdenOBjDr/wxBC3G+NdxgxdQNupH4S+W3nA0xHJzZyogelSdMq4
Ql+hZPjIHZOkIlnkThA1c/Tv+lvt43cKKCQSYHg4ORNwok052KdwTTDaiQ47GCmW8RmPUl3JD4B9
ZSiqVjbT7G3pUykYXvOOG97qyw0EFwHzUQLCbTINyZRPxkYwXyw2MMOhnFaTi48DGyzW6hsFp0V+
jlHR0zWit+IK0/Reavco5sxZ+CcKIVTEZ9j8ezJfTF+sGyz+HzoWr28fFLdCqqMWLKNgGl7H82iL
ZhEXvuek+UYQZ0+HBa/mXePlLUZNfV6Jy9O3nm8/7DVq8nK0EucGW4ktkoGGcVf+EAI2jVW+16by
90AwARxeXgOQFS9ifh+IhEUFBydGLAkrDi53jsKiUdhtcADTbL0buo9uJQQfcJ5nyGfrOXnYosNK
FJ6lnuqgh2FTRthINqHDF0jJe1wxAdd+MyQTMnz8udcXaYERNzKiSIAwSGPJl6krhI3o3c0JWGmB
92oTbDi+rVI+0g+rVev2BY5c6us6Qha04/6WAv+sEJhNWI/IeoekW639/pA+tfYNSYjHwMhxiLfO
vnD8r81BZNPyHWPZPIOZV4nLofrMRp/PMYs4fwFKiBFL7vhjM9IBYVmGsRJs5ZjiJ4uxMjyENYTk
S2Nw+yLl8K6W4t0lD61bUmI8GZvZ1sbiKGVt/J8WXOdlsrnY6s6b/ghGmC5sVDtRuWJDf6WrMp5r
dis+lYwZfQE/avhaOUI/4NjP2T9mKrxKypgP8D84i9lCU57WbYPIAVAJepD4iS5L19Nt9K6XRN/b
F+SePX+hEk1oX62R3Yo3lRJ8R+hsw+QrmEMV8RyU86//xrbj4RQgtZ0YuqbCIhQdTFVQqOKMSSio
5wLRoL7O6IN+VLnhL7H4H1S99ov29sTzxmafVxmmM4iYCW6bfgIMlDRAsh5aQR85egGCDtx+Tm6k
4YItH4t5+9gwpsNCU1VEiqJl4kIWdbBRJaUoJQcvWXQp48OjB5wARjVo3NIG7R87DuSjVaDDibO8
/a2wgZgEuYIvfUmN/yYQd7PUWQgj2URTAN/jBw+PnfmfacFkg8ZRnhnAZuh4gmJMsvADXyP77Axz
a/EFzYsEUpFvBpXeMjfro2e7o1f+nIT+ijK2bbSXu9rNA3FZaSZTnTQN6DkRrIEnpE0gT82Jihw3
eO9RgzyKBzfJRPKsEKGVZonYRJM9j0EMwA281Z4PJtXwoDvC5WpExumYMfxhrVWu7+RXxarYEg4J
pEIDiRLXY/luTz1KbOvLjDq8U50v26+mxNKqVtHOMjEyF+FyfqUt0evZaOhmzsMEFUyrVuE0Ol9V
+xYllMpo7oztuUw2jr6zQba+9tQzzDtWi0qC3UChDI/2QYPlth5pYtJljKqcbTVRV4OCtVyWZwgU
ej970mgPZOZKfamvhFVPn/Nn+y7UNv3ye0xlRWVchbUfEExyThIMO1Mxtccfx5rELYdvRubnpmKl
JymxLl0WMWYAafuq1d3nRbWTEJZeWCZXrlbPa/cB+dAA7DDGGPVtGYNdytzXuTiRS8ildLkh3ue0
TRI1GLdYmXx44kbrJ3/IUMbUBMov06bLEePSzTphVjo/STumFhaGBp3uKpjW09as+70aBf8ljnLe
gctw1ThL5wBbkA6O/KRsuSos13VFtfy8nbkaIxmH7VfFVZW+2IO4b8BgUZWaKbROEXCJ5NPiLDsc
ITO73iD8UoxHIn787hbNUS0LjKtn8T61EbOZoMseNLAN90Fph75b9iwnooWa2ZHvEJzMBEdwCN7d
6fMLLhdkED+jMAjK46t1jonr/czSiCilHeOjG0LN3vPtSGT1hbZbXvw2dfVfV8ycgpRfO0sFrUfb
b6oShhMV+fOH3ONSK2ntkw1TMXeiHFyR3qQcCp8hr/+n3i5ILMTluvhkfwYJd8sqWTXdn2xIIJq3
dPqYnxrOLdpMY47l82xj6H3/IoyT01IJkxIJb7gLvtK4BhhAmegD5nSLa5nwwugTI69vbgrBKPQq
jJn6CL4O1rIX/n/Lz2A6QtKQdC7v3OAPxVRoFkyPkRylPyK9LuJrjYOCHVXfjjpgJSnQXs5CUAHY
CmTxvi2ZHpzJpIwGZmvwvKLAX0PXvxwM+3XdTym18PwUl4c+1Hf6G+6hd7xGmv93vcvtNiJDkUvp
huIOo4lrVWUG7TYQzCBEgURARYlRZOuqfjhT4SmsTNOlpStWxiANWLN6Dqiu690xYJxncoA6b6Bl
Dyv8PbhTOj+KaxPX7URLZsQlkB2j7DgIzXakLzAJe/qayjXQ1Gqg7ThGeO00hRhG/kNWTS/231yF
jq7/DEvzNy3AJsts85wNzjOCYhQnq+bC2OooktoNyRVKrZQtstvvY2TgY6nnk/DFfBtM0pbQWepl
hOHhA2JibB+3yScqLQqO36xcjTaHUbclK/CVz2ihKRXzFwW25ObX3UJBLkk5XIuyRMfmLgTa/VG3
zysvgtMx9s0kDeHJO8F8BGr8nt1Dz8PRGSiYKnNwl1elN7LVzGzLrdxRbna2lASbd5met+CKNV3z
sbuRObuC6eZyyOHh1nh1fAVzfqD4QJG3//su3y9eBMkioUT205yR7xpaYYMfiB6tooIOqt2HyEV6
LX0YwFwd/duvvxbUSSQJe215wbxEKASMJ3L23DApIZ+S/+kn5wBpsOVILXq25wZikF6J/iZJEXK9
P0GLEQ7ilpdljefQe/YwgugpW1eV+eYraRan3nFDyWlv6MjdhD5jNLK2KE/21nc+GbdEOF/zIZBi
wu8902suSzk02tmIeGVCzi3jUDZSzjySzBqvGQsttUAx/1v6X79Q6/A6+ihJn6wl0JEYkoJ8yy3N
w4STwf7laub3wKcgmObPdlxh8fts8XAMBMgKDAfAGg2Mbg+PP8Qq9mRgMk3vAwfb6g+9ZUGlHxVm
eOU7YXBbP0gYox32E4RHJCI6vN5NSqcbm9yAc12/IPE2Z+IsH6Uzj2HPfG2bhx84C3sFLhBV+fOI
xTaK2ZSw5M3uXdddQZlra6qN5MLADNH8BoVdCDuW0lwiQRFlRuStKN4Cjk/vg8O4RCyw03CLGwYD
6hIf00qOa3QPh4FjcnSabmsUlhn3Bl9HF4E2oHL9afq8kUbPoT1oMDXfV2XTA9wvZf/qVt8iev4S
KilGK5i1GGU5+bEdHBALYR/rb0F/ybWANE82vP44Yuj9S5Oj+EUe4ykAsViNMNjVuISEaCyuitIx
irrfBhuPhRxeygB8bL4znGvUHfKqH1ZzvP51eVRBWZ8ZA20XO1JxewldLxBVksBCzj77EVLKVFPC
0d/KG4wARGwemgIQa+3pC+9k+j62mQ2nrdb3VEQE2qs+iz3ZnR9Zj7A9bAYHzDHvXeHAzYz+b+Vb
d8rDmsrH7P2z7BEeaNjqZglAC3o0kjZPi6m4menHgQAJbjW7ebJb+mDwHF2AwhUD25GInmn3l+Tw
OhTnF14zcQcW9SQ9GXuZnFloigXBeQTYCEOpEnxIBjy6KMM/6Zhz+/oEAfWPxg/U9Mwvhn+1GsSJ
U28NlXjMKBCqaSz5vBS3u//vl/3oAKtRxAVUmdPKttVEsjSSJ4xiyUsm365BU3A7o32HKZ/fCWsO
jl5FQ7D9xh3rhMqbeZP6e14hgGZbOABzKDhRY9NA/cPwZ48XEq8BllFym+7Z+N5hiAc9yaYdij6g
5jRJWKzh5kj3tb2DjhjugeZKX0GSrSwcpaRcWcdbRN5bK7UmrUh5afCqfeu7pw+DF21F2UM30YHz
JuSXk6r25qIbiZuJZ2sAhBsEg2L27IeJXaEPeaIslxc/xKqE0ryoiM+nE2pcfDY99HE032bXw4n9
86NgG9T4hWHVzTuLkB/+40WVBEjvK60g6NsUaR8ZTYOhyeHTG+MtbmYQmH8JKaU79seiB1rC5jeL
emUi+aEZHH4l+QdBySpHEe/pTuoEfZPzpnfBYun/wx/CiOdgoSLElLD5T7aJJSjnd0qaE3S6VSmx
fz5pXYjo0eK+OderAhNAkLsvaZ2/OrDNBiTr7YxNzrzQEGxaqDrWo0xnkmFE1AeGwUDJVrbj4jE7
UDR1TLjPYXlvjJfIbIS4/D6dzJZwZlsEJnqnh4CZ4Ds+RE3iqBZCpwE5uZxyQIVo/XAGsxWfq4oN
tzaCr8cTEfqkHBTkeqr7T6JTq+b5uHD3hugvr1Ky2OVREyx3GXSa8lhCACiuv6PcxmFh4Buk1Efx
H0rXaAS7WvhbVugtooSFDdZnaHjuY+seMzfB0YZdhCfTbIMXQbmp6UNvwf0SjCq/8uLo56WeMjZO
cYVpIspqud/6l96jIfzRhMlFSpBR94QT6rNHs7YljErwxjyU3LIW2X9MuYQOZwp1HMy+Z4uluukj
kceKXpnW1zh9hOw3AcZLibPyJX9Kz7ZHe/RTTSdZRPTO2IOdj3djuucWOlAGthYKsq0m1JIEkznA
NzxO8dv56HSe4Axu8CzOthczdebgA1AWSuSotwE6sCpD47FnuQExDiYWDHVJSprmbHgJEnPtMqFy
+tLxJBbbmP7v0XQOAHaAHS1UmnXoIY94Htah0R5HnUQ6OVWViqTh+u7pWH720F8dFB37OGh3N02f
U1gsLfq6XHAf3MIiTObGyobTjkD4w6tLnIdyzGvIAwoOKPWv/xXT1vB/1t2kJ9OoerYmZmyM5MYC
buY1ZQknCCFhvWfPAToCE9oPyeMd3LGjqsH1gChLaEaRG3lg2Vcu1jMdLFqRECyw9N2N7vM5GsOT
iYaN0KqTOVoAfWW/53yYHHAxfXG/ZsN5qhHGFtC7rgZ8kVfnq9UnvyYCgFoWxu5Xcyka16cP6+Du
F9T+JeAKXp3v3bcZi18Vt05b8R9NgLGlkhomnRpSzkEPheXUuGbgLjt03sBkGvfw3jqLvvkDSAms
XxU6t9ibUwwTeTwjv012HgEjjhRsFty2m9gieSo69VdNFqaOpSYi4o/T2i6QIShFMmqyJHRbJT2Q
n1wfLlmiL+/4ROh89j793TJfS7ZeQ4LcFBdkNBERxhajzjpLU0MRK9gRZq6VnpWasf7jgbwMO3vX
a/TJbpVbeKbXnX6/jxTX6VE3Tn92ozb6d4/1EAUb1UsdulyKKFqvGiXn+bOXnEh0J43eUAwVNgTo
e1SvSQgegQFMp1G9t1fFMGD4aHHQcCoQ0LZr564DRR/pjo3M1l46nD6VeosnTcqZv9PluncSq4p6
NPLZug6vi3CvRzjzOM60t0BnhzLxOP8pRMRX0c3ohDxkb3Y+iQLSkX2xlJrEiIna3vG1U6ij7gAZ
83/Ltyt1mKwtBszU3Vrt8bstQno/VFG4nL+FDrJcGGwAq0S/MbN/BLnVBDOd6a541rSD70HVb3OE
yQwWCakEqqj2t18LEG27CzkbF+FEXn+pcvzuwaa/nVVL/ZiJvUV0/xtaeNDH6TETHfG72obb3bKy
P4HPZMM5/fvsSQ8pok0GywGvIGEfllvEBnlbuGR8Ssn7Pz+UNEjZZ5X2H0wsyD3lNXxWj8Xlvj+t
7OHWwUW1L2pkXuv+21Wn2GTywlLILjDtaitJmNvcUjrBysAW5dfCNEv66q/JX4/fX0v1KOPsBlch
ZVpqGRmuLjgYzX1biqtmJqtehKZjsX7jBpIpn6i4p8PKLM+VCX3D8v0j1NQeT4TvTrU4CCMJpg59
M7Brywf75BVc1Hhs9RQSWpJ3wrksbPCxsBsABTH8u8RBRMNerd812w98A8pDqMFPTUAwwRuJhJi1
fiUfHLBB1diZ78KC/yQINc0KlC4682Oikp2WAUB5rbvS6DCdF0VOnHHE7o4ty2Owqdfu1ZYf4j5Q
GcgOYLY26K0pfp99u52MkrbB+QkQs6p5vkkNCu+RWqyL7Raea6kB1iDw/yogy+SP0ntdH1GoyTqQ
l1GMp0ZkM8YDjZdE0jWSBh+9dK+ivwFT3CiVetsNVGLmyyjArS5CIE2GfBfoRiYaU4gjxGib3ae4
ok8Fi33axlRXVmswqpj1s5Xeg3/nWccyRjX7KjdeKgH6emQFB1mTTwOSYUW8V8x9wJMih9nUeS8t
Wz/EK+P8rwpyHzNUohmG6NNIiJ8KPVLc3Ke+Auy+F83UdBU8F8kh6hsWY+EdCz16dAUhVKG87gcp
IdORAdqlLkKQK2EFAXaQLWppwXQzqDqqOXze1AbHMsWlfVbSkamuyMdp9/8Uven6U+dlWscVAUIA
zKzKsT9ZJ1s+uLxMgc0q2vHaYA11FqwwwFSGBzU/V4pb9J4N8me70ymtrGzV5Wes/iDPZdvA36YU
mRa4CHJWvukD+tVer6vgoAMfSJS/JAOPI2N4USP3vSIaySiP19T6B3RVC8nOXM2OD3Xj+fPdoFqV
Ha1UHKvqvK5u/dCFZxzXgJdySBVwfmerxSZHiYpzmNycgbCmqG5CQbFJzYYsflJ7+fwq/sPR3xhR
L7sxvYVzcfHUSZr7UkmBoNohB4d5iCn2BJ8DO0zJqeaJ6Lg66IU9V3KSskz85YQCJNzM088KO+05
d2nahk9QolMTZpjDdZ0Fi/XXrUu2kAlSnvzHRcsA+CcM5QsCTgCcyoDVrSq1Wd1OjKu6PTHFSHCD
vUFe8thmHJupQ1f+JdECKTisoe9HBC1Iylfl7J1soFkKlwbdXyyidJdPnSK/q5gfUfWVW2CRPef9
5MEQa73Ipti7u4oWV5MP3ZjxZ6WOMwYs+Ao8pbfnDHBaeFZAFR6Gsugx4gbqOCTiSJPqqSsPEjSc
Ca4x7H0ZP9V8QAanl28dwZ9C8zdF2rX6MOt3gcsY+y40Fj5UZIdLqEfSzopS0JY7foe9498UoU8W
EjpUBCsAkZ2rsdD6gwz6KvITkTXln5iX0Z8UJKFCnnAwUxtTlBHcDMckEjQkAqf1hzF8dBG5XedO
eEyEJI97rusXwcVqXxmRvZKFWNdrWKuBEu+jw1giPKm26IEhOMLY1m2D1md0tUTJtjeLSEYH0Yak
e71VRT21dL8g9Qedkh9TYY4zuOFDproHYTzjoG5KcCBrPgJrsBq5oD1rRRDAs/shfpms4cxL3lEH
EkeAHOYEWQhSHk002LFSbL/tGnIy0eUz6W360giU2LuYRfuSGLQM+/4Spk6wikEEs8f77u4JDYs6
9jXmOQO7GrNDtHN5nUKqcOdp1NSn6NG+ATBgEdy3J9no6w5UOEjJ5KFXZ5/W8yV3lu2Zf7JHvZyZ
jkpqWAIvVjAT1krn4m+UD7dz5+zd2UN8adrWs4IhceTYWCobt7IQdyV7O6mixC5xJ7bgwZvMj+f7
fmIwm+4B3DZr0XRKLBS2n/OGMzyaiPo3MN/hD/YB4A8wR4sZcVeRHyN54QLtF2MmoPbZ+UyjMW1k
tpX9akNiMnYJXXH5xExWN+V7BcbARoWz3scXYgaLREPzDUvUirEOrr3WXU0gEfUNgIuJ0w4754+Z
4OPKH6XBCwv2kyGFLpaXRSNCdQ0IpcSbBwrfQ9oxgQE94V+5zDvj0KtCYSAUmy7aQIqR4RnUKmz5
S7J6n/gz+VkWHe3/6ffBCGO4gbhbtxMO3VI34I7WREVj8Xh5rSiGgLBL+aUcgY2BH7eVDsCqFLi6
mKD1UrOFW7ldYsyGJYqai5UtOTNLVYqX4LRF9lnI136sQUNAcMFTlo4eNxG0A9BR1NP+R14XoaF7
TIlsKfvWfW5nYuF3l3nfgCtr4+b9nZQ459D87pW/7bPfSS2YeB1MaTADRzuBxg0J8+D4l2tSlQZu
NeYp0U3Zzp33KFOFVHsulQB31YcUUhSQ8/f6fJyB48lM7tSn4B1QfLTKjF09KzNRxTDZowgusRsw
FlbL+wN/MjHXtQRZhaGPIksgacB03O/chAALRkpGrb3PWemWtkZ7A4YhLwk7EGyt8WWDACTG7tKE
0w81hrYXhNA1JJzlS51aWKZiVmlPbkoYnEQ9+j5Abhqw1nqiLjxjgkK/+6XT/AgKau7mdYbulq1A
w6ES7Ru+M9TPyzsfUyWql5yBza07yvwMsEVUo6z8WpyX6pAwOfCvRamv/ZyvwzRohXiVU7715r0n
bENxFkOZo+GFDQ4Vgg/vnUJGIhAFssOo+L+ykzf4rdN/k9mkpMMdqgtYXxIHY7t+tiCfshMoq/Mx
JPKDkAUxJwBuMxe+khGfRYWU0tLkJmW9DFMPHVyPSQss0Wfioje+kLyrzLWKkZMx17ifXwTvjHg0
/8zRXzqv8O7DXcODN/jyZFvn0W95nmERKSCzB4A9lcxPlORmTS3CohK2sZGaZPnGQrkeRNHM0IZ6
lyWCxSN4LfW1AMCOdHhRUMCFMBL1zlWICGidPsqw3XaYpfUT7QR/Ig9AsdyBV8N9TLboPIYv6P+b
FObdJ//pCEmhyT39tyDtoFgEbJvWg+9aIwh58PMGeLxVyTD1CU00rj+mqZImjf6FRAyQlpHC1QzD
DIJGKUfQDQoBhmjarqETDfM9NFPLXlJ+eYl8wvKPSoJmduAAfNI7j+F6jw+GqCX34NyUR6h9XcM8
OD/Vb5H/weBjP06jIeOZW4BAu21Vc3oeMKgyGLhfD+ariy1FYUkIyve1HtDi27jHCbYdLcRft9pz
rKXfxg2I+78jLT4b6EXugAyJpowQggHg08+FBgw4RlrshZT+7UOmlTl6ykg5EqBE1yCdKbIUaqF6
+SBiVLUvvbGowtyEJ7nLTBK9LIzIZaA+KX5lCf1MflEiBnFNHmaD8jBc53aof7keUS8F63PIgZx0
Zz2BHvYDcrOlYPtFcqDh1J0/09dHXWNMIYiN5QUXtjMrT+1gcH4kTl7tEQMauAssASPaehViG0q5
9R1yk+u3ECCbtFdGlOr1DTsL9ToWVQuGZh7+6K9P/nzo9gUxyweOaduugDK1/ujHLzF0DoCGDNo4
qOrXX81BgVjOtUJtD12+ROPp5VYBZNMXPA6HeHpbf41WQjdrhIk8q2ItmSAuHvkPaur+h3/bYAuy
f7IBiG7TYG/+TQ06oEzeUpQBy3Bib+bPTBQgRRonxxte31nvqk5qLGDM/UsILol8NNM+0H7cc9PH
xyt81MWBT4AmE/K+TqYvpUKhbYbzD+mg+hYJGp963eNlglPdCNrrvq79PsrzIaGEAi+mHfNJ7Z8l
W8MPbqlfn4REGTY5DM+UUJvkgy6nwvjUza4Vgqw/Xk64byRKcRflzf8kE2YtHBkIotAghrzcM5xv
Fb5kQHYD3v3+jRkMsky3jkW8squNB+aEx5013dYwsCmckIi0IdLotocbdJ1QKvzSJdBnUo2Aou38
G8eL960K+6yl/+RtWAeGBv4q2cSKaEkWcGy6MjPlYnqFiULDSiR3iILY29Unk3XcVre2MIw5+jZ0
bY5ww+k0I8ZzaBamio/M7iloDiyUerCh9Gk19jLlrnwGRpVHw8aOvCFAYB8GBg4czcPpCZvLCWj6
v5wmas8W2BUPsTT5C1q9RhjvZ2zRrOkkaJONR4k9dNxoe88QZ6kYxK0yEtLQOWuQqz9GHFJPy/6u
wnFhVOEEsGQfeZbv7QdCFWieVy3fHl1GiyzpWbinj+sqGriUg1XkHsW2AFQHDlwH7On38Om5XZ/9
/EhNMdRWQq2qyDTPqZ4KYPSyh/+f3ulMQ3+/pR+RP/T/+ApwO7s8LoJPHeatJs3JmpKcEFoQZv+M
CpDY1r2zKKKV4a2RxF9S7APGKpI3XQH8zWYnqe+/V7QMi8kNpruUUy/kZBVEJ56s2Uvzybtr2dc6
wzvR7cWWneVIAU/UOxROOFlRHSDsvGmLu23T01+uXdspKy8ZmiR9ydtMJvr+aeub00/4+SKGKuMi
XpzmYeXdmpcyBAI0FzQMHmYNbzhqi8GJea3/79Ez5k3YebRA7i3AuqWCcwwmiF2lnnfcEcjJVEp0
muWDf5Hw2em1EBwZipS5k5harjdwskn7BZ2Xp6FFN4DzhxcI7kwuQ5TqWZ2/aaZYcwejYyrBIrJ8
bbp2VcTl3vvy7GHiPyOw5RSJ1YQ0D39lQN1NUNVFbMb2B52uyGcfakBE1LavKSYp445BAfNN61/c
UOLyTe3/mO8va6v/dQe6VrfcDLSJbELu9NHGTamEh/d8VaU1EcOwaoEJObaBGP6dUucH5iOEneNL
J11Bzvtadz6inNU16J8NbtPfYHJrIB77ZGFfiqL81Chc/Yvp9U0GWySsm/a9iaqflDAX/nTDnWUU
ZKDbMT2wB792hCGg9XeIaPNIdwcLjY7Aa0YDffyQ1r1pmx34VvHfDVbNbI9zfFxo/nJxqjcnNKFI
g4t/Qz0ScqclFXE5BRST7sekyvhc3LqMEDHuJgytlb8ruAa8f6KyJ+ho1EODkMf/+GPFin+Wmi1y
b2vYqtjVC8lm8f5kK46TYtcgoPAIBIJR0s8ryWoTdbnxX7wUUhCQYBUIq5eRIbH3GEKPxqvmoYSY
oYM6iLSv26qVNBrKJijFDTXihe/cX06/+vHlDEV8249MTfe7m+jaClR4eNlQDEe57rtqoMVrGlR6
0kPyqYRqORL5+FL2OT9zCvHyMIwo+EHjEbfXFBX/La8A+Ng6LzlOlSl7Zlsg4woW0+eOe0AhHh+i
L4T89I2B5BZRNf8AOkzpEySM+8a6H0ovr6FjBrJz0+gj6PxxJok/arm6ejgSY3hNxp7f4XOEKUtT
6ofldHsaOcRVQejE7AYKRfAbld96pEmzfd8Cr4zdLQROmGyT1PBYzs8OY7ChKw8FHzj4dRe9khdA
Jp1lmOls0PFmNzDfG1e1ldrlGeUOFICLojQezugXdUyevyqfG6d2Ilp4q0c4rfkpEsCighZSZhGH
8loikMmDLio3PFC6ZnwrsoZuBsP8D0CSrzZM7A22+0dTNlt9k1Rc8j1EkJn/bb4WUXVBbrdeemxc
PEn1GwQjwQoGlad79tYJNaySxrez/GUZbX6iUvduuOff/jItPnBXyvW7O/XT6y5ClZiCC/o0/tvX
itPiPuU8RvXGkiKblXdM74FcNwq3NDrvAmoGQTr+EKYUJFIavv22vBUjFpl4bzWmiVLg5hYSj5IZ
ynlGedWYxAinpZtRJKtfWmAgwAwPMVUv4m7FTsOLDMvdiBJNV+A6Q6Y3axbmQbqy8BK4X5QKzaU9
DGI5NB3PmeB1iOI2bZ94hpJrDHVu2GbB+3BtvJxgbmspuvhYDaS0v7slT43/+PmpqntxP5DRGEy5
lgVkIKPh/349wPehx+ErOxHUdYsC/fc5KVm8qG/RIyyk6k/lWKabVPh9f9HPjl64yeKfk0QgqIDc
RHrkj50M2qoN4UAHrXFW6ywzYbpBFTf4gYEkT+/0MvUaRtC93LoQabuL3saMR6n8dt0JkUxQahAX
4bxVQCHzsv1uHO1wpgxWeK7TVdwQwoTVGFT6NoWt5cpI9tXwgitCV2hX5rh8pKKmgSPOsaxMpWV8
Fo7Gjtcn1U36iD+0B0CVGl1kjnwpg1Yze2Aw/U0nMg4phovuQtc+9hmPrlNSiyXQ6hH58r4QlbUO
/G1YsKlcqD+xbw1sckSncuOQhWq35eZTTyodVGE5NFQFdwGhCaVcvpuphRBWnYpi3M17kiTVAEak
44l40zkCRvZA1Nrf08sBvpEM9yVHYsHliRnmQYusZFojqxECIKjHfkQWkEzRNwYpzRJP4fmTASaZ
yaOSDltmHBAJlF/MGewnbb0csDV3fG5sKeIWizQzXyuaWYPh8rE8tF7JKmbs3JA26n+3BCekBXFO
irCzWcgBH15hmikOb+f6qAyKhmIpywYRSmHDbBVmq9C7cTc6d8DUblvkGQZTwhNXRI5yxDW07/m2
ixIvSUyAq8XJSwrzaSorBFFPstJz5mcQspxqOVfT07KjdYX+YfAMldQpTRFxtCcSo3kAjQ1giknl
tybIxJRjc3GGIU0731c52D9DMc4pw0DFV2R4kJLO8X1yAMza3khDZcNStMV4uePx7EnqmqLJ4Brq
dzQ71JL/T3fcNx2/Xq1sNFJbJZZZIzM2qA72Uy6Cs3pJHk7VLjcE4UnZNK5ZD/WBcEUYhxuX5MzM
NY0w38KgRdH4/d6BlcnaOeG/vDvv7kHIkbUIutN0puQK+Y3RpJubZHuzHmhMG6l2GW5QjGdfa1Fm
JjHEYvbis8Fqc+85JglnXfra/lC6ESXPoODvW7Gs6gMiKU+tJRdhULE/txSMI3kMK3i58UdG2ODQ
G7ZcFYM4mjFR9MWaOhSh0nv7z+j92OkGr+IanFW535p9rpbCayrl/0Qcx+3u2P8RA92HztzkL98O
x1RqYyhG2X/d0Q2RFKtxaoX7I16xikxKlfjC5zfMQw82q+Y3tEZFt1XucYkZfjeGn1def1V7jkaO
r2lNVMAuvDUjf9CEknQAlIJtZnffBL8kYv49NVTFWBl4udxDtx0A6R5TH7edf6i7a4bmWSDoHqQz
IySZ44shJnbUTaHye7M86gkB0is2vbUq7QOVKMeZetl4XzPiridYk1QU0yVjhhDwQOsjnxjlf5eo
uYTO/OmI9wM9xqo/n4fPphcoK5C/DMkmu/Hg089/0X9cHX/XplQsSZtwna/SVhxoWbI/P76oB2vU
QuRwOJxk7IUpDLOoK1B9Lk0t44ItSBpHq/WS96hlrYIC00bdhOwaSDayUXJ7ye7r0vUzeZy7rP1Z
EXZxYiWDjKDQD+zKciL/p490gKbfODCjZGbVNSRlWKmDBIg+W/JAzGYPkiNH+WxA8b3VKUXsOH7h
tvAQXmU2JZQX2BV/ua69jQlfAgnkHja6hQNoo9inAy+LwOGBB2OdcAw0YGIeRGxgU9KZnUTnu1BV
7FmdhOIF91fzHpv6NbhkNv4onwpw47Xa2qX2F8jHW80QD+XqWlonNBPVRsnncIbzF2umMOaRBgsR
Zbv5Reb5lwEfDPNW/HgUVkLmyxPXTsMkJEyTsoZxUgMJtTrJcIyF5F02dTKWgWKroJV9CdPJV28D
eSrSgJHLV8kjxMnJ36jfAElROQ042SpcwRUKbkPwsnHhcWyNbggaUen29cL/byDBKiXvoIcfHnP1
ALlINPz+WiILfJSLvzf6MWtPNme2lNjDfQCOEKoRY4ur2f+bRkbaLN0AKdRAD1gU0fDx6d89/crP
ulQbaqG481M+VpsGt54eVTHKT5PG0jx42nH/CbTNw08Vwz3x4LHkpP5aLGlbBWhw00Z5OZctZXF/
R0wtKbJwc6Ms7ubUXZ8lUNJYX9fbCLI8cSiwfELjmKFfZbEq/XaqeI5T9ZBIXz62iPVoex1sPAko
x/PQepzsLt5BH2AwfE1VUr4kwNNoESEfbC20WHPEmLuMe2+Qh8ctYW8/S+Q2k5eqnklKunpp5OUO
d/lFvldsUo7JXAC9iSF6b/M9OvQSYiBNdoK+srgOefPwBFQUHtTuPltLOnZhAEeOs4CnOCvnzujt
+y73U0P0IpTyOyZWYchJpZ26n98wG3uM29A65nkSI5HJfw+qfIaMpYSpXXKrGEgbpQL5Iuqke+uL
q3ZqEx1d0bjHZeeLAPOCYC1ewVYfeMZ6G0cJerP/sybKeX1cbG48kAfGgl63cXGuCeCCgvnxlD+t
stXpS7tUHpd/trx6QijVOVpez6A4vDDUDjUgJPTp6aysoNf7fM3aoLOdhiyJUoRtqlJXufewL8ej
1+gxNbFIaawZxXBnte4pmK8fcvReK7LlpvvfLuGG+8Pfi6xjkJBvbPwo6/CTHHWsvI9MUoXY7gC/
uFBSBR7fwHvd+yo9mZZrCdCa1HgHB2g+p8xns5muZi0/EXPCLKt9q3l8aqy8PatDKebHJzhwewvn
GbD2vQNtMHK77CQo6jd9233NBEwanNrOk4Z9CZxfHH8DdWjtsOCOgilx+5GYMG4srgqLMnYGGhrf
HkQFbHHnMyrDNWg9TRECmc2w0dOALQ2DciMbYZpbptHqWkRQRb9Gdbkm4cJSI3/eUk8w9BhsWzi2
3AgFnH7/fVnA5GGR92bMnshvn4MJ5pOnnevjpHHXPF0Y7nMLnyvCn/YFCCA+U8+TbtScYiL2ltSM
p+4bKa0Vm60SnDxW98RuLWv5SaN7jtY2yhiSSJvahbGbn6koJHuTtT2ZTzY3WnLFIIpVn1585VGN
J+RmVXk7gBnyZ5nvv98wqHA8yVWil1v7lMKU/5LEox/1fB7FempjfYIh43hPy6p7hwPLAnRyf7kW
DkQgQK3qhLplTPS6aK0KGL9+lyIimQqPwkvA9c4jiCkvx7Zw5uRy7JNaz9EsMDOGN+C0PO2++mwS
p3t/25F3xCSJqr478xshrm+sXooG1zAx1DC0ZRB6+2rJIq6UubKGry7QI40zWr01uuEaPRVdI4Gf
i6Gowd++FS1vZmtFLctnT7I6BX4NSPZIrPHBi4WmVygvK6cTg3l8dqNyPq8de1Z+CJLZXV9Pbhb/
1iRE0oRt1SUCyKuzGNaLl+VPaah244S9R0IbwDPPulM4ubQL4slpb8q9cYOIgQ+HS+1y63aNhQu+
N5XcZjybCmJhXlbvLztmw3U22N1z+qfh7TlvweOPJyHDXkU7TY7g/NB0lynKRObYOAqWonm+xZgr
5V5JJMfZ/mEIv9GbtUmxD+LdVrMtZh2nTxrJNGfzdrG3vzY8HVOmYeLJKsbxpLEtjewFaHEaOgQn
Du5rbP7GPybJg2lqqwaVnCkFBq8jgF3DwqUlYBYHwrIBhItMBrWDqQgce26orrlZgaduxCKSsjsU
YYmEbvFTgyURau+lFqVStkR6mYk1Ej6rDLAzUSFWLX0MROJM9Wl/tCg2jl+CPQoCArO2DwpRCwMF
Q6CwQkF1EQZZBJtwDUjyVRLZ7PwD4Mwui7CoMi468fWxh+z4s65GR47QsQk6faAwnB9a5IYfzEks
LoKbnlhKYsRyck4xI90FlpnrsILLBdlG0HutjeqGME2H+3IiH7qS2xHwr+c+37vqIk5FzqnWg9vk
Nt9hU469jryFwG1fhReTnM2Pec1L8wn0cL7SCOY3LsLqd7YnHMpjswrZhfgxcqicF/gQvRIRaopl
atuEILhyWPet/y4UfGZu/60gLuNUZKQukjFvFwRzdmpSCyENdi0/r2w3/vIH9p3IMiaxqhLzTVSr
lzV9X6Sun8XqgxutKaCnbUj6UMsePWXY42WTj1w5fM5mbo9hT7rf84r+QLNGOjMq6Cop4ZH7SZMl
JbdYH1E0J2VuwcesGriZ8oThqTkaxnAck456IofIt+/pV84ylzQYck4PNifHfijRxfSqT6T5e7sT
YsjLf/Vpv0wlYYsPYbqNdDbNpvKTPBIZ5x+X+VU2/ETuqUT0nrwdUbLNpxOlapZADd0shVHTxgor
f+Uzf4JyFtzw6ezqAbdP8OHoZjy+b7qoPsZTCU2oOulUcuOOQMI8fayt6H78laRIhJA46XdlVnn9
miPSN7NKkW7qOjnO+UFMGPvuXWuQH1A47SxllP7QE2Qnli0lzM5Zov1w3+c1rTrpGDnIzZap+p1t
fjNoGuDKg5TkfVM3slrlm0gZsr7DkQjS3mQwb9PbB/ScdoWO+pXAegofvol5tsT0sAsefdOp9c/f
auQjstUnj5rKnp7CIdQbIu3uZ0iJPU+uEcyjzt091EiqJSG4FucYqlj64AkLILrmx8xBQhJyEUz0
42oEEGWw3qVv0YO2DRYC3a4nkfXox3LLKSjeiNMf+9WLh0nPqO7Dux4OkSlZnThmCj0mub+jEXJD
MK9e6jWg2PsESG7KmuGbUL/Crw+g5Ntq/ubFgTYex11Im/gK2irtd5KzfNs77cV8b50daeCtdoOt
tVlBOFuglN5sLvFKtion8scxS2V86FiYaP6DGrpczEKj+3LflNypUNF57xiV19QreIiHgWwCRL1t
NlMj4Go5IAbs+EVsoaILoA4SD7vi4CAdHZUUkWpHgoEU7tEsZP8otqrzCcBTInrePtKtNQ+P6bBE
RjQUpgdd4f0nbIrbifqAXvzijcM01ci5CEUd32oo1RopK6zoUiUOVQ2tde25Uztzx1So5weXQ4rD
a9g9tMniTVyBstTsBQlF72pXi3Rap1SZtIeCA/PowOL2+5DVceSJA7iy33gxEFA/NpO7LlC+Xl9K
FYv17KEMkquAqlYkIwV7lOzlEaBCZMQ5mnwUG1KMRijgViFg3sFx5MNj5YpYOA2Sd8xiiwo+FwjJ
rFnF6HVC19layy87smgw8+OKh5cvGhyMKw6RynO1wE4JVccq3pbWZVdfWVSaSYkGVu6dPxcih+7r
JD6Qx6/rlzG5dnjGvz/ZhELZ+P+CRSLIRB/hxrNRrihhm3YwCzozeFzYn3fopk53aLQZF1+916nG
Q0Ss0oEY8KXe0dzMWiLwtWsSbDXET9oj2RR0vWW9KASuw+eGw7ejX5Fmei3RMezFP/DxnsF7pdVp
qT+ZXyUkWoJNoNixoCj4Mnn59wmXIZRqcpbxwu+1dWuIxTydxXOK82kKRv17nV5OVr+YU4j56Im/
B6XwbGlyxddxtyck2P/GPS+vHrB1yZNILvsbMsfS1e8daJRUABPMTArX0gykPPKiMRHhnruwAfBq
++IUuJOKg4UI4nF7dy8cU1FdMnBkPiTUoZ5YvulLHVbblZjXxnadrcjSDJXAoceA+xZQyoth0ruC
0K5o+EL0K4XlCyT7/DzR3mZ7Yrpuf02S6UDxvlmkW1VuMcwdDRc4ng1YP+uslAM/3MnDqBB1mz4o
gGrAJkdIT6vchhlPrCFEu3y5GHAdQzvLqNDCajxX+LuePrc5Khmid4IXJFucIFrL6hXUYlo9uGxH
lpqtLju+LTTA/EhXdhrXzkQTLAdl+k0gAZjfqfEF5/i7ZJY6yS0bSwTr5RsW27qVtvNe2Jr7thC0
GoFu3hfoRMn4oFZmMC9rBJ4HcJplggIwP579EaHhUPhyJSJYYUfr8ojeKuyky5ESaLWGzEIU2HJL
NBzvB+E2Eilio2ql9DbJbpx2QuWDX733c6Q6FK/sXRYqj81TqdrBdB3En0+ZDsSASNoQFTAXHMzX
/6VmrW18aTprcm8/11Le5mgowEqQbN7cj28Gwy+YLaODj28F/TQIYy9l6X9/bcWD4XnKD+2xUpiG
GssibOqU1wW7uyUt/x9UZCxvsb87Z5dt6SQ4Kqs1HFpPieZPrOyKD4XWbYaeLmx8oR4vuvGIjRPa
vzh0b1ua2efscG3V21upaaU0/BfMu/WpJ5H9aZJLjycCdXOeY/kBI15TbuqAa+U0mgtH8ZQpR6yT
27xSoafHuo/h7d41X2hGXr3Z67yk80YaTYFt3ndsqyRwoNOYWKrqafqjxWAymgcJbbbiwxLCzYPq
zjpBjAQ8/UkMfGA4qb8X9f+2mZKdRW5jJ97iiHOSJOdsjLGIPy4NTz42sxr1oxNyzWZ7qCa+Yh7w
mR9YR81dWc2toMRNdp4aLZoV6R21Ekeulqg1uEvuaESnPiZnT99Y0B7VlAU5GAcndaTHsKDYq1U1
+EvEgIQuK1ONlkdFH69ooMnktItJN3pjEpu2VDLh0KxSyfLhaSo4noDiJhqPox1KuNmCRTPfkb/d
F5fKD9VwodN1j6TpmgkfnR7oB5YoVJVawnCszLakuv6cabWQWy8y0UeTWs8DyDRgDSrfQAo+OX7B
zy3iILdq6xTmp4JD2eVV/htGGr7fC6Uui1+vXE99azqVZw26ge5+JDxfU/cJkoouu+DV1aCkgaTF
rCaAfImTNONY2wZvjofWa/rKcsEleiP8OYbBG2mzdK1jBsHKFPYmlmhbvwNarU5/qUxZn09zVdO9
n6xE5rsQG6yacbRhe9yUszFjtgJnKyZ6Xfp/IQ/JobKBsnCaSYS7hbRj8Q7a76WKzks4757X9y6A
3LObt3dujAEYzRHli6/hUTDnM3aArChXkDUhdTNQJHUjDypuqeGkk/qTtrzmKCsZkkKzRRR+ldCa
4+QvFHueso+dMg01vBATbU+Vd+iRdalykatdTH/OWAF0srDHvzZNM9O5aTz4miym5uYtFVV0B9xo
pkishxoFmee5QazeRRDvpgiiW/cpLgKB7mjAD+hDA/PmDdJ6BZUbScakauTiSHov/08Q8iBHBTPE
gn5X8LggftgEJZez9+A66j8bCiHxo7HSVfQ1/USDBfkciEfTwfAKjhezA4hCcOpObsimEFFTQsM+
W4wbXjhQe9WlSukP6oRn7fmW2b59uzc0gRWrgc2Z8KnHQhigYsedHlIMV55CFavyoIGuAZMhBnKF
j8b3oMvmXQGL1HDt1e57Xbf7L/tnegZYgdc2l+BCVoMPvOEHcvbjjvfGl6kQIwMBxbAybEBNEz9P
4Zwca5YEHu3TrhlVZHibG0i7nJPJhFULBCwfKoRx3Gt/6OXvyBonMrM7ZlrkR+bmAKFfMLwKNCGR
rfvn5/sVtRCgrrNzO0gWiP+MKJwQ1n8k6FVMC1Sng/M4mkyvMPubjW4QTNvgCL/4yDs4yrrDdRfs
a52N+iTDdB40Px2Q0y187bmzza4bV0LIJLQcHLuLPzGqGqPeK510UXkNOGgdklnTxpWkJU9lt06s
HqySzW6BGHD9GyLrN5ilSaK8gt5H/ebU5jE2OnIzg1PnuTPFQJ5sOq8/Q5x+kPPMcILWCZek9fFA
80mAFo88FdQlrCDa1zLYiHpOdIiH4Mz+6BfR1b6gbremRnR79v9B75yWheh4Jh5cfZhYWyA4pQgQ
pSOlWOQO3R2NMKvZyZ7ChUgvEgOjWUTQNz6d8rhceROSQXSnx8Obv+2z3x1Bqmo0jnNhM2KyppAI
/oCe8R16w4niAI0S2gNMh8PEtK7Hl81MiNEsC3Nfkw8iWzu56cIfmpGrpJHIkDt8uYWYCm1WFdLC
ykIulG15R8xiIKRMj9DYeakEWj3CqTbrhGca/wbmt8LGBfHUW+hbYNvfIOLyTZL+Tscfli3u5BmT
IzjmBqRXdCXr8Kud7QmNpvK2CEeYWHqDlosfEf4KY4Vv/Bt/RhZ1Bd2N2wUxFsrUhnpyebCxd+qa
4rfteQPbcj0vLMMnVROadiCxcYbiaF16qWaZCTt1qatzKk0jhXsQEQOSOOMpgWXogoELifPygi9r
0QeckY9LBL6c4BhBoTT6h0glG9N/Y5U0i5QN5McQmULLHO9WjXl832aBIwr/G7XtpDON03TKuWAo
Hq2rncchthLtP1xBtwg39li4MFTSO+5bpJ+OGKcj1A9mM1YhBxD4Sg4/F1xE9NvAwOgPXwxTPg0G
oDl5gPzPVfXVinyHYpnjnPNEcNxRQCU1b3Xl5gCpc4Q9Geuy4GtwSm0vbn1nBhyud6FyOiJNC5yw
820wbFQTH7g7kKZgziIEz4huAEeJXGdoKyEU0ntyvIQpCs5lsj/+sOCpil12qtCFxjX4rHysTMjk
G7c595UO4bVFw97Dr669ZnSy2Ylc/zu7eJWVHGIyPyErkhiPGp1rTsFPRBAe33A6fKUf0VBQazuC
UznT5dOTE8z10gzq4kkDL3LLEu0c5uI93oYSoBdNrIxVogrIywhGsgldu9nflPiHOLU89LLuP+AP
gHtZNKSoAoUhwbCXxmo0c66mPPfjr64DK025Zit7uOzSOnph7dCnsdu+OoNK5ETM1+p8nyORHfRb
0NPjW7wJC55RwKn+lBDK77CUukGZdcpLog/OcdhD1B/AdFrN9h2tJ9Kb/nUBJK8RIshB2BRXKYnU
StLVmkoO6voJukDwnET77nvsEcVlbYThYHtaHQQQxxB+ux5Ba4C/0JDG9gZQ7nxlg/+/mxJ+vPSf
qN0L2+U6EL+yJz3zN0ZIr510zbozIWl1GIGZ2fpcQAK0A0655uJvDvF0JJtvM9vD1NIqZ/XYmuU4
JZmcEUf+M4dJLxyOjjsyf0WUat8Q0bUd0J/cb+bb4JVtY0iIcSLAGXbzPS5gMwqoyimOT4C3RFr5
+qcXHTnSMtIVHaYy9YnDLg4UI0FZM1b8KcuUXBa+d1RwMnFQVUhPUQjIygvHNOi4Lxxi5+WEIUdM
P2GQp5w98FIMLzZPWtYMYpcUBrxzu+C5iJwLxzGYBqz58UmJIQAq4kl9F75gzW2//P9Tcv9IvmlB
Y0Tqlzr25LrfWu9H3hxjHX4SW9rr7MUM2tQAjTiDEzD0t+prnRR5H5+Z4oXChvoWnWwfm7BowbJ+
CYUwhrV7FIFHKPCasT+UZHe1odka22CLrRhF9O1Cqjx86rD/k2tjYCVe97txWtRaJEJnjeY2dr88
avx3xKe803DcciZSxkD+nIEAkCf5z7rpH0+4z2p9rCp56u8kS+9zzE4vTAMUSCOLAjePU5YzfKQF
AFNaH1RFE9THUvXuRxDpg8L2bwMpB06jMX+cEmRFY9ck/Ugcu7ReY/vVHmW0gc4tMIiK3tEGZYVI
Ots1uu/eWHgTPv5Qaf+HR9p2fwMJ8WAwqVhXvUU+aCeaB8SoZoeivmZPJBG99kfGYh05Z0gLLq4V
hssAazGgQVPeDeckQT3KHnvJpqcD6zoAeEa5MVTLDjWxc0nyHHiXte2ZKGxdrDbGeCVAcdtpy59P
4ZH7NIk/s9xOZ4kmXCb7cVNdie2Z7nF3uDqQI/7tfq4VKfN/1SS1mFO3wQf49YXs1MKRqgotYWWS
qEmDlbuFywKVxBUb6dmergEeZrfr4+Pp0dNAvStQxEDo3qnru5gepwGJaXdtUx/IUVRUsHVEkdpo
2765hR5MLyG8Wcs4gRNKGvWtqE6QDK1Qr+OLa9IaM3gBhqFJMCzEHgS11Ami/yj+AGuA5f6xTSAD
uf8+Y1jDdjp4PUVvbpJRIGFA+yWH2dQS2RiYS4tACXteyoh2RV41dJTB4BzEDJ/B/Ar9erX2WV6J
vhvofNcEzlWLg8lUEVvAGxvxABy5QPRtz3rflvfHFBoL0gXPRlO+lg7UkLUyXwx33G7ppO4pFfUu
vujOTg5EGmn6KnHqJm/TGvOsjaqMw4tGuKw9Yb9sQuUzLWWvL90Oh72BCunxoL9kW0E/FvJIgjCH
huowMCaM5AfC9jEfwIfLNM0yi8tHOJcW03uckCf9R48Y6oYJvAl6piHrlt+5neBDqYzkcjXxVMF3
DbHcOWEK14nDg6w5Y7U6nrkVCYN4H3nVsnasjMIbTTOfT1nqLcnGPMjIHWfbe/boTy7Ed3MrIfSL
xYiiFJRF54iRAd5qXwRfQ044rLstmSrdutTGo3fel7UDtXWMsG6A9vzbDS4VNnqceLENkOZvoFb3
e7xQkgcesvvAfIadpUUVbHfu+sd+H4INUZ/kFGvfpK99gmLaH1R3ouK9F/ImxW1wwOk/t2rHE/Z6
5lY6jC+Ec69/UfGJq0RruK9ZemXM8dAyPZPdtPlam3QQ47j19zxCdXswF3SdKJPRR/auSjIDQFAH
7YFxn5+WQ3jxiherpMkctBn8cv3qXRBaJNipzbscw19KtRQjHaYaZjUAX69mVDM85lSRs+YaFcHn
BQ9Dh1K3/Gp20GHkMhjQMD9xsEsdlB+jP3dZsUGjNemR4BrLjCiu3t78n2shsmq/vMdBMK7Z7kIe
zXFKhEaFD7SfYLv/QapSEdvRVXvaUO8vOFoZn440pp4s5cC784msZrwzGwIkbI9bUaQL4VrwXiJe
obufHTgfDUSZE3jJ8HEpgwgafOXMKXw44PcwpM0tCe5ViiBT9LKhuHPnRfY+quiNGVA0FY7pSBHf
EiashtM9gtyM5galcpdMVBGXTezoEWh5UPntkI25JU+7+sSSVbz1+1CNc+4mcc7HK4Hk9orKm5zZ
nUbDmOobkfNt6QbXjH6604FkE+MkI/FgRTofHe+Htl8drPBqtwCUH6W+hGVmxv4m8uhU0lg9scS9
4CVvUswIdNHNK0EWrauvJqiUEIkF67RrrKoyn3AukFO0+5Vrhr6zk6N9Lxq8KcjD2fRp32V0hnQ3
nU8LS0gYkF2tEXFRtSVr5EQ5JcvTX/z2W2NiVI6PvAUt6UVwAIScGc4IKiKL15aQSsLTy1LslZ3I
M3Q6ntUFgJ6CUMYZpApoyljheoZZ8s76Os6lWdZ68cmI+kLCFEPAvAd4OUP7Sf+XUgBlDGr56lVG
sB2LHolMZLqlLWG9iy+bpxXF2VPrsAA07yNCNfWqD0UAW7oI6Am5cJ8GVwy43Xvxgzm8ipTib3cd
N3oXYXscr21f4qub7naeanJr6pUHLWBYATGMAZPfam+843G0Jk0/CZEP68ETtWuTq7M4S72CXmra
3ovxHd289dYvqsGuloWvXedxrv5K/JJJ5rGFt+T0TwVJVapa15aRksLBUQ/PssVf7qK0iGPer8J6
zjZSjwPCLEW/J+W8vrZ+WCBvYM1wEvgjJ8AJoXJV8iiD6aUOQgr9LJtjyCJHPHcws8Q2+BRnbOSh
JTZ7+gWtDQLULkgXm+4ewyheovGCd8+lqMThTk/PoUMWxI6B6u63IESqq+i+oSQJZXybx6qwSkOU
hGEW8JfLBAVP3n6ykPRQcLn/GluIGutfD916djMNCZx8PSYM2M4AE8TFEderC21ElfNmEHGVZsVD
HIEarbdCZbg2/NPjNq7FwMWRqAG0wLbvx2xkurMMcqyk5cx2WnR3qfarytlnv045JE7VuXaT0OEh
HMnXyicBIdwk6a6ywh8OrWR84aEC4qEJNTLBBB8I3sec0h41zp/JJu9Xy3O0DzNGb3FwIwgADJkz
7S8aJpNyr8mVUPZi9WopZo8yG3Jx12Qg64OsiJfwV65dkxn6yXSOTynSzgi/CgfUL/PF+K69IOIk
9TJl2NV+dgHSrxUsX58R9JTmSY9bpm4bBS1p3v3183HoqqMi3pNfZy7K1uCtmBBpyaAw7tZx8cTg
hrbHDRSmrXmghEAIhGdx4vR3AB4HAlmfd6bUBPlwRwNq1Knb2njnT8ueKuDhylTCcxrSB20dH/2C
IZeTRTkuvOcMA56SukGVbRvbtRXEuo95z96bhTQ3pw5iLenAONEWlP23BFJjkrZa+MDUCPQMlJhv
otYliwkrBXkC6ccnd1d0v5ITVQGhApULYIJQ+AirnDEoLZQ9+pNwGwgOH5P/F3VQFeVeIrpFIecW
IGiWngATA2ZNC/ZXoWFCBsn1gdF9IAsT8qLFgfLO5czgpcit3JnOIFK5pguReBQkCVjHNTn9lyh2
hvgM4uCLHCF1mo6jms41ga4/S3J0yqQ8tP2+ibOnJsPIcKSIFvXXkHyl4ytaWpL2tx4GqgXXELw2
JBxAMy4GNZT2n+6RnRxxOjo5LfBzI+N7SykgzByedFRtO6xqxltqMoDiRPwGlthUEmDlAjfRsuJi
YgGa3oJsBsSzIEj0nASqNN0hzwe1uANrc6bCEUJln3qqbUU1JnTgVYKHfw6Njkg/yKd/RDR2DMAt
cwej1ycgp3me2tiqSc/EOZ1YJRGvMlvzEckMgeIFyYw6w9rQPTZXLv8vTw6FwKc3GCZfDP0Av495
GJLD3KL76ykF2QLMPuM6sk5ou7AYEFj13MFbIvWOX9wCNULP9rajGCi+3KYFni8V+VQiyr+jQAtN
Q5sPSTa0GtIlEj+kg04TgwxMfgNEjbPQ6/9Jik1iXvGtUkd4QrxauGxlRjSEPfsYlrpZFJY9cROv
S1yJmZqLKhBaPsGp1YKdlCxRIwYyatMptYPm0UYEZhMDiUGFE3Sikbi9o3BT7CmdGs5GL5QjXYYw
lKl1xTu3V2QbkG7prPvIQmtCFuXGjIvIq2w87j9kfPJKHV9mTTZC8PYg6LYUfCSZgR/6Dui0RP8I
Rsh3wHzhTNyeOky08EYDMO/o9axEdfiWx7bOW6qzS+IoRrGCadSyZ8C2VLKa89afmBjX/19iowQC
oUNCs71dC+Zj5+B7jq1qdmmxE2cO7giG3OehytMJduJzxho4wvjyTrS9jQOUpqyMhfKp81+MzM69
aXS6oBUTwtTL/1AHY2oZNpXMaJ0+0EVBeQcd9bwD5lTZWVLUow3hDyFXvJYrEQy/IN2vsND8+LfP
aP6LrGr84cV5PqPv6717edVLs56H59TjoAemD7PV0LY2QbGPofcT2umImA8ttJJkexiEburHowAj
eYyRApgyQ8i4GVCXZM3lm4DtYMArQieFXvJd23/p28UYQHyyCkuFIrGIn1LgPiVvm5vHffiI2EMf
S1x43e9qARNjFuqqfxM5ByTwh54HQ4pTRSfdFHN0H6dpekLh2pwqh3DDFwL7TXddLlj/v5lWtLzd
XbrVW1ZyxCrBq5Vz1BmgzEXwMqy+BKRJJsVcHg9dETJFHFC2g74UJ6xeflGdFZwtu5tDocWNrlSb
5vBylxE7dcSPBH73LRrwp3xx/otd/ojwfkV6NJ27+npgsy+lW2e9g3C+ZI9pj9FQuyfKb7A13yPf
468p8+tSfHzqCFWncV8x7rKMTZDubAtlS/OLD6ljOfF+lc/y7UDTvDLOid4y+zPQrYfRSfyYqvia
giu4dlkKb7fFcv5eMJYeDgZ+dZdBHVP8FEZEfYHEDwUdQuQ5siOaVN/Xbru5cpAHyzwV95Li2wrt
nt0rqJNEbzF8VhXnyvkzvM/5H5VYZBqvC5QakDKg2Q/YBbDxnWukIutZnxECcqpgQkh/VbDV6BVq
OhnIWMxVv9Oq2IN25xq/QRi5bit00gZ9yTGetCdQJeiYjcAL1EQk2AFX2aquQOqb2KWwhRuWIbIT
9SxU/fGVSm+hOevWQfttS1ix//h7gK8PdDhlrctmrcOcqxjKaGvkM0Mtwgmt69oCJQ2BglzqQxRc
G/nnHkf/Aheih0Zrk18nnkzKhSNYXIR1qq4MumDwGAoSNOrPp/vLHmdjgxleUaSUnfiIwBpqUUqH
gMJXIqeC3IpM5s0+Wn11ZpQrTnS+tPnGVdJV24KM6qQXrUrObRSXom0xgKE/x89e8WkO2BOTTzIp
u4EKqRXgCQ64/BbXPxvopwRJELlVFk5M1wDL+7k7AtSK730eNFsJlThcQqhF5KrGDKF1aDt0gV0U
0kKPfu/wblsDZR11cNI3uGinlJfvFfitYf16RWaPTR7Xe2YLDx8BiEAN04Q95XoS47AWyXni7ovm
UbArbwln5wJw4LEleKCnfq2wAZnbTOQQEkFfC+HvC/Fpp9Y67fUjYyvGNV+i/JYmTvnhFCaNpVxL
xLCt56hVDJnckxjwXkndI5bgEpv10+9K/42Jtf2VyJ6wNN9GjVSHJ6oNGqmaQmHP8jSVcGClFzAu
k3YWd8rIkVf0AC494YuM7fT4QRz6kDpb4XMy9xYvSROrqlwayxp30DA3koMLogYwvT/iNu8+pKKA
TTx3LI1I2z5OWk55LdRtsruoHgKWuSHIPfoKlqKiime5/siLNhcbZqsgOElSn4K3AuhlCMlnk9LI
S/Zr3VwrWZMMPJ6kDBhaFam0VE/ZD3iSJV9sneVie50bhvXIVAiKFGlU2wPkOqECBksIBA0INQNJ
a2L+cuoIGMWYkldkfe1ZzuGtWxMpfOtONDsQNUtix8dF2zrDDv8XICk2gOby/mEq1OgkSV6cwG24
UIRDfnxN38EdP2bJwCfJifrVrMM/CVbV+K31wEMpXmR8/wN+hNt1q0CCwozCNa7V7Dajo/JwooqK
pRIsCRnuwJV/3bwjmVf9UICoME/RGPg+USLTdepz50AdBlkJDPY/YpFTdXcH5s+TlUpPUi31xjD0
+qqV3Bz6SDCHfsZHMTm26zutrFcupOE+YTsjxWwGFIDJEMeRFr0bngu3dltYwlNf2cYDnyqxntOh
dunz5z/QeKS0Fwxog8bGdHR7pp3iPWS1nJae/OPtm7FG+uSyJuobokyBLs27broOmm+R36p8nkdw
u9h34o1SNOMyeBwBG9Hd8BpUHz3zmzrmIRztQLiX9M3mUE0CyDObbM7I8BNBVVhl/1mQO0fY5SJq
Aru4bm7tfHITQTJVHv9en8GGwLltQL+8dlMKKFpIPJAUmuGCPnfjXMz5S92iQmwcU18IujL4QyJX
odPSJa5c3Onau3Lv/F0d6PXYA9jGIFUpDML0LmiY9nZlXrkeIB/lLbJwvR8rzbOUJ/IM3ipQYS2p
G35jsE+UuTMM3uRJngPGByrNH4zQbESXLXaYD4IeDhmhPJjcNNFmNjLkxWYBf/8v45L8RCODAciQ
hwjPy4Ktefreln+WrcV8zOT1ESYlpNb0dOsjxifF/Qamud++mYfeGm5GMgZSOTE4OhYrgiBGpn1V
NJTdqZqn2WObfmbHCVl7tBOTp49Ca/GBHL3gaqToqFVi7WcgV+Tlb/XA2cl5/hIHy3mJfg/IC2ex
uf4hnX6ykrfwhxnzcVvDnPcfzI+acZ4JC1Kw4GYrZToFN1Dfu/3A7Jd4aU2LXV+WSijy0VFzjkfr
aTeE7tnknSzcZVi2G9zEJ8wvDkjQHPuZf6IRVZnpuMAx8kWBBK+MbYiblcvoB1Fv3nIT8WMgEP6q
A4nzWIZfJQqSMyQ+lgJVr7ro+9mmVBVaeTa3NOaXDcGQ+fmQUx7LQV9IfaT+mC8K8TW809Scz9CH
b4CFpFIRqmEve/ztPZ1v2EktlH2zqEu/7uOjsDTOxvTPKR2hQ+17UlLOwqJsrSgk8Pd8xxwgrF8X
OpBtyK7XgjucDaH6uidIDDh8CpolaAXcvxZ3V6KTH49Zd57ZRgd4vGsvFhPU6x4I0cqA5ku2r4kT
a1f59yOENqUW5cabSk2ZvMR4g1Vlk1wxLl+l2kubShxOq9D8yYguexioY8LZccH9Wmfk7rwbNzwl
kzGLswLf2qznFQ2lmlPqbo0t6Zne+VpOFtjCXVL1OaQfS8fl5o3nuURE5+CTwcNHdgnazu9mvbSd
3nesPGe7hX3TPu0v2D4hOE43FGn1arE88cvmCvJdrTgDrMUlaozgSo+DHCMVyWM7S6N1AHBCxyss
btb5gOPR4CZ+044XERFC2dmmPLPSH7wNyEmkncnW9MXKXvw6rNn8nHEBEhNjHwfPLvxlD/HEpIwB
ubJJ59n5E9qfrEYaH7de/ncJtTxy044xNU3BovTfVZ1Z3GPRJ9YRFFZpPgDVp3AF9N41LyEjJCtK
I9nOt4LlE/RtamuP83iFHWzZdt/iz/+odtPH+SZIijSSRjoyeC2EkxZSjd7bFtjkBdDCjsc5yzHy
6gWa2n+VjFqnnOzxSJLzYKY/0fv06ogfWa5o8WKrkChjJKZoIA5IOI81e32qF6kxioDjjwvH+7iX
Iy/RpDJ2OnmVQDTP7eOAoh5uYZy8sGfqex7Gu26uwzzS6N1ys8AZi91nDUpqnNTlDr67NStC0ZKZ
LmYqTZLQbBJywTZh2lDREKa7OtAMIk9F1pmPq088wDgPNgrkLoPj4qs8UOqNy9lcWV90TfqqPrQ+
HQqaGzE1LsAhHd3RgNLVnlnlFxyPeX8wpm7T5Or8oipBPQLKn8h3onKM8jisC3XON2K+IkyvWlSK
9CClb19hwnuctO63B14skafuRinEUcmE/xgR3TjBHcncAbqyZGvg8f817wy4kiKTZUVKDWL48hxx
aP2AdFqo/RraGPZS2djfityphA/Oh8kKLH3BLCt+XegJpeOy3Smxkm0YQDTnbNLOkR3st5JQidK5
Sr7Qh11eSW+XVVt29sR5hC+p1ZvsOJHiskBUtlMdWdA0NpxRT8CsVEXaYUto/1hQ5UPCJEFkOEF8
QVERZNK3txZ64GPsk1xWTE0jLzauopJHy6+2xZtoByd7V2dyJU8LB7bTkrNInRqwu40Hj27W5r+0
OfxcaJbb4lpHkX2SOqwdL6FvzVzPFlIh3VmBUekap/2sh0mRxIbwipmOCoI1N3BefADq4Ordv4iY
WQ5T6PjHnwvMVZS8OO+tmPx/aumSnew2S/bHxR4O1/4iQf9lkXlIaHbORmCR3iywuZ2fvs0pjG59
zVs7TfxoJeItKtdMsINGDhSbWHbHg2OOaSlTPxIL+lSf8JrL0J1ydWnqPXcD8senZhwkWACHu1V6
1h3sqGJuhf3gM7FOvsBVMGK/7BBlkC64WWSjxcGV8w64iDaFguqYFLPEqzDrKs5xhvLz5kBWWqH5
cT1ZMhNemuhzx3EN1nsggtuwbD1EO4m2PeBPeKD2hRpdAP3RI5h6FDXNArhRV+J9CAcfGaSZByFT
Pgnac2POABNODF35tNkNnd0FKedxvPxwfIuXW6guI9kMoh3F+HHLbxiYdTLATtXM15157kS5WMIA
/Wb62ME8z+pxCR02CqRnAkNxzsR1C7eLlJrbOdzW4iqVkubFP19ar16MpQWswXuPVF1fnHUe7FVW
E+SPft5X5s0t5YIysQXZvDOICHxFzyowOfZRZi8ca9BqO1wF3jfbA0g8xts5rVz3l74fwZINHfiC
1fVAYQHRxg4IP+X/N8vSAXLgAmguu6eF21QJZQOEaPZv6TxjQqzp0KdUPXRO5t5yUTxFY3M0T1/U
xqTk27BYerVheBPZ00H6D9zslFiLdV6Ooiit0XSR/jdd+XmjH3psfhH80CXm6ZAqS4YjNeKgKniu
c4U7O9rBgRTz+0WUuuVBM7+vvbPWxH2VmejRTZYE/dQzgko8GlvQCcpUfrDgK6g81509gbO2qng4
4fIjD4rXyuZg4JpJLXYmpuJpb+K4Ad5H38Kv2fd+557CADKzRYI62nd/Hz3Sc12+YPQB+QOe0vKB
rB2ZWRIVDUL/PZv4qt5sfDnzodu20TTfN98G6hBmHSKB7SGyJdafxva0lYht6COURStMeq+t6XO3
Pt0m+rIpVzfK3UIbVtNzlOHfgD5VSx9HDOLnab/EUF4U1HZkRaZ15py0dBPtqLztGquZxryxYf2A
oOZ5LhhTSrAmBb6uf4Pp/8uLgySFEj8XvJFWOWcSzlSCwzw1ONRSQaFZb4OmVrEzAl9ZkIcog0D1
dksqHzRzLPH0t0BTo0JktkzI0LMLDeSt31YrhtiFuhACw6nYTQKWHCGKDHPccssQqlxTFr5Pi4Pa
oEwglrFWbQGViuFv/j5HDWcbtGiuMxDX955rgS9KL7CnmUViUGpw50wEft3OmiVEd6Zh9oYVqOe+
nqVELCjpQ4w+6aqeT2/IuOLQsWF/HrJVo7ms2YQxUyQECEQ9KU7Lh1qoSuzUUHQkD1diYEk+y6E4
kPxATo4MAqBLupWK21ZgG+F2BbiQyStrsgbuNFvC4Q/JYh+nJJH4+RFAG8qPZUKKkrhE3ThikoV6
RErrfQnZoR2lVIi5GCAj/QWgi4WUf8lsi0ktvBLUL0VgkFNrJuLBaiXpcpnTzRXUZsdZFUxkhvE4
vdh9RpvkBFa9tEDV2n+FOUIJTpO3MbV2AzZevhkOgm9PJPNp7DLF2DnKLBywXAe8IF2qbh5BGet4
KPuelOZVuA571hpZ4rhYMzNIp+n+JCOu0kiLySRkxTfG7RFKPP1FYmz+kbzMVu6jLFOvg3VNtl+A
/Hn+6RQ79WNuj3vU3Ze3AuJbkCy14/rDcgbsfMiQxsFZvr7RHJTZmlYucSYy8YxtzrtzxInu1xu6
1YkIr5cHBUV1fpUdKYUx/HjIb4bmw4Yc3WBFkFWJDiX34k7sZtqYPrKsT2xNEnqPhCwWKuV0hCUv
uBNtOhMfXEN4rLEttDhUnnQyj4NiRjf6FcXM+gpmyuyQ5us0EuxlMk8mK6FVKkzGNpNZ2xCuHj7X
5FeTB7epXHZHsHtO+l0oqliEJXVsG1chivVOogLm6uhx5HaQPxBepHuZ6VGlM3H2fyEOj9WGdimQ
hJgAJd2DPd5/uK12jzzNaUtoT7uk6T3NrHw6PVK3Ite36KaocLYXD93Dk+GuHGm0YC/X/U9dvvZY
FA1xfVjtMOlhnDObyHm8KM07TKKXKhtF5uMfALNNE4IPN9MBh9GWJzbqICmJmiZG/R4/2/4TxZnZ
hG+gmYTYqYcjVVgp2T4RcGC3VGwhb7/Rj27+p3Wv7Re+8W7E7qRdt8WCZUATj8PTjiNKCYL673qW
xPRPYPKCd68NuEwce2SjnfLsK+nmvc+V/QSSsXbjCYEvWbaJC2b50hZW21nwSc1LBscxajtWje4C
xbtuLfhk7PgzmySxAjZiM5+D0paMbLpP88mAjI9Mp1yhaCHtijtCZDtDh8tnLl16C8BgL1R3wd1b
ZkOhnrK4e1LNSLp5J2hug81WUhb76B9t36QVg5uArD5vgw4JzzDSekRsmIvmfiidXELXX+4DhtIB
jhokeyrmsC65HKlNRRb5vvEFNuwlyiBWkKRCkn/7tN9oDIxtHEhRs1ORRwdj6/D8xjnhd/k6DMAb
PcE6nDI9aA8YxhUs2lkJPqP7z6JpA2rWZmCOKNZBxqCgI/Em3JAJa6kCkRNakoK47SRfcvwlLMML
XTpRa497uijgbHnyeuhpDurw5GJnTCuAVtQdBLH4xscOECMW5dKtfY8bToqlpXecWvL4fIioqxDE
Ma1Sawh4YdjyPmcR8Q9+SQ+mzpGNMbhcdW1jypsAbHm7vvGbDDSSN3vrCCjIVWX0IUcyMEWQ7V5X
Wvf+JeFi+pUGqcT8OJZ7zUIgtARSAc6hVQtrNnFTbNqnMJEyYxSvJZ2oJ5ST5XkjU1LJSzsUc+sw
Q0q7OHHhDATjk6D25PXIbQbAcv31KdBLUozEYEJm+98Pc1mw7vs3OwLLdwOfYsGAXM6KMwZ8SAis
mdtjxKrhLxP2UQ2V9OJfwvjurcD/pujbJAyoLwKu98OCAB1jNp1VkY8obLvO0h3dkdNM8leUXICR
ju5gZ6rKgfO4dJe4fsOmkChbCdABCkOC8NnsT7MlG4noIxR6fp659NqKVZMueO5GrO5hw79Du2DH
lYPe704lWrNoJn9wDK3im4rxfV4bL5lMEIyHL7ushSW2PqUyS1CZHVQU1rPzIndeYhflJNHU8SDR
JEaDfMvJew2kz4QWOdA/Fvi6b1RiAPDWCeELXN7TQDMX5TKpmEgkG/Y3AQjozGLL1ZEn/AL72Uqg
+ho2FM3A4QmVCNOVdMTsH9BhYXcz4LKctJfmTM8FD94H04jyA9BnYKsAyypwENXRr9a5nDR19vqV
brq5NVi7dY61yJKZjHEasHb1UsW7ReMRUQx0yIpLCunrzDygnlEBlAVHcASAU5Tl1Oy0f8pci4T7
y5I4dUO+lDU8/izzW/yD5YC1Ir+rgpncC4UbudwLp6WQ5sSHMNxBHq28jtl53/KlIJZWdRD3/GcA
T9nZxKKoH67oqX9sMT7/0Hg6DfiWWW4IMYeJ0SOxcZeo7TQ17dtQZaywx6BigxoaM6WjtmZpEYDj
OF5FXiYk7gva0q6z5N2sfFpTsIJtme+B7B5ADbwn2EP2G0V6GM+047xcWK1ieTvWmlXOnSahmZaP
sTGMUuLCxa9bHgNAvpHN/Efodcd3TKdHMmMNkgqXc+rlTwmla1FDqhIQoSqvJlZbE6aHJd81WRHm
rScY/gmLw+D3TGvJX+tntrS6PJ9yenH55Aar9V9eYIvUqUwy4i3vZ5XBlpdxzPoQOP5G4t+pCu6x
9CcLmS8sw5m+OxvJ3qqKjRj8M+XayUrQV7hV8fJ2XbOe7C7K8/cb/KUfCZO17F3dVa9BWtUt3mXF
O9Yfo/G44kxCJQWBjoxtl4QtQ+t4xAyzkTMoqGybR8HFhMotxqZ9GYlLCtKcDIi6p2o3jdslsQUW
ipnXZiOJgtPrgDXyLOb+6uwbaxw/xID1/CnNgnuik3QQlucbf4T5PG+5m1XyJ5T23kUy/Eufzv3n
AKr54CfkI96BZLzF200Bw89pft5f8EPuK9Zwu/v1vBRenTbtBtOmrfIVLP1WxD5yEj+TetVN0vD4
ObRaTXldRA7uoyxzSoa8DFG713jQUK2qScPXLoZNfM+KsVPy+4UFZ+ax7xyUSDjAXaEvfkf30SDJ
Qmawpxgb08zxrEGPNS8rOjb1gPZJZDEA8jwTC0CXRxW8jMD10LIm/ECenFUBqosQljoX4q2StfY4
8dCmbToMrjkV1LVEKxM+RnC7aU6Vrs2+X7lHh8igb6fQC4HoLLtNf4mqlDh5sSznK7DQEiOH7Xys
EKzJJga+RLcpdkgNbspcVVPXLS4Wq+nDpZ3v+B4W9MHiCBnjK9hbgjznMQ/jRF0pDFieErDucTi7
lUsG684VGCVoryeco5EI4DFMbLEb0rtClZB2QoZ5Dr/3HvAiAYpdMKn8K6DWgQWz40m+jkRhtBLD
DruKFQKbw90J44KI7kz/Oyi/CCEHywb9bSI8A8lku79KU6788i7sc33Ggh9D8jK8haxUnJDcvSFu
RswnP/GMUya8MvsRsUBUd38p8rTS/RD8LJlVBWZWrb5mWimnC2IsjjoA7q2YCQ+5wSvSUOoEWult
0TR8fibigN3mpDGx7FGRvRDSMH98WbtYFar6lGKjZR5Q/Q7HIFN/gIbtH4I/jpxHTaCDsR/7xLw0
NXuzhNJ93Ll4qilmtlR2sGatN8W8n6YXFJVlTHvaBy6L42SDhNTDMpjwSbNCIeR9Q09h49hpn8N9
UI+6iv1gbrqSuGYwLbKl/wDxDULAH1fIRQtOEfuMJpfY4dAEUx2CyNEoorzR4K+gKRAlK4ccwwI9
9mMkwnEArw/2D8g/3kTvzyHjfyGeWSgiJAbDHGJQCMdKbb//Wy/bp3al+n47NOaLnSGP6UhH05kw
MeIUwj0gcA/5feU1AyXTw5jq37Y5LPCWAcCUWYDnVKmdHvlAfespJEaMDrTOq8sbuI+NmUIxJ4Qa
MbFH+X9h1yA0t3kLD8ay7q7GAY9fh3PAzhil20bH4t66ENG3XckMlOru8xFxC39POQ7ATj5tBoQr
t28Lk7OLKsmerexyMd/igkOnEe+TSclPpJHsz5U1DPWu0TdzSDU/C0srR+YpkDiVRzQS0WYg8pgo
jJM0JUGm2IaKaiFiv2SXMIqlXWigFUGXYgtqcC/UsA9xgong5H9dGGGOgtIaVHSUnCLornmcEitA
kIKW5tgL7qgOWkxwyCZ5pf7PyJY84B2eAKuaKpbstm3j+0hBUj91c7ci3UiEphwBADyZzz2QzBJc
SwbwLMEmR5I2KtEt18xllF9yzuzYJfqvLbddIdr9V+LrkOAXqrzecI4kKmTmaPi4HdNbaJCoA5cE
7oS+Qf2cKrCAU8ISAViPJYlaL3A4KyYK4BkeuPL6851liPh89pBCYMU3se/gN0Ab2d+G3AfcVnSR
sI3XAvc1H70qF3lPIxLL4hhkWnLaptaY4WJ3X+j8kHtBf5tqecYVllxOk1TqvvyYNFfPktQBVFfo
/pkddd1uYyFPpLnrxCRwGrI9CjmFr23doo3RJJWymG7/36A02eY1zj4yUoFaljaSSXC6KvyPDq+7
HYrrg9NdXJdpZWwADAhVxDBAJ1W41UdAnfMs5BL/mfCp0/3cJ0Gg7MPZUjOO9J4Lldtty9LbLd1C
kZQ/fvbLg7vdNFJj4bOm+xv4aqsRQR6CRSqL8w9g5OoYWf1AYRqPPvNLn3nreoGuMFp4xMPM0kgF
OIQL/Is1RnUL5svyHXiF4nOo+FXZsA7OqrMuJT/bxwTV3amHRvybdPrSkw7k/q/h2e86VpA4y9eS
KeOO9HqVyz8R5vrryeNSFpTFG+HudG8WbiI0H4HEfj+uvfT0wlFRKqhHy70029kbQzxxKhX35toh
azN28y3FdV+HV3mt8khO/bzSCoDfvoEgeeNtXxyPkKg3lus0g97CB4Jl6rDUU/Kg0x84EGBGA5tG
d0ftL5OG2U7ZZkop4XtKn4H6Td5oE7CMflmXRCtsfRZhlvg8UsphRyiNoJSVI5pwFcmvV/lmWCzn
jh3Dh6OLS+UPeAUkTwKH8UFePW56CgoDs3WxffK/PlNZ9VZD1l6uD9tOwVIEvf35qLmtxzWvYtlM
bKnUsXE52aQt0BV2smtVjVC9i0/PmKpuWDdo8R1nX8L43tWvdF82nR54eL9WdeZEB9iCO8jkonlj
SgiFdSZ51D7YBcXMAw2+rn5PtKYKBH3x5u9FanvGnTKfCuZWey50GUdKbnEpch2GalqyJCjEMzIF
6whI/Q8D4+bOZp0iLNEmf52LrQNwwRRzxDPcCdmx0ThtoVCdzvbDvNQUuviB4bhTcyHTAyu01rFC
U5Y8U4PtomGurCtT7CGOM8UmHtKk2UAHG7b2QPhjy2aMHYtsLc2otrLe94rHoJD7GRk/g23lv3wv
6rdbsSrqoflTixYKk+EpGFE3gKTsrXpMyyQZWXNobU951gQkbk/Cnx9fN9xbzB37OUfySd36rOcN
/3nVbtxoj4b3Q5lU1vO833iQSoH4lUd4CIR7Mnhn6ET1Vlk0944yWpjygOw5ipwTABM4Lf+dJ4kq
9gYa6R6p4yN9K0EApmytocrFBVEnbRu+bUiOffpzr6lAXAxCcBsmszG9Xdx1rtoII1+aLyWkvScf
2rYWoiP/D3bfYWwZZCfruJdDQFeb+54eArrrUU+H6nvuhFSALyN2dMN4RSwDUstw6pnI30dnuWAq
IL+kh8Wj83GhZkZEJc1gBTdJ/hg5SQZrYUoTXBYCT/CF88NCR8iFA6cw6VGSfUudHhsVvdM5GXML
eIxAYF2WvKBydGwyOa00LPvd8roWOvaSxJd9osdqGh2rhq24bB/CkmdImRPNAaBAlcVY4WszkRPo
3UtlB5zlx8sts+3FgLkd1bmrShrxmHShmz7A1IOo4KJh/b+kfGi5zXOQ4S4X/dNk2rW1ozgyWFOn
fmugPZMtinkOMcrn4KFMgk08yy6sRn1HemfTVh/gsVLRFPZYDwbrDRx1SfEvfXCRCD6MJ/73/iRH
u6/B/USnA+0KTcSdq86hgW8Bx3gws6iySV6wC194tzP3uQOCQZvDt9ze/y+lZ35toKM4ql3GhsBL
6uO6Hlc++9YDNOdHACN1Ga4m8UxtlD9wb8mLLhE9R1p/+N9yY+4K9Ppv3JwVzEmY0s36WhPcwGhD
XSWmoeR3spa7uWNuoxJK+lCcf9cHXBvTwBVv6XxM2d92CjUrHzfd5kdpw5BZ6p1kYxUZM3kafVn9
AAhZTIhGrLxRNUetQxoIyH8wwYduLMUZf906gQ0x127tzT8NVcE9A7qgsdz+SzzkEph4YAy2ZDkj
fPyUJUdR/A09L26Bc8jprVUzTnxFlF8f6aPcMu4Kit7S51LZJNkPI7Edg9eL0DJ/QUD05nUvZK+e
hfXDV3Ahsex6UETh1kcSWeHxyweTJHIGajZoSXg7QuuEQ0NRCPOXNMBXB6dkAzj9Kcq0rvtkt2IC
XvoqmuVI3xlUduDhFIaBiISdgV5AWE7ikVkrHsDoByTjpMfe2RpDhvHnJpwvVcF2LFurNwJYegeM
0PNZ0nswS0btlLVJwtgsfwXIPF8BJdE3Nn3+nXY7zG9sJLKS9dYEgxyCMbczwGc02nJ0mrOqGQJr
NsLDmgc3roxiuBz/P+nOQZe+5KrWtaHKhY5wPkY/5lY3JAe3wKmrdFrqLgHaGvI61i4TZBXw0NmL
akiL19/G+T9wUPyUGEzzzkdcra60+MnHI/sf4J9V+I61/68J3bMyt4FDZpp9vweBqzth+TEh/eMj
KF/DSYrHaCrCAfwKDUYjluHasm2fB+6vgXJioEuQbMA21/lie6gfDrQYejdqpdR9Ia55e+PLWyCC
0D1kw7FgzI8DODg2g4s1ycp3SKiAHRPPtPAfa257Y0dSo1t85nTnawzIPiQfA3v6+YyX69ahERSY
k8u5w8gaYIug2zLAhkIFisCH4EWHaKKRzw2rCo8jsu0p285q6xrpLJnmdpNXnowZ9MsMxbRaDaAK
UDlY8s2t+Pj3w6zqys2eCEYB1wVt733CXJXtg0VMf+5muHwMzYrMMlIDZB/4pCw+9k8ZQk0Zx5cd
mp54HPPURhLGvabsl4CGgxPDQQbI+MjkmsAlfG0Be7s8wUq9bKgMZw4yNfUEF0g5wUVBasTXHTTR
u0xXhyrKXRXUQ283WN/nGOwcbFhpzEMwt01XeRcH+DykyzPCo9MNmiyrEU66MpLQvicE27RqU+lu
afSZ3PIEDZAOEs8tWF3vGiEqH/ae6TlgBQTMVofW+yB6arf9yDNyDzC92brQw15zv5CNIuyjs8xQ
QNfYUs463OBKD7LtcS8xvsznQaRDOOJq+6fsX3AwWzBZvBbDzXW84WHtRtwwWRicCXscbldI6kTb
C5wcjdpovGxSb7tcKJk/87pzDDaXUL7v6JmZxUqPTX0vNt+WObHsmqO5lUyLOsY5CASmvI7YT7SN
K9nYwwTeHpxdpnpTeRT2qSxy93M7Kz303uyyxQfl8bXr/yST8jLKvzqkvbpbh4WVqh+0BALc9wMl
SxbZ+HOnUY2OZi6hqogU0kss1H5VANe8uHmOs8h2qYVw8sBZbEn/8roV5MnPwhOhWQw6KV47xqtE
sQ1Ibtq5onBJTu+SgX2LDGF/IqhERN94pBPW0pdBSo2C82hkoTgaylVVr8SkrGVKWetPi6ML2f9H
qhUFLfVUCyE8MIyFOPnFEbv0EB2LLKgWoOg20P/QSukksPjQV0mCk5Ex/ppqj/Om3/KK5qilaMbU
OKkUsvZsTLpOGwrvwkjxKJ6yXEHds6F8AKLGGDRQNK3OhXznv28ICue1ptI30VcKx+C0lJ6Ajy9R
QCyc+i3cRt6JGSOe6qX90Zqyi9PCEFciyUMYIvg1Uloj0FIhfxTc/qzhYn5edDCVnchKbOwq77Qa
V388NBkmoB8iPbDw7XI0o09FPD3mw5paUZYKGnJrT2KcE8f+xcQKorDMgKcy2oaR04ylq7+eGCjR
PSBhLbLC5YjaN+QFz3QqZBuF3oQ09k7VuPbeuCKB/7pomURwu+HouOxpduhc3X6q+MB5S8PnAptH
LfGqcjI7l9L8gDtH+dJssvuIsrod5YKt3m1ZjHOsprPkCdQ2aQVAb9b69cLHILzrlZ93skrrqLsz
CRiWScLu2pLvlA2aY/S0pamQjr/HzsYY4d55dOecRJj/KNaFsXowkOL40DotV5NpMtghTO90ihDM
MapgcV9PNMoR6O01Nr/0v0TCFEOtRk9E3PN2K1bHYxkfnCuWcZTw8hoRpgIhhyYvYuZ9tuqVZqyz
zV5g+2a5C6CndD2WsStHTDeuCKJakCVVmBumTZ6L0kIiS2O2cAz5IqQcXG426KEnhF+WAeTV+N0g
tMdLsq12/q5Oms5Sge1gx1AnBI6G9D/btg23d9FbxT9YWM64IX2vqJgxtOYVwybMKWwbhAhhLS+K
n7YCWcQovKAof2H0EeeIrfE6V6l0AI+ufjJVSOif47Cw5hSiLEDb4Brb2Znfz5QQaStbbgWaoZ7h
kqXzfgFM1LGotrOfq0ye5LW1tdZ/JOX79i2TuXLETrBwKTrMGQQHUFoX9xagTrBlebYtliAziuCk
wErqmkFhJpEjHakhNtuKW9Zc1GEFZ2iOLxTw60Nebt2fgW33aAyourCoeYUAGU0QecOeNobAKP4V
HcgGyVfixiPvpj3tIG7+l+K5aGR5DKWhXXz64UEZxzmF2ftoNPZ1OAf9G6cG/12C5k6b+J4ty3g3
vJ5NNYGh7PtU7dGZ0RQzrMQdec3HZRXP4E/8i7J4kWHjMfzJAB9/hNjXlGEoiuCKG9XVZuqpBuou
ipOLZTc/MxlO/Jayf+NZnBe9sc2DJRCgc8n/EaaFzujiaPvjUqGS/0YG9t8WwKzIFddjmOzn1PEy
XR1oPvDWqvq/A7sXqvtCtdXUBOy3YvNnYbX9bO5nQ0ONE5z+h+q5WzQjVxwL/PeXfHKc622o07JT
dr1D5Vhglxf1pM+H3xrJgw85GpnYQuXlkMZuRaXdw87qJcfT0YLnoftOGDqrymf25Rz8XBsWWu5x
WucSlstGIsJPkyQyvkZuC/+jdnrl37AKSNQB3MxzCRWCfexfgvNHj58sU4XlqxSWkuIc1uIUc8k8
su21atwK4ZpUGRQX6yc1M7ka43W4T/ax7pfbdzIKb15SvVRNQ8ktdapCbKZooACJUIQ9DYW8BSB1
yGY/wWFxvOpxELFk1ul7rrum/yi+NeK+RDGFC5CYtj8IIdBIEtE1kdlOeWuFCP5ho4xRRnLVQTMR
Pnbo58fhHs6YzD50fjTJW6rDmoL9tXhXxdeksGXcywdjWMdZ9UvmK6f29yc3ZE/8kReeEZIcvrha
5vsQg9AgCMN7nfKOzZz7kZ7taRoR01T4cGKU06K3G6Hx7h+MSk0zDE2yLM5cauq4ZT1AgMfA/ABX
MNbjRoPeNChwjKCMcBU/0HRllFxjXTCTQgFOQWS2Y21YCUxHfvPvUpqG4zRfB4WzycLcdpBZHZyy
A9y9AiaIuCMb/kEjlVTFki9jx5bRWQvnq0gEmtqLe8vi+59Yq8DLSLzFFGz4HteY8NkzzXUTqDKx
LRWrJZUhWxVQecB+fagySfCCr53tlmIEVbhHMpDdfuzkrOwLOW8+n8N7nPU0S4orHBJrW9HDVmoj
w+nGyFfecZxWfTeHh4STrv6ze3cDXuWK4HIhjnKMwXDHk11QTwi2NP5hRL6U3IQ/iWDyo6Ee5kdx
u9xe9FxGulnMxvNJbeCJw+qPCZjdLue7Spgvt3yuQoTcw9SRtzQT1wLfZr/WD37o2l3uAaCC7Eic
j+IXMlj0NY1MSwfVfqo87SRyQ7Xf/M6yXJVEli2vEFKh1kMxqVLxM5tueDwTEMx3cU/iAzkGEBEp
LEQznPr6VoyozITvds2QLnMPU28Pi5+RsTyvWMmlkUOtSkjLCOezOWiEHpHz7dw3ROSPh8GHDo2H
4MB7WMU8QY4rWTxL4LWdvoEPktv23L35CrtLV1LQUwd6bB34uplZqRqJPec1gSZ1cpBkucO9Lttw
EYHKtmQxp/84ZW+BK0OxmcyjwEl/wHzeDZDIGslLkVdqMT/vDqR5NfpWdPFJLVoBErGqFlBqXjJ1
OXhdVxjsAjAmPjQ/sbXU/M8INcdGwydbkg1SGVnQJqjpz2T5yrh/PBOEuXA8Zm1EBk9vS/f/HuY+
Y2dJ5zh9Ud716Ng7Nw5sh8jRjJKyc1tf4oKbNMI8y/KA1181adrDV7Dz9MMHMQB/rVILXhSp28dz
bzeJRXTQqgE3J7SIBTxN9jSRBIt28xAEXyXcxcpdC6eWMINE/jWHxrmwy5cHYi+hWYeSLiKVtECP
9w9TzWXC/fSrBTBWkW9334nJpfUiiCyXyrXJj7023u0f+is+bbqsoegDAjqzu4GRJ6T4ory0lTm7
obSQXgQkelttAiKjjoiNn3n5pja56H3oWxGVI8+3tRFnmtQTv6Ok1OUM+CIUOnY1AtXQe6lMta87
2w5Y0SLSmYbdto+I/8XYzf/sp5beOjUt+QxPEA+DGBM65rZE61MxQ6XSvDd+4eH+8ebuROMt/1sd
7y06tAW0Z5LmyAZE2Xm3i3tWqPjLb5CoxmlFmF9JWl/dJzGM5QfV2R+iTcG/L+Oa0hQC35AKHQT7
7APLJTa7bbCcpiNGEqLO5kPOGevnnDZz0QBXMVgbIzT/EU2UVVoogPFzPI/EIue3SrNwOwL5sepJ
6J5FKuJ0xUPdXncrQv7LL4dCNOgymSMeGCNjjDi281Pd/6/8YLCUZJp4KUcGnhB2QtP6SWBNl6pv
jIPyNOtGqk8bq7L9/p2JP793bWKLH/m1rnph3p9/zYlNE4S/wvQBvnf9YRLqafb5uDek3tqj9wJO
Q68xQPpe5LfRfLx+I9qqBao8SNOwGwaYq/zr0LCfz/1Fsx2NG5NnD4FLieFzqC5xVSD53RdhykdT
sMrKClM+CKljUtNrpphxyWk8k+KFpjmdxABw4gReLO7tfJJi9sQPcjQjCQsy1mQ2OrVy4JeBtZrg
cS0hWyITfGVtr+uz259grqPvrf5VwuzJlqFuIbGsw2ox+z4+B+S7OIJRj4umTid2iP9lJDHG3RiF
+Pza/QYPm45kFvpnYAiU7L2wJssCrH7Rpv/PCWPtLNCmqPksTpe7qZMJEyNWGTzpCeEiPIND18M9
n/X5IJpHwBl2cWjaVJkHxm3Zty4DzXyuS9A3Dl5/nGq8/WMJavUaVRJTKD+/tyYTwvJjaTNsa7l7
TIlyvUaCMohrMyscHSDHhWQjRdUlY/FyD1mHywyBfAf863gITlHZ23oAZdUAyVk6vZe0u1a1xrU+
+uU+8EASpD0XPl7y112ZYfEon7fq3y0UQVCTRod1uBS06ON0WvuX4jjCMv8MLrcs0o72xHvNhUCk
K729FgJH61jGINIt5BeH5lPVd52A+jNroK3sNXGlB4QOSJ7vniWuCTfAFthqt+FjqlC5LVkXZk7t
9b+4ujlaOtKIMec78bPImQrK4o9fojrVJTsM1KoKH2E8aGKePBWxYb0GkDmgeMUseUe9nhKplDgq
AOQ7bQrLJSOK5AkDtpMfQIttIu0frQ178SDoxtbB6IBYnuDeJFUwHXA2L+gxp7Xb+gzW/oD4+iwJ
1uSygh6gIZnZOxfvP9znHSuIPikYCpcSC5BLuGgaj1KTd53CL2/JSjHhG5oBqkPApixS6Ins77tv
HMHNhQZvQIsqK9G6Cu3Xs5TkOW7zrX27u83FziD28vjqERcyT8XYayL557qGDxGMxKPABH2jV6m4
1KNs04kXy0lKG9O/bZkjgtJNf4bSdXix1W3vY0JYfjB7/YocwdyQT3M/BbOqYAfuSR0OGXdHL69j
pMZUFQZYiKtvzPglVPAtMTB9quAIp8VzVv5hvuNyhFgMRntwCWi98khf8Nur42c4rJxSU66SlTx1
ETPj4IZj9a5vRxFBQAlibVrC4/AeMTdOugksFjn3pNqUKZfeYCemQoQ0dIeMk+rP6WBrAxpOvE3e
194nSIftNBmdkB8ZbDqODQ47hxthsxNccKJya3VSiWA/U8nH9GO0rmxkt4FjTVgdsimmxUnZWP8W
rwTKkc2XJKLunSOl9TCFP7LBcHPwdJVPJYDLlknX9iMO2ubOTOfPf+R0F5KJC5IjRwOZNVCmsrmC
gp7cMKMrh+NFsT2IIbd3JJG/oMX19ak71XjB3pc73JFJuJGozZxvdg9a0luHHfv+v42SbsTFEF0r
B8R7/nvdAnjKrNciSid3F2oisBOztCRBPM/GbDD+hR/Rk9ndJHVY9umVADF3QKAVpLC9QQHyhMmQ
NEJtyT0kg717GD/5iUiCQEPLPUX1Yig0jUbV0qZrGW2JOSCFPlSVxOfVwafeMkyBb55WxkjjnMZ/
NKg2hmuBIT1K3hNPkJc6+HrMxi7OpVzyCqvj9IfLNokhfqMJllDUhNFA7kLTFRHYfqASG6Nz/9or
bOizqT71KWjG9MGbo5h7Q0W3ofOA7XBwUd087CmaEVHDqSrLAZFk4L2Um15moLJWz2uaQs6+L7eR
eKUSnJnFeLBwfU/+gn9y4d2htRZyrZ94Js/INBFYFvJfCxQD0O6KOtSWFzJoeH4ELziF6qecRvMB
9yWiEEqkVfPh7Ufd91jWSpxFp1grdH8RwYzB+vhTQxKeM5Y5R94LH102Epv+UjOJa4XqWKzUiW9b
9YfHTZ78og++KUQDGsjRoii0M7AAVC9lhXxgQOPeu9SzykiQJ1dJ/JqouluDkgjdEy5C5nD/tSG4
Y1vzIIp7nB6ILoMr4oKySfdRo1l6aXbUu4aWUTF/7HGaX0LM7U6uDHHwedeHYi31rZvA7lIdq3Zv
i9kH2vhJyuQo7NPRA7gt2uBFnN/73ELjIdxqddgBX6xR56rk/mlPysc5lITL7OqISeabfBoFZ9Zj
1gtl1giX8EIyOtUMldDL9zm6+/c7F0spo51LT5Y/0ng1gr5sOqLImdEGJP7vXCZlMYEElAj4/oZn
Dy7CVv+Gn7tC6AvHC80mZfSX4ntQZ1HVyMutcz/NMJ4q+V2/LB7lpZV/UnW/5FeKeQDhK2w7TVHi
8ntcziYybQQKAbnpsELhHGikuNbV1+bkJJNacDcojb1ro+YomtLmdI7B6iUD5/9N+wfqx/kCqutF
3lyTktnSaNspEvj+BLAdY4j12tgff9mDoZNqlbJBqyyshlyLvZspFbD1ZDmuw7ey3yVHFSGD8Ar4
iR3SNB75zejyei4WQVMBWxSnYW0uF/ogFCAyEVM0Vho0bjfaytGBB5+2ilyjqL4bGSg0rVt4obe5
xjpHkJaFmGV5mqyc1koj3VDs68TW9mkQF+y3KKReeU+m+RA9ZryKzpkPKXXAfPX5NfREo4BTw6Wo
3xL+Y4pC5C9FZ6PQaQkGw1kLfMhaYA3YycpSkPdaJavnLCN9HuwXQHsL3X+59huINWSOsBuZD6BR
GV0QCJDGoiMwCsQZIVTJ6niA9ioQRLnzwgIeYH0jgxaJGyEO8pTOkIhAUCCuIX1tH6M/onhgKD0r
hPi9BzogtptFj2/X9bKoitaTBn/22kx88GXHUXd/VwPtWlASDQ8JVk4SBr7OR2Q7tckocpKVzIOv
kpSeAGqvwt7LyKCxZoeIEyI2uD1SuXmy5j+Bova0kJilOzACl5/UbcfFXANMh+kRPUQtKGgRvFVB
0mr21pB8fdP/1EJbCvdnc4lJw8WjmrexfS0QXG42eVBCR8e40gqxfgKBxtSbBCYH5Qvq9Af+8CUx
SIvTXxD8pWvWjdijMVTbaOOM0/HlerIRtjyuBckfV3PHGGb+C8LC9y/fhXd2hur5DUFg9VtjFw3+
J/G2mS0q9mqbfCHGSwvoGEuofQAIiv7IB/SDulF8R1cNfSKaPpg7ve3TyI2ntP5YwLu/pCmkvjS1
qgeMgli3nk9O0lQythu9AOxLqk+rtI/CJZ/VQ7d9UTUvs6YCMLsE5iB6u/uElLYK+9RCT2205oa5
IoqcafWi98bDPy2Z+kyH03m9/uOREsZM/8o0HPLEFZhRi3We6vbMBOz3GHTUD906xH9zO6D2HWU+
nwjYf1XSUjqVgNZclFU1vmlC71kb7Gmh8ZykAFUzgrtBC8iGNOvGo4GHa7Oyo3TtIv6AN5DytrY0
z4q+b0D3rs+RUTGLe88861WbFb7HLb5Nnnglhwngp88Xd6hfC36TWhSpRN14S7lUR8RbdcmeMbKV
SY22qMu6bZeDmt23G1O7Hrr+XKDxDMug9QaFxGXbz/AXRLlWxGnXLcer23hpp14jOP5gOX5lTUFX
9aHbuOKyeQJFqoLo6hhsMSe0MGVUIXUiB8GNUEfswDelK32WYFZWClua1V/EeBpvI0wSfffJ4948
TL0cE35LQJF3nYvf/3AH4cMNM+WuBRMOluCv/ZxyjqQPRxxgUO1Q9a/KgXwBBLG8hAHj0UKNX6oT
T6bs5jtc5Zp9CZO3X+pD0sOxJPybYlsFmOgRaptJAIuAw5qcSgksnodzZ9Atf0oPyUhrA4KcTy/K
bZnDfB8LWcchivodt8zq+n+S0KJT6GJvrHArKbmxvNYYNUo4Ci/smp6mNYWVghvbqo9OBSidjmRH
sBuZIU/MkBefXOrrGnGS8G7hD/s+8J4OoV3Wb7BSIHnXgi2KfRFLyZvE6Edgjj7wD1G53dkawpZ8
gfykQIOUQabMqp5v2HrsKBYVWarAjLqoBq0oaGJ2WdQHuiqyzjtmOe6ijl6NH6fasHoW8zonDsz5
kbGFRDJyg3yWC3/rmUdF4UrMrKifnmda64u8zM2vSDcWN3HMSTl7PyBA0n+L9NmPjokDIon71+SP
ZgGP2wFMcKpt+r43E2BWuABquzbwSEBqXQRaPVn+N76prAGwq3GlRVqIeqwGYlxbc73o2t2R85h7
KbFVeBpidAdLAZ9QlQSfTfDhN9lNuHdK/bSiLK3zMwbjVkwukFEiqZpSOjIROEI5d6lv+WdR+AiB
klPDZkHcqJyAHzuAFBPk8Pt8YB5GPAT/drXp+7VEWcnfMLe1SkxlX69eptrszZ0ZUWHsrxRvJhLC
xZJfaWvrdZXlpaZb16XxjiM4LVyf7y4DVxFZGX0iNb+oUqiahEYARJ/M+spRRPuhFLXN4yHRUU58
4GxhCDfBXln7lLIntec471SNAt/tCXeqeTXLpBfd3N4tIuvBhic9XBNXiUUyyhdUN5lJoczI2glz
QoP1lXVk0CkSFUreK8S44LKghtCHSdnwnhFj5XRVqyeghDSXcAbHcT/9gtBNN/2BBFghyEgpKjr5
2bnB1Kazhg7h+iF15oOXPp4WyBhZrxyh16vAx5sHFXdHZ0mVOasie0H+qNRPIqdIH8VxljNl3YTm
HH15sz/U1QHDtAY3FwE8q2vXz7g7fYpYg8IOqGvSXyPwgWId0MubguFMfusUumTGlX4dGMCV53DH
39N7aub3YJfJsrAhf1mt7rPKGW4NiAwDwB6vJhGGztUvv/J3DRE6tjgMgVZMaCcrgUhr1N9po2Iz
Nxh1RjxPDW7FfQ9iEgLLG11w3Km6Qy/XWhHDEnY14ittLTivDEQzGWYLDeVYiriLl1he1mgv9y1s
vurGN+d7nOe7ZsHBPkl5qVzuQdg01Pyb3twE0xZfRNUDkgB+grp6thY8b7inrgm56LpFLWg7FYb6
jehKWf3tncwkuMiESDZurZXPHng4gY7Ixc44c2hA2lm+i32deUygNji0gVHZQvWd/yUuzl0+8qeR
DbZKy4k2C3e3Sfclh1gGK2Yjflb5wBTvine/30Ah0W0dbiSBb1yhOiayF8gAIw5Dk0Jqf/tit5Ba
9gYitcgMeLKAcslN7uGO4WITlCBDUiR6Uo914E88WeZYtdAUu3M0/jn8S1y0N1FJQR+Hixyu1XLO
z2HNCP3noEF6yMVCahnBwbh9HNt+To29KKuP+N15m03pSTff2kylPCBN9G0mobIhLSbaeGc5fWrS
vMgb6homajoOHxfkJpZWB+ETfJtwR0duP22EzmW/t8PD2CyQZTzLxajG0vidsZ/Uo23bEa7H8QEy
0vePw/q5J3YMOEqN/fR0bbxF2mvnUzP6wDpIatGo6Wvdo0qFS23U2WJVRukvBp+WGE4ys0WOBmCx
iMYEEq1thUUOhilS97kCp2A4BDjzGBPvoakdfur7m9/FLoZRxPOah/jKSmPJjsJsSCilT63pV0R/
UHgf/gIEPeIURaaJjD5Btpa1Yubs+SMwPGHbj4X7QM1uFM6u3SIkDRKWUQJCUndCxbfKWUBHX3hR
chUau0TEU0GxRilO/9j4s702J+7RfSNcf+0NFJ6pbT+uy6fD6AS4OGpOLGJZWjLo+bJcOWVaZbAr
wb9AFlH/6twl3cBK3H2Zfj/oMwSet5n/mQGwlBbl/aYSXGSiemVnqo9szYuZ6+gsQr7bmT4PAkqm
7/Keg+/kdtgYYH4UQ0GaMsQyGhciqlD9NEspY8IciF0w/byOTZj94qPjMw3gmXvwAnu5vNU0nUiz
khJ3JPuoaWJKOvj9MMepw40+SCgKx3cjSTH1+sDvGeEZDSbEikQZuXQHCrCapqL7Xe7KaLsoRrfc
QFY8biJQE23OytMmd3+Ac+j3floGK9QpE2OxRtWANIk/WLMmojUgm/JuH/KF0Vh5uBtvhgvSa3Oz
9NGNjRrNoHKVQoXmKZQLfVBVgKt9KiyrOHNJ+jaRzgb2CsMFQecvF6q9T20NsUFOtRBDGZ6QAfL6
Xt+x8gOmhmsjwjq0o6ysznkiif5cWWsMt4+5e1+W0l3v+EEmDJQmr8JTtOia5OE9VVkWwaEoBxhv
vu/eXtPTDY2bnzVyj1smVx1jZ2Su2peUsCjt32nBkdclFWfCkV9wywIoNGBom0a6ayWeOlaOzGad
Fs1Imo1s83KRk1T/c7osRhcvcDpYqz0mQS7X03EuNEInp1afsbKEeUEJiD7xGhwtwsgC4IxmGjCU
bpNyrCVedI+0Tpbj2AeWRsxIXQ6pLGRoxj7Tvp++UfiACFIxsJCj8CDEMe1yGbycGlLpZtovolqE
OO/Q45c5HRs2G3GggUYPE6cXEoXOqj1PthXqSHumlGF0KgjM+eL4ICPckHa5K8fx4HghchZIUmc6
9fna5nn4rGXmy0zx3T+oWiVAhG4NfymiYDD35FwYzmJHnKcVBRPyHB8kZkhfeDWO/nXLdb5pJdze
uBLxK1RAaaU4QUP4ciGRX7LhKKryLG1zIfTFStErKAdan9ksa4LyQDdxV6jI6isM7wW3+7F7WnX2
luvIeNfhAq0XludMy1ei/LwARZtEWiD54x8X7hukgZCwjNQ1b8mZ73Vk/gyC0X3oHnV+W44DOpWG
pphUduqAHHmV8GiehHHFkRQsxJMG6yGv296MBD5oK8LaFkoTRHCnwTioEkjWEw9PISdTHU64WqMx
YL8ar1ku8ByRB/8/3Gnf5ObfF9hus5aAUmgQVJsEyYYsgJeAjyyo4Zei1LhdsJ0PkBIWPY5kRMAL
VLewCPOQV7lLXowa2QA+FS6eOTGRrdR6piOWMNWv6R4geFRjs17b3F4yuazOHO3eSDNg/XA1Djka
CjQT9kd06RLTAYK8zO7Iu5HMUDNn/qENaAHaIdhfUEOHGfzxhrJfFUr+GUZrfOHHikuSWdM5hn9E
CUqCYt4x2QgV84T1plnnd5GSz9wiz7Eo6qXkRQjxL4N6qBRlMJ5nYU4mY+M9LhWVjCj+sjUc/4K/
eL3E+L9vz5u6GcZPDP3zbnvsrqnOYS1iOvrVeLypMVLTX1tbMu+GbnNN/DONS71DZdynrxuRzo+b
Iuz03g6/gVDyWzrKD4QXiLw6Y+bGVfNNuzS8/4H19xdsF7gphjjFvTf0BgARFjrQi04uaIZJVmm1
IU0m9u1LeTLcxG2Lgry+CVei38ooKlXH3ef78cNbHRimy0Z85Rji9BcONgCNUHSvJ4orTrPDTfS5
v3zvS+XekRW32CBMKpOYEQIXeMc5Qh4dHhshCsW4VH3TANxX0d8/cyrvbn0/b+frMRNcm13dzTnD
OvefG70YNbST58DYeDdvd3RTyZtZCAw5vy9H19o662cBTKRQHLceDubepqWIgYobpYx2zYxyQjmC
fw2AnOXUfL/5WLBgV2dT5LtrhPHItPqxDKvLiOX+qTCfXeG8f4d3ra//rgLJQG2ViXvNrSpfZ9sk
pR1fUEAYC9eygg4khlv1o4ALXTl6n/82NBPTCi7pbVRT6VpUfq6QqCMjC+lAmvOTQpzCAXVy3SJh
DrmvQrk7t+dfhMPJz0uFq15PY8xsGByJOOS7Nhsp2enY35Uw+xKtx11v/OPz09Dmh4/h642VSfbw
jdPbylZqNz70D9q084BL0sjKj0ZBj5DNjUL3m9jG144/AYGWf1M9UkKREgGcQqbpc+bBQ3ME9Tnb
O31Oy/WJ3L09pDLFEKksaLeVN8MGpYM8H5EooTlFBQCa0TgCDwhCEyqLhCPFhH3WJ5LSQkxqKt9c
9r0V3/dOPpwzav0R6ZKFeRutjcsbQEfl1Gm4df6kooSXnEWJKWXRYnFzmJnCoJVgZi+1abTMDhpE
hbDJN7gyOuLe12jTfn5zSMVsUX7lYFePAV5/YFEVV9bX4LuCvGRwUNKoTFVtTvZm4UXrcO8Zt0Pj
726yDMlCWreOtpwwLY3+JqmSgMUHN+W0RzFKUg0PwSOQ88U814LdzTmSsQWASXHLrpdf10l2UA+4
XcoMnTPeKAraWTTkET90LdTPVu5CAhTv0e4waGoyxn6O2Xr+l5u08qQQfRhiLu4zR3F0jcKjoxtP
J6IpzFmeFf7SGfxN407GKyEA43dyFobEYQOM6L/NdICx6COKuLyiWY9Y/OipNQnBiNXbWhC6xeTV
ay+toRZT3PF1X4JtdJPpSsTGVfy8SFey5OH86FOWfCE55Pw+oEo1i8DlyJ6UtgywZtVyxY8/eHMq
V35shmm7PW7VKSmEPWzrvCQIjfBtn4PgV5FwPZIu26t1Zym/oCRHwrx8wdcwtSOrgFQXW+1uXnL+
qdsDkiWdMI/PsaU1CSkZFfBNtMa/8WL6RQIPPiNZUCm3mYt0FrQirTr7DsN2OdlP2flVShwTvT55
dHTLL0MCdx1AInhffbVbLeddGGvClcfzlYy/DyHkep04dHHPGEWpDzMvVlcsH35CDExTRdMw16CX
psCdEC1Z2bNS7twCygf3252YvQ3i2lb+zZ3JsQsmqoOWu4+qtV81m4ZySH4qV8mOMt28W5d42Jc6
Nac1Aoyu7o8wdhnsHcNGBtm/cf8iwAxbvPv9Wl4yhMHPub476h5rjb5O6tP96uopGJz4fqhSNmJl
RV9HCB/p5LsE8oz10jau2Va384vTUeBjyE2qTSAAXzECNjxKsxAMstWuxrwqGsJu7qd5U1YLC+fi
qttUnSL7hHFV+mMma4VcC+p7KVW6OWkF3JkZnt838xtIjVHAqvBcsOwISLriCpJBC7Fb1XvatI+l
LwRzXQYhYgybleiqYxxM+VTHNwH9mbt9t5C7Lw5wHADcCFcre3xKVPR3dW/9O1uFjMlRrvOla20V
0v9FK0jIu/jQEmCIyDekSQB7MauFmEulV0YiT8Fp9e6o74nE9CbdZUONK3IMmVtM9jwX4IQl0e8p
l+6Snmooy3neeKIc97SxIyTTWwpa/cOfnIcNp82TKfk0jeNmsd0J4HX55MJtqznHTS/wBU7RPT+W
8FkUjKo5WYFbD8aI28x2YEVdsuyqOmVMGpjimPgvIVzfdf2Ds9/LG+mpCa/oJ/dV8mxMHhVV4NT+
DeNg4rDZlMwa5jmMCcRD08kqVMV6KkIgM1oMwSfaeYrr4KdAc1BmTSA1sy0gbcqnl0s6uNrlKPJ2
ZnrMXv/snC25c5iDLqykTBw7fk0tSTurlqALHHPMwkYLXK1csuR0eNd5VbNqKc8N1lT/6s5jnC5w
4DrLw/WWnEr8NRSVXzZ+BjzrHoyGuIOisLy8oa5uNk1VzyXWsyUvMbbTUweqgna7//l9VxfgvO2Z
Cwvj3M1cnVzwXKlh0AfQmqL0X4ydg8HIdrhHv1LUBkP1HYegc4AHE89IqBLRFl4IFZWKUffpf1yC
cN6zitQAgFoJJlIXpL8Asfv63hAG1gAcH9BcQpQ5u5AacyhvcB/f7g2+TrWoA1zpxXf6m24Mq+Qc
uq2FxWtgB4C+d5fBlhNJzMQZp9QrhNcI2jjqv0aGS1y7iJ2FWskO0PjCv4+ZZIxJbi44zUyMUIGY
KluP1ksOskP2jluEI+x6jIX7rYjmVrOGI8Kl3ZAeVR+CRrXNOgz4unuBm1dSYPn/Mor3nUBdUDQA
89ETUKSuXSFVY+wAdhRB2tIYn9W2LWMjzfBPeUZ/B4tdUYQBgzJJckCej7Lh6evf62uufewiUpS3
Q9TQqeok923sRdhOA4twiDoYFfktJK+IXcnHztgKdso6xQVTMn4YPaz3jkp5cAymkHM1nm5QuO4o
XMJiZ0FfSM0aZhv1zlNGYc7pCZVN0VMYP6jnqbIN6rQy6kdF9zq3jk6vfLovA7QKDvfWxx8U9ej5
09OKMeEjemVwLO0b+4b32P8VBpBeMwY94mjE0YLTlY80ulJCuex6D7ytzoXSLlrNXfOS8DKvcp2d
NRYlZD1W5pD7lTMGokcHNWQ3gnBpRdarQhiWPFP6TeJo3uf2Bm/i4oLP3Nm+hR5N5Cz16gQaaRzB
WxEb8jeNEkeJM7tP07SApTcYCELHviSh9j/7EwMyOtGDYbhuY2uGplnyZHZDudvlGR+dYUqEsPDj
ZoIRiCyQ6LF27cJQJCvjp6Kg5CS71jpGFSbGIizs1WqRNLuTUAt5AMIs5HAUBrgzDmbUAJ6V2UvL
FKXdak9CxvTnrWeyLEj6AWTvk2+9wgLJlYtwEbiDUnJW0k2n3GjT2FxJ8yGquLp8O9lA/9n20nUg
eKvILKLiJ/eLBXepAnbSfJBLZTFkuIldKx7tifWVevt32nfpQvE5BuNTvsJ/38lTCkUbXto+3G5g
8aukXe3vVjxJddFRaBow4lr/w1bZ2j/xtCVF0DN9J3WzIn+AKdKq3hatZjVTKolkHg35jy2HXryr
IJAhMODR8MZdmEx4vegw3QzuAwyW0FY3GnIYwdmKlLLYhqTInQt76riD7/5/avvIyzpZnh8gKtrJ
GsKSM5wnf1YPezNzdwrWE8BPi+pBOQUJJPeMu8rAU/YC3IdZ9f0f8hadX6mPq3lcHpJJJS6EAdel
51/6NH0S7PaNM5Raeglynq2rHRS6TsTSF98D6p+6+UkWM/bmGRLL+0HpBZPv+SxEFsOfZz/RAOrs
gNL5OhTShU73oLfYWEdpiYxy70DjvUQS7GVEm9XHBMiohyj4oz3EhjTQSP1/Mm8PgK8Tj5kgqFCB
/PVeLAH/Mkns3ywRSDlHCx2IWRdonLBGvW4MYEV46Z6Mg7NKY8RsltAC7bH3EPtDBFXPEJYqO5At
7TZL1+DhvKVb+7IMxuVTHL5KH0No0wJM9BGWuzjWYYSsC5U4qCx56n7bDk9jcaIfG3sBZbwtRG5z
6MKHX/SGDSblUuBjEcf1D7R1hsZUidFNUO24caovanoEHUTSCdpn6NktUciApyO6E7nW0Uwttury
i+klxasTrswAhH67HzCwm8/xKKC/bu1PhJFj3G9uBCiVCWNl8/8oJ62APdpF6pqxLIbiduFxCnDi
7NleLliYCkW4JAOYOSpi++IFHuoSHjCqrFUBE93T5hZMZCMvkNnyO3ZAnrgnPQRwdJjVTiTFDpp3
Ham7uY9V6N5xW4eFpZwj62Ml2f07aoWQYCBDxGVw2CrECDE7DT6oqSdTMmsgOugthSNNKWZIQLDo
mlNrOyDrIAz3TV13/DfInqH5f4oCuaxyW09tOLhLz7DgZXbAcPKFKAyqMNlSc4Mb7mHwRBpmX7mm
yTcRL/UkWZznnmBeU6tfK5IjJPlg71Odd0x1mDGmGmRx8QLBVgmx+qJMngWFCTyr2W5w2xWX+N3p
imUfBs0LUswsQNxiPTORIk4N5pZgLYlLIjvJ+nXoupj5yUOq+r+5XbGkmHIqafKB4684ZSTK7PIc
NiSOb8qEuuw9JVugiiCcqXNAmE7ORl8VE1FQOxvRm5afBYSRQc4RPrZ4I7lqS9MtbH7cFu8dfMZ0
JBpho77OJKTxvnmCDoF4l95VDVa1JOf2kUVmK9V1PAcQ0vo78tVNlgczr//ax9AOSl7EdJ7e/AiF
ZGu9er8YYzyqPqCXTJzMU7yRe/rESkWtToEjW2fcui+CB8TvbxvPhXu1vWTHtAfogNXrjITrFDMB
gBkaSePCJhOIwR3Dkr7s/ENAoSfmINgA38gUJ1aFzxUuW8rzKjwwbFMKBapFVT4D+39sqfmFHHue
61Hi1pW+TiUq/pCT5UJdOVguwxzbeAD7VRhLUdSyOzQMj8JALBGcFgjnAu550ZkBOFQaQxLezU7U
KSqajplw0auXHbOkZZ2I9xaAawZVCTybRsranHQE7njFSYRZfIvANL/WBrXznDl3w8+FHZFQueSi
sy6XImwcTo8bSrL/b9kE/gXsaXDa27NjdDQcNuGggcGIbDwZ/R4/G9pbfHQ7vvpN9njuajfkO0fw
sZW+J9uZISux5nNUeYdfn6S53+EKojYVbRDdYMd4jrRl08sdUs5fIPbE+YgVzUwu3rZfkwppnzRN
eL/RYHKnfkcubdcEHJA1ObGIiLcWQHpQt4A2m7ml+KrLhnL1a/dsnCQL/6w/IggOmoYQZJVAE5Rs
jXaCR+JZlDS2DQUmzPROawC92hqnA+clwdVgAhKf1DtPXVUUG7JO2+N51wPaE6hBh/rUDQRTcG6J
ndnZa+sR1ISFhtVycgWJ9HOEmZUVksng8mKmTdGol4nBeJfEyyys4S7Yy0U5te83XdBFyBeGlOF1
JnY6D1w2XPas5S9lhq5zP41OkPpPO8tc2WPFoyfbfZrASRTNfxiC/QJJA8xs+aLhskgYiQp2GMIE
4mpZxJZ6uo5PG8q57kr8YkIR6TyfwH0mPZqew78HoW4gdzzWOQYvBz4YgYLda55eGCFGSGEO6oMf
cOghZNnPfFwa46SdWkgnPOESlEVTZRxa8gUQ1tjVyRaT4JZh2uqIBGfVa3MV2FpJEZOGTup53czB
c2z9K+T4v0Rg2sLTbAfRa5XWGSzO5G1G8uOZjsgclMtz/RGPoTGg3Ufn9y0MpM+WaVdUpZGKB/b5
gdlcfHlxqBwj9gsbMkjjhDNhIhLOqG+DBW3vZHtKYw5PuaDJJAuXx6dJF29JPYZ5+/h/AFBc3QER
v+hmI8AxnY1SPeZWzTh7RFathLolFq1kyCtQy1n+P8feKzBfbAib/R2jrjjd/vbIq8R5rUMH57zx
r0u5G0XdmWBWtViLQGafKMaUe+RRAeVXXjiaGupjnTH3sKwWpBP6Z+gdGYn95V6hXPpbJSb/Sop6
E3A9hk1kHhsp3RU8AcqNVmZCLNQq5Tu8hPvnHXqOieyOi2hFkTU77m1lacygfn+4r3CUbLtbCbEs
muVPZ/V6ym3fWj4pWEG1NCU4ehyCQ2GCLxWxIGsr80mj8aUsWD3LzzuQoF7TvYTs+E8WfzHzcWl0
TnRfshoqb6/Pc0Cjmko/5imJVDZ4FFAE4hNB5OEALQoi+I+UOlEmXm8iSBe8n0+5MdEs8Kob3y1j
UP8+/mBkJoZhCnzg8U/lQOVP2nC+lu43kaMo3qgN7YEhOfy1duqp6pvCzlvvM+pRAN/RMS8+T9iO
bSh3t+qLBuf2OyapD9C9V7fYD9SdqfhsmgA/IUNKZFTXmnMAnjWaBNlhSF32fjc8Sen11ZSAc9Em
99D7+gpmCZYioZ0j/xdhlBI5VpHi27NxczQm25uxjXgplCrnFinAUTtAP3WMqsnoBoh/dg4NgXKw
HfG7glih1TNL1qyL1YbrFiZCIRyt2lvbZFSkoMWhY4KkhxofoBSC1XXpVoBRl+h6WsZ9np2Z2b8m
i47pbQLOobcu7JKHFVog38mdoGY7RZfyRyNj2ftRfdW9ZlV1D1v6sCG95rzBkWHj8J1FmjXq+PAs
70jSWB8QEZz35gJ3JBkuuZR/hT+CB8Wuky8MXJoFweVH7XkVYOJPBneItTBWaOtZ8hZ21cAdrl67
BCF6RsDvClPurWl9n5h4MagVbvZq4rT3pYPdRgP4TD9SlS0KzFBPFV7gUJCeOkLJnY2q58AL2wq9
zBhOCBjhVirHAvh5rZ6c2VjoQYPNriZIdu6WHxTkYdVWCD6tkekqj16M47QuF3k14FWP4LU0PBYg
BDzBjUNviD1imKSg19pcPFbApEsoQsdgcgnLNEU+sQsUU/NsIfJHGJV+2rBBk4op9OaUPNL67sKA
C6kn8QyeAl4lAt0CsDwjJsdfrS/BmWfbznEuCMsAOqR39vLnkT4Gr211gCNZuiGyS5A3Z9jRBYXr
+ce6RfOnzM48ke6eGZ6VNChhKp1tzarM/WV/noS9mvXW8UY83rUin+RxhmNrfek+8p3cR9yHu/3L
HP5zXlBEbUP6l1EYfqHK9CTbCQ64sKDvpz80RgCQ4zsO08HHw5VWB6ksQPNVsGl8BkiGCIIPTZeG
wfYYgC1HjqXvZ/cviyJ4WKQOqNwOt+tWOXzsgy0ps1RVUsUSFDjn64oT30gmo/0y2SEpztJ5ex7c
Sji1LIPIjLhybeggn4AK/RlqaWrR5TfwVX9qJCup+0pYEmCREsEBvgqtIwkiyu68vSe/0nu9Id86
QDCUVLNCrgBzo9NjZfUPFnWeAdmcj47v+1OVtK3R12lSvM+Xtz9hmCUgiwRK4K34bfdf1MA7ialZ
ETw6xUOmz1vYok0+Y80E6zYjGvUrEqdZD8ieJ8FqhJeB9uV7/Rmr0nimeAll3e9X1Ja8YgKXfVzL
YOfZ2PzbUc4Y8/5DdVX3I87jBEEE3ADfPrZ4oyNHLh3qu2sfeZTS+A39P+L2WY3cuVqzMONqCaJY
tJiP1i8wzANa5YQGuidMe5tlDjioYL5emFW56BCNB8EXwdDmTB7p23lllAXOGUxgRRrh49YpK15v
q7J8MC0F/JR3xBXM/q3Gzru3ANw5khcJO6EZdl1Z72h717LuKjGLVU86F8Nsv/Davij8eLeWfAyN
oF7u2m1FfQ7ibx6H4yGXrcT3Ml6lB18XNFvqb9bS4y+5arifkcBxSCshRrzVg1CpNEdJpfASIDXh
uXNhuT2fxqQLy6WeifX30uM00Vx/qFJdIcfpxZURcSDyCCWZj55YSuQgqWdAQ7Ia8SlQ4BTbEYtI
Zvtdh4385YPyVaVFKsNYL9L/SYMtRF2mxSaSZ6lPXCQJuhNPvHq7RMy6h+vS+8LUNogz95WzP3Kq
P0k6MZy6ifS1cfTCKcVAdhu97glKW4l0bOlFBSVCt2SQxSEm+zo/22PN1YMI/O0kfCDiOipQVDGk
MpwCAhi02RSL6QIie/HpG/clR1sRfmakQooeviA6LfKJsQAN8/EWrEHSdj41AhGSCNfzu5L9cjF+
A3NNvYsbY6F/hYITWb7C9lN1yE9+vfgZn8h7gAaUp2NVKzBq4shHG1NEFvMfujL/LCCgPOC27HZP
RMkaDMniLsPllSA81ByPNBvkxcY1LVI0InMkuKSPM8rBQxTuyXlLsHu6Jc0bqxnoIlHHnlo73aIc
qGjbe1oYDAi66i0qEEzex9KcC+tuiKIwtumnzIRmACHkW8W8K6PUV9AyCIoFGzZyOQ2EfEg89T5R
v063YNwMR2rB0Ef7dCr0fDoRGYUs1YviVznr8Gk2cfl7cAYhea9w5TKLr4Ra7HNHxQtGs/w7skUp
5ex4QkUde8AJbQXUjESuAyIL0Z8BYTFZwHpW1dNZemRV6B7ZPs9hG9j4q16eeDTEhseUZHPBp1LF
Ls0LURdr2T4HZUxn+IkJgg59vR5ldZGhhW3JYmi7WJRCs/hrrCQrrrZllZIsGFyq2SfVACmuwmER
oY+U/ayly/vSlaG8xyZeJcSqdcDTIs3m/LQbz+9/F2kXaPqTfrJyhvbdwGqLrOuxHE79olfuEZ9V
8HqbPBOeIp7FNuti+yz+vynA9ymvHJk9OfPO/P39qtinL4tYT2ufBWqjtnS7yP3DquJmUt8T6vxd
w6ceVBKwwk6SdCG6LGHACaPQQsnxHUk7rOYb32eeo3pXl3qmQnnBxEH9W8CghFkzCms25a3luRfg
3PFyeGtdTAsY4dFqnSY3WX7KUVh67xzKK6yq1f87iEOXJgwRAYlBVSnOZYpvtjSVpoaYViHBunV5
Mpnx9LurMLBk6OSIqXHZxMtupiPuWVmoHLE/JraggO6Y2sYXhsLnqucDWrEj2K7SMPvxK+0sSJVR
dQjpqFaBbnpkOKufU1DGJI/UGykRR1TQHvC9N5GaDS+RLmzug99Fgcdt6qkvV4y3zTP8wSNNy0PN
O1PYqvRsMFmjY1Rjq6pO+7nEs2I9bAYPj8T+fd52pre7qdxt69cQJvayB+fvirP21fUDz/oIKIaC
LpzDAP44yWDcEkP5M6TjA2T3ZgqNKTQWLJo+BMzX9cH2oWd8j1N28U1y+We8vSqjxd6ihm/VYLXV
O7rybAADEgIuBDyP1uWKpGKHk5IHO/4ChTDG51YCbrDT6lsvtuEZHq6lTqcZKVlvEA9vjsfrhZEY
uLzFK1EAMh/9z8asgFoA8P82XA8agsD/hXYuGrgwKGyzQTzlGuTCVPIrrt3zcmA9c6AjL7rQLMYZ
o21pp37/uDl246XHrl6m5bCMd7ZkZNwdN5+yzssdWvZ+cGhY7B96Kq6at0u+ZHJT/gcTFa3R1ilN
pbVC1GDMgb3nEnt3agpjemV1HPIrTBjGu9MhvvotPtPn5mRr7C0JCHdgQAuk08GQnDT0Q/1f1Inf
fO6ki6qAPCON9zJmdvdTexrX6lf2ik3W3PMaSvqSrgzN5TMZkV83x4vyETtWVDzUEk/DIHBxXEwR
bBssDl+C05ALrOXaQYSwI2/7n083XQf+eQl9+D6lCJ3TleJp6GPz5S+HbharDFteOsOSQRn+/vZI
PZ+C33rIsv/xQJrpHMSXg39zzCKpYY1Jsmz9LeuXNQxZXY54N75rGxoLlWqwOTDvYVoXIo45Jg2Q
keVtv04j/wGVrhYGxmlOqx+XxO3hdxICPtbWwNV6HQ4Hbo2wLJZ1VwYL7Pylasan4aN+24FAE3LA
3+iiJPywn6Phstwrk25FlZolXojMQzwzioSsE1CqRPZq8GqYzX7oX34Hv8bRKQEiNZKZLNEH+63k
OLbqq2jhxj/uSF7rBk+9C9yxtni2M0el0X1tTmH+kK1dPXfKiF26jBidCOsJgCV7U58+U11Z8mFC
sv3Ectg6JwHLSEPrVNbhMN5yU/whGXN7sEUoICYA2TNzUkLK/k2sXp04YpoNiW77qVQPLo8w/tOM
WVEjPj+hBypTOM3w6FvdJ8SeGKW4vmhziq+Hsk15mAB0I+dGC8RvLc8fMHGR5CX7Zsi2Ontxrn7W
MEqiCROp/eA/tMO8JlcXaZ8fo4N/p5zsIGFBGGbMsCNdDsiquzpMjT8xihvyYvxmSpVlt0d18jwq
wnadWQTJVzcNY79PGSXFw7M4zIUBZ2s3tCi7WvsL6NAMeNMwC1afGvm065xqyoxciQfYZjVmTyAx
Iqc2BHwOMX/tq4VxUsn/+eKENv1v8Ys9NnwSDZSOfGLI4uTy8ou7imMGiWiD39X3Ie8alQCaHnKl
wd8ZEk0V0+CXyLFKINxJ/IEVlDw2m24Nb6dyNa/0xIGT1zHFI/tUiL051erMj8eHCMSWh5PDWIr9
tNLFaFiRrh7pHX+R+YTibZkq0+BSmgOWM0dmufw4Jm0Rgdcapx0VX+cgRBZ+9vkKyr8+FO++ygpV
tJErutGG/4ELoR8ToXtCRCM60YmN6hv0HaS5rlYyFlWggT2Ikpl7oaq7BjHtRYkY1w4dYKRBNRJk
lp3X4ck5k3rWMykHCtzaZIbTkgrgSdQcuYs3OOWbc5MMv4CcJ5vt9sZm/DFyYjYm9/IjDqA7cPlt
tA3pAphYpKWY+w1eNql5FV3N5qz+7fiS7XDZW/bCAnfndqwpbMcizhPKTm8vYM21ltlwkGT3XYq8
e/pjef15ZBej4pKd+xq7zF0KNlVP+au59tkW2cTAq10E/oEuo95lm9YPoqi6dXMK/TK+8rtvImtm
6zpH7Z81i23G/QjVRrfJUlvOdHP/BtUkxBPKdGpbs5+yMf36HabhLGQFyd05N0sugA8EYceYffzL
gAO0A5j54jIeUckp8n/1mGIMNQz81y7fET1I+PWL4OsFKCOyycWQb98ZvyAvnsDoSFkF1LEdPKTa
HE1rIinzvI5Cy63MviLwtmmcKqOBeMD8c5W4SBBbYuElKjsImRMwqvqw1gayAkgG1YMGxcMFvh3z
BJ5HItWEi8IRS9wQdeDmidaVQPgkvrWWb7y9yOFdfuhbdqfC1wIkToelIVDdAVNshZKUGGD0pVj7
ehSTQBUGqRCXEPSo4wBnEpHBnK+IY8DHk8k0ySVhS4ll3Hg+6W+QrvOgKIVD30/0IJDIHNID4gu8
67i3ncZCfHFBVDUj0cEXwjHmaTDA97LXoPaz5jNzusdRX9SLqEFX/k6GXPHzvTwHEPwyaWmKBf2W
ObNrp95xvPcNG9LlXgkQagovO36/S+0u12PaKzYWv+iZ8zPwfk/ypwvwDcZ0OI11K8dcREO+YsGu
/fE1q7oM5t2p4o49m4/73m9l1a78BeCM5gWQmn9YyQOZmaY095lxn83ffSHjEAljkz745J3H5GjD
Sscu9y+VsD7JqHe0sow/BhyzR7QtAICZzFP0zYSB82EJGTjglB7v5P/+o2sqmewMl93fXp+oZjs7
fzzn61mgtw0xkXTd27VLUs04/t/Xkmg7avsE9J48jQyX14GWvcb1o5WXKSSoniu7AeFiY7b5U/F5
Ty/uG4oP5TgwWtGdBk1xxxcO+dp1H0eaqyLobpk6kMMLMc4pD34E9JfPfBU2E3aznVT3xScP8/Lw
+GdVyS5mxtcClNNr65yctpBJ3bROX0yFTZut87sKMavE07aURQDN5t49GMNy6VKbLIrUMyCAqNDD
HrkfsekA8RoQ73uPeRxYqbP1l4b6HFoO0GxCpp3trkrPeYFERglWHjV/zXODamHnj0Ca7ff0uFfF
F/8O+jjj5YqWWlKAlM4g1TXXQJOYy4bPuhTmZqajYu2ogjn7IhlKfcfVMRJ2GxbGPl/0GvKeUPTr
Quqczs6KySSxipHXEHZfwMEjuAlia0VQGHOUODqbj7hBlA5tcvkHt0OcNSmiNDchagRLa3yDjEUi
xFPEx0SSrbscYOlIxFK5bOMbr251gUIH5s6ebwOyRDrUk0Z9Z2cSmFt8PaMGKCyvP/xVxrNFC1Zr
xniTLY/FkYF49Bb7v20x9ULKwaK/WFJ8i94qsy8Ie+gLXY8/SnWZ5A389OiQzo8DcIC+16nK/D5O
aaAw0s9ACVbs8wrjC87bE0aEM9wQH7fIDORJ7BaPuWXfmZqREsUHreUAbUebH8WKpOGZU1lMIwJq
PJvshROodeVXgh7sEzTRoZFhdp9VYrpDe6nk74afUS+lfLxbAIJbkmJAtU7w5IGK9bJvUb1Ki6km
W35YHQFRO/cuF5BSx14R5/E2vpsCtwH3zaseK5d5BwaNvKTVRm1wEmFI4+4tyic/6hkZAZUf0NUR
/wJsLkOgsqza0Vuy/FTtUw8WUxizoxI/AO8w5qUtF0Z33FFDW47VyUdf0DwlzXk0fL38P9TQoLqW
6JyFEZ/05YFwHTfBP5CIVJ1KaV+zrjRO+f19Z6uIJVabIaaZk4snV5GTZBBro/ZiIkfjn6QHRbXo
cCDyty2jVLMx7e0uVh8Hj8kBJW0WlXHVCnbe96eHpbfu+qV4y3XT8DYlWO+sNOtgAdKxd2Dl0PQj
J+ewmj2XBRjL74c4tNBZhGXKecjoPka9HeTbNqkT6ptIa/F9H+NtTd7WQ5OshLY+iXI0As7E4oVY
tB8Vll6UVi1ekPJBnYVhD2baaFeXfUzve2FaLMkR8ps94GTeFi7YjKXZZ/HJXRkfkkiYnmMQMnkc
aWL4S8hTbJCppzdRapnbbWdFP5IWLa8lbL8bG3mLRi1Gdha6D8VXZwD1Wn4PkgT5//xehAi6xmKa
Lm9soaC3+TK1Rgu150gXRsmN2K45XQNP9hXbJSojtrjAhzVp9+gwbhDcpKTzBnehGfBQrrwVAuMO
JUR8MuSLqIUi/sf1lVWYij9oMUudSRc4sZoIs/Bu57Tn9RuzLQycPy/U9V4UaS5BbDNtTRaH0LNA
eWltHxrIVqtc/NUW9v/F5CTONGyeeOGPgG2W0gJIWjs0WBi4cJHfPuOqgVm3/MJa8g0N4VGv+36g
xWwDzxJqvRscjGyOVuQLMiGqGmfjJ0dqMpz8MilqYwUiIJPSlpiqQj9A36ucsdEwDi37XrbXGTYp
aSh7JoIsf+g+YCTo3xebEFrERi39x00VcNUbhsGfLghG1QGd2g1e9ta8lQfr4Q2DTg4R9ztdtSIu
CZHqUOS6BEXVS872OFk/waXCEl3XsUuUjefeGA3Sw57FQf6D18dFrjSNy5TYU6dmDAkahCo2ddTp
9KBOFD5zVaCUOZo7OyKpAnpDrovcKM4SNrv/6OcOOP8VMkywX9jTg0sfZhK/OQDJMMrnPS8avBLy
mdhJ6ImZOMeNU7G5nsWW/2ZTd3SmNMW5ENKM7RRdu8rs1AxWQCH1AYWmJrN+BFbihYS/ob/DBwPX
+0J+ERR6zWddTpvN9sUnF+LaKaGJ8Rn5HGz2cdmuK2yVb7ChsEHh6b4DGSqivjTbL1rmO3xqg5Gt
YaxT9IZOv5L1NqBcaVDdmB6L4orG/46K8LFwtHx6cYwPbUbLpJ5W062+RDnu21GHETEohue/BLM6
pyxjUNGGnvcKWOKlREyheuyeAWPvPKG7+7GtPqDCmQYuE/6PLF9994kJh5CNPxxTJt7CzHmPMibv
F+UEUY66yfCpD2+s3WGYWnwabVhhQDz2Vey37zIPpgsa2T1T/Mv76uzIRpD3VtM5nXLK5YnhtakU
iB8y1buw0BETfF4sykSHJZKnzDWLoF0koHMJgRysvoikTcuwsvMoWYzBijYmo1CDtDuORl9EjDOD
U2iLQXI1r7HuRb88MrcPUOC9DGmIrLQc120/VyOn5ad8HAmQpJcVkje5DKvY3cpQDd4t42oX8Myq
bOpofqiRIiJdjWLhjxhMqSWyg2RhS3g8LjTwGz6xvgqu76+05u56FE9iFV1HVL7MT4lYFCB71Z3V
seA2qU/NFQHdNfzCCUhoURXQ80gR9q8TnjCBqpaXNL4CftmXWSO57fcokai5UoNyeSu0ylstbavp
YTibMXZf0s36DWcn6imIja0GNXs5pfHifhQVTycFoIHZJMDZpFPRD2dv4xb7g9pD5zQbt29HOzvT
4utNQcTrG3MHXIAPIKeIE7JAPHBWuLS+R3qbF0yGbp8MAghjNBGQ8I3jJntZvy3Ho6sXoDTbvClF
/TKlAAiZn+NLPyToqBH0wNuEIjgHJ5jqdYx7ELtSSNA7byvHi6w3JWLCTGcPdSx7GMYHa8TH6kr6
x5CiOzox/oe0Ec1MhSHb2vtIVU/0m3OLebYpmPqgALZZHWi7sfjnVASuxp2bHEa9uGMUclOtSLLx
EUcQriQ7Ia+TYJaBYZzq7z546Q7yagM6W8JrSyoVt4tNDnjYW4PIDCut3bTYRz3MNXZCauJctaOp
e20uvJuLWW0hzTo92H7umRZajATrfOwhs5GTYIu/ORciOuHruUvX4Je1HHijDC6tWWq6OYI0irOR
Z1J91sdqbR+mo/f7tXUxgh0BF22IZeo9wn/2KIBdeEG/n9RMBxkWHsbUFxmRby7y3sUAOA1ZT/1V
P69qWVbBP76NIIjch6Z2pQL0ZFOW9J0LhxxMunu/s/8NQiJIff4kH24cVDrlj7Xq+O50LNgIVYtI
+7GSrYtjYle2Ri43MqqGFqhICp+H+4zxgxJNexdSppUtx4tOCgIC7MN9fENQ91UBGEnAc64tA8Cz
YNjfSvZ9xJMXTVtwiIesQ2melHomlwJ73eV1plFKlqsfYNh5WT3PqNF7vAqpCMe62qbhuWRUDDvf
wDUooDXUrix75SGREAUNpOhPp24VT4l33jwSKNWgYXvAi7VxG05GZ9lATASZzcrUOM3bjpb85tNW
Gmo6IYsr1uaUGpevmvCp8ZjKYYeBbpjIGpakWiIIe6qAye/7fzbfwRihH+TzNaCRGEFOrA+SmeX+
R9NiOKaWOp0jmHsZXB2aGfKLh0Kn8uwd2dOhqSTiWNDj6prr7VJlq7z0xWFF3eJesalV1t/v+sFf
UG+dX7Dz7K7CZEeNgeGRk17vs9oFAdEavCxYMW8EiJmmc7aTOtnqwtLwnFGtSaCFG4UZtnflmCv6
vPfV5/Abs4hsclO/lwccmCY2gEUrXlKpMOBPwblJR+IwJ5JBsnYmVlE2gaGsN1xH/sIM/ZHl5xfh
Ews1nbKHVR5ijxrbJYRsMvsA8vIT02uAvLtulF7MY9z2SfS/IOx3wmTbWrzMmTGYS8+FkOv6E634
8ctoJQXq/lbC5VGFQc1m4UjSPV7zu11NNqAJDs7WqPYMjtbUJ17J+WmftXEOWmNjxTGvVIDGY6Hw
gm0cQ5ZCzp6giNYMAIfRpYh/P8oBLp9/IkoCjuW4iDl1Yxr/Lqq3IBcY9fQB/BTxkRwJhdJzr8Ar
BjMjE5uO2AWbK80dH3Tu3m4ZkRQQGi3qL/9shTy+7blDMTu0HWdfdBkeIUdc2lTIRuI9c+oQO6CG
SK0M6wDA1Q2gxCvhKVSlAWFMusvflnbOlLBYbhN5V0D1vnKbqyBakysYGJU0c2DmhcfF3YIC9HHV
iUgkYemP8RFhvTkpVvqGKRIqyp7TfLXlCREEyL0CysPeV48iOTr0b2KGnGY8iHoDzGNU9BGQZq3j
Y/AZv1Ueg4pkIaWRLaawz4b7alJURmdD4gikGgN/97RgOuyMUSBV6HqHAF1BshZC6HujmsbRg5gS
oyMNCP81xCpfhBWYtq3p5syNUNCA/XmDlf64nj93TtvVy1i9s0DqRUjw3g1px0YPCuzV2jZlSQa2
YFNRChbvSnAWPd2IMHgVPXdLO1uKoRD6yfvAAzIqffqeSkmvHsci33rTk+XFvcWQtzQMf/AJP4Kg
Pv3DBIw5E4KI75rN7R3jfC9P7GoNXoGWVMntPaaeJ1VDmUF0TVYlKL2XkS/lDHQTiJ19oIuvdpF4
0vm+I8GkICtKoHUm2BvDb2KyW+zV9+XnSTO8tZWiC3wnqANt0/4CrSggjr1pvuK4kaxGyenX0FUW
LUyCGIvctXklqHstu6wWEKCemnAvYLXLg+hB6de9cJvpe/41K6DDDbHrJfDmrJdUYJ7Uaea6hBMm
3YHSEcE9oljD7k9ba55L+kXlP5PhA/CU4Ob2obY9N3mobLnjGRAJk0gyRiZarZ6WG+0/6p+kKx/W
aWnoO6aXJNLhQ231noLJlElaaMzyIofd8ia8u1ZkbR/n7a8gfnTQq7EGszZDJ4q+mz+X+bVUYw/d
bydlgTi2t8vw6GtptleODY4V3BPpOziV7qgjK2rUpDerPjUAORsgnflE4jiOKzWcs70Nk3bFXH+F
Hpa5C4z65KN/gneEbqfJu/1bxik1EEbQ3xwtIi7g76cDeDZ74jYtVu4PR247G9g5kHjaW9q/WFIy
rMm2svdqIfUi23VUW/5WVqXNCYvBmyT69fuMZKJVDterWOhV92IAl5wiRPsVgF6Uym8hiG2/JMpj
MPDLIIAAwNd+54+Q7BsDZ7KKAUHayyf9ldH47cy2cH57HBN6uPEiZnoXdMlk8cfqm/C8eQXSdEKS
3tZra6WGJHPOg2gyzSNaXma92Jnx/4L4HreVdEJa2x8+6Si20eKdxgTGigzzi2/NtvS7YMcge0Wb
JB731hNKD/3fDgdmKO2Uxzz/9hfll9IocnQBLU3foo2Ep7EPeZT0kx+HLOw1M8AZ9Fp8ZjLkMfc0
KTBOTIs9Y+4gqkp5ishby4+9O5l1wf4flmjVAV4ILweF/oUGD0979gQul6lT+5IlEfRx6+o9xSV6
7YSgKXbs+MwBSXS4K3+YGoFKM8rHMUKaJ6gVZdOOtEp523Up7D2cOODyG67GSK7s+G4Mhc4gcrOR
L/U7d5+5/m9pj8my+RnQ1jyfboQ8eQ/kZmafUzuu4bqfmqItPosh4NNmYJYUgMmSUbYnZxTu5w0Q
osEz6m/5iNIrzO28d3PlN6v+Bd1zjvQFf+Bflg8vo/nTM/S6T7I0y76nf8/f+RUevQbMub1m7rvD
YWfPkdTt0VkQsA1ylhMApAKcOVASSrQ0DY9uJ5ocPx3pQTGjLL3vn4zL08/izgPSPKzz42YBAZVU
YVbIxavosrhvvXHHa4UKf1e2I+PH3eFBUASb1yyCMakJV/f1gDlKK1q7GBArffivrCHiKmS19QpI
BSzghW6UJIGdvhfKupF8gekQL/IL0xuz4JuH2CsTVVhDfnkh2kXRWRLIpngqHFtYIrB0FN6aZ5az
dmYaNH2U14Rcq/n+wvsNEfVrRdCnV4qKTrL973P1CfhwimI5bUK5tEofF4ZVSbgyp4QgJ7MwUST8
bWXg9YVbnxgDUerSkyzieUFLh4I+G4bBiW9vn7VTdtmyD8T/TYa9eZmOwecOwPKjneKN7DoBh1Ti
AacnhuOyKzOoBYMO+cDxRreFKslbifVOS7d2AHg7C/nJiw0qlI/YANx7Ab9CLOkqtlhBMb+VCZfo
NUeKl+JF9c7Z+sRCXL7CKIbkwl7XqbKnzMd/KESQCUuyeMbDMu0mcgVKCvHIaNJG3J8hWmm+z08h
Wg/H37HmPbgNUUDBiPp9nEAfc3Ub27bRmH2spQv5mkKsTOO5IrkmqivrECQWofjaCEuQc58zdAE9
k7APAAO2RNMZYU2P7X5MHieSptGdXvCMTXXvGgU0utWwwxvpzsQR5TSnTGy8yuKtt8+iVz3+YaZU
VPbh+Son6MwIQc+wzG1sQke6/aqu5cW3uR+iGWEoj2A/dvVpQOtHi12j8KKr9r8KoLchJ4vyV7C2
giiQvLSMsnZ7i5BA6fQPkp6kOWo4vu4t1H6y2D2rQ1ZNIYg4gvcyyYH9FdI4pRN+loF3wrDKdmm8
xNVyeC3fL8uEb1T9AmK1LhgPM6H/EvWoOOuHIhmr5zvh9bqsVzYNhzw3UEvAW1pVkqoaFOAC5zxL
yBom2F6GrIdkPO8GMMtDxIGCPL80bXL+oPEEXbUcggNsmTBp9nkTEX128HdH5dgeNKBixM8CtVJr
MUypHwvWuNWwreKzhuI76SEBJo7BuEhmPkxX787/rgq2zs7kUQP2HAwEfI1mwy+dBvC+zddizDNB
WZVNJNvK+FPFUlVdzMpns+uEORaqAhDz3AjquLKs8ZLYKlfeZQvjjAeBH5GfOJJsm+Xu0kFRwQvT
UAGuJ5Bp5a8iVgpi4M5VETlfRh8bylifWgSugN6l0hCQZ4yFN8o3mkkPIkKZnHm3jloR3t1vqd7n
lc9PfnnxY2rLuhTMsei4L4Hy647/xq2wDfhehr/LvFl4VIeBFAszUv351TOcc0QHWirQgg9OS3y5
rNWdQ1B8mI8hEGlMb9sOed7R1wjkr/RTIEAo3p96JQKqV+2OkyWWv7Z7vIJc+EDJsScIXxzATOAx
7Wb1FuqP07NPugX3WTx5+LvfxFzDj0pLcL59o++iXnt/IJ//oLJJfXiagbSO83BvMLRp112H0UcH
hK5nit7E8GxY04/l5P0D++Ufnk+d/VKp3bMiwDLpxJdPZTfDuhpYAgFgyZhfrUzva9yX2Je72Qy0
C2purvQcH1NZMoKDaePz4lXEpoeQtOmYWVG+PgiUlrlvV9esN+dP5IVBfx+gx5KFx1V1IbbtBwCN
nQhpAx5yz63AOjXHMZncI6+gOc2c9Lx1/35UaZgxfVlHa59mxDmn4bUa2bNoWgF7y2Zon8Vfrbqt
yOfGWdskSJ/7AD9heIWHZbt+HjuTDuolHBBnE0h/w7KWmgBxHNdLySbW7cETjjAhJbYJExRQGXhk
uA8NixohdN/eWh2fAyePs1k3+nt3nKW/7h/vBAY++WBN8FnCQ8e+5qqz6J+7Rou5AQ1BGCb9/ODt
jjqZmmdrb8NZjruxjK6FT4ctRHIxXKylkXvyehz2hVZJDLf27njmBwTlEhrj732oTxMqBrFRyI1R
rNSEwJ/HKpNcNgdiX4xbNsJ4c8PIAcdKdIdMoFVtaKuet23imY1VBUHDbiCgfPvrTzdfzHXMfTCZ
3mZ0zqLwoLJg25y2t1/oWzB/g1iNIUho2cEW+H+UMEJm4Ii6wzcOOQ2hNKGHGYmeuqNDrfDKJwdc
Fhkz0WDoBoInwO9vE6oUi27VatI7cgN1vN63RoPdN19BwWshm4APgiec2Yb6bqoTK0XAxmWexgyG
SF6SNR9Kj6pnIFYTPvM69PXzGizaWNgOi8ZbdLg8Qpr47OjD/GovGlK04EUu0H9wOFUwU5y75gzW
N5IwybLDpTP2QuP6nRkQVQlYKo4c2qSbmXP48LzXq3x9BtxMyytHRskDA+7ASBlYS1c140sLaC+X
EwiFIGr+CqC+yB8pwC0bwlVy/Ql1+c+1gnqoMNoRfv1fsUsZzoCA/HeR/eyCCLHlkupd5+mUCvWE
r7cHLLF+tVH7QFIJJTOpKucEIjQYXrllge2KSdhFhdbpHE4lIvxbFnykUy+cgLs5xy7UB7pxHVb/
WoasfCoqzwoZdCPIlrD3AS9t+aZ4dFxlH+j945sKb8/SsqFkzOb+WD8ia/g7Se+0CqI3OkFpKZ2u
X10goqAxrMcF+1gvzJTas6hFNLIKLIwcUzld7U+0FHw5Umzf6zE6lEuaDNB/nViBvfrIGJ2U+66j
qssLvxZCR1XD0mzrHmkkhRZxKFQ43eTQCKJqj8U+DA9ngZPz4n5tL/Z5d5lB0nUyyw3uGEAHHWhJ
uLfefDWzk10pZDGjiHQLcNyDQ2pV4qt7eCWdFlZQhUd/7Xs7T8ki/vBOwOBQn1RpU3Zy76+0C+YX
V+YnDDkcE/8Al3LP2lt+Fh/m0r3Jm3I9KyZp0PMM/LLnP7rfRWe7mf9lOhzsR3O+YHTZN7FYcMxF
JB1rbSuDklQ9RMHqYYx85rT/trbs+2YHgwfW8K5/BCLXv5DiLpykMSJ6Zizm4gOeuaGLiSMlVypx
cTiZ2uId0fjmoMkkI35dlkdAUs+NCSmpgl2bEc67aDKVA1KsLXeKNrSpY4oa79s4vNzhxiXHd4mf
7VxsZzG+H+ZCFnUn98k2yN2IUHBASG4UthJ8GGYgOaw26G1YdaixXn5FEhNBsECK/+lVsaWBVdke
Wfi5MkkZpGjQVtIFsDYuO83Ve2f/z4EcTDMqe8k/eb5jUrKAInMXoUHdx2TEi6ZUkuUvvEyUjTOE
3izxPjz3oXRh+t4Mb67JL8mGIjHZt2Wj0iTgOJ/2Z7aJL43GbhNCzLMrHviYWXJ5ilc+L2ml9NM8
vN30eGaPuZWopXh+q4iABWMOjJYyhr+2XgVv8twJ0HtBOQ6ZJ3SLswpOKg1wKYE7w5TCgVRStD8a
6apTLOdiPYrVVzyKbrhutn8vetjp6GEHJyUmHusMsAbCRD0uwP4nK0x4U04F8yGLYOXS8KgKkc2F
U/1tYGOdLSwt/JND+Prkr5VeaeEtkomORk5B1ieu3JNNNhaiU1db0+ZuvE1N/tBdPIb1Ds5UrLlP
4cZPWBe7cchT2mNqDFS6Y4um39nc4Z/XVUIjYQYGOQb+TPswe4wL1U2DS6TwEjcaSFpcyi0zwFlh
FPj8nIlqp9RU9/z7m292V7qKhMyJxuOKRYu5p0PEHpqu8tqXWpVplMFzfAsoMJp+jARfQGqucB2a
aPJ3ZkpDD/n+fsl3ibGoPrM09mMMyW5AQwidwuhBjnmH8pIHvXOocVloiU6u6Vw/zsyfuwdNG1Mu
cskGb4oyOA8T316HXUnS6nzI9F7DFZSHUr7bifVf4KRMoRLGvrChAu/Rrzdx+J3tWYoeEMdQJTtw
007fv8Zc7zwBtTtg8raqsLN20M1+lwgK5h21mBz05pyJhEVkWIm4CmJf3iNpG1Yx5lslhxGAD33w
XuVAeXIyyZHLxlXZTP3zX5qhJgAObWtIoIOvgKiGAE32eWcm0xOZ3LpJ2F4YoKDeeZSpivt5EhqD
P+ZPT703lup1R1/pVg6StVq8TmUhJ/bOJei5dXwM5T/N0K6cD2O3RvHKu3pkZ6zD6cgXliFJ5BYW
XTviFvZfQlbj7WR2Jr4wrFYQ84aTq3NT3/4I+0vVqq7xkgB14qxgjSLYfPtLcpUXQpuBPtoQabWq
dU18Ci88I1mpA4Tbr5ultV7v5bVkT6wYh89rk762f4z1NKwMQksAixEHhiMHfs4n+DzxrtvByfS6
7F6Yi1SI3WqHTocMLr46PjQg30AhFEwH2CHue6kvegIzCB4k87Yc3vhshYczlPPuqe2y87in0pmC
yoGuNaFnLhhSeh+xSsNISScJ3XYJhWBv0aJfoAU13HqyEUwN9dVLWOG5SyfpLLMzUOfyZ/aSKSEA
bYtvCaqBzp3ExYr54pS2SdhXNGF0NdQIvcVzwi0fcObjCCq6ZMJLIfgDvaV+9ktFm2yQ1TF5I84f
VJkgs35RiNALP7TU62t5p4PtB0YrlE+TzsLpLimKV0HJ8sXmH2mxz6fEDtLVyxQcyZ8VNam5Jbff
bASAUPYosfmwtQ5lgKOoU8NmdZCU1C5FMUNRPCdjeqiscfvmFr0M1QmGDw/9moH5Qz8sqV+a+ph+
/sAXqstnRhLhsp50MobLZl4k5XtTVj4/bR1+JVgxik4e0VhXvSmhM1XDrrz83EiRIduhWQRQnaVn
n/6xIXJ7nh3ZRdCOePRFehZgZz0Cn0pOaNvw1OO33B6mBAraKco4NKPsjTbfIvAbUfA7HUbhvZVU
IJo/+8lu0G7PdXSBjjQ31H22WyUJV7p246lbdtxBVH3GSMQUhu4w90ZyhOhzvWKfdYH/QFQlnW9n
d9r4VCwQcGrPhLTD+/g0pscecYCO0okxGgeNyUdDcgOPAHI79Ya8AW67DYHrtVPPAxeqiH9vTb0n
IcRLLDfeBLUaizWiYh4ycqpazaYO1vM1An9Ks4Osm7BlwQhcZ80Rlg1THwXGig7osBvpvDt5OOb5
O2XfpU1bqJz5pvcb/I8T+qGkiLWpVJXlw6OaBGkrIACTQDTA/bD+lTre7uyWJeBpGVBAWNaeIwJi
EHfjcS2mgWOl/Mog1ebi3Nihx1Zxn7WUpz8NjtxHTNg28Vk7L4dHirQHR4CNcbZlH5VgbPIe+B8g
/udE0Ejp9HIu3Hxe10KeFTxTqpWR/IhvDyzFwoPc30hR+oz2YHhd7ki91vmhifA+/10rhJqayULs
uEDfaVoly2OgE2GtoM+xtPvpcImh7wp7bd2qe3E76vMcg30HbxdJt0ZbgUOuR9D6d5NSFr/37tEs
2oEXVz00GsZLbpwnLV4kFKoUgtzc/OON9ZQwOPWkcRaqSV/lITveB9omlzBJnmx4DeDJFTOS7ujk
s5maslfyvYNrqK7NZdyij2ulWATdudmm2gX8LNWfFkQJKvIe2M/XYSPD9HGCwfbrl+Vke0HgYaj9
+wWrl7nKZDBlHhdA6YTCCkLrD07xaMSMzl+CrMf84CS2o2Il+vPfZy05uI6THXOmbX3Ngeq+dizt
JSMM7lxhapyEFkxqNUdc68eakt+yimw1ncNTslhpNR1muzTtZLw2z2wjwkni0rMwjdjPoTxyj0wR
ugkcO4Y/L2Fw2ypZuWKJXqq0/TBXfoivOy8ZifQY83AI+hMIoRnA5cDhuyUtxRbicWDg37BQpBc7
YzKxbnIPxcQqax4TJUVUJTxxaGPEZz+Zg6m1MP6OHsx2+tiovUx0nBVRe5ebjAAdeqvkbDiAUJsD
erQmDIK33Q3pqhm4W1ZVZT8RBiW5GIMmPyONwi6xEI5cY1hr/mzUTLjdXF2dZp/AwzqL3E2rW0oR
hsE8gJXGoJzdhsfpuXl8ElEupV57v+xw+FOf1TsaGvvvB/cxLB6vRUxh0cdYSbFoiDiwZTE1mn8f
qI8vRmIzC5grs3uOw8udnBrXOkBroJQgzEmAEeoCvDjs0XZXJbZRbdoxp+pxxtEtwZ2GgS+uikNQ
GY14Mo6Rj99NIbLjb5Ge8NTmUIQZp7s7HRtUgP/r6vbvX6pXTvpIoVRUNReQQdbbpA279EQ+YneL
fcxUeD3sIShQWh55XVqz/6pWK959Nf5ACFWJTZx2/4Z5OY41hTwE9GxIM9dPV8o2GjfTl3sJlJ1m
z211FS2uUUs8NLdrkviLcG43r8SFQmM2NZvhJZUP+NNddEAXZc8fPWzXt5QpDkb5x5iKTscSXU2K
OwFrwUmSze+WxN+6yzZjnYQM9B2Tr9ox/bffk8sxeNV8+lx2vhFBa0rElGaWa+jNFf/x1zO0VSo4
zBEb9w+tv0XCGHzQQYoepZ/9F25QQXz1dWtvMlL1ZpMi+LutGggXt4OE7TWau3lBneUwNWOE43Q0
nJeArb4FsRDutC895rAuGVyoKxSCF28RJz75iiibTGK2HaQLJXD5MEkld3m+Byim1B9Lge+X2ke6
Vhsy0egRkT9oOZNg37VRzXIr/l8LRuVr2oOTQPU3cpDN6fbIIbr12+fXpBSSms9tLryhPyNpL5AZ
CHYsACai7B3c9TscCdkx+pMtDQYnGK8aSzmzCSvYJWH6n6XDZaKJXbTja1MWVkUHAe2oyubf873a
9xL+q6drzuCQcqTV4hlrf/mwi2BewsiAceOLiedcRLpHJi7ypMREhGNvBwjiX0RhR1FjR187nkWc
h8EpMNoe9F/DQ3ArXnmPRMYTQUwSen8njHpjQfubANFh6dNMsEmA5R9nYU5Wl+N1ocMRg/GalodQ
xAoYD9KMoFOQM0TJZI2yQ8eILsGhFV/bJtQy83krytvT3ue/nouXZkUNmghHABPIoD1hSYg4y4b9
1AU0EGq5RWazcgbXHCJS03tmtJHQdKayO/JCH34vZV80rxRlGHP9j0UvK3a8JvuYUuBajI0Xk0k6
SGj0Noajwunw2SLyUkRjmOLK++2v9QxPUaiOgZMwQvhCNwJRNFHSQv8WbzpHayp1m5oBiUtB11Uq
bFdzfrYT1EXotzNr6hJiF+1WPi+cVAdlz41fAIKGycKMM4xnK1CeJjvPQ7s+5qk/UXD/t0qrhnEB
itQJaehRPj8dUSylvJxRpvBJIfmxH60sKoKPXvpPqY6Qwl2z8pnPw6BSSfPfrQpCHp9E/o4smhMh
lwbC2UWMzK/1DuX6ITLUTVYowdwrGT+gF0TVlQ39OUXYb47ZQ4/wZ0Gk4D2i02ARTCSAfEaYQIHg
kyH2rZIEz565uUfMZKC+7uWLR5UenzKFqF2mlrNVtxb1u9ulozN6gvsUwxYVC9tjbmgpj0fuDz/Y
2v47+4MP+fxtEGizzLNVd/uDZRNVK37IUCAU0UybS25BNjjam7/oiI23IPziZmkIJYbF3Gf0E8LM
ZUM/vyQ620HlRKCpbmIm/CSMjfW+E3oUTIV+MNpRWwr4hCRAUrt7wC+wkh+NWdzuK0nASIUvkqjV
+u/vYojNGbXPAM9s8GTQWyb80jkUqYdnFNxLJOjqEw+0MgQmUujZ84YfEJN5yDh1svJ58ve5YTQ7
6ttK/xHCjSxNQBqdnd7HuGIjcTt996RwAAPD4PTuukY2Z7qmCpy+KSXlq2Gpctzhf/C/rOe0nXsd
MHN2GrmPrYCFYqAXh2GmPZk4BfD60rJELDCehBrMSS6H6dd/bllur17Qv7IZe1iFb3E4P4GxCLHK
ftHIMNDLEX/E3ISyAOwBGwk/cN5wwJkuBfOWn7hotwUiHgKFCs5FpObniyHvLA6LU+KAw222LqXW
497vllQFhnv1en1JhLcyzkz0musnUb0ZvCi8OoJWLuXlwhqS6ptm3DAgUPRiN/ycIh5Ln2yFZaQo
loX34Ok2t59l9GoDQQeNBV/BrYALlUviHsBkmx6V364oZII/Dvw9nIhSuuCzY/qBf6voXAgznAbH
aliOvslNdK8U4P1ZeufmVb5IYWByRK+eyv++y/HB3ERkcIMg1RyRbhpoBSScUMPcCietE4vS8Daj
7uMpApdPV44Oj1ortiMzO9VvOXmLSW2C+XamslVqQN0oQLvREzQfa8DLKO0cZWDGsKBZzvXfHvVP
SseVvUZ103kxGoJxf/k4ydgkjMM5Qng8jNuO5oEd/c1tD03DxJbYasg1TOfI6xfzgkr8Lx3MRNNh
VLoVLiHunpyFewCjHlKlPJmcYYxoKJ1dGAoot46DH6LmW9FeVbXBYiYTSpcJI0l9oSarn6kYym0m
JmplOLpp1IhYBjUu0zMM3SLuCI/tNxmAlf2vU3G5ZRnrRpIvHLBcahFt5QV4SO9Fk65JYPlUjPb7
Mj2uHGZcHyan+VxU0XRFCIiAAcNHKi6Vc185/zwd2SgFz/SM/KFCipGxoGqXqySUvcQMqd9YK39v
GXmFkdL1Kfs44RTcRUpPYLvRhZM8ECg4vz2BXEwS3CF2WmmGlBNoafxBukGCuQXcOHLaVNWOe5sX
SmoSo22/jYlblI1c5Mn9ZpSq5K5lXVOSMBOlsvs3FGf5pQJYuWcSLdz+i5kEN7OW6ZYmjk+oA1Hi
slLkApb0o6lzzNXMUPtueVRaQn9q58vnzy//lUQJQgMhCLaEk8WrFBqkush9dt49UbfjkV06tKCU
ZkjTlp6c/MYfsOysOJ0rG07TBiXpyHwlN2ztvlOT5fxgrGF8aUgZHBmZUnqeBusuUQPrUArUaj2b
92F65yfmqctjw7yG5BQbbT+naofPy/tLs7L1nk2qoVtSycCZyGRgPEF58GLmIUP9uHiPP+ElolVF
R32uYLKqq6DmwgzuMXS8xgCwlJacuCVGaZX/4bRJQFaJzbOU7Mb6YbzocfLv1bhvAnMb+hvJU7rm
J+9by66M9ac18Dvq8FvQjC1RD2MDIHs2y34zBJ8+YWvIFR6B4sgwuosRCFY5zNwX11Tp/8eaXYrK
L2F3CGkM1Bl/t/QWdiTdeCW9q4JFfK2IC1bPpS/SEkv0qL/Wy8O5sP9ZX89fhhj1RPDTy8N/tZhc
AAkVhsnd7xHwt0NL3mmI16FBgROOC25M0Wf/P/Svjgawu7RFR/1iQx7gCwG+tXtwKtIhHu65JNAi
SlXntEuHgjXJMn5C/w+TNeev6wwo9B+aeo1qTnpEuNsO7rtWsPt8CAlX6oc97SiLFn3OjFpeXdyv
nWoHuuuVB49Y33kB0R4NyEZVlQ99+dEI1bHqRRMOQMTNXBMPOixeBzDW0UsESZBHc4Tvy3L7yjQZ
nmCYDavPLHAmd6eW3ulsfCv2hqT7oIKZhlDP9K0kVNbBlXGdv4WqxqYsYCiG0gzh69ZxoWqUfAON
hgreKjzvVnYnOENLG8XTG9PNwM27HvyzL1X/hEL22m9HMcYVzXpFwEZyjLA3iH4p9ykSATGKaKZ1
u/qE8yK9i7P4cviNh1CK1UHrmIvobk7P/vbKZA1Itd/406tHNA54RCdSzYl7hTtT7aagYT1X9Q1V
its83n0mQ8xFhq+lRaul+OigN/iEban2saNLbaVqc/0QwANkPXTayNKxbS9xzi+VQ4P8Fx3M2P4r
WM7rvq1woezJHClY2juGLt7ouKuNoRI2SnLfOTIPIt/HUtCEogwBl8Z5kx1zWbiYTNE7nDFckycM
dNdUCE0ayMxufpbtKeBDTB6HQ7NCRFbSzq2+S8VfoLShRbIuzqMYMOwwqa78n7MGdn2WtwOE3qOY
RXgzCG9W+VvafW/JN3S57O0yZg/Xxa5HNJGGOCmCYGTrAeniGNLK/wyWTJOfbkvnC+oj9uxRnobR
QcTI6pPegLxugGqcJrCzwslfRxW94yyhYNL9vL10IS1W3XeszMIfdJyU0ej3FNPql0v+YXXcigRN
9VW0DkZLhNf6aWadJbHyheOlVI+P0WBzENo2VscJlhAvQ/r057QRLotBgifLQ4lXZ/sEBbNonRgB
39YXXuLYMeBZoijxup0wDxFpXtRgSxGv+rFuT7NIuXu0zNk7C6SpkW0PVeyfwTRD4jr3fi9T4PN/
kSrfOxo/2FIHvMH8ExP4nhcISbO97H2F0WChBLSyNMLWyk7njSuOi3L2VgKbXJyo7LSBZ2JdZD5m
l/RAZaSM4ZVDmwqpj/8KrhCRgvD+q+oeswBGlGbrX/MjR2dZ0Ag/B1wTLMADvZyGt2e/D+LXnrFV
fJ2yN7XJhAWq3JUqTX+NhHH58K8O7jTM5VqDNYrTXSk7Pwcb9CCxgTcyl3stCYjjCd0b2aARlu3w
ablA5GXKiAijZf6Lh81eFX9JGNO1WMj1dAPc/d6s5wh2cnAC8zLiNnXXdEMRskbndd9K8KcN+aKn
4I9gzSW/LGY5gDCq8cQDZ7t41jW6A0G+hz3PUq+AYcQ8f1xljOgfUuzuLKKdwIFB2ZpWUpyRF/Zb
qFJK8MPkmGJ4efVkdaEcgpvPk4a5P+CZ+gKIYhz7ZOSZKqeA93f4CBZ9Nv5Zla7uOyn2x1GL+5+d
27CHiyp1zQ2pPt1yOz5XZ+GYSY2oF9KLdL4o7+TVylAD1vmXNX2+vMy9TB8+wbirt1y18O1R9scR
3UZZHC7SygS5/RK8+g4osX1SOYpvhljkM0WMNdygWuLQHYbWbhwL0jmg7XbFS1H088m+aMXjHGWe
zw6UmTMY7LVM6vNaUPJQHJoSbae4Lbrb97rYms5M1Ku+iIKh5rLb1K1CQh6f3FYSL+6e1rVXvc8B
QtHAzMMnVjKq0cDm0ZrGhgcObDBsU6YBXoU8YPFPpkGDChv7jZLBSv0DY057dlh7HBfWJW4PcWbJ
mTRjOfrQsMQthp9/23JeP6VECCjqT79Z1IO1gkH6oghXFN5UJ7qo9nqt7gqDaYV7JTbva/10qOEw
TRodXv8SF9zPgoA8bi7P+nfyw0w49tOQJwm+uXBtwk1jsSpLNT3cFTGL8mIr3Ru8ob9vCJ3YYzIu
HFIBY8WZ3tEGM7GVTaLZSiHivdWN8EUbvCiJhBX0JfBXDbOp1dr1XFhrQYdm1SSc2g/NgFAWnGY0
w8PfpJy0wVEy0ZMOGg8KQtjB2t3ZEQvF8lB97yJimBXAurLCIGcmIEyfpalCseqaY1DH2VeTfj5R
BKOgyzi0s2eSZ+bTKt8H9iBbiOsq1AB/xteIdLR2YMC6hyk1En+U1d5e7SeCeM42xoxkHTB85hme
nPgGDQZk39w3jIKci7CNx/GhumI0b9xVI/cOOXC5BOJk75z3DvHEWt5QhOLs+6rrPJz5LODhBYEH
ZXsSiKedAZL1Z9rJ+2iNy9ICPZBPpBfJbci9gJKRELGaKole1x9AI0APQUaFS96pM3aolhT/Si8q
B2hmffKEZXmH2BIKweLyYiKWi4Qb/5ZzZHKWJV7zwK7WR7BNo+3nxqCqT6zx70Wet+wc7NjvZfih
nbwhPm6gWUYoeH+9zC6560IMBbngCtouo3xOBZl4BxE9aPocW2/QfYqr/26yb/ilh45I/xEoP+gR
M1bMraN8ya88YgeB4UxyL6ElgWPXx9b3JV5LjZrZIFD7Vqi7B/U58eDDXwMkJWuGZ8hYWB6qsaEJ
lGvOxt0kPlAJeWBC87WAnqedowO85g0cR7qTrzopzylBziD+v5NJLrtfcmyu18iK7wkD93IAe853
pasALrc3QBq9qxmPatipwqu10jT2/O7aBZDGuJ48JSE/GH5ZbH+LITSQHL3GpXBuYK0ziWNkwbMI
TW0pmTACWYdDzF3W7qsHi8raQgPw2I4VBC8IjWVQq79jPyaAPzTnmjMwHfDSBGyUE8YPBE5Gb2KV
YJIReNMSxcduqKHYhuQkHfb+BL4qa1v1q2O/FDX3kAKbgJ05yzgs+b/bQ7hG0fGKnSMRsSjn/FfP
rvSrfSS5tY8mBD0r/GP9SB81HJXEdZ6ht+McTlgGfhVTNIjcGzfIgVui3bd+2hg8Zx/C4PL8yvXO
NDeQadBxhS6E3PK/CkT35dJQC445uwS7U4xZwV52wnBDZcqWyWhyyrUWW9mQIHwYOT2JfdLyfNQP
do+mup/Tm8cVtf0HM5c9fF9GNtrIcmJHr/g88ALTa0n/HZdx6aRBJQq2SEbvDEVIzoTYNl0jOqYn
/fRLjLZlIDyKlnYr4drSo6P76xb5ACbL7aR0YBzUQEumxsVqCH/5eqewV8+gA9r8ODw61yWzdwib
tbP11Ye5+zlgbPXoxMvoHumDgqUicjkGhyfvFdsjzGMAgCUXmgeeMY+aAQN8LgNj+CyXJnnbUo5+
bWTNgzt7suxuuhK9+v+Rd0kvKlOpBuiVJbrN6XPVCYkTQ4GL6HXshgRHbYwjmEI7+GhvvQR2lFTJ
SdvmZTY84Co08tRO6A1gWu/FhO2CF229WZx5AloVwm94tgCMA6TF7Glbv+0gksqrSyOtR1g+VcjV
Y5XwU6dgd7Kze00HsC9Jynh3xFawy+2yxlA77ydOaUWElF2PqhIVTnI+GboxGiEYYQgL+SCR3VpY
u51w5H6TqNamT7v2biQkhpP7+T30V9yRkQs25oPRk7G3vFgJdYJAKFUvwHk2isq9in5BeqpX3Ucl
+R0JPsMX4O2z/+AyTYgxvwGZO0vGRydCap1RTre5j6AdleWe1KDdv7HUhTGK4WvyIeH2kTJ0+Sce
56S6cPiWg5O4+2iwKxqe0OiQ2He09iasAB1O3ycI9DD5RqME8eiQdicPH8Y3p6xZTSI1rluVN3dL
XIzgvJwOWBC8FEFfvWwnS3W/c56PXJvzOEbpbzn7OOMR/Uo/0G/EtLw+BvkY8loxSN2yzbTImVv2
io3wKAGucQqLH6xfu70Tq6+AhW9U/Cgl5vs50qJY9IucOiXwo33Akb6/0i5jjT14VEmuxZXWefSS
7C++uoz2Dnxn+lF2zeB7tFZJQ/LEdkEyUJaaVHbZzR9NEdVyZm6hO/nZWSbznmnKImnYuaN+qJBr
YA8GZIxo/gIuvzQnT12AMcOgRGU7FBOg+jdb5VSxdIp3JtEX+s0YcpHo3BggaSzhcqXB47owILtc
Ozc6YXX+i2nnXM+3WxSybkHPnNVMaug0MSsV0rmijOJenPQnDkUFl+RKq9aiuGKjc/423Tz5y7jD
+wCiZovnM2fL9l5J3Ubz1b8grdgoA+FN0C4SU8gRYusWVj7HN3eXdcJKves27rnv+boADI+M0T4c
roV+6zcaKTEGbxkfjg8TYP4h9Vpy6fYXnVCIPcibgKABqNzKZVXPggY8QrRKoU47JABN3eVWGyJI
/zEEa/Qf+wRJfydCEau/VfD8SgBEwjTAsYA41o5g7MJTTSRc9PqNEMQgBPVQOXML663JXbivG8AZ
o4SbEhK9IkU8F6ETG/F5HFaqKob0pTlfxcZst5alw/9I9ASzWTA30mCW5P+L0hvE4ubHcIuFuJsx
yH7ao6u3ZzMWmK6WwvtqYCK3BkGzkno6VD2Nbgm4JuwS12SINBzERnoy8YIkUVJbHwnjTnf83BNX
DG5IZKuesdd4qsPneTtpr1YtCnDTitIJPi+0iTYlhBw5oLaTXZ2xgxAwhkXM6/5HZRAL5BBThxHu
kH18gZ83nF7Hw4B/TGiRf2yJ/X/pRk9/9pl28QU4KN3KP85SpNAqO+oO3uUSLIOpK9XNYZXW6S5Q
cAgTDzzrdy2n5aVOxcJMonWVRVBHahLqs0vUpzjsd3XtgJAyx0EA19mWT1C5fRulZ5cfNyRnVlJS
4t2kQjF5F5T0JUvPt8TLB90mA4xmx3OJVjsRnABxNLFS+dAnDweQiabP5d/GyNwe00N8KTs4LbUM
B74KNr2vHZ0BMDeINmbhe+2PDPABYrO6/ghC3b5PjjsEtkqg2M8z3AbVb4c4Bwu/HKymduRY5nZu
revuW5WTIFF1YXA0C2ejpvOMoqHOPY6s4nGNapFaoQ0CteV5YESMglQljrLvnHCrAKm/jVyIo1iQ
BevY0Wj3xDyXizQFd+weBAB1k2+8aL9us8aflicER2htYZIDxz+o4NecC73F3bxvUhSTuigSeU40
G9PLzBoPv+SOtiiwlTanjqvKToGw8K6oPEoVq6/0sdPc1uEWHXYSROVvJor0193okJebSBVFo8H1
32AWZb7hqxTw8DN+PtbsqrJ6Ndv+pP2tP2hg1D/eW4fA57pK008G6YqDqUFNq9PfB31QSWwz1zs1
332/B3dYa9yKtvRYrSP1HXgoN+ciGj+pozMdpiNdwj7rDdH5TTIfI+2KVGjc6JOt1dCinkUBIbTT
yL0aLH/kRF8HVTDN91VlPdCut9g/Ltn+1ER1GgxfCGzuvoz9xwcvKlfsmHNCgi7vD++JTmF72aM+
mXqivPQ6XinclARZLIKV3JMWJzPfQAwhFJ7NigD58DHm/EHNHS11O/pj1cBRZT0W/CR/yEVaz288
hMjrEVRi49GGCwh7oc6SdG4wGWXTr2eKe2LzUXIGafV8xbalAXD/HmjypTDpSiGnf6W+D2xBJ4qQ
XkSFu6AjWuKk9ue2aAEjVDHDpBmkUBq/SeI5SbISioKl0Mf8nSrbvA+g0QAlQVNRgG36U0YEi0X4
WHeYUJv3ntlTXF2fZCIIR6ejum03/luF5fwaYEjVqHHlkJWwbTvzpvEnftLq/CfyEvmlyM5h58tw
O6fjrZrFHOzMZLALAI+1x1/Yr8c4LIuD0bYZ2Cv2OUxpoP6Xrf5hZEu+EXHpj8vMlcV6G/KDpcUg
trD+T8Wk3Ufn06FYe0mWGqdVCzjt0YR/ipr5dCX16xVTwyk/2q0YmX9pOGpXIwQPH7PlugoCx+5I
cdEgdDCnXskmc/ecyNw5rMIfPcGtR7eg6M74AQ2bTY5mgNFOK9ParGhYyZ8Wd0n4tKEOfHWBiCbB
oJq58EeqFXUuBtykgDfGBsvhi+PZ33fIyOkW0ngWaAx/aTOSqOhFWm/4qCtiKsU3VEhTQgxDUVp7
Sl9Yy+zM2weOGsWR7ec0vKSYtCKln1KSar/JYCq4ilwbV0c9iA8RGs8Pn6o+WiJDPq1+ho8CAFsW
TO7X6rUlrXrhjrXHpwg0vjEUYhe34ftQ7mZeVYoX01vAcJwGuXlz4iFwCl1F62hKDNM2PZ5VYtms
rWEkrmQroFyyu8SHoRxJrLeZon0CMnRSG3FclZFdsMBTQzE1lqD0QUg9QMteh53umZMeKEqDe3a5
/zD2EQUH/YNOVE9nSdt0S5UPGcfkG4aZMkNFa0B5oF4gCYZiZAV0dQSRkBcBZbtGNk8oh9bxQZsM
gLsD8w4T211C849x6Bf8/9ILC47AHadNZYMB6t9r8eOE0c+sLSSwrCu7DE+S0gxxeLgYhdBpxB7x
pcfe/J2FlDTsQ2owO2u/iYRJfq3gW+zsr5kype6siaIYpCkYCla1VcYikwPhbiMyMoEPL5/H1hkI
vbpQufxJKES8j35HOMEc0h2/OfMNccxdL9e1lDm+pOEX2VlDjGp/GjD2vNhy3SMlTTQcKEN75Wug
e/HB8WOYzzoME6Adag/oji7A240nVapg4U6lBm0drt/gHyS4pjAjyf+TJElDt2Jt9ZlmpX8rG/40
V+gjDxExKgKGFQDMYkElhGdeIjvpnPJuuxwNmOiSrkonlDbPfOCqOZnZV871l+yf9beQa/GKfRnX
RWsx8OBove2/W/WkgcW6stSTHUJiTVLdBfqmoJRtAR3csfbRHJcFhxSJYC8fddnGVBAPNuWE0Cay
RPycfPNbFy/PniIH9fS3MZ0YtJihI/RYUMQxNfAxiyHkZECbtdT7v8dQ4R/u3CEOAvabvyjq7Ouo
FnGfcqtmET1EiIsnFAh/5lsbpse4340/YIloZnYM+ygpvCT/4rMEP7aKU1nMHqESxjXQNYx674bC
r+TxK86m8cNeS15za8OBynXH4eMFgSJJ1OOhdD1Vjoy0Ub9AHzBnefkTvnSw/d0XERQNVEMZS/yf
vH1O+b0yzaNgm4r2cBQZW6Ot3R2Jbn8xa1Dow90OzGxo9VrK/d19BiL+EDzc83pgVUkzeVPpHRd7
AvsqCg6iwn8Keg7l2ueFKE43N2TKPtcJwULh+Rf962p9YA8jKXnW5xylb+7t6SoupdE7+ZbnZ3gz
oht51sffZzuAEwkana1OKVDLAtsbmxr6RENAvDGLYb8nkvkSsllW5yaK55uxiohGOtbqkCcVceKu
Qkmn8mW5uorECC1Rlrv0MpEMhQ9MdhsxOi2y2c+zAAPwS2ONX4lAg9xOIos0BeEZfiMqBYYmzRRK
INbzEMCg6yomGhd87VJwroNEJa75GJtKAVy08nRTdW07LGqYqLi/ZnAml/Y6ZiOjBBTg+/SU1pev
v3clTIA8m0CLS7nVGCCqCu5mx8UWpXWdN3SjCvj41RqORsqihvyFOW23j+pYVmg10RLNleOK4Fgr
81quu8/xEiw7aEcJOc5JHUic7r53OZEGrWz9YuhuctC/sCEkXVBgVW4Tul/4pXZSn2HVx5WHQT06
GC4yahtK5T7wPUpPNoqrQ6geaNgjrtD86VZIJolTjkY/SXuPQfBwLSN1LpWQz4rAWXImE/2Qmrei
QF84mxuPR2pwzGa6R/cL/gllQxES0TjdklK8+9Zu+MUY3+owajF9dzxsaLvYAUMP+SCnBOWCOWYa
eBRQ41DcP8iK8/8xZY5TDi31CL+CMSPFoPtXLzZd6TdzM6vhg9/PGxzlveqsfLPY875w6Pi+kpYG
wQe9kSTi30XQ0N4tOXy+dxtTjeVFR6PwE6fxL9XdtKTCZ/uvHP4mGNukOEH4hU5NG+Cc2EEnkzOi
YlqRrgGVzGFaTYFUJ6x/yQyVLb8kkhSrgAwLTScjv1/0Ld2NwpWrPMUtoT0L3fnNp9hu+pjTlph0
2qrndDCvzmQXi+4mhAgbhCZrtqmsrJzAEs1Nm63FtZjWacoJfSkvuZgmZFBl1pU7xFMR1jQEujSy
NRQjdrHzyijZjcXvEiPa7HO4jI8YxQytrKP2kNCH2nOOIdRmPWD3376t78FxzFExd5qkEz0LSB1f
62ndYbNXx+mjo+dSloshYAvyK2o7ErXsggVTmbJI0RQ7uJYdYMVGsHNPNxdLNhXNHuOHbJik/+eP
T1h9CpvSz5nk5eHVmtWcvqP3230hOfULfCYeNVV76yVqVbSHy5ezltUJIahroEsAYjBPcZsBinRX
CuPCy7gDvqTo57sVovEUvjPL/XGufhVCv9rhqx9fhNFXgrDrNdxLmPzjpQ5fTFveW8N9lsqiWQ7h
DIBZlhN2m735g/j5dJviEz8NfY3Ym3OFiEGDqP3S3R4v/gY+UnIXDwAuoywLfpOT8BUVFQnq9ups
5AwrTdpODRZsnNutnHja4lgu8qI4a5j3grOQwzI0gKrwkTJAn6RLa+LVwft21hgcjxuAQ4Ez8GYA
JAVsWmCJ+RQyDLkZRrbu9J0g5J/DuSeVz3I+IwMMbOptc/MIukEsKjdZdu7C/GHw8l38I/ZYCjHZ
gPtZejg/mlTCS8CKXOWQ3FAOKPNS7PUrrFwRujikM7pM+LjeYACL0QDPgMLpp/BBig5GNFD5kuhG
wRAW/IkYMZiPUXg20jfsw9kD2Wkdy1ItatMTyhU783rNlkv9q6bdPbZT0sECEfe8Ie777ATISEAU
6EZWP7827pZNq+ZFTQgng2sJi/BwXHng8gNR14yXCKPHYDqGNjZsulDuNDNO2C9P7Y/ASld0DSX8
TRDZB3BP84kgiCtRqXZPvzGQPEbYpRrxW2yZTIbxTdeMzWaUsfvGdzhz6UApjIf2Q+FDqfWsoJxZ
mnV6rGxNSRaf3ePiEAi+Nej49GwsTY1hSfURHNt/akA6+2/EXuwrkqFzFMyLnn3Ur0u7V0b2SZy4
GIZLpOL5ml+XMZkTXfqXkK1QnwzvlhF6u5FgV5cEFQMHBG4uQvfH3QTF8bUlMhjLah7FWLpzOPxN
uNTW9e2ZZDZCA7JpbXzEUANvANvlamIMsxQLyMiiyARslwD4Ob2QZ6IEBIlVaehnooMoAO+oeQpl
sum+Ds2h1NW5c8T3kQf7VxFCkvZwvhNDk58HF91U9NSCdLO+Tr728RoovlF9t9rgs0NkeQpgfcN7
VdICnL9pwDT5DO4AjK91U5lxjLFI1BBklpZzggzKV6DyU8ddvU7h4X1NzA7/Co7ooX/TzAjZueoR
xC8PZ+RzMMXgwDoN2EgTjDrcTMmAutTzVYMm6NcAoiG6Wj+TufCnXAHcfuPgZwWWgstCdESjaQGy
lmqHkRB9UZERTa63DnzUZ4RSL+otRBXqAKbyaYPqBCx/vpUmw6zekVQjiVUc9ti/8JrS85Bnp49K
K4fVL0G6QAcdx4dL4u+gXFi2BQBMdJjp8NGMwPAODFaMzmNVUik19yMnnDmuf0DXOzXG0UyPjn+7
Yn4rCKqxfOuFpadsYQ7tUvmFgZkmRqnNhThgWelo6GyaGPhJHurXpmKC0hfgzp1zg5AZePN6WLnz
xgcAXjzV7bv01LDaj2AmTfpjK7Mo8i15+pT20J0MGSshtLonIRuvMRM/EtoOfHmAmG2K6ZaFF9pA
Sj2bkLOepqwyDCg6oTWuwUC0mD11e0shegALtYUjSkHpI6FNilJxSUfKyMBZqG9B4X9JZCJiJEQw
vES0ZxX6c4uSBIhFOvbvms1lnshp5iscw60XqXRE5PzznzxDEDgy5Nwp5/7cFzMVhtBrkS0XG6nt
lHWX5yD27KOVBTcTCy1E9/jzL3hxn2SEtTY01WUz8Ybbif3qsIDXnJ3GjEukUGm1TG5qPlIB8WgK
v0jqfda3RUmmAt98oWFP6joJps23VAvsB0VkjGc9jSqjXHP69s15qQUxgapoQ3xKmlQFfnNdOTbr
VEWhL1fMtiDDEm5i9alHhrj6Li0xYJJSSqhVMpV8zcSW7/a1Mv/i3X6GoDjUu7ucqkeAGHzrDow4
hldMLp1/56Xj5mtr00LwpuNEwx1GdvRHziPK3+pR8vX/81bRvxvTgF+TfkzsV1ysC9gZ3/XWGr3q
4yyJbYJAMSQykc8E59k/G7zsFyYZbxCbMKoZiP9YfULDaqIZivgOw7eZejoj3jqCpdB5g/YhCuyO
kWtn8XKYGN0UP1edvGGyYcNkRwg69sZo4b+KsVsaU4reqMKzzIDubFyJt40wavuGutpscrd2MxwY
Cxusk4PfJyEMs6UcQet3NRDZMgQAGBmie1uhS47LCWikfAG9py1yZldpygCV9csezjcl6pcoRgWn
QO6aAUrHiV+nK9iVfX5eeZKYei51buZf4f8JHR8na04gbNi/CSXSHhII3C4USRLkEPQeWbHYpi2s
MT44pGkJH/z5W/1gTW0O4gm8ZtDZY31xyviHVauQBQ6LFso8T0x8tHiZArqI59/pdY6KXCOsY3T1
c1FDG5bRmqd1NaCGYNFtZ6I+/QsTSM7hdwqUpiZF5EdXMDUnIZ6DBUh4y85PfideaZsuXRsH0Qty
Q5Vi9sf4Fr+fX9OzJZXaMOstmmLsedIY4E+jLHoqzQy5sOq4y4ODw2ZPWn2+Vuxe2wF3US3hRaEZ
ujsfpvdTC09/RkXOOX0uepsrVdNafFknW8j+zVMRSTsOKMsv9+PZJvOYc1GexSuGMm/M5uqiIeFN
wweOHXV3wfkgoZfkTgvgaFiRxZSMxCGqoQfxwPSzwp/pau/tS/7uGVLPel3CjQKSkMDKrHlZtywA
yrRWURy7pkUko7Fa4QozwfIvmJlH1FXt2cyuiJz9D//XKDWj34+89O1frg1jUghSxM3InGmAq9hS
XAZRbeIx7DpfFb6cjI5w+o1xpiCXjpQW4V8/oNTUKgJyyokZXQBMYrq5TsQqjvSB269q/KwprgKT
3XuIw3WPxN4NWUyNIHwrdIA0m03e9mX/JWaMilUh7hk/rzdXweghYWrfx8hebFMVOb1wrHg1wcoA
cj5r7Za9Zk/aF8TBS51IIiUEzQPMtrS2nSdboJ74SjNSeA0XCMeKlntDQKdjz6vQ1yKzEbU+gGki
uMzK78fWd0J073OksKDCbB0zWlCyf4LCP0eRRUejq5VR0K/o9MeDLsZixGFfFn2+YQdx4q9gYaeq
vrSmjwiW89Kw2ul7Ewv5LfhFmBa54nU9xWSUfR7XrafPI53h3T6n+K3QdPLLs425oK1hzBzaj1Sc
WSP64dwSYKhlza3Zz6DMN+WrFGMq0dYzaOU11UX4PSUIGMMtnfbq08FNRZuf+dYk3f5vuK3POl/3
3LpXl5TA6/onXphj/IvN3lM40MQ3LtPCUsA3fH4vHhsTHCmaJ7tqyz4Ye9aCI0AvM1oE4V+QEYLq
Q+7K20TZvOOZjKuLEh63H8Jd06on+jeCeIFHpYpsIYf2S/tgWTc+l1jbG5++2cjVIE/RaXBiirOu
g0DAFyuGhO3gmTzDaD/O37zPs6Gk/lbkaREQfoVJnnnThtDzKJLrTFK/owm+N74iRvzGj+cKb++H
xX/Ic0Xeh/iwR6OSRmrv+NxXS8ex0dkzW/zu4fraufM/XvAlL8KySXiL/RAriSK+S4d8iibXU9cP
fgPOcPubUf3AoQ9Q6YCZVveESVHaQILq/3cc0mexJqeNqEoX3wRpBLLw+FYdhQQwK/e9l1y7SvZD
tcsfmI54MGlPHudypU9t+cFSKwJ4lnF0yu92D9sneGYHuHwyHPgsM2lSiiFgC1Lm97zM9tUEe/um
n+zyj+QIw6zZSBanYlvegA6WSSHnrlOK994kU+0qRCcGQi83aNRrhkze1XyLk1M8nQh+OtoA3zjO
RyvxC+IcozKbiE2VTkpzeu9DXwMKnLG1RCj+DYrr4lnucNddIGS3sDNVaHrdH8IwVLoaxA0EhFTd
B+r/FTG9H+a0hTbyzuha0ZnxxvBEhsjW4fn8CnL/NxH+bb6/htI2Rp/jTbfjCq7uaoWoCm8y1m0C
41/OQV7Rc6BRTUAHIENz4uh8XiQJ2ZuuGjWrecU1aI7VxFhclCh2mAxV81GlAQPW9InSI8ktj9ld
YzRHROP5AN2TQfApJrqWRIrFIu4FfNlNE205VGWDka/JXhtA5jwoNJ8Cg6IB77xHPGY46dP717pn
yB8B5pFLoFpwcTKVX2A0Nq45EZvbpFlIFrojeTBMOB18Jl73vsM4VuhAifFEneTig/tGlbmCCy+i
lyZpNzdM/5luZsq/BqsTaNsnoC06ytc2/8XhzMdcsbpYp8oybClhbdT+LwZKaZfSXRqh14RI4Etj
soPOuglydIqVljLy5bUieBHEbcpUlCePmoukyxVKIGTwupNa1BbKCum7siKULtr9/cJ6JNcqxPS0
cmi6yx4xC9/F7eF28Tawc97t24BteJsKl7BWrpebQB47YdEINMFdYTvFH/ia5awutd+pt6mbqkoa
aqnkfuac5Am/p/b2aN0Gcv1BukaNsY1hVaXP//0nZjB7Xb7kCfpplu0NeWDJwC0kFKBjoAT12D16
h24czRFsyN9AQCNQZARRr2poSY+lb2qUCjW5c2muoePz5JfXEfFw+V95+nchSS38rNzqH8uB/KiI
cIf7R+EawxPdwpLnJLAw5yf1fmY5iIX9E0mOurAXarR56rYKVUQpPvfjGt9bQJgjo69ciD1A45DG
sJ+5amjmCoHGCQvGWkzTEshe5tGLcGzbX/cLm6b6jaAMLKDH5I3tdtvqC7fYb13siu3eree7yaH2
K9h4TFJSJsBhs4zEsJTq5UG5pYZ2gwXZFFC3dSZJ57HLC0aU9f1e1Tj8rXxD4lSb9FBV5Vg2oTtL
2Kd4jRVN2GJdI4tJajU6Rr6cUKI11H+gGDYKJFc6RioyAgVKfbb1no3Vl8YP85MeD/Uu3jlNTsno
fwrq59jwCimzGGvQYjsLrkuy/gzYwYiOUf9h10QpygXF8vrxdbb2o5Za44E7EsSYwLaoHCQSb23r
S6LgdC4OIder40J/1nEl78b2WW4fDnf1E1u+NBmWHRs87IHnp7C0tWvbYZhpRls+IiUVVeE+NePB
d6R0I29lrnP0tzS/iDVgkjPvmS8U6r/on6hp8mql0bO0toM9MhVZ2nj8AmkxxarL/DNqVLQt1T4i
XVNYOzuQVni+AVOUS4OYJ/dZUarYF06hnyv3jwzoWNriX5M4G0ALNEyHBvWcrCU7NFIJiYBOh7zF
qGAjx64c6jYnQ6xOYYjfmkOJETvh2m/Z0LJ8j9pStZz1sGnIwlNOaF9P4OD+tDnDSz02cXrKfznJ
w36TEd67QPx8nkJ28CV+UeKI24phk2SLaqDvwKo5XPIqPJHfTESxu2+eX4W5WMLp1KEJlADdFy/z
0AM9Me/XjiweBL8b8KRfTL3TIC8Ntf4HR9D79PvBCe06zgErjn+/pQeigBgt0K2qNpDkpJ856ZiL
wwFu4Qo2OZvFVJKf1fxgTs3d5JX3b4CdMuLnaX/FpL37XaMs4Jnbi+hf+f6FAlZGXGblxMgOlgG0
Gl/ImfY7cO1+NvpfuhLKaU/HqDZhVhGkwmzfxvmXFaPtHL3xZbnoyPR6jMpWUzivcRZ09+UnGzMc
F4sfE03gcb3e9lPo1fHCPA0dQqoNRzvwtkjwcrTNMFxCCEwiVDZImRvaqunR4/TgCA6ceJ/pUfHJ
eF500+PHppli58hEQHJzOy3y/hIDNEIhlTDpuBMbBu9RSUXT2yGAmmSLD0UHEtTbC7Q9brXVNCR+
QhofMEIBx7H4SFfzJ7bGtNGe40NH9Av2gUEmr75O0fYPuepYIh9cGnNUbNFgrG23TJxZLnFKNmM0
RFM5MYUWsV4yslxg7uV8UQhGMEr8bkciILEcm1MmX73gJ2dp16x15uNAxOb3e/sWXYiV6i+gRmuN
yjYdmp03vmzb8rSQirSo2KGjVUdYNZQ3AlbOD9bgkCzr72vCN626N88c3nDLB5NR9OnyIJlOTA3Q
hKUM71BRXCSdZFkbsNQBSBLopK211r8fFCinnFClMeIoBcQ6++WB+30oCEkjEhvNinSBD5eAvjF0
FYieC3fXhaI/DDPK4gGj/AR4TZi1ksIaM+5JDtSoyZcM96A+/XPph75DpmyI1WDPMCkxeUVxh5MM
80UUpvoS9NiQuBZwXjD8Hz9CvEzltQqSYXRey6v4Tck/9Tyngf8y82rMi82QD8G8pXPFgZbcTJmF
s0elApWiFerfIhcqp89od/FEoeVlH8bqFDoccyoWU+pVaIUTg7tfsNAetfCa6fE21C69IhhxUB2l
Aq5MKrHB1BGFQY8zJwlYH7F9gpVWgUpmZbXMNJEEddFvjAKeJMYq+h2gFfjnSfXKpyDIQMk8rPpo
8ZQm/x0jGrgoeQFzZjQpaLQDAE1v00JqZmiFLDhKtxT5Dxyy5gWN0YTN6IM8P3OrOnEZNBe/7iel
p1i/yE8xjFMBqUFXrX6yb0PIgOdwvNspfLi+N194RaI7diglabTPR3/3gbptqgcNlLWW6RqGtq4C
ruZHDGP/KIi3Xlj+Q/UE6W3BmMSS63b+nd/tfcb7QU23kUxDFEXGNmyjIrwPaQ8nulaHbuCEzmjB
001M25pV1HOgtH61Oqsriy4bVx+lYWIkU4ET4fEpn4+2v2an1t0Jo+h9JVwzGeoefJ7ni9kHBsl0
A+QmQKV8pIe/f0H69OqvWKv20cxSU8JM9V8LptU85tF3g8/eymx0LFySL0KRH+8HmC4OCX2hU4wL
q6aC56kyxo4qJqRG5IzlGfJLK1sb0O5V5hddTcceW2AmJ14EUF3AtoZIrV42FUP/JxVnvNScX/su
XRt2besu2ZTjPql+h5FmFZTnu/Yflhxs/TdWG8gTfLC0OqbT9wHw19zM5XOA5JuklTBLn9th0QJ8
NFIaUKub4Lh/SUoaF4vVJgKa6SSY87OD9Q7rysgzVhNg3ItuXH5GHu5H/HZUsPGWkiebcPAKq88J
Y0GOE3nfwzAyItDrKQvWJ6pjfgSphIMjB1Jf/D5W5I5t5Dy94kxcOUKD7E665Qh0j6LRcn+bgUyR
4+/C2iDJlrWOj6q4eogQ9w7DGvbPvHIgSamaBPCvvXZN7voS3beeZZso04diyuU/grsb+fVcqPQi
JZuTd5d6DTBtkiWZjVd/ZMIAa8Q5tjWGu4SsgIWw+GJ1t7gzZL1wAOK6weFa6MV52rqs8XjwaSTy
QPKLyPE2MhOAsEeyUKGZ4BcwzKFLu/PdtV/dmUjAJyzmlpTsdhC7KF++BYtqhHg13Ahm/3Hj4pBQ
SKRlVz05GGb7MTbNCGgz8PyhciL23FrwMafYFT4SWX4203/b2kS05R7uVSphOKkhqaGwOJSHeQIF
YzzT/AOqlpTtq0uJnrCFMSfG2hinV/rQ7q6SWdBH1ey//SgjDKGJyPuKB9w9RBBTdHsKNyyQK1c0
GX4zZW/sSiTS9hrHM/Tj0YdMO5++3qZR7V8mEtmWfVu2xIpZn6qejC4GwSCfXPMM8NlQTiBOuYrL
XH6mnAMrJ3wKII/yNe2z49C962KUXoV8KWUQ/Y8X7t1SLYJo2zfAlpoQFuWrHHlqJGYugFoneY9S
dQj9IoEB0iAHVnCefZEhBcXBS2j3RjsAWr9R49tIMrvthY0WYpOE8kFp0ctLTGs0VS23gMZw8D1R
f+lAwrC1FA8xTpe1blROvjgFXCxzNhQZZul6AWCRzoi9WESUL5Ek14EtmIKj7PZV7q2cUQgCSsW7
SbrgRKIFz3WRbTdDR0cZUNaDiNEhMoXDvsT837gQ3qI6/H9kLcUbG2cqAdSA3XiYvhpuRy6doywN
umV9u/j/GOGaO9AtZPRR1D4OdyBtlbhdhs9RW/ItbJTNnKCAw5oNk3slhfqQ54rfo9hIRLt6EDxo
wfFEHctKGbRHHVVzi4ksFgi/GkQKBgjQ2pdIZust0+nk5Fxr4UZOpSZ1JqOWUM0rzmT/ybKvhfgI
4ahZYAxNnWTdbRBX2IiEhBZZUFV6bYQXg4+68f9bCGU9WibrRwCg/XRXfINm4ibQSjf3C+ITbXQv
jXy9sPvtHAvensskLx7X3ktEdoswQDTLA/R4R4c+CpZbqeU+Hrh4tb4vUSJwVmYD1gntXryHTeyr
g/VnboJaf6svoZuVMmXdm+u8RyRrh4r9u90hW/NZsb2qsn4RDwNbI6SCQeRC9fHigDwQ/kHd0Phe
aZCs1Em8X4caIAk2Q5zkwtxAp6Rr1Il8VEX1pTsy9fR+cRsupGWR4WrE3imXnJmaEqNmowX3SPHe
DOwMt1DNb2/fodF6ryJoyhdWtCtUpK/CxfURd3HO5SscRn9cGmAGBoj3O5W1vA34Ac6cRK+tKG+R
AIgGc1iYuzApyYCzmrb+ao3exmMMS/m6uLMPircYsZBuY79Z+iB1+Y/3YMB+6+deR36CqR4uPA9G
DpHE+EI0j5bP/IgcXLd2vMxrdbDFyw3ROYfE9/gZ7VRVBRxFtWNgv+fgc+khdwFhtEqBcQjscvyb
K+vN0qiybUkmIgMJN0owjVMSxwzK4/It5OW+HrvfzCtCx7bQJCVnEmA1x2RWzqfog3/JJdy43QN8
xX8kpUeV1q6sLHmtwTJMzoJUoXiN2K88joFHFw/AgutJd+rI1UNcZGWZ9LbxvKmApT5bzT51Id9A
KscL0BW0muqRcWiXuHaMkoTIQZx5u/lqO5kT5i225MkTdo4rdGRwJzeNYZHogn6pyyjSN/FuZeSQ
je+pQ5iZYM4F+WEO7O+8c58e/nTxao32tE+U/TDPZzqvxzLnaipJWUL+OlSIEC/1nUI3OtpHKfWw
DdQyN5RvhW/pSeYrPxBycRPqU/bocLfUtrVeX77a/J/IElIATyYDF26np5rPh8/pmjzoUq/AH/O8
qM0KOv9FeXyLv5vk6rcAEJfoJzIQscPW0geL0R8bYTKyLL50ONohdlvr1Obx1u/LXcEM5d2cE3TC
ATW6BZQHDHwv1/4zMLm9+VStp+pqc47B8bh0oTBsqXpaZzyJNtPfW/WB1F6EoJaCGByv3gGo5ixj
120SzOE3jncfmxXa40yaLint6bRaIRhqAdTU0t29yR8aI3X9sgbjeW7pseydnBoKBME690uAd3Sp
N/I5N3r2ko5L1GJYvQ1+VuwjdIrI+tZLQZ/WPYmQlhfqP9obziuBYkltBWRoTzYGv/03kIRY9FvA
IOGNuleh5Uo+NEsl/dMO28G+K/Asd5GtLFLBZ63oC5A4W6hTvbFT9Vpqs1BHiiR6CIjSuQxIFITu
jL3ARuirqCmN40xrZdurxcPiHDLwYiKvHuLR5kNd1eVP+reQkqwo+4Q8vwRwv8M7kRYQ1bzlNSqg
Brls8LU6rHmZGVd/l1lUkKHVkiHJCnwZLMYeKffaa3Dgy360XFgIAwiYa8RuoKKnbto6NGYhVNlF
E+0ryrEP/Ykhv95J+//9Aviftj/pWiIb9jmKbhpHZsytX/YMftgyAmO6l86hu4wiP5ksPGUZT4jo
5M3ZaWh6XkWtKcXSbF/iTp3DQtGNN4yZ5ENk0AeN+lzYWkCkkGO2eFviRvTSiYaPrscxH3v6TDm3
730x9rplMEjsQQZSbyp+EVDkJWsbFBZMw52FgvpR2yB36DcU3rXRLJtPIo583nMsGZnoLPXTDFBn
0WPfc6L0yxDwKQV2MskHqkoYG59gB2K09xXPPzwLn28Xub04cuqVseLZktgMjxo5WWRcZNbuMIuS
C5sxoY/kmyVaLKUWq5bBp0bm1o2eezKYrX0SFi7P4YWKbcjXNYLhA8eJdcTjRkf9c55AMCrON9nq
+sNICbBQI1fZUpDT2US9UfCzxfECrU/B9UfZsx7u0jJH41avJ04qBc+w/zxDxR96ffDKgiS1ujaU
JLxUhdPPjaBIge4iBdxRhHUFyY3xtOLDa4aAPmR7YyGZ1dBU5O7w7znVLwOx0pz2l+PE6CwsdYBE
AVEZBQIVPfbG9XYCTxysCJ3Ax1ZuNC+RQhM9rq0GDDKPliveFmmIh9c2cuqdq+D4FmVBvpILCnNk
2G5wnNJ85rcLdMiKljHDeErI9wajg/ptGlWQA+g8PreMEFE3SL3okUWwmdYHPTrpN8MsRwTa54Hy
Bsq3vehj8f1cJx3o6JWEoaqhYx1yioaRurjER/1P9v/AfySzdnXI9kxVulXk/nQkAF2IITjr+QDP
+GLwPOJ5pcvYlPd/Vi7Lh/GPT+DQBWp73wIq9IQhKmGMGjdiXxvt4xHmcrMKn00qH3QCzqXo+6X7
pbn5BCN3i4bCiRytjzvpJa5tF4dgSnluMmNjr6Qmu9bcii7TcksCKkHi4TpKl/RzOmQHQsVgmB8R
jicvOpe8dPZECTKRH+aTWSSQw+Zy7+apdXT5iMeRvtgN5YUlQKVv03LJQFFsAmnli0Ak+jmlGcQu
ZbKNwb5H/rwOrUIBOvK+Fo9rpUA3P8zhxzrF5HE3lV5DLowHqz0NsKst/pSvnSNh2gYOCFUIbusI
L/TcEm8VPDUhj4us2Swc04ySk/Iz5aACD0JKs/nCv5mXb9WW3hxqCGf/hcn/tKWIfoM3vR1wycl5
VNUXpq4X2LlScoMBVgqJb2Nk8zacO92BkP/mwxVl4pDoB57LxzWx9bl15Nvx9Tzg8a1YuB6MLfzZ
5qV2+zsbFUEEnTucu0hlEoDx2lioO3U/geKQ/6pH3p0stom/ERenUzLnbxf8tB7/Wism7XmAnN5O
pV5JAWeUq5aXa1051zZXPWDB+uL/o/NRTNZup99BNZj62ZOrbUazVKZs1WnJdzdigxOWp3TtRbMG
jtYD3K99aFnr1lh1i9YQMfZAQ+NDaaeldQBWcS9y4ou7uO7fYt9X9abdMqzXjVGuFDx9h56blf0e
CjTDz86lkVEqHwZBA0SxEq11aeR5SacpDgununIeSRqNSwNMe+66WfK6Iz7w9KR/pB+gA4wVQvoQ
LFZIzE10t64UCnCgWEnY4QhObf0Aa4ARY11ZIv2TV0ReR359G5p7xTRjQlV6wTurIlF6Zt92lHps
216HF5UPJi76oaXYhRTX2sJHEOR9v8QKY1mjBpErsJkWjZq81wVmm0I1higiRVCH5qjGd/9F2pox
ZpO+J5B41CVbwzpja0kBe+wYyaJHRDZyZUWLNYll3agPUvux+iiQe6aSo3BXX3H8mhMwfA3jBQm/
Nu7gUZccrS+jO3kqZ6YMoQiNy9hAcvT0DX9uIrWaWocuXSVbY1ifup+ZK/p5OoXgvJaUH0psfYCQ
uTt2Bc/0jj561ybxmvANcjNf5Ujk7Hb/C2v9K6fI4mGwg18YJjZGv0ohuAJIbRO3/OQ6hDTXjCWQ
Xb55yl7e4tc9n3kkAzl2dXMJdOBDTy0EOWciZJ+t4icIYAKQj1eahxDH/5+23vfN5TauxzuEL63A
YSjGbYSjhjDRkpbYZtcjRkLnxWrSzHrVkDg7XZnubK7XB9E2ckhf+8WYwQg/Gkm8Gojl7uqkiS/H
zLMv6oazSHqs/aqRLiyNMX5r0j0XEq5EArUjkWtPm44kY5RtxrQW/rf/ml6rQh/Dh2clA9hf0D8f
pD2MH0h8408ezV1ysmsdN0+oozBXWUVhITnm0K56xOAK89F9WVhLyZdLrSn4DCoLJ34BEX8kr4iC
5Upe+hsQOIapeAzIuzo5w1KANijxn1a+MLh+XyMY0RnibdYLW7U9flLdtGjgeYDi4GaBE33PjcUn
FEzdx4Ipw3SVW0ndK0h8dwaHUR+ntvyAlVW5RWuUgh1t3VjasiMlni2PXfkZ28njDtSXNRct+uSY
Yq0hnckQxS4vW4GtJhh5nrB/KsNkgMmzq3QmMg2uJ2qUtt3UqEd5Tpqs+GKK0J1b8A/YcGtEjwae
I6M6795WDvEmB0uWDINfSQqRWHI5QiEPe1buKntw8Vl3Oa1RgFauXIo2UMyJGvsvAtlB+I7OwpMg
P/1UI5QDfeRi8y+Hp3DQBFUGTZOMVxlEywg3/XXcm4xjB7Z+IJQwTcepKy95iUNu9hd3TeeYD9zD
xqLHH2OVzT0ze5SczT/YZhZe96+FmkqHfbpjhM5bdu9bo/Ppe4lXOIjHek7+AQO8G9Clmx0ybd3p
X52H9Q5K/4IMnRfBrwFzpGmtMTrwL+dW5VjQxZfBWEg2MuQbhTh4fVfr2oGkuq9KVByk1S3EX+Dl
/SNeUkoQYVfSSoGDGsd1REHBEBjeJ0t4hstv77rt/j7Zwuh7DUyZ7GzQ0JWOTJ6Eb9Lb41QFDYyM
OKsCa1MbHSotgbqEkYw/srWmFbhg5TJ/EkIbIlK2ulj6cti32v4ItZt528gUDw42DIdeQvDBsRz1
bpF2wq1FrZbXICNlBsa0+Sa3tM5isJeJbSE/+d8uXNnxgvGExZosL9Lb/HTb6UpDGRiuCCAos8PR
SnVWNZWuHN8BlntspQrxZRUyrFzD+4oXmjPir2xZpMvSUwu2iq/MpfdMwj3bB50jaUmHYMwlOKVm
aS5AELXtkI7WXd+4o4cD6UVi839qVmfOGf7v71c4E68PK7HQTTvzAsonBvtI61ZsZK8+s0LlMZlT
ILOP6cQzsIOR9I2bOZzMiR6Ie4MwyWNLhBzPb1pGK14AcNd++50FWg0bvPrVJT/vw2pVytAyeM0f
Tsa8QGoj0Z6STGcZSTkfmOgDfsS4IlqNq/gp4x/Kkw2mmDhSpVurJvy/2ZTWRDf1xfdEFUzpzPWX
jCMRp/0Ua5oyuULhlW85eWxGf1+4/F6SCJW2579i0jzNNONlHjo02ZmfYqVzz2LL0DfXXIpiLDLI
X+bT4s7gPdhVbnWc6W9pxoQt5gIrxQBUi5Wawe48wEykI74jyoskNHdo1CEcJ7LU7GNze7TdQazo
wxfTAbW8TbCLF1+87MQqGfUOkxmiyOwKnWWwR+x05Rs0Rly+fXfJRUQBNr25QXg7nft0XQDe0t8O
OAy07mPj/i4F3ddHPWsoj2mMjWgm1xDOSmEeosLS3Nk1uHf2+tvn+qHR/eSjMC2l1Ua12D2Ti3Tb
ANvEVB/AGcgPc5gIQewETnTXupCotCu0GqHSqg5br5x88R1j+x7u2v0CPNHKLs0YyeNxvI0PLe9g
3qP2h5OENE6Rf9TZ0rnnNn31USSRMytAuTAoujYOudzKwDZTTElHI2u7hYvN03NPWHv3cq7Ak5Xf
1s819UTaPTXOpOw07TX0LKJpoWTcGXW9sfRBGhSWtqIn2IgY42aqHCuggs9LYPvBSUMJ3egFXuib
se30+YaBft50M+p0xlqlo83xL8KI4Shdmk65X2sIxgsTOSfnICV9TC4DY6pyINQyRiSHZeBTYHpY
hy27Em0HsOoiVmwNeMQ8i6Og3x/7PexiXeVvgoqKfSsff7TigBV7ZxqvtYN43Of0wCC/N+rMgKiI
IJrUTd/dx6lih8dUpOQILB+h0vx8CPOz4NW2t+VyvNC+99ahzrRQB7T29rvB0DeKP8OW+JoINucJ
Nnj4swGxTY7g0rIykYJOelrU9J6BxJm/AFitWmMGjPXY+zzRgclS0G3XDNS6y9YMznFPl6LNae/0
LGhPw+oluJ1DRcYVOarHJ3u0t6znniAC7lvUmbEbz3hpHtGz+bK/nD8+Hd3VQKs7+b2ShUwJwaDs
Cenbf3geRD/c8kFMReGY5R9cmAckUQIlnZBFXvRr5apsVMle9yzm38WN73jBwhNlsk3vHBQ7mX6N
/o1i1OmXfvk3uJ1dY4NIOJ8tGicB78GMHIU7KCGrnPrOLPH4ugnCnwuEKuTV2YM9YwRQ5VC/oJql
OmqxLLSZ6e3TIcQQukdQXQNmsCsDMryEZeWSY9n/Q9mMk3vhdmoyh646XI1Z/raNPMJO+oYxEruu
aqJjR82/mavAx6bBTtMSFkfWQUTvZ2ruRP9fWMrljYy/h1SBUTBd68GfkpVwByepBmwMdIp7NUXZ
ksdlPjoV4BSXFb+7UnwUxwNqoz0EkXK1zNF08X2OPB9A3Aeq8N15dKiiO9TIU0WmlGsdVMh6dFN9
SyzuX+UHA7fmThaV97whvNLCIzG+mJu+cv72ABiJxyZDDKuoTlwuklJTrLESqmruEYpg7BJdosAz
wYaRJpYjGp+lElucHNhVNekWC/b5VdBCeILUAlefj/e2FFzEdGhzHLZn2cA8UrxHZ/pJmk7JTMAb
LyMQVsqvyPiP8cu8wCPGn64TzwUxEvB05dFqllff99aqaHigzsQUX00BqYvUKxHt22zmHvEjE70E
V4t91jtlnXisyqT52ECjpFQq2Y9uPkVLxzcmMZ/gAzfyurFqnKrlcHUX6IHOwPDhWA2R5yrsIJQM
Dk63ZhRc1e7X56fJzi/v6s71PnFNwzAFgrDZlh4Q9NumcWHQRblS4WrVLPLxxAM0jo0Fr8PyuS55
NvfOy8swvTQrSITFXm27OFzPH3oD0ll+qVzmL0qs0F21QJpAknl/Hnk1s0eS3W1zIFkNwbtBB7CE
MsZ2kpNa/8AF0xN/CZa6m5EKlNcgQJ7aWDWfTIEWxEvzQrPC+lgDAgs+ZZftCvB6bxQCNytkJrOq
d9cWty34Ye7FbdbztTxaNx6E6PRTHyNftLWaUrwTqiVc5HtT0esq5L//ZE52pr4+NxKwUCdN85lj
LFuSw+PpNOPf2VEFNQoJnsD3LpWg4munYV3/qSJ7yyb+441YlzUywrc5CXsvIwrS/KCLEHhJ2L7W
RYc0sxge0rpVukyjTMt3HD3hTq+YZ4DR0DvINjergs1FQTYAfn+5A6m74tPNmfIRmQLd5nB236dH
M3LiiBrMBa2Vm0eU7uL5Rzpm5xV4MW14Kq56UZgVRHJumiujM6C9lM0eaekBQ0Ag8gUc4K7iWD+v
EWg2MD3lXpxLa427R/Vjw+hPdmwwcU5SpCoiAUPtmm22UIRNcQCnnW/65CrLuZlpTsN/HQMboadu
pWOse6Gvv+rhuSLHHVOb8gooBkvDKFptlUQ0VZNg/1p7zk/hYlkY7WSW5i7zOQqiOoZTS4NgzIFO
FZgfHqu3cXnKdalozPY3aSLFEJxW38lHG4CcSMg5YD4lMYYaDbEJmOX6KQ9K8tsYcKkXUPsE6KuY
UsLXt+7O75yWMbSdef4sp57uH8adX/ZpgbgKAYjw4JCZyJjKZl11LTKGK34GDGjir9eEh2JoCjb2
GFq0bd1tzhhc5AIzZLZUswe+WEfiqIHgQEbwUdHNTBuecbRvHDBssxY/3/8iZD65bsTiVQtfx+nY
V7a+J0jMhg1n3ne+tflbtqaNThNRL1pMloBn5BjfXFcLO3FRwWdUuil0rI6f0F3uIoU+Tvjk8A4D
64UFGzQYXvvMJUVs5RaMSSpcsUmpk18eI8NuWjm5deShlAqjXYYFEl8RwzSHZnpcCQ37VsxJajFp
uGYSh35iUrUt0k4wc2N+geXysh7BP3P8A8bgpLnoYCTV/J2M+WPpIciHzkbKvC3nsximPs/hkmpA
B/hujavGAyEvogGBgKIpRJLSeRvIhZ9nuHOqMkCO/5+lBndNyN4OXGc/I5r1GgVO+WzIxMr8zaCc
fg3ap9pXtO5XqyIXcawONgO1kRWzN2fCksDsWYH6TbN7ok+Y9neXxm1jaoJ7WRujHqdqkcx30b+G
CyMKLPVSjia8qpxbfdCMJAu1hnIhx4HrwN5ksbGrMqgPvIG+FdQqdnkz1yFfE7nGnNNjSWItPeGV
hX4YOarX3U8KsAE2c47FvU8XWCq7JTx7R9QsMTFNk6Dp4gUt9VmWTAa4uD5/pWaqqEu4C8PevfS0
huPRSUZpbCThLPvd3XPg+cmEsW2x/D1xQl894AVj76OzVa3RhuRp+JCFDhAVWnCpT5L7+knygX8G
G26n7vvYBEzrZed23er/bNa/jadXSrrJx5zMWy/iCVNHLyEPBgnRsvzO9hTITD15IK4+gnFViTzZ
VXE7/zRkyiTDUuGhOtfWPRf1abcFCr/saq159LeIvrdlpSEryMcrb8hEgJY/dcRIcArLRO/bb92c
QcHLsg/83aLsrL0EMe6pgdnicC8ZKWZYdx7kk0kLVd+lI9a7zJOz0Yv3kOzp3KJEIFyCDFsY5Skj
78jkaQu39pbGycs6x8+PRWrZVCM1eBfivriUXoBsLaygQy5DOWnQmvLG0mlzLTh3GxUAN2SWpSYP
0qIgAKQf7OR+7tifBuxYBTPjwGgST3JcLmLgwqxu5ZgfwovwTU34IV6XtzpV2FDrzcQ1uNnki7/t
0m/FaJalhU+3kwUISOWvfHnul1fuwBYdw4u3ql5PJ0liIAj8AsRMTSkXhtzhu/BHN0YcC0Ni2DoZ
vY1tmo1NjeXr6VrMDPRLYDRqxUwmhAXnnEsD/Ydhb0+Eq7sV9KelA6UikUa5B5kLH/93GAGLsOQo
aV8pgC6nDTitDq3nczs0oaNJIIffIl0nPt5If3BS8Y3Jv1eZIysD7xNDI36Plxt7DOs8KxoKaMF2
lzmJ/YGQ7TlOwsblyKScBnaCgPLGvMDUq21lIjZe8Ipy0nAVnMNKuX+cEr++8po3LYhjaIlNNIul
ZfDHdil5E/zKT+oSmWnjJToOTPNT6XSIIER9+1BVpwkBhyu0FrqC4e6qJdTeqWvM2Js25YRnaGvZ
3kz9CWXN85Nx8QHBMXneA7JA2JSJz/jNGhzc6lFcOi4boIu0/H1VZxvGfqDhJroYaZQOywtLpi1e
8vgBLf+LF9qb4UZ6gphV/68NrF6fTdo+TxuXMXhfIPTlnW0qqTTOMtb94e67/JT5xuy16/E2jJVC
bINSXl0AV68U3LQTXXdEIj5LU2wkj5TnqWztdJ27Dehg2IC6hP9sZ+0uFGKUh/m87EBUgyN9L41R
NmZtphpYYP+W0jhktc744ObjaGTU6CL9irvPwBi/7HRSJoXvxE96Krut3fuwZDaCLAzK0CJ4V1+P
lb7m/icvjX9iUnMyHWMPkhwihWEKsfn18mWfuov5TYfNiDqsE2eAZOqbTQr82MAdj8J9tL29MSdE
NTvWKUNiIaxFZRMY83q0pcoUH+z5aIjJa9BFhzLwyyP/oEnLO8Fpl5GlKxTjX8Nude319HRbtSie
GWGwzWYibc5rWtnFx6gd17YDc066l2oZa7pNLbzugpBy1ol/s7eNMfVc5mBEdKAueHUaldrt/cbX
3dSL97uc5nbSfQFTjR7aJUn3lyeCC7CCs87JvpExPBn5BSCvFMoRWDbVYJQDwe9ahQVu1NeYp0XE
wHhkQLQwN+ZtQYlAiRY+EzXpQgNAVbh8aWRhbuowp8Tk4q/KMIGYOTc/vf+WLziC6i6fVWOWseXB
jA3g0HZfluQRUq1WzWxrU1Ey9i0eQFFuomgWpDE3m1O/SbOdrXxQ/Ju0mu4iKXVG9EbBAKk07Q1b
X88zGDdfa7bjdbHdP7SER6snl8dRo6pNvSUyOalWrtDmc6IeTLyxngcqi/II2fYtGe34aSpg6jjV
3rRqOTmPYwrnUWahHRyRvGvwNdzsWUrqwysCuWUUPWrZK71nDYDXtIz/eH7JJ4y/Ns3Sy3UEEH5r
giACd3mZ6Qp5OKWsoYG6mRdOJ74F6pJupMW3wdf3XkoYefOvrNVm/H7uAuP/KTV6N5b7Ij+rpXs5
XBuwma6hfYCbdoyrBSwyCnXXybCylBQswG5IOTis5lSgsfmERaebmopi5Wj8DUPK01c+r0YR6tXY
wY10T4ToDqxCP30laRuCAZ1iInEjFzpMhZEMT2IwSa1mRxbhJnT/JT2zikzg54cNBYe7D/1oxO39
qtw84QBeicsR1XguSm6G18/a20DwDVOG94gEZ8PnFtrByBR8FkKi3Zi/gJ8BsKT6JuD8KvZmj0Cq
VXw0aXLlT2xtHLHFlBJuNLgUxHeuel2mTO5EhDKR8KZmPVL8HvoYg6vpyYShwKW+GTA9zgc/lNcT
Gu9Y8jAEcM400azwmw/oxC5toJWc5Vg3GecbKfBaVv313gPM5nVMBpSvdfRjbDbaiATHiTztQLB9
qqRdkLXSJKfUtEr30cVNH7f+iaNdRQztMkg6r6JgU5YKYJAuLsX+EA5Mw1uldPjF+t53YJbWyGmF
bfPJUIuP6FqXNHGqHQbWx9nEHZ9zth9LeQyGnxynU0LQd5WYAlL2l+bWBerunPAJ6Cr8ZPzqmPOu
LMc+XttTZv5SdhyttJgrwZprY/xCTozX4ffOADhvNYIW2I5axST2Yn4jNC2Y19KNBLMdGpiJMb/l
NGiVaaA8V5tdon4pAQO6jvLYDytk3Ifx8k82qUxh2EewYITkk8B5SfHMMj3F2mJd751p/u26BRJW
2DnQwDVIhxYhHkWcHmRfPUANksaadSRTO5phwrsKR4wAeT8rd90Otsl+yBbGq3m5LuVdIOx6zFCe
YrTAg2t1WkHysNsGF1r9v+P00EN7B1d5LwJk704DW47rcfVEiY57lxXsZ7q55C8DZJp+Q15ft5xn
Z5FyyHNm+bpfFGJm3x9NQ7d13/b6RizqYxOGLdXqqpQCP09UoMx3JUdoVuHjujoHrmSMtunIfpUz
JwAWaNvbkkIx/hvOK1o0ONzX/iEW0s2n7yu2MPZqIXQlbiS8lZhoR46D0GIHETN2MZ1JuBPZuBoW
Hd11sGnqqgitWIDRKdiHgvibscg7339KA7TRZKkz6HW2EA5w6p7u1Q9zI8zXljpjiB+187xFg8XQ
E1to79SZTq5hFNkXjPWBqoMii0VVsj1D67tsF9HHyjvDTZ82vtDlSykVipwCVJ5Vjo7fYzNnWqU+
eCeT8r1EcW+JzZzX8oTb9wiOE+i1D8V2tx2kYs/1/ADNuRLVucy6YY1kBRGOaBBwQ3mFVqON16uB
+REDorlKvAdqRi/2UUN1jnN4laT82ERK2MIR1n34Jhv4Q7sIQ3pGoz2zUoxsavGEGeHGRPM0FOqJ
6N/kHVVMImaGUVTi4/yh5XelvviTaOSx/dJ/gmU4Naj/tD8LWuvux2U0NpzTEpbocYG1ozL8joZP
pasTXoCHxlV+7mkgWnR8z39m/CKkKSgfzbjG8/uzQIsBu8uooF6eitLy6F3oVxAmSFhQT4hyAnPK
bfQvNKPxrhY2d8T6Mvo5CCs9Vk68wFWZpfFxiLNFqUUYY7CwxxxzD/WAzUwTnK31kvWxPLoFf6SW
YQ8ZhcwI4GKrXB1s72sBibiGy6a++poL9R/WRCmQ4COodIMG+MOVKzNrnkC6mUB2ByqguOk5mbJq
pwMnnL6zSj6HXWxtq0CSvEEQRL+BqOZNlxt+wF8Lq2nyCLwd9zRXXJt0D1PfuH6EetWp5PzGdMAa
C+/s3P0UlP1w13PKtgUx789m6Y7mTccfaTu8sTLYcE27k6Q+T/VGjaMT+kArdGIYCUXZfksjT1qW
wnwgF9RceubErsUwIGBA4XpeTfGVjq9/2crNX6eIIyH1L+uzkhLX4CMJB7xxqiemNb3nUMhIRchw
nLRwA5YU3613OVg0kyx1nlBw093ClWCiidIwN8UVhCpy+09nMlAHLth32PjiCJZpgAcEbjw8Wzfu
Nos7ydXf9N5Fric6WnKtp32Ewhd1aK9npWutNz3x+q+2y+b8aySlCDKmF2UfJfug/CWoV7k4Tr40
fSqeb7F24H/KEXIdxT/WJSCxqD9WF4Wg6vfNwlN/UWBLJ3g7TbzZMlhxvBVPr2QExxeUHhu222Tm
ilg6WAo2i5Quc4DQZCk6aLaijYpLLP8vV//Ddi6wmEs/1700Gyrm40RufDqtBz6UBpD2aJNoH++4
N9cqzuPcFmxFT14XWjIeI3yPZdFjbYnsJ4jvUXyaQoiBuaN+Gqu/nONafOHNm521+LrrL49t3w+B
Soiti+sVw/m0Vh3Rl7gzlAkmh4OFuicM2kgkhE+zN9qDBXFxV+0UnNMZqsw6EQQRP6c8KzVImgeo
miSwgUvwNupa5p4W0kBZPQ7oAwBJkX2BGEsd2l89eGohhUWJdFh2cXaUfCL69/GzJheHnZywuTQu
woFOOgXmbTTul4nAM6z9DhOL09k+3V9sGuV8x4kmAua8NAme33jXCfu/ggb4WGJMDTGzOuuUSUxw
7Qcq6avgCqKCKJkc3FmEgc00jLorjFdr8ZfWEKrtJLtDhWHVRbe1IJBn9oUwUDd+rQaUlT4lhA0l
QodNyWVNyZB9oIIcjcT7ko8twOHIst3uNUfeKs1PEnuFgKESZSwskgyji0c7yN3i0MkoybveVz7F
HNIxLscZ5XYq3p2BJ3xThj/zn+d0gLn1M3R3pZKS6Tzln0Wc1/6gMuiKVsr67O10ol0FFtkKmX05
35Y6gCIaMPYSpuWl8Ga7Ri9ImKcpULMpFRZIEkf9Q/psvddeuCW28ZuGvaJHGBVJHKcqiZ6vVdW5
/src/bICOKHatxjfYwnhYs0aJQ1O2exrDPR2JjJfE4uM3ayrje2r2/iN3zidmKfGRLbAspZEI9Ty
r2rqwdZbRL9LS71NTgKmhkHwyN2o6k3SuP8klSVeiw3rPi2enhwAjLD/TZ+cKJVcrEslvTWY2QZ6
M0lCAPA7FIT06sCipTnI0vLC/DrHnffpKtPaxAuU8BAD5AGGKOdL+Yl6wDInvn92gObHels4LFcf
MO4urD/JtILfE4A5239WT4D7Xtxm44WHpZThL3RV4tn057d54/CP/Yq5BvRZO1si87VBfHBTdug+
B6tDqEYNtz5FKCGkS2AJRmOlCp72NrhrCgP4qBqQ01vkyYYuiuGDvrqsBMNTXB/cD9TNfXFHqh8/
qiD/mGe0DG8/Zmffe0qXcvrTKCkd2xwey2D4seEiXhc2IKETabtj24QFHExR53oYvIZL5OiwsOnS
UwrlMfRtjurzGT2EonoOwAv9K395oDJJxHOhers0EF0O/HkISxFNiHmdydYpNHJzR6UmtqZ1yUSQ
C7OXMq+SI/PPfONmf3xiwy9l2Vd7BkeOM385WucFvSfeQRxWTrTaWK2VqlshuCG6kciRKJSIArtF
zedI3IY54I477dJth3wt9kftdO04pAIrzUpxqC3FWHOd0tkILc5p3IY1qRahl3T98WtuHYq2QAzL
Lw10YGDq0fwepj0r9fBpbEQ+eQ0Nf6VrTciWberkF0R7FY3E5SjpH9l037dfSPbxUB1WwrN8YlQ1
GxmnRHrn/pa07Nc02FV367cJ5mX+TnwS+2AE6b3e1MOJc7ZsPG9lePjo/wh/mRfAOAxu5nFmgfvf
7/CXtLg0AD45u+ARRx2IZ31JxPDaRanluu8nIdBBMlTBY4B2QvuEsw8/01hxy0eHdQggBcSwRAsK
gBuDEY9qj1r2tDCF/SYmIpKl/9SpeAchxDwntG8epi+V/eBvfK6CziDYCKTexivhCOSACITrNiif
4gz4TPiqlEHSjm3v8R8RbvUrbXUcLMJZj31i0N46EI4q6Ewf6UprUNcnJtngTPx+pVg1NVYBWhuF
BD4XoAJ9mEp64K/bFYgBJlFlUjyvLy4eXiO3/uaxuxII+lu21ie/tZFsLZ4/kPP6P0TggOEBoxQh
7lrsje9g8vuhOM1jBiwGWPLWlGi6BfCddnGpywxPBONwYdU1dTmbH6ZxKFj3AHcULqRIWztaM1pp
PuUDzzCvBmV6fhFdZ+cGqqXR8FgEB05wg1P1bUFm+TupC/iyvZ+g1vHJrd6ZZPThzbp+a6HAQi/E
s85WP2YTx08rB5Sshm1Ehqc/1BbOUB6jh+3ZiV6rQmJXLQ91RbbJ+WAo5lS1rTFolVLuDHEob/06
/s0Y4I7WSNE07F6fyK9dw63AI8kAYl5fN9AeqLDyzSPSEfg5l/XWFE4wTTrwGlB8VN2NMInzYthH
fvmQrRuTjRSJACW/Ge1HKkF60CW9DQuh8rusgVnfBKRddtwjSe9zoxOdiXpSMmigApQDEupn4czC
h0BKk3yYjvvMmrz8tA+YJI9e2kbjcWIfKSJu6QLuF9BurUqaoJqveK9eHQM9jmXnaChHo0Xj/+el
j0RQGd1ojkG4+Ngcyg1DpjR1RtOo4RDriNLQI/35cyX1O7+zkTsjwPLAksktJ/d26zfUhyMTO1qo
J0MOlrZQtBEL/gzDf23XE/Q5x3jctcyqfO9vgsrPGBbrTUgE7e8mGV/cGsz8EdqlnL9/lFU2JRBt
f6OaBxRwEgOlJY2iJ1++p6zR+KAZpqP3+nCSXcRBFjBnoEotHGVJ5yenSf8c5yM+H88zy/d+LUDP
IK+PIJVEs6R7LhfkuTdmEh+Q0w/TKG/LksnaiE39R/9UzuO0Stm8ponVLto3OEKAFmfu4hlRzI+W
IxnDVjWZa6nvYzYDKHUIdoDmB2VuinWqUYVBTNVkPsGvfWNz0V0rqC8hywiWNfY27fXGGI7xkENV
KkX6C8OGLPDVZcg9GiHVZEEOlaola6Nya+mKpeS4ALQcfj22yjO8ubA3uWfWQKYvFTvEDOUQY+p6
82Ql6iLquSpfMo890zLF9kpeLPOMGxb2mZiVlpLI+wcgPECdezvA9BE8g381T8/kRPSYEwLq7Jzw
pxKvkqSR+X02t17to+DPm26B1WObse+aOzSbGfI36iPo/G5gA3TDH/tjNknKmZJO/wRHyiMcBr7l
T0UW2bA2D8VXkQx0C5nE0mspUPA5SZ3fVqzMGOQPxKxMm4K2fgwuCe48vqNytHrUDPUjzy2keXkh
w4JhFvZm18J7Dildn6vveugqVsiLvDzCEUHYymGlFoQ7M1Ov103syBCOwwvSApDYtx12r+SeijYN
+3WyYfD8fD0hWyUKIuB2e/tJFa/9K4Zwg5TzRbQXt6HHGkk6zTliUjI/5gUWWe8LYvqlWkRJ+Inc
H8qaNYI1HtyzdPkFUlSlHSBL/Ma1Bxu9T3vJXqVNFNKLm8y2zEKeP1/DDObC1Fm6danFZM8qrEYQ
f5l8AbWxp8D42JRabetrMND/qeSCBVoAL5N+k81JCYiGijFdmbFoAmP/0S+DvzYoidvUc3NI0EsB
TdVCW+KRxH3H5C2E+vH942ImB1xBhlXgDcGOI1Si0bsnFPznaDaov1yD7dROeZM3O2Nyaa8P3r+t
/PU3MEHGKLHS3yYtJGNCLZuDLG6I0Ij94tOB/VyR337jqnXeqep6diVlSkHTpFQkJbQzg3Y2Jx+i
mht1tgZbVMrzBthupMi4w5LiuYDuGhcTKtjVSTZy+A6JAf+X6CBSxCm5nPw55zzgGRKMia3Nsm6j
D1tQQsLgwoU75/CRj50mphbKDvKyDR5Bfe1HB8sn8FWWn1vjlRbbrjCBimopOyxlZQDQLN/4Y2f9
6zBy4Wwlcthm85IjsfOXhP4K6p3P09FMSi0lIbRtOHg2Y2zcanGmccQ5zlctYzXwjPajK1uPqvc0
J0x6CrNYRt84O4qaaf36NSh7QvWdxnCMZOL4A0+DFo90zlj8FQuSGRGP6BTDNjYpTjjPmAiploYR
Oom2g2yV2MsJ48RZ3rCFQx9aNNg/h6nM3ysSWRO1PYSwjFnk4tdlaCM+fz13W7tZhZUf0oWhhGEu
O9E/oPPfBhSIkliC+8fBZ6lLMNF2uWiMFAnU+H/FLY4+N0e5N49rFIj5qQnmJsi01VjM7hzg+LTk
n0D2E1bEWOFYD/aN944iK2qVU4TRCu8/KRtvKYpoG8sDh/cbsF4+qZYUiv/JqUFeoX9q2joPjvSp
lxHZQrOAMZSNOf5ipbp+FOwtG7nTZkwst2zVuLTqmU6QGevAHBXgd8m0RF3O1NCAWn7IcxYYdr2R
Yc6pW4acyfoQQpXg2D/m/15ggXYNMrclJFi/q/+snERcfcqAiF2X94Yn8W7GeSd/zRfwPzf/fnRI
JWV5QzZSGkmz08zBL1wJjyi1f+WcgW9zMhm4IGo8Gjvht7GEg9MTXS3rqLPdEHM+jWfkcu3B+ALt
Soog6pzzhAXCVYyYrlD0w8rI95i8s2WCHD0Dm7OF11VyNj2VjNgNsSPvxfnI7oU0Et7Al2Jev+Ap
n0CH6RS/Sj8AUaKrq8Gg2kRvDCoxonLF9Yc3DC+ZpCnmJoMH8nX89J8U+sEUKGNc5N4G/hM9Fw/6
lPy/CuiV8nqXdBMOIKyHOe52OJWvrkLHtRy9ocreClVfcM3bEupQgRy10UanOkzpooMInuc8R+Vv
utGhCLuKfhkBAxSPoRzwp+Tm0Xme/YK80AbnkrOXhIuk8Zd0s7WpxeS0KeHZSF0FnMqKduELZQpQ
GBOjN/XCxA/0AgFVmhjPUymPF+WN4f9YNjN6YBLK4HRX8llfPiF1bBdJEupeg9PkvzuqOm+NJ4hS
UCazP7mGqmEFXaDeJAMedgABb2c7ZtBIWJRYfqpuisR6Y/7jadKhZkhWdYPFNDrwrHou+evdzH22
zGSFAJORlQY9I2VL3T87IqabJ4IChvwFQ9CM8YBUwBQ1NEHqzVMJK8+hW7jhZNmQR4yMSQsl9bpR
grFa1jBv9DUHWdrS2VNcoPJOAjlAhjpv3IdAJzcGNJF6L19/OzkvCRnDccTttqJs3ejw29Jetd+t
RzgQu3s1xVDDs1dkqhPkPsUnDvEc/6koleye2UqOh1h464WJlE83Kc+B+ElEbllyFcWxlytr6Dw9
O4qsiR5vqDX7ROVi4Tu9/E+VYdoHdcth32tJ4zkXJHzJ5p3VL2vZ1uIHBaNPLGP4pxC8TEcnmsIn
D3O7aQMg1wi9xCjXZHzN1bBu0YGISK9T7+tfwwbjbmg8xb5ri4GT9Ti1CvwYkx8M7QdnKKyFFuIN
dDPCKmB2XoP9LJ8EG5AToKqK5ZzTANKfsB2wxVKONbAVY4cgTrQwv9z8G2PIfmgBsWZU7+IC8Hzb
Pmo5ZxkrPV2mRrOcY3un0OEuZUrNh5u1jvYljZhHsLMKfgbwt0zmBEhdIPVAy2+F7yJBX+SwVnZx
zKzRMubBSGQhxGLk9YApYfNHMYtwvNRurUptrw3CyE79+inIxnq7LEfHi7RGzI6h+qdaERdDAVm7
5Iq0IlIbXShEPM5SN+iuUoblpJOx9PRgC15Qgci7bEej/i8anRg0U/7oiSrV95exMoCWEHb7+u/I
IdUNabdH9qC2wqOroUUdyJIwb5KhgMgDBRgqUZixpXIVKNRHo5IUToNwMPTNrCZWjQhJMnZKAkGX
nbsjFmEQ0h+BDM8vFW/9ANzUQMNVLs5KUR8yndNa/qCknumLmjFQ0bD5uZ5LQ5mmcTFrksfOhFxK
3oOwrBlJj7n/tMqDW4v92mGUcqabBZeSaXPmzrfFZ18/spvShvVGcoPcGuz1fOJgvoGS552beYxV
p7GM7978b+czjQYBRB47i439R2oI57/IrM0GaDXP8d1GinWi0+tTf77MiZBtNa2tlzVdEEDUbr2d
xfAUnOtWJM0fmrhJriikvYfQfB7SM/OHhPYm0yrU6oQkZBXvbjzg0IKFgpUBk0MkSQjmQxerM/jE
O9Pj7fp6/IY05q5PMizKMgurP4uvQN7xmK0vUAxSaVU+UCJGYcCc0CI9TNugU4IAs0Sc+LLzv49N
UoTOf2Sy49ypycehb1B5DxeCu1DP5dnMxHCvQAHvj+KAH7vfyOxGppifg08c91NhbFmTd5I6GQy/
eprTMGzZ0COkoBdhnSwo286KOsJGAhv2RkbuoKl0gYt+oZodgtBTOjyX9M0bj8CogfBRdxeyhO7c
ehtj0wvasmt4VlUL0GwKTetoecPKdY3Cwgf2JHTcy0LRE4zu6N9D7K4ucuuZKMXOWGtQol5rbg8e
DZEXOerzXIftmh3q5DMaLeswZotLSxMS08CIcdx6y8/RmwIgwrfbZ0P3WS2O2sEleGHD1CwjF/Vz
9ggNbS6MXP+wAsjMANM34NSlqd0DJODGc6wzNeI1u8B7dyPFusP71vXFQJXTSNsBaG+y9qM0nxw2
vVZWY9UyYLM+6PLVe2+22Hvto49E3+3st+lSibhxC9w2wICOJlaFtHiMCTZZhtt+QHhDN7ni8PRw
le4Gb+qtVw2tlw14BHaqTmkfyLR4Jy12Z5k39smP6IVlYou4Psh49HFPYWAqoEPCT7UoUfOtKH6c
+OrQ7JUmZWMvmKdDJmRbIjOezvO/EYqtG2liyznWFA7O3A6ovbtvrf777maiLZirhflHGs2IP7l7
u/ytAolRRcpsnfWFCaKliLM9Gu5Syj6dxPHq3kh4KLL1pCYhjltZt32jPdtXdvjyrE0kZEBUo7kc
lkSzD1c82VnmtPed1DevKCv4FbyQKF9HPoZ+qynWAy3YgoTn1ROFOd3TRUVE3U6C108pkFOAyoM9
lWYc5QjzzLuSwkRO2q1zkn9wfIPzIKoaMv9j/K7obR6L9VlVxlGWtlkgN3pb6azx6aX2D1vkUisC
Tnn002Ew1tbrLYTzgjMQCUfOnaqb6C7TZtw7AjTYUBzjjTia+syYKOYssjeXIfHNcrd1n7UB6cdj
WR1hvu5685gFqfBykGR+Ecl0qL6aqN0v89KNx+oQWwkwc8+SBqJ+fy30KxT1esXqanJYeHO025nO
EACSnfQfm8Aq6BEOSs2f3Dhs+PWMzukEw8tdXZS76Fk17S4yPJbGbjcJ457HrlOv0GKtlA4zYMt6
EfhmUn7p0GrscnbR5bkHlzWQvnJE1Oy6cMcfFe8Vb5zF7WfNHz5bM51ZYgYfQDExBw0j428oN82c
5jLDAef4bGpntTI+dHTm2V7tNnxt3E22x3zOj8TOxJLwc+hLVvCVPUhtnMkqLtznmDEyzVvACRMo
gVgUnmzNZfrroCQ+HDaykmF1R4KQ0Nji2/FtYAec0O4W8HTURPY6Ib6Sqhr3+OyuPQWgRxz9xtE1
w52gPoHHeKWy4q9nGydurZR5IFjGrM0THmvTMMiKAtf4RSBHtiyDv5zqiIqNg4Le3aqsmIjH5fR2
WXUyocawLP3AGt6A6dO4f4tNGR9izYnugskfrF02yK5IJ3xKP3DHXn9TcxUSATqIbCxmIUR7i1I6
bnsl5DN0cGIFAl6gGCnAUS7MslMqFD9wuzAppI34L+ebnznxfKeOsvmpjsawo0eC6D2vDJCgZiqG
nm09gqQjwvvxe230avAYHoAHR2w7vyj6GsWeSkAuBKYNFkbXmtjtRNB2xYX3pOuheCxXCMzOl1Dk
zlVeBWuowpEbSOjOJlK6/I2t49hQPSbhwULAxlzKGBOkMu7KtV39MZLCVkZnb5oQo9LX+uU0ROwD
fAPT7MQFVBRgzDrIeLobJjH09Nqi2B4tak5xaANVAJDPk5G3GA00wzYhzDvuZCJkMwEOjK3ovlZ6
FsP6Ds4RpOLeGX79a0GZBtr03HRmqyrdzGM+y1iV3VZPF4V4TDKrOjwW81KtL0RAXixW9hPOY73R
WcHljw9bzkvu3POJN0txQMQK/4QkYUPXdzB1caiJnzbRuSRPnI7WpnoY8Cbn5HEoD7AbgSTPdRlv
5XrOCyGdzhQ90LJbGiFcpb94l7kZ36s03AgfiStvUpMnL7h9oyPsdK4CLDejIZzkslwI0XywrZTy
fLL3HiIjS34SRIq2ZDa/wIgeWM1hgVA+yRo3RchPdE9tje0T4qgOdHXuCXoonPP6VERGMj45tj1k
/R6gd1pc/DZKsXoe/ogfNW7ArfYUd3RDOL0WlLHNSm9zAOo7/8R/ruZo00dUkqf4Iz6zp28tecWW
ZSm1/HRkuQQ/RvX+JkrDJ8+iuORCX9QrBTudrJ5lcPlukIB369FpYxc1E5d5TvXRWZWyVYnCljCd
mhQuS2cZ4RU/oTjj+eI5KBDhAVQPK/6YpGsAlWidj1+Vtnt0oyVlQIGSE1RM6mdE3761iBDOsoFT
QCxN8hnBXBsdi87g+wrupvfGxLyBSdu6HjiLYFoDDQJdLo1jgR/KXiG1FRaNn3rlhfd4+Lx3TYJr
EvdmmLBova23IHVYATdF4FnKDbfgeP0aW0K0qxYnL0A77rJhuQrLqzeKfKATMksYk2+bLuyrKvX2
0mCvAFjyX0i+aS74UjwBPDutPUp1uchFhz8E8zO5uX/2ucAYk2fpICLhmQ5GoDShERTKh0C/CWuj
F6LEdzBAGT9Dj04sY1DZ54E2ExPe1MZsMeyhxgKmOSKUTJxL+uLopchzLZ4hHF1oc4I8y/Lr8ANG
ahqWXSD7wQ+IdxsxCFDZ3ESG01ocSEJr3V/w/jPqpb7RG9GD1dx2poLq39LfVoE8N4KsbX8Ilfjz
2mywbpgeLVvFuAYhhMekt5SSMol0ckI3wF9nePVvYEPnvMdN/01P4VOEX74DJqTELrpGOMzN0Ogi
iRStCDKY0hXS9H9WUggZHzJct0RqebvvckgusA9EFtyIb1Fsz0qUmgKawFxE41EWaaM87+P2Dr3R
4yYIPDgxqILhWuFj+1A30JWSbWgVDx90ahtawrxwDWzDJLdzb0F+ESCJvZ8vydyMzEvT9D+B+kt3
mVWMdxrv+L5eTvhiE9M8r/uMA+Cs2ZdGWmNGUnAHcV01dCjv+jFOc21GD+mDgDugNqHwXwxI26lr
vwOuwRYZYt+OceJ+CF/n3WCtpQRGE4csBEprbRncJF6Hthb0vTxfF8uOP+lkVp4/9F2ZZZnAylTm
21kvKclAI1uENjQDIga+dME7wCP/PvCP/ONvjvpDnr+EF15X9OlHB2ILXV/9Tuah23V6K/GjXhfJ
NvE6wkbXR0i5DO2vQnh2bBwPkeTi20c/z+c9Q1ElLhcMbiTeAmUsUJzo/C4p+2H3Ldz43l1v7hUz
HwaqNQtuyTVJ4/9UeSmfobtgHKiXcw5FzXy2uxyVTuugliwPc11W7QZdZQeIwmSkE2EmRFcijGlJ
MY7XlTEa88p40A6ePZzNL5sCKmEUunz6qUnh5nCUdfuxis3zboe05v3fpL8s9kk0VKJTL6qpoj7q
N/XlXbDKDzkQAg6JAQfJNXYSY9azxI0Igp4+ln1FxPU6PHqPYmDtd+ZQkrIxHOXPRJr7FMN/fitX
NrfJTcdrWDlHS7l/N9NKN2rJBbU9m7zV00FYbU7EQbAYwTAG8JmKcjhDlQvThGxHSxDhDJogP1a9
vxsEeYjOuXr4ZDLkQTyMxxW2kJas+twUFwsn7AQSSp+13LaIp4tcGK5foxqBtIC6VNp8WQWhggcl
XtE7nYNCpIzSri/AOAwA6dKEA+HQbtLLaCFOJ0mZiHjU8HqoJoF+7yMDD7TI7wegssBoWNwylS0Q
5sZpmUrXS2msuAmx66QwzQRsc2Aq9Gzc+gRm71jnU87pbk/Wto29Xh4TAIydI1IfJLNnt7YTnage
AoqUmZyO+ZiTUf9+bMvDLOIcosVOtntN/9Sjn4jk4u73hNf53cIRq5run/QjSXyZ9iS+/xSv9kZE
hGTpSuaiG1AcBjH5coS3I+y1zfXugHNbTn6C7oSEEKnYdqcNb+hgboPz54UXzmi8/PxFhwwBx6H7
JeJ9QL3cIpKeTsf5vIV2YM75Kzz0eTJ/+40LzMZoJs243fMeCQxntKuUNn1BDiBoFM4nV7ePdbju
criYHBXG7JRNR0Wd+TmMaQY4k6miEdMu8X6ZwOU+exk8nj0UaOXTcRxnPuCVY2kE8I2S433WRadN
mHh4kj+7VAcvTgeXfqoxJLoyRnf6J55Uh9ns/q/q8NNJbBFC1qUHA6y9ysGMq8BF6jR9jSeIyhOd
5GM5aXAG/XMiIMh/snDuGU7UBxL0KZKOCVjVszocVEY2e0SKhBu0WqGIpqecVcUejktI+9d8F8bT
xEW+2i45q8fitnd2Qrp9u9fpt0cO3tPP9+XWROMjqOfe5TtQyDPuuK1YkJzZG0YDXKGbk0XuKquE
S2eoMKz/ISNk2moTXrYH+2iDHJer2FX6vabBadJAYoJbvdtT7yJtej+wpMV/Oy8sGQOf2uvNodXP
HK5hle5Dw4o+M6FixIADuC5oSKBehHP9uULfQofjK9bIMmDQZsLEdsPnWbm4MCZs2NQURvwLbuc8
/3l+ENcHi8QCEh9sW0ur3JxVIMvb2kLAnv/29uZ1twNqPPp2FejEHWGfcfzXfosbjksQm5di/NwD
gXWQMw5yIVE2TNevm65v3TDT1KFRFNgjVUVUx0pgJCi/eaab4cYXRxmjX0tx+9riVg/+tvQjXHlO
oHV8gAzxDE2M/ZysKohgzUnTo6Ek9+piIAyDp+3xRt1wUdpuNDe8AYq61hhWhN5fSInzY5yb7xem
QDxbO4Ir71HiE0yky0mGenfLvDGsJq6YXFY12LEbErl1/bj5i2LvYDcjq69zY+uawvwJomz3d+yZ
MoxsODORu0Yo9ngv40/I50H9IIKgDMyNSotHBBiVnEmdUQOlMy43I01kL4SmHeDN7qawQaRhTcXY
IY1onK73XRg/0WssqXlRRgJfdlwwCBjImXcxOByidPwNtZXo6cIhIo+yzh7OlIZzM+VE+Jvg0Md2
3jU56F90OQUurBwO5+rjTCYIWlurHPB2A7EkUAMExfVrAg2tDfVvxLBls7s6rP3uUZq8tiOW6bal
BFN3M5Yb3QH21u3GyQ6Lb3hbXbBC3TNHYo/xmsw4+ozK8sHad8oAh9dRhqKDFmmZBm/eLp3+7bvE
yDpe4cEOCDGmyV3IJTV1/Acqgjyw5XI6uqcQD86uPEVWsvjJfjUPICf6RxlzPaJZWgt1qOTXIN4D
DGCXS2XWXOLuNaFlhpqXOI5Rjadez9PWBhEtMPvQh8V0cGLHly3bAV/Om8uDKFa2ZrPpaemkGQv9
BXxCiRDEDnd0GnQmQ8uWhc/iEJMfb5dDSWZUsXkQYOOmuEsGIzJWO6nb6kZ4j1hwCTsKcvryX1kJ
D2jLE11asvUdyLUwEcrbI8z4syOzcociDoGCxu+PDlZZx5XAqVxoVbBRmFQbLQJU0Fc0Ukrc4AGo
mkstUp/IvsKIIWqZmWtPyouLBKubiCNh4TuBcM4dpcZ/7cDWC7hjiGsPHJtScHv0YIeX2f7+wmxC
MajtHQG4+WseOq0g3u/4S/E2iaaWsK7qeKc5KkB8kFvyPDdpQH8PnrjG7pBvesieSsKczMlhBH6M
6Y8HOU6khM/7+0lMDEr9QadHNKIaU1nW3/rXwWtudZpRQpmDKUSJujPvTA6eWCZr+6zOP5kATRGS
mmzrHtSB4Ri1maYkQZEUrNGuuQofgqlersdK9tvaop03ruAx6JakzMXzpJMCFLzmL/Qi/GRU4x4L
oR9N8ZLPcYoak4qC0cZxXrKF/vOXRtbQqp+Rs6UYzlZEb5k3HikRf4XiwKKV0KjohnzqgwuMj+d9
gMiNshNcICE2FR6x0pzxkHacvGIIX2pjbwUWt4QDFIXPuzZUMR8h/ZPRdXi0r36EIR01NbVYgAA+
8zdpQ5maXeaTWo3QLwN7o8bLym4MCMB+JtjsxPyP/cd19GMqKlBsjxqekNSeuGJ33ZwGfP2THYKO
m3u4NYyism7mD7K5uaoUOidpNH5iH7IGrPLfqcXxalUqK6O3IFCdOJ7qEFTvhkS7cHI6O4aGJ663
LbwuaXwCNyZ6o7ya9x0ner0JfLuCgTEWBjqtdPQCQ8AWU25fOEt+T61tdwT1cD7tBi7XlsdEM9R0
xM2e5Bz3Rj5nmV/eR8Vstb8DuaqBhKfWjOtOiC4kLZEeIO4Y2VFcBSlBAH4LAEDADjvnHQHBH8UQ
v9lh2kaEsHpvB3wCLWQgvT6RlxLUwjB95wYjO2TsT0Ks1iaMptE844lHyRPN92QcfWhzO3gywTYi
+tLoLxLDSyZx60cqYOqjdF9Fbv+OakAsonpQ7sr0r/wUzfrEOJAKDPDRRvv/H9XQsmD/Ujo5QLhG
CDcnvWWY8DKcRV4EQDJ5RRP9hNOsM0aYcETVwxv8kz+DWCnE3WJQ08ujIuNgsxaZkZ8iDF3FrIgI
aXzzJJ5XytiMZXfkL2wWOnJmgQuf4wE4kBra5A+wD2+mTK337KnW2XYyFyyxch1yi3nNguFsRKzX
HBOmdPS/v7zeCy6wD2hfJakp50bjMlH+kZMeus2bKrmKV77Sj7ZHtNg0AlkvBaup+HCbdR4rN4wM
PyXMeN6ZgBL3qxeKPG6djPKn3xxyXoNlPMSpCyFT0W6xibhd4l2ivlrk2+V8emquPzzZrHZ33gx5
c7vWY64H+fBIWr0k21PM0ZLTWEQbVXxaNMeCZ4nPzOpQu6w6I1wC5jl4xjuBoxUcgY8814jkuLND
FPPBdu4BXGioovaHBooKXzLU3/wHZpRNNbclRdUW6Pb9UeKu+5s9rbZbg1H65wzkf8Atr+ERzY7y
QcqArD6018S6gb4hX8D280MJrWCoEnZiPUWTH/uBX6zacZR0ylpXZpWFBf2lrBVs4D0LDEj8C4Qi
XulrjdMb9nHv8ZPmF4dStZC0T7y1Y6sK1tV1FMUvF+00yY2+rL2HswERAPn5JB/iIY3c/ZDnR763
0Ou3niKbSYzXovXTHF+IWP4ooS5PkgG/BSLDYHqS0MmBuGZAtErf3NqbQQ6/bBnq3YfN7eSeEP1n
2ydSkcOFjEEJACvmSYXUtaCwLWqyWJ/bjfGzuEVAuzdkygYkgNAPsMHv3WAAHgWCk5ltTp8bjzxF
VGb/S2d5/gWtcDgZRQBjtuWkiLISxTCF5OrQR6X0ZSW49JJKPCqd5tHyErPNVPT4TTfjekiretjA
T7C0tSpp7ndfveDObsf7p/e3lB4QR2IpcuYp9C10dVBAStI58UsPBfZ0Of8z5y9Mac21vqPDlxTK
PYfUbK95L25aXPZNJQak7pLDgLtaQ3oDIzt1++QGmDE2kY8k7NK2alGcmt0z7Sq4u98Q6E2lps0J
OrXxiAm3SRzY8CtfeikHbmIJjRigiufilf7XCPz3HWGzmBwnsOrhB5uRjzuNnpH7NdpCesewJOTO
wQdEIrygViXlNIbuNpJz6d/Gtsob5ihthb7OZCF9TBhVbUG5vg0WHkCazH23GxQczvDKO/lEqTc6
QkRJynjZMU3XBjuvvcgxijRISUGgoMt97pzJkHG7KIqa8wj5baDQt7eE3Z/kCfdPdizAKwpKFyh5
6iHEa1NEhVMToTyyRPNdxAlEqK18BNGQMIOHLn3lfPYgnQwOAiE8gXJUvudJDsvNTdFaNnEvHLeE
PUbluPBVzibhE0v27mdV3Y1kXZsgbHF+BmUWZspdu/qGKbWCM8kElHUNebENO+sfT38ZY5ydkS7N
vD3RXAB8OVTwIvXZhH9eieE3FuYuP8S+Yu4/YepHxFpblGJugGLzJWIW6mUfnleXBAShCMZyqSPo
1zSMcAXzfuS7AOZByDQyxIqXhkf639rhbYchB7Lpgv9oJtkrV4bMQD7h7XocK1VTIDhzjZsaF0t+
RS2tDgS3J27HSKP5MVeAoufYuKrUqblFk9w1hb6bijgXkh1WMBJa8yabqrhmgUctda9ycWN7RGqD
XVM4ZGsnBNfKJnnYDgNfSq+2YkdO5almWuYsawbqmOwyMs4Ws9igKJ8lNXiLJoT5ptk1uTuNsi8y
BHTJWuEyuDzdQocyy2398y9fvQsH7z1mDulp1MAorDpnANdqQunyH2PScgYZ5CgK7dVU7hbz8nOp
xD+RmPjtY45UnlWYIvExqGWR++6xmzVMOGOluzFD7ibpF2O6WrP7ZDBg5P0uct6mOf9dSJcuHqhS
hU0kOPecc5oKdPdj2ODemW4hzxH69jQ6NOWg8aEgpY5A3gB5BqMExUTD48m/DNiUKMfFn/5CaPVA
ZIXbSQSUTtWYtDa0KuBnZKcLL/SZPAH7ZGvW57zHjFldbethkf08zdu0g7ZjFlu5ux2d+X8S1pSy
KxD5Zg6tzQkOjMZfk9u3bSy32yVCRAMwGt2koxwn/al3WUJAHgGEFOC4g0Bl7aMoovccBCIc71Zq
G21woUCgDKrxMjyvRnNI1pbY/vvXZHFHuaogwKDmks0Htp34u2R6y7YKa9YVCkcrMzphbxs0os00
C0JOi7RwOUBlWhBvadSRGB2sCfdy+cGUiBHHNQuiT/LkYl6dS8VAs/ieHNl3v3/YhAGUf1bfAdMT
hD2nJ3Qlj6/b0Z7uRmgf2OCEmFJVJt6BWE+P6wbUYYWU/zZuwsnJ1QHkKYRseW5FWLtfML6MnyBF
m+N/2F7SSHcph5jOJyKuVeuN9ee4m4J3v6+yhC/0NI7a8AaDKZSBAoURBCKUzLyutP54JT0s6evP
JU7Oaa+I3gyIfG8aPIJ7M/Q+JeapMdvAwfq7koYSh2B2abza22ADwZ7taicIXgLQ8eJq8kR7emXR
7ChNK1r+g45paUzR7nfgLNSb4nEGuW0DKCyWdPk2TCw6HKuhxuDuoxP1YFbxQfJwDl6nj5LFOhvc
kUDGa1NO+Scc1ho4YCTgCEASrFYoCnR34q6whQXxZBLCXyuaJotKG3xVk3x4bFBKp4VALuFOwqqN
x+TGPTKIj0Z2bGsamboLLBbaDx9/TIFl16e1UqDL/ur9qWo8PlKuivwn8mG5QKs6boxT1aWzFLRk
nLv26wLWOVu827xAn4Y9RV9dFIfHmHUamB3s1MmRgro/0ZW/sUZ3os6inihIBVy05nGvtEVGN6EH
Z/YcB8Zw+4YE+msfAaIcshE10AcwKYekqhXCBExtkTlEXQAqqwYcLe9rG4H67GBTGqKJhEhFSotf
h20coEkDijC/HZwl7tzKuBgk9h6uZL1kYJhye2Kd8TxNK/IJmvpHJMj2K0bjYzLuiR9t1YYJM5Rc
OqM/ob+izR6eXsCAle63izKurDaDsrLKjEfzpxX/JmU4CcOZE1a6eQINtC3CaQh8zWkPrUjtPZNG
sSGSGK+d1z5Zv1qyZjnj5hLxGNFedDfQpWcDEx/jpDL6PqMABkFpkBKGFCpPFzxKc7XIUqYl8W19
6ykGl+7z3aYGCtQK8KGDgp6cVDATXDzhMS4dwfejSyyWH+rtMcqJrmJoJ3J9kIRgFzqvaErQKc3v
NKZgQNBWXJBfbDCcnLF63xhVbCU3yf/VycCO39WLBYJVieO3XUlUdMGacNUcTHM2PP7pzO8YDH8s
v6POnvCgqWeMW+zpgCYAGlzGiKX9PkYSpEwhTQVYrjIFPkETyPtJvK7iokrEIfZbCD1e5uOeUNYh
Q5bim7DDKntfkhEVf0gAdB0kdzZIUh1PqisQw7Y/cow5nV1+60VrE2gw+sGU4N74IdZrHEOxX6DW
LrhfMo9IZBy2t6kR1mhe9xOBIa87wDvZgvK2lLAlrhxjm5218vKYOo8WnKoUuDNl6lsiSVlJhMbA
XFpcR3wZmEfQVobERRf8NB4QD17WTtunxcbD5/wcilllvzZT81nDH4+hffSbk9T2K3OrYOnBh0vp
2JprR33P4qdMHRfMqN7NOq1/vgsIcuSt8whWedHii02zXhzWq6ujODQB/5LGGYW5Y7AR3b5l9QFy
zduOC/Le2wekKhmXcR61ZLHDQYwKcY6cakFT+Eq51d1eFmP/KxtumJh41WYBKCRA78ozRZQbTKyS
RQf0XWcXkO20BlYAAZAUXFNC32/ylYdJVO55EsDZ4hrr93C7i9xJ3trBm5Scl+ilT9NUsXaFmpUa
Y9fcEQMGaxLa0Wb/9QAU8ifFagtvplSo5kKD4GI/W72CmMacmhgtrh0m+4yoDTWWUGA4MIkFwGZx
nqFf4tREjiCG8u4rYV4eC8CVxiRksvECq27hAeihDi76fJwr4voZDkKgGRs89hI6Lg2aHutfrnRG
KUa8hgurODwYuY5TD+qRnSVSKnarh/EwArQX+5rBXyaAVj4W8HJFCJXD/O0m80aJ7v2P76TyGsL4
JBZR28PPRwCyai6R/umh9o1YSvgd7C0f/Pl2fuWJujL3jygdgwqHWvZKfkL2uk5s602rDNKrbLp7
ZgT9ccPxINEKnlCE7RAB2+a4Wi6g9EyGEZMszDvqHyrbxmT76vCV7pPnN3El6GjEqX+H2X1liIBJ
lUnJQc5cAFJIWRZCOypg/x/xKluJi0mw7H4DL1KPHrj5hFMIpKzoD/fAnfXNoIsBvzZuA9dlLwiJ
zcCaiD8B2ifg44TdQG8MTdnw5z0l4UDjnrkoI0/ZecXrmoHPxnW6vQ3rXWEKj8jsU1MYFurCcuut
W8aQo13Hytb9Ecz/sGkWdrcAikSVxMMOu5XNoh4vQewEymSGsGtcTDKQ0Jzk1uw66rk4WJzimShO
me/dimh5zTcmx0Jv2l+k+qcOorl3IgauT9ct0tnZ37Q5OJuPryke8UYfd7T9J+tTqn+JY4e2Nflk
1Uv67usY7vb/YkI5dNMPSDl1k5PBUNpEOiHiVw+uNCtmRvztKZE8L8HXaU5I+Y/KRV0NghW3LaDI
52wW4YBTH0t6/INKj2Mk6J4lXQBFkO95GHUfmasZrOvEPujwriJ8RxTd+1fuqazozMGR+/4CRlEX
1Fx7lZFly8OnFdPF/sSaoXG0CjyL2Q5N3N/iOniM7UDQE5SwQ/FPIs9nYXpWXjwRw/+Y6RQgMTB4
tkowSFVZRWnfB5XDSrCrr/FBlE0fAR4WK4R4kAao2CbSe+t0uKi+jb4eIggcBR1bMB+zasBlR7DD
x5AQVXNns6zboM/qrbX11crY/IPPpyYJ2LCcyvS7ABWPkCGw/ksbR9ehcNP+HJ21/CUhIL/i/g2j
ULGvpG1Nq1a3r43I4Y6BSVmNZMnFImqaPR9nYBDJlCXdu1tP9134OkYI/5P16Y5xC54bM3RNIO6f
TH7HikVAKECsp/b+hx1+egSV/N3m6T9FA0ta3kSwac5gFDukfRmAvVxq0+YMpWmjoykGUNrGTPWg
aP48MjHTb5Enu039Ph61zbBtumyOcFw1+zw7X6Wya98aGZtzE2rHgsSckBXGpp25yaduxJePDvHd
WMERNc0JH7Z1L9gAtnDF8lTy/P4G4HTXVUqLdXKJG0m9CB7d+FRHU7sXR3hndmgcP4nzJLzJGQvs
pMLQbN/Q5jqb0EmTUEYAekDyQF3zFpxgc2ZiyjcYg3Qg9oKKTAuHJl2gN4Hf5sLcQ3kRsJ73iaxR
MjhLeapGlfOciXtHjNGzuQOlKx/Sfwaa76bCAW49Cw2+qFlYGsflkz0lsTGww3MJrkcf1+P4g8MB
MIEvW+mpOoWoVIS8w1XO7rUabISNGiJca4qbR3CnZrVgKsUbi2hwY3UJCrepfNUxlqPWPVWhUlsa
+KnifOniSlmkPsUOFfl8pLC3xjIdMuFpk8pFOfP5RqELcMHALTKyyDYhSUJDc9c6oxpDJ7OqzK/4
YN4NYIbz07vgGcWtfXwAu3PKTDDdLFjaQepBdU8ncBE1+29/JbsFjg0wDq+afE+xgyD3Fi/KDxe5
rVIGk6wIhNguYn59Pc02inn2+GIAFPLbMLgfcJnJGoiTdXVbM/Yp9BRaSnPZgQf0Cs7KxOUgnkhl
N0jqaVf3iALn9oDRzcGakzpAIM87hJlrMEWmKOcZ58zQqSwHl2zjEyFZnFaV7lWYeDkOs1zO9bIG
zitEg3miG7BGsZhkRljWz1fjMa7pxoznj7k6boH2ZazXDyoZ2bN9hzq9bv64HY+SuZ3UPQ0VDgih
7KUlt9YwLzhvfvsKSnvW5MJJ9r2MUucp/xHTX0nVIcTm5jRDdlkiDXmFqjD2ZYPK+MCyFznr/XDd
azD55CTMof86AoSbaRrFpoXSmkvnkgS7IBFghEJunOa/3oLLcNgO4mA0w0OYZnw954e49vrV7co1
M/zR5wEkd7qC2nEavZL6c/tHFFKth6dNtVI2zFV94aWwyT4Q9ErNahfc78DgVYGxWMYQ5eLYyzA6
1eBL1u7+sSCLa/ihBAwoB5ctNwngCwuG7dU3VOWCa6jkDYjvS6KxiajLU3JHYNPUfXFOjORVcTKy
TUMif/yS56QmV0EqS45Ul34p5Tbcv/E3Q4p4zWNAPhHoVNPtvqXovyPkI9lU/ia+WgqmDX8XxbA2
x/az/xaMwQb3U31G+cu+5bq/ZQrLrly0lvPuphkvl8zHtKVKkO/rn9HQqZ7um4pcRx4e4RjgkpZe
yvryEbPv5HIUyWubLyPL9siFxPaf7OsMKuCHkkcllFs89HKpqk4buFnPRSVuwTXqcTg0IfI7j7AN
UfqZEohFjP57hZB3Q/09Xjfw/Z0gf4W2yGtCDZZUUf1t9Ze/aYbwypxlGOruS8HNwdIoUUuN4WjA
WveKAf/k6zPShWXgYLd+s4i0Rv/MCUP7AxaUi8nGfx17vpadcQUNlXifljfJ9ife6UBFdDTL71hc
BgViWk7/Qzsx3Rz4MxpXcLpJyRZwNAneQft2fKC/mQJuWut2rcJzAwVlOmsoj9e8hN1gstO8v1BU
dDE2hsGE/ytfKdR9DlESke9qgz8JQw1er+fxr7bO9cpQkJS+/3DZ0+LZAysi5Y0SX96TT5ZRZLxF
ABMPxwk+Gkhzvr403wHgxI8zXjSpp4JqVF3y2I5zAHh1xHybc2K/1n+Dsm4d36GfnjvZVT0TethX
x3IFxb8Kda5QtbRdYzScDWaamDl2VZHKfelhBYSBdeR6uGcsIwq5NZ88JgrqOIPwjAQoG4d6FFvT
ZyektgpmOK844wFSaesnWoy/jE389gFodHK7DI3KkresgH/C58uya7UX9QyEA+dUBP35Trj+lWNb
D20XZtih6kamp2XyV5c7WLv91kjEn0H32xkMjrdSUuMHfpy+sgQwdI3enQPLlachwtOIIrC2lqfK
WnlkMKJ4gBEu3c1LWd+YWWTPF1BdxIKHA+0flZVolExiUEoQGkMlhxlj4Q8fZz4vQGJl8aAaJZ8O
fBqubzqq9G5KEURpD8zQIHYR1h3CPPAFut4XTORAxnFjImCqib4q7aoSm9juMiaJRAEWMcfwZIZF
HBKLuwylhIrUxk+MAEXiUzRqsvw1uhUEtNEIVKV44CZBH7c4TySOLGXMWyb0pfyVJrSYGKPlbE9M
gN1vgDT8tKDlQac221cYHxJ/RZh2F+rITqMMLwK1tP84STOD2cntN0528/u6xXEKsk23ic+MqLV2
23z+haLAql44W4bsuIauBqBl1GSYW//RBbWU/Os9i2LuKVRj+V3tUopArKN/W2FsirvecGGSKcfW
6O4AOj3j9AOnqJ63tktQ7V2nJJwyRiCUCQqKvjxPTErOg8RwO7e4VDL6g8YXHcRQUeoomz3VrXJb
umP4MT+p0FZ97sDRm8JNXaEppJ+BPxhK+bk9nKdgnM/r85lQ3C0U1TmSwpSbKtucqyjfttTnXIK+
QpJl00V52BnSbuxVNBQ+ztfVEzOcLJbv8eYV9qI+9KtsSnVPCAXKaHPiqfyqV2zlzMiKqjaQDXiB
ieTgMxf5UKEMjnemJppPgazIWPFfNQ9QeSgxzlSjzImE45FkGz/Y+PiF1IPHFGrnQpVa9V5rJm/j
y+z+GgNY6oRakiDcj3OnGl/kESShWVLWsEQEyFvMdel2QyFMTUgCCcyZ1psw9dgN4S3jfgxBGA2N
U0LhRrJfUxLvlSffnnXPpB51DyfrGQakSQ9oWvGqT6D60k7eQVKEI1KhvmMcLh4WBdW1QvWPbr3H
YDbvngfiJhnx3AyE4peieMWiLNUAYHp9TTxQlhiDAFapXRR//fcqFQjsvkrW5t9ua4XIUpV6n7Pi
dmy90RYtth+bCVEBMBdgZRfKkcu+7fcGp14S9dnoewZIQLIdSpRGuv6POfRTKXsgdaCfHgjn2/h9
+LrgOrklpFdpPmMCzGDjvuZQRMSfoZikaXw6mqpLwX2koCZ42cC70+NK+XnihKZcAy8ZrQqsmS2w
8Tf+XlcK4rHT0Jb9Zl7pyAUDeUzcHNeJ0DPlOAdH1370OztOcSOHmlOl1mTk+8oQ9IXq/5M1PNTQ
FUTHDtNDkwRfFh4kGD34B5jtJqCmerqf9fzjLb6qdFjmTJBC5uK42prWsPFqX3HzVxeLRCNvia03
fbkZRNtNVhjCMTO0I2xutJUQgK0BTpErqX6mlHXgkRYouaqDsR5/lSX8qpFRyOAcEw5CiIMpyQb2
L1Z2O9PPJrgmheAyoLsRsIB26B4xNYY4Reme7QEXJUQ5HZZM4Aeul2JsN2Qhq0rMYB/tovWkivAA
eeryvrnHsflBupgOweI0Mf4xAkHCd1iVeUpb0JsyCY6d1NNP6nfNWVrhsxOpllGPR/I562zq33Qf
HySnk/1BlXUbX2uRZi+NOIIfXn7MKy/O/yJSRr19uvDpjtz48/QU47aNQ4TrTkkIJLmXCN5dWKVP
Yj3ws5KRSGKtyryu8z+Qj0hoxqMGRovVehtDoJr/WkN9pcbjAP0Ztjh93vctRuumrXjxwPTIK90O
6tQZZ8Wqrw6SGkD92fLzAvPfV2wjn7snB7SOmJeBd/L2l4lpZ5SXD4g5PBablcIZrLjDs2+YsmHC
B4fD9w9lsrNLA+0ewHfnRfyP7KOU330mcCJnhlyj7pR2pz4a4yVRomwgsyVIE/BLDYrhv/780pBe
ymqCwis9wQVqZxxHRtrozKIBWd1cUJ94SOKEL5/hcqJqRf1wLUCIaOZIoO3vjZU7Z0xhbWZbMHcH
/vZmsf3FBqRI01GGrIhOMLnGCXGfKP/Bki3C1D0J025ZZNUzdGbXTH2/jhiyJtmmzrrP5cZQCF2X
k1WLnAzDGSn+92yhZ9mbEwE56tZEef5YZ8nD/+Bzwrmt8QkEv4IG4C2omLh6M2Pn5tRkd9BIDeHf
SQRhwuuDzZIpZ48+32YTk4WYoRviFw5SWhn9Aooje8acSl/L3G+4zTnh3YMxCEyiBLSV2fjlCCjU
1GcqbdHubBxg+4rcZB8HZWbZmTl1vNe9id0/ADQFZR7pKyRNNgSncZSsgNTI/kMe65Z0oALcN0/D
+2JRs9aucMBUGAK5MGeKFg8T4c6IAUt7xAvLBvbT2QJlxbSwHwaC+fp7pgXTuqaM/5L+4MPua0AV
kuFk0Ug5uAfK5acb3/ZcNjilQhG9Gm2Nc1dhzQimKZEUbHwKqB9Wi2ZLEYfQlU64WZzbtgzy6tE0
+dvJjo7Xe9qYhpbsWIA/f59RnvaoRE161sY1T/TDmGBysHfgQEKqMCfJs037fUtjTsecAt9MOAJk
Viy+wZ4AT2axbaw/36I08totXJd9z1SVxYnzGbIUJmEoig/O5A4p9ZH7ID3sf/8nORzDyPZ3FIuL
PdeB5WWQeoMPfPXh+vdIk9kCanf7X7qCp9vwmxb/j0jji8eg2Ysw7LgeHqGPNOG63RcLXxyhbYaX
wvGk33Z7az92cUE0q05AziWqlwYP7FNsteh8FQC8RB1fpUn78c2GRhu/VUg2ZRLKW37J2K23hXNY
XPp1y+GBwowajavQ+gZfCz2FsTFERNhTLaBjAiSrn2WpbQ2fBLsXqDNSxHxYQafXXAGrt3pjABZz
jwGUOvZg3oipcWd6NJmRxV3Ca8ANtckGJB5nAjB0GCd3PVzBQsUVtECUZssZ2gwZChpVYD5cHzps
edgRBLwXqA9GX4P8gF4l0dgKwP83Uhp1KONdJayxEdp8oAD0VTBsrwC5usc+EmE4ApsTFS8dAtoK
6Foj8l1dHkwdIdlJa/5Ka9GO0znYdxXy/kA9+DCCJ+077gu8H3td2TPYI/60hMAY/v7K6YwjaAdU
1LnjG7oBwJtznVSRoETU4Uks2a41aJ+SypSeDM7jnrgFUXQkyRqMm70/PaVuGjOwfMEWDtS5ZFin
Z8K189+OfPQPlo5c6Zzpu/86dcxrn0L6VmTz3BXJ9ON5mH0+aysc7KkZM1+/aJ4H2s5Eood9yPWt
3C/sXAlqaS1DVbeEsav94E+9YeNgajennFQMUSoQUccwGPYmWDqNgSzaoOfFBFbSHMcTKbJWZPl5
oBAbl07bkqSLqehrFb1v0Gsjpbu2ih7UB7qQfaMrAS4Pxmey0dp5LeNOk2WV6W8ud5UUyoOvMkca
tEg9iTSILXwp+e5mKeVpAJMFAaxnJIU753We1uw6CQbd2fpuyYLv7hnBvvslprYxOXTiVo+az0WY
cq18ez7yCy5BuStHtXrH3XJnElUD2MIKwH2T3YsE68y0WMoNeHKC0zck6Bf00nBwBDA5JahBvxfT
PN8A1EQKR3jAR3W+6uGfAmx9AeG94ADC8uf09dK0V/EWx8rTbAsilcQxbKWqwYHxfXFIKImbEf0c
Xl2Wx7pWaNA/Gsqckw63nE2MPpypm05aIn1v+fOQD6rU+je/UYsYUwveUb/OcxuVKzL+Tsd5bQ6G
2gPVreZTx+KUqlulE4G6H0AUjvCKHGWhnvzNU8+blr3bV5ZJ8wvAAoHuoDryMQh23Q4tKwCOpelp
5s1EFgZWGHg8x3W/KiBkYmzOnttPT121UGJHL3RBQ1ESYfdRwQNlSj2cXTavzXbdRTRUyVciu/gd
Diae2zlJQqVQGp5D5JG886Zc1foJg1qztpU84lHxtaUyYiboa/XeRqjMnMfYq8ojIihF7YKIaMPo
VzDRvlxQmRZqQW/xHAZnOIzKvqVWaw0XpPxbwyNOz7ObfHo6SIABSCD2PldDfgA1c4Uscs9nyrxP
xDB+9cdYUeX1jRAegs7aGijYYWeGg67+fJXHxyrlmNphFMH/aqSPuE2U9mjCiURjbS0gwy7NwmP2
JRPUbeRBOykyd/bJ1HtXQY5FkkJZbZ5ItAeDF9fiykeowKLnZXZyL4LFq9AJ1hWZN9E1wa80/w4c
nv/+2mjvXQW+MJ6V0aYGpfEhSgCaesIEFHg51/JN++qgUSs3NeuDTJ3GWzjlqTgImCPkKPQUsH8O
fR/cM1dCFk+blEeAmeeLCTfUniFB0Ik6Qd0+lNXZWvPTnlqrFQvmQ5re58YFYfNFfEIrGO4MekGl
ydqL6cO9wNHQlz9/XtdsFNTlbBpAdLf/43nJpx+RbAT45SO8bxA8mXwcRvShb7mI47zcSVblE7Xh
R/WbacnjxpErpVF9gP1qlldRTprOVIfbjboDhkPGFA6git9UCsG4HmwsJefGxQzycZmPqIBNKy38
WgrMfc8LvTynVkzcXJwf1hp8bcLTFZSxjdkP6CWi8uVmyNe9LUY8AWJ3Lxyv3NXJVHsXdnKoYbG9
wB/4LAWgWAUM2AaXQ7gVyVEGi7roT3zUYiNYwfk+DysnXIVQPsYzqV0uEOzeqTu6ji0NIbN1I5Z+
BhPAdMdkf1x9xFNjEm0DoZpo5bRL06mmf6uA4GLULs8ZSPijvKii+qYHnI2iTUMYd8z0DU3af/My
Ic14FYg6nur5ytJoQlltfmE8Qvlmi4LbFYhoRrIttsV7vp7qLct+i1SDQ83KUbuXOpj5hmSaUu/m
JLjqnPt3ticED9gLGweIaqxTmvmBgyjOmwAX1YbSYFQK9xNPs+xLlFw23x8zMh33OsUBVwXejSP1
KsiGBIMrQ0VcVooMH75CccI8hZ3EH+TVGdPw75OFeTvb67kAtFcNzk2CHUFT2ExioNnrTYBtszS5
ew8XMZzlD92g22CoEpTML1mwHGnYUyFFdmfMWpRC1kM2+suVHVsSGPaJ1m1Q8HB8S+a3yuRjvNjv
uwzyvd9vgUafepu32oX8jo+nqdA8GcBQS3Glot3lFvW4i1dRkHgIjC5TrgaoD55YvmN4u4bnNUwX
6uGGdmzYiw3tLhn6Esyy2YgtbvOE4gb2huYYBM0BClKFmcKfAKltqIdlrfzwY1clr+LC97X8qGXg
QoNncluCaNA750s1JUOTDYfQebOqFdg7/5yb3gMTMhpJJqYfwm83SkDBDMtT8N2rOfFiw/6ZqOyU
ETUxJVMm0TF7UH6EZ9LCg2rvKve3T7R/1NkFOSPlEYeblnBqMIozLH8aOOBfysgvFkj3vqYoNWFW
QeGvFrVziALAEMDwfDyLwwGN4Jx1wgIEp3BQKoRi3RYb9PCQj2MfC3cYE3dpflPLvmLRA+bI2ygA
74YW2DGXzLwFI+N2p/csRvj4nF8Ucr0I+qHcCDJfheWvz/U7SPf0uDvR1ixjVSlyleTp3Vchll8l
EisNof6EPWFCh+z4MtUXalIFNP15tZqm+cuzt9zIPrxUPuACHKnfSm4rzSgMw++kdaQNHdypg2XT
mVfXxzFK4ds7pfdKgal+GLstYuj5mwYV2oe8QBXq6rGgAqoThqIXqDbccJLCbrDinL2/FaEcoupv
ebBwiBdsWQ/Qog+L7OAfrrQ73GpEw1Zn7g4N9PeBqMAWhTN+GDS+FbLJBxCylPTK3QFDH40+0Ndj
lDgS71b/mX6U/Iznx9xvuXX7+H/3OU8RFrPyxWnMsFD212FiWUzAx2z7bt55l4iDDQYxQv1yVTkC
h/j+O3/54yIpp5duBV0nSqDplXwCXWjKf8OZPHYEVqsEMwhyJUb6mB5uo2rCJ2R2JXWOGZKeCbKC
2SMz7+UDX5+Z2HoN9LDj2/OjVQRnH6pUoF2ZjgVM4aZPPUPfXN2gwx3EDAqv6mOqt7R0yGbI4mUV
fRy39X0xB4INH7Wf16WRawdABmg7fn0Z/FT6Tt6e1kuSyWgW9nLUfIVU42HBcIjbofqOyHuWez00
CjbmzhO/2ZVQYKPTDC/OnLkh1ne5tDlMl8N+/aPN4i9vX3lTO+/p7eyik+z3E5sDZsMs26M2+RV2
OsEiuXP+TXKG4sxwyhHSYWVTvmDAxFSpAfS3haMxhM2t7AYLSwXgbW+1wlZL40GFCb/YQdJvpS+Z
ea5nOZo/nczVq23kuu5J6kb7nChTK1tDdZO4P1giDpOMr5Yk7AJhyvhskQNChpZbfmgO7VQFHqVG
ySfMxhr5KfVB7Z2bEAaONFY0LcsZ4gcp4w8ZWC6+6kNxyCSQ9d18xS+eAt22ynRtSWO+Rb9TEvsS
KQWqbIZEYmajdQSSvZyYItAmtseQbvmstk42PJ3yGFvhCXG1gtytFf5nWNurjJcsW4SIQk+iPw0O
Xqd/BjFSq/It3rrdMjcqzPH2aMAd2W/XFx8yTLOr5lC0prglbosEdO809fOUpTG4V89D4Ae1AR7u
S7CL9URfUp343/iDKT00wZSso60M371wGjVOsMzDCM1vv29UH4mMVRkOf7eVbXcLIWGzQ3Kd96Ih
a1/pJtsPpp5eJK4CI2dRf4VUIsyYq8DqAnwyYHR42q6jJ9V9g1E1lWWPTJN+axLrHdutHSs8eY1x
QkO1AaeFi5DbO6hlqGpkFimVuTIivDB/8+fBvS/4909jz0LjZESjECcbNDjBVhoxncjIKcmq4MMB
i33msDcP3BM9bivpr0Aaz38RGY4YDpnBISL3erv66SsEcXy6hcNuFl0s78aO3yKhJfu1AbYeOPq2
9BWu07NaS2F8ZOU9Z096aY9KCCHUTB901AeY4i5DVrYxW7s3jVTDrzJ0nUbRWFNVY5Id7yFnTva9
tJo9xUGiGU8m02ndQvEaTe+rVHLWaX8/nJ+OZI1y4vp8u4+9OwLCZr6CNkD9hUFd+9pt7kq8Hzrm
bddzfo0LMdPasy8Yp+C249ovOzjDRPIR0yr9zAyMO/KDxJtzbIQ+7DZiDbe1XjpCbDT9XrzraL6C
AYOxVITqcGfW5dWuzRnXFgaW+p6yZ+Gk3xBCHDVwSEy68MLOiN/Cqezucv7CKCC8A6pc3XIWqVnt
aIzHsQsbV1wKlZt1FFYEgucGRO1XIn9FayP/gSMY27BTjmAKrLEBZBTV0WII5TMZfFLH5TOXZggA
SvDfhwjfqBLa33DOZqVUz5Fun19zb8fC3DLDmaZrZ56kwBSlbntI4QcilRNAz9Ab6aIeaAcEj7am
O3zFQlNJvoP9Nti5JH5EKQBnWZ5WXtaXnQI3ersglU2rW4kMd5YyyePWk03H09NlwG6FdVcksKyM
1TRFotaJfpXPOXkqYh2beZc7hHLV4WN87bDeL3J6JD7Vy+oKWohvwvEKJw+0sjVFpZQ9cGW5IzOK
eo8SZ5n6KPsfuwMd5McSnvnWBV8tb8HPIPtzaLyHePGTmIgTa5NxmK3YrcGPaZ/gIV9anCj345Qf
nnfCaawVzma2EghxLMRjoBvWkQpUTquWjVAZi+uHSYIz3GpsruBHNJ9+4ZEnj+BYt0BHoVcmYbQF
FPQrjJScUzpsjvSS/UVyBr1dph8crB4jWP+/85YVUcbsWknSd6ei//3UlPmhlq1xWeWhfNKZZxNA
iKjzHKSBWrNMf2JaL8PJP4Gg/VdEuKgLwZ/M+dH5ZHPKflkHk7fcruVc8JX+dphbdpd0AQ/xXe65
7VhT/f5SyKbIpeWBHVu1zlR2C8DX23QyOqKKwP1Gx/S6pjzJFYl9/YghOS4jdxOlCo4F/sne31ko
TGHuFbGm8bma11pIBanVjJnMXoGY2ECkzr5izS5S7EvNID8WnAqalaU/uek1DXHcdNutImGThJ1R
Tf1ElI+xoTfE7PQ9/rHhA05CjwSf9h/Cn8w7ckmK3buulsAkYlUg7e0yZKM0aON8vrQRF/8Py5C1
b07dNQBeerpq0sK1G9pCMX9bgPVjBcCmOV7KOwXbBSPjfgZYOjEW4IalRgZHPlKsHQqNuINh/CBF
qtKlAtgEg4KA1mcX7gDQqSl2DeOiUxuZ3o9dUqazOGYxu+CylA5JAKRL9efUtZyqDojdcOHKIQD8
BhKMKHygOO/SrV9UgXT0s2vkMrhX0GSyxaLKG+GeB43845va7O9FEnqbMOU4n6FHvihROSlgabFH
RQkQQhQR7e6boi6ao6zQyWHn696/LPFzaEG+etppCQprDuIgFhXnN2DNE+B9U0B89JDyruf9Yu0d
kTEbiJPrnFOo1AQcq4jTNNrUngXAuSCkKZOY5tIq4x2HIYxpMlvgwJYsO/GaG0o0etMyST7HuXWi
n9pfh2QC1QZ69SG1johvCOboMqgHdv0jKAHF1wn74p3lnYFmUgexOpY/Ki4pg+HoHKcmceDsXtcm
8sueSvGfjFQ7Rf9IUIM9B8cpv4QjMx+63mfBJMx3uxon7/57JdLrDmLuKCwKSI8uw8AjTzwkosNG
Va816YrW9qo/aF0CU279aWXCnTjSTZU43Abg5Q6OSdVUfYB2oNMC0xw7jpBKCoYSJL1RNdAnXuK7
6cSEJVy4wmZFjnfjlHMuyHOMIJDv8zDH6We7EvEFvhXJVcxAava3L3207RG6AjEYTDaVaPCg/qBg
8pTwlfr/lzZLtfk0G+pjhkUU9fx9nD9a747KffiEO8c5M99RqDGd1qFDYq6F6Hqe82HI/YVoSkvK
LGP/BnXo7IkfdgFv3NU2wKdTRnwHpFdzfBcqoudJZwHmzFl3sZfz8LxeFe3gNJ3M2ew+ngcpb6Gj
tCFYDeYiftE+WkkCGyEahGpnxYp7QLMq3wksxuOUatABusWGYy0C6eCc+hvgk5RlTNIfljsQzVn0
J3IdcaL3xcJX0jkrJaXkzKM1021IzMiSiGb0pXNmWfw5n2jTmLevUJYByi7d0b+a2gIRwr4IDmzn
CCwDeleyRPjAnaISZoggql7os9d3R+vqYTu1MytPdVeLE1AZC9Q3ce0nCF/BXoEI6nzyGVTt5Kxm
QMjwvyKGNkDg7J3SoGRY7zNc9GT/uHRazsvjz1wenCmbRqVaz/WPmNju6D7L9zNKpvBgPJT0q3To
RJ/0B2N7a4uerE3JN7+NvNbwFK3X6y+P2NMcfzen/K1gjHHHuXu4vRk12b4kwZXKG6sR3v7tt2L3
+f4lem9tYz7jfGtmYokqytAJI13uO3FLfzuNxWD/X36t90OKeRDQBBuKpaOa5L4J4CBJkmyQ1ufn
aknZCdRyPudcQQTYCFF+X3N/0DLzFbSD6e19A6s1VHHR8tcFF9C2x7XqBIodkeGnDiKfk4r2C78Q
evTLmLoLN9oq5SmdMTEWBG32yKc2vynDwecn/zT/VROkxg9x2nNc2KGyRra6B3//gqVQybMedO6/
Hhu6bmEtkRqhrCOK/KmOwF4kYgDgBWJk1HAdNL3pE4oGcb+j/GxW0a5xpvNsl2Q4VyTeD1HMOYs8
0CQAg2QKBLjfVzpP8y+u9GXt4L30DKSszxiyh5Kp+ktYfAUeB5J6xIJaDRqMPwk9rcoQu9Ts73S3
lvbm0ZXUeRA0OBAov53kdUIontnmURBa7cAToeKfNrmWDHYbJ3/y3HbN+oBhwK3knjzyBnIsRUnm
HBNlHlixTcXDQIUHSgbayXaAa1XyEJlVnuxPsoxODIymK99TbUwYhZrCx1NmZhSMJ4VeeslXNE3A
/E29IgsvW/AsiLYgri+f6ykLrAITZH4LIGHrgQ70pyDkEhlg65nyHQRExcvOKdvVrwtN/5Kb3BCs
2mFR7Gm7qsumxSthJBpGkUHDO+JOCrJMgewv+utKmCBYesOntXja1xJfhrcrkq7cJq8rawGPgLmE
wlhxDQwS6rwhgQdkxByTSDsdlNz9LWk/WRq5M1T2xL1mx47cZPQX5o7vTdN0PexwkJ8Tewg3oaht
G0g9qBaMRZhH0e9hD8xvcP5X5pTvJEQbo79iRpM8GGFaa1If+3SMubY6pWUURe/qCWE2rBzlxeb2
XZ06LKHxPGPUehXGQvJEXJlTHkTVnDU0aY+9P/Zj8azRJtUwj9ju4e0JS3vKvcBLHeG+YvCZngWG
BY65K1KDFKabvQJlry4QdCGbZGagUseH9LFxG8OF++0bZZ3CAiRIe4luRzvWmWybnhyFxOYKEP3L
43Pa79vri1QL8/7CBGudFzuICgOG4ugitDV3MJ3i79qwCcr36wm0gBXVK4bUvHx/BNuxr5cWNbvo
9Y4a5tyyHp3RbpzieSGJyrEHyFwJ3zjT85UsoQ+zVlvtggroPb8ZZvyQYmZ+OcuB2Z3OS2YbdJVn
RIMKCA6NnHCL4lVgABTQdmYDMyehCmy7L4mVP3ulLnvdcTjGtBSkNwGAilp3JDrf9SO9FBUWk1bE
21Uk23CWGlXNU0yFuE/T0SWiLNaU56noEl4tJnkJhG0sLf6GeZ+bX70M9ggEJuXzvst7/SP76cRo
pQesyRionbIM0hihvSNwbnT3x9/rQBJRdYGrhpexgs1uHlFIOM3PmeJowaCY1N5SduDEIu8Vex7V
BOjKhEAikG1t6qIS3PX3EIagk9MXdb8TbIcMYjdENVQkNka7AEx7WkVzUjmTdSr22WBHl5SSVjmJ
Vs96e16neZt1AlYVHiJvtSyIlczGpf5QOuoa33y+9sYehQN+inz+tQN3PxS0W5wkc6TP2ktxjxp1
uKDOAYOfoYHZxt+og7PRCNF/o9gM+s1WjhDV3YlEz1nHMzyWbQTtAehAaQeR8Q1ZCq5akWhf1M7/
K2j0tWv110r4sI5W+XaN2FUTULUKFJooBwaqjHEryevP64HzyJL2GVxd4rohGhC8Bie8WD24tqO2
im2p1NbSYOqCkAHpnASJHSDKcnM/fQDRs2Bsh06TIthgSXgZC9BiWbyywC5p5ZIan7S5eyhBqSGi
fhYqlWtJD78wMVr1Lv+3+WZqBawRqYMr5qx1EMHbk+8d8ICXAPNe9IE1Ww9ZcyJ54bX0kPznRnFl
du0KRyvJFj6/ebqnnzYAC7P3K5lY3S+Gf3uWpCM0+SkOGrQdZeD9aheuljZUgmJwhbhSIH2A168Q
omGEfrshIeNqcrONKsoP9oaewIaZSq60fdXrb3U2d/rqfV1oKwgDEqEOv/wQz0cTBxAMcVKX5d3d
1NRT5jZRztU1wOG8tpQpimjGQcBC1VQo+4LiQolV8VbyEMn53IaybOMYaF4gqWWb9bHyEGmArEXQ
YnQBoiHFfNSXrad8SYb6q4M6UaRWdOc73QElZFo0yjuCg6s/AKbkYbmzpdyjxZe44aE5jgDGipLx
iy1p5hqpvjf8YUuFIF5unVy+D3mCBxBWeA6wcvX8MGYL9MjLwRqL4zyaZdHQnr5GZFvyqY+HRmkg
qIe6Pwu2sitXAgqvbBgv9uZ6BVD+MkVOtb3JO/P46tChtOtFmUO5Hn8WxYrjVpQo01qDcxwECufA
MV49rc7r4Vd6BcCFxHhErAx2g3wqNLLExU6a+ghQoKjTnNr4zp3oVMSrzlSU4W4ZR9jYiKVCuxXK
LdIG56gLtDysFUPtg4sZtIqOEY6uqjFyKHCCM6C55wGLoJ2BDa7L8Hw8pEDbSU6YsE91dKPiQTfK
HffdrpmtuHYp6u8HCpwymxDvua7S6oB11Cg/9V99Z1t+Wt9X/Cao6EETFPIzKzpR+j29wgi9p9Jr
l5gXRrwBtIrLbAUs1tMjcabKAJZO1dKmvv5a7RBEWTJi10TkYYwmAJr8VQ71FLiDYyqeSj4TMvcd
F+6xiQw8J8UUufy1JwTAoGX3EJEm1fQ80Bp7gH7s3Ixu5uW+gvLsuTJIj19bk0a9Gem6Tk3K2f6B
f2bP+8QK7rZrMC1kZHSYU+cK/ho9BmiM/rwCdHwz6XINsiW5cVU4aJRh1V7fqAeeJNkGdJ1c7a6+
8T3bANM8nOSVQZAq/AJZxyDRuRo4aDwJww2KWsRudmRzYH5D0I64MzaQDm4RVTVRaslXSoWDv0ZT
ZWIvXNWqIYi0p7ZWuLutnDZpUt/9p3Nb7/6iZqAZL2Yxo/zUcwzqYhOh6MSWVW3aTBVHVL2MnzB2
EQcP23HJ2DMYBWg7hwLXy1ZeYNBgXWO6aqSqGLRZgm2FM12m4ZESU7lBGLkb1KNZ4ECfsIhpEpY0
ZkTW2FH1OpgFgn1g3psPrU7WiPcmf/leLbZkkyx0rVF2ZeazE2sIDiW7tIyhe4x7EIB7F7Jec9FO
pdIhfsZPCdO6EegrQ/TOUk/101nHnlgowfUWEcmTgxvDVlBbedbvzi9QaT7shHuzU7Qje5DGsMfB
5qO379KKEmFACDOrfXkTFagHGoeSDDfcggNMFGC7B+9TJKZVG5SylKArT1M2d9pPl3TPkLlmGfCo
cncy4/v22P+0Vkb5BSLorSRq7oZBOnjnZ2EZvPvTZ62UYqup3BjvRcwm5cooXao4moTfw/gPtppv
avuDmSxGL1g9v0bd+Zxsl30Kb8T1Vpjb7dxcntv3xE2wpzmglN7dV3OWqTA92K714Bw2LxPEs8gD
mllEZE+5d697lLx/EEL2Lrpg3wJkCu00jAFxjE/XsgpIUTBNoqUjAFJIMOIM1QcDKQu9QR46W997
tqalmJfktGFurHFAcMO9f/DxhfIuK3GgAZD13xKAzO4XAIRMXi2vfjiPMXbjUmz/cV4AP1wiPYzb
TON8sojCjSNfZaXQW64nM4Xko/lqwGEgRD2mEN3SuV6i0QIu2hmeNDNC7KdHKip+CHFil6tA1yrr
QMPFSTZk7cOiTafjjX5Bx2ceJQNtJrQb7bUAx3LMUwWjn5mEMa2nQAU28zpZhfG/IqcVpBaTnvmo
LGz/Pa8/cGTnFoJ6t08dtrrsWSZ8xnjfz1j/taE3WcfTZUhnJlSPEKbyTJ/JYaH9YLHMP9iTrHZP
laoY9MTAmsafruW4BjoLNHkJCrWABmUOwqfk504grz3LyYyUsAzAiA2wbxaFhZTpEA4QinKRBM9n
JW3nHZHhJqFPKgRF/ugxjc0/BSga3334kVlQXuMSqU7CG88fW5suqnAtBHavUHw5FRAsIrhObiRI
/WnZ+Mw88qw5Hlc55z0NRgDy8W455SNCm9FvqSVpH2oOKmKNaIEqCQ1qMWckE0MNZGtngZGzBjrq
fuaTfdkazHTeeCunrWtrE/KCasUvzK3cE/2ezPuS4Z5uXCxZH3BnsYGhdUHLdZVmJV97ZyAlcuSp
MkCLKgAJ6LPgXbyc0Dn21IhoDvzdfWungk+7ngzwlaHRjnR9JOTCc8BOVBpI9FvMPqkaVwJutebc
7mSov43bUAZKZ5eL1gyqkmfB8J8wpaORKBj1GN9GtnsFgDwOKEsEBJFdLcvoPtqTOnpA0r70a3JA
GsEw0edCyR5NWyViYxuuLTOTuK75eJ4jEagLHwlmtvVdHORLUfMWwAbv/8yloQ0/kQGP3pw2pCOw
haBm9Ibl4mat45hG7bAfbMk497/l9pBhGBRbmJ/eIfggWPlEgimRn1rzUXQMDh6AbkUAPBe6djam
gIfrr/kulGAFceyw9oxnwwXWz7zQYVgwWEX7/RJPUvWm4MCCq2Ud0ep8GT9Rqj3Y0GjWWJm/GI/l
EObsmUp0tEW1vtYdPiBgJDJL5kIdM1egnIGutJhGN0fVqvgzKp6KuG749NAsXr1a71fgEcw+E0T0
nSpEkupmUkVIVwQ4Sq407iStBnFAy2dJxb8rikXdK66euJMuFmLASnJzr61Pv6lbzU2KXCFVp3F6
PUcCOGxwP24p3AsMnYIdubtdPbwEZrVk3aTF/8ErLxSGM4y1msZf9SKJ3gdsdenm5n+1JjRIUTV0
JjcxaQZmjNfS/+uBm8ss580viog7wIMfzeQ1hoYXHWeRxgianSe1SrSxLfCUBr6/t1aX8Ks4qeP9
GOeBmdFpw3f496gvC16FHgg+JXUGYyRcH5Z0nKts02LOul1QpVRMH0n4bE9UJFsNKd0bzYevFeo0
kAUs3J+SrfOZFzvEP1k1r74YlVEGPFPP2bJ/E+v2dLAsAQnNJEAi+NnLkLfEycYhN/buZdUaXrva
XE+weZ+wyTHe3+xCvOyMIq4WG5BKoKw8d6BVXDZqOWxWEVkYnW0ldMjxcFBA8kTS/prRE8+X0YVD
pUjC2OFsu0t7dhydzfMlJeIUv5IY/WFa8sj1W7vaU57q4LPfHKpZlZzLX1SqN9fmwJC/QUIByBw2
T+ogKnhA6nMUE02hmyHU5OZVZAfP7vZVXhDCdklk1sECRPPkjgFwxAGUHjlUkaSsajlcJNY4tiPd
b2SU9ZXL4eGQaIi4qhqUdKK/nuZ4n3AjvVcv8s100q7cBrgvQ7Sy54VBnt3Am2bwWssIoXinf8JQ
IAJhRq4JJcyQ1/KyC3PcGKHv0LaRmQqMdgyyG5qZAGDFno/P5JowaaEsNE7C8JPWrCjbmMh2AXuN
GBefARmBfZ5rOJkQYR/i7oLzQh8tcyL1VyljPovaFD4ca5/bfLy1HE0EWC5zTSdTGSMZwhsz6+yB
J/exMg7C2ASiW/MjzP3LWpvJq2o78HBLep4EkFLNgtXgrYqvQdFdcpJrDo5e3+dEn4x+IY6cLOyr
8BKhws4FPkbCMqDAMS04jAYVjfR/3ABuckSamh+/mIZFbkwhDUJ8Pk/ZKNe2pafHFNnZx60wwbrB
y5vpSjfjzKuFsj2ccW55NNtonmNSie1msGDk4NX/Asr3IAZgfOJpZPajx0UGK/aFZqavxjgSf8CD
E5WySCnCR8flF58vZ9+e3EwDpGkYbHajiXeLUvMV5HgZh8ap6NgBsh4fl8f5wrxG17HvuPy1Fsmm
9Y9WTQDG53XpERCFQ/KQyN0gncT2D92Cevjdl5D8Q+MyniXBIsKHmEhNcsbe9qO2vle7vnsfP+3y
usT/en3TIFJy5q9Fs+ZbLDzz+N1pRmZg/2PNXNsL2peysN9P5XwoFWNeLVEYEMf9POo23mRmQIxu
9JFYrLmFaZlDMEc22kRqA2t1p8PckL4wOPXMK/8rT9BXU+N5HLssGZQfr1lLSdRtQU9ARDTcjGkb
WD5ds1yNQUtCgNjc45CDVqxjKZ5z2eSl1G9qMRwmfASY/vQHg26YIHC2UB/xdR3dLHwjVFmf8oKf
t7F36zGnYtr8qO6tpGYaFuby9+A1DK7BFsOsauKVRYZON3v+Xf9s9WadrfX5JTrkQ6vwlY1E/nGG
Z2Z/RVbzYjao7jcg8etX5/BM1TB1yvPvUSTcwgTgbETLLOEMAXMkwRT7pveBYPdF8uNtI+fX5Ziz
0tbi+xqE01HsCqQogMVLFx/M+tJDVaLYSrtnA2DVTxyXxjvTYzq3B3pnsvDMthUBzc3WkZ79pcfn
i07a1K6zGc/zxCqgztbUtumbfuvyUfX/9vOV1rBxV871aBnciGpMPpbvHa+c0cxvN3ibCIln/FPC
ZhkOjVKAi21ItOskEAy8fj5Oy2qufvwLvWYviiDgaYck9kbzcAQeMhWmQKi4dlPqmQruv7JRmAYv
EFcdie4/fq0xDw/bJ3oBMNZZVai8fdOsll6+zkLKx9cYlyOH5kLlidWDwLGZhTnUkQQl0avjK8ra
MNYC4h9oGEiqJGZPHKJgpeIXMev1d49K+n6z/KwWT7W7MRyxBDO8hGEZvDu6RQJepL+Vo1UNbP0k
o5cN2yc2cgCyG7J8zbYejv+3fU0KiMdJuXXZkKgprztEH40gvfq+2tftaCEvmq1PxLoHJGV8K0M+
x27cO4kztiK0hBMhjh15tiz3MDY9F/R4uZpB1ZtQVHuzK4Sc31bHxTij4FhhEbn6UgAoSlRrKiFZ
a6BhElp/1jwIdmTocm9qPAZFWbO2hEMfYJpQk96whYvRthvUkxK+git7SJh6qD+l5sKwqgkXwI0u
uN0Od80NjuZt2uq+gG3ekmenS0lctPOQUJQHx/bLeHxPJVacoDxfqSUkfEvfAwXZyF1DwJeIam0A
NdjhuG5+9rtmuoieI6dm8MKVTIT20dy002W0y5qtOYUPU11smQOvz3mjZdpHT28BDRAVLU7ISCRG
yLZnO6/waHdca3ihzV5A/OpZKfnKsn3pu9IyXn5FbmEVuan6xIM8BIxhkFMFlgt6ptT4XYNdYtLR
OfkIS2A5SYi7PYeBi/EWDemIlRd1s/qY5+PZLa8NdWxJmqdCYHlNF6K/wp1eMZtUm3vduuzDTwwj
eOzZj5xfseA770MMYRTf5oJ7zw4x/bjno94fJ1nbQFfm9oNlj5QybibbhkFl6NBkUhtKYUvCczNT
22PYz46JmtOOJjFmt04/Xl1NVY4T2AtRWMPOqeVdtOMIq0D8N2t4YSf/OgXlTEVZy2aXLXFM2ZYU
pkWwlE+ngSx4FsCn4DrA4kdLurS1PA2seyC3erhyt8H5noEUGwFIoMfqIBTPcTQqNifhPd2I3xYF
TwteA2oQF6Rt/O6ej+dTpsSxbkZoqnweHCynsGV0XwZsEK8z9uYjGuvPczjHTKKgPAOf3yN70zEM
f6LlqX85YV8vWuWCl5h2PSR1f/ZdiVBY5j7oiC/6X9QzyILvB9NmfOyCQUm41jBVIaQd9zoPLVP5
Ek1vHfPdE0yAuaOtSIqYsvM7hBglmenfNtXluK0IWIfWS2JnBFf9OtPuypI0XM1ZHFqvxcG3qI+z
UveCo8N8/GcVP/wIWYAlwn324CAgkBJ/YPddRrkY6VNVYnBgFJuyY8/YUYqPTUBSMuZLlHI3g04l
qF2tPk6WrRni07d7wmDYHOgUvCof4CxVrHo1aVi3dRb/ATkIiYAq9TsTjiyl0i2Yiw9KrMQXd38y
+xZH/G/b0YveEOn5vEXMgAuPnBbZ9A7KNG0nte5pLMVDFgYVAxy8r6aQxVAfUQjuhcs/lbGsQThm
IFnlkUzRiDAbReyVLJfkssEzRPMZe2epuc3OglsmLSpzA2pF4DYm/dDO+nIH/RW4k+R1WaXHNiof
GT1S55Pt9EsFKXSK6OxYTsvk0hOawPsmS2jJ3wVAye+r8CoE5DZdxkzwtzg3GX6BW3w9/3VDQfkK
fDABBVv91evM5mjrnL0+M9yb+fcjOXxZkcUZxthdkRD2CuwkIq0v3eCAjxkJ9MmCZ6mk0NBl4R4x
wJM6100WVLM57kKT+ZgmGFWyjnFGc25fdIkd53FOAL6v65wWyTFgLoW3i5mOVtz/qYDu/hCyIPsF
g5UzERh7XfTKAA9hiWUrNanuyAXT/pkgFyMxjTp/+KwWTveKAO4QST6vQhRwBZeIvwA1RHRhXVUy
I1pKE7GvA2dFtl/4Jjhb8bJ8XhacbbBVmDsVX4veJ+7PqZowKhcujCrzbG5fuEnH+j6CQHTNFwd4
v4SwwvyXkqW6jCI0O4Wyn/KDgor3iaehF2REtvA4RoPfNFOQ1KrytRrVOGASYEGOvEceiVkw82Sf
pxvuWbSDNarGwK2/ePk4oTL4jPPXUkQG4s66Q76gKVI8a6m8UIh4oo6LJG2ZrTj3joXtIbW8GZYO
tDoudwg6sHH08ta5qT7JBC+46kWPaxO06KEKee76RwxI7sun/WcadBSvLIPaB7WEdyPG8Bpau3vC
5tGYxde1w4FEF/UMerYy9jhuAJg1SRmtBEEK3bheyNPiEO3/YoCUtg1CccEaPZUV/YMoN9TMZZiu
riUHWq8hIyu5oqqnb88MN3gBE/k9Q4jG7IvT0FE4cD5evXuHTMWFbc1/Ff1daCf6+3RcRmZzTKoh
+gxwgNFOXfS1QYxKLEgwH2Ap0GId4mXvta9hmP2303PNZuyzQP9BnVoehGR3nfpdZyliK8Zq05jO
ZQ4twPD/LbL46u7Gd/1w2EMrJPpdfWeVs5yOblRRBmTbw+aaWcoSRxwfz6ppX9QRnpLt12laD9NC
TD1uVaIbZqj0FcKUnMl6pglqJChJFR9N3NB+oHeWkiUexY4YXE2OWuYVTcRwbISIr+/tLFt1m05A
CpvWl/bVURNN2l+hKiG0Hwnq1hfNnaCe5Gvn6QYb/V0JJjM/dJd38omyh0ol7CqxPxCRnOdg3ADJ
jgKF9dCt/3JNkmY33IJYVMJMQyUS1ePQLmhmnRSSLOGb12jhoRfn0AK3PEH07uPE9Ir94/aocdMy
lRKXU2mWvQ4vmKIUva77ZMxtBD6jqBbq4Hu8bFm0Q/OjA0OkE2O2tmrF5LRGtv1iRl8AofW4ZNHh
I83oM0oIW+8EZFjYZwOfzr6mKxL46lDUWosx2wieCh7p1kQVIm9ZjGeiZFfOYWg9N4cIKvdjSqMb
8n7Zlm2YCa4aMP5JnheyG9Dl5bBsaAGrLYdXLIsWTQPGGM5CMfOgE3D9UlrzDhii9RBdKVM4+fG7
hW+i5n0FngrQ1Be1PeUkJlh/+x86FblZM5PkLBhz9h2k6cTe1/muCl058OYWfqQ1X3U7tfdJfXXk
XdEPqbUhlYC8TcMicZ1L2SOU3DgkG2JHPH/epCERVv9hEuEkifb+6/uA5pWnTJO8VtkcQ+hSXASf
bcao5vltcg+eHOiVM1fIFQJYXr1PNzHl7zpvSoN6gY3ilF+JxL97ADwBvhh5L1LLF5pT2PUdfcRd
JW+WCl7b96nGls93JcV+U0+owUu7lICmUSvxQNztpo095OxEDmguu1ZPc08yU4qs2Dfvowv5SyM0
laaKcgeftKFS8WiQAZHL0i0LUalEvSfTdFac7U6TL168dmvFix4FP8SyAhfBHMMiWGl53R4actPv
vnu+gMeBWiptfSRzHdJQ85qvOv0huWzv4cUutpGULTpnl9t22OSHgrPppyXxW5AFCgzU2jm6K0Dd
aZat8hWdR2qHGT7si1tqYxEa1cxwdcuFLEcfBrQ6zcqZet+1+dEdTo5ELhAXfXgvUZfpFWIyIE/0
5BCbzGOJByeyWT5QIjfNZvKJ30YDh+DTjKYx/Tj98W+pi4tpyNQ1qlqyKLAG7iScjTQW1qK3VcuD
Y2rjMSl0bp754Fn5VxqzOYFWlBqRLyizYo3JbI3NX7wonwK6Cij9CuZneC/2KCO2wk6T7Q0tGU38
6wY3efTE1tWOCkus08DI9uov0dC72xOkCXLfc7w9ULoKyybZ9+37BrQyJWQxHTQh9hLc+194bMTL
zFdp5CS7lyFGXYOf0UW4isq/40x19WIumDAWUBLWzXWuGRbfbbn/6/Gecz/wG8sEu9gTDP/9GJF9
ybITKplOqkF3XlvnjBgBpSpGDoedfJVIPWg0gkxeIpmOVw1qL4Wvs6LKvlmCWo2xLgMkn2o9+Tye
E4t4DMZyj7LQv3evgkc36TJW+BmcPdC8XvsnesYDjxW53gS7rmiDm6qV4q1X52k1UWhTDxMV/asf
mT99824vCfHYhqkrjIX4NYVPML7JfAwVbSp8LwQ+rXudQiYlBtQVBarPFNWD/tS2jvVMZAqxNhuU
WEHHGdPvQjmU8/Y4nK1ccWY1POy7ii8N7MvnP4sBhrJuysDVmGcxoWF8ctUA2wUe3jb7m0pRaumg
h7M7f/E/eKRmA9xNn8gDu8yv6S2pu8uhZXY6GwioQMhF/D4EKhJ8AGL7gjKwE6iCC6pzjkLZ+wEU
A2YXa/LHUjeyOZ1oMzOFri4vrKAGkQlmyhb657iSUGG/6vxJ4DN5soRaDycN+Wj50Ld3zJS920xb
77NjFGA++64BKtvLOhrw8BCNkChd6nPAbZNde7XkyYtwwSWCNGlLFtSZ9qI/HVlmA7ZPUhDBMQh2
THDWItEBPS+AcZHfQ5LPG2XZV6XnfhPcdPWz6ar3Q4DebL5+R59suRktZDmrEvlbJee66PCi2J6z
/OdFKospVdrMJPzN8iPEul3ciPSMwdBOXJGULjDM9K5uNqTiFMdSHsYCj4s7fUGPHrF9/vvk1Kou
T8RLUWyLR+SzBFoSV+DvxQGKr9KHH5svkKHI17+rO45PDBp+thWJ36aeLNU2GP9j7wM4mq0V4Hid
BtAHV5PgNglwFEymlyq3S/q/89s8t0mKnjP/cvH9T+h5T2iGqRBboU7zRo6fl2xarTq+WLQYVifi
7GKAqsnBjnXWrqefVkTyb83I+zwIFZUGMUH7BzTBuYVn+EnQoLnGJiJ7ah8xNmTexFByPACzv8Ad
el+nfS4TqzHemjLKzGp3zoZFEfjSHiaDFFWKxkei47AG5M8MQ9s+uXX0UswdDcrDJ7a5O+uxbJpj
LdaPkats3zpzDJ7wTjQU6/xTGQJbJH5kalqUI5GHGXs44H6RT0GvwXDvlMOVY94mTJa8kj0TFNiq
mcYU82C6nA6XYPMYWSJ3I/sEhGHcGG2cL+4uOUSPw2HkFmemFLnu9GFIVdej+UnPOxTKW9hzeVVz
Mum27+ZGxkGe4mh0qYM6U/cWWorcOphS7o7sTNYYxGHbWMQd9YWcq4yiG7IL1O7KFM2SzDjj5vfc
/LZlyopAxPz9AidDE3x/SrcrUSgzZ8tZztJedA2eBMdlmyttGOdqmiVf5tGWAYwlfKuq6VX6qJiM
QTzlX+LcIhWhB2w/D+hD//rejtjvBAGE1O2VLmIuM10fU1le+gdHk59bf373obh/e94lZQ62/67h
C3ob8BTDq53bYKuQO17/eDvvl15NZkLb0FccY3fpgeUFF58MiCBHH3KHBq5eoDZtHCVwyIZPS/tt
735Mi0bB3SfMZKryc7ImTVMKLfVJAhkjIzG4MrN5F4zYgGbZGZdTEBzb5Ifs1+QKnuUUSRdPRfh6
e7ChJY504JHUYbKgFdHsHVaAPk0SmPKfgVWQBSV2YctHtzPEYhPc3CZt6IA6Uem5P2nGeEVOnui1
I0mJ3GuOv0sQXtGoRlVasR/11372KtmfmP75GkemZnqGYlfiTqUnebWy9MEbBvCk0/75k85nFs8Z
N8JibcaFgMxrfwtlzz92i8T5EK5NwyvYx/oXT6Yvqg6++fKoOKhSGTAvOhSP00tYUm/Cw3n3h0Bd
hQQt9KhbThm2YZSPfVht7s0eNCotHnTCZlUUjn1AN6xe2/xTWgDx6lz9rbY9vdJr8BtGHarNwNma
cmRJTq4idzG3nFxxXWgS7GPAsXzdvEbRXiqa+WwGZRRHEeZGHbqvEtTwZTI0NszzGEGIMGVQEArN
Ef5po8nJF2QHzMp6gSkobwcS76WqfDKAl1lSfaXwl1/Rpml0Cu8Fn/RI63F4jAztbfXNv4suaxai
YBGTwtsfFIYjcnRUorC/6o1+yT5uoVwl5hpKSOHOVlcSGOULNCa97hYEfLE2jk+QNpuBZEiIk3KD
cbyUzkyLkTTF4TGwE+phXV1PmpxnJ3eTPRfFYkyud1lQT9aVu2rEokuBmzYoK3RlHcyR5B4hay5o
gI+q44FDhxdnxHlnOsQH3munud5o1/U9Kg0/BlhiqZcclW2lpRfL99tM5YLditu8XCBtwSO1loyu
ysDRz4Npbe9b8yLUFthRwuHrW3gGhyPYx8De5d+PCWlbU8mGDaXJnL1aW788invbaluqs31qCSPL
zVTIOcz2G2DltW7Sw0HSpdLrKVfeVF2oDRmc4afwTWZfmwqbKjmRmf9y9g4kgq+1c18SSPiIBY0X
VV69Uk4wEr3via1sgN0wTtK2LY2oC9CLKDUslZvtjPlXxKm8hueblJjFOMOWUhuJipbhd3YxFx+u
lEk6Dg14ZguJ9jtT0SBjZIMTNqgs7qOM/KnrsnY2hZjRFV7hHwpIiIbMXQY9rfHsSTbo9z0SemJ6
G6ubuYU3FMNqaAUv5CfFlZZY8gVcB9JSTZ477Yl7NwOyFIMEHUriakmWIEWtCyOOnq2EUED7N4wc
v6qoVm7gMTPCCyOsDccy0BvFP/98Ax1idLXmGkQLkbpUlQNWN2605vlau3/3tKiAEDc2ZTg6XOx5
9AfyjeQLrv1WIpd8UJsoBiV1XNqC0bxCsynkqC/7qpcr6zwTUis8e6h+Ut2bMft89oEo2he4KqGy
aRxRYLioKrERUQkT9BxJTobZBsFLO5rpwOHJSyOjVyXLqEm4jLBtlSfhMHAZitctn1x8CmfsxrbX
VvHTMl2GJBucM8YxtbWFXI20D6qtdNvzwZwm5558qbRO/rMn/cVaKUy4ImT8pD/RBH6+/8dT4ABH
tOaWHiVgwVwjf5DebVI+fyubvok3Ck8ibcH7ye449KAu0+bwFNaQSA0baX3mLxus8IT5g1rq4sU5
cif2jS+lxlvbkoixs2seknyGRnLByGvhuzujr5Z4KHNjpbQ6e7dHyM4hC3KACFIQiamTYmi3KLqA
sdkoj4n9Lg1lypdLl7cSdH9a9+NZgUNTmfjUnyxPn7FoMY7WKZHVM9nN6JWvNTRVQWANrzXOuxi4
KfspyTokFRoVY7JEIiV995ScBLqkObgCbzDJhMDNMcPycwSZP2133rSh6naUDzkNcE89QSd3V7tR
1YtkFI+JmJCCqEvKJQk40H7bZZdteD4xY1vb6Wijt9+VVVjU5KOI09G8AvU4ThUQtGtBIHLTV8C6
/Vzcg1a9YHAGe7wFMkIy5P8ZrZA8IRBQG5e3SjgQTD8gD7VS8wWW3LnRigGRLMJ7dbOOgaukWRKa
kw65ES6pNnolF4bEmhYJLdIGgqXA4aYGA2geS66FnSWjeP0chAW4oqkY7ydjFZ3UIy/nMzZ1y7GT
7fUlQD6kimFO07cLBUbvSN5x4oFWd45A5dfnHe/KBn/Z/xRKZ/bsR1UbB6BCuPpRu0tmpkEIK/zD
BY8sxYXmpK3fPq8ZLy1nKi0m6jIq3NgqIiRZ4dc4IiQOs4yb5fCmPFwgJOgz+WcJrdEfgjnngpd9
PW9oRCFnLnBT4eyXuV3xgF0dgyMBrbOUsaH2SLw4p+NvbWe2U1BJCYgL06DTSUIyCnWcwPKtN+nP
C257QmQauhqNtWeUNPJP2A3ZEvyu4Pu6ioVzbNtrHdnHU4A2wSOyCdeuRI61pVNPpbE5dFs6Bepv
eZ8JN+LsjmUiT09e8pRI5vT0yugPQcmGLPb4ez/Yy6LdBd3uLEbxmAAAGYTYdRyXCrVrxhNmJsnC
g6PJf3Nfzbupp7lvZfDJiq3F9kd0wplKfQ3yQBngl3wOf9x+zNF4XgYdXZ5rw/ACztA4IWPL/dE5
RPKemQY0pfqqau8pm830zlPobj0SbpSN9x+I2B+0b/6/SC8MwPT1zRthi2oSn2NkVLhR2gPfNbmJ
O/4pa0RXSPe8cIcIe0yJFoz9OHbTTkMnYGGj2b0qFzs+/FAuxZUyykmGioo0GfAIXTup+QAFQYgQ
UT0hO3BKmYivp/Hy40eL7zrODu9nKqjRQ+7hSXFjTazSi3DLGXUSwciR78/Pm8SaMbPT6zzJ9k14
M7UXckijG/guTtVhzfR8SCRvL/BiUGp6K3gQTMqzoAdHI8QV1lEBWMybUtmin63Tj2HPWic+hcxH
iIN1zIKh1G0AQY1bs/w7ksfk8UCWnUXXdzHhwCQ8bpyV60SpC9MgtTrcIh87totesqbxVQoo/B5a
jMGL0JkPom2IfbkAM6C1p6od8Nv7F1f/goD2dfPKXT2GTZiTYj63tImNOzNrdae40WtibD65FPfQ
mMQVJ6RJMbdZpcUXnGXKzAFKU+ZfMIP/sabeh9y1TB9wlntgwYh3fup0GL82hmZMcIsDo0ZPvDH0
QspdV8rGqZ3pX6AMvxLO0g2oApZhGSUeQO5yY7blOKp/xhQ4W9SNOG112yKuMIgp6Ft2Ecnm5Dpo
Su3X9GQcsVyJ/xvjygtZMXHF1NXDXfNReFHAAA+aCYexbd8X2OZeAw5wedGeUZfdn1/ZFgfequpj
w3xaGPhsqnLnSaPdGPMxbshnSsOGcxVq+VL03+ic5PUpDm3Hxreun350EjEmvq4wVXkJIsDcKbVo
xbH617G4aCEg4tGJSzN4FX3O/lgrpKzXnBLv6l5kzIRf/OAXaJQ+HRPtJHexq9pCyLVn2jtqXS9G
Lwe6lwm3ExDM2z9IQp62gJQjdyBS2o0hh5u4nKeITa0k41U+aeh/St4P53XRpJyAoqLBwRN+xe1R
DSVTnSSshJv5nPwU1n9ibvr7u2REkzXzFiYHhPRU2/eQamjB1A6krarlxYf1HbX7e46iq2m8f0lD
Dn+pOz+J7locrX5UX5y0KBFDAnAIw1h06cIWzmVq5V5380OgUub4dY+RwPpW/SzdFuU/nWrgTwkA
V2+URvGHsSdydAomEi5q2Z4FrGfDJKt/RKsu3E0SoLvTXKGXdzLGY/nCOt8+DH7hmGztzykXCcwT
IejoYAUAMk6nhy5BGTDX3IrEGPW5ysqcVTYyB2gcN/czgWNLGEVy99nCzCzG8XOusU6Zq8Dg4OGP
3Y5wpphgSDBIoIHEI2JvcvFHQfvoZ5DJANEk+UswfFXutjiRAsg8N22HsRidLnvRu+3swWHCebm5
NCaDPxA0XGUvi6TfD46QWZbCTvzcTjxybIuL0QMkm0eboMHYeGnnrhuoCulTfyzjQ6oykL0JlC0F
lwlQ8XCQ/F0MVWRJXShhbES9BnNk3yTU5OUq0XvD09p69fMqOc1XlOeF4IbKiG0zrBsaE9FVcMAb
FDESlbOX76P7vAui6pBmA1f82U/+/cLJ8ZrOI4PZR0rUApiTEEqd3fuOIVomWSjbI5T78JFG9ZzX
pKWDlNCyCoE3F6J/cyOdZawbEvA0M3FDX4/ZX99Dz4dt95m6eVkFqSxQVQO+3zTcMGjYICQ48a2F
vlpyjXFkFSjOoS7PlUJp7+tOW2UL9XObkk0Pc5FU8NPznPpwp5Et1O7+UYUrJbSQv+FV2GNysGXe
cFhzPF5ehoJ/xfLl67MbvfowjGgqOtPEQo+3ydE1j0W3JGsxIk7Ey3JJmWaIQghD8jSdGAPEfg17
aHe11utLqTaXsEeLGr6nCLbFArP2yyxZ3idPTjyleBzCoh8s901+CEWeW+REWfr7nQKi8Z07fLZL
IRcMc0efx/I8LIRZLXO8isL/TeN3iS8681be9n57URiz0tn/k0c9pN+K2G0ATapERkVOH4zEukNZ
F1qDWHOv7dA6xIBkNYc/gMxmvPshPKn12NO0yMY6PEJtTdchII/NlartKg1+gEAQ9TIFKIUVxCq3
vkF/dyTe1BD93Bmdozm653d5s0zjjtwEHgMwOKBs9T3qLa5UMluEtB3jTHh8ISPIE1RObX6mRyV5
+rY5n0A6hijL5EgqLM49uK9Up2wlLRHVbnHufutxYzLOi2tgHyzgzue9e8N7DaVaB7EQrJfdNNJ4
2ftv7J2GHbzykdmk7KAvzx7CvwdbzOBfEAMDzw65tTX2NxsDUu3mqWODu9aEbfPYRzNfLcXGUQbK
4BajBrJFvJRwOt3uDRgW2WE0lUPGqAZ9nn2aBZwBgqpELBd4FjjTw9QlQt91JseMWMP5/uGomrPe
y7GN3RT/n6MCovGKvZDN3n36dsmUwGi/ckE4KO5cDpP4El2VFwbLuJcCTvha1CKm2jNW6Kddiid/
yS+cey9/Hmb1EFfiXIMK+9byDQo747UhEl3Bbcgh910e0AYQNwr09ZPNy82KXagvnoofV5ArU3av
5iPvl7g13UCUHwTrIGLd41s4R7IxRkQ+3kcpNXtpy9ekjTJmGaLb+WZGPhRGIf7FUpDLx3ESIrKP
vvHoAsCOZQPDhTTLvhSgw/WXh0r3nhZdCyHdVnwmWjILcKtcl0OIJtROLnmWVNilKr1TtmU9iNyn
F7ZusWY/CLOFco/vZtck8UnBG6si7DHJ8rl92J4Omx1nxgfIpv7YFBp7+OZA0I2K6yftiNahB9uu
oWu+UwZoMNXn3ReQdhWVTJPnU+Hox/DKRBkXAywAlUIyrcR/Buh7nxpe57Bu1Q72w/SJqHvarnbT
p/tmHkqP6YYN6QlXvvj4JuJEBBEkIkFX/C7UEhVDgnrAqbRQXQBLdF1z4VRM6vzRl/THu5aZALpC
72Z5nCCglsHcyLoBa7IIIsI+CrkLt2E2K9AZXJl6ZrR6wwI0U+vzR6Qh3Bu3BPhDHA99qJCOiHfs
70QMDsovpgTYvwFaYE+9VhgKHUgUriD9tYk/eWCV/xIY4C/QAVGI/3gWkuZ6OXblMmuaf6ccNcSM
ZAzHZ0cUmhmt8kWTfGbQoTVTEhtX3qD6oxAgkHWTUVS822U7DCmhhapaTWoZmDhQoqIZ/d4tFyzQ
FmMK8x+J54wCzmX6zAkQ6i0LhO2qZUrKXxigjFXn/IADBviPHizqetvspHl75t/+YL0xlT/h1sOq
CmwPR3N4luKMAc1mr25+91t/poXYLXgUpXL5GjsAwP5s+QIz5tuFPJoUVP6H++L5OU9mPL+NTX96
p0AMycff4r86T6kcsvanIW3VWxB0UnnCuvQKlUf8C96xZDY+lzDAK5I4jfAx7yhH6bKgHbsDYyXZ
stPalZK7cyhuJSfnpxzghp5JyrXFlhUGe7MX9/TE+LMQF0nx2kS7pcJi9t40UmKxmjdlHyjEZDUs
4KT9EvUahaNo+NTkZiRK+TvjRb9sEL62Shp7V4eqkLuqjfcG12uny75KOzxPY+/z1Phcvua+Ctm0
ku7ZRCJdXhRt9Lugx4xTO0yJ1FxUVvytSMTpC9ERPVCBwIsRVAfG8EOeueo5807HZjjlqZsud1eZ
pWGqni1v2xgV2ab9JCQHI2wF5ptoYLLsw2zCZMosPAl2osbmfwNL6XgBBbxZHJPdIkk2hoNENQns
jZyIQ3gPKSa/uM0ko2G21EiGr3Dg0WeW7yE4/+QXLqBTMQoYZt9hbm1x/iS+OwBV5X0xlyQh1JqH
QSDGaN+5WhJe4OLFSKKdAGK1lqPJZ58V7BlJl+PN9EFEd87X8XHDVKvRkG1TzR7aE/+FhEYKzuZ+
jLINbX+zxV93olkXl3J/m7rUeRTv9o+ib/Qpd8+QC6iwuwBWHG6pbMqcw8N3TG8lJSCbKuQjlsZB
+HceEHKOqjEKEV97N/5zHw97WKiI05ojP0ZddklMLrrwDBykV0cykn7NxZe7behJQdmluNtKyEmj
vcrtvTmNFVxvIfSnDOCZlIUdo+C6S664bg3IN9yUmOdLbl8VGOuTd0gJfEqVC651qbBM2lsU/lTa
ypkG1nj38Ynjp7qc2G0QX2z65ro4jVFIKYrcYF0LWzo6Q6qHFMDCHX9aQ4C/ianGESVZErpEUuRP
sxpvhDPsWJT9Sm3ryu1y00x/AOJtgT2D7GGrEbFVeZkehxmWa3hAc/L1Srivgj0Tu2MpYJvFSHE+
33drRVj3izn3MHNpFhHFPg16xRqBY7Ql8S+c5cQgesSc9C8BbL1PKxpCsoDahYU6RRL34tO1CtNK
3cE+hWDdSwMs20ZTMlcEaCNXqpMnGvg2ixpHcSnqwaJhUocCeiY0phg2SVC6G8T5tdl2mAmpz6JB
XLGB7Ps0fSp4B6RdoZ/HqphXnc88cjpsfxQ41qWj8WkINCIvIk5u9FUpOIxu7YAX7vTeV53EKOvj
ZcLLxOVYfbwdEm/chLZgNiQVRlqknsSSCTM3VevBLxCjGQ0mWhUt+mkVU5mkoFSCMFwi6sqCx3Xd
xv08pgRiQhOaVD2y5C8K8NkRe/T62WRYZhepeosXTranimYaer2UdrpTsYOdVWnUvdTd9DJ4ZgVH
OgEcJ3KfHCrC6UZrBJ74FDoIcdTpib7qiRr1Bna5wZCB6WwL3b1RyZLmrOMhzMUYh3z+hX32P1fr
2waOAHHv05grRhW8KSELXBBgfwc/Q3kctjkS0VxH8HM2wRA7lBhgyFt/I/n0E1LAlfE3kdCWxpei
ebp9jqsBrgM6Uqb6PFFHTZNyMN4Z2kiWwqylvubhjPZsEeA3I3uYPRV3+1MERORYyWCepXuoRaAm
uOfmgZ4ydZrbaBFEx2MG8uRy6ZAjDuv7R4o1UKqQ8Umfb5wAn9QfoVLTwv0pHIVlU8w1VdhzNp3b
9giNgz6gUDhlc12TVw9LfcBRkA5m/CTlrS2jJxe/qAP6CEQH/1f2O5nWEWe9o0eAETFs0baUimZx
8jnfDsOGraD8BEHMFOx5BFqdaWJf/1PD9X4L+DPE1Hs1NXQVunMmgnAp4j66jNHKfON1U8GamzLv
1JME47fNRReG5EgQGCutOXrlVlWrbHH/KSONJLJ0Fe5xvG6N1Ih9m2LRP5fF4ca0oQjM+06tA/Ps
RcYbTpTP7WJI3taWayb/NZjHv9dTPsuZXsL44Dg/Ow3ZmhOYXSa+Kn16YDVPV0BSlIv/P3I+smIq
pmt5DKLwKLJnTEbO3CqMQmDfFrEXZD7RVt424+p9E14nauxmzlQbO2P0tZ53kHQpmC6mPnyCqefR
Mu16W80rlDJm5nQO4ZWuRRTKpbn6sCZ1HzVM8TM+2CUxU+nivStsV1RB1C1mBCqbMkpmo0R1otTc
GghSdDIKZzv2mn2PSAtOoVEeyZcwq+kJtfCyo46cxpJB0BR4tHMXxoCDNTe1jLL7eX3q14UX/k3f
7OED9mrEYCtsjvRMrZJAb/ZdVS0bQtC/Upm4D2zxmEJzhQ7smBVU+eJ+SFshLB84WPFj22hLX6Mg
lYLAzATMrmwovSjOJx9qGsyuvobdapgwWkRXqNPIfKzaFKDXlUdGp0ZJ6aNaHG/dX4eA/E7LJfJL
Nd62/77HKUgENTvh9Xg9aOUI0fBPI+6fQYtvOweULhcLLFMt7SY09LFfd/btEGlM2XdzxCNg/2tK
E5UiO9IRzuOpFhjRQ3wQN2gqtsHWI4oRPYdJnpvCHhBqzQVpjwoSixtM/kWfxcwP032HeBRQ6Pi4
9/69FDb840FR/NNnFCDX2oPU5lqZ7/W1s/0yTGF6sJTK/a25fvwIAxZ2YAaiv2KdlTh5+/pc+sZt
jRrBtkkhbjM/eVV78ZmuaPRnIEHOUPfJFdS+uIBaO1SzOonJ6fxMJXOUQAyzAA8pxJ4p0RtpnvRW
B7XwF/uCHnPkPkXnwIkuQC63ugVhHj+A7JG7/x7Yis0nejIau1SZAhr+Di4U6/g+PGVU8OVv2SB5
TKuZ3ew410IcYZxBIzTcUb5iJ2MlFd2TfGQ05qwrt0ma3JREzgEVcjE6eDjG/vmHLJmTE5dbj4FG
z89Orknbr3HpDQ/VqEuq+1MXFNNMdqpZsUpxq8Gh7sev9MrjKWqOT6KQ8YcTR/4IVCuVNSV2Lo3O
0C0rxrRdmaq/o62xfnotJ5kk1fFxmhRL/tWmGILIZ45Z3lKCKmEyC6CfF0jY85D/3bAJ1aBjW3B+
kQkZoGXW7na6Kxrlbm78Pz3gsCOawgPrlBEcSc3rQVtmDIyqm/Tp1oe3cCG//g5swcYFCNIQU8t/
U7RZXtvdGHCCsA85CMbLlTEtgTIyNG4F3oYYSWC9CaOxEqo418yKAmBBqsQcHnt5Tni8QyovfVgb
FtaTi24F2G4Fp/z41Rqs/wOqgo4VYuEYLoa7wtvMp8zVtAf/73LjE0EKst4nN9RQQXvY/kQ4obuZ
/nrQw73tlaTc0mOF77N3hY8jgYLrTUQ7cNJK253jv2I+dAMbkEGz78wQa1hp7oQmh+FKvt/Xh85p
eT3ZlhG0NTdX/x3gmz8UdVBr410r23ndeWtsNDwL8XhZhSXr+xhSWCM/e1W14UQqXQDmwforfFtt
gRHuug9roUohvHZwzQ9rQ7X+MURZWh5r4mMOcE7x8S6auseYVB+3JvKAKGk6JxZwIWb1g0S3D3kE
nIy7Dw4zhE6nnZEj1exoJ3/B3MjlLuzXr1zS3QM7cMU0Xg9JHd/YXBx2+lYBH3tc2ITqcfY6ykMa
nJzOX9Beykn1f+GoLO40/iYzBFkSnsGlii/fHTKqHd1lApkmo4R1sXnNklhNYwvcjxtmPUFVrS36
mFOiVPnVgkww6hyV+Wz8OIU+WrPACqZJvdcZs9oV7oapE6QOYXt62VNRYukAEr8BTk5mmNiNjwz+
p61o9gFjh8ZpdFyli8bGFRp7OdnoXDZyo68y317K1xGbyO5x6zyMxQKbg7eEzR1WQ/Rc9Ns1OUxk
FbSNYj/fM7/7ew5eb43jMk8Y16Jqv8YGbp26feVUX6ZFAbRmYuTNTKuGwhwN3bdhihqkprXnI/h6
pTZANunewc1CkdlSQQiVrE7C6zOOj4HbON7J3ukDiD2dbjm8zloUKCypvR7kRfrouQlDh88/gzec
W7BDOl8margLvTpxXrwkOP4YURDGYQTR6oQR+F9QBrxacGpbLUoLD+jS1y6rv2LlbD8Og8HdVuK7
BkxWZnIUCyZTfdAKfRyBbIydbaJP4UefCPspQRFNI7LUqxF8/npxdOL7/BXfLl1yIuv2EfUSeaeC
Apbr+FNf9U2hZjgmBor+uJoqJ1uD3QIfMw1nIkRcSFVblXHvQoA6kQisuCOdL6rvo72f2ma4xBw7
2LNCdYDXz7rS5+wiyfQIe91OpdcjnPVOwp3I9a05V/aUs+rMfXt3XJoHKkgEDh9wapcLZl9Fj1/l
cRzvk1JB2pzoibSraye6svtiOYlzzj3VBtYcCGT28hrh9L3jQ322MIXhOGAFv6tJWDUbVEpF5GAb
2oW9gRwoYsEFh2t3/phWF65KgyIsBn0dJ0MCskk1Y6a1u+pEGFJtXWbrGpHqqWugCKjjfVTLUNmZ
f1ve+3he0IshS2g7/829YzF1vbUfON+WWgaKUVP9//ED6443ff7U6hxwePZiW8MMf9rYZdQaGbj5
LYBG64LAFO+Z9TDA3YZQaETCyuf93lO+aFdcxRM1LjDfzmEBEWVjsjlI3m8SV3F/Qf5Or0RbPSRb
6DC3L6gq61CWYbZt3DOBUGZFLsTDzAwRcLxC5rC99QKxBxtTnfCwrd09slXYw4n0KzgOEqO5U8O7
IBA+3PIZaxUqZnE9aX2RkYyVGeOJANMRL3kVidcQeGDtTjxlT7qDEoCXSE6tLyTfC1Bo0uDTNRdA
aGrw/CdCKI8peHHqLvTaetAjPpzBlil5x1F4NzY7wJbUQOGgGlNxLi8bATNjrDUu2PUMxDZ/diR6
PwzGGnDns5SSXwOqdXBWCDkbEcXlrQ7yLAIny/jBZHCMGjOF2c+9jN0vnL7p83YMiAP7risYjQ4k
m53Tka45MmbPWEn0DAbtSHs3TQYV94knn1nS2S+F2dlAOb7JUrV3m/5SF1X1NEkYxmQ/3BmXuQlK
N/ZG+8eu2cRcfJZ5BG3K3lyNHBR4pjs/LfC/8NWPIlak/qBTn6/OQKknMIAfMJSi2ZuFPuSiDZHW
PNAuCmn5nU8B+Bysy6kD5W71dyElvzYKphTQ4z5G6hE1FapEigrMOW8wvP7M4qjsn2GjwcG+hkF9
Or0qCINwj5+g284jetORQ1bAEX+jAWii8AEmiBa6wObf89IlrXiXEOhycllRe6TYcDERP8MV2hLG
siEs4tF+Ly71nrUkV3glmTQe6ctlkBSU/ZrV3wf8vEtPVHWUP3j71IGvToQAu/dtshOAgdcpqBzn
0bsKfbBCIyLclVes5rmkL28rm15UHeZxgtE4iTfPCsIrmMiYbiz4/i8Tqm/BU1G9bwosykEH+WuV
US0YzD4JiHxeZ1tC9FGqNQf5JVvZ1bYhjNGstzN43Njw8gnPZwWKfdx1wp5EuOY39rRk8ycDRQrX
2c3z7nLSEzrtfNWA0hIUvG9wvumMgQspcmThboPRqpmNOddPb+qVn4CqLhRnC0Tb7SQmIh9ZWQXe
rUTGy4th5I/eAmhLEyzwzeHh03JAd+zFixqA1akSEqMTG3DtOIa+1xisKmdv46Q/4U+cQJgEbxRM
HmqjinXa+fHctfGPGa9P9D+LUs8ZmSoruAcbByP74fS1Yxwtl5dzkqN2TNs8jrIl12riaFTCqXw/
wM4Lo/6mPrDKucO+Sm9TFaVXDyLydIZJWVOYFlvHIK2m9RW/L1J10yDSDO3P2z5Wdrsm68lWCtoL
rDxPLNbGoc0ZFOAYnQ/ke/+jccOYNtd7uVNOgqJ0Jl2XnBcO99I0y2UGFhrNWfyASL+JAgTMG/q4
dzknGpPurX6gThwML0J4BZYpTsJ4izCWloSIaT7XuhLu88mIYDadz0NAhzf487WP7htAF213ofRL
62ZliP1dloh6F7Bg0xeImcEikY/YtMeiju00d0qCrs6jpEZQpvEtIGLK0EIfL8vlG3eEJefYiW3V
gxi/gfTDOaC/eDI3guF9NVt7OUNvJEoX0gHpQ6PmaOaz0bS7HHfy167TOtNez4jiPClnar4qHzzK
k6kq12ZOhoWYpBnneEadoYK7ULHxBi84UcYoukRfH3wFOElg8b4VaLEYhi8uJkXRZZ+BDjLjwP5e
bOVUWJE1wY5qM+JnZQxPQyZkuSGq8TPAq/+xzfN8Y2fc7H+Ki+rbK5wGSAib49W3zYJCpmd/AChQ
fzvYFwl9Sk5k4jrtaF1dRAzFKwKZEokYfhiOKPFjyKCROrPYf4oAaQPvILPlvV+zMKjPRAyAaLtE
POhmhL2XGEgA2vhLm4SyG6nSAv5h1F0I3myv6H9PnnZLt4QzdzORltioa4Aeds72w94nzoq1Heg9
p8+Proff2d38sTvQDNmVI1hoHS4kA0yV7Arp5L5VnH5gCEVExd0dvvKgbNi2zFz+l7Pyj2I7M0x7
WYuxF+yTJX5Ms3Mi8TVHCukAAXhTeGQ612WktXr51yUx7QlmE3/ZgK5W23NS10moiu7I9sbgaCHz
ze+6GYgn8mR4s/xvaDc1hHxu4ZwP5oiyf909Ef//XhLFZW42X6eT+jcvnMGZjq1SlA9bKL1amvcX
hDTvJSJqBYkrrdP8BO81Gu4F91xrt2o1HDG7GulM1ettEnyxgzH0gKK7UoEh8uQmbUCEuP9fQfaY
6Bo6cSC9m48pJoWPcJb6KcPjB/FXnLOzq1nmhaYvIb2n19nKSA4o3q71AgNfRF09/Oc/1L58bkXp
jNn2bGig8xo9RLinuw1/Q6rXkke9TXo+FBgoLqjX4wO+sDbV9Iok8CV4VhM1MPO4x5gPok7/Z0Mq
XXsp+JUA+pFvED0GcN/C7mL5WFkbSZIUY4yoGXBXhB9YxVgpsb5CO3wSP5fJ0MQ5JFnBPKxiAXRh
2RjzfbsPtEzxNIKBF/xlAiTZ1SDbf5WTzu0Ohn0hL5us621r6npoygjnZ+WSuTZ6BwW93JSE/5IL
r3x1Jxlio2dMnIdsbXgYLRJgS8lvXXzpWRZ+kcAWAXh3kvlQe7MC6gUZJoc4rDt37deBmdsBBOja
YUcKxEapKQqNh9lr8Ew5l6rcb1gQF/IYxTBcGzmkMMa3AaTvVM0bPl/zeDx9ErRSO6Y3oQKaKXBF
9JbdQ7M0BIuQk6d12eUTRN4T2LUepiym5R1mUn0DGX8SnviUggcwXu6GQRR9f0WQ7FzFu/gSUIyy
gh00uXQy96UJVjJiCbYJWwEBDsGkz8kWEeHzk6Xn5uqcd6IoNOUhQx7HWPhynMWwliev0o+mciqI
RYdDbTeKup/+6i/fmgueZ1BuXcJzmb9Lfe08XubkwzEUulrp+slcf77Pq5BvgtZJ6QlO47EQn6Rd
XCyioKc/BzysoXXwti2bFEZPqS5YHQfTeKt2BEBwAeznwZojm+8AqEga7bEYO1WOmzWMABvH2l/w
RWzfK9/NmXe8BKTvXjl3Dlgu8Fl8EDZRqNVQN8oR8t5OccFkSOKB2D5R4YTiiJA2NRojd+kEMZvl
yd26gwby/EUVFPo8iXLRTgDRzFA52x3DPsyfLpJbfeG2FydXB1gAVmelwxyXUdWjn9oARrv2xau1
rFzd+JnSHkr5GALz2abzvu6SydsavVBdisKmlSautD9D7Ku8A/vQ/wLPuF+2cor8SA2Nc3lrYMtj
jureZptZjdZHmqn3zUb4WNLpEUs09NvlgS/5nUwuFvT3glFryV0khQGu9U/cV14XS50rHI682kTg
gjZjx+m3iGvydij4AZ0zgXnY//rUYUNgh8fNRwynqcDhJTzDXeyd/w6XrKgLpGl57X4UYKgASKvZ
mN5mIN74cE61/7V9Jdnjx9GaPlisSDYgYZWhgJuXvGOZfr763O/S894Gb72IJI8sRjMCSoSO/dtB
gODEdTMPJgWUzmZKr/y/QQw68YlijLL+Zx2n4YZbYcfmSE7k/dcbQpHcZWxGV1aAy71SfZiGzxaN
YpE1bY0pYHpiWOortzKxMSy9+dzgBLgABYZ4Cndh1LtWmPmZYGUn90tcuyhMoF+LC75XuGlWiDg1
nIMrr5tNVk+r0vb3/sj1MMPANwAViYT+obA5NYVk0MDuMqlilqk7bjVzqMpYZ7iwBouqoNyws9qE
yidzBMd/vRw8Qt4+FekS/Vhd1idzAgcIUnaULrcF7U/Yzjj8FbbD6J1B6y6OlWCjFj2tMKILxNc3
50OFh8Vrio+MaUYiifQ49wYIv3gwENnhfIQYn6ksfOUXRndTKri6+hk8C12xVAOPN0cRWqIenaEX
mO/YQbnhMpjegswiDNckaiXJGUMkLqZ2o6ykt30xAYpuASEe3ZDTXTTZ5z+YTEnUkU+VByLli9SJ
W4k8cG8ZFW3rJVS6mwl9Qn/DwU38pgYjUNdtfOR5IRr6QXOLN1SeLC3HWmWMc2LfPY+mMWECh2k5
NWPBepirV4OS0QpgLCOWlwKpI1F61vuA6OE8dGGQnUakbx3WmDuhpbGbLfI97aJRxFjEkdjZEdhb
yWmbVhIgBDA1gNYnnqVZckie+3yQVYAuguSENCHG0xlVsSP/g5SRec9manhf1i6vheQJeLo8mFcB
8I9ync+XeEwluC2VOLhMw3i5lVy08tHjLL8ALHshtM8KJRZN9RwCdGqo95kvF6mZxvJKP1dRLKx1
K63iXzKqQpKwsZVVUO5Du6gtJ8OMdNe6BwOc0ZPK0N88BLlpS/2eVIlq7e4H9xSD7y3U88ScyAEq
7bIiqhVRpB4OLol0tbtO0Iu9Oc2n317qRQmm5K0kwwFHbh50vlDXp5TnbgQR6EMVQbG72Gl1OcBB
BQzUcmwXb2Tio/cNr9ReqCrwbPtVse9KxSYbm3FXTa7YogQuJ+2PsNwHvZmh95cgRYMiHosnwC3g
ZIpXfIDLwQ0A6rFdPt3wFaXhBNlji04uE821+3c6xeMdjoeEpk2ApSAhz8Aggd9xQifLij4XouvI
lKmLrPV37PQn4ZbkAaiFfKbUTjRbqHFNYfPMnL3oD06zJB/okZuwUO2JVA/ixqcEH1SAuQTxo928
JFVHsAbITN3xE7mA4/MGWUa7FL52wuwEo/vrGdIeq43rFkyj9vwYgjvHYAVpIV0dVvovXbegF2gm
3chgJ56wPgmDt/RPJT756UA83xnHj/GNWmm+FfEQEnlzLYK/c0NzaLuiacK3OqOCfHEaCjnQVWlW
jwH78HiEIc/c7Jz/vXFXrZF2/VL6EwRK0n9XTyS/tv6EXZ3/Z662dJ0H0DDwGq7EsIgu/M/1kMCB
qJMd5a1x+N2AKxHjLqlUXjFwT6IpPAIh10a7DXGIniM5B5SZJk3yoZAL2/PzINdtMHBl4zHbNV0I
cYAGapBgP3fFqLQbFWfvEZknv7C4YDr6aCknHbby+YgToggmpVJ72bTqHxfGvsMnCljUD+rUb4Lp
oCIUPwxXe1qXNLHMs/Am6w9x9iQlQKysW7uGmBazPnc4z4YGkoJfYaVBVnhA/2L9TMMvFVaMW+8y
2sE0BN0oBIg84ek79+kgW9GsVsYZHey4KzwCcPciRirF0nYx7Y4wQFxImxl9O4iF+TmBh9socCsN
icbyAim1b+LhpF6YY78u+QFpQnauCz9gdo4OCgQrjgbEy7ryEiBzgl605J/63F3YICnqvEZOafgZ
MKEGvEAeHAhDuucngiXFImLeR5ucG1IP/xfNGvTmzPc+jOI/3141PY5LBj05veehZyfBrTxr1DxZ
pPLUtEmuqGlRLGyosfgKkWHM8EocDwquXHpebYUsu/MnvY+itPcZws75CWBqo5zmNV7jjVGukJ6h
TG1TCkYdrFYxe7onbYO5eIokCK7kyHSAATT1mGAnyxyeo4OqYq9LMjxuHHaZ42MZ2q0Z/bgBMSZh
mKyAJpPpBnxSBESpgYxSoF1eL7wXSh9+l3lxAbFNiQgdkR+WMwh4eSIqb1Eo7yFC/xETDm7aAYsH
79mZWGuNy8kSyhgR5aQBStFWXi0xTFpR5Es3CjQMdTkISFPPx/uJp8JZH2Y1nsn93OU26WlVBk4V
mlnQlSQwUv6md0dRDvW8Jw8/rnhzrHyXk9r4gBBobYr/hG68cRzjGJVyrC5LQKKsjlTWNsS+aJcV
qOe+ANcVQIPbME8CGYbGF/jpR7rWQkgWxjZgCTLtb1cKv14G4bGIqlHVYazmYuPyVwxhr0hrkprM
4e7ZnK1dSdkl+7Emay+cVQeDXhDYhUBnFyfPajDnG1OslGLeYp4D+ZSGhteujBm6UmBWuwErYxe6
D4fSxm4Jidex3bdJV8qojL+u67tZ6JW/fYfpH9r+AAFGPVuRiTJg+I9KGJm/wEUsXdtgT2j6+yen
GeU+s0fzuJi3x6qpFmuZMUUvfqwxT7qZqDhCsVSpvWAoKFGJFIsQzLgquU+pXval6RSh0DGQeu6k
OGULURPz+yvuVTH5ZPsmEC+CULqpKy+JMMohaXkuz4TeRVkiizhTwmhWB7KNnpSPtuOB5i/EDgiz
IKrWEYbOraIglv7ei/ZH3kiM8gOLSb64SwhR7ytAZm1919fOVSMnrkjSG71MXp1appZO3fS2cCo0
Gg/xHvnczbW19RU/ZLYb15H0Aw7Oo+7Z4yT5dJev2OCmbcwMbgyLDKjp5WAsYpHlVOlmQvThfoS/
FyBLRKyU07GLKyQbFhw2h0CRRwNUqPMFdlLhCdk8zR6nQy8cEKjCGS2CcOlLYL3nnC1OdlUTCdm9
XxhPl1pE1CR/Saj53XehXggU3rV5549kSE3I6BmqQlmU13WMaQv0GeReEnax7Rj3fRrPMjm+e/jy
aAOXPyyS0RK+1ttvw/yy63RYAwprF2yFt9gsqBdCNAVBEBZCKwNI7gKdwzz7Kw1/7Yd7grbmSqiO
SdT+3h1inkRtM3AdOHGPpoXYEYZISoBCXGe5P8YTvMhVbA+H07gtFNKaptAKWhHeuoYqaB7Myz7R
pzQ8DrWmgyGLCXjmR4Tn5p1iUrxno00nBQcE7r3ApUTN3o66dNXZEzuGV0ompk0Tn2tjRQJOX3cX
z1B3kPOkACcFDBRN3MKHiW11fXBCpM85OoDOivfKykyT2Drnn95hp4ppmDhpnGCiMUIRaLPe4vEo
PFBJTBYxC06sA2SfYqX3GtTIs8GJ0qe+xh/dhgWaY1Zzl2SvHYEkneREcKmuMwJljXbQT7HfQphP
kRKSZimaKkf6PQdHXOuw7CzP6t1zedrZlshcCyPXqsuALCDSknl8/Xpu22OG+etTa6uWQZNSJY1O
7lTS6cL416TWGlPgi2CIyvsa3Hnp4DQVXfYRd033IoSrICdj95t6elbwD0QOe8l+jvW261cDgoY9
acH0OP4yNgCWsh+9JEdMVQhP7/AgZgj79QW41f8sPOb8sicfOgwjt4Zh7c6sDqvPfnR5ddWoA/kt
JfmhI/ezvFMfd3RbRliW1dyM00pinZV4ZwhARdHUy+cVzZVmZJBTIq9exrcnYA/TxuzJIZqfZUyr
1uXy1twu8N3jKefWuhqNdGEM1g2MvoIbRR5ybNnPE7eQqdkLwvze22RJdONqp8oxXgTG9pDaDEIP
VKUvtBkixA8JG6klMRcjvbJShVPV83JwLvPhBnSLHLh/M0ERPdvKy6c7LgOcaQdzQl4FrQ76oKIU
li49ADrEhKzXHcUdy5bVhMoR70knoZBXKGaHN3UnFC0GUd1yoL2sGf+Hnd3FcDleZBQwDffhvskN
BA0J89UEIF26e8nb/dXuJYIeqJXz9DdXbqmiOTOsMxC2b+tcohkvGqvO2D8z7ghVbnlAOfm93d86
BUhjsMjiGZ94p96ZYEtBSYLd0E5gvhm2ViIUYejYwnROtryUOfEiN3kjhp0MMNG+PqDfl1n4T/+D
Rbk5HKXcgBe9WsI9Zctc/jphX3HDKqiuNWqHNMzFF+9hwmXeCMz4aFYW5dPcK5MRypT1R9fCIAso
63TD1VQDds881xK8m8M/5kDigwY1wvb0t/IT5uvb1CqLaIDzwVu94dJOOPPg/XQGuUpIeTe5OSqn
M9ncmJqy16xxH8fdlFCHZuyZt0bSK0VHMsERcVKk9JeB+1abqx0KWwizayhVsxOb6lVZ7jKFpkIe
kcrkQCUl9mcU20ZaU+LznY56RqfScwmLD9+iP8t1G3KpuDlrST8K6TU6nfee0/aaN2mpwuMVqps+
5kF5n5MWOK6r5dE1eUIT3u2y525eEkp4PylsmJIr5vrZfGtccOc1DcU69UyjkomeH5NNGsf9aXLM
v3UFOIMOEWxXTvvSWa3bwtTjzySEuU/Yq99DK3ZYzejDqpVztz+g6RQARcVqUGg7o1gnjUIDW3Yx
vDzzsGjvjfzoKIcXw0fQofwfyEY8GHWyZV6+CNv4hDCeBy5FgoYn7wzN1xCwiKaEv8ufgxTocOMA
WXsCCmTU+qqL/KDmIiPMVxT5y+EyodLqlwiSRmW0qSpn8KOGcHvQJwTJyLwd7Q8ivD6nom+IbNp6
bMoWTRAh1FRC0+7xkAhM3++oJg7a4JOfNe+YUgvP/QOZhqrTz7ogy0idicUdwHNQMi0l5ROOrl73
DS3JMynL3Ht7H+YC9sBrfxKWUyBnjW+zsziNRGD3KvLAdk9MtlgxEoWSlssN9Z7CGxg5QO1LeOVy
67LwlrbGf1pzk14vXJgbBLpsVbkN2daCoctUS2FpBuq11e9d6g/ktXu8QbZzVte+zWZPAY/wQQ4t
2zXzSQiziohz2ioLqt+PeKKTDmVnPLxuwbVjdx5U8G4tswDBfb8yehQnLKsJzOwogzFfCC33Vx30
70dC1QeKmUJ2/8rKzlaOgr6iHJEV6gvG8lgdRWJh3Qg37xxydR2VfF2KxyuN3oLli77JkTe5PcXr
HwF7z3twAWlPo6S3kD+++l8UZS6Bdxdjam5aUobGrMnPzbpOJJMoTIEKJF+rL+C3Jl0Nw+q+CJqE
gP8k8T25ruLFAHlBN86x0ZtjpAfSVEhxkisVsk4f643YCUTueY5bvKyLraMH8RJr9l/aX5t5nWQ0
S1rkqcT0iBYY6i3p9py89LK14ltb7gqDaATIJQZM7/6opnEiS2L0xZu8cS4Dk5ntjh/UdBYjOemf
mH1CRd2IGXSy5hPJw/uZPPVtqnsxoIYr6exCE4h6dNN0f6vwpmzs/csxmNEPulCGaieF990FnDPB
l5FSS/nLsKzt3Fla5UPbAw7A11XXqDNBoiynHIJZP1P0W1/+Sw2he50WfMsZrMOI0rgiVgtcKBfz
kziIlodmfd9nVoimIsfvvi00fHYafpd+jvyimyjGqYmNeMbEpA/qLtYHB25KShzYRbaKjpx4mRoJ
4HJzKwzHy46kXc1wHpqECvOdHSzH7SVlcDxo/zmvkjKAsxPZqKb3LVid4ZA09NT0FG12BL4GPV+h
AxzfW2mcZpdldovucMPW3Ji8XrAReWNMnjrsrQ8uX5LnR/I6Xvl9eRs/mQOwWUnMipeIuBw5mTKG
OT3oDrAyh/6yJQKmwq4/T4P1IMjjMLzH0mp/At7FBT7h5+FtgVFPr9f2cPjEH/Z73t/uDDa1FHTC
o2ikbg3ElGaw9sMwA6dJw7QuG70i7U900fGfYD+A8QzLtKt4GCteYna6GrvWaAMLrMrTVDuCTQvX
1SZkDQGBro2Y62LetVZE6SNV/K5kHCZGTLVwOOuDAptAOgs9AzIhCA6hW0cq4ObXwNnJNGuU5J90
rdoZdjrpgVkH29zkPZhvH9uuryA/s17nRQun7gpqGPzp7+WNQBmTyOECzGok2JGCSoS70qFmVEhO
k9n5Ct1HPQgTwZYnjZgIikiRehegvo1NzW6ijLlG5V42yv6zRxS/WK5hOXfEeAmECmAH8BaqIFOk
C5tB+z95gGG0TOjKD2r9gHoMwYGnAhRmSERGtOz6FN4tcQlPCZCe2sfTXNa+4vTq2LBtSwlTOrUx
vyYpniYv/v/0H1IJOEpBoXbAia2oivEzjx1lEpup82iJsIoBldcK24MsGrLGx+aiCrgRSvfom9bj
GKY/EvzlaAxdMhbW2us1/OFqXz8vwau54gdjvDlW4hFWzd1zmClZ1jlEOiakzF0q9wnNApFsK2Qd
FWxYfI0lXJ60dhJULNdLV6W2Y0mcCi7ZlXwMEkhcs6qKJwdcqFtSPYteQFp6DPQpLi1rCsWKau1y
cl8O3ijeeY+n6uIVrcQFCeOLBD8UCRrPtvRcMhskiGM6yskPzG6c0hixBmJFd7NKXdrP7UlSjzPV
DC1AefXYKAZqaV5TgupCUlE+kDu8ExJv7W5QWUkQWMnOd6oBy6Qa5uZzl1kUpFxw31WH522hJDDd
yBK26gIp0V0q22RGTeo1FH08YPicTRRp+VCw/thHxzYsQ1J0KmKfOzb02TvgWk2u961gju7Snlbn
mLrFamztE5p8zPmWts7ujSljT8h73PfolI5Gyb1Sh6HRJ1pxFejhquaf2sZY1Fd7JxlRBzhxgZ9f
PdZ6ZvoSK/m2WWZCWCl93SdBjVEgzfrhoVxU5Ue6fY7Ld1V0j3YROJEuDQG3Dkmrcq6F+N/uZDfL
Yh364xryI8GPFV6NRWixOACbKEWpeiz5DMMkjH7pk8lqtknu3JJ72hewgQMsMDe+Y//foeka5qnf
fmpr3k3bAJBdciT5MK2Nye9IeHne/gy7Ch0v3u2qt5KIo+09mgyYz9jaPZOZNHM05pfGhDS2jxRc
NH32ii27L/jF+fH5Ca6b7kDdtsYb8myG6+KeJM+RMZ/76kLG7662XKbnmV0oCn46LSFoTJ4eu8uo
bbql6ERHkz+9NWPq5Xw7zGS20fK7X5wfKaGpvdzgladQNZumKB98rhWcPMNr3fZQAa6iWq634gM/
9lTHDf4rCyIhHBlwQEACve+1z9XR6lx1FwDt3SYhQOkNBiIsi4SvENyhtchzw1XsfNEWujsJX3hW
d/BttOUij0nbjllV48Fwx+qgeIopdb0ox4odtP5OC+ot9MCQ3QJeCf4XvqR+NHgKfbx3ht91NUxE
vG0prmAewlwqvwtFtSqQi1TLPcWZHFdQ2j5t+Vyb+3zgD9Lyj7spmCDhoQLGXc/RxnKfUjwUU/bv
zfRCzwHy8KfWrxR0rwgYN5+1GDwiJJsqZp99yz0/Tt0NHebGWkZLXqjXKChjbvDdOp+YlJW98bc9
QG7d//hM1LQDzyJ2imK1UPWlaDcIrdj6JvIoSI+zlrL69YlyXyQmd83ZKQzkYSRN9OGbijhZheZW
qmN59VgGgK/XR2gsN4uZDBn7VM8O7ftztmc2dvGy5T4lXbnh2qGEzallw8me612c9FmmeHjP7/g9
+c+cTutr0yGSHA3lOVLFulKkpu+zI3Di/XLHU0vJElhWD5ilIeVO35msUJOppPtruBi/7c27Hc2P
DV6NAYhIimv6kTM5pifbc2oER8RH0AmStYB9SLHsyHsSD2V6g8RWP6BD0g6ElMjb/1ShFcmJ0LgW
gptWMU6TwJlURLWsO+PVVMZfdoDZvkBc6KGUh2mtB4zRI9P53gXfn1A3jvCDlOnHZTrHsnE2fzxF
GOeR16KjHLYb+WaTfVU3ky+HP7GzcZYfKPxpboQkJbVgUZv8HNI6Ph7EdlIDx4qYCAJH+ot7d6Go
yB/hZLnF6UiPWSBv6jrID2vPThHwBQkRzSNUz1GcgiHkW/dqYUhmSLv2ghOQf4NRB9Olj4qE75ow
lxfiTFs8H49uOBVNps4b7TLqcxFZeKKAhcJkc2dXAdlLfGw6pv80Pw9fWEUvGtpN9wMzQL9mzYg5
HnQf5AN0jMw8iK43IXilF/BaZLLHnpriVH9htfyoqjIPrSYz+IxDvfdn5aemL/1yk6xJw89QA6Fl
vktJdq66bCiwJEgo17ueuEl8vD1gewkf7hgxFM66TN4OMqoP6jXR1k8yHbfA5zF7T008+WphTn4C
w2Ho8h0H/c0ALF5kXzoV7NQK4PZS/W6idTyFKBWRB2AomII9DqxQXSwzQ0VOn3FcVFRlZ7tuX7b/
8TyV+XVT1LLMqzZSPOssuwt0deTc8G7KmZN37JtXd5FoRoI7+hC6IJHOtnsQbVJynXxsorewTSZ+
TWjCVyDMm2sGxesTXHqA7W74eI6yuPQcC95vF6zEAu8wIcmqRaPw4DlownLgcfJwaiPyuOd5g2PO
PgO3KVHzdkGLSlnjvSl/+JDtTGXw/xpTDy2b8sJlqWUXAkRUi+AnaGAaSHF5nTBejChTWybmI6UH
bJwzeSVj4FNOWlaqlZysIYugfEOMNdTqd32uSRCHiPh8aUQYZbtKiZMtTT0d2IWdTA21qwhxQpBy
g0Fu4okrzb45fBbwyi+hoDltVfrAOxorXeZ151X98FYyUIWhuhYDEo2ciXbGUK1SAEM0sGoEukal
sZgIniyE3X4cmdi/sk1iuTqj53CaRmDYD+CJjwUiT1O7Tgigz+63hS/kiHMMk/hgVSdOaK9dbK2b
KtIbHsc0s7OLlq17L5ckjQnlTSh8yF8SgYBHKPSUfkwjZY8Bgo+DnadAKxvRkx0NbI7DUAU7peoq
VFBuel6sPFgz8AEpdKmnMj4g4vMUrmJKHYB3/IdXE/9dtoZsMjn8aXDeU4CLxNniG9qkKU8zPZD3
tMtgr1o03E5rCG/Gz/xj80jHcOmX6xf2NLE8lsmg0qpVu4cmfIpgZnIMYiKrP2ggFXSYeTTsgB//
2w4Da3pB8H4Lgat5WXhphsDHnwvr9eKkl8vzENfl+PuQ2nsns5WbMce4G6x10524r6ZpENIjea/p
4Y5b4fsalyRFHkQyBbu6BYKukhW2Fcu+umroRUoHZHbKimvgAqdqMPnSEV7ibIr168kU7gwz7WPE
QivQAoSpG+WC3JKUCRq5i4TDJD443leA3aGlRC/XUt09sSLUcE6wDdAqHZoLbhaQliJoESx+O7gY
CpxzMsozMZC7LZFpXqejjsxjyi9WW9WpPekCd8Q8Vc67dA5HAJkqsh9kOfMJAuzSXjNGVXSX1yVg
m2m2s+Z2ArqVj3SYvqxvpv9aIuiOBoRsi6S8TqDiRh+JIuCSPMVOKjjnPVn/xE+O+y/VrCpu09nt
gPN+H+kuxPJjA+t4HhuwFBbK8npVkOxE9HBA0kv7vyAHI2eTyoUXJe3U/BEorpLTiY/QVhbt0Om/
LNx7ReugU+c0guy4z15eghOqBmyAs2XEcEG9W+PyrsWMGibilgLS8I+5iDkacIZ5So734Cz6FpPJ
VKqEZ1wWNWmY7t+r/Sfb5uqfL8Q2v7VWrw5lSWx9VtYDX86x+r+FoK+5FprZ0zRZC3PkJSZtep1p
TjQkjzd7rrbxSSNaqcVBsJS9jo31aw+wz7QZVACwgGEf+Ijukb3U/nquRxEL8GUnUa7qV6XfJ59U
N93NGld9OdGEy7tjSLIvuS0ujfWYq40SkH5j4cLpaJOKJGiZr0hNnkY8dLr7YYfxMeMwvj7SbIZJ
J6/rffkN1qosOMiaH0JrGrOWYfAcu+eG+QclaVitGIrmIxYlj5The8v0Wo39WIcuXgZl4pRhhUta
zWUIYN9VQ7dJ8otX74DzzPKyqONu0TB6xaHvVYxSzQO4wJwiJvFp0wtl9NxMFFV7Ov76WIXVOJRA
VKTmXlTxGvDjI5wPy98Kw+7s8kf9QzKcVlusKwjIulwMUtjm4zVrtqNQKjoUKviDfsFdzPK81b+8
uQ8czlEfpC6AkccZQFF9jTzDx4SuNGfRElrkgdHXrEvpDeCJZi+eUst6SZYwfr2MXwIPlrkocSSX
B16BqDZO5OCnF3ND5Q08hdOCa8dOnrNqeLY59wCmL3lyXZaHrMnw32OSt0GZXCu6keFe1zAzxtt6
tVJptnOkEFMU6M+aAJDExdu+sddt2aeZ13P52Hefu1DvqQGXBsnaSN8FztMXOXf57qg1KW3wQNZw
Nt+GUnEz92fL+4lXkW6tqs1Fm6lql+U93ckPWoZmXu9XZHmlPol2bl30uEmXofaG1Fa0bJne/DYd
FzV/RmCGXDVj1rIlIoDlFxFDDzjQTgUyljAKP7lHPuWfDC01a+cQ6Dv6k+dbV3mwhQf9xoFdhyhI
6+u+813BmDClm10SJGgkdfT97xbasffD9cyXHfN7vSIDE7avBp+Dit7+lZh8fxRdpiZ9WVoNYZBn
fpfmp+nv1EGZ5E7WUfiQp++85IBOkEB4wKq6rn8cEJa4hm9tk8tgQDJ2/oukYPtNFr16CiXwuNaj
BYc72GKY262/1JP64sxdQQ5GnC8+9Cz5OLuLHBnEUtdqKBlOSBUeZBHSTN4QDyfeYIC2/7XvxamF
HvZIQVo/xr9cwcOQXTR4Q36b7a39F1Q/HF1eFDwZha243AqwxmX7VIvwkR4zbyAtY3VoPoJs4N+D
OG+ymi/fUxTUcXDVteE/fSBREQeUuReelqVXkiNOg80SgH98BGTVg0ipiZi7eFwivhpqk5mh6sWR
WltT7IV6GK3s6QKrAZc+S7/H6gDa0kVVhZfKFlVbnIil5TbbMxwcgTCYue/Z67rxJo443Hl7JyZd
T8DpWXZFsv0V8wyIZeuMCm25Gz2VHtFyMen/hDca1Mvrw5NfldWrxk2TQiwNDN0hNpWm2TfK0pqP
h4NNDMazkcnkmaU+4mnqyQBBG7ucB3atm58mhEjATYOphx/aEJswL6G3sGAFJgifNCDcIGEQ5vee
Ikil1++r8Jjm4v1y+GH+Lgd6HlwTcsivGYnBgyp07+REU5DEY20yqu2wkxuQsmaQa0JSvKu/PCL2
WYH3CrMbglzIIgutQGD11EgQwut2Jtz4HHpEWVTENene7ghC0AkKnPlRjAaUjjqHCaISXFB4dKDF
TWRgn66I6b0XZvzt6NZ3QtreF+BZl4pNMZ1mEokFuLa3frtnEa7khus17Wx6tf3kRbZmuargN9qA
XOEPhXAoNPl1wW8k7+b3E/S7wsQyYeV/mSzZFzX02u6Ml8Vd3CQZ32MoD5LVWqlj07HLH1iGceN+
H3A9bEleeUpOvFyVmk6ZfbPjrtQ2CKpoZIyGTdMFN+eNtqrioj0nppdz7FgbDG42/uV5J8697af/
ZzCnlJYMaTYfQM9r/RSQ5b82MDsZIzC206Exlg8lzvdj4bavL9CQDJCwHWff3mzw4gHwZdVy+/fw
Rih4cELg1LlSOy8Ni6rzei1ecp6dh5cBAL609D1Zmy9e1Ys1shEgPSqWrPJZcLKqO45VGwNvoh0h
dS+XyDp1bw3K1fDWN4V6W6/FxqBOKhLVV4Wk6493gXLLxW4F1fN6PFVsRcepYygWcwVaokz02abr
gZbnjIiyYxPh4Tw7x5wLSdc+gG0DGvXwFxM6tRCSnZ1Mb/GrqlcqTiux7Ltt9P1hpdd6zW7A2BFo
9V6lUNPhscRJPg3yAUvKZ0ukpe3ORakz2EgcMM/8a7ytWjT3HigNBwMIXwEdeD3brpNsECMgw2nb
ZFZ3wCoozMnyEHJgCAz8SuU5a2T8PhfJezLQ5Tohm7Dsv3oxLzXgrRAyiymJMJJH6cYoM9+QTUIl
cHTv47DbUcwXEpqdRV2VwVnNrNiS4NtSmXwlxRWV97vgn7gWqYd2eRoVsRC1Kofw9AFmgSX7XzD5
fjUyUou+3kEa+p6Ycqwr9XCfTbTvy76HYdQI8Ht9XYko89QFZLzhFZc0fWkwmbwp7lGUKQBGbzka
ASl4dEdkf4XMUJynGRer6q6mfcdcTqF9GCPwCwSXFEM/csbQmwsES4uqxcd600u5mI9GMaBFoBSw
aLGUzm2ayfyc7rp7nB652uYPPKRwKJfQdMh9g3aG+MGBGebnerguWATlCNq8ApVH87AFKJtEa2+V
FIibCBn5EvaW25nChtSz3qnmHNxiBLNDIFVkvrJg34jc0PYT5OY+U4SAIwzYMu3XQtWc74E+cdN9
YthW7Js6xvZl2bqoGJasmOx4/nm7iz8JusqCNFz1ZGsqTvUwfYKFdW16hLH3dCFY6gGZAed5bHU8
BF+IbsYz/x6Dxu8x2PiRFHwXsOvxcqy2RWxG7qck9/X7DuRt4/26yzKoMjWKmQXGJyZbS/iBVtWH
6m2xOHAedfsr5ac3wZ0ZjFdVvqvys3Yq7aOio8Cul6i4hsIx6QFr7P9SI5uDc0mDtxjw9NSvW4BU
ByHIOmUmbOm/W2WTEqplEVHihuaBOYNacYJPOvD558itijrBKwf6R4EItr273rQi2rPzk3a0waIS
j5EKtUuU1TkLvEwzStI6+GiG5cDTnPpccxVdnp6iorgBVJHPrMaD21TdBICtXoYiLDYv4vicWz/h
szX1BFSNygz3+9gzKB5Ej1ckgLoqB99//Xcl5fJkNV2DWYJWZZioR9svvDkdOsmJGPD4xDMLCy82
a92jynuO24w1TjS2fndAfHz8PQ0GyX6ZSgjIFM/wLUKoRXkwFOv3Eeh6VS401vEDjehkq3a4JwnG
Ry6ynf0x/9mJNfXbWPIrAaJtjWhmVEWCVBdtCSavdPhyqf+2rPNHw3aJf+nRodKKVKWbcXH6QIb0
eMhz9V5is9GluDdZS7g2fV3EkZMPu3jSMnbW9LnzE7V2NTXx8xwBTwi0EmwVwlkgqXiHPkIpoXQ1
X3EWbO4JVbASOUyFqWBkmCPau1mPXIMx2ryK+IQWI+DbHjm5Sb6DjXn/LyZi6byTFiq2W4RcHzAg
HaGRqIMfke5J6a3fwe5E9T1sjpK3GAsQzOLQhi4X3jMZuzm8zgXAe1BVQVM9KxfxAiWCyA+DiqWy
50lJthVvBrb9oanB5nQmiV6IC/cRlveXktdXs38v5s+MQn27VCfBVStD2oHXttxpY7Vkj/KCgelU
LjkstHhkZAd05ncvUyHeM/aWn0X5P6EZBDC9T/Z8v6gillfWTc1Bmf3QoySW7uzWF14IompuxOOb
80vHzmhJmZ8NYS+Bovhfz3HrogP7h0B7RVhKgopROCX6hgD+/P3AvqOqNtuDcsoAbq/zKC2RtyTp
eZpkULIgJQk2aFYbo5P14GFUQpbe1xi1dj6hy45GPjmo+mehN+CsAtZ8v6CqNP4l4gBk5Q2m9uwD
GoC04WMnO8BWpM8Ko+CrpvqAfyzS1LNuwBobZsR5NTYS+0R83FL5tMGNVCbqTx6TESvp63X1UkLT
uM0CL7hU7eCOQjFvyerdGpODobQMVeMK4wRM56i3oWbwd2rF2sCSpygsXe7NYe/nL52WiHuYQnlf
kyNT5i3mSjFcAlW42Cmmyj9PpvEkxwwkzgoZ12fyxKd8fS+KHSeuklxfxmLIQjbzbwNCf/7RIKW7
v/53Aq0DX96TDw3Hb/yjiFpzDHxcpxQMKBJ3h1Uhl6/em5i6v6ptybAJWL57jx90zaEREBCSWb4e
n8CNoZcKA7pt31o7UZ9Kw2mT2iLiyXWnv5LHEnigJaGGj3I0yGiNs3xPv7xi4EJ6hVDWA+fQC/l3
8EjOFqvVStps65FeuvuChcY3H7pJKDv9C7uLS0yZnieeOuhRY0f+Genf+PvyFicWAwcU3dlEEJDY
RnivKW74MUfk7/gdYQWrtQburEnBnrPhZdviy6IIKAWGdeqnwPKv6MvJl44623/8C1PIcWH0b40e
HK8STmPqioJfCyrynnUjQ87k7uTJyfw74B06kVYVlGGFFRWqzhTEus76gA97oEbScydrmB9AXFc3
M9CR66vmS5gJ2S6N1D63OFZnBklJV4T3dXASdn2tZIAUsNlHGc7PW/sWwJTynOXGOtUiG1yhuoGZ
3rf7Wp4gQm4PSjv9YzpUvLf6eMe98pBZUH1YXwgYgHJZTnUJPhnscN93fHK+P3gC0/U2ZyApORKA
SIe9+B+/QSt3Yjf4IsDPv5i8Ge/4914axfYuaQ77taPBiLAbYoRfRnRVHnaHwGN+cH50WwdQJfx3
D6J3jefK9cpM9XVg0CbGvc3hsYE9BDR9EP51m80Tv/QmAsv7SyWLid3W1FQLw1J8rw40uYRbzCNu
/dX81ilcbBAnj3XkTGqrHayMkYf7U3mbpuMA95JW3V3qKkHKFfyK1KmqA2wwM5iBxGVSMbI0T73f
1vlG1EyyGKULcRIOmXbW+ugSlggbDdrkv2Mtg5kG0RjNimFLAiivq19CSuT6nM/HwgtzZj/9qYj/
NZt8WuH9r1qq5kkDQ5k6Sh1CMH2ULZJeli85JO2GWSFTltPoNboUChBj0/HmuQ+uFWjFreLPNnhr
mghR2hdbnwGLvBq+Q7HvxXmKwWJCeZm5pGJdLxxCY2Al5rE6AUOB26rp3nwLn2M1ukBfOEoIkkKY
n2jU9Jb6QdwxoKdZT6Q6YAylJ6TtRSV2jNeMLmTVtcmJA/mbz85KhKH0ZNN7jfJ0hgJNSJ3PHr7X
Rs2Fqj5I3gnf6dlYRqCTzOoIamiyF94CwTQvLGll3Cs0bOLN7mmDt7gScNIV6azAN0/xt88nSW+t
kUbnbDUKfk3xeFMZV1cpJ/Ec97z8WEMQ4LAr7g6Mw/syokv7ByaerDai0xDHku+1gWzYwfpmDceM
y70kJ5fES6CWReyR0dlaWEiiiZSULMT67bckyl6fNCRZ2MwPtPaOe25aX3imOuEBBLRWWdLMzaLp
WX/OVPqUp69PaTyN+C8Q8iQvMdHht7bWvMbB9vq+9icINcuV+EYt6VKS0KEf/py7FnkdT+zcHDpn
dPlslzK96bT7fyECF4cV4AJ0+rvOC72M4+9CTyQ/Z6Zl5uA9DX601UXjb3KaBT2oagzq6g5vKKfb
FdrjBEvTPumw8HRbib838wcJ+QTSC3pVVRhusCTGXJOlOj11lS9bSTVjC/xL2HleSrudJwfG4k/B
qd1Y1UPlMqOwlrFIGWBh88/q3+2fDc/KYEeUuX3BWBtJhOQxy4bHPofG0ahLR6hhT5Gk4yjWCcAS
uU0VgUWHqdTieI1YULpEuaJteSrSIf/HCX/0X5kFrZttw8efc2wJ7S3LwJkvHeHLn3S7HxjhIRxc
gy/OZyOgVlQX8O85kJunR1Xq9Vfvvb7eIoDyI8Z1MUgHOkYEStzLWAQJGpWgz22ZG1QsBwSMQPD8
R+gpvv+VJkZYMmiWs5K/qbXn2ge+Da+GvMPgHgs1Gr3/d4zJzdDcq7dnW4+mUmTADpjO5X1EHwKl
2PEzCP99UQPPSRIl8uqVy3aHAFi+dY16LG7Q6P0cxyXi3JrKemWIo/8nzD5GZwNG1kSnVgCTFOe6
YMEXkmVs2HgcAJqfrp8BKqUoWzhbesC3Q2HDTdYpS06hf7WOzuNnrwx66tEKgQ+wuOyEH+KWE6Di
P+B6c+kO3y+JXIFlLBEPAyMjo/k0+qMua6TpHpBIq/umMM2MFLh21+6gkSw5uycYd4zAlDFGoXpj
6fWaXKGQDZPU9FzbvlbWuicyvcXH+inwhha1F1PkksXEJGuE0/yoczHAxEIeBup/gRJsw36r8DOx
mO1h+y9Zq9DpyjFSPfC+YZNI/bwnws3sKwlkGZqOZEWEUXG1q/yt3vvjPocPSym+Y9bm9LlZyAQm
UPyQMODBWK/F/Hk9nWmu+Jcyy8vEG0TyMrsJyFgjEcmKk/Bw3BWwcvDcPvMtiC5M9YAockz4G4kY
n0yST/a5YntCvSP88OmnEovcPmxyguxsOwVMaKQjraeK3daDIgOjoeZ9WIHE0gm+1IxeQRc0N8NY
sSf0DsS+Z+BmfQl5sH4uiScHYKlKtp0iE6d4tVw31nBvQBXPPKa6R9LmzT/Ge3utx1uN4cMmogeB
wHjRWeGFregTktyvzXdsq89XVSRTKWfRozXVg6eb5Xq43BxGdJ/pdJ6eeq0eLi7jYvtgDBnhyEk/
p7mUbgHBgcviQQqv7ULKbuAm60/Dq6Njgr77Ss5KjeHAQbnbpaHrSmAhR4pPeh89rG9tnvbviBcv
IKOOEEENqT0DpK6W7sqx6/6U3FgorNtWkGRnt4C3VxID/3QcgvLbPVF4GlCSclssq1vDg1pGYJHL
k7zKCWZXJDxbFT90rHQhT6tnEYSWae+GZzRbUsnm4DSN2RmylaAuoMockaUvbTk0PTKuwpjcx/jo
FiHRK9MMw2U0wSZuehS7aONMMp12l3MoC4rnhfy5FipL1mc1qo9SWXAXnVkgThi3NGQIRe2UIK2L
BMsEZkPB5QTNNPHr3IlgNblVg+8cIQbGBfb/8qn3wNSE8wmhW+d0KIQsEttRptIAT9+NAnLM6yW1
A5b4PRWV3uEseC88xeZPCm2RYXYJL4jalGPdTPxEXaK8hFi+VoSD0QEGcLF6b/Yq6iTofWtR0oiV
3f2voC0/amPkC/JeXcIkDOupsJOUFkJZ0Mm0u6pWgClwYoseQA/CjfpsxDmnYwsERt1yiB8MwNnW
nEid8DDfXZ1Z/DKNIDyI2a2I/y5vE7hlTQnnRtG6NgLJeyb1Jqnuj8vsY+fvbQvk5YmHrvyptCO3
5AfNrviiB0/00R52FAIGxNzRBIlz5FTHoERNV6kcMR5j5Dfrg3IICIiMS+T8BsqvUBtoMhAi9a3d
5IrudpCNaG8dEDY+l05h4fu0mFC4raVSyAg7uQneIjnSY6gkfBHG6PvOwiO6Y4aZndu+s0jUsqhz
OgIp6D/r4rqERb73H/GUwM7YdMRz0jc9na0l/BY8jHYQnpLwyaQOVHpIQ2kfc5TnsuSHR1KYjsUP
MyTof8hckYc+N3CUs4EH7fLiKYzCUTXpGdVVKwOr5eOkj1ZskMUXX0mX3GSYhr78LSnBItX3JDSv
jY3/cyPJAE1Qgq0frsZ0b3askJMDnhkgt1r69ZREECxbl+CTgx0ajXT5+TGrGLEb1HBEuD7f81dq
kf+g+BL/f71WPnqQHHI9s58yW5EXvz/WcO8VnPjLcNJyZKPoL3Lb0sdRS/RVFB2kVhQcWi6lzrgD
PWo3MceE+0lXn5NRHXSCvpZoa4NyI1bRqMxSonUgxFnp6ZRKZq9X8SMUEjV2cH2Rhq0Og6HCcbjS
g/FcCiuj/KXI0VusAG4nkdrjYWKOcGzuBNXXrnFmEykQXOwy6uoz39rptuZJSBabFMeALjNU7Mz+
2FQB6GCdZ6PZ2ZXIbGMf8YM7FWAWCfS+GkEIwZMrDdW/olDTACR6aYaP2Kywzki3Bf+udwEHqkEw
gJbbU3M91/0fr47j/0JBVgwVKTDcY/kQaDyXwWQm0ipfavLDRpfXFPJEuA62a5kzgxWBzbyyMTl9
vz8DHN63f6QOIwFw5f2mA23XwCHn6Acl+8pytfCj6Urqpz75//TBr+Gvvrkdh5/05+kQEU9xVEDc
4s/FMrSQmnIxxa3J2W2SIUFRMFSDeFLrf3kQbfkxCJRm0J6vd54EL/yq6TcYEul+4nuRkH2qFmoc
Xz/6ksRmJqIJxciu6XkN3sFwAKrU3jD2DfZiJDWezhfa4UznsYDE+rdSGkLaJuDR8dVHPd8jCblc
QGOHaMFO2lTEqG64OxsQwjBlqUIhBgGNETsnYU8MkfBd0YkkuJfjnZRiNH3OsmkELy6NQ0iCB1PE
8aN/teLTMYuNqQczB0guw3i1o5lEjpPESj1xJxZvEIx/dIrtUTx6rNAC6UrbHmQkyiE4E0ld2k29
fp2UYOJj/JAM0dYS9u+XM8f79Gu5Isz++ItVMABNmbE8VcdNd5su1wWC6KpRHtzQYnz+GvsTUTyp
hsCKMFo6NMGoIeDkecFTLhiWOGsr1V3Cu3+AGj7rO2dC1QTwXRpqyTbhozJVFJzw+MAoui6MaNAQ
4dMITWWxkeYZ+wQvIlfCrg9YcnmBZ3oFwuFTJVmc56hbQv6Xv227wTmHC0u/8JbrkiOsJy6uR373
VjzGTYoo5Q0Vs7wDb86p6tYZoMIFmNdLsybO75k8ckx5R/8vb8bh7XnWZURU6sb16GbmJME1tdoi
N8wP02ks+v1v009Nbov4cTvJexj15rmeMcknK1b+FKjmBU2ZeNhSi4kfFCTmTiOMafcFcW1Is1md
iAiUMSdxb0sZNHJ9zvgNF/kinWDu+60qoKD7NtczJzEsvwZS9aIMer2oIQ+RY7sRZylx1f1R7jET
7dZRh01T1fDYSNI9gsfay7WBTL8tcYVjdl0IJiMS9wYklNdeav4CLQMNdzyXyUvMXXBv0iPgbYLW
FU1j/H9Vdf5wmAwsQelWOerJDeZyzMjZF0eXpcmEiaUNa+oj/j9Uh42+NQzWLKUEdPCsG+wuh494
cydYofiMTD2zImEoUDpjHZyB0boRxhY83wzMWTxzB/OENzhaM0Wy4D84ZWCEOBoM+HgCI99MnEQY
faq3Tb6SLhkiD+mgZyhZgwvfjrjOJvSxzKBoXhhSFuwXimocZ63P1sw6Mf9Bh5U+2VQpB0cVZSyG
w11tNuzLodm8HD9rut/VN83HjYEsRAAJ/898+rm9jgcPouXS17ARBnwl7I4E/Ec4Viy+6bptLaaZ
KDkuRCMq0c6nujNuFy7/tSUSjShvAkkTuiXJwAU729Dg38G6Nl0btcMCYUktbNxN03F+h+zs0L3C
LtHjpe7/44euzsRrW/tsfa/0Vs6YU0fhjW8M6arUKBj+eLPEUin6gcgsh+V6COWNYR7+9o6oCedv
00yx3qPoe44UJT8LYovHVxLXdRzfQsms/qKeFrRhgeeLuGC2J75VR1zghNkxJk/cz+bZceRisC6L
rIl3LV3pMTXW8FRndgidwj5AVW+IkFb9cB8U3rWbqY1DId/h8sMP8DOqiEuCV/T8nqdjXyZ6jOyi
T4drHm6JdLoGG6RkApIDBInM+qxKPzB/m3YQfV4abVsEwG4sTbahhB1sh51OTFZ2N9UhrUIu59f6
pR5sHx4AmJXBk5/KkieEia3ZEYnXovwj+1abv0dhiejRE1S4OzIMkn8ULVx6MjziOJGtR00YM4wa
mMS+Uo7p88NpNUIqX3pihE0alEFXWsT1bux/UTNMh7oNCe9IlSnEy0siM1QIwO/8Ts66J8Ycp3uM
vZXIknkgw8FzzsF/bnBMwhiMutLKREroROayUgAQCSaMdbag+7+IZcuyHfqvPjq7gIWeUQfqREAe
Dp1dit28cmzoSu4w2WvztPlAIxaq4LO5pSxOhDX7zqmytwMNS/1LEdYmKfKCaTvB9MB62j9VBMC0
YZONIV+IJPI9nWExSkCZSdaDxCZm7huiCoFEnbtYrCpPe8tnUVUOLruvLx3MjZGZHWEiQ1h6pFIh
ia7ki3QNwJC9MtqUSA2F/2nf/AnWipJYrCN/Ayovqz0tnJeHmvacwMbp61ORZNyjDTblXXRk4mOK
3XOC0QNWnz5nS3auRMy1lljty6uE8gt5ssFmGAtIcUSvgANM56mBVgVWCWiH86G/S5hK8zLmyD0I
sYRmIg7gpWVLMBnGs1a25oxanRQ7RWQHEBUfGkyF8GWfd2VR1rTSjS2ZgDDh3w/8tJWAlKi4bgfG
FI0jAa21o/mYKxnJf9JeFoV/1l2C5xEwI4zMrR/4jto35jqP2Q4bc5h4Owm5B7pYVN3o7uk2f0Cj
k3zP1jiwkU5BObx/Khg+f830lF5kvZSYgmaYCHJHuFizs++69weYeEchzO/l++lWtfbFc/mTn4St
yk1NlDxLzT/zILWaFPSmsqo1Vxxkcd8hIt1b4l5Lt2NNuoUIh8GfU4jCxXkujMubCrk8R6Qs7J/F
JcEm5vgFpsxENoquCcIWW2fwo1n4DW5BVPYjVFG2WcMBbOyGqet6re48WTO5SYxZ9yeYQ3I/t7dB
+6+au0w5hYeE7K+HbrrN12HJg6RpLXpl4z4ArGTkyYXBURHnEbMLAqiY3n58XfkhXzanqU7UNNSv
LTTpWAT3QoRA3eQgvb3yPE3B8KfXnxdimwAsQ1PYjaRyp9MwSBkcN3lwElgvqiDPsUwlKmPlk0DB
8BxzIuQgw31QDDbwmREqfKtV1x1cFDg/id/inCdkXg4bbApBzwMPbmg0szWr8JBGY75s1YwFmTHk
JQ1sQFPZOPj/XPw1xKu8GMjbPLDOrgvXkacYzItEWyyYZyDZP/nSDzrnGjOa76UFKLBonR/29rMJ
iADFnJUBZ8tBP8nIXxINPCBPOIP9jbpUgiLOe1KgEm4uaImVzb1ABWcI0BllbyAIjwkB4x/Jh5/r
v8fXIKuS+NLOwHWm5hEc9TTwMzClhssvXQl/uxpFb67XyVoqh7RXtwutpGxgzxIU3DY2mriEl5ZR
D2DQ0wBZMTbZNcDpZSswe99PjqI+/MjOUo2BrfAP9g/RpSu78Br73HAFeLl2f8PuExmSezbl5Knr
KTUpr9GcrtRtTp3THtM9BUtyqC71cOFrxb0j3EJEjRS7BZk2o7tUt9T1tWE77M+3xj1qYN/DGfTk
gRNM9Ubfc/jFSUOlC5CWMW0XohGBlZxbGrTk26825iBHHPyv2mRezk/dkRok7PI++3A0e9lLS0aC
ve0i+1FV5I3nMrfIKgkMR7Zjauo6b/N3XU5FF9MQKtxDm0j/40/Mr3C+HSk91sG9p8FV7dpmmYcT
w6b6DJKMkEGZY30TeVvOBZgi1XyinXfBUJrHAkVfCiM6WlnM+bJE0n2jPd8ud/6AKeHdwwrvD2Cw
d3xSQpCXG718qd1rDqC8E+eEA9tFq/tuzJaLPjSD+zPzKFWFMjOWBbIIjOsz+TEAUKNiw8gJ9ZQl
oGHqQRp0fOa2XhsJ7ULvMeTMiiVSDscsmrykYYuUTcrSV9Cmr3zWiEc3xDL+KjiEYTY6dwbEcAQW
6ojUAbFWLZkzGsaIysx0EfytuI0DvRLCEdvCTiJq+BwcoGrhM1UzAfAjtpvmxkBTxJIXRSWtxPyB
qiEtunR0UTgC4NpMYkVgJhwToaQ0GJVlr75SRYRYEPNJX9Ezlm6Md2509WcPgzyFhtahOkuItD8B
dtOo7rQcG5djHpJ9U4GnioOAOu/Jjh6dhjOIPU8bWau3BU3+y7ynEgAV+utONwkphnErs5g6+DUR
/hYAdCmzgbGOF6y84Chz9pABEewYX2DOqCCKofwSPSWM4fLKW+UV2G9xJbXSubVEXsRbKJYy+Qin
vfJQg12nV1pqkWGPFnYCGBPaeIrqUTEPLMfA+2VIvY74U0jmcTmhUHpcI058uipMYpyGBhG9wmEx
Uu+jKuX5PjMlxtC+bdEprL2MiDmLtX/vAvVlAvRd/jG/pojM2sIy8yujcYmKTNJT0kj2Rm9CFJWP
XF3TIsNNZTIpRPido4aq1PRz/X64O4KTAPWz799mL294yRpYsAJT2Iyj28TDw6klMpD85aecyg2s
CCRLVknlP0xx3rjNwYzZinha8JZk4ClUIBCA571n1HGfqIxJm2a25viU2J6Gi1zqCIc46+p792N/
eCZn+39NZRSw+X3/hsBiRvAcSxcwVqQO+7ZIQGAIP7Ml7GyfBwLcesvnna2WwtCVOM2+E0MEde6J
wfwXJdAe4k05GZlnynxUHAAHx9Kc19DZB195tdpSgz04t4Pa8aVxbfzw60YDlFd9tyNqhnAN4jlD
HU6FPVuEzQn31tdXH6URnFyVu5T83psDEgll2pnoxNCVQ7CI+9CV1h7OVnXCW2X/cTeNP19tmf/K
phxawfQWs9lW28NKYuDIX6uOKRNiwXOHKCYwXeeMeAVTT/iwK4qe3S3bWv+zNQ1JirkxDulE6/Bn
TSiFEl8N6q8icIbnDlp8QDJbAuWCB/W0+SnsxMw7NpzR8MPUIeNmnNfd1xTlkTX02THq3M94EJEr
SukBVHwkvVhRcCf/1nBUu+Thpr8MmxHwth57jeGdKncT03YiCM4oN+CpyP7OEup/+QzHVHXe0FUr
CPYXrXx1dJzI7ClivWFUEeo7U+4PEVDZEIMbLDnyz89R4ih8io9XfjtWEpyKYKDT4Ol38xdPwwp+
Ml1uhHk7iYTsHb+Iu+QuhWACcibtQRlhRwVf3Hm3oT5wqRvUTxL1c5ikJCQ5VV9en99m1jxv2MYu
30vxXgdCcaGBIJk2ux5tUbIwpU98AUUea+OBe69Pzbh8ScOT1y1EPgVpkmDu9Y9zUB1R0PssjiUi
FLCy9sjA4YHSGYDKfvzfl6YjR+NIBgQuNytD2BedzCMbPjMJH4vtu5q9DqPqNZryuYh5AIg8TAZn
Z1Gh+64ifrYRJ6KsdkWZwCXRpPqg91X+PENubWchKnhvx2pcXomzF19mj3aJiKYIYdmJW1hXmLHA
d+Ly3PSoboUIWeUgErzy1YTyWu/q/5ZCTQ2Fo42CQW2r2671rPbjFNEwb4cIshUeOR3/4vJl0p/b
DU1Tkg4Cy/mBE5vQjWTCGUczA9u1cvoeP4PE40eEbVqGH2SrFo8voDC7Ad06TKfRpoz7rQDhW9cl
XV7FivMwufzFg/vS5V5v+NAywL8Gt4uvxfXRWKCR3n/aBFwoSDeNLexozlb99vNl8/zlrfL6OI0P
ZPLpv54gwZcKxb8WO9ET5aXirk5VnRBBP47JivV/QfbU3iN/2UxwwZXQRBlZRzjFK+UT90kqBFbc
EoVnHOT70nITrsNdM9Kb0ee85vcCyt9cmVQRV7KA+IIy2cER6SRGr7950Jz8pSspz6cG0uyKO92E
m/1DmnQYeWcyUepwMxVTK3L0ozWXhoI3l1q/bzL555etNw6p8bmC7Yuq0JbMJ3shk0Jpn29zXEDn
xzSLuikJjdEaiNP5YfAWzUYXrjRI18w5W0SyGcokbFpCUqLXhmjLexzyUl2fqQbxOSUNn3UgtqAS
63AGxGhNV+SZL81j2bu26B+Z4hi7qzHgQb5HltEge19JWpoMpjsJM+o5qQE+dR7KKOG/W/c8WFoI
AxplMurONkcco/m9Mr82M7W7CQ0PMXMqldrGVqZ16bOj8FQ0wWEhCwyXogVGNC4rAYNKzX3M7Jfh
D0zj0mwHoBD0jfzSZ/3lbGGZ1xO4kKx//8YtYRbmzJC76fNP9CkDtn3DuoeK5OjM2rLcqEx7mTJA
4hr+08PbIFN/cUOABNSdhFUNQQSYZuA91P4e8WQbqMD/nX22lqEA8BCVfNp7u5zWb0K5TL8ogM67
m1HN5JAy57NLza9PRARS2AgRNCj7/JlxMuTmbHpqIluT+7MzXBobrzeG+eR5Gbt958oNn98cDV8G
T33hUyhHpIUHtsRhPIin09eesC991ACyM5gYppssn+/frrWp8ZvoaD6l/WmxnofVnMrcNCirvGd7
PUBzoGVBBgHuEEe6hEXjAodaNxYJXHmjvG8gVDq8ATW5CMvIOyeY0URp0wWgJvCphZkWAKsFsPfP
0xx83Z6XrkhKGEsRbMR7SDYRH+SrHAyqkGtCI6hssv943bF6SYqZal/Z4HMf/NZfd3sQUF+FTFw+
QvPXKeWWAKs0dvYCAC+3Bsr+2iwB8kqq/2wR5fUYYJln98O7zTViFu7QOUC5lP0/kkAJvgt4z1WL
30TR591uibi6gGYiy+yK9btPKTaRh9thYqHNsLMTpM2bjVGEzdJU6IEXXnJlcdgxHz6FvFpG6luN
WQovpKIgJ+pjLjnJJ2Oz262EZPoH1sh+epdcrTWfFIC4lWXCq5o2xPmFWgOrlUJeJ91IRsBZo4id
ye8ayMBkLRzw1DfjdC6pTywhedb5kSteP8pH6rdiNujyyKM4f+dmA1epZEyaJHKkC0jhVLWc5ntM
66IMr4WrNGpldOHmCpe6DsONVfXgXI2NgYXypaXYK2H5g396bmldy7qXb+Cxeo2ZFVHtCzcPc9Zu
RM3xQOGHTM6q7w1nVnajsVljky85Vl/G5g5rvLuLVVibHTW3u6nhFXGqPBLt/bNV7QYPP+BLSrQs
asrCkzs77nJsTbxSC2R0SysDUYqkNjYGfm+aDeYHSPJIVYUUHJzauIq9ZVhCMyg/UdCd6C/+sbel
X+VDc8jBvwZ1Un7R0oGemu2PQt5BdrL8KoKotNOPTH3e0pgGYZ3X9v/NbX7wHugSdYYGNNGY8a+F
1yoLl9DWD4z1CDUwx9GpTBdBg8a9dt1b1rDd/eyMf2k1hFj2jJImacGd+yiYbN2fKdTwtxmgOF86
xb7VypwxmneVCAD46/wjnSCEKD5tTrZksMSXcHvuqbkFxkKzyJNz1uI38I1QnkSmCcPK+CEOlh5j
mFihtfU45COWEVRYAL7NN559X0yBmhFV/l3WhfmZmpgZDcA71+XfJvicnSIvoX7wHmGY06m64qq2
750l6YfCJ86GtfYkkRlq8FjlaWcuRbaWCpv3cdJYhjGPRyVzS8kUlAzga5Ro7vQFAMgI839664GY
OxSQiIFuSrvLSlSvZJo1NQFIUbyfZlCkpil+BvT4cumZ59VmHZCUfyXPgDzboV2XcJnWB84f/6uE
lJPEG8bHpleKK8Mauj/Es6kjNrTvzWa+Tw6YUpJ02ZAbZ6Y+3nJLHYgDD6EGWOE4wEzxeK/W5m+6
URe8WDk0IvBBu7QUxJg2Px0RWwHzjeX+q5Sl+5Ty4Cif06UbAF2FZgRVCC3eNHOrRVnZH7Ni5ZTX
VaMKKy3NBbtkHC0qFerZcADpaDDt43DJXjNMlW/lcDNHcz4FOnxYiN/oKjuPkVIQfrbTkkibkIsB
pxX2iJ7i0kT1g5j/Rgm4ZO+YU3eaguiDbXat6cctOFRIOrGwCK8aBN/UlHegwuV0lW29fWrSdBFd
vT3DRBBxfpeewI2wr8256I4CI4OxrzA9CC21tf6Cqi2fEFKFmiUNAyBtQgMrPXjZ2Gi0BFu3YoxL
2cfTfuwePjiKqPeQFppVf/2oHZSSjzXQTAM02nP21p3GS+THEmKPP9RQVKa2IFnjYd/PB88VxU6/
YoME4c+Z8kLtEZPJ0BGcz88/T7NO0fxyrzDTbyVnWdjycI27dk52ZJygch3pZ9CzESqgPkrZvTC2
miu4A8girNUtZ22afH9xq9blflUJjrIA0lGjRpXME9pIJiiaqO0LObRBBBtPspSjzE5Zz3SUuPZ3
RPQtS/OMNWi2vYvgCqXja/j1i8f0AHWmAK4xQDuFEYE++LpIUFcnlrcc5Oa3zBk0jeCA5rlM6lZt
oEEVY+8A6WVD/Rn5mF58O7Xo77SQwCGCH81ombwRtRGz8Cvd41hEe5gQWWzNKwbqxtzObsB5OXOu
EkPsrFgYmKH+3LuqM/FCShTnP7JMo+paRG4Z469AjM/0KIgpz2VgDYYRyCAK25/kBonucilEjMpA
XADYj1m7y3v+yxWUFPZA9stv+XHJq6LzzJpjpVg9rHl5Tg9ZFZOheSheV+51vE3AeoY5ujSxIevf
aueqMknrQ0zljT5v0JAxGKSiW/G+jRMpUGK7VzCoQX+PbDTDGg+C7W02PIZ4VNKxWy3dLOyQVWE+
CgeeXBh/63TyhDXr+4dFI1CHPZHqa6FWsARiePnzAxWNUyQvuIjTY5Se6eU45qjciXtMy7tu5eom
9PDv6n73nH7ZkrDIkWOciF+np04okGg1cohi/KPNjO2fuIPT0B4xNDlF+GXyCYFnYtF3AXR28ahh
bk0TNO7u2a6ez03prK1sB1J94LT2YXJRkrd0YEZ5W8KQdm9OmcWy2txW7jYv35lWzFRx7aUgGOXM
V/caxwqMKf0Ap8At3rVdycEL81+SniXFxf+OGD/Upg8vvACH31VzTfnSY+eYL9zFYZB4359ZkgSa
s9kcA9TVeIp6e66vBFLA2w2Systk6P18ntVo7S4xV15gW83omxYJ9SS+ZIGctW/YCxpHZCfjtyFx
uTvB8w5eM3U0/Dp/UELUk3M/4wNt3nqwVerLNZLcb5/jD24KxRjjn0LZwatsJKigXfftVX49NoG+
CXQWyAJaB1NmjCk6rUKn2u7aT2Jtb+3MW0MYGyLyw/OgdtTNBDXDB0xnW7zYjLuWp4oD8YYQxpe5
asqx1liK9p6Dvy23JxxH1jejKUOeITFX1RjFfin3Ju+wgIwC0aCCQCuFDXOVoeNkCaFe7G5hKPJX
5tiqAT7XthfcOmGykfbmjKpToVrmUEfiqTsBU+KQgyWzLKW1/DAjgJGeE6Po+4gUp5/tI/wXVNmv
NbG2qWK/3U8LpcHM+VgXkPP/ZZpxJkRQuciURtMp0JGWlUXCbxBFMxsxed9Ddydw7ZDECHa7748L
LChQYRPJvVryaSDCARb02gMb3xxTu0ErVttKPne6sVt/wi0qRfH2pIvoqg9ywF54cuhTdmemKqg+
3gny8j43h+W62Vd8MTeQJXefKp1zqeHc4PgXts1U5qRUr8K1PncxKq63Ck2UDAF1N46ch5wkNwhB
iOaj/sgWZKtVaB9c/UUq1CSlqviunBcqdmHubEgzUaZQDWo2Jc8c3Tq/b3g0bGnbzTWAh5yLokZ+
QDtPUmxe66ks5E86ynjg7HclUXx1raMEGx3OnsskQeFWcSC3vP3xS5OhcLw3f8ZTs9OoahIkyAwq
RFf0wm2is8o03qB5Xqtf9C9xuQf57WxuYpLaB8KniSMuF09UDaVOnPR2yh1RhFRSXmwNjqI7vLnf
pencQQX5jEHwITLz/FCAg4NKUdFe8ym/JqMi29MSh3B000C+cTSdBuerYGUJDdN1K4uDc9WsPbJF
5Yuzl7djaAP2dQMpBECwleCd/Ux+e0d8PhwNPiUGTR/EbE5Xq5NIH63QJkZmiLl8jHLMViyP8yxR
Is4AzStznEVhHce9OQwiRqdjb+qHoLrrLrzckpyN70dfxaQ6kViL43187DH5vOYYWGekynTREYTq
S5uIiBI9/UfG8uRIhUvLOrNA/phaXyVsMaSoIcvjEuYBaxyloNMyU6rb8ryf0oUvKTiHBdYSVIXJ
W5qzvfobY9Ak3qZb8/Gp5dQROPeQV+iZWZZ87lnbl79D0PFiNk+QnIdbzJr1gpGWNlsm6FdsmwIo
NRlUeNef45dCGdKkvGmj3Vw11sT1wdyhddLUcqSzp71zo050OwXzNPWpHkAgnitWnv24SO2rdYqR
vubR/Cp9s2kzLVMnHhZcGJNr9rIBxhvgKoeSdYJ2un/Cwd/heM8VRXbIpgRMMR2ILW0bnvEhCDJi
SZm5Uo/uQ3mKNtqNs31oPrtxRIDzcxLvZR+f/n5O6nrDGmHVmvC2EvHkGLucBq4HBdW6tGe7Z3BR
qFfDnDsOj0HzBgstYVp/VPuOskpFpDpELMBRrR5RYksfgIGgdufyuaHbrwpyWoG4brG/bov1CI8h
ynV+2zXDU6Y5HKbkThsLfswqqBi8ho8bJmwH5gF69qmtDhL1T+SR+hpDiiFkkQWgmOBoe8hSkTTz
GD5J/JLUhrWsN1O2O8BO6wP8O0BJFll6T3bUZL9e31RDLnBinhqlISCUBLkO0b8Pawf48KYshdb+
py3nyHhgn9MGjb6kiSBiYutP3BfwX51GFkvJApPBiw6hzIDTtp74O8WzNOeyQh4KNqiMRb6QPs8y
9DTYmWkgdJc/WHHhN6O/C5JPz9FA9yXyXzFoHKIHr6T1B5/NgccT2K/InIC6k4ZVWXbfHGw43OWS
H37c6163AkxSzLl+xjTxyeiGKh+aH8Wp0Dm8YU0tsvIBsFHNwlLzQ54I+N6unGn5+fZ+8b39cA3c
uWreJLp5nI8lGWbwr23zlCDdcpPkPYIiyUFBgMAGyivtyj7Ykxyx7AbQk0+PtJoa7wgykhhu0YWm
HmfREp+OsMLq60ri4Ki0kXecaBYXoSVhcgtcPR72tcVX8QQUZ4V73hccFgh5GSZr3Wx6OUeD10TO
dpmttXAIsntnf9iimeLkXYrWul32o23AR5/X0ilb5SU7LyVueyNo96OgVYkAC5QsGcygQ7d3ruvI
ZWIPSGrFbVS1fg+cbSHUZnftK/my75Cr8zh2JpDupGuNaN779DwPeW+IXBCt6/yqlneqa9Gjjv2W
iFzGclRhImXjCGSTNEsH9FyI/fB6ndvs5VZ0DIGUKQo5Jhyzeyo88IOB/kUzU9bSN2hk8hVthZoC
y2rpIFYXkT3OITDZA5/Zz3w/+EZ0RfIIEI1TPsxl8Awp6wsFxYNqSX6M8H1GeYGQlHkXc/cDP2dF
dusfuH3g8kOtIRELs01B43cnx0sa+jGzS7Q4Bk0bJu5NMLJQKm+493Rhx0o6RQcx0ZSjA9V73rii
Zbbom1ZLIdi7/U836sC8ADpAAzrwNtu+8bMtfPXJEpkMgnyGhNFGvKUoEkewAxcnaUB3gTA72cAQ
mHmJAoK6hqv1ocy2Ddca1etBzruSxBvG9T1fm2i2mMJ9+YZmfvcRRg6RKUAyU1yRUKaoxUMrRuan
Z37/m7C33HnuJtL/h6X3ia/mTiXfJh/dDaq+otpQF9HhjWeaEvx/4OOvJkzfFOskI8h7gyLEgEvZ
MsoTQWYrefE1WAw/TFzPFF4syvZacLUV7lKCoW7QxNknxUp4UhjLa7qtcGaoU/MNIVly9PX2K3cw
YiYNd4Rdvh8fd3vrRmVmelylXJnZxJ3BY07pndWOBe9bkV0dqrP3sLao/VciRslhDVq9aj+97mYi
ei5hdwJcl1gudEHvGWAqA3uxQHqrMF5HFFj6zM6XOugD4JwakJrJvcZ1U7HVsirqBpkEr8pPS2Lm
7HdxmdBOEoyhkQwsHYaGsFMBR+/glBhUSlv+eXLZAixFmta6NEJt9/waKjZ8YtbfffR6Pfl0UjNh
/3NF1zrcydQQP/ZgwJSnPH799td+gntMwb05h003XPtSo3ls97E4OzBPYoiWlzV1wXy9BS1q2fn+
Gxwk1m0xDdQcXUG1/T8PwobwuE85LoW1zmyXHWsmx22RlaPKL831RWYnEeaeuWs/rWuiD3VNqUXy
FofwgqdUzpFw1vHiFye2/1eZV93EfG9zwNfULY4ayAhOhn+EevSA9prGwLxH7jA3godNYFbGFm2u
6nokl0kpQbkoz3XbYjlHecMas5z0CAOjEFaXeQFZduRi9/nLfbHEillfjGlz/qDUVglek2PQJVly
goz4m7CmcsOMp16Y76L5MS7p24mduNCfCv1ATbFdkViPvExsZGX/SOGppwaawAbYAhsmkkWY5w+h
u/weYLQsn1Mpo0fmLB2HjGzennFwlby/MDgljCmiF0UtFZBsPkMUkr68rF5vik0FiHwLjWHoj1tR
nn1qHtNDKQUWGV8h92cGcM5cyfQod3HdEUXqVb27a75iJ2543Q6OwYHV9JWvLNYFo4xDUBRlap4F
cWmNa098ltaYopeVQBbSijN1JPy9v8JBJ75ne/F4Mb6c3Y+C8siLaIiHMVzxjpLcnqw+RHBTDk9Q
rgbBlxE3IZwVXYEptKqC+6PdNqJXNzUGlmv1XmtH/nMTg4XaC98HQalnTyXWtwXTGHa7vk/uoG8o
ABq67sAwNzq45T3SUYOoo69ACVRsNQW5VzbdnVm97XWw4otQchpSXTGWMJhPjUSAfovVpOBcKKGL
fBX5PdF1GU9FGcsSOqJdX2Cd/j+QnqagIzCUvCqblJPLbEOzYYpDvPTcspTyAxuPArCnfDUnQEaO
5xTWfE8V+t1BSgtQq4puDBLWc0sz8/IZMo1HO+qnSgp0Fy7y2gn0M2X7pKbMhuHI4e/FyQZRpDsH
VM4xImyRSaAaEurJFf/26xQpEiXwtuZs+82l1XzsroO6fg/R8qpMiiOkl15Il2RSo/kbwiePYYgA
xIwnaFsGqBMDbhZ7OAwGwW8zyvBlQhyNc6nrIdPTVdZPRp6i26ZOSG7GRfzUgjtuL6gpnFLvp0Dk
oEqkJNNqK4hl8GhRSoUG/7qa4mvbLhUyDSo+HDyIGKQb6gkPyHQkxN/Jlu38Poc4X7ClXMQKuXNU
Rvvx3D7aSGrqBj43iBILtzLCnZIfghhGC4EmHu+51D+6l0G1s288OasseHvzoy4S08zAqLUQVWd3
+gVnpyKnN+4fX/5X/s3G6yY+AoCQ9OAGqLOEkbfD+mtQXIRuoORL/AY8s1OpHnr7IMNAiSz3Hx3B
aLqhQmLAvBWtNy92rAC32W4w6fyI5kUdURWJHTOkJ3h3WUK3v0LI46HbAv4kx/ZJYMskxtVujl6c
Xl/gQmmdkmiZd78I9WN7/3WMd3Yt2yh6/PDLhl5jUwiU/zse5mcNjLposbExgrJiNCtjAwBdVy+P
wvLQhdKCQ1aOsz4uQZpVU7rrNHaHRbPHrWkLdhhRIdpkcODNuW3VEzEJXWxFn+rc6aEC+qpMom1C
/oJqz07T0W17Nzy2CS1YSx5NpJsLU4k7GcXEw3k73KGA9GjLBw80kTv1kYxclxN0FzyUuNSvGmow
191mIgiOpilYQR0Ypdr1HghUtY0sFLf1K4JugDubrc+OKdCDD/dt2mcgvHymfMIn/lolm8H2WW6g
MaEYstP3MWsfpyK9hh5gADLdN1sBFgcbH6L9QxnIbZXqkoTcy4Dt/cXwY2ApSXrcI9V6i5q1wCjh
eEH5I7LJtVZk8eEc5ZXX+TesdC0p6zNJv7HlHVhxosrDgNZBsWfhI9B3NcP8qVAe72Y/3HHRPVK2
KU1ylLT79SwaU542LY1TSX9qyCGx0h6CdBC4ob5QYrxnbJ88AzbdMI7U1X4NErztYpdSth1fjiVE
rDe/f9D5G3aI+Yd+ZR2wZElrhe+LZZp9uPRTVqe3BFTeg0k4GoNPwegx6otWGbNx6bKw26FpXFyd
rSN+2NQhndbXwe3zJPNrtgwiTwvWx31qCVkc7TpVzrz8nyxqJNBL02X7WXBH3WK4szB7oC0eRRn/
APXH6YXk5nfXOb5mXewAKLjC3V+qQM9bB7pYEk2+tu+Yt6G/s4IlLEWpp3m+2mXjZWAEjtfIuuUH
IcWRlQwa2sAVid5dAlKPsD7P8vyXgLy3p2YKAYy//f6hyMjiNdwLg9w7Zyjz/dKA7XOgZy5+258Q
A6SV8ZOmHR539dvzGj5+s3HpKPbQntfsxkOTdwtyc5uvot3jru+zpXe3CqHKO9rUB4nRmmxs+Rjv
4jGr89dyK/wCwXgPQjvXttRGBjlmueKCR1Vur/n/b9KYG0ensS0AZkOP9PXoIEybQOmCQ76ujq6g
OXTupXBl0urGg27k+Mev93VIj2hQAp2s0h20nDHn4F/T6lVAeyBbR8w5CgdlyMNJGCpgc3GByo7o
cFMUhNr5S6FWX7R69ION5tZsYBGYUOVeFP3liQHoYEpGN7QLNssSRGvlTLmSVbXDp4oPh92ldton
wTcAEWfDQnHRkENQU4d7fA6JFxQPrQB0iJwZUvIaMilPR0P9/W7PW8mcC/ZKSncg2TRqgZoowdri
SKwfnFNiEYfPRxWATRc1LAOptf0A49f1cuRVJHF359DOtsZoqb+JqbFjlBpbQ2PjcX+189P1Vqg9
pdZ/yMSg3NJQkKNj5qQXsd4he/TmaQzSVdC2isjsA+sIQES8Vadox7QwIDXRoU8vPWcgpGp4mu77
kaMocMM3Eg+DIw1RVYBi6F3UuxC9tBDYBLGpSBPphvgBkpuwePbjfPuSkg5PJTrfpf303CKm/+qp
rB1L9yV0Mh16NgMxJQwMPHA8lHNnZX/KI1bYM4EaFH5bX83otYA4NIghsqD9Vyqn3sbgTEdgAWGp
eYi313NfJvpxpIJqAyEHunHxC/umeJDbgoLbX5PHZn24JIV1wZ7o/BiqhhUaXUVvtel3RDpfdpy8
3785bt9wDypD13qN2zVYu6BPMA9l7Lq25eJ2js89IgU6/fQxG9n+gDzNctnxhbulhkN0nNsUsL14
9uAgEIyNuv/6Qs4HSbw3U93IBH35yVQCr1kmstXnhOwFVYy5b+YhOErR8LGjLMCi/CYgC4Zsun95
m3hq8T8thQoVPrI6yk4VXU+KiXqW3T75GpFAj7diVQmUmTMH0ihgB9rixSCWTL/YN8yOBL21lwi3
r1uNAabt6GAVftnX8zM6ZG8EY8wUP4MklSLDM5LGsCwsghXsqoVXh2DWOx79cyiVf7xpGgG4x+Bz
Xt7/a5WnSVqAUTpJrIZuicLSzP5C5j2NFCIgrN5j43KBedtoKnA/pPkrTOmvxV4ZHFAln//7xDaB
itudJ+2J6DvtQF3e2t4duMLeFJb8xt3eA5mXS8lJG+e55xoZTygx62usombj1vnQqLlL6TNP7TrJ
+7REGSLsQlmiSDNimpqN6wBElbTgwUJCaHKOLKZ6dso9C3upIl0jhs85SLnsQ84QCZN1em+WKy0Q
a4rw/9R8abMu/PGhU0tO+nJFXNPQVOw8i5jh3XMaDAdgfHvIpjbJXoYyvI9xaP9A9E4KCJiVHK8d
JmDx4ZDg7P7ZjzkJnb+pzZFYStW3k0E/tkAzZPjDO6Tf705FSwDSl4po9yYsUC0Oyj2B9FMZLgSl
618WLia1ESYmBne9r1i4FImLEXaO0svL6w/q4lSAPZmRrCwwga4vo1QPN8+3eAvbeDKS82eFGS/8
qzCiJUSeNzCKUILLYHmpnnO69xK+j6iijLjETzAUKsvEPhGEH8nhkvakEbaGmnfvv87Jy0JgBCDm
7fslw8ct58MQbVnA+RAV94VoA3XBZ8nOI4SGpEGEJVDtGqJWvjTS3QD7hurJk6xXpodtaPedrT31
qpSWGE5kSsPITYgmADZnRQdBc9hp3Vd7ccXxb4hqkaHyCIFQfusWVjj6pNgLIWX6Hcq5e7aY8Del
p5K567DAZnUPUG6wXie/6dvCYlhyIlz+RSUoEle7m/Kh81rNPK1rY2EoEeANkiEskLwKsYmyIJN2
CLzZHG7EYec2wQqLLMBnPJWTUBzt1JgYgdADTYmj7GZre5vZr1mYaBKr2tcAuIQJQ1Ifty/V4hI9
TTTILkguqXZz90fIwD16sfy38O+qKsBSpWI02wvZiF8V+lp+QW2t/WtlqsPVb0Vgg1cCDoWKX7VJ
jEKej6iyJo15YXK7cZrDeIbmQMlzfbHSdiR+p3PCvChgI7BK7STxSO6LpGG7AYe/sUCATOn2wsjf
DHRoNf0Otjuy/hBUWfOHFoFwKVC1lhgg76CwQgzzRhpOespUgkknz7PFwTnm3Z6C5gzCGLWmfZ1Q
qKtD0uyqmynCjObl5mNH3nj3qCoJLUW6BRhua+Q03TdvgFz6SfwDenoMfpp4b5QPUaZLPM6y8ZRZ
a7dvjnZXm2gJAqTdx6HnowF5iMTkCTtTmPN9bI7Ew0BbR7Up7pzLRHkX3wf74W48aoB1NCkoB5M5
sCFcho31JYb2u8ItkwM/6ziFSeJD0AFW1xSn/yZT27TxRJcOhoHfzocQ4GlYpPYT8deaFhVkaunQ
oUiipU/MfGNgAuVsCCXL9PWu/tFN1x20cwfzcO9fz5/3vosD/UhLSQWs+4lIi0q9yd0s3UJ5wVMb
pr6KyplWXSAPPn7Cl7SI8a9G7mmfv7lxiZwK2x4FMOkPiFl/0o8xMGUPv/STR6Ea/Dux3DSk2f0O
/NXcF1hKXGEiQEiUqjgqUTcgAtEWM3RtaNWw3PpzkdUVIlyZJu9fHsCt+tNZ3V8/9Ao3dW/ETjmc
hbusHKEt18rYSRgqQyHNe1ovrOPmg5CK74VEO0JROV3c8sxDaxUPjB5fKymGSPYpLCPbyi5Oqi/Z
wUozsajWyqSPJvGH99v2/GSeKIWxof5Kac0+givxJfUuaMTGCazq1AneG1sO2xWytdLX8/06L87W
A08BvffCQGPI2ug4gT3ISbARunVv6AYGh+zXgED9VI6A/w4cgMB+iRTWNi59EZVhOLBFOjKf5UQ7
BKohjtZX6Q/gJF0JFjOaK5KPoXadn+fdUT/cLXOkQOKqcVlMMbD9miRQJr50Hw07DALLxXF/VAI4
DXfCtzyNZcwTfLaGJHuiUSmyH7VyQf640CYOaoSZGH0IGm3jB5fPqliRf2rkFyv8yR1nRVn0I+7Q
qHVkGQCwXFqXRhmlJFccXfb2iLEmLbLlwQCRXv5yOx21Pg/bZ1iWKM2GyIzAmpho4JY/lQAUW7aC
qA0LlrAZSoQALqeZLZWQORx4mHlXH2II4Y5BK+rFb059SpTYzOB8S8y1BCEciHn+cBn8difSY4e/
0qRHLPLclubq/HyP2wmpg6KRmEk0p2HYamTiXXqxILji5GVbjBqM+xTSnJMKcTVz6SK0a/3mKA8+
eFxYexPc2SM12ziRZtlPaKnmjjwvApc+ZBt/v3TbH3934u497+IWHo02pIW/VcfxXuet0B6ZJtHV
ACpKMAtBWzsdYkSpz7SYkcwvEfRr2iGpeEvaoR9MQKCWlZ1VVamY5mpcXvmaLfea5PV0e0oEg7XM
FHtbg6cdO58+KYMPtpWC8/phAiirab68CUBfKbGnRIu+6goEOOtm6FBFDfOgCCp2P0HibaITAGEo
FwiPaJ0dtvwKYqnKTYRiA909IH8sJE25zoSLlA1Oegy2pXW/aQdKtuc6iE2vJOStHHpTFxdxvgt7
kmqK5OG7OBUC3ThPkdJxoHyoo7W4PtE4480Nee0ht2bzq11Que/T3f1wajDnMjTXjugksps3bt54
ys68B3dB1bDNCMcMifJGs8nhh//ju8mpynQzJFbbVmR214Lfaml3LTSQB3gn9VmkN0fJ6ir0vWrK
EDcg2SNHo6j1L0XmS9HEpFA02iPh0IE43hkK7NYgWJKGYouSoTPJaWFw07vRG1NaGBhlWCeBj4OG
EgC+KM/KBKjTfF/8q8AdSbfoU3OXQUuWM4KoY35FHz7uFWa2bsM5RG5xzdfxg2WDjDJgfgG7xRpw
SGRsP/KFlLAUzqzWbljym2PWJKq69BjUEyIoNi1udqMZ/WSBLJ2hFOxcrJ6MrrlFxMmF6SOgHVUs
9nJpNOOQkvvc79FFYnGHeRvJvWjuv1TaaKqSA+sDAqyOihCu132aiLocT9lNwTR84PK6M8Ye21NF
aLeRBQt/HiUNAVsVnfV3f5VTOb1RrN4lRxikUzwvH+S8xLg0L+qdBKxd8p9pywflV8IJGviwBRG+
VcvdmSpHlKpJKwL3RToPjPGkyRWsHseDdkf0M+ifh9hfZQbC8nkKBrYkoAu/E9dDdUKsDlfKXNNp
43g6nPwqqVS4hKJ96Up7rlo5xHinyynGnDeNE/G0WBU1EZUTzbpQtk9XjV6aXH7vw1E4+vxkTKqX
SMhfgxZZP93EW858e884B72qg4hSo7STHleq+8YWkaqJhTfBacAcxHfhDEqnnVvD4ioffTmdg3rK
IcB7RKCGE/jFcTAyQqWTm9niJ7uEIHwDqa58Iqsz2UTSrA9CShDJy17CObM9HlA/Hq56O8wuwTF4
IyYRqw37OhgBNz8vxxlRPgLkAau0tT8xXHa+ETnS3uEGQjVefL6fcljKnp9Xm+wvPKxRZ/UgXnYz
Rwt7v2MiQ3B8jZH6UCNTvZhBYfWGGRc/igYWKts9sB6MGgLblsG3mXa3BHPuGHLHLukfMkfsLfnx
jQ7a+4ZrSV/juW833+C/5Ta45Z32do4W9jMLYF/L1f6OLrgZSNnz2p1bCbGoO5MTDGOclydq0GR4
+NZb6zKOmzVwu5M46rSRY4hlw1tGRpGUIk8yMx7BOjyynTelu5pCQ+1A0fkEj29/i0RPxVm9an90
C4c3xBMjAmd5kQjGD0m0xlwO29RPwFv2pH2rTrKqfQkkE1nJVIG/cfIjpEn78Asesxd2j/eAbcnM
BETVr3vtSbtqx5ndieVq5eHaXbtRGAoM2CvuOJFQvhLTXDazFCUUrds0LiW3F876WJ6nybOfUldt
I2Et97qk0yyleGhKLycEAlPObjAjVjyUT2r9yhRcS/jwHiWU0U9dtQ8CjqiuLmZirDkd0lX/EoLd
oqfOYChk13cyq4XHVD60LOTp6gj7cIYRUrS8jvytXGadGX1QXtovP2qyE8u2wWdV+7CYZlb42KbN
1PrWVQDCrs9pidwkinToGfutUtsLp9OJUrSf3Dg6kxR+50HB/3SpKGX/Q8THlAeW8ichsB8GF1oM
9mbofEGqZylD5fRpUnyXs3HTtyU9J1qscOP1wWeOU9AzYBRHsMHS9nq972FvhL9BrwcKa/ApETWj
FRRAiINd7GQ4i0+1N/15lLi6YlODIv4IWzuuW1HzWx32pNByrU0i9AJzVDfgW9aC/O4HgbLM59qf
WEK2h7UmLxDH3fgtaUTVTWlR7A/0JoCCk7VlrkYmyeSQyGyH+eW8cPyBeP7PR9XqHtDOj4MEzQRl
1oOrk3NkMMVSd506VDH0sJ01uI10O66XJhxu1f5koONhNgWvnBRu+pbcG/wCMkMbDo4PRsvoHPzT
7s+7Peg+RFv4aDMeeeZjwDfff7TUJKdMbdeNyaEVVrvGHOm+pXbQrfT6aXvndbnAK3O2a5DMO4em
Uvslf9qqrB68LterEW9XcIiGlmLK5f5RYd+4afkSOWTD8EplqdCNN+TwpTKHX+2F+xyW1fTFY3UX
8layWLHD4DmqynuvLiWni2Tw+iXgSJa0apDKpYpbUwDN5amWJYRa0rCtvZfokAKnfnnrVZGmw8yk
WADktbIZKSPIeDEADHEVPGJ9ySVXKPl9EBcXTLk9xT1miaxh1N/UAWTQAzLxHbT9ZtHKpjRPyJen
dNEAoVVz3zl9bSmnc6GOJCX8eOmtPuEXadhembElaKuBxdKN8qtChuwY22QHxIIOFO8oNI4h5hbj
FF3NxpKdRImhWsGFjoIRVD8yBsZJeKBAnRV1kY2iZU7KWYbp/GR5iIBOk6XxM6Pu0TPmzAJxWCOi
7f2J60OQJlvLuZaTmw1od3xcq/7hU6RwDJMV2Dp7fii2xhFc5/TzmTfwtCQ98853d5BvjYkzKO+N
KMGzS0pW17JETLaWLYIhfSUJGvJaoeoabu2NiLY8V5z39MNGfWB+etHS5kdRtXWG7yTpTMhUNta/
WUMNnAJaAfga4lS7ssAQ35lpiodCOJa5VVhDt4nq/oEIbv7H0p/kx1qaI1zshiJMt/3PjkgQhcX3
DKKH+K08/0IP4Dkj2wgm9wO1Eb27WDWzSeSypdS434m+blG8WlTlL1ihh3/GquCStSk2URnk8Yod
VqnDYy8PlWiL1qlRj8zgb4D2wd7pF7teCF6eSa0iKboYnWhnHn5TumYEaxiOHJCmlm3vUQ4K69GZ
Mmqtle23V0W1/l1LuzVY+H1Xo0snfk9QB+4MCUaU/JwtxK2X8GdzwzvAz1pcW9nsV7s6x1W4YOT4
J/tdJhzG388HdinNYSLN8JxgfB71Mv/2E6XFABwlSlnaw6GoOkN9ty+v8qOB2oSgB6tt9e21Nn8R
B+Irk35fwWTqMhGvOrNldcpYcW8837ZR0UjxilDpMoBnHv784brqA8zKj0r4WYEhC7swzOxje2J2
di9BbR51SuqzmJtkj5mFL5AX+n9hSeo/kYuzwgX2kgGZUVmqrrAs7b9ikFbdcdjCa+pWSBQmET3b
A1/Fwg3azYWfocKXblOo3Vgs+EYyz6ufSRlIISaSdtc+th+v3JrnVugWSP/ZlQw1mEtNYdWBECMK
VqqyzzXNzbWc0Nru2K3HPyS2qtcVpuOMxA+9jiIt0l9iBHbF7zryDveCEF8FSlpOBJtvb40FP+lX
L7qGLKJuNXA0Z161pzkk61Dtk1ds13wfc/y7K2U1VA6kOHJ7kHtQux+Vz2GYYb+Vod2upsiPOzxE
bxVUBOInp6GSEZe+gggJhUa19jqosfiFLy6Qdrs1HQ+gUlZJV+tAoWbpD4ki/QDAiGEPAO/khZef
UF4DKxhji4qJy2Hvv3Td6o/gA4GiZ5F9OnhgHyBYnowxGmeXSjVEIcDysO0RCesPuwYsLiyHBD6V
/+FO60/eVjbSVcbxAKz+hWynX4O5QjkeBnHgDSWhlMWThzjAPVUyf/gJdjjIUqoLi1bFwziGSjE/
eNOKDZa2nxqhZGoXBFzNj1q5gjzZBH6M5A2E90PpQG7QpkH1pCQ5pXj7LSndHSeKnA5IVpHD1CZz
yfih1V2Sy38C4fGp7Rs2JMwOeEQRHJkoYSZGL6WBluIBSp7xmFoznFgZEdNBuG+Z0j8Lry2ki8DY
XV7XWCiOHxGXxpMlFzloVE/24mO19GqwFXeEJ2MLiRZ8v1eoGEEFh00/VmDCuPlfx/X/v/cP9Gxy
3EfBcfiG3j9FPdiPdH1FQ3Djt+LPxOSyw45mnixI5jV94flKjU1zKrkfrdAEYTGxYWIUTgqDK4ZH
cXKKJ2qZnq4690prQWFYwZf1GaAeAXAyB6Nxu1kibKkXN51HF6/UzHz0KM/JM3s7VgYlnozDnVqy
mvgS6Ae3fYkeQ7OmQhelfB1Z0CHoZd5LxRc+hqK0CDXmJsGQ6j9zuby6vE2lsOhafr74VAjcNpzH
5u53H+p83cMWRhAx01VRum017Rs2laiBeDw5Z5Gk48vViunBSvA2DWABKYLqjRZOBMH+OmOvoQGL
S7KJXiIqngiK/FR6MAEjKAbK5jCORk8GCyYIHuyFBuOPADbajbkKWurmUcmaR+5c4s2X/SCqjFzr
MC4l4yFYU3ykvceFDPB5/tQEHZBGsBpAcfldj/v7DKvtrqx0spkjbAPzxpVCcVh096WZURPiH8Tn
jiSEXttaR3/WBMwcFTM8Q/WJowkWndNCok0LwZt76yLVHoHTh6I7tKnM1cQntUDd54ligVlLsJN2
n4yN4LjTW6up6cWR039pTGSnfC6r0UX7sy0BEYaFCZ2qi8S6hC1FtxFZ8CPLPsj405L1NDEBqUdu
fggKZf0IcrhLas/JgadG3v9fObHTB2bioTnhxKiRoAk+x5KYNLIoFIvYp8mAA71lKaMnzoGnnaKF
M5em5slKhzJuvr+pyZOBgxQnhp0yK/xxKJBCrOj/etLhGfNCxXkZFglpFtYlREB0brGQaLSswOfm
AM3704J1Vj38P4g4WPSW07eOEcDmLMynhEcfULvgcYOQAroMYGmfajJnyCVJCwl+uaF0kpQl97xI
4bVmgvJoPxaOHc2xVkI4HWKbbwN/KsOq+wwH/8fqh5C5GSlXn7tjV3VPt65vfwtpvmgGQgAvEVAo
l2EhrLg1yg9/pt6IQEpc9F1j23ZEi9LtaUrbUlYP171BsTX1HMbKXYVpyNRW8qlTKB0jRHVgetCh
hEU78gXVr1aDjkyEQz2463Jt0hayGOt5SLbmPSkOxz1SOPpdpxcFihbHlPxlx+RfAR/usqB9vTV/
Ge6X5LiCy5vrD8VojSVAPlIwtxhVfH0CRNtL19F3kgs1yQ1Pu5aEItA2UTpWqs2zTlgPgu5GhacN
vaLGEFC50HcriZIMf8EmsAXgHwFjLEucXca3MnJddYwAcBVkDfRwXzPXvFLDxQoKcexVeY07sr/H
tCZoBBss1tyDx3X30Y8OEBLAVGX1ztMWTRynWrRBKqmyWjH0RPVOGpIy5wCT34YTMwon7uKcaYgO
ShGXfcn0WPiaEtxPR55hDi4HqPhJb5mLxWmpeSFEX/T3HDOuQyKuLArlDe7Gp1JQmuJdwYwLbj9L
FH6O9mKYLsHnjC0XfNga6KMwNuujKmsOLHFVyXhAtKdB/0b4+b6Bj+7ADNhu7E9CktMSgK77BdEe
ZnBqKPxZIZNTsZcb2evApALc/dWi5lT2uY32OjIvzLNtK5Zr1IkFiNKmWf8lAvwqVUWOfb31ewWp
BUAyKgEmc+34lXFvwLVyNupBGa89vqvkTxuAawjWzhCOEgwj0XkJ7ACz8PBEH/fl1m2qyRqC9Xcw
Cq/ZuoIKhFfzfAi4wsYdhIDOJe6tyZVnwa+jEa9imcBTPm1rOgGqIxshEXAmOZKPUu2csAO6ULDd
eyfX+yczkHCvNekzSLLr0WtScGJbdqK2MSBhMrXbw+w/xpEwVAnAd2pTKeTf6n4f4/vQ9LBiKbQa
0dsHuvEbV1F8LXuoC/HEUQAYTAGvSM+auXQKmm1NEoyFL3yBOpwfuTST+URRYvdSMYrUgiUYAnUb
/f1+Z0B0KjmJTVO36zmcimm4qNZy1gSv4qZmYVfLN1MOWoZI9PDrG1KTYuFA2dwFGj/9RecapYqV
15psl14nGDUr7nvRGTun1pQv8FJ40jjc17PblpXW5jC4VBLptPfEpTCBwEelBJP83sDkEY+jKTzj
KnokAKorup6Bs5/MzcbMRuxv/z/J2jQMQsEk8deGVncvL3xUsnqG9HYXAhRzwd0SVEMlnlUWJvXF
rFBCNGw3uhFyENwAMtTxraGDGYEumzQ2xdmMJ3kh7wrUiT/cg+UimgBaVIhSPO+Nz/CHkXs1Widn
scikvDpEVQBUyvZmazQlhz+x+IUZF8nUYlKTF9E0D0nNvAvI8Myd4RJn7zituyOiUydo4DgUlyJv
WUE4YTz82BeHFpAq5rUr2zIKH/eTbNg+2tY8hT9+vRf0I71bpYKAv850ozRe46r5Paur3q+IUlU1
P9TNbb1Cxc6Tv2YE9Ruwoc9cu5cmug9Vorzbek3ugYnSduYVxD6BoKqWoFNNQzLYZ08O/R9jJKyU
bgNkboIq4eD6FCg3HyiQoPJHhTCJoqlscDmSQTSmx/Rqflnr3kjIqGy0yiwZJB3zdpY8OkgqUR+A
PWY4T2fbX+uGHwmSlgOgSBP7VUZKOCVGzKZWQZAhyEHmpSaPIDMNGSRH6kzq4X5bujTD2w2cO5ko
P0Tzwy9TaIAmu8Ka94cZWdrX0T6nAZisjS+JqoYCuvT6YdpMCxtNZ3sWDMhFQ8FBEYU6sWRUaWsP
B5UmxA7dc9JJHa0IjX7UF4ihBEKYMjDnkn3ATPCA4iNLGygsBGds2aNoq41VNGwrNsIFew4DkfGr
QgMDfbGj0ALGM6EcJiq5IUi8rzD1+t7b6W9vgE+N2pbdCSIz5zrxSoIpfQxNDzfDpPUj0ApCN3aJ
7tPged8h4wgaSKJezM4N+ReMBPpzPkuajqU0ywAsok64T61sDKmYJdXpZnmxMQ66Lis+ZWOOxUW5
Ge0dLIU9smenduPcIMkA0ilfqyP6TA8klloeMxvgC2PniSY09wSRGmexgQHbVezwt5ECeFVzUYux
rqi3Bmd9jcLbo/zsZbR+ChTexdSXSrRtDSz6h7RgBV2+v40QEjRLSmi6NZjUsVBtNcTB2BImRc3w
77sn0Q0jA4oi+0BUFfErfmL8x+Gi+L8AXwxE9VAf6C3Xdmb5V+9EXNNqXvJGsmuzx13bLy/rqnQr
vH1FkVvqBdV5xiBX5AH3kCu5yXDE+bPKfH2CVTP8nWifnnSa2KIhN9mjALsat1z9EXAkNK8F46DC
SfNwDbkK9B0w+ai0JVdeyccjrpRTCmhd5xwOTmx/NQ5Yel4Ugup0TZIHiAk/6xrRHHaY4HeK20Fc
5Z+jQ6IKVI/R5HKN3sBDeU+s0zcN3bdmbn4/KN+GdYNUEvAy1ZH+AZeP/C6u0/DJUYvR09qjpUqh
QUFOp4PRnuqIskdae46qg6KZzLAbp5FDI3g8w/ISfX56p2uA4ljY19UlaV33ZTbb3Ul9kAphRU8Y
aa7y8yyJUdI6D3Kb2pluPtxoxge912HYrkHYukFRJGhZymW0MtVlVq+DJt7GKCXt6AlvoiIYNBnY
MgBNUF+U/PCMl/unwqsxf+47BF53k/96SeA1g1B/ak+jbuKySZJ1r06ZUED3v6OepFBf3p7CHi3/
16fn/SukI54VYDkocHhLr4ig8kA5dNSP7s8HTH/iO3V/X1sViKHjeHI7nbZobt75Gg/IfdHlwzdD
SFyN+QyhPMEAGACIWDvb5HFhVwtqjD2UBF9CkjoSDzY266gaKG2opqyVW0htuEaxUk3CusbHLuSv
1mruQ0qwngwCtlxhB2uN0pru325J/+WH2C5bXqxfSrjqhS5U888MrKv41t37QLFOt4cFuRaD0wIa
4Zi3bx6SI2ojFRIDN08JVpaia/Iqoue3C2si9QNA0ppI0QDLzHbZ5UmySyvPJZBmrxfJPxj/JrCw
NdYmNc3wiAHdoH7Mi04wIbN1Iasla2PBQMvI0hi77CgJ1Qa972/v46FPDXysKkryooA2pjMPMp1T
sCx9ICHp7d+qpxnjiolWQ7rJwVbJ2/zolzMMtYX+Icr714dqlXlVbzOjKK+HfHzfMPobhnEwdUc7
qRhPpaThhfDUtEK5ddgZlmtAK0w0Yj6/C9NYoClmdsI6yW6IaIFK7WdCDe3dCIvB9BhW9iMEj+fT
kaIcKxoVGuifMddAcBrZdz3fZLiG8vOcKJAezotYEMFNG+4pXdVkPjtYfAjyqE5A3mnNUh7PF62e
RN76/JFpplJ1luoHQ2p5s6Co4wd9fu0ja0sweMzwmNv7tJBxKZ9qUTQY+wbrwiSv2PleJooEXgzK
JfQbJoatreJXQJcLVMTyPQVK7F1XFCJ2vJz+eUlNQBEfbOmMI64GMTA/yAFT/T5S8TSIB3EH5VTq
Tk6iRtpqwJf9/yTg2bR8hZgbsKaaYy3kaaJZsqqvphytyZ/oHPS/GTLskdSV+/Iozj2owrTsBonK
h6sCjRXKkaHKJhQ2EkE7ymG5E38pEIAUtd00jQ9DOOUORPK0tfCTWgBUfNh8s19OmclnFtXkyZWN
+jt4lCzrnJVqz89ijGRH2wOobLo+npJa7S11pmilNFvuewBV0nElW05BgkXJzox10Ls211fb0VsK
b3nfaRdKzzqG+KE4LWi5a9Um7TTQz+VN8QlU8I86jU0tB3r/fdYEJrFbNVMDSY/9+lzEzwr7dUNC
9Nt4rmTr/VZCgIrMsWhDJI6N21X1oNeBkOESoxBG9BaJ3+4Fvl+q0cA2V7pJ+iAF5sqz2EuhHcsK
yrykb4PRbIz+C+WpH4PdYPG35co4m0u78D+xRFqqBaBBulMGEwSBRv8wweo8k34YxBfKSdaEW682
37CgBDKDmEEm/yO/vB5mis+trTwdIGWU2fgMTDeO/QgCrpdHgG0K3ZAion/BpeXCUquR/QtQCbzr
0JoqRr9ASUM7dxbOC3hewhNMD7qvMje9gnTUBvRdi8mGbbK1ISUrTNOSLRE6II9B7cnZZNVk02AJ
Adl4+4WSAUNLttZ3V7jyaezheGd3JFpP9hKGoqoEZFZCFDrS0/NhYl8YSk7z2SOMqx7UonHzu57t
47hznEZ1vbgDTp7MGtdR1qaca+ZwpPYD9VF++TpmzetC+tIR6yIo532unmQK+lLVz2ryCjW9yMXK
lSBb4koGXDT4IWOb96ye4AjeLO7jhYqYQhRPY9VBuYzIQfiFnCjMAeJVsLB8vo/MWtjaY2NzqAms
Y3igNK9kg37DiqzJ8BFUKLSOAr9qLU+bC+T37mS2SauEsWZI4iU3IRh/PNmZ2jBSP9QH0sw6Hpfr
J/orSyH3fNoETS6HZfxsLWoqL0B68U8f0RbQRViTleA/RGlBxI3ogfw5EfWcLf69RItG52giJm7S
a2tOoZMSTc439abNh96MmvNJd1D8Pj9hTxVK+njoLY9dZPx+81mgAkfK+L9TKChSTVGPZ5FvE/Ds
+7/4exw/kAu24ceCI3FpvkIujkfTXQxtkk1T4DaKF2UhKMPjnEgSiOFGTztKtclc8z41WMmqQ+//
VqvR7NIuPywCiIC9Q1iACquKxw1Rr/eFEhfqlZRxy+EttFayEFKyIFx5sS6Ds9S2URekue8m6zlj
HzhBY/x25iFRhf6AO3SY/y0S4tNM2tMLWLINihHdY7a0FPiQe1ua4Sk1djq8eiMl07aaPEFGZX2m
GjJKVQxQJOoRjeYT99p/h0WIkb6HEEmFO1CPB/Zp/q7DfVPDBeBbEIDMeb5prcaSLhDq/ofSvGgG
cnHSLWFjMpTFdW38XW3e1p+rwfqVK4Y0OQppKhICmwHoEduhOtj4Qoqvaijb2eSfUFm7ssu56mw9
rpb8f8Izw2Sq9icMUn7PQkvGwdwwl5AVUpvWP3KQJ1fyCNi3wwjczM8oYH0giSSMnL5TvADGIk1i
AqqluFGhRzaip8HQ66OqhEk9UOG5uhJrTNgwDin1aAhE4Dr4yXfsCfLb9HfBiBPHGNaEyw/eqfrU
Ivo/B5qGGBhUfxhWMPvIJGJ+hO6PeHySEaHLars/vulmi6UjAyESxG7l3EJd/faJ/AXDoPsfCFdw
MRXEtDRg/YDwiY+3Ta196Q8IYvwTvYPPDKB+IP8VZD7pvmeTBTl9e9mp6GE18KsmMf3K6FOAk8U+
30cZ6JmPKGC6N98vRf/Xu9U3HHz79SkC/Iq9q8CuYDgi6BEdkc6uoehQmZkIq+loGUA8jEdgUF74
Xyy57PrmxUsiaL0LLy7KnUL/nig5faGOXo2+7kWfHBakZADbEQDnklmLFaa4mZ6DKqk9oyCMNu3f
HVrg0N0x9YxB7KUr96Rgz9Ix4/Y2P1MnJwX9tiIkq9NdJz3GbVNvbIedzXIZP0kKx+uGWUAJCdWE
Ivv/ZikFO2ecU+wsVq0tskPQZ2rA9y/Vb86LjkiZ3ceoB/Qh3vQDtXpH9iSkVCPVXNXSe5qcpNkv
NxNPGtlEg9kjwNGtJKNzRtTAn59rutH2cVtDtMb3dLt45Owm5ZS0k6CylAY2b7EWUbdmbihveips
HLL3ERnaegxxwAzrXvBn1Uj/YzAdmZ1M12zgSEqbdSG9S1hzTJo/cfxp/eAaDu+dg8IZmYRCtDNO
mj2IwhiostGIrYWGIviSu9k8QmkJEGibZaiNF8vwUBrAwaRKkBWm3Y0KbVqiOokc1nlqqrKRLtL6
olEq2JeWQSKJ5K860TA5JJYKkdCW1X5e/hS2+W7WjLZLs4F1oWbGBcrW1/9jw2gE/Ut42cb7NJc7
OgupKnkD+mu8mUxeUuuy9qW7kX3snC61FsEdrfpaWHOJV0t/89AUF2vN0eWrd0awI0rZS113PcJQ
pLF7Xg4e1oYkCjX3uaJI0R2K0kmVsDRH//c7jNyhYuzqZN6FEYMmwWamECKn48Js2uy/P8K6mYMq
ac7laVf4MpzVRDbzxWdqPJGNmuwl8Fsp/yybR+HtEZliF6Sys4CqoeMBqmYAAwwF9+dA8q5kW0Ti
XyOFKIE4B3DQSYg6rtlZ1EG3LczE7bPOeOgLA7v2QOn/lHHx2Ha2GLKyk7v/eybNdlHS+ccasbUR
+7ElPFxuWL7BlBmcXR6jxE/5hvYWaSK0rP6p1m8MuiIK6eoCnFiEwKfrGMVpdjVu6bc+QyXfXr4q
0N6fPA2Y7KojdtUcjzofmP/lREuUNCTRT2ypTRUgLZBn26vq5dV2eMm0cbGeJSVpc5dxozwUpG/K
UwOIbjTb1h2cVMvEkmoe3ocug8cV6py3rH6AnXO7KC9J8My40IbMch4tdJVQY7hdNOFW6n+3MrH2
3zqG/V4VA+86js/GIZg+5dQbqh62vxMiPIXWJB60U0TZP5CWNC5goM29xj1uSxU4pL0ysw6CV6nN
ifZFW0yOWyiN7fsHemsAO8nuQf/CQcRU2yAyr8oJ3rp29xRWqio2BGvsZHn4WJUv3tmaUFY5RcQ6
4654HqJkAC0qBxZT+0JlEX/5mm23DQjem29LvqlnNr4Ek56o22tTw8tAXeyfEM/uDrVcU6yHjWju
mHL3JJgGvePbDq4QNJRjhhBVmAZSLv47iXNTwiJHFoo/VosAk+jhzHEr/ow9YXT7ZqTKfS1Vj0Yy
Bgd0mwBg7exEDzuum5Ur7TbPOSPeUuvPCQk9E33Oml/7vyTzzNLcS5+VecvmgsmhaXhG1dWcFERk
ca+71xW3lnYS4/Me4yxPYqohT14kIhucsPhXd+QV8CKrQKL276Y9cz/ybWTGi2JrJnf041phLAqE
NukiiJcFXhroCKtfvC7RrvZu/eS9N6x5JMKatrejIZKYfn7jYDR/H2tHH05bSqy5MnAaKwOeORSU
6ZbXmWwUgPB7dpMv+ZOT0mz9QRqiCm6ei6UimwVDKakq/Iuc4BwQfGsHwm5piiSJfbX5z4c3nqQb
tdiiAG+eR2t5nGFf/C6Tu2ozqJiexLC5morMcQdLuj25V0jG5dR7szSmREO1ihZHD5toubQ6EH+E
z9AGeTlgbta15QkWbp41QK3tswtSh+1rvV2+XLEuhY6CJInGO9SinYWH8f7GQj8dTIehHzVmRong
eHP6HMEd1nRQcjKHqJvizA/d38YpV5QFxeGxFb9aCV6fGujIBLzmgZ+cdUhO1inmGcXV7e5g3I9H
OWUXKy8gCOSW963c4eW4m/ImPkRFB6eWbZweUayUno0gD0bZqVIrJOIMwqyomWOfZ1Nu9L2iE1iZ
UJ5yPyG44Atpf9xrwLO9G20W0RE9+WwcRo3i2H1XYs0TQwGIt8GgZjbO6kGbxHnDoMfzU9dlRzyk
pHnqhhDHWLjgsyLHN8lcvg72OeF6dBpVPvVISz6QPts65cIb/VwRHKczwUATMMYPrd36gxI4A+kf
mGLYldR9O4z/l/Pvg0epWw1+POWGMzIYnt3hvcJ/TAKCWJ7+x0KV88ZDLEUMPXn9JnmJ7utfahb2
bhGoAIybR74sG2Pa24VE8Ld6ncZHQ9xywivExAZlSsItAuzuv8/QxUo8pEAehOTRd2fVhPY6heSn
LLGPCuM6kiK2I10eEwQx0IDleXScBg6tFzBinYmBp/AZKu8kuMVQ7se3W9JwsH4iCnPcxK2/tMQ0
aSIP01etAcMDmV3VKbYBa9wbosgBMurv1ODeN8gO3l++vKrwQ3Agip7HDU6Qzi0V1lI8iYbgJMa3
V8vjV5VWLK1k0K4g3qtRxu06+RwtH4pNwn3YpF7IamNluAKg7T26au+LnTZ1lGskmXszvm2IwSkY
gj21YOlzmGvWoqr6zWfQMZz81mpWBZicVcZAz4MMDi0yWPt/S9XmyYtXR7ZNeRPR2mTYnF/CfQtV
a6Z7vHOQbtlv1Z99X//qSgIyDGNWZs4wtuOrL0u+3QxI8+eDuQhuZlIRqcBSDnrCT9irAZ1VAktI
1uJH8qEZ0TSgaMlJZg/vpdXx7uDFWa0c0k3yUwZWnIUS6L4Ye5aYbFJNITnM0zypRzxxkL0727x+
NvR7ICL674YAs4L8lgGQyJupE0J2QLpEbiYjcEP6Ten9vCjvhqrg1y6ZNxYdS7MJvJTqPy50P0Lf
D5Og9h8jIUiUXzsMxYDdcSx3/em7SZzDN9M84aHaiCV4oQLCviPrjnVWs5Y7xY3/s1k0XhaeKIUG
0hQaF2cER9Jkjf7yu1lQd6MQ+o9YJRjZXznnY6ZLpiHC1YRKFqB1F8g1Mtf1Ibdr79uD7yHW2X/6
ZSpKCghaGvGxBT7lKp3e7o0bCtnlI9eId393dK+BjtIBowDNJFI2/ka15+1ZnfCkYzmtyaky18N+
6aUrVcJnauxCO2IGi2FCyanG5WV60k/O0XkhT6Paa0mgKZueIq6KtcuEXETYPfkOZo0jZiNfB5l0
iBECp8qp8g0n/j13LslFjKKQ8y9d8jNDBXCWsv3cYIzYCSHEtRXbeBjAPs6ggEBrOBX6WjiqqAYS
ndtYeGFBBRBPovUodCTGoTQEYZOT9IdEfSpOU/m7IcvyM+HaKN4UMeT1/h5ynwWCUHjfLvCGPsqs
dOxZtuUp0yZAkT7Tv+0t1TA+kNT8A4OUyyq7c0yOrnhnzxQk4TurwXVoYTM1l0nMjTk74Sb9BJaO
/Xu21T3mfAtap1rFtv2WmyzfkAK/2+V726epD+RLpkGsSORX//01BEN94m7cdeLqodSdi0Djqoov
PVTxasZiLyPLIrqiMXP9WiBRT/4WyDX419jRmdEn0fpFxqH97QAMJ+/R+euhYizsDbOY7mW65SL4
ErnhGZ6z4JtR84W3d/6IsfcTlqx1R3x+DhppXl+yqPHLXcmoj3Dc34v/+qsTZRTefFgQ9bUZ0jrH
jJs9eThkt2Rc5lXAi3TKlxhR0pzRispCkFFc7fghCL+wjqXiMCtZJ+/Ay9Zv548Pf68v0ft+dTLC
ZJiQ1hDSMpi0P1mP/cOZp4gIWmAsz4QttCviDiCmCYpzcaprGetjLCKSoCadsao88hqzEHTW05gb
xbw2FOopVNPfnWr4t6sQ/FQjeW2X7VFH1gfF5dOiBOO8eLxMzTw8F4k3lok241ubtB/Bv7VIAbGZ
psq4jyHid7Do26xc2WDzKpFxClu19XFyyr+ldZaywYTmjMl0rznlL/qsQmfANYJkZalOAmh4NLS2
aHiI4a6q3Nzg8bAlgaSoj1qec5XyO2nQnLLjFF8lXH6oY+rFjV1lDojFepdxno8YBd+2I4dHaoHs
K8fythcKV8fyXmQ0ZPvT2jMPr2Y82mH72yTrM6CnzbKAB5Bnc2q5grJgdQmhMX3ZKFS53UWFjpsJ
GQXw/wrM6dZM2fAXa0IY4D8DfFJf0+KScZzRIyxk0F3pcsaok1EaOb2sX7pAitWI2RuURBFl2i8b
e09ntnljEEMddJskitIrdRmiBc2TljaV6067r7vZxVJUr6Kx5MwMAVzgAjpOHN/UQqozhmBwF+IY
Ou5WF+9OhmUSQksXoC4gYVwlGQJHPx3TUyLuLsBbPaceJOQBSuT8Bza+niA8ZxheEvcFZ8mSf88k
RfohaWrCeV1yh3+IP6MOiAaqgo3JexfDUpKCd5fXy1OAG3iNgE05m56vvc0zu2waQz2dy4yhqs2d
hwuriCu82Lgeyj3AsuFSa4qHNw+dfSOqE2sTag2xClR/LzjJ46Sx98AdpTHCSHH+35tm3HTPSnZ6
8omHMNhIZ9G5Dn09IeCCozF2yV3841olD30WG2ff4YcR9xzCx7j9gsHvjkPHBuNIJnYjWeU8OdAR
kMgku+RBcEf+ukLagBBaN8zRRx/FjR8H59MIKDFptLnTAEESVOkP4M9/WSEaYBoXZ1K3+IH2U4QT
epQ6th7NH/CgurvVp7nvN6GEyOJSaXOjTo4VmTa0SpchZsVawrVAk7SfqYwMObjrhsYnk4yw0gEt
4lNgkjsmL3ZR904UCIB3tIuxzYhW8TAdTbqe8Acu3zW76DtcQ3mkP0/BuyBn6Hk8x6Icc5ffZ3pD
oGfSu65/BbnMqfEIdeqe3mLRh73kGkswkrCiHVTS1PG33/rPxVFgDyerflIx+RG0/VVM9RiiRTWe
Pp5vv12M9t96u2CzTHJTKa8my8D8cfK/QVRrnqhyFn9WxikoldBt7x5eKtWN0wvB2JvUhBZT9RGy
jlfGfV1BJ/rKmbbkddCkBTj2ZLF9chDtS+HbhuZnnAU18zMITaiHMmPtG74dQnPtXWwiTUOOcOpm
S3GNGMph43A7p4Wp93nBdQeTlPrmNu6eWRXIK5uhF5aqcU/tF3HivR9h2PnHzJ48JWTyeg6+74u+
7diJXrDFGuLSFDE4gDCVRJ0XZFxZfckaXdV0bhgEkX9aPL4bgKuYytbAbdt5EvVm5akZ7X0L5JlM
7YHesaDdCm4tE9tZSLC7O7QHlg7ZTxz1DALm8RMPyUH6NvibOJMZMcJyzrMbGvHcz3u062IfS/6V
YCpNwWvolvipmoBigT0MMQkVahkaHHZxAQQ7TQV4ory6Ye0qkvp7B7FiGsxzvsiBqa4iew+GxZLz
n7E6ZWJHald75Gx9HmmT4G0BO5fnKZkTd29TxEn79L2wEQ+y3cKSzu4Y7nb+D0A9A8rYz96JcnED
F56sPW9o2o/yR2QeNyhRLbwU4Jc16jrq8ptE8xUBmwX3s4ftL6V/zXVpuL0a1/fp4YJ0GLojbZDX
dND6LXspzubD0mA+WpNhhSFGBMTJAhXZKfPaZ8g9Gpgnwb99vO92pvvguL6SwG53LBf1vWIWlOBS
+JH0TZfxmeeY/LCoqhSlcfKYvnsXko6XgH0QggeHAurNou6Hl5hKIqtErrM92vBDsl/vFmNQsD6Q
whhb1/SJwNq4lMR6Y95HPBnSgasXewvLpQB/qZo5Zs7Ig+kWojfR9hfzWB7o6/NqAX2kd3vTX/z4
udItGNpIkB41V7qfLZcGSFaHds4CnISGLE+LD66cHx2sFbeSgvGaTS2QodSxHb2iXCTh9Z/g/UNZ
CI8gyZa9+2guRRhALw6Uc5FiqB2rq08ycaH9irY9VxPwrvtHlK6jaM4aF0Y19i+V5qFKGEJGfSun
j5RVepylZoB56RaJGh5Es+C9iZPO8y5WyOnHwcEtoeLt03xvbWTW1wR1t9yXpwjSWpTt7koKpoOL
39tcHkCSpbAtr7dD9QUEsM73PR4us0JkE0Wpa2KVLDLOC/kC1KqicGwb9BZntAAlT3am3djWePYg
SsCw3NrV3lNt6ZI+XhdnaVfGQK47j1sFWpMODKpIpzd7Lg7CePysXTkHitlIn5wLr/V9K4YKG1yO
eUCTHB7oKwHkwfs1qRkoba6MEQ7r1u3jb4P9Xr2z9uLwzTneAI6sw9j2WSzqZgHQ6xdNBG8bWf9N
cYv/1QqcQJ4bnuGLqH4SHSXBsFqELnnyT0XGLx2JKsh6py70Q31r0SQOv67/PEG58QO8HojNWG2y
mFEAb/s7ozcBhJSQo/Ry1woT63aCBukAdrH8zl8V5gzXcdfU+f6/UhyLvSWpuUgh8v8JK/9WlWzE
6ZmusbhLNlc6fqwlIejkTMObbm+6bCHeVWwQRgDuL9WzZ3I1kcmUR0iiFO83RRrDkqutwPHrfU/5
NyGMNCZ0tN//r2mk//3D1Lx9xWEfsi0toETfET7Re2kNtKWyxDnZF/ykewfBy8C6QV4k9tl6cbes
oNLTNx7XqkUqqX7dMjeYr4/mD/ZVBbn5lLRBMXdfAhrCigHeMLFA4yREjvNG+c0ZamS5m6qeFRTH
Cz6E5qZf7VQyJu55NS8BFJ9fur3OGwx7PfWHPJodQStOexCY3LcLBgqDDLnA3wzPtJw4kVcderom
qLKU2Vk1JD4gpWckVsZcBLumxh/unQUdzTRQIAjEmfgZPOpZVm85Z6KJJESce+6jDTARZsJQ7jEO
Z2mwZpblNSb+uHPy/ODKgdxnsweoY5KmRqLSFOSKRAFxUtYluIvhVna41CZ4Eq8I8M+lMkpRYg5o
s3oqypwigybOvN0bSQREaVGoW8mkkg1ceevw7SK88ID89PbS9c4bqOfqxwkT8hHUSXVv8XLEsD7N
dx02LqjSqOlFIlG+pBiSTPXWo3XSrE+0/LtbIU/FcfcvS7Ssg1NpWQnoHOQtVpXBfm87ByLHlQVU
QnraVgmbAvFybPOXCSgRidPUVizuuItsSJ2EXQhBe4YyOnVInJ6UEN76n81uv2k0hTdmhiLhkPqp
udb1ZvAAdfYsh4yKpoL2HAfif8huMv1tAtrZLCsUjHhPGF7MgwZqee1vI08tJp/LRyT9gMaJIcSD
fBspEA7H5Jk/IQ3Xn/6UoqM8ZnA28OrkY2pZb2w4dANOBcKMfF401pFt+jhLsfxrmxDRH8uzCm4l
+LRbdZfQxcYZ7zj5twHgo/l6FWWYo6FecoXpXAP2D7AXCGvKCuR3yuq6ul0JowtSaAMMSTE3Cg8X
Vm3Z+EMSaefOSBjXiz3PAeINdriJgG8GIYmgS/y7+VsbqxjwzFNv462Sk9lFGjkcJmv7Xk6wW6us
SDgpx4W4O7Jl4lMzP4PIdbMbbBYj7q43qorVNWSPlVQWgA2f5uNro3PisSQvFTWB0zV1onGbLNbN
5MGWCWQU/xbD1/iIMLw94s7cqFWTy5U7qKBcnVuXalc3KcRDqdMVepRXOkHFIs7p9r622clAUu0y
IK3ddoyc750X7wZQkknOXB4BnEhV67mvJJozltPT0UKSMtprEsFfT1dS7eUII4H3BHQLuKVXp1ZD
n/N9u1uEKGPpQIqJeaLrogsi6av1THkA6Q/Jq60plaSKZ1O0TkQuUD7vlEKz7tVzkW77B+ytGa7v
9ZuBd1rafoclUiEQYIdxjsH7yflN2b+I5y10Xot+Tf+q1lsOqHjjTErRMbTvKm6s8d5BkK/0Mzuf
JuAmbtwDJH26PxSaA1YL5+cyF0zx/Un6yVlPx2W8ZT7Xryyho/2NV1T3iKUOtg2dn1m8auuGsJFP
eabqAgkgsnLZpdVThi4ZYMAuYkC2U7ZqWg+WFZ42bADoWJNDtoB33zDatTN1nir2G9heFJZ9lUgL
8B12kh0IXzMzDdpTAjiaciLNSCBqjtOmqS5ndE2NoNenhROvcchSvDKZZI1SylO+TNce6wwMJAQF
XljkEKa/Aw2zipBEFYikr1kBb3SkIWOPRz1yOPDMVsfMhtxelt6NUYWIvFg8c80W6k4RiO4a1Xgu
c2uMHfDfhhbqdVKHHMHlkxfLCRAzJgA9b833sM7dAfBxmOL4XwRY2+KVdg8R6qxscGuuuMqg+aw7
pwJWwQAllJ5Zt/JMRKOFtF+50tjx8uO5zTPAW8gDZHOqGE2qGMDlGmjsLGZ4zrscTTpNmSDgm0E7
Xvn3wPy9aDl0NEVpgDCuq7mmd+y6V86YTnSrNlXeMhur4GNcqtl8y4wWZ2v0GfUZbzG0nBLs1Zmp
tzA/DF44bQ/ixSKR8QwU1AjumrJkP9kKxjOsDD+tFo/KwgOQ80to2N4BcxBRwhAyTj8UY+Ko/iSB
KwB5Wm1NjYDFX2RplqGgFT80CWz5OzX+nGBFFSfWjkvTJqT52YBmY8IYgHmrXIkF3LUISyMCwK4u
qYzlcN5PgrxMytePei8bdt9ub9v5lqkm80vMyy8VgeRt5zJIyCwuFUqFqO+LS1aiwPZpRGMjGwPt
PXSat9RwgQO1SqtWsDGCZCZHJ2aTzwE6Dr7rSzz3M1YZWLmoa8+06Dmbq38SVvsPn2lzw/i7U44Q
hl5NElDB5qkG1+/loCIi45r1ybttMkjuKy46u24V5v/SrtrwaV6319szbwod04jA3lpcg0q+T4mD
ewm1pueeAWl+EpwVHOkJS+ErvHjFzsqR4Stq256AD+F6admibJtBGPF3rl2Lc1bhjK6uu4ND6vBp
vYehop/M7WbXQiPWJEboIsCue75qpNK0yNHY2iQ3QzdVtVIcLaspXGb5xMoh4jIzaCu6KQ3kJQQp
1klEa1UxFjPE9FoDcsH38Iof/oBkm95KELbEvCvJogIU4SVxqo599yeL+iJkP2M9R0Q0ezd4/oae
psxf9niuDchjUbZuNlb72lu2an6srgOZIJeOKWnHhou76INoFdYX879/lYDrS6632uHIZBQV+MPZ
lBWWovzBPM2YNG1OCXepNIGS+rQpNWN0ct+xdkUvllP1nfqjx0ELWGXgvUEDLPyDJ+cTTZBXmliJ
zIMIbq3lUlYu7eb0uQT6oo/eZ7GVOpbtnylPsvgDxiLpibtxTiosxZqmjU0kYiISUOQKd3dMAy98
kfLxpYfLBzfnjAEyTS13gXkfGW/SNHu2QO8P+Z4cWelTpiw8TbbZu7VYok4IImuH+akf95L19WPa
Uv8nNHAFobgJBAt+w25BL39Gy9VynzCwgF05F2fNLhzVp81Dt7/cxThcwPvO9xu5GHDOGPEkZcsu
Q5ZpYGGm8qYWprQCNrqzJ3Jnxv7Be6EXEXLbRRs9hbb2nyS0TihQWcZ4dkI4qJTaKOYT1c72pZJZ
qxXe0K9QKlIED3B6dDg1HFhNTbBaTwOigE8YYpWscI++GzrvVWONH2PLvOHTN1uViWDclduhGzfd
MzSSe0WiuXeiIETb33EQVesiclwm4DGcQBpIHLaV6WrUWn0EglvSpOeYMY783c6G8QelUsihrivY
oXb39c17o0r+xvIlLNAIA/S2szmAS7eYTTWVf4rJw2dMRja/ZS//gjQC/jQXwuUi+YHhIEKKo44a
iqUPGnioaFNgpz5cgcq6N8u8/CLGp5YPVm+8WbT7vCwfEcDzYKur+VcP+zsx94k9rWIyrBnENgVH
mGUMtSPk90I/0eoPRjtOL4ll4td1F+y8KB5hR5OHjI0DoFDSJFu5M03mJwMJ+12zx49qg2tL3pLb
XfdDsIt6KTJK/4a02O9nsJOQu8STJdANk91lTIkgHmCZttZ6LXMscZx7y71uQD7ujotL952GuI9A
4c1xS4xAMsXwT2M+th26kIuxIEIKTSMGGXCTe8bNgekRAUQ859BM0qqsyp1oaiUMrYahTydElD33
clhIYidyB0GnrW+fYB19DEuA9ZlY+6LZKjRKVGN2XH0fvmLm2r6MbtHhnAnQ1ozw/5sdLQtuFPOm
z2WQPqpq1UPUfdrM1g9nn5dLTYcn7mPmC0eCYgmBrGNGKj82B94fj1p6NsmITrYJcIvYBAWEsCIz
iYVQoReeOlXUo8iNIU4pWauZtI2RBbNxNUfLFznMUlmfloOIYOXt9+rLgLGEiYlyxysFHHzB5c/U
kriYGqqHSPeNwPJbxRZhegY7Itr5WHk4aFzWXYQcZCrZoiTJnR6LyEasKjr7n+Y8743LTpNlECQH
SL+s33MDrDz81pVnr/IZchrhRfPyIKOvjDNdUsYdvhG7zJ0ceArQT8dFiVtDu3L+0DmTIUXEfz+X
oYf7Z7vi2kOVPFOXtKM4ENyH4gfgS78OmkNVPnfj85ycp9ddS5AeoPRZs6sLHvVvMt5GW7LP/2Kk
KCnGgLMVQHv9S6BGr7/AtnTncGdpKiWaIIUYaZTHSPwI7ZZH3Vkll/tuiPVpz7PrWTbkVVkw35gQ
TxEGuwUQUd9XvgribyVT8+DCbzzLfO1XFri3hTrv9k/nETnLtLsaNA7ZZSUXBqK0ErX6WDQpiFLm
oDUjWKwylTQoF0Qv6BZCN7a0oe2mM9vARqp9DMDu2o6BfdoVVlEFj2EDYQph02JqQrjPBqFBz2Ou
dsnYHW3AdSxfHlYAUguCtIIKSelYt2a4yNEQYR6u/XS5jhlXEUSPvEI3tjY3NbLMFWtauoelWhBs
k4soSZBQQl5Jkqc2iulEsKxvwtBn37Y6Ht4bg9yVpEfcw09HTkJOaJuAXOyBAkcqrAwwjlR7nfUV
ZefVDfnnWRAVhK+bX5aGeVxbY/D0b+KCCOR7Y8V4Lsp5HwS/9mMfqQJZvp45R4efCG+lxo4KVXi+
WdFEPYUSZg9WkdNNjw7NG7o1eqbLo7ADmAsX03K3TxxENTs3L8H7UP8h7SMKyPkP1tmlNd/B2k/P
sVda+M76tKHdWSfdAeGZSeadtKNMbP2RFQmZhEe4mRNcI/vuUogecaw/S/JaZk32NQRDa8IkSEOd
C5rR/KC9mM/7e5q+BWS+WWPxQKTd4FUeT8Zou9wm37i9TPCMffUBeUlgWOHHjv8EwfgvTszTcjhn
OCrUXpo65RXkvM/tGviXUO87hrYhcD9VR7RmVmbah0vYyS0jvPvHqHJYIksoopRThsHpAF0yotA/
J7J3Ky5i3DwJ9XrcKjjbJ42uJ3fMQ61W906sCSwHZYjKKnVZ77HyiJyeRuV/kRlVCvGOZ15lcxdV
OkVD38dw5nGL59kpzrZ2bBzFnD4Re0z3sxCHhVJb31vWxPgPgUFJmTBti5V+LOP/xJq2WXMcf+Vu
qG5pv+8JutvZgC5Y2ZmAPTlFfpLSOUv+8Lu2FaiX04URXvjSBQDwMeNSQ5NM59vX82A6P7O/vfI1
XWNYi4FtBW0WuE9UbIwEhDbnC50gM93uNL0ShJReNRP1K9lFm+9VBpiYvQtlcg+2cJNmSwxI8TLT
/vhJxxcMPdyIftAZpES0MCX2NhsMur2bzPzEORKmRigzyfo52lJFV9JaS8ibZ95JVUeEELhErfjF
kEku2Zruhfv1jesWtUEiBA43qUZbLPvTJQgbGcCcnQYqVDvUmpaK4F6aYpYAKXg7cSkjdiyM41/W
foXYUxqQK7rCV951sZaSabR+KS/m0zEad9j/IWdmtYIYTdBbCBkTOhbcpz7/41SSSFXzSiZ9IVGG
ydi+KiGsAgjk2txsGRrt+jKezuizp71ODe5PV8fcH9xwTOa5nvkRaianA9/pBiQTp5V0e942izS+
oSaZx2l46YKgnb6jK+wLAAmmycVY2aUxa5qr5IxyekAqF53sEjvGETyez6vKMqBCr08m5TL6tHyo
kiONY8x7pScTfQcVSxwX631SAulj//DOxr2daOiOOc9mr0Ny7YGAmnoceUo1oaYePWu3YtgGPDps
WKDB9P/z2ycLriUO1rkuOJuMyuW7kraf5e6Qf99OBb3+6/JCuDDj1bMLFO/aURouM3nULeVSC+d5
6Jz3p6cVdcD1sOqp6j/2D+qBpldGrRwfKR0qOtcAz7804OWyOqiuBRVNdotmNM1IQF7BFXk/MEXb
3yWkTkYaLd1Jv9PPlLUDIZgVKSwb7WTnq40bksh0WbYxoek53sDPWAB1HFmoUO3dpYx42qZeLnQq
mzt/LwFktU6RjNHPXhtd8W1NOAfd1tVBzToS+JMCsohfzSD/3w9H8bwaETarFvIVneSIh9lqCGy+
ineD0ycbJ7W0X6s5MGbzBwz7HkTeaQk6PjSpz4LKwriE0XbPP482VO7eP+Tmnr3NvsVgL54KNgml
oHEyW6nbtPSfv3ECCemzLTz8j0wcUWNKnEFnZTZQoRV/YAaKp2GiJ6MtsEjsRaNWicYPc8p+DCJ7
myIfx3w23ynIEzfPriRGrSM9itVeMtzJZAXr7Bt2c7q0OLWp2O6QPyeGMSfj/16KL6Xp8KKAzpPz
dn24Uo8ubwYvPbCHju62zRPIksaa3WRN5P5cv4ACQIkSqeR7aCiKvdFLptCifOgoIQi+Ew0SnMM0
eHMAGX/1JPgZIxPYWn6YtOP/E/cio+mwbsYhDQ0JmekFW7Cw+P2VPSncyFo6EcNKtn+vFDei+r/e
U3Y0DAzaQCXgs+Jqa6wbZVyI1gyqz3iFDjlPfeYSki53e/RrtYjwaYrXj1R9DravFla3G1gEaBHj
36hbs8S/GoaT9cIoe9waQCFFW0VwH0ubhh4TJal8hdXp+LlqALgOvpWoxH04IUDPgIS3pKSlN9Hs
h+SMDSoFaXHAjXndMZz0lC6kK4+LeRlsMKzz4+hari/VII0pHrYgmmqAJRbYKsOm0QkGIg1qt9GG
q5GnEdGiZy5FnKzV70d2TGi2g/aZYsgnO/4WBpg9a0KOH2Z3Ta0gclEPQg7sjtajrHEtGO1uqoFO
PYyY2H6G9gyT2cbGy6W/dts2fjMMGEeQSB1OndHt+3ikDSOVss3xKddOy1ygDvsJo21ZsBj6fX/e
Sqoh9bF+PiI6hJ6VMcVIl+7ufSnpNAS0X0duh2TWe/qYgOT0rKfhqxbseLR6qovNWd7EdNxQ8oNm
p5YR20LqnxNaCMu9psZPnZdW5CWz9ysZ4S404Chi5M1KZ1HERNrpfBncF5CNYPHz2NUF3Cc8WorU
T6b2JEsHLVKMUzLlqV5N/GE6Bqt5umewwUea3DyVmFLeqH2ED5t31jNo0+kgUco/SEYEk4MgxuhM
tbBeHKypWUaa3HItGPuYz5oPlHNOC8lmdqsLtkjLTTQnNFk+LvUx0SqHex6/aSCiInAOMkhS1vMi
Jdpa1eASh6d/nKMzp59T7BkqGXEU6oQfatVW/A+BqexVwIiHkQG32YdELC11JvgWKPliEBM7L7pc
JHpD/4rtNtNpievroIVd9+lqt3BALsG/DO13l3MZKuxCypOETMeMM9Lvwg5rDZei1x30sf1tQQmN
ZuJn+gik3mYM570nbDy7FTjB2RfkOu7CscwaTtWItwcuGwvxkhmtciu7Z1kozRuNWB+O/RIJLVO4
psBzgfgkQ1PSqXE/1BYFMnFkmDI1Hw8AdXvCDpkydwEUCwUdc5+rYdc/IuA7wo9woKOMBFG3fbp0
T7FnukrHB2HTRbqulYqQjlPVaUh1uGszWvt8xJGvYc5kvEQSSKAmX1LNPH49i7JztoWWlrueKjZl
ijhn1vzzNaJvSGc5YOLmfZrm1G/HML1V8DfKPZRD5WjjkMVy4sxg06rJYxL2oaLjik5xAU26I2jc
TGsx+3BaLZ5WBxuZJLofIOED1wxh3OniDibGabWJyaeXz1H1JcWm2nzENyChQyzahCVB0gdAvxp7
yviz8qrZAiig+4IAMxtnQw9E3gXDl2cTY+At2H7eeJC8Axl7VrYe9xpjydod3B4CPkzPWCSoIZcg
xEudy19YwVIh9Y62/YL3v/I6WKz5kuEUOTQZu6YMAd45NxePjWpZSIQnQcmB35IYP7LkQ4XDnLM7
VQkrbul51oitGZgLpN+lKKPvIGEUkcPP8OlGwj7QroFarQGVORcsAkMyBjSngkZSS9r3Y35KnCNs
5MBtxixSquOAc3C/BfOnA1s5ZcHSlqf8gooRsxjjGI4v5ZQi0+z+719sF73uEvfYcG38TF1bDCV+
K/5//Z7Hmv/Dp8GPw2Lhl9GosvWKSb/tQA8SQaMwOJY8LRfT1YxLa68WQWOtFO9qNjgYKSOpYn2Q
7rg+hUoI7ofAupsQ7UFTFHvZabWxA49Cc0t9JC1cJFyQYZwHjbuzis7uweaoR7fLS8rx1MJwkuFD
7wfiKgzPvLATDX+cGPojWh/GIZlkVsrnUd3tUfU5J7/3eaShrsqp1rvLcSMTY2qyg1o0KeeHhPJ1
3v9OQ9DKqcicR5EsgB6KJw1l+EoitSrG7QVM38Sl4/MME6hUq3XONkx+QxXtuu9DD2tp8q64031V
L9Dm0YiJvMIZ8nS+opjHTbMGUR6j+FsLHG9+vdhsxiBX8fLyMtuLNcl9LCxKBtPjzD58JMSoOYGy
hMMoeSaAEfgtgyPxBL0kGQCS+6HGd1vy2/TlGCkriMP+lFTUCVUBLF1I2F3p3KuecrW6yTsSbxP3
R9D7rkQhjern0rpt4JId8ZaptLd2WUaPK3kDZ+TQ0ndtEejseMPBJrVrGZ08WctzR2lkwN8xnten
/WhVrWbFB0x5G+Ily2lfdapWzU0sy3N0ogr9B/Va3NHaxzxM1D2PpLxud4psvlskT2s6zpyOJBPR
4rXJabuUHf6ITXvyMbikmLZ8NZSt1GqyIYMPc/UKVorCnlO3hQj36P67qfX5FnNsy+knPvf/yb/E
QeReGdK5AVppUtmh0i865gXXhUTsqikN/9mdZuR0BjDdDITSnQHqfIt2Ga6lG+6be9hfi/W8OQRn
TcbPd2fxwk9CEOTeS8SRzsZR6D3b8Jh2IKobsK2xHsweNGwqa2rqIZl2enLeb0bTn3i1nHMRqjPY
fPhVWHkdD8+tqSx24zlpjZgTKADEaK+xhmotlHhVDO0h7SF8IQJlQadZ0G43hMx9oTayYFI+QaNJ
V9gwxidZCdssPmXeL2js6EesHTfKEitPgoPlATDel37kiaV5SQjCPs+uAArGT4y4R1JTNCb4MOVH
IDPNjkkXgAPHA3o6AGmnFaoDKra5YmHN0SmdWGqs6CfQHfE5km56Rpr5FbI75ziFK0m/oQdyUjp+
ql0bBspi5v9ilShSJXoZYNarAjx4gfsqZh34by1K5ZEboPlfBCo5sy0pDGbhcBoawIJnpHJnHoUw
jrcaSAQupqAOoS4UVPGYpx4/wAzJX6sd6/pMysOIk/PVdfDjJ/qL/QqRx82yDj2SUgW/7YuZE4wq
FtSb/0mTiOvG4X8p0Xb9NVkeWZCASAk2ZynkAdr9VjuYepSk2bQ5zadvfszar7vui7zEmjSOHCkP
pZN7zr3gp6kU2AsvbpJK3o18W6YJPW+WUapf3IrwrWAtFfH7QlIgPTjhaes0pG6FC/VpNORiYyBJ
clZmO3jF2i4/vbCXvPAE/hVoGajzs3+hPe00fyCODYauEXMd9P9nEAwS2FKHMnAMMEEsp9HkfDng
7whJhfUcYIpTA1uZ4zKGCc14uy7p7EphDioS/QX7lqdNzA5FmBJQgAQNEzpbYfay4JiFHrlLrmds
CZ6S6Zo55lbDFTWIMnGH+D4T4ICFTAl7CAaujtDV9YNrHY35ZZWKgelmsG6cQaJwiHYgQQADWOJK
N15NJ0xdI7/1+RokyTIw3658IAOD0LLMXDqHj/QMYSbuA2QGcpi4rJNmLy8itL9rtI1ZQI3eXJ5O
JOYU4zwO5NFOlrmmmo6Qo/e/v4hwgh0irBbn4KSlY1JM0x8eHhLtjKMciWqgqIn4VgoO5dZDnPUI
ukGR1nTlJoGXlZgfF/8KcxUxkL61H3gPiUr/xXAWVN/FnDNlPjD2lJTd93hfIGTfiA7oJb4YlwvX
oG3S8WIn1fcHBLQjJUA5lRQnbcOLDaBCRC2+fQ4Y+tzHY9BLuOji8pm7E8SurQZlieYrvzhe2L5G
S2t9Wj1E8oymVFW97AqMVGpdQpL7ZH5MSgDeehWYOU+94r2Ftizw2qnnefShZQXWeeP0b0GwgB+H
uqUCbHbpFPt8jkwLghr/2VGxKdswmjcRZ30SudCGJA2x5LiIQzAyuXXOoCHeBn+DvCAf1Yg5kcOF
swR1oE4x+8l+PwrZdQ88wroSmn4hWaS4fCzCjHHvtu4RRy8d9DUwr+Uy/lxujNNeQQKOp+Fl30wC
TUr11efdvnEgLAa5tMGt4n2QSFI0GX4lQiDBtm/6HZPcArfRf53jGZwGUreq2/akio+5mgQ7t9PV
e6EccDeO/Szs9h+6eXPTSj+RVbs6C72gAK15L67XnxyI+xxIJ7lC7X0xBT1FczFLO4fLVsFumC9M
rgDCVfDkr4eLujJOHpLjicJW/Ctzqk/izJFlMzRfwkF7OelCfteWUYpLD1bxocncAtsGyodst2tq
Wf/GthZ00zBep+a6hoUKh/qjzvf5MOifwZV5Uy3HkhogBimjjchizLL6pIByCMoxRYh2eidOQCsd
AqaQplI3/AkL9Wne04OKRf0TO+Hsl5Nx584+3vynSKMuw0dLMaGF2YXKqdJEIFagEVqmRnaQ2sUZ
ptMz97qbQWtKveJQSzcYgauebATrirQ0velfjnUXB+2Ixtp/JM7DTsZF1gH8h+xMj70GOM4YHXuj
d5dPG64VjKnwxzIdN/XJMnNbq7hkOCBYPjagXAeTGMFV7hWg5/HJjoxJu9oQpYIlPYCsILEBFU/A
klLUh+oSoj9Hjtb1dzuScJTsm5h3Z9WDYlkuJ96nlqop99GJNuOxWZg1LlvHqaznFvvPEMJynz0J
cOttwHXE0fKOL5X4mF5j+kueX2ebFyTGIIikvLsoQLTgVXnfcwafKN5Js6oWlDPG3f0Sfe/IOu5/
4uEoHj946LISmniYAtYabGirK2QhlbFCvW2CkFOhSSO3MHu+UqhATGZNbpIeLYKcJrR6oM1mE6Vg
HZEEdtXaYD274usz04UInJmm4MlpdbXmZIgWhqaeFmTru85Low0Bb7+PVWBD5MOHscSgqghY1H9N
3h6i00+e9BPh3tgih8xtGDDF3K52Xm6BTVsvHuHmw9qks6UamfaHi9lA9WNR8F7UP7ntVZljcmC8
jTaDbpZnrdueaTEiLOaGxYtMUzg4iRxmxNWrDRrkbDguhks6BncDItuXY/IVcqKtPhaiVuyP9eZc
59pEhLn40LVnHtAoIlJHUX7cZlapfQCgfmg+uDGJCsuW+8APpw8b4tYbKD2Lk62Tast39dREXXbW
DSc/gyYHcVojEdhYTHzKl2eVeujv1UrEAKzdftZK5lBkoWRY0pzyviDZV+7nSXan0yM2Licjg/jM
KJhdHME+tFb9cOHecCkkkb7yO35xP0Xdzsw5byj0NLlU8vMhTSLNaD0U/8YIRbdUGJoDsBtVvBBh
gjgcocksovHo3DmXR7JrHbcsDcEVnRY8SWwo38Sp1z9FeKpg9hBZf7ElrHYOjyR0mn/ti7WXQ453
H908P1tdaMgJiO8miQBwv63RIXiaHtBbkGwuM8IR/Tku3aBfU0mEXoVbWZ+kJuHowrpTXPa0s206
65ZxLXKD+pg+zSNFjyJKU9ANgGNsTnq1cfdStUmRW9KLgej3u+fYOPB+0KHEAQHEXvLlwW59opyX
uFYTiDdZiBbUpp9nTe9qbgswS9FQJTWuJWzzDMgPInfKWZgRIJv/YYQzu9/vQHLaYBsiuqu+n/57
VkuXvy30I7IHiWzT5kcrTJ6+nndY4HB+m9jAeCOT0DjAAwjC1V5dNDhmfIfjxLxn40pLU+aYRgW/
1U1Xx1ffBwLs2wjKTpAVDB8+CqdazKGmK4+QdrwnmwDD8s/PHqu1YHdYxh+y+MN168bprREQ2+Oe
hi5uGMT5/7Hn+HePkOh4SHa17UoZHoZHig0U4yxm0gX09yKEhBDr85tHrCerKGQtRiuOF9PUGYYv
Q5XsnGbgSuOkDBYrXmwED6mh4+qzdnhPA0uSZv7cTimaQ3dvjsqPXxXufBMeR0ONJnC3SqvWG5fg
14KM8wbhNI1f3eU7Ij9ibgt0Qyq4EvVfKqRovlSS3+3gsRwqa2SYBMDjciLfePyzAiH2Cb7jCYrm
ttcjoeV5uCW9pRJhOm8LAhv7oyJoqTxNsEiSJCzWipACBD5njBzw3MASD0fQA1EahL8hxphMDEZB
OKErxmSGMdv0/dDd8QjaZ6rpE3GIQxC44v/uh5nOWEW/k6LSHkce5V5tt7LjThzlml4SAd3pGRFS
Q+9weyRu8ga1mMWoL1ovkS0G6mtrQ8QCfzHL1TiPvZ3981b9D7Fft2Q6CYUY//o5qxGyEIBeN6O/
npAf0LRyaqiFkO7aZ2yq2BUQZEK4imf/mRfYWLTgaisBsHkd0XzEdQjNptf8rRSCl3E5NTDwoRpo
X4yr/ZagB2y5H3Fi0grzjTKEfjwdhhhQxUuS7gY4vnDtg/OJt1nNQx7dWTHqhhiD6zFuIwsoWNOL
Qz7yLkrnhTObqRI7oEsbAP5B0bTYX4K6dUilmZu1eSaypyTBzPW2n4x1UVAEquX59l8IaGFZEk4N
WYnFD0E3ltja60q8eI9mxfkuQ0U6DmCyHDCp1X1pWoBJwPDPwhrssD8cenjlcrXX6AOQOurcxNua
DQuFYiuseMThbvTEsQT8Zyt45r3dKQtcYIulytdY+KH0//WrUACJ+F2NzhFVq5voyMMeAy3OchMl
pwwyvJjfLrALVGaO6BtLoDGNhZsN0VhCdBk+wJSv1tW7N72rTRTivyKiJSxZ0dYSSzftrZyYSJqb
HWZxdmyXP7pLrjHhMffNUvlR0ULS71seoKz9IEH+GM1ujtsYVPV7FtXjkhCIfD4ipA6cgdgE8zHF
UUePkxxOlNDSvZ2rH3DnsotqCY4lR7DmnJRsqA6ipNut6T/mckAdiTsRchB/DjfE2kcVdm7ZIdif
fDc90Hc20zNggU/mPcwKaDw+9SO+oqmokhcRSZq6IatS6cKBUcB3Q+6hjTiyuBQerCwsAsqyII32
7b+OomowSjhheyD8tUUJwt9GKlknnIFjIG2VILXnDvdg8zaydT77quT+eib5ArOPhjhwZW6BH+Aq
UU0D50rcZwbicCGFLk1Bo+po7YtoxLXRLEJoBTVo619j2aaw7pFHudnMJt4fhNHrO1v+NkHgUzH0
iKNbuPVjzaP0hDLw5N4VYQvzXchqVGyByhubmKL9tEFDXm5WZZ5xtlkxcCZp+B/yl/o+Tlgb/JBq
loXNS+8/BuYC0IphuAYz2t1sag5DFtttvHmIA6Gq3gg9y8TUClZwb/OjdoUTxu5/sUkPRDYo89oN
JzCzdHS4PQJ9APpWpEA2DLChLDjqvrsPWQdNn04JGM7p0tGwqWfvgei5lmWYcpoD5uWe3iWmSKJK
oi+00yzSGraL4pESn8PucQayToMUSjLgASNgYXp/pFOu+P8aPy7j25NvNfnTkssAkB5O5oyL8rpP
+U33Yx4vz29GE/H3vOjYo5l14VEd9QPZ2y+EPXbc/Y+YMlIxUr+r8x4cmMA1R1NN8vZjOsRIo1tY
t0qaWu9MI3boE82VM1JGfU6p36MP1j/PAFqO04J7EjavZ2JU9deXshLK1qLE5TFok5i1Lfv8wd2o
JUASj/m/E70BWtWXSPC63THPr3jDNkW1ber3Rel9Sp2yPwAxzh7itw3gxxc0ZivPRnYM9vPEPtF1
gljcUyMwfBI/uKATJXhPYpyddC5D6YEaMPtJfpaB90bBadh3nfPGNymJuabh0e98yrW8RbsLSmWk
RUTBw8PRlA1gUbEHaYZuL1vmUstXFRjDMN2kGatxyTrPU5oqL9hRN7/mWXoquaSM0PO+fy55Hces
IFkmyIo+08tsB7QgdcoN5IaoG3FnihRtvOHSvAOmvslG4hJ+yW6eX3ruvda0AQJXqFza5a8lFrYJ
zIaciMeayo4Ikv98/pMTOBEHmiip36MmbIN7LIHCQ1EUMdXe0Y/qaAYh3E6CDg3+jBbbVhbqpmNu
GOdmUNyTvSjwdESD5QLNVND4IXA1wmLbxuNmScKja9J7/jxNydcMXB2yTDpnxaWIekG8iGSH4Foh
glu8J0d0lsv6iGn6/Gd6/FEge6qBYPiefplVfbnY/rczjWct712QZ4MAVLV2greW9wZWl+OKNYKm
xtMP6UiRTX20IlgbgxWKYMi1MJ+3cho/x4p54euITHhw3DjJd8Rd600HfPij5UbDkl6gSgSEL2cQ
92u5zE8WvDYNp0r7ghRlUVVByD1h5GE5YxHxV5ne3+WaeosfrofjNbsnY6H8cwaDC0oO6bPri+cx
eMOzNzvfLNdy2+9rslhn99dpiwZq2zyVhLV0MxGh/qgMWcxl1c9xeyg4Bq0ABIrPXteR9XaLFLwV
KsSFZHZKNND4KCpHNSxZrnZTRLIdw9DDQsbDMU6gvPhU0u5RQbg/YNMA7QGzgWQpDYRVKxqx9gM5
Z7oiKyKzHeXKPNtSKyHpojlGNjPQ6CftV3wRD1jtdS3VvcxiClY4gkcQwKe/9tcqkn4qMmt1bLdL
m+KKDjpwne9h2rA/xl+IEBwZR1ixeqLuwfgDkQRzzK5Rt/CrenalYG8nX7BqAULhtz+eljDtQfHc
OAC84v24/5LCmebJC737FhUGIIb4Jv3V8RSKX6LNrNfyPv6RQ/8JhG0JhPzCOBrWQRqFGSosYxPk
4MsG3Bhpbcu3eA0M9roCn+0So8TB1dwPz7W0MSCxZNcmOlFyphq/Gg4zf96rCRFzhx36lbyAkG/g
jDF1/vO0rEDcDPx0sTqsadx3Jd92EP/OumuyzJGkswema1JaTYsCogYIIXC4+xOQIT3jc+5OYt38
7nMF/MFgiHvRUsbbAgoRV2N09MXDeo+V2pxmlfvSCUprqwbNkTfierTdZ4fzMikpkYrcYBkWz0K5
VTlTyXwNSk7gT8n3xyAvJd6+RiE88TnuLEoj31DHBLZMfKZ0hb+yGEw5VMMgmhWI42A9H3Kcuz3H
DATg1dkpfiqduRrgZ5/RD6WcVRpLMg7tRa7VZvS9VaE0lMZp78z6jSznU7E8y2ukj81Vj9nmOBwF
pjqpV2aGZKs87xN15hswNp7sRTgVbdr49nB8kqWumLHGlZqTfhjJnPe+JdNhNX5nXK52LOX6YJDT
2tdbstiwC40famt1SpRUse8qmt1Yha1v3Cm/zpK2wKEqHR35Leg4LMavi29Ayaevc/+lkbfmdmWs
marPVcGjLZbSKQBiLEkpzZ10+b/M8tZ+UMB9u8NmihsfI6LtwQb6Ka+mDpxznZ2Hc/et8JM8qRMw
C5IV9QLMzM1dGZczbSy/wO0FXMRwCVy8h2CGMpnYtX/EE+Be0XnumNH52ZuwfqyQuRlbp3OtGtZ9
POK3V30KftM+oUWrIz7nycCHuTq5q1Xc1Zou2pDEJHLeX/bqQFlVlqPUwQdr1vKpk5ljDZLhA9GG
Qu1Ahzq01ID6E/OJ6k8ty3Rk+J18yrKLHcHkZ6yDD/diXxd9zwkpEJ2zOqkLJ1j1z1MrSUbtSeR9
1AIOmDG7N7LGiMGmhZlbrBa8qOnF0lk2urqXjfYd2PM17vFHvKzLqNpapCY6ubrTTbtk9EpAev1g
X+XhOCaBs6/CyShPir9fDMLYzpw6FJz8Wr25SufkSMUhUTFPlzoCVap1gh8favOkMh8AmWnmYn/L
as4Akp79Jv9Bkgvz6gadHaLv7dQxaQ/DdO74jUDMw/CZM/aIezC1MFQ6c9ALKerRzOwON3Pnbxm6
6cxktKZxHMsLzv79HCUnpXM6v48YSrMpXpHfppvt9lqeSgMdnbWfIqFOmDauF7DUEMNbA76w2SNe
IKYlnRiKBMWVQvQZDkpWXdNPB1qwGiLGaRdJfKnQgaBq5tGyYw8BwjmNp8eKT+Jn6PzjeYeZo0mT
GMvGIW+lFDQDutvNYVRwtpSZpcLlgxJ15en14c7XcxOZmrv2EcOES0adZ6pcEvcvzFcSw0G780qV
/bHQgJ7GPZB0OuquW98pj93pHdsG2G6NXb233R/LEqWY9olk3L4SXcYkWbaQAXEjxLSL6qxmrlOF
/ny9qi//md3H8a8ysI/1pAAjYR1f6vS41OxsSdmIpn+RF00qhwvhi23OnzS4Z7Hb2+5DBKUQZxna
ErKFGsNYk6PRStUCnr+b1OjklanOyj2f92Rzne34xdM+Bcr0qhihlwTQ0rZnA2kBLZ+CxFZPykJt
y+zrihaSlJwu6J0KQkjvw9Ax7l/lR4gQSB4stjryGeCAQbfI+3MxknT/o2oyuOAdVVKaoLw1sqEk
DqK3/MtMWMpPZ5v2bI58D3tJVEw4H8bxHCZweYOzDd289b+nfN/MXl0QZ5HXjPmFSSKzOE9EXlsA
L6Be3XvSjjEfHsoNC6grfw7ZBlljuO3cPlTQYBQOZDn+vIEvzc9QZkmouhyRdrzPr9lLdWRlv/ij
qMSL5YTzSVxI8vH/N5EZeRSIJ2FSX2wdidwN3wf+l/MLyvKKwcUe3tIkJdsk9HzT5m+bNsxToYjQ
mNgnf7/UoPxBk748iKWXGR8nNzkYCK40QvtszWF8xJj4xIECg97Rc4CUXVTohSr1/4o41oDx/2yv
FicZ+KihsSDZX0Po6kDO1H9QaPD0vOn+YEGRlfJQWNaR9kZ0PGKgoGa1O1krRhw+cgAHAMhP2qjt
HwFZMrX171xI/VZPnB8UyYczd+abVwkku8Sp9B2F90MvFZI52gWgrUHtQTIe+TL29zTxiO/4GFl+
GDu0L7AZ4c5IkFtnHY+zife+MfwypZu3EsvlVqQMZt6QShn10TARtehXbnbm7M+y9/by7sAibY29
uNYPxukgZp//YVXSNQlK3HKhvy5/qyjcMxNaVGcU+tBrBytZ6XUn7e1QBqDQ4c/a+J2O6U686snU
tXAvsanlxg11QXRmH6QbPOPESaU3puTNgRywB2SIjDdf7r6I8rK22iuNrVxJTJhT0EpnteYj2VUS
OvlHX1qqlPudqYvaViIUsooL/RcloCfEcUzMJL1FU4JQIydxwIXS4Q7xtZpCFZWeXh40sV86mdRN
+BemFau3CncvDaqCJrlsinbGuUu33z34YUpbBApAW0ac5RsjaPY2HorsiwE2d4rbhhjN1J/JMXGU
CjrmcRSXclpR2O/8TrMDxecWnSlM5KAGWVGuaDbwmpwo2HxPCpYzV8kSzvP9GE06wutpJA6Xapvy
41U1lYZilNMLQ1aWVBHq1zTUpktwGAF7PB3b9s0hTip1SofLRhiHs1/upUV5mRX856P8uURoXJSj
ifoScl3kkRqBe0Frsj3BpWJ6OY+7FwhgxLNG5e2cab53nMRnsfeq8ej1rs84hO6ua39/FN1K0uXH
duuUO/IXPjWGr1U3PEZuMVwlsvLVZZSapFbUqfmlrfLSkpqR9EvqLlzTV/ck0OuQxuo2Gf8YhAVX
4BcxtNoDsnBPCLrLwUWuU/iIgcxIkd/dQVqqCeS9WrwFy3BU/ELxNFohjDDfD2Yzdws5yNy4oJEv
5CoZI6Cm2jOpILUkmFo9vNExo/809rf+sdaPQLKDc01YQffTRhS9LiQhVJRIyCpiVCmuPRZVaL3O
bJ1Vpb4dq8+OuySf5L5NGR5ZilmwOWpZoN3pXGRmXg62/VJnRWcTeB4tS13k5vmKPoezh7NuwIRP
vaJ3Ykx/uv25mVFGt9x9zWy04G8Oc9fXwv19hl6rOgLmf8hlZ740oOIpkXApnRU4cV65TkHfaXSX
wvF8oyv3SKGYZaQeOjOkpKyV7LQ1eNJF4LdiDBvs8eQkE4POtDP+jaailj2VHQNSFDqwYK/H6zSZ
CG9PXAxhh1RFy7yyhKQ6qUShgwHMmpybAI72VOFUQDpOYvYCLeBRvDRZmf3ldqOb6PU2HDJwA8I9
EIeyP38teoaDZ0cOCBC0lS78qlXJGRDYqJPGoofQK/tfXOt9H3hKEKV4gFe2/807SU7PFeVaQWWG
aCalulxumFl/mab+R21KtYMeyBf8OCN9RfxPGqd6Y9FHeoBLOX6fvQFcw+Iwrl4GLGXpgBHueBGI
r82p5rCdqsHklRc3lq1eRmgccEkYJClYeMG5stij5tfFH5pjegAXDC4wcm9J7dYWurgLfg4gCkAB
gjA63JBEWdIVrs34Rd+rIfawwmli49pOP2hxpg1GCFVtzv+nikdOVmMGRVkD5KOCUnjEARvFaaeX
fUFy4/ooUVkq5ZbWhE694VocPW9a6oQYE8C4J5VErAf/9fJUAR62I2AWdGffZaUfhH7/OWiN5FqJ
ZAv4UD5x3LhXjAE9frPwFwZcjlJKURQZrUxs4kcNwnJEV8e13Fft9Ag+MFzyu0sgP/wqetJ9i5KG
R/n345WlmaMH3Y8sfuv2wWvrlcEE3kwfcOgVL9gQqZJjYxzx4UY9E0y1mWYX9kyb8DHiUgU64W8b
5Eza1V8to/4Ib5pRikrMPQSD+Y4WMFn5UUOc96b4VGpAlgSVtY7hT2FVX4W+tgawzyA4vBMZh6b0
/C1bhwvUS4BNGK4DpUqBj8GmxfZY7GCPzInWqFduGdMdo6Mv96NpHlK9ll67Gvzx+Uy4S1i+Kxba
nc53Q5TrgZT0O41VT7rbhqmP8HKaWB/fWeXtC57uHhGA/dj4xm54FodzDHo79Ub0zxnBSO6NdjOU
OmmbH7W7qOUxhHyv+/RcMWUoRiZyURCt7otWMRgQGXXZ/YYyRqnYgUwBrJfhqD/1QUyXnpRUmt6A
AQIgNkN/t2+qTV/Hz1BT3OborGTNH7cJ9UGbcbo7V05WxY29AOmpEC1hg9MdIVwcqUhQogSM9qMo
SNR7vDJXBOClak6cQ9+ymkmajqW7rjHsNZoPtfmvp4Bzl3aN90TyIq/PDlIRKIir9R7NbYwH6Nsq
4pvsU4BvGLPIbxBHPuE2GPFX4g1qeEttV50VB0F6mzaeVbTH6r8XMU231QpiE6xrzEmiM1QAdb25
lyJCqO5uAHlGA0204sd12snaVBTUx+vv/H1UxbKBbRfxRGfY5zFbmw66YQBKn8CAl3XxuEhVXXeN
jUradumfV759aY0540v/lTlVEFarskDh47SqgjC8x80BKT/jP2X7bRYWS64WuFVuy3R6G57b8amC
uTYYkskKr2ntk3OrT/HwdPqFs6y8TJ6aTg3ERzBYp8AErsMqyRtRt3WVRI5hyZc7d36neIMYqgEY
MUZ1qWvL+USGIkaFv2VXnIrDG5Dl8qkxr1b9mUcZIIiF6FyWkRMDMXQMeACyAKMc2GxVdqXJ0zHc
8cyQm+wcBBvx5rY4w3aJCBGMUg1HsDEW9rszrYhIjeHG76PQ2kOuUovkNMQCY60tzGGo/8KxNyXv
lteVjlLJIsWyoSr9YvfXCHoIFk3kjbFazTlAYlx6uoAFBmaS9Tn6e8dSUo0680LNYxw5Wsc+Nb1Y
pqge73RlRyn2gla5+RU7MSVJPmvaVYNjeGk00BmtTC8nulXODgfAqNEzzKWkUE7iXf9ttWPTs95O
bYuKwnbP8dpd8MhX+v7RP5B//WDyFoRDyBRDtwE1OoZTu+hEN17RKnihrh1hhYu4t3a4gRoZKL49
jJWNyb/TeEPkrOKozr5qhN6tHfJhiE+3MxAvG5/ieoT+tamHM8c0JV8964Oo5ioe5XtL1c2y8BFt
YUX6I7hcF/ss+vCxjdELNptOFRu0nmH17hsajrYv8eBwY5a3Ie7yiPiS2T4xkVmNN/wfMqf8UjuP
R/1dsqldtXO4VvWOTX/ScupjUEaYlBxmYPrVIzwNDMeUm10tWU/Kdih3nwsg8KwngSMk/TDgyUN/
UpAt6Mva5KriUT2T8mFEPvv4aSbK6S8a4Jl0L+EpSpTis5OEF0sNP3EXu8LBeWSXTHgJNb+tsM/c
T5b1eQU1uDr6kQ/k1TuF5NuWa4UBLupAtrC8V4yNmdC7HanuNCw0iNXVU24zxsPMPXlE0F+Acf5E
Qp3wP52Iizw2X+sQcmB4n3bLC42vYkFW1KS5DjYoO+WQz0yicUhf/UvANQfWXys8we9rzB8k3z+M
stFw48+D5lPlY8VrG3Kx+esSXyq6DFKIAktsraUURm7PfX4ocE2kPJ4wwDZsZVAuDlPYnVs+mfeW
kZ8wKr4YA5JNH6rfYmHnF3tWNK9qxXoaGB8yTRupSOjoityQPRImiwBkBYIxrBB55+j6FT9e2z8s
jtHt1GnK7J3JGvzBrRdzrYOtN6+ER7V8/J5q04dOZIe27+6Ofc7BvVbkEpJIIsEzXI9a+DsH5n9y
ol20Fx0euAWqjlTPfdV+gUSWS+djaJXSS4SvU/lnEgST0g8LocOdo06bbwlbinPJ5o6QbG0Nu6gi
nWyuMGtQSuBWp1dqSzK13ROMDaxJckFV/CF+31JNr/m1gPG3XQA45VsDmCWR+yCw2Vntjxe+aMyu
WKJdpY3qv/uI4KVgprCciJ33vrQXXkt2JSiX6UFBGTmcqnlhMVHx4uRY27VCbvMf9YMwt/dbk+/q
oOuSVqK6GGod5BbOt1Z/PKYigvLgc+UQ/wet7+VsPxo9jQsWp3pSCNMv50qaKI+wqww4JhD4ed0h
yC/2QyxjZvBD7xL4ZDf1k+4tTqjxnYNSaqvEueF6ehQHTAdWqj83sV6IsSw+lZTdLtUPmlAUqz0A
vV+uuVkCQ0AnWpsN5d1+sMMImQKuXRcNSH5+9skI83kT235JhedyiJ+TFMJ3Bq53zLuXnAjtwixp
zj26YlJwAiMU+BgM8vCz7apM1c3h1g8J6xfcXlLFxGx3x6UZ++GTw2uCfIVphBrsATPNxI9maqNV
sg90eYtfxtx7O9dSNOi2E6Gqbmf68B7GwzPRV7Se//XjFAG5/GmMGIHnacBzVLpqOVMoKye9B4Q7
lC9uF4uIOdT5+9OfbUUKboTaMtXumzhTvPtPOOk1qlYrrGheoxEB+GRuOdcAF+XusRjl9v38AZy6
4Zzhav+eaeR37nBOh9PahhT4TSfRL1m/5X6WgplGSX/eA/ssXxB8sO6pFWI+rpackwgFxb94rmtR
mXwq5l56UVCEeXjG0uh1yDB5YVPDaZOISknXejvi1sEJ9HHxXaKTX57p0CVG7Dvv2NWteVXyq5ya
v0tiKYAW4ZNQapYqyrEn9hMA88NgDw6Y9yf69se0EkBC7tyOmctDNfSuXAzGZ6gJnJnXYkoiK90S
AUxnI/oJkMR4gAwd2awBIR6i2Ljw+k6e6c5W8j/bLbeRvu43Wt2FcyNoSdHN5A670EuA0ifB92Lt
Sac1V/ngQW2E8FK3+fRD+0AdfaFwGyCWWKXw0aav7LeZGKJgAL5begYsx1iltIKbZDNR145PGD3l
XSmVrBynrwxRW7vZ93aZCvnb8VtVcvTd6HteYn58K0Fmq7Kt0KVk/DlhgF0Z9pXpedc3GyNPq4kW
MGrRLGha5tlVPQqRXiwbcgXtGWJU6wK677rBI/ApFGR0vvWJu61qWA+L7GtWjKHe20Rou8ygayFv
9pVul5nxbDt/FX0vmfCRV7f835jclXUMmIjFSpKEQAvq0jQRwWXFSJZXB1MUbaqBOvx1SK8OsN2i
LYnbdDjGnmZhz0cYxaUz95oLB4Li2v2/ao8UL9vZ/+2/1Bx1X7c5fTxemGRDHBjolSmFy8IQ+50C
pLmBPS2RrLqHasRvGmUnraVCDj9EkFC7lbxmLw/fMt50X22LLD9qOwtBKP619p65WSEbIFnPrgIx
uhev20hc+d3pFd5MNt6W7ucmpoFCmdT9GyvQEt12Ct+WYO8Sg/5Hz26JYK6ZGGsn6PKAedIVLvy1
OByZ+NMIToSfau3LivLyUaY7ZHCTvd+9SAOQcKmbqwsdp1OcFMjfKCdtDh3mHKrrx64Td8uE5ljm
+Ax0DShBJzk50BAlWtN3BC1pBQHZVBu5/TUGtlvE/syQ9VgXcJOmB21lLRSeA7gOCK8kxN6nReMZ
yaJp7otgEtpO5XkFly+WJv9rrgoifUSIcYVEHR4wmTbnLCA5FqTaGokaGau32iBFfSjKUav7r9uq
qkyjnsbbVWv8hAWArm0TOuhznGJPETvSdUHezkXUOkDsvCnp1Fu7khvt9yf0/WuyIN00ha3DZEUI
HA2LGOYp3GUCNkxFW7zMyWlgj2eDJyzwHYRVTjlbWJHAnksnAS+G4CSFj6BH2c4PNk7B1146lcCa
zxl9ObAVSjgk9G4dlmxSUvRRsMC9x0pnobVgu/mYwwIotP4CCvKWK+eoCO2/XUYRzdC+irBK80dg
02MG4H4kQS9SKqaKAfTeGGbKYisHQVb2w7gF36+6kstPeCSOSLrd3ZYHi2Rn0ntBbpCRzk5Oi6PI
oRfvmEmNEtOij20hnjVEOz2axaP3im2zpC92Vmyp+hLhVi8PZNeCEbqbLC2nm9t3Nbs3zYSq8RpO
gLg7O+FEax3xFrzrXQOyqTAmCbBCg5Zn8QkPWGbbb6mwQwk2dWP9T9D+hbDr+44SLrUJsOgb4BUP
c2ApP4z0RXMHUHtzkYw45oNfzvXZHoiG0hO6BHnQ6FluQCl/r9HFquAyPflXNoMKi4Yx7A7PUtpK
3qqNeCzZPbckLXfUvd/fv7VL8GrHfEJ/Kb1UFwEqMKrqB7qJjVHPi/s6DWEk5ycBgRZtxHP8kXwf
IR+Mo5GPZWzcRu2e3SBYO+p2tbddEWl6ODkHcXVHSTxdwBODeqJzZ0haNJUCTspeDUPKaNKGfIgp
GLUJzRSCfxDlufNLilIoGKPgugmS+rR0Vxdu+1+utNMqLq9YO43+DiJD8RCRvp5ACAOVsYn3iHXu
wyrOflasfp1wZawkGxJ0Ym0MnFuFbdP/AugE1cHM4Dx4vEtm/GMUlQtoCZ8bb6ZKPMDgGH0lg2Wx
zZv60WV/SeTjWHj4egnw2PHohGRhsz8TLmjgEr+xTW6m3Q/2aFma+wwLrBLzwnA1PsBkQ3icvn9d
Vz32X/2+Haz5fsK/LJmvTECsmlkgD0eHCWInZNU+OgNJZvbq0g2qE9O78r1Pq2Ney8Xay6+GwrmW
NDPZNkWRnEdUo62kQZxDb6A7fzppVdPBVHeBaU0Cq3I1tX3yeY2t+J9zjcqywYuFUBDkESJJPOUp
SLpMHKeth3NCwGW8HXbXHAmI/Fh4Kcr9X0zTAEtIOa04Vve2g/h9X7975sj8fQexVBYOSxDBpWXl
NrY4mmS8xVv10h6Fbg4eM/aSeamQdByQCBfxyZVEFuP3HyQZVnmdOXLA46HLid36JDLsqsP60hRG
Z25T4o4I1d4dAmADs+XK3M4OFtnm4EDvcQoID7FKaghwyRM0EDYogI9NmN8zP7U+yps1X5dHkeT6
exGMdgwth8c5gQFiZiMS2lrANNYcxKjB9Z8pbmHxlfY9qWUlzbrzF+nXTPjUk9S4Ww84b3bpPfk4
UtzL3YsHDtyJm5UMn7cZoIWvUZlGTvBq74ISlZ+Pybb3jDjBVi/+SNOBcXL6EoJ+dQ4DKpeM8tSt
rwGBYDCfpsWkTY/IzP6hp4iLNpv6ko3RL5sO3c73e2LKiLz0TmH8yzgqXGiuSRLF9WFZvMXwQyqD
6dbCy7go6NLxWKx0tNMuKF2knI5n0SRRfxA90uZ4HDSEVedmpZU9b2VWYF0e+PdSq3ZnYorshKPA
z+w6JZBYXS5/fEsaLO46EDCX57arDWh6ovdLZd2GGcr721CczODesSpe1VuV5hWu/d//DneJ6MOM
bnEQyRppWCJy0gtKxRjIHA9KSYdiIqT6Rc9sUPifVUxwv2w6xtZh7vNCG2K2J9yC81idYiR2Snd9
oSrE+8DXkK0c33/DTm7VVj0LsWsll4RB5/EolJD3Icry6Z/rGn+KPMR1gWKmLgMizOHZtU8BiFqJ
7bkpjvULVSYHnDFOWCIlXNS1ClJAVzrvnVVHIvTyzKhZEb2yAmxQ04CAbBCCxG2NHh+EsFbfE4+w
wR6hQBeQ4TA2az473L9PgIybBcAcsAMh3Ir+wjaxTmYKgSh4GqRWEdd8Z59S/tlW5CsZGRHF2iel
NKJhLPcpmBljPxZeQUfP4a8ZfhmjV5StjSHO/gIr/907CtT+V1ENJGcUS2iZgyTQUTI0FPR9D0e2
buOd7rOqixR8N7lQsjgrLSKXMdsW3l42vUVhYk3CzWue/JCVCPpVfyIftR24fmC7+B2h6PoXkbMH
FKDfDqdwCpYR2TxtS3Psk8QWGt6Z+THx6l4Gn+SIH9iaRuU0UgciWI4XXCyZpepnBbVYXGolvHC1
QjyNdnp52FKfR5dlWajgL5R5O6ZiIAoy5w1/nEIHMuEyr+BuPTHVAVdhTxUTqFMRpempCZNgUIgz
qS+ViGu3kpiAeyJkzNTGBFdQsz7utpKFsuVkfEUReotGqrneBQRB12+ZPv4715GEWyvvSqC6z5dQ
q4GELtkz3bddmo04L/jJ6lP2UeXp4tagI/Jac0Hx1QFqq7IYhc2dgyvMv6raGBsQyI+AQfRM5y3g
PLLEXYbbXoho+nMk5iIMKxArVM0puFNVbU8idqg7yjMz+2WBW/StmQpKHAx2bzp0i99aDP+ujQlB
XmdLRTDTq0yHfvQ8qwFvt1yyadMOAbE4gtlXo9IXasLmYeem2QIRlQ1UqkhgblH7UrzTvo0bnYct
6q1QUOkdAdvLvWYLj9Uzdm9G4bw2qUZmh/75yyvMV61uKIV62WjU68unKHy2fqM5GpAL9Sta5FfD
giP+huVMp1xyesLlvo1+aXjj223hyMYi+iSHkWRcLaNDriTGKgVjwwbmDFKm28zguFk6tMYazOzL
rNjygs0Jj0DIjZ8M2j2lmKeozHR+lsm9CRKyXlqvX6ro62gm9KjB38wnbq7l5hnns3GG5svgRsWt
hyg0c6nCvQVZaj9Z1fn886g+RXgEDdgZefj5mK7Hqar0g9oS1nWNSI/VlLLQT3qjLt0MipRTwzbm
8CDxWVO/Uzob7W3M9PlJWlVGIlCIkp6B5BeuhX1sBIdG+bQ28ENTMjYhmZHaO7/83HClualEpz/K
tYYt46UP4HKehhzVnZzmo34DBgs4WhmDoP4gFEPuDzqMftYdT2Ls2zyS+tm9/7J9CKUKp8j0THm1
rlhxeavhiLt0+o1wvi8Qe2U3nP/4Yaz0zBAAhA4usY2nDvGtukXd1vmHgO7IaGF8vymz6idtYcac
SIZNaPMhLe3dXjiJxReEcO+CLV2NAnxA5Kt8ecuLvKy9uOne8o3NaJ6TT+/8l3CKIdE05SUU2D11
Jhwr1K/ntrjQy+dmsEA514n7s1fCFMqZtOHJ7jM90nG71j0S8XVkFTv5xMwZlzYnC5KRzSEL78xa
WdTcfyCWOp13a2NUHLfPvSiajcqVkqyATRINmOGKeG4lLDcHXK6DnOEbSTtMQCZRid5Cwepkx9/p
PhhVZjZ3nqp1IXdchWlHUHLiyytVw2D82S+18c3eaokz1Pv6t+TtrTOvdY6+hqPLO/LFc04AGpQi
X860jYQ9kiiiryAuWdoW3jrbkJsSj8wmJ+ZNy6jE3foLzVPZR7bJQz9O8cq5qDezc9d+C8Pmg8SB
dR6UgKsdF0/EV1VnrSPhuXZNN/a04BXJTWI3SWhC5As8nitcq1YOsZ93/QG8tWgjI6qHpkc0plVq
CNsQjEeUY3ckPy62nsxU2H2FJ2UnCDWoithjvz1Szs8wEidGC9fj7kVPeTBO/ex71N9MQU2ydl7R
ZeAwebo/LsCKPJhHYAu98kuKFe7BcBuLhJIjeiOC8Rt7HzBMG7ZXBBnrF5tfv/Z/E652tLHt4I7C
rkmI/txbH1LmKW4aERmcgkGWsyEq20JcPGuaeEQZmADQtO5OwjOSPn0m5pp2AosfzSAJq+EjwSrK
z/xU1rjuc9gQLsLq6KuwBDZYq2tsQOGezQSu8nIvSNb7cUZjg2Rt4OUnnqZZuRFJsHqXx46OCCcd
A4Hx4pZZaGZsknsoaDRh4Ec/Y2WeDkv3obWe+Lgdz/Lf+KVPSPrLS0QonU2EcJ1Tp/Mfj+VT8ZXO
vLSUMaLRKjaRUi2agK4kZG+/N1Tpb0CYjn4Rm1X56NcWna94HiRhxEHLllJESfSChBX6obQgLrsj
RQYIVjfiHRmTkfNKigB+IELsGl4PG2/urpbU8mwyi52Fa1+Bqdx8zHJ3kNXrs4GgRn6j45ZgxnbG
/w2U+7C0LSnlBteUOF40ZR/6x1uOHLNAzwHArLG1J8ltDTkWcVI8A1Y5RTTrbeJYZhGoB10PVvl8
IfqzWU+bkreDEti+0qAUsJriC57Z86tNHbsRho2GUt/gPwFpm+y4et8GaDaVYGmCVwUv/mqXxgcG
EhhAot5bljP8NZO6SU7nEmk6hqwO0cZgSQ+SKz1j21QCwCvRFExUr4XwUoluRjJdZgsgZeVpyby+
5C33i5PzZ3w6vB/n+0gPcgJjEzh2QrF5kU0m9fXAzoADGwkSs3Lqw2Vah9vux+xOsEOH2LxmbbgH
ySXIyWgsCSUVe31QHesJfRNzTCtzz/REZB1a5sd6t4I8LwgQSN6lKrv6pSQIKpI2WP/WnBskh1S/
vYQjzUQCAkRAes2NEZ5FkLtPivM/LQg9mihxsxdHpOzgoG5w2M2Eylvc/YmIgim0rCrWZqDdnUXK
tt2WfBgBQCsR9S8FX7JR3XSQvN8rz/HLyCCY4Nq/R6/Pu3lBpofG2DZBowTNF81troH+YqnxHGLk
MMJv2hkwsCsaPTBFHauHFC+scJHtlWmKCzGSUnumSu1s77eqZCXocV3ZlHn+m0OxNcFH0ejWNcxY
6iZBY/J9BSAUo9jd6FSgm7OZFfXLpyJ8mNyIC6rQDjNvLjE9frbOdDbs5XCTwz1LTSO2/n2Qtzew
cjcMS1PKhjUqxRboHXi6p38sA28ei9qoFofWTuOVcE2pywD9S5uXrL4tDM+oPvjQWYkPvHsNZvNK
5iyF2BnGBp0iGMbcxY2hko5iubUqz62N7/A4xu2SMxFcb+w2CtlQJwDv2BDsE4rSKso0oLcfa584
62IKe1gG9fURwRQ6mskHckaWYgxi+odnATNWuGSJaja0AlHQ4nqRwQHynH3l5S8VIv8hKXZ3jGe2
9Cg9l9MIzWo9AUfHpSalkuDZuuPY0qMJBMQML7UsNHDWUiRdmGbVeap4KmodFupxB6ubAhZ+X/v5
0UCKF0q3vBqdYF+wSNQk4ppuCcwccdz0TtpxXmQL2OY3z4NuYudRNAvIleWhl6z2aLmNj5vSfqvv
Q3JVG/ZCMF3nzJlyg4Tw2AYjROvsw1r3hhVlMkFsxnvMOZPGc3GoqJGrUH5ZYumRjuXxl9rrYoaL
svc6kPjfR324ispvmwWyHvgu71nFtZj4U+S1EQjhDetJvjK8L3QRm1vOJ01MprMrYebThdLWdXOP
L5LrFy6210k8QHRHXiS5XIT/znx3JzV9elWWN9tK2oWYIgg+pjOUAB3Eq23UIKZlkPcp07Lujt53
l4MKSTrtC2ecEI3aCkGcj39zso9FYqehRatxvA7s0MLSGkaBROtCrOnTR94YfsFah+R4NaBdV2QJ
wdIvShd/b60RylW0qeKVg3vAwZlz+C1o/zlS26RyQGfWi529pZRRHbFfwLeQNpTRBw4yVRzZ0dR8
e00Ianh0l9dAP+W9OZjxqd5M0ccW78b+B3GN4UTfVYfASpu3zTx7l2lyP79oNwMqEA1hDfJR9F4z
WOCbfPxN19z/sNry7LX68BPwb4EtWX3qUMqkjJVmh8Lm5snKY2HyNhJ8WEdtJDH2ksXjiN9Ed3Yj
RsUmdacSfWvX1xgp4xAySKROU/4iGem9ArKq6kc+d8/5vOoytymuL1zac/XpUAFeDARtelFL7hww
6NrGiolkE/oydt96Bh50K4ibUAhNskwXDVqWJrqJl82nIgILqZbp4u0ooyBk4bhD/bnL3eFI6hd/
/zylw2pvyk2BUzlUxQRVpMV8/w5LL+16+OkimiHmW/8IDJKGnTwNToCPUjxxT5+npIY3mgPuYYON
2b6PrNiV5mCfv917fnqp2Km2k1pPNvvoLqEuA1DqPuTgkWvO215ohy/8kHaeFiTpuWn/7lIPoBfy
jDpHfkwWEojdqXUS5w0f9+xKpLZl6PPTJpOAA0Io+vMHJuLpD/5nx7bk0KWMYZoIlMhnqz4xnE+C
JaY6aCXPMzq1e8wc6b1CDR+uuh6xYySH3vO5Beow/E9j4HqHFW/OAT/ODTq98tVY86NV50H8nKWy
3eXprTnjgbwopWxbOR8JgROjWyt38L8AjFzxW601iykW/5l/ed6QtjXOjt2fUGEZ706/EW/wgQb+
joefpXR46W9xy5RyW9GgkSt8QG7SISl2lnPxAvlbc8GPBynj3vU4oBlwuMM+EsH4E0HPcUXRcEE2
LOGCXEBh1Ytn4liVIloHK3st3Ne7ufBQvCwpPuFbguYqBuBrf1e0Xw2ixci8URuYpz6YK/Hxkrgw
y/66/zxxbNrgYSSrhWPmYLNLhNNrfFBW06/EuhTRhWLtqpaBgL43Cjk+SeK9ltGGBx89tEAWXNVw
OF1VnToJwsdgJu0O0uBkmjk55n0AsDrbjo1fvdDC3u9BddqQhvH016QSHkJJgsgCCIdOtMEzWhwb
n9XgPVnBkVjUcIaTT5p5N7qdrn3nQrY2FNzZtONoDGTyh/ikkAC07R0zP5n72qg93Dk879pf1sEA
tneZg3zs+0EPCoUBUK5YEhXn1APK0y9ORb8Ww3nQrZ4vd+Y2MrisnbW0jwEzCARhO9ZwV6UJjCg0
Hsindv+gUg0KZiXgfdcNxR5sTsVArL5EaG3bxQETX+tgioYx5XaQG0klA56L7y9wmi8gp3l9eTz3
fO4K+NTgT6w0+1bV/kImzdPnay1gKPOTTkykHh/BgMPfFn/bgpqOvEoz9kv8CsdjWaB3MHKAF8SB
9Ik3ZG62v6VWbRS+ALgqLkK7D6TRtqOH3K/Z91YkkeLsenA7PuKincUydlUwE3dpYUIv0a7N35sd
894muD+9aPn0d3i5n88JUGnsZDZOrSB8Q7YolleUmMLoY+fvY6sPflU9grKKDzuh8Mao5TNB+/7t
02h1OoX2Y/Glh0ZSxCAc0B8YoqzKJIq9wVvmMiUERhXuhG3vIQb+JTqZPbhcV1rE5lhN9HO9LlUG
/Ehb5D9SxQhrV4LWyKJQrWahtK1GDLnJYKDjieDNsZ35eEKeAA5/Ot5bk0wDP/ELAWfSUaNqwyYP
LneDlnzR8G6NiBzPou3RCsky+qO+Jw02gEooW3yiIm8mdE30MoPgyhZpSL+KYU4U+cZRTlQjUQV5
HQfwcu7HwLdxpfpqX8TiwE2XXQpG57v2Brov7eD/st0jfjIh032aNwGc4rJSmIN+3kiVse32Ptf9
X2pGHY08z0me0XJkK0xCGOHOouaR5i+dZ+WeakA58C4Rh76OgjlfHbbXb4iGS9LlqNDROSwg0vTv
8SFIB7oQtLRs0CLfjWnxz/Pbrb8kty6Y6LTdwnU9xRvqCNJIcqon2qZqBQZmYh6Mf6k8EOVPz5FH
Oed9q+VIqgKCJ5oYsZOVUDlx7suGjbObDbA0FDH9joRtZq0gql/SDJJMcdc1SFHPDaDC3QhXUzOg
yvj3TrF2NlfLGiZ2e+jLIGchsaONX8ZQelZgON6xdJgEzJQ/eIi/jVNbhyIE4ID3rqDWTCBAeOBv
yyIiQZKMJqwOtZcbScoOZlb3YdpEZFqlNreW5aepwD/nLT60nnZMtbtuw7p84L5+t9RSb7/gkoIM
KEejlZJ4nHvb+yI9jvZqUaw2S7Nl1P40/jrz9DQqoZEy8zAE8DbBTQwiEXu2axt6cxA/T6SSikZj
FQr6wjGakh0jXUdN+NrKXAW/UpuML6P06hYdM13V9vNHcE7GZBc5UeHOsJH8df5anxUi9wOqKXKG
VGxPmxVEIEYkYgD6yma+Lw0PN6acvpoq8tywnqoef/P38Fhob2/6ECUlQscHiDVMxvyL32xz661W
BTMcSifyhjq/hvnnWiyjHHFEuBx2ubV5AjOU99YQ5NQNlmx30KzrzS/t5xOZtTG6GupOU6qXI10w
t+BbGpqjMo9JrN6DTv1LvPRRi1AzR7p75n/tZrSRngQeeb4323vN3PwdtyQddKhBV1hlAF/SvztV
aLRLltVwFbHH+/9OhFjWYIX0mJqyFVGtktQoTTTC2Pk/UKEff/A4ydSOvAgqFrVPh3q3klv29G0S
GS2rAMaWvtQXY4R8SstOj3/JufrkprVSKXpSNn6zAp1i1qOYY7SNLBLKGM/3tIDxG8K6CiuxKOnI
a6uuV5fsMrgL6D/YLb745zKGBXdtscOqpYxKHUg9wWrSFg6rx1/DKAkTp5LM/BHzj1Q2H0yhd533
Y/8/D9GDesED2dxl/D4nhKn7QnICl8NZ6UFkn/jhViFHeOBlW1/lxxD9hh9WxgUxexu0RJWSs8fY
mrFuRhLYQyMgXFpPZD+Tbc3xt+o/b8Yzp+pCqWeoM1rOeX1RhrEZEm6zHpr5kG0RQliKJSGmH+HO
S3pyMTORmdWVyYReMzTaJKLp9tY6pMV61yYnErouity8zCxTAcnSc8L4Lxw94SaljcTml9tTzWZ+
2giDwvFCNW/wi0fSFcVwxm6zfrikNgzRJ2rNEY6lIZG0LP4Bis+ddi+ZhUOEzuduS+xRQR2FqlZj
iO4tIZsoDl913n0pmYstBh0tWjRb0RlGAZ8pjkKsFQdJ87kaytcjWDEQ5oi0jySpcFo+g9PsaSOG
AuMO1AuW+qbBsia+AFQY2CzuRRmO2mvH8Q5MmGkcgAFslUjWbws18RU9bsAW6eJdRdK+LWazEzTN
wQijwhWW8TWMjvfdDTeTHWR37n4M+QFzfC/gbTflqHMgBeC4b/eFKxEwpzg2kAgMqMQNeH7IVYit
SHVzYxbAxAEFcotMWWPCDEg8PyljDkj0CxHhMjra1Suz3fxSS4xQsznE/l6CUoF1YulRE/a1+vLt
ePagTWRrhgi+/8dBKOapHCaQGErmhNc9Y915PUlRTUjR2h9/KusDUpQnO2X5vVasLOnjJSKSlJfM
k7aHyVFLa1RS5PZrq+ZzO+U6Bz6XkNNRSXU9J8QazYNu8ETV5k/yOQvfRsEaF7vWDAUIY1i0X/Ok
xPb5nZOTxYU7ofmAN8+lXy5gwjM420UIldYGurLpJeTR2d60jTbGffFipY3gj1AV9qBH4FykrlZq
2pwXvDv0/CXdf/1TIZUA/QUu7klo59IKg5kKm3B/pO29fplUSCdZcR9XTyDbom3x219LM5zbw4Et
kZF2ZmPi1J0MJprRDabqv/9NWXR+HIQ44TANkD33nmy9BvUc/bpyvaAUomNttbseGzIvvz+x2pQr
depLzsq4bcKad9gn+3JVH3lG9XEXIS+EVY8kifVFWEObhDvYYPlwLNVwO5Il7bJRurjXuvzL57V8
w1JdwPM8vP2T/+abOm1dwnJ+7XBaoV8Mch5+YW6zLIvzQ8bcW2i51YQlq1Lw5zbMqFzWUFExv+ew
9SuixvqGH+xd1c+RrgJKuoL6+kMUWJwT6lLrCNl3Qvv5pPhux6r783Fsmx/0cPJ9fwCSoTwfKLk/
/87C26E6IkdYu0Lpg08svArdwp5GpzdTkYw41g7noZCcysx4mE4lMbHwmn2o5EwcQIOzOxgb8XQ2
PD1u+UmXTYw63iZ/BIuB3uNwy14c6jdb6ev3ZeCyGi5bkDaaly+ACh7J10o7XoFszEPxQjTxt2GD
4pXx73nN9ywFUYjHnMMQx1iVNDbMnUkObhFMTzBBPN05/NT4YTZ0gJHVnGA7xnzN5OLjwRwZmr5v
GHALIk8sKRWszXvk1BPcSG628ilZl+nWSVTpdNLnEO8S+jCRT0R7b5iiW/CqwafDfd/ULZ1qpeN0
3QGZYu4pN2TT3AEmGcC8T9I9sJKoOyfz3eaYcaEFXimCBtaO//Mtuh47WaSzwYpwsZQ4yNfvHlIK
W7IVFPfFzqtdb7adHrs8qTbVOLlucXPGAjYEdIt6ITRmt70E7qe/PaJ6qwACM28twqqJYG+Jrd4R
slBXBWLBrmouXzIwwMNngkByDQiUJuk+EhMuad4dZ4mAyuhiUzeL5NmUy7cgIYC2D+dsSwJFs3dR
uoDRFeAnHBcUFDAb6J6mBHdi9veFXd4amTzDnttS682VKY8Ejb1btX5ChZGC/onVFkG2M4MQptQ6
h+5qm7AQm0UGWF6RnWf7ZTggB6bV8/4liQNwxQm8R1Hn13HinROC5LjwnKOLzs137f/2R5Ls05tJ
4RZzTmkroGpNlScYo8gYt1V4sse23B52nIFVShaPjmS4vWkawGgGm512NACwyRYXpYHRSdLzq0BX
ZZNASbmhoOTcsX1nyw9T0c6dXScI0td3C4S6jg/6hRx0Cm65lSdvLgdYyUislJ9m4ELeSsHpiOmZ
nrQ8Fib0O6FwmJ1RlwvRQW7lv1zVRDY4bK1urqvyF1CYPRwstSLSVogeWaP1VigKKBTwqMtumXMf
ZQ266vp4ExR4/7Z5yBWWGPzbglb/HyA6rttX9vnk4yZZkh03op4G5LsO+UJMn+tcTFYasGtCdcuF
AN+MoykwFnxA5sVWhJHHWhinNn5di4wxLXKhrcr/oTp8erhINkUceh6I6evIB4d86X5vsm+4G4O8
746J76wnM6dzoeuwE4o7dO7cmlXJWmBXUlWoUHwq/VgPYMcXJIvcJBoq5/2JfKwIO+RquyPy/Dw4
Cx10a+aATpWSjVgIdwKGJ1Dp+BuweQRGDTFaVzcNx9GRon//v2IuazSjAF0G9+Htgz0pjcgCEAOD
WR5FGY9TcTMGk6uWQAbNCO5iVyMBU/B+PXGKyTt7YH/l4WUIWmzgNyUFZxntHCS0D2YQSIS6RuUQ
dhSb9k+dTrcNi+m30pr1CUB50/SFVC8C1JpXhaYJxqIHBVHyyiWWD9Q9hOxjBmip29OnvTOLRl9N
pb8WAVWHs6CUzxh0xme3mwnS5ZF8mSsL3+aTjKuAmJFiUCU5CZtvwo4zgpGF2m664PBth3U5uXPc
RyTXmOTDrbFP4keliygbyteVnL6YYyWRQTGHn+ew56nQDDaAhT1muXCWP//EpVkI17OsORNkeDzq
X7Z5dWq5GZdpRcOcCGwkCmMbKY56CU6mBsCltJGwQGOEzdu4XIsdj+16BVxBUW8n+ZSpLV8vkRm8
O/kVJe73FtzhUqmr4cdOODvcKFBOicIB5cJ+L8jyNNJT0zNcz2QIKKdOQY75qVJfUnA+8JVxhIt8
vhG8HT09t83SdHdrtfl81s4Z3ZRMf3z/aPtI3wMRpOfb0MN89MLVD1zRi+6MwEXdRDP+9d3sAIqy
ljRWTe7tgb6o5ghve2FtjAJRYuSpu/eSUC46m0ZjAX+xa7GRm0teg4oBqW7wx6d3DkHEJ5E4htQY
3H5rOp9XUbAOq3F8QkP1T5rtWH9qRbQYEQLJ81alNkQrkAFTs8AOFsUMjFJ2iOJOsQFaYhQgfzxG
YkdQ3JifRzEAIfLeEwZADicOG0HjA/zZtLA28xB/VcHW0uVPk2Zibe+IoYyoTrWcsdCW1l0PlJL4
X/sbbeG8ReyRgNBhyGYzBMYgZ/Q1HYKnkMJvpl5cGb7sN4Gm2LzuYXqsMHa7fPsnVww1JEf+HIgF
svZur+VMNNq3XFDnBUh1ZV3ahOTzsEF6lSxxipStLCYMMPcE7U3pLgKLwc9nh2tFz5d4/xt4O87f
MPm5nIXPMRjPDRSQSuQnz7aeRh0yK5Uf6LxX+Z3yiP9VohgIvbSaAqR+ZDHRrsGpVRi1a1DDwG4g
Wn3sRqVUyeV+I5FpO81/f/voW4Z+iSIINx+UoM+33e2e79wzviwDdeqdipYYDUnnY7W1MAsiwOuO
gG/eOgdVYvNlwY5OuDF0umj1qqs5Rs2yA45aCQgxxV1gE44IpAeME9QGZ/44Jn83HJkrpTmwhlMy
BoNeJ03QY07ziHTytHR6Fc5z46rxozWMTEUW1u18Zigudipyc0IStD9Wd0ZEsCLvTi8lDWtsz3dB
v1NlfHTMQjVsZXmBXxiN8AKWPaA/w+NO0Rtot0IVdECPBaqc2OaMLE4U32D9QIa0iCC6G7qOODMw
gLLMwHYt15jOfKDyNPkf1bgf1Pl1zB95AWrhCTXzflaI1fNOEXg0qd2mMacGxoNMf2Dof1WJx25J
v01mpG4wnkCOYRjS1GdM34uFawncMTCNtfR2leAPiyRohNukCbS0tLmuFWzk2XgP21YX5LRJ30yz
0r2Hmook/72g8nDWO5dGu4/0qRhqPF2ypAdKkL/9f7JIAj+OX4XF9aNsmQTKB9DojEHUv024Km1k
2LQrSZ2mVQV5Y4PlXMch9WGSGX8TIxrB47m0QzaH6Nd4+FcQwJ1rRO/A/HDBPP7HF7J5A/tjdUnb
+V0jLjA6VbZRNfrjCTfIG9JhQNNlTz8X1E3JPO5ZgpaZIuc2N6tDdIBx1eh1XO98djUfUo2FagTd
nirp4TIUw516MyXAAnvt7SUGpUb9PYUBv1W7ziPL4MAqXCWrVDTWMkj2Kls2jbFB3w7FGoFGIM3H
6B/E3JDFNY4SSUL5fq03fU1q+vDJ/5h6MFuUWEJ7xny2IZ1+2Yulgur9FQeynNW0EBdwHNTMsKTO
eMbFt0xfZJWWx+NIndNhguU4qpCPpQzSqQaAU6nhvrlU5I6xk4smeDv6clytECEc7rOmSa/7NFFS
/s27NVXXA4451hM0twlyuaTwf2C70oW6GTKvgFgMfy9I7l+/QwxEuYP8zKm9ZU4GcpUpyJFUwPAX
3YvHJC3V5MHP3uGULbe26f8EMZe4C0ZZF7hJ6QKz56CTGTOHW7M7ym4rIw3/3tZNqFRZjwNm0MrZ
UZeNx/vv7h6jjsYUPpftBXnFOGmuLq5C2yKfOJb1WZ2UU5ZH9fxhN389ZmoewjIGVnWJrib/L0//
DiviMy9uaUMPiBaN/3wq5GIu/gFJZDBsUHzQsdVspLu5iqmMoYx4FZHGCvsWeqXc/m15RcK3jjoV
H6bd+7MR9wbMUM6jcpYNjWjHxS9daU846lL0Ia0BtBX+9c2c18NlPzwT5/L3SoDNsU86jz5VngQm
4EwmPzTH2PVE9SUx32dTR+4YPv3X12g4LLBH1+YevhjWSWo7m3Fzwu6dH7cRVXejD09hBevH1bZJ
uAk91Oh/iR34eS2wX0zU2lakvuM9d+MknfSZLP0UXyEWpZ8yJO70+jTwVZL10F6jtYQQtVolXx6Q
MYX4e40Iu+WYqGi6ftx6Z0c/bwkOC2SrtUjefLccQgyKNrOCX/CsxadD8hMLJWL4M7BENqOhCbmy
FFhq4etm1SjmMQbvbhOOhDS2oLvEKbVIRNWEe2VHnC2BXXBV6N2emBcxC00AIF/olI0sILK4EzMQ
v3SHKjfXWvXHktj5L/LoHeEo0oPg9bjesoLwsFXeI6hxlPwC76seLDa/+0yZ8QOJhIjffJHnT4XV
4iA3H51zq/XDkfcw/eQASEi5LS4wxDd7cM0Js6u4tnZj/5Bktjt0Ba8IpQWEav92dKLiiYvfuot8
dRTMtx0byT/4Cc1y3Gmzb8/sTNAQj+76rHDdfy6Tj8vt0zLAh/W39g8nYCYdB0IBMhmT3jMLFQ0g
RUy60k82G9UHo97sOpWY/j1d21kUB0uRCVhu5Z6efZ2eTlAMJz8fhvfD4G6JU361xbL/J48nQ9Lx
IpSCg0AT11j7VrEYK9131uvTSITFYM9fptVQmn2ijMatOTM3iWsOQz51hLyJbGNrbLUp7WqjWtcx
wyfeOv74w2tIQiNZCf/KAUexMvx5S3dpC4L9ImEj15cEaT70ft2nWlO6Iz/h802QK3PGc0stpA/4
cJWMK/C1h2H9tM4ZC7BjGhUes0ccGYtf8X6RsxTWKkPd57jZWbAKmr424FixMqOUi5Iysssr9rSZ
amI6oqzNp9jW323BCZiJH+we35/I2AMkHrjh+IgwCdhvveBUJndwWJTd9NV99GDa229eNLkM4DdM
fwg1DFUoSP0b0WTn5nFuHYF+CH3sWM6U26CcFh9KNcvKz8YdQpfk8Dk8OI0WDp8Q26xdm3Vkf+qM
yQl9KMCkQNCFv7/XGLHaAwXupg0xck7kwphCzuzAJFal4zr7Hgbi/YcQ7zs+4HCFsPIBd46PS2Cq
kRvUPz6kGA8lHK7UHp7zFM8ZIlFx8mQbzEK+0EPvV64uUowiMssC2G6n8uMcDWRy0JNUmsWHYMV2
vXugt49I472GDqIpsbW9JMQSQPt4KXg5UqHxKafA5vQezqdvFVYFlz3D1pw1CmGiz5lJSLzampaI
1OCqP5C5geAIIkgOam3reP4Z1N6lhsj2VLo8bwDAns9oP+NlaL35FLYvfCoaP0t9VlekRxbgFsld
HMy4lMCqtE0FQtCwhTn7RjARzQygZJ7RVaagZQ7oeHKvkplr86KaIuPnjZwNmfXtZx7rnlJ8YrzU
s32qyKOBVWtWh64KmUEJk+oIa5pMN0Nv5wVY6+h16CL4twZao53yvzEQKLpDfzKw3XQV/BRCKULX
Su0eNCCsWVSSEJCXwWacrrqJPz9/XxGRps4cEyHPOCHTjBn+XEqBsXI7xSk2QUgUQS5uebBVHcBJ
bDmebmMo0EjkYsT6tlZh89YJndiMY8qaLG0xbX2zxenAC7TxXnpRJh7FyFe2brJtKIwkaMreexXp
img/J7Cxq+a4zI/UBI1Vl9ofXnSPoyg6/mpq37qESFHNG8JaHug1t89QisCGZrvqaaBApMt37Qj3
EXwsLxOsjMItcR/wRKawqA1OAOP8OlpQyz1FmTn8ZjyPcU8dHIkmUoa2kb8aqV4/WwPpcXLjM3L2
Olx5HhkIyWZVcLXhXYfhBKc0XlGwUd8OrIQpgVP/wCKdTAxC6rhetbmslaPSknabz6U2itHNUOXy
PTSZfXGDCnkPueobNlHHq5VVUE1O4imlLFXf/K2x1FsgvuCuXsiY9lz3wwtshG3LnVHhSW/7AbV5
vZ0U6xMC64vLrNtJt38JG5hokNE0zbOLPR1ggK3gGUqiRXVe0gSTIox3Qq1Vp1Jr930j+PlUZejF
2KpyjF3tA0YJwZ+/34I92VnU68Wc4J7brvhLNyGuXw75H3xJr7N7ij6/xyjZUK1JvV/wtgm1EBnp
Ybx4/I4KzaVW9Q1EPbs/qMiY+VY9pxnvqGT1IrwFg6ogBKQJuZSH/EzGJBQT2BHYAUX0KnLZXTC7
XdUlGL5smSMMbottqzY4dM9V5NA8ZStH9ta7Jpt2R6IJ5cUP8KCeWJLWwJO/V50PT0eso3Xsdtlt
vqQk5JiJKV6e+/9VJOBFhP068S0Xfr92YNK1akTEumr0Xp+jVklOw9u61h/zpkQkRXMhHa5l4T+K
ekEZ0FGpo6+khQc8jo/9JdA1zJgy65ap8ISv7sMzydEoTEe6qlGqr0QKiIPH/QlRziO8MKy/0IeK
gd3oE/W96M6AMRE/JGNHKE2H+sH/g+gf1dTWWLZmDuCsV4nIr0s6tpg+iOBmlAbnXC2mWFouTYNU
GBzQiKsgm50vmvJzo3BU9bnz7xH2v+rIL1vmIS3Z/1/9sHV5JdWxog5WKFZMW57p7xpascNGziau
wST4Duo8lm/DZTExHU7Js7b6eFZQf5YNCX0NVeIGVHbxIQu5Tru/9xsNtOo6HWbmRJsAWX1cYCQa
MHDqoHBwfBtGhzo4i0kTpeQqjqIGnnS/16GFrbuCBChT5PiFnxJ39cVAajbKKjJhCkHLdut0mh4+
2Ahz60PDrcD+E7d5Sy0rkB96YLFH2Uqzmhc3CnJ4gdA1CL30VTZSKYbKYIcn3WRWn/hkuMdmVKvg
wWmoiuoefBxOTvk8yd7FpKxJPnFfllWWHL6ZHXm/wKAAHvaqHTIDgAIUsEwodvUhKyY1q3wwGj4c
1y7Lp31rv7UxX4Xprpcx3DSSf5O8GQIM1MCYnjHLNb/whMqT4RaFdOXsWJzV8t96pHAy+0/NMu8L
XNMvCLb6JtOdhjlZbJ2TknTv68BaHTXrcarjYvOW9JIf2ylNxrgyF0WBMu9AiA7mWo/Y3bM9R/R2
uqLd+2zNcJvtzjQVo2L+n9d7GN62FalxbLgl7KmAZs4WhW6IVRs9DDYVmfIrH3DotuEWt/nBeqt1
ND+A2uNVW0f0Iy9ME2HwSALM/mAShZYiyv+VSvB6WzWsFUND7BMC/ZjQ6EBMfk6KKZmkdyAbY5ME
eH9/W1uftRsMU2qHTMzAOaEQw2MHLruUb+TNT89jm3cSz4nXVZ+LS+Z5mShey505jP9139Wwi4s/
n9p7tkutAVPrTs+pfmQlwuRNAIRXXkQSCjHMh8BkIcVr/Wy1fbV7drqwJa2kGDeK3g3kLIFaAMd7
t/5tsg1QxA3vu+r3xjwRv7Etlbf55OSVuS80trmB6nugxLXSurypS6mXkgZjvdykHF89q/ZIuzrr
53zSdB8ttRej0QcbyfQhjx4eB2Sy5A2quMy9p6oFhz9pClVviFoUiRn37AG9+rjfd6P535TWIDam
PCdsmbZoydKz2qPAwyxPEbmrgkgS0vw+oXV588kWPF3v3zZrJtTZZSjWark7dSGGE1QOqsey+2gm
W8dp45b47j62mtICv22h+A37iu813POkp7hDUlzuYMx4jSNvbHcODwUXTm31J12qlNUcdsvnlRl+
CodseJV/Dv4PdZUgYH0+W5P2H/DiTNcUQPU5SPP7RUABcbxrEo0wZfRL3J2exp5ckRjgoqWlQZPc
R3e7KYnzoBr5aPLZGJWIZ81g8CQaACLy8wxWkbOLQhqus5RdbE9B6em5xv3+HSuA0bRBSpFo57yk
9kITjVrGl/36cZEU86UK4YWnIC2sWjY95jHN94PBWr5+3ShJi+TZMguD36oTLikPyTnlMTsGXBOi
NjYH14EjBKwkdmvPtB8yIDwtd3jhl68r25FDS9h0X3BU3p6xRMUfzzL45QlsSkyiTaAdypKOdCQQ
h7xvSho9Wx4awV/TdN2hEp6RBhP8D6KCr5Pi0Z+h92NceTXNUk1RB0snBlOHSNZdy3mDbY5QlE7Q
AKAnYaEnxdpVRyPkheISjcbTjIKMqZN3RjELFCv60FjiH2KomQQBQL2/Oa4HFdu+Ao8baXEa/dAl
1aeZ0PKys/wXivYjcPtdLpoj5r/1n6puxtfJCd3QW2mRHVq5TOVNWyXUkbfBx4ZZhXpCXfc9Am0L
/Zhw+Ihxpdc71fL4ihFbEb7IrEnnSUNTT+yRLz08F52ZtVVJUPjPy5lnp9yp1pCi9z8kZ/8vnGXn
lgghxI3TaCz60qjPjcVdxehVFx/2bBzw/GBTPW5MImLANQVlTEF2eYTuhnZbYBV1Mj4qT+9w7l0g
qJNOZ/qwcn5Jf1B8snc0qSJsDn+v044hD9qwefbN0sSckeFptdIblxXc+11jCiDyGpGm42nO7uFz
meBLPW7Nt6HhFJpVon8+9vKYS0Rpd2Q9/M+dOwP7TLhgi5b6DzqGnx5eMseCkbPw3T2aL9ajgplw
A1WTmeKzn4Hk+SFTpqLosClmizht255u5Sj6ElugMprI9FWbTP3dvuTjd7PZg73aMbbFYT3b+jMX
rGwHc627YdcngCTCWEyxui3xeqwNzE3XaM7yrmdNPUpt2Lm8JzoAjjQfSHUtM2NmtJ19EubQwepk
doe9q87pF9hicj1seHQV6vWQ4qFD2tBpxfLYO+0hOieChAmYBRaxXpdc1o6ffeUyoTcc3l9ekM3f
Hu+62qT9+JL5BYM8ShvwPCTlRWVkbX0Bq/k1bC4YIU2U1QY+PVC4lzJuto7QScFdHD1fo+P7q84i
HkNKl1q/fKo18qjOlZRKgEiWmEH9TnokrHdRkxCwLLPlFwhqD6EDYp8kTigJa/CaqZ2nsUaGceC7
ZCvVqkcNuwgLEcqRKdcuyCgaUK80hyDVt+EhhRc1q/5YLaMpA5fKldnUtuVhnx2nakPikidSJ3jJ
O1XxYrFvFQ4XI6IEWHeFq+rG+4WC7g+n9ApFCiH1MheIhSbua/xop6GA5lDlpJe3yVCPZ4dITL1X
kTow8/DIqmf0s1RTkxsSMrmfG6dp+B40+KDi1dgqsgSYt57phZ0FlxYBgRF/AE7NdQbOIA32fl9v
DVGa/4ALwYhW4geBuydgrvjIrBiv0HL375srYr0OJzHfFk7Ux6D6sm3J/h3TLQOkOGKh63raUz1V
xGA0uSk2e0Ygr7Tznx07UlrHy83boU6tFSn7DhkSpCqqnhe0irTOjy2BJnsKNxC9jMdMdU1XbLfj
OqWp3kSSCDIymIQ8XKLnXEKwptEpZIune7Cf9hNZ1hfTlYShyBsLT/17vzDdO8un2Auk2GU02uR3
MKRbKXjgfdfi+dNaueseCXfyErCZyPnruOtIhXouYoXdIaSO1v5NRBp1V2SIAxpx2WDnsfD5xbmp
zsP/olscOrHkROdTFlJf5IJVxO76Ggzv16dlKDDhnYpiy26y9sG5AFvpw9oTi1Pd9OfXjssrCgPg
xqTThwmSDnrq9n+IcWdvV9uTb8De1Lqm0m5qqoqWamysx6oAYJKzZbpsDzLJpl0Nj0joaK1gkkCJ
Te3Fr0SLcLSrqSP4/EIU0NEr/i+3VfpjW0VvJG3jFrMwUxhIPPZfQXtr/Yh6DdMhTwFPn58QbZ0h
8rXHkmKUIH/pHquLEGVOtSz3EZZbRRFCZGyAURHvbG9uH8w+JscAI4liKnxEK0qfkDhA6UnnV8Hz
KJSMLWI4suRTQLd1g8CA3EnerqDl+w/HUR7lh4BTgywwEPBH3oD9KmklQfJ/P3lWk1J7W3+PpQHU
LJ+JheFn3++Y174DL/nTyQSoaG+uHWZ0yS1ZsLw8JGAsI4+LSpetaRkRqfphwVKJwrn6gIdelpbA
8SxETN7rLAm/z9JtgHFnz6aKNS7QOCkbuytlTilnKniSqAdpMpCxKdefREcqJOU0kk+5hkEUoOtv
IWgp3L9bL49vA4hXIRNM6KvZpLcM59P7FUnyl03ua5xabWdQZARu+2+dJtG4qYvvh9i53BL35EF+
+2wx9r+ZF9oqX10Rpd1XNjJVGdzMaoSDZ5UegXV6zP06ZvdfiIzp8kK22RtXkNXdmToyw6YrOb7B
TvS0YQ8Zsu/SHjMGFV73H23sNeHExr7K7BSb9/zOxlhYVdyJOjVhLWIck2qfAm5Lj9FfeHl1mQHx
u4l+veCS2vdQaKwjqE8f9Lo3esgjq38y6pX10RyVC/rIdP+Hi3pE8j1z26XI2MEn3EOKRR8EeEd3
+73B3/ah7nhPwEUqQDHSImLB10Kh6OP4gmHtR7HrNjY+NZYUvtIcKUXrByNtrEwt9gIy5tdDNsBZ
FNDhApZxLCJxHhQr4OA7k66+//J6NtMex7ee8D/e+nwC7y1TdQXSRSX2i1B5ZH4ydLqXQV+JZg2i
aLxFYnBj+ySUBml8qxf+sIP4pmu+GFoQCdKIPQGkYzBd1YHsLKE4gZscmusG/jRlF24m+TSz603W
HAHZ7pRmf4yufzpXY3lPksKlpyq4oN9qLA8uTDXpdP7SRIFSrlsHiie9/sdIJsbv9VXo0pKosfbe
CpxrIHI5l3Y0H4xET1NB4mIdltFGkRFM57mfaJPCQ4QBERIfhyoz/CRNoPOz0OlqTAh3ZCxyf1yU
Dt0gAyYiTNP0deuRqacStFHR1zmvSByV7QnB/3VPNG+lTqav5fZrlpk1361HmzbOxXEBqoNfzWkI
R16qgzLzLGz5pUCK/cKqXLHCabjliouUjQDOKxzvFtHLYDfv8CcWbZDtBJbstpnYM66iGll2N95U
PVmzJphBQkaoc6zw2gSvqrJUNU8suZPNwMu1uRctSx/YlxbXMorXLKpiFFoOdEdGQos9Gd8tD/js
BG58yFUmsphigpjq+/D8Fcizfp1X3f9sHRIT8A029hDzhbASyPgF75XbtQEjLkRqW1rwkcfQzzBv
KdSuwfYzwgFkh+oQDRK5bdvWXSlv1xwhIvWnv/rmy4VGKjMuSajJsO8xZZdUajwD8fkYnzhKEP+F
A1G3blC8boIrKHZiVOcTgyZyuaho5XQRhrfB9+g1rA+d+5MPacoRPyMahXxrGvOOv7sVamvBP6uN
k4lxno0Zx8CI08wANQqApY4/uOrG5MG6NGV1utyD/n8FXmTO2q2+VcQcwpBo0wNgC7LZk7E87hRU
dHm2cQtWSGQwDs2e8phtATqFlOgx8aqBybxMw0WQGL3nBTTxZiHulbMmIFbF+wU16sZdLO59iApp
GUck1gSeOvCrRQY+/w3SOdR0271MgiETL6fPWrOtKCgdsHRmYdX9yX1RLPrz8OPX2rnlJQ6rGqqJ
UArJ4xRkj6TuHbVMakgYqiHKVbZ8z3vBosyfub56WtZwH/E5tc5k39x3M6C44CXKLKR1vNF7Lbik
9t+SuvvvG0OHUMBcM0N9D7trobAGUDWkaWHN9zaqI14Lqc6qHlk4vqLY1rb9zQY94kh06pWX1Cl7
hT3DqZLlggRAuTU/0m6pmkyKVzo22sunryMeL2yNtfTy1EBP/IYvmqFbEXgSPy32hohTe2aF+ZpJ
D2j4tj1FuGOa4gVtuEl4gPPR2IsD+BUrwf/AxHQDWp4fiiftb0vVUblFEeOCjvYhOQBTlyyl2w1q
B1D9O2Ha1B2NOg576BoxSGS4VJ71vrqc1zFxdBbaou1+BfQNfdj1jzsTETRrLCsEuwo7lqJqY0SF
LoqRsTEuuSMBowFDpHH9HwgUdtjlvNln/SBBQRE2ZHVXL77zGyZ1vPoJ6JUXhOnTzHwYVCfL+MJS
mcI9Wguf6310oaJ8qwyjmU4uc5gP2ehMN/C50CCNOYcnvw67uMTDMjSScSyxSRpLzB3LyJfaoT7Q
ECA1RQrjAXthSMGbLkJhIJ2SPGZ7wDriXANWFsfyKcX5uueYgxoLu9k2Zgzi9NiJI9VJ2fAjoNVr
GeBHuUBaf3jj/sjM08Iih7F360mv8Kc1Demj9NGYvSC4g41FfPP18LheZd8qf+Cbqcm4t3YNntw2
H4bvpYW4n+Qn/XbcEs1/aQcqJsIPe9YztebhX2dmH8DTh07w5enKN/UL8+dXQ7EyThSAtg0jklI1
W06mw5RQUWBjvVall4LJTWUtHbZ2ThPwwK2kvzEi+B5wAGGAEtxPpGY+CstRDzFmHe7h5ZQ/E4EV
bQhkxxOi5tv+2B/PplAuoVswTu1+pBU+OzbFr0wIzoiQabIabG5zW0BmRiLQ9hPWI1C6tntqgn2h
CTRkHkxoncKVgBq+gzfasyjV4Y61L2w5oHPKTi1yJ+XYBfPA6U82DuMqS84ZFJnSsWATDIKX0PI6
1M9htaCCeSuWnaiIFRDNkxxzXX3dQYWWkJY82tIjjmT1nIR1HOyX4WK64eZ8cx4Q9o4Pmauu2E08
RisPuhRJtNJAY8R3fxN/s1G40akmlnrHEMLdZiZ8kJ0FcN8VMziBN8oxyEcSQKaHpFWnc7F4Ll49
9Q9Oj+3Tupcgul+go7syGErhR6/LKPCiLs1uDHHlAe8nl7gnhH93ael5YNaJtdKrG1MRpTIpzusr
NppdFaAjnM/CT4YCQwLQzLs/AJtlGSrH3w/l2Kz8d27YZ0TgxYmKoZiD2FdWLox/yj8BwOAjKumI
33RGVfYQ6fnYmEx80q9VlfwRyb3iSUV2fqzMY12g8y0QQLPmodNhvDB3lngo7WRs0vp8IME99qbR
lDPWQya/AAMkLaTh76rxSMHxiGT+hwwHi2De28kf45D1BZWw+W3zugdsFpTWIbotlv1rVd2lFICr
tZjSRQg3RSR8cu93C4lPJXeR8oysLLm700WChIsoOkzH6Lff4PjA7j2jrPNrMWHhIuYRt9VtX+Vn
wUzTUwoS7tsNr6Sr15kiegEmC69ujWD4E0ts9hjwchxRt0K/R6KV2wE0g2R/jLFw/q/XW5pPihpL
RXukXdqG1N56ZpU0SBtDpL1HAM6f/1P1kup/gkIJ6+TVjc2zQpn/vQbtF2FPvF46HECYCuUKNQ/x
0BNsp2y0kC9B6aulkAjPoGZUeNBhr/aM+pFSMHyqzkFZKHnTFVnyACzcYjBMt50ziTom/qK0Rooa
WamckewArRXnCslwqATy8ISepa3g8QonCTI785vh/7TfcMX6/BTFEL8bVakyUCPTSan3SF1KBwpD
6LxJc/y9fJ1jIqkcSsR/TWJ3qxA+b7mJ0lk0Ff2dStvqRO1m+TtB/9G1Mm+uhi1I3XQJnvg+MnCL
x2JoiVrERVWzH+OsD+FHxkVjUS1eTf4WyACtzM2xS4bMj/xXyd7IyuOdlK7nAlSBYPJm919RIMqi
PS6KoXLYBSXlH5nAmy9rpbARVXCKqa2o/VB2ecC6A8tF25FdXwaDIzyUWHncdkwzoYV0E7DTQUUT
HUD2HJ0jc7h7PG983suXa94Bi3+q8OwgYb2CSx7DWgnTNSVUVdj5JOm2iNUGqja08IAJcvpU/e73
NmGMMy9pIBA/8sCr2ea2mrtrdZiF5ojRB1ypXvG/dDwTdqpE9wlCaCy4S78xq6I/2+J/ttKId4Zy
mqWu7ZrTvgQ4Zud514b2UewOs0sOo0DKkdi53PUhgNRzTcujnPozXIWGNkJypyHGicWeBAsfJGkG
8QoQ4bCqHjOJlTNbUL1DoQphAnxHw+Q8Lt3Kj/mM86NTcM0D8z+P3xlg/Hux6nA0Q9Ifu53MSivE
u+Er//5xqQ19GyiSdsf7G5Nq5A3JnPL+0NxQ/wuGKFhg7B5npPb9kEWuHYM6T7u1YXh9m88cc9B8
4K3nxd0KscaNwy9N4WYNL/5x1msuOPeKcQQwQLqsLZY33E7hqI33veN3zVqR294yNhhsbSjLoyZ/
HuhnVTrtmGZsUWVbcFs+lqy6jZEHBg6A1Di9ahYO0aCDrgem0y93rWivHZMnghdfjBZzabZLr8rE
zNulDcGbAB8XbUmkNOcxFa33TlZAbLG3tJnDg3zbCfiBRYJkoYqalixsjGJNoGslQHZUbKLMHMh3
tFUPvn3N3DjwXLzeEv5gdPYmRHD3gjdusgApyzsGtKhhQzixIGBFVPPzo2IPVJQ8oznkIkYpZFT1
p6As5z4SbnjOW5XGLYtnbcvdNor/CahyjD5cEVwZyL5eQSj5sizFQHof8IgPlgsc9vduCcWkb1Z0
W5B2KQVjQWTGx2gQKu9Xk62frMBSICSrO68UjEPdkAKhm0Ek+3J7tHxmEvE6LHiV+ZN7cfjcjHog
P5P1zw9KuRCyjiCL5SOIwnk/oSKrz+N4kw+lAJY4B9fbdYiBU2u9FFL95MNQTjQcSF0QT/DT+hu0
4tXpQSc7wjraiWzYEa8FnaHLRaGYlyRmmyEi6wOUK4Juub982MJ32f2DOjQqVBpxhrz0+D9haHvG
y4a5jFeINylAYTakZ6PyTqR1O/fjZT3czYoIBT8UcqoR/ZrHO7xY+nP9Wp7ANnYjuGuwfFRanBmi
p0nxFgbiAdSclJPgt09rdnSQ/OM6r8nnT9siEMe1+XC6zMYcZAOA1V0ndecuSvoGIhypCDM0Z7nJ
SPAcfTS1ztSBQ9IQ1Y5Wb548JkfawJmPxe09z1z1A6KQnepbxQI7IY+yurw4k0ncTntiQptY0yu2
9c69ueVOl1RkqTlGnEitjGn52G4pWprgwJ/TMF/MS2vtU9YYeirT6mYVHfvmg1M2I9Dh2SwlXBLs
3FFo5BgBpul1j0EdNOx++p7dO4y2G9pBx4XNa6UFJJx+GiZZ4GVLqMuXWqUJpzeRMQSSqW7mBASa
9VF+ow9XS7YrLbXe3HS0shYKWbBs/CfxmnKQB6OK38r1153zoxnkEjmQOchL5fC8Rj1UN21Ouigx
Bta79sPwdyPy1vHOdp6aSIpAWna/TkH0evNMFqjCad5mXqYYQj0puGqmkTl0ZAzk1yCnz8/Rp/Di
UBStqiaF0yJtxdsN7hROHxzkMoWFAvlODUPIhGgQzDEM25lo11dQUbnOzN2Cp9FiRVxxZHVZlaGD
DGptK/J1HPxF8bG8WBl8y0lvVcTs+xfudreqy8u7crsjMtzfxyJT7l++uoEP2WtYcGDj02IFx95+
rGPsQd5He+8WuSBbHgLDdIEmVCTGAhvZWMNVEk9axGQdQ7TPzFY0zTOjOqt4pzJ9PlfskCO6rfF/
+kvIMG2SDbdLGjOZ4v1ltw4dlDCw5kLBW9L0G7HRMvhp4yJD44kP8NncHYDle88MLy0eztfouvlv
x2hzVnxQtjKRB4BL086SzbqQXScE/qUvyDCzPhaDAo3Dxru+KyDHqP/pivrff3+uIs8y/ryDRxfi
78jpr7syzGWqgdtgSOthdGV7C7GmAWf4H0ujSW1di6UkgE6GnE7gFllzakh4XQsoxMjsPjUtXcSv
55GLZ2cNbFxxUtaDWsSjeDoO+OqHQM5LIniGq3h7tO7OsXcEkv8/mPpIqMHCo4wmQFcJibvH0QhW
2zNfd3W7CEioPp+tY5M94t6lFYVP8uaAYqEBc2JpimvbGdY//3K58Yi1JBUSv64Mp0aPQfHp9145
71EJYcDMvUELZTL5z7kWisEL6apvg16jx2onLbsg9xV2hMCqW165OJZiu1GvzSEwX+9fdK6jtXvv
5jZnL9lnfQtE4XOH1wg/KYStTfq7ownoZGzWArAiU7BF1ZLgbFHyt95Afpb46zxQhCXt90/PdQs3
WKhFJnX1LcUSJhRItIpGyGGwAASvpNOKd9+b2hFD4zE5ub2bGWBv5sDDpO84U4xm2WA/s4JuUC4Q
tTPBOg/IRnm/3ug//qHmSazUlQ/elWzT+gAHFqcRD17RSxOxNhBr2fP9rhfEqz59vul3k7rXSqdn
VfGbDqQQylmoa+XiAbcuaZcsKF5Jug37CmIQyS2ICwbs/hm9VyZXALsI9E28lelQig5bgZIgxtSm
IBG1OphkMsAEseELYNi+A6WElUX8MefblMDUo+RlikCqVRl1LF0gU5iHPCSheplVoLDs9RR44OgC
bW3A4yen2IIFWSDYFqakHFrIWxS1J0Kc8YOCWGspvD6vRkoduTeqrDXGCGl1tjPn9zp9xs8bST21
CAXq8348m6vip5lP+oaZneCCNKbLs4qy1VeAU0bAptKUf7IHdye9ZezP5z3lMAyrKB2XEKJeJL5n
3rdkhVjhVvLCnT2LL/30d0KWE15k7zzX9HcrsJ9d08vkLOb5mTtKO+G9xCmX3gjTaIAEv7opjy3l
QRjp9pzpD8gnmM7PNCA3jDtw2IbddbT252u2Xn3dgBXDnJe1u8Y6sPjoedS1+Ytih4muQtQ9WqF+
fNetp2GyGG9G4kqMs5UHmTNF5qjcQLb3EvFrqawi/JUCBpf4o+zvN9G2OIi6DMImEhkNQ9BwweRb
/5VsZE6Vxxn3GxmNxr6avYq5DFJDvS5As8Vc6oTl062Fr53//N5qagGPH3x0AZ/uow8wu4pZo4pj
8oHyO8Sw/8qb5Oa7ttU9EO7i+ea8MIKhx5358r0k9ZVQW/ZNvGBev19+iJPaGT42tdM9bhFN5IqD
ImCETjEFKMDCWynh2jb8uJp8oyQ1nzzjmGUci5c1kyXNE66YResjUu7WW9KDR1sb3HMUOvEw86OW
xAjRMjAITMTBmuCckkW4HW8DUxPmruzvw7j/yz10CyW3mKGHXG6tMNVkIt39AkJwiLPmDK9lWbD0
M+MwIhpNAc0GU4ipClMIyHf4wpOSszsunifbguvEi+v0EyRhfDAO8kBWUsbCmycNc7z0kEivN1vE
64eE8Wf7CB4jjKC2bV7u1FATHpJeHLpurqL+9D1Cv5Q02UtwCl6BK0KzIAGWjuNpV83jgEQ72pjT
TDDEyuXjdK92f8uwbCfx/q9vmANSBx4NjVNtVxYQHSJb2UenTDdIkR2XLKcycYQfpiSbWzEfKWdn
Olkz8SwO+cD5bgANjo9k1Cq8ZvubUDS6sc1cv9egqK/ktiN8S4dOtEqlKPddjzssigWOPxF4Qg46
I4bj6rXqRoPfV6B71s/YV5qxgxrR9DWjJJNoU1+TpuHv9nFq7czp74TU4dALEWMabEqzunTg2GC7
fkOP10OiSNqbyt1A6vdUp9zorrekIhe559xJBfVKVEZhOC3MJXrxCrpjgy7klkH27rP4+n55yciV
3ufz8f5JqPcBiL2Q/eL7FGy2r1EiwcIpeNphYOzk3Bfza+xpBRDUnuYBOn4868BRNxg6rB+RZUxI
/PTkSrFjClevX1yRsTJvOpG4CqWYBU2MSLcxWv7U9Wp7gPHh/nIYWmwazK2ElzkATKbJ2sZzwIuJ
LqY4hqJ4+5xKIzKv4db+8MKq3bbu0jskwZHv2GHciaRP6fFwz02/Lu00wSkZzi16mb10vjYvRWcV
2ChL8P5wYgxVYcp+hVmyMgdhcf9W0HiiDOj39q03bCKMJd02ojzM8UWPMhJLid50mhmEB/DWuXiF
0qw72VlhoK2mHCGOvO/WsQB9F5+wZ2D+vBlSdAjIhdpuhcVThXD2KoN+ueACePhueTutTDvd3KCR
NE/qjVtAv9EXshPtcN2yUrAAqEwNaZWqPYKIGfDmO/1RtNT4MQg1HIUw+eAB6AQp+esuodCEYV3t
YB6lpB0qiiYuQM/+NJ5kqW8mR87WVYSpCywwBpPyHSfOOotDLUwpa0x6BpUtnEyj1MgbsYXGuAHR
Z01+B0daPEeLPYt8IJ4v/h8HNq0BYMXyGJE5hP7knObkOxXg5SXU16dsuJq+y0HsVazdubOWblNS
y1j/WESrg3qjbTk36Qzstv9NihNeU5VHXHB7acHP30AkbtUBzPL2i4bwYIL6DBoQTu1mJcEqs/hH
bgbk5nIb0PPtfPso0dFQscdMkO6JsTghIgrtYDQqvolcLyNSR0rfOHiueOr4dALslDN3wyWnlglv
M/GJELyXegusOgcz7xj61mCBFzw6NgCECNu7ETJE7XjlcHYORmmVEU7FEfo2B1qyrhv0GZktBSyK
Ar7v+JLX4UsioH+oG4HxEjsOz8nQt+kDmEv0Cfvr9ka3cpItNIjoa9708PIcMXZCKRDgvYLnD/+W
T2yhv8bt4HyiFz2r6esml2N9e4lPWCjnVh1aLWac6IvsO+Hnm6phdFhnvax8f03BM6BJMwBZhNzY
6ZJam00EY2JAnkD3SJG6QHO5pvNgtbrdxJoSh6Il9Ee/Z98J2mdmWGsDsE35kGMxJDkBQwB+nmAf
MrHpTlUjztg9RKiLGybdNugQXGIGdInv7VRk0zmDyhT1x+Ccv6tTro3YrVJdYQ+pf9ShSbN0hpwr
CFeUGwExnE9u3noI6kn2UjzkdztfGZIoQkhirYzDwcWCvfbU1mA5/jTm1nzT+qoFj0eO3YYd5EUU
OFehxIN57vCUqsbOYrG3Z2/1Ds3+1m5iHuNoo5QlbovfXtd06ip51jVTtboZ9YB3q5aX8R+LAMLY
G0eM5+LjfYRYAOHXawHml6T8TkMZS4/8+rV//aW0xCx1v3s4LRNAtXn25lzr83zuOYo0fTBLeDhc
/IJi1ttNzQp6aDg9koUNYBozQ9/aNOCpN6BML29zdMsIxUNBmz7OWf5vlDgBXblo6R6x++OZ1p+O
vM7+qsqaK5VLEYWauHBO6Z+rcJHdax/7Q4V+pY8qvQv6Wo71f7/BzzD13BHPqBcPMW7ORgV3tWxe
gaIcUPCGSV7xb/olYf6MMfUmkPy7YNfQSJfrizR4OMofwHioPuO4+WOIqYZf2iU3tGu3vqCBRZE8
3KVS+NooOXGsILZY26v8F68FR6YLm33fIzU009XPpDxv/UDIQS84teZ5gIRWmSjzBDngedRCp3Tw
rravn0Y8i9LQMVy1gAikq7hw8vBeH3JsCRO7UvdhsFAeVBRWDLEEhQdnHSR/T7k1lCOTrdYEMHw+
jEpxR8QwHFcKs4YcOGqGEDicJJO5ljfLLG1consKQQ5YzscaMqRboosAPWSrMfS8r4AqO0FpZC3S
deEUX67uPXVyF08cNxo71uxUqEJFtelXvB4fa1Tdp/Va9O9uMccEddOFXVvaVUhvHz0fw5ZEZAJ2
2f+7S9c9bUCvZBvYlnBv+3u/u09dX1+qbZ70FwK7W9iVxrFpxs/MHA82gPa25oU2tGB+qwdF5c9U
qfvR+vnLz+3CIi0mxRBRKEWdkaQmF/9nghwGyTi76QRUwA5oIUZzip57SvfXjUoW0DGCLSPXlAPz
KBKmuSiUmR9Ccppk62UfHBi/ApIpxAWWbIVOWwydWTpdyE0h1xqgCFoqXdzWmTSczEojvcsBmd4d
HNN/Dl2Lvkg5M71xUsGivs8iMqyP7qKX9u/xFcK+mw2PqZzhe2eQfLFwqG4zzHcJl3pc2RJVrhH9
CuzzkfPTIlmS0Vr49ZwDQmyvWvEKBe2cKFv1EHVzGPPBDF/GtuG6ejMMt3LNK+HZPYFzfdGPFgBv
tbmoDAai+DvqMVk5MCif5ceZTo721ko77k/xJqJ68fCbD4/vYz9LsTarlO/9ndL6kIpcBPfX6na9
OvuW2PNbwbE4lQjEL1vupsjYkZvQlBP77b35fIw2oltLwIQ/9VIYtjltWST5Oez/Yd3t2C3Q8P1c
PYsxyAs6PE20iOv/rFshJJole+KZDXE8sjFJ3MogVEDtKV8tFPZdu+n3aUJ5glBLyCSMWoDsh5gb
feN+SugHvTAX02KvUt/p5hfPJUb0Dsk1o0byyrCrYz4StTjlKskHZE7wYSMBWjbMS/QiYf0wUWd/
J70zTnr8+sWWTzuTkSHUg27/9aQBd9VhidIidTkmG38dNiUROvC0hZjdUiHiTk3hIjO4Js2t7psP
AV4WguUg46CgB2k5NeuQn0yv8//g0YyfRjNx7DxJZUL6IF67j/NZ6AnKl/9ottoCSb5DO8/aix25
9UuiE9/07NJZEglqPyhy2f11TukAGTWhpvzNyppPAoOUoDVTa7sklcvTp94yaxQ64RVj4GmTs25a
ZsGMpwoxYwdKwOaU2mdPn8gOh3ihOODqCpQ/Tju8LY0JHH2rIYPulA/76WB13r/PX+faVnxzPB0N
xlX1fFxgjmR7wpi9QN7ezIw1HPdFTPIU38nukaBQ7UnXtIZfxRpxoSnlznVT7vtoZcV+x1cSqWN0
d5sm1wsLISTDkPwDw3V4ccZ/ImCa6deYTuQg4GRt4rHOBLnGb+ezj6KCU08lPOVho1s6n/AWL9wi
eoD90UW4RNYRtoqhqIiHGxACOWC2/wlAv0EqPqjiRu7z4/9t4ZWUEs8W0E2QwUsMmgtiZw5t4cW5
brnmV3JeX7N1yY5s4yY1Qd0J6sDBAsqB4LR3OMMVbr+B/HIgqsG/2V5aDplB5mT/JzsLAEy31WsT
xpBwHQmuIbmUaKMSRf0042cT3hiphQb0MrnkbDhL6TIp4oXlp6XBBKzp0EmzRG5PQdTsZo7MsTlK
rAmIJFLdiG1LGjJc6KIp+mMak2/gfeyED/G613OlZ4OHn7jaB2jaetP6Mqogy/4A35yEiU/LGd0G
Ycl+G8rUM4aynSADMHqB8bUszt04Ax5cBxHIHTgxSDi8habv9LOW3RW0aik3YvU7hfCmEFVyrjKU
WZXeGNLlqbjLf0DgAkeEqYji+K3bIQXSdjZH7lb0/yLoah5XEjz4/MjK1d+GpPa1HgOkGqIspoUq
ZsLMdkADRMyUPOvog4k5tq2/5B0QqFya2qMvCL79FUj6PN1N4Ei++M7Sd894GbCHnow33WufTASV
+/OJVEDv1IGUboxDIGkpFe5Pd+/jFzDYlHy5SFpYYd9zrI2K1e+m2rONlQSvUE4yYnnpWltaoIaZ
Gl8kZqb/ozbI5aCY/2Vwdhvp+TiXIYBxGvOk/98HaZ64K6HEhUWEM/AtYcbMnmDqDwmSgDQCNp5u
w6OTfjyM81156fzRHlRSn1SQJthNdVdELdcaMoGglwz0EuKxBQQ2Y4w9U16V+eowJBU/EYukZqBe
HmBamIYYxE8bDgIvcLUkWicHXGXzPScLLWlKpeqSoMPIaOULbhsm1W2qqBvkuz28MAUtUar8fshC
6EafKlYQkiBbvzhst7kzZT2QsHc+9KuUwIJrawe6LM0/loUnJfbq41dTGL+4+tRb1hHYJV6Cdzgl
oGUwn1zmcVcRpAehVpsGLlcQWTq0cbPBpEqAFwqQHGECv09fpr0tRa5Zjz866TzVq1zK74RPPrcy
F3IQZpdfwyk6LQChayqUbpGEep5eYH3VRfwCHzRexH6MsiTZWsnSc/+dp1qaSiHM1LwZLveBld6U
EuKfXho7rx/CRzDw2C4zjs4jdTOYxILSsWxyT1iHZtPD/7S592VgioMFTBOVRFuJVQzGg5LNSxl7
L4weIWp0Dzr0Q7kkB+bFK0Ky0mzKK/pawcYoGksTK3Y0r6rBrri2SGgKhinwxraQv1pMyiKgj2mv
CR8TMS86rK++ZtOFPnOkxwZW6Ml0yyFKLF1A9jKLvKtmlX/dK64PyxT7Xwn/kBM1ii/+SUjdprst
/5gZb+kPseoNzYdg77O6srstnZPhn5CKtN21OefekRiZjxVayib0uGl4DEapqdNZSsTE4lqNOHs/
ScYAXs6iPkcVGdrA0pRJ5W0mxzy686QhywRvY+TLtBgW/hahJjCOPGV09eeFdy+z6VspqYzGUZy/
8tU4/9HQ/8QUJoJDP/7kX1LGwlB/JiYi/zB5jlwR2OsMaqUf0G577DPXS60zVwrDPCDoSIslAvGf
yB35ueoN6OEiBJ5RzUrhUfvCB3Wt7UkmgrqPSvQchCS+kOH1cLMr9eBZQXthNzXfcdeIlUhW6BM1
J3kGrnUWXBYPdAqRuG+xbM5jRagKWughxmsXQpb8ERT8RV6QMk+PPaI3r3RVoUiwf/QgWR3JuoEH
+2r3Qgqp4BedVuA91wl226PFhC4kiEhueek2CHqRJ91mr0H6sk5WoWPjcnYsPJs3/uKFm2FYR4Ks
pMM8f2qcy7A0YWf2f4Gh0KpZbagJoRymhk3CPEzugenLdJWG15WzbKsMqrNyqxcT/FFeMlncqPOg
x3yHM2RpRblyh/g/wGqTC6/WU28QJ3bVu9oHIsAF2P0P7QxVFL+j8MoGhqWu1vWbtvpKr8GyzyJC
3DG5dh44dBsE0+iWZmJTnXtO1/RkJcPmR4LbgDDUeYoUZQJ6xvUvaMbtE8H1kbiQaR33xDQqjAlx
6Ee+8NgMWXLW+wMKYR0UPbn5MswnlioDkuFC87qQRwVHIRdHE8cHaJ40qpUEEpiT7D5LUpO/VfuD
P6KrrEchyZKfqF8agbs5QHwk7ZCr36oBfFGNgQAdE00f+5Pp0tc15GF/iJcFX03c9EKee8pKc6HH
3UT0h7RdrQFhnVFjpxG3Fj5JjR2sFzVKrnQce0Z3kD5IkiYOPhHn4tI41mM8fYmHQ5Ch9vMGO2Ri
bCCgbrhyRtwFR8LW1RmhsWQtBuYui+asCUcLTjHSl3GYPgotiHHg6QaO2ek5c4EXdzv/UgaNbd44
1F7Rv/Vw/p5tnazKM25EGIX/foXwQ6vNvpd9JstFX7rnQPiOZTUiH0xI77kTP8VY9pgUIjDXV5sk
zunwGnXGOGiLBc+xYfjr5gV11beGe3B8Imt7nmvDZpnqgIWdPIH0kJPLzeVVsk7hYXUO39lbZgEt
75bK5gK2a082Eb+GKvkSIBXmwe67CyEcQvrAEjAyM2JlpQ4Et15cuc3+X/4Zl6PIjdjgGb41gN9f
dg86gl2inKvHb88vyYkTS/xfuvUKg4b5L/WP9CdjLsq9extqwtjF83fgEHCYtRFQ9QmokuIdJyTe
G2O4jrwauSjlWJkFWvuaqtC24AphUYWqUuHtqNHr0om1dqdm5UQaS9FsGVvSA28+fsQOjqMoJ0cS
UCcL43J8JMYXL04GLD10SpNLYupT4FP3gpT5N9iPqDH7nDoUV0MqjXIqq4WPxDmt0faOrQ1j5PPp
11eT9TsLlzNolaJLGTqwGirntD6cV83k0suoLFN+QqPcXc+7rqdTfBn6QsOUyK5dwzHDdpUEZi+T
05fOvXpDtxdz9PCGn4HD3/mzmK9S5/Vb9whrrTsbHjEj+dMza5ZFNMP3hLvhuBEo26i2/YKFwZWU
Yk885uE6sCelt5NBGCjtX7ar0VC1nyjDLoPR/btVg+amtBCh3c5wBNxOTxaofYHjWo20lQ/T/62E
YSVbxtZZkJUs4mM0yqwpyhe04t61Gr85gV2/XvSrF8uAd/jG3Y0UzF/86zOS34ai64BObjQCnv9A
UtO6LaJUA9jhycj6MEYS50fUYgjWenE6UlLtstnXHJW7RvYFa/5SioP0Bha1yOGyUjp7Pfq/Ihis
RR+9Q4EvnIRa66rHttN0qn4ju758RoiQBs5iicq+es1hz1KV/UYfwYeskLbDFPFb6gid2MPScSS2
kuO+oR0/VNcsjhdbdEy2QM8MucS60ykM+tyDTGvsvE5hcIB3VjGqVB0qXv+c7HLUOkqK5Rt/Stuc
2KZz+HIkm1LslJHt+RWpYt4O/CDmykst6F56rrBM/u4lnEdSAkwyi1dURdZLznMzQUl3XNpWme25
gSoroMsGzxE7iCnpfU7lebjZXK3DOU7bog4kPIw2C76K/Qhj+cjgZAt80YiojO2s4jl+Qtjp5xJn
cIYXpUCg0sAoQ3gFIbsGut8Lsz8D3e2nn3838+v8M7As1fbyNrQKS+OU4WVyOIfTf3nQ2z6Oro5+
HiNTIWzcoMCzomtrlEdvyiDTTkZg5vtLv3ZScqo+Zn0FkDHUc/UxpoXeznwf2Blepg8Ztoy9VEzt
HOh8hc4j5OEnPhypsM8h75Nk+AhwmjlD3SDQZzEKNBFNM3CPpIpfgviFjnJwD8zQREi3BMntXG1B
x/QL6wK632YLiqFDJX76qHlV1Fm2gZSQoRLisy/7X6LG8K6jycnbdvK1D+Vi7vSobg+QywOG5xRp
hndzIGwmUWm9Uyx5uBE/5JP7IwLhiW1jF6qI1Pcwwa4CCpdlJO0t8egfuVOwMBcROpb03G3Vq2wG
AZrtDOIBBWjTNhgXBsrgyDH2eYfaIMdo6pk5ZJuatYHzuMXSfjqqzT9NVeJ5UZOegEyfcsfiz3V1
gBkv0b7Hk6Q2AOxr8B1kuVL2yHDthp7qpuFwZcmbATNH8KM9zahSTfWV/onzp+qOF8rX2Y3VgFzR
v/5YQTP/oafHryxwWZ+Gnb0IFBC51pq2xZMlMPAYVVNNYoz2nv7iEZDT1XSkkynHJ7cqqA66Lj/E
/KRhPFRP61KzsBjuLe4ee+3KW4JJiHQOHHwrVZZzNflF4WxXk3SFJsloF/+4dUUgrRmuKduQjGRi
0X+gblW8M6MTSNiw5kdUzNP5ySrxO15CB75uGXj5b/xk6qdWn46eSog9cd+yzGk9npT4xpTkkqEl
2i3hDYlGkPO7K4okYJ6OXmi9s69cN7R+7/2Fh4LarBRKRK8XogOGL7BRVBXsvCVxL2pg8Y2+Uosf
R0dR7lJ9il06d8G3LzC/jXEJDvaX+QcGbchQwG8mcEZL/dc0lxMcwYc6CzoYipGJ8s0u1V8pXhv2
Vd0O4wVXVKiQZ0K3jW8BQliuaGhbMpDXJ+NR7RHUbmZHlvAdpizgSYwBRFq9WE8g4M0RpD+GAjqh
651VR4PTH8HTGoGpCfnNI4TAMQ1260QAD0us/7IbZDjC2j40L1AFefgmFdQzSl6uwhedjn2jQ/Vj
jsxO0lV7LHiGnSyGm3zyoidpViidWWP5bWhgGVkDNUV1K5xW4K9D0drWu6fDqVs01K4dz8EEDBvQ
HnoD9CCYN+7pDDKveF8fUe/aPu37UqBzVYxECYY7C38xVldX3zriNmfWEtMye5t2SNZfa3BxqVVy
dcfo2ap2/If8Pa/JMnD0fQ+6SF49AJUjab8wu2AIpjim6uXC8onxG1zgzAoelLTilJA3Mn6Zbt7q
7HPglkT4XfztuQW4ZR0HnL8y4vanidT2ortlYn+clpjVlabInDDq9u4vu5CY6dRghi3nhqBjGLCj
hvC8dyFH9KPeX2arVImD9ail4jWSKSz3UdaRVOv2ajn0iQipmOrs7X3T+Ha6j+j+vOcCO8gcyYK8
esqLVoc0vo+ILNa/Q/Jn3QUEdXzMaQr0Rq1aY/jWrhZwQPz+Ed2AgWJglEqH5OS5hDPfFkn7QxXO
Te7Tdw1gYKP8/Jb9Tn9PH+GUx/9QG8jQmHK7kuqASj+RcOj3GUoo9zbvIU0zgAsGyVz5sLJ77LOD
Vmql9KfuXvxaNPTTxgpq0KwlYug+EWQbnWv8pq6vemz69MQ4+Dq3ATrbwBUzJBtfHlozZPTud4h+
TLf1Yrp/8WjDqzt7IRZ+5XhRO6yRSjxgBH2/I2+9R5IAcVI6zykN6HieMS9NOzpz/aYnwEj4Dat2
gyZyleygEn+KxCg5kb/RSgcN5/GxKUKkFp2iAI7MZOiH3qQ3oysY7C/cd620GrwOgm3iKCYbNcED
ZafdF3CENJh3gxuHOKG1dRUEOW0BPmcP0Ji4PixnD5jL6w/bc9+l3GP4KKSxJ+SRUzs8gxIMKmJx
ED72OARriBBULeUVGiQf9o0U1LiEXex5Spzz2XhSXvOTOA/bRxwP4Ka2VX74XGrqzqmc87icZDYd
nNwErUmz9czWG6QToe/EVxd5LuBbu054xXJSqp83l8UXUhjvefNmDVz+s+OWHeUBrZDH9QdhTr89
W4Q7II4CsbgRV6+Kj1RHdlWdYF8a/jOeKkufssIXFu0mkgq+k1MGiNljQl/C40evaJfpMxSNfK+8
FgVfFAqxDyC427lQS4x+i+XiLBwcMS2qNaZC7EzlNdUp5ZCvcTVdrEepuBz6Lh0EQCzubu1jVfkG
kIMkNcc8/T1ApBUvJKpXsJNZYSZv6SLcpa/VTpx1O1U+Jh5WuLUsHWl0pBlwdW+5AwFj0d66Pn3x
7wi+LbyAq89vJSV2NJ2AG/kKyAqbjnYIfwlFHOdpB5ePoBSuX4rbonCWs+98dZvgaZ77vOJxXSYD
k+BjGhkSuYYimjbPT0ynHmlFuYgnV73ttUyKKfrwq+tS9uyql6ZAvTFCBgL6TyWgMPaPE2MIhCM3
Q05ZZO+6FLRKlTYIya5KF/wb/nSx4ufwzCvnRpFc2yoGLgme9rdySIBJePwbUODBl3g/ePoIZ9Zd
4K6v7Hd6SFewFYG+b7RBpx9ZpJmXQrLzlAQtisrXxizrgC+QF0qJmTg7ejKhoY12Kmf6PhPAV4U1
OG4F7Tr+DPW+mHKTHpiaOYPa80D0KCVgyDglKxW4Mn18OtuynCj3K4oaCrIVnouFqskpBGTfyI8m
r7ybgVCZoN3psgUMN9vdZXReEP90yseou9qMHX2tU0YggkgD98cMR/EOJsS4hAlU1JK/EaZpkksD
aPwAtwQSQBS7yBPriHw0ar1Z4ahSAocv+Hw2FvvyD6M6RWutmbj9e+hAlPu3VPTRvw/YVGTl96zK
+q3Kuo6XO+A0oeaFHi2sqIL0C14qY7UjjnA+DHVxy8CdsKVHy4afMG8cy6DVVfw1jNEZ9YKdhurF
qObYsdVzOGJ9BTCRLEDdE05xiMjrB5KVaie0Bri2TE9ykl8vkJiu9tFkbjEv5Xcc/kCD9TAMHCXZ
OvmVm0AHlefE6rfHyb5NCrze3WAKCBEd8G52AwS/Whl0GXbDoeEd5NiABeEaEJX4AgyW15KFAhyL
gn1MOwxctry7LysUcljqg/WWZspcLHCq05SxPBlmz4Rzi2eBu7Cy/XBbJl+8iGH7JpVz9V528LLE
c63AbtuohBEopuZKcozPZ3okFs9EUxlDln2sGSHp68r6+jNXezvlWMDuMIQZx5yPbTAF4+qHkoQo
jqG+tm3c42e6CzNvvSdF9W8lq1OfEQPC5hxEtElRAjXvTPau+MKggPh8KA3Gszq4TRxkQHGsydpB
GWHDVoAbHYLalKdJghlNrjX3GiPwnfHKn2/+ERQhTAYm/rTFskmbhkgORM7jRGT4gk+O2k75fZyU
NYZXQPUZAA8O8Ff5n5mxHYVgELoYVa9dO9TQjxSl2ff0v5ATRmZX3z4m0mHHGZ7IuUphSDVKXqoE
886X9TsBgUBrs0a1T7BmYJljgHfXpxWwdJgU8PQwhhMxpLtM48ZtSkHY77UeES6hcW98TblwXGBe
mBpQr0N4JoV8BTJMl60vz8qaDT4InSK9CFwhJ16Pigk2bO4/xtVz/oOrIIbmEEhXBO7q9WjnrG9F
4PgUZXAngsS+eQi23D0FZpZ5oXvOG7GroIozTVZBhChnuGNnhNpWISrbP85ARyfTKwWIvBT+nLPq
KFV5c+nuyuaMMpFGJauyBiQpmqenu2teiLvPYTFdBbzB+YSBXCk35njKmo2HAf28H57Vz/Ivrz8Y
jW1+tgJdKwVscuCEUtfWRXTJQtB2IDJChNC9zsfMEHojm+oMLayHt65q92aJE35eXhQJ6FPC3S9E
tVbT3pmTQOO+53k1ZTa3mWpej7RrQ2XNCpuJOGJ9xa+vfiwEi7AlDNfI6W+1T913RyT6ToZTuVK5
IlleFmqT9yP3HVc7JVaeZ3m6zxOs+ChQY0R5qpmohYFPUmz1UOa2KGLdY0gSJ8ry5SocMTqbNYBS
nncqCxCwk0YfqyKkROXgzSM2vxfbEESHY42VxHdOIPDWfZpx2DSeoUVAmtyYixxnpY90nhE7UJNc
DqFwtj6CbKSUgV3AbiEP+UBN1mIhMVQhbF+i5jWfRLnxFeQZkEottL34/jnSAXo4jdQV6zMl3pnF
M2xBf6w0yBZiEEOnqdOz8rm3rO9NKdepz5gIa3Va+7tXhg1srJkgJRb48XjlmqkjMPn74MoffO9C
PAknInj0kOMA5sgXm/us1LLceX+OuIzoMnqTmsOwiLiE1V7L2o2saFaUnriIhlZMAoSAmyveaen+
fCHMDFP5baNV1SU/QtpoN423UuQXRFjZxBsYaBvpq/H3+XOxXx9vzqIm+IjQofYlYKd3ot+xonEc
Ir1Ab2BdjVtvviLiEslAX5XJX+g7eaCqxBXYrA2TD5NtkvyBNaS+r5NEBXaIHlwT6En+BIxljm4d
TfTslH6r4MVPYxEsar/ouRcgWAJ1Gpv1ah8Z2vJLZ9XnX2h/rTFFrBbj4eCY4SS0l7FxlJgOLjZ5
Ig4avx0hiIBlyHugGuHUdDmlX1BQ0WJtyFKwN4e1/K0gwoY4YCjB0NmL+KNbNu9LQAtusltci1mn
B+kBuvV6IdME1N52hh8K+ENip+GS333x7WcNvnnCCuEzFHr0L9zQDC+5Rz9aPXpMLowmQYL6Zd9K
NoBptXlgbPxhuZ7oSSSkNkuJDWxdNKvKs2UYQQs2cpg5ZCkgjdXYR+eWGUItCH8C+/J0s7JqA0SK
ePIobfjKlX4a7UXnCyS14kjUowWEwaOvXx59Ihbn5Ph/U64qgx/WsMUMsaQf2ukXT0vnN6QKy+4g
J1fvF8XiQpw5LoGyIZ/cFNPrCQL+RzynlilQNMHvFFa/wJliT+PK4tNVBkEFeHZlPT+6dNoju2dO
4f6vUAuOzOCkJ8sZyenZTqoa0SbfmrSgGsSivJEpeOPbY0uMacqBTV47a8GctMKfh7gLhkyjVv3w
T3J3MNbCbtylCzep6He6kzMD49x+Mxf/Ho+wrxNPGJnd0C5lY4pjUTb/a21dAVKINr1aWss+Gn7k
iz8IOQiTmV7AjlOTOEZY0EwRY7u8XOfO8s0y836cEISUgQp9PJFPza/k/KypQOampbCdRfhy2vuD
6frWTqdGqDCfsKEWfN+obAvDXIFI/SvuujK5KqgTK03yW0FI6Kp8JFhIo96dCa43838/C0momnf1
Q8RWLQuro+7nTi++6nUQtqEW5pupy8MZ+nMRkoq0Qnpqu8QXhxLK20Z7cyjr0lLw1QBmJZ14QBc+
eZzeQk/y6b88E7wf5j91u+ov+bJPTyIs/vu1srnY/wAnE2gyuOg48EhPOY1R9TjKejEzSdZTH5+2
cEuhSGhXcYnZZQm1wPBZ2v22hdYNxzkFIcCaW6dXkt6XTeTnygMoeddcHYbHHb23FGShPdcDhmO4
NOdnIotNGTrw3gsI5kRFaN4CcavCvq5zyEcALXYxssQT0WssjaNtztziw+I8UxP58ztK9FjFF5ic
5Mpj1LK/2xvQJNZvxTksleGQwrXvMkVsWYlkiN4nEgY2SBg5oDKwoeouwBtUXtOPu6XAC3ONLhQQ
k7Wuf93y6gHgaze3t1b3a5rxwTZvh1lefSf8X/DisEWM4Xnag83p34pQzh9QO+L8xKiJ3bR60DWM
eNgeYg/WW9iQ+Hrcsdqvp0UHc2+thWE9w5T0qDLd90u7GD/4JCV1awUDkW268otZNhLj3Q7VJaqc
Sd0MN3zU7ZcMiCHFDjeaTGjqmpOD1zK2YMjDOmiOL8wl8dAFR4c4JFvHHJz71STb8uUFhwTZjWPl
EgkmKvfn8QZHsySD95vFleMe0m5XtTwgu2SCfE/bmcA+3DQq3w/TVtpCv4lvvb7n1hj8NDx95HRC
4w/QGAyxZlHqSUiL2DGroFkfYgV0j5vaqS/IfkQ8i44N/9yhJfVHNnnHfaVQOexyXvWRqhNu0ELb
ffPOjk/p++VDpSMvZZzuJ7PParEu5AUokT3RXv9x03ZxR8o3KIflD0dbQWJB1zQh/4hkUZL+gkQF
CwqDlMVeUYspGotd/6fwdhn0YwXqHI5CwVlRx8W+gnbvTOUncYinDlvXoufJ+TZek11/O/wZepUM
dIptA3YkXiZ8ijXg4imnGEbkHUNNr8FngikM/ieDmP4lyDAj6uoz+jVGqL+UHmohyDxd6/cqUjgd
yJT8ekpJDqqRiKP6MlnEmrFhAqwCOOOdgwk1HRzSLca1tBZl5WxI6NIGJxdFc71mZ6PFMt1sxjYy
gt0GJyw+OKbLjRgkI/ewSnhgV9vdXTpsrWS5sUtPhvGIFK/T7EzfLbUG7K8ynEs6HJZziYlrNkdf
O8kFaWJvpB/M5ZnOvzLlpTm32xcZCD2djFqjhtuOPwb4Mdv1NT1nurXr2oVzb/zwjCjSvrsP8V2P
kH33JCTrp8fRe+NQu38zIw5gFB7mQNiAQiqpcLdU/7I9adxTxRzqX84G7lzMHyXM4AslotMrc3Cy
e2Ah+Rv0rAaa5k/bTEAR/icHhNg63ipO++NdaCql4kPch6f3ngbinF81fjTfL9TKYLo6DqopW4sU
0prKdf9/5IGrRy+uY0gmsId4lcpfr6jputU04NaJ6QuRkUY4+6tp+x5R3Egur2EJ9xFUxylJxwud
2U8WnmIC9lfuUKQ8LgiuUsTEJ4EBByr9u0aSpXA1mGawZUiA5DwSRasm8jJ91F6HR7lW4zpy5AFw
ym5C7/eiaaWpuiVDISbN0NPV15m7A0SRHwPTMwAmUCxZYxjWAbm0VTz7YJaEFXMYHVdVyvAXaJj6
+3xUKHr9+fm+DHtFez7pKaMpIBAAzkxtSVOkXCAzC7sLLUI3MV+IuXVM5laFqCKBu7HMw34SNJbT
WMhNvreIi1f+BC96uvad+bNjhZZYy3fDNXnRESaDjs0PTYxgV6YpK16YKF9iMJyz8bEq6mTzIGH4
myV5dsIcrxGJbftdcORdIjCIddaNw/fwmUEbt/Bc+oCxhCi2Otg3ic7qFrO4FYBLFehuK2jiV13C
xDiCkrA2opVG00/06MBR3AO+uBblbwvphWJddHRf3+yXlIKtckOR3c0gs8e9KNsbd5V59LzWn032
9ZVV44XGuEP2FR5iEO3x5pC9xpxSHn9t3psbtMT8OXwvP6bzE4vAj1FBiEvxiHgobQX6MX/0pkoq
I0MSktvpztVkPD/fGEXJB481+RitvMyw1EtRwrCzHtp4ej2cHb+Q6w7DFld7dJ7UEQb3/dGidKpB
iETXNmT75Ftvb8ZpraQQ5a33uwTblhJpOFiP2VG9SUCzY98V9Xmwuehp2oFsEOGwgsF24GrIXIHe
SQeejvZAqcpo3c7K9apoILAxTYB79KUh1XRElN+9CJA+tD2pifJdHa5XFn9A5rgjuVdkU5D3QWGh
ELzEevLy3V4ijGUyyQqByLd4DnMmvjW2uSyRMPGiPqFMhPD0rD6man/wb+3deXfbCtI6gCLp18w8
/RJyixtKFo/ECNbK/usCbVXgIZylRCYvDdZEWbZCl+2+eFmUPnhvglLGas9ySf/cOsXFwgvlmwep
iESKbsyYtFD+hQaLRkIPtVYImBhSP2HSp9cEaXo7YXAeZ2M/7/knSvrcMJ0rXSOPV/Jm6prA9btn
oVl/Dsi+52K9sV+6f8n8OgFyHAzu1uqiXDMFq7ISBi/bJ7wsvDUwKkebccOkDS4hAmahexKdm8dQ
bWbl7XB1XMYYtF1Y5gd6g6wi/ZXKIVX6yGIJgxTMUQY/QQyQMSH6hhgkxt6Uk9p2f4pBXittkIP0
HTBDNsYe1FlTXUDvcreHstrAE+VJC2RV6R+USabfYNynwVUWopGHoKMX7JevG0lc2mp1SZHg0yCW
MYoy1l4Vz9yPWQ3JgCZGZEcL6W+5O8A5yrMvVSloOBHChoPGZm/oDCKTZ15EGKTXU/U9sBe+L2YP
l+7qdAOPxZjO7XfdM8g0x/dy7jtACIm5KcmOcibpcAP7fZMon6+e1OpBCTMxyjAoQSxljsioRxn5
3UAx4lRNSmR9qYC8Cn+4rIC/i70aAlD/J/9fwKFZ2CNMr+OvjT9Prj39JUtmdvF2Uc36cPIalA3r
wj7mUfHs3NQe8hSa0Z9V8TmBz+ZCqtMBzxwm1f01/qlcNwOr4+M7Ada+SyuXWqzT7P5pdEloqFqo
jwuBgsWVcD0dkzKNriOJmBqV1ZbU0vhHMpC/j97mJEqcVuzL5snlDjAftEGYb3rjVqysq3w6Pd3d
Zht9hXQQmMxWyuOUXxHTIxjlkBMGXbXoYM3dX6vRESdUnwyOAqClW2KpmWdpIta3ui0QuFFseHdj
4DuMIyyFx3njAcQZFac0XdpdXTKiUcL2dWMf2Xl9HIbOuP6lmnLGplvAoWrBYI9tXfvrABiz4wpo
ynWoJaO0Kbdfg4DmWDUqPs/1ERLTQdjG2p6gcyusA60vxJUL0LwETCv27BRnK3xEzNfq3EQZ6YKV
mi+xAke0J5SoEYwTRrnT/vTSD30LbOUETD8wuSkQrlEXYSKJFmdaEgIRW37Dcn/tPhrhywWQ+RbL
q7fMY++U/ngLNIEgiSHHaq/9EgGmulNy/6tb4rKzSVXnSSPyrr/zLBaXtLLXfPr0FKkoqQDVzaer
wjL6S+k4eoa+tZryHyNonmAbfBjYLbI4gzHNY67AlUfpKdX5JWKN4EYZfFaQxzj3mDH4rb3Q1iZy
3empJZc+HN6Zv5hB5MmGlDWazkSRYMk4CdW5X7cKNeG16nGuCMI9zCee1qXEbP5dmIxKV8TlepDB
5gMVT2SP8984n2HZHbMOuBuM/k/Zb5AOu5F4MdYP8QeJr58AbK+XTlpV1lgBWwqLw5eFyaB5E+Pa
dVa8QODNYFNR5thfw7ikbcB/oMLlr1rfd+AfDcph25I2iuzYIAS5Gp7dtCF79zx2Br1eumKJIRCW
gfDkDkyyoZInELgW1SpwMAYL0cZ3RZ7fOOkqKCUYxG7oprsSxiBekiqtBlwuqXj/5BsNcXY2YaCN
BPGqwUh2yuuH8YxVBTqsZXI2qroXhmSBnCmTIt95YbLTRPXNe6SeIAGvsS3iHw7lPk1ftlzVu17Y
ky1KGzmPsAtkAdRxRJK3WpeTzmtbX0X0yrM5Vo5MbMXxY3dxwFXKduaAjgvwdiUtnuQoz9V1B+J+
wr4yv4aOu/lfOmEQrSbgYnvghtaVuOy1O93FJCZLp7hUNTx8FjtXPC/xFEu3DBUGT7dkFQlgZ3Y1
T/5QDGUcmMVz9Lyty/MnpIgzfwrHcXOEO1vKJ9g6epjXGWi4VPyhRT6FL5yAtaC/bTnapGNcbW7k
uMpt2SwqXHbFPWeWY4pfS9foETbfAOHR9Q4Zd9mMZuoHb0Gt1hG3w78vdB3Z/IwsOal3SvYMFCfu
jUbTRnBxyqe3J760q5TA+mvT/C+se7GA0xdxojs8YSfqV8ZBIAjivk1SdmXQZaxWdfgwbB6gejNq
3GWvidsWJ0HA872+1ndTdopv1I8FxyP5VxGK9czzLQDgX4dDVo2OxB1sT1lAkNqznA0eFrzgJYJN
n5oyxlEUoMJBkCvqlBvzyKIA3nr3WNFCmRYwTJPx2BMuI4ff5E5QGzCBvMWAMCoX1EhmRArJNogJ
587xycM4rDLxCElpaI+wqeDij/aDJXrvAv5+STBx+9cDKDnH4cW+BLxI7NWZZAV74JSz0qtxWVGO
r6fPBrkrtKkbNoSgqcxZR/b7Nulodyp3dGKuhTgleuZwLxV0r0ctfmYmGvMNtbXHbresTkCcLVX6
l5Joh3rxG0d56ZmETP6hrOhv9ru5uMI/A4M43nKgXWv589Zn+5fUzEMKOSc/uPcqodbhmcsCLlh6
MHXoB+8Cr/gYYo5eDVRs8RBaD30OzMKzZLenKMgkD9mI4BKER/GPw+XcuBIqXM9/yxVikyfFYXLX
JKGn2Ht2HUiOa77kANt0T2kX6wRSRR8bETQs4+NY9bGEeL9+uIi1uCIVn/rCKmpjaxwZmawvdqF1
p7eQOCSf2EKldqTAwZ+t2DNiZz26BAj8XOvPZzxgyPYBuvoj8heHZ/VYNnbhOiW0Cs2Co9aEBAE6
FYphfCElk7aKcjyXtf+Fg27KQpO+TIVZdJruDQL6/ez9lmTIQH0shurnz7efXdT6VNMRZQqMjzLc
nE28Hb2DztMJHbAvUA66bTqvTXDGJtj/NVBWUE7G+rhCPlonRrbTN/cUikkl8Dnq4VOoEzGdpqKo
Bmz8uuWsTh3tc9t2f9r5umahma1zbmQDk5ODi+SJM+gnY2PxLtgFUvE6uihpcu929H9Vf10FMoqn
dsUXMqfB+AXAwcvuc+XXBYCRMbBQfjFZPpigyMs+Djr1Ch4eNQgULvsE3SGSTaT5DEBb3LhgmUB9
FSXZjc4O6HtKnGsL4f/wsewU12JZBxUqo5cA9w5brWPKWh7jjIvR+NKcRyAUra3y3XZ1VMXka0On
zXtP3Rl2nKSS+zUUZu1wd0aLTMi3CnO2IF58u6oPUCWSM8La3+UsR3K99YpQQZqmZaTPIhiRuwvD
JrJqrfriE3unjzA9znxBFiv7Z2oUWRskMH8Hf8Q6mfyisMWNNdnRw43rgPOFd+/+T2NFWOLNZIbP
59L4iLjPtlqn5n9xxCn8l056FkyfVTNo443IQ2nlkFEzIQNh9ST+7DicZVT1jnGLowXWedOyQ8id
LmF6NMeS38uZghG5wJUmIKX+lZazTwSmJ/hjaODQo66B+Cj1P31fWYX3U6kSD7iewfC4yoyoWNZW
C8gDMela9CIoZT5lFGIwb3TtmKyg4jBhsUCeGb91ZwR1mH56b9z4TBJdG2gy0C+mxWHjNUwOLPWJ
Gh6tYwgKzppzI7QEfzynSxOE2UFQo+ri+WL71XkNqf9u8RrFWN61+ve08XbsP3cBMPz94pm0NyeU
cwCZTJvrO3Msd9DdA9uBnaxRk7YdAImA2xf1yo7oEnRKg7nQxFfB8L7WQVYM1iBw7wlmOqUTolCX
eo4B/pktVESx290OzCJ6FrHjDCalSHH620YESZZe+iHC8yCnaHirD7ZmSS6rHqoRkk+XTX8IO39l
5LuA/ff2BBYbvdSHoJvyd1orATned5DK6yzQVaSV5B12+32cUMcgFNxpTRnP8XHDQAX0u719qH8u
MkGQXC56RmB/WOuVY+7FZV2EniZl+djy1nlkLNYKIsSyEZLSTR6JWUlmwc23rkbUTFHff7kbesnY
K6d+c/uXH8VcGJ0/8kYKSJllAFAUSollM+ivIjvbkKHK83q92w3/0s6bIb65ghdsVaW1SLwoyHo0
FcsFQHFBKDRPWnHrGZnoynPfoVALUv+/jqM2ks9mrF3fa8DwSy1KP6iWTacNlo/NulME/m5Ej81H
I13jzinn2+1HBmktu410j6Ng3eNFrmLHtmyDj2XuACdc6tEVcgZ6jdksOWK+zXIgub3rlmQm7mOk
M4NExoboT4vyt48fkVK1EjreHe9JGBaBV8DW5fGYVHQSFHmJjJpp0vBoUpsWp+1bIBangGUIJVo3
OlIfjVOrUraMhk+mZEM5InecEyn9SzNXLFL1wv9TaGv6wFs2AtMAWkapheXWhaz+Mz77ecwlbtgd
hULOl4LrsNVbKc3wO5xxJV7dKDNYMtNQ7oZyZR6LaD5tFqZtCS/DOFHQA6b3B+DFUCAn2cwZsTTR
2bUNhvxiQk2yYEHBHKHnh2cXVOGN3u40Ix8OveJbsdyg5v/0a3TtayhzqGDnbcvSZtkBA5Hu9dhQ
swUGtS5TUoDMS1X9VyeIAqZtMo+Z5FYzjXHmPpgdzEvdGVv7lehkDCsJjhx02VrGgoO2+r3aqp9g
Qd5cqdWzt43SnEVWaGmi1gUPzQSLaJiHpB92iuDSIU1oLB2f0DdqxFpKltGgVBHYzHjllifUZdO7
jiCYE5fSuHbejoKa/Mj9TicBIILcDbgm37PSQnxxiAg3ebJnjBcZO0gRP03LD+M4yle7pBLArdZs
0an8P+rkDc4KNELQZ2Y3RNnndSS16h/VXcZzzUgWGkCblTWnvGn6E8ST6Kyg1OxI8srivR7Obho4
GW6Jqs91H/eAW3ln0faavI3xqCsNRI7hWO7CzfO48s0D8IuqP/awiA7++B3BqAx6V5sfevdJ9tud
VARBLjdT3sdpgqALk5/L/YaqgMn0vCG1+u65zuo+KV6TPIBh2yZSdB2TdlsnSKEa4/rE2Wk9F1ps
gOBaWZk6q22/RCxIRQPY4+x5p4v4Gw1BwQ7f/CZeQr1Ag8zbzMOAO1pd7b5CspPherHBOXFAMa2F
Z1OIZpviK1PLUGiiSe/2KaX9K5BcivIkZ+71hvIar2nSBnBZOUrwyx2LMTyN5CeP76pFS0kH7NWw
9HaOkEUoaPjGDfPRoGjBBXMI0gYWjPJBirQra9q1Oxr4mdQGgAZvx8cEcndhPSEx2kF/DdS2ZC1E
lMCymB1jQ5C5lXwOFNkYddEUHGRqXn++f4tt4R3pztfOIX4/ivV3wh3CuvRvTMUeKFlqnIMWgKXb
0akTctseHVoCy0LfnnBR8mYj4el8Qn3e/jXwQm2fK0CbDlGrKXd8c9qPs9k/6XPC6NFw6BDANf+a
usSv8iLxrt+OiJJlx0atlHQdQpwZTrNGrMo36ZZAiI/jS291P5S/S9RMayoklDujSOJHUj5gZ/Pn
5oihSRyFL636X43fzcKbNNJJiJgPGE+d2DDt9TlGt/1YGbboCm4ATcgQ1sZ1IwMdK1jnR1IK3ann
G7AgyHcDyoxnuI9HE7y93o2To+q8jfD+AHbuLaGMbDYi8op8p4oo5NFX2YYuquhkP6nD00Rtc2PD
ahFYS/FmMUL2b9zDo1jg7XYsD7ivn8c3xGfc+tbyqZPzwR8nerhexpkW0SAViLRMu9BbYp2u/l92
o+xsxi2pPI2flfHEVZBE/vEThQYc+lyQO8VZZNA9znPbAGwoljQIhJY21TwK+EYlrz4/x1k7tq1g
xls7AFrMSqbcH4ONFaOmTH8DMoN3SUGhYH3gyKuRP58CEEhatZTwwvA4WRMa/EmQeMntDIyd5Oyz
2DYBviS7WgOLHgXOGs2GKJvvWSIUYF2F0dDrF4cYszccAO9VpDt6IhA1kYCL8GZ+a4HVfF8OfbqW
OtdVRd6q4qMxttSW0UCDDQo9iVEBSsU/IcX7PVRqLOMPOawDS7r2ph4MFCCqloPE/QAySvMzBx91
quQ+FE4gca6QnN3PQu/bViXtUd8FgDpEPryaCvkJvwyOo87f4Y8HMK+r3K9+W0GJy/aiS6FtsZb6
abQSAIdX7hLysSZrlPWjyl98TtoZSJ7stk9IarnGGYqfhaemdEq9nk11ZroNFvKPlP5YECkzWPaR
JcHJKmx5j3Kf2PGNl/6CyWLT5mQDscBAgpShK0f9NeEdt2y6f2HywhXdLWi9IBeBEPhFHs39KhzT
qdPOTi+eGNJO68FqhSYapu+MMIYpp6qC19hb1kcR74lmXE9UmrRCugQv37RNenPjtkZ1Dz+N5WJ+
LhSFkEa9jCkMfbwUppwVnQxVu/afLN32u79E0BsFpyRz9vgE9EE8xFctYdkdLoJNRG8oA5TkKRo6
k5QZzmaAFbykFMdiSAyH4COb0dOBJoO5SnrHMqWB2goD97xiX6IrgFW7XwCNlCWXg6ctOeMC1UYN
c318ctS0AQEfkzrUJxoSr9ddvCY1UM23/M41q1ZmnazWwzYt43ss0nQLZnYGbUKsngJyhF57JpXx
R+EEcDXm2wBcsgf9K4RGb2Vj9VO7ykuce114D54c226hT36lAaVtJv6lansPAM0HMctqDrdi5Z2u
14brej2vMhD/+CLv/dDd+LoKJGWkqJjx/qMkOODhkaEA680LT1eVFW0KmWZcmCk6fFdvXnECYNih
zhV4LSAfqm7qVMmO6DHQ3Z2hNN3j/YtCTYOOAISAL6zUfWDnuvLHN6Q8IQHLeq4pZGb5MStZ21oU
SyFIUgK3voDgUeGdShakDZtocUBtZhA1S6Ahnfv5Lk0W48TZoeYtg49rwNUgXs/Ztos/ymWDR4Aw
mYvDQYLILteNfe/XnITXkAFbxtooexoRAd9glUfQtNpNQBzjkyOA9xYcmVf37NXYWVm/tJIB7jUX
PLo6o42DeiIF7MIQAKOehQYA54mz83pqZJynb4N1mjjer8/yQV+uFgoBQFYhcdzdgxBIrs1EMd0T
phfFiT4sD7u0Nkz+p83GYIA8G1df/SF6+59jSC8TtAeQTnac9dbzSy5LZAsKSh9StbiPt0DYlSzE
M4HDAtRzA3p0h9K3znFk20oaglOaZRmg39pRSbguFsBGnpDeDXQKdUR9AOV1Kmm0bT3XJn8YA0Ts
kWGWV5fgkGrjeVkv0n4y6wS5SB/v1It0sBx9AjuD3D2zXMf+/+7Etb2eW3yc8u04h7Ej+Kc+4OCM
IpoGm0gM3EEvYWQ60l7fpiJebUWvqHWqXxMz7VdqB3JG0FnVNiIaaYo58HYUoZ2giRokuIDRDBaK
wE+WF++oyohcv8ukZ/asgiJrEtp9sIrB51db7+3BFY3BLiz5NwOqrCPg8dHaVKPFenNOlVkiKLOj
kGwIRSfOgK+BUTU7118Z4SwQltAclC84Cgf0fGoJv/ZIWb4SY3FWnRHPSbSb9AdJDSFYk9Ealmly
zw706/+loKaeXEyLRst0Ot+CZMPNJvZf9yV7EUMEKKgG1/IZNrdvhoxiF18jEgybikPRdNNQs1Yg
pzm/GCZu/GRLvmNYaSd143Fb60a1hw/kBlpK8DXUOGc3VLCFNLd67yDkQiCc/wQlZ+haJ+5ODxg0
VLCzge6q2RKaQl4bDSiUfge4pzm5Z6iQPawjuKaJ3ayvfm2J5Jx4krPsLOc+XQv9d3zYQ/rylOVR
QKN+vgZCuj3448ZkdbKrPL2nO2SZKzsck7gBCOEye3EX6YLRXzps+K/KgAGO1c5g75gOEVx1HQNK
thPpO/ZwpVMWoSHJp5ePoiuhOdMFf3NeOhphZ8GfRPDrYDT6854MWiONdclnQj/PJPuLCxslxt0R
etbi7kApLU+z100yEAphXvEwQQ+j3wYjwcllZ3ABpVZ5yJCFapzikgFe8UuklWyS2vPfDP49kAnt
bg8Pfn5ahZeEP1izZpv830oRgYhkHD3f5BwY54tb6uy95GTFlYaamC3vytlO5xMNpW3BMyADQF3A
2uSLkg4KovU7UBVqeyx9Cb5tQIY+WPV8j3LZZ+1SU5TbyYy2G7NDJpMf0mtIHofCjM528TC1N4FS
oDor4nSTA8H+je74nTGSKXYZhypTsvJmC2LRxm+XakoYQoIeszTg5dODTBILGUc2W3B5n29nhGj0
hB3B8xdLJN7U2xH2z+n8DbX+eTCwQS2scn5FQE7OWEnyueXl/5VpVrH5i0b0fJhdYs2DcUocGk5e
jKrQmG7cD25wx7mIPn8lbLx7Cq2LlcCkQkNsJBdeUqz4KyUDd1T/eIVFio6xUCCz4Kdb/SJArC0s
UzYgReAgESj0eb83UEf6K3uwhJrvkOBkYvwyUBsFbQRwz9m19WtgNiv4kpIxwKJiafUWoLf8TWKN
Kkk9ex+UhO3VqXcFEFmYI05sJf4V8XSiGFYN/kKSyeQOIMxNkGameOEB0CVQGk/o83TFuGYOjAFT
UxOb2lpKcgL+EpgeMFBwBUB8Ew0+OXesKLbhfhQU3EqyBAuUYFMhvCOegwYqQLHSuMkLQf89nHDm
lkqjTAkj3+8joqxMysGG1t6YpC/67/PHD2+nE3+PjZ4A3ZKak+bcCwRtHOicQbyKGk4yecrmNp25
TBg7eIY21p8faSRQfZvoWbO3S28Y5uvUU2XT2TfNYNHFl7L4hqayx0gW9Eh61nt4Y8y/00Q5Pu68
SeK7B+sSQIFJroPslKHMjbUiFeZMS0fsdBA8leELzUCV9VYqTHZJMqNXRJ7GH/lClAkJ0AOxPzJY
VJMkH7ipX2f/i7YuwxZdjxE2bpjnnUYDphJl7yoqzoJmWcDzCvMJcA2U/50KVN1MFdR1FRfe55lp
awHNTgdK/BpZbkEBQvBXfK7dRMPTzapChRcsSiKRrpmBUKZNKLU44ONRFgiAI588Qj2AGJ2GMMAT
Ws1loZmungHi7h+uSXFsImGK4JifFlAyQFd3I3OuFdOHWll4U25ysOJkKJr6WNG2+Yyv3HmIAQfS
9fBlXfx4/OnXowStdF0sCCAoAidw04A+axFYsEuZu1JM2UGHXTs4bHllXyf2OH2r1Bs7O1eNVi8S
5sLOpRU+J4at8OkRtm/ajlj1kBKYEePY5m95obr2cjvvLpyJqB1eAtB4APHsvFIOBYN7G7zra7Gj
AdDp0seiWuOlp8s/8XJOdyI60p0wPsMls2ixfzRWMZT+sr83u9icJ9O4YgZwZfu8rAD2M498Ik5m
kCM2ta1fvKAkA+Jkursp5DjYmqumpDJrJXkeutlwWIubyqnV1Pdzd0FjFxyrcd+cbJjHt+3h5r4D
WKWNt7pfDF8FRkItalX/+SPV6q01XjwvxY+IyCSDEb1m5dt7q5xWIjDDXJpNGZYwGjJq1JVQQJGd
lxjtki+GbI4UQjNpHda8me04q2EffsjT2CVI1DOf/IzIw8DstbM23StYh/g5+K+d3+dE2Cz0dl+Y
0aryqpIGGQ1cvKDzfF4cOeRcrmaHbNx9EI+HseqK9fAsZD0gclZ8AMwHZv2NoAZFjFR5xo+Yx98+
8qYsgWhc7X+UDjEvKHPda4ggbYBZNry/0nt1LQkex6Xqw1gCZop1UXwd2m60YMDtCMXGSEbEej8K
die1fUG5BOzfDfPF5MtGCcuWMGWcXEYomcEqH1+Bq8PTP2shA1baDShLB0P2X8FbXi2HTkFSqjrc
ooZ21/g4s7b9w1dJ8wpDYK+425k59jvrvDyBbDTV9F34XpQ0ozHUFWOxeWnWxFPvL5Rq97qw9SSk
2olkbLHbtpaCHdTIKwIY9ngTXq0/7miEooTbnAODNaXX36RpBwjvPlsH4G9F7Di3JHhhNihr1GB9
KwbJ/LYUkORUW0sDrDzHlPazHqucqQyaJmQcpZ3ielgawQ8L0JVbcWGmzwsuf3oivyZtJ72fuv+1
YaR0yRIv3vSGFWt0sRn2u4sGg71Z5V99SbyrOd++rpb4gbRi1VVMhdKIkAVxiq2nm4MS/ugl+QdY
FIv8bhewiLCb6LKMa7x/PSWNHb4GtP2YUR73vvHC4rAMfU3oqYWwkcXnMRI3up7AX2D7IynWCSrg
rRxC45j+pTaeKvvhoThcEXm99KDwaXv8HRFWGbcUA7oB9KGvsEaVRUKZPLviz+NQoSpLi4vwAWPm
XQN7qf4inEtrwfClZVb6+sR2abP4A9fQ4R9AYD9FWlX+ZODnMksuXmNBNZmIrTAyI9wUUi7Qfyx2
BqDy5LIvjQfNwQtlnHDcyfxEN7FaTi05+vAZRPdrRNF/vKqYUYUXDv4vSmeHlfsvmEBVdsytLcIo
hRXWgOScmR+4CmX/GLUnCceOKegvZa5/NJ1IX0CNy8wGzlUjc957/jNgx4U6tVvZL8DtkCR+1J4o
ISqY8cgwoaI6yQuzKtyK0DAKLBxwqUYVJhB0MwM3G2exHfCWNeaBhfgNlZlH4ljC8OU9js2jMMQu
LVBUJFVDWurMr4kkH4EhZDJKmOX8cBa+bOTCBTy6BLOrwXskfw4p59OX3PLbKRCN2Y7lSXbzyrYT
BOao8Y2LAeKYYZi4eqtdj3sZcUjZBSAt2MxqCM8KQnBeu2TnQRSq5UvevCBlwGWZyNM9wdfauKSs
u48D3kQImMWLptVz3Xn5ELf7PSlUbAuDhL9F0JQ9EcqquR6ttynAbSXfSg9iTfVjiVhXGlE7xjih
xhlxP4P0lB5OBbohjXMWNQDEdMbReqAGGLiAA2F/d2sG5yTP0RXsHhsGJAJffhNMiCG9I4Y42fa1
XtRSUtwXYMQgMqRs2+3jm9k+4mvzlvvLqNLAV2m3G+Ng0aaKgaRAZx8bqgjMlz2w0cezXH/Flvag
NuhzA6AkB0809K5/+F6i3uT/vInNRWE7J5FQLhm86z4VMRvn6ekge/AQFT8xU4h6wtdWy/29iKaA
YI3kvqkb4KuOuK8HQpxoGsX5E5/EIR/3xFlF/EN4nkpMZ8r50hAqrDQ34k5liU4G89hHcU5kVVaf
XQOE46UgOGDo85H8/u9dkNenW4aIL37vcdZ1CcRILIBqAc6PDEFhsryAc/LC1gUhayjFllAWSVC4
zPtlpcdeQyQeDWO7l175meLL52op48xoZH+1yqrhBv0hZjg8RVwJQBLvQFe8NMjqfBsTaKL41Hkd
b5GVJvgQh65HieVPIgX8OaeafjtGRiKYyULVhnXoGu+zZApEQRVGp+tzDFeuRgTcWcnupopyY82S
FmN4mw7Su7aK9iYtvbBLLMlPJJYZvM8Ag4M06jrHs6Sz+4ln55rdnfzTnQf9NuiuAs1V6nxGoS94
QUiPa/fit/tiMMHxVODbDXP3UtS84zt1pcOPanAmQOZyFVRzjrJPVvRNB5oz4hBP0iGIgrKtjfAo
C8ktF3EXTMRprNxHE4KEy5ux460bZTduqs3vQ4kaw6r+jhmE6BGJsirVTEiM8KmoRRj5zzZtFM7y
kOxcWektyPntqx+gaAedBhJZG1uv9u4xIB6VWWf2kQNu3t08SeaDcHe8+iNFYLbjoxLVf8rtQAPN
/pY5ml8Az35ioNL3cYLwtNgzbsXx5jrcvRofeVgXIUx76BEDPnzpszytesJwYvcZBKX7WnON8KpS
/GWmyjvR/+u/kUZgDOd4wOy9gHFA5QKoA8OBHAar8oofXAoYAjC+TgPd1tEAsE+psp5gaXnIk+0E
y+IJVmBZ2VZfplaXMupx/G+nDy+Cexdwvh+UDkl8PvbOhj6Snxr0hC4aPNrG2DAVv2N0+p28TXfD
cqSaHJaEeaaoYxtiKhwyx9/8hlYW/6FLBHmmeGI/xdzOI6h22X2zFISlAWxn92aOO6eZTWUhGWHW
nEXWYpwXngH8/BlK7pat1DFv0PXt+pe9e2LCuQECr7oL65Pzt/hVHGd6J9caZ7OC41yDkfptTf1S
mPXlRysTTnBp8fRHhLYcYHZClN+2PQXi1WXs6RSRI2R2Ac3TSvYcGbU3TwrXQ+r593ZV2zGpuxfz
Yey9HLrKF/7Qa3foKU4jAXe9c2uMAxEhVUFmxu/Jzw/mQn2dW2oKpcgUaEyt3nuPygr56Qm4Tu4W
okhV82gIAb4Ts1Uur+7mnIan4xfW5oJ2hG7i111VGrdUIaut75kvR9qajNF3ox76H0RfSZWbHHjk
UzHLa4W/Im0TI5tx0L8BprWwzw0sgTN1qkumcv8yBq9aS8p2oqCm6U0+Bu/MoJ4I+dSgG9nmBacH
3fdAd29D6XAJdnGnb5OCMIrWYDRzzPP6UU0SCoHZ2QRD43f4C4B0bhzH1nMq2kWByPPtpqUozpVO
LJZZa28gt6L5xeTobAD//ItUZlI5guNJ3ldoTu7/IxXqwofr1TCNFA8qys7zzWJq9Scyu1JYI+GJ
uKBVP4V5ytfnJS2dpHJHfLL4QT0VTUqyshTFw2qzL/7PUzesiWpO/QEdcLAoGAZACH2NUaRSB7O8
1TDEdbF8pxz3CnsoyhMHxcoiXf9ni+EAGt40A/jlWw1t6Eq69/lXZld8Fnu+UyAAhvYwWdhchNXb
ZlBBP5TngrsiR3cdw/4wmhkf32OCJt3KU27b363e7eWMHGH8s1DdValASnl0TJgklSRF5Vz5CD/p
sUzSsMj/IexpQEL+ZqUk0R58nthKhqE/kJGeSX2XtThz0fPjOookRLx0oXULKm7wFKduzNmmj4z7
XCd5If2MAPw0oajilloKPHhvJIBBC6kiBPJJox6o5DlQOQmmSqSaFuSFSe+VEsx8taRbzVDm0JbU
43BZL6cX8E5m4Ul7cI1KDIwT+4gmW2qKn5z1tPxMW1/hhQUzSp6f/n0GVnK13net1CORvUs9jyqm
uYdwMO553FyIjXdtR5Hb+nFk3nJHqCh6bE1U4CtvK0Lp5J7nrHiChsXkAZdwuPCy4GFKHP9Q/7Eu
nNNTlB0yOA2eOKC150czlO5zlXO/kkr2cS6nttBOr5HidcUDNmGwW9iOQQ1vL/Z8hk6NE9uwgGoL
JpwRdzcxuyebNPyJUaAQG4PoYMLsQzzLsZk2JusA8q7Bj+qi+hLTbDifOfF6WDgI7XhnNdrMNyc0
HEXTq6uUelC5uCr9L6imYM0obOETA01Ybss21lmiCtEzdDeEFdnFWptC+xQz2EHZJFOT3mYstmv5
6ifnCBVUj+R7CvBeAmVXhHS9j5yuQpX5PNKDY6Q56qVVjWTa19IR1BxvUpLJrbmDX0t2qZbSCS8i
MUHOO1ai809HahqJldUnspGaOu+6Mgcm9CM7bvfqQDyWrzE8a1F/FYnUX85IQMyUxUSDe/VZid8k
8aHZHdeJjre+73nAIhLQGytti2Fml6qiwlqh9a0tjwBYKi8HkzLteIqb4LqgMaL17qA70mI7zfb6
b9PgHc5mv7Ua63ylZLU+yp39X4VY0RLM4dUnyaeV+e04yDiIws7tLMBQE84LAyF+Xa8eavhS5ni7
Iy1ih97PIUNnxXWu15GB7hNDDnkJ38H8SqeOfxf2JJxjblqkJmECpKx/m3nIs5z7XmkP+gFqnfqj
XNXm6Dlp8prRcLIi6Ji7Nc2GWaS+5uy6MWMxuaxIINcpOtYIzXIWHAL1nFEYPdUp4Rrw14A+KWlY
uzTCyOioOVoi4jATRe0PcaR52tiz+f75vvCjlVzgqImMLSm2QEC8N/M6LGB9y3/zW4r4xMJ8CtrN
1UOVjoVuBQKpjL1QEnZ73iiw2PKHCsZIpBnEc/iQD3T92Pi5ZqLKgSY9fC1mTL7wPm5P9jb1qBv3
9C96/cvyLhcGEDNEwVZ+7Az4eKlA0SX3Gc1Luj6erKmzasRgIxwwOOAdhaDk9DQUjB83Gmn/npeB
ncGLz7nSi4HUTD+CedQrAoZlFKFqQx2zZKNisypT559hYrhbbpfVwCtHJwcwymhDcXfgLjaNYspc
RDwwFEytok8kVgXqd07LBrxvfSa86c0JoPh1qPp7WQYkOH5474DsBKx48ISD+R+SG5QN5Q1qeRRU
fid3g4pcIqjvhdf/txdfad9kRqKVc0yT3X3sPXirTmyiYpbesbOHP6DLCN1poipMUCUgPS6BxbIb
1727aefit18DTFQ0cH5eWDYncYGt0CMr2M7Jlr9p4nEZA6Sd3ji+9h/Q1EX/DulcK7e/0CxJTPEF
esed0b1/9eck8pk06YtRv2+KokZd9KA9uWsI+kLw5jcfo0q8lPOWR/IlUfDsl6Vj+4HdNlYN4uEL
t/OKpacpA1i0dwguHy2W/voPb34clabj4ylEbPzGjtTq5f1SIuiJrs3J7No7DDwn5K5TOd4rTUcS
ZEdG6VuhGrYhpkabuYZlObPn8yGX69be1J2MtIQyCpvLlCqdUD2eCY1cvCGb4gzz9uxi0Vj+hbxr
PQ0CdsnIB0oSJJUTNBoPsy7omJspcSmdoB/t+G94/vDzGt0YBFCGtv41f9TGRzSLbsT65WH6jDF4
SZQi09n3pqTs6D8OjLPoB+YDXD/9C6ODbBiYJVV8dJAY1TWbRty5AxNV4lIrq78CBogtWd7tMgOG
R46AZI3EyWKJYAQ2UQPZIml8exkZqg4XugYp187u4gGt5av6An8lzCVcHRiiOUW/omTdoaV/2t4i
f+LdBqjBi1gWAF/5vhf33KqdNIcgsEe0G0egFTclFGDIpbFbbNJ7FR1zuAU7g8qOwtaenr+GKR3K
zlDancOGLj1/8A5S9il0V5yLvOie07vGUu6ErfC2HPgsy+izGZVm124lGpSr4wMQmEVVlsvDsXRN
p5ik5sI/wMteWWldTGC7LHRzfsWDW0FTwCkznudsedLWc9kSaqKr+auOuze+tKF9kv2y976WwaxY
phhC9249q9BH1GaJhKS4RbNX3YWajn50oLJGi7s+x7QZchhb/Ou761hWLwaMWRojSV1A60OZKp4K
2JUMHPn0rQ3WILR/+j6GurkwESRYAYH/oYjnHnG3s6ckG8SqzxQPCUe1lfRqLemBYgWrWM/vFw0t
PEmlPJHRgkQSfwxGQCc91VTDBtJXd74xGbY/SIGsRVQCK2gHp2M/Mi8hq/QD6arWaxZbU8sBX9j2
en56NPujM6TUVLTx1DMfyrzysDgMDAGuUfKK6LH4yTy/sOfI/JAPG4cNGET9iijVPW8JKP7uQdms
vcOIy4rtnDUvCybWLyg/MSqGykFbYHgTiT5qxCnkxr6V6RcsIlYidwnlAmqH1cwI5QV1czmm9UFv
R2OE8Rsiupd6kwIedSzYA5edra9UAQbIR46RhXnFDa+3rgWyOOEu5Ca5Hw2OBBY/gYDY+/QiC9EE
ZTEieySzvtCyQ4hT0B53JmMMGkJ0XJahCM2MtRO1QWy1QwoK0+SYZavoA4sHMtM2lHW8BJ7MEUdd
cCovVH2iRe/vwxIKEFrwGLbjFfNFN6TS/ahTl0uoSGhi7b3PZk7EugVfv4vC4XbONsezfon7Kxxn
vueySoMBMI8KrpbdjQRMilOdupyS812+T512nIwCkUXid+0deyXBqvLVJPzeeUoZtsdU4s4ZC3QU
8iJP2DVEJH99Mni3XiZcIf7KnulrTSeXdlwdNGqyEcKcG2OUK55VB7Q/X/6XzVsO702/TwCJgbcZ
xsdmB6fVr6GTNieTS35BYWKKji85Oo0JAO82cgcBuuAnRNUWxFgpHpPCL2lhPCgUt2wsi84CYonm
KnpsMo3pnynPpYUSLedn3xZTvSkiEpV0P7KA+xcNgCdyT0sQCl1icek1G8vye7sD35FO8VXn8JoG
WFHuVk83ncSp1iE99jEG3GgYklg5XEigwqXQtUpXTWiSPy2zLUj6ouzTg2Cc/RKI2LKrmIHkRK24
aJEHROx6yAeG7NsYOvG/VvOTbos/vrDQnhTgVvc+iJtzVZOPXe9f8IS1sQfztPeQWxxO51N8rVHB
KKK2Yh0Gt0yOhF2vmJz7DYKxPz4fwV2+X4xnA9KkV4n/zxJLEpzMP+rDHLD6ATCKeRlg6F66yTTt
3I3kuBVgZwfu3rANj3c6J+NuAnlitCBH77GQ2xzFYgSNPBmI2S96jcOWZQv35LZyikxZUagCa0ko
8wMLIcgBxlvjV8eXnsX/ApH4Nff/ikjZ1Jr7mgWSso+S/HDJuZowgLiKeJmGp/Ki8BNQ5PppvhMA
OWgkwFYJkZC/zyI7745ZkaV1SD2NJXv9CrB9xZFopLWRuXHASiKGR1QuPlKNwhk4SVojcSdxainy
OE4UJcoaOaj2wBFv3OFUewhlmjVuuGbY5fBy35BqssPeuTuqBbmdkIy0X35a+mrtK0H6XQg4FDMv
vKYIh9ZQdG0PFOhIfUgJ6wL+0pq+reRC1Xw0HNAC3un+bPGZoEGtO59rSZUSf/aMPFJsZ63OL30t
Q9AdmKM9XLji7/XkThitvLT035YaUGmoPzYmqE6XUciilmFcSlFM/xSegebYvtOQ4ozROqvWpb/A
UauMkoMNyewwNni/rETxvoZjbq3f4Crso312a9BOohR3W1FH//sBQdfjJpGyCehgZfMOfePYjf47
vNr6D/mRIIN1b7GgjJeuHFru1Zg3ku18sFL215Ojs7tHVzHEU5ovYmlX+ljRNqlrEoupJM9UYuQk
Yte0yWPyjl0ic/rnXJcSCxFYhfm7pY9Lml8JX7OWT5M4oJt3o0vIa8zYEefWB5qlU1VtvsvP000t
8Tu8AyahyL4KDtSwZ5rk3my2RLfBUNEjMaTkTIDqS7tD825ig7Mei/h/4ApMFUb4ymx3nA5zbeHO
8pBpEH1GY9r2PwUEbSQuZ9WV//bwtsl0OBliJb6sdLorG6Rb/4IW73EKOgvDif+wnYzeffsDwfP9
Jszstbe8DoHgIQkue6a/8XB27D7O+pQKqt/qo8XdYLDJwBYM3UPeGDOtAnixAj74Me68UZNu3tRx
PLisSq6NqZ0u+aAKZW4sFyKGwx+8cUsUt70H4G8urtJVHv987WKD8n1U5f711LZ/C+T6jQijX+H/
3s+01nNhTYIgOJblf8hontJQljxLCZUshttp2DtHAYTwooT2JzJNBrR3LnERTwO4t5EWhYI06tOS
b05OsksetFIvVzwmKT1EUhoe/787BfJzzsQkJBw7jypwaMw52qb1L040OqzS1KSRfFNgO2tOyStA
5sNq2zA9gevIK2DYOfoUafGgR0y4pz1+S3+dwn4EX3SCTEcsSV6iQM+HjpRb9U+lqsugaykC0b3a
p6dSrY41VJpYFxsXrRGng6GdxmVTYvWe8cCdRz8TEm5cFtvGaxXw5g1A8rMPBBm8G6ZZ2zSI8RsU
JIH5X9k4Bgv4fi7hPOxjs+ak71U5+gpc9uKfHLHM2XEW45dTXCOxcPyumUYhcTxTvEXCQ8KJ+hoI
+pnsHzx5/9+GeZnKTedTzobzXcgqLXBzWDkuP2gzNZ1adf5pofCUOcSJNVT0BWX4K6xEdk7kh7dH
8IQUYxe8J2CKd6dmebYkUxn4YQVJif7J5AoCxg+rMkWNsU0OSTvzarZRecj/uin5y4wtjIMQVRkr
m7psRGgC9PJZOwpfDF9DKpZ9/MNz+oxEWjGcMlFm1Q5gLEZ8XtPWjrXnzLSFn+Vj/5ucYNefFON0
MYG5CX7duhiC8ik+oIgIN2fFPakBFQFGJm2X0t80RThcXb5TjL92u+k6Aje36gnSHSsRva/qNd+M
wyv+zFNDQvXKfu9siep2Ydy0rjsxvh+KcrUSWNQWn7UzeyKS6LDTDGQ+miVtsGOGCaQOUd9ejdwU
AdqJQZYYBZ9FMvQKEkfKyxN5twJe4dxsItlPecZRejpX6tE1pg+9w7Xv3W0nAYjuDF/vsNxFqfgw
BjS/kOHpZPSHZaIO2FszF5i/PN18iS9nbWIR/gbcX5qggcivzaiDLssAPexZR/Ce4ELd/vTlI680
sKMue4UzuUdN8R6RPXNO0Ejk0Mxg/bdsz3TeV+JS8CgH18V6I8U2sBJ62orgpqOB5gUr4yClnlDC
rUozwZbIZ10BTRrnL8gM7nVejtQlEfMRJvKDPNXux+BAYswRcMVHt4IU5qLxY+heK0Z7Na89j+u2
vdMHO++nV3VRjcsElNdLf1jxZc1P73WGoWHpNEisIgxvTSGamdsxA2YUGKftFVYD11UX5hVEXdHG
S/FDS/4TL9VaJVXggDCypO+a2JSROwIAnyZN8hQ1DTBgYPs3zL7fF40pMk+DvKq61EZmur0n6mbA
YUeVVyFt145IHGX1pgvfgLHcJk2GV1syFEohwLG1Fi9vP20iHPsrs8PP4rsY8XRqFVSK1o3xSTQO
C+4Ri1Pamrc3tiS/FP7Te8Yk4vlAB5rVpg4qaC2lMqPM6OpKJdgOAZx2lCrLtbt9/fAnSUZwBMfN
8S7rlWjobIkBlpaTlq9xDmcAf7tKgrexFG/sQVz1OPFuptAxqHWhb2JNr4wMz8CfG7wdJ2EPH4xl
zB0GiDg0idOYGGKdwlSpuI4Oxlq4MUBbdB/mYnIqa8hxSQYUmrHeq5iTlZHJwqu5eemT4IHuZ0o+
H/hEZX1H03FRhR3z8lQSWuI/UTNN6zf/f9xMXn6xaxz4jBk5u7Xbru12WHXYieI1M1FKRihzqZYL
faTL2h0qhqC8PW4apLUixSmD12vKT25KJFV+X4c4RwjzAUv48dqI+N+dwqLupOMZ1itq/6vBo0fa
lqebP325KYMfRA2Yhslyj3n7K60JvzsPKb/7IKbNngqBX/VUR14XcCKHAMc/knPqXJxuE3R7ma5r
SuQfdD6qQZ78FEYxprAw4iUmEmVw21KFeK/ch6KwysKMDdMOhVUzfR46DsdwLn7oCGu74uybPKe8
ZNZfxellxtArfTNxADCI70uZOcEwuh2wUUrArPUy1JGzsKe3Qafysu3sBu5pb8RMOmXqOTFBOHA8
gDB2yuz9TdBQU2Qxiw+CDtdzh6nEc8xRrw5DP686M2CL54FzpEs3OvEZsorND9eVBQFuyd050LY/
1iInuwF3bx+EaX0fPla9dfWZjq6musSarG0OVRbmue1aSmvrGgkrreoWbLL3kIQiL702wRmesytn
alqZLb40kDWoqzzG4BcNKFg0sKJXyKMakbC91d1/t5bvTWj07c36RL6/HbfL43yclHC9miP2IYbt
/xwUMLXYIB8LrBXR4Ale8hOo0aPk/yx7Xy1f1qjsCCqV/yCJFHcGfmGlUkdvIwm+fSfH9EE7Ki5v
i7XXDTMLl3hpJI0tQNeQ3c1B5ZwiUIyhCeHsgjsMKKc+UsK8J++MP4MOi3athS4P3J4wL6LcdmF1
ao5meSbaTHKohyMomsVlyGH1z0XOrcxXUcTnsFAdiuXDSNhBI3a2aJUlejSZ/5OVE5iYya8s6aST
a3MtKpFDO4w69JNHWFsNsuhnM8ipSmPssOK7Azur6djQkeZEcCQY7QLDv5Qd0ZMO8+3g6AMNCPp6
oK8YtdLSUzVc7asHNFRd5bUupo3erOB3c1iULSzDfZcS6QssvL6nz2TVuYcGiy9s5n5Dmi3sJH/U
0XJQ0VRLmbNVT0rdBG3N3GrWU0gs9S2Td5iO9NJxLbwdb+ooFMLy6NhfdeIwVz+7EXJ2OpiYj9VH
Liq3m7Xy9Qa0zSMEwjqQEQzShfllu5U15e819lmy7JIuyLNKKsZ3802vFVX7kdIJL7VQT6P5x25p
NpAr9BM1IE23ilUDrGrjmjf26v0h5P9zqKNRNJHf/F0Tp8ieCnDJMqEZY8VyHyHgV4PZal7sK81l
mcFJtjjao+WD9bAw4K+iicVc/lcYrnOUgOdGzNdvbHjkh7jX/f02E1TMy8Pbq/5viHZIdof0Kwm0
fvAGUwCU/Pq5zD+H7eJkJI8Nven6kSLsByA0AQmPbGEH+qunSp97iIpZG/7NzTnLZSn5JUfA0BNf
RKSmkbk8B6KsW32Ibm+l1/9w/28DP/dKuJWto2bwysa0h/4hYvB/9b9uu59OB43YuAw+olWJnVhV
gUH62UFof27q18QH6rRjPhUoKlImQQSqtoztcs0MJvY+kVwdIhmDp8y2Oj4RBol/oY9r6/LFSYiu
pysBKbsD8YSz1x1RHIIuBvAuw4+gRdWMYcP+cPz4p2YGy61Nft/uCTKtH9BXajcXY5opvTXppKi1
oXHN44CtThb8caibHMeRxLpIjb/ytV7FgAWqoClFvRb85O6VAxAn98zxCGHI3esbSCbqal/zA+dT
MuNbnjiTXU6ML77lVfT6cpoUIuag3s9C4liF3lFemVrunGP9Ccd6OHzbV4N9TEB+B90TDnXCtZIl
0yGgXz4y18NAB1qTEqEOcRUE7WdJUsD+teyRY98GcPWKdjN405Ru3/ejpjrNnw0VvnurWD4t4+Ne
4teklEhGcN6RCtbczKndeH8J7Z/QNO/wo6kHAPQTqDQij/2XVe5F/i4MwjuyaKoyByQ30TYbIA1o
ELP5jO90+b8bZd1PuEd/QHJttTc3d/Oura52/8uyThy+QFqvIth09pxiegKUlN4gciks+Dx68ts2
F47zBED7ZeKAz2X0a1hEn4hVLop2ve+xuUk36+VakdNux63tia+JHlP4zhxlWV7H6+PBNiN6K+Vo
ZjRUxakE4CVr4/ztM1KChTc5kg3J+jxlpwvaSlvwX5bu7nMhvKGsYzBohOi3Y3xcGZimOOszLMl4
riSCwqPHuLzVl3CDhe1m6ZaQ2RCDU6OBnjKfolBHZbY8uHlJ74dmVeTVI8xLd2akKiHJBrjydWLq
RQDRMTfcBRjc/7P/dv25cw3dMqsq7MYa2at39LU6SsggNyQfHTVZm/EtUKLP0N/Drn4P3R2uXnm9
BMFHxMF0h4wU8z6hPjH9T3AdUS/mCQa4OEUGt7kegAPw4TCqguNCzU8cm7pCOwaF2/F72B0aSXEM
YUsfuzLa9V2LgZ/IwTJ/a3invNsiKBXus4Hkqm6Ie2aOjCKREBRLRR4jpLSaw0f1fX42eXW+ML/O
LIfRTUip0tI1MP1NPQS965fKA/imsLXnC9S29mVwbIOYNkQ9xF4Hto0Nzu8Be0dFZpm2jcKAS2fZ
f1pGR++kw7uIBID/UuT7Y28nf4MEBylTyINd5VN76fLy5he8AVqXbgRha70+2Z46N7sE3bw4+K2j
6rxM/9TuobJ8ahyHrQxIcL6DlA54V823ot+UEBvoN5KAxoxbn+PNpMgNbQONjzb/8LgzVzXVfxwG
cUecCym5/kjlg+mnzd5Kb84LJjsOMUWaHmI1klOr19sFpTZZqvEKzSR4NQVueq6iJPE+eAwimsWC
SClvCiCjmqt1UBTjV39oS7OTFTo9BQnak/MZSxmfHufQg2HLsJGs6Fk5rShH6I387PscjrdYbEi/
xw4hiy62X9BVKxhv2kZsfgkxWS4Y10tdLaoGNr3wky7lrAAhJB0OxlsmzjwWXBy6SORWrEsPY2Os
SPOKLprADik0E+HKvg/zPaHFSRejOfiVVywMP/8OYTn7O8vWXtgBWjczzL0H89mLgzlnLgM5Kf+W
ConPDBQKVi1iFsn17RKKDSoJaVXT9c2tFj7Rmt010vTlbphEmRKLClV2Ttt7yaQUZjpgwX6dp70T
odW8D/GotsLsTUNMBIn9U+I1PbA2xtpY/a7uqaWJhaak+0dQVtU5mGcdEgO/uud2wvEikR26F8wk
IzVSudHahXq1anuuvg+A7T9VrR12yTpXClTo+rWmS5VzBavir+a8uvf0feed0JQw2n1S3m6Ekkyy
VQ8C+zNi2B0/yQH1z5B7AlGj6M02j07GrtcznNGnNHM7SYBhQwFWhGkhwWVseLjJIO9h+lGHefcz
g/kgSEzeiocNVp6waPEfXeCfc76oMf2FcQSPIlcafhCzg7ROCaFDn9fLHfuL20mAxLF/93MzX4z9
iuIYh7goLMY2IgHKQ0UbqIiG/+trHC+NTFdyK/WgaMSrD0xKwxROrHW/UHVE/dM0GBCIii+qiS0Q
H58936vRPBVHBZijp5J6rvWHsZ5Y6YrLvZEhk5FxcLpd5QsQVtK882gWVpuECHHlMJ74hR9KuXYF
FVgAiJX5k4xyH52yh4DtqjKDfqFp5HSXYrjt1HCeVY1sPP4WhEDfm9DO7T7+72pTyja0vZuzo36O
F/XbMKocJ/EpFJ9+emy8a3/Tww4XyfObb+ewCYDQMWMcVsF3rv2rjya67ohrd13uUGSMjVjp/QPW
P6tlkFjoRtfuhxMYRg0VdMCCx/GTvvVgM+uhKTf7yODC1x67mLCggO9gCwrWPlHNDl1wio4jTyRY
ksb5P0ftnf80BMSMp1ivYRKh0ovsrXmLOt65DSqGNvsvyAMsqXdlPI5xK/rbPPA2WM/JDIW7iaEp
0+WzRf0Tsx2iKA0UwMWc5WTcSH/Fx4yRitW5Uw6Siw8uTQwEX5F7L9tjDI8VxOAXGz6WiZ1eUWvw
HAJGfGOGM5xFNfTBszpbqqVCcUmi94V4frUGeww2QbrSqZHF0RxMYFQDHGSXogRX/rDAEf+kLbVv
PZ+hkyckz8AuZPuQZRMjZVoQJ5NyGZ4AUpW6QxTvUKR04wWAXZewvKqUrNPsEAQgsfeW6jK7Nyz3
BKnpgh/Owp0UStpLa9ZnO7sx7Dqi+t7DNMyeKSNwdmyG1XsjK03F7175EpUzCY+Tc+++oY91kPRk
1YCnfU7o1wEDZSh/HQiZdsX9nBa2g3K5pc4c2WynynXcupnSt/sj/eoblh+9sE1VUEJmqcHrslt8
IleaAcD40aAx2TDUNAT3Gh6yr3L/arAiYzsdUBuU74a4A5tfpUaTsrbBAvPaMhEn4K14/zpj1Gj+
a/LzF8efASs8S1qyqaxJA6kGUkX2dRubjxfWzZvCBXL6/gdoHWp/Y6r8pA4a+Tb65FKkpC8oknkl
eILQ6GibpaP3vosxL88Vqmb90mHMDgmhUySuU4/vbYfjgbju3EcwfX6o6bOQEdBX2w1pv3Or30Ec
A9eG+pJMqXMEyyUVKXrRJTFzjER4HJfglMiAGITQgqhcFa218SiCMudMw7w/txmGziCGnJUFPxkw
7wto59K740KwmEfz25mCy3s2ybk8gxoq4HllVmUQpwesyRL5+tC+54La/QZjcU06+Gl9IIbrJjeO
5j/Ern01E1SpU00vj1lSD7dtXZ6xV2uTIeAfTEXxHxbWMMwLWHE0De/eANQ2EgJdyfo/V9K/3OpY
pBBgPZnY1iFfjBcnRPbyU/2Yh64sARrCAcWT9yKkgsIIjVGRuO4WGhSSNr9FbCV3BMqy3+NIRaix
pyojf0/oXlT+ipLHm1e4Wo9WS8//Ci/naz2/RjtVAwvsshEGc11UpnHcjVmv2G0M/rjYNnRrVKne
6xDIn7vgfmjMlfU5utLtkSVmYHVLlKITls7ulNsGV3evXDxccFSlFXgvpdjggdxFkrtyEvShr/Ac
NsizgQ/T2xi8GRdFwpVCtzhpw9JmNCk0ffp3SFWZU0JVPf8GNgh0LoDAdmkOVHVwybM93AvS0UiI
w5wuHza9AvINvgcXSYuhqy3KytIlnhFbOfr6UwpWH7MPk3mm9AACh/lg8+P5MD1/mA7bHnBGfc3o
vDiJhMQ8kBKFOF5jeoLpt/7ftKNGRt2v4yYux4bxLak6UokPUSr6CmWW5FDp7f7CGf9Jcv+x1yU4
szSUwVXfilb4LjWFX6w1pqOxDnCSf+6Ma03h4QsQFivQM8XHTcfUiMZ1Xh0hKoAIXV1aoVBN9HG8
j8d290M99v/1/ruXx1x9oALqQv/sJlv8jJISmcuPJiu5JxFEtuRgjOO71YZ7DzBjye2vtgtAJZSB
GHyFT9q4ccgHZSBJlXjIULW2fiDTNCV4998ft9qb73936DljbO8K+O4CpFB1XQCxrbaTZioq9uvL
YCbi2aq9pCFGTEFOxYX9Edkm0/LrLdVUZQTJ2WTjRxjKIcoGP5/v1Pvigqxp9MpQDuielNqH29Kr
AlTS9cYEIcNieGDVfBsvo2lf42ZTI9NXf/umWUsZLitAKba543bo57ZiEtRiy1Z9BrWPE/k833M6
PvFJhAUXSEQ5zgjz2W32TiqNUVXD/XpLoLik1/Oe1Ui2Q6sajNcQH5Dp76VkfbDmQ4hpS6R2nQcY
wvqICiFfhKc3z8xOWufVARafvmu3u3Hc5huCsrbCQeQxEg4JI+wemhE25b8gKIG9VBsPDAoOuW4u
qgRs5UvK60uRHUCp+ieeFkVADsxjgE3UmdXmpwnPIl83b27DAId6dGXrtk6fjhR4igzGbtMWE+ED
AwpfjWazhasf/9QFWxYP1fZWaOubsAz/cKfqaibRer5Os0d6qvKRQoo5bJJfE5BLMflXG1dRZB6B
iUrFiPaKIe7EKZdOXxPjg/u7Yik50xw+BTry2G0vL9+QTXWXG92O3DgQ85Awunt+DWBhRByXP+lA
DQ4R2TPv71Zd8mDWVMUzZ9XmSN1zkR0xA9h5Fka9KmarWkU7YqaTvkJT1PovgzaDBRdantiB+NnS
abaV/JoXUgdPMJeIEySoWHRtgmdxN6awvn5Zde9wvI/lzIiayqebNUoWng8nxJO26uzMJ2+waTo2
bzkT/zaNJWKvxoHTMoceYqTBzb+DYcL2juoLBhxy9vcRUX2iRohtoLUzu1iW6rOlXS6sXiKRWfXt
B9x7iBDKehDPM1ZzJpDDzxPKkuf9GeWpBDMz3GwwlGAitt2rx3Gy+StCP8qmqaHNIlQIXB7rn71/
HDkKFvrUyTbXu4CuqHB6Z52DX2X67o7plpZaO2BWQ669oJwTmy0OUzix+2zHMoR9WYTuK0sn2wtP
hJYuJfdLmKQjBn0cFwT4Bksq33N0ZKjReOUTiMKCt05qStdS6/rC1QaXBa2qgRJ55UGbY9PaZ58/
CzJguIPDzR1y2zues6wCs3NxaFfRgUHLe34MYGSE0rrdOZtAeyD1RHIBXQOMuYoWc2y/vBvpQiKm
wdXmP3w9RJqRLZG/4yVrQ1ZPl93s1XJqEsGb+2cB/7Ufh0UGZ8aAUIWCBgFdaSr7ruHwX5LrHH+Y
tydUzDXXbuud649UFRkzV1RxJjnrnrBrjELEDBKDpuwabTKcJf1N/SMm2KsItHC+/TbNdvmGkzl7
7dHedsbsfkUzkZi4UpXYSo+7RXzCYA73G36mpiaw2/nWC2fxGoQziPW+KcavbM14oB6HfUQtj7xb
LGAFby7+fVsgjuogrbzr5d7ur+zJz/pX4gAGqjIDsS7AzdmVBmTLfnpXgovPwdkEC+07BCe3dqAd
NCBi3CwPpj898ne8vldaWb1i4sX/3FcVVPpd+kUDRjgLSHHuFHWANCVz1dzeyODJoLit3i3SJTs3
YYLfdlzQtBq5AQouATbDr1o8vkZEscf5DBwBM/0urlRPrt9ZaC6bRoLtTZS97MiJRWfpkin7OpVS
eBxIRW50vOgG3w+8zXLcPrKjplCztEmATkLCQkaKfjJQD3Zjg8ryW8ET5r3mTbJltVNnqpQ5xbac
7nvemYqHLc8ajboChonbdCid4/zpsq+/bGOm2AqHY7MkOSubN9M7j0Klc0QJ4dJRAJMu6oUl92uG
7ZHtoGQe2dWp7WMRe7XjCFGi3FhEJhZ9XgCuCrvXT1ikqfkydERYRAeF769S2bF3TB3CLID7IFfx
PfWu76Stmww+eCge/2j55Rx27bRG26JZ4tY593/2Pw/U71fljaEaUdNgEwhxBRGIUN/8rNLMqY6M
qg7SoOaYMeefbJo57ZwSEpZBdGcBy2Dk95zwkFoaqiLDWY1TzI3JTssjH8rXC+wky5a/Yu7mf233
dvqXfxEp9HKD1B38BJS2cFwA0tZnbPtXaPbZa5Re5Fe9uAifrMwT4RJMAzgnCI6dAoz5H492cX1I
woH7AEDXUVi65oR3fRNfuAKQ+9GfDYaGM8rnddip75h7pBPOPrAX8ph97NlYu8CeI+XCebITnYEB
teiz4gp0+XIBCpRgaqTSI07pwR8vgwciUFK7SIY7eGJzReHpj1D9oIkN6Bk9Jz91vkgIjdM2gC4l
2B3zvxYf8uYQ1ZgkzIFhIz6VFI5St6W6Y6dFUPIPBtR0L0wjqorCEc+PYVgj4T+wHBkKsELcJ9M2
hz62tjZxdlaDxreQjVZISSTvvNDqm1cjtHEh4746Jk/4U0ooK2h2Dts57oROpMBsLQsGP5CWMSd/
v4KlIpDW5k7WFvexZlyZovTpPZl3/Yrtk/3yJMkQNRfduxsOEsuvaqL8oxw8p8Hl9qY5Jn90zfI8
6VABff7jNUqY+rCTBZ1SFNsUJ8ibIAa1P8boSRK9JUrpDDe4v2ZpNTgfOfDuC4XlNhiHb3IDmRK4
oMSWihmIvdUIxZ22dQIPnhaHbsh2q9s+P7gaAPD6b3ndTsIMwp/K8vktl56JBXMwDWw/IzxwdUy2
lJdFd76bG64pcKXrJfcBkPdPhAwiaMZUrT7+WIDI/UDmZeRulkQmKAauOQNMY4VXBBwynkAc/4KG
Ulvf4LmSFUSJtCKy+fujVOK9TC/z+3pW7t3VsTJR9KHmmd2lBvQS601cU/KKX2ojG2xkeHQpqtcA
3szyPXda55e2OQ8i+8MvivdJk08W/yp2/rq1YQonvXNGmab3NoX1Wfnd+i/TFDqhABecI2CQYSqQ
Ap+JtmAsE2XV5FeOvTkQPsS0NtSe1XJQceVYkKkWKgGRb2TkQZPF1NwigGTHyVEdgU0iF+jd9b9I
xzQHn2k/VEP66kyv1memR++GWAnaJbTW7T4RDruU3Cm9a++Lq2uHouSw17MZMg06JZb6gh72bzEt
WCNbRhPQlDBoMIGgPMkfamvNRB9nytjNX9/xQHfpagvv/SU5jWT6X9J1djhAEmlB8cFsuoBu+gGS
gW1MkClm5UkkO4v9J8qWpRzi3tTkneTjWo0JdWsVI2Smr2VbZYf7DkVQGtfcpvzv5JB4SIrZDl2h
KmO2jIv6ELoUC46rf9aU9owkbACoxr/hGIWG1utFjOpFFEfozgAtq/OKv9IcH3/oW8thb9CDru8O
8LnOtbeYEwh7jpR6WYKE7ccnd1EBdWQP+N6a4J1dbCmdD3zj3N3EDQnxjxtA0OTmjiFum8lCKkOK
N5k8RpaiOybf30Gvl678+nl3yXdOxSWn7eC3ZYFhNXEJfxEFiaTxzn0TeiLyWAHpO47lRt+dJtOy
PTj8WisbHBwFL+UqwA8zrsWJGIbfinxvz03Bk3hy8NA8oCFAthxG5Ye4WdAb7cLJ4Esp2UcAHzJx
xyaA8OKBb6WWZtNa3ssGv/776Rvf8u4nQ+ma6U+scnNFmHimOjO2zufVRsp4dX1MBUiaVDoeOwG6
WfCIz3CxKr4jRB9iB2LPVKjfeoWoPNN+Vd5DD54sERU7O3aTmmGwvEDNirg4coOJC1/FFlHjsG11
BW18izGW67JmORtEFfNtD0EZQOTgAXDgIU3osGQn9RHSuacEfJaVOIqaATfoMj/cUf/BygCrbipX
HWUlpVIz0njDXUHkiSMXWjjyVX/lgcj8soOmDGR1jmn0T50et6ompBOJcy4SosR9+ajJN0BLPZzM
nyQXLRyKwyt9XcjW5gJ2KezLqhkF64nvNPCf+34FM8n8O6SfAjT0gMoe5DCxHiKChxQuQ8T+NlJt
CAkj8Z2ggEZZuGU4Rt5Yw6PN/LcMfULds4WxJXH/KgSsr9WuQylnqvmkRqVZ3nKet+/mHvChhrxI
pioOXJMAIDT5iLjXninasthnGjl2NCYAVrcXZGGhqvtkGQ3zp7X/V49RO09KMGxoymWeAN1e8ZnH
Je71FtTbgqmpk0Gog947eXuc2I15EWNBtU4xqzl+c0Cs9WXcTYyA7Ss7mf/mIHcQ681IfWZXIXRr
4xiwWx4R3ItVwVCLppTz5hReFaQ1WvFxD5NIFssmYOI8qqcNiXbRdAde5Gfdv58nuJ/sVGxBuQiq
fN6jy4+/s6tcrFL8URxOagWdlV0lFLSXvXjp5NFTv1mvypywXbEM9sDPjixyxhDvzxwbklvHAa5u
A0kyX+AqXInO0+F4Xw8irWALurvUgZTXe9pCKHWjFecNyZ5bMVeC+a0RP0FPP0RRrNIVxYx+s1Ey
DV0HlXAvz4xLLBPiYJd5DIHBiHNGG6tafIRqkipK6VJGSZq8z3m+2VMZp8rdpFIAo8P2oBIYlGeO
ivFq1j/1HDME2hyKCN4d85ElXPXwWI7rzPd1LF5hR2HJ+y4L5uAoU0g9WL9q1Y+CY3YvjZrnIU1s
ZGTtg34fRCknjAxeYHpM1MEWOGX1yKzys6d6LckRIShUVOC7Qj0ymlAFdJaDZKLiHdO9YVtPGrLZ
qPci6rKXbgvzLiaW7rAwKUO7/pDCnt/OvFgk8S3T5mjy7GJ0isby5GIRQSs55Y+ieCRPzJ8ee2G9
YUUeYwlPFHRTitW7Me4GZfbpYhnrszbl678paxVJpJPHICCCgOxYm9uhwpLyyHQ2i3miIbrqH56e
dLd0/B7iIVMR9wJnPXls+ilfW9BDqJ404ZsqkJlk0kcX16Vu/HYcP5AOCa65cHqkGdxhADGpzKPV
SQP+x20UbBpdlObhlaj/tVTC4dE7G60zqTsCPDnyG4+r01mrT2qmOVENbDOAPh4ybfleYCSB7idn
ZcxFM75WAcSlvI4ccepT1adVgtNYWhzrEFwN3wDhs2u07G6PoJurulcLXjBAu4fAwODBvoUfm0wg
FqMap8DLaiOJfkmfBbSO4r+eq/+KhyNpjdjAunPSQRZ58pFZrs7kIdn1UeYWCvrdYTI0X6nfluGV
0eXLpBoBYuvNEqF3sabiJIPCW0k6dJ2qzIcFoczwoRoLLenPT3uo9zC8Vzlzww/Y7djCcNKXGN3k
Ks8sqE9ZeE0CPe1485z7aYX3m8CQk5LjZVIiwFMYfWMaEpzNVeJuIDIpN7kGrGTinmUSuTDrcHfj
UyQpScnFT+dJAx5rrnP3sIuSmnJ15wBnqgKIwTcH7zQxKKuFP/eURFlEoMKx6jB2u/003QqKs/4l
EHfpMzmf26dfXazNPsJEQ9wLPE1eFuf8Co9JMyt5ETNvwsZZER/6rp+KajXF2Er8zM0HnetMvZe+
aW98nZxJtVm5zu6WtwjLLbmo1QoL16KN1A02ZFGgctZ4vTyJzWGW10/toBrJj6n7fN+WnT4QDiTG
3ZBo+rVsWoJ/nGqvUcFjXJX7ITLdfDwXpyVyajSwLc3XJCDPtha/Dh82HTVDWAGA5k91V5EJIuKJ
A6hag4p0mtTOz3dAWppm7am9wQxI8252qrPzpQYH8LzONWG4LHZc7VAgIEIPSdg9ORHmrXEwOpJN
yJDLeIgk8slfXUZ09fO5zZ2xH0Qj1tP/a07iXHIjeZt469Ag/hVLytUGwvMtA6/os7ewTTgrutVG
TLXB+4Uzk4bSeLmqxbqVsXyJhIhBqo+rh+bFUfwHtMXRbV0WBu39NBs3iVj930gU8je78bvmHovX
GFojQQoB2NWmIrlCLxl989qSs2mvEqGY5iuDqG5pd/Dzxbv8eW7djIzNT3I6h9ixqTSTvkGHId9u
sGXBtmEAMM2gXC2C2Pfb73ml870u/Plxddqsze8xuHpTqoYf/cyXXrCh0a91zVGduBPTibJNqPXR
fse+hVMUw1Lupt//7vBI4wIq7rTfEYgp8etfGoA05wO+LEEW7SEPt/6h+qWFomXsap8ecZQzX5Ea
zYfinZ4Z/3uoVowaAdsuDkexVK59ghYxd6i2vIBCUEDU2JD12Ybc1wXbZqwyVTNru6PqaMuTwUjm
hJNO12IRXa3YJKYdqBRltpEUV1n6LJBC6Wp5+bEx/KKPov+f3N89oZSRUg+Dn9u7NJGc/FgHKPMX
hIfj0eJ7aXA24G6RBIv4TlfYRdavarkKtlXWgAK7QiAb15ZZC1fTGYu1JX7AZB87jyGyDLKhTbvp
Axh74DXpFnQQUVb0OZzsNu8POb1DzkSP9BFLFmQZjz33wzdRCNpJHZo0+bAJhhtKbWLCChhHVR8M
YEJ9/+dfa1XUJ0ltWz9e52NdeHcLO0oJxy87RNFmv8fzyjpvMOXACGNFw1/ON1EiEWmXbDBt0L89
5kp04RHAoOlYLFqlh5ZQRrtt5VxAU4oYDckpGW0I3aA8+QUhQr3lhuO/4hwBbQ1MlmwygpZYlgzj
vRn5pjHXXWK2TFmiG8bqxEVPxKaJWF05l/6XoBT6ZIRo7F7VqKG+vPwkk5El1CziOjSLUx+S/jKi
0KXkbcdtUQ+3slvPt5JvvVPmBaMxktHNZte/+YCPq6W7U/ZyfgMzSn96BwHvwCkuE+LfESZfjBj4
/uMY+ByHI+oYnGBJ8tl47Xwkq/MkBG77tRekZRTNaF11NkNIEPdEqVE85v7xa20vp4aNGudlpEOX
YVU84vAN34BBY1c0HIVtvQb1jCUMKFmAYQPRnmI2er9flcfZiOVHd492kCF9LT7lfSW/cB+MkSOd
vi3+ZEx42c8vV9t7eUnyGKHjPnLDqzbVtJTXq1ppFZN/gLvN3cYqoeCSHJLJlevZFqhMiBOgc6QV
VVBeyorblz27EEPXTTVZJzZytdky5JoZTj5QdPHy6sDMYsYEgum7+H9oLH3Dg+f+WVoWWQDFKrqh
CTQQY0jVhuKk5M7qwAz832Jc9jeb0CKf/p1G6R2yqm+EIiqTcsfwxWWl0NBng/OmyyOXyVVQ9TT+
3Q4fSDKliDAoET+Iy6UzCLFNRfp4XrYSF/h2liaUA6464Noc9o2+qG3de6YvyWUpSMWvCZ5h33fm
06yJ27tmRgMSek5S/Avq06qnJjSqTkb0I0ljaHYJZ0FTSq93URso3rB/aNEKLgsJg/l/nqa91oxd
JDldizrTqxSQd2CuCfDYJs8kcT1/x1aiz2zkZNi6iFRcycWuLQXBa2E52Qiyy0bzZLEo/2mxz/ia
BtOlQpZ6MS2SyWFVEiChmlX19ZSnPSrSsXazkYp4wA5s6FkO8Y00IB7oXY9Dxmp9LpMUobiUzxoi
eLZARAOOEwiMYJdxKkjCJJztwQ/pe9tShH/ImNBJWYj88eb/qRaXm9yn/oPo++eul7Nlj3F3mF9G
3voYOMA/1wIo+v85FWjrAANdrAGG1VIGhUzywTuuCBo51R+YAsMlROxsfkAk0uST0mGY4AMSMRHI
BViYhERSXKxUOAaUljL2a8+sSdkdmZQTQ29Yc74E9gehttJ2KOAfGo6rXHH7hdtXPv3CgBx0nhYQ
A3JY4R99yWzaI/kKt1BSsUryJEMK/33zDq0jvbKwQVB9H4aIy7fFmOaCtXnYykUDR4JRE7JHSKAm
b39zIUGBJfJIWxOMBTuHZABJn/DxJkLcH2zQDPK+bquCCvw7wlpc5rFrn+5BFzeFTZmXfd8jrc/X
/jUvjqv1w9Lc/DJw683N+dRFKki6sgLtpgohYnW6jv8sE2eUIFG4BYWHl1WrsJkKJIMQccjPf/Tf
oBonuDc/AgBXVrmmGdJKWpGAFCVgoawUfdiRlRZ+Y/6rOpElQ2dnCvYRvrwA943vwiIARRhT75Fk
bUZfT1UCsNEapLw9iHlJyuX2TchKdazVjgB5WgYGDHQrfYK5tfu0+bUfs8gdDT7Dd6BDMAVVD+a5
J9djxoXKFKn2odG5a6hD2r4B1btjkSKPgL6kJid54yLdCAD/y2MK2BoUipMAnCt238XAv/3eMvTM
yJZuvUTjSUR4tNoKd0+qRp+jvenIyAVTcEFwSoaOYtroS5mZ7y+qDha+V3rjFzrBAZaKHOV4WV6/
Uvrh5pgS8SUL/CBFn4oR32qKOawPrS3SU/6WRHz6S18gN/iH+f1pFSBmq3kX2ZXoqpSGT9FZu8ea
d+XGvW0C5PrVGQB79fc3ya+rnDbVWM6l6l2VE9phKkmB5a3pSLo5dqKAnrAphDESECd2Z/UWdfQ/
k/wBWxDfK9i6HEr4tYH80NrdlG4hKCycofFrl0SecczbZSZ/f2xiRAOkrgCqbAjjb6TrNXrUodlZ
8A+zoFlRm64HY3l0fievmnqxsMG0YPVTsn/zI0TZGxrslXsGjqRb3aRrXHHsd5DwYomObIdnQHrS
8BmV4c4y+6eE9KmXkgdEsFd3tuWa6wySt3LuCIPjM9SEm9vv3OK14blsStZztM9a1/VMEnc4e9oE
tF3bbeNZw65i6c0SaMb3StNEG0K6JBcz+6OFVqpS+BtMY4d6zDeVsZ1urKCBfYuc3LfJWpEKFtla
2XmYtm8DfNGlXNt+z9tOlsAXFTQ1l7ZKrutI8pr4J+W5i3CghCVmc4KGCGnhdONYdoTljUroZ+go
iSezFKv9rcSP1rcE9unHVNqxAWIAdW0socNF2xQLPd6qpMIIZ3mFwhQCh026fALt8OJSvqdLYJiZ
gkO3kWV6fcR8X5q0sg6N8AwqQnEruZeT/v7/og2yl0tRUfc/qP2/vaH/jpnojRjY9pP0b9UgLSM2
CEcZ6nuvVVXrF9xkrtbWvjffIPPPpJeVm43QUJ6sohU5TjoTQjtntyOZBBQLVbOJm+t4DmJzN7Km
eoEdgjQZpYbJJ0QO6tmMZjVzCJOWCFPwnjMzpaGrm3NWQCV3SaFaz2/oMQUJ6fSMle6bubB2VktN
Hs2i1y4rpHmiIVlSNtiWAzm3lXmYIWGWTNseG5+cbOzszNroU/5dfQMffN9X1xSeYOLHNotUbL6K
LGOu3CBwZUSG//P9EEebGcx7dly0vie9OkXQLEEh63fd5JM/GAY13fJmjW4/bw5dr6PE7QeppQOS
oPOZBwcfNLSVzSW/EWiNPLSxPX0vvEqP5o2QH6xMh6ZppGt154JvnQknOLzH2Futxdx0N37QUmAr
FiLnb6Md2Dx+XPDpQHUHce0Yl2wocLMBd4XIH4q6K/24/yKYjN7otoLa4i6O/vBf8/AogoMskXK0
/EPKQsFp0LeW4qdmnfvzH2li0LYoW52BG+XNSnzyxVwmec+4NyhjtofU4xLs1ZDw9ujNkYqtke4q
oGQMidRaD51JuI1+7LVr5gjEQI4/evE8G7TbeCQhqv58d/jRkNs61JX9YQ83Lr8vSsmjMHTn/u1u
f7pj9V5tqtTFYGKKQvS2OpiYl8wbnJ0dc5egTRW9xP612muAuRa2t7GzUuaqKvgt3gPFz2XP/2f9
8i9lFLVokTU5iHIR9mRw3WnKunbxiozIStO7j+lyMB4nFODyx5XbCH3+GahtmfBEryoXbVgMUjx8
xEMGc8VWdPYk0zCp2A64wrom2R+W8mlkYpBi12SCp73SJNdv+fOWIy2Nr03RLLkd9C7HBMlQ+lbM
kRsaFfsK33wItFZoX1pXdCklOU0XUEPUGojfRFu2+JYs2Gmazmo0WaediRB+McE7ZeuAYX7ku2fz
xZbZssnHdDgSEV1c5gZYpKZuvvIEHAKyHxWDg0aezM3s35MD5oB4M+dCoVo0QMxKS7CnL6ONNWeF
DBq/1353fBFzQAmGos1CoEArMiCy4rPbjNiLhoaDGLUKfHAF/KszFEX8dNbcN75wEnTkKJVw4CHL
mWUdQW66D8wC7FZ/38JJFfiwjUrzgOCOEqNApLyGIP6TfOO8+LL4f/xegxEDNT659NwWVr9F+JUk
yxhIH6fDm6AIwClk+5k+zFgcW9A5sGaY5IPXo4FsGBubHhYzy4kA92Y52imDtv80jUx5eD7NvK2L
ue9BduXFW39j9OFCQb5IQ3LE/Sg3o25/l5QHkJiaW0rHE7o1ylYx2qe8w8DQcizaMvBsAs52QjyH
/DOPYACu2MedKT3QcI319VA7r+Gd31Zl8MgftoxRhayhr5o4uM84oG2V4EPLTiulQkwwbd4fI8l3
5XMuBIiQyuT9t2KH5Z8wqPATvEOOhAI+WbYl2koM/xjB6I5+AxMTVR0boMbgadh/KxqGRrRp7odP
LRdGFfSqjLldt4IU7Ur1KpdDU779jc6a+DxXdeavLP1kYxEQfAXaWo+MRmtFWkRu0KFyVsPWORik
0egPgC+wGNUN1KZk91WlDsG0MWztv6I8xSHKGmLBAL2qPxlToZ9aYLO+DDspILsajfXFmOdptqMI
plOge8iInUNK4wUUgXdbvrxsrKEK+I/iItVFE4lZiMI6NlbyDhOY+EjlDdiDiNeKubU1M5RTnj04
8qiooIbJJDQUQi5ntgMV7fkiTN6SewSicBEqaH34dr5xiEyQdHrXb9SHZWYV/TLszXSCSewkPVbx
FS/0kniGKP1yj3pTf/+d3iQY4i7hj0PxnHahkPb6nbi3nCQ4pa6La6CvtvAXej84nxhy6x+C9kIL
UNW23z19JO3mrTcUwjvIiiphIQaMlhAvTvBhWBG14E1EKuyd0AUAqyaTxxBRIzzEmKN704gDFapa
S+Uj0OCcfcxLY/v038r3D4L7IHLYllF4J3n1LcOKejb/EOG+svEiwyONe7PcRqf591oTwP5NU2EM
FmsD6waeIz+hOx45eOMvZPSwbegwJdrgrUZi7juDp1+a3EnfaxCbJ58GjjQPJ4QAp1Ajvi+2R7uA
+lTef/32dSZbj84QDV0gxCqjDuaIaXwmB38ZbsNct4WMFrpvJW6tTBQp+ZE2gwmj6xxMAMwU5DSK
TpVVViHgMpN/PBRTJp5aKojlyRf9ODJTQ1fLlWg+CCQgiVZrt0QRGtOwPRt39i19fmCV3XsRIneO
/8LoW1FxGXiRQEQ8GiqGRxGIsk8bNIskSBkBo9ZrJ5KMk9eHTBWRVBHcdvBT7gw8fvkwtDs8v95x
70hf8+Zmge9shDapItqRZaonuG7D7W1bxTeCoVT6OP/8kkIA2hJI1A6XKaqy/VcuTR0msz+QAXG8
bweBrMiIJ6s7ytCiOAyaOSwBJ9JQS/Y2qv/xAE0ZxpF72yYONAVOXn7Sv4sI/b5vN5KayVDBN2md
vBZV+nEwy9NtlHHSdp8E5k3u/ZyTmoobK5yl1fhOXcaTfKVd3cNwy87Tul8+JsLNc0O+pZYwuswQ
qOjpIalLpoNDgptZyxpri+06ztCCCSinRN93BbzcX4eXao9ze2bvCGD2jZI+VNv1MNklNSDM29Wp
W9rceacw5NJhCz1l7JeVlxwfpTnEOOaYUgvrCnyB5SwQtzecb4+9pGebCugdZr+wOOA3pr5vkxCq
5ycQLRwAC0FvrOCMYgfy9s0BddsQjYFU9EzMG3LT48aan9tHhTiajFLiW40pFAK98v0Z+TYVEAJD
iJJ7401WjpDQZBLFDNhzNURTP9xvFQ02X/+iuXG7/lCZn+MbCmoBcyr9JYNLETBhceNIoUUFH3tu
rcVAU6UNded4//E3CI+7PE28GoiCSnqy21P0Ekr8BkGjgnaFkV1J9h74BBHCaulbKUI1ANIn37uV
u7LsKnXTPFdl1mZxuwRF2LA/aWa7dpnrloY3fyr9g8lyPlOrlg9sdgdQN5pD0rw0BaI2nKOWMbsY
bDBLQcT3Sa05TxamTOsZcGqysIhsCAlvdolFf+b2rDBq4zfYMSCBDNw5uMb7l7U6A7XGRz/qHXLS
s2b5yd8J1ZNhPDRNf9/btf052ip9SnJ8DZ4lU6ToNkPbafFOGTh8Vyjx0byS7ahg/fCJOkzSe/Js
gLYWKyhzV5Tn8uG5kRoQWNbzWxrClVSfBCN6dVmDCHGZYes4A2AUMnPliXjRvBaV39dJ1mxk8O8/
+HsgH4YOoHXnMtl1q5llEjKExCYgBtxWq0XOUqxHZmzSjAoAQ0MJxRaY8d8hQZMiZGrecLKCfGEV
DRgW/d6oWuQfH8L0PZnfmjXBCrSvLya2euB72M8hvKpyfX5X4WXGCR0OJBjyQO7QNXrTGq9CYQpO
51aj0v+++sdn1wDlD0Q06tlF684ZfGIVeSllcqaE+Wv5xhT2Lev+tqgTZL9LFh/TBLdDdZeoJzI2
Co6d1jwPmFAeHLCRmhp/QQ13GpK77H8Z20FIVrVkbY0omVxVckLnWpMSB+oKSZ80evsDCaZ8qoc6
Va0fP21BCtbo7fnzoPehW2iwRbQDeQ8yZ7TTBXWlEAanG34rqb1cae/ZsN8fMty7o5ZyQFFlX3wZ
mJbRqfCjeSxo+cnzuljqUQZG4aXdVKJjic9g801AztTq5Fxc6x/LcK1pP5qVSzyW9MoWkdjkpGU+
E6IAaTJB+cGECSTdEbemPhgkWCpydxEmYGK0DXg+908WH31OCLKPT9RVSBLqxGS6ZzJ39B5YXT0h
H3kjBxE6CG8JB55ouo+VQpRBuBr/pf1fPTcM7yfzdIlt1Xhdbn2IzMBkRw0txtHfA/21FclRG9/W
t5z/wP+NIw0/OSwRkN117cmBLMvBdXJa0rjykp3/9OcNPQDycO5BSG9ql9YZLOOuUQPL/cjiFdct
fYUfZ1W4dTBsuVLd+u7zjQf/dPVTsETCPBceVC4tAli6/X6kzcWdXeL6K9ZngI9qoqx83CoMOOiE
E9iW+pIljmPHcMlh6Lzx8sashdKHl9kv0xHZhQuCNOy/f3fq7rbmtT+F2OYdn5r7K1hBcZK0ugZ4
agitboU8J/DG69XRP47LIpmtD52K57OY28b/4ZTBT37u4FGJW5vJDMtHkHRpmbN0pY92nuuAAGTa
G8zyl7wathReyMM5itBM6qejrQbVFF+WwDqZKvbi4dqIHbEmG3sM8buXc3UKIMRBtVf1UnQW3uZW
PHDCMmgsqc3Mg4dIIvs6l5NH56y05of2YLtxOVn/UVJgIpUn4A5yygx2lGiC7Y/Rap6joa79Cwj0
Cr3hFScVNNujTl+GkVfhjRvoOSInoEJ7IlgOJbN1hYODT+OL0sVhVclA11bW8SoiN7NFOkLOQT7O
siFTt9EwRQnWJro5zkmrMgW0nawCiAvaZdBj/PMjTXkscAVHAs4Z5qOrDqeMdeOZVHwme7E3IbvT
rpKfGU7OzzrDW71q4wIZIBrW36xi3jQpxhVDujwFVSZL+hh07goMZEnl5nCGVcTmvyckdpdQtnNY
NtPTtFakNIEBQmVbedGSLLySYZ4afr8XY0s0713DVlk3Ntf/NHMhI/efZpCp+ADVrSWIB4avhbA/
08ds5/yYveE84HFqX46Ca8m3+yxA3UGJzScVeTt7q7BVmGL82NcWVKza8VvLWht0SX903kbXSojY
mHXThbtJjKpqnknjxecz5LHMwpl7fACY2ChdR11D0uniBLMBhNw3TdWi0gPXUTl2/WI2BR2vFXS9
6LgcpRVwgXeFw85vVUkrZ1Ds8PN++n/txAEyHsJXBVwSB+l/rRVNDli2iEu7wLeg3BTjNUs6w4e6
muArrQR32N5Ba2rzcpuBgrK3eyLKRqk+wYdcZcPUnmr+AHzNSdSIKtrqUceSTX8ZtuCNBegoL0y7
2r6XwaxSP78CvrMDkrk2CI/XNCsQI4lWiGyvjSdnxsqWA1AdD5iEnKeR3zqjmRk5q6wIGsU7fWJn
4jSUljjEGZlPriCPkKVKicN/GnwvGaS3Qa2/pioo35ouMj76h7Zgw91DiV51nLzMU12v84WdNxLf
5xBqnMczoUq7XMhkxWqGxg1uxqgQFlwG4PUBrjXtNOndGpHd+HJNCXVx1/4NXdDZvUjY/Q/18hWX
AK3RV8IFC1y3ORKhzacz992tS9QFeABhIBZ1/wUcgDCRoc6ucLliBalCsYcxpSSC3ds+OQGLb1lo
s7QwCZw62NS2tSJlRuSFQyQe4fxYnxVYHYswNDSRnXgKNoltsb3UMibRNhnHGsNNOo6cuyisqUqL
Gz54laJXFfmYt3NLZG6lpr72WIeQ0eBEP+pM1YktNKZWxTR+I7nSriHkX7MBCyNRcquTDSQVpb2R
hnPtD/3eMdU2HV9M8wMPk88316yplyJflCrXn8aBOPQyTYW9jowALjVJavMaqe52PYUEx+fw0qOs
LMrYgrM0OiGZBJpx+Ic9VmD68aztWAdjV/Ce/SZJ7pZr8DadZo01XksfARjsKO4EzCpm0/XSnzzr
NwFouqdWal5n8EUvhUlPKZBOjWNfcm16qzW8hc8baREWt8rMwWIvyI9w0qyV3KEQ4+4XpdVXW8L9
iWydXP4DEAcuwd3V2B8GQrGk4LrJU88Ybl6baUCr8Fac46ELFsNE5rr1rVPoZ/eXSdH8WJktoQ1j
T+VpJXIWzEMhqtNUb1h8T86ZypcJuZ+9PEKJcpyAedE26LYRTNQlUexKGivYqyamV5GTUCNogWeF
TyzOa2uaXipz5wkyOGfAknUcH52Wqm1z2OnHfpIBt1O364EVI3ws1Tq+gDWKYmcdsMC28jKjQYHq
9Zq1+2oh/PjpxhK4JtkL7J9OfTjyBMyye7vPKhHBtHVmhv4ppGvuYFuUmxh3xKjb+bfR1LK9Lr/l
i9q5K9meQhnrVbeXo8KjTj8kKGG2kUR166YViXHLE5r1vWeEgzCU8SMKjxhYAC237YHySYc943Mf
sRzQZ5EqiTGMIScoPRgk2rMNnBnacQwP3orSPfHI1Mj4yKEgjeFB/BkVQ1vAqDb6d2nh+8H4RhGV
PKknovdw0QrHd5q6yKiHSv8pc/xM4rDD72QWwoYiJTD28JMiRMymBcTN8A2xV8+VPeVsBQJakjJL
KHxJR8zkLYJC2pwFOUJAVcxZa12OLZUlGMWd/jUzKgqWPJxcJDKdgh2a9Fo4gjO2kXBM2cc1jO79
WPW8z9jrBgf4pCxPaB1cslj02igbPKQDO2qpdJMN4K5DVWxfaZANC3wPehdIJrpzGTMlKHDr8B/G
YYTU1ZYoci83yEFwlmmgPYvJkiSvS9GTZoq8JZnsD9CVcZ9nu37YX2k358Yr7jBOODGhx/qk0+4R
lsGDDR2Uhd67INGSlEvIM11SvunW5RBZS3tXANcsi2mTOPgeccmi4Hbj+WjzkT1RHm4hICDmkj/L
wzmo1UkirijI1k1YhgEfTsSaxDd8rpHzU7b/lFLqmres04eFeV1La97l+RH7ygvJIZ96l+XV8oGU
3Sre5eUYOGlmATFH4iGZaJCI0zXjZHWqv/wGrQ6nI4oE811s2/zEUulNT5p4FaAhQMXyzPdieLF9
lyGChUufud/tchSwjL2JQK4CsDNy5R6NPCxRaZdgdYKQ9H+weyuczj08X3TW6oVg7UhSf3jOmd3q
w2r33LayaKbe57Rlnu6y5YbXBo0RTt8sE0zP7dV1gyq2+9e7HC++3iwxAT7JqELa3fuNDNWTCkf/
MLwKERPRT3aZs2/ZOqClI4yoiF4ejzo4CKPY8hyGcUeZjDhEpAUPoSI0fS03ced10SK/iUBE/eX8
4KnquAS7sHySyW7CIw4sm5UfFbrUI9MuS9HBIQgapnigaUJTK/6j5EHknZzuNPZas68779d7xj8H
OJGy1t1hgt0OcGiHapg3zvMVEhvubgTrSraeIgdIWCD+A/8Td18uxxj9yNZMXCscItFX6j6oPs4G
JPr35zK+36l/O2jcuNBfanRsNn3ZfEHbaPOnODvL4YIVl9leIVOZntmMYImyd5voxRX5myXO4Ozy
7LOjM1ML252tm4riGgqr7mBJgQEWX6ci1zQcxTXWTSdx1uojGRYN+vOwA82o6hRbATFYFPhNxa+v
e355Q+eCcBuw6VMPGYbFSATDU37VbD5IL03Po4YjWhKfuo/vMgfLFr3D4wyYrBCHrv64gb8ad9xk
aVoavpFv4FQJsZY7SefM791xH9sBl1VFSyUEo3WIMurX5NQFOb0HViT82JSa73MzDP10lruyv36R
+4pVrgoNOmHLKzcS/JfSB4Ndloo6fGP+H9sWLLcYb4oYrMXCgRXkATUboVcAfNsKB09Q4Oc9T3Bv
4iTQiH1M1TDx2Ye7GowXbZWCPh/OhATpQ+Fuv56iRk/SEUBqHCxp9sJYzBn3lZmjyd+OgdKv2c2G
rJ/ZGxCL4PI0NuCJgPYydge/aDtVgDkBAUhQLa/V7OtYsdfQCOAg7G9tYdYcnSVQ3JS+u9gdhqA5
jmBRMe0gqNhe+C6YgQ5nQCxN9K4hZOWbz9TBmlBdapSkwJ13CCemogfpGUeqMTbFyYJlPdCqflt+
uQ/3T8+++uUKhFxh3RET08I/z3IYW6PIaEi9/wwJgV50MvY5sKvcSWXFl2CQ77qS4oSWqR2yOwgk
j2oZsZfqw2IBHFHXUG9aziIMotdafZgWWYJmT86ST2fwOUEI6C11+HGyagEd8Nldv/9zOyxCyoPP
wD0u+93aNeglJImyGoTeQ73yR1FgFS+x0zj8nk/v7kM3OhvUgvw8g106VV8PH52297XEx2JkT8XN
d97clWRzCik5RfYQ/gq+bCMHirxB572tYX5s0EQEoDFZS8PFdrANZ/VidaMh0TokxHYN1ZqeC/NB
g5e/XNnhREGXh1RtXxUwDFiuLAp7tOuMcFfi1jH+dbJ1/yRBwbrFGFaNz4kM0OeVPWIx9Zre6YXs
o8PBHewEsN1UfW1UwbH/iNqJvMSqTNL26MBZRdpWCSsFcrS6ukd0D5LsSl9RKhE8ch2IwbY0epqE
YePcRPnky3GMAun/HHr85BX5xg/j0iGaOQ+yc9Oq//jTZ8nUPQjpMF9Ku0RNLKfcwYzubCLulnBS
V4lQAHYkdnxp5zcCNcmkjZ93T2u1pu7JXM2KMDRa2RLFEnol8rqVwKFPaESevM+pcK2ndv86NQvn
8Ogxpa3wvPbuiBu4IkNiVlAnzJ4LUCMkVm+KM2EJHPTQHt+8pFNjSv4mF4ZhysMuLH1BYLMlQpJ3
5WpF4DfmRikZyv5XzATL+Ly9JeVFYpJB1NLQXyTFbUz4LgfzQfHo63h5Tdu7sNjDfzmryXgOyPN5
JVsoE3NM6k00YArCGZ4CDaCIxE6W1nRg9q6BFj1D/kNGKqChWF03lBtJ+pZ1PoQYXbqM6VqGD99H
0ggME1Ek7zNrrzzjxd+YUTrT5qQ02PVUPam+Mf/qh8JwwILi05f3dp6KLpAcgexoRlGwLb3ILagb
elxcDuBoJ0vNTqyq2VykGtisa+q3HdSmBoPWc5qr5m5Jrc76lTBPuOPP2MFgPBTt5HK/kaMy1IUf
DGXqeMzN11jaMMwk+bv9izM1ySX9FMK3z9vXSskk5tp2l7yr5nRUdKAo/Uq4LrugIW2wRwlL7NX1
BjFHBwWDNkmxENS3ePPueaIQRtfkx+ZJQs54nuRWXYD4Pc8GFmI+yAleCL6DxcFAnoLFPiTOp7+c
q6WNfT/JfWGWXIY8PbwfWE98EEyZKV6O0reJ6k+z7f6qEZErCyz0URyK7rs6xzCgjCzY8Ppdgu3v
P6taSKXBZIZMOZYWzvQmm6h2tuM33r0HAImkJAJ+KdfnGoRiI6vUqlTGeY3F6recG3nI2bxeYI6n
VOywI5pQooHYzOSdvWnAdIvQ0hLlEMBz0dolSi2cYL5I8qM0yRKxtqQF/yUyKIXa4uq//6Js0J17
u4Co0vp+mKIiQjqaRmkIHb51/fhsLRzEP1QVpdeQH+gd/IRr9+7fE3zQc50Ex6346ZGFeO7K+7CQ
7Jr9s4RVvtsDWpHFyBlJ/Wjc+fDFEaV9JmNkMxl7N/TRMuaXElr5GkKmpOdBqv1XVNLkN0qUu3t6
jFxBUZ9pXqT6+jQfmaIAySWO7UcujM5zNlP/hM41VXjChNMFY5g1bh4JB5NTf3eKa4Odg7ohVNQ1
VANNhJAgkUu9JL7vgXd5NBi1fKenyJ6Hckr/jG2p0+hT9vRv13UEeoGad4x+t/HfnSH7OyaXXiQB
Wu2p0SuWULop09Mej/ObDNz22CIcqhrBHQy1QdSSw/79LRUDDXObJBUHuaTmk5e3ClWXuU5BUabl
rn8wv5citpoY461ZWjyTBlhuS+5s7h30fgMjZAfkIrnbNe1ZcAPpANtwe5UM7fLK8TiGmQMfEW+1
1NA2y0R5zwW2BB6/IbYtImQZYKCuqd7JSKE6XqFF0nrl5MkKb2LbK+ZVzeK5zNOVKKqLzKIdP23z
atlkAn/QakQIITu7GWgqUbcIqncoHmx51wELw5FkfEvqKuY8S0Nec1TKlDdKU6tMsxVEtxSXu8sX
loR7X4r1pBp6HLWLkSSjNIfhN1Btvv+3VvFirRO6Odbg5XhTUPh8baRqklIHEHe5lktPQ8IL1QBA
IwY96vG9D93TXILAfoC2eh/hoAIk9EP3Z9xzEZSP3YtlIprQgpSqVzlFf252GrlliPurEahRaBts
0wlZnTEpzheib6LJaziUJj5IFEJm5NedtJTNlnxR69WvVHTkdVOrYekqqtpyivN51EBTW+WvZbSc
PEmE2cB7ct6At1Lg/DySaLfwZLiiwyFlW/cAoTFdHwE4sMbwe/+McXJK+/JHz/28s3xlhMC9yrV8
JWvOKA7es0jjyFGjjiCV80vK2V9JmWPU+iYcIq05yQs7X85YdIOMVYlxDDUcGtKu8DMY9PbMz9pP
SR3KkBJLmPtqT2ZaJvMHbg3WB41bSSSQkz2w+uVZPzYSZuxaoJAoNG/RYM7fvGGlDb3GUD1y3hGT
hG4G/b3EFWIRR1CBEWQ0f6p447jX/QuX4BdO9QG2D0UCdZ2QWuhcwb155d6zd63ZR3SfP0PM5h0E
tyCQqZgRZLXBBa3t46cvIQh83PJgjxIKZeYdKPHdVxkcYkrcF4cBDQmN8/Xex8yJPtRZRF1NUsYF
HzuVjArdLi+NJmlZOt9/nQTC85AtPtk5mKFUpFQUZojFnILyV0H+1wh+2ZfJ6/j59ld015gvFrEL
rysp1QiEbklW4aLRzfADnk41/JaDCjMmq/hSDbu1dztFB8oQ/EkgIL25NHhT/qlkFKTU/B0D+fEL
CMMRDCadZkol/Ard2I6szYvBycsJdhC9TKvEG/UJj4E1Lzbt5ygLEIdMMICC0tGRdBgn8lTh9fIj
6CLPSudARBaIj+cboXM48gFVHpEbpr1hDPs+tK+ao8FAx5SD7U1b2Mh72BQIvh2WvEDE+KSBVCOp
+HnLrc3K7RaAA4JO9g0Mjna2UEE56UYBc65etQMo5ENtcpQ1MdIyJTA5c5s5NCT3DNHGUxeaQqCy
d1VfQHRzg/fjHqvHnPC5PUtD8goA5Q3xSy9yKfz1KbYegeFm8Rw2Ht2rqT8M1YZgWiyWNJr1FzMj
+HUNV7qJePhQFqmmyjDcAp6v/MM2hVlVt6CCV3dcyqWrr/kNtTXu2WgTAVXFzud9q42XN0HnRG3M
llAN89l4CIXupRty7QN0LBv2TbaKWms7np18VaLjCHsK6q7zBdc1D3CwzhMAfnwYQvuzbUk2mVD/
feEiAWQj7vteyO1xd1dMrY4H4zwpWUFg6H6fJQ2ILSSaHRD5sb++FqfDnbl7ZPWhu3hufXdp61Pt
n23i1KDvmOsA5ofiMSEzpp727oTegfzUg6iDLmpGjZZttUQ5Y15sTwvsKTl/o2t6uagHgQycp4df
ZObYP6t9csQ/BUndhanC+257NtoW2WqBv5at/qAUVN6sWnDWmfnsFvrvXd13SdL4iQjHaTKKwqE5
PdlnTNLGsKWLehVozKO3a5ddmPK8Xo+NLt/OP/RWcinnzMJfrqS9kqa5213WojyS+nZaemwVFkT2
bbLT/QE+dTj6LX4ZOGresL21UFZRpldz7MRKi02m13r89bIEawm4DhSv1qWt38JH0VeRiTfSTEiz
aYZEp55sw/0fCoVh3PCjaLoHEMkDUomO4NppknlzLLwBmnZo8gSh5PZ8wkAMuXsMEX77ToWfZ7PH
T54Wg1B07YBLQ2OSr4LllwnXZkXmapLcXJcRkJvkfKHvWrNROf5PCToVZ9EPWfWxnqaBMYi3Tq9T
8DdkajaLNkBS8K797McPLVxY+1a4a/Mf2PQP0bVCgxpup1p+4Z61mWN52Snu52GHN954vdJGAHBj
Lge/VRforA3Znk4FR0IxhqD7pZVqSLspdW0w4tBnL/R2Yt1W25/1U/9Py2q7RZysMgUjKfGaDI7I
M0tDO0Qqlua2TboCl08aP+PwHKEiyCSrk+ICsGSBpMLfVgkHbDeMYcelGjVigO6pmgRolNEyJiXq
a8TX+XALvxmAw7xGEHp3E7oYg+d13ztcC1PtPa19vIeRgRx5zVQNvAm2p+hDP67iqLyxxiIQA2f5
Hlm5ENtrgO4any7Y4n7lPo9aD/Jk6RGSt7xFXj5re3ETMw36AGhP+Fr7oVKKZ9oaLES76cG9ktdA
yOLA8HkQvJJNrgGigfIq7es0oWK5btNoAn73/sjqSUaOvHhSy/YS7Cr5NUh6DhobQ5QKwXIvxNvj
ahZNeqRMlEQKVudLUpb6yf1NJce9SrEtCUFEHuFmCMGAIbJg4nmqZ/MFF3O4MX7IFNY1Uil70k4n
K7nBG/Pw5mRdKiai2OYa2KZH2NgQguG5gKRQx9iilMkA08rP+3vuGl1tK3IDq1QoOSbQ6KBrq5i0
zYZN1fw8fy/J55HqnPMuofrG4ACPXW/XXHQhrNOewC9rluXL4oN9JSjEpLrskPQqO6ZNcAu7PWqH
EYo5BjlFqS3dFrcq2z3znDNFDTC191+xv8K+j9jvlmNZnZigP7scl50i0Eym6cyexkHvk3yoYvJU
XH2/itQR30wWHrO+HiLTDmXEFxSDdA6t5fJ2L2vKbWxRdneHaOWesjpJEyrK/hFyF39nQqt/k6hu
vcRn/vNpFLU2RaaOzg0jHIsKP3+Iok58NNohI5JVfJjDQLadh5it8+2Gx4nEq+7+YWZs3G/7J9qi
u0dpAQ++8cffj3vwJbf//hHczNImFnh/p3HfWMoHy3eIc6NrVVLrrwraNNXBQm1seArefdMc0zko
1X44po5aOUDpaus8O67zArKjHDQqmwVSpd8oN+S6uBIodcZJYl61tw2/Ude/RwzHQQZdEHpTVMED
EfF1FDRM9ANjv2TGUYAj2qE0g9lGSMG36Rp68wiwkzOrElRkQ5AYH9ymzqzbBln/GMwu1tm0U/Jr
LL8TXAhkQTtLwaig53LhTuLwlTyTGfPlJlZ6nZWAgnf9zWjtM9YR+V0XpyQiEt+UQVwRzHVzMmyH
mVqdvICDsrMBC96Q6gRY0g76hemrdfHYYPSiaynfTLA78ZWMn+zeWNzN3tCsRQWbB/iu6hfwyRZQ
1AniV6RkXoMePE9v8ZKnGkVAZXcg/vKK8WuVLmOmo/UHpddCgLe4SJHX6/ulBQV9ZSBOBHPY1M3k
D0LzyQ6Hm5DvJk2g80aPiWd2sg7DoP5v90z0XYei/W38aXXI4MKxcBM8mUhup/KP8mE9ifkr6tbD
ECD9dEqoj8JgwOE14fC1V49+LFm99DeXP7f8HeGI+SrL4rhursM5sktXc6FgvYqUrGcVWFxF593f
l/7gndyUhgH/C0Ueh15O5aCEag9YsEcAf1rF/jfJ2tl7GhRWRG6xTwbLaOaHBr0U2FEU6wRQI25k
yA64AgqN1XznrschpeoaZSjSs6VxAJPppOePimLs7mGqOq9+xO7lxnEfTs6lxEqJwjLj4JLE/Vng
seQMTORtWV9s26lGlkbRAq8zL26VpsSzGPl2eeEqaoje2Bbawam7uDafgi63CgPW9g/bL7FLe+/t
L35DSqZr7WqZ7V7hwN4j2jqZ5H6FjqyyL1Dx0EorfGjcAvKPm0dsdBiAqMuM2UgH3r/zld6eWFzs
Ha7+ro9D49rqbQCQJfKBfE2ADh6Ezpd3W1VIK88jt1+3nwhIG2JveZGhjUt8aYkce0rnRiUI7i1A
on33fLy498NPjAyYyuOF5w6uYWMO6ANFN+wAKS2kLBgDLWVTaqvwpP7QOgkSOpTpnXNumqb6DkpT
q85/nFYMPGpocWy9LL5OZUrYtmjjofJkoB6/NZQrMroLSzjoOCHcmBYTGSf3crGBxJId0rGUqY4s
VCG/O/ybKYHXhz+/tx36OU4RqTr76wZ7l1pApyVbXVHBmd/nxF6MsicH+wW8MCTzVViuB5Zub/xU
PfaJIapToK55K90lszUL+Vr7HfMNIMI4ImQ06JCNbxXzCR6nBrAUAfxF9bUEVFHP2eBoZjrV4ALR
sW4eSXKHUtnDF0acU+qIBknD1DvQlJrZ1cXoIlxIIjjAIbMAZtCZiZ6GEBtNDddwVSjGZnQWvl7H
yDd8y/kOI4RRBWghvUb57v7nDOH2aVJiMHKJnfjp8Ye9Rtqod+cNv4seaY/e33oka1G73IeCUtfG
nmHNy/3GKzMCZtbGjiIz4LGD2tZ18aTFUvVtD5xaBg50KJqBOY3vPooMm4tuLPwU/SgqcvI5loIX
5ozsBwzaZMkeNF1Ejzvj9XaAC3uOLTCvzDyO9/4LJYxHJ4OE1nxIjVGChmnfQkPZl9S/X/z4+CMX
4AoA2/IKxbpcjAllK0EMM1WqyZ92R79ZusV3HKC4V8QJhvM5R+E5WAK/KqpUx4+wHiWHVja0U84i
EOgQ3RC34qwhuVhQ9NHQO+AJpPcbMbWaUB4SKZjKwRz5ydMmQlq5+doVK6Z3ykGsn5zY29dOaiFn
9TeqmLRwp1ViOFNY20gA9qCXpgqZJ+YwrTqAXg0ccXJLGRbRaubvxQ80L7E/3n0/V6+1EzfyiZOR
BO2KwUbRY6jISCXrXr7RCo3/eP81348VuaTJrJuXIgxauR9NXzcUYXMJjuEKo65z4JDYbT5YYN/e
gomDTy0dDTaeNKwl2mR+oR+gOFHYuJpeLrS9VRxxUqur3gNm8AjvJdvMau7oaaWjAL4HTybMeXyF
jCr0RTiiegPGipBCUuA5wNZaesorRHkRKFA+WKTeCawZEouJ/O3eOzlmkyhjcL6RfpM0Lez40IJA
2xysXXHif/OrOuT+KGpzxcaCCJ0QYX/qsJ8aTShswzmK00H2ICnyBuRuKYHWrJHg4knDxNvRFTSH
sSRiy8HZEIGg7ESOKpee7FEM21AVuOnrc4AyHXX2DcwoTkZ7cZy6sRcgEOKX+3HlshaIm3UMjxDi
fhH1Mz3rwqDksvVzuFmIBvcIrS0Tb+I/f6PnQTpHaI1UxWShK6UUoKAfVD0wXNIygAVv+2KmrbzG
rPKCR83Qdz4tO5EZrss9SqYBiZphige4+hVL5lNbEwJF/HZpk226XbfDET1eghHg4EBniny6ZZPs
8+TmdWdqzgINMQFuMH7SDIKe7MIORtjlTXSbLzEWffwnqCrF1ILRYSPzONM970dwFEREIBEbqwm9
xTCmPXWDflfU/bMUojbPRCzC89YWXZgj0QgeKT9/ZULsW75+ekkNRwZwRxchEdHmjGcaV4d3+m+0
Tds5Ys9sEoBNGIwDjCWt6D/gSuJ4mFNFmtykaoUZyqZ9q8oGkgrLFs8mN7h9/btwQ+aebRpIsRib
11aMCb5EUEn9hWrYf22VLlDxqqaAhqIPHWJ1O0JkI3/urooBb2g6R6Mi92tAP3PmFI674wfPv/XX
XgSRJSPpTz4X8ylK1aIzsMj1aL86xfq5eCTK7Ni6PYzPRIMCTRNAu8n0nadOEtlea6j3RB8KEJ51
QITVOQXnqllkSC2y9YOVNrH33v6l8sNj6DLpVRIWs55pELe0HHGngWwEuYNI2d0s/EIoii1CH0Ya
GzG9x4oP4OXGPihQPI40tO1W8TiAA4Fst31A8jKnnG4Q80C+VlKAM+pJJUDbkhb6weA+2qCO0OzP
V07ohfw3TcpUPnAerTD0rrEcSw/PagzHP/y7JHCITErD0eXT55a6zR9xydrgWtDEB0yxovJRCI6s
B+NaELgxeGO8+x7NCeGSCt9NhtnGuI+NevckMbIH9a468MVvhKDQPNBqeBBB6g8Xwet+6gAchbAb
qh032YJajDbusxwBJXwMoneMkO+FfLPhgjWLmWbNgfqe3CtjVChVjZkVkxEa2tSz/hGMJIezC3U/
C0x2Qao9+PrvDnYUWuMFDJKwUhbNX9MO7rSMYUWZPsl1tYllNXYb9a3bUN/FR37tR700kCayYXq0
62Nuo4akozJaIx8js/zhWq8pgglcHL0B0dcKFWLuLHEt31X7t+JGTw5MmllFi0m/eRU6s7E0Bduh
mA8Q3ERcSfiv31qGY9nqPToBCWAL/VSHDs1v3EFfjbCuXJBK/SyYHp4GiKh/IJdSKELi7EsyOnGp
r0/asqsXfz/Hln0ZSx8jZaf8Ch8rSQio3yia02Pb4rrS3VKCfXuhLQewP/fA6jDoCfM7Ny2o7eO8
A+rUzs3mep6Nk6t+9/lOy/JIkStakBpZYooHd6kyxRgC6igv541LLste30ORGwGwrH3eiMba8/jp
+wz64WyNGCtZ2b1QsIyCG7Eyk2P2U1kyR3M2I9sr4Dvyu2Ck+HtqgbOJDQPF76hXcXYfwQ24qltn
v6laaiLrqUcM67uNXwqGfD4TZ5mOgHmiHnV4A5P8MFuI10LkqZU+f6+GPqZD0/QUwp6cQfs6OrBz
w089Snase7nSCbt/Fh7KCCP9MZYpYdw8lIBKL7vF2wXUhLEsxXzPcwJRe2Au7m7nW1kqWiQRbSn5
SmJp26dGfYjnXV3mwGP4/2oNu3xPERY+MCx1TtAt3OKC1erPMDuAlLNNHj3jUXf1ci2EhbYY6yNn
DvNOTcgLFlRfxAVU+7ttCC01rv7/+yC2S8KR7OxHMBhBAbaXb1POAUWsxNhkZ8EoCGTv8Hd4wQMe
i4ZP9SOL1vXL2Wc0N5z8AB8FsGy2RBFRG93fFPinE/DZidAbGHrtG8l02csVzzOo0zcF0O6EWWJe
DFSX3o6czhLcuC7eHW1ySNrIjhzstJskPYkJWzla8SxzNMmzS8fr7O+yctewLX9fJuLuh8Gh68mL
oXgkwDVYD+u/ZkYGUwmJQVqZrP+c2bHFougqJLihUAdSr5EofWWetCCObpa1rSvkujE7TmQApDnZ
1JJ/yr9K9G/LeTw6MdlL2zOGcAXm7pBNcLKfvkGGu/Gnw1RHfwiJ/u8LhnrM5Nz4GyHZU1xaHzQ3
fSTfdsLhCqYTEmWh8A/RIrD1LclwHQjXSzGGj1ycthrEo2bg2ksyXpHzRPzSyP32aO2NxHmKmRid
45qJH84HV8pcXtxnJCUbx1lkudmwxdI2w4DVg2CQKUQIqJIMCbfy+0HbQe9JBdr16HETurybCuAk
4mCyYantIoqWXVELwpjVcO8Mi2jWAXMvYvG/ksoBNBjp0De74hEtJaxpmL8ZVpcPL93aSF8GCv68
JqFGlqCMOmGcyrvqT+Wiz1ZHQLiBHSNOUZHjcN/e7uO6nZi4UazaxsvLVJOhy5caVsokigth/8Fw
WS56GISYaFzOCtk3K3HLdiEau/gwVJFkBwcHAOnE67TWquG2lOgd3ArSoXofNn686KZDBjKzYEBV
SSJXN1Yo7NI1lYDXm3jJFyMl05Dy0wAGuC8MtkRCsATZO1psoleP4CKhDOGyqhEmZ7x+nTzogyDo
FLRi8N5LaRbQQKyVcvk9PbSG15oFeg/wVobOy9vCqoad89xUnWOnCEl7p70s1qZYcGBlZfhFSIJ8
oGr1Lf2fjsSt1NFDkreC33lQIwrUNfsjOxiP+VglBN9w4fnekCrnu5WB6xfjzwBLQLps3jbTlLFP
vNMvBaSDPEWeBV/HCBBcWdgVLrkvamRMRZ8CFkv29aJCIplWwS9rzcK0zocVBmEAgSH+i83uEhxj
ETdi/Qt/6E0ddPEcw5zM5jfXlkFUHkfYFV7ZswSPF7MlYKf0xzhxhCLyNxw1na7UBqiZUD61g+mW
cw6+OGKB4qjUf+Mle09ZFFQEPEn7IAw4XunNaDZTc0SmukwnuZ948D6j8DmG1h4AIVgV2Idpb0SS
Nf7Fupr3njgzDZwmRHY+l5vWk/Se+sMz4QYlJjlfQMWsRVvDgXnUCmBxrcVWzDehpvjQWQcynWX/
eC+A3/AbITcsP9EME3rHl+guufxBob8HcgwrjvyLZctCiPecqaXfcCriZ2gAIZgO/rHilz8ueZN+
55+wemzr1aZ2Y53Y/dy4gxCtSoWM/7mAAalRTj0kuEDFCnkXsWqjonHlcUSExnzzR6dDmCBep9ji
cYqh1PyBxnehvhfyNWJdZlMjgtAsjfC0+l7vOSIdSwGnMhoFteEu2xFhQ7agpGCmk8kJuwhnOKK5
nzeItIYMIrRbWxen4HolqsD91c8vXbg/u/1HRZCRi2s3Mfzx2uJqVVEfEXUinLW4ewyPU08e7ol+
eEraf+oWf6Ds/2TEOTVosrSmTG6a/WPoDJ8YDKlMhCzzH8aVEAQmLBTnXRKHzS7+U3oIaMGDXlUg
Jo2PxKvuhsm6063n6BMn57GjbzONgh6wOpDkTJ1Dh9hpMFL7wgXuQtn/vR7F/a88PmAkj0/Tq2a2
s5hb+znSHItZ0TU1zzg0BQiFkrDef0qlG/b4MbU49PWbL3/sjGjkvw+TYNUozvXXW5pW1ZNss0dz
crw3OSCFdb6gF3/tkp77GwQZs3k8PFoJYU5qsp+d6q/b/chGOtXjql3aMnZVjorCczaBDPzDUQQO
HWDT3BKE1NIuMbr71X5iji5bSBjHkZyic9iaWKkU0zVdMAlA1rTOTrpVi494XG4xkkL7B+dydRkg
iuE2lMSC+7c51cR3+DMqM6hRM78usyUOefVU6DZrv4VEDZJaYjLlZJzynhTYAigQ5kSAWTwZygoh
p8QAJ8m2TEaHJpP8u8bNe4myHL6lYHp8d+/wP82uKi6zw+HqSxqbaFIb7aZ5Z6eNT73Vdm6GHL8W
9lYNmSQYxr6BXzSDOyT5/08g7I/73+yPuzb5UZ/7h+O+AbSzPzDytj7V6Xaci9qfknSMTAO0b9e1
tlyRfKptfgTR320xNRMjYFYvp4wQN3EGTUz2a+qPfbZgu7duGs2paemiTjSMuMx+uB7zfeoglAyV
R85i1D+Mk9nH39Rey/mfhRUantLFn96soQQ903Ms0KW+AdYiM1zmNPo+Zi56JnzC/v/hdjZ3XkPO
dDcvvrQD84mkB9wyrFLR8yTynyXWOnX4W2FXoFr3Ibhib+xqOb388QdxXGfINgEwp+tbx3F8DMGw
7QfJLGy09gRaZFGgKlpaRlxQvBHlPRPUSimH2ppDMlrrYhYuZ598TvFYMRUe+TnUK2/rxGUH7yD1
PfawKzvXSoCB9D3LR9wxl59dH5q3ERhEP6IIfAZL9B8ke3DVnyV7jiukIU3ciJIl8PXPPQXhQXk8
UrDWPiweJVp2WsKtUMJAGE3EjxEmWS4fzCKqckalwP9cR0U7JmnD48w0eFTIovKACSk0lz0yfzRY
FyLwjjbxyechK3LL18Te1m+/9LHlAkgzHEVnHKSm+ZRi8LP8b+PhvDk6oEiNuJ+lH4NZcJPteCxb
cQqxsAVhANCGCFyFaV0Vxv6iThVM56ZZk9MkBMKDjhiZeYF7avYxMqimGJkn7r3EvI1gZUdOZbt9
liBuBCgUfF55juCk/+NV9T6lCKyYWGv/RRUdg98ZDMXbFmGXeODU/rjAIyrASWM+ejmBOjj0Xbxd
/G8gjcIZwileMhJn4DgMtr1njxzT8CM0MHAjn6Ui3VD5smQK1lE3YGsD+AfL/dJsqQzjflWyaREZ
TnABGSOrzdzU1kk+PTHfGM9SYDiRLZ7DEYfzzCTBONUh3G9pQ78TrOLtbW5cYZ2St7S9MEOepkIQ
InehgaYDNthvdG5UjSS8u+J0/Oc8IaQSNkRxE8mfc6d+zs5z0+vaOeeUFgSiNi+UZmHLNDpMavMo
1QNb4JiW94ilPrECzZsEteAqLCCM+LJWYqPwFJjBZOqgMHVvXbkGzhU7BxgBDlyEVyu0+V8Rx4Ut
EG4zr9tDX1XsKNNR0AEyxwLG2+Xw4LaxxfFcqSjolxDcBXZbCGoJVQdc2KWNvE5wk0MCtCFHwB2y
pbxQWcXKXQpUHzF3OJ/nyZojQXip8aA5X5c8S1RHLKHHOn8q9nGvuQN61WudoIl0H23VdN+ZkcOs
FvXvK5SVIyvPYkYTYaCoyR1Q/DRXSGC78osqqszN5yqX0aHX4KzWhEcvJcXj1kM2xIayzVs+Hj5t
TH46IiXBUmthFta4/zsGZBun/ti/7irwLTDTH2rn8WxsgAewrhDU2KXvUHs89pNRVP/3MK4YXhg4
nb0K3opMC7j94Xp3VT3uVF117ujaJyEnLG0jI3rvf6tNU0LKMMS/hFTeGnd15suAbjsmqzdH2Rlo
pqMY6exC5Xntw32DOhMZz9lXz7pPI4SWgUWrBEOmDbjiJqa+yc1gHyh1rusiVMq+ZeLyR0StsMOs
i6LQIgRXA1chu9/N3xdmZa8QYVxDJ4jMbEICQh3NAe7ifp5aVHYU23jxgQ8vw33LJbfFUCgs8U5n
/NRXZtPaEujPs/FEnHxSWw3kDXZuA5iv8rbFKLLy86H1nNl6tQ6HflY/HH+uAyYGm/ZEBl8iG/hr
xNbLm7f4ydLtoeZ+dQgs24ChJZmPnFWnotLEJd944vlzhyTEgZJq9za9obaAR0bhEmGX6LChiRO9
89cUx3DyB45eXh+YYPAOERBgPuKEtAT4Tq1oi/xmdLImLVpdGZ9r5eDks28WLMgqH1+CCbVk9L3M
RCPY/hAW1wf+3w+g3gu6oX4YR33iUGsW22rOSfRuK9bqWdSfUEPiK79sqxkhw+IlNH+1WZ3+tR5D
hcKEl0kg0+uQhcxWcMDxZedZ2X2wiHQ5uJHz6nSwLAUYb6fFkTVA3u0zYJ4+PVuGwKMNaaNHsohl
y1cHtprkN2UtwDLDj8B8ydr5uP+XKxuCh+Qyh3ngxB2S0akrCJ/YcBqPshucrnT1+6SfwXHthVuH
P0BMkXx0tFDKblk1fcqNjJQbQsghvt+jJGocCPVOiBf4pfrGRAZrJGb0qaVmSRFXyyOAn29uuQY3
dSoeYyTusueYPBl33cVdU7zub/uLf/R9EBVkBCRauXyruoktQHH9UTrMc4n4oXtGr63N4rm6YHDS
4RfJhkqO5eXxn/yB1HxlymQkINTmhmpTfGvqVkNxF4Ts97kSFNdOduz94a7e6LuirPMH+5QPtrJ4
qYYL/zIaO/JE11CtYLuep7acC5teAh/3gV6Tku+6Ze2ggFsvb/VkmZo6pe+CTPf7NENbrXWXBNbA
VrHsEvsrkzGSmKNQvV1qbEI2lBccKlXpdcwrq7Zf4/lg9dvRZN/MMfF/NK4k3i9lhT8lxmqT0xSF
n5P/CxvhPRXTznVuUkaxF0eAjFIu17V2opkz8to+W5AcLT9QNarXYyJuPIgT5/ebX+51tQ/uNT+w
7WBMZIB+JNRsbNTj9rNWtRPPALL730ZaRMYLvs1IQXk4cnvLNFJwc/HMrQ0HyZO5LHVPA5ryzIH1
t03SwACrni3cSdtG0nlTiTUU0Sh7kUbyc3MiHU23/NRBnuk+0TebvKWvxzsxPErOBiQus5MCYGaW
Bo9OtdLCWrI8dAl14JaQFsOkN5LdR1Xa8jQR45jKtmte2f20XzTSc7JPgrv9VNS3iFlzGffuHFRZ
xngAe8qLkUoDh7CLET7ZQde1Wk+jytplr4s+r4QkCVt5vympAtBkP6/9BNqUfWemV7WoWHzr4zib
PjgQexITpAX8N4c1gQFFc4wdWC7fKyxK2V/nzsaTsOFzpVCZwTb1aUtbVMYMmM4vXWF8s/QWrVPj
YXVwSCNDfVrarFRHm7ZtudFvdcK/Oy895DbrhtOE2flwoEZZXvGBxT6yzSxs6DC05K8sonURfOUO
IhmPseuaF9dpA+OZhGuSvqLHVvhiqLnf2a0qytYJ5Rg57RrOTU/HSNshOK0WdsHeyslpDy29GJ2M
Z26ioyYuqJX6QfaWshfKUlZg2nyAn5neRa49EYV6EtT1gmJySLzlk6DrArw12pKyYyaMPcTLfIv8
RcJZ5/eblhtYB9AFhO7Sb9CcS4piR4duha6LsdCRBQwbaENstxAoEQMcMOZZCfg/a1l2o8NE6IL3
NLUOSurkqCH/NOEAk0FOjlVUiQUjgsr3F8E2REa6thsO+MwSNunvlY2qvucyxSL+/SL+ni3xlITU
Zmm5qYnILjENqRgXrCYOZx/WoLwfIx16jXLJkHobfxVPgITiSSnkYqj/JylErcYaca2XUkl89PFs
NeMdmsWsOqYAJ9TyXKPh9o1Xk0bu2dkS7htmC2l5FWt24MAS873Rwo2KlKXFMMK0WQcEIPnvuj1z
d35DwXAIsA5Vvl1HElY3ZxwF3iTVQwxLoBuZJsC9m/PiE1JLvdKaTwZzOWA7fvUh1gjWm5D6gOJ6
0ZnEgBgrwbDWZImP90zyX4B/MLpdMvChEIj1AbWMb1naqy5d46clDFyQ6TSge4mGJvgaSv+rrU0b
x7YmGv4GWulUTSYtQ1KVbARuD8sKyw36fEfbpqmud9rC1dEMHUZkRT+IP8SmvbLaX4fB+TVAPSPe
nDmANzvdNzBZsce7pwBD80zXRqdmNb9+kpf7yH8m6iSMQkKT0lNDISEc/ltoheGN6kPUYmJXGIXI
uiZ/b/U9jb/PsSWNcti4I6S88EHWtYp5xzakRu44TkBhH8A3RC2ooA+3LVMPnES4X3Q+l0TxH8Iv
ZJu18JU6OO7SZC1hfNFz6er6NUuHzGWal6X3xO8C44iQUmmtxitarpbM8nw/p3LURIXEMpx7woNt
cAASeVlejcuVk0pQBJYRGJoKfD+MxynLSCfSmsPDXEjLbNlUgEPFXZm+O0FzuRHqe0Wc+XJXqEu4
oE0Ak5Clw6tuBQPl8EP0+ubW+fz+UzdOkCvMxnI138/GEuFgWAVLuDD0WDWHzxQc82bHhoM7boZi
qS6YwU6WISjNmkIPksYnEsJanPMUn+DTy+bJlHOAblOFAI/zL2Jdm1miCzDHDag4KxoR9M4bMh6A
jOFyahx9aNrcPL8alD0Pk1mQNc/nT75uF74sjAhfTIPsBn632wYiXQ5rFECCo7foSyo7bxCU0qBj
dES9qBgNIlkmDhR0w2JqYJgwLpn/Qmoy9x9TmhnnJBXVAUF2S9Q7MGEagCaUy894zaDu4/BqpRMl
5/Qr4DZyhpymKdeoMMDGK6WHdI4yoJPGA5dUndAcvrT1V1/jYwBlwr1WvfWUypUc3z4f+r5ds8FQ
hP088WDBpwjTntSy+suFyXOqEkD8NWMa3d49yB/CppVsm/Pu6CCk/84Ll4E0d6LGLvDZXC4SpSZ+
qOs1Py5Df2S2E8olTk8selWlMHorLZHqJvqpJtcmWHQ1xMhupMYtHVSXtVOcj4L8Usqs7O7+9aRm
0RgrJ/kORgkkRaDJZakWp3hXiIr6sfmQOWsCuKB/hEa+k4OZqurrcvLEv/ZKYu02VJle2ckoWTeU
wwmNobgIo8+j/tYGRmcjQ+ievg2jpXvUm5pfQoG28TQsXUH4Q50TRvIZirQyR6+Ai5JunEoi3sM7
4p0dsqveLEtG2v1XIRQ4AFk+iZ6zUNwTEtDXFiSA31sTr0bN5y8HqdRvjTw/85VghOQK68urjNym
IUAXzPwHAhb3I1+D23BbH6mr8ZCititRDC9kluv9n19QAtKmB/2CbaNrxwZAky5zrgTn2/UsjLZr
J/kKsAIh+WtD00J/Qe5e74fri0rrdFW276f7ecZ7a9RjfnQwB1R1CyEFZMmQZznUmWdMaFW/N6wA
pOpnlDjHmZ1w6J5RqTy80JHpdAom7B0yibXdhaLjoA0Ct9RsoVOxu2Ggvk7pFUwQHN3nSOmykO8a
LC23aiaydgYPdOdbRURAIz98mbSHmrPIxVE60+QgRAnUhPPqDXYy1KHo8Nb1ofaaCiV9Z5HnnHx7
X3HCbs610AKMFNL8I8LBdY4MC7AYFD10xfuKquF0wPfttFFT0MvXQp/vGuU7cooxoIQVBJCVyAhT
bzsGHj0QC0Wt/BsDu4Q5v9qcu3y0lClJ9FlF/3kN1ggDVLgYTPQR9Q9Wuvn5rA5+JHg2eSK1nHMb
y6+ogxoPFMB5V1toZXbbn8yX2LDJZsIZ/TCYbvwB9+wZKkvo8UQc8NPvAJpQ5xIl49EmUzXB/r9r
XtNyEyr3SnNSydPV8Eqk7G895jaxyuCZbnQzpNSzNkRPrWiX9cjl5nOjYwDVxICWvNjjItv1M9Z4
9WoRirjBqmAPyBn2JHNYYSfJor5lt3ss0aMKH07BHmFV7Dn2hLUxbzgT8d7ZZqdQmgMLDxIvwncd
8xXqsN3St3gn8QLJjMJ3f95fiTgnNwjNdfQrcEGoZpCPGUAMkm4BNIBf581QV8tJy7Vw+lDHkYo0
ByXY/G40vRge3RbzYVSQKF2CayWyUMQaB3hOKkj/fsygFwkEa+UtYzQIBdoUExfqdisxC/bjaldp
bJ62KZcPmyK9JEfpP8/SKjWBDE0OzLW7gR3U+IFBvu66hBZv6Huj+w5+prCfyYPADPuBBhtK3KAx
hFvjLE3oH4jb5q0mC1W2CrF2Ty1NCqJ3Ze5Y5di4wmBZ+wbvadmsTZH6WOqSdBJAOrQZ+MRidxzy
kcLtG0SqzRm3Eo/UwfiAFjU+5emCsOIJIIw2h+twgIGkA4DBq+Xa/JZJUmB+IUQc1MG5DysUS2s6
nb1AaG2pkkmqP3O+vzGZdLfl/gtBGehxH/N70CiOCCjCmCiP0ztCwOoY549MgvyZZJMtMx+lUA7f
Fl40AKIzsj+Odt80q7XSE6xxlz2eskMn4t6RLjAB7txC/0baHZtovK4fgQ+bbrSZuCJ1Oq8z3Yjc
y94C1LqnGs8TSAcjoyj0x8xd7Fw6F1Vg7RLp9ypxKluK424AIy5cVSitEHQFiubTnI893pCDIPBE
fI44JNx1gkz0NnIkj/b7i6HYEGOpz55Ee/IEfk3fvd8RBU/2aAMutPZyqyCao++D9j7dylLlQGHx
omHUwgVmjhMk8UpECn3CkEDDKN5xPLW3T/NK/p4LxUFqZZiC80/FC1Qeu8uNbpgDxRyw/uQgSONf
ShPpVKmRq9tg/IJTNjhspi8jHdESJpMgylWY7kMKBLTeaohSAM0kJZaRec5dLKlVlfyQdeU5Dscn
fhn67gjer+V1QPkzKTFp1yI332nF9RkUNgUlvzNrl2CARZG9xMni5C8UW9bSwAczHt+zvbzSanDI
1ENqraTgkTEl9O+0ZinlSCxIsLKQhadAu3pYXHGCZiadKcydddMNXaD1IgpRd6BJIhmmiJHVG7w0
gFe8b5wr1Y3z0Nbk3tk/TOawJpGmA2pDTSiS+eKKb5EMU9nqqV3mc7GEL/k+IfdzCTpJGECmLbOZ
KiZC50bS56lKnUa7SRaQBdaD2eFJQY4j+Feh6KS/lB99UH9LkqInqZ5fu/19N3S9Ox+Zn6BwzF2u
cy0U/53PcAmP/gzKwghVp3GARP8rSPZom278/RDqn6kHrnJBrzjLm/gT1Pq2KaNd3tcVPUNZmDLr
H+xzn6cxNfufGGTebjPuzKHd+Hak6HMNOV6winPKRyxKb5A3gNvUfG17nTm7krE3GBGYQa6j1GlC
cHcPsWaZzYIjUrfb6ct82qDsRMjwsJI/O6/+SnEMswFlCTQnh6IsWoojEvXTYB9m7NB9fcL/TIHo
TID7f+Hm/6z4+hIkGsNfCetgh6D6i556Eg7Ae1pLwpfa8IQdk76g9mGkvkX+42FM/p7PCd9gThI5
K1fIY7Yz8JfSgx1AduMQ0cO7k9MyCii7tzE3AER8sZ8C1rmqrGm0Ww4w5gKviQtWzgKdeUXyUdvw
Q0YRVHD0iu/DM9Tel1ts1TI01yd9Njx/BDJceFEpFxErOMI85TeCYDpscg2md2m4UV6t5UXBv5gB
3JcQNL9re+hiMGgIXYRUiXKVvAQDpw4zY7xLKJuuz98VT+9IJa2elO8JFwpu3O1tYWAKnvdwCCH9
fuk1elSgLRCUULb66+ejlI15KlXLvLoF9Th62HyrUHIKWC6Bbg9Y55IuBRlXT+S5/df3NMhcrRaE
dfN9z6kiAJRUTT6mPHL3MFlKqKU4NGA+/pScgPGTwiTOyVfrG6WvgM9ccvmqokgCudOAh1dqhXa1
a+IjHb8LizMa+o+IlEjFR/ddqnjG3FG40B67fwzFCEu/sTuia9JwAjC5K2CcF5/AENOf5lpiyHaC
YoDL7S1zYAnwG/q/Q8oWV2y7Z6ns9CGm7v/4mHwRnXJMU28ZoY0s7lSVePl+4Tx6SE+DRx9khBi1
4MxWGq6eI871ax4+EzPyqFfZw4lgHfPd/ihfPc+gC1LXNMovvEDC4GL6EL2j9HRsaA+gTwGgKASB
Nabm21uspQIDdbNKFbKM1UCgLmTYi9T6b/GOK4bpWy3eZcIwFY4kTfFIfoj6ALV9/U5REsV8XA0+
+O0F5S1D94MAe1N1JFSZF3+tKoDkz51xsGGR3/VHsiC1/Jvk0TY4wvsPrFA4UUHgO1mvKClh12Pe
S3u9Sp0o+LsDYdH/7nJWvef1cZ277BDHXdXpfKnfLc4v24zn+wKRVb06k6UHtu3Vz+LQhoUrcVkq
9/PCuP8vvp9yx4P4W34JwlFK2s+s5PriuROMSV2+bxLKC7vVzijCwOfSwjtau27pz4Tnkf46MlgT
1bSVzBOjm+CMsQEdNFsPZ9c63XwJNhpw6S1jDxwJ1xGhli6kF3rp/b+bfyVowDFSxPC10dPB8iXD
1CLGH4hXJJ0K1U8ia6Vs1UH0YYARsvBsS+IFTY5yYvz/YDhFEIe6phBfWsisLWIa18C/xQTk+OmU
N+Xqi4uybKcSNgAmG+S9qt7NN7OBMHtofX0ydukYxbZ410SBbZsoxhzaduHf2eeQBlCO8laqdeBr
lEMjfx9s9JASi9ekYPlsxKrcOj6d18s00gYE2ZP8lpRpkRu6KvvHhu2x+lWtAC6POuUcyYwxNbjc
vyMO/hbD2+akdkewPgTxZhniwvvi4Yc2SLmJ3SYrOhmRz+5eQvt/EqzPjsPIzMr0FwW0L9W2JG7v
MZdXwYaV+6RmGklXJ3SAEmgKid20eYo1xGX0gw55+5i1mXN2z+oZE746AcYY8jUaUXU20/pxyzE5
tIqZwglx/Hm+tWsXLVpADe4obzJOehhwL19MgHoFW2cqhr7RVcdBOvXEYTSN7bomuRLSi5lmxAVz
Z9k2FII9251r0upWcWmjYWRkDyUCsGmZtlQ9qdQIJEOYf7sepgoA87/T7ysPNqTbCGghjoq+4+M3
ti8T1fDYAKM5I+jDw7Ocd16Kjv8yM+nQsa8M2WYpbf4MS8zwXUtuQ4zTYSom0Qe1QCoXr8X9a3Xx
Q9m2Eti17UmDl8+MOtXkPtz0MjyFGGGS8pb6vgDuii9UpV3g1x/FMEOnxtF7C1iDl0DupBsoLRac
2U6BmluSY1a1N9bpF/KXO6imLfDbfqXvndOX/aQQX0gWZFKYMC+4M99gSwFz5WZFY+AhNqs9DTGd
fFHEh+YZC6FgIUFaqjSE3qB+8eVYRt4rw/KmZpwLIjjBc2xaVkJZ15BNFz93BjX+qNIdct8SCLIJ
Gw2W36pZ7qyGjRx0NZgSfme7l16+XF+WMtZvuBtBUxa+M4mYyLUfye+ahdzxR2r4HddKgqUkD/Hj
cyf4zfYeJ5702AsznP31EyuWHHScAPm1IB6RBSzDq/grBlfqZ32TDa7Wp8XBAbiWHH/u/b++Kw3c
W8exx7mkojBfvCGKHl/4usn60gVfe4jEhOWCwOZOUoBWEXNrfD9jXqI4SR5c5H2HzkprVaF22lnI
CiGE+ZFbailI9/w83l5SAYKZ2YkkqF5uTilX+zWKnajuDPJJQpZ0evvU11TQqtvbG6rFlhihCUAb
Nx8iu6znDNQvOi9FFUFW12nLw++M65ky15ozRUipCnEpmiD5uwou2Mkj4dmuTP6C6xeb5iyrsYqb
HJRBa+CGosSFx+MrusJsOIwNDT4EYhjxqs4TtnA5GIoxoQmwQRKmYJJb1m69PkPhbPfn1KncodfA
YuOgAj1Xj5jo3h5CLb2/FE6Rhk25tRPsHR7QsVp7az1Wzt9hV/QeL0/sw9UfGLoO1aprnPXhWMHl
z1iKhZXKbBsPl7tSkR/LgDC2Kn+tvl+5PUXTWPXv/qWhcLvNKT41yIErQFWYdeGpsRdJkVerWyKJ
tzS8tewZyxInYoc+Xbe3hIOCj6nwUn+ZG24J9mYiC5x3eD1kG1vPyxLq2YqBYKwQFoaFEuJoXC1j
lMwAKK3yxSzsNkyE/1SVtcAtlk3LsKwkB0kMp4T0RlARgBGJa2Wlu4tNCA2A7KAm46DvahEfVO49
BMi+YBXjkMz0N9kRr/0PNxhy31eL7O7kqD+5hz4JkoP+KqqIV+O4Lup6vDQyWTy2iDs8fp7VmGnT
HNKJP0kwrhNNS+2vzYhVIl7L/7eqrgZhqBcNYPR+2dcxyPuxoCBU4XjtxouCKeuc2C5Td75kJdt0
7EqbBtOaIWNZUa7gN8zbhTujoC8dQQuVysRRrzhf6HlljZ6O4rhbCihjczhmKCFCozX+hC6X+Kx5
SwJl6qRWvZR+VqymZoW66SEXkapU1aUtiV5f3MXf7bia/EhNrVrxaweWcYRSACS+WKXQ78bSnxxp
wFFvThpBn48QOHKc+ZOv82hOwbk3PnMRH8u3kXz2/LApjHiiFnprw2JGjpuEyTpg9sla+u/jItRt
JqO6tRYpnl8u//G4+ZGA4lvSTOS2ZxVq06e+/MJ0qHNSXNk32knVAR5aBcNDjrWpzAXpMWLrFH2N
8t0Qj4PcH9IHZFshW6qCIuzkV3A4lqQ3oEzxP6VSwRPgDUmM/PdMk+tknR6Os5Hvz+KFUScTl6Qf
9bW1JmOYaN0VYM4RoBfMLWpA3AfcpvSRyrIm7r7ga1oSSpuZlOEkwOJjrutiL9XU+RH1OM4Ty+vo
pKipzP2PW+FCZyFhil5ejCHn35kHiDVehrq9v1nbuOPZ02L+T0kdct9ywo4MkAXIW/HKV1Y40VuQ
DiKtQy6BGZYoP3uTsJU8DurcA1IqOc471CKLrmWNBYqYmsa4RfZJsTpo/a8k6QepZGoSw7GT1l6T
hOZs85c88tOpw4iCKiSd+ueQZ88cmmVqFWmn+yZZd0/hUtHmz8ORrt2Xsd+htXTvuYp9d2Ocvl/f
SnunzymPGpLRCjILBnfXCEWu17hBccW9lyfD3cbzPO7uSImj+T9Jc1mMJg0fPGegIeoMUVkYWBW/
lsF6e6q7hrWJa0oXl0mmuxED4alfT3OdVGQd+S4BJFt0I2WWSTJwtjTzC7mRe9qlk6hNdluz2T0r
4N7kuZ2yLHcyxqgPLyYKxAvEGNRhbiNlWzRmb/bHrf2zowfxdWA3E2BCORyLSWAVefZQtBmQxPNf
lcnhkP3JkCim3XGhytR0dO4CBwJOXlMEtja8d9iF7D+YIea/8SlNE9/Td3wlrRQ4Ohb2LAvhElq4
7ku7e7SPygeDW6268RFfq/3mtXznhb0mBVc68jI+zZ/cmEFivIjtrKhTspdOlATe5Vj818QalcNt
Lcjs1uax1VjwDZ0OYqbkd+0rsKdBm1Eai7etugaOt0gLQW6ML/BNbjzja0DUidRHUbyT1uw+XbVV
z/WOm0ad1F9vb6/++6PnPFJWv+9/E8dIVmATuYZ8/aUK29j7cirmR/ENLTMGjhvTjamgn+rk5FIk
GtMpjCy+obNjGqdk+Ws4JVeW+egmBNo+npNDffL8TSks7oerbEAnBTrXrsyAiInkNT+SXg2bRO1R
OD/p6032Wb2wsHCsqCYzVPjQvkfs/8X/I0U8Ab5O+BVedjAi8aYwepO+IvpViJqipF6sLyRhzTSp
UT5cLRYB3d0oTPAbsPeSpirwSqFyE7XhTJisletoE7gR9clt7wMRSOiZd/UI+Z6Zhj1ukTj4jJyE
ge1037J8vN1VYkIeFXeidkyPzqM2nwjYIfDr3n025M7pKqlyXw99z33IA7GDD9FmNMwc4ecXFV5K
N4WOddQPyTbSa5yNCppItOpt6uvIlWFD623kwvNbT1wk8bBAewq+QeQ6QGiDx13OqzeV5hAYGLwy
CNEVyBAERd4ZRDswARFxeQ+MKoaFTWp8WM5UIAJnULgQJ9RZVKYv/R7iYE0LfX3G/wC8dICneUCU
XxBsO7V/DB1O1VYujcvCdrmcdb6kZ5lxPp9dSywGxk2NwcYwlgEuz6jGs6tM2b7Uh62lNWqj6qs+
uf6PL4j3EuDaWASR6LPWQ67I1z+aLgmwNuFzst01EFwHbrFjvgbNdOGCo8gIJZERTcBQh6pjtbDl
aNfuMO5kJZ1p3ndd2hWDot3oTUYzuiA9boklBT3B4zBVXfoBeFj3Ir9ctZSXZF4nEXqB11u+YUaJ
uIre9BYS6tHRv9HuInxzyxas9nLAo2lb/WfRAdlUK0TbQQDVTZ5XugDBxoLZlNIz4E0vqYXhFpgG
hXCqFcaJ/9UZOOrGDQmU9WAqEvXquZHffgWjJzmq+WERXaxiMm75jtSJSxkv41c2LcsrfaIwrT2x
8gtFX6DPZuxFSbDb81emH61YvVcCdhs3xRSYYjiNpiabhG5bpD1qWkljR/NwVrYEqUkizVmqOG0v
hSKZXZ2bew9isrCLuMhtkTWcbEeNYInhVsx/E9mZpgIzQGqxS8mLw0tMR7F4ShBrgxI09lWHqpLs
ZHBlkKU5/uy+LtlMYcJSMXHO67JbDFF9S527AqPKY1wT7Fez5b+vTidzUg1e6aoWUd/Babg2tJ3Q
VqlJKvc0LjJP+4oU0IRdXCr4U1Q5e9yBWGUWL3U+NeQqGU362TGIihn40MQAvNXDvKBX0jzFlIB7
jjGxxTewFFppOyhWQwn3vYSTPQ2mwBw/+q+X6IwxGlxdPWiMrP1NWOFAp0UKIhQIdnppc/AI2sW2
3N+ICiRifbPl3I4/DrLA16kqUexvYjvnSqZOUiSA+onVNFmqY9Qy/8NJCyeNlACYpur+5wg5r/pa
tgIEtJG2AJBgWculu1bLeoJDFULvVyFROESxyGMCjJ0z1NokPK60IrR5lh90xlNHjPg/3b3OtNPS
/wKCxNHIA/2TDAHKh31SEJv5PHlV9XpMZBqHkduTa4TzGS7AAT5PmDZRoGQQnbAcCG5oR3aGMhUS
l3ztMqZAngiX+1p5mD7aiW7iDq85EQK+gLCWKsgLtYMBjaIgco/bL0KMFcFcUvGDh/dO9NS4Jd60
HLbZ+ruY/dVwTK3H8UY32BjD290VY8j2FOHKoV16hP+6jB0WMyUnUTT5lajd3FrlY9kpuPic2tce
2vJgAqY155QWYp851gyNxvFJRzouZOSeehSfEKr/hKtyyV1EfWzlnyv9cLqf2whcjICKIxC7VLuk
Q/MBRMXy/LhDt0ZB7Zzg/PiERkALFv3Sndfkmls4CaRfSEpaMqXvRXwpEU1tkReZjaXEN+89I03L
7bDLguSQoa7FTmClonyxuEGl9KWpLdRwwUH+Y7xi0erWezRW+ir/blcKMqUcCT8n/0X39veusN1c
NvE4oEsoDnol9p1rzSG+viq5dSsZNz74iz6QMG4g7KSVkLYi3ESPePE5KGdYG5BJ3dZCUKYsZDWx
WKjL2LACOLdPKQWBDdAAm/JlL7VEnzZEKOE/2RCETRfFYOyFP5LcKU8J3peP7QUZxwCCyijimDMC
TXEwbNslLbat4uXQiI1J/d9s8t0vEQxb2pboWNBduKVnzl5ki1/xofBSIH1j1+wZMWVzz8VlKdw6
FH6b0FKF05u0b3sCrUmqxk+NEH0uLGRRXyLfsbTSqUMeC75CLRI53fTbj9pzqG31ecyP/4PGhZXs
1OSTaEIK0wYOy4z89CmhdaSow8vRacEAo3cCgOScxc1Q6bJAfNbvI6LgoJW8I47I4vpVIz6ElNW/
9YL7bSRQOE/bWI1KljSRfXuJ0hL3EWG5opoFzk4jvxdleWEiMqY5+y39VAYbSt6dj7bQ+XJ+Ooed
YCrSEy1Oaw6QC9kCFp36IKzL44f/OZGXiGrY6oBMCshYgX2S8HIoYkE0Psrk5k/FDRAm/tf+/pYN
g7pzurQ47MR7/i4RCO0AZJgfjxB0F/J1SmSta3sspULXVLHp9oEK4g4Qjrns9wwDGTMn1N1czyif
xDPYoPm9PLj4v3x037yfdBJH49C77UCthfTu/GJShYZJncKU2pXRrEojKHoZ4pAFtBgpWIoJVo4e
4Vgv06YDthhXGeq24//MNPZR7LR3huFLEcVXGXAmo6cXPyUE2HQNAL8ePXWrPGYrrCL2zICUnKCk
otLAD0BoY5CaBOXL6B+uJz3pqAAnxsABlDePPhvijY1H0BR032jmjtx0zbyFuj7/iTAaWDlkceGg
tx8wjrx1tdx1jsfczKu6A4WyELJhiJro9XpvkhuigZ/sQE9be9Lm5FiJqv0y1ug6jTkZzsfjqIbq
8geLPsqeBXzgChYNzT53tlQfFphfJ5dnXRWD+ugm9Cq/mKEQEylRO+pI6N4pEECKU3ucD+4jgWnV
X+GKlINs2d6xvgD/160HEW+rM0lcpgXzDMsp5c7lEGXIVHSeS2jPLWrvg7z/J6vJhVZkNP7w389O
PhaHujaBrkPMGlGOSspJzc4wf87SMMyhErRofRr06cyyYsKuIrNgKrR7Bs/b9lEheEfqQ3eoao3M
PoIakuFPdLOdUhJF1HWE7fEm/WFUeGru9gELd4tBsA04ogHSGEc5HPEIGRzb0HbQQeZQkCzu07lP
w6tfO62tW2jf0nqRYoTZuakXOLrE7eVlOPTQsc75u1+7kouwFJJw0vTNVn0B/xaseU/wCpZQ6+oe
ajXoQdkCM86OOvRG7ghxkXVlvuEsTgqEODaW6ySjCYXHy4eNRHqG6qWvMPnPcNxtgV8Fc0RKP69O
9SJLRXeTq5KhgPfy1HZXYRsU3DSMEToa06V/ntJ2XQltS4EW/jIwtSnIdk1NrudteT+7RRCm3TIj
L1ZF2vmeS+3SsWLYYOZMeQziIa/RZuFsRSI0zQMGHiF9rgeckfeM7rySGGcLV68nnJm8QDg7hKNZ
fNtPVDM+ZcN5P3R+a3AL4h6pUdgkCTPTMW0FULZsNJTfZJwicI+1u4Z4sad4ZgRhgU9DSgvBreUO
EH7kZKDKSL3JpBDCYRkwjrIrFRCWV6zpYjy3KkylKhikGCPLTE66UCGyiFM/8GM+SGJYdTDOWJqB
XVYxjgp2zKHS1GUz5uTIPZZAnX9bSRfYSodTpHsiz1OThUn89YRW277/DD6dh74vzRtbgYnDRWDQ
z+fEPi9OT0yazlOQoFH9CbC7VOGmBOPNLZCuNMW1LwUUZt7/JLu1IOALNJIm9d2VxMaYfrX9XGfc
rxMBvqsHlIbpZWWTlD8Wi3yE+eKstbC1CWDQgiSqKbeFBqKXaADVOzv6Csd+FfD4L+GaMj6cI0et
GW49FWhbfnlg99ePQ5RbyoCkhINwvaUQ5ErV/j67rVbKLVXrLGNmwjwfecF4PphyjceCkY5L0lQc
rar4MbzEU/Ey/cTIvLfjj95ogedbmBwyu1KARy9FYykvTLT1t6hJDVPywt2gJ1ugedjaB4hJnZVS
ImMec0AMtQtT/r9KkSfP4YtgEZjkbjOOQWbg7sj5J+jQYuEBOjwqLx+RCG5JJFbo68FDDXFPi21J
LSG4ADnzfVNX6uZ8cTLlquEpfwVFqdSTI/2hJrZMzCkSZyQyVj52mE/WElrahAsmpr3GtT62JTcj
75trGXirjyzb+dGmGVCB8aIqu6IOom98NQ4MpvY7tkXzaQNYCcE+nw5G8iGoWPC/+m6aHpCIKc8E
rilKS1ZOIfqfQdRN7Q7BPRbHNflWrlSoamlmPk5Og0DQuoQHfKoFI8EL6e55Uuz+1s5AiVl26mZD
AcihXwlf4RoFG+PHDkYxnqDYTMUxCrnxgRfatDSCvfFcKc4asCgkK/43QE8wcALNvBSe8y57r6Ul
1HpEfvL3xuUuJlw5rH6fhgPRNWfAQnc1iRuapb9gUKG8P6GmddkyJOka1wK9EjfwY51+14wdLr2W
KHfFsJB1HvHAV5GX2UBcl+RVvMN3GvnEORzrzBOdU2dC+ZuzLP7Erbf5xpT1tZ0ztorf6g3vaIs/
q9oZSaXIkJskIRdlhEMO8N+qRY6bnHSm5TMjul9D6GwarypxfR97kCoRlOjRrp6s/nBmwkshd/er
m+HTykAmN9RzcnhLD8qZ7GkcJ1WSoCRNjfQEElwdG5B7rtc41PoPk4QM9VpbmllZZ/qDt0fq/rLV
gDOJm8SrSJjZIQ6Giax0YxPV9t3F4NEQGpNObE6LqofSy749cc8HFCpJKwpFqscY6nyXj+gPRu7b
xGDhKHhDkABaajCLhQkv/xakGl5bjYi5wEe1rAN+8nmmE8SIjO9GcAvz8SOtBGQa0jJYWsLSmtBf
WcQTUJ9iGqskOPW6lcjUtxkdGbt09+p43IeQNxnYacMXRGEf8EfYr/W/b6qF6uPgk0yehS65QGVI
0O0RownTKoVMgBXwQmf9BrK2MBmZJlMjb7KZdtZX6dLEJA0SiJJHGCDg+V4fSQEDnFW/whGGGAgv
aZ+0GYkfiWXXV+5GU4RjsfKkBV7AA2znPRMQUC2f7GoXurCwyQ9HGtUVpSxo6IMCqaY/YwZn8MKd
QddRvOZxQf1+ys85IhKEDWxYnowGvAZ3tT7iTcpmLT2AYVZfRle0gq02wT9b61l0DwhsQWrmxWdR
YDp3WJIJhztjF7X3M8HIHG4BYYeJmODDMJD1sUrjxKk32TcuHrY2WxUmXmtNcWfu6bPN57x17bfX
uURVspYfspKmrcE6IgsVuP5vRfeXk1aBhxWGIzYpXUSzcTFAkmcQkNOEnlNIViPwJXMlS7k+21bN
oy+V+bJIfbRg9k1Gwjvv1ttGRdBJOWdXA/Wx7bfLXZC9l0ve0NFBCGBsbjYph+tOOWsXRdvXnFEW
FGeGJoMfrrO0rkNEr06XG3AleWv7YaHGpw2aMPX0y7LoxRLmIJfirjotSmt7kDf/iRu0Q4RdP7NB
d9pXM0XGlD39fZ+mu7N6veQsgxoLKcAaBCdia5zGn4EGj2qHyyWR/FgM2beWeDKBESeQC7r4hmCW
IWmDWQAA79gzKsYytvkED+tj8voDX78eud9ffQlTYVagTaMLf+CXP75VwEildHVz1TyobvZDY7jw
F/8OVjMWfg+YGO9/Db5S+fEz1cNWBw7oE4cCkBSooS0eEmz/8UQa2KSFMYO0Dnozxj4p80yt6Q5x
+9rmpNbMKWQ4EV6CrEM43Dx9sBDh1iPM2F2NrmTzK7/dmIc53bdc8Con8ImpnvZAmWifWnzy4vTh
fXgQabeQu996aHOLjgvYgvJW/jlYc3QV21Egw+Y6siUtU2/0yW8P0V0uNQvsi8kcjVzK8T2+xwZH
H6b1VtbQzvH35IH/CrUMRkRzOFR1Z+eQTSvhk2lZT2BVDKl9fJRifhx2LrHLHFJKKpepVJVWX5fX
DwIHLDsV6wUFwUa1hhyiYMUYbDS7Oq96Dsy0Pdh3ye0DZw+QDludNhcwP/eyVVatok7TJdyP5jzP
Bp6lnySxoEkADOYfikBXYXRckUf6Wf7za+Q9wSOd8uqryaN2/KruYkl8g7g/IIKUQEg/Gsh+5Z59
kyuYFXDFnQIJrMe3Pma3lj5cuRKBEUzANkgG0gkpp7rIWeF0wk3cFc2h5yOpMGVUQRL7vPDSdEFs
SyGN/Lqm1/bon4bPuVZ++9b3dkDs8DYGgFZsLAbuXWyaiTzrJKqVkJUi+GWd/vt5f9O2/UxYm5Sa
sfj71MgUcYJrcJ6CZA4/9s4hFa9WvJpNmDoejCCAQ1QBbckLSNi6XqqJ7pYXrP6Jw3PA+lZ0ui3s
sX8bkCkUrH1F041QS4tPvofgGqqnyY2lN2D9LBDR9+e70wrSV/Jw7p2JHcyKwSnibPw5Iee7ygkm
b/mVYZT4YyTqkOiGTKJTsjDMlUk/wp97y+OgYbOsxC2MwE94bXNkeqDA6HmHZfgmQp0wK+bkEFIb
gc/LwWbTO7SMVLsDLbjhTnijXtiUyYQdEvFvJ2WQUnnFrdR+s3OpT85jwbd8C0bZzmGFThKz4n2K
Dq0NpIvyHB9sTeEvRVtnW0Vusl5y90KtEfe/k229/UMnOIrqHzwuAx3SYlMTyR7OEyGXBrMu3H+J
8TG+w7DRPKMzMB5//lU8V+I3Rpeds3dOPjzj5lT2t/MjQhCfX7RXGaz1vTeBl1W91BQpRKy3ckO3
buQK6XZE1IeXzKTOFm+q93JJ+ji5rUCOtsSgTmAGEvEH0ReoF1w/p4RkHLRcAfkGHON+uP6zcme9
97Kg43Qs6tBIyrhy5s1QducIwPSM1ez21fve73UuEMJh7nDDGxCNAJUz/2lzsyRMMHklW1GQ4Il8
N0w8ZdIa9igXSUvtVL9w13J2VIzb7453hdHl3/j6edeeU+jhsqZjjnY6a9hhffY+aapYt+zwtgcL
PGNQYjKe9Oj3dc9rIg2Ji1cHz7u9ht1GPnbacOTmJ+YsFKWKpAxH/iuvr9teE/3K+wl7pSvkTPAs
AGEl7M8s+lee/BDv5QygDsfgB2EnRctwe3ONKQ0FR/1d3ieP46Z1y7AjEL4jxIf/Hm7oz+gYAtzw
/hji5RxeTq8FN/5B0nkw9k7TXK2XK6kU6goS7UO2WHrXb1MUlZLb+W2xSAoFJKpfTPcl0U1FPiPp
WLbfhoCwjU/Q4ayFJsnGcPMS/BBIwBUcWGukYa9m7bjRdnrLf16PYFuBAOHb5QWtcJkwGGHb8/r6
mvcrKydqz1ELcRRapY48ixB0yWbO2dAnWM1Qn39g72nu+HEya38BCyHR68e97Rg6ZF5LjsntYY2B
9iam/c1Dh5xoWNbADq74excYbDmEtaI/Xlts0GGOd3rLRPE4OTONnB2uJ/3hxwIEEjsL9+09MatW
azN4H1FsHzWCtFCKuF8GneDo/0Jljx4QrRSedqaZXGomb1+52lUxYqDIzm7kzk7Bag9SoQuuHc6H
gurtzqp+pSUIfAqkquOm4FllO9g8BzW8Z9WKwVzL5vRUX5EFftn3rgza2FGWt53CWzwxWlLB6HLy
CMKDxblyvL9PNmXtj7LzUcFx+FFh/yO1S0FBa4JH0XDTm7VtTLY7/+6A2gtgctld5JiFWbnnls5x
Md9Yudy6dqfclq5dWmfykUcAELQCgkTpsBQNrQpQswJqpSpLu6SFvZmH6bix0DX/+zn2YmEMz/lo
QcAnLeOpSTi/Z+Eqcgv22Ms+k9uHuMcCWMxDvceMeq4NphHaLGtylMF3e/4rH8WgjEmqykWoyYte
2NYbVRTQxF7ZHCgcIQgw0vlKC0Ndavz3c9y/rmwHSTd3v1LKCoCpW2wttzlUuOMMj5vWq77M7jTz
aytLppefQR6nIbscrRV7VSqiF60RbJEvgD4Dhi2ocbj7p69Hv1QP2e+f1T8FZi8jaD+PzZRORSb3
+UFHT4wr9envNfLSN1EkiIXOSNnWS7eFQHoixWsqraUjdtOo5/xS0bT3AxYd7rEPimEkOZNxD7eQ
qyEYz32oa9JMdC+C3OTDWMA6d1JhsOTKmsxmwYJ4eBS6GTxd3gqhKpgFq0FJ57hs5t5e+cCY0+JN
UEBEq0yqOY0kncbFE+p390hG0V+m0wP5J+kk2A6ySlN6WfCCHiaiJByJDXH7Q/34ieoYX7nSBL/H
cejoByesZ5NdHmwLXHTAriVFmgzTBhCrbLb0vfZoEFZVBzRL6W8m66xJijb/A7TaS+PfOchayUr2
oO+bnlt3nkD6TB8THHHtyjdEkgPmYmAl+0LYb1kXZw2KAxpNR0NTiUQB+xjkRLKLzv2FIP7sR2St
OYXK3JxpBOoK3TEjA8MwqshlI1N0GWURiV6C1fTFNIykIL9uunU2/tx2Eas4pBieq9xA0Y2PaQwC
FEkgWzCcbgDVJxqqEt5z5wS2PFT77epGL5GcV6qIjBU8UfPr3e2x9YdEAd/fAasgbFCfjW8G626k
f/gDGk1sIdsJC0o7+WH1gONaqOOGTqz7LOEa7ng5qhG1hjoUKj723vJtpy+Yp0+hjb79JToO5VR/
6NajtrOuC2xu/PPWCURkC0iDoIthHfztRkVUma15yH1KfjoyHX8DssBDP7ejMUB6eZ5RLM7TFez+
2b12Ts7Sb8eJuSaHj4unmQco5oOwQu/SGnwNX3vGu0qPxusvONkxVIdwyjLsjAZ0Ux7/oFs/7Ksc
h7hrqKVjSYWxMeSi53ZOeT6HjYif4vWhYNZB4bX8pjyr4US6F1z8JjtncjfWLwBeGQkfpxMLL0nY
1wl0Tq+40XELO/dz1G555lL3QAn+lNpPfdFkc7sdae+ZuBwse5aHVQq6jiL9EL5darIPXJ/bXb67
1ErNFIryoaSCN5nxz35506Q4W8gtDbs2cn4asqEwTrYSln/8B1dF5gZCMRFQjjm/sRYdS0DnK4Oz
2Iuzi9R6yqzBTBVafuZJUT80jps/ymyhZB08p5DPqtTswIFPboF8Q1b6TcYFz0DD3k6JQDtefMwk
+/nDekbLrLjD0aMXbZsrENhmrd5bVBgAfNTFPkQOpE2uxjKLxFkoZn99yxgZDpLnsZ87G6meEwY0
y8ivMqpzlr3xHgA/37/OCdvxlTOyDgUcZLo988EH11qfLT17PbpQ3zO51rgiTUXNHq1SMbu/Jugu
LfysRv52qbcStaFxyuVQ5Ff6eEDkkt03jmcbGcCwoVFa2ioYblIausqNgUZyySM+wS+6eMpcbBrF
DaRjOZPECe/9BmekFCT6jXXYOnBu5ropu00t1z+Sohj2SYe0EGnBoxAXgzudiGlz9Xy/qwUZIu3n
mNqc9LAOOFL4i9sX/F4PGyQxaFQvDl+gS8mnMyyc9raYMFIzs/5aqkmiMjBCGiM6owUHFvy6GYBZ
G7Z9XNZBCiQYceYK7umfES5Gj2EeCtrG4U1IjXkGcN3Ma9/54ww2yyAnKBWbQRp+bUyhFydtCpGQ
RvDKE7aygqhuR4pI+FsQ8e5CTIIpSWBhsGnkpT9+q/ylgpJbKoylL/DLQcjQqmayaR3N/EHqYG3G
ia1wJKizA/U4Ekp4YhH19DtnJtNRWJw+1xAAsYjH4jn5BTFU+VKy6GhzDbJqzkqBMkFZ1FhXtQNe
9ilhCx+UqufyDlztX8UxCP4lFetOYSUPl0ynmAKbhvlBCNA9aU49LlagSINAXQjMlABC98ORETBc
hdnCpq01qFMkQpJywZprL8OQS4UsktVwSLMk6JZ71/FVjDzN2spQsdEIQFjeQkUBjoMsYumCaClL
OQJqAL6DbONx7U7kLMsxJrHWkh2sDbgFo44NdT5KdpkQPT0ngU4VNScNxuFKfGUpjtDdOC88Yc+j
OVi/XyQvpw2zu7pLYpozwgYY/L1X5VSeHdoAIcbf4PBMLlerwEQwDffwS5aSiqRUOUsKpCNlXM+Y
cna0czifM+w6vxw4nAEmsCQuF6jA8yTb7WPj12k9gdGQ2InZ8MKL6QgME25a4oPeiNFDXqgh3cRL
wUVQ1KfhCKDI9edKjSXsnkdkajy8Kkn5yWZ6PPP8OreDBwwRPdfxeC+yujqZMBICGAAq2NtksAcK
zl8zaOTtvdbXSBO+oVq0lOqvchPBKmMjm68bYQudzA5xud8zepXO0HBexpbAu3nuAKbHUOfL6PbB
uG1endU4mr6sVV2bG7GLMN302wh9qN58r+ybaRW7T5EXg9JID2w7POYVX3U1Q3GhPMQjUgD2fPYY
dG1PGtxbVoSpXLh3yokbWT6FxZzkCu1c5ZawtErN2WTMJ9QgPQ54KdKbzaLFoTHy4NolB1lotCXY
gvHHllxZu6fNQEKRB7FRZxf9LuzjXTVH9bMDJAxikGi7jtQMMxksKrmjve8T1kLvXLo8XMXd+Fnb
QgA+zHv+diA948kx5JWdt4QUUCFjhpHhid9xRqVls2I2GfacAMVL2EKzPIfL0UnT+hdF2YRxnp4N
wKGym8j/HFS9fN9CrEXzRvZ0CL+HDfVjZf36t/5TyRKReTuvF81OcyQEMlMBGW1NrCuPdnmJzqoc
tf51dkbS6cyvUlXwdj25tWVnlPnpmT74pdY0LTnemdIk6ieKMgDUtdyZIQRax32cMFilNSsa1/fy
hyDhrpnqgAmASjQTPkHMAPDIceC7rrYLB9fRVV/pTaPSWfwT/FXsrbvwPGT/6v79XED9FxjXdZix
nSt+ZNBCmQLH1zljmTIiZDJ9PDqhXwXp+czCa71EBxZKxK0o9czeC6b26NOGXyGcEuXCmaUAoUh4
lmFi6pYtfSkiyj/2dN6SmzBuYvJbEzatvzxRCieHy8xq4WhUrMZVD+E3zJ0d8iwMxIZ+VrMFqpWE
gCz6BgJzMx3xtpZ0+6CHhsm9xehNF7U2qIqlq6DBjbp1TXGOD0EZ5nXyLBIY/2Yx22XKSvCXYNL7
IerxlbfNMsuXLTvh8BvP/AI2XbiGXThR9i88dHyO/b99YbxNz6dWTEX0RS9phePBBz1vuV80Zp9Y
lga74CXIMxESsJwdBU22b7ocPPtbjaTFi5UKjlWJxJ4YV/Fx96CaGFi2TGTNm/fUIF/38+D90FAo
hf5R6aZQpGHnf/lYoFOsPaJdmn666Ouf5cApO1IdFSbFe9z6FgpArOkS88A4pPYZgqcDb4VzEAEm
1VtFC8dFfVeaGVIo6+A4jKzyCzPMiGf3ozsRiWTVRSiDuvzyVCkip90LO+ygvUmlK8JBwrx8F5Gk
xwVizrHcNf/SUrJq1XIp0TNZzERSq/queYzu9fHW0gsD/+6PmkdfbP+7mR3hoDQIkfdfTFTCKtNc
Zy3iPdwa9q7/zF9eOR5ZSsjzg/DnFFGnXpxSJYZoQ8PD3eTfdFGmi1PN6iK5vGhSA1Kj7iAOlmaP
jNGijCyR8Khm4sf+rjB9cCZyn5X33DlsklKfSFHo5dHZ7FTjSapKWPiojBsCvNff+mG4MFUMlZWC
yTii/jpJFlKToMdGCs6YYijtBSA7kdcKdsaf1GmboOCYCovVy7S3ILihVUzG2JeZBWexKFU8Redz
2AJ8PuhhgMYEAlzlQYP7nBz6qF6KvGLG0q5fxeP2IfdWk4GvtXwudXXr6fEaKBfQjGOdGIpMIGOD
Tx8teS3xvd2McUxQJxJi897PZnmq66KQkNdfXfhcLCjYTJvxedqeOBnTSnFDee3SlXLqhMHc2hbd
v//odj1AzLXDNSXsrc4Pd6SjKq4xwM2NiTKsw2/paFA8I3OnJEZIlrr5JC9IZVK74KVJUKOEcMML
c4P4wDIaMVuK2zCJWTjzgYUitzpYN+8qp31ZTl40tzW8OZx4Avufaqq30dUBfpBL4U7BLq/92rAU
HviGFj4EAr1eLtFeC+ZQDVbZPVODvOm1UTU8maex++faaVcbPdz2VUtANVNflsQYPob2v03/z6Sr
KB2bR/qcS1xporX3BtC+qwsigx4BxL/dv+712O1H309KKRVGgpukagnhwSV6mb5Vzwq22Qh2itvR
DLGyMcX8KUGDa+8OxVuD/bEfYeSvJnzU0z4XA8cmRRfdjRpcuITNLbNc7MCgeWxahxq5Cj2zOfzG
wKXF+k8MWw+R/DJJvedcYlpexNdL5yuxoYIVZt+69HNjAX2pyNKM2vp65cCWxYdmdQt/JY88eX/k
1LJUUECqR5UIrs/qEEwCUyNygumSJaeK1Ep4al93wVb9SmPbAetN3lKyzUPGVdGh7aS7X+ozvJBO
FlIFRUJUSWl6HGTmDaWQS6lfqRiNss1ZDa5NAcIC/bFytJXRQR4oU7WsuP7KhQe0l68LAkyvL8p7
jRG6kvo94GaCU0Fgv11qbBRDbPofJSjGXXFwuK78znM7pJ8zQoRwBcBoDuiI6QvoLEXFgU9PHvnJ
X7bRCErJq6dKdNCm0KPAgaKp/7NcWJ7BtzmTkd1MAqk26F5dAsx+Rp3OLyc6gUZeMx2hOm3Ws5ik
juz4kwJVnjQepAHQ2YI/FrEi+IqdY6g3woYsNIPDyWeJEeF+B1Ny/yiCqDmQlTW+b3jPm1PW2urS
Rbw3TooYgwni9/oqMpimPm/VW2u/1EcLlb9a6zy4EzNkxndGD1nNI77VPcS+tI7jp2e/YX4oD2e9
kWrMgXNMZC+myTDpvrF0wliSxRzDB179QxLsQ/d9Wo0sKW1SQVZ3FcWRKzTHivZnR2+NYB032dj7
yUdNBP/SkW7bKZ6mF/bDrm4z+D3IEzo47kjsO2gKP2V/Pi598ZQMfU39F6sluvXcjw0p5wzU051m
leOZClTUKFdvFtJRsSxQwZN7C1sYUrwtfxs9ihHYcM6mXw2rwEEm1zcPKHVNubZSmqF22tjiKYK9
BKqfvhHE2ZmJJGJkONU+syn/znknuSaoiyfghd8AP500x4DqnrYc3jJa3atQ/ma7ubPvaX2KXtoT
zNflkLMIRVJexHunmS+KgkCm0JzvqNEgYjP/furglhG02tbyAHoH1YeCXWdU9HiW7zNi3wNT4+uw
BDBYKSLNIUYBffOte0WEe5bfXhIUSn8eyEZiXWq1r2Rz398DIAN4ENTZtpZKfM0e0rQi28tOV4aV
z3oWAOfie7m1xRtP5//gt4HOIFrKmBLyWbjDRk5Idh3oCWaqZbPoDli4klH84/OtQ6JbxUi41Hxk
kwPp/VxWNhW1oL9GGllIWzn/cVey8o8rBvjw+s30rKsh4LvBWPY53XJ0BjpMR02Wd7W3svvnWAKJ
SxDYcwX5vRbRyJGlNuVeCBCVdBTwGQ2uoczCMoXmFgeYhgN7EISyvIzfLb2s/t92LcqNeMjsmSQn
vJB8WoOl7X0gBAodnbqTjl9jSg8PxT/V+Vfgz2KYP93T9dsyui62B1u9GsE0/Bmk5dsT5jX81I1L
Wwvj8SspcluxrG/owaBctJfl7E3n1ituwsgYKtxxt+3olJNP6KfJhPlB1i80sm6RrHvnEAXbIHEg
tgFPlGQPXLdHwRQcnAQEmcUlP0jDGysYpMEBDnj7UARUi3ByHbM3tpE8ULzM/wzdw+tTXjown5q8
oLLkZCmYN6FesVQ6rtqp+mj+yCYOXJxOwOIeyfJdZnUvRDGQt4m/TUGWIRyPwRCsOTGJAOjWFfM0
/h5YM1UfaPPprW2GfBbqY3kP307U8m57yhw7zyHeONWo0jKw6NijSkh3Mhf0fLwaewbvUeE9bAFC
7pYQBl2bb//g7P175hbCfSaSYLdSYbVzBSExNgEFlNCGcAtulB+BGWGhlNuFHT6OaMPGyQwHEfbl
3xfSH6Nh9/G1zGcWUJcmaVI+/5ns/uwziTP7MI5bxcaltiLXKuOBGci3ClySt9zyxOBhGUh6avn9
aNt59/xq38FxOfaW12HJ+DqKr3QVTOPWgTqJ1uATCC55uOO5Jse3ff8S0ulRFlb9pV6UX/O4HMSA
6IhCk+wcgojjlIVuv0yicuVHsosFagVYa9FjiHkKPv3GM3a5sl9yE2bfgzpruTMI4/YQwxI0qauZ
5lbt3mqtMdsHtOvSeITjM82PfZKmBOcrQYp41U7imxsrKHWczieO3EGi3La5P3W+OVm4szLIqiQD
6gerykeKXzXYZs+0tOy5F24mBB4XKpUMOwvsFCZ465uXYIwGirB+u9oeTf0pG2SnqK3cj3drHthI
JppvOMQxGRS8DskF+bRC+VzN+mSQeHKY+Hhd6Nl+7y7NGEu+vPmU2N3sj4NiLSpIAykl2ZRR+Di5
EdE6B5IOQkW5E1+7hXZkS9K7yYpVdt2CJS22hZiVmGq4m84auN3Dvi1KXQalLtCd2/zLLJ01tF90
0yoYRxR1UFW1OU5u1Qmz4t0jzVDDPrxynvwTBq+0dTh8vTOl9bQvMb3WZm+GYwwnmWZjwNRoNpS+
sXT4A61QkV9EppPZv6h6MyxykzPqKtqiRCfAZ2YK0yRobtlPUxyo9V+O6kFykIh0wMj9uqWpYwnY
+Vyc/JVBEgYt7Cm/YpmEmcYobCdMT9jSKcYYy/mhAD4S5lezJbbkcT4AZd14mIMXK4hf9G/y2z/6
vHSny9uC/CmkeF+yXs2hQdgeWOa6sdU7p7HqnZ+GySaXAQH2jIlfBzQ0P3il9vEURtUQKpL1rZy6
NV46xOKWHIvheSkmnbrWvGpCr/WToT7GgRjIpvFR3Y7nZh/Yoh868Y4fSoVxjX3KqNXYl0abWBhQ
uwzXZR+kdUQ0oA0oYjvH8LnlfVt08LQ2bNbxZzBG2a21SJm1N3yBkfO+Oqc7L2nV5b3kkTAiuyNW
4H4bF3P8TwCcqV59QqIu/vBbS5miC+/tk6jqEOM94XRKt2WwvAsqwF7YS3ylUzhTx4T8w3r7Ac3f
7h2725BYpYnvEEMTP4MzCzi+6jx9R/LE8csDH0zPPMq3QFNXHLJ6zcKQAwJQt2B07f8xfA1SCZ0A
uy/EDy7WdAwYkkjYPZB4jTZTeAOXmSHdRly7sZE78bQgT0E7TwUSTenQWNYBa3QqYJ7uTfshmYsX
Ds9AdR8OSGB7dHNrGErD94vU3IRcxnJsBo7mTUUO5tBdHPgmeCBr6KmAbg9Uy17HHfBE5CcIbXH3
Hp9Cqnf4VsKGDpaYs34A1ADEx0YFZbvnDUyjYlTbG66RFN4ZdrZH1ivhNSE3tpLCJ14wLpg+OR25
IHNuueV34Q5PqHzrd0AhvOlE0rFEnvH35WLIhpUt+kZ0jlbAV8UuzvjAj1tno0W0YfAzh4z8nK51
8K9r/l4FQILEl6B5kANh0NchZqjRxOKJ4C2A+0/iu8sLsP7c1KTD1AXsJwNuUnp67PvaqvQsyGV0
DQq5kIH0UPDfjN60hjtozYhLB0xyU2JBSNMZSHqWs9XFqkigzMPOkCcZLlkz8V2K0uVfdViZIWF2
JcGYtpFsMQoCau7GSdwa7Ve2MFGk2hgX7MYZ38rzNQWGus0Cg8CdVMALjuP4HRgbmuI2nqsDI8bh
8pIF9XWTVosxj9gI+M9Pde0hrC3vERj+GKZZ5UqLMvisj22Jclak0j+MZYkvAAuBRdVr9550wJHQ
T5F1DkSDaZ0VG+pAm9sM9WNA1yjiZIFl/XREbeAwK3i+TKs58QWSXj+ElX7bOCge981Exes7twh4
/om15ZbOqVP5vCu25wP1QkCldbnnLoXzMXwA5v2+cMB6XZhrrqpr/NINyugMWu3vLwiyXufyctoH
cU4ailBsrOAQnFXVa/IPuJlZ1JWsfoESqXl5CecfLc7LbPLNeOqV4njO8JsmzZALcCsQFInxHeFP
UvcMqVYwexYt21wmj+X7D1Zf99IWWmv1oTi2HwZmvoM7g8wwvc5InOxaoI+SnHOHq/LH8ceB7zG9
AY28GwfJ1ZxWW2IZbCEgGRRpPmWnY9VB9gdZ+YeJhFOMs6lHhKiCTK5G1puBM8K5tKjHr8Ysk2bp
PftvJSYvyixMRIgX3zmnpa3ZE/DxqdCJBBTIHcRnSFYPy3b0/UtdQ42rvqS9f2zVf9KzmCXkm4me
XE/s7o3VHmbWqqT/wbJlwtr7fOrqDnfZElwQ3SDYrznMdkCC4rncFzT17DJm8DpY5N78gWNj84Lq
20GNaabwqLw7IuDPmF71oOHSQ3747noO5Qjs8uPWL5fStzphymkoSEyZZcAFiLAFh94WU/ciCB1U
HTp7Q6DJ3+z28PO5dOn6UJA0w2Kg6oFmGVmsLcbjxn2xbpW+sLopACq9jYK8Ar15kmW64mwFi/Es
Wz7zGAHAcvuaaIIkocMieRSumbst6t7g874yKhg/JMLS8kHqBJ69jAgAT2SE9zagrNgVUmuWylS+
YVYHHMH6WqsBm2M4gNsoIdcZmYQoQzgIqCaGM5e7mb2yqtWXW0eMIRFixKHOit8AKxWheQNQY2Hk
iIEaFmnLFG4ovAWuNKLo4FNjop6gYS1lbMPiGD1Td0q/tlnPoNhdFuUqGyf5yQLV+j+qC2PAali2
OTMSRE26ASq90AWjBkYYGA7/ttYIL5yigmOnhyFEeADExJvMNx5If765EWvCNCZ905jmiD+lGT43
iKrExj/FeP8i719ihJRnqiMLxhp4EQo82vzZyF47QEDJPAmD8rjkezErBpwxiF0kexBm52B71Wt0
BQutfqjlA2tel0oeAVuXv4RZW+IutnkMnx/Cu80EFyrRAwkauXp1ezrYrukWBQiOUN1KMpRH0CqG
SW6E60ZR7BlGURt4pOdEa0FPEX9oqXWj4pYsQe2asNxji6mHycj2sXs18ICWG6e20BzITODjlcUk
U1u91LQ5YGEzIjzhSdw18MPnhGC2MQZAs7YJ+86r8uMWt9H6lr6edmNH4TYd3R06dvTSyS9Vtrkp
Rhdkh1/W8bhMh8sVHbxLYj42rX/iIPRkIN/B0acLqaPyVFXYpoxNHtH8epkLp4QrCam0Vk8Fh80I
WNZbrD2SOvdaRbQ1LUXuCD4keAVabjZBFiwuQLeDzzfOeqUuEY5jblCFHEzHF5PH6Wk5jbcv0Jnh
YnxzUYxn7MCwIrl1tPcLdoBXuUL2AZoeLZymJeZjCOR40cQPo/0M+ZV8TcocfHAf2oPqRhyQoYCX
2P+AEL3XohWVeqERVNmlwP/zLn56NMS/fClGZivy680O2jmdj+S4bTphBfPi7xbMwYQkUKrYFvll
kwKI7YKm8IsLFgoReyLpCzyaLc/BJHkxlsKvRaHHIGzXlZx1/ndGViPgbQokz6j0NRrUaOn4EPWY
ggX0HHmtRWi438IZXzw20zo78HphlITmwbYdeY+EfmhJmqh8Ci5kTE+wHZLn1aFohQ5Z+ClUoLaN
NRkc9LjzhwsSjXTMdtaZfpdkiiDsB5SbtWKpDu8kdrNbPhtmMgYOnPWBFgYoIF/QYW3+29m+NsQZ
ebwESI+oWHt/yyYhl2azHPOf+OqJwg1mTLqt0gKZu6PGzYBB9aryqEPjhUq6TocOGL0CpFbe+kUf
F/JctqqEgL6GUiPA6ViH/4yf4Dxrmq0H+bH+Cq/cmZjfX0O6R/P4GK2CCsDVeTuxpcFS8XrnRyPv
pMwnfWGkPeWnkiA2Vow7eoEXSQdlpshOzJhg9eguP0dd87BPfMl4ycuT3S/id+3fIqHgzqB/hO0h
p2BHssIGQmVCSo0kRNTC6yGd5xWoVadfY9m0fOR+ahNyBD3CinDaw041YS3jH/FKLCD1e4CWPsdT
1E1IEIWie7Z8pSjjiUnx4L2k1fICVsPrFCdaqSjrnw0ZrWEQ0wIGmE3CV8zawF5VFWH+NOYs1+6G
/B2AYjleIAnhWsJNNyn0bleVNA5SYx/lIPjXL7Gz/GR1BaSx8oOwguaUji+o3afGlDg141UQ4bkd
TyEeHJ+nigREcgOjsXVf6uIWqBpPrLOdpkegFWMbRTfxy4I4yrwJJ03jJ5T6E3crwwyIxXnPn2Jd
OiaGdNa5UhaaMoSQchAfKqYkcLi47xCEa2cMD7jCk3v1UR7GPaVA+l2KpyINAnexNkQiwwUNoWc5
02ew4mpkb2XaxmnZtKMEFoXnc6o3fyeUo+c8WPBEF58T0v+LkFupXKMQzsN29gzfOhBFeoT5Ji/W
xQ+/sjvz2wzUzfuzhDuCVJFc2Rb4mnI8ksq0OPvb+EYIq9DOtGI3Uxqy2O6etIGgdhNxGbRJaQ8c
NJAmZHYv0E5rdO6OHPF+PWZs60tZ2gc7aAfW2TzPdWrjRO6V+lF2Ru04K/D0hx0mAIGtsDtRzZhw
JXqX2pUJjua4GEuQuSzXLfJwx87RtuTom6onJS2G5NWDhqMkC6Er2jnW12DZxYRRv7dIyl4CbxYX
CDXMBT4vADtTPquaTswC23BmCoyxb9DpQz0HiEScHIDMCkeEL7L0SrW11yhx+Je6il2kKyQ5CoiZ
vjg6SQmO32X0dNrwBNQyGC3qDLyuGGsEaL4Uwm4eSw3+y41HFYcPtp+0pBn1ha1yFUZ14g38v0XO
IITKF0Xy18wQtsmvPlou1PWprfEW9AoRycvmvm29CxAR88caPDDYS+RJDl0xDlyFr/MZU0RQO+Wt
v2ydf1tCDqMVenlQYiliaO8xCP4jiHFb5fXj2dK+HKhIMElUseQWeWtvj5SOObRdW61fPLhi9FRj
gtoutvmEy13c+u8oLmCmZZa7bYTqH/RqUjJlbyEpcTCUoNQSKWPddFgPBsH/4ThvaAGzdm1++1jo
rJRTGMSgq6DVvJgBx50EIqRJPgolNflVMjuu8VjbPUQYv/Qr0OhC2jbKTGKCCVpKrIviMsJBKf8i
OoSqtCLmn2n/7yrDaP83nZ55+cYBk6bwVvINsUJ8vx4J+Zpijb6EWGcqjv8qS61ZnsdEuELWHiqp
pcB8W/QWeC8ViNfs+8LiOfNV+X2zhidC/q1TQodksoXHjU7zNJe8fWUVv5NrPmgzVGS/LpuvF0yD
8Ptgh5TK+XzY83LWcOrOh+MdKaQ2D9ld1AG/feDc+lswxu25O+kgJVFg/rcQZMyB7lNLCr9xRRUi
8sHK2jwMx6gEZTvbYoBFaBOH7km4E1XnXz3e/0trB/QaaASDSZdsDu66J+IETY+1hJKZeDb95pkC
1ZpcofX8m4neojlgm2tIbs72OGaiilwR6kPrxKV3iozJHkdezpuYq7O63q2vA0tYH+cy3Au8eZoS
9lXD6iFaecjbRwGwydrUeTH4u1NWlAIQ3cDUc5OraAoVBTxqGubIgZwROhnYG3DYGsNrpJJzY9fe
ImHHbV1sp+2H1nBRwYPEwYOG/ATGjrkt0UhaeDmEtBqBr0TrYQ5KBOcglWeq6cCqdDZz+1POn3PR
w05g+fTVShWiQqeuj5iPOZgr2/hhHz8iZ3Sk6ljW4FunsXyDSkbV4Wp+oLUu28KTYn1biGHZq/6B
OepYcrtG7YGIHh/HD5shpPyPBrrkA5/0WizY/9d8w9tlDAZu6aygVk2pDznhYxJZsQfgMBkmVsQ5
XNHGy2vZQZ9gkzMOoxBdChcCBaXrNJ5rgPabJvwyo8xiMf1ML4vtlyxMsZCvhIcyuX/lVKnRr9lr
XFxhKQ8tfs06fnF4+M+h+54XACAoLiUMbB6HbhBPJrpZVcELqmF199JkCkXVWvZ4xceYStEFv0bG
Mo/7Qlv8P7gmqk4/U5NVUyGod+60KxQNM+BdMg/n5wFIuudSCKn9jvYoqm7Ly+y1fkuoqQTlTTEg
JUPJJbZexEHeClILjc3Vy3ymIAP9IfYJyQMdknpLFdvXBkp72BjbB3fx5UdEVeK7JeMlLabzMXuz
RY4Tfxi3UD/XIoJ2C+8ExPpGC5eQ3HJq+VUCqUfbJ1igSF0o6S5fpmtSBoYcC8iY5TPvP8FBcgtk
s0CdeW9DR3eGKu0o7VgkvaFUdOZPfP3EOdVn7uMHTmRSJ1zNxUkSDTsynqrZJXDDl+HFjwvXRkbb
u2Yeyh2b4mk3DlxS/bvjrittOEzE2CN+ptpnfm3YOKKa/vDcmlA6Qx24IjM1440i5R+XaGDRZGzW
OvmMEDbiuyc57MtmoRVZvMi1mVaunJNYhyM8mD74MSBjB4zTM5aMeMM9RtcRE2ngxtJtrAzKBM6F
xRpNZGeGcL29lIjfJsPIA4mqsO055c6DDecXjtwMpJRARvYqUSoAzpPJLlWIzSiFEAz2BTp97gZf
i8ir3B9O9RKGtoSCGKXVV6oNauB7/r5O7BA+KHbp/1hQE2z3QBRJ3pxkUTQO89P6uSTHYAqi9xtx
Sik+LnBrNA7dU5voGjdVl/GmzrMplWfkbcF7fFGHsSH3LplfLPUMIJ7yCDSrpy+9vxBjWC1ZLF12
7UHB9fuCmrlDdollCkDrTapvJ2Bjkq7OUDWr1c8I34EfEqGp7oMikZw/7v3iTDrH1EXBK5NYWi3T
NEd8vJgkw7MxEvjV8uR12puKhCzPPWPuakSp/ufeC3I/wD0Bggood0YRUVBnjSAFWUTeZofW6iRG
tPxvHXW0gSids212JFrq6b1tImu/NzuEz/HN6CnJWMZJhNch8jgdkZEq0lqGlu8RTbnsjYt3swMy
AaGMNvstU3feI5dpskC0gI00NonR8cVVXb2u7VGRkiYDQ+7ll1KltjizUhIwQkX1QfyNKoKraP15
JpyFaHBZxzcdxm3SsGPjEPH35Ya+EUZ5BWvZuGqjPRmUvD97v7l6uhlnYBnlUjzGCNaKwwkweI9e
u9zZVGfy5wDCe6Y01KHj6ESsKZZmGfyMS02B7ICfkx42aidcvK4mZdY9nTMgW2ZrPn5qG2NOoru8
PmqZPlAd1+nb2J2hujToCXno/mpT51zoMcwFXQHIGl54sHX0sM3otYQhFI6yngERMp3DK/2/Tp+y
kMynufMHmR4IrnWkNgzBhKYJgxgqvrSEgGDLv8OtfDn7AgJPnMN3QPdhvP+o8s0+b8P6A1Q4E1oz
BM+lhlZcCp7oCxDqJs8r6ELY8u0zCGyKbQlRPkBHHMwKjNvmAm+chpDwTpTfswqT1NEba0oCGkTq
hLOcE/D04clMXFA12Hbwk3YF2kko9Lzcf3yppa5JCoOlagad3zB2lIBQ7ls/EOM21fXxgU96Vxw1
uYhbmFIwED9FjZyAupRAStAHfotUSDEbjdxrmwRNJIg4aBDMw9WmA2D1YMkWBbR5WaeYb1cjwes7
iqkNvwJgjigPZgM/m4gTr9mlQZSmGCVyyC9lZ3yJm1NGCnjT/LLBxs98nUrK45FLld8V+v1WgVgo
hLBMLop1ZrjEdaAQAbV6VhEsVK5qmlxR1MV/VxUFotGxVw7KpW6xPJeTff4GQdULRG2/c53R5Sb9
THZGN2Ip+BcFWZPZWIbo0WnK/m4450H3QTYLAqjTcBNSsg/FcROiZYG8tt6fe8MyZYlg0lRHCW8n
xD+d9WdZtwER/bePvqtgTPYVQ0o2IiWqSYp505Mgd/ny6mftSrjEosTfeH8eOONpOyeunB+1WeI+
oUKp458+Mj6Vl7jBzk+TICwwNJHPP8raGx0UqOI8Ab9zI3NtorkCAk7n5ytZXrMnHhF2vlYbQNof
EfiiuOh3/AkXYTnhqsy9lRqo7gxAQ5kdpt198lrsLycQUbGioOAgNobgeqetrLhXpfl6aka4o13z
HRlVxpFAi4yuVJfkafXJ8ChwKDFFNeJdNQz17Gc3Qg4wVIn45HJFUGHniuzy7ifAvVOrKyji5sAt
ee91BDIHH6BR24R2gduQM+wXWiV41BpYVTwW1/lY1ipx7BD9iIU/Xa1X7W0u2i4j+02eNFGWSvVB
qL11in/C+rv6XaOzj6CRSjArbR54J+98JnPMiZLOzHDzu7Y4pGfJ9/1pRbwG7FYQij/kC2jMkwnh
bgcSy5guc2qvW5SdPQorDpud95tsntRif6+FOC7rkLKi8dMywjd+HF35Wq/4+fw841eUZnwjLE8f
vAfCO5nrMGagtrpGEBC+lZQzDP00e3E8R7CLMGQ595WhwokSXF0AXygkh4C9tg18ygKanCwPkIQM
VLD+oPQeIKNmV5O5uHYSivYBgn5YmCwcHf4fTky+cTeUKQAMCcm9hw4FOjXsVbWtdoVvUuBiDSVB
jBB2QSvBQWefAp6kSSicqaKbYOczZLiAw6JJysDLWrCK3rXByuDU3cM6mmv+qWBPUAl3S1kfy3Nx
CKaaEteCu3s0vExLyC/cyCqIOpLrqFhWYHLYh6rU+RYHAvD+0Wo8i3oaP1f+d426VRrEkmtkVEGX
i8I/fH4QvaoKZax+hq90VyG9q044N2kCP0943y3BiXx9wlsqC+e+iwuMYmRHP2ByGbvOI4aiqrxI
lZM3JzKKkrK9oUhpUz8ms3wZzkH8H0D8nTfJwT0wuY2hiLN/HXCbuFRyooGxTHBGXN9R7V4d+8lY
paYiFLPFZzrTqFXFA/9/eoAEm4TYEN91BJ3oWTzvVAH9jh/dKw6FarctehREjBxvRb7pZuHBgySI
wAj/7v4Bflw8FzZaZpeb0oxtAgBdoizRKdjJyLVPEjtmssxKzykOvXO9G9R/+rGsVd1Z1rZh/5j3
5BbxhPxcLjcLoct13EQrLFMPWpBNYHSdMkiUhfjbZ6XSD91YqYsWX7uK+6Q1d3sPMihLwtIE19mM
SX6bGk9YRL3xV8VjiusGF/fjhBBcXcUAjrBzVoq/xB3CDYwBduFDjmwRx3y8wOLXPg5NBE4HTvBD
V1yrpN0/MU5sYAKjwhT2M62h9MDE7IdmpZlOPJsepXkiZtDhVx/nf6wat5bEy6JmFFu7EC/icYPC
C6FBmxoj5QLFiGSMfcAioHtMTjFAhSE27sDhNCn6C3G1OvUdLaGY/pB4Yk1K3wklqpkgnK8Yu7TZ
rQduK0LOlXTXTdUfzsQ547V1O8x4BkwrAd3l/HfUrQgEmGvZAm1mLbwi+ZuBM1/fTu2LntAiILqV
dMBPZAwKpmh92fab4sLc7HHAeGTmLpddvQ8h/mJjZtJ05ch3o9+qjS5bohCOJaJEHFUDfE2xxwN4
0F0IJ3l/zA/M6FvhIx8v4Ko3aB2SZGyrVgEKDwL4uY1xV6mmukpYaw3bwnpyK2vCIhf3BdfoWeqA
OyWywzApzomheW/8a36M0daWYq4xuYgg1cQZS/K/sI8Y3DwbWtY5aCZTeV1B+kgQL92TRWIeMgPE
3mzlOK6ctFmIrzAf50xFMfQTm40jgtDIiV6ex20EYDGaD48kZHXhAo2Wxhq//RkSH6C/Gtsf66C4
Zv7GHBI2CLrYTR/6WuRYrST8g7TPKIU2hnQ349Z5Qvv7GGj23jvW/rbF+gEp8C29SRQRrTGpEZjp
7V/CbQ6Vc3OUPQF1/qQn2549Ocelfxi45N+gf6KIwsAKe8JJ2VIY8sSbxm+IJI0Ucb1cYdzsc5Tf
QZW++KqIrhcw+pvx4owHCcQDyB8wLcFOWp7leIrdaSfQdJsLLP+x2GHmxyT2OY0cU2pcLpSVbOkl
Xbs8zqfZo1tpq55V7/MaauMms6++n/n6yam5v0lWGEO3rUG7XsbRpmWbqC26/ruwTwSDthKnZqeR
G2/aprV2bSbiKTt4/0W2pcgmpiYH+b7JXntonhAUavGNpT8J/nJNqVedB4hDoMMnumz0MND1+t/e
QznM9ux+7JhGSfbfu3QDKn0ETiOB5ODlayUkOR8ZXxRbZdkPTTmvpkA3he9rpvMLLQXIs2pFCeYB
RhyexiizDEUzGo/E0O1olUrk3fL29+xWrMKBA9ThEUYw/sAJbqYaVy5wEsBbtK8f5kV5yPHtHEsZ
9oYXny9VXcD0eHsW48NNP1msyXQvB/KKZaeKW0jS6t3uUI25uMtnkS6D2iViZhWsLcZg6g+vFEqn
vt2DDEsIdYyQ8Kz4l4DItDF0+YhmWOITq8wJPODCBSgNVtWRX2d59goj0P6tcVuJSpqn+Olcj9q1
i2dlMTeuF3C25KOOuTYx3N6M41UlguiEQFslxQAlFet7bICyPEFebyvZejvdF4WDLJ67y+qGs+0X
ApFZe4dnYV7msDB/D2TsQNBOcthvWwDPZFITMZjEJ8NPM9r8kTZBTlHPC20wwx4HJt5l6YeX9bDh
ZJvP4oOA6yPCS2JVySkyPKtthbsUTlBYdieFix233eZkPiAS+JhffSlUgJZCW1fKVZTq4osIrpkP
s1CpCmZOXZFcznVXRkajdYWAcNW4w0weW/8Rqw4glCgE5MpEIPHyrauMY1yiwXDzcR8zHCmKMt/U
EJSZ0agGIKvDRRZVB/GzcVrWem3asFhXfzzTrtI9chNX7Z2s7zCX5BCc5UDHcs/2aes+mw5dkpO0
IqTZl+AKCWgBh/fhmdbklzOLVcdQpBE4VCGrGG0ImCEoWMyNTp7aZE0HT+zNxWA9etyscbTTsM3G
Pxz8F2oWgiPRzQ3DfsHRnTqu9Ee5SnKwBq7uNh/08xkj1D7bmfH3ne0T41bn4sscDsGU5fk5nvi8
CIfxg2nAA1ldcd+wx7W1zzzlnO0JqXWwt+lbv3ycmzc8PcIQ+xYcke0lzyKJ9wBegaXqLyNbwkqI
DfFrYdlJz23zgJqo+pQG97J0cHhF5M1qWmLzwtnBu/SZWA8+g+tI5QnOWizA/Ezzcz/MOEiQU2eu
vbG6zzK2VwtNQigtINz5QniiEp+qf0JLkRjCFtMK+zqo8ekJ/LOhkvcP+TylANYXtgL0M3FHt6Vw
zx7iybrkPVZ/Nrd2qZuvEQaA5HGoZBGlpa19Yjiu1GAZv/6df49wm2Oo+zCfiUelfAIJa1TNqNXP
SeagWdWun6lACZozAUdRxFdDBbKxWeIJF8Fxzqmcvwtw/W4qVeJsqVJXpDKqxuu3RHNQbFOHme2W
QVlY4kDTGm3aQI+QnTbJ2zownlsbQwhlD1kQv8AYax23pxaer8+uKc5JxvgNq5Ebv8B/p50HqCVR
Fj2SSo0v7camyRbp7ZfOX3j1HEQVEnXYtZ3A8lcbY4FpGVPHGABrJtylj8ZuncOsVPv7GtcQS7dy
NgYUJaQu3Kkl1W9Lmn9PFpYLRBY8LxgJXuvTmn3g15/FLpBaZFT7Q0MTiRpeqpc+uOEvjYSIiQLM
m+mvReYpw0eZMwej0ORECx/MVvjZW9KebMr4PmGfcr4Duc5uU/e1G8bCVNL4uTVtymAuaCrHYrQt
l9czGfcEZDBIpisrmHpYGrgTSd3FlaBT0muyAjCPNAYjq3NKoUOQuuJA7vlEbZ1yWL9FQNzRXsRb
OsRKQcusvnF2pIbB8HWI4j6JjQaYXycqcWjNZB8XZGpynb9TqN+xIG6xdbWXivROrwi4tuj2wQMM
1hZ2UfnqtBKK0XhQBZZcjuiotKmnvyJgHYaZfq4uxMogskXNwWuxqUzSaM9ZqP5sBY/xV4aWnrPp
9Qq3vp5UyI4gmWC0qN9TCy5YtL/+8nW2OlHxE2YhacSuUxir0IoeWAFkMZqjUfWBU2rHRNsoIlHJ
+81/uc/x3gJSqJmOFd5LYk+XlBhVy6nBVCJnp8+lTdW39UbT56J8A0cjx1Bdef4qzsNDepwL1sO/
8Ck05w/wG13oJXM+7FNlMkqHgba2oxswaZcjyA1r9AUBV7p1FeRmD/VlcF5hFdE62izjTxYHYDdS
iDSUnDVPbKFAifoZASzmDpS7FkCh/W0TC4ouBd+9QfazXtUu8k8/YU/RZ9Yj0thpbJqc8vy3ceQV
cCgy1VxOo4N9CjnaMpsQ3xsufrCoJM/qvI3mL8cIdmgViUADuY31vcM7AAzb2EK6GvjE9AKvj64g
QWLHmXIDG1BRr/woSfqswLmGHiXsZwYFxzQv0hS4WwWEVGV1/pVFs6FgD9Sp6FDWT+U2UKsIa20t
EhSPw/X8vfm1DjTNM44miFQ2fRR+wTElpa3ZaaRd2Z4u46FCrsmmLgsIewbGSYfUONc5BRvEBfBD
vG0kRfq40YdDbPdN12bqRROqX2iw3xRlH5HMqfHHpUd5qYOUYjdwGvfpx/51idT7f03L+CAys6w6
F0mCSvFthNbfF0ip7yJ8nnvl0ZPOsbqwbzJbtkUjE6KLPHlsXmiwNP5IckZW+5K/N0eJ3uuyhIv2
Iq3IyysuqzeWIw433AgOYlJxY87OaefE3CpyrK/aU91GFIdeiaUgclHtMgGsDoihoRGgIykbpKRT
7kz1Jv+Et8Pa72VHF5G+DFJYpNm7X0v/cjonb5dpbfeMAdNeemhlyNMDyM545xWYozsbZEPyWQln
x3TYHrwIi3tYJNQYMJR8Y97ghiqvmUkV6iJwIHQkU08I/l11w+OTxGpdMtUmkDrQNx3qzLxX7Rrc
cdWOE6WYxD0g15Rr/CGiaBo1+5Ev8hkmZ89+OhwatKd9Tn2wzLIq6/sfrim9ecWRCBlAkufQmwfj
Bz5pz/pdWEE40L1BYv6hDDz8CDi0vRFyaPIVIyO8sW9/9Jn61NUrQ55KEZMEwBDtkCzdPSbFgwIK
TPrtOmwlYsmMCUJVAUeeQiM/Fld0rdf4MjcqfODAsTJIKZHC452ieaeKGTNjj33OcLGUtyMB7lMj
HE0+GT9lf9OX+U+3gSs8hL2HCz1iGWanuuT4hDLgHbps3LYtSajZyU1rIqbuS2l8jVSYEXR7dXsI
sK+j9d5Rn21MUvgBj7SAsCgQMI8yuXlFFkCQ8wqMUcCE3Z37TdPuqvIzyyAA0rpJkbtYvirW6mHL
PYQ5XZC8OsK7W82CRdVS6bkG0v8WFDDJnFlCxDi+YAEON1i9I+eevMv7fKEGXg43YSzm9hTLKCIC
qaU3zixqSlSMqiSwE/+PHs1cGr7pqsGzaJUtiD1UHSvxIosCrXLh/TRQBWXueaHeDRfwHFf7jXTh
4oW1mUYUoUJbzsp9K08jeX2tBBlaCAqzVQKRsn/citbOu5QOPh6kbU/L3+y7cniwFbwWke/Ehc5s
JsZx5kNhSnVzOHwMbdmopINlCa9/NiGRtDpN+v0qzvSzFHG9U6ktAns0qrNYUbZXzM+VJt7ifdLM
WveJV2KZO7/GNBICsbMUT7YS2V15/LNGf1kuMIA7OTFih6lwf8hC+hy74S59TV4/hAtgYgiL8S4b
ANmBy7rmctiCo235M5DkY89Lvn68HXI86bQUtEQjhstSqkP1SYC2boS9iTUq/vtms4M3h+Lcxta9
XlckOx10QODeseUqlZR4vZcp3s6BpzOGkE0hL5NsQHIp7tIaT+xJxn5WXLg/Tf7EwUHPFYDVUncN
Rk90VqMyX4rWrgHegy3QaK4ldP44Q6AfVp3fIMf90DAz0zIFfzBa0VddnY7hdzlnGUx1kwCBkg4w
hGBO8vZOTPVAGY9ZUJi5rznEpwa9ZKBxFJPbesfjy1hxZ9AivYpnPRhquN493VTD0o706Puhshyf
/5i54/Gr2NoD9PGDONFPkx7yfZOlhJF3RXcVaUBxenLU5prXaASSl7O8WCYCc2A6XlPBGwWumKWk
7z7vmCDVqKz+MYL57ubibS3Ii6TxNihI1zcyy7RXu+trPq8M/DG+rASPMiC+afr78hvSAohAp2cT
20oDeC8BPIgBCZLJMFYKC6p8Oc3HtR8iKjZNVRKZ/ffCXV/6KN4vSWCy4a+aLEep50HWC/WFr2nZ
qadRKDhbtTXhepRptd0knd5vk5gwyR6edgbaZBZIMdkM/rlKpQb+NNoX4JPY7iiVqwnUbOyER5WH
Ixyz7KFv86nOayWeIdW6m/NFaNKIgCyqpBKJQCEX8cqdyRP5aThhMRp+vAj5AHIDyLwfQFA0Cioq
GkWAEgiebhYt6Yjltt2o+DyAdnf4OTMn4Con3/oNZgpzbjO5fniB8aRdkc9H6IpApVakeczejtUi
xrqSbkvHepTxrouk5m6H5UmSQEFz2r52hkib81nAcHPrgf57pXBjhS/npNEtdvtFBgb8pZRqfslK
cHvW9LloTzbtluoKsffX9xPuJ1yA3KQ8tgU/7W3LUFSkTwIx8zDsgGcHBNHNfZEVfdfdG7sU0YZY
l1Jyrmifu84574piPRV+mp0+edgRWUsu3iYm4WciJp6tJeOlAIo1Igh3z7xXbgnx1Ci8RakWbaef
fncUiq0Ghrh8fBz4aHzN7HE02+CO4B4+EO6B3nuExUVYoEjw7zpRg6KXNaQO+aXiRvNb5XOALsbO
PVWwGbx0KpFA6ktK8r7qlKyjUxn6vfdI0IeDxpf9QOw2HyWsRI7VmyC3eqjBAenUcz3pe9AcW9GJ
ZRYuVxiAI6tixGPvq/sJ5oo1hsEW1jB9sm3A42wzmbRKTqxIf8tHM3AtYZVni5i+Wa93euFIFTIq
2Kcbf1faWc5IPHqFtrAFKxMsJ/YOCVcbzo2gMky3yAfF/UqGs2bibedxGbSwWIf5R4NlXGopPw0Z
Wb+4N3ROG+pyX08KQZDVADBQYVxdhMBF0odJOQuz3BldC9+KgY/VTkdPgbFSYo3lC2Ywta8wWMAf
u3xU4+D4kbF0t1QZlPrnj982P8qeXjXlyfAlLTl7pVzCS7yqDWqhFWDw4dL9MujqzzYQM+xj7A6L
/iiysMrefHHxT/TOzpainlQEwLjwdM6XqGuqKCK7HnQXrowTd63hUadRCCYM12qBc3TFNpc4EvFq
f+NMBDAmwu7l7lQLWIQJWrRxX6YqybkwPib59/Iok2/aNSn4tNOi3qv1nEqt5O7mT+8aowm6eWMs
r4dvZhgeOsa/gEbV0+3ebRA0t2WyeiCLnxP11NQAmZAHfS+TGLwGsQ+YQM2yN+b/1aT5T8m+x1jR
GJ4Ro/mOzMbAinY4Ji7u5uZSEQsb0lc/2qDBfVuC0UCkjUuYO8bCH/JDp6d9KHw6py3htbuFdb7r
u7jpyD+AEtpww7WETCulpR/feA/tqic2cnXg+vKJtgXgg+lFrRcQVTuccIE7Lhwfwj8GX8YfqUKB
tc4ug2Y7wDjydF/Eo78g3EkB7fECXaDIxZYTOCyRqFPpJEI01HFV3uvESsWewlna0GY008gcWXi8
jnHtRNqCSq6fdcWkbYdMQWCgBgV/jKWdDjvPvvpsVHb/acEStZ3hMPc2d45WyW8rvrwiodv+Wslk
FyNmSoSJQmr7eC82f4qHeKiz2M7BjWQHtOMQWbd2EM4/0tL0FtrLYAQB+ym6dTuKuB8EOFuTmXoP
mHz5f8Pxl0uFV6m0tx2Ro+OS7UUPAyDlz4w6zCynU+DaWo1NKAm7DmZshox4FeuMWvjzBsjdU1Gz
hPkCvqsitOKTbpPBulYWSK6Rei360FXcTXwEkPih+VVd+cAznVlQHzuq+mXqVmVoYPHxBZyzgooL
c/Ss+scRn3xiKPV5G6qQaCzfr8tZ/fRLnQo+BNP3gt5gQ7w2TlZ27fRpA6imRi33F+1auFtdKee3
KSfujHzWzhArjsykXIcLvfLsYvOIBuhrtHPkpTWiscZ/q/rOwRhJ+jjzWecZzqiawwIuuvepsXkz
b4ocJ0Tnlguf1RMAysAMxbDicfz0iN6D27nNdVO6AptDMqE2J3rnU5ItGuAwFj3gdXa0bbN438XD
oVeAdiJlAZXCSkZ5/Aqiey/TSQJGnsinvcPXo2/9lnnQtbF+1ZraLSWmLQPxD/ty1JibqLHgT57U
eCADNvu1cp+/h/OAh/LbvRhtSFTQAYKyJQseZY3B2S74+CzuBj8OzQkLay+mCT7Tt/vqGdr4Nke4
3MEGws7e6ZmjLjrDl9dLd/G8i3axKwcF5WQEF3j1+hR+tT2b1YaYlqot1yWB0Y1u6AleO2zEk335
VyQzLfGVVycr7b0TZFCdhY5bROBiGwqMoen4gb/dtxmb8sctLRm9b0fnct9d8s27i0gy3V8r51yr
6qhnfQVjMdYHQ/IYJ2XDoNLJgbntFZFpL4QJ1XPfOX64zM8tNfcCo+1HLPjT68utisi5gRrz/KyD
xi9zbwFfJvvh/Emt34tEJBSb3Ikys7IGcti4y/PXa6M2woueVpxzqk9uhKucte1j18FTtt0Zwk0S
exNa52E0xGlYu9zIOrIKwDsvSDmykoOeW1sapkPM7fOkqfa5AiC4Ll5PcOjpJ6s5v1F/npmYb4Fq
AKtrx0zdtASTI91rXZABdxzE7iHybqECMidFZKrRH2HUI0ltlIPrb72f9kwXJewBZ832dz5V95Sq
JhByXGxKFABYirR8iQSqreC375AqR6GZYTuskOGjBNEPNPsyPzGG2FYMabTWlgh6T9yDoRZugDie
F4Vl1QantT2O4KVvsYoLIjzozkR3Yl1eNf/otcyoDO5+kTsfRiA26V6CtY9yl0/fy31cvRNs7uN8
V8B62a1V3SBD+yd2mJvVbMZGO77HB+kezgAOppDNwOCFfL0xYOM2jiHWpvVtDSimPyZ1NbuwX3wd
9OaQtafAKG3+h3dgoQOS+Feo2NLH9Hjyaa2FXlnUCd/xjQf7Va2Vti90gzIeTcXd43FUnSKB0BTZ
rI/vo58oYDqmMbjZgnDr2gxY7TJTqA2KGz9B0u2LxMD3S9YNKWBdm8GdN/ojV6UVvITBQcNPkGd4
hQKJjy4kir2Urwo2KEtnz5qLGWboQwgjA4Co22HifzTbzbl6Sd11Uik/O2SbDbuQIOzPrcEKUNK4
94EfILY/ZQ83Stdd70n7O9L+8kz2ubHyYQC9NsJ1mO0kyIpDje6rTe6BBQFA2w6OelxK02N/dojw
DJwupw8cDZ9fWa4+SMNAju/Qr2B80V48fzos/QViEO2N3h881Q1zTAQbnSyEFclJDYGx6L0qR0sr
jQXqnRZDaACeQqOoiZapE+TEeZLRXnRb3SK1//vFdm6eHV8TXkQ2YyJ31ayVxfTEdODAgwWtlHTU
SUBg9vuLcg4RfwoEQ2jd+ZRh+cMEZA3ekWtYUDsU2wDkfc2kbuSZLjqyDZCUUa0ELFnYH7sPHJg9
UHcmDqqmFP7t98XzCQGbBgo+Z6kJQ7OO2JhrQBgKGmXdZUVw1/d3xEz/gA2s312OaRH3arKPBMSF
z5dEUQbHO4Sn7ESqbHJ0ylM+rfDqJ0wrqCcJWRPKJoJCurvfY/FsDn7cUmvuDaxWkzDQ5ZnnFvmN
yD/O8j9gE10xjiesrm7axQn/oRea8LMPg+EV/CNb8yIlBjF7fil/nsi6KTe+44ArLI/A8QWG9pUI
wagZ/X+xbzzyApjGJWGpdzDJ3NZSsGq+I8VtdObgjsNOlgnr3QBZCtFMaTExTbu84fTjjaTfbdIt
TBWpz1gFQIMUJE7LVHVfxRaZEemkcmdWZCLSxRIz8bMgnmsFj32IW/KxSdptojhIXMCvBcN2elH/
XfDLQ+x4BlkJUyjEQP5iFEiCwXKsSlBKpHJ5Vm1b06vEA1/RqJjj46866RthqXQ26h635NQlhWsp
PpdEWp25pzZCNkFHB9E8Qwau6KYA++7ubHJs/q6x9HsaH6WsneLuvbk3TyFmnXUon035J/ppTPIQ
QsIRr6SAnKGcyKQfgRdZeI+ZFGbkH0jiq399zD3hMbNgiBbhNNQfx3AMymDrP5HTWV0QwWHHYkxQ
L1zmYNEvHTiszCq9pqHiS7K/mpD9szGirdzbRV6CF4+5AcMwPCN+LAVeB2odourF1Tmj+rTS84TF
n5SDIKCqSUf6Y5dTDdvcURgJAavPG6kYR/RjGdoisoz2u0TkT0ggEprYTo63qwL03XH/iigllV4E
QvPHXOrTbpVdDDn3S0SZVuouxPHLD3K5uxbo+bkQ4Rkss/yAysg8L3T61lMcVZP/3JReIxVcoa/B
Qb6hn1m0c3EbZffPNkA/eku6so0K/zOmGGVWU1RrPT4Cmr8QmcCZYb00Xe3nZVHTg8on67HHBnXu
rFScxDGkJ/hOGOt8f36+fDOv+9i5siV9UvOZngtqFDZSFrm/37O/OlD1Dd2jitW2j5Wbrr37q1Ks
WMuZwyF/6LAlLVPzD++sNkvnkWVRj3Pwc0UVTUgab8EK0EyLqMH98J/rn663qgtNOzv/p41L/cDb
K9C+WFOYRMh4ZdDzHoRI7OKAipNmNyuAUGbpkv0hmHAp8UTA5FiwlsVNviaoqbQrKAl/rr1o/uzd
pM4ep/fkWcU0o5zvMF9cBvWNLvEHEx14YyKkM9SZ9vhCgVw50oGJqRYLxmu1Jo7k0E8ZDGZDjLjh
UmHJP7VHTgrcou0LmYBxY812Tm3yrvVtwjTczHckF2CFVIKEirkLIs6Xp4X9w3Cyei1b+YPZI3xH
JQIE/sYpGDVitv9vkB3DFJA/ITlpMp96thoSOD6H62WXvFjhSSRGrivWF3o9dzlZjRlL1kH1muQi
PnlFffXpw2DCPs5ECgawmnY0mCmgWHXSeR4b7hHQRQ/e1broo+5FyOGE/VqxbKT29+T/p4X8rFYr
FSyPQQnT2N9yjpxNl4aEHVqNoXNaWRBOf6dTmAQWasCHU0DkWaer9uQxc4f+FtgiGZGrR0wx4qEK
ULnWuKCJQSa61FeX5yFep49t2Ka9tKYIAAaVO6kkxHLSlwUuXv3WikmoVCcdVULnAxiczEFBvX2r
zIVAZnrjbpYMsg1nvVCVCAHzoZg6oqga22DPXunge65fUunjlDRxi/Wmn1AWe341QfNs0CJLJIZk
09+6pEjzzq6uY+5DJq78Ukb5QaMPsTeTLMKh+Cp5Gpb8WV0o/3CLs1fs0OXaDfYlSrV0jH95+erZ
q+DwxzUOd0o+6t0f1qIKAyXglmDm3m0/KcwzSx8aNpz341IYlfEom7sDQqhE2olvpBG4HXnKuU32
obxYOqwMg8OhWUgqAshKWpkVb2WuNIONXUFm53pzsShwUhhaqOmQMUBGQLxkmh5PvXS984wTeZmB
wd1cA2f0ocjG+M1h5jgWHYGYvzp/FWCEiRJVnpVOZMrGRj4nGzHCMLlXwxXuZc+RO6nJoYnkudNa
dnX1gkcY6i/gLCUH64IxhVxOJfzdiVYDgT1QxwXG5m0jspjvM3UGzmCKzxo9OaOSUd+UCl+D6gwt
EAk92AvrMxCl9QHEobhbfwxTGS1dhXxZRuRtkfW8futc+cUHRxsCqNRsytflI9R1OCrhe96hiblG
uTJhAh6cf3Sjxwotah9FM0XRbCeZxjfGLy+/7xLkkMm3I2lHmq30MWSM0lh2uPwQ5LFS7CbnoAWS
rAEBuTTMhNGNlMkqqkYOduOPJ23nJjUmD18Odm+GH08RfzqTlFr8Vzij+k3EizqINMFu90RhoFAC
mjKO90qRkxfAjE5jIzVxkbCgybV0+7a35oCPnvufsvU9FPyII8PtW4/lA4xryLRuzNGISGlw2WbD
g2JT2WtHLW3i+ESywHIu53NvPFaHYLCDlzkrI+0kQ4stQh+DnLTdcEjFU5P5K2vRveP6SsJat3WF
Xl8N0DcQBI6c2TALiD38kL9OhCRT7dzo/pqrZtogKoSp+/QmJdcraUnw0z/qdJWL6+batke4kEfV
/6LPBxo9uT4OGiIfJT/zIQ8uWu5hGUrSMrno8QQw2YqeaB1d1tvsr4qrzgqb88PdBdg58+YaQXsK
Z3fo/4Johv/vk5caPSkwECKL5C6zegsua2zUZmUTzGm5aQx9z1UwfeunjxOeQDhMHRTISYNm5VZS
THZnv3pfTYeHHCnlSkrTIfyWsqzDHOuF43XbuwciuS0ucUwKkPwwuzdSkqeChW2/rtyp0VLxiWWS
UnqMUkn8AU2qpO66pO/lMAiRfUAU9H0LMP3/Wf77vCIvIH0R4TfpPd7tcj7pKUeDMAOfbu1LwMDU
TnLRhJrPovFB0Ej+oY8VhqV5yRWq0EufYT1qSeeqy/bypcKM0EmoH7otVWRqfFWy5tnTLx9dle/Y
qpanfhBJB+U/m5B+1knV03edguz5LnqfD2ZNhxTbVONufOgSi2WkZuMtXMUGWTF3dh8TAwEpA8Ip
mkiDXMgqy+AClR2KWSa2r/gg0dhZFzgqPBxI6+cjoyQihLqtfZTb3ryrs01DhwdSqCzjhHLlx6k1
vnyO+HBJwRAlATf0Jv0S8gXozxcSiYXHeCB97YP2ti/gUNSsoT3y/IX64P8/aSqEBKr+qaKqY1Xi
jE5B0ho4BG7I63+zF9GeNbtfs/qy59obnFlE+6LHJbC9QJT9GHO+jqwghCl7yndEPk2+Gfe/MESJ
WnaEIi8sVnOdja1DIRk7GNRXXRtMKCbmU6RxvafWnuhJ+OP4m102QF/2T8OcOwK6sm2wRhQLLP5c
yMdkLF4s8QmoUnjxfVsMYUcB0L3hya1v1fSsQ2NOdODL2aDNwcUKA4CLMaglFLfqJb1bm1dKMZUZ
ISvj+m2vjR/VGeTalHgBAdnQAxJFWo84SkqA0IzCuxAd/pNqIcHVsy9Trq5P+8+v2ufDXBdxnyP9
ASYwzNjeEG4nV3KpDqe/95ZtoYOTTHR3lv4XvmphJaSTaoN483GZ0w5dDSpyNzPkdp85wiIDhtm6
IJfEdGOj/1BpGWkMPr7zzmsf74rH+DGXoUk2WYS662S4Ug4a0IVMPVUtbfMrqqYvle8rwbvjR7PQ
GRbPmNu5A6S+y2D0yiyc1HXqVq3yaa5xU5/0Jmfq0SX0J8JAA1QMJzXISqKtYo5a7YD8bBchO+6J
mUpxcnXDLzRUwroB3ez+FFYbWwehqkLRcg/MjNWbDadIF3AdRrU+r4tigMRSquNLLWVUicOLUUip
PlFcH8H933qBv7fKI1eiG2P2/EcND0Fl4hvNRQori8F8bi3bRzLLRpQGFuTkneOFvHX+V9TVsLN7
Ow5JkiHzPisnXDM2XyK3A9YLIl7hMySrCfn7Hm0XmgLLcoqkjAp5ARTPGyRAKF9UApTvO+BXykgY
3CJh97wHk2/JphuUKo8KQOS0tQ7Vhfd3yL5tK09jdg2i1T5PxvYEEOj01fFRCMHUfXcUQQviNNle
0ewDKn4XSq4Bfckvm5NFU+ky8pzBg/CDsDnWzVyFAZL2wUVPGDU11L3eArNolojPESX98DX+7DQS
f/9bx4TWjAWiERo9zgQq7t3HmA/ClIWngSrJThhR4nQn8CDpxADJSIlgKeqv5v+qR8PIyRAI2ZI5
16Riqfxl5GAilld7vvp0Ss6K47IGmDCZmfdsowIBXSB/+6fZTXtZXXjkzWPb31N6XcFEJHSEhtn6
NYS86aA4k+zTONqXbfhsTPZMeboPu5yuFrtflelBaSWrki7LnmdHf7q4cNJqR39xNua2eGOyLS77
ipcy4AOeNZr/TDXA5a8Wd7z28HUx0WQ/9x5KP6ji0nun2ebzxR1X+iuPdxQKeDttCDtkuW2quBAt
ALq0RQ7XbXWrhw/RJDpnXCUtg95xLuMkr4Em6+XB5g4KJzyBvCR+X90cqIaJTSHvmGjnzEffwcsU
IJ/dxq3b9n15CTPSkvAFO0g3qZcKVovoc+vdifvOj8Qf+ob7fn3sOmff70MR2+fTSHrovcC7RDcT
JaqUN++LeRW5o0Cl4O0UBzugu6kR/UL8+0CXb/wMmuIBel5v0p6Aj+igfSbRQu9LwAi5GYUMa2dg
+Cq7JjuPS/YQ5GFRB1U7jB1c9Kd1VkxqM8Ln9tshx9ph/HGesIVnu/HHAdLrSYvHxMsny79FrI7o
hBY0Cv643wf8LOMNuCqUBUmkRZs8IReu5E1qGdyknwdp7X1+MSscKpYbYZCU2IZEq0MlDL076VhW
cHV7k/v2ONRBL7cPpgxbvdyiVVXHvy0/ZBinp+Ox9mF6KEvhic45LTrwCfI4Uach5mgcET9x8RNS
hPFICvFwPs3fl537PPY9X5s8gS9aFpixuv3h+zu07H2S+LIETQWIBpW1Ijsfmtq2z7z4xZlFaAyO
uRqjaMvFm6kJ1v/CLN8XhY6tt6uq8yEaH3mp6RSM3gejGkUyw9xEgGb47PFu9QkV5Ho4QHLjH/xQ
YMRO+e1LvWp6L5F9wkeV8QUUuz4Sel4wfO6SpG0mC0VWVtabLmG/E32kiZaiuH1R7FEoEY9Gaw7y
LneEO+6nTM0byakzHK2JEyKfEGjAzZEFmcYjFNvGkFUahkR01t1YjNGYTLb+44zzDQj3yTpeTqhz
KoXUHhKcb8UNLgc1QU7u+K+1mUPKxjs18XZo3uriLYTOYKkhB+00EQHtSWPq674ZPsGNhAJOzoJt
OZylXXHlaAh3Qgx+ak4EdwV9QALUOEYVrtCBYUy54aalPP4ajvO0R45CtcjDQ5Nq0EuUUmx13eXK
rDvai2knWEXHhRsZaq2FsPoj1T8bvPBc65NikzTZwQbazGHAZ18ZvhKp10BW6InL2DtzJpj6bynA
lp2WoSosqO5kth7Xk5yan6iVvsHxd/ReCJgESdjbToodtqn/BOZUbOFyXSjsMYuR+VcLpThD83bp
74XCTpf7w48jHJacgv8c7vgJQDKLuqKXB+uJTd/O35GfzUZn0JosVybaYOk+x2t9sy/7s6ncr0Hq
fHbvVyoWDBo+f4WqK9H6etvybQGyWJZzukGopcpGoshNr5dwphfgdUcHqFeAfqbRzoAkdZOYtpGI
KjdIgNrskGEdLNWZcQ5KwkHczOgiN88f4TJxgNVapmNYKnpf7jqoKOo3fVhLlq4OPdateB7aZ3Y8
ZaDi4g2C+muUlwCxnYzwrDu2xKwRijw+ywLCm93OOEkuOrZRb5G4frs0Bj8ijtmZ/EsmJp0ujgp8
X4Q80vXL7nWOddCqPYmypYtSDpTwOrSyye2jSXwZ88VGYT1C4mtKjzr82C5n2GaJ85W0OvjRlSLX
tNmQI7xLni5cUX60Nt2cXDOAylyh7mmf3tJtbILD+2ijQWtvOzg6KQ8uFDi1QdD7bZabB2gzHTkt
kgatKKDQYej4/hWLWm82UeylCJsmxew5CSs7reg75I7Y/TxF40rYe3+/sAoA+LzgZnsO57sr45XA
p9kKNPNmhfB228OgAcrFpqwd87A65ZEIBHpO5t7bj+mIRUIUSU+YsAMtH952kYu77nlvs4TQKbjh
YkJoAso//8W3oyjZ3YLgJhAKx37DwPX8pHO/mg3plphJ+9BopKdDUV3XGTRn8wDxkPGtWXdjgA5K
Y56yQeTgm+1e0eBfgoYTSf1yXDh3dKjwre1uBV+1M3eKMnI3/SH0uDobVuhLyrUv+Sou32uNqleo
/74fA4s8AFMIIkIhY+21OCtTmU+xbOWlNNxCvfOj885VnKqWlft4PN1yDbBytPSW1QbtdHcH4ByH
hP6pItqwO/JQ5Q6GTBCRMJScTn15VrojPhgYVGL+iThEmC19dG1TAniYPdFZVnoFVqEkPkcZpAtO
5+Lk8R1WcdlHWPu2mokvmHCyc37SkzMihF4vTTJsIQc3pUfpcLY6SzSGFrrt6eWJd+eLVLI29cvd
RqVA5AfiFEKGoKi/39UBLwvUTSqMAQrgMjOQJkndkfZkftyzTa6OUSRcta6Hn4QOLsgNzNLpjQJy
auniFvxE1eSv8Vo4z6ujEQi95J6TY+PuZluEEXaCxkzGG8r9c88lu+TdwZhxBGxQE6EjiTgxWj9x
JMLDZE5ng3YKLesVaUKQTBByXAozeEGmQj4TSurVtcTwNqFqNOZiDqoqm9OBB4ohP+/FpnKMI2+k
xqlPfRTy/b3uErLezltSEz2q5ibwjFJ7aopR5XWQXvz+TTb7G0ZfHI4JrQC0lfmbuv9GO1kiDgzf
g9hNzAul3vEXx0yB81NqCDGs/GPGpvvY+gLDu+Jz7oEfolGjN7etXwZO/hWRjisdtg2z84dZ+KpV
ExGCJHpzltpS+YIkS2ABnNgMOTbNxTU1whvgDg5GZIbUwy22dyYdli6MFk1s7ZdiBeAmzhJUEzeX
6A66V+WgkvCe8EGpiozuI0opgBZDE41bK7q8EMpTxhR3NagSBvHwwO9cMwEy2aHHB9z5OD0cNEbg
MdtRxYYDZ/pOfiQ0oOPBdLQZO8QOrC9uWj4LNhgELX/XuQIrTB2UnsRTDvv/4M0rpJwONeUgXTRZ
iI5gEqzNrYwFDbqUaXZ3eUHUvzRZ4wbN9cNGiDX+norh5WZH8GaS+AwZ7VWsTToW2KtplBY0gCe5
4yBACxlDZDo14ZcXhlbNeRUAoMDwnDO+neAMumZ7a14PbXix6g4x6mFipuqLLPpraSwu2P7cU9AB
kytJy1sbTOCdqwuekVsrZvyOYhjObjDVFjg0qykfLaUDLVIHYWJLHbXKSAdp7otV/d4ntoeUAHqk
r+ORzZ1P9kQ9y3145GRKVd3KLMMb6P/cqOuXc3CKi3wShh+PzQa23tpFCwprdC1VTGY13G6u7GyI
7uJFs4lphwZ6xDEW/KdUR1NAtxJt06x/z6+c/cSqF4SOmNl1h+jjmcsPSs8fT6de49MWL2H3WCkp
kjTcqahIE5nqbm58ODklPNW6QwSl0STOQyagjxiyNYxiQW5WoXOCXLbZJMD8W/gVC3fHaZC1DMIi
NvYJjGXjkLIaJDIVpFbdAdztK+0/HujX6klIpEGXkd8hNbRk8+iTX1bwkTgTU0iYUcYzOkF1hpRe
ywGQfxq1tTlTfErCftJ8LqKH0SZNgOrz03+/6qDly+FmPE1HbcjbI+2z7BWflhvnevDipaLFDqo2
jpeLA9ocFz86sgd4cClduzASyPZ7XH42L01AfQBLA7IbOkwvPj4eZEShTSm0t/vBmTY/p193pNUE
jGFPNF064ancgDwZMDV3kQw38UWxjM0fp1z2rcepe6YxYZkoKdVlWCk70lVCYCgxHm7QmXRWP2dc
D77xDEV0oLpb2YfaeERdGWeIeX+tKNTeX2NLiFiEGoMrooe0OE4iDAfLzDpspx6KQ2osZx6uNMhN
f9r2hDXlp6FhqDywHV3kXzcWEwmZavftlTdBhe9WP1GNI7KLFNb3dKmd89RgzlVvBGvLdu4pnMrC
Y/m4b73kTYy/1+mFJHAQgpJ4yqTfirBC/qGdC1pxn4aLw4KcI3b8MiglO99pa9xn5YOmnqR8Ai/O
G/yrVyGoIsGnA1IlCeDmOgfc9VcpCEPQyMcaqWkO3VAQ7eTQOeh2zJ4HoU7P6rNuBrQEEWrKqRpq
JX0q/Pr0gn38FwdWzqgrbHBNv8pkZRfSpu7ZqDgTaolJCCbhxT+csIkuRWTKASW8fQKua6MigM7s
49ezle+b67iFj8y2Es2rTc+4FjMy4OHGOUAFKjy16IXKVDO8DBkX2c7UFGn9yA+SdhaaRcN35gLi
/x0atl05YvgkJVCc9raEVYvwNnhn6NWPeJqiHqS/QIMKVCQWvCpc2S3E7Yf1DTSMWWD1/jxPIbtA
UqQFkZSpjdN7tFzG9stCis9puEnzExJZw8yCeeLeGJf71MIAeKc+TXXX+xT8ALFDZLWTZOZYxZ28
FlGyPFT8uTUD92dMSCaUMrkJQpp+1t5JVnRNH7GCXXgLBMBzwYIl74pbC+n6mYHBDDuEE/kqmYC8
gn1CFUZEk4HBOdhZcCxMMCTOWPaaPihj3m9fSBHNedTafTslz0RmunePBM0la8WOXT9l1yiIzOQb
Zk5o6SylhV9oDU0k3b5rsp7MK7nVKWlLHpfWZ91xxEZzcW8eW8QBLCSjxY7y4JuwxafPdIBhRII7
Nv2t9pOtDtZhPpT3Z6IKQg0vr7mDohM9XDRmwXttAvtl8EUTw8QNkZ6+rz+1WBzew7/YNReJYe0b
gwrsJICfDnElRD86sz/Li3lSs5qNQMNHtXEhffYtl/WHKgGr+Ehjm+81N3X/v8+15CNqW57qGDP3
FkJgrKwZOq7LPrN+JM+SqpibrgrKxyY47ZbHsaBdklfog70P5frvMMzEJ8EDEMZnI1fQP1ebuFPm
+64pw2PRDFZ2s/MW2y+mD5FRTqoOHeRThSYKOEMQtaY7gcBB3qhnEMb6RTq2aSu48hzjdH7G2Lh7
7pc7CGb/Euec99qzAnt8fGKbss3PI8WZ+/EaBeVHF9H7hyk/Li2GBB1bC5rPSmGLy6qqzOkPuN0u
2o6pw45xOF5YLFT70Z7DTTp3HpWsIl3IWv7gnAs3Bff1/DHMep79t0itSg0PMEev2uFLcsPT3ErR
fmqih2nBWU2XOGNACLc/lR7UfHNneEQtBsdqHV6J/m1PCK4dZk8I/gGtfhD26m+kwZKwTx3yZvBq
d9X6YYIsoRJYFrh2ZT6X+JeyBFR1gp4heao/dxO6dUGygQ6JFN+PPLgWb9dA07zBuQ7P325E0lWl
yqUtfhNVSsxKakh2OxF59CHB27vXcSQYjN0X00DEF+i+HdbqNhzrWTClu7gpvE79mntn2Oe+txaf
2l8B0ixPICe8qyJgXcs9tQHCUQq9w6jqv3CfhUeosG/uz+cvY13lxTbPjVV2tt9N33OZz8tbFSLc
1mE1OJwhgKHgK2vNOVsCOJZYbmBQYxuXSQJ/dn2Azt30aNQjbAzEQeTAzJganU1CBYA0rM234wdF
jVDrWGAOiTKdrWZ9pA4boSXs3R02DPP8piAQfosNTqbChdGVW9xGnGk7q8dig2Pjvhci/O0wa3CO
G28MErgKFQED7KL7tXZOggWf6CtSvY3mLdL2xlhRWSvcxSqspm4n/feqnuPrdyUNP1Lu6Z61lkfL
PiYF58HDsX628c/gfMGOLwBQhsSG7xKzlBhgW0uUcicOINlf18te50TkZNuF4ebLvRoS9wKTNaow
Hgjl2egke+d2uYjWWj5Swzb0qtJqAOSBHJbTO/7fC/5qzv1sRsZc5NAw6jmphxrkdagJb6mBLUUQ
fjA4L+goHL6ROlJDX4sxp36jatjqogHGQjcs3MPi0C4pwAQVMLUI4sGwFh1VyWvFIASnrH35lSyZ
Hx/22HT/uYB3gS8+sem/yk6zqvDLbFFlPYn63vmb1I00b9Cl/3OeKRLoC0Io5eAo9KObRiuHdXIN
WK+r7rGilXtdYzORjEG7SAPNCdRHG0MQkudkF6MerhFCwtPryHIGc5JVOYDDagHA5jCqY088bILw
lABPad03gMfjor49UoD7JERRM9GfKyLLI9wZH39MF3gZ2BoOPFCg6Zai54uv1DJJF5G7wlNPapIC
RmbWEbMh3R13Dc7LfR5ejBQVlqq/RrV7vbJOcYUXneRZaLoHH6TH5DhGP5CcR770ZdTttEx9yPZS
e/nhirpFeJlh9ypzV68i3BB2JNawwZeU5NIy9nfw/ozVF8tIDAaEi/1olMn8ciSmYn2+7S6jW7hZ
tdTrvql75POIj8ONa3BKMuASwwmjddwjjLfd49ZO12kxbt0Abm5roi+oPoDgOz4pMyGvsZCuumtu
6c1Xia4RVEt8PMwXqPPI+/O6NvQugloIh0EBeOhw1nHwzrLF75nKZnPqMWQIUzdYeAjXdHsv0k1M
e1+eGvJdTlpLW2vgLW9zM3DYjGNUmCvO5/pZRtCsZCu49EBO1TX63GHMIIjCryRWs6FMSTKlwBBt
/Ov7xm7neh6G+ShOvTZhJfzll6ukafL7rD0ZRTSI8eP4wdIoZExPlcA1AqOQhR3gUkQfWpYhX37h
QqwmlYNRU8rr0M/5NUWcF4eGlRFD6Ryd7GUpEu8eZmaxEK1KK5z3CvQefLQowlzEcC0h30FQcRir
vgAdSvKaKJhcBF65MWo8BFzu9KnravVNiuNT6h1I/ngAnuXNKdQqj/FAVQ1phwyvBJsrVE9wg6U3
bABo+XgxvEMD8SI3XH3YT5JQqPqSRaGC1NxvnEeE974XMd6VtJec2nV9LO3eA1IWRRO4m/wp29b9
EaiSr09mHefJeB9RFiCMijhEbpHXarCmRIXS4ha8B7LgUw3aHi4++WFc3azzcozOt7kYtrLzC8lg
T8MPDVcDeHTkxMMNxw0SMFJdxnYJSO9Yd/krvFJXlO1AKzHIAlSQfaZPaJYk44pZbcIp6oL0vzYj
JwoMvrEC0EPZWvm7NGWP5i7v2yyOGPiFtl2lroJA/chQs5mtaAdESL4t4M/INBVgNwKu3DJ26LJA
PVw5h+VgkG8bMK/LKhf09dJcJPmv2yxYOfZhsNtQIhXdzPlDEkERahYylLaCxXoC8qG9g2lPnGTk
V9OOrECrN4kHgoyYgkN7791dtF8tgMjsIS3omf9j5j0YpUnpVENdLkiquPXqLv8wxBemsPrc9RGD
JmUk5JnAv4XJawBKpQp94znOYQeyxYuSgtY3F+gvu731dv5b4nmlUJXq+VN9ir8SCKhLue7nlRIV
TqHtfkA7C9clVRFWjKZ/KCfcISxWF1nQVvk8HfxCl7Eh2HuNDs28y0GckZAyXyM7UTsh4fCpLpbQ
rf6W+YevP1Jyp1DJ6Alc3eTafmacHdn5dVBm6JYMVeITNxt+QtAz6fKwSMzkNn2TVvcT9HP9tTwv
1wFktz4W+LyR5na8FEfR8tomOEwIMAKcLVLwFPNyFPcB47uWgCcKsIBi6LRBibSr9XqqZZoWW25s
FVF4M62jgrSQgVeFI5BNrHRr5PcBjuJBAhQrNKEGF4sJeHF3GjETI7vwZj39VPlhkkDjTrOiuV7E
woYTC3/yyev3IuNm0qQu8nIKEudWCbb24Z7dLfe3JzbcWViEQs+e8ifVOdP9EH3uxLdzDI5zAFCc
3hTFeWAYAk1rZgddiwT/X4KVtMx/FbrPRBMplrLSg0YSvls3R4BGNP3wwexCguCCrCF4cX6K31LN
0+kE7TI9TcAb0VWIGKmGn/8A6v7jodg4BT9GMGfGR/1A7B88NplsGcg3jeyFlrNPGRbluBzYP9xd
Sm11WHaTtAKCuigw2DKOfqiuuckG4feEFj9cyOG4QXxtbM0MpspP0L2xEuJG/o6J8v6RLqsqiDYq
/bU9V0C/xXxHebRezk1rmOC8RiA8p2KtGyrORvgjfjh6AzXOXA3jsK09n2/yHiEIZ4UdblbMcVES
nBO/iRuKngualvh1RDNm5KiyhCLjjGIDP+uYOXnlE13RyzxKFtzas4t7spQ+Th8yLcETcCJRz31i
WXeE18nyZs+Ey3Can8/nTxxS9EhW/KvWMwl6jhakg7KUChLCZX1aB0jk/WfTzU/FXa4O6OAhj76r
CkqqZrIli6CPBu55/GBOUPbpTaWvRrdjZkN5dT2PbKZSXEg/H2sRXh3ep4eFzGfK9c2y1wIRVMoj
1ygQAs/KX+9/oMAsZF3sE+8PLHGgrLG0QUpKTvBw0IPwsm601aU/denmIFuW6M0qL+SuOzK9KfKI
lxk5iTziAz144RPK6d3UzLNSnJ7gqQINutwJs8IFAd7/UA/5TONs1ojqHsUOHAwaTVRItgRdmc6S
QEia512bmK+RTW5kbs5PQI7D0WSXTP82BhkJTMj2G3ulUgmXbTwy9lV5UIm7i+8IGmBq6VkszRbx
lVIIuLgyTRoQXmCX72yK6eBT+V6C/8thiiJqLXKm43MRr0rVvDHegZ83isp6LGfh5+n4k6YP+meR
Wab1PDRjfRhTb3SlY9378I/qbgtzmJQRVTwQYfVWdZVOqHRxjDlaeu74JxdHdWkV+MXZK96uAiWN
weVo8AyMVVnTRSl7GgyQmk8w+H/oHfD+TJQ2pMpGWKjwBqZylEYOzjdXpqfMVyjAYINSGtiNaVmF
0oyvfa6fFvryWNYpQEB+utnsGIjq2iAU6xKOTGWNHQkOVaRj0Ja0d7HA6eLGThMDdZdouwBA8CT3
QSoZEHM3hcx+3cn6Vc2W40Q7BT15DPhric0ZL7jfvbPPyvkoxSxXMRCX8FNp69PlYLQgxaPcosH5
SWsBCa0kD4LHB7+TxCoFoDNgKOcCbnIMKVuZ/i8EQHw2WJPD2dp0UbaF3lcPqLCLwkhvDmMBZH6h
dO58Itpqba1L9YZaTWn0eo+fYy3PIavAdHW+lVHRqcWvjsHtTNadJ0cO4m4IZctHHzCxD0/D9OFl
PVnMM+a20oKtvqWl/6dqHsI8XYhPF7FDyTZQAfpSPDCNazMRdf8yEpHOuX3u5EXSTllaQrbzpJ/o
oQCfD7jCiAsm+rqPiynrQT6P0VrS2bRiPL2i6vDfnI1orDS0W/Zog7drgrrAz7Ytr/VvmEnwAwPm
2LBTQ46793emXIbBVZ6UArnOAiALEV4gDXxcnA7cWJVItYR/If77mB4GGHg8c5z02khK5gW6zTFI
NCAQ7Jjx2J34J5MFtDMf0YTeh8Men1Q2zgrtSRQG8vgh3vywEDi8Yf7M0e/rOm2SizXxABsyvVrO
v/Q4deBeULD2buyJCCD5jurb5EAqbbhKaosifqZcgjroveI4ZMQYR2fgKDcYgDbbgjFWnFM7XSqU
+HEqKbngCJYR2tAPwdE3MwmIothxEcyh9zKrEGK21bIlMuXAWl7+ul9wdejcgkWfaVbtgXZr6YLh
l/v/Ix/ewSsSE5JIcjumONQdWStNLW30VqyB4uwNJoJtJNU3omd0IgLOoG1nDTVenH5gNJ0zkC9x
6NxpVVp+x+Stu4aKaTYh6alOvSzkLPJI7Ews03YARQNqU56RfUV5dGor3eJpPGvM2Zzg54qamAQm
46COg69C/+bdPI7if6xPppFmq1FsxNVuplRuLMOgjzgB8i77taEZYiztqyPFzQQuj1liATfLPmfY
hOWPtm92++PGzCu39hMJi8GZAreLVdBTzRm5XQ1MM790bKtj91ADw5OrxjpV618885fJ4UbXfInR
XzsD7z+9ks/Yzi2jYLY9wzRxli1IVFCVHj3qdo5UKI9l4xO/bNjzAUtXZ/IQmBDpkR7MIwn/X77b
n3q3Ft7zxACdvmkiXWwhuZH7q9xWXRQo+X9a+DHfdQ30a5hxV6+93TgFMxFS8OotMMdD03GMSoG+
F5BHIR0lRzR1HnzJ985hMLBe9v3kdyx950zRhk2KoiaxcJutjnurJuQcO3d8DryUp6g95v5jvtNz
3bLlo3LJ2Sr38wE8MOaNhSYu0Q6SltMqsSRM2wYAFnohCE3qwwWTfLqqaOTjWb7tFVWExNinbSUM
pkAQrR1zxqi/iHGCsoW15lRRzTnKTbzSI7YaDgwc7gKxWBtbbmAoCgXQevEVJexVR7ylLRno2v2C
n4bGvyAm1VG7/Cen8QD/gokcS6ZzDSUNElCuPHJrMzQP4RiGwzonkFUTV5Xd12GXOqK+cLqbxOm3
EtMw9DZL6qRq4ZGiFJgLB94s7pVSGAD1rWgFoiwJkXO43ZCpAE0tu2gwiOi1SCFoA0exfAhOAXFB
l/2Iio4N0+UU9yY0jJcMMuntPuoqa9VZXsMrCZq2yjJP+krsB7UuIvUz+dIxPpY/P92c9wmCwQ/0
oQauE6XLfiEIKQtYzzMNcNcq0eegBOmPcvTaz3HJcUtcjuxlTex+jasOq2qLWD/tkWaRluvF59Fr
H3vNGfqe84t8BlRA48JTIYl0WMBwpfppve3CvLiYjfJCoamRa3hnjMzhNpMLjszqatJDZJ7RQ+js
TrEGbVWkB8jfCQ3oCUjaa+SDomWmBdIkXvvNPbG2oFQf9xIaMboCc4nbIb0FyuSzeWx+2irblVW1
S+oVf14Ph2WlJdCx3qvCRXxfTBoK/O5gXJpJj8+UUQICZWtbY9Tdb807Lre1uGVASoGvvvze+NOO
VZMUb6sQ0IDRV9Y/75Hh65DHlxySzlWXOciKwVjPkqgWkttRU1LdpdQ+694+skcD7R5mxjDGN8ka
qdNCAbvb+YVAdGzlauux+jh/rtaQOY/Ct7PWLbCxZqZ6SSSY3nc6txyeu49IUiGUm5jTgM7yZ5jV
2sI8rhoudk6+Z/rbh+hol4u3QLKwXxU4egPZgX/iGioQXmRnB2v4z37TzsfQVYL1z4UWhzloq2MJ
BKTlY+qhxUuL0WRrkw9Wzxg2Rnwjgr8JlBymg2A9CKlllT81RTVNsWsOl49nJW6dDyGl1S63Z61W
fpfijev+noPBJHzLbaFGbHo8bcQ23w+e4D2j+1nBBnF+V6f3tggsham1MgGh85tIH7pwxt4ivEzs
gceUCxoTSHsppJKmOHanaYpYaAVdwc6tKXNZNASwA2uyvWNszYRKRAkO760OP5TPxyI664M/iTvz
sa2eQxEEr99w0Lx5FayL9vzS+bXeAqj6USom8a9nKckOkRFOirH1cEKK29zBBiGzqJINWmlWaFG/
XU0EtzwqPR6Hs+N8noTiy3y4xVIi3chaGu7xHR8xvsBXW4Waueemj+DT26Zvr4Waaf+JQcgzf8iX
Es8xbutvb3u/RVjJ8A2YglFNEUW+2HIGEbnzjnejFM4tRC8dDtCxmL2PhNsvteg9Tu8F78YlJoGg
eMlAdyCa8za1bp/VoSTSGexrvmmBFUuAb8buH7gYD96FWpTb2zHK+sIKVnicf2ibM2jhtJoTi67v
aOsutYAvoDahJGaphZZj7LvroiB8kjT9BDIGtYYElAoWpSvbhCwcMCe9kniveLrMSKEtA2ohl+4L
sZdUubM31Gy3I0SieWz4kYrzfnPuqMLTMANCs5jVfTdDzhqTxH5ilrB/THqa3MIH9GssyoRwEzpE
710a52K7W5/vpyFgcrDQo437rgN9+LaoivWO1+SxiuieYmDOONQtQjFtMZhyr5o8PNsqj6d4qxsQ
2nsC44qh/VNuQzVL40T615+/kxr01aFaQfCWVBQ0r3az5bQX2PVhxmxaJ6aMFfBdJ9Q2cWJcT+ch
KJUyME+wul/7m39tbE0OrDj5s3GaOgudUrStuTNnMvuBlDegv+YSvGzgtE1u6GfCQAuZoO8tPIEc
6pLN9hEZ/Ac5s52oMs6XxzAS+qm3WoLdIZ+ylTksnek30OIqgGUaAtkFQbEpdl2PIiDR9PuXLAy6
buc5Dk4aFnPg2GYd+sgnoTNfKvZp4wL5dXl1HuFU1/dsiOXQRqR+XObGOejRW1whJS08VYNmNF3S
dENfVNIr6VmGZ/qHeaQpT2MYFQxWqmJ0UBbzsLtU/+TG4BuAg+46kshwe6Sfgnpieafd7vARwCFf
5HUMt+54FX9O68GgTwIo3SFfcmU44NzBdWt2LcQOn6IdAbRYzMCcK3c1bKfnGcrCKIfEmA6IKcMp
qg4J7rLy90VZLQA6P5p2DiV9BgfOSHyzGugh5QvKIi65dw64Ti7ONE9dSCr6i/IB+R97/SIjuln+
PCNNE3LX0JtYCTGDybm8mP9TgRb8hUk9CebP9kcR9I6IFAE7pXwy/u0hFVAnu3jMPIlQTZOCwVza
7f4dQj8sN66oIgwRkDDK9eZAE1jjA+kOdZnctoVV5Pik9+8WXQh8odiNkOX3CojpJ/UjkBtjmfGG
wnudKQLHcJdKzX92JBYAt6Dmq0eHdeM80Bt6IIibRXArr//VcEPQG8NY8WJXRrKNekzmlKPjrSN8
FHQl/xdBENgF0I23IA7Usm7Y3toV7kRXxPhhsaHqRYlP0GfEnXF9jrMAtBXRNps7gzeDdAiq/XY6
+mEtE+4wcoYW4nPYB9gs1kXulF9PAByFgN1gNSYjhpZqRRapa2C/bLg8VxCEgIgkyhxERYw4wFAN
Jo5R+wUjOoaYznBVsev53PQ12HddikB9kyLGpGajunWvF9gehI2nsNeICj+lJ7jCLnbN29na2Q73
l7jWRRgDddetz64N1GXQ2u+6J0LM9HFArh3TqSgdYZuxPyZALvvzYNNO7g9BKDtzUYV2gf9/jVUe
tJ9ItRCouRyVYS47jFURTX6BOETIqJdyduwc0c7iki2Pq4s26UoyL0LdjqdGpQOfKEp2JALZ7qP7
Q0/OyalGp3bm8c1fG85pY+4YCxmSZ9WRkbROHWirhotY/KW/JXu+P1cebqgmFK4fKmSB/0AF32Xi
nC5SltiFvtna5XnIWHHS2mvmV14ddp+yU78ubtos222TtqeUDKQ+y8xoGV2aFUyRGDEvbFyteXvm
O6GErkmSpRN+rCwv0uJAn+2YnzLbPP85YTJ48Y4Z99spdOg/nVEWm8VBmHW3JUiu63joIZRrCak4
WRkDEKXF5Zwymt5BeqXUHxq8vhGove3RJIxAAA9VTE3kOEwHDddorfY7ItuAbmzq7RXM/PRRjcPb
Nks2uTu6PcNH1tlLF1ngeXGGNBdb6uvhddfB9vVfZgi6VqbqTD5xQtTLTasgO75BVdXuRK2wnyYi
SBqVCjzMkUuv0nVgeqmHdHFTEnU5YVYi6NfiJPx/z+m2O2YVLG1Tsr81UUYDEdYyRNdxs8fn8M2G
ng6CHyPA6ApLZ9LwiFa+KS5V6qCFg4Qxfyol3WZdhWv5ViAspNj5GPCdcfMU5Q+2X6A6YbEw73BA
bOc+3m+W2sJxfVaEZm3Njrp0djHFh132a0haEWpoBtyMk33n4mP+/p/YeR/98PS4i8C7HPrMqfJK
p91BQraFYtA2oC/2Dhf6PNlY6CaSHFKf+Ab2Ng11h0nl57qkSMa0szbpwIhS/ePAKh0RT6j6ct8d
ANR+ya7gxPWPyuoZXmv+wf1XhazSBbKE6xj7SfIwgjWrDzMp6R3dJa9rRYLOm7c/WKlqZFYZiGkW
09zNRuubdA0DKh+yTTDJtQrHON0dWpthIUWNtOtCIGBhk23QCGAuGkX6JxsIHuCsC6PKDDUidR7d
2l3nbZKBjkl09UmxHavNMyxJZEAzqARo6ZAzWKe4p3yBiYrF7Qy0uq91wxt+cOVFpKPzhXYf1rla
nenVJ3Fh17Mj3tiydJkdFWI2nfhRGMyyKj7Buj/GQzoSLdl1ov5brrHKfiimzSmkXzJF8wAJZ5OJ
0KeJUG80LemmWM5LC/yWiL5BgvGgmtu6fFZNWzGX2gpUtedKjwa2aLuCP3q7oKZ5f6X3RMmojFIS
/rq/iXIWDrfTkIz+vT+Dw799jh66jI6aSXnGUcbx1Y9y/6fWZ/F8H2B02CjkB1Zj9X2TEPZ70qNW
xwAREryY7xgKMa3TGMof0G45u8IP6I0KUPusKyqpaQyHgpEXKYOtTQ+6/DCKYPXzZs/nSPeCr8ZE
GBXEXdadVXDJMhVEoi0sQW1cotVQMrm/mzQo32v4NJOijG0T4wKiPDuONBK2SBahU1YePeQV93U0
fsLqLMILpQTVRDOSOlS8zLNspI9nztVGDNRR5a/Ltzjmj7Ci2ih6DkTQqs+tv9Af+Y8MoGB73j0j
kmW7y+1nB34/uEwm83YtQbwGd4/XcVVJvwI+zZ4qhonQWYpsfkvO5XrXWVG/GiUyzWRMC+TTR9aP
P4auArQDLB+aFQbqbRqYN6lxxpdvZ9FInTiVOO02qWz++Zni4K65ddElSRcrkClPpMHknAG58oYv
yTCZYcoXhPuc9wEvKA5w3VaqjGBUDYDdvbRypF6QhGkHFCajQVTmtCu0papbVQaukn5+CWHlkH0Q
OLjYieQ/4iH0haHPyS3RnvxEhATVDcY3HMnsdSCt7LWLKEYrAv3c6pTRTknc/wb3Ha2gNqQ2HDRz
ozWJG1l2kzXJ3phP3HgA76QYDCH2owWsov4/ndZV1Cps+mu5wHAtsUuihqVQLvx74qxKcbKgFLhF
UWF8ve4WqzX0yytbaSSWPQZnV38h7izvj1Vc1o6AcM+qVARmcTt0UvGQZ1tWWr9pLj5RN7+bJtWJ
ukYrCws8hG9wqopi8Bp1fzGd2K2l+h5003LQGmMWxJ9QooCFvft89sivZhyHMUD4+qZSyyf9ogqy
BwNENNYAtSzYDRB9IETYijwzg19tT8tEued6L2Lx3nAJoSz1+xnw39ak2xTN7+x6GoWvtszysT7g
iyYnFTbwlXxMQgLIi/uCws1TpJNgPKuuRoWwercOU6Sbek5k+ND1f+voJ6E8aNbdE33/xMaKQc8k
2NShRg34/HXult9hFI2xbpxzsNzoS37/tMAmfyxLXdUdT2NYO74vY+YXKEzq440ui3pQOGkgA1FQ
etJT5xn8SuUbLyn7HPMrl5wWDNo6U2aO56kHvn9D6HcmEhvH8wHzJL3kEEVjMuN83z/de8BVp70y
jiDkj7KFjwcwHAxskq62pgTm7bvB+5p1bYNwy+uZ6AVfVUUdQDkhd7hZSTwC2GbvxDJt0+vLBvUu
tXs1geWmGMtcBQo2epXe443okq98E96B852bKaixZL2txmfbQFGqTuScGhg9zOOKNXKZhC+KYgNL
/CU9ykRFpGv2MZUZdQv3SH1/qXcAcEK0ULuJMuAwKRwdnCDlV74jWdcjiexxIELkrMMPiPotwmSK
eE5nZFGz41v+I5+FzlFOOnYjtueLZaFcKxlIejYv/SLZ0anxwhTb12eMpU5EycYYJv+qLFMNaPmr
2shzk3ag7acVO+35I/qVpf3HREfOXw+Vo1NUOECFdjK2ATxaUkSV7dMVcYtYHUkrpszkjUiEMSF5
8QBDvt9MBup0vd4wb+Wubt9w4DPH+YPkISF4C/x9xjHODj2DftGyklXPZLXlm14S91gmacQV/bgI
Gp75kvBJp8Ycbm+nzlO9OERaeG6YW+tSczNipBdWNMewhqcbQsKCvRZwt0eIe2ar2AQsGurrTQ4J
Qb2Zl5n14ybTtDKLlgGb/gkVyCjsJhhm56hDswWhHVvCTwFz9lbUY2T15roH5ZfAwF8r+cdxD7mQ
W31TBOo+z3yGK6OpP1uySaDQhanKRT+qWvU3TPzX7GvWEJSlU/SZCO4xXFwU9Ks52jcU7WDy9/BC
/1QbL1sAGdPJkELIbqUU1xCsO9vAx6bCNKsJTQJSy76mji0gjJNADpWysuctn+E6r8DqyAGNmKFw
LlYV/7lGPt+An767FuZD0O6Bp1ZBDqds+ZHqCF+59K1NtznIhfdEJ2Q0wjBI83xeKkO1oLvgbTD6
2MPvMprec1xuEA7lphr2GNAI1/d66WBt/qiNFacJAWF0HeF7C7YGkP3TqUqY7MagQEbD5Ua/XrT0
k2rHTHJYhNO0sP6bXTRXEF1mqjO3A3sjoLFMwBjkfxlGByHt+CUm6ku2tCvNLJQYRhwfbgEbOlPM
uyDuYZf3kD1SseswXzjmWSXNaZn4tKpoE34ZzEOG7igO92VDAoq6fEsxVfumg+Oxl7ne1PBAAJxJ
D48v5VKj+IDhDecWA+9p7BO5s1RuNThNW8B9R8rxQsFateHUwTxzIQqU/GPWT7Px4BQ/58kHsDON
hDZpf9Uf2itb6HdsPE7YkxDpfEMxFDS3fCtkErOPFuYrTU9HqfOYT6dCocjUhFJuPxw5KCGhr0q1
MAk7m17zh2Jvpu1TGBS5uD7gts1rmLJ0yiXsiq49nbZhBf0fXznjbFbvtxc52ZDkZSN9nLFUGhU/
US3qHL+AwCRfATusw66ZUl49AC0Bd2ei75V6tOgn2X3Ti/JwKWNkH7awv61gE3fGUxD9ZFWjZWgl
PELzwvCNNisH6/tqkqwYuSaLuxNc+2otUwViDsPSXJoc2UhWakNe6nBEWEdfZ18yzL1nOikf0e2v
SFP1KiEoAdiCfvQNUArR80FX3VeD/6gLV3CrybZgr1WAzINr/DsMusnFotKrNI2ipcZZx7tjQKKw
TLX9MDSyAhtK8Av3Aoa8FAQrvAafEQywAdmPAaCtTujydz+mDDAaQxlz/agbfveT9L/733U5mdNW
GkPtpAas9ualZHv8lWyb0TvdO6VYsF2HczZrhp7BNyFCrLMhoRzpof8pn3vS1HhWS1/T82J5w11m
sr/ZL5hu9W6IKAWnbf7wKBCPJJbjLx4wyqHNSCP+z3s4FYzhl0CJHZIkurzo4hIoseOKR4bYiWRc
enCe/Ld1NZfmbGQ7shfrT6v6adW2Oi3l0mahf3vu1zaoRZ2FAaVX8wqvQGRgdCSJvvzYOIF38A7n
LsoKHKnHndDb25YEQm5L4d8yWxr+sd1uNqJExAMwxc1colTKhoKqMc0CzpYu7256QzUsj5DQCWln
ugC9EUOfPfodEMmE2jnqz+sxJXl6Tx5c4Z/5QuCxpqFG/MOq0kMV5b0+w1I7WgVZPYZDb4vUmOVU
GR/md9ZaH80CLEnKUzBEE9cDJOKv3QGrD8eEkHgo9h3wMwbuWQR9D26uG9Fny21J6jzgM/SVTfK9
LVOaql+x8HzdDSXnx4OkI61GZ7b50g91SbsJx98tX+CvyZC4Oou7LW6h0HtgJmmfm7+5P3svAbxR
1BpMDaUiKEB6YZ8M00JLheVek5UIzPvX3qrzwAm1ALHHtEb8supFof8+CIl2VAI5PQVYWTcivHqX
bMpWnA2mAb4sNm1dJH6X9s5M08pzHjmdpFK6c1K7kmOA1ygVOmN5dNPbkJEoRN0mgwMSHWi4lAQ+
e+uiT6CmVWRYp8bHCjzHKkVvzDz1LXy0g6+FOPK4Qp7jW6liWbJ4k/3QIOlmwlROG84xbdiHN/rx
aBGUh5TIzpmsp+ZfxEgrexKuH8cp+AkDoR9DYLxs+BZ2vPyazkIw5IyHbuAt5l2yY6PMzqzpm/on
vRJtse2hlLuy88ciYADKAb4ZcRs9R3YhtcFaTn6j0UCbB35tiY+UW7S5I/v3nGzyyKsDkz15rHvA
Y2YTHH/XX+z7XeqZsk+Y8mZZ8Kvs9gjBTi6162fWnLCjIOLZGEdPMRz/Nj8ENqhC/520uB1i7yy2
XUx/clD4V2Uh69tWt1KnTZHz5D3JOf9OVyLqqWvojpAHv92jIYr+rKIF0u4303Yc2oxZOBa0hEiZ
aX31eO8e6nN8DC7j+FlCCWRKJwrOCbrVl/ZYNz6VZx3f0eUDPzcHSDL60F01owZ/Gu0DlmDRI006
I9MpX5Ia0b0BhpW9eNOJvyoiWO97VCCBvbnzZO+B8doMt6V76HzNSERicxpL2pajE+se8jqwr6HH
gK3BLQqyHxqnzHhkdUp7aVSOxoHVmgBHffEgb8D0Ly2pkFNrVK0q+nZLkf/6H8fRpui/P1VFcxNN
nWWUvpxi1NsWIN18TV4/9tw+K4G+Lje+ngWb1B6oxHwz7YxFM4l27h963CR/Ny0zQC7lP4mtSHOW
+ZRlc34ax22arQVgdGAAzDSmDezbVyjGSJuckkKkj0CEcEtSid2afX8uparQTPZppXMfxWTNm3pu
9YEUvUs2bEDYxFjneOeTTNGIvUcjr4Zj26py9BMeFMr/VM1WFZT9+j0L/hSNReC3ey8SIkR+Nmym
xg3iY+ePTBn5l1MvQaFXqm4xF2eZrwvLmMS5BsjatZaHHGsRAp8/Wq/mIpg4tT22sX5ixm70BMwb
bupLbFsao2TTAFbf5r+DmGGEohSN7IUytvTSJR8LVgu+PwzSw5GJeZ3Bw5RXvoqXnyKBdBBpzMo8
SccSNo+CUp45kdvVdID7Njd2ODv9Fbrs5dUTKbADXrctIguLsuL8gqU6koXDS+BI3MwU/f8xqm0Y
ekhN8fmgWiYLQiYHqO/JDYP0592zjFmYlvtO2p8vRu6M19iOZDarxG6Zgr6fjegaAss6NFYNuD30
5euFQg8NL1JWwtpA4n7pHJgWtOoj5g2abq6nIEY2s7sURsgvqsFZVccdyv3fmXBkTHCtRgcfQe4e
Zd7tLpe7+52kZ3glK9I4inVqk+KMy6XC4sOBrhdZAIDTBQiCkIKfsi2xVFKmQjGJeDg/teWbo6fa
4Xe72FNrS6IVURBpnwoXpl5diSk+iDRX6ucySVFXm/Ezu8f5CVSyZ8n5kYmlOpP/0Nm8hQq8isZq
oQGh0m/FM4B3Zj3rWI53f8YvDESa7iBelb1MW8JtbIAztWueBIoazxn9X8y2nvdxXvz5Mqm5bps0
Or7JqdN7ox/w35xheRHs3gbdWcOQHyvJaFNG9PngyxlQUrBwmMMgem16orF0YJKQd/20KhYTbv8U
28RSD7ZmwVIt2vrG0Au5rFnfqnMNvzGD30hkKBhUCai4lCtEwya5lGHLkFam+GDqvb4eSmgtHb8C
asCZzsHJmZnnjOMKxRggj3PGxbLpoDKxVsjNyLZ7B1mQykItaNXWU/t4PkOqXyaJDbsbmvtdtq7a
Y8wQ8QU+PP5OJRm4014Q/SLCPtFq5I1bJOmehWxIEiOzylgFEnShgbQyihqFGX+mF+GFWq6yQ7gY
ylDIBZs1FCieYt1jpBiMvzSu5cotWy8kJMGjGrTuORljXVx5gRwo15LMfYKr09iBBPT99IShO7D6
vmJ6dcRIzW9w+7MnVcatGLujaaUOsptaE9MLSz/fz3IxY2RsTPVSztLkGqoq+us5S742JlRsCOd5
0ntb4m6CkIZsE8nyaiKiQVNcdwapR6KfSTWD/EQc50dcOfvYNmLqWXnic7rdEr3WLd7BZtyT7X6O
nd+ztRayJ2VpYR1pFKhY6KV5A5GQGiO9pcN3w2d6joMpBy3XYZx8VbA/mKgEeyNOp8YuKurZqLYs
e9hLe6Ey29anCdlGqNcpNeIUigh4SJ8lEiIKSW8g9IQKXy5CdpGV5rSwxDYZSe/Mwb2Xr4VCFG2u
a0MCZZAMMbNBudMfNBqkR3eGZA/GZOgHGw7TI007BPSr34SkYolQU8BfYcdSuZrSGeoHTWXzWDOc
mYIOOQiJ58y3YG3U5iTWE4MIgsxr8STK5Kp/uAB9ECPh1Lls0l4Ki52PpPayLHehWZrX+COTveyb
uBL2aM/m7jiGdsj5WvpaG8KF0Ktgal4u+yGnTJoJ63xdhDCqHTPq/YvDEHu0KPTN3s5VotAG/+Ei
f3/+P3vE8PeRP48jxyip2ordjws3F3dc6b83nNQKI0nJAXjjnjeHxA+gGceKUngB7G3fZpU1mYzK
+8lQ7oL/spJ+Msj8QD3Mjx8r82z/x8Qda7lRnlQGwvot0Fz/g1oWq+7uu0BrPIeY+rP1fOkseEEx
OeOSoo4EPDMdzGAZP5D71xNbl8F8o2PSHzSCk+EUwnSNSeWAsOwLUj+EXq4yGwtA2ZMxuCTvlXxP
Dy9G9L22idKBpuQkQYQz0FPioO1iSiyUxNAInWJGQ6/L5wd2gbDNddEr5Nzncj8oT17Pyabg561j
I4uRHUfddOnCe5HAkQfzQUYI4YTVoU6dsTNKEfs9ikvGoD2eQOYoemy/L33JPnURqlBcMsE578UW
H8lxx00XbqAqjbR97jUx+7x1u6cIdodxH5gkaKpCjpp8Q0tFKKSOjIpK5xXq3I4+kbOYof/+1gj4
MslVKcIAx0+MHa3Hv3mV1LG+DQIAWT1QnuVXl2Hmf2CgLZiwrBBWqq/DdCAn1a6PSE1y5pBmPjzJ
Rgeotpm4bjJ+OfaUqWSc0j96xzGrzjYDmNsUGUtlCP3TwUhbqIsjhbqJJdLglUoR5KRyNRid8qMv
Y1pG9O4MFgE12pw2lyuj3fqc0TMYncOvjjoKxRVUVW0Yx8eY//rhZr3vQbsaREa/YwhsJQ3A3C05
BMMGCC2tdguykINSeHH4l7me3L+3yNftiLAaHnaRKKuqIZd4W46BO7WMS4YfNC0t+BkndM99CBuU
LKT38sI5nJa76gg/AeujkEMQCzKhtBO83+4ZRXlUHVb2Hi2Tf8DJAVHpPy5EDQghlTgXO0NdubTY
miSlRAWvTKkYCvj1cFNv/weTmz4kd4VKaajT8sfj6U4NWm2fiLuZVJmvIvcCQoxApQntFPvNW70v
DAGtANGYW5WYS9AxUzxhQlsO5AJa6p7i7m+8hPyzXg8OI1Y9myUNoWdL1OBH45l0Cd3rhJJJA9jh
v7y0Hqm+iEdWT2YRLegMclblpBO/3RKsmtAnfKD9UAqS90HFGBoN2oyV51jaRm0qOK9VmC3pKaQI
/pb0BYkNvRWPDVAjTrMvc6155SdSV98djjReajaaBYiMd7FT4TUqFjB0vwqK3Ylgk6ZNveYniBh0
Wt+1v57mNMjhHfL/Rz3P/tqYO259KReRimyJNIDDWb8z+cH8nSpQgTxiz0D6n9VTYf3ZnDhS1IbY
acb0GylkbqyqhcKVKsUPKXKMCAVKHCJH6OUJs6Ec4LQ8OPsVxNk+QDVBTlSqABmBbB0t4WRRKd9G
M3IXMsUWzVrs0J4z8bePcJiK+KMDwlql1Y+WUXe2NasnNOelMhQl/8TQLirQsI7CyR28tWyc6fEd
grl58HLeRgPShUDaTDvLgz6o6LiT1Qi9AcuoI1FvYeYNNiJfb7Jww0NdkcyVcsXo+lwnbRF8ISDD
7NQrpTVnvEZ0YVJVfYgg/YWJgLuq2JYf3I9S4iDfRk41rCTJkLd+ZxSeq4nIaTa2988nvt6CLNbU
psGBckE1ynZnKeCsYhFIJ5SaS8o0AkcjKXZj+ywKLV58JARI8jnXSVhbYWwsMXlkY5Onm6liorUB
B0FD4CpJwXnexGYQhpc9tNriTwLGR1W3PPUdDFAIQoPCmBPCVg3ZdP1dHuCQTrZN4sfyupJlKVQD
9MXcrENr3OxchBu2tT8lS9XWKxldB6cTCdQPAoQWKoS0FNmZw71bYRLyh41O9uo+zYlie8T07yJh
P8ewvc69IEm4dSg/2tdn2+L/t9QJhB6vuF2R0tj0yJmMfQznuHYWexCCKbBPiXlb5A1dpijvDPqY
Xny3CZ/iJfJyrCNWCOG2y4hFjitFj5UZyYDvXqxX08SAibrWCJRAZjSCN/Q3rkntputYkKgHcmrq
5mbMq6RR5+jKsocDnWqUDi5xUyPT5GDBKZ3NIELMbKYAFZL4hD0OCEd1jenjEHOcipTPhoeAnO3t
RVj8pQd1q4kkYpvjQbYC4IpzdWt7U4VcWhEsfXHcAo8u7zHX7iqGI6FtkfkGzkIgODHap6Sclz/w
TFp99fIciqiDQNBwazzofo4xfLxC5MH0Zrp7Ce68xLaYDE0O5XWYNVF3/TiKMl/JYEtUUzYf6OWf
IsQooCZNzQvDhlAaKQNOoUvVMAHpPLyDNANqWN7Xl1keUT4ADz2NN31N+o7tgUSrYnCxVy3WLbg0
Xe3yi2KW3V3yt0J0yqzHrgac8Yo0K9/hnaplJo37yPWOTIo8vsUvyD61h/h5Yn9G3jgTIrTCObIe
UarD8uJVX8VrkFirmXpO0+5MzSqnXXI1ORNrcF+KLfdW1iCV3eVr0YCBGHgmDs7OT5FMraKkbiKu
QkgkX4HKWm0UCr3hufkL+wQ9veqjA96ZDS2gGwoFHQ4dMkN50apfoxlcpCjNCwqzp3XfeHq4ugmh
KhoCtxHCi2L6CL9j+P14zxNHyQLTlUM2brudPfrvVJcL7GtYi9PzZZBo5gtsjRST0dBjTqhGGvF5
ieDZIzYmQJE1yKad6K6y9fFaahA7qgPAI6AS1WG4VX+JhyChSN0ZKjxVwiT6J9LDlM+u7CaNxc7z
r0SED/4yxc8CNIFApNTFhMXabxvsWaX3KmPSl0JnV5gigiCww89iT/P8RK0TjwyjGB9Aq64yIUvi
OWnCDELBr+jdrvnXXS2s1vUewrffw3tO9tYRRUnWQwaiduDQO7BKNtqXjD9/paCF8jfRakgXTyMm
2C5m1Kr6iqvTZGhDbJMiWEjpJf8yM/qU2SQlmNIJBH9v1MRMdrrPknou6+Po+UfcDj0MDlFEJBQn
u8aqZCNifFFMvsaDuMsrmO/c18yOC9f4zgtaex+ct/qNjhIZctxK+6q040fujK9rm3Hk8Ph6JU17
UPRfz5DMM6JgrFp1htdvMV+ywQFQE4EYRHGD79HLxkyecReaRWxwYkckFJvL8Ih5PrNqBbDleiV/
Jbi0M5MwR9a1yU0vLa7d3seIggMmEmGGZLTIbeBbBwgbYU4PO32WW8RVr033VbYU35HX5rf/MK9J
T1ZG8m3YDB66UoWYDmbUB0ofKnJ9EgXtXMTOtwy3VdFwjt0Qul32iJARV1Vnt29+ZgqgUkDeVgca
e7/EIWHs/jSjUERl3IELqsFGBddmRJ6yDMz7a5OFKb850g1erSsPLB79/b90ZzLCYpjKFSs4EeOs
GUHFIMz/aOdTLI+NZjkRiTlZ7kjWuteK7gBYz8mkAW5Y717vP9ieoy63ve2WBUpLXGmo+muqjDwR
zDLgnQLoTwz5HF5gucB/EX+vLAwaQEWX1UKChAcnqxhOnGogFe2ZAbDZPp4Ye0gAtNCeDZkB6atx
QiLubou6Ygv3sPZj++RbXIfm51DnSvJiMu9p9+TmjWW/1IeL6502vZpDhOlNRMhFyPK+wocoPxUn
EiF6exfyGnMRnKOxN05k2K6rCB5KLZcI2pGvbDP2DsFqFZiWA/RA+TeX0d0dFZ4KtezgwlVCqVao
SvXPWiAyMwKTkoOZeXUNgstu1zMGj0XocgcQgpaFal8CiCVD+UvjAEhZ+DZnoBum8zzaaPne1F1b
B6ziXqCNmvL2zSAUIxkHhhKq+GpxhFmW8LrwJwlCqUtXkaBy0tipgOySy2PYl6z9oNKMTVp7XCji
glYHhoyv0GMs4ehq9JteFfaHiFF1YVLSHv/8n9grUxiJ5Efm73e+FsMr39FO02z2dxzHdJ7x7RFQ
ptDA1U/eetQayTsneR9iesfy4zbfOeLKj5iPvPeKtwy4WlyJ1wRvmssD/8BMZHWmn4S9iWCrAyBM
Kq5bdnju9EKAYtmV1UEXK+Xpe7I5GYlugJTeR7R9V4O1tsP7qgmIc2B+0R8R4YFKJU1y57kfBJk/
nJdJvNtmVM+rvzf4g3n9nfs/FwkdnlvtZuQHjpOSCiXaxE+iHwYhMcEwdj7aB7L8Tx2XfkEnN+6T
mMbWbk9J9I1EHovs+B47rXtwRgAYlIU8mqOKi5uMVIbm+S+b9ksQp0nP2ak0JnRc3ftIUrfB+Hn4
P9AkqJODvX9qeuetH2Yr+ZDzBqVbp9lEQszmn0e2mmOKk5Uip/7avzXiY4WqfSZ25r2pRLM9iwaq
1fJuRjrKXqg0YdvnzPUXrd1XxnymGvAH4f6oHDd4O0w5RsGjBwwz411dCgnYpaThwyyhAcfWre2B
1lxK6mcbktfUAbjdFWE7YpjlsCv5rf0V49g7lzRpIxPcanYXvD98QUyUUnbl9SLOGo3YzbKU88KO
so1Us4UUpIPyxcSgA3AsftOuhucGoKcXGpGuzmy0lwyEmRyHnF3ssjaI/8RYS/rg7gF2DvK8S3RU
+XeSrLQmRCbMOC9fixbJUW8gjKHH1PW5co/eGoRDqUU6YhKYQyO5ILTl0dj+P7J5vR8YBSNBYowM
E9pFMVZUeqU1YA+c06YxZ1cgt7yjx2G2odwCIraMSvlUqm2V7i7htuGSN5WNKiwD26EMHCPEb9X+
EYGiVQe4mU42sNTk0S0WLfqtOxIMEiJv/qIJ3/CUkAaqr72g5rQ9oauiV6Lr9j5/XZYieWs6OVV1
mc/RyK0UG8a8BfOZP2ZODxjUMKnhbF/c3SIWuBik72TJSOwCBG6MMpIkTHV6gtciVup6eBe51nyr
hJDI2MQMkvfe0IYcBdyNFDcwNwt29ZfW1d1IFzGDx35WBKLYb44RjmGTTaM26uxQxO0ombJaoV1Q
8b2CuF1fue8LEZ+ONXYHQnorkREdUh3+e8dlXbipoPgVY+wO+b0sLvLvwfIbrQvLp2N0fmfLaOCx
XmjwJ0cUKyE6BS36F+XApDRimfUIWWXeJ73jyiv55bQUb31t7zp+lXQTtw9gonWXv1qMoZ9MQvOQ
Jxec7PXr8AgBTIeTYCs6B3zDpGOAzmV67BtXcO9pnY7BgLAavkkHIkjlk3yCiMZNMNZHb4Hy8wCx
ohNk+osrWMQBc8apVjgiV3bcbEgPvghHQDrnY3Y8F4EsHg3M+Ciq8ZvysLhNOdqEacFq6mPUBvuO
38mNqge9PasKtkK677fj09PCtneOiB9tJ6AjM6rwBqZcv3SL0OIMXMqa2INK6F0pW0Snd78jnNDI
YOu92Z8M+waBwbOTyRzLLDxX2KWnDvwqloJcVT9f6ZTUdduVT8B44zkYkoLSNFaT2Dcm8XPRIQrc
ou6uXi7CgxuPHQ02RrNMkpnpNl96wjLcpwUnEz+dApg2QaicEQFb+FiaQIPUxfzh79rKkimlO/t7
61wnRLJ64M6mzT8mbgfbLWU3Nuso60J1ZPOYllJTKTtfJgxRoZoV+nCNupNYBWb9wzUs16ho4Agi
IdfxfiLCizC6paFBtY2a5AIgDKxK5eZFGVr8qfSMTPsmOaPbjja2f7dV//pDw8hjdPcMUPRzsFb0
5L9YscSZcLXtW06AfHaR7mRCD/pZsK/diPXx7u05bwoZxzWaEHfqTlLTvShc81fu/UvxKGAluW22
5pGpl01I0B6IQvG/1jHbL8oQ8k+sSxt0Eo5SG4Uua4JEWp5978CTy/weynuSa/8+pYhFYdQ1MnTp
kTU5QS+BG37TBLufpRzLsFsE2WseHX1wzXRdK1EH7k/5q7YAbhCgk1mOPa0HXaJvAP/z5NMmFCAK
yEadtoSPpEDzbs2aebdjy3ZaDNu/rLYeLme7dbMqyxZCGQD72QiO+6ZOhh2PeapXZiVHe/B3oy7H
h+pgToiWCNyiyyL3vsaVIRbj9jF5IUXGJuA17c21WHsa6u+RL41Jyyh1EywmnYHaU4YAfoRSMgMv
6N3D/BhLND6/3uM08C5FNudDbPK8cgtdUp/IplywasXLsgsVx4cKkPWs1OMclZLzOtRMDqS7R5Fe
RSukxDdF/YCkh5Hb0FjfzrYhNJrpucJWTapPQrS/zHv7/lBs5Hm5NhJhkAPZ/8/wB+EeG9YHOr86
ndujaXH+f1yoZP2Vyc+2lnfIxcSO4hK64iiVodQ7raJMfx9arQ4+d248TX+rpLZGhYV9l6sktTfO
4dwgSNhE+8qjbyVW/VipOBPlxdqlz5M/dAc2YnwNLs6ja9ZLTTEOzbFyFO/seGH8bbxC2oksV63A
hbQcHL0HivGxboH6oLBdHanSS2Mj3Jwf92CxZEGMIrTRxutHEmR8aRMk3JMGe+ZtsOKzuPvCX65U
gRV+3fL4SI+2BYphlJPuefST3gzN+2uLr2PV1Sty9yiOSl8h1UOfTv4I+2OS3zVkSNeK0KyKagzh
LpXB2SQuHV+fbHOBQWs3KPfHUBsbMQ77r7yhdx+r/yY5xdguHggLAOU3cHXYrbDifL0SQ0QMUWXA
oM0RhzF88xNbBluUz3CzMpMamBZ4QwgXDlbIR2+W4MG2f2fyb/ZBaveqefRUlofN7Gyz5Tc9de/A
8c1cCnYPngAdLfwUMDCAuRtSK6fd2s+amN15W3dq1FPE5fxAHmou+f3GH/ufj4X8Oi6TBeduN3hd
i+hQZfutim4SjSEbubbQrE3Hi2+v5eyyzQDFyIVnxmhKtcL3R0z3p/FQO/QsYsfrQEcuD1S75QOo
8YVfOZdaXMM9kYbLXzR+3PVm60VG3LNOsUEOmf7GNOsSdZogbsPE9h+TvXWAK/TwL6bAjIfPhqUS
f43bhsBoj/gnjUyQf9ZsWfk7kjTb1Jf2By3conFRBCJyZch65k0cZZSRjzgyPQ9bARXPKErhU2ZK
JrwBmOJkDE6Oh5+5xL+MOkkJCNkxovFPA2azK7dL947QmNaovMQ7x5lQfr5UD03P3BwBaPEI4nXM
TP1MN/hLFLBINKdwgFVW7ffF35OMZ8NMprN385hQys23rgZbkNaAZK1Lmr8pkEhIQBQ0VSAq9Pxo
oLmsRtZx8ODBIOpLlpoQJ3WOhIz98PUpPgMf4jXoJRX33vHDBcGdjhQFigwxrmglAizsvczN0UTX
Z0MrQjDUap7RreKDTRgblLeGPYa5xKpRhlpUwG1GmNTyZXpT8RGkbafhJUnCr8cqcXnf+xw9uod6
d50REzeQdhJEpTrpcCqnLQRMLrAvO+y4eDJik7EGa26OgI7d117koLaOUQCi7fN7PksFVv4wsT67
aL8wdCHHxzOrLYKUWbf68FvNQNAQXtovGdBh2usR9OK9wZ4G2o66/6I1zBo/qz/Bi0zOwRN5CGUm
8pI2DrW7PN3kyz8I8ZfBBFu7l3Tip7EmQpiwxrseTjZWih23qxASdbos+gafEWP5PovtCt43OkeN
EBFitZZRtr0aMdZbnWCEsTcWI1tCgt28rh/l7jkQcoLPvFLcfEiWctcA3URATMdcTdZWvfhMICTj
ySyQ9yTAaK1uu38YpAo2SeLRrPq66LKCMnNCu3lUuEcdpablZF03Da9M88U1hmxmePT9+trjcNHU
eFFGJNoAwflLn/NEQz3oh+QdvtwEM89xSZpYjUPT/Mzgk59T2t17Wz3oaFqMFU+PCqu2JIKvSJ9t
XXWFttSzPJ1fKhi1LUnFnCyucm8VE45u68le6iOF/1YJcGakMsyECziHJSuhuRao4XgvodiLTDEa
9Yz1vdrvU/jORA4YWN346yVl1wrs6DOLPnDnxSvV4AlchwAk3/ByA1ZLUdM/x2wFynZ2UKzubG/U
J493/LSiqLI15bNRAFE5VlH/g+UkCCK8Lmnb8+/8XZWdn6Ud7Pxa4xPyepr3ePpxfVNPgo4kLR8Z
RXVD9wTv7tG36zKnUtG2CfJ08U0E2OiWWm8qCgLX0DJjSy8mfROi4TbFdd/gsRho24qJJdkhaVcQ
PAQYiFwVG5rQV0mpxkkwe7U9glojceUV9IvjbpOKmTu4Y071ddX5a+qG3FnCcgAfHSL1Cxou45IR
AINxqHzBIHeA9ETL/9qxNTie5cHe/+HViCvFdxQ/bZNfetSMSySpLwbYLeEEfgLTz2ncYH2pVXJr
wtmKJdrMZRcW6Anx4XrIwPXJtNKBqb0FTZDL5QpW1KZdM+w7Uczqj9rMxexXpB8a7tgGxQcao95h
p2cLBlWdxXpSyEPBn95+druGNw1D1nwO+WmqHPqUXL/XxPV2lOP6YOpXprUhWf9MSMIWvv+RPyFb
3klxwXs9/xLxqpTW2yyuhrSSrK5hXH7vD7S2Jo4SgOo7Oqd8p8OuVjs3LL1yVfWg1pie47NjUHxU
RP2tx5czYwJNtqd39m+Pk5DW6Hhs6PWG63kfoAgO7byFP41puh0tUr8PDdtBBGB9gh4D+q93QIWD
M/QJF4HxpzT+K/Cpa+67Zj9OeGJ2LXvSC/INY+D8d+ucYU2kxRu9oSVEN+6E1AR/35nKAv2+gfUi
Nc9DLcBuvNyRoiwcBV3e5uhUyz9Lio+/rBERzgEantqZkM/f05KCFSTBMXSs/zYezttj1iLTz4op
9+Q0Q+n4HwJsnkiZg6nYEUMnwunk/cAKcFzCltT6VcfzmHtkBQ3K0YMK9VWN9Tt+T5RjqXwFC7iH
2FDtGoCljSnL1TRGAd16HidSKtK2eY2KPLpF50cIn8KIhZ4KLLyA7+zrf3Xs5ZhHgbEHSFjPgxqm
JilrAXlHuLzcuaxVJSHG8kMDi0LEtpU00ovLqZgUUyz8s4WAU77OIzm9S+Lnz4+AtjuH/KWU5Vy0
8EYZ+f2qh8HlLXZ2VAksTOPWGFW5Vsvrd5jJjfVZw/bWz6ZjYEW2n+aXKQ8wYEuwL9rengeJUJ3I
+tbON7V141ZILO7cPVzejltotUfgs086WWSJeYZTdz3RmNRxbqiI2Pt9uFaICHQmCpqbuOmDa0aP
xg2qG8dXjw2N7DALRLHuH8lkAG5aOdeIg2uLGLXnsw1SDPgywSRhAHh99gX48IQqqsWjprNN/uL8
e+RqG72kRs4h1rAuLt0Pl2mN/dmI3p8S2y83I5oItBWNTr+w5/PnaRT68K3Q62Nbl6bDBn07nZn6
t0kL8VOvFurBS97J9Xz04JtE4BB8mgAJ5xX9L6fK1dz8IhRfEPv9tViewTENXqxhhd0LGKU7e90c
/6zZsUnduZg3DZHWrsH/z0yed1rcGwkui0y/vkc+WyrLVfcHQpdCUoZuhtUctZsxnd7vOzXW6bdK
6SJna1eBBQAchK9oc8tf4yfBHDHLGfyuO/y9RoviDfXxATX1qzRLmlr0nSXg2u1B5FeSuGfyB1Bv
lbzlDAJQIDmn+ncwSh7SR4rAOH5wANgShsiIMCJRpcTLYKlzmQOzW+k+F9Jmmxj2OyeZkRkuuB+h
0RXVpP6gEUqq2xPd9Bt/G4pJFtU06qAnCNpPDI6+A7kcZVVaUO+TTW7sKr4iXhPg0NrKNmuiwWmj
4+lwrkpMKE9VzVf8UjMy/ac5Bq3qF4eWOHw2mDZNuXENMhSyNFh7ZOTfPafHngscB2CQ9lXdQGXZ
xULb1h5BgClrgkyQjRmNPHqNtOLVLM4B4r8qkuVFVI5Gg8p53cUYHFRAfyjzBh8mwZwuQiCCkusu
0kLVnY9sb0OPfRpaRO6QuS+ypfkVEG65O1eM6qzOp7bXGvTbgjYh3sz8ZEdkX7g+qJpVL0OxubB+
qMLWrVHQpq5qq1k06Lo+LB8G/xW3Bz9IMMcWDyvfFvlga3C4nyqtM73E1ciauS/Zo/VcjaiI4B96
UYAuhlcaTAGy/gmyLWqj1eDbMM+SslyP7+zxT8Il/CT5eZL/GSXpSQZJpKRyC1FA69SEFGJUHWwy
+IegMGPr87+2TLYW7oeSO+5GM0igT74oZuSso+kEUCjf4wyu4Bi697o0U1kwR2k7dUedIua2lQrl
ReX/8LLTNgjRae7lrSlO8T91KsqOJxsG0nsh7nHoS1MVzZSAm134omEBX3TdSB/LlZ6hu5u9v6Gk
DhJ+lZOJXBLA15LfHJgsr2JSJAvOyZ2J8+Oae2dbdmIJH9hb3YPFmx1KBRC6iHKnchIrD8ZfC1F8
voBHx55JMXwaLwSGO/rf2DF4OUiUNh1HZhtir3xRVW/40zettnRbCA+zBzQLHgv7q0DqWIdle15z
AesqeLVGVo6UlO6jmq/2MVfjxXEvXGtiIq0KDp8K5pQPXCNy5Sg8zJtKQwNn4I3P0aFGZUxnXVw2
ZyNY0WJp8NNwk5Fwf7QJ5KK4LM/PkaQdHhm3m7gVFQbr2g/Bp489kYeOdw779E83jNiyVygix9yy
z/8Vu2gsrEGUNh7sK3mNJO59Go38mSKsrXZZslm2A+jWxSJmyhoJWk2Th5ahID8A4qXa/fiH9w2X
LzNFBY70GFn6nKQGnNzmhAenKESQTtvk+PueC+vv1vt0vZeHYfxIkugJSezozfUHqA/hK0L6P+kw
9m0fg6h7dnrZYd2EdUzfS84oQ9brIZfsob2APqu9atfGXWs3T5T9hkh8UTt8PWi6rbw2siP7z9F2
msI3QzxUeEpS9qwMOoGsFfOg3olwKHENslfrZp8YcQ9AsQYecpMJK0ygT6Z3BGZqXGCRrF6D4Oa0
0fmSRwAdw8gy2jLAMf4C5o+BrpnGD1L9GimwbG8mF+hpAP+xX7iZ/yFXVuhr54U6Ng2q47hBVIm8
B6hbKM6gZMEsdk3WTSICGX8pc4MbvuN+d3YjV2K4rgRq2ies1gosH1/uRLld0YvWCwHDzcIpdxkS
jE+qHJA+7vWY5jsHVwmtf7j2Pb1MCMnW3nrg8DEbFUg+9eqBs5cF3Hc7pKuYzV+OVGJm+AasvmPv
Xsz3uhXk1AwV9KuTWwHjYi6qHklclpNT53g4iFxHBX1xCQiMbMhHP+weDr9PzMVSfrnjj5ArHTBM
udNZ7Gnn5w4lXcPo+wUhxRKGdx77NJ5ftQOpCyAAfegT2v9TGiEuyDhQwTJvoX4pc2GnnxmKBjZN
xy0XuUcg2lcgJJQDcpL6090z4QuWSgR5UHbrFv19eoPt42aygVphcBXmfWcUmMQU6ZbhHu7eNBJt
mPHT+1C5Dte6gqeyX8yQsyv8Hw31XZt52a9KsMM963qjkGAkT/FX5T4v4TZ67N04yyCvM2hoYEYO
TfVdhObESnGN00i+tRXTcDMRUkOMq1OYgchG+ywv7/HPeCkYcC4aIP0dFau6H31VdzMnAAw7mgoz
roZJVVk6FeThzgKyxI6zv1rRqb6wSY6o6GQdWMfcFqQRRye2ZL5e1BXAloJeYPZNDIdRlt8vLc10
2mFFfWiszrBkRiCE+ALs6JHLXRhH6vweyWX8AKZGT+VjJB/Ljjn54h5TbjpAJsLFMsZ3xcmAM3p5
2KoURhl432xbJ9jAok+RQzcZpQfJgaqWfv/TuJcrOHJNsZxjInfFQRGTEOn+24l3PyrPRWmFGlnP
2hlCvvLQZVEFeSdcFyXKekCM1yAIEk+V8mAY3N2FKbCUgD46Oi+AXbt+g/80w6gRUzutGQ+Mx3Gj
u1VQZWfrwUyNHkmUln0PDALZuNuyMePPx525AUjeFC4nImVH6YyY3YCEpAfDE9i6CTqHFFF8Rq/F
4T9k4S0ZGpPcCr9UDVT3E7myvZPkBOwarmr44EfZQhVFeNZ1SAm+jVTik2GkK9vzf/baS09rbEig
PLpZ2ZA37KLpBa8sUor1bB8f+1xrLVbwfgzzBuIp4bpHqpqXkGZg1AzVzMfJwFWNudBOsF3zdBYE
jUn9cDm8HBddVFMXOMktQkqaO2qW8h9f8WgPo+C5k4DH9e+8Txvn5zG/rBi9zxl2H83l7s52rdrK
IGy3p9+evZwmAiJ1DA4TsC7bAdEcAKRVnmcZube5rMMLgpAUnGia1qevY6u89wIHaV2hB24JOGY6
CYmqRuEGOPX54tOIJCuDagAvlS6kKIisy7Vh1mKrzvqkxziRGQid+Zze7+Xv9DShFcCTOCsPrr3V
o1Bj/CxRI53PkMSe8mvuBn35lVoWxv5Nf7rvS12d//bM+qD7aRY9xVNhX3A6xxHRjGWJWufg5TKL
FMjykRPaT4VDIrh9StlnnWZ3JVUFI6lw+2SK0HjVHiJKyiWLazt6vnKdmSzd5uOMxFRT3LlXfy34
jp7Ed3BBGe/klqFymYUCPZaODcE+qjwW0jwWAyBwD8GFRmRhOFD19fOYRVyRcmEgVyUut9MKmrBj
j0UGeuB7Cga6JQU20G/+FpWOn+DhiSgK6iX4WKs9vSpqW0tx5AD1ea+LJ6pbNSIb/kkHFYY3Pzhv
wz+3ieGkyHQrgJboO+hcu1jT4ucxJMllpy+qVCZRHQNRKcsCq25uD/psPSu15hPQsrG5d6X9q0gX
ejWuDQZrfJ85NusFffYyPlfiWZ2XIbeFm/qo6oUOotEWrJRyZ5Uj2/lYFG2Z2AgRjDWtEFMgEdN5
93kZr3umG35lx/2LUYdStM88xGfqhi1P14Yw0NzlWMuEAeYkhIlBwR82bGU260pGFRkiiP/rO3Rs
A3uIKGnMoJs04eVu/CHip7PfvLVWPv8FwMqb83Zcm4FNVCHHjUKbOdYpV73GwO8wZB35155ER6Fh
dlR3TBid8TLM4eZcqjE6HtSz0T2JZ3NSWHRyIvsuUF0/n4zfrK998mNHJBD9ZuDeszk92c3dsggu
SoejoDKNQpu1VuGl5EZ4Fh8KtSUdpi1vlVJ56Oe+EdaT+2mTB5r6IFEjgYIsg9veaThMopIzNtiF
/elxW5V1SJg5IhYKEX9PrH3Dkugrmjf/TR8mBFTDXDGV2yswDDPDCZy+rVa/2b14RD+CpV/9rqsj
YnXRlvXGdWk8WXiTK7pR56WMIXwM3sACR8sxGWVhn+M1lrceceVLAIk0vNsr5J9pxkqjv6e+OFxc
tKldNtm0wtjgwZdHWrrMXreAKJ/zn4/d9YXXn59rIELLKv+KFr3fb8aUFt9T7sXIVztxTTodYV7U
ghLvnfbJl/clwfVdjgMg8IVzC+8lhVpMdrt1PGYi7MstdgrYK4SziFVPtgGWbIlsZfNdXWQ/qfgg
kkPWyl7WgjX4DwUAFuaCWaZgyHUA3x/WjPFSEJDFrKcK6DuclK2pZ7HxnWrkSCDxuP+8+CIMfUtP
oOlIULmPfFW8uUnAM+QRm4YRfaCNtMlVn7vA0DFjmpbqeV25blgfFIaIUA/O88oc4A+NxPzRx4FJ
6dtSu9LBJmCluoESNMM4SfkZOMNJUnC/DvH4oMViQE57IFOkZB4hwjwHUmGuYAW+aufODVOacsAz
lE7HSjLDFO79q4RisHI8mR5qkqGRvRBUjF9q988s7aQj3qRrFXAW9hdAAyZxCX8Wa3UrdUeslEcW
e/t9SPil7ka6Cc8DQ1RlSSMy0mcVKNdTIsveM7eV89pPVKlSZTyY90nqdrY5ehIh2CSVHNeTyAFB
smxEfpXZQ8Y3HeYA22w/T9ek0ldJAyNYHbm0Eo4tdvKPFkQ9mvl+Nnz7DA5+0OZR0de2UkOb1QGk
ipqioQP8p/YX2IRSkVey/Lqr/X4fAfrriXowrFNl1VPvXh+MdJl5/E4Q/5ZlWAI6ZKwi6vx3yKzV
mCWclvkZUMhi0nt5K+2/bxtCZBUWvandRlpV4WUjK0KV07hgux2vx9Ld9t0t8kVClqpFGq8rhKMc
rzuSBCO9ioPp3GJkCmDjmJZhFR250ng44DLOGPJKBmxhQzvkQzJXz0HjYdiiiBr4gM0/5uXBwz/v
9nxg7iV10uB0Y9IvNhXEoi35ptb0U1l9V9UHmlB+3Mq//cqBtFuokN6GBHpbYU66itP2F1wv8xyE
SsWxpzH/qf2u7OJdz75f9VlWzecmcdjuN9eJoyIfLssDPocPwzsWH2cdsvbTBY/krkOFGV3xI9zi
SYb8TwoGlZjHtKe4DvCfyw6SMvmM5JR1YnBOwIbXIwjNCLbpCHuhuCuIc8AeJEU7+6dQ0Ihd8jpF
RHxyj9w54iiPiLozwu+TRTYTtBX9gG8D5DCkAKUjfqiWJPoYVqC9DhlHYWRQbp3cUpy14GD5B/Jf
ANUDfbzNCB31lvqv8OP0L1aUZINl+ewn7/5+0zWZpE62pdhkHb6KQAEvACmM+i03BroZ2uawPQHP
TSGQYweA+pfte3/x3pqsre4N0SbKwahs5Z+ppOP+zxznKeo0y/qU3Jl42EQiD3Maw2eviHOEWz/J
nCS1l8t6kwmbTiv/pOSoI07Cc4TXqLhQutwixXtr1MFWoACIIgJ59IcCC0MVpIcYd21wRp70HSje
DXougAL5385GzyVrMP7E65SChADk04MqoLSjdm572p/5sHeEpz34wyMydj3ZE5BXMKjM27H4ttue
BS7f4DiXKSZIdy8n5Jl7LaZ3DxSF2zFfYcYJAtVnh5mK/1IPFMrqw1ntiZ3f3U3aMG/J3ltmw4Wb
yqOHVJdi62hjgrChuO+PNXmnTFMHVs3B0+JYd85bpha5t9a5oL60+dIrurXsrOGDexl3qjarF3Ps
lz9f9qm6GtN5ji/cnnuiSyTSgW1Q/OjjoVKf7opnsajMo7K2FzYegEkVoqpnQSTBwB8VLAZwrC4b
hKhfm9oE7DpR4Y/47CaF4Vtz1+YmU+4Hzeir0Y9s1wJ9XM8gACRLsLXc2lUFZE2jRx6zkE21QNwO
TSKCmSKgAz4l6WEMUJHCyRpKieFew5lq1RxVuO7Whsw5gUXS+W+xcxYWc/o/jnOQYLm4otBViUJA
Jqb5MYAmQp16vN+inBdDE/ncHFXESu2AeKl6Zt/44z+MEcRYXjvKamqMywNdk9I9z9xUMtNgCfmV
cPEW23EVuBFs4y2RSoPZxgI9+iunuqslV3kyaYrh2zvIDoP6H4UfJoUe8VswNmETjFusF33Xvvkf
7+IRqb8WWhscJUy32LItyRE1+LMgrQCFHQIazDOcEVSYYjpaMAsecJ5xXF9iHLTr1bVvt6lRXzzo
cs4xOExBdjWXD025GWMVxTY2hf5fwG53fGu+I0Duq+vBp5+k0JZ5we+e+RTN1TASk63oeYlsPOAU
V0hS0Obc4wNPbQoEGVCjl7bjNGe+fda4VoKfTUc/cOBLKXWuF8FjlzNe5Wnbe7n+mZUnwh7NckED
zOT1Fg/Z0CeYQs/+6+rjI+TQ398dWDb8/9ia+wG3G3zqgXU4dQYNN7oGtgT/Ws7nsCGoshbB5G7a
Osz5zu3E+VxEWnHNhrgbgcnY7JoLahoHvyWg448m+Q8JqEyl5R6wjWK5mTgQ5pXMotjBLMdT7W33
ZzKIrkBmOnGCPt3SJukEst2vBzvwFQYXBx/aO8WYSrSXOKBzjo40HwwJgsieuRjRQQT4ctCNyczD
uwqae20BZxqvVuPfwJA/Y3tkFFCehPbEakcqH13iO+qFrLU4CDDJwK4Ft+mJBKuqHOqDGlGhcGui
oQBs33h3QDko4eSSUA3hA2GOrfpBJEjBcH2lrIQc8qxV0t1hw02YilYwTo/rLnMPcJkp2bs3AkjL
I3QE1jetEsYdeU96WmVlDwLWaObj04+Dod78/o/G0ZixnuOMgCGDbUIsDDYDmqshKBr6gNtpQZzk
Ov/Zk7ggSFiSuQryb37x1QLsqSoQwHddQNiDzDf191i6knn4lOgJW41pB1Av31g0dncsxtn4Yc0S
yUEom0c8bwkzhkimaGO7YAjryKGUfrfalXgA5GjNvwlvO/FsA7zKWaPE9MVtx2HCEWl0WjkUn9RC
gc9MRkTTyoHlTIgqiXJebGADDB+cxAlXxPbfINCGyTsHnJGpORib5uRDk5CsL1Vu60eIbyTgfFj+
1wnCGwfF53mCTbkhga9otlt11Jr18I8ar+8RlvDFExn8HOK89IhcYugdUAXf1hPLDPTD9JZota02
THw7yHu/16g5XVVXsxqPzJfzFsutM63uP2QRBzi3kh0P8lqCeCYe9oOSTF5YBEX/ipGp7Ie7ewdW
lL9QFAsbEMJ+AYwqh2j/sGYfqZ68DC4zLiP9u+D0JlKBbVeSxi7LSj+KsOM6vPKghMc0n/t+U3Wv
QR8d3w1XwWDYEkBvgALmpJMke8Qtzjuu27CHEVWdU5Hgq5YxeLB8zsYQ5qCJ4KwRF1bGos2urG5T
v82Q53KmMG2oq5Y5/aOFYl5ohB1BJx900zETuG4PaoWvAVYcoruHegCM4tCzUTSVFKdVsaHbm1U8
OaGN5VEJrXhLae7HC3qZ5fZmGpfn4876qxyehC9YF4X/EG4zmK2ZWk1WOENPwa5EwA94b3R3P03a
booS52r5CdRSf9OewAu6sd4Xe+RRM2LDClvHausqlGhiLRVDcmdi0VZ6I/VeUxm5cahZ8S8w4lpm
4Ngp+p3RZqp5EBxALph8dJLy7pTzQ1ty1ol46Z5i/zXRd5IEfjCF8U/BvfAYEnEQRNdjFXUw+CFd
Imv7lFTyVG0BLO68Nsln7pE3H5hm20lbPz0T6XsxFR5S6FalPPDqIcBlyikTLZjT8ey/2Z5kfPwl
GeitxnkiWnXMTu7RvijpRIKKALyLhM53Q1DhPNTdmlqtFsP/VfMIcozmuuRVBDhJwzTPqP9BV67M
Odqo/bnSMCGn4H5EGGIkpemfiFuD6fFlZfPxJOuY0YJszDR6RCWFeGKk8129apoNH7GG9o0pvCAv
3fIrvqKjTWpeumIcNtcZDhMu/inFyDjtjvsR11WF+jxQ8B/Jp062aIh/+uRe+6SYfBoAoOU3LDrQ
kFI4myuPUXv4opKLHraoyv2gAMuoJVm1WgxuiI0tijdUmpps1rmDz3clvrZWOloahLvw4VLPWf7H
vZ/AlsZ7xKbpr2e4G4gQQwKnSYuBFSe9fx0TF4Pyl2QUhzsP0veNOqazEvrrFdnkCly89KYw1SGw
tmadYSHFAeMsviDkdjVKbrnahXh1+R9th3Z5081l804/Ke2v6ajrOvMy4lxKMemBdYH5SBL0+iro
WgIC5T3/5KuCbmZRWR0x8I45paWglhG+GwncTDr3hrlAki1n88vjQsmHArpum0XYDxPgoHG6NdCX
0+R4VhgKzbJpJYm007nl4n5LZ9ehlSHKOZ8MdKqhVFkKNCK0YLSIc8MfNRNOp+UtVg6Pdwq5nr1u
kn1kmMbrrPSw8Kk7LoJMV+KhznSKXCwhq8xjcSD6PfT15jqIjvwBqx/CoTF5Zo7/DFVPvvVt/tdl
d+0lU5oKRVjAJ1YmCUgmPOpJjRLhn8HJSlMGv/A20eu13XcR4tYR8K4RIwY9ZeqedDqhJR3EQ4QE
11whY54Z1gJZRKTBPMrTB3L8ifhFCcksiz0Rb1ZNwxO7HRUJto1PuhFC4iaE/DUrGRPo7wu+qZbb
jrLjuG/Vtg6URIxF6Oxizccz8GAohVLxUA47XFgwIgvH+WOKl1NgQo2tQBuV86PfpgXWj2bHhXnp
DMp8iaBg2OMi3FbaQA4IrFIrzdu+evSNOihzznC1x9w6Qo2kxlvBhCMkLvSHK3N6PKAXn3l+fadj
vRhkTSBL9piz/mMlI8D/4zBR+byMcJCpkNjOxlnlQleNO5ff9CX9CjrtILTZaJ36sNBcMYQIrrXu
tMxtAMR+fNODwdNq8qb5eskVqjuUVed5QG9Cj4XC8cmzqpjfdPJoblfgJ+nVXGWkfftnSL5ITXV1
teIll6XH+3CwXreE8KC9HXVwFUNiKqK9Vgjcn/Px7gg6d2y1/VdjkvJ6obXFIX5XF5Wb5Qn/60Bs
1FPV4JM7SSDAbK6eDRu9I4TXmqt0xbGf1LvPRpr37wj9slSdZQp0fZrOUq59sM0bSlti7/En88gP
uFMthfl0WbBlMlWHfGGbjQiHQrqTOW/8/Cg1QATqZ4qbx50ft33Jy7vuE7Kx7008gkyiHT12roTK
iuzrsVeRI8UD6SpiFMeGviMMx4o4Zv8/b7+RE6s+/JaBDM+NijHLJtKs7kPBA7eVRaoOBfjZc9CT
tLYYGHdtPVljADohhP4Xia+7SNEJ8PXef2OIcPDLcXdNSXEN0l5xmda52mtuQls11gJTi/HUlUcZ
gmZzXDKBbWC97VOJbX87nrlgxxOwzo2x16oi0gjzqGCgxyijnx6dOVx2HiftoGoe6YGznj9OPswJ
srZLh4LBkTRc+plFMkh/VQ05I4/aBZDC08IZR7BZJTHk0vnFmY0jYWK+Aet5k4yqs0TDI0n50n18
BMh6x4323DKnvfdCxJfgzrViP2Z89sias+MSWGOc7LLvswcx8CA7GDCtDn1YwpiqC3UqYJuzIJUp
4r742xT3oNWPBjnhReqYHMnLVk56bsq2tddJYm1TYNPOWc1bm/JvsGkgGu8Lvks0AdU0nGyHOnad
Brk4vJa0s9mef0QtzBP0ELE6h/UrmbqaWHpWI8xd75J/0lEbzngRudRQ5UrTeZXagsaiaCDOpWCJ
QF5DJc1yTizitVxyUGoio5YmvGtr5iM1TRdRiUl2vm48UrgoZktCayKZhGi3ddRKSpS4pRAWAF/Z
tTFTCAqm7QlWNO6RU7BSQUUVf5hRZBuRLn4YglX9JHDAWHZfDE7/klhEgdvB+fFsIOEHUrDU27JM
YdxaMgCvudv4tmkmg3MDs11cDYLNu1VQGGBr+zc+fVpNQJzmlrLryCQCyY3UMD7ECY4BoRQyIxzV
ODOSIPEvnb8M/Z8mrthj6Ev8AyMV8KjAL8PmeWqYmcGPdLXt7qF227Ph2I/u2ux/DSKZPlczy2h9
KUi6SmfsBHEVUXZg/VhojUL0jmLlDgAbj8pO2zeL3x2RMaiwbLHdyR2Mvm7vYeOm+pZ7QZPoUB2F
xPp4fLM6Ew+oMPwYhbhVBsu+0lYh258BW9QILdGwCl/Y1j3jEyzwPdQnrziIAG7dqPIxOBiQmOla
UlmT/ygiSUO4RvngleMyMDBbJlnUoQFSL5u8svL2kxydjJ3R0L1Umltn/Kky0Jmtu41/o0sbK5AR
DlFfGg0V97vL1tlPPklNDSCpYqbcmn60/8rqx8SY1+L8+R/SqflvHF8gWlD9u28W5AAL2H1hNA/Q
jkMnBU5HKR/xuTojI3DGr7hAi8I41pQt312gh75/oL3ivVM01M1fv0aWOPuIyh9u6xRaxE+EFqdi
0IhOT4U4pA3Dhz1hgpaYCGY0IR1aC+WTg9PGwCnTuwFyaQmuEWBTM1ZmQAkzkBfOc/U6jCPWvNk7
66W91FCEvpo8JEh7vZJC1DcZICN7kZqZItmfFjGj2X7y+Iwa6PohqQtgN7uygVsm7N5Mu2Kwfq8t
IIrLxWG++py9A3bGYYpHy/IMvI0WKORv33fMJgGukG2hUsxDsolNj5mt+w5VmwRD2n2Upaj6ePQo
ELN8WzCy6Ir+gAR+ILA5vqZrS/SZKhdWgA+GwqrvwPhZUwmRH7EXbwA/NoI2AlW9ctKq7ExUOYjV
xEmDkR1LX4ueqW9ZZQkpUN8YBSOx53/ECreSwFlWw4GPqT87XM3YM+O6QRrnWsqQjAk84THpCwz1
p7NjsDXvXaXpmmu3mtX9+oOi9Niv3DDmahzAO8/mnrLc53exnhF4Ijw+oPOCsMDwScaOZyNJ4ly0
V5XdZzXGN5OsL9gBBZ835naUzGw9wMoHZhoXHnhoUEJL2xGZU7R0qIydACyTKBG1zprxYIYtudmT
jneAdDrf6PV5BdZFLBSbvvUN+PDitycs5tc61LHqwXK8FLyXQAQazYNzyV1MTd6h7LxHPvxG+B61
D/46iV6HPQaVSyKbfHtfe66jt46H4LCrq/w6AFrfSW85efSlUTWXDZrvHcOHF+UYYjIfYDLbiINI
qoa1VJ/heh9D8k4/5Rk6zhJPeIaRhCw+BJJChsOcerZKBsu3Vs6vKEpL1qTRLyerJp1mY80oO131
kcoCuAvW/Ttz5DqK+Ckg70JX1IDz8t3o1B0u1+lNFzqBW7nTDyfAXE/OlGQ3Vytm6cTpTKIxeTJ1
JxFw2bwg5bF+Wx3fY998HRqiDNS/r3/deotTNpGI9xQUYIoYsRW2TfGKEkYa+PUq7rcXNdKhlQCj
Sv7cf+05D4FZFrH3nxG8iXUZId6CkYGywJgsCV/xuclFmOwS9YpKzovwkcXvs6OeAw9AmjwWyaD6
xCY4km8V6wm8Vc3B0n4R8N2EeK05TmZehRpP4Hirx20tzWCMHVg8en89UaYaWnkJYUh72AqSz0Op
R7Q/IlJKhcK3mnpOLs4Mz7ada/STvMO9g0yVuAgBMHagLm+Z/u/GdnvGbT+YLVfke0KAELms23Tr
yetZFFkTg9re9UT7nsaLM1hYHTaqIlobUee/E1j3i2N4/P89ZdbKvxpqX+fhhCbe3uv4WNn1j+li
UbnTuTEkThduGa/pEo1gB1WEFy+ZHl05K9sEPf4HngfgHUJv58lhFnA5sd5e9Fv3Erzl7cWenwjW
X+ErlOYh1fUSkma9BZ45z4bu7hA4Ynaconqdgqh4/DcBAbZt5rWISWk1ym+W/iotfgh4tHUsYyDc
I8zMiQBQv8HXfgBJ8FcVabE1Mdgy4L4WMMlclGZHLSBE11F2GEtqh/dIyPUVlV/VA+8sZPT1jIs7
o+8nFvH7O9uE7SjQBjttAvFRm+K1B6Y6cSVioXgYQeS/JB+eHvn9QgL7aeS05aPaq8+Vw3DXw00X
gBMqrH6tWy+Sff5cQKVX6o674YmoWkcN4sKYoyuuXW/Jc4FcZ4Tnx/m1HHFzpiJmyjso3mdOjAmP
dJjAiFQ7C9wNb37g6crNohx4+ONxrto0CejXCfhJKRS4XlhB13Aig25aIWtHZHTkRSCGClirQMDP
nxSv644G8Zbfy5mDaoK+TCGMZpCsiatNUJRrJzqvMbtSlWKdEEkNCHiVaTfUQDtpzayuMleZRKb4
71EykIaU8A/pNUtDjLHAjSqik70ZzguP8vAbow53e43CXZ771558jxXJzTkyedUkX8zGy2BRNrJ4
HvWZdXbZIRVjtEeJ6gt+xjkkqF28paozsTzcBAxy8pezmaJDigCf/zUg0F7F777aCRW+igV5LJX1
sefeblfgK9W4bUCi8Azll6a0dKO7MJqFdoIg1zUx65pjWy42uH6TPL6UCWTzkNLLNxiwQ9MayTGv
7l/UCFpoChb3N9h1S+vKiMHRAjcQhQpx2TrZ4D0rOKiP3zcTcMIaLnyC37smgO6foRcHpEeA2ttQ
HVZasr0qpzvHqBn82KbAJvon1BJWk5MFxXQkxgehIU7FUGtTzSkvj1wuLj0V8Y1ewoUM0i/9kSFx
Y09Ak+zH+tLuKZ8b2k6BQ9vbg57lFErc7fJxc7AR9r5CT2C4afSVBa7ME7X7QonabMiRoXl1fEXy
3ZBpyChl96mJtvpAi4bIZ7csxoC6XPb8cg4m5Tlnk4AQlYA7DUxbl9QQ0jX8qojxA6flMmD7cLii
3syDp/bKnN7ETUmIhFt/tBZyjMO0z4ZsWjceM9YPow8qeu2fUzNwAXODO/m+NZ21/8gydLg4qWPF
vArmFWnM0KWLfLZR0k6p+XNG8jdzKeyKeVD1TBZR6KVr/h9AJc8oWScfhjVxhlIWcWRvth+bnnrG
77Zitzn7Wkvmc+x1eBmSmRJT7fsZ1wxUTTPcCFY2rY35UjMpHNFa90VsyZizZVSQsemrAd2eCu80
M4cvRp+fKAHW/PvjX3UZBRAwZ9EOfYdFi8A8AVR46yqTMgeD1xJe/YyziTh8+ehA39UbqWDeAk8K
YfK8z+ILoPlehrwCIsh5/uz71nDGQtMI8g6dkFMmNNhrekBpKq2Uv8oUbMzs/Wjwh6zF6VAxg703
hk3WHV8inIA/ThakXGPQqUnjWlrLdsBhsQGW5d0doQVFVd4R0XYrq0sLXOeBgFUqGGovfNRS6pJu
W+OLmtq1CzEwYg0dssFyrttOhFikdLzz60SWX1i1dLQtfw2IWuXnV9aiSD0YRaT/ukqmFuQZgT5N
SOovhnNgqdGit9lnhZmHUa2fClKSY9aixbG+/DfoZgHTLyf/zOlRHOBTlVQ4o4HvCUrK/BF0l3l7
qCUEWh6CpNdZkN3w5Uk0yMwZO1I031tR+E2IOJWHMLekPtr6xw60/E0WERBh+gcG4h/13vNoCY8r
hh/yBndN7JPsiKuQPbaQB2BZQ83ATmS38Z4HwFEf5A+64bZO7xvzjYXf8VMgDHqCkwkZOPrkQq3Q
s0TtINt96GrCMhGXkxsrf/ucsjfPe6oPg0FatmD2qma302xK4fm+O+CPn7RvtiM7kxJrUA4MMhxL
HQe/7CHIR+RGpoFVPSwHvCaGMU10szWZbIkTtKp8x4kMdbu+8RiUKrno2UbgEp0j9I9kfaPrTylp
OYEYU39ZELDV6MRdWKRiqsXQLkFu6pFak4vAe2p+DUrUpqCtyBu4d1pq4dHKPyzWCGKHyRIzKTtr
+lvHKJCvm/zmGEqp+/wdp4CbNs57lyEMSJ0pinIt/b4FtdUUQrnlum8T7gXtItUsQu11E7Z5OLeh
cppjxowEjiB48z+nrDvtSm3r5DGOvuaiYZacIcND5by7klq1t4GGu2ifZNRX6H9OLGJB3B08dK3y
yPfKupBsDXisS3Zl5DiWkBZZFCRZdGbTnc97gq6YfqGtZVr/OyZF4A/KiDO9EOqMrfUM2jNRNogs
galWHrvEI3VqvLJ/Ex3KmldqplBJVjluEc6x3x6BGfYm1JKsueXLHRHEuvZqpSZJN/5Z46Fe31M7
PWufyv6rNG2eFmGJnkdJBjVzJhMcEEuJisiK16k7jOoZJsnOLJPA9ZNvjoiW7SDmeWPY9iNEIaWp
kWp7jJLoQeLe8X+zjzp61lT51FUxboeQUbhuDKvQghMEswNvgGhH2KJQvWb1rHgBUWF5TnJci4p9
payz2bndb939XHtGq0Dtbeee0PVeLYn5eOv/KxtNnhYgO0ZM/ct2bit60FXaRCrK2jkvmjesrFkd
aGARzerTrg8DZq6odCqo98Q9vuNAECBf54dxCX/Ci3b25UfN2Njp8os3y328L7GHXBZDZbUvhxD6
0qYTPUoYzcT0oDJJ601lgcU23flxTThFOU5dS2amo6zz1wRHGflo7/3YCCYGleaycCGs/85UaMhc
NUjWateZOmE9cJoYtVZJo3EK32BnBwa05N2CT7U72mRvJSojzz+Z09AYgdmvT/SXLy2/74ABClIC
xi23M+JsA94jKFsMP40pGZndqsO61Wm39YK+BCInedfQW7o8tZtJxisokZKr0cvCk681Md2meAdW
QF+VSOx2GdWBMdPXnwKLgFxpochoadGM9p+YfBUObUUT/EbFbRfXYuPX90HST+/piPYxfPpSo4zF
MtHVrWX1kr3d1/GLiQMzWHDntKuTarK5bSyQdDNVTCXvv5J1MVZIsQa0SNl3H2xqfI5LFQWvysvI
rNFXrRwKjhrre+ewDoUeANHcp3Pok/Ymu8/CtoqSx7e8sqb7cSKZZ0HIvgFtFccxShauTBYNmBVq
4XKaHfyMGNg0hDHn0GJ2b6oY2CR3KCPNDTgFw9lbpZqjdS8dVKCBz6m7QAZ/g8cdeIo1KAg3LSmL
/DgArEIURnyi5f08XI9axOVATIZVwbQA/1v9iv/cuRVpVQ0BIG5CovT+2wj1jOCBP7V7LnTD1iHz
NgGsDCZBLoGGeKbuohAx/mCKp286wopquda/Ui0Jx2h86v+61FQ4zFeya5tyX+SogUaaZUTMZurT
5F9huSr26Fox6o/fd/y3MY9WwwQIPEtUoc3dnFc2mGzk1DjkpoZq8uxqoVzJhpZBzFdVN8GFD2PR
oSV9saDSOe3tzMb0r2O2djJsA4mfHTIwnPz/e3W8r7S2wa0h1QC5Jpyfsi6Vet1hUHSSrHwiLdQh
K+FSUDv4RatJXPxzzdTAUNSBWQi65KMyJpol34MDbSwsYVNMTvNFOGhhAxUPPrRLht7gYBt1LUsj
4/ks70y/uzsrHfKpdHiyeMnqfbFYOXrnXCc3G/MlgvU0aTbi+47ahPgJYV7H4cPGhyAsAXv15LUE
RIBmzkG7vvwMWak0ev2cXUaCFa8apMrbFegZqEhg3cDgQRsMMI9sFddZguEZrMEWEBluG/2iv5M3
9axO/YOnHh1dfFw2pu49GOCgqweYqiKTBbUXWnAvtJI4sr9cp6cFYAeLsOg5uz1TQBW7ViyuYlKG
xO2coM34pwlP4cm9xy5Ib4zQcfq3yThdhWLPbA6tUQNuIUT+v4M9YxzfXWDwvPyUvAgq+OLZYkpr
oJC0gukwTHDF94cj6oNApj7ZnFNgDl6dLFw9ZaEUT8zEEjL+3NNO7IvQNtLIUbysXkcHHfIArF2j
2xdf0e5Oe05LSpUik+U+bLGqo2pd6RiMqPSZorOC8l4ymPmcsMk/U95l4WxFXcX4wOWsIG1Jaf62
kKNEF1NgeRdPK95sBQjOsDuGVSqUGO9Y+X+euvxyYLJ0b/x19Eo1NS+9VMBH0w63IKBdscMWKawO
yOTviqVuG831u0nmRb/bUDZVaYEq6EAMGR1KpnCfBjbqzOcyH82dO2iU8qPheyTZpcd7Sj3DMRsw
d/dErm/1gh8+MylyMv394vn5NKdJ9XKb3X6D5I/PDQpLg47cHZryAryId1U2+jCd8Dbrgp1sikqA
f0UU4/SJYSlcKMYm3wdDHG/cch4HqN1IvUZJFi9t2GTtcW8+W59nOL1LiQkqCUS7JPnHePoKLkPp
J3Y0OztG/a4Ci1cqoBh5ql+eW7npYV9v12OkgTiKnhHf0iVe1AKJ71tLe1Gc512k97OGxKHy+KKb
rU0bNS5bYG4/Wo4+otB98vD5QbVWGKixK8G3advnWI13/Ojse7rE95HKpBBzY0mIBIxjmfJokUvy
RbnKanEI6z89d3lWvDs7N8IWqBMLgWJcdjeweVCoOxnz5Yajk68dsWIWNoGHt+3ewFVm8Z1F64Yk
PGxupUqsu5J7rnbvw0R0CZiJ8uAWOoK93QbnRWK2btDOVXr7G5/ay0NChKmdc85031TiIX28kQ4d
utC1P96zweyDN9466JUsjCzIadTLJrlkurZeSFCN9/vr2Yuv/FeettwBG6yCri9zcBS+Ai483JHn
+dyHDH7tGsRKFfHK26vMLwkFcbx5C0McxQnzNj6E0bbuOTKLg3QI0EQKVVgevcrO4dgMIGEIbqnh
GvfAA4U3hBJYqInxoppmcRnkgRn1C9SJ7EQqUAb8gkvlD2F2TzhF3AiFUnOPi4rw/YU9im7/ldTI
QPAKRxTu9nL2VfRKbgXpFvmazkyrtG1q5OBHUGbQKUfVKGfBzbp/Gf1sY12gGf2j8iK6imDnTkl2
9iQDaAeBK2iYsJEzm1HXzPZv0DmKpBUrdk5x5JBe5TBu4I/MR6im23GzJKxwGvYICf+j2EJmFovH
1863yGtjXstJq5hw0jsGopUMYnU8z7CtXtL6K7wa5414SYfjauH+YrVHHQTW9uybgzNEY0vjGOQe
cULkGuXrWGtKIPIMAI/Txk7cS6OHZ2/vC5d0xFrKpUbI+MzA3G1MvVc6Qaz13y7VutD+YD9gJwNP
iCBk0f/a5148uTqrUu7yFe9ZAvAU1viMlstXAxZHOl3L7kxyHskZ92k0eGwJYcQdRPozxjTnaZHT
FWnsw2RlKEUIhdZObyzjj9i8SvjMXndNDxiCr97dcEfDg17mWRdBcWZyfRI+YbX5F8qsPnnygPK6
1kr2vkWN8wBI8Su4OC46+oNTsFmDPsdbjQDZrLWRp80GIksn3UadTuyvwRPXm1otojWXFUXFFEr4
cDhroWWK3lsRA+nikZIlUNgWTY1HHvhPjg0lM1Ium55rnMC/fsv4Zz11aljnXeoeXvwN/Cfay1RI
DI6f1j3f6ZHVvoCF5/TlQnzATTnrLoSh7h6Y3YAFblAAK+2kkS1ygwR5xkbjU39hoNM49xSY6X7m
JQ/w9ZxEQ/W2VOOSw23HK2/z8amekxZLc9dHlpFSyPtuDGUJ7DA4zq1SP/MbCEwUKNFgxyjDZ2Nx
fETlLiw4xYPPv0nYp1/cUthnXQDAJm+9xKyQGxxx/u56U6azqi+vM/dI361RAIaj2VofQxAKol0g
5Kb7yQl3QOs3t/gVWuIWzPS8Q4JZjC/WqFkRKKU7V55NA+Vh89yiLqo8EMUF3A0JJph7dnf5CYp/
DKU+QL1HFkOfZhGoJdWQH0DGfYm2skevgzFEoVXzlEA9wBAQTTXhtb6822qfoKOeqxrXRmZ7mBac
qqgo9TTav+B4dTqcgWLqYt//xIbqjcJOoTHFc2GpCxA/Dph8j2lWgx624TJ42HGQnBkSOBP6LRyK
TVEL0zN2bHgB/elVovtI6sAye+QkYCzB44mkZn9+4atmJMUtRsmyHu3/x8uHQW/qU0NqtISaw27n
mPoAgHUMBPyCZZXe8Eg3fnY0s2Xp9Yums52E5CNNPwbB8s2u0BfamkdLPSUGASDSJbFHOFJJLrR9
v9NvE7ECGxdpTN2KP9hIQc9dd+I7jz6Gb2NVa9DvjMdHnK+wb8fdOgjPlIf+V78mVsAzYHov1bjd
767wcITOcXtAqmlQ4WNf3xWZr0PCdgcl/x//HSeq8OuU8iOt/8eu+M3unLVdo7rosrrN+pRBPF08
8HkQ8w8+ETM7lD9sWMowIThhBH8AdgIvtgdntJLaMD5R2j69DHfZIATCtvS4QAuJUDgij1m0NAuV
pjRrhUCO0fhRP/n54TEZQI/cU4XjXDdzOp4c5noTv8ZyArR5YWQQ1j9CmKbkjiWuKh3z/YFq+7h+
wdffO+rDx0LfeTjxTjLUKvdq6kqZwcNGvNamDfCP0QiuFc7BHQ1d4jTU+N+9KM6cKlM+bhOv0VbG
JNcsTdjdK0qk6vWFgZOvxW8e+IDyiTRj3xzWahj4X0JRNX4/g8VoUFvZEhTH374JHPTZKeCRdhRj
YaFKvL9rx3pRYUQ+itD9vVCjAuc7rrTBm1oUwkDpfj+ZvMWRBYfVirGtSUprdR/ubPFPHf3tAHbO
UJ+cE0zmI+gL9KmCX5zeTcECMI/wDqP+H55WluCR1GoSiWe4qOi2UClQtVFC6exh0WIMob5IDxna
ojl+OBHJeoaQtSZY3/b8GARZ1xpktdZlO3m2a7nIjdQD0FNhaCmRmnA+UsifwZ9P+fuyxFdRdNXM
KQ5kIWiz1QZzk5tpWiP+BZDVcW0Xb7GKJiWKP5AZmMdx8pYPDVsVFQMdsO4jyj8X1hae4kCgwKw7
TFA7ZlgBh45sz2Ebi5zZ9oWoXt1ImA3MFA1RhQQbjmUIRpxRvCNESfchsmRlWO2BDhBfvF/k85V3
Y5Viit2TiLa5/dQlWqycRumu8tlrulmflSod2+ERaJhl/XqBtvW5zI40sOSTgJEjMVOK+yxZgWNo
3lW7TIyV8hx3RzpdhMPLhuMPLc2noyHm5NJ43TFuEWivvoaIrXewGARqrYlv+PC6wdW9HgEi2h4Z
M72d2bhiqCyodL+4Ti+kxZ83a6kdjFJw/jGBVs67VBXj7qgLazDvoa5pHC0ty2OwmnkcT0QqnhRS
4rdDCLpnJr4BkaeLSkmBCs0KxDzFQrZ4fVOJMZlEg2Hyepq94aIEDfV6PDjhP4FM0HTqa/7o7CjN
DZo/DvnkQA3umdRbIFUxxMuDV314XWNkS32NpocyJjX9QbuJVJTgsFgLh18qWYOVCQ+vUcbLo3EH
mdWCajG8aITJDq8qm3+b+fAfXm5kZ6icHigTiQDS1liR4DHRSHft93RN8Hssf/cL2uUabRZe98H4
41qjymUbZ4IBcbV1QBbt5Eq9neMDbFMSKH3d1TDHrmrDZzE5wK1X1amLltqhCFsH6wfg2Kon+cuA
1iNmsjITfqyyePhvS3xiZTF+uPTDWWClFvP4+fhCsrcgAy/pASLsGeAGXUB4ZfwTVHH73B6fvtmA
FQa9XHn/vtAFYS7zZslMsrB9KV4hHkp6mQdP7Rv5GC8j7r3A2+sbLEpUv7EGQK3X4ftqLCCf9+ip
hDH2KCEas6Cf0uN6FBfdBD2Nlzwsjbh53K/q2j3PTY7nzWbMrXPtW+umrM/fAU5zisEbptJ4t5VM
J70EzI+KCEefayyOmpnyBQBQc4XflRHA+pHDOxk1I9SQvZhR7epI9i/hUZ0jE4PB/P6GQH5FFyfb
X4ptQX5mzhn9isTLURd9OLmDynTZ+wnRYaiISZTzRnEH8dQLiZvZ8bspDmAJVuSnyJn35hd+DM1d
wvOVm5rQgHJUglDy8pXHUWx9CkLrJw4uQux1EstxcYi3AXG4Hw2kt68UukXEmjV3Lu5ynCBEPyKg
VZVig669UIc61oSLtBF6heL7u/WI0gRNi9QlXWm5WkMmwkILngTeJ9NnEfoedh3/IXEjSwPpYMei
QuUrey5lqSWc4ZSdgl1HQjowXhfYc/2skyBXwv2T9kfuXt5rwopGyy3x+9OmUTON/pA8wtd5/Jfu
PjPemFW9wdgiHrzu7VVq+YDutZgePAzOOGsONOypfZvcVoKR0QUZLI7C1+dtjOZo73LhVAhNHtG2
HldY05PjBW0JQh8Tx1cZHrQfsGWQN6vrJda0825JhfIat78+TSA+RSyyCydpuJ5yen0TY33ud8e/
Gv3WBQ51qGobRy4hrSF8J/L41cODl0jd0eTAqFnKIVoVMWrDnAnpFGMoVDrijJvR0sUOcwOORwY4
bWvzNrHn+Z58K00smylq0dVDi+FZM8OpJ5Gl2Vnw5/M9NWEFXucjIfnBYvb2z95Xyi3IFvYg1uzE
CrcyHKDO6woHQ5G+SwEv2weto0sqRTP8hgOcNCiFlDHnphBvoKvdlQ599VgX3B4hG7xnnI+RAq3F
/rYueWFo9+uhN5gycJaH5O31FqR5fvuNmI2INxH84slCe8AzNpSzQF8AdaGlFpz+CPz/WanZViP9
K6VXJV/vtHG4wWYYzWYpVO5eonJSdqfkG+3uYqLgfinHrVonhHVCdWfxqbjfevF417+yHYX/mQol
enbm0NaGZQDLZoBvqQVttFiEjK+q/DDgHfHZyWXe2NfDUqWmkkLDDlTU6YWVHB1ntIm61mcSMCN6
rC91IIp1kSWw+UCy7tFcTLpoieLNNf+XAOrfYRJEPDXa8bux9CldxKTnSookUQ9Q8vdaKEUVeBlg
NtsxInPfOwCcGG5GtA3j26orTjsLF3HD76o5uEB4OH93GRNoirz+yhTH2NKLT/ialxseWXagb2kw
cHgI+W2eANhTUsykpPMcDF/sys10Po8gFEB86k0o0fMokDMO89m1cpCmjFuEpMoIkDFtyvabHbK3
GB+3KgxCLC6qHe8+pk9KMKb6WlNuLEcZRQqJordDxeseF0cwdjTD11RVh94IT9sNn0PNDx3wPbyS
e3AtXYiDgPQx5JUPktRharXXKFM09UgV9W16GHPg960pk7Tl969zjS+8Z8QlEFGiWNWcapYFBTXq
Qno/A9Rm/j+xLlTyaxWl9nW0R3V+tCEE7gpn+OcxKyCnnibwf7STaU42vynAIu9YSD3m0kzdxIJe
7m6K6XZB0y7mZ2X6n73yMfrfQTX/QI7RavsiByXkCe2XeDlUQ1ER8X43+mKoOnlgZyHynGklK5oC
NnECd2jJKIQYbQuZZ79qtNSwCu2HBTzh+cDJ/IwkX6eOHKcPIOClSQWVODEI07bmd0nyD7RaZhHW
kIHdteKyTOg87KpATigyCohb22jex+5jhStgk0m0MdJVUlYrTDBzuZiP8CrHyl1SM4O85XjKYAr+
lmWKtZjbCrH2D5KCtr1cF1A1B2h+C7EzhzmJF+7uYid5OPpzieCJfF/UCsvfDQCXHc409NJLXfyN
f+4E+cbX3C6tR098eYor2fdOFoTU95lHowOvA/6tU9pqm5HNT6HwL910n28Y3zWYmDhLSZ/q9XhU
pnCLWpVYIimIg+hfwQ+fLIqCPsBQK4xtJX7WkA1VCrZTHnikUs27mSYvuu6s0gcOHstUOMEdyDQ3
QP35Dk+JPUTLNRmHy1FoAjgIdZ2Qa3dZqiUt53O5Gadmy0QJYtzwdq9B+e8xC6zfuWQrnZJrexQ/
pzjwvVaT74r3YP5GLWvXTHcl1wbLC0AnOmuKAY3+Pz076c+mp/7M2agmrQitl8EvvqejeUE+UgbY
bnGibRhtNxm9ZwhZ7pYkDtdp/DKgEA4QBcj0AMifKw+UX6BogdNeA6otllufUhkVmIjs+UbH1n8P
+yEGlpEZW8y5akp3s4NbcLaNXB/ju7c93FhsAHObuqM9+gGjW0dkg0110zKpI+SjL46SCmruim+p
LxUqH7kVl801oFXXIF2Ijum7llO++TQof454W2XkbnZxaDT8Wfeb3BS6moCc43f5azwM3Noj0bXy
Znhbbfi8ob7Y4B9u8guETua8rrNUefmn8g/lwcxl6n98onq6bsWdS7anQbRs7d8X0hViZLDZFRW7
xioyoh8yBt/aTbeHEeonGi/U01b1FixdVTydI1jvPcbRRADz2y8ASFKC2wImxY78ewGHdOf7+nfh
HHl1Gw0ZGgc0CJ//JEkvRapyeK13AqLKuDmxpnG2WEZL3uZaB7DYz5wnFreoW/oVUa0TjvjHwxIs
dqqoFdfpqs/WI/Zd8I+QMjIty5XPf7oGJ7aMGkrynBAkrWF+Joe5rqZAUd7sY+bWF574uKhh7VgF
rpWVsS1w6b5L1nS6dpXpdjQKSihic455wO/7BbAvMFAYzOD9KENny4ty9lovQjI4sh+Sjn/054kK
HEA3a3bZEpiXMkBN5YzmalKvLO8hO+MsdglaFxGX+0Ra1r8TUPOxKLo/j6IjJ6nlU5ckkkKcBB+V
fOfumnxqiDq+GRT7qMpLtVmmyTVBDBxS9ER9Dq9KDSpWgep/Qx6GmZjDPwQNPbhngK6g9NmyRZTy
IOtxVljjxHNEU39F8yFmBYOEUWD8bTax8vvsNmt2je8tD1g2yNoep1lKH7jDffAZ9L22gGNAwuKM
7G/fZg6N+3D5gUp/exzy96ev/P98xZx1ZTb8iz5vrX5iQt+DXAQAyuqoA9Ns8dVodTufs9NA9UIY
JnqgIO1D18b2ZChW04TDNDSelIpN99SPsvC+O9zN6xPd3LoEMic6ldIQl+uX548zR21R8yN3dQfe
jhz7EdIvfD9KDhJE5at/3fVaxxxT9XmktPwodDLnMiOrBqVojdfNQYIztYRdU6iipAs4K3LgdRZ8
jltyApjQ9h1UDF6JxoQrM0Uk16pIEsrE84cPAMVXeB2VA6Evt+bG9BPHwUrNEmJYPTbP/EDBLnzp
fvprpt20l/DUB21wZ6TIuqxs3kNVjREZzgl3lZ02qlcnfD4iy+9GrKpoCRL84kuMUx06qODvYaIV
9WaUZ9blFKRI8ftiD3BE9UmJUpQUomCHt5bPHwhATbzPjqOHIi8L7bU/+jvYeqluP4uLqU3MAUkO
nRxnM6mPzZoWvKjRwN0JjKqMY5RUYS46yjnO4/QPfTsFqUH25QfHTZ6lbdPYhGPW2Q6NYlo5bjZL
IHTAvS173bcGMrmhBSHCi98TO6PYWcqucZt7XLajv/GExeF5xLJ25UldurgwfTzjsycYt1l2hP45
IpGtSIG+EteeeCP++TdsYMgykWJjDfCscussQxG9g5vqbVMOylWRjf/3xjhcCavlJiqa//lkjZS1
FjLTOKfyhkQwb6C4x/ohTS3AVhW35mnfivTLMfJQhgkQXSQojeO7atYRLya82t0Ch5Igg2uFiWDl
4d46dvitRsDDr0lgIcrKC2U0nIkQb8uokdIxxMWJ3WbTrtXjPFxEqzOoEQ/sH/o5ksWQ4dePs0HT
oq2kSp/TYY2tb+pT+o8XUglxxR8uWDtmBQ78c82adga4bJPaMxpOQBVscE8ewogShivsd90NLY5f
vqAYo5k3WuNUCOqHMiWIlBRt5N2hPS9CtsCGC+tgh0pqb6v+p7AX9m/4F795P9Ed3naZMOB9cRNa
Yf4GCCwcaFTDgdO+di0mHAaFLuEvvS8jqdiKKJ1ita5vFfZhxrU1XriUFPg7BcsHmyjtAeHnnxkI
fWKYnPQtzZHWFyfb7dm9v4aARW6mcP05j9axJJPEUWdLdkU62SlR+hlAYxSY/NsfQGSQI7lDztce
xLwFXXJFZVPzmhCLP1fAhvItic9oKJCpKAjIrJdvkmIZpCQJXnXFVQJWV+sYoNajat0zegDpuTte
aTDNtTkYRhWmAxeGEtYJa+AfKSEryI1jNfzoShE3+dt6MUpi9fjj86JC9c4UtPBElje+7KETTPnZ
o6FAWbtPUbQAdmqlXXhqmBk8pjSTDpfjvVREbmjCKrFlKVu3VD2oAfS8XG6g7KsZcxYY4jFRIIys
KxoDedhD6rwh/FcpOL+XKak5eTSCk4CBKMITZKxHm9eyhDdi7Cxai860ljTiqTGhksHwN+oWPaNX
xwC40WycuFI0DoRfGFVyT6a47ArtYd474kO3Kr2OYuXpcnMbaEdkiKnIJ/DvHFaJuSpzRFdzzs1F
43UJrKHMaGw6gY+k95xmHoCtvwdUUoSxA+xG9wlSxPS3EJGMtBh24DtubUit/dzv+P9VBnAL0q+J
sJyZXVARE+JfK1i1fjmF6k2Np9lBmFMTD6EDdR0hsANlmskY+g/uSrJUmmpQWpwVlZ9xPJrNnOx6
Ec7DLT8M6ibO+rqry7MFe/2z9Nf4Ha59E21+ndKwa1OStb0XtFBqRs55wdGGmMO0IrbmJvwl6Gri
zXLTaAig+UKizq2bdaWYXm2RMacdKpN5NZdhU8jedB05Z48wZA6HAQVCex6a/XPkGMgV+QuU++ww
eJnhLJmHz/kztKUUlLQnDvaGJFgw9bo3haIwpT9LtFBh9ffGhpIA8qG5z+5sdWDyFUHffwA+UcmP
xN4bQXsjtM52jtekjJIIvbJfgI1jPcBLUkHuJQow/WlLpDMgFZ0uvNi5uSCT3DTnvrCZazkhf125
Trw/wQAUtkrfbAQ28I1ntkMY3FkcqEr05vXNqK4QnvqfA4eS3TwY6YU+xezDxdzFoC1kb4B6WptA
BvJwBFnHDFeT4QZSHt+IuBB8GJC541iT3h3bnFfIp1yzbhTpBHMpP/JGCXVG1e94yz6bJgny+j8W
YWlEGm1V+mYHrfdNGuH7wno8DOOw5Q44E0AJJ2RVw9SVkwftVnl+aeWa7Tm6AmedtyoAyR1mphnl
HNPnf1SwpoZet9GTpQkZlYE5fePi6s1JUkRnbNj8ED4qScNO2wJdKl3gA/Lib0KCAaOSIBzJgBHZ
0xz4Nr/19aH6ylofjkapzxkSQzv7nDtKn+IQ9ZQTgE2qOPgtZq84ElBF+kBj2Re1LKjrmJYh9lnu
3EHqou7g5+2sWJc5tP7qc1gc4hrc32X1p3pC18a9fNZ3UfWbqvX//CDnMf9uIB142pTNFXtyaaT6
hk71GN68We2cuiLk9q/d/mL8gKfzm1K3bbCpYuf2mZRO+c9Y6MszF3QbfAJMGoeqFh5GF5BnMr1W
xMBnW66GLImSN20aqI3X1semJ140DuKnzntm7Vj8Mb0S5AdivFdyAlbq/UR8Q6cZOiP0QzyXIn95
W4xAgMgMdcq1cPKLfYqa7rDUDTyz9uI1WZd4KEnD3YOOWTN9qUGbrrdlkjATAherbrqd/JlptFYH
me44rp1Mzf/VGOKFirW4rzEDuNHOrLxfYtQ5FevOr6SJfkO9LnbyYM/tS2/7bdhFfcUbr/PeuWh7
UwZwIDSgCtwQcdq1VICv+9kVzi+Xqs8gWyN6GiEs7M4FxUdszgs99h7lK5SR9q6v3cD48yMDjU5H
Sp0Uocei+Mzd28F7QSjIy2lLAVewNzstDExsEA6IGQxdhaeVuguSeCmFZvPuIxCCIh5OExP8It3H
vm0cqbMayI0sQ9mJ2Xo73IxGAqaXK7k+NgCAxkfkRKONASzzFZHKZELCXwY/w8g3E/hGrtHpBOmS
7JPD1cIHwjGL1FdBs4jzG1mB0+kq7Im8AO/06p2jBt41iSejj3fKVW3JCmuvTBdJEdOX4q8vne/M
tYqKl96dWb4NcwlwDKf4w1NgzZ45NRHfLdqTYwtI7uKqmMQNdOJLBVHWTOZThwzLRFcoBGFBQv1y
Gla8iLVBrLWS5X9I/JAGpnMaM7QPKMZsXU70ZadWH7xy42xF8ZA+2Oz03D6e3RlbkQKd2jUvfN4o
Cie4FEfRu0YBL49byXGILML0ccRJWmfilAZS0b99XedWUOIR14UynUTkLTU8y9K+3hE3jK3wbjqS
wd0IZDMjiaLvLES2hl1UjtMK6vZqNXxW4T16R8d6AYeMRPQzcDu0ss3DVoh6XP+VjDFlwmmGwL0K
3MoPRNpPlYMMk7Yr8zhF9vtiLTQg3b8uUxb2v9JxcKtx6RcrCdrgvPP6Z0MluxcAjcf/SQgtxYfb
led7XXX4J3Sk+lEjIFXxK9XGDQWeAKQ0h/Lty0ILCel8bfgJ6BRzNc2NTqTc70fPoshcSZO2s8gv
x606VRVTPjnN0uc9157KslHuhFGi3AcGr3+b1YGJAKQgPQas7iaJzqPagd62tqq3jiaUNzDL0ppa
UnQgWOC3xezBykRxqMfjbRhvP8i34+81orANRHdL1XJkA3qnt80yDdrcHLMc1l2o9pMF8agpFRkU
mErd4qp5FUzyiFgpafNbFLj4b9MaGys+Wj9Bfak1P1ynAfD3EN8graHhXWZC/e4Zhers5nqO5lE/
eKLo21j5iY/jFPNoUDGKUGWdHf9ZvK5KBTrPEPn9Nh4+8P1SK7CptIB/7GY5UtJMLf3OnV6WDgMS
Ck93MmjtQUoN7aWhXFq+fMctzjQMLFpHswe1A9jBXu8ETWLDpvYYH5awr60HpSfXGpkhgyoCzmtg
OYcc/vum0jH4sO3ckqg335TAIrRiZ443qCqn6c6sbuq4MNZZvq0gM9BjSQbfhqw7Zpw1Jg3cMCeZ
TdEH1HFiphKtcbbiwqOY3LmUiOANhCfO6JDykM26+Ixj9tNwD6snG80YtamLaO8IOwcW2wPA7V+o
d+efQcZZ/qncC4Z+JRaunSSHqLWXl3UM/03LJnQvyGlGANhvbbFBghONP7Tw1geVGfanLDGKXYem
bPVaFnMILylM+Y1sfSVCc+6gM+v340ff/TZFZuwmqIvNxghKj2pXS0E9tRCaPaJDFkBuGk1HA6oZ
WrVzugn53qM5VwCMTmD2k2ovf2qf2leT7htv93dVQ7SuW578QqqN/DMmvQAnAB/lxmO/B9WNIfGY
M9Rd/MPOf/JEvBoFXM18Lz8K8yUuP3rYCFodddrnw9u7MZvwBlrsyhgVTzADhZpUuVGwOMt+76Ct
Dhi/ArjMeDtYD0SyM/1KxnWtGOf4sOKRnOu/2gGhUQZNibcU1hAYZgWxCipTJT1+Lm6hEXeu/uOG
TyZdLTM7Ey400KGxVi+WkK0otedGwMoRkCcZbykCCwOgHFEpT118W+6SJ+yNrb3sAZVL7LSHaaqy
kEbXRo91k86iggdZsUZvy4zoLqHDWLxRkB4bOcuU9mzTH1ghf27RSNFoOrtcWQv0JsWS3KV7k1pM
+7Zq+fjQIE15AjiES94Z2h8uZfNZy1z5+gKuEA/BhzxyJ3mgJLHLnfq2fh3TInQavTviPHVf4imh
WzqwsEEvBVHfDSESFIblzmbK6Dr6ZlHMNAfqHr0i6n3ymZfrnpIxbFnXwFcu+Z30BscHW3BRgU9i
Vf9Bg/3pg7vfsXQGoEnX9UG/D7FSHtw3Pe6wL3eWAq1Ym1SCLrVAuUcEwl/sjFvVI82UcB7aEgQR
9fcyX+Yi2+OA6K2+oMtNTvYf5mr6cMiD84NMNILXOo9kiulabZ8C6/FKGZDYCQu+gN5PTutUltos
HINMb6NnKwTDg9PYdMqs5ZPS1g0aDd/HoMOTw7jIZjJLI2cn/R93x4A6sXC/H1dFAQTKvAqhP1e5
UJ6dZzh4DJmtM0eiOwp7Cruhfg0PeNAqJL2MbdaEe2DKW5d98bqCjJTkh1n0LIlNhPWvEVqsunba
yoCD4muUGVXOz6n6yQhN1YvIpT7bXOeqbtXpDECSJMUs/dCDd+2FsqQbJEaRXxg3oxNqWIRILymv
5DlxOLI4cZKoY5RowijWMI35OkJAhi1XK6lpxsMgM6O6JhLD+42hSTmZoxbiQAyBSBTJ1RAMcw6S
WOGdgQXGSjXilieAreIp91yz9bmUey95T/QvSLRWGKSWry3WmLL5Y3M00Oh+DT9ZybHZxaeQPj4r
C3ifDKeFcRoCuiDm/tnDgSHaUL/EAJt54ukPgRIyDW5dMCqJkjwjBFQ1M4egssZ8xmorOwnJxOzv
QQx6fUpKpeD8QiWlDkW8Sx2PIEbHI7s4m8Vk9UmkIB7pIJAvnmvh3HvL2Vd5yFg6iTUdrUOYr0lU
9Le9PQhaPAz6ud0f6lSYgv4IfZCkySNoMbnVDcnqEN6svEtR57NzPLOGvnC5Uzv2GSM8Zd6ymAt7
YLUpjVpu3VY7dn45yGXLcPyk3o0iQgBNpdBUnqeyqLfBlnS9s9Fk/zkwYdnXYwdT5/9ORzG7uoPI
sGd7ribDtzZcciKqiMMwqzml4akO209BHx16VrbQRu1cBDXK0/5upG80e3pEBpIGGRd5KVaDibtW
Z2LOPq87Dme/Fnoha1WonPYt/dE0LORmJ3qbpg1BUrldI3dQo804uTcDi8+Cbd7WaRE/b2CWd3lA
Bm5GOg+XzaCAw5TMvk0rqxbZkSBsMbadIPD/7jKJCvrQQJl83mZRvVCEqoX6IoqQKnTkgY3UnPlT
cSFVSvKn1DgssOV4K0ECTCAI0BaEV34gedN5KZVu7BWz6UNAL9RhMxz5mIOPFE9fDGd8dfUExmDw
7tB8bvmE8oXhTAH3hQyOxAxG2ZJ5rB3gyxIlLthoguhBQ4M48h/Pm9avs3LD9yE8ETMbFKbTtNi/
K2epAapXcUVkCsZBJm29qx9dKX6cXHABFINRMhJandau/ogosqBjgjOzMshF1nxB2NBObNsYMfpC
znuNj4thtVit8J4SfKmE+/0p4y5AenNBSjt3qqpJlwkuNZR9XsHK3WC8dWnZXEAxBNE1seoK0Fgn
JPkYrTQH+466E/at4uiXnKM1UBVgcATXS564iQ5wrKFe9MAlobGaBrg1NqYAcD7ONw3LB5p3vehR
/6ezcWbSVc5eRDoAo+P/0aMGMNEO5vd6G39i/ReGXTbQqBwFIuXZDSTyN2B404SEbqFsualjV4sg
Fm85D/wwaV3ZeqvgD8I7+rE3u93ff1CoOlu8moro4j/zW6zXy0Po+eVU7Se3ajF7v9oYXfrNs8w/
tiHGWWb22s6qlyBtjomX0dF5ON43bPRX4+SBGwRXjS0QMzkDnZ7h+frMhzpc+J4tA0ExWeTsXl4B
OA3o6L9VMoMEIs1zvEv7GqtRVRZJohfz0rt9u9QlKNdI3LLMZNB4HAwrHpRqaZx6mhQwr74KTbV8
iNYxwhs86YLnNi+bZWIeR4zNo4lO2GSKUuOnCCyUx23fecz3RGFtAIw8SSHlq5nrLe/lenqeYTKe
Aov6bpqaiCieK3IR5ygI1XA26Hdg2zTr4Q/3rqPkOec4Ie1DmYQQ8Arefjx2lvIX9/KkwsNenus0
RSOG/LjSvUaeFsRYwc77RUw5sl6eq/lNUJI+WsARSQ5b/jIA/QXNYDFbVRcmnnYeQQHcy9TyS7DU
Bi28376oPngG12OlaIpJSr2hRxfJAHaswq/DZkNiYaIjBTtblN1jqR+NT8h1TWchzgoSnqwpaiW/
R3d6k6jG6nya5Iib4N6yUNvwn+L/N0lzyVtWRWgEbc7WQZfKUoc1sW07+TqWiJwQMFPNNzdvxopy
3XVeYpmrsSKy4eKNSqE2l/T/DmbOSA8yKTCLeQGf9bmvOymQGBswtuQ8TLWuSZ1ej/Xu9EK6wvkf
FJNekykDMbdySCvFYSww3BpuE8DF9VUVuzOGylcXzTZ0ugMzEOpcL1ArhFeYzoxu6ZM/eo23NXrw
KCnjUwWFA4DfF/LhMdGdyEcG2xSTHTdfJuh2dq1BSIH40BofSrY5tQcOLm2sMH3R6hco0EThICmx
LuSvSlYwHR2yMbPb01SYBLM5eRpsJ7iGnBDNUWRQKbfFqyXqpF5wHlhEZtMwmARLTlbuFupIZeXb
InnM33nBYO2nEHHDYO+VfZLzf6QORdY+cKhghnhoKttfjBO+HcQ/j+ylEErDWWt/JtX9p1spEYaF
s0FD300L2nMjCGFxVO7NujqVqhFBej7njG+P//9xFYEHCVnGX0JoULNXTTqj4DKcxcSKtnbaoY2i
VT3TGdJqZmEBaAbh+JpAd4hUDXX0MyZVlpPTu4Of4QI3u/D3FDvln9XhbWWCEVCQ9l9VJ2aLCrNn
zT1foIXXuI2kJ0J7VKv6gfjc28FfQU0r2upBdrxqLdov5BG3CLyPS0S3Un6UlNNkHWDSQ5ogJTvg
EXV/gWTXgSbsmRZprS426HGXm5YfBlOtZ8AZK2WzYxIkEOw+1PVjXuPvNlPZuL9zFws8BJmp9arF
LF2yIcKxPyF+Fs6zQRIYZwKS0vNWgR5YN8kIQCK74e4/0p2q4pMQJ1ZYz/xtQ/ZJarkdDzrHhUpF
+yjBqAFkSFF1wP5BnBlXiXgnGMqFIrbz1NUDaDLGPaJy31e6sST3nhYwR1adBWJ0RtatFDuJqXyH
VkE0M0A1HnKl4gQr29+32/z3//S+hxYvREv9Wo595WLarEEWQ8O/sPTn3dN16BEkKajSeqH0qHjg
gliZJX/FJeGGDG2URrbriYhDVFEFmg5hXJt51feuduwpfy6fZ/cRN8+Wo95LSglUonYhO45g4ydE
b+1MATXWX46kQVVOR+Ut0eZDNDXSc7nKqJJcbW3Suf/urCFWeOw2S051eSCGnbO8Qxi7tl7gY/jx
/YwwfXUJE36m4KYRxlb8T74c7Ra6RMJFvE2CtyFvoIgoVDG1ycyCS8GOHBqFPDb5zOO677A7wxRv
0UfBpySdqV9tRpWne2YmohKx6J8wjRzgj7V9M++6HLX5rcefV9Dy1FH5d1gVen42/r4x70LRyC4l
xFjeiUOHUrPIr6iZarmKF1wytFsD6RUMrG8YNWwq3xb3s44+iT3g92fxnCmMWkzb15/spN2+JOXN
tyzQA/2cb+iQlcWKnctPjHin/YOuqH5aj3HPRnsOzyJMxQJFYnaEBP0ylm5Ti/zhG12prl6r7/s5
VAaObiVHq/nDaiRpy6S/Xmx/Z5H61pBC3GepipIa9vqLhZNTEkqyX+oQvQ71vgtBrHYbSALGHuul
NLcZQnfrQ2QePCnY2j3An7y9RCbduJ4zPYxpaz7de4NTmvWhqvItqvkF6EnA8EIWkHfV5wu/5lzt
S6R6QiSBkS5Aqu0HTP+9RJ+986PAS2y1Kn9taYU50H5kBjRhQ1C+ji68ZPDIhwtOCEaHTSWJrSxA
ax8eVf99v6rn6Fa1ICt6tSX74v/si31ZYMmZJKEYhF793TTh0HoEYFv98IznaFFUKxxwf3ngn6ZM
wWcFDoOfxOB3jM9f01diXqOEg5tdQcfqmY4zwZJyMDwMJYdsk6WijdOeeA0Tuh3Mkoqm47mBV4yV
w/rYGBEYQOdFjshV5NLmrT6kNHfiruae8mszve7IfQyUJt3/7r6wzkQ3BVEfXOke3f55twOr1BCv
V8YW5LRwR/DIRNDlYyoMUl5VQsv9cTJiFbXginmAAtHax0w6+h7Fveb1CvYGea8fv/S0Z3fqS9Qt
VmZfjSb25XkJDQORRbxzyRjPTgZ8mWg0RwHn6T5s0e0IO4JVaiQm3zY0xqt3iUZqu2XCHheh1noC
5qtEweGZqPyc7QxbQh9Gep7Lw6AbllsuYkMpH+FRqrcgjcQossfCn8nv9SizKv3WdIzRu+9sSnEk
SBKdwp+50mby/ot+gJxXvj9QsfpN4JOO9D2XufT0V2hKygVU21tK93rrqMlcwYqoeoPeuGvnSVjW
PEFrwvRO6njQM6s/x13eIpd4hvRoqUhDRACfpYo/iCq10Q43b0vWyiq3kG8ryfzsC8jBpZ3cdd1s
2O5Np6mwtQpNLAReZHaCErUm2WWljFXH2qvqZxU6koTtRBwCRnMGSAc+FGiFNWY8h3CNr0QQHwf2
rEwV3tG4SN5KjIN/v8UX23ApVJM3I2cLGPlXQfesuLSoznpRSt17OGropmZEGYc5GnwlZ1I+n/cY
+YldsL7PdmJfh/xRUie9lM/kdT9b5/NRafoJdBk6GVezt0BffbuSDqD3JUnInB/F+/G6k1s/5mlq
rWF5DuY70P+FyMDS7ewTAUanAUVIM6MQeWhJlkv9t3oYYNRvALO2BxErmGBGDjFkdeIHIE1k18A6
8MWc/7S7PDUjrWrODz9uDTLgqhzmcIsW+pOoL6m8/cF/WzL7heYtxz4z1CiaRojdnCtrVfy7/I47
95hATYUFiTvd97RKzFvDJ47Sous7ypTHg8h4bVkprwGCnbb9OS3gWWnROOYhuS7z3wTjjQzFwIap
G5KhAPa9YXdX7PTRMzjp5NXg1TBys2Smt/BZPmNcdonbiR21bPIhgTqhSKpNhjBMgCH+7+Bk/G0P
3JaL9TH+1v53K6r+ibGs6m9Qx30ykdlHZBUfXlq8zE8rTPBTdyGksyERZEdny1vG1cw/Iz63iSOR
d6EwB036HdSBYXJKs1SU9usWz8g4m6fu6i+CdLsSd7KYDpuSIZhHDpQI7TEG3DthWFAwYjbb2JB5
f7dK3M1BKvLQV3UP97ZwixvEMhXJUFbrzlor/VhyT0jGYxFJJU7sPfmZelny7669WlQM1AFuNUI7
YP2uXdFos22lDUYJ6OLmt+YU9BJUhRFejf3cH6EhKP40IfFw4kd3Hvtt8mS2F7Ss6/texvvh34BG
azNawfCiEgIHY/gkq35xbniQMmPuUg5Q0i8A0QJwHXQf5PntdDT3F4gWYsUzrAErcMoPRIF6iVf2
cRawMNN/Nu5mloQ8756ypQZdSwdX0cNNuqzEmEXa9leA60f4f/X0eQsV+wUOU0dO+F8HHJal/tFf
XmifsIm6tS3PFDuQnCmsnuAlfdrQvgttGVOyKcutBAKlnkPFI50hQ6ue8QhUo0UJZTb7lmjx5qo0
02tKrK0bvPdmDYHDhTs3tf5jbgKD/wLG15pi9szY8vkIJYe1kKdLiTOcOclZma/N/LpPd3nT1FLK
m8RwKnvnfFnqarRtY0uIEd31Kt2YxSb5apOfciKiNw1FxVGoI0vQ6pCalqxJ1fQFNskylMbpM6jP
PvG2mrEE1dmqc9A+05qKfDHRnk7/Iw0dWTg1qpg2kkOK8jhsgu7qnNtxaSftirW4J6CxvPdh0o4P
K6bM2YXG4d8UB6mz73nz7XJNO7yfH69/dmnaeKNUajnbsvNR7BAhlGRzO70pWhAK19U3c+40AKfC
C6ixwPr4csQ9cf+Uho7YPlkrF4VBpy9K9mo2Co65U3hW0D/ZlP1dqDBqJVHRTbi3vVmaOwIRk+Nr
pEpEf6G3aQbVr6uZapqoTR03usLYq02F84OARx5CKR0xhqy7CpaEJw9joSxuebxJhcbjxBW4DJtg
RRXIZqabaF5cJzW3hSxTmRGJbVO7bDkMGVLqYvrKaTECT2fTwi/C86CM68Qvf4Pbrd/DupDK+U/2
eOXuFXfqpaYtQIWewbolbWDR86vEn7E8qbduHBCMuJY0hf8CPRGB6kb4T+TUqsh99z332i8rfc8j
7rCvtyraVF6l/rSum+HwlYBu/Yqm6ywK4z/EQKG4Dk3pBunapmzi9XqkMUK1vaw4Wnl1fPAeZdA3
uoM7M7iDW4qC3JmTsYt8/rOlI6Q7LBao5vnZ5ZaD/1jVcZqdfhxtIVk375MTYcayOghV5AxEHE0S
fOI6AnygVD5eMuTAtXmR78RgxtlaHHlT4p6rH/rWCUV4VONjmd8v1b025AycSvatn+qAz6PERpgp
vJgs1Sx9mnbIbVR+3n+9YNtimz64ZL4Lhpe0vnrE/2wzbzYz/64NfJsNknlT13PZhlPN1E2zcQyG
MTbUqoJ71DQOGbjPsgorXu7Gm4UJjmeUnR4g9LHGRJQ1b6M6D+cJpUbQsE687EnN58V3CbRUg/Db
lq691AlUtg/Fzdg+MJKwlriDE+PXeIbsOhFmLfR9OILk2EVU0bch4Y00UNssFIZZcnfVQCSr7uPk
YfYvKxpDt+P7IR0Qf00BNhMFF74TZ2RfhS+FWUSGA98ePI2cNSB/LtS93yNXuNrN8RXotCAX+3Dm
uaAgmVXcSjrBjQYhGqNoszvfLApve0bENQ4U6TDoperFotMztfbKNJz+Yr1k012BqUbqmHqlr6pU
SEvWnKG2RNpPlWlkIrS4xgVOxBJ5g5gEfzjoz96nUVcfnTJfL9wsOq7nPP4igV4Fhk+z53DoqhQ1
5uFTBWaJqqqIh/Ax7YytprHfcqRJ+VXVaRrqbtrI28ykIarTjrBwCDRkcBfI25rQyEwgXQMTzbPL
eHJKT7pV9ZEDUC+XRJwd+WFMS+QLNHAh2JjrLBRJOPmddfRo1+LMexio990l++6lIF2HH8lhvkV2
XFwXXZgmw4f7QfW6XVEy2FpBbmugPUva+8B+1asbWq7seB+kaMIpEFl8d/Q/vW2e1bDg5oOtIK8B
7KmmWr3H77z/8dAx17DEiVeXezxznHu3irfoWlmuMX5W2ZgHhc/kZ0tY76j76Orhs+WLR82mxAW0
ATO11bABZzMsmEUdo1s+GjHjB8nxmmMEH5hPDGW0J+c5qWH+puuvh7MCvTofKRjff95iQFtrMHzC
OeJQPEPkdPZ4GsaWH1+WPSychj+d+FUlzlRBmaICBqFbVySDGUql4HazFy7O7Qnwxml7mcEAA88A
o0DATAmfvChBHNaRUjftIrIMPPfxCnhf/mrnnAIYcj2qrsXyw28K0y9rGeBbGsrTLeDgs1x7OMvC
fJMqns86h9SLmvxOZ20gYEX2SBuczXcbhujDRa9mhbAlvlSTccF7cYYCQdIsVC3sL7/6KzCYHZid
FjXB6R0bJbffjwYDbkWSC7KHPB4NgpsvKMwVgwz8v57Z5zyEuKqh+9sCE5oTnyovlGKpMqyT1h1t
QDy8io3ihbxh6IVvZbdUoTb6uoNvQR0qt3QE7F9SmFkAimxOwJb967ouisnr0RgggPi2YNBKr8kM
kAFeXD9HmlayNv3NOwmTH++OOtNXZjsJHGLogFdOxWYOquCyvymujw355EqWSnPLiJKcOUq+6kLp
0zcYlLqKGgQy0DlWcgAAcrwKAysItDLoeqIOBagZEW5VVXDhx1ygbhAXYnRwzRK/IQxDllFR7+Vq
BS4DwRxILBGhqgL6yfdT4gJLF4UC7I3f2m++5avUfNQqJZ/HWQxl+IDkoXnp+/WCCLZekGmHxHNh
0Prwe15NJibIYkzXHsQLm2wh7Phau363zWN4I3TbSufu8PiKcqtPHSE7/5O3J01FcqDjWzoUYEjY
5YNxpbey1Z1YlzBsXgfXH4NPwQ+ievsWRh6dlexXjBWrOjjUDzfCPFOSMGQCjolSa4Oj0wHzlqWh
ysDrSA9NgI8KqRhe1kVL09Qqv0Tfz3COJKwl2vgTyJrMnE2RaSIG8M/H/B9j6YG3hBJroMHRmE85
PYkjWS45Px2CN5CtXsuwPYObh3K0ZlYVzb95CYp4IKg5BgnfHidMiZLKmbtu2spbHi6VyWCT7gsk
pbIxxE2wbYbRACyoPL4AAXTeft0nTgum2AwpkwgK8vH50nk/f6RD2uD+6MOGB2CS3DWPFfBUf8sV
R28s6l3JPDU2sUvmde4oxC1PIeSB8ChZ0sycrcuxK5rxhdGByS7Lan9ljc0WzaemcXUEDA9ryYQh
zrFRfrOFp0EmGs/J/YVBfkZ2s6G2fiZPGOXUKIQT6YZtyQ0jc+tyOthsafBjtV0Sf4+oCD/rIc04
SSti9pIP7UQ3kZj/LcQjhYOTg0GtymOQHQSTL84YMn2ARFrZhv8MWNznw5ojgPOwjeXZVI2LH/f+
iVBxABQgaCuSpCJ8VcLGpixD5ACHcIR0OsaoMYkT+g3M+YXL+MmRjfmXAzOrSkqfbS2s+HdQR2HE
LgtDM7cyMCPByYDImjXABNu1KZ4Rg/Z0QnjKSkKp1RKiv7MuySJUxw/vL5i8mGiS2bSEUNmEJ48e
8pUDOUKRC/hmUw1OQlalnt8DKxHVZkmBzsNs1Fcw16O6fEo0Doop1KlyZZy59ycehdI14KdjlMEH
1GObY7o2cdKRit9HqU8SS8KhsMwZMfc/c4k4fmifNUyncFjrVOfzr+rzv30AuB7txwCAzD2+ibZZ
kJJPY+L88iztxw84AkTEkPZjf667LOTIDh+PdlR8ax9k1mB9U1HjhULpZcAZ7WxnM/+h9wSpzn+E
3CtuLQwREli59MqojxqR95lP35Dt041QMAXfPLAutO6noe9KcwRxh1oNpUuLhL4/KQgP7o5Gu4pL
hadMa0KicyEfD9tkUvRhSVQCHJBn/ViZRkTOVTP/HWxScpk+bCgn7UMJR96iwqC/GsdyMiykWJhX
//lEZuAdAsMHpEX/P2pu6rHNE707f11NKspdLwmF44j/CE2WIElkZRXZEKCG5hZTwooUvIPXz+n5
M0lrWYPYMNQBabkbzg9KySTlciElcUjR0PvFyP7WTSdNhjlnRZqk2Jfd4eWwMG6VYkxUkztoT1oc
Tx5rLxLFS/swOQhSsbkhcuyjsgd4VLJcD/767qcgDwsYNeJy7oGjydOjWLG5GbUlR7zNFTmsxH7G
bBt3Ub0Bm7W0AD1V2owJXtJbRre2XbMglTsNSIeKJzz1nwD6zMGQH2kxmcmyvj7VahAvndUvb78p
aHbSq1WWvCL7xcCY3LhuRBo/uD3CxeNxhyuVKZcNbmNHCd3LzEByzBOwbDKtGH5LRtjA852o/6eW
Dgkg7k02S35Nzws2TPDbLT8lr0tHMS5AEERa2oOjU91YkZgntk5H9Gwp5LJI3k45MzzryWVTh4O7
SyyB2V/CGjD3IKLuc+8l9jynBaRzN7q8uaKULc8Ip5uY3zjjNPOKa7P1iMdC6dy5oQGjh3NyHo73
wq5ORXDGhE4B/iuX1Rv91TsrubrErSHIX0gtdBUKHqNYE3+8e0AEZjU+jFib6dI5SrATg76Y0tbB
l3E/3Un3Yhp5ER0Mb9r/YiPqMo8OVMOUe3TyLCnFvz7MzZIYHmcozUyRUgd4h+yj33JWhp7vnwDU
FZ9J+JYXLRO9DyX1FWks8pU20YJ/+tDXluThdEBfbcLnaJ1fHf7tDY+djP+Fi+Pn4G3MLFuuhNHd
GM0kd+2TT8XsAMyUoyPgb0y/PZAuCha2ljYWHBB3oALmtF8kTj29Oz9+sYb0ycU+KCyWRLHYUxUj
iwWSO7vjGxOgSr9t5S/taDixBsx02fl0typZXVm8dw/UFqJjmVja/mNWbmq6pG6iV1pR0goa1uZi
bKWe726a9/JcF4Cs8ThzlpxFLNLh4thEsjkaOtOfUCzZLe2qnbMZf5EHlnShqvL6VQYnyelFQKLa
mkGgONsLpw6YtmEK3zMLFkhWHFsCjTGOtm6653UYXUWRYNiYSx4PBP1KNhqzwfYiH158CEGKNY4A
7G9mcS02iwS6aWHMmEZ/+sOGApFjaQayS2Vk7+OWdKV+yOlZz1FHzDYoQDL40ya2+yypthdhV+zm
UnA671YSBSvBm+c/fIUOENwql8+BUPAgczhRs15y1Trxm9bIGx/8bRVj0l15RlDy3tEedFgnDwcj
9xu3tW1qM/UJZV10OkaYRBb/jcjiH6AN0X5dopcGBdmXAsi/NAXBnFUdBaaPNuUuaVOIkc84sp6n
0QlP+UBFaqHOWqae+qfG/L/c9fKrR8l2Z5koV/9rFaumwSwguljsPDllI4BWXIPeZmKV0VPVfdeN
mvcOdJBEmwhJEeBzauDlV/oI3+n+XYupeBrjlLOGHbamiMJYNTqkA4xFsGlmd8wJmgbxbYKRnsVw
5q5aScetRP1jPJGk5w/SR8fJn9qMQ5KUOMKCcZK8c5DdOAfZ2XBj/253EKJrCOyAoj6Kz6B15LK/
1tYFpsMiUyyIHni00JBvVdK8otHjrjslm6ZbnOM5b2EUGBjl2Y3zlWwW5bkMT5AVdNdaeiCcZUs/
AlQOwonONbZN5mufxAddewTc/iNhkA3KoSRaxVpREMTDdhoFRAkD+7B4xmba+iH68l1mAyJoHZY1
BEp9UPla4uoEItVWMFY9bVwtRBUhTMjOJVJW+vKUMZ6OCpvuVoInYIsvnoGRYMr+nbWqtVOxP5Rd
Rs57hHMiE9O928acTwVgD1M8M1SaGCCVkRgGxZEwEipiHQ9yzB7TrfV/bsm2zEJD8LG/Gqko1S3/
yaSxJtaPUz1Zla8nhEJOgnFHQ3x2PxfAd1dLqfRf2qkQWkQWgwZTYasVQFrfARq2iE8woFQ508R9
y0keXUHZkymNWx9blDoBp4VTz9K0UFXrJFOE6ljj7eJEyBLHMWPPJ6wI3+s6og3Ozz2vQubuAxiW
/5GL3jmvV9GuMEMmQD/+0aVArjlKAAW5HyAIXAUCaLEfofWdzRyxFF8vN+9sHJl7JbQlvCpWpnSO
vBBjDxuNhXI7g5zOyeFqYmZHUidfd4DmM8atHfVBPz7GZ6gIYekSnwgZJkXR9MNUhdhcOVV6aZln
nwM/CJgqbjePa3JKOitRbvXM2JUmLrvnfKK7hmlBD7w0sxwy/jKYIsbjK/2YdvydDIgA52//+s2n
+FWYPUekRN1gCKajjx2Ake4KIOApH3I92xhjXElztlLWNgJPRAHnq+rYcKnUOK9+juVTyWH3sC+R
q0tj+GDEUF9bXlHUdiVj8AZ6mu5rkJBBUSd66HqyK2/3pkUHX1rMtAjCyozT4pOZdrMgwxrIOLLS
zgEUEXGUtULM1NQVIFzl0kYTe8Xgq8mhRG/m1jNX9JB5XfKHqwaYjhASzdYp61i0gX1d9oEgLOC7
fbmWC4elt7DFm++PeLY1ob3eM1ugQHJPkh++ZkWyJVdoGY0Y0HbmKF8+4wg/eQvonuDYhIyGDbaJ
ShM2k9sH+TtxVBhO7GxOajPiwAK+nxTAbj2GQ6Ev5rxfpeQZE7LSXk2hdPc3bF0ZfEmyJwx1Ib8z
fimKw/NETA8GDFvQp5OXD39mipUGGehCNZrvqj65Ygf603kn4klHt14qoy8ur/P7CRki2jZ295B2
YjoeTUdCqWPf6L/d/Oh5sQtPCvunzi+qFADXtsaaS8vbCLp4czOprQ8hP1npQWbk0w3noPPjpMNt
nIceSg7j4P5DJQrOVy9zgvlNorZLkG6hSoWsskKICL90VYcpP2Iil6gCK0f5/tACqF1qQYQGRpSu
CRc+cRXz6fcdXizebNp/YxhQZ1ir6Urza3aoJ4Ycxt1arHNfIlcgb5WzW0J9vAJRlzWtfM08wdDP
KBUYQZFkXVxVadM9pzP0KFySGBop0N4X0aBJ/MO6hnc5TXn7TlA17qxwUv43ymyd9aYBXVsR2de+
i24pyqqPqj2neYsI6RbA1teLtQ0A2yfplOTutLh2zFNX2zScjw6CJ//EWm0A0lDFOZjNxUNMQKzT
yl5fYqF4kYhLidK3D/lPyNbbKODDLRxJCj8cQW5O/Gw5BoDr95MzrsPAEzkrTZGNg5M1Ju7zDDLD
4QGVF3hVvW3Yml00Ht5i8zVgP345xHpnI8Wf7ID8cgk3D8wpz0UHIG8qL8TgHBRusn4dbZkd3HSG
pbtLys9QI7Uw0G3KdePrZLN80ODkrzw79dLTrPrFUFSC5X52IalAvs0HtJ4+eYWre86vGOfC74+l
rqGKmjjThaz0a9+vkipfaFHetvbNhPZ5IbzGn1w5Gf75V3Hyad2FBpAnc7Ejs0GcdXUFUj4xc896
4thf6H98mPJ43tojsJoKg/2ow4W2U5y8rRIYudHlHBP/fuK+AQU6D2lvkQGZCNvlhhwTolTXiYr1
6RI/5Tp6zek7gGqTCOYpZEmqxlI5RPCOfWB4/Q6pkQxNY4ozWAhx25yWE/oU5JpFWtuPMLGPFIKz
C/T3QW8t12TdLQVE6PbdkH+JlEN4k2dkig/gQ1yXJTmUP0uUILT4f4szfBNHpzhAg3u8LxrKpTI5
jEYNl1Lxg89e+OxzCGESe9heYn6JUOX5rCJDIMY2sb95O6Z7x0rRJfNxZC7qqwF9DGxk4nBJ+Gi6
3Qox42iJW+nAgmbk8I+fyZetA3CeOJVCJIbx0nllU1DaEnTctsDJl3asWYh7gAKnVx93CtJoZDQF
5T/eIaeYzGUhr8lTYoNnd+zFxJXTqmh0rMeCr0JjnbBf/MNPQCHH1eD5D8tNzxgX1eNlZxbpmD3n
ShxwZsEcJrIvyxt9eI4EB7ZFeoTwCVOjO/7KdsE/S4TuDsn9206Af7r8Rj39MYl431cFLWZFIRoa
lNIDzanMmmn2yjzwkREpA7DZfiJi+5AAH3YjEmgN7gmvUxcxSBh35c22WGhyE7Il6q/sRgKzPhCj
+n1U3x7rfw/GuMXmoFOY7JHsOOFfMN5gRXae+zYvhqolL3mvb1ZNu3/jVOKBn3EWgcXKJv94PT0U
uhZ/EafIhQqAkiT2Xq1xM/arfWy3SRMg1EKE5Q62Ol209WQfm0N0dB2LM8r+/fk982eSlxkL0dKk
1rb11xUX2bcJzZss77u6dXJ7mkkR5dKCf/CN7/QM/ivof1V/694YcgAMz6lg4z3aJrA1HR7pEuVG
hIGN4MQ9HJl64nwbRfOWEmSJETL3f1y7J9h1o3xBshvfZW+HvxgjmHSvm9nBjoheZcErYdmwtB40
yedzmvuFY86Ui8waZtQ3KyP1y+X3a64t28QXtuz8tQqPSFME5bMqQRyeg9maI4orPsQ+HblvBzmi
jPKjTFBXeEX/x4WeJDA1O3yC2QBW8zN6cBPWPK2E5U4USthg3+UwyJeSw/N9IslFBqS7Wavew4Ep
V5tvB5z5jodhb6C2BbnddfhrbAV61TFjRDaMGzXwId1SkNiC3cvZLApKBbjQbvgNxGMYxwVZsHxK
EAuQpTZyWxxTwD5gJE3E5S9jPq3+P9zwQaOitOx/KMolEkxhiHaDo3y3JvScrLeHBKHT54sMR58C
LdEN1s3bPMwnS6bQOIAoa5U/TZa1/XkzCLk4SxUguKFDxFu4hrquMxT4yMwfRZUfT0zn6SL7jPnn
37D965K3iIwbVqCEh7DSORH3lPL0qI33CTrTp3aQ+AvEYFvFKAVB9mFcTU4fvbsHCHNNA4+C4E1l
ChQDXzGt7ah2s6jlRDFEenev23Pf3mRDyDzX/h/Qp0kXw1IGVMx0jO/s5OWx9CzPUZwquwZX+xKU
qYp/tw3P/KyHw/22FNc9tHuLDzjZ+FOLwjDd8aL7cXxjR8eT5iA89wYJc5b94hk7Ak8FzVYArg8g
kgmfpeGCzrbsAcE8gHaRUDuhjLL1OraJoYVVsT5RcckA3N0Ml5uCNQPvSU1usZXiXJEavzH7sG2u
zBj84hWFuOWIe3MTBrEN6/QqwUhfBQ36LGcb3fYs/QGcwdGZB80+Z7ZgSW189aBHHeRc8bLKVQ/0
Duj7DBaIYb8o41Q5s1kYqH+crvFThe0WxObps0YsxuFfJc0NgmVJPns1syA9pJO26pei0prgjRh1
VszGq976arWa96xj5evvGmCyPqBR1LZ94Lzh/9AawFhp+ZHL6l+D9aiVTFmnXyAKroF/FhL82t0D
k3C1uVqCXOoBVZFdLoJH+7K52J5RuFGKBNn9jabXP359XnTKgfOW2mV9Cvv4Qm8VCXl2NSyyuqpY
ED8MT1RNa0NG0cdbWrsx1XEf2/x0WEtnBeZ73yI71MoqYdM8RBB7QkA6PSITgrp3MLcDSDyUOimG
Y4gpsHP1gD/VIpEDjlUtp98UQeQz4uFY6r07vLNXOQqPSJSWQeV44GZdyWY3AX2fOKfv34YSCsft
LBVNic/q4eogGvRQTEeeldBwQxTdD9PM6C4P1Cg1fCpbWdbyGjBf9PJoYTV1bTun/fmbDeypWlVX
vL44YHymxujlIXK1Bmyhe3PYbw/g8zbOI8rRKVnz+1xess+tbM6/Nv/QUsUnInbo+aEIpfKKlzDt
l/ypzHrLL5qlFFvRF1AprCS9FUmxkEQ1OnKK19VMWHBjz7+okWO/Nz+8+xUa2W6GXZBwro1hrbWk
A6d31YbfsYV1qcvh/fXz18M4xu9t1D81XHbOn4swGi0vaq1y59JuvNBHJcEbEOkYn0zyCkpz/i4Z
uWuWXizQK4DNUnfGlAPtiJjVyQ5IABGzOjlmjV2nzsbhvlVOKKRFNpnnUV6dogka9mQVllV2qcsh
Qx3bkwlpHulqoherWdailiMh2Z9VRdZH5jEwNvr17+jySpgavd2ZtdyMHI4GZalIkCWP1ySCv4Nq
5c6fW/xAGt02VzvGwC+wob5zeqN2PXqw+KWESKI8jxlhIUf5zZ6MNi3RFcUAWctKfOe67D8SBG2h
kGGGSG3HnTm9R43zXvXAREFYqKHpUOwlnBP4znwNFYHYLUZtWpm/czp+j3nQCtIo4U09CC1L8Hap
xIhpHktwtdLKB7DaoF1qH7B8lMvC/NOzJgK8prrdk1r7lm+5Ar13Pg1yuPKgNY98LEkUFOnU77pY
QjFPUe6gdsBoMtG37794oJcaFXDTxQgL9zsrKkOsiFOS6U9RlGOhpaYpRqFb9Tf0nv2RGSnVtbF9
iNYZ4bSNeI7gSLZcN3mpodR+VYP3IrFk5+B9NAb84fmCoEed/zGr9EZ36ZhEZrRomn2YjjKpdS8B
slrB6SR4mFSvr/YEFSgdQImpuax4PtUwiTgLSKv8pnVchEM1aPBAa1ZE2cIy7S0pXorFgFriDQpk
54kyB09EHO9BibJFw4S20KSlBQji92mNJAvYDOWKvs1MfOWV6whpwVB1Kwiu8Bq7wVu3lgrWxLwE
LTssI2j7UcNSQygIbUW1uUn/mGw947fnCwKjLjQXqCefQtJTPDZohZX7IFwH8chHTID7mfZt/tRM
ZVR9qWriI+j9i7Cq9vY2gFMdUzMviMawQWfnd2vA+AKBepiruaIvIuGu0PCm+jGC7HN7Cppcq+XK
scJuLF9BbApJhND/ARQNtdh/YhIgA8yHaRzOhfAVXVs7Ilgtu1QpJ9iKexIZsS1IhnzNHFBUY5Q8
auxXQcUz49FmCe6Qztit5kqfwJiLI0HaOYiU3VcwFSn/sQTuWZwislzSiGWlF9ojOC3d0ebB5L5w
pdP4ruw0hu6o2/W09Qnw0QeI69pVO930OoEBSYFhv8STNOsbupQxggYtZeb4IWw6p1zsr5VEp+y2
Em3fF0bPbwRq2qt+gC7lIO2B+9uIPR1y2GEsq1jVNZ5rKbRUnvrVHa+EA4EY5ozpRE2JA1jX89ok
khOM9aKjyQIlIn6OiFklOkvwzOaLjiNIfgrXNO1A7oiHYQtcdjPtQMifnGVhhuaSJAbBq7eRcR4T
TKOIWgUvn2JV89CqR79HEIFzZVQCmM3V4SAe6LSHdBxvknLCRjvJgyXVWNh13ftdpC6MA15pEH9L
4SJ3+jUb86jb06hsEKcWM3NRKy0SLwRszFzABUNjWW2MsnNeGPvik41s5b9GsQW8Kk+ZRYkdBvsi
Sy1SNaxtTNK3ONQw4fue4gK4DRxBTmu6LEdEUSWkrSCBMkT4wzjbQMbzvV0oN3sKuojBLokMv7GE
VHYCKJsJZIqEyfa1PpmzZdcc2QY7tv/uO9RsgK3vkuTy4JVBwb4q77W30WY4y3mFkKzdPfBUkm4S
cu5KCCZnHh0CHJaWJRIIxhm1lIx2XSxj5KxYeZpBg2R5J18QY/3WMGS3puCRbxOFtf4u0ZWWLjtR
FtJhRI0XHB5/FR5in333kG1AvoT8Jr8oict+4uLOCC2AuKovvU7HkHCI8mtRV3l9Gn5r7qb+FVSG
qQ4odX6gUI7bb8Jrtc//tCRimZiIukGMgVNwoEYmBKAiyBH42TqiQRCA4DqbklhogqV2gayUDVC5
MrVyDkzXfb+4aAaSh9S+qiZjBFxcHPpE1O/10rl7HZ3m3riBkTY5B7DRYO94XkSk2Y0g2BvQNg/L
f6v/jExoDYog22rmrCXD6a7/m+rBGjC8exykif22mAfRNvf50qpmnWjBhLEGPmcDNynENSk6yokC
AKEu0kjg5YQy0NfJnDuz2TWStxxb/3hIe5jLye/67RQVb92JBxSjR630/NYqTlNnY/YLEMSbd3Eq
0H6D/DgXjkPiSZZ3wUnWcz3Fj5ZKkEtbd47fi/VRCu+hBpSHr6KHOkmZ5vNzfQL+il0So8jE8svR
a8O1jkXMA2BbYfhh6Xwi+ko6ZrH+oV4udyMxu+pssa3TbnA3nShCc7FzGAd+E0mcQFPVS9B9C9x2
Or+HUo/3JXtKGFDMgbfDODSjhMFtxm3BuYA39eVq26fvBw4a6LvfB7lfccH4OaJpGoUgzCCggsp8
I3b3jVKKEJb6RiVL7eywxES2UIJ3/U/xHrkUrMIDxNmyEekMEOMvNEKdY6kwPLQoMeYzQY8/CNsg
7hiXgqiks02rKV409QmlZX6hJjXyZO3LnZW/Ng6dUDqgKK3iFOv/+FrlOlZ5ZjnJQ4G7NqmmblUo
Wh8YYa6UmW/Yu5R8Q1/H/nEUmF6kn6gRyqSWY9S4q8BvMeBPt4SLM+WB5BAYCjcyux0dVWWttYlt
5DOUQ4dGHVetrQ/9reww+WBaJ+3L9PkHYwUjUaonocq82qhJ/UlcCiuwhbiSD6C/GI02yGwpl3mB
jPXBCSxHr+DGExddLlIPwTZdGlrW8X/9BCoyyGqAV+Af11knuTVdQlzUQ7Mb+LGQzfssq6NsTUMz
aDmcrtBHDGI+tGKmKmkNykiTP1bRhES1Lx9r8E3t+H1VIJadUrtsk+VyA5glgAJoozoT949snFLY
djzKZp/YNACSo8lH0mg1JDALigvp4sMfWYX/Kjj8CqwuuUBj7OV3s4Iix5NNktShzEpJuY55ZJTh
rAurt5lSOnqJvfOlTZuacreyee0rPCGJzHLeEiS/FZxQXyigzLPMj0hiQp6gV3VaGdZwxXjsr8QQ
U8UzxBFJ1/GwWI5DEaWraFX+K3gNYv4ilhxSUraJRNcenczhFtb1wYyMUNbvf2OkW0OFx9CwxO/v
2OAE/Ul4+2nYUNSS/GMj2FWBHngzc77lis8a62pNaLccu97NSCYOmkhXr/+Flsn2DBeQ57cIJhkg
3vqxk4MPTLEYG/3geM3nHvUMo6WTkPZTGe0PNEdcZ9IdLUNLxn2Vz4m4K1QnuSnytWrVMLuZj1EP
eCCzif/2FErcY+9W/7LQkDO/RdLXNZKvGOpOLF/d2JsbsFMKVfx7Ew6i03M8x+Fh8sYiL6+7eJ7I
hgwnEVDZpo3HMoaGdjz0jJyFHsEio62XNV3lVSp3U12jfzIa/g5J+b+w6rpxsJt7+6pJJQvonEYA
8cV6CJW9If6G+U+pK1iUO22cCovGBetpZXEbcgf1mMubOnoKhKp2NAoggNJjj3VhG1QLWD7Rx0gF
NqloD9CCRTvlkQQm3Hu5NZB3Jb+fbvJ8PCfMP1FPW1mfWkaqHVZUD/hv0JKE0iPYlKJiIlPizwSt
SukqwNovJvNMrBnUwMuzuThNQf3yF3ijAChivF5Mi+0EQ0SMrFeRZNB3oZf09LBpv9d0ZzezFFFG
5BQbQPaKm0niRuV8os8GikutogFsR8s/eF2k0V+QRvzG9U+C9X0iCa6C5mMxu+sGH+DEgrsl1zxo
LxZrBZJ24hhNm1E5QX4rqYMKCXpr7a+r3kbNPt7tAjg3Zr36+nWhMGalVFyKLik5dJixmB3KahyO
EJyDEwJjL7XsCU2RQa3o5j9uPVjEm2Z2Z2oH/Bpf5XOElJCx6qHe4bzQ7AvpKRkdztCdyUX0C0I4
KG+0xuVW0F/VhLmyW6etF2SH5adIObMz1j/yQ04HsOM9jQDZ99wCvDq1MPi2mclOoAV3gASD4jNH
D5YxLNQ1amoa2w6aLGiYeF42SJgQnvgPnU6x1jzI3OITCT3tJsWUv7nwfA6RpcqtUhZGmpK7XVJ6
UnsFQwHQjLTPeIsEOTaMZDQbu9kXBHbkoRHoFahn4fK66ouV+fX1hQgLLNvhxcKJNlxYjopyZA8g
t/0hqpWI2hpP1B5v4RiX8+m4LRBpOWCjiFpLp9o/Q/1yIg6fTe6JO/RVHalUTBd5QwX1BJGlbJqd
gGNIzdqrt9P/8mtP6k6Yx1fqDjD5Ea8HMBN4wd9uOd8O4u7yDFWA0iNdyBgiT5vmZdnUX5RQU8Yi
dN7H0FBm0/6Hkdr2a1jVCswFihYBzXAR1G820MJKl1Hw20dnEpSjpOfRmCPmiMFGlXSChdAJvCa1
34J2KIGAYyZRWXPl3bjYurRrHirmyZba5w3aatZDXBELGd1dk5CrTHj+GsXnLV6J/F3rQ4fjHB2N
hdFbP0UBv7tnU+/lidbBBGw3Qu2oNaxCFFKsFu7+Ydl13NPo356Uf5aNzVPk1buRBieIFQFMURfU
oIXDNSNVXxTJbqfcByRVgus54UOHvwqNwr1Dnl6jv2vwF4Uu1p63jgzyVvf7AQWhjS2wPtMfSxQ1
TrX95bXRLYcXVfyZ09FoCr5nIufzfh2wQHIWO32Ss/vl8LTTFu+2IC/L95pKrrFuemCfix3ilTUX
L2DaAcMnPz/QCKsnUeM94V1fE683XRNi/3vfqtHpIamXbDVjzV6SQO3OUK2rocCTZVuEJh+/U6iO
550Ahy9AdfUnlVSAdNlZ01BZ41AJSIkO+IWFiUv1Sbbuq3dUmp8qGny6v1C6zcSGB5zKtcI7JYvQ
HNItJ9bBqizkS+1PlAFShPnMAy1jxwLUaNiCFdrqsg+BXv2lgeVmCCZWBPFzrC/a/osFlhTUl4AZ
J9wWluCVkUi0DVaGyEamqWILfWJKfoM+rdNTJ4nHTIpneZLpz5i7vGtO6uGNg3kcxRExsgYRbfaJ
6P3kyRG4+Xnm7LUw1ZvQ/EPcLyBIud6u848S742veD9yy3Lmo385077MAKzLtLMs18sNZyEsQ00T
wqTfCsFidT75tqeH+tab5+ImK1/VOSByy1nEHtFGEdeJVhP+/3gQNqbf2m9u9PHSzaBccFE5+8TT
X61b69sIvbBQCdOvzwGLd7WN32Kf5oZ+EFPBNUsfbVamVhx1Tj5mGa4ajpFcPv25SjHXBb0EH+HO
uKjJ4DxJbYQO4uwiex3DJeD0NTVyvybKL2yrzsCA3nUSk9qziG6bgqvjdxOh+mv+0v3svSv3jiC0
KEEv7IOVcJvPNkGo2KHsOvVhK5g8O7KasfodvcFvonKwm02j7kVZ1hsr1cNR6GgXSyLLiO8jB2WW
bUoyZX4ogBBWGEKtgRKimy9o6Fy5UkU6dHKn8fzGbDve5MhXckXrvhPgGn+txZESEsYnpMbNSP0P
Fh643QgeVQYR3EmUnO0p5FSXtc09Q36dv3mgiBBT4hVyZ8cuJNAQg+nEfoZ4iRMz4JMBxqPahzFJ
DERxxeea+C3Rl0eipawk+w9UVzemjJ48B03DaHMh6yUdXwOhBEMeZxRi1QbKQnas6aBgjUvtWFd5
pKiW47eYQg+PPZg/kb2Ox0MfWRYDF+EmMcQtnmxHKzWGqzD08swlSkQybjGZ6V7D74yhdsDMSdts
y6RCTx/V6HWAuyYF1DI8+UhrfXbYdCUD/sKvJ5vvfbSD1fJsP1UB4xt0HOxp+9HLPdz8aadtdfGa
//BqpO8T5sDr1/nMW9P4GGyRV1mD2CtET2oRb7bFiU/VH+fNE88QbkIw2/xTLWqGg2djw30f8omA
iQpXNejg7Cenn5m7m6DBJxUvK//0RJp+arXHLErmi6wYTqb9Vtsp13MNvRMmBgWlLBCiu3Nm9/k0
wLvIoURkiV7ZJajESXrwfM2HkN/J/F1xrA6XXPP8NYgHT6on6Y+tOkbL/7/AgRqXIDeCgb4mAalQ
oXiDMj6jBeYFewyWz6npcwmhpHd9ClH/E8xqW922z9pUq3q5v0fS8GZ1Zq+InQCAhk6PNzsflNOi
SnHip3+WQaWLhviSXxOkrfCAUQ5+xNVFd2R3sd53hbNYdmZGw+9znfb39DINeouxZwmgDr85q5m2
sWYwW6PAZu3ZD54+4wc2BZcB0si1o+x1ygGFBGaxecpS8bgGIF5TkJO6vL+gJoCPbz45cxLmfsh+
L3tCYhc96knNozfS9yAcU43uDkcccbPyRHx3pXbeNz/r8H8ucKDZ7iLaOJAWjt0qNKwhuDAXwUXh
45xXBmGR0ptNjHp5vPzxCYqN0jR6D0Cz8MmkcEjrvtwZ2A12NVbwhkR3c89VC/LtAy5iJ872kHpY
A6qcPVQyKbftOBLyC/BtvXz/rTPxkC4HYIAGci8zUlP8L6HK9HfUO7mG65PgNwso2TnHRomov+2n
/zVoMb2wo3CtfW80ZRg0bf62kCq2W2LjsBMbK4trBnnMWAkS5OeZdFl/mXJX1Cez5VxdRz35Wwsc
LA9ks6AYiBzmZxLJiOwHM00zW0HGm007zBGhrYQ6B++10cm8BKa2UfMchyRQfGnXPSTYfqNK6qv0
W7EStLnNaVWv9IwPyHnUYkW61TEAsjVNr6sXkIQz28bmVQ8D4JTR8oTLj0TK7Vy2DGJkLAB7N96Q
k3w7j1YGkOFMwF/FWv4l2b8I7BW06ILeq0SPLE/Ebg94bYAE0GmEL0KsRrPbupgiGXO1U/blPlIY
8PC0CXRUYutY5hjJ+rFIRxzaphxfDnwusW0JRh+7QyfA+7WgkiuYv/FwooNkqXZuBmBXvtbaKACC
lJb6DGlh0lqw/dfLbW7SdgilWSHWc4I8MS66Ko+5fcgncUybhcXgnGFyJUfOmcvo0yl+d3HMyLku
J4j2HhUxACyuWQIdl4kYJjYe+/KM39obF9VPuwYcGThVDb4rHltxAkdgC75r1MdeV2FuAImLkBA3
+DLyIZuR+US5Ol/LRtxNY2P32pVgQ8nZElrDH3chXQIfZUkKpx+GNW0lNWlheNfygXkhxN9FC0sN
Ip6vKSytpDucX/xqrjxR3tXr+TW9W5BWX19D0Xw4+FnISwGzsvmzgHSscuD0jYy0w9k8nPLY9boW
lUMZXdTUgvyLEIez03nsa4brMAI01J44nA3DmkByDrj4D35r+YvBwNz4d0GZwhhorZttpNK9asPw
B3+4QuAM68cKVvyxqdLOLnu5J2l5aG6KPMGvC7PUuHo+Zu1NPd2TkKaQHfqAD6bv3vQuNaXKWtBr
lFAZVVWSODeaQgC7mphFsLyonwxcCxXyiEzyGZUeP19Wn3XBC1uB7lmRDoAzjEFOLrW1RQS/K/d5
rAXVOxZRnTxzXmUOTCi7bF7zFnlPlfESdFNFkVTLbKmXYW1kmj0BbLJiXeShf+LCK4yTEH39FlaD
N5r33F/+Bv2imbprgl/tDNyNFN9OCo98Dp1oJ0YC49DMUzp+xOInAqm5WMzd3in/N7YKYkSeGMaR
/dbs5n5klvGF1otC6Ug/uBwr5mU+MoKzpuQo0oxO9j4w4WQi46JvpJuJqxNCGx2JmR3wbj1m/IRw
N401GyWQ7qSkcx4GEt+flPt/YRSlycfGcMzcj9kMKUQvFZgUCcOsSFMNMR6MJPHz5u5pjGuLBmkX
D1WoLHkgDvjHc3gu2qa0VWGSouS5/wT+d9II+vSX+M4gxMi3qk95CBaAjJg9hnDnIaMBqfuuuyR0
PSnN6PR3kqSF5Ss/AV0c9ilPIhuSrTTpwX0Lr+Vn0JJ0Qgv7IGCyfn60gbcKSrWKIFFCgcrrR4fe
U6brMZnUSlfpjBumwavdW3eUSFH8/xdMOhrkGKKpQmLOjcpbbW1fZjylc82HN+47iCc993J/AvOX
RPcSlOP9qBxLxJL24GIIrILef1/RR1xHYou7wMyGFhuMMtXoxPs6sEF4dph0+uHYRfrcl8mHFVYc
vXWhQWkTMYNWOwnL0a3yI3lx6/bASvDCaAH6nkiN32+oG9kPcxTxYYQC7jhIYU8sQe675pRO+g80
Eb18z5mCGYwvFx6S3KfMpP40x6TFKCvtamJJLuNnuZMkJ+jz/Eqrd5UHf2vbsIVDQv95fAh2qxM7
OLxqPte1sdvYM6HH1uNf2J6t4DrPHB0M8QstCEPUg+zH+NRlpdNUWf7h7akAhENZHlDldID5oBYS
3FZrWZpb+KSZ6JTHGzFqPtP6zjp1YkP7EpuENPAzk/YHhf2Z127kJBlIRyfERhqVKgbKjEBs7VIM
YkeI5RZU5wGidfc0Td8vq8acmxa05lZjIT1eWATPlx+Sdz3qzw7duIKh0Rd8tqpIJ6vY5fCrbLDH
Yu0poLBeccV3AXYoHedtDfoXm/Lnw/rroornxJywgFfZJ5bzLJvGnap8hlhpgckqsm2ATpnBU1af
S1yo4Eb29q7EhXxyFl62CJ2KbSR2+q3xKzKdHUIS156duKFYcSvjy6b4F9EKkJ3mUXRiAR7b0eXU
y1eHV+IG5bhIXuqYt3Kp0z+qM0SYuZtvq0t2Q8BmSv6boB6PGVZuJOB+4lTe8/qA5rK+Sj6cWvI7
d3PO4Il56CC8vld5swL3HOL0tq4Sny1DmRhbISyRJnS7cXWN6K5QKKtguvLPcGu05fvV73ZLNjgU
EcD+XEp2bq48ygvKbF6J1HCxQucyrIZ85MA83qmesgaE0M34XBDXRIkkd9GW0qzQirU6uJZTZKwh
vbb7rJc/kE4Ee7Bgr5/rVkELjDAQ8XdIEtZRe/ZX4ZeSjeHBiDKjG08KCXgHdC75jSntnl6G2PqR
jU3WPNYB5SBxK0AAtk0xc6GaM18nAOzWKHmr5GAgBnKPg8AqM7xeE557hKAqCZN7taocH8pDXKci
Yuz5Bus25Y7nrjp6r5u8nJNsSDTIHx745KbfFuNG7ySu6ylpFK22L2EUkv03Bx1dWGnGCIuc1n8T
QGDa1PlPL+MzlhJTRfqDXUHphrs1X5ZPITFjqVO8571DfhFq5hL2tv//K2U/nNqpqAywXc2WEJEp
sYVwau514o626qvjZ3so/o6IC+0iXH1RZi4aRWhTypV2HwFmgPM4IcQfgUwfsfyWz7hsUr9Q/qMF
hel98Qn25WxVbfUZwdVfOYC5GSGW16gsIs2Rn5iLrDKwOA+TTlmlqg2TSaHEpgNAkXmSzOr66pO0
Z36quXIrddDWeDrrcAgioVDesHNbHH46juNagvfhqvpir9x/CJEBbVmE+iC1TbOhdyMldp6iM5sx
sw9cAjRSCMMUsWOmIJJYJtPXLuh1nlvzVlMwJV077sTGVnGX347hsrmL7T4bdVNFke1XL9603DkM
dWcehzwcft+8mfH8c1zwaL7gMUa3uhbNYOQQqOFbI/rg4VAyRkmh1aRMj2EiS9VTcQhykysiI5Im
iSsM8YszgzJRcrl7aEfag8GmNP+QXtTjXty0G/2npoqA6SOJElcCc6WeAH3rY7eQ4FXPCORceFHs
uiOtHsz2JXeUXOrRWSolVjUwGxM/mXxoS24LbyLDXFuu9P0oZoXvqTvUmgMBopLSGZQzLWlAoVsm
Lj8KHbeFKyKf6zGoa0hmcxLLVn1V43+ynOvjqAifSADq3YkkXlgoiXr2uN8uwokcRIhniFjFd3A7
HsM/oSsQBzKFCZgmdYkc1KDpYrlls5vdYUTpXoPwqm8c5y3WLGEEbT9vdwjFDT/XrNg/W+FK2pwC
s7l4/uXhD6JsYv/SY8etQ0CYbwbeTvdFwvUHtchkjSK+fnAUdb5zqFG5uOTUqas53xAEIVv6FpYj
VQzKhdFaoEGv3fVEt1C0OPjiGw9nkFzanO50yEDLDes2YfrcC+ChkN8NtU+Pp6TnaJeJ89ZV3cZi
tgamuG49eltlzT/KDvsEQlwbXeOjchG43kS3vJn/jkrkYuzAd6kDZUskBhtP7UwG2ev/u98LUUNO
PT1dxiAdVPeR/+Zrdha9CGm+GicQdbVdboQepZsgjLCXDImwgloeBioB32RgBEwdpfs/VpYrbCVm
XFhkB7zVwPl5IjgnCCE+yCROgn4VGaFfsmFipFvkQrb+GopsTvGg3j1Cu7QOrNVmn5mcepHl3PKu
+aYTMKhV8aa2vb5m7EAycZEuim+tnZpPP9km/sQswo6v942awL1lT0GaSr9kmt/ueA67AHpD6BCL
Tmixb09YIVJl2PL+2sUt0OQd6i+wiCfjwOwAEvCG/1jF99M1pWWL5zgW9js2HSVrNjWNMfkrE7+P
GhFxiCQ317D/iLu6lZYjhHadbo24591E9ck2mtSLaZGKxj8WIAE2cTpZR700CIoBgHy9cwKY9oNz
th931C4Mn5HXMeldpZeEqhSi9CCba7Phgk1zPKNJJ18uxKQCmpGHp4Oky9qLkLzlc5Vl9vGTX2VN
vt1MBMlcQT9GhOigcqLR+TzPrIIWNQeAKYiCQjSIJNYq+l7NDnsrlGuNMOPzBfjGfcphU+1QHM0o
qCUJHwWSp4US0Z+ejq9HhvJpKi52AdGaqgrT5dz9vmQfCeOir2Bxv1ksusQG0AaFVGoN4etoXN/D
W8JKf0nzWETT7YEnA6gFZsXb4mxalN5544kvwLtWfn2JUH3kvTXTM8GtlCj86t0svK39OwLfCcG8
627F/OOyY8xDHo6l22VLul9R5fcV48iQjMGpZv7BORwmHcnQQf+ReKUAe6SsiDcuVQX0izNV+wKO
tSAQjI5wg27Cu5IBfmDkPuUETq/DwF2+0gp0WYfoJUaMKMimyMx33Ge1INlJWIhIhbXENOOZ5dTF
VS8jmsgfPXFYkrn0duH+W14fMV7uV3qx5ugcjyGgG3YVKiYSp680/11VQWmO5Dzo4BRXJvCzIyyd
mru/R5suIfqpBRT3r1XSS8PyUpUoY9M1tm4Gew4s4EvjKi+RWjNiBAJW0MiCnEFqbP8SJROInAZT
VCFZBD13F9gnJMCRF1mhBs0z0SamJEMPJKR5uoNxtF3aIodhTFljw0x4YvWK5p5sbleQ5N69Bpy5
yYkEbZ58xpjkvFimHb1KkK++RLFWTvfW8up2IU0webXwMAkiqyQ0Fw6im61oVI5MD1yfZ6IJc+GF
ffSQjZIZ5+VW4aCYFCTQLB5Lt+0JSSn0MMeeDV44QSMYOYLnGlPu5Rk11woWBo+Cl9EKtsVucXNN
wfRCBk0+sKIYl+7cuxTymlZLx68MKjug2RxmSNM5Rfmg09wjiXYWrWjt+EJ9hUnMv+MK1GNd1ByU
hUEHxnzwWGyb4KrlOFD8YlOTtVt0IDM3AZKruyvv3cKaiW3XKN14KyZRRbM1BlrM4Y0LvjNQ+JEa
Rj9rq3qeHkd7jFoIY06k3N+ef/0Dj62G4/TGVpcLizJip7HcJHsmS6I7dnZJJvnRMP2dOlcb1pD/
OizoIKzm/DblqjpbpgXS9LJECTIXSR/Ub3dm+UCOZJ+75un1lYULP1tRi/6HrazgZlQTysfcxVGc
7lrasj5RsChSR9mCdd/QcnIh7XY1utRBL8I9BF/V+RLzJt6btUOhY03pEle3UYkET6sqGytrpfWA
IxxR7mjNPStqTfx85BLGShEnbVxlfgZuNJKkOxZ4Uyk2R0jZhohho2lkTsZiJoh7Eezg18KH6rzE
P7ArUDSLM7iAeb/Y0R1xMOEeWNn0UsLF41gqSX6dZVaAyrIGlbAYz7Aj8FilwDz7QD/td75/+iCb
kQqP05RLqeE5RJXhZdix43hE4dXUPGdXxlAraUpV1bqyLBggZLEX0QLcF2VODdQ/Y1LJ9t+BFi2V
NricJBAVxG5h3gvsqxvy/nlbaIkLmmb6PFzB2isXjZFLZq1tuyulsUKN51/7tIR85FllmoKvRpBn
vck/TZ47RvyihO8HT7201FICb6hDpRzJU9OjKYL+uv/j+m6BBkFKLapodSofkeBgm5TK116fNN/r
UXd9EYV5CCpHVWilU6g8bv7hPfsSOukv3FFMaRJviFm4tJDcCs+mD6of8r2T29gcM99bPG3ZxZSh
gwy3BYWrbA9WpgVsWDN1nyCKmnc8qirg+ob//EA59Sgh/3FYxn02LnWJZlSMg37S2RFWFNQ13u1m
Dccrr7VhddWyHSaMYAU6j0ya92hNcMNNlTryMiXxD/N8MbJ0cdSkjvYGRqVdWqExS6zYdt9Exvy7
pIjWrdkaTk3QkwnZSCYdJb3SUNlQozMzEiBaQeGFXW5aXiyKNmFBefhxzmU6uoAqEUaF6V4oDaof
mG06HnW16G1lR2xXq3hJ5xMUhxStAgKWFOiIo9oGCUirAUvJiR/fg87VhZHLb/iQHBzbzg9G/yxs
+elgAc8Lv8BlLnGmgp4FTgzRkMHU5rvsVk4Z8ZzjkXbvdVJtGzMSJJ4DSewqFjtJGdCwJAGPAplf
B5/H9rb/uo/wr5ItiC5y9iHU/jc3lBNgcyg5WYG2u//z23+9U+RCZqXpQS3yV0sHtucjClZKHoz7
if058XErlbkkoGTTvnU6n8tX/jF5ZXt+yywETS3IIvrbWXCmfgnKWrXgBFaiWsFncSMUmE8xD2dE
LcACkKlB3kqotxxOE2hTnHbA6tIJa62KlWtgu8GdQhersh9W1h4+Qvzk4OaZnAQank5+5s4VQyE8
HCAkKWk9aqD90vj/etgW2Vfl3tqcSP/Ft/2yrjbvMc6xla2nBvNuKYYrqHkBJAUvedDCbOF9grBm
VFFNRW9V00mPQqr3frDjIds0DckcTZMDw2buhpYsXl1xlK4B+mqykHgdDMmZMLDtCyLgdHxwBLuY
TEf9mdxVqnHXDIuxIv6owBjN7qqzqKHCsnxEH5t39D619fVsH5t61y9MJYe1DkRdLSLhywf9HGPO
VDwafc/b89gFznEKitf4QTvKoUftujLlY9fKKnjWgodRyXuoJp4xLEPahgM6YX+OacZDVRry+Viu
280IGL2BTa2Aed9aVkFATyTVJ51PGSltAmLhKJyqzFRYctEJweuVoi7eCOk9Q6x/uLhiaYqIaPPV
njw0QnQ4RBscAql+SyZ8L9zM3lgV49812cgTZblYZq4DGL4b4c9zJ6xCiQt8trN8+LcWAu1AoOvW
lJeBKYjXkuHTsw3fVBhdvEZHQavzm9c+UgmTIU/Q3aIRFDoRiFoZvY3My5dRH1ApquF+4jrpiaz/
EWdxo6cau/2/dB4Z9s4f0Gr8VB3JmMpa+hvFJ8AbH30PGEB0KOcgeg2aDalMzNgMqrBBP99GqtJ+
O38oRbjUDCDLWWk6/KBDOepwKTkQmXTtnbWNEavvPh79xblxTUnWtAs2r11ry1+oPiX13kJRQhwZ
96ecCysGfmK9elnM2iTnF9Kez7oP4mFZRhZbUx/9Rd2piol2HT44VgKmXLEOAXQAR10Ll7xmS4bs
o32k3mgSJF6ixG6zBuoq4Ys/MtXM5OsMJsKd/4mdCOPR1k3N2pE3OjX2PPnpeGje7dgLAlw876Ci
Hukucm1OzjFypUfkGnajIjGsN3OCzumqYP8SVzeb9PixC4NjoqfH1U1g85wc5GJitKUrNF4CCo9l
1VD15n2TG9ff+hmxp2xmtGub61FAZmmtiCjcvsqpDYf4Gg2ugHnhyr8vZRKtzEK9gcSNo8J1UyIi
xBh1QnASPg2Wm0T85iEaoa5kaDtL+CRIS+5Qq+mXxZV1BoMEhQ6lyTZUXXJ3p2hGiOQ5//x7BSMu
fAUGCUqpdFfeMMyi/P1ajShPLpw1lby4UIIQUl1Q1aMYYK8lJUzi/J2AvQO9LFF7n0SHlf+6ihq0
hMHAgavTPI6Y3hON0JMx6RI+Wg+6LImnLWoA4uvWoqk1l2lJR645io+2e/5mrZnjfFJ24Jy3qe3u
T8oBE1ao+i7l5dILOpsNDRR+SIFH+qWvh3Db7sJLfAMr7oVyinf8rzkLBZURBgak6u35a7ss7RNW
Vegnm5eKJMTd0TOwDw1WRMRC27fDp5Pv59YQQpdfpSfV1QncQwSMRaKvv9OhN+UGgNu9wIcBUeEd
XHnnhCal34Pm3zLVYZM73miM689RoDX6nr4DNHfuxqcfuhWwnbfapjN+jv2iYcXk8dT05SHSV7Js
UKesf7VMuNM1iRdspqozT4DjXgbJ39G/Qht7Uupxo8pRPIWy8OqHAafkuUENLVayPul+U2HLXmPQ
4P9p3s7bwR59MrieIn+UACPOiCu8q3jlcpW/DdtysTj+imJrBRFu6c5KflaJq6RgxC0Vtp1/AB24
FzetD5RD4CVn2Fc2IloK4kgbi2IYBWyxQfVT68XGdGCdmmGBNZpAJ3qJIYS7QKJJOJh66dQHsyLe
nweiO5EfNevhCcGO8rsYzNz9PEKQvM9i+RzSLas80xLxx6NurTEx3nRIi6hVJylU2zoBP9wWnk+S
paN1K9urvYTQ+Egcl3ykWiMntIvbA5M1jKBy11d++G1I1Qmgz5Tga+y1sPxJ8sEIeOu+USDOkOCT
K6i5dfPt3pq9e/E1FXImMe3k9OIrSPRQZdAfcTFbJBmOq5agETBo6UEVi9hlRAuAn+f9dCuVOEvT
ujyaoYjLz/5lBVNM+Nt4CQDS9EMIYPX+iSaY9/3fx+MhDFOP8fqDy0LgfUpKIf9KNPLnfW7O4T7a
rgQx6QDgbWoJhqG0Awzij+bczOgZdGWbB87UsUIA4N4HjqWR7jPgH9uic7ImIAmUo5feYDkymKHk
jg/K76wajXEJ51j6CFPgRQ4VLExboazBzTeUNmkGst7R+YoYTAfpDi7/h+1E8GgI0k5UGUkZAwKC
3obD6ao7T/N/oEcSfrogdtaC7f9h3VFGygSx1JDK+c9NMgfh23by1EAv/rGO6y6NJO8Lg8aYdHzU
n44eZxTHK9YSo4VZEjFdeerlE6Ke8awDCPr0RcNq2M2zVKzkHQiyLzhpxcK6Tn+VwbEmGwPi+8+m
NwcxIu29MZRONoRUfZhUsDEXK+p4Roxys3+P7f+Xo7ZDxknDakCpDrF5PqSjniv6b0GIvYDyGKXv
g+6YGq+XqWJeC2DDkFEQkZ5+su4OLcdBoZ8AgPiufPmRkGq/9Ef77cZZ+DaIGtD1K3HWi7pXLt2f
nTzrZ+N35tHLvArwQTSN6pxNVvoY58Gtm+EI3R/V27zZ20f8obDiFSXQNLof4uwKDbLbfvNgf+0b
LaAUZx6QAwoFbHgBzkaISDKYAd10/4Vvx8m9FCcdciAI8kzV2i7caZb80L/CqHtgVKw6kQ9ith17
Oa4md7ImocpIT6PLRcYYP+jrznSm52Qr1zZ709ygvHUqfDFQjWLScZbPNlFYy4J2G2B1Ytjyc3Qk
5C5wyOw3TWjS0Ze+Tjl2msQa168XyConIVPjch65k3F/31cADBATlOIOCCA4PEqRvM0vPUyEM5/G
9Mk62Mxj/0Xod8lh5JqM3LJ2Nw6X/vViH3T9eImkRoI0zRU92F9il6Pk7orZJIT6EnwJiJaYW0eP
dXyuZ8TIcK+a0Cf//GfEL1olCZ1SIxdw/C2LGoikhed3GSPV4h1sJn4a49HJ9G6yQ3bgJcS0FD4I
VUnac2V/k3BbhNPNVLxlSavLbEUTuxULV80SHY8IX70fa+ifwgDiOTMcidQVpNMoEzBxiW3cKEWv
zCCXbXwGT9MisNKOFCxDboJI8nial8kEv3jIRKUYmf+qYymI2FID6t/1Wn/ApiT/lQlUaY+ZBzxf
k70SE6FgbG3/kZP4XI0Yy55Ob3YNOxrTADSb4xMVlgr4coXLSp81t2BlrKLgbp63XS71E/W492W6
6R1YscsDcW+h1WQ+LSlXxMmIWQgq/JMf6Xip+15b8dNmzwWr07Q6lGiyhm1MpDxWTggRM3rcROn2
9f8+qNagruXPNFZ54RXkiNGERCw2ENMsGFSQt25FHWsOp/03SIqeEJMSBcxnuEM6VpvhP0qDMvKz
ObLtCZ3NG8jzStjVig6gP0iX4//1C4vL4ZoJgXB1AMBIzvAak5gVWKT3+95qeWlG5QkpNkimcxiw
RZeQEFwQ44vgPI2+ZvKLBVLqrsxM3FHZa/qgNNUWH2x5gH2I7OndsJgV/9NADDIrMq6lb8jQzlnf
DeBH8b12N1TqH6QBLphJsgYWEGdScrDrdYMpEAQx2nh74Nn0jiwxWhqmDCfoMGURfyMbW1Z0Rr7a
y4kYwIQFp4bw6EHVb7BW8LLMXLobkASfiKk49A2lGeS8GKvLe/rJ8W7sN6NucpgZhUyOp6170dNM
PFhx81QDKqYFD+03RUbwMdoqE5q3R+Z2YM6Bi+goq/N1Ts4y93iQN3cPPfCcRy/DriLjuM3bmmP/
Mx/LvJ6EAY2a0kcJjAFcbxZxt7vi6wzt0uvHuDgQbeE/YaxbagXUeyT+CGg6+BjakUdBLLV6i3qA
RJJQXgR1v66t4I7UblqSK8X0dn45DDn6xs4kCNN7lIrN055m5NyrBTiWW50tPCJbGcZqIAfk4rK4
04dvnZe03zUb1I8SZxmaWoxrW6x84rgU3c7xF+IfsBaTK5uF3yPRhf+4kgfTRyGo57Sifv6Z5eUc
ytsJXqntLafb7fLw4pLGSt6mLvwa7LcJwT8EPTPNh5LEIEFkigwNWUkwjdw8IJjunEnTIIO9rF29
9rA+47SgHw3sw6NJYSUozQqWiDqrxB4r0BdaCRWZkNf+yARqsBivaQRQKlC1hB99i99A6ZZzp2p+
wsnHCYohjbkcyXnuT4j6CTU7tlr+PMPg06ajWZVrb5s2/KUKPUsw6pxl0KDZNgNfFGCYS1dO3eFU
9FalE+dzpGXyu7MCxbTR8abyMurVKWv08TlDmejyWbvlpY7vwCtIHh/o3OWlxhhr9fnttwM7fYTq
MriEjDFDj2PdAwFqNKvY1CwEAW8k277K6+G7kBEf9Z1gpv0r8Ht+TgsISYuOBZ60cOuNjG1H6TTY
NM6WBcsFeP57J9AxhgpDNP5+dIzLSl5mXPfVIzUd6NuRfM3xU0YLqiHr/jqtje0D1Bfb9qsy8dDf
71j0nngPUexFIXGaqL7frbWNq4hDYhRiG0KvaZ8Ja6pWEpcKwuMT5NEIDdkLgl+M46qqoFRqFNLT
fWUXjxSfLvvPEy+gFvyl9VzNvmDfcZO+r55WdDUmJFWR/AkmWIZ1ex9aH63NQBkPNlnP+ApOILyH
ZlC4rK4Qayga7hUqGGMEJj4rcNq0K6D8UkcOkI2sh6qQaOPCi1/19VV5tZpsBQDA2uxzMUzgdAFL
ODb/aN89gkC/hRuWZEPo2s3n2X1OiTar/fiBoSOvL3LA5fNBrQ3hRAkPFQ3apEex793t5qugVR1h
gBhBG1Wh5HM6oHZJvCOEUdk+ERvVtw3CkjGz+KIJAJOC23uUsOogZmEhu/qB7Ny3Xlr/wPsIm1nF
ojk0GB4IE98zOTKUM0plC/kWrDCbUlDezVqI5obIeDNg8qzqLWjZhpqGYdpamii6B+USXNKB1YK6
mJOjyKEsWqzeL3q36xeiSut3dQtLeMhfurejeppD6dX5/YGFVCwI6tFUvULFpYnm0a6uoHQZOYm6
nhLV86o1rZuvPjvOwFF5QhorJeZ+/rUmlFWzURiffTzOZcTB4aW1AHW1io2gFPHN3b0KaN1i3mZY
RxbSq7mZM1lQPG6KQ83L0U/hxjbbmb6X2uAQ6tltBAmndSrWTq2MQq0HnQ1QmdDMtcIyKZCrVrHM
6oozsiwMTVXWC+xf2hcD6QVSeC6HzQVGX+mAlWfKAccDM7FCdNaOgfpGEnvgbD1bhslc2WWB1oxh
NbteHy4izMveFvVEHdtjgHaU/Nag7IsySTlSmRjEq6BpoVLDADGVYG4An63cVNWplrjQ1svbl3Lw
j+Hj3w/Ig0M6Zua/nqL8Dowf1AMcy1wyobSH8v06NSnDdWXqTK74Vl7JUmRXYl1mbGoxcuzO78IX
8EvQ3/QsKI8QzpTU7Cp94/ztsviRp4bLrvdWT6PU/kzmJxw1AcYQzk+pYNrfc0Z1MnuVXoOZUe37
kMoWksuEmaSsO0asj3c/t6bB9BMhaWVKQgIwUVJu9zYFFAhElgUri7ZRdJ+4wcJm7htrlJp9i18T
Khl0M9uFNZBl/Sb0amWBwt7KpiCC9xHcMxAmnuUGFTLR1Qiz3N22dMp6lLYTbx4hKOpGjF9L/3SM
/LWd+f2e3j41V5HUMMwY0EcOz9Kp1LvbwkQc/2YppA6VRNoasHhMlHBkZWyG/Zj9pMq/ZxRGtjX3
G5mVWVHNO6AQFcExgCEUFpmahSoXy/6qNW/8nnoZ2tJK/elouV7C0XQ+n6dow8/M/TjqcKx2+rd3
eL7QN8PX+AOKPwENslgZ7A7o1iu0zTA1Tydb0wGm671gRzilDgsHXrBaK5Kc58ih72cuXz4nCJNC
0n3FktL/5lFoQc6LdaAmplv/WB4dUtZmRsiSXpWbXRNbLizqb51Lioz+jEVJebEppQNOeMZn6Nxf
iCyDV6F+K4SLKFRKz0+I1QKiv+1VqZWUEgJieLBYCmow8vrKMUssiYhd0gJeHRP/bKxqiyZ7cnuJ
2QDSwzQA0Z/N/85KWTiRGOWUDH12sb7ARg8dYZp9eD++X1tmep7vFLSaeY00mutXkRPpIvYOBjNB
+m3nZ5zINttb/nidzxEtZJQLYo7mpWIQ/4O7mVb9aIBqc+cqx6bMixixt32O+bRItei2QiYCz5Aq
gm/M0YccvXMDGXrc7Tt3MV6yG8w3YcWUMoxW4ZsDQlpVJIxgvHpUrAxuba3zy79YTb6ZF/AY5JNn
/6Ecps4KB/Sq8tUEGKaKxKnw2eeASijj0kPfNnpLC4jlePpLu1Piyt7Q/Fb8G/Sv/52RyJOllSqM
rJoJ7BpzFNhSbPM+7pYAF26go0Eh+8FVshMJFaZh+pnSUGs4E3llb7MgiTW3RMQeuBlCiOrpDAZi
NSfeBaBZN/PSletGPtZ6yA5f1MP3Ci5pZWukaKjYDqBXmxrJu1zo2IXK+6DhePE/Wt2j6HtuniUL
qFJfY0l8l/zelqMDKfgMRSap0Due6RBKZYjiStWAR7dRaCbqTwYSEvYpat2Wr4qPm3cFHEUjMng4
ZcnbkfKKuHsOaUEGZul9xoBurOZf2zxVEH1+tfo/G4fnncPbVl4l+2HxjKOqA6ms4sTozHWX2k9z
MF+Fj7rE2Vg/OcEIPjN0Ir+r04IFFfJ8yn6Os9BNExiCBAfH9a1qnzHIeN1CHUL+5IoMHxRu5M6e
zUR3ti9ANzrOA4m/uveLWMXXteBYHiGZU1NbM5Pug0c72m7nwyIqaNk5WxzbTy3PW6EG0Gq9bZe8
dj3ZkERpG9JN4W7REoZfGRT6sqUWcvfOmcvL8pcmr8Pmrg2llSROxutsO2ar3LaEjc4mme2S4KbE
X+pTRfyriIuXXmvR4XedlEXWFA4Eze6R+ZYweE3QCTtXSYSnVyLlvTg60Nx+TDZg32dnPqiBmyKg
9NoM2vs9phmCRJf78bZ9WCv1Xo3HoZ9G40ksW+nzzVnlmGE45ztGpFPBTXzbfFk+uj7qoVGrz6Bn
qEi//ZuUZTt1VEG2wkdFuco7XbDrCIieu8qajWzC+xzJjrerEBWWs74AcH5nMsahwCKQs8+xDcOt
QfRdDSY8lIVKYCEAuD5C7MGYRQnWfMbyx8q91UqfqhdNslX3U2tQD11lYxcgDe2Uqk3XNOk6sGtm
uIbYz1/pUd+hK0yX4QErwWiD/v15jMpbNKOSPX0GJd8YAb/OjY/5yjq84epsDgkmpjoQXvGlhFWH
UuhcwO5lmoo2gwyDmyd32/pShXHYAC7JpgW2B0mAO/p5AqXUu1uCI665Uwkgm5ZPKbzwvxfZKqqo
6mlTKcwi+Fii60Ub6uJKNryh0zbwI8TsfcFSmNe4sCwRtlqzGZYNLS/i7yc4gA6gvtg1o8MXIxu1
iHIW3/c4Vsg0TgaKAW/gxB0NDGP3oEz1aN0DL/hqwFybt6NbEkpVykckOjPtf1fNXKdN651+hDK9
zso47IifgIdz1GQLu0CLqb1DQ/JwikkAxM0qvZQXD0dSbJbBZ8QAKHOqakdtmKxe/yg62UKE+pxL
R0PuHt2xU79GAqoRR4pDAxUaoadNYgM3lkafDS3JRy6lnxC0DUOFXQK/PGCSk3Zhmx+e4DtkbZkd
qm84goJgWN86RxuWI46JeCy+bteYS5XREPKNP2H41GMUOq5iOh4+zw5f+TTcDhDq2CiAWIbQ0CbR
RsVJF/xahpe8p4DXmr1xld3wlJl3PXvh+gIcKe8NTIzKOeQu6W+I6DJxcHNbDYUON7bChpbokBQ5
CdbmfknN/a/KhbHjQ0cOLaFUUY5jzSdsi7aNRqV76nKhBnI+fdSxxsMCC5rOYiz6cXacncGGnf2e
TQyWuzlK7guN56x9D8Q1n5EKpN99WN8HAPbajJf1yyMFldbAkQRNVbfOjnF2nbW1kte+px3Z54qc
O5Fs7SiM25Fk9/uoDQuDaENam7mjAf0tEat1T1uUbcvVvdOhASRW9e0Lm1sodae/P9trKkLZV4L8
nBQNqBgFQfyIasiiHuwRAd3JR/lDgVMIahE1v9zfNk/wPKThnIBlbwcxfTTy6GC/vhF2+jPvMdFw
vTaRC9DODYRb6BvgcsUWNGf7eLouFzU7b2yFEpZFqmxiW1R/UtDduhDmWEeKZsTSEf7SBCuik0m6
aHjUSTmLXLfXeCrREPTiLVJ9AeStf1jMJcZw6VH+Oa0VSzivElNt6atE8XoMHtqvGnfPkub7W/3m
pJvwcJNZInMsIpdpzfbKRbtkrcMQrXkXKIF8i23Ia9vXViQOxPhk5q3Uj0BLeirvEFDnAYMzYXyc
kE1cfvCnqKVUN8aN53IyWjMVHZJ4dBQWA/AqaD5Wz4aVWZOV4+ZORczDP9FZ8KeQAOh5Ub47Qz/G
Tx10NXvZ0bmCXRNM50R7EP7f8kRpZxGYnpvT/qBQTXThlN20Z+MLn2QvZTZ58u6f4M/jR69hlbLq
9StEg3yxY00pp9C7D3CQjDjY1K2Kpn2Xk96lGqeD2HYyH46sfMev6c/DmdW4DX4Cq9weSqaVnd3a
FvKEJIM/ILk1MKL/xlfDyN71aJO76OTDZ5ZXM6TsHlPDb0U/ZF4LsVNHEYxwDq4UYltf4hXSzwX7
V+H4Qit9Z6fzpHiSh+PPnwqGyXSFyoKzOEiESuYp3rLVBLf73Aw8hhylI3xo3V044DuQk9Dzyqwm
ZWUe3QmeVZD9sCB4vOuY8RF1xLWIXD/RkywBsrbL9VcZfiMMc6UUJLiaIzzfN2YYklFk3/mCf96v
QWOUEkS5u/BI3ZO5LW9y+l40otUc2JjguOd2tW9SHE9DcyXxbe2OSbyPuQ6YmIkshVO9W8+80zuN
Yeow2eim0q0FHPNC2cYjCK2NQkeX9jYi386eDPFjqF1CSUhzUm7P6pSMFNgDY14Kh9rsOLMP720S
seu7v8qWNWmMAJROFM/eY3KuJsR2eOB+9bOEBz6TD6i5/8b76BZw64WL3vXr2KOU1uihR1AFuCkZ
WzWgrKNfmkcd0lIPoE7Xbou+CUk4GAQdsCPg1VpJLj4mRNlVaVf1wDpKmxG0lmKLIoCu96U3V3it
lAMfVvV9WKiZf8I7xIXkM2euUkym2MkUt0+zVuuQB45P+i5ygbxQDOhsYGY92QbVG1UCqC/JUGoV
qUapmtyWzqwGAsoN6v/SHYm7JKtQIe/qdjv7VL04qvqqsAGmGy89XEE8VJBL6oIC3tKpEuETkSi2
vZ6u53Ke7ej4RbzdQWGJQfiW4KAigRv2u36+klIGOfLjOb5/hv+P0Y1tB74jyEngoR1z9KaJn/1J
pgORWt36hRBVsy9WG7BeoCz0s71z0T1OiZlOBnDTIWVGBmEYGDBz2nxl16njjeZTDU/mnofX2AwB
paTijhwvF7NQfDrL9HcPzGapihdfX44lxwyGrPwruCWJCVnKo5F6FoyMcw9ydjKzF+iPxXbnVDlc
OOr08Z9R1Ch3a8I7clniBFMtU/xIERm7SiGAC3Q+B1knQ+NauZlYj3B3Nrm0n5fPy+wGz2kEpzTS
YVoPioJwfU0hr26zvIUCL1GXTsObWWzylA0yMYiwJgNhc4X0cf37bUIOYegcZosBFd87qBrKmXRV
XCm6p3YsWqGn4kDW3ni2tbUlmyiHVScPU+Tfx3cAkuW8JKwQu+6Nkjlmv0Cwc2rXi6BitnxXeCAh
0xTrKeYh3fhTu/LCGp+xqdtRKNUX/TPjpJa49DwwH5PN4b6aDDAVjvxOLqO43XnaYjGSpIef1b5l
tAtgSkw0xJTFJTi21/FQ7Vx2h5j8/VS/qHhHB1eFQqiT6iFpyt5aqIPoI+IFbru1hb10L3hE4NCa
2Dx8kSDgUVEWtuQs3oS6I2eh9GvhWPzGQj2lM7TQAIRYwJRSjYMWUwACMgxOj++S5p1zF+gM8oGi
oYdAWSWRD/zLpiiCAwnRWSKNDicLkGxIT9ZVouZ2tluP/MrdF80zKZCpO0YQq1C06a6c2mO2O7ys
Z4diqZFogG5iY33HFuGyJ//jexgpxdiqoumW2jxX1vOGqEcJWaFVQPyMgLEWB5iEVQ4aqCt0zWFV
n9tEVmEZn3DCj+tRT2J2u17G5qv5gvK21ubAXgL5aQC3rBPLmPebMdXTzqTG9JZDRH5DzsC9Yj4a
mseCw52jU3FN3fzYgKqR9ZOJhU2Hp7XvEWQUwuOPYTk9bIaNs6LvzjAAn7mJeH3bdYC+h+R/Pidk
rhEvGvrMPexjvHOgdToYlvXGIoxjkYU2/AMQQeb2QoqqYQzgu1DZnP6pv5y0sPPjX1w7CpndDzxa
rCPFByg/ndcG3A3ezMnrFQh2ZMKreNrIlhA87a62a3oNNq1CfB0XiRqIA8jB58RDvH/KD5Dxqy9M
DMn51fzLw/hMkinnK3KJEYq0zmY/rZ8fX3ocPLoo1ezmDrJDH19YaV8TjNIrbgZqglheWbdKq7ya
xODOVeeZQvseztPI1XnC/0qCid1JBV3KfJrm4AwHi3W6OQfw/A0ZwPmow1K9hn3XWLUYrE/VcU4i
E+Rcr8e55QR3iDOcAOm0iP2JrfybvAv0tpwDyzf+4vbm6vNwOkFy4R7+JPKYvQvabAfFslFqJ1q5
iK7cnlTpBXeu9t3RfUhhy3hrEYepbFmVBbuCTK9/1pO5IjpPIACFU+7FnbN6jPyqZO5nLswelFcP
gxHTRSDoFh6zrWyFzQegED45DzRVvPSvRIWX954E3PghGkjpIGrFjSNpKa3Z7Sq4tSF8ERoAVx/9
OxO6HGxN4/SqxEcZ3ACgn2PrbNvRRqqtJD3GLu5HPun5tnfZ5hACqBV+45dTMjUdI3EBCQuBD3z1
J8H15iaVVZZIGX7DOt6Yu/kRUs5+XDtgti9rhJMGI/ombatHzu4AjMKQx6pfIAcB/b53tzOMal+r
vHLJr7NKnjNPyQJAAeqOQFB1zpPog8LiVX7K/gUD7+sjhH2EF14EHGLEatmmNc1agM5V+WNBtFQD
YWwYm6icKxS/Mb6lMbsrvPrh+T7UkUO6VfxWvUXqA7zT6gEg4l9lu46KVLfcEULqQpJrROQqPxi9
H7b8KEt2o5xAcODvsL+y7GUfesGKXmbR2jP97pikvfPjw5AjkYDktRpDiqYZZMxIIT9xPdlofU8Q
0LFHFz82LaR7JK4Kk5pAPXwwfl3fgT7XnJ2fY5+y3/C9B/EviGbHMxamVWhjcci/ucPRQZxNR7qf
lVvkb7eDjRX56hXLsN7XQT4T8ALwIbN5hEvGCSffms8cRAWs//YKO5KjnDfr1gRdMDIeEUlDlB78
+R1hdJd6tNiJOyXoi2DVpsMhfM+t6m/hUsGmdw/qg6OpNHzowV3nuHNN3kfdPkZ4TYgzVEH3C9vB
OYN4zphpXbFCFjOToshClrr9lSnzRVnr7fhVkIvwJfU0OrPTpBjnYJyux21VOAOc7f/PIKHWQhXH
YgN1CMAHu3VxlVcx6PgBRYIjNpEOzZVumKJH0GrjNgGRIlJee4WC5TDcynnYf6PzqQ290d2GWyak
9BFtoYt+phd+vbHLwc5e2dzqzWxVmQ82uHld+jfHNgSvENNGUsd7ej7YWLP3/1xXqaqp9hWh3142
CfuG3gfpVVrc37u6g6BwWL3U2vayKMNo9VJ5id3uzcJopuMtW7ojQdOYiTtGfp10SBsG8Bb6htxV
/pphOArO81p8qJ9oX8uNAS+yejHfJLmMBuvAbzr2+gouZfrC3hesouUuIXMX6tws1BuRFWwb99xV
xmYpcxDZWfV/0QIrXhRddMngu/P24txKiVf96vWJlKVvW2x2UecFh1dcQkZUybJeGARW1CvH13S3
Go6ss61vyq49vy+UHBEuxZKYWMCHW47N1AjBq6g4mr3+icNfX3MGBGhnUBfXlCy3dvVDJqPtCnlU
86XLLddTmSp/+Bg3Q9waLZCmIvcSCZIreAt2v1ccxY2jkHnn3Xrzh1PCUs4UPGgOcHYRNvvVODzD
lLxzYbGVCQLR3eOOOkGWZzSjFwPifu+XdHS0Y5sPt3jW2hbuJ9zpQX/1zp26dWHkI6c3PsfMHDRb
iuT+ki949kUui58gpeT+GptFlkx/1c9ogAwWSS3CNVx5F6t0D8UHyB8jH+aXFKG4zKd/JG6trXZ9
h+COQGr+M5iOipyIjaBzJMfOe+aRvE8T5aV8xW7yrz6OmE/T1hOflxvqT3qYUlMXEPrvfPOLa796
Nz3ReirUh2X3SurzX1tXpPJ2MQeKPq8ga1CN/FSwHGKF/fbBmY5lJpiziPtdaIJJ8EsDqQ4mAdk/
0uKz6XsEtnskDmQ/hfBEvUeKbJHbDVx1vmrRN8le1Vh3tmfigTr+GVwDUu/a/fM5tfF5rDigkWs1
l7hQRDyYIuFk3J48HQLrf7LuaFM/Cj/W/CVYiJ+xZpoxxmHpEiGfbGnj8rq5UHuozK8J0Z7xrm/S
Ii39f2kzoi4n0+cJmMqa8c6bFGnCag4XJ34s9PNDeHy0h454/kZmLIl/yXpi5QlSILT417TBfFZd
HOPZ9aIbcpFPr4g2lBmr8ZfN5iQaw+byG2fs0Y9TpHE7gE+VuwUL2QOfsis0nc7ByAWS/miBjo2T
kEHNX7QPsBLnWC92vF7gcUrz2mrMsyXYpA5nugq48LgPh7J3WcuLXl7xaRMrhfhJWQxiGAkaOB7Y
lXvek5C8mr45Yvyqp9uwLQp9FKsmX6TS6ps7ONrjfCRoAE33hihgoNog6vLgCSfJ44+uebVCf2iR
cQ/qh2XzFyFtw25tH6DqpO/H3r8zSn5n2xqh7qO/mHfWMTfRM0xA6T2e5oD8MpwCD7A5tIH6GFW5
3D2opdTfRZvc/z9wtJlvnZN3jJV9m44/5JY5Q4LxjTe4Yn+ldWTb+AdFua8lTr0wGzhcPPY+s334
8AlYkdHxkGas52q8TvTY4ebJpgSs5ujx+6BVH9mqxQI3SwYGaNcJ+LdD80+I+VikclDo0BJr5Xig
a0bjhd4HPXb38mhpYBKnpWs9oddRI8o0GbFmjG2SbFepNy3S+ueoNNZpLD0l8vtA2dIsiIKmqmue
f2Eza91AcRhLywz6RSqtfY5AP/JBc7Wz1D4299k7to05YWPfatycQFNHt40pWT3BhBMl5dIP5bTX
dmzXMkAvBMAS9TCTU3IDIL1ax6MyIJZIIbZTm1/lErpZBF2E/cvQGeCje8fX0KD6LzJSuGPeI9KI
XFB3zFqTUqf/0cMzglRDhiwyDT0th7mbnfnk4oKejETPjDJdmbO6xNzZw0lUUi8LxgTP1U2Lv0w9
1LGFnH6SHCtw+1veR79YBs6xziM/RLS4PQVWkyTP+gElcH27CLFEO4gQCtFD0ttwlAbhDCt2DCme
brwrksw3asIDhf+qm7qmD6O5y8tSeOiydQS+qFOVupXtfMqPn7iaitWu805AUwvikILTneDqn69y
i1taNK/inV6TfydfHfnQVa34fO1rIM9xz3T5EFqK+Wh9xBLO0xf8olAduYwq+sBknHFAqNGUerOz
jued735KfMP0tehLo0OoOCdSiT8lFwvUECGYbNrBxaRAHfwRATHEzSmGg7bj+tXX0x4OAZ3gkJsb
k3Fo2FEj2Eepy2xEKHV9s0wB3C5fU8xjPXpStEUxnnn1Grq3tHf0hoCHxDu1zQ0LmZ4VxDVI7Gp8
H7cmMhyageUPHgYAbGAclvoGDIf8r6IpMHSCBNDzklaS4e955jCeFMHdO2KGaHTFXURYgdsb4f11
VGoOcGRIdTD08VHuxYRzZl360lT2iJt9nxzfMIaXPj9SihW5I5aN6xwNmAOSEawkFZ0AxNwaqYKa
VT1kKoERxhOggRqFXQF2qB9qYxiGrRseT0a8PozLFo0J+EXPSDs0uS1mm2q+qPn9OnKW/YgWOEwc
CU/LITfOUAgbN78QaRH7F3GEFSNzSA5b9mIePioIb/j2GkYWMS7yBfE8gUvuslI8iHkCZJXCpjCT
SmPfMca8siWwJJqDueU87gG67oYnmpWpD0mZq4MvzjKxicNvY4N234pdVuts23RKLTMExyQX7G2n
+rw69yOy5hdz8xZQFA7KqDmeFHmpspOoDjG91P2t44bTNW+ahi3Ge0mVo9dRQp7EJm934WSchIL7
fpIzQgMwt8DLzl772lvYL7CV1MLMP7JXFOh+YeL1oKR5vtJAfA1+RDgdo/z99E3df2tZiNDG4p7o
rGh41dfFSy4ujjSjjHq0vtm78F0BWJPIU7bFGYoYhPqlyzqNpgmDk2+NJIzFwS+v+Aw778GWC0jc
cK45MgXy1zvXh78q1SPRSh2kfq/D6QsG9HxlfOduh7f4j8w5U9aP74KIO0jI41oZ37jx9ZDDgkvy
TSyaEfxrNexqsQe1cTnjiRac6glhbTJKZwcibEY98fvVjf4tmmYO/3ikCk3MRmNAJ7yT4ju82Ja3
KmpFvm22Erwet7hF9Qq4BI3PcCJKW2BxGBpr/67ydkuMvaa0boC6mHzGQK1AyeigT+fx4viMH4e2
eyk20lE/pyA8s05mlujcrvSSkK+7j4J1Ci/Qgq9w5uZK9tcd8/Jg63vUQUdvYa4sg4UdUOVwxYU3
x+PkHGoudOJhr1rooJ2GqfA6r6sB339qcUha20786Bj5ofxjJshsJv12iAVfq6NwsWFM8KDHqGHK
JpCXG8leOL7hxPQCiNaca1i35RP0+D83h2Pi/pujG1XNuuueH0B5aoNqoWOTYVARfh3+tBHJw9QG
IZo3959QY+hQm+Pzppb3w8yVI8CBw6bDCEMC0PiWrKdRRiyvO0cHp0DgsLUyx1PqIO7ftWG5vQMh
K2v8H7z+tnePQuK9VaSi4yFFFS4h9/SdBdKcUqjurWL8XInUSCyFTiA9QIPmrSWYrqcdIhE62dpv
RCv8SXV91iDd3VxYxE4mSwzZfDc/f3TnQjwP+UaT01CJ0r7QelIZghAABlKUTOri2rOX+LJgmaxO
GU1iPp4Djmh52tE35DuG6Z5pqCF2NLohv8AW74EfM5Q8PDku5lgvh3FJXKpUZHhOwHqVFEvS9I0U
5lMB19ueZgzE3kc17/xeDKm254croX/5EzJ44/egpMvoIgaSCasXPf7mCxVrAKQNy9Gs8C6QYECg
4+CugsU3GEL7MROgejVIjA86WMUeUdiqfkZlwAIT3lxyRqTD/S7QBWUmALZIxrGRAmfNFYzdkHvO
L/N2nu9bqg6213XO5lWEfWI9h/hA0BvjqaI+/yJnO2sCItBPdJR0A9HeKcwll90sFC8+o/MlNpQG
RUeAQjvI5MAeOxjIllKxZyVNngdIW9n5w5KmXogxpxoxqoO1XKDaTHD7dSDQuYQnYracZ3QeXLYa
Jsz4Bqb9dMg6bpy84cWUY0XwTKSL5W0Z8HDrMzVFqzileV6mHu6lGIAAv6j5kn7pVnfBBDmniIyX
dacPl9MCQ3/hEr/+nJQH7G7RqVJGkHetJbaNkNahTsTlwzuezQ0tZNHmVENLfsnvefBX/SYO5jpg
wZnBQ6fYJ+b8K4/sTuIUoFsY1FcB+FWUIeV/O7XnUJUlzpmSW5yTcqjga1fKqAN77zNT5D+s8wkS
Pa+GDjSf/Tn1PIiNlTPWw24wNUOJF6cpX72BFpdw5YRQ8JmxUMUXLgivRY4D9lF309ienpzXCzid
vhV1U7NteTn0ZxvhkOf/0NgVSBTxajt2jcxCuC0rhmkz4C4jbfqD8NgAXG7Yc4MHXum/a2O88jcj
TwTuFkWIEA7Nn2phw3A21tAJrTSXM2eD6lHacIRfV13EuE7Bv2kEs5ywihNw9uOi9tiyW79KGDcc
e7xP18lHRZaPiarqmmAQQDla6h0HvJ+NpVIrhBoxbDXG9JCRYJ69aX1Se93TLnXy8PSY9cFa9GAh
pI21ce6VSbn4Oq1391QpMvVDGsUATXX9QUceK4vHG50LAhrUIgqO5fd7+pyJKFeTJojQRLwoZusM
ZiaX9O4zHCfal3GoaRJNRuP5WcEdxqPh/ihNMPYRALXE0FpJ3LP7+0MaIhLqg52Kp+LC9SUmCuba
pKapTp4ISqwnzm4eztKTnpoL6EvXNPMKTDR0MXyA0DP+H4dmKJXIXahSLomWPKyMemcYO7kZ6UFs
qxCu4+/GWW0MtmVDI9R8xgDHr7fq6KFINnZzS0f2WLNdq4rRtb8/Pnib0HPUkAWoE8M4daBj/W0E
euc0G4iVdD9QTHtkV4QUADJwNUwvexbd9WV1AN7gANZiO6+sPrDvHUmwWAk+DIV89uHYGE1l383E
rQ9AFLi14XnOX6cQCCz6TciKdvESiwecGrI2Avv8Rejw25TCmK0f1iC8djs4kR0mWcebrsxhzVeG
C6xVoXkft3XoYjJJQ0u7XyCaUAdfjqjj8CO6dAG+AQDs2G7mpb+6LhNOAz3KI3/3gcg/ooqlBt8B
crzUXb++rCu74AS6PoDvxZFPOegFV49suixx2PiODTS1BjhrO7Iuctntid117P0SjnKKuFBjJKDv
chV3Cur+tk8pZ4pY0g/3RwjoVzlo+o8dU9qGKZWrcRjpWdM/hIZGutkn1Ghod2jEETKHCi8YHdsg
h+NLj3NrlgvtoUtIu9Dq1w9vSd5n48LBYLOXw9ELYZ2Nyd1jZIzAxA0N3ynF77dX/zIkwW+OOoyL
L6euf7zFewWWf+KHkgpJDgBCcbMN26nHg8HkIjIbztmvxEZKpTZ/Wikvll9ntvnB5aqeAtVKZUhs
BbRCbzuIsRnUv80pg9c2wCrfjEXa+aTUr0v8oe0eBCG217JrRF5WQAmJruOhaRMrgZ5Bl/OD+Hrx
IVkw8LODj5NXSMZzqXcIF72atXUdToPrFHJdps5Q3OB3+GA7drYEYT2+Bf6WFQ5eGqlxFs8cMKQ6
yD59/RRhZBJlNcYnGn0s/dr/Vhyhd+gCiiX7J5VXpkvRFSiP+O9wkoSHPAGPjZ3+rjxcUfpWRmBG
WruWchyuBuARNLlgEZiqQQjWBPjSSE+o+WreVLrE9Gvv2lt1jeO8EEJ4T7ts5KZpdqS38cQtGTqN
2WBnl+CNH5wpBE/I4meqzfhrgWXV6q4YqFSnxfZKKhDACBXqYIYbnhXs+5CkdRx4n8VhmWXSJAB0
gTNscYi6K/C8y6RcxoVC9X2/85GvrdtzIJMhcgChFb0QQdHs3FvpHPqw1dQcHupuNagX89RKJhF+
H8+6YwasHUzBwZ6RqXTigujFmF08gro7ynrIbBNB9q+vd+G98n+CFXIyV1Eg7HP63dQIBxqqUKNp
MUjubOaKAncfvEzbwn8fXV3Uoa4oJTelhfgpegLyuiWBuYCD5Sy1E/n+GptEwHw2ojkN8Q6FPJ9h
wdnyOw7W9HESjyMVSvB+AMl8FSKuyf4e7KVpFgJac2Km+NtjwLbrXZVx0LZ4v3eY4N/m/q5zpUkP
dQxsEEGqIr1G2y4CWOmjeKDwR5xO5lBlcZ0xme1/tjYdv5CGXypWBeLUxUlLc6bOHJ+jA/DRP1kD
yOrtWPgtUULjCKnmxZKSM2mJFtcpqQQEDLbOW/EUU+YCD/jSLNzdxKV/KesBYbMgZ4584us5lw58
4YVPgiuDWbhWn1zLdb1ZQ2P7d5OIJx2ps/0JoMduugLNGglhr6u79R2y6gvJ8AR6shMxdhuqJTq9
zYsGoGEn5TA6bKa85nhmY0enk+WG9OABgsIMmkC+nsAR3mDixYuP+xYWt9D3yutO9UijUidCoZM7
SULOBsv8q1JWj0pJDXCKaJiU51ZRbsVFPlbM1Yku5GFEyAvFYO/VC7t8V0baaHC3ttfkcnevGszq
l0ProHaIeldXSXecIRNL1AuH1lPa+FOSgiYHvzsODjDo/Dy2JdsYdg7oTYjbwJLUT09gLXlAzPvk
rn0reWvNenQ2Tl5HdGYevjmMIzb15xisv/ax+Gtls/oaFi3nkONbgEw4+hPz1h2lTDlsIo24j47s
sni2d3c/xyv6fEqRs/FfHHlOwxTBenIWPnp8rBSMMpo8yVgOO/tW+zuyk6N0uLNvWwQzBChwF+os
XNkeNMkeRFJL0u2i+IRStnFuN0icam5PvdSlcKcwLNwNO6RTqHpn5NGOww7WRCS9U5X0TpzN0Pzv
3ce65rPhozkFlOXORwjm7Xo2UpOLzpE8z9W8lirYifpCF5zKX6rhDRzyHqi92CE/QXloXuyploRr
LsprIz3/bzvvMily9sM983pTSAW3u8GlBlnhNKonQYnK97sk9297lLVh+CnZQoF/IgrZz/3IUsMi
fvdlyNNjbeloD6UGFuVNbOrqpm748wtq/7+06d4G2wyQEBNkRoCFy0/yJu1HT8NBqSzFeCI1dm9B
NwHUnUAlwxuQj33o9+16Rza9rIDhaKtuBrjFjyfZrVrEOpZ6kNORnsb5MXsyLx0SxQ4XmTLmH3KN
zzybISCVDrOFClm0jcoBwn5TAvf9jWAUE2GhAxw3c9N9C6myl2ZCSOGJHJpKu1fzSN5cv+zDbziD
sO0LYxrNHKhQylzwLuK7saaNuidZNr5yhSJgsb6g9kRuICefldJOES/EvV7k/joJnBf0jRX4yMZz
8K2N5V+R6XPKHDNzs0yvt1ukgXuehMcIpxTg7cPCoayFa3bRPMDcY1zBEJrC9SlReiElkve2bg3O
QE5Xr8dnMd8MCFf+cQ2hl+cSNt1yGYNWFwIw8DfpkTzE4XAlkdu1PMjOTEpAICtS8RifKivLjRUr
lYJryPse7yqIXH9lAkDGq04e/2UcZXsduuI+yIdrdaKYN+NI9soI/uQ7w79WZ4gKERSJk/+qPd2J
MFCWLLjX+2fNYQH1Dcr5TC26lSHTTL+3sUJI2cJm1f7LAZNTjTpWl6DH4/ocoG7YrjhsvMH7gmFq
DHlGMaXsKgybfN33LTWwAfgKrNlwCyi/b9Y5XkYBm+c2xowiosNb7LEH49Vtyc/5eB+XRqOxmq7r
pv5bRXIWhC6DIr6DHytEnCvuhdA3b8nNkxzxHn/8cWzqTTA5Pbfp5KpAxrUbkhQzBUAePTdf0p8K
RIgKBygJ6htskAiRpLnPed9n8gJ4uDYfUjnkzicplGd9rThnyTRZGoeVSP6L8go/aJpl7QNVdhJb
x2q3zjoR42bnGZoJu1vpLI8GAFQ4wGRLqLhOFIg1frAxe4doLrzLWcX4cQ9FoawQDySlCqKaMK1p
ewTy+CnTehaDJ8CeWT+h7zYICgqJf+jLh6bZVs6o5MsIztKbBHUqeQ+FzTnlBfSgw+LDb+9bYGFR
JzUBIyEmHPuDkzcyf+UXit/mmibeERZcyIoufOGQZVvlCb7Q/+7BlAI9EOHCNjjF5LfSYz5rVylS
7pShptQTcV+IHqUL3+eE6AJsgP8RJNusUuJhtyi8LrXY/1W3A61zFSnlU43ImMfFWvJ+jEnQ9ceU
neB+nwghWk6V9g2/8UAEOESDCMzVVJO9bpdQAP28fzPhTU20b2hXAptXRqQD/tIKVVWnhGF6pzs5
rEvnj2vDFqZpHcwVTktXEgGKAtWQoe/oyEs6PnW37CeS2MHIIcSi0QQaTg87wn4s8Ht6+hssdjDx
IsVXYUvR829AXKpqbkUkffKhIVF7IrBcLxmguSoJMKYC4p3ZCNrYFwlYQg2ezjWs7MtKyeJMQ+an
AWZ8kxHsGxJAkSCHbsuUpJeg9gq2XdEpDuAuzlF9VjNSL5wEuKUq7W3zS4skxiK6fXc6wuUq3X19
kVzWObRI/gQGqH5/aPcrDLtYhZruf/FNWGSI8isE8vXSOBN7GTc+i3cL3MtdzpqrUVKHgtvmAM46
cua2cixKcEaMLDrUKGf5prcD6XROd13ex0buSSqBt0qPvRMBawl2I24T8qVTT2UtJrA242S4zX9G
Y30fpksgIZhFH1kjgeDlLnCkHrYvXU89mRussR7GS5k0/A6IUc7H5S3QdUH+YHDxSgCv8eFSdh4E
wr88+dw1U6Sn3qczzVqKIqMuhzomKM4PRNXN31KwKBAgbSLUf5Zf3//AoCo/lQLni6xT/yGQ8kn1
RmKDqBfEUVGlgyRu4VfBGdDotWr49PgoXHwg9dRHX2gBBIlwiNV6oDNHi1BMAlQrMsGx5WAAIUBD
WClM6yIcMqNrePSxgyX45RwN5nCbeqozL0xfXbXjELiSCpa9suSljx7yeqgZ7hU8mVGKzKwPollL
JtkBgcLeHquEILvVAcJEXcNNUGsDw7zX29OBPlpuFZ1RvGRf5N2jyOX90lkiI3fxvZU4ywJ7NJJy
32ey6W88SAJ/UviwFqWBikGFskzpew1bC9XNMIFxSF/7nNsnQJRJbGV3QhCo+6DRylhMCLU9lnsv
Ia2ESnVqz+P0ATpDk/OW7+cHBhMoxXnJ5Jjqe/bD49Ytlz9Vw1nK5kYbHLDKVLKc4UOXC4wB+m73
jNZcnynVwiWxLUYfCjP4Be1Az6ke1i9JnCfYxPga2394YscG6lpVZ+XcvyVxh76NkMM9fwEcngEc
I/Ai9xd4mViBCnL89G9UpE4511sc4D3qT9oUcdXAbu3QVpTQbLHy1IFXCkIvmo0eXhimu8cDbw28
gktJIN7WlgZtOOzxFOJ0sxqsGWJKZUpyz/jFOeshmELy2JcQWew8B0aKX3mrj6cTLIWw2r8zf3S1
1Gxgw2avNnBk4SjU470ZaXH6lDJvSqbUo/2AiGEYcgT5uImS9qisCrsGXvnMbj4wG9P6l4igUQGD
QW3vThR8PS4Uyk2w9fPAyjtGj0Pw8mxN3/oaOtTI9R6hy9huRegfRFscP1CKgY2T+VYjSb+S4pCg
uGlTGAbGSz00mh0gVD7Jyl7XqLQfBtRw/eV2aAIS/qBl+YrEbPisOMFVRieArjP5rG/CjJHwSZxU
VmTjxegUUofJAfPyuJSXRFcuc7/QwzPlDzrn7RBWjGi1RB2MbPr9rrdm1GpDmYyQqZzqH682ALAA
p4NDPp2d3iFQl8MfizLv6jJdAnd/HlyqcnV/fgpz5bGnTNX4sT68Y4jsGnUwIKRykpSuPIfzgSPt
wGk94unRHoyUsUI6j/jHBOPWBCqI3962MT1G9glwpW2/+n7enFz0ENV9y64v3TZrg/Vcj7M/YrI2
jbOJ1SEyusnFSakqnqVsW64iY/OnAr31pboTg3n/7X9JD39E+366VORXaZtb9y47KX168pthV0fG
eIxj6pRHGnRTSmOIuRs6X2uOalV12aRusBlrulJ+M7lTus5mXct6Y16YdSUSWZoogmulSbAC1S31
I5i7CV0o5on303GT99qbQ1Iy73We3JJ+OSHjAEG9/AjVzyaVOdxND5nwKt5GlSfa9bIpz6UTKQXJ
9PXOlqIHgrVIrwng+L+COJWGAGPORHyeUxAx3zsLIiz4HNI6ndw+Rmf7JhtrkY6cbZ6WaaP7Llt4
ujqUxu8MLY7jSbkDI+Sugdc8QVpoDYAzaRL9+JLqWlKn7jNJpz+YAGCf7pHcatcLyxMPLeYMAtCC
Ff9mFFgsMm8jTtad6MEwwsSdoO9MCoPxd/+Up+cbKpV9i+/z+BeLMj5R1idtuctalAbYic630w05
kwKx4Cf4t7wcNSgEuH946+5ZkXafaR6PgqJCjd+8UDXeljY9lLI8xeHboPKRtJGu3tXs+1OkIgg4
U8ewsecOzoACNUbFK4qCP81uI5ks6kxyq19M7HZdSdrHndzTfMOZaWRNit5E8NG/DMq6RsNo7ZoH
Y70zimyhI8/Yuyz/Y143OiyNZvLzNs6GAQBQtyer2gMW6UB+WYBOjdFIN7MrROTtp3Z8krRRQ8Pj
0pUCXpDb427DZLrUnea/QVHCC7JeMR76NmpbtvUIAsPQD0PSgq1uLJVnbjptaBfm0BC7CRLUG+wI
Nml8ruTMuEfz3chHFakovpmgSuNC8Gzx0drIho4tb+PtZE+o9ZSdebuMZ2cynpU5oqqf5Z3i4HxP
qiPOAV6UjJ1gAnikt4F7Sqzw8bngO71zke9DPoyq7zKEZN4w8eMFG+T2XUFvB2bMepSnRSZVICoH
oTm4D5NVyhImBEvQkJZeFr/g+yRe8JypXZBANlKBZlXZ2dZD/1cAUF016ByHTUxDzbqnDOQDDnpT
yP0qSZm4oQG6jIdzTP6so6aSL23RWqZ2NsNwL203C6S9xnlpU7xTzFmyc6nQB8TiA16Q5aTzkBaG
mJDJl7va/EyqLyNBzWkEXp6V9y7oROi7Cig10EHVNJNE9oH9tMJi7pBAWcI6dd2HV1GXn1G7yiMk
xg8kIjOoMDyVr+rp1YdSB1mtsnz3RlMVVXEl+oT+tYsgeYv4tak/bkubB5h8Rv+zGcMv2UajYhwk
4vH+wg6nyeRKiUReeHU/V1Zyqr7QyEyYM3zoQPopzVVB7PGL0z1+1KBKNxj8cDFOS4jDAZN0r9xF
Dae/5lX5n1KG7KnXIM9sU5h+EmKUt67kGxAJwchXRn1MQHtwcefzayYPOQ3UU2uh/wekn9Jt6tSm
pWfpcy9DTg1txWZRXYc48l+l8gn74kvlTvrNChKyE4M/5MOcT0FCX0D1Rla0CbnzdHg6P83cLlGC
qtUEwKqSvz+WtsI2UzPY0L/vK1yNp3aWxGQFHPKn4/LviwZyaF7en4ggRpXsjF65oSi6/0OmLFmc
tanUETrUnyW5QubaE4VzaqkjOSZhtx7QAA+HxIXFOWZnsU8OjDJ28QvO/d7gi1bX52HejJueN4vf
2F7v/qhP2Emr/UfMzfZYsmU9n2jfPa9//Rt1dozWcJ3A5biLWjtTafayNVTi+Hg84Cv6QOl4uWq5
l2V2nGKUTRvMysoXohezuBPaMNq7IkBnnDXzWTQ+jh/cz1PbpqjnSAiEbL4X9bEXKbSaa3tLlfsd
+e3HCok16ksOGf7INkZ/g4NOfeSSGDDsYATKLRxLE7rpHvS4GVhbFbJcECKCDILTptfKk2//OS7N
J4GXwzAWGCzt+AF9MYMb3QngJUwPw/JuQIAHWpNHx8cn5iDoVCSHCTpY+tiuB/dKLORo1F6inD8M
pjRE1ZeLOj7v0qPE+8BoiJnpWZUTF571pSXF7tIvhIPfC82VNOlOcZZZSNqQKSpszlAwNjj40zB8
dxiUDw4U8vhJE+iqK1G+nI03FTrmkfHF+5ptB3kN4iFM6FPi8nOg+3GDS55DYXzHK0UrohOIT/RU
6J17N0+mHYmaWpxXWaTMhIAHmxP0tbNBtMGC4KrQ/bzQSIBMsHaSvOa0jxAKWMFTofscpAeythu3
fCS1kGoa4zWyfLuumJ12cri5LKuJG0FePh/EgzB/FdgQq6n70zmvuCdR+qEd7QS9ISaBjUzXfbCk
Qs5geY//2pEmexuCGj1SgUADx5NHMMGN5NfhhqCrDcGMYpwtQ+8foGLKr0a73pa6jvqSDsK36mYN
mYCJt+HM8CrKJTErLPjur/cx/VtiXmtEgf57fpxUbdrol+mHZXgvzAX6A1NxTeAPuX31d9zZ2LSo
lPgmkUF988UnXgxsocByJJzbK5bw+5YYKDkrvC9IXxrTrHlTUkJV3RGJMPKwQTpnSIO9OCznBC92
fl4/P+sMlw3JT9Yyd7D44Rc+jAR4CAnnLAH6KTVTDsiE7rLw9kUs4qCy3wwLBD6RCXwRwO1LZqbA
p01NMsauOQ8baKjSvf0y5GyC/OnAdv2wEj5b9DrBjPrSPCQJX4VJjzFk2FUjhDovuxJCYAfwJn7K
p6cQOyZcBg83J6+mkEK4h+ryU1NNmoYowdfULY1IzOQxXSWs7LvhZ3I7iaeFeKsc/GlP14WIWPqn
xo+Q3SgZX1QxBtK9ljeSOuh6DjWOHMZUJDHkgUAs973j+/MjMjQtZe6oxufkb0ufXUTybXLoHUMl
dQ+g19KxwfTOVmTVYGgDQi7iXcas58U1VnmuOa+bgZuyLPyRxcXP45ILdaI7G67AlyiQ1+e1eltI
TJNHCqj8JoOmJ1QQAQiFJK3rbPsrcHk6Loau1LVToVkcFUL3K34RND7frKBSjNcxxgK5DKZOTJSG
qhmq4vAT+q+5Jq/oGfBIOE9IOmiCrDXLpX3sjgYaqbEbGzICeZAAqwy5FHb55xCT48mbzA+izoCq
BeOJDX/oDJgXgdRtfWDC2Nv3coQNuVe4Bne/g64MPXXbjlvVqWUJ/+H6iztkJ/STp89PXFUA/Hv/
STJUR7d8GY2PhpuNctrwqkJBwMZWq+KKOid19FN/qBa3kVsvTSBmPIaE3mArhYckIrkIrV0F32uh
peM8pzijXxXskZGdf6oU5cQ7MIBrLoAwqTuix++WFDMYzCwWG1WEWwFWNL7osZ+v4tPixSxEVg4+
2cGXd8JTIe+1S3ql983lcrY7X6HFTeXyGOFcSOZ6Au1LednW+ZO1RXnudqanr2tJ+ID5XzEAl7DK
QlWlJZ6Baj4xgal/RLajk1yDF7123oSyhSRsoWig+NKY+UntFL1+m1wgDYRdYqSPRahAYBBTqV3b
xX6k3q3q2qoPe7zHH0NDIW5Z/sdWoob0Bpz+lzYhsR08RI9TAbl54Io8sv/01zXGmdwurPsTOltJ
hgaKBMA0BFwsIQkpKCJWztP7W57UBe6304GvulFdr5B0WhFCxjH3mWovjkcLIdNAGtnes7sDKYQ+
B5qyLSUFiVv7CmVjUI9oYGb8xMNf6JO/lLwIP/94SnqM7WKB7GRKThzJM4JMlLcFt3vdgCL9NjgD
82hUE22zH22Mo9/oSFVbRNMaaZSJgw9xeXClEVODSoAOe/yUZ8XFOPUs5ovNCo60OXUQHv2UuxgL
ibHVUg4FDj+uKbKN4evMaRee6eBKMgJCD+gHRNzNUTdpeFuq3S4p9cMLIJy6yPguHyyt3rL7fMtm
NM/t162ZJa/ryHzPWiiXJcvCrHYpXC8BhX/cRo/A1CWU27jlRayKMavuGBH/YAuZVXb4YMDO7oVM
R6SRHf6c4SxblhHc97zNYFUY9Lot0EwD/mXcwMnoRbsrhrHYxaqSrsup2Urr/qmyPdWFxMANIZSy
njzUM57cy5E7pwYqkPy1SyS3KoRO6fsYue7989iD0jmk6c0jBGpiGU2XaH5DAl5QiTjybhBEMQ7P
Limosz3lEA3Or0leR0maZTrtFwCS9gB5urbSn27c3J78zkIunWbYeubv3luI3lTB5EqFkiVUiN7D
sAr/LfwlpaU+/jWRVaYuhJQj30IGfwGqm8mVE+1tNrfyLqG8had81m7KOEcowVNlkzCJ9ECmEzZE
T8PursE1/RP78ic74q77kbnDsbxJY6eHBXsk22gZmoMsYyUQpz8moMvVy5cGTT6pafrK9ysmUJvo
ew7vpDslv0Hoggfwhcw6/jV4yN8TgsKsmE49aMRYxLEeR0BOjma6iHDqkYsfaOcXPprmoMsQfHZZ
Kq0RVocU5uAlDCILURgG50QzCYTWhO2WVCyvObNF8jRPV1njC7dvQKGXHEuzOFqhY3cbscUryJdU
dygsXNfMcqk8vSZslHQrA4yHriOsJhnYzQIrXNvJNbC11wwyaP25KYlkAT3Wu0hZsxeUZLOuBVbZ
ExQktzG7wDk/SvGha1qVbGUVkIGyqf9NQbIXUfw1mkE+2cS6VozNmK7qOz041gzwd0MJVx3Xi1pq
XXXv/pl25NdUbSC2fNXPludaeg55kYxZpXjdCUoPDgqdVVqu2kIUjn82B7NCCDjovldRaPtLArV5
KUJCqbNbG+5TH33W8W9CtrSxttygm8+WOpMMr3c58ad/AFEnY6hyHv8gBlXGgSlvISrkxhzBdFgS
1qERnsE+J4BzOWus4xnUmB56tyrpfRcPsRrMHe4Q6Cy05ZWHqkHzwIwjPPMKLAwlQWrbkOdAoKQm
tkloikf8zEqnMkugaJlhbc6eCNe8eKrkmkV70cWnHw1jevgfnp/xsj1HnGGninaZzxKg239QQAQM
qwPzJTt7BGxFRJjcYCpr+UvGSr8EgBP1bLb6YJI+T98b6DhMgDxwC2MkyfuhnxzaUq4zNEHKm3BB
DM3HWYagdWRhMxljVnwRyfOAw2mNAR5xuFvCNZNkLAgt9y6zE2gz0ZIKzFmPkJmw1jkgqrfEGli/
yGxUDiEj+m3r6GfdiEmR8LGS0HWP33XX99jHWGHTxlJEzRLJ5uIv+pz21uplKOzx2ndSboGGx9Ca
WoFk8lumId2Fv74vRe7k5X1PAuZohIw2bj2JF/WO9uJA3qasvC5cBiwPIL0sfn14cWIe7hkHMN3V
mSeclgwLFNSSFFf/oM+KGu6ImWJ9+tihPBUm47EzCxR+QJeXmQY50/PcOxJccLHiimndmQyYB+eu
Qwj3D5lVThw8acuWzyW2kbRw1aK5Wdz+fkdwEJKXHYTmJdVj0oVOMFQ7fuE3QBfbDGWJRnyQn0q3
YThlyuZQwqSLdDtk0WGhzOb3NFK0Mb57zZUiyBYNkhSb6I8kRyhM8nN0QbXLig+tk45H8TMFIRMt
JOTvvqMRE/x8ztojIQXZj8v6v4vV/U/sPNWOb7i2OXQ2C0pYy8E622LYobiKyTtQARbK8EzJupnh
1LkGl7LkNJusuSuTsM2vCEZwZNjCktOupm/S14jz/ba90067DQ0PpMX8XAzmbD3Norqo0P3bhB7I
2bwIlGYm+hhFb14Pls4hN25xYSxGy4cW0mOy/U8bQozxkVs+9R4u8YGkpECMimdgb7jR9lc3fAAl
fB3cZVwt9oo0kv8mDe4mMnvT01JOz8HFfqmMWmI5822NvRHZm7RqgtOChhxhgCDMbBRz5DUGnAQa
4LiBpFKR9gejuJ0PqC8wuxqh4WgMKR7Bs2yMVntVXyBaMEyi0roIkCiPwaV4dh5XXdHWlsV/XZ0s
8UP5sNSNIb++cKDt6FiHOaAm2IH1tGJFjO0B4fQs2B4aPPXLIU0GE3/dVIiBeeKFA7xkVmD/L3tm
7+YBCfh2WvkofmQYHLKavJKvQ8ngvTToZ0dlzneSUUbU0Q2kyA+DxKEwg3XAfQvHqJx6ZXy9AcuX
zkmEtcgsaovbDZoFlydqUEFJ4t58W8JuckbzSuHI83h9pHgs8d07LGQ/iChcLPHyAguX02GQuSzo
3XlZJZ2pAHplw1f7D1fmqSpCa6KhYlHt9tHEB5seYqwprgkMpPXJcOzEf1/hPo+KYhgYiKNWvFk4
rilzA9TAfHvNPLmigGzz/OQPrmhNA9X5ew2ma2mEQt8EQjlsLqXg1Pv6W0ZUQ6trzKzbx2VBECwY
+pRQd/TjCAE6TA1cD/pJcX/G++qq1wpOBJQpGvyHW5DiFWZNUBRzLdw4LPq2rrMzO4MPEQkfETtR
j0m+wBUMcYoThThFA53biddFmdxICZ5d+QRAXnaDxWN17wL8R0D8QSU1xkWOnQecyV2mXLJnGkKW
rQ+gbUCiIP/vpKf+I8OjnvrAywmZP+q/7mppD+s2D8Qtdfg+/GjQL5UDqgVeoMYK1VxoMasBhPrE
OXpFH/lQMCKCSa5AODc4TuS+g13yLMmHq8QKWyPeJta6s4bDrRMjS5IvjD7FnM78KiqqPfmSxvrS
SphnuqwxJSgVOdmmpZx32y6yRCjrnbsw9OdYF0dRO5S3IeJSTQaWD8mCsSKRoYBdcRdZ7nuEhB4a
+/DIE5gP+yox07BJIig2UrNa/W94TEBe8befhhuzw0gAkyGGjuNS2BXyQXPm2UmbXCMCVoQDiAyF
I4nSBbceNwfV6wARFH38V3cTLurrwnjdMhZdKhJKLAl74NTrldLOOqHkb80uUUBwq7Olbf2jhNSn
1gELAYwkrc9LqKU2HG94X5Y+KSA6+ASqlOphnik2DVj2iKr1DaMsmPcfWIqp99eubtohDQATQpcY
DoCMKQO/bCYa3UY4+pe7qpv/M/amrK2JkCs7tEokOnyZM0lEwdWPREevFppTPjBoLNPDsn0UpEoT
cDpzeiVdu050gABU3pwUztvNFdlfg5Knt40NGReqQryCCtq+C0QVZwNYI8KszyJbmHi+ZdTfVUhE
jioyDCVKyP6pdBQcJfi0qvh/49Bl+H2R0t9S7LCNzWvHS4etixd1aQ8kOPfI5W0m4ZN/Q6aLF7Vb
RiOFimJlr/wVmiEKubNggxan6wMiKDKJCgtjUBW6tg9nlMgqoPnEsxHA3iTt7CEGfcOCOYxFHqEd
KSnG+L1c8PDzwkub50VJF4gxdpPg8dn0eRq4GAPlSu72x9S0UH+PP67uQrJ3VDpkVb4x2U0c3oX5
mkXNj/05JShv4/6lUbiwHBWJzp0D6hNdrTsDDNUVWdxz+nZCgjjmzfrNNBKoAmDslDKS+Y1I87VU
o9zTacU3I+nLNqLjd/A9l2e0X9Ho1A4VwT6EsI8OzTnwEOsxL29kbRLV9ki5u2YmcMCyLw2GYAIL
Ymd4+Meot/SbKKBc71kpYZtfYIZdW6UZczWW0ss6JStpkx4rgwGBQYdruivWUI0E5Hp629AgLFns
zWvw0rHaMV+uV44CTUuN0cciCXzeiYVcIYSHHbhUvKB0H8b+wCpVxiPhBa+ZrnLO/BvhnjsWGX9l
zEaFq6iWLfbgg7/724RsC9ts3cA144cy4CshiwyVXfH+UT2o7OGD+bQ+RGsovWrvlPMFmy3+CkOX
gj5/DexIcJOIYbyPmHRZvz4h5ARyckv3P9pbQRSMJf/XzYYQNmS1Aay7kDyAWYFkxW32oHngpaJx
bCJquRoy/X+zUq0mMMOTK0bbAO93XiN2j/sLtQzFcygzjsxFj1v0jHqWO8DaVx3FXWCiRaLvFurF
witfOi2Mwb3bXOO2Voi0mQg91LZKYl9FPno4LNHplfbb/yL8bIOA7xoUyRmn+/sWTnY54HFd75u9
47VwC6R7fI2KKAhWvqaAdwUZsan0xKBaMAILEo91SS6wauA+Zkj95y62DDPDgAd+hc9H8chsJBbU
viUZu6X3lsQa2sMdh6yeNxB9B1ygM67NDQq8uKvtZ+tJLSxMvSSOSbyg58sW2N/mEPKQTWWfKeqU
TMys216VH0/oSNhxHl+3j4X79ZC1sN8vwxXKbCwBq+D/hdDQNw7PXjCALjxQkD3i0thAWb39+coU
BzG7gBtaHGzNi2W+Nfqh4/vW/yuO+Y7galX6CCbQGJYmyiiZZZ/hntjnh9dZD50PZeOWOo4wEusx
NdinCUz5y0Uql/pUAflj6/bCbhMbbpZbmfvQkYhOCNu+puS787Yq92LcFAqE0sGbIRmHgeOwvn+s
VL8W+b9j5CBEVZWFgiq8LB1okr2oJYHh4w7dYPgLbpqN10CM8Ki7b8EXV9qbx7yZIjA2OvgSL+MR
x+mJu1HyvHb9JHxgZz3D3JVjMzHpDypka+nRNRfp39G2Z2Ky1hnfwDPL3HSnFaqP3OB+WZwG5Ew8
6pPsAtbUNL2DPR/pdHSSObBnUVVFo8BsMp/DmS+ZevmTMP/OpojNrikgXigYxhWK/mXhhdzTYwDb
KTw/BXXxRtzlSfyk7h4y4LMpNUaPHb3VxQzZU2mM8Nj9DVK+0irxW/w1+DHsDc25zqGnZmHNfIFY
KcVWmA/d1eKa7GIrxA1BFIbwlvXJKEqvTyFCyqGsmi/mNx8UJXlXeirrVqaQvNQ7qBywPGgCuYK+
bcYumAgDw9mZMV8Un8gF8Eev8A4IQg5aGqcBFNqUBYxNegzhi6TCrg3tcEgaewOQa4isWkQ4YlVS
0K47n+ZsfkHTthIf+iB2JoGyJRn04U8tykQ8wYPC4ba+KbXV/zpDuGIqqZw0LHS8B6EfGEh7s7/u
C4Ozx6qBi/ZCnDNM8uhIAOH7P8EeIBTgGbx0rvk9THR9qaD+nQxZRMEo4niGyPftXZCso5Lv8pO0
cxvd1z11H8EUFf8YgWCet0QPYoaUsy8hVo7EOQlsBn2KfU4fQ7Yxe7IapGXb2utKFmsdPuHijB7R
YHu47bIWxporbp1+nFWPSISsY7mqDoVXT4S+a8h5UofguKF3TpLCBXm3VhBb1+cNkqomjdW/yn34
VRlWJvwOB2CxZpklgoGt0nVbUTu6g/Bduhq7KXllcRzu3VrxkCAXWrVAvr8nTdxaOA09N1d5rZY3
FciXVCajdoXEkJrJszKRtq8xkICrCow6EmN5Go5DOqP4UQlgIkXUP0TvNsjXxfmrWioiKBrk7cJP
xQkRk3AerVEhq0gGdtQbmi4Ooq1O2x0brRRim1nHlbynNpcgFm53ffhN5MUiknq0rrp+fpFGh3ur
gzxZI4zsRXN6EIAsxM63MFD1eCelHlgE5ya/QynpHajdx+PM5RhunWZlOKVW/SQH/lmi7CcuV6+g
Ph5wSQA3aJCK1zTDx5aYk6Q2cnQq4ekdTuQ5Lip4I313nvULGKX0+BXWNsmt1/a9xA3wMrDKF9rC
6EQZIXXF6uWHNphL+Et1/Ev3eYi2qgIhTq1EVEnyDdq0Tl2vThZOxwgypn6gL338MTb4dmJxgxu3
0ibkxXIZydd2yVWxA0LUY/TbBOCj6nbRzh0Pnp7y8zeQKHY/kyIBk77r4bnEiWae7F74WXy35t8J
UzBF6Qb93Bn8RqJ5EN2BSCFCYPly5+ANkliFguQcRecc+RetnvMSsyXaCeILK2Jt1GVio8DJ6rfk
X+CAqbOMOX6RzqehIoYKLbaT4fbL+9Jgt8EgBSYY9xrUc8NdWo4xSJN3cQiWHchYznoTrf30ENaN
Y3AjEdPNeDx3b3Ij1ymQCXWx7fpG/F7Loyi5a1uokdXe+IMdVVfS2Xg6Obl5wuj7EJcvzUv6ais0
NLBsN/BytXJfk3P7s59LMR/4dINYo8+NSShVm+PAiOqd2DzG7KgDV+zSiIeQThC9JbuhAIMrd3zH
m6OSoQ25iZdEH42M8weosqwMr5ifa7nhNMItZaefMN3x1dbb3QpaaA4p0X0Plvr8ZSzjE2I1j4Di
t2q/lRYWwMVFFPKCgee7oaukn55LWuLCreSg+uZpus3FErSWR0lU7lmQZmv8z5Oe469MJ2/YOu2B
e805Ppr59RNpRjUOzkv5+DUU0iU307RKOrmHjFkgFjqTSza50HJLh2+YMnTF4bDTLUIZnntpzl0f
eiD5UfQBH/2pHkbITm75MGg6P6KJ088O8R127PGGCDktbI02xVdk1EhrSkj/6pyGljzLf/Euiq6x
BpUi98GTxMQxRNFPs3su20JR2D5Dsm4vFQZTQwvUWQAdnQuvo04tVoz53nU2Dr5lfkEH3eAsOAuy
frdTmf8rb1ugYK4DoLCOOgnQV6+ia7pErPJhokC+PI2yxu4zl0Ffe0c69UBxfN02vQ39zUUAlNAo
VWQK5XhAD0TyfZFXe0oBzVPg9/9KKfvuroaKMXl9LP5/Ln+Tom79ALmXr6ZgV3In4jNGpQHnnw0X
IdNpUWGuoxt4AqWYjl2ia/z4aec6iAiyJI6D3R0oxxgfm6n35tWU9GScglOkpDmU9uYh1cZkFbzm
l8bDC22wB2GTFicGdQXjolK7nrS92Cqs8b2XGq+jNK/6dErb5sFl6tb0ctV96GQcYFI2/odFivk6
F6m1/pFBSSQXq8FO8vvTzItrI5/gqbJ4qsQ60GsgYLPjit3JOuSEeq7t8ebWPpcSXbm69Ov8wV9B
s/+y7ijvyNn4f6CGJloKq13rY9+HXIHhjo5U8CKWHYoJK3UmrTxlHPMxOCV+UXah+NhTw+8szjm8
zfG/SMljhoArhizIHGT3l9Tj0DQ2Pp4gSGb8iVKUGooe1ZJwP50HHKLM8fhhXFxppZGgs2KeypYb
4dMkVmfPZ4y3FSy9fsf3yyXXCItTSm7KfFq30CoGw98ukUk1TtoutnUWrLNqWOIsSDKjrYuF7y6N
d0XIO19KJks68l9C/35czWBTQSzuD8AJHsSEqSkiUu02Lqt221EfF5VWbITMO8u5VwAIsZpAQTda
7BYSygRNQcBWK4J/oUT6paNZNqtDOdImUD8Or9UafhiyqVqBnawA55ePbC6eqVVEUay/xZK5OeZE
K84KQ/uiSrJzZh7yLjvTyNKLcsMUhX4ZGlGkMHRzjZb59Hag7+jZxR7LkU+js0htuYBbkFk+APQ2
SOqcUima2v8QkMvpEUxMvp2fRLxZP4D1XNfJhLK61LZlOBbH5CwjivLeljW5mxNF/ib3XyTRQ8Dx
E18lnT5Mwjty4b3I5UGFw6gojrDQI80CJPdJBriVEuU8gRlJpgfnBFP3BYNUY+Kh6RAKTcomo+LA
o/ndIBI/SJcjiE+7SWOi1GYmyaq2qXaU/n5dMnuMw3JQH7zgJdFi4SBEh4veZyUW1BsuWtsVLX0K
qAO4vYuyUwwMnI2IB1IJkSlEr/8zyPNWS9imtrhHMrPmFx1/cmEb5UaWte5r7NEpoKHRyqI7R9BK
qjA4FeIi1G37vLBHbfsKHHVIf6oK2R6YHHHhR1MP1GbOSFGJf8MxijzsVIRt/qYivg4TolrUUXxa
oqQRPnPtElRWgeUJp4gKLr20pLk/ZarszXzdjIXE4VbrszrS6KIcoak3rtyVSMyPZXOTLQFx7D6W
F7K9GTfamnXlckHucDlThDorTwgIg1P01lY47tdp8MnQKoILMnE0ShJJ6vVF/n5QCudDVAGLOzY/
84M3U8wwFKFUZxGiSWMonv0rxE8asFrivkdpn1BN9FDi8tXOXxqNhOAH6FOuGskt+ZvZdzWc+Gqo
xCh4/eVRsFGEM6QlCnop3fuu/AA0e6FX4x9xHApJWuDja3HBr7l3dk7dm8yJRnwLExZIbxzEv8Cv
89BMNlCn5A/eiahpvSzsFX7zUtOYVbD2NZ9ZFvN1szeYb/39Mxk8EIRQ1sGKFuM7RCL4jEDeI2iB
cMU2/5opnpai3HnzXoVR82ZzmEKQ0nVKO5gyrb6EhbNZgG4R02FrYwNtJFeMEmKnOmD80MUVDkv7
R/y5v6U2O/yfvWABKAdRyw9XNEGgejf7YW41tBoCNwyVs0KXX4AYJQawe10/FuzvHvpfuSlYGs1t
o9GxO+Bfulaso0jN1JZLsTk1MbIH/+nvL/SNQdRfgj8eDekrXvxrfqyp/dL/FoHAnGnO71KAzopZ
W66Nw9vTwCHmJr1yiJ3JwGDwxVPebdq5Io1w3FU98eOK4nd7eV78AcV1GwV2ohIZZ/CBeqnlGu6Q
nb7Ss/kAJddZtaffBykGXPivZhZlM2OQ+zMQjYiqn1vZd/DIaUs9p+z5XrXUrQaN6rN/UYIYRqE/
/WAgqQUy1cVyUWcT5VhyozAeQ/ZzbrXFjZjEVP6ALaiP+0ldViPneo99YPLLZei8KL3bXPKGjoDj
sAU4d3L6HBx7WNNU3QZCaJ93VN+r1+sLdDmLbMB3NKscb0f5fUGZj5dehKrI8x9BnzIGJMO3Qa1i
WNR7y999gO0/DblkwZ7zEMvCl814xHSMGzfo6RDfnS548QfEX1XTx84L7o4CERaPB6fnO+A1g9Eu
Gqd76qWLCS3W6s0XdgMYXBd6htmoYyjLK71A7vM25jpHICRZ9l0gIoXFhNcN0Np9UkGCFm6ddDYw
jLpAOEepBP73sFVyhotxmdmNs9G1CjWpUnZerKWi5lwNpGRO5s+Q6XK8R/5mULSF7USc2bbHJxRo
pfOhAvp3qmBarhJHj8YIN2OKLuJvXqr9JsaBOyId/i4FLb2dlMqMb8bPUdCcwRnJutqdKvAYFvEx
d9gfDvhySaheoTObeMFMKHSQ0cvAC6jLoLPWoCT1760FgPOuOsAdCO/r//GVsLujtnJYgZ/xyMlq
5hMW/YfH82f3KnskourydJnXthJd+EH0MEui0aQN9/vBrLBkYPpfYaKC7nVR4AS95WkSXEJof1bk
IJjmCvZBJRDkl4bQ2F/XHOQr4uplsE4EoQSCeCp1wSK5/+b9dpZ2yLA3tThZ12F26FfuiF3UXcsM
lvovx0hPzCbnQDCNmm3WRnF/3cgOaaHHgYe/6oKmyZYgDgny8ZrnbtdkQiPdgZWK9KBP5Bwo7Ub+
KXxkm9RvogFtVESE9UG0tU1HXL6n61of3GrjSojsrxGt7PXgdbRCmz2jZPkLJlEsdwkdcE4v3Rs+
Oc3NuMNYI9hvHDyD/X/HnjMqm62aml/mq8OVjBAzciAvCPPFKvgCyHyRUgvy+xxFp5IgRaxzMekC
aolrnFhS1A1N//7mZ8Vm+w2xzs21gnqAs3MVcB1tGLYwTIt/FhoiA1pqu9TI5UgzziL0fR35wGwI
4LNGn8hltlfBmj0sCvgg12jiMlhzCXIFiZsZgKxGa0MhIJpR4iqWcCEi8NVZuv8Zh3TIDo6A0Vjk
YRV0D70QUswR+PV1boTsqA2MPFMEhcf+Vh/mem9zQb9chz14p21+UyrYtdrwjnI6r456a6ydHfWo
MEhBFx/0shnU/LeNX9+frMB84pBR+2+83oURPSp8gUPmei28VI3wMDJfnJXSH4ZruaujrEdEpt70
R5aZvME0lyO7Wz8WeriTduQaGphN9QBgbe3yKmKetFQ94FpEQmwVDYnI+xQoy3Sc7qLpM+Ycpeu6
feQlK6bWn5BLg0FRaSF1Qa1s9+EwBDYrsdtsXMnijXBQBRjpO/ERkt2o27btZ+FqCDCLah5XKsUa
IjLmYStWQR3O3cLQPhbT4xBSNsnyg/lV1Hk0cRLLgezLvHmnlEz2a529dCLLNTu96cGXFJ7hyrAQ
f8A6kGrt45aa36kfhKJWQHg73m5wiL4Fo7HIlxOIeX9a28UzWO99FCB+XzYA0dJWVv/cPq4Hxjte
XVMR78NgXkwvABuLgR4Mb78wYhQOExeX5iaHdMPZsoKEXr8A6q6g1R1HUC0UkmHqzWFOUW/pZvkk
u+xUW6b5ScQ2lZxQjZ++7C47FMFjzX6vSZ1cUunuFCPWYF6GCSog7Chg+xA5zTpKUi07wMYj4iQS
h+AVXyeuQHTyUHtYqzh9DxvqLOHo808NJ/BgKYjSAQb6/Xs2H/V9y1Bhpc7HuTp6JSXGvFoSMh+X
GlYqaZyo7T3qSAbE4au84Zxd3Aif+F9J0ZLCrux/VOwyTVHlSKvAeHcfZ2FdxpWGDDBTcyUynP/j
BBIZ1875rzoQsB1X1fhFZG8DR+mdy3HrHau58qI20rcyGt8ZtKxaNCXMA0R4Isb2T2/dBFBwkO7v
np69k1SWtjxVzpNrexeWc52H1RjyC8FHLNLk01m0PSh6z+bvQhc4HE0jINRoP/VlR0aa31UfW+xu
g97nUIVyJtzNiugvpkk2xyQW/NLZVcBlmbH788LtIr8Y6rw6hyKjqnfSOc8RZtGJ1SOlu8cbLMAb
pysXsoF9qOiewQuF+aCQciWLAiC7I9FZXVMA+xg4BETZ+Ko1Ghjoqh969dbeewppmXB30XUGpnkD
pDXOURwR+PXh8Uec3Ch7gehjU9Hw1ReMtnqP4FKZNcjMtevlMnVOaju7+3sUEWic5rv8vsr3Cuwo
E8kiWZgiFI6O2rHjcxQAap7R4erMNnQDLIN7UGVwto18MLJvfCvT/78grtTBTjIhT7ClfTQirUtG
yqoFtHM/cgw5AWOFNjo1WuN60Np+6qEJAld8sTeewtF51aUI/UR1b5IPje0+WwQkfgzIwtLzsiN/
mTZQnJQm3wucrFL5U4RlksPiOq+w+sFHFLa8aINjk+KB/WUaVpY1+j5dVoqCmsWdW1Zuy5GpKmBi
ZBbEO/f2kKj5+aie9UGdHB0zwP7ol84Q5KQwP7Ts+122TCuYjy8CgmbV3fkKtHffTjxOh+Klia1V
JLa30pY0R5wd4c7/Zes+wHTj3FIPBJcbFgXq1G1W1IrKL+1vAM0PXIRgnjdKgItGIsv/PKRBxZd2
cm7PLv2okGJ8pORIy7tpLJ5GrpZ4jpjWlCS1uQOiYSXmxx5E1VXotX1alm/Cptt4qUyq4IulD9Zl
yoQXrQymNe4BwY2xv3zYwAQM6/5QkBTG/YNdAUXkHn2C9rh/D5hzCVjQ+qmTCSM9csi+ZZnAq9cg
mXWD9LW3pFqb3BS7H1Fs+5mkDnfgHX4U10/D0kvetHM0Oujo+vYFqGVoHNJkKeVWBjkZZnnNPGFX
YEwgr2fkaHD2aHMtebt0nxdJiXp648u4rm5JRJ5MsNDgCBDu/edNGfAeX8gob5TBt/1czFaWAtdX
BRYrAVHzjm+Qj/DhBMK42avjXN1mNchCcS0EZOpDUto0pTkvu8EDn9OyuFdLzidf9/NbYjKmu8Kc
KjY51A/meNkRuIAxyiUhKkC2BRs2CS3UYh8E7M0vqMfGHlY5eONnsgOd9oq9Ca/urPMNlS9fqGw1
UEEQzu5avFSX9iTpP/YCYTlpIrEnTZ3npfWVaJi0OU3JbeZRtTm8vqFgseQGfhE3OFvp6H+v4Kyr
YUeyEGwDlqcD3Ap9pQLqH3SpWdeFX35zp8RSNY2gnFIjYRtK/Lb20sC3XFOKpfBcgplML9qk7lPI
R3j8lZnc9YDIbwT5fa2qpV9/P9vhHVRr/GmBMWOBA26mpaFy+gV0yiSldUOvuVLawYAsvACP1DkT
F/td8lFw0NQZrorDUVXT5HT/gFxWmTrVeVxFEzt9ghw90G24o6dGVmGfEwU+bGDm0wZov1BCwOT/
3xuuB1DD3GQc66K831vP9liZpa+41TfUsOKw1nTT/E2wkCa8Lwofx1NMKc9EeLu4QTwPGSEUnkTj
bZl8KmlJsBpJfZBIg+EXZ1tC9bJNIy1qLyAKyrP5FQUikUxJPf+sOtQIqGpYnQYAjIbOCUeGPMT/
xslcGyBUZAeEqrQIGl6JDVlixywy9Q2m0XfTQeBd7rBZxn+aaYdCJdhf3Jn5cSumHQl+JneSJFk4
cQelhOjgtHQCHMAv/gBY8A5IK1Gs7n/4vOnlbSDqvTDo0byPPtKvXz+uFtqHHZ4nrEPbb6KfZiYY
iv50ubZourWWxtlhDk2A+RULcUhOsBeKx0d7H/pgVHBce9VYF/MTrF7O7j0em/LrkPsStcEtLiuO
yIr9Ahs8/IQf2nncJndZ4vQWy+fusHKmHDuCTWtqzSa7UZcD73jk5+HLroNcLZZx4nmvjH94Ayjx
nfGPqT/XNZP/B9t9QjeGg5thIlBARq1x1VnCBtqOpTbwYM2lHh0UJtlZN6FEw3L4MoJgi2TJ/+NF
Qqd6bJS4QRfN9KMApZFBFUkUYxTqJC8AYMR3DYpT74rS62zGWP8C5WB+b3K2YBhP0UWtVGuPF22p
xTaYw6EdtVoz80zhAeC5d7PrbrUBDndt8vnm/YmBk262SMoUF16AcYabydSfE0Whu1P+bBdy2GZO
hGbOFmV8K01fQW6LaRdlMe0ui6wrUBf1FRTCUNVNf2gMXFUB9zoh6bcxAWRWitIlqL1VDXsM4PWv
qqaXUYoVSEV6/mS2xK1F1syZSwZeTAzZpaIcWGH8sUN5FD8UE4ZwYYyafTJbw0Vz6nODUFnNoavA
BtpcPRp8N0+ftv/FnYrv6t/lo+FZCybKO4KuYHvXKuU/5OFYXr3CBKKhwbWJ6kMwZP1BZoyf7kD4
MUISuZfYjTcZgpsOmQO+jnOww1Jv60KC+KbFYSUScj0BhgazaSk9w5tQaM0lUe5pir56LBAaMP4o
k8r3YC1b+mxh5mU0UEIUcn+Jh+KoFy1D1LWdOaDgUi8AqGpPcTLqscCT4HCLAFqpajR6PmJU84u/
k2wHm/Dravl1C1FJcaUVr0WoOjOj0lgaYnBXVznd15LoN9mQ74rgInI9hh24geRvAdkFMbtGNboM
nw2h1Lj7U9XyYUIHV0TlmDCY2sU/aL9j7QlTyGnpyURZsEw5vV7m0coXddEdTThhrh6V6Kxd3/Vs
N7InUwrl+wWVV4gTX4Hr6d1DrtCw79+3A5IHjcVs7PZ7PUyb6SHLWaehQBtFXzqecYm4MgLlQp72
P0UtKvhsZX26y6ww/a75caH6O3xBTX138UkFxJfBIsCrQj+zWzxRyuiJ0pSQxaTbL1EShJtMs0RM
G0Ny/Nz0d+eYA+u8iUvwSVW7TW3CfWNbzBlydqSYBXeOuhgaxjFYliHFRkLNsIRRc1FokFtJOD3w
IFHHZcmAlYaxr396/gzBAiaphibYICxEScB3PzAL7gVmPlCiFL/f/Jsir3kPCzM/su17Ou0Vtysd
DnnMaQRWLh9QQrCM2uKZr5nXxpYQ85k6oPo0a/0dC05wSm1UfX91/ludIsihYI6vAYf8qkf/Stvl
NQifuvXySa4nVOe+nuD5FqG7YgIvHce2WlX3sfZF+mk1Xy/dtqOcAcOsdpZKwEHf35JQbNepoegs
FHH/SnVY5vWDpvJ1VwnnQcTveYMMEjXs+8oitKqcW2IyhRritKW7kPsX/i2p8yS4QzuHgVJIS8Vh
u/axowa/3thXkGxgUQq2C+iORP9yA2t0S9h9MA1bElNIUqN0vBeoyeaHDLWcvYvrz8FBS2yjB5SI
4rX5b1+LksuruqZ6vuzPTpCkSYFgdQQjNrNvUFqKof2xuAt5iEM4uCdGPRFdjevVDmqajszWuKEV
YjI+6+Bcju4n1IBkGF1TDedDOn+nOalnGg20QPOHeFwmSKlaPTx3ZrIA83ZEoW1nc7b+DHAOIVph
KzTuRGL2HvbuH18xmMdIaTuTo3Lnz5zpZ2TwuBw9ka1zFFiZufK584cmiadjET0a2axQ9tprrTIh
K2lrcOeet01lJ2EF7KqG/d3FDL9wETiskujhxausi/cXB38DhfHDZdOzX74hinPR6uM7ab8Vmhdj
28GXUPMRRVyLaBHRzIPgnWkQtN1LqebY/rtMxPOC1x97C9BYZP75PUsgawxyGoK9NjMGhglM1bYk
jOcDtCobdkxsU5oZ84ViCf3jCjiXUnXbdcMUG3SE2K/Q8TA1Y85Kpad1tcMjMPc+g1Hiqy/XLJpp
paXWWVpDItMpSd4ZynI/PMpPtSfO29Dctk5AQATtDHtG/ZcQDwEjqtq9H61D7tkKpFoJrcGJlZnB
qDCMJiFWzw2Qc+B1zYNR3IdSOvTI0qwpDsrFjIlbvPgZohsSTZPZEizznjlqayCaYzwnsPU17BSN
mgo/mQ0R8n/q9Hagy7ghy+chI8C3zITqW3hNZoaLq6Y0LrbKCv52okNc3fSQOiLx4ur1MLmgJuvp
kE6wMY5B25qubT1xZvBQVZnJ4SquhASJkYWZsOJuTvnJlCOtw6/BXWJ24kJ1of+rAaLnKlBqu/DE
SozLX0Mn+u+TiRiIOWEuPhGC7m1xr/CCdkIk9zQ7gZCChW+Y9ChdqB6796rBTF5UQPAnb53kvU+M
sleDhxGa7MjjYlMxjoiIjT1sy2+N1bmsj9jsISzc5v8oUPBdvP9Aa4VQWR6UGcLSD+bIlRkJK9KZ
CSQ8ifwvzHin7cA0KZiTBaAm5uKugr7ay6AaPdhtkt3Iw43V/8zB2xea5xVjtP8eChA7nYDK5n6x
5vKlcK+9qu56+TXhKNvXL0oM95pfCcC6Vi0Sio/IvYT6xtnpyWdbEGD6Zr9eWezoEO309Zxliscz
9PR8uGGBkuQOft6jcPuOL4+8vnt3Ipt7PJQ1+0GpzrwKgb429VpQOiG3Bplvk30Ch8BnvZR3XM9w
n/B3g5XxzhYAbB2ZBEM+5x+k19/s83+vCEfOc1N9NLXbhRB3rajAhWEHdNIjofpRJZcS4AjTFrAZ
wbHD+7YB3DHx9XyiqY5/FXQ7ZeeW9xA1x4AKgzPdO7IIGpNRvnsTIGT9Nm4+WgpdE5+/DVcKfbHC
SGMLsh7r0y/LvdBM81oS709G67LmXgyki0kxPWRsnqFG9qOpZxctlz1SMZTAWrV5ViXf4KEAeCjv
jRsGJJp4/hxuivC4+5v/t/2qNYJDj+VbMKBZHOemwEkPn6mixCAY9Wy32gvhqHtGzbFUDQBzjUIb
euxhKHrhI+M6FsN85TabQSqQrqaMmHEJNZSbzyWfIkWiisvBVYnwB0dEzMAdM2Thu5PPiBGG7+Li
daH9uxZExU16LxwVQL7uDNisobVKJKMLgovBQd4FTnkNZ8yB1wthLDQn7j9/ZcxujPnItT5KsXPg
E1YIAmsFbEc+U6MscyhJVv5ZD5PhqngWFSQ+UepbhPwtjZJ8NhN15TBsu87vOQcXrVX1XCGnCGPE
jJ6D8xLENVUMUqM2uMrV5SD5pBZtC4kvbXNLy9cHwlpUKJu79qpYbU9b+M5qJCG6YHXpzFmB8QXj
4vCj7kA5VMFUejPhAwobYMMptR5wS6jNl1TU2+3fm0xNrDF6IrhWitQlgK3VAIrWbz8+4HS2wicX
BPpTZjnNXPvhU2ksqhEOCAHnSZtOaFU5qXfaZZEvRq4M5amWvo5ppbTVriXgikdCBZQh20ft1T+S
MorIxyzbYYsl7IzBmPz7UQx4aunsZAA01J2t8dImIRJxU5a7awOsIhPAwF6hpWY5TeOJBHVwm7+Y
mUhKC3AZh2IjTDBVlMBRdeEzEcTpXG1SbqshzDvXMGJxsSG1JHHeHmMKhJbiLns6RCmRH6CxmRaF
euB5ohmGxTlDNp7wQfSvv/BwMp/j9WujAUY1d2xHSglvgRMA0L6/5rMJjfrrKIt9PF9TqyElOipv
aq5mP3Qp2fe0ij2Uqcjei64xH4rhJaC2XSKjdJzeC3ypAFJikhUZf8D+mU6p/hwuam3n2/mWIFNz
8Y0dRTKCo0QB8elMsliC8QAzTMEZV/Ewjr5PF5w9nJwfVcEsGppAnBIQ61np0mwqqJGPEpc371DM
d3nasMkkkIvi1NR0VeOjh4WRQbVACpY/2YUwGaPPFN3RZn8m+vIAht+4QpAoGlCtXBHrIROvv3jS
AQQSJmG2GDQjGlWO7NDmpYCR3YlVyxai3N7APl8nlf38jdBzuc2BqGbhmfykPiJD+pHVuQDwtf93
TXmC19EnrbHvTQ/lrbxYvPOg08en2bbxKHXTJZ0wurD8ywcDxeLhCf0Afoa+M8UC8LwM55xfAXu0
3bBB6iQPVVGUu5VJStmL/uL5FCiMLXqI/RTF6zi4nE5h7ackddmpaeAxAoeFWEy6+1vDKXEzDizU
2NNN5CFA/5IqdH5YNRjIe65aWXdMgXXSPSfj7VJbD4C5B6HobkQkbuS+Xk5yZu5SxRdGUAk5GAjD
+3GGzBSahg5J4dy2NFeqsurTB+aqrJs/0vZpn2mTGSMKYY1KU4WfDawdbU5Y9d1pEQhxM1sg3c5C
fm5mOp5zUV0O6H7FU49S6qzff4wP7sDyACts4W209ZSaBC9PefQdg/1KhpBLTS4gLVxgqmpmsXXT
BJDQ87RWPMc1Hs9QLgftQv/wSbbxtq6OgyR0Ine6TxNxtYF5qEynUrRLzaXHmLnoF4il5cuiUWoz
8GRW9ToEjrdmoMZr3XKHHtzY1/b0rn1AABiXi6F/q1cCinw+dwCaTvNsLJcFvXty9FBzSLjBMTTQ
5a7d+SKK5G1vIKGolqjzL+2QfWNoRHgiBtwH5dRXT02mZNo1glZbPcBdMeA7LX15yk5nR6IwMn5c
kDCnzKGoELWOHGsHJm6NROjAJaLB+82HNrX3MdG3kQaCwVEjfTpmHU2n7I+U15Aon4fr6e7sD3MA
2sseizbqsl5UP1osE39ocvPud7XgccyWKinbkrttzZnK93JH6jHcgBDZWkUtFno3xiCOaVgTULGg
pKmtNfqji6yUFAGWN8yh2ydOkMmQEHOxWDpvqpSxNZHfIp88teIOzlui0o3B8oQdgPRxWiNwGASP
rtx9L6eg+YcaRBa540brNCy9K+kfHqoaGEP5KCcSbQA2f8dQyus04+ffam4XPr3X2LcECt9xZQop
+QXi0MLdBFpZ3+0Nhl21giRsNehkgYvOD3hocd/C7czeVUeP2Xd2cei0DxH9oia124riLS5XIyzX
+DxMv49BTlnR3SosZcUnmezxX3W/xBgrvALuQCpHci6Bll95ArYiY+YSgSVCR66nSXAFvaoRefGV
Hxvn/Y3wGm8cfZfSR3zhvy8PlH1T4sEO50K6ZJ8R93fwoh8vS+eW4CaCl7gC+e5JY4PzI2X6QZPc
yz5bS3k20gc0/wHBH74jaPXW23GqOFcuwn2+bl1GP3xxwktvQII4ULErE/nALkh3UaHda+q9DbBn
UZN81dqIbKaZgSW3hT5tDkd8ExtpPIPrpU0ZR72UHWnYbI7yl6muOIN8NaudR29VF+AORSblIT1U
EmB1y2W7i/h2iK7283+xj6xEyfv5w3OAeVjzINURswF2hHDD5XVQ8XSKVGFJFMFU69S8rzY8A+O6
fMqO35GNtiA1cddfsdo2NPhEbxCTmipu/Hgq8SOpmsVRRecB0olOFdQn8yFayqUzYWEuyzavmFLQ
EcZqYf3sH72mMwuQ0d8tG7P4OKouDY5HE21+cUnUoeFkaFwatlpgvwwCgElCn5x1UsnROUQl4JN5
h5WWUvRoNFebG12WI6PCDz3CTxjMq13gAy/FV/orlC/i0NSkW1eMfzQ0U3p4DptU6Li9D+6tvfS8
eBAmFoOzHqtS771ypiKmTNcJIJKv33zMAJE1+HQ5g7ClzGpRUTgryJb5P0W+ABttY5dnTjtCKN2N
MR3KEmOSxk3GM3ER8/nF0Sd0fiqOwYgiswGeZ0T+la4ZzRyka37e4caIloeEBgCP8oF80XTCYRqI
gNN0HdSQOROzmL442ixqWaynFNcCH23JVIqEYtBYVr2mc+TURyVCg3hfxHbEb+yJ8ILIWjwAJMKh
8N+imkEEYnTwvP6NNQE6Vcd8FyVHif1ZNFWc3oFzvv57VEzAffq9zE42rWjoQOTC4RwWVEiRlKdM
7eu75joUOsdV2KOxh9l58QH+BPuHGiSHYNDgX4bOxvcLOm3rz13DzHE7o50g/iqFQ33L9KMY9VFa
MlXwXiR5IK/oBKe1ChvODqug1+c5PcyPfUfdDo0CQy54db0+/mTualdzziMeKYboNQmfFPEILIsd
OtbfeIN6CVCIw6OL2Bze9dZt4HabR3WaQ+3Z9VxguCOAAjXD+7Q05vUeIak1NmiCHAIJel6NyCsD
ld1Im+NiZ16TbGqy9JIWUeKc9hKcsHvmbPgC6oiBhqd+v/Nk3tXuNroamZnuiM/uqyDQqze834jt
TozVaC4OnR65fKATdO1Pk38if20nT4dgoJsrcxxAsxkWyMikI7XwQNyzafoUXflCT+VLtJa+DRmO
tHNrhAfPp2fzg0hWLFr3R9Hl3saFYuBGVXOs2Fdv26aVGECANlMSqZE4x60e0uQG4rS8LcsSmbkD
5Sx6ZlyAn735yAG4OvCHX7LTbwjsW2rPeuV6zevzhldR/r8OIUFsmWWouKFsU1m/nD3UNXKCL5A1
jOY/ZKjjCDAhjiQ6XGaz7HwiewlIF7yfM99PuWPt5Dnrp6CWS0IRe/MDUxS/Xg/tU6pFm90VDJov
SRdN0RTab4vceSWEUk2ylWW8JnDeujQntWn/Wdj3LGJJLFAIsTdj5jsoDXViBJ0ViO3Z++tKO2Q/
0RlC+bJUBciJe0TDlgrwgbv2OZURoLqbwEkBcS3NRGO1Bsn25XeeoGLBWxE1ryuZglQIE2tjRQ8O
CPn5zEhVebaX62OLodYXuejh4DCTL2LFx/v32yw1EUekjvYqbu0QhQFt/bPQ5bZwCQdZ5cDyCTtM
6l8C1HHE4BCZA8Fd7SV8bbTfcOHeNrlMFBcg1TV3o5XElKOMBscya/HK9N2mtIDM370QjT0hnGYQ
Z/9gRcUdOYQsKTh9K4+U/f3MyxfIy4b87hD3S77yvoBOB0HM4cQNHhP2luFVZ1362awbH1ZG5kzB
MAJBnZbw4SigcyzdstvXEXqx+ktUyirlF4iG0+d9S42y72sMvxaScSGhon+GHf/mIuwZ0olnTlIL
gZrx+OSDT4wPqdRZ6NgbQeGRoqsco5PoY5s+0jEa5pvPwQJ9Z08dRNASpmU71MuSSPxnpWQWrPXr
ymrx5NITuCHf5g80YxYpD1xxCc1OvJJNDYLzsVUBG8T24z5gyP2IFBKfDvgHM0NqwDnDTvVxM8Fj
DaZhkFb5c47HQDoy6E7ILcGuWCvvpftbhof8wtFOALZ+RBLzzvp85+AsXVFzB3FiBiwocfJfbxaD
P43kui1dadfq/rd7Tf+Y2Ue5pC4zxqRLWmtcdGmS4q2AKhRLEKjrLli/xtRAowGR9iFX2GR+EExg
JlqsgpC81lqDYlhT+Roj6p9Pm7PmD8V80UEPRCy8VfCPHChIPnMOUdFHzl9RoisjyyUkad1R8Sre
HxLcJ0a3U5csy9fiP3b94gJNR/79UecQAbHsuq8gCV+Si/1hf45fLJsza1Zat7msVPAuhhLRKkSQ
OVxNewk77haA1MkAJWnQ+R7Ise7Pfc28JwKd/bOxWkcFuejUxG/b/gq+WDb6S9q6zVqXFUSY+naE
d6xyHXZze5FLTc3v7ohrBl96fmngKiSpOIdrC6zdzL9FxPKPBD+QwYIbv55tNCpvoW3IPqyRkfcj
3e4Vy1zCt6O9xKIykj/kITRTYZ/kezMxbYUJXefRQEScaaGIm7G4uxmRSa9JOcAnfOSP6KJ7mb/O
6GRZfjlk/d4rZH/CBKXtmUGDx9zx3J1t05qbvgexurTQ9bYJC3qSNI3KKl8qwY7sdTDgrXoHbn5K
fEJXrzyk6zcYEwndAz9vaihN0cnMImeF038mehoIRWNxZvbCfQI1kSPwpZa5J2bjsGov6J1ve/cD
bpYauoCat8S7ORnmYkanVbONaM8yrCPnAVcmI2+AuDYSkK78Jijr+bQqh7YPjGEMaSIZ4WbU6s7B
2CJ36JoznOkO+Z81sU+rvDP/cNXiwF9WmSDPOrM48GkqXtnH9t2Qz08IBZrJboLFBppu+URi7yjG
HCIAn6igdYKEHY+7csQx800t80O3QRWx40oWhriHFUFXUf+06+OYltDXkVsjDsQAqzQQbODkh9kP
i6sJkshwOc2Et+8mkFfGlXvCQnfhlhjFiSX9cR8CLNd0ZZK/zj/sH4Bi46yhneiZZZjzDpyR2jbJ
gI+mkAzLtElP7FN+v+AqZ6mWOf45wClTR7qYiiNuSvN1EzVOnjHlRrHOcEWQlJQpbIOD70D+yxeC
jpZIsUA4yrO37+O1QEIlmbRBWB3p2bo4/vHSbsVUygWYJzjK5IhsGjkkXfWLT/hSKAUig+p0+nGb
dbNPBRn/8LpbSeaN5G8bctFAt82SuuDd/H3bbjaZDd+1e+fDbt3Fic+VkXW1aD4PPtshPLYH/zsr
f+h+Hc8ndaFUiBE0TN7Fn6Z1KxMVkJecAPyarALwYPWX4S2enIhH7CQVn1XQABgdOA5GWsxPqPn8
xMewWrV+LN8NSKG3N0rBeyw4wcUVoQXdBTGBqt8KRidVwX3sTj4lfYVzuksPW0Q6JLuQJKYrSZya
8+f+ziQUPrXF9EIYXPePYclzcMiW5u4Cpoxw6wxz4GjUqwi0i9iXpY2OlFQDFfXKd9b8zssJ9mO2
w6HOs6ikUkKlxpwUjSsTqNxygmJOx9nveoZmbZPxKhDE8ch3QBzbtGTMeOrNfQRG1Z5C7kYOAXDA
DcncxjNJeTdZrQVZJblgvdvkIzyy6V+w+4WvRt6qFczR6d1N20w3LrklGQM2UxWc4Jt/vqA4rJiF
FlQtLFBmWoekPK+RHyK95kd7qMTdGJVSCQ9+lTFF2+rG5FhmU9dvLbzkPxD4WV6RVww9v/YwK9E8
n6pczW2xfRMMx7yowUUYKKm8RQQo0l9FaRx7qy3tBsCgQz4bbDuc5q1DL1DXG0Y90PDrQdUYK3zG
Zibd3ENUUsR+X4uND5d1f1xpHUv+4J8klIaiyOU4ywbUDAJrFnT0PyQz/tMiqgDwbZogwI6Bk5wz
SFCO5xPQJeYL4jBcTApUzDuvp2LXvp3bbkqV8B8iBhouYlzVsVxFRQ3ZYtNVJK8uibslrfWL+3PK
aESbskdWlRZQ5rj3t6yAFXwQn68NKLMKHszc6uat1l3UaMGDZolZT1MDTvCMfzbHW/UYFXGH4yOE
n2Pri24HSo9w8GgTHzzqZOT7sQsLGZYtgdl9oLXYp1GURM2NEoqitBMUoxX6DyvQBMjfUdHRmkA1
o2F/Ikl2OE65H05Af2doGQvN200Dz6QV0TpYNH3Tuf18mdKDWU8q4u/VM1MuUfPhmyq/zjXf4s6t
zWRJQexTlf8qyYqsaZoaHVCYS8SCfBOFXrprg8pH14587Qar5B89BLEmNnRiKGF9bpDdShDVAgIv
wkKBeMX9FSlTygpwbqK6BmZSoWoblZ56cB0db5y3sbSwu8D7MEfatnvBhGB72wA8eOHdwU0rMYtX
TRf6xUtTTXTbhvfTAWRu36P+4DS8Rq0r2lzkrIhKJqW/9pvKrouOGK67Q/wGyMe7ceqCluCSSn6h
sC60p0cfHr6ule+WqsyN5fdm3ndTtpubC38JnV8ziGlWJvITHToaLfnDU8iCQ6iKKBT6/IGHyQJ6
5LWuSRb+L3sWSuFlS0desbW0Ru30xhDujwYnoLBaeFt9orok79AkFH0SkyZnojIDtow9cZYaQSNW
xYkZMIdJm4kCZlJ20joGLkW+u9+TdpBaHo4MMgAmYMr0wyzCRV6YClv3EAeqZUT6s33fBrnHXAL7
sLPXFLspBzQK2V6QmOYMzOK6pQmTQJSlkdSL8fFeA7qu9uXkmHq/owAkAu3G4dimyxk0CEPbVc46
w5yBWJWltdcHKKiZ4D0YeczPv3c/7dR1QQN5QU8zurYRuf3NxZHKkV8J6De8qjLpROvAhuIjdchW
2hdX45P9FAO0awHnBP7Paea1xF9NgdDPmAnQjj0Zb4OJgNAg0ppqQY0MjXYiUzYg21gbJUNyMfio
RKslrW4JQ5JCG48I1FkhUbNR1AnU1AxZr1UyoakGC1rf6ogLAiL42J3XnDzF1uJElBXW0ujLqg9J
ZqkdlXvREHjQc8iiXJAWdltcPIID7lJucH9RnTciMAx2SLRxctQaKJgVq1WkM/raH7o03xwfCKpH
HNN4sSaOUUrOmQ9BIyLRFJxm1W4KQp6859lqG2Osujf3D6Qj+BS0OXLzhLrNsvjAGLd6AdT8y+AO
jZAwYCeh1oPJta62StZdTTJTYv+YBn8o0tA0qxdKOJsNfxG9bZlOQXoJj5z/rindlfu6IbvCSe68
B/hFHuoOilSCgUCRqGS+phQIlfFS7ElazbxBwKHqZ0x9tbHJzFKm/hKPcP9LgxpBs5Q6x8gWreoS
eeshTjWESo7tl4ErUv2uzfsT7H4bruf8HR+l7+H+IWKC5fiHGbNnaSuHs5jb8R7MAjuE7ew4oaAi
5QmjXVhXpK/0fIlbyQXmcNItNUXuNtFRMcz1YTz4qgezz95p3HeDE4g6ByHmZInvPtYyrPBG24Dp
HDDOCO2hmVZFd+h4gP2gMbK01+Wzp+T2yfWWrJCT4CDsoLSTKDeyNRO6j4ZM0ak8WngF2p6HFfY2
+utqultF64S261mg1qxAuRF1OJj5iKyuYrPz5fsG7D8Pu1UM1dFJ4uQ37wjOoWQTu+lxzaV1n4bw
ID/+LsYgQNdzYhogsw9vz8snxoI3768fdKJJZci9gUVKB4c/FONvYvEzq8xM57YqA3Z3cnVp3FAw
Kx4INllxruxkCPMp/mZkOx2NxPqw7P8LdAMgGhQ2opOtcIj8bBbEq0uk2yHJcDq1aYPeYmV6cIla
Esw68phcqdlMHiFDYFJePLp+sBNvyG9uLN8sAtk4r3Unz6CNBHshO8EueF5aNqg/qXzT4V+eDMrO
EHehamhnKkBA3K5veWL95EAJwvlTidm9age1S1SOJqiMoiVzIZpp2E53nbOPmnS1oPE5ikqLJg+s
wstyQNgxoKwwAIohD/KvoIOFoiZd9FS0H1CbgIQwUhMCSgjSDdyHI4oIymn/l1iXKBQo6Be+6slF
RtuoOyq+FErEUj5CjQ7KeWz4vUtQClk/m0IHMADqljjThtmBy9IE36Iq5CBdVVQ8mZrKUChNpHqV
kEi6zgWfj5NyJ4XhPxbP0cN/6W/DmvPm9baZIQyv5DjYkbKfDCZG6615Q9dFgTSE+oqjUrllIq85
4Phpg9FclU86uTA4FsbvqUWZPSmBM613Ul+/V6bXCPp4xR5FXxeu+mqBpQ9ELWqJmsIWuPzUGfSX
MPq0qRFxezbDKfvNceuWDVo4suVNQEuFa7vaaJnNn2TxHg5pQH0Bv1C+cb2LWdZDdLan10YEL1+P
4tyxM6+8OLE25e0Uyaw84YchKh9x/gx3W44QggDpJobBEylF2Lw2YlZrIRLxtAR+Y0Ey0KSGEbaa
ECyqgyTCZ9E00vqp0Fk53s5QbKVb911vpkCqMxRrDzQTTcObagTEcIQd6jGuWVkPvnSxRtRH/GIZ
KLMrmaYGAiJ02MurORGklbMyR+2fJ09haa1rzkf46lM65UUx+Fj71mGNNzZwI6dnY+qGL/TXtxDS
8x0q48Avy+PE7pnWcmLbVKmHzd0Huo4NrlUQVYKC2KaqVJG2wc9kFqh6S20s9GJCnpIviFpe9z5E
9yMteIY+rekwvIOZ4+BXS7xUu2MjdPa2IymYXuf5/jbzz2De0BUlYMsxI86Kifld7vp8cxH+EYVG
FX/0z5GJg9dWgyT5dSm4nbQbKoBNIpB8zCHZuQWdlPZr8GmIqm2A6zfjMZ3CrpOfCwU24+Z1LukP
2RW9AUHo1ypOOxzguMCPDDMyDGKCgJ1/vBiUy+IPrpA/xuuAYW/1DssWRJ+cdfIfqXTqDijweFwR
3j3vtq7vvFgeFpk6FAEvRpP4ZQUK5p3u5/V5o8XIhtmGXoVfZfQswnXvzvpreIqR3+LNC5XE+8q6
PkebA5sWB9Yse+SzA7zRR0IHMH8e34nPwryUV+LJdCnTreROf77QppvPS9l5JZyH9HvW5S98qRpL
lqdaRl8ulhj7BVcpgZnElanirjqeeb/oqdB0nbY6NBUX06jtgvAzfZ3bOwl7R2djs/pv5eJbx0SK
IAtda4gzGWSnotiK4hhKMtTk09392DyXMXGHEv1hAl3wWghOFOWMxCI7m78CQ1d2bG51Hf4WhjR+
qPf7v1BFgeNlsXOpjPuRsuMSwhzHXYX/xWcS53ey6LMJJD4kP8BXBoACt3USiEwOp6FN6REfkqiP
JmqxdL4S1YbWajpOD9510tdGaFi5AfGU0kk8+FneQ92q3i3IDoWcLGTFteDHML0tnxnJET7ulhSt
gV0kztjNMvJy89QUT8PgMqRdeOJajSkd3qADihEVHb7+rCFr/ZTxZxAysRZlYlhT+wR53JFA8Jht
CJznHiqG/I5hZGY2TyPpUmd8oErIwRCfNo09b11OE7daZyu6U8NWMCJpwRH41bhEwGvGYQbFq6Qz
Ia5sbdOPwCR3ZTN/KEoE+mYoEcpR5BXffWCQH6TrDqWRmvsx5l8jp88ExHV6oGqLUsroicFuWeCg
kEfHc+/gBoGMwci0dq6dOF7ohd/ETfN8IjauX2U5/mAbR0ia27jTj+pjgAqAPzl1dLj2CeSZV1Nk
pzRIbu9otjI2v9lGGF0kU04xsxFm11H3Vh5RRLQY+/adkp1gr2bfjIddlimfoH9gbfUk19S/PEA/
OSiEAknIYuUlcmfeUafJC/CeIIoqB3cXl46O/fHue8EkvQqRRwrxX+XLM42Mor/7xVMOiOKGdkEO
J0hHIvWbUZq0kg9lHi/IKgB25/piRmDBH+QcuxXPPiiJRGaoCeji+g+7jZMG+Do+cd8X92BwLiTD
3uE4F2NeK+GRX+XJwTcYzgECePD1bM1+C0zhKqmXG1YbO+y0LDTRhzV6pHNQPY41VFtJ9hulOe3Y
ZrkOWTQiIxP/9iPn0GnY3fSkrHQdKXAN+l1ArCiICVpr6456Yg0dbV/F2dQo7eM5XYp3ae4KT0Bl
m8YN2xZBSi94uOeseZ3SmS8tzhnd4xe8bvJ7rrNtvD4DudvJbUQw36akGdL/4yw5dKK7QI9aes0Z
JMIhbhHKA3fdw93IVQSoK0lJFdX1CjUHBgtUfqWZA6RXanYqVI9BhHbXxQ7w5eGbfUflBZbGAv/W
hakSHYEWbx7Tc2oM7u8TdcPypHCFMvFeFfS3SzIrw2ZVmF/ilBrSVi872N1gST5sJJyxuOLzffpS
xvKmmFts3Lg/ei1V2EPChT0qSr5AgmYzvtHHvoQcKh0dlMHi5xBhhqdSW466WKJlB9n8Z86wFo+Y
/u9L5lozjOutC7MdHr6pZWrKXFLRRHWwJykzby64TPVpvlHAf53r51JTcPCGyM5wkzCldMU48s+H
aEeixfjkHdAxCUgle2Lx+Z2lsQzjgQWr+OQk7Ov6+u2CdW878MHaxb2e4JKVnHgqFt8SirpBTFxS
ZUYyHkLDIg8vtLJkWl1iDQSbJd+irWE8v/dSva6KxEL2VrIAWyYewH9TdezCWt32zJ+NjOl1Wk+B
ig48dHSWr2fT7OYJKgmLjoOlglj/Hl40oFJ5otX22CePqOojBwJjC04PZOs3POqM+lHmXtc2YXjM
W2l0uxB5EXz7sjgrsPlLelctvKanTvbTmJr8A+F+tP30xcT3dU2guoEgPs3XQ2Ko4pEN+AZUQQIt
2XXCscL64BwgbOlikEStVCVAXrAXQdrMDk6BSYji5wjInoDN59DFB3hFDlUEUFh148gEOAFafKqj
Um1Hfoa8MzmV4uRQcCa/EM6yV3zZCycnXp/3VN9TQk/uEDqsObUQGygRnh43tZQ8a7CoEm+CR2q4
a2dlGpTxiOF7BlZv6iSQLd95z0gwiBB6+pr/uudomQ9F2pb8dulBGi+fABFYCR/a56KQcG5wTgWB
C1RNp6FbPTAo0tFbaT59Nph8eEQKIseJoWk/G8Kyja1pQ0ueuqJGHff/kc20y3KI2ZYWi9SoMvns
Gp+wI+TVQJ7YJo0WTG7aQK5jECKpiZV/DJkB4wjyOjTguKMY/4eacYSI4EJAWJZ3oZCIYY9yNQfF
sRjkIc0iSMveUPYD0ddPwnQxcGB52POenNG6K4MVRNXJJb/iC7tqD4tnAd3CPf1iHn6asr2PG2PY
v63C7+I0uN3P1GSYtAg4BraRmbc52e3dXiwd4SU8GBuVRJvXPL5A4qhg69/KwvpDIg8vFY2IXrMk
HKKC2xj2ZVJEyvagSRuYtxs6Fw/xRzLUuLLnu066tg6jvh7D0SLxHACrcmitn5HS6SgtWROaPA0W
vRoKr6Ei4JMasYlVsR/BYFYOnaY9xwwz7pzCHa/8mNL31KG6gVNXgAlMppwrH9A1CLt9eZBP0Yyx
3OT9DeLhoMR9G40mEgqZwCwslrt+iMevqS/TIAuBhOA28PnobaLVH/I4zYzbWgIMW0FfpsvvzIq8
2fvrTf8GwQVu/nPyxggoGyNNMFBoiI424J4hbVc40EJ6h77eODgUk0ovL0aSIKhDvD/KbAZ09d41
caisNnYuonpnZCXl+ucJRS0LUo/PbMVvMpk0qxreh6jOEsqQxctecyk08lz9svNM4qkE4zm7W7bF
bAfwWEf+9KxuLUoyy+jbXDcDrMyzxEm3Tp+mfAZCp61/AjqLOfjUjXhTA6Q3/14roE6z8MiW2S2C
BJEN62VpciE5rumnSpOnRVP3qSyxrePkLraRZ5YINSXuRc4ce2c7I1cShdmOyD7m02sZ9cqli+eR
rAxHcPllbYJknXWerQQTglalwE+2kaeiv5gquuvOxsr9tvOnSPqafne/1MYkcuy0CylHjM+eNghH
2SWkZuQtIn69RL+WXOktDqEjRixPqUBfWenLiGdbD23jUn7e5kNBaK2wddNkdkicx39KMec9Thjj
dvkBee7mxFmxRFUJFbpRJJeoNko+q+uXgVTS759NGKJvZYjKB6sqXNg1dKcu0ROac75UxBFvAOSh
O1k+6fc8BXkMsdRpb2BSWegnWIngC4aZu3x13uPp8jDN1NqefuRPCTI8OYuDHmWTPa5t7jHJ/WKG
j0gQH5FrsX7nER85gXI88xDc6N3y6RvzbnDmtCMZpUZjzz7SKAr4tH5ZDb4izlGvpaxhgnFEvhDV
KRnPCsdpq83cTMf5XydhCxPa3nAe1+PjIZ6HbiYvaxm0az+3IqQVil9MEeADPcFJw8/b0SpOqDgA
YJ9708vLsmbUEJfdjQWkmASPozu0vwT/TdpvOlnVas+QQTAHkVF57Q2zaQ+MKzmOYBGfAA/zAPAI
9wSo/q87POxGiLbNTrIq3Pw2JJMO64mvHzV4AAJ4DsT3WMM8+PTDMfcsDcruA/jUwl/MnV+gLC8i
hbgC9Bo7+n81Q+2fpYzpG7QMZiMq5/YrR2viYKyai2NVzCpaETgDFmQL6XrD/fwzG8A6ejQZUa0Z
8Wy0so1qDJQnTmUlfSAgmyUuP/DyKatiFS/C7+TYWK5kuL4cbJJ51x2r5+x1y7ZW3RdEYYotGJmG
zZsq1cZJuKQbsyQ2eVEurDw1yhPFKaBXA8/gYmXrVAXhp7aacTC64PNvFeL4uo/JTOq7af0C/nVU
86qIOnCrBRKMZgRnJCTRsyrkVsgpqzqJ/hCmNZLygyA6uIRqzcK9wGYiqDTz6qWoKcDrtVYGHg8p
iwkxDZ8stQq0tF0fRLQzEDI3ikebGDvmlrAVkFICDq7XU7rPUM9MccNSRpxJ/khy5SSKb70e+HBN
Cdsk/tqGg4sopnAQrSF2rSFg5aPVUbmUojV0JjxchaPj7GR+iIyG656801oWTNiwiqSRoFaQuv2K
/nJz8VzAwo2EwWGuGbrVH6AQKYqokctBIg7gZECWI9RM+JJAxMigxud322tjsYRojR2pLJmxnSQm
N7VvrYh05AC7tqane7USY6G2ZONrWiO5EKXvA36CKRLEJERgULkNaOuelGQ51JzM03U5z60+gRbb
ubiWVUh8qrX6F1bPfMcBD+9hdNgewXPEQAZ4oPj3v6OTiGjCa0wt/0yMd+Ha9PQ3QVcIBARBgHdX
nSPclo63yHymQjk4bi15pwCl4FiC1jpdCB9ryl6OxB/eP8DLCS9mRmIe6Q0Rfs/s2Bm4JxsbJf+E
NzLQK1DYK+8MJ5k3BIGz55UnG5ZjHwJL8dv5c73Zj2YA89oYvgW2YSHywOcCcCvS0Zp1t0oSPOo8
LzGzpDf6WfzWWehjjWX2oWqZXQTl+ltakRxheG5kJyxKgQTlcrNJCMSAaTAZM1mGOzbjP6T+TOAf
1yZP0drVPSM1DtTs7oKwVmf7NftcyQTarpMAWxSfKF5kdaqK/6GxpUlYMO0PIL9hjvgb+IE3Bgod
0XUPI9fJh7xrO9++K1idDw0B4XXyzSEvxJ4MaXpdzRXefHlbYkAyp1HyYDh8rdeozDUg8/N5Onug
sydyP4x/grtPozJ/ezRCzsJP6nbaJTHY9Y7Yto/5nCOOEBiDJ1wbp4aGuugez1JLCP0bBcLd8CeB
p1VnGXLRr8A6+hXWhfCdcBVf6Qc87c7jQSiExgUOX9Glve8FFPFsX7KutP+vLXGaS9ri+lW6Rh9u
atcEJX3Iio00PmubED3y/twlUaZBPnASjeotWMOak40JBDlW7o1g9xZlONYyCxQ+a2HdSMPIKzC2
LxAJ+8jxlrzISDo0zjpLUohjcUMGGkd+PvjVFEXcgV3dc6Vdii5WqgQTxbKsOPooifaILjPxCopE
7nDxcoHAo49FcI8TgZPbpBwS+kehB0OsquLFeiEN5T3dZKtubw1v53kLtfYV/61jN95UaJq443uB
1aMbEKQ+ulv969mt/TvCYNLRZ6yVtQJiNorpLtqrKrlN0PZ5HoBQA6lZG5TOsj49eO5ocJRNJ6hs
WV78EgF62nh2tDvjaC2lcNqz0/urb5Zlpd5DaiISMkRLpP7lcl59gXfW4HgVN7wlQMIVcgWw3PQ3
qzfcFGoNTECXO5+IfcZxwrQfgSybumYu9sIeViGXAgGmVSmKC7oM6n+KIq1N8R3j1GZ2eNK6dkwG
1hJeNkKuooRrWkzhW/qUFYDqyFQlvORONKL3ArJyWVTDT3tyYQjpS6hOEY6O/l4Gpeuqc5vzAqwn
JMF5afAVC2rH44g+4SyWTYXrbuApQ0Afjl3ILED34XYtH6l7RyIkNmj5BfwDRpHSovai1HGnZd0C
P0U8zVGj25UUgMOLDWyrv0Z5p6nTG+Ha6xO38KzRUtIUB73EB3HEwGtNt7lzG4s9hp/iEDtJBbbN
Jfg+04HfwMi8VDMBTxF9ge0sdOcxbCO/APMyLRoeMpFuDgftqjAX7dXeSc80oGNtTv8cBwvFNnta
cglPIwixZg3bmeS7oliy/hUQlG5cIr8PmZONlw+oA0RsSLo67OQ4EKKIxmr1uNAu6BaqvJn6n0bU
a/48e+aivIt+BCj6cgDp9oAisuwXM2KnuR0pL5QnKOL2/BZRy5dez49ie6uj32rNJHJtYnrtOaoK
y6H3xZ4q4FbU9FR8GhIbXzpeVEY3/zkMsMfYecFLL+Xj0n4hRh0uQMrlHYB+hZvdUBl2sAzG7JWG
7woY2E/PXooSmsqxQus2kXWOycqoetvB04wktAku0OW41gVbjxrtfr5GTNQYpn4d7JKxfIBJaPGA
BeSzxl+HclfEBXWpQRtmNOXglOL/0QM2Zky8r/VrtQzgPWbeavFJnNWMJzWJnTO/TlpvzOJsX0RX
HJlhpE5Z7UUxDcl2+lNTMr4dXMn3Rn4YgP5RptO3yucpcGFHxx8N9RE/N2amgpwj/Tm7jUB1ZABY
zDHgdmZB7fS9wpl2WAh6qEqtm3un5pAY4VtOjjQsSAM2SKUNf72yItrVM3oln4oVT1QHC/obFr9R
gsey7rJgzPUhcv/oKJog/dLwhFk7ft0HU+YPzBTqyRlxr3mEkZoz0VyPQVgW7moSY3/LBJo54tTh
aezbR8+JWd+Y/1bSNV+Uyao7rT4A7sd74RHGPuxek3Ahp2ISE+vlvTtvAHzHvs5zCiIYEH7spRxM
wK8eY5Z1YeGKpuTyqy6bPc5z8u6QCyFB9xq6KcCGx/xhwuiwyF70fkjBw7aHAP8u2GENnvAfTrXD
HMu/7kC+K9uuSC9+dEyjuIQ3x5T7n9mpXHt89TBtDZj88hLaVV9wHOOp3Osse0MGT+/UHDV+qcxc
Z4oXg0syqBslcdG3xFX2YJTyyLsV7xfvK2ZAWNUo8mQ5T2j3tUqS/SkFt7xVTcqb/v9ktdGe5xN/
i59WTjUj7RJPriP1UQ+UsMdbjgPOKkFrLnAJzPeB6PfLJQoIxDD/XNZOXe4+0cvcdmKtcw/kAdjc
RCF3qJsxjSlZLPTNtp4QvSKudDTYQ6rI6J+b0VllV2DqM068byxioa6OG/CD7f57WnnmxWdzMRwk
6ywuOhy56WEegRYXMjYXjt5IkcnmEQr7U4YkkmPSWOgKsmw0HsmCb7hACIrb9xQJLqfGjzBdtZwP
VeZ2Vi3LFbc9yID9+kIFuruMrYqlReNH9xnXjn124LodZN+L4mgslLRTYhbzNB3WhLRdsggbBv9q
5mAeHl2tOgu3NOythAT7zBmi+Oyq++SNQz83v05cTVg+PnEg/2l74UbUS/p2GHXO0C0M8z1m4QGm
uiAH4tTiRpUBjkhEv/P3rHxtCioS+EVhgkVYHOaofoR8QE+OSGX4qFbpOFW3LezcYBCTxRyH/G5E
FD63ddxHMJVXG4zc6WI/CKnAVWV0HkCTRj76Na4WWNfQMvs5iXub+CYq7BHgffQiTor/nwnZAbtz
HgoLvlrBg2R6LDGeQ0C7MB/y31iEkv70pePBoc4TpIVR+41J/+vi6pmi79Kgrk5FVDeHpu51+Vxy
3bplws0LDNtKdWLUs6k8jRs3hkEE3VwBmRCrwsenaTwX2Ixz4bc5BDsics+XjiicI8WnXFY6x+pg
WfgZF4JpN9Kc8DZw6D3GBVoIIcLt6pDtvxlSB3xr4GR/8S/7A7M0lI/NR5wlWhn7666+mzEiy6j0
rl11SWmTL+G3q1BtyNjPl5P69DZDS6BkT/h/3bmaZ2alzjYIZ13hgNdg9CDtHk6Ik4cEl5hMS8BX
XR1GhRpwb5gcfwQig9bMEMGqctbJufr7Qb3qxMFK6BFnJQ6e6rqlUX9qiyNU3ddmkuaraCE2j/Yx
pB0IUytp/yKON7Zn7qT/ZnVy6B2ZKiljMH/hcvdAPclOWR/E5sL/46STrP3oRLFeuOs/q+esVUkr
RNxQ9+5YrvvYRq6EckaHzYrZhg3bYqIN9Wpt9/oXS7DgOvRT2ne8LD0gHg8euA75X/EGfbHQ6ChD
RKCKn69pPAan8etl8AgNK7PkcJ9RhZnoewRQCeIUbvpX0U7xK3x4eATTbakKCIHfwTGfzA5Ilp7A
erEQFsBJW3+8z3wUmzABk9tTdaqwu18NjOTxv8ZsiOROh27dBrFXODlC2BtDYFBug1a8MF5ircym
3vNkl3UoRehPh5ZKl1AprYGuFAKGo5PYCIyIUrfBinAFjepoh9dlBQOi0a+g/cI4hyutnyn5ZKgw
LrF+mU4wwn5LMsQ4nrSmSkvbOi8UfEyC1HLUltJ0sGB8x0vuKkNIHHbUDp40dtIccqK3qGD9mucj
HPxxBs7BFVfixmhKydQ74CHYPA9MAX1wbMg5ox/sOXdJGOWNOErn/k4wi/t+I6COwE4syKo0MTXW
uFiHfLF3sfO/A4I2VvyDIiPMBUB0IzSIIY/W5UXYcH/lZRJrF90PSO+kPV0MAPMsTZM69/mCHrSq
atat4c6p+FWNgGVpLlPhZ/xRS/jNTrdnozd8bsmtvqNO0ocM+dvg/CrnLhQShQu6A1DS6Nuyakhm
kNVfMXkBMyJQGQNpK/cQEqgmE1Fn1N/jxPGQqMemOOrIKVpQwkBPDUuNJnJrhOkv1nLEtzNM8/cd
fhV+AddjiAnjZUkTvnO7KgZewi3ansyBUWw4rlJqf5e0/57ptk76X3QUmHAecBHTTzBrWoBPKdhz
yV8ywERofiCkmUkyfHPpK7+m/B/W8i5mNZeEn65s5Ea0E8xRnRXRhpk29+PHdT8wPUKGWbzhpl6D
1y0y2XEeCRmusOnaO+FDIziDLaBz/i8lAJ9DbR4VHOJBg+4DT5idVAsTM1PEP8QPgLpnpMRdsBaR
tP7Mr8DK+OqdUy1lDEVeC05t/GwceU8b7HISmXOe1X3cFju8xKAJUQICdz6dAlNX8U0Y8lRLLtxH
3Guy7tytat8lTb7baa71SL/KWydcfiYXeboUSEn+w/YEpnWhd9l8Gmuk/QsFZ8ct0X16FR/J9phI
y15OiNI4Jf+tRP/gSBQnzpalA6ZuGzHw0xRFS/4uJdpb4CNLiAlkLObXcvZLWuSRpbEfMdlGWbdf
jKsgZQmfiF5umKywRsxm5P4x6Uhj99PH14TkT8IcG5/otdQRbGfGMc8Y7hQ/Zm0InHZUFVNy1GNM
3IBvhIlI0pyo25DIN2Bs1h6ODm6hbhFv8uiaGlFbuoADcXDB/wfi0b/eTtuAsmyisSSMqGcNXp4j
WEpcCPGSglVJqC4a5zCPtByAjRVSeyk9Czraaw8KbTHKjxpEokCZejGY9gT81BmL0v1WokeTyyLR
0Nbv1vDn8C90Y7Hrruor9U16oTdvyFvuLHEoYQGc+8CtMJTax1pPrvy+78UY3IXPQ6aHjr9ud3dZ
rB+xy7dApvEExCDS/KC9xXq2YFYg69yF8iNVdEhXwA6vA3FLep8kQ1t+TD/B6AzJW7H4CVTlxvab
qkbt3nkF2Z4XFnbtXEyNaSKZaM3Yocq1UQO8WfK2xw14D7Z2JYMJvPolW/dBBKaUfwm4I3uuLi6v
ZxrM2PJQYIQVUzgknI12hI91wihDOVidCZ96NwlAZjQWo6JQBtunNx8mbkoPXsnif6Qwr+5eo41S
yX++VeQmEJBNh7nzVdlQbFdTZf93qCFNSrFOkuFz0/pCDLl+CYIc/tpx7nU/97j2sPHe7SAKJ9jF
5rk5GicQvDOdHpNl57up1mq/ogLGwLrl6aqye05faPsQ1btSL1FTxIK9cDzZxYX7PMe+7aAnoapZ
QJLDMBCgOZEU6iCpz7bH1cH2Rza2TkLGeA7z0zYY/jqKRYfDIkvdxeuQrGZ5EIrND4Vi6KAi8ahw
nNrOmpfogdSdV5sWuL1FyzHqpqhnZ7vgQFGAMnTCpQySRsWr+ptyoB7oNOKZ93trMtoNYTMxf4tG
RTATAT0wV95veMq5J2KTTVjigYgMkJRb36R3KRf+rjNhyzFByMckCJfocV/K7ENbe2hP4L0RLme4
uQ8IpE2hHk5e3tnu4t3STxkLeqmaG4CRF9jEavg0AyGBug7fbNYRFCo/q6xVyCSAhDmVEIxu2RxM
8TAJ0hywg0BKwWzmpxwjyUIjdqlNIznfVIISg35pIVOuPxxe0A+d55uFDKLofg/8QheKP7jUH9Y+
z1Ania7zZwno1RslH1mqc1r1LuoHe4sD40LfSGo6jzHdlgSOPiCSk0eTaiwXBcdc745A+rVtNLkn
lXr9D7OgEiAf4w8PXWmKOuRrcgdjNNRkNcuRZxUTWgSxmRBo+6MhVUpnu5meoRirN471njE8D98H
Fdrv5VDrZerMM8E0LHym6koo5bkbO3aiTLZLnq4Wz7QWIKjWChlA8KatJEXM73oEUNfVbXoPrMM+
kSYSCYSdAHuBNQynnzMibrTezm6kKegaTtOLfVvVmcBoFbyUWpawvgHpqGs1fjDiXsR8PPdRcbKk
TYF66OHb708pvY3h5EpWd2ODsMUVt/EXhYz2Q96rbGyLbh9pSi+5jHD2crUtPub4iC3ggm+T7FqU
0z+vWFRG4vCB1Vdu27Xi6aoDySU5E7yCc83bx3XUM3kfWhZKIMWd8oTHTFut8PPhZsvHEkV8cm+Z
bUAdCjC3rAtI/GbBqznckOZKBICSIrXZJM84SDJYo6V15YKMLhT/A3BHBOb6emeGfW+d6k/WZ5EX
tpmcO10LnlgmQYUJVda5uszj5t7fr27NAkwd8UfQh1DNBacPpU+Xb5Qx++AmEKXgSHnrP0rMXiUp
P9mhzCWO5EqXSlpPo5Zpj14oagkAGvkX5bCUkYaTC56dtUnu2lxI9qg+c5ODkUt0Qz14qbhCq+mJ
j3kT1JagPBvwkcc5BVZKslP1CiPt0iAQr31Gd6kexO1WPNdAQDzTX63EsIUbTJeaY9x5VMIj09EQ
h7XbfmUDXaFXybGCPLsHTEkxKUMRo+Zfwj/upY8LVXtHJ0PjUKRl2hVxtoGVM5GBklXAOrHZb3Wb
AH5FW73clOBl8U5ObOvOzN9pDifYjNjs8KE4sAA/Lu0mAanCBYcT1lIte0HRKnPwIfxLvcttOLMM
oeTVKqDnuHXbKGpOgogl547Z85aR4ZqTk64ALhJgHKWGGrfeMMXgmSy+8FQtli0xX4JXQ5U+QEiJ
see7NGS3BrHzhCCbE8mcvWRmzli87uGbJdxSrd5qoL3xF4i/IjIUTmx3Z0XrE2xRBAH4YEeVpRNE
n4ls4G/2eTA4VEXxgwLTSyycTFdaxg9ME0jcbK/V1xloK6YIoVJqkI8xOKP7FNDXSP3H/H2CN3IH
RNiEyauRrRSyI1DcWkz8UhyAZoaLGWhg5X7vyL7dPlNV757yo/VzqxqWno8Nzh6z8FYXZP8Xs8u0
dtgwavARGZtN7VzuCKnt2RyMIjlOfv/4TFGAIbbh0o9CbkQhnOwW9gQaO9082koO7uIsf9qsWmG0
igNcprqlubuIpjy7pdjoLhw13C3dCDMF84/h/PoLuXDN0Xe2IQwIEq5+mxQjwh1E0JimVGWLQcz6
phJvaaSbhEkVhnIBELdD65c0FK8LaBve2ryxQDnPNDgzmzvdmBCXtCkmecc3zejZIpjYX9A5HFdl
gPNYv8lJZIkISGLfyJo10+Ud0FlCdOHomEqB1DY9ZqtfEhriglBOonDfJTNqWlpy2kX65v5UuuhK
MC2buST8WuBHwzf3qibxyzFAvVcLHRreSiRNq4uuCud1BWDcEttnhiRy4lf1oaT8ZbnXpQsY+3/o
WiICAIuvk8LfGPc9E7d198JIEYbSJ+5P/2+AByRJebBQAWFQMvfxymt4VFOothj/Mk9d/tVd9Iye
F+ua6bTveb2WCho9OOb1leENDD8Qrdl1LSjnQYswGkqrFv/IHd8vrXWdlpnGfgAPNQHtGeLELsCJ
CpGnr56UNmTv25icUPRzC8/JGdi5neimcn2bbTnUIqSWkeWBKtcBx4BdlOUmW0exiUKpza7Z47na
bbn7xh8kfNLAHHndui5kvwFzAwPytCC/XJs7g9Uf+2JVJM/cb1h3/oMJAWkFjQ9zn2dx/VqeVGIi
vYG3ccnO1BPHoSXdu/dwaXH4in+h/ismtCcPwpCbWqmUzFIGscKV4tjlC20ZkiRm5+cBp5KfVv1m
FUeR2u07uwhC7ts8JJPFiwUrosmPHNRXBp+Zo29bU14Zos2C5KcPRYL6Kr5lKrGFx2QX6zUmcyRD
2xgUFaOI8VyFVts7vAy+cIcn98wUK5lJ0T24f5rH7x5KIMKnig9nzGdoubF4jSOStKm65OmWnsJD
UL1zJYijM79NLwS3RVWF2Rb9rnzkJmArMI5hfmAuVMjJ6egtzpdXVvPGHlpA4kTPMXC0P2xsHmxK
7/z0AdxlsiHWx4K/fn67jyCdOLAg07aTWtn+FmahViI/Aej3mMm6g8wMQs5qyZiW+dX2xwgEhHQ2
xeOtbIVJw7rvrVKgCMKPPxqJQw5jjF+YTMM9gdOk51Pk1MXffnjc5oMvS1J0eoA3n/WkACuO7dtR
MttXZ8TJ4KlU0tqt455ZHdPWcvSzn9oZZLh/EWHrF7cLz5L5i6B36GJ/ra+D3nXbbjh7J/FBy9tJ
QKX48loyiUSx2cmh01x6kbsmGv8vEewMCiLJ9GaPFAHkNVqYbtPTLfC1Qy/53fgVBe1VbNA1IPlj
pJMZ9a/7ZBdKGSpXq/k1Mt0RVugc1MmvfdfYlWcKWsfBpMbqddKYc0ni8BrmJfh13t3XDGJafWNQ
+ZDWeFAiA1SmIrvMXGDrWYCkzHATMVt/s4niZeN2OaVy3x82O2lM9XF7KweXTn2rRWgD6qwfpgXv
qT4r8kTv2f/6EFrpz+6Gq/qjj/RzmifgFW8p7nQhYpuRDpfWmOuI3JT5cb/TH4XhoYnQ7kQHc3Jg
4sfa9g7Ois3cnqkatfwmc8qtEH/D7XWTQKjoCv//HI8B3OjoCBUTz+CCF67onNxXbIK2vKO6YVdD
kHUVNhO1fCikY9BADamhh87NPvkf0YhHsRLh1O9TDz1z0u0lfrIBlyEe2YFi7yKTHYLNNhWYPG7m
H13e+kJ6uGLfGM+KkMGjjTFZL/epA+oqWLPqVTyzFrOBIcVoBbGP20GfBUkrX+W5pLa0Kdj/Phue
VBqW10ks9JNO0aM5VYO2j9QktoLHz1Y1GCE28BI72fdJjxMSIPFEyvSqWFsfFKEutt72mFkD1Lj9
3j9UwMuNr5M9BTT86h/UN02KfNT3jVR0QzwVlNusrGsxrOZvUhYGh5zOPd2p/wh2GOPrItSim5EU
9IKUnPoXfenCYQRstGHpJckhvRKoE/3UyAp5eVzfxEoOPUgL4mXHtKIGrpWoVpFhUfFVGPkFr4qg
S+9Bz8XBczY3xYQdkI/tnwlxZiQk4E8KMVp5khILlWvAj60tJSBTEcpule9JZBkjLHHJJUskXHEI
eqwIK8HFSPpayGgREoPxWS7EfmWBHEb0fF0F0OePPtjwJr341X8X0r/644Filn7yjvAN7By42Mji
knViEzFfVtOreW8VrhuplsOr3WH0s6XR8IhPJneRQWwNkN/0/XpXOGhzrH/1qxgGYiia5pB2sr6x
d1geJzOqMwU7UyAmmObQoiQ51MqmQVIm7Ai4N0ehrEkgkfTFDaAcuPu7ZPk8WsxO4qtS/Ri0EL7r
Zj0fDh9a7yjXtcc6YyD8kx3flPLn0fyNGtjuYY6OQr5u6kFISbTroIiMSP/kDScExAYYXG1O4zIx
AQKkA0CwTDDb68m+AjDNx03XNgKqvCSi30k/DWN2o3IksUUjTybLTsJWVxQ3VPYyjrVqECJZOFnU
NmTfxaT4eQaPdOM13Ts97F8vabWQ7E6C9ctS/g6EXmyrNNrI5PE7PrDzSlPLssJOZmWcPHIK7CSx
LsPP2FqKQgDlaiY2ZR0/Wkxe8K7wIrX9yBmVcnkXcg2oOLdhcew1fSkmIE1ssYq3Pdwvv/HJmD/h
Mw9wZZBATBvTH0Y0s3Iqvkg09kh7z4qSJVOmHNdPSWD5UnRRf6xi2A0R8ZhHG8zKuXIXASEhBSYr
moy8iyWM//8KQ2+D4kDQLdifMEaJ1ru2THSKGXyeUFhlD9O2uQbqHnR96kvADvBcRdNtjZyN32UE
LtuYYBx2ah1lbcdbNoRjkwPMOIyL7Y4Tr3E97vTVI5HSFkNv06IaM+cLcHOLBShUJDMlWWmsseHN
KdYHaWCRtKayyxWh/XULspKCluPQoj03N7O5qkdibP3t8Cb1KQkdQvwfqMt/p2pfby6oZrEe3rJu
VEfHnT5+UIihx1eXgJNQgevmPBIqRnxpUuBupmMc5Kg0inBLO498VlLv7nnKebQrbbJio8zrcDb3
sX1g8CksEwn53YubeytsKGuzS4M+NGwT2l6pxUYudwg8ZDTyxwOOE1mCoBrcx3VrxOAu/V1zOUN5
uSn8txTwTj/yitAPWtKLA/3JDyRMZZnlCHbrlqTSLZrsy99L0Z/KeVKS+6d4G0Zrnn5QNsPhU7DN
K9qDwYyudqHQTtozj333Z9vf6qz2DjV59MR2oDV7aCXBQYfIdjsfVZhDHngeOgErDV1K3LlQCMJS
EtTRo0zCFK7qqJ/g6k8Jifmodvvq2IhURMBFjfrWcFic65pwREoK3jUmHcT4IwwXT9+wl2jKDc3p
DD/GB37U/efq3OzOLwpnpHNg4MeZhXRSFhj0vq0trMB6X26sDMmQsIclAB+tTKMP3OXGixZ1VxpF
VhPK27cXZeNtxoXr8xt76kTOPz3a+IrfsZWK0NTSVKsgEz1JVtRHtbPVTKCZb8DsFyZg7GONK4lf
OKY3iKtR0XFIAP8kDvmda59+S/hj2bkdu8zQM53NhCJJjT4rFy5ZZffKY5r4aPQ8iC2oDMlbOIfV
eCn5ZI03C5G4Gq256vmJmJ6sQxKULbWUu2FoJS0+0SRxlvzoN48M5KWmQUfywEE644XrK1csvDHL
2VH0SxUtCTOqvVi/xNOg6iL/S48aSbFFO3rLGpF1bnHiW7MO7Ctczg3vLbp7HwVOI7Bg0aZR567k
h7+jAb8bGDL7/kQgOD+P14vyeIU54cE2k2jn+T0wH34l4IjfjLZ6eFWkmpxIv6/XnKzyCIHIXrj4
1YMIesvwFYN2VxS0lpfzItxsNWs7Q6+TzsIn/9Mxvj2Z7EcKAxvzzETO/lqbdruWRPkX/7Nz//9g
QqZCCHMzVopk+szUlD8aHzaVEfBY2zUIWu60dvK4CNTb9qr8bAHTKaBrQk2RgDecyQgfXqCu07Nv
XGMNzD02HS/wtsnI/u6cd/wfSyqWCHcsUIlLhKkie38aeoZRdZ7lYfP7jfeFZpLJDxyPDfyzt9Sh
AEIc2DVC8gpfI+GZ9o91btll8S9tWbzlaFeM+DSlbtZiWK7j2rK9Jw+qgBAYr+LFEMu7lx0gyv1o
0I+E8gXw6RdzVHAJcqFnsEGy4eYU0OAPwM/HUX2b90BF1oTZD1kNe9G2zMnhjsca5OktSh+rodPb
3BabTUsjOS+6BG2NJiRL0e9n16nLVdTS3Qqpecn7QUkQKo+NtJK+bacU7N1zrF02G3ZZQXklD2I9
9xm6oMbq4LXop/diNYn2u5ooRbM0Z5VJEeKp6DT5443PPm0b7Hmv7/i5l8fYQUsiUOsJjHpjBgVG
3o7o5m4n2cgiKHG/va2gnPFUNE1q0OmbhBJoWOAps/fAGoyIDpIYXrT+7KONaPrt9Lg4lru+0Zr3
AOJ4TMOi5XcU3z0AxSdgW6xt8GWCLqZdvQGRRhYGMbYobBC9jaFIvRzGlOBrHTARX5py0YgQ1Jwo
tFanf/YYc7j41pYumXcKEWJ5cN4uiZSa+g6DyVRc5fAtk1ZvF+/JIbB3A3pdQILqQChrdUOQbXaW
L8JjIRjM1R45t+U009385yngcmgquWENbkojqkDbTWP6cYaSvfHQCUAI4MRmufUELC8JIL27mHRP
0Ktgn/oE6DKe9A+Fo0Fr2rEIDlw5T7f5nnDScN0HtHZqqEsjsx5m+E8uQXEM+BEAxPYcyT3a3GSy
FmR/+AdIqW72H6Ztlrv72nxD/kHQNe6gaO51uOJiScHbL6QGM4lTTvjEGh6EhQyRZh8XJ+IHd/eO
FEDWXHPuotVgw8d+M8I8OoINZp5qqxAcjqea9Y4r1b0EGfLbySUvzMxec6bMRybkNEto56k5gThB
fWsVgkU3HZ7sOiBpwdhM7GWRTS93/gr/nEVM8F3Src6mq1fSO+6/DCQ1Co4YWiADQUc+TsglV5gp
y2/PNEb8VBWz9wFlcbo7b76V8q+LooG7SQbRwFhi7GfIUE8oZDkYGd3jUzm6GenWYnNQCfwSXNTP
2fk7SWrmqHasn6z06Bn2onbd2dQCBGnIhnyYXzFZcCjvlAAKkPACXPsZPLrzLNqBCgy74rNsR8p4
H/xkBrI6T4iHsF82Zm3EGtmwpviMy4ZrQ4dibtJyhtlfKGSV/s959ZpMKvW6JfOkbtgbQLm1j9VL
KxNAv4nKbsbUL/HspbYHVix5WxUM6+lN/xvR8Xoo+SwjfT0AeV2WWUzyCFD6KHOa640EAEZkHyJW
9wKlSYUttqwbGRHTEq3NNbqW9AOY/QNukVuD0Moe8gucfhosPMl35WIRg0gXbxk7inw5jWqkq/Xq
TMByidTDqsmNzVV0s+JMARTMDlcROiA2Ye3vhJbqcy+S7NQbUHdLN1daqASz5MX/e+EgAJQMNpLs
Hbpq5hEF+WqMcjQ5w9c8W7X3ibbWyICZ6LjUq7s3y0GDIWxV/VyumXKcuThHJEPm//RRREfd+XS1
bwXl0vwyMuyPEPf3u5KEDuke9l9LggFS1x/IsTd/nl+HVPu+ZCT5BfOh759fcISSA2ju90vGTFZ5
vFXXPL7z5++oynPEbubhN2lCA8+iPVcqzfhqhRNvJT6RPjThMK+bU//jjzqer3uqy9F3bl0qXF1a
nRV1LZGL51L25uI2EFf9aqojBzhDJv2fLiF23l1X5XV/ywIvNcXfx5JYnQs9cPx54o0jJ8gqA2i+
kVkiR5RcrBhCf7HqfWqAEqE4mwbd2tO6Na+ndC6V9I2hwKE9NgHvFatFZdMIEpPcuBQWN8xhW6xe
aTE50n6otPL/yr46OFdW/Tjrt6MEHAH36W/9CFo2OztikK0FuVjjgm8VfeerfxIV8XTx90DxHuzt
ApoWK96+GPXVXmpIr8xKViZfg+cfn3MEvi+Kw4lUvVG7UiW9Dgmub38/+sXt305LS6AsNRqLqGHr
zNEVlZMyb9OleTo4IXSgERYdWvfZ6N29j1yilL7vBwy4W6PLsH6Vr++jbnl1sDi2n/S+G6rVpYzk
dMoYv7Nt5vIB/t7cTEp8+nzNSzOYbRjuu+9YpfrHjOF7ApdPPb8u+AHGK3Id6KCtgM+WO2QjFHw+
SylQTyV6K6+MBpvGayKINYpdE/fm5KSMEUAc4DfbzdPsOgw2PG1kLsitqvF1+vF++uzaJfzEAhho
Vm2JqL+9mGTVh1CwKpL32JHERebOimI6n6yquyCCd4Jp8eY7/7nfjwoCdZUW7ubktQfKDwNISFJZ
kMTOGeX3b7fMtu2EjuroSEKjf1UOgrR99sDlfpdPPS38x8g25qb8LPXIRQk8wNnq93ofcveMJ99k
/s1PBgbQR+uIxXzSc1UryrWvftMc8/b/UKdXii98IzW5Jv+hD9f47zZ8kQTIIFQNxnRE4LaSH1Fm
Vm8qRC0bph1Lz2eqcq3TXwbz3M5/YkEUq5jDcmxEcHWr38njNx4uieeq0mSOQsDaig+u0I2TqyjD
3rZdHwKAjns8eW41ik2XRrCPpDnd+xC9DU32VHyoYnwf5xDz9zhQyuuN7G3UtnxqkGgDm3fTPQV0
4JWhRnfifBGYf+2RmqxMtAaJ4Ydvo8RNCXmj1HUKXmd4qpWSXSxz2gWWDl17dtam1QrVvfbuKDkt
NI4Jn29cabqSUwOkxhHHTbMZsRsNNDQrrsbkKa7Qe+zzcz6xiv4xvR4jMubk8aresa5gizS4p3r8
hnRndeDbw+IDPbdMNzbWiRYucp/w+EehV91iZLEJd/zSEi37rM2b6qfdx9jF3g8I4U6fnzGuwoq2
jPUb+s2BzRen/tgkOCXd6u6sH9in9RvPKuhWuus+cI7dMFlR7xVhWMeZBYfgIiQ1DT4AJSKS+HZM
KNxXnHyWDu5o6f70thC8kjticc3AI7dxQWvslE5VXPYjwHEqV3oslK9CZXUM2kY7gjI4bG+ssFyX
ZSZxf8uAdbMq2gYcoZbrzRf/HylDlH/QVZWHa2b4QDRvJxzdJEuNKKSBxqtYFqYTlbkr/8HlY6rR
gD8V7eiJH2E7ti9BBTPDHpmI+4/bV9je2tl9Mg1ACTfwKO++a4SOSbxqf7YRrCN3hwdooiVnazRH
xqfEXQy2Tbx2x69AdQOJSyNB93uSZgjW2cI8Y8UUZBZv8DU3KKYs7yJpKk9fM0ZIbRsoPZEMHaCo
5eHAEdmytyz/r2a9DPJiohhJ5HRXO0dA1dYf5bhlHW9j6BevGXtcoInLJ4vubk4/MYPpShg23u+4
mrLui80wPeMB9nlnXFyuXZ9VNdWE6Yglu+sPY8vVq4wL+eU/WRnk+jqAqH4ghhTbjrYxDjJBysvZ
eZw1Z3RZg9mI7B1x1PZ/StNCkkhWSQ/UkJZbcokd4pm2i8YO+GUpGILtlwqjdoyTNluOkpFgwfCH
68CtgWH/OaDGlw1rX8zv7+OpPMGh47aAdcFN5dHUGeGn7QXxMg8SWP5wBO7us39GJJzMk+bpt3/C
TFLbR7pNLR9KZXJ+TB0zgGkUEFizLXjOv6Tn7p420uPWEBXKpRJ4Cm2++SRoOk0GiW4cMPxv5xsp
g9Wg+zwKd5L3hytZQfsmLISxUuBgyCiZFJ+qdApi/CIfrUoWxStxylGXamDNUmHh8FuF3jAPlN9c
DhEcbvEO2q185GhoRFeOJ4bqjdF0GAs4WIQ2sETYM4136uoB6ng8Nlmj3DLFZdALdIHkun2tWUAk
JNiYoKxXwhfhOwMkRjpbuBq3iBDBwzxfROkKVgp0HVFBccKXRrj0BaqEp6Gf9OsvMy/q9YxYee3V
UGXokXL21UPUN7fhDRbLJql1cGKib0GSIGIfLCTaOp1SC760GmN21/YcFiS16y2hfWiMrmWV25sK
FOmmXj+GmS0b15wnueAza09N+u5WqFZ+JSGwD0zTXQTdeBjvtuZy7otz0AFt0MqHvIgeMiphTXX2
uT8J7F1Y/3RSXMks/nsSaL29mxauzjgAd3UjxrHAyWwcXca1T5Lkg8eMila7YiX7ujlb3KbOn/4u
tGVUX0I5gEpXJhJ4A2fFjU7zZUwKlz0EI/pWFpTVzq1Zk4bINw++KOrYN6Y1P2X0Pz/HuUAYAxZ7
fNqAVJOZJk/s3az6+gxTOUGXK6tiu9k2FlG9BeT0bEL+6gZZc01hC8qA0KOR8vmjfaNba95eys8v
PRT/zYyH07pYgDIOyt+KOgZCqkSbEnz3IH963Q9S3dNG8BCT1EsGLW69cblZy65nzOpCcgZCD39o
7fFD+7hRzIKVFwcqpOFfI5nAPBIueHYm2skw27kVc11zxx8qZOfgytVMtrk+lTz93L1yWhkHe71S
WCfPdueHCZQvD5k+dNGkfaLGbKYjDGf0HiEy7Nx4CeErl4muFEOOeHSlziY6uQMOkbFktjihzp89
rrXJcFfuRQvRI7+lymQtxZRinTxZUcj6R7e+oeeWVKyCHiyUwO74Aeqj2YLRM+TiKPVl72q3fw46
oaXotN+hDaYe2Mrk4j2oK7shaOXTyflK4h9xlN49lKZb+Fi6e/AaoD2MuryN7SqcRFXlaH+FDHJr
5bEuGjXL3AripLLUxc+K3+IotWcYhZYuvlJoX73CyUAMWu9gvDruv4C5P+g5ownGvDT/xMVR4yzz
GBSiIExiEjX8qobuzkWu7ilEiP2dD+mxxF5wHYuROX1nZnGbIdgkVQd1w1LJ8GLN5bx/OxwIC6zz
Yp31S+zXoMWO+6nsdGNM1YS/ScpiVIFWJOVOFvIjuHv/EXVOZf/k5i072U78EXXCNsTU7uhjTy2c
AgXQpqI716rzyKv3SLVkX5kDoLZtErE2NefqJsCxdRrWd5589jy4at09s5xtdoXGvVmzcPXp/TCP
e354Q3TVcXjlVz1iKD3sLINL16wb8PKPYOYC23qgRe5RgR8gOJhVaZdco6V6Dp8y0uECW2U2RR8z
wwa7Y9fk6SAM485/4sUL1qH4U+DRkQfXpMGYqg304ssoxJY1kPXwOU2hfLGyJvpRZ8uL42mVyR0m
bcVaG3orJur5BwYqRWWVxkEviw2FPdLW3gVeUNAZyXN50EAhbLWy0584JwrkpWBlYdcw+xbSxGLo
yNnr4umDDypr5ajPm2jaRYxDtr91Mln2s/av0+0U+BtIZIYes5YSVbfqX7w2fnT5SVSMSUUCbw+y
4SquO2ku+t61EAEjXpQIBLN2vC5i0lLIHivWFMa2/HhHbwwDptNockDnEvkiu62fTMM0yhnFRxxp
y56psZogfPYV7koJdwNtRQ+FDeTt2YkT9GnLeqbbd2EKVQNE4J8ro19kjohZ5Ig3ws3sAT8KyGcu
ufoFbkujFJB2naZS22Q5Btx+JAJFW6xnOAoQpo9G6pRguVw8HHSzKboYjFlM9puJ15wJii3ZxPA0
Okbs00e43a+RnI7MJuh+hBlTRgjBQOwE3D1cKHe9ztv0mKNj1uroY6hxhi8XJHkzXmIRwxoQL02R
zJHmWs81O05bYQuHnAGuWZY5PT5h9EFajHeEKCGsHrmZ4pCGJQ0DqjgV8WewrHMfpfOamrTE6/fI
jWiX5Yhm3mpii4os6cvLOx0o/jiDW7kayMAFQg6AZhCVq/xfoHy2xGgVIkSLymTl+piHQIBXnkO/
WxomC2VAUrRU6cNI0/e/NETNUjHQMsBIPtdVVxbz95bH2F2meFvudSdOdBofs9hKELkQuKV4SVcn
udcmWYYnXVN1tPRXwaGcLv1Eoz49PCmc4M0yfivD+zf1FAy2F2i19HuIAEKijg424/h16sMNSgu9
GdMwXBifGUfz6o23MpvAbLoK2du3cFfyNQVHAQ+1iNmsW203hUlFa4BA3XYT4VYwVnP0fdTtdvlk
wYjGEQLop85d1AGeFSFRAyRgIbQxSkXIlcStFDGiEcRvMhD9jJS0CJERW3+/zW5NOM5CL1vhZgmB
5lNq3ukhOg7vsLh+GkBR/ShBG8LbLi+e+ty2M6fifXv0a9ojpTyPIiONv/zywe1+mN+49OhMG9+O
XQts3laGBSLcElVu0u1eMaK5oWkE+/mFJxJOKPCtJjJ8dZxwahoiLN4vEB8oNL7CsoQt6q9OyXUQ
iOvFzhGiKsGGQvlmRFUmCQ+G7dhPu5cLnrtXb1s2n8sU6+/oXjaopBc6TVm2esdJ5U4hLDrRo49h
xbABGkvzEPpQxDE/ESy+FquvTdB4bJ3l9zpcysoXMBX+JxCMDrZv/xloH7YSoIHhso7ZUzuOQKua
1CUPzC46Dd5YROa4LqARjqRlO1ATI5r1D9PosMea5y/YaC2uFONMEz65IYhoDv/ekG9HwGAkywoQ
pdTAXVgwU4ReaiNfdKboSRH9Gw85OfyBMF7QPGHG0LXYzAFjtOoMhm6W95VPAhq0R+QEIIPINZCW
D+UPW/ztNEAN1nyP0dajTWLlzJfhFI0ektmNEbp+sAKedzDZvcjTo+oPakazzmDo70ESQ1QGH3jk
sbZ8pQuduESTLNNw4JFY2GsnPRK01pU0V7Ui5cbRkjbOE9pFX79qFMnAMuN68z0S5V3T0UVigy78
s36Uk353bVvR7lxIfuGbCEoKVxJMwGv4B2infbYFlqR43T18UbJQOnss01y4k6o9XwGGstR/zDOH
gCspWQI9cX7wF6CwED4VIGZMdq4DsVUGpTtcKeZoRtkILDWGhLmGvE1hWyJEBGEJ+0hVbOloGL1P
n+5Aq2MDu6qd8Q2lLHcLPeIKIgI+YUET4qlNFU92kU4f6ezbRb4m6UB82xJmeslW/u7RB0O09J4V
V4pG4RYNmLiGUOKsdsJv9fLsKoVtgj7nYCosgV44a/MnO6QZMDjceoTcXNac3j/gmcOfiWDTvmIA
MjotAr5jroTZlfWKLG/mM7Sb/cJGPxfdY7XRhPv1/C7WNZlmuDVh5N+YL4z4YwKy/2R6gnsvP3VA
QIeNfn7+ihuQ29ItIocbkViyfHG6/HMkn/EfdEQPaux65BrJ0oENKdvHM242Wd18urN5HkPy/hea
pFpPa25r2tc24LeV+umsV6Yax4i5+rLWZsDWuwesTY8CPKk3uOThdTTN+585JQP4VMpw+WApLaLo
kdh9f3Zda52rEUAcymQkkP+P6XUJog7FCHV4+wW/2ttiQRunKr+KSDo/QA4g9qXaaJpybbb4/DIc
j2m1BDoSrWM/WMWyRKTLcoe5tH9ELIcvMiMo4PHTYel2WIUdRuwQLdtOIh8871iJ7hnmw3PVIjjd
9mEG/u4JyPtbaP/Nx/Ggzgytzl5E8gFgXStCHT2VPuKTfYfduuffIp4EEjNo0m7/AknDE0cPiWMU
q7yGOrtZhKBBi15bM75ajyVT3/18q4QVHfg75zZNw8ekVV3P20IohBGp0JeFDhbIEgZBvS1qg+PN
jAgvC33hm+oOWrZRqvb7DBq36sIaNNbZdEolm5Eac6MjJudobrAdfjVE8ok3HTkZ2B2w5W6dnjrp
8r3jLApoSuCOUeI8zieYCTFLeYhLJzQEH9fQHc4N/jcnBynblLfLIv0TU506VrDDeZvpSXE/73zr
pW6MktzA1Ok/RJo5jDx6kXrVZtjzJyuJpOu+45o84Kfb3+wBWaIbWStEhrpyeFmYi6uQSpwUQUPz
SPGZDvJQFJPpvGFKVR7FdR+wD5EPe5qRSsehBuubiFi9aUBxhn3UvK5EAT+OjGtAjInML0z5huAD
GEj96xR8+bmSNmeiuF5z5liiIRJM5mrb+AiwhDIxuQvDq9UKCdpPpx0NaBBgynH41S+O2jqeiH75
JqUtJ4RcSrHT8F7nuCQH9/zbHBx50thhDz+dRwmNRr2wYAPcD/BVhvilIfR3koWr02GkBDDZc5Bc
VEEjV3jP7udfW8GIk90bGN13KrgCqpUQKLKcs5Cb7Bb3TpzVH/DV30GE5Ppv30AQdUD69Q0dN7yJ
5DWS4RhwZjWVeclby2eMPZZqt8cyOqq9M38lzspakNH0lA+LfwxendBZR3jwOZ26NCPjpbhMY9av
Ci0VIKqatw3+aaxxi1isjMBHz7WiY+D+hUzzjwOL4Y4o1jRBGx9dIB0xCviV9ebWUpu/8t5/tj0b
ONAyZvzADcqt5x8Ch5iunv+sxQLNCD0bO9KPq4/Y8TSwA1n0Sggf8zCXfLpL3VXBCWTESFM5wS7d
1rLn/1FgHX+bJwmBK6rucIViOwdQ19G24ykLZieiE84NX6ZGZlqzqL4XvDWqW0JKoECjSKEFaocK
Meud+upFfiuS9rEcJLPn911Bdgz1SNIBwnXKfkNwWXR0IyWzUVCi2NQoINfFiLjZ78LN7flmyLVS
AI+VSMIvAxmgsDi/tSqndWZGi76iNxUgsVNHYw2k5JWHRkFexrgJgTcXvKxs0W2mzR3nD0D72Oyk
zrWqjKcWYwTk2aHgD5hQM7S9k5lPJ4Cv8UMZtObSMsXX0CzhFe2Nqq52qySdWYFbVIAXSucDDK9J
F1OOWUtumTHj+Pv18melpeqq+WoogjsF9CrcsAdimeAFxWb+VMGsgKPNbwOtWrAyFidBRbOQmh7j
IU7q5WvrR3Z/oAryOw4KbnMenLGcIjvdwiZUqQL05KKTyWBYijtEHz2QiVv4SG8v3766yUg/HyDR
rClhVgJOlSgdjGlwOjM6feDsiHyenfdf9r8J4GZylsIpj+3LoIdbZf1As3usqMnXD8TVo7YXh6mJ
tuk8Eo2Jk8NW6TCIs6gyDcXQyEaQUxYD356JQoHxp0AGGylaPzbZ2S2XBmToHVfu7U9lQIR+jsqF
lsZIapOjesBrF/nCcd5ymNAv/tzaAE8eQcp4VoyZar8+03PGdvZiJXxGDNWZH0AEU3+NawSL60ml
Rlth0XSeky2CUmgkV23IQqUki0ByMbEKa6uYavGKd6ReJfaJmsyW/UuCsWzDZTb05oq2NTNeksbZ
zh0+ToaBRIZ4NvCSAqqItObwWe9yQjckZ7GKFXYPh99DD30mPFJX48yeXtS9dKRCt8zSVxGHNO9e
+uY2FSR3mzC/1blN5A78xYZ+hiPpl0FtpTTox1Pxdt9Y/Yv8FhvSfFsKUvNZ/RossltdI8jSXXeK
RzSCIvIuJX9IwWin7xN0TMacHKZccSlWX5QNW8g+qzUjkwcig+2erk7SzgaxDzlaY4uTws+7MIto
QZE144qghgEi9THwsGSfMmVloZpZYY5JgL1Uvs/iF9F6Be2ldvLIIohNP1KliXBC2OxzeXuUsgce
4WNSXUnldK/zOfkvus2a/qnbL1hUfcCYaFzW/MBO+zqnIrhExiJusWxeBED+PqbhWTdRDjx7WEkb
Kao6BDMLBaTjW5GHnSLXC9J/n+8QiE0pn5wJLcl6/caVr6XSo2YHGtxKIkuG+0xKKhySwgA+ZetA
Kyf9E9NhLIYUEsZ5HKIu1K1OhwKV/7gPk534VwkVGFs7xNiyXHSCTJQNDYAEYoW/03iHtJvuWobR
EUU1Ysn++mAUr9veaCvaHDEJ0Ihwz47v8tFPWbX3ixb5f+mMjZfT8PJgIKRMhIiOQmKJkWVW2HhB
K8BTisaSmXXETsuu1C+MenGbXmOE55hfof5wvyVHJ1zDfmya2NV6b1LpJ4FH18J38Vap30jSC3Lu
MXjONKbUL2Zu7OXeDVxLZ03UKU8kL+iLEks3XNt+uT+WNbw6yIZTQgkU8j/CcNvE+eNr+uWTye4h
Mx4irWrVwcq58DyWD3qCG0hna9W9PnJW1UMuP7UnR47/TugorcKWifvbsISq+izk40NjfE12ZKpZ
l4pdc575G4YeWB6c5oo/T4qmt5oVZ3cO/YscPtCNvOna6eURIRakJwWJTk6cJlUGaIZrF+2kd5RG
/NuwHwzsLW/aHzn2KciG4IhIFljST3Mb9CxV6U9gEeRPxVTmys+zxEsf9MITIn4boU4w5nowcz2x
axPC+rSll2WqIKkWi4pSLVUFiyvy3qeTENx/L8zC4rbFHY61WcSxXlsmyiLq2RESq03PzzTie4EO
UQ+tQ8jOyijKVQtDa3LBp73evNxa4JXXWFta6KWlWjKP2zeFZrOKBdFHKEG5VENeAs73W0Jh3Mtx
odyAT3z7jhc5gdcbiVnDkkJIVPVR+FTQjt4ZxQcHl1b/RInQHVpl6jKP5atlWEujWEQKNj1SnhFk
AKkrA130CyS0R/bNGqjyG5P020zeoxnsgQa3xv773MFGXw0gKGeLfM1TOHrCSPz/vl6pBe+HKvLc
RK6VHxowJRyw1vr3b2377XKmA2pqK1udAY2O8WVMZgl2/bI3/MW3zIPJO7INoBshsxTePjWHioGC
c/FkYKQ1kR+yAFHX6NxxBD4znFAJMwQhX4wAEbetrrAxTa5hSxId7OF9/wGGpGP6EaVUeAnTc/Hi
YgkQzgzByVod+UIJtPHesS9ddfI6/fWirjtbPpy5sPwnaUWYwRufErultxgLkWOLjLs7Sd8YT11d
nOwzRq7YQsf14WVq4tMawy4kvZiqASH1oraPZKwEsG6wWYwnVimUZnPVrMgy0DBHtzI19tuQgCfg
8jJbJMi+iN8qTn0yt+brSq4dzuXh9ufniRFWRbSDusZOBLMdZ89Ys0O/B0+D1Ld0nNcpjd7HoAPH
zWYY9g2U7MHv4JvwvW+2qeCu8O/WC9I+sb37elDIqomZpgtiW6AruWp61cQ+/BGCott5HvmkCpKM
SGmv51sXmZt2lyrugy0eSi5IMKiwi8YQifLLqy7fIQL75V99TRP09Sd/AFnMACPy3NOHb9k08dXJ
NY6SPqEuKGdpJbAaUC0g/tCCnRNYr3rq746PPuQ1iqTABo6TJNNK1waBpSVpT3b1kj73F5ElUEVo
EZ2jyO24oGfMb9CNjmUXGmCcQ8dsecOL5oU48FRo6o2REzikpJULuXfVS4WJ9a7YaTIZ1ph8H26A
T2jDw5qZ/RuGzLFp+IY6IBuUadNZ64t437v9qymrYwBb0cRR303K3r3NKOs3a1ML+5Y63uBog60c
5NxDjl3fm03CGMtqYpXfE9oK9wnU7hu/yTkfPFUVwAVQ0ar4bscy+OSjWlhOoLEUyRy0S/EmCFXE
xtRIkKa1dA3Oj+oJxz2rMGi4C6w+lVb5CQ1N+njedKaBek19n1xtW7yXyG4Gs1mBHVuSYX/xvrnF
tPjnIRAHnmctzLMlUNMfeK7PrG3irhr22pnkJ9u6mcwi8bNf4iiCiXBCxbaZ4TV3a7Narb8Az3Td
DakWKPTgw8dsDnY6YOd9/a/07vdq1lE2Tflk7weT9QP2RkBcIHsAmrqWz6oYFiOHxDoB/GdIerF8
rC7ZhTFhpEmv/AXW3VHm3NAU6uQHJYI2guA4QbRm1hbBnOb0mH+sEpsuaV7TXbTzfQHxwFzbGDc9
JYYfguUrUXEQq4ogdhpYscBvZtPXQYcgVmIlnWIYH4KiPeRZrVfCrDwfL2VbkfcVmOB5AYyTzgJu
cyFeT6BtB5LOKxeVB0beKGGE/VjXUmedsVcJTYt4bWxSQ96H/zcjky3XIz/ozyd4e8To2k0srWdo
q5/5UMw6qUXN1EF4A42cYJYz0mmyRuUsOGub2EO4oWwQVFyhQnQ4hxKgvc7bbFuQSU8PXCV7HKCr
n91GxxGRLx6VwbzqHdPJxr+TnRPJepEn1PexA3/2y1Vj3OsBqi/q292LFX8ESeGF6oXmQR9Drayx
rNBGnEyDSXbYnse3FjJBXDmFfPi5jHDW1vfTud1WIGyJK89gDOE01auFPKuMscOyYKbLkVNnwNLS
a5AioyEeVefuXtHs2vhGmPPFov+vLw7xidoyZItVUhWOTWNPU1qjZVCzK1GmGdzdVPkIITSSRSJH
dckWxz22ughKCSqnS9wnICdGTDMlMQa+LwnnOJ7WOznWMDzFUXSaRKZKcuoZnlj3qUt7il+DV/RK
+4LFV6l/S/6OPyQX43AnVE8xmQTs+oVViFk0yZSxSbnloEQk0rfZWMi7bD0WDoXaBitF/wFtbqkH
dxj+2qlUhbqHj4YszmkdPhgH4SEA3t0HFAg4AJpOxvTuezvQIm+GRvZLkt5zdZapZ9Jlekl0zQdu
PfwL4/3scL235eScGrk+WRxut/rV0H1Emy34O9DN2hJE+6pJXP1tbx/7M3w0JQTn+nn215evBCGn
JnJY4x7gXHQWEC63+SJKTiz78VaWCCHFZBQ36S4HMEhdfSeBVonTteOJ5g1GmStuOM0KWlIJuEzZ
V/Ci5gPJobA6za6R8lKH6OCI3K56+O2fhgs8aTlqdbsLq4KZsRWlWzhPNfUorrPaJXqs8sGUu8AO
HllNbm0TGIw2aRw8f9KuZHdblWYMRlerOxQkgBXVwgTvx2OuPqe/AIyfn1V8uuKAZotMxRguLXT+
jhoe0pQhUhckDMZjJN6GmYejMdXjF98OJcMPesVAglr6xv5MqEXbVeqGCOR+XZHXJdY1mxCSOXQ4
PcyrpaT8hEwR/ID28MQ/4xbZIq6UgcdLGckeR1dTWm05cxpCvcsiC3XwqCd4SQae4U73sARbm1Px
jcAUYerWaDeKWndIbjYvjj+wNuhmMPmQXENRMvipet8zb8MFfk6M7hofqM3xd1pRPdO6zIFQc455
EDBDGhKV4s7Shhzcm2JpmFHD/dgSyHyza3rPmCCZBYqWBCM0lZp3Z0QYFkMA1KbFcrR+QxWa+0wQ
fVqmfDTtS+c/1gZfoEkqNtgCE0mmnpjF83Je5VVR6SuR0zxh6nlJExZjdYYArjas3/e67B0ldEMH
EOldarkfIiM6TIlKUPAVFLJpAgjBsFhWpYfwZKApbP24nDCMloaJGloP+3B6eGmOMxHG79BgbvuS
Xi+wBJZuSPplJ0r3liCMbhqxjbVr+jQNrhqHeIZIskrGzD6HIHBoT2fxG9ksI4SNQNDqDL14NPIH
5OtBO84sVLcjpC3TffAdXufEevi5Z5j+90+J/5otRqovvpVpI5FO06uzN3njE2Aw4al+JNA5UTH/
CVlIxGxsStP5YjFENG/TErYIuecfDC6MmtEfNFOZGbc9RnJjWfI6ipnN1XhLC3mq7ZqT98OPrXcm
bhJxVl7PwxG+u35C2JRCKhHh0ex2q0YD7xOaeFRPbtkvgthfs1BbakBKWm4eRDp63ZJe23j5u1Fy
Qdj+ATq8qR9AqmHJ5qHQN3sO0ypKwbMIALI6U4XehVTMx6u6ifsebt76BC9voHlbQBhG6BAnK3Il
mwVgJCbNOcFZTg9XZeanyahxDMCqf2j+x6x8bWxpHWZoolgq3/R3HBxT5CRK/Aacnr4tyfs9k0/D
pbFaVPpCg83NphaxSSNo493IMcrAbtEnWry0yLaevhSER6IydbcDsGWCAtegFIs64auqYYZv9uUJ
CjdDLzOk8PUFcbUZLPbyFgT6Os4k0degMjKhAgLBVfHnSF/jW2ehmKOS+/hGS52sDihdRRLwxtNZ
uPeCN+30/Zi05G7zWmzoi+4o6gaDHgee4P1wYMXQLEz71MD6RAQYEg6j9IBjWEqrdBJeBTjNmPXA
7Nek5FFav2zr+Is+Zg81Z8xPjerMGD78mpx5XjCD7GVYl4VoEyf1o6BxXroYf1047nEizUt1mKOE
XChucpy6Ov6YRYykecr0v6evezc9LJpwA0xWvdo4JVnrJoE7SHN6NbeZA71N2tDy74R5yg2McEVH
Psf5iAChod0lVQC8U68rM6uGIMFQMSDYQAkM5yuzIFGm6RNTZnlD1L9JxiY92eSPFj+bzwWWrE5C
dQthyyIeW4W2Mu42k9EbHA45vGS7eQA0o7JQYBbu1bHuhnwPXfDKu4sujUdyVq8N3j69lzranIBQ
lVq/SUyalzR3AYkd/IpPEFbkHqG4s5sGNfYAsp09ks9+6c+uqE0wLUJsR+KavqL4YfwJKjOSFJTc
XhZyJm328fiZ7TF62fagZk9p/8SFmfd54MYhDyqPtuSq4ttpG3dOvzdj2bHdTvP76+N3gwI8yq5t
lnYaj1zrm5ofa+TqqPG88IgS0dN5nZ2gC/yR8f/g3A6CwEWjrbAwWneAL8Y4CSx/+E1DqLDmr/KW
nxz6KVOvopuRbJn5K9hkn8UjTjAw1tDg3saYGtAOU7Hq4wcmAluhIImTHZ1jYEbmVcUeOoobdNYW
WHdtETSnIXzdqfudkEsXUuvN9VQ6drKzluVlbEU7ez3gO64CGQmrr0RXUAa8+TX56zuVm43Ho0QB
oN2wb7/DBZMEy636MU7ZBnlnMaLyeVHvL9spMwzgZVlwdRh34MvX8WQ1U9g5hC6H3IEPCgO+Mxht
pPKiyZmg4Of7e7l4fjfmHQIVIEYjzHmaClMU+JTq9fP1t4IOM4MoeQjD096QK9W07iEZDGcp/43T
fy6W5JgMfbAu7NJkl/1KDE0rZZ+OsYhK2aKtK3NPKTIwI65lEJ82wX4ye+ncGH8Lrc/h2bMsHi4c
DNRJa/+d1z6HgSlSz4pzYtNYRr/9MMiJxojQrXeWe298CMy6Ho0/b0Efi6e5o7hnE8dE9vzWTw2H
3BJtX0qeUP9Jvg+/+medxNhs5k+lfuqvQYPFyMDpplwI7MDXBghZCcirmGh7ydBh4QoItJhofQNf
rg10UiVSzyyq4qje7n9na/9BpeJKkJZK+qb9wui7Lg2LqryAOklV9SBpjIJPbp9iU+lVfz5ceara
gYt/KaMBJ+Cuxu0cuOrtcSGGw/KI5QnCbbEfhOYgWo0sPZOxz+7qOEldTU0QB4qgzRsH0iRmzw4W
OilFe0Sz+u7DS4C6glJLmPGcGvkPNnaCRC6NrbZMsV2i5bNnRrgtyeNEuXMGItj2v+cEMZMqMnq2
xMsZiFF2pFILOsOE4zEoEHgxJRijyaDH3nmgSRY5hwVWvmmyAYUfUjtqUjyE52YJt8AeS68+isDy
JXi++XDExvHqHCMhTJLK+qwZarj8xSBMCeQf8Zqh7oTOL11eyf+BK8WYl1OSA8IMEQwjgrh8s29+
9SF7ss8PkPuDJ0wUniHUSWX02V89nfdz57QzC2PNmtdXkRQ1Q0opD5wEnjMd2fIxxGny/RnWkTcy
7B6zIRUMntEK149/KpHj//yS7kDkkuzeD3POn+CgMLbUywysu0MgHTd374TLiPb8UEpWw63YeGXU
8ydoqfxONpmfB5XMMgUvrjiy6vtKyV4WNRTaJvsBVpCdXSnKM8Wjp/rKv2bDXWaQSeegNBnqlusy
ewiQan3XZTbqHggAJMOg0nh8Y82UEwWGYNeK8cs0hbMREybl047k4gGBLW94LxDI4dL6D1DiFDjB
RlPgQH44dAFFsF5vX1SCYFv0gCaEHkBURKJJQfhnl5DBepHS2k5SQMAIwjdHkaCkcXo+dwHgoHOe
C0vk0kT+r2DuflBhILtdflbYvf6CTHXDSGUmUi4PcVpHqm5dpjHbvpb4PQhmoGhZDtbB3onGrczH
l+D0H/NuowhQFKfxjx5d/d3Pd/ye1aCeObYCcwdioUlkgOB4QP1ZqvV3n6k32eVZiNQOP14E95hj
Cgle+e7iunVGrpWAKl52VPKRMC6gEoSf5bjjdFbf5SgHItNrxgZ/NjwGrVvLlL2gHlpLH6a078Cx
Xa18EHvq65oL/cjEvTNcuOnM5vW4kAFy5NaSU/vG7Se6dpQdFc5oBhWcHgEnK9LoBEa4MQ/00dxB
10mLyoeacadydkwefUWJmHqcE8ELvK4GfRCeigNX+dorjvskiAaf7AECUQxxaUmj5bytQUxcsL4C
DPTKzzAI5dO+252RfIt5XQCtlXYqpJyXkU6xVFAsWy5F0L2djy+NGUwq/0aTVl/js32jOcP7NoBM
HMQaejOoum154ztJ8WWdNKeT8F7LwU0tUgFLoXUeRFhGUOhDMLaPO+Uv8AqUCqpvTFiyewbwKMop
YB75wAlHIf9ugnwar3u6na4hNteCEnYsA5Z0rBNXEhRrJk3JJh0+6dbCsc7WoEKOo3sRRVwgE1Pj
gdrsu/o4TfsFTJLo4l31SeVoPaxMzlpG8Vhqh/4igzB5EHicssRL50/JcSNWtgxhOz+hIaZWwNen
wKpGeMiUuFuQxHLKIzoAThFbpadfOVJzSu0z/dH9QeYHijaQlliFWF1poINAvxmPRYOcdRNXbWNu
YBL49FnK/8qB4S2lGKPLVuo2qhqnDUdsnwurqOQN2g1Ca9Qf6yFX9Cq/0CN1v/GEq+gXZOP1AYtf
5EpNn7Ft82eXOF5B72TR4LPfRC/Pnsz7lmqA7mOeUuhH7ljd8EiYOZ7XuAKIMkpouM0MdqQ9EyQX
m4OUapMyM+fhejk2F9hAQDmqSBVO6O+JNv1MHj+hpmjO4bohNwt0WyIDD5nCZ20ZA6qqR2YEvghT
VgrT0titEa+HJL7EBLJPd1KHgGMgn9AkuIUopcdmPgvEITthbguMyCCTwD5eUYrVSvEdYX4SLoCV
4ONSCEWT6D5/Wl3dFZg3ih/GHfJ94sirpnsd+/mVr/wPvtnMTRSjrr7xUIrLEWnv9ZWvxOpcVIUI
6HLfLgag0pkkkEgHzqo0Faap1J7yituknY81SN+pAej9OernwebkX+jzO6+tuuOtKK9hXBIBiY3L
PuwVJuAneeLaRthVPeXoNnjbLYxsLZdqOIGWrJhma/8vVwxLREl4Dhdph896QrzQ29dpQAIhEFjq
0DSWn6/8UN9NDOaaVMABxSDh2u0T5qX2qjGmQYxBXda4EbeaX1Wkr305+5MB1tUbh4iVE4aP/aWE
5hfMZnbWD7G6vnkA+cE8/x1g1OGo5lHi0hw8F7XhYVI6h0Tyefc9kID5WPjIyTAPrlwxkiSmHzrS
lUdX5/AbRU1Dx4Tr8ZldqgY/E1HJdq+0bWXA2mob4uV7P0zoe0DVe+GgxkYgRqMVNFDd2s4N+Ow5
mxefMdPzydWIV+L8UwcFH8MG/m+Rt2H6Gpn51WpNXLsGkguOotaUHeOG01wNBk3uz50LEMGSCf8K
E9uTpauJ/YbFrBs1V49PP2Bp9K8U5ECK+aBOdifLu1EfGIgu5LGkvlqNFMvwEaXTBTJqbgqDViEa
928oEH+P0dYe13T95QeBTNxQSxRWTs5XRO7+EXqRYQnAebJ2vYrpWfb5ovce1zfoX9kLb5RqxLm9
G/jAy4R/WhugynYiZ6YNLxzPUxB/vIJEND15HUDeQIyzFxjiroJ/6irgqj0WWhB9TnXaZuHXoYXF
jfcix6+pJSFPf44ZK/FPMxUhk/EAiY4E4Bo8zbxHhEYY49ykS/5HjOawG7N5/ZIugcm8Pj4yVgDR
IqnNjmFWA99cQ7hb8bpaL/cYBI6kTK6hqHtV5uaPpaECjG3V76VUzTpJEV10o1lKZg4LgglqgdAS
RRB8h6L2MSClxaqa4KlXpxlrTn0RzyETHAkApRrrN9mN9jk2aLNzKynvnEopNw6/SRUVVCuUg5Ie
6w70rM7snfIX5goRS2Ge3AqRnCRk2SITdOW4VQKsai50QXvV4Ns3HwKl+qCIe0kc35VuzXcYElgd
IWEta1wGi1TIec1scCrXpINeQBp/Ypj8yyZeOiFealrWWkgNJhUtdMMBfXco6ZppMZaoKAvRPSTR
OAz91QaCcWmKBWjVimUBFxNp0BBC+A650QUowW9HhS4MMhzvH174v0MiyVs/v6hBdfsMZU2aE91J
skgRt31U6XQUkvHKOhAxPOBGG/u4kCdYUY2wJU81v0WsUeJDp5Pxn/lIzr0EQjGCKuTz8HhdZZ3w
gleVxvPBLtw3kBQy9hNwIXZU3xDHIL86M4mgS+Uveh7tiCEDi9N3XUQkZQoIsIKyDbkIDXS7g5GN
LnDQoZS/bjwrizifQSRRLm15R8Aw8wxB1lenjutg3TvAwX+c+WJFxxeB/7e0ceKBDXn4vhCV/gN4
lZ1C5S1t+/M/Hf+zgPkHPhyXJtT9eTwi2j3qgH/AZ7K3DDxfSPCG09g4p6UGyieiZMIH0WAfF9Iy
z4d4CsW3yDYw2hOVQ5u8uTpZCPT629ZrMga6kXNeklmKTZ4IY4LiMvr3iA9W8k7qH5xJhSdNXVZC
DNN0ja0RB5gcw/nRXQctjT1eAGjO6b+k1GXGUFDLnV9hFGrvtP8Nx9vemo7u3cmw5W0FQVcRajRn
B2pkqPhk0no3q2F74qHnSznZqS7l5Xccpyqcn1gJ3MjopSFaYrsaGYSm5wpPO5Ac9fDzTuSKYnzJ
LD1+12f8uEatPaDASIePF29tDo/egAiCYX/gtQZM8R0KyRfdt9slqIZbrLudGRcx86QRgze6cO7s
0BAoFwg65GygZLHetIj74nYsZ0Xhal1mxHNMdYuMwy6Dba7Lxolt3ng8xBGwGQoisLVFzFClXL+v
du4cGf4KRvxb1WwH9EMie2gmaE0ZQaJQbVxvvNHgLNYfnW87pRXuUOv+MWAzJ8NluBX67q52vdw/
c5Xncl/OYoGNTnPcsHw10yHqjCBPRHbawy6JrYyWy6xk3z4u9Br+M5XOFnasPA+18pO+xqAdh13i
1guy/m4P6Qo0fRgAx8DY9nGLoPxkK/WLX8QvlqjGD97erHFjknfFYi2PUqe8gJ45kFWee3pywsMN
0cpk0K7fhbSSMGoLApniyFUe0mjmWaiblMYVUlFyWtvUPusE6HZQ7jkaPeaFiVlqFrO2dQdhiaoQ
xpCYg8IfX3zhbSrf5HdqPrq8pWtgJJr21oDDKZ+MVd11MOwfGbCEZBuYKEOOUR1hcHiVCN1blYe9
LwkEQ1s3fiMUZcsUNjzW+Wt5mR3Cf3CMsnSojHHk+qgprin/zg0po4sU1xq8c7PvvmtkgUsT85Vt
AxaQIW2SxAE/Y6rJwifT95qojlowCYua5adzJQOllLTJVmp+ODavtVnhj/HDdJbM/apZUMs6eyWR
SwN+aiXTK+B5nqLMTdiC6VSZ73XgD8PvTXowwqZUC+seLcv3UjynoStNC5PltX2qNBTLE6S0qSKT
Yrj4Y9R5VF19wb1Wo67vsE2NJzkRAZUJ5q+Hx6YjggmrKAs5BASScuQ/cOPhvVnoOi7c/LQm3+Y1
xi6ZBC2AL6JJksbrOVuwetSCVAsaustQKEx9DJ15LqS4Vnz88rlN+WvkSXEE8QYaE1aWBLi1tY8t
85S3Ot7Uur4Wqq2LPeMVMLD/rH9TsU/ASxY8NpXHldryprR+j4zKHnLW9ZswOLyyPbq9OaCgMArS
gHGdO+Xun/AvDXQkU5uGHJcEbDX4LQM2aFA6Za/HqoAzTXYKfXxhNzxNBHnREaNhw+hUPde4kDKb
KJKSG7b7Z5RYk1WfF7R6W8la04k5MKaHwZdqKE52KMGEhFRGGWqzXpI73hgUYit4HrkcHjo/Zsoc
uOby4I7oM9WRlPOIVel92m8ka4Uwpr7LBxJuLM2EVOQ5gkUiPZtwQlIXcLZ/3L8Xyy4HICVNLNlO
yul/dWvhJhDhbUfJnrVDxcFhH0sqEIggW0VI0E7eW4UMXWYGyT92Ev/4+/MMp4/+owmHtpd5PuFm
y+Cobm2hqGckenAWynSWMMCYACM8GbgU93y49SyI8RwhMZueVQ3aUKJKcTNY4sIGs9digo7Tv8d3
J4JYOZdWGBQBTRVIoH3JeYtrolASfKYrDdXpWaJJV1rgowQSomhNqZmA8zCN8dcAjAcrG8zuxjTL
1+upYw+6armSWThQqrpb7rVsTpsp8agRlcb1c+I0YZEAsrOUgfSuxqv4zUhM8oJg5Vmqjp74uLmj
WS2tQK9hSrlj7BEwnbkhclBa8oDyByTFghk4cbxuic5ShTqlDJE+e/RyyVCs+uvbZDI3SkRB3LY/
iqX8OMyhcYe+a17c3IbH2WrsPxYttX9oYK2XNxVapVSJJOm4wyY/m9i6pHSmM37Aiwj/oDOG/3mG
SrHNCWIptC3MXcq7kxZrkmKgACCYt198RugKT4tqEXeEXmfe37ZYEp2AB9PVwTw0p0O3JhRwXNCa
lCSf+YKM1C2wq735w25nnEkYtMPmSEi66Ew1qWo2frVVuSFIWroLw3NG9/pe3YA3L5EaKv75wrJF
mZv5kZS0Q/quu2B2q9VSciyemBRHVjHocLdmiBs2QkuvxUIRYq9ugGlD2FlttnTP9E2GOgnDbVzO
wasB2t8rOgY2KdolQu3QarWG0w/QcrWZkUdf4ZDEwmnHP3+jEkdJjro7nUGUssK45c7X/4ICDVgP
PHGvxHeBGCjewn/O5YIZ772DhO4Gfe5UGrSyV27XJbmKHl2f6nRo4GMVdlq3m0lOdUAwG5NmsbQB
evZe6JaSMo5OBt6YMpskXIImPcukoP0ggRm5S37PaT3U9dF46IuqCYg5k6XNNtw5muq7gwAgZqkY
PZxauTLTrxnXOdEBZKChGbjRDjVM4baEpT60pdVP/535WW/ujQnigoEy7XfyGUk9fr+p2xLF+4d7
rtZYtkYuopJpnN1PZkT6TGnM7+Fvwany8yNxQ0YtUOId9SmepDsxpygeX/UEdk4iaXdq6Dv7uGi7
q3cglTc+mgLRJWXqiDOYzuUXDO/KDfuHUSmyPLYVn1sJ8ViDt0xYi9oDYEr3h50R9fUM3FDjMWsZ
TV1yK5hY+8l6iBiATt7LcoOD+glmj6QyOay6OeOk6u2TO19tLFbed7q94jmo2QTUysZM+J+QndGo
Pa3o2KFWKvyD9RcXfhtlcpcebpzY23BxcdvM4pSTu/CvEvyCFmIUJMiTTKisnWjBlJgcwivy8Ez3
llmRvjSBxqW/xmBLZC9WHJXknQhY2lh6lUqwgfNfMZ0k4+4TUeQd6mf9YdRCtNZaCPJya3piorYL
UDTipgof23MXWGAnmSWbYiWgBfTygH9V6d6HAWNnFkZHCqPsev0opGEVa7G0NCqMTSwccZuXuygs
OQe5w9ODCnQAboukKma6Jduh/QYm3ZK3R0PD5EFUfExfWvHT3GykzJCGSX6O99u5mo+n0+E7ugM+
tOWBp3ZGrfjhodJA7acOpUwUfP+e9nAaMPZKTZJYScJNT5NOTpaXSnJup+ATyudGWfDJp5gJmBj7
zL8NpCux6WBLqgpzRRETdqGgMEFK0kiCm+2DzbM0S7Ngd8MPotVN8bq8ztCw8KYUdMDAVJkCGHVj
ul+nlLv58zi4ARkgvveQTyLpREvLeknU6jtrWrZOyQhwKLsiLkkh8WTm6NINOPJHsDgY5VZLN0DQ
Xsl8XCAv9p1D48tc7s6ah/OiRyc+ebL3bkw5oZ9k5VitP1QQMToLzLWZihjk1cEtPm/NiYIPzGO8
qXCzB7OVNgDVTT3fZrXHbQj2u5oIu3tp5g0dX+DMS7iZ/KvJX68LGAKnuocT5g2zI6qh93AEZEsB
uic/AuNkk6tbRpIl8oiKyPrUN7oE3645rimtihph4oMNAYQGEVGhb6xcSuv55gk/cSsrYilpzfPT
mo37Nx+iGl4NLQJlQZvj2BMLx4wYXkzXQ+LZQC/6bQgg9UIGCb0KOiy7qCv2mWhb+VV4xd67mgWI
PsqjIQ4PMn9C4D7lnHoW4GysnENFHyD5xM3oZ8hQP/6sfHFbTRf8UbHsaSDK7CYiniKmiFbtWEku
ij7OIigSyiWiBmeaULOsJjl+E5+IRvrEJCqFROz43B55uyNks8i0mXPivomKBQvH7pyI80x82myH
RjFEYVYiSbWm86/s+vAG7q9W0RR9ISzXYXNifM9W1B6BB1WgUfytVahZAwuxk5MUlZc3ysxC/TtC
WGMmSyFxJTxWXndahq92m3i39oj38IHQwHCCXq5i7p5nRvKIAFShAhzOu8+VNQfmPjB10DeDXmuV
blhx6PgcAPwQ34/xkkcC+8k+on0Ntas7qPBdCaJGyDccm3KtH6vY4NAq6ow1OUustdZaTB9O+zgN
nzh+izluDF3iRS/ggEoXgSIhVL/rCPwmGAZFpmMwfvqe7EtdV966lHIK9ROAqtHvmhhfJecCZQuS
r+8WkeDBXgm3UbZXmCeALGD6KupwK6Sv/ad5uuOwdDRSi4F1qCyTz4K2Pd//kGKy7G2UzscOzgi3
ZcvJ+EoDWQxlme13z/2VoM21Pf2fyjl1XuwVyGMhdKjDZGbE+QaosMGCu99Ia++CRA8qk3+sejQY
Fz6CpYzmu6uYpv70C1j7b9jZez4HWur3cutjFz+UbCRWIayePKzjEL6K4px9X97VtiTKlIM5ytb4
HlA6xXvebos2f8wcIoVgpXe6wf9b4FAh79s6Zdzrx4iviTMfbR004WSTlj5/7tcobBnruK3kYnAD
xBIVcszSDWainT3WvZKTBqVD+oPMKucHhDgU4+vKZb5nYIIzO/ccdWd1r6KwG8X30QWYpxZqir6+
cdicEPgYGLrNuEz9J0v7FTyYnH+80HG9c2yaW79/m92lNyMX2LvN9FahJkf2w3dDo35fvQCV+84f
fRLfKeDMohgQ44LwY/M8mAjd0zfGYte93BtdEbIuF7BUIVgpMD/4oU0Dt4St1Yz5FREipbLTOwOK
fLzCAdJtQe3EuTMZEe1PGrTt3U0/lHgm5dNk5GP9PdcS7NYuT+UpYxvzZVDkr9rjt5PkaJHzRtaS
wx47wQ+HDvAaEndyJ6Y9Obh6a2LYiGnIcQC+x098b3cAqhbByNlKA7d9PyiWT7baaMVWgHwLtSXG
XL9Of5iQR4vSwAgrm2l/ih9dVDCnPLThRXncMrNOXMSjbNKgY2Qv1zr11slGoKkhlwKVVsgpRn/M
h92pfsjhapH4HO70w49lZNGAKXDvX2GitGHW7qDseUkvZL6PM/SGRZ3iIAtK2jYumYnhugIexJXH
sSrA1LyppWNCnmacECaV2QR9DJH/+xgYDr2Vn63QxjSUxp5iCOOADf3UAY1kWMopkFhW6H3StOIu
EdEppPKIRJo5G9DTcMQqWUQvLNcXMngX4YFJszgahGWtfRPHrtWQgBzTwRG/jrhfv/B6al+TTY67
q/QQ6ALCf/adO3BOqPZD++dbuMWRS7rvSaV4zI52IVT9XBg+8Wlq4qPduPRT9kx3L9NjLSE55kMP
Yc5gR9egJaSxbpeGxxf42vAugStfL8rme6iJT9+8ZFq0f5RCz3FBosELKCO9jRe/lExmdCSUkUne
NhiQkrmaHqBBvCmAdAmFaz8Vea8k5MXAMfjS/h2746Ufv7E1UOeFTKFw/9RTmMzPZPFBENrTE2cJ
mPo71IS1GRjHM9RLaHX0TBBWg8I2Bzdhq4oPrWnhIhM3wZY6i7czGFCxm5kIUCXSjA8jev3rO4T5
zjYAq9bnFfZDbQSeg8vsFL9YMHPuwARKn7Mb8hynA8gmTyTaxsrA/cOj8kPoo+9nbChf+sCOP0ue
kGbQPEdCMr/yK5tXwJ3+p6loas/8pvOaO57Z9gdf6LrSdZfxnHd12JMlyBAAutWdmwh+9Hdk76lI
+qmrujWbYOIJhN7az/QARAxZNFBLqszBtYmietHTwKuIqxqt88uCDmqQk1cny5Ek42kBCbzYbswA
LRjnGLm9y1CGTM+i5HDJoNcSScE71WIyuu6bdwc/lVeSi6c+svzv5pK5F+qa6FZg4DdBFEFSWZyY
UjNT6k5yF7zrSg3J+Ui1GhBT1SLHDdH4XWPUa6NNtDCfz6d57ZYCjdxovwEvD8v1hdeDoAmo0TGX
K7If7yz5cRuTMwGaciUbaRvt7jtqBrvppVlrPX+tEyMTZzksen4zyZfxisLMaMnTY1+yH8zzciWS
RldBExxDmydbt1K2vj/b2uvK5zk1GDvpNVU+3DG2wsGlS8+CQHfeCI9Mr9Yde6ReKKptmK9EQGv7
R1eRv9FNDKMmE+Vguj+MbcP3rqHEwTrlUhFfTnzPadLbfKxhGBiojJ3ZKndH1QLzFACLPvZrMQCV
N++VW8DQfXo0IVydG9IrflGFVLH0qUldl8GQRMVma4EsEXYSPG14Gwmg3w4/iAKUWX+AgafiiS2r
9KOwDlPfH2kynE4x2eT7isspt5AnjmXqbEi6avocrntk1n+vzyhxcVIUTG2PdTsT3PJgzGdJOZtU
w0cthxI8iTkKcPuIdEoF73chi6vPdySvbsN8kQgudltPM7y+J2YTjdHWEH6C286OyisYdQpNsZNG
FUnmlLhXAyktcMW5yoSlcbsLCZ+Hi5QAp25b6naDTHJsXs/Tj4rF523RLweS26ltP/qLT43nOV/Q
ufC/k1bjrDiq0au9pNY/xHgUj3G2Ud94OJz/1q3qmsTqhQNLhuiHxt8GL8TtmtbPZ6ZI63zOVRUJ
rAC9AcDU6s9XXgsI0mSCbYDD2y7OxnHf/A5Qsap0PuxPN3hmTYr5VRo0UPr9/eCvbeagvNtS5YvE
2cTt5Ia8HG89/4tpXh4qt92A5IjAIPMZhsmdiiWV2DyTFgQyZkJSRF7ftPh9ahpXLtbwmYq+DUuS
AZzbo3KbIKNotqgWjO4+e54hj96/EUzfsXf1fXpqmaJ31FJCoS4P4egxjoWh6ZBpb1PZCD9pNZUg
lJJ1VAbUhzkuPLw8c+jG35WwCN1QYGiscBGjDTbFu1i40MJcvSQ/yvVjqpmMI4q7SG8GNlHhlkkx
lzghJrGngZD+aS8/ju5b9rlbg5lY2MwTz0oKw73f9Ex6AnFLgtIhYCGkNUjWiWtYSjBmkJxWVPgr
HgnJdxnPO9LaWNDgC82VLdwe78aZFOxxxkDPNoZHcT+N4d2MhPlt3vKd14pSFUHOwkiBi6eYntmm
QYvdSNkR42hVeBIPvrmPzl0NLECruOP1QHMGXlxBGGCjZaPRiCPAGuJgxsuut9aLphjdWiOa6ztG
2gv0xP8UsHD+wUcC08llgWwLnJpNVC2pBRByzhvLppM3hGjok53ycabQxN+3fyx7F01ImCr/cW0g
nxODxJiUu3goERtQjJzJnGU7TEzH7jCg/0Gj5c99/aml+uXs2G4A/Z4U9EHocfMFO1Tdns1u6VqC
F+ejBj+F77Wd9WeYkTld2VYIn7T4V0o7boVfvzmnWj291zHc3e8dWu6flR/ug9Q8BH6ql3PR85J4
PZckGXae4Wg1HxnYY1bk53tsWo8AT32kbCshj88mejTrEfXrZ/LHlldXpY53NTkqvrJxaLneugP4
Q18or94tl0I067sGg0qLOuz873Pbsj65cVMqVJtVugfOmnB38bQC44aCqj6brtWuV6mlBBbOmOft
OICGkd7/GDXw2y/9jqhc2jNUB2wz9TabCrkmJ45zcRvKLh82882liZrP0GViIbc7IN9g9To1D4/y
McOEWHn5nw2Td/wHF0CpSgeOg7p6F9B/qu2bTV8M+by2mntBffdokYQZuMl+XJivQrOwECC7S3w5
wiAhJexxU1WkVWeeTxzQyJ9Km4lh79oISvOGgrAVA/SDNPM/wF+ByYiglsArsURyVwngLboRAt7O
+24Cs/0LO0ZiAfPJCmk4/PRdcNUyuBHkaVkg5cqa0hvzQ42eca3Q7SEmPV03ZYouderojcq1EkSp
QcIz740N1w+gb64969cWAzMGIw5ieunWHdAumj55YmQaI0Q4IGo8EwbNdFXiazkHD8jVO31lRRJX
SJFCyiu1EIm/N/R3YXV2eLEIc8seOGBDLM+bY1vmsQanfdVMUySJaEm4LtfHbxRLFr9iQ4vLRDZK
RDsWDuMuFKv1ALD++a85BOqU/shLztikwQqBaKqUOlGACylEgeQF7mFReiIXksEpoe8rhTJxbANo
5xkonnU3F3Gs3I02j1iJHm00xXipxp2KAxPS902R5qahkcNDukUUeiQqATVV/6mp+/OOMV+ji1vb
3BIkh7FtFlmZDniYJLdx3/cWv/9dC2TWKzyU6btpU848SZuCVEcdvEKBnOCuFgZBe12bwNQ6DnJB
uSJt2poXH1x1U8ZrxN0FuetOCTPR2Q8StTZ00k3I9M1s5yy1DH7MfzMGCEo9bAx2M+79GfbCDYgs
5NrrUDmgI2+eQbvwa4orY3y+6Rmzo1+6A1XCfyyeRz8feWnP4PK6uoGoa410osT0ZWoWBDT85k44
Xmv04vsLYsX/zuYmXRg6AekaWLhwRv6Cfsd1PqmVsfmAe7ktPtbchoNbL0D2DolVbxk2iTOkQ864
ZpIx42iRU9kipEl52w8ZPzZ9NvR9HgIdFtMIDdl/1pGFkxT85IVIWoMsVGSYGkzR7bV+44N8AHRN
kSmaVEL4rRgH7d1OPMcmLQZrWJz9SIHedV0cYqF9gHW/d3SDXaPzShaIo479eSc7ll3eCOYtAzgU
a+zNi7xZkGmifsxjgwJn3ElmedbSwGgqCFsQl4fzh08BE+uZp0Fgz8tFMk4wg0SUBVNPCG18id/a
ldzr8vR5dX+71mE2h3VtuODnJIn8i5Y70DZUAKNRTMli+9T0m9wXSLiClqzHQDPJBsAMpkj+j8/T
G3MGYhKI8AHUP/W18vGKMIuQrZ4Nuo1CeKiPIWePyRFoaW/qDYy88LjPk7fJofaDjRv4cXWjZ4Pr
mIplF9gZclodVlD+98RGuFBx5MWztHxxpD8/vhZEXRTdmLOyY8W/7RAC8Bq+x0nybJyUj7lM5i7C
wa2ZCsjNboPzzg8tKqu4kRZYXtnx/mR0QI4oe1qU1H+HrnYUSPjSqAEEjzjBKYq8kxNNo2nANbb+
l/qh4mctve4k9zwJfwhQgaHZiw13Nx4HjT9/+zgE/S2g4BMDjMeYDx5EjsH2V0mMWqArf17J2fon
3IYh9959d2LjSzKO4dSzzzNQ8rsm6nYvmcaHcDicyelgNl+1Yz1mKClN7EPakz1gyJK77pH/DBJ9
/mQ/wJss+sjWlXJ3pSCsEJXGprRPRMpTAa0Ejqkv0Dp/U1Wgw7Tvssxzn3yEhXXio2hF+hssyJ8S
R1km9uc01M5v+xSavxCp5CtIQaHFM3l+aUQkijCNWkJ13Lq2iFawuOINL1RtJxCN8RxDgnSDiesu
ceBYtLBLaBM6YPxiCD+BeCiq3bcfIg3FgsKekSsmPjkdixeBtg+Lsmp2aFnG9D69jXHRslmQMoNF
Tuu783PjWAn+9ur/6zxFZC5DWraak1hUJwrpBtac46Yi9DZWw2zKQpWq5qPgGYGeNvttZqIKK1Wf
3cErNXUVNVXFyJTS21ove49Nf2ikpK48aeHClMM4gYmuPX4EyRnl1P5auhpBUqenqb81UyPbnVDI
1QGcEQyce3gITI3os45N71f7rMYkAFDaFJuJFgYKyFEunDoh6ZV8OuyKfmHSzc01y7kNyGkN9xO0
nnKWcJMWZm8yPXoGpJJfQg92cccNNAIJppA3l+nBYl5SGwig9IuMtl0ZT7tFdzi3b1UzQiBhXGab
VvtEGJj9JMjGLy4p0kVfFcmTsKKNx/RCtJzmmkGPU9qTXoxjBSnMUpTHibFLhL+2ka7bgvuwzOuy
2GkwvtJNmrl1p8Ip2CsGEtf1/LODfTNkx257rWIgnfTHinMQrlEZkpPXp1OvOdj/f3/q+IyAXQEq
2ZoOeJoNeyy1+lGIizL3yH0a7x0/Zu2PagF8PRxvwS1BGrQiyErfDhUr/iwyiZLjIaBqtQQuBXkJ
T7720QXJBLEepOEk9727V59vgStVpyqXRtYaK0Xgl1cwnWL/t7IUT13Hm2uAfe9GqoIN7votssik
NjBgetxL4qFrt2zo8m2df2m6Ki1lRolGCsPRiX3qubMqOvDS6eem3rHYSXoqFKlNsQI75FAnlr1H
6TXGxeWUgtIrceROxldjtlOAnNZQhKjZUIyZMvHjMGYZRzalywkw5n0SBtRatI+1fTkUJEIBk6Ma
TWoQOIhHZ0kY9g6iP5CHnMkDY9QPXiV23CFJZfNArMCKIfZxweJpXAW58hPJWybYc5a12YuF/1Am
gKMP5eJHzg0+sr83nxzDhyj69o+zsMoK9fN5/lrRIt1VgP5pB0ThvTm/7QxPBDEnO3hPeVPM5k61
NCvw4H+s1sz97wAPzOYVXzdGKXh7a7oudhh9bbgZKyi+/t6z/rXJ656GCAlPe4bP3ySidPf3D1qY
o129ewrpuVipAKnI23YS5btG79fMyzGy/GY5AXSS4vKsbgGj/3/n6dlJ3gOdpgaoHFFdjmGShi2l
H0eJsncKSfUpGXz/tiBKfvO6aiax3uW8E6RlKQemZJsOz3yHjwxFCltmYJUT5CzueOYS234xs9vh
LRz+g14BZsWMwa6Y8TeKwuiHsILgN/fFFFf1peTbR5UF0mDkuhW6+rEjFh9U1PvxC/xzPPARM+rA
ol0kMvEPsO3iLoIQS4WYkQ/KVbhg6O8S/KlYvvbM9UT8GdOdo6Zd7MbcRFZowa2n85dL73CujxG+
bLwkDKjC/t8R/1l+x3bQVWOO1/aybYnnODNXIHaejVDQcXPeFRtU/xxmsWtMFQtqeoI9TVLdHe9p
8MBdj1g6Hgobs6EVMW0e93eF+DiPZkHxrUL36snnODu0OGQ07w+KFYajMqK1qTN/sGEUDJ+P9lvj
dFf6GB40xWBdWiaZornHUzkJgov8tJhO5OKAsEW6Z7uSxRLQscXiTyGALsflhd0EtmhULT58LBPe
W2wy/oX6HkrjDw+HGLftqz7Ub9SmwKwR4Qj9Ij+xHfYkdF6/IJbmnL0hR/Fb5ZkpV40JymjWbMu4
j8IyzwjekNkaDTQkdTOm9LONN2Im92fmwUAHS8cxNKMJM6gX4XZLjjZuOi9DBPLN9mSTxdVCxuQC
PbIoIuARYFHFsWStGElvb7EMy2Vbdvx+wayiPiCCSsSxwE3aMyFNLXeT1HzTQ3wJQje0IDkmgtbU
R0bBnCBUIYYmM+eS1st8+rdHC2EvzVMIaRitpsJm4eJRRtn0QK7UoriRx5J2w7mJ9KryyId/1G4L
ZDMm4z2mMGIB2rzmr3hxQH2JFuNzcr1ORXj5F9cEhbKJOS3IA9BAM4hGeWzlFFYfC2MRNME5fAh7
pbjehnbWYPeSu1SqYIXTjmLsgA8dTQ/M2HKjlzz0gnNUS/KXIt+A1UQwF9XjkaZ/xhWfZi3yUeDG
SrarsZQ/j/siC7q7bgdypUyC17FfJHh1EalsWMPGA33jeh3B8MqIztNdXqQyMcvsyTF3ZfI2Uhog
ErK/ZK3epgwr1j/JbGtNsQyCE9veDkkB7AbZBobkmVy423UFdMvKgot5grLGotRMxFYDYvRYwYnq
tbFuy15ll0Q9pjwbhwHvmCCwJWtuTiNBACxT8q5bPyN6C3qPhr+Nsa67iLxH8MZ5OUi9ChcF8cJr
R+Jkv/HcX69h2HPNJ3SDf65rjmoHz8bw9J5MtxMbGegvTAa+pQYt+F2WgYZLBxq3rpCb1tKV7KK6
nwochxbtxKxemlJwEH4uFrAJp3Pmesv/bpax/aYK15PavpxwZnCJ+7zliT+2pUKQtW7QF+6wuRDH
3AEksIMBWjtGUP8snOwc1srmKRjS2pBU5mL1akzYgnxaKtsQJIYhbRokEk7uuqi8GakoEELIiDw4
KApqceYuZ9srYQCDprpRN86zpVBzgr1zAWXiqHxd7wp3vD5tf9j/Jl5I7IA8bi0BxYr98Ibpuz9h
oxlk/Q45DRtcMYWBccVV4fyktM4/f7DRsK5iP05plTD/gFZJvLwcINqM7Rc63uxuoOlD5CzFvuBh
tkXmZ9TeeNWEtnVFi0wR9xtIUtfpLoFn3nKREYzLmM51oE8tVXzfioxep7XvOwwQT3qwdaeI7azE
y/tSmqmfMNpFgm1RnlMLemIPqCu7Ql/kgxPJ1XR5lt1Nx+5hmYq55P5DgDXqvodrv3K9qO6+k0XY
nuTF3PmeUXOjK9uRMmPlA0J+kHXXV8FOXsGxuJ8Wqf2zHe0JBuWI2GDE7bKNzwHiOCaiwCOCX20S
9euZ8oUHMSBBYAxwptncACrqP5GJNyprXY3BOuRO+fGNix+caxh9srwYaiDT2QFne1CDqlhCb+aw
WldATPfBvQCvC1JiTUnZT3Vo+opy/fs8Mx7i1OyEWsProS8OAhuO+FzVU0ORJIeGFgt77A/rB2gH
idhZPnnkbgiQELGdScoOGyUVgw+eHSI3Zr980QLddkMpPEGBLbHdScVFPIe8ZVQ+58PbTA7zgplG
FtfGyIW846LX5EQaw3Ke0R++4xo8lyo/OuE8IladrQNG1psYJ6GMHIbApgqOUvIZIBf165WXyxPJ
xQ8tu0sL0V+xaL338BFdT4joyaMdYUVBztTax9bjLyeDeESPXbVAJZYOCDiYdjRfx0Jf/dHzybBw
J6hSnuvkQnpvZjg9IGQBXt8SZnfeVlyrImYSb9cgkffMPuTk+yht/OGT9s8IpPtTXvc7cdBDOzkX
XlGYmS52Z4+GhnSkQLreqlJyz9q8aUNmFrLuL+bv7IdFDQgL2L8yw0mQi1DC2SvTaqnp5PigYUZX
Jeu7mnGiHOCl6FKdgp0jVkul4idQmMj7Ua25yv4vRwQ6gc4fcjD0j1PrLVMM+SrdijbJJtoY6JBo
/b+cJTTskPNH8JyyAz4SeCsd8Pfl7z5SakasSoSofMDS2c+rvX+P7aBdWbjKTLbCGxzlsTpwXaVr
PpLNFHYQUpT6APPtPztXbppWUS9NfQB4aCatj+Ovc+KhNVVV1TWbvhqhCctSZGrccH4U1fiH7V7Q
Sbd9Av2wYosuWCxKPEg5ELGNC8E8h4cDKP6rPzj422G+VzVRscoxKSMmRx66GQV0cV/pE5WnXsgk
TJJONYKhJmXYjkO+OsP+/1TcptO/R+CN6P557Y7Z4shq5z2+PFXvWY2EcCpZ6Dne76KMBMBDZuZC
0mDXuerJGJdE64MxndLz1I5WyF6h9C8tMTZPWd3RfQgxQzYveO7Njb4en+6FGENRGf3KBzzkKNbU
XCAOxjrANV/98vmDNc4vEhxcir8vVaDFf+2/T0R2lrOt9Ft9TxyM8++44rtJhVQac4DfIssZu4+D
GPikkk6qBfLCiR/tTmcPCq5pczARvnvCt8la+1kNty7ImyO1XR2ndSRrKuznwWYfpV8+sowHeJU8
wk0oJpRQlsqecHLGjPCNzd/qrNJ409yGcV4o6YYvXvBBDaFZtbxQCxMQW5UN5GumSCIrrwYJ/hHu
OWXjqnPqQ/aMfmnukziJXXFZpiJaGmmTEMavIDsvcRoSYzmudO8xy4t571qzN9lt1zYVHmwBwJwq
l7qhKzxbgCfb8gaER/nRE9SIrc8DP8+Ef76Ab6e0QK926KSU1AVCl7IdemO+kKHQklpslDUA3rx+
XgO4gHBkwyCk08/qaeZSr3UjgKVwTQ9NIA/2uQHAXqGOUUa5ejhHPX80BxHCPTiS1SGuJ0DGayFV
XiWBnCmFspCJ9BdPn0ViBgqoCfu0BwZQWNzdE5CXCBkTj0UdTLol+5Hn9YniV2f5hOY6KZ5ChVFq
WwS3IhUSAHBeQoSJYhyA14p4qkA+iC8OvExneaCm7SRS9xBhSZ4WVHuPuSlyl1wZ6pWWFT7Ed1Qn
Wc4SxEWeUHdBkgi6BGslLbbvNj/OD4cLR3yytlr7A9GbM+vQvxOKJUTuED2PsfCvqXDGouZenIhm
lg2265tJFtTrrBAriYtfgkwkCK4y/57yrMRjalF5nR8DXnfdvyGnKIghPEgypQxStwAjRjanAh82
xWeIldG67lmhKNdYX9Nb8cNLu23Mtl3CVys40ritVZx/uYJzR/Bkj2+8rJ0ZlXs6Os0y3HSu98Sf
T5iDbLSO5DHWZVtSUWQBa8JEDDqStH5Tsl6y0vmBru4s1UYiMg/cDVeO0QQir6eKsdEPjGJnX6fS
gyWStL619SItWQ57f3JiywxXbCzzh7P+JJg3wGEMZqwwSEFX/M0Z/qjQLLwjbGfSdvhJSCmU15z6
5oscZ6supOXLyOvu0yO4gy6AUpReYf58EKQMznyM3yNWw8pz5ZGSfyAmoX1T9mCAjQtHFhQc9VJj
xCVoFsehUuzXNX+9HGMQ7oxDUQhohSf7xfXMJRLiimX2rVdDaDr4IdURry2oTfkUfWlu0hci7kYk
NsP4spJWGdQwFd5ShbhoDu5weMu9sVD/1tqt4M0KXRToQaFsq0jo0nXeMnYJjyCDNudTQiFtNIof
4MqFk53F/bkYNtxOKK6Y9OB85QiTFywpt6YH7l02+LNUQctXdaZzLYikc9X0WwXVWK82jX5Iu8j6
eMrV+0i50xnNDw0JT8z/VLlwcrH/xbVAjj0Bzg8k0ZPLEHy8z8Wtd1jY1R0mZBrfpBQTkm/VzTtv
wmYrT2GhOWeq3TXZ9VH31QKwWeIttqFDoX+/4wjPiz48VaH8H9syJAPxV72LuJ/Bk+D+M0R0w/4Q
pJV8IL2XjWUTtmDqO3EYKli1pwRMJFbpa5po6BgEQSgCVwybfwfuw4iO/E4VIDEGwN5zPQAm33yw
/pgVVncaBP0rZZptdV5j1T9KJhBQol0y0xITeA0PBdTLoFHglHrnSZXfzsvSfPwdLiMB04FU9W4V
0OeID5tKM5T2uoyzKzvBJOtuD2HmX/MHxYWZlnwy+Zct8tzmbF4xrqsswc10HE/BPfrXQ2zZl4Rh
BtbWipWYlcYg8R/vgbO4sfpxN7utzcT24Kb+0TmEULTLmCc/r6ACAY8M1f3hrzVw+by9yMINxLU7
8FZKKWit4Y23PsMx22REQlXAHba4rBmCnlS997mhKooZBvvfhBEkO8jXVH3zFrVPCsRJvmVoDiBx
7QtRx/XIYJQhk/mFbTYbEwiHIdWu4sebj6ELSIq6j6bEq4tZ7rymgB3BtFmLxg4msFGWuq/L7CGp
JZrnV1jwhKGvceFYw4HAkC9QAk1rCNPlJjotkKgVcBk4t9XC/z4r+R/wwNnULo4UYJBy8HQU4r9q
ZGZvWaV93viMvNJS7hVrAkirD3QakFO+YFF9z0enak5KMu29dtcDJOfqSc+ZsY95TmL1TpoHVPK4
iXYykzREPJfQYpT9ZX5T2DpwodqQ/H2TZvBWaJ84qgFaLDok7Y5oStIbE59XR+kmBgulM13jmWkp
QCyhoUvRIIRoZu2N4xLNja0Y3LK98H1FjAMmgFFBoUNmFYjiR1KqDzLCBIA5DFOkSm6SHM3aCmQy
qeV3Ts6/zHEhn0EGrhMeYKHqen4jAAcwogn7t8hwpYYvUqBVgSgWaL7pRpE0gUb9B9wQ4FypacOO
FJRPVuls/Wg2IW8D1pwDJSxZRb7gHD4MJQEHsOexhIbY4O2hRbHQN5SiKL/ZzcNSYYv6TgbL9cFP
lo7FWgroJi2B1XlmNn9EYBgHTD1Thn/iYbyuziPD84RmydmcYZohfx1anWJEyuibogx7N9s/lxnv
RLGaSFZthqGPmcKS85Hpllbo3tlC8/+KR7BpZ92zwbJR6W6zxzJLruHt4kQ21RYsXczRz0VMzox2
JHfj8pShMTJ5cSvgWW66ceygDzHHvetfyP9PyDTyRteErcP2PDZp93TF+DezoJZD+bIt1fE4hyOc
OSqzVIzYxbh8dp+Y8xGh2nAILnkvTQPTFUmMKQQwB3E18ik1DYLvQ86dYVTeFwOK3PdJpYPObq7m
z0TeDkSolLjsT2JQOSZhw//him07R0P28aGaYf7LOj7950f70XQnYA5l7ubVZhV8XFXdcwxfp6zL
1FOm6NGcQml6K5rI7M2rUMZkCdL0mppMWjmGxlRGBgSrhVeRYWftckGc6iqJLf437YvEZSfx0qEo
0caZH/JmeVbOzFTqYZB6O3OZC4rDOegr5BYt9R6W4feSESIAKf+c/JAxjLiyMG9kOSB6a6YAi5UO
J8aejfxV+pW/fyVpFEM8iH4VR9amz+lR4IjHZlXpwPyXtXUHnVoYcxpR0bPHkXHgF5wLHq0DouuJ
sJXCh0pruuPrkcaH3eoxL+jkK9lQNYEkRF1K72e2n+p9AWMcLQwn3lZhmyHFzc4iA9cygg4oWKyw
SS2ue3S1RYpzu5m8sZJUnwYDNcl64CEk2OpsknmyK0pzZBiehWegQR6S+9tZTnKGTzUwyJjjiTYV
eGigfqRCYaKML4Ku5iBNlH9rkDjAonNZzpZBBY6M3gA/KzDknTliKWf98Q3yT7iegovgK/y7wYZ1
ak2WtEp0WHTxNZpRxDdDFS07FqgFV3CCy045WHb3RIcGCXOgl1PzqOwm1fzQnmQPDs8zF4gWhNFc
h8fOuWEFdWfDas8x4zW7YQpPS4hScgazR+E1QcpX2jYWcQAc8I/aaodgrZhYqPvSnJZxLYYRiIny
+AeXWXVZ/KLti/yChtEiHczuODrc1cRarw7l2RdzI/TXZ8o124JdCJs7uu8wzqlIeQivUPiStpbI
8kg7Ftv1oZwymOD7bvHAxWVFDc0oQzKMC76Dn7FQg8oAYbUCRPhEKubkvXJO1qQxYTiOOm+1xgbR
zg2D6MjLLe6aTKoY0ZMNXeQQHuihsk3yGz2juDPVOp3q3p4hQI8EF9zXS3sq/MfFUGJrI77738Af
rq7piX2Im7UK6UxcacRabfwS0+THOcSiaw442MSkRe0KFhj48a9DWKT1aZB/w1zrWWQTazJsXILk
DYxTAKNQD1p0PW/BRKP+dICa+OHz+jc2iQ9Eij9Erd5XIQyWkilYE6z62ZQnmecJURAGrlqAhWbU
GqJMdF1OGpFhBzZFgdzRT/x08efOIle5Iu4LwIFIdYRIXInTZVQc9DG0hRY8Mc3FsjrTZMcoLwXv
hjl3nfnRvwlbEXhfS6V6D9a92thU4Ge0MCqiSAwOaMMbw2orkOIXa4s/EkBCXIK4BzFP2wvVZpSA
5OLbae/OGnDFeuy0EW+hT7ID99Wp2UaPbkgNH1WdycDTRpM6Q7KjIsBx/hiZ7+h/A15hHwmnkf4M
TI7TXlgV6aOMh29RFSPGRPB0SvHADlJA13WBlZ3PRLBsxODbkuiNf/qrE6flwNCCxlfHGpzavRWb
6otE8Ze45qEMpsqvUBA7arnbQE7t9g1y1zoP+kUYOZxWEb079AmEkBfoP56B4WPkCsNB9z+NkVBm
24Ea0zwRfjvgL4jaEep2wu3zYbLCKfPtaWgxn7HV8tQyRm9jdaeYlvzzLFwSw2PMLvJQyuoQXtJS
DTXDBmFhK9/S0r+b+K/k+C8tLYi+rxlygdlgh3WXoLT2NYsOLiZJnj9ANCSKaEEScAcg9KV9kPFx
BPFPhjytW36HacDtrXeg/fm9sNR6/k/vqfTpraUtBAOuv9tG3yiOFgbqLvt1Mp041JHrnrz4TCt/
wljN5Q3si/MjYaSJjJsp79RNNdFF9UeZsH9Y3TNtdAhntATkII0w8XU7Tu+wmZhBqtHmDthBdffZ
9JyQ8PVi9DJGIjOwrd/zC18u0GHrlZlyrbNPW9/b/sodMaAOrhwVptByYR4o5qtQTPCsi9flOANN
x0nGpzF0JKtBPy6EJ/e4NNhb24nx7IIbDcGfsY+0fiftjAyS9y8xvWXfO7in+NjqenM5rTxfi1eK
eD5MPQwWjJxSKgoexKQpGwVu8oTgsifFqLEXw+/HwEsGUfF2F+uwulmTtWssgdPVDNoDLOUNAhsA
9SRkr6p0vTETWjj7LJSD6+05T9ubRYJDcl3CB++qJ/PrQDDYeAiCgo0RTYRApotCTnSf32Fj/u9B
xE4VhvOI1IkfK7Zi+3OvbNoh910b/qVa8aMyH8FeOxheRKir4+ziWS9z6lWa9fSjoTO/3QtqlzpK
4zHC6n8WH8XWjW6LiznIxTMo6FZ7iui7GEEjepqffldbF/dC+Hoezr7xzYwR/V9Pt8FAZHo6WQHB
nRtAOwBqBqAVhCywQP69dsMLTEVR19EShmE32kiWTeK3TosaM+2LqARgLPXtiilMiHigJjQT9Gqb
iKuJLHg31sAu+caf4KTeJm+AZS2uy0IWW4jsQq9cX4KkvV62cCUaf1/DtHidVEmxW9N1938T4U5P
X3Q2u0RyBxZaZ7RUs8082XetiBaQ86FuI+tdoUesc9rzZ0A1UrM5DHRfJn2IWhmSkMk7JwJfFjNb
drUz/CGfjrk+1szoQc5l/7vAdpVdto73IU76tkm3qXIcOIGKqybSufRDDCgcS46yA7Vv/FW+88QS
pDeDVt9ohhr8dgIUxStkIe16VGQFWJFpvh487DyePGN1JQOyTCf+QHSA/JL/+H40RkQ2Tyh000HE
Omq45fIW6fCBf2MAVjfUmzzXdZTF/yNaogYz7UUFzWWqVB7c4bkCaffualoF033Lh7m24vsiwBwn
N0wSVgohClD9iNoEof3tp7n+Wuv8mCuCpxtmLAXwx/EweedVBMEdHvS2ItRWquSy4+F1KOv5LW8j
prKyY5vtzTX9J8+CFuztLlWv/SqTWYaXJkbIx9U4zMryy9JB3YBR6UBZnNbp58aYlDkVoxuUEfwG
hMJEk83NL+lMyD5xcwH9NapoZyqsU8GVZc9OBlk0IaaMKQv62BEePBaqvzkYR8zqQtq0yYpI+Sxd
hvvAuwtXOdHD0HAjzvrOQW1ehpuKrRIyG/mbq1UM+hb6EcShRn+HArVJ8rBh/nIte/JKLIS04fRQ
0zdlbykdu0muOLifFQ2hNuqzW2bJVBWMWBaDJJqsI5n2B1L1eR0Y52Eiy3hoY8acMPkKdZNIWUgx
tuEJZ8LlXGBvNYBZ2kPyW6RkELGT1j5/NOp7rcObW5rtGL/9Z1MXXyV2CK3kHnchY+asBiifevvM
MT0CJ4O2tHYP0lSsYGU/GPHHsGjk0+bjRpr6AvFuYnsvq3UwJKe/BOcyvABTPPeLbllY2R9BjpBJ
dm8hKC9WOl/LuPVgy3k6sp5Z6996q0oqXASqvfXkUz+3bIL+GE4Z0x/a5cRsmokLCVSEmAdZCr7Z
HQ9v/iq/05o0/GSernX17ikLKSPA35IRbqZRLkEL4cVyr9JirYtkXXSwhBpyErqGfX/VQ/jtD5jR
Qwhve+tIg95QRoGlZ99SyugJTBK9uFVeUxnI1OISxZyqeY4Bgr4DHyoRJOe7IYrUGtIJGFT0GlC1
0+83soTyMV200Qm/MM8nNythfvNJpZizRDmb+L235ReZvdDxhnS7qMqlL/iBvPEmWUbcox5E28mo
PjpteE+tszSWKEezTh0AyIAelUtYHNHpHozozm0DgsX2BfiVZ9fJd4iNbc83bhhy8xQNtZ2374xl
xtoEumoxFaZXc38qtwqFl2J0Dg1VrpIznEiac2z85/MyZZm3d6lc3tBwlWTaj9lSe7LZH9jYX+WQ
9o4By5sgU/7jpuc3vLZOfAQaga/ReCUcPaGNrV1aKBIqK1G3OmhQ1XpheNz/9+YAAuAqAZJirC8A
CL5MiDRNgtze30UnGCfZFQX+q7k1T2Kd99EmmQr8wukTzDaTxqIAS5oXtE80E7sTLPGiC3I3ZPen
ISrBirXaA30EsPLPWCkhnsOKZ5R+MJJx7kEaK98tJPZ/qNFmo5BfxbL6t48GDX1feYsZfTyXjniD
ssew8HuaFMGnbT69spzbFO6iU+ZXbDxPxYewhHQY9lNe/c8cBflCrYZYXBQq4rgRrNPjAsJZVRyk
/dZgLCVq+qS7Zs6vl+BFUAqotM0t9gC+gK4kGR2gkAVFL7yIpO9V8SYGeOjJSAm+tsV524Ek2NV7
CECT2MQAN2Cgfnmt2QnyRh1gWu9aAJ+ir3/mJeBYYBxMUi7l6QEUyzDcvrGrjIvkylKYwXD3ovIu
cjhF1ickTKRiWmTK7UVlUzmbvvMypOpUJlPYhQOx9QiPke5jIrXTIuB5OmbZ3s+MYLw/JxH9Nnrh
NpQVrM1orrXuA+L+p7XJCKgj48j5eXwq9sgap+8w33ZJxJiX9WY5Z1OM5/tz04b++YZGXIVCN430
ELNycbJNyaEydrWHoydNmGrD1PuBvqJY4i75WJcKFasFBqB0vG7s9TDISNJkrm/7JgA5A3c2T0TD
8f1blsFbNsWQw0ta5SbXLBdhbjtx+bulC3PdMDelcmAvWOQCsED3V9o0FliVjhMKWg5ZwiRu8MUU
S9fixEV86AJmqPnqBSei03BDGSMZlyckOsIlRQMBxZj0V4v00JaJPQk9mk8QgZgUPFSKXWOk/U9r
hinxJrzDDH0735/wgxh+And9ljrkkpfR58KC3zUyvdCn51gjdkb7gueVuWJcyn7FZvyD/Wf7QOtF
CKmecXiW5yk2XpfF1+IQ+1ca0uRHRV5kQS+UKJP2Q1WWY3xLTi3N6aiCcAlVMZsVS/U1+21ewpr1
4ggOe3ovyrDD1TO+5v0SkTwFjxE9TeNAN4DCRyLmb9mvH2IcE0w9+7grHadIf3ABWTYcdc5zvcQz
vzv26w611NMDx5f0I9I5HG82RkANCCz7hO9heTEdX/zVipSVt5geDxLHCMuFdNb39guczIcGPME5
c1aTqeL1sNvxmKt1SXmsAkauzMgOu6llmF1D7Cd9nvk21EH5pxAvcmho4oZLkWxm25l7/XMl0Xf1
cZ0iAnrmQJJYABLPwB/kpSs6SQlakhVT60hQMv0lq6RVuLfUObtRwN2UCu0i9jBPjolFL+Yqpeea
B7+haaKAJIlmpobHcXymTw4+Di3ceH5B41lFUGxlG4DOCAljbNz7mwAf/0T0Nd33WdhYXpX7MOY7
qR7KnQO3YZ8C1tzRhZtuVegEQNlvdTTF5bZOXSC2Qmopg3v59jbnTiHJZA3yz+Q7C2vX0FPosesq
Wz5AI2LOEu5UR3t376rwkfR7N8EMzf0x/uwTgJ+BeRe9V7Quqr80Z4NL+faFOuFRCs5wi0oxdco2
JtYJqEO9h+yU7qZAC8jH4Gc9ozyOPwlz3eUGfyymDUdZepbtAK9gQcrpnDrPOBWjePkeZsKCygVo
9PY2V/OtwdYXPZp5I9OCMR87jO4enJPW/fqy+9jJyLdxFBUyKs+IsvVKMTyTgOhLJzyvyePC+6m7
+6FtHoTkFaNdlcZlbME38jhUVue6opODr0EKonoZ58+tmGo1+mDZVs1uLkNUiuhO0z/ZIaqRgcS7
uZqNPfeWgtH9Z4ksP6ZxmSzHczjwvwf3f1mcf2cMkCQhD4N8mcA66K1tSrwC0eTEkr4Zb7ueqVqh
kDY+B07HubyVNibXvbY13pbcQffcAvMELVoseK8Z+DQozvRjQvyzfXUCwEbYMysxRZUE6ez8Xq8Q
PkOcdSNY+yrAujyj8x1qwIYtJUixegRHk+juOWTua5PiNLZtJchEHBcYgqLK1VG9WqzzYau8qqAH
ap+K3sKyoTfexxFi+HtbNg99qDcirVzizNpkWif0A9hDIdC0hpApGrusQFW5M0hRcS2IGPPJfRCR
blYVXV7uJZTeMBx/MchylXYE7+4ty3VkXRmFfOrG3TPvq5UyJsJaSNG274SNoB5eIxmL/aDCLdSm
4bS0TkDZSXt+2n6sZHA41aK7RF6MTPTcdax7xpWnb3Tv7X57ffbqOhEx1C0dRLSbaSnHmaezGLiR
rzl8EbumEtCYdY1N0kSfDu+juG0IUhddpaVSzHYQuOmTuWWVeGMiQ2P2Mb8Wx9igoCsOh9KBs4C4
X0rwYjYifFihfqy0OrelPEA133ABdwqfOVKplZPhdNSvcMTlyZnT5cNRO1rN6ALLYOWoPIKrHDDG
udwNuwkq6QmJ/5yQahZPiGvl9UIGiKZAdNcw8O2R4xoLiOXUBwXnjIhmkX8f8S0ZxtULtlgNJPG1
fv3UwhuZXTAMRLF8Co6tnCoCl1JGR96bjA6HVpkZk6y8txm5oe0iNkuNpEMb4hADkKqoyoUpsRT/
ZaNxzY9iWyhkPvtSoCTYLuELPEdeLtkRLWLwYWcleC8vzRwE1oLYvb4IwbJEY85lBnH+hD5eW/2l
RNHHreMFjRZgsdSSzAIE1lR+Ld+KPfV0/Bn4DOoEGws7e2Nqvq76/FH6wy1+TUHigmqWU+RV1HaT
eg3NroZKbQzA14Y6tz1Us0QC2BAhxgbcejoEznSpYxOlTlMz7OYclDAp5B7q6mblGj6Q1adx6U7U
thuCwzazlZMQ5DxAxwoUl3ZjeW7O6NIi1KYJ6k/AetlZfi11q9t7dE6i5RfEK6hqlaTF2I3mC1DJ
fGbGbWbdwy7EZJX+Z+iBz3ezdQ8PraK7MdWM3mDcq/PTXxAPm8bOcUkefDVmqY9Oy1XKa9ZjSUXI
oRWpNYK2rT/j5GXL0dZz7XtMt3sC2B1lgFav5rRInJ4GDIlO5ELGitUCJyZ+UvpqiU6swEIXYRsd
AQ5JkvkR4zzNX84SKFwE7KTtqRlOPej61FvAyZFP/7Y+j7I+bLho8hsbUMUZTf4pXUxNN4oom/zH
gWVhLAKLSVOst3dPFtL9PIzTztPC2iAz6FB52inSWJmqgOmFCVuGu+NH4C4R60FekfmWf7Adlo6+
hynkZaffIHb3LF6mL6rUFjxhZSmxMZYqcJwCHj7n0jrldjfUujzcGvc7Na+SnoQ5F2IfiOcBuu16
C1I4hDG6rfPzK450tqdqaI36mxbHxyoCWgO4AqefxGKCL8fEdLTUHnKZODGEnP77xZHvZhwx7AaL
FNx9u3y3gVjVEqvaHzKpexhHSyDcdho0g847eJfOgynlMC2KxtmOMgZh4hGz4ROmQPA7WhKXwuG7
hDe1BGFDSUvS8dboZX/QJ5ZgOl4R3dZbL7v3mOku8hYc5aUjiJwMGvPyBzjs4shSpzDR9rprT+sC
rbJ22lVmJ2vx6im0QounzUXNSPjfaa0zTBoMntgbwZ568QVF0gD4bh5v5wlh+g7Crg6Q+r2Nanzl
MEEltF2uBHq+wY7Na4HqeIyd+QKgq49zYH3aQCuclZvcuavvi7tA8+aupBA44phLpcJAQ4eq845B
W2f8rUhY4uD5h1frN2IKT5d8xt3E17swyVX2OR50DFuNY+2CNnLy3qi3Q30yD4MptklWhxCL5i4N
40W097CvR4c/NeAsaTP7/q9rdxR3ctoit41wUWiNblff7uItbJmBS0/5k25QZvHnjtBh+q7ATSNl
wWI7YXtFe4cKBp5M9TCTatpe/KwPclpiefjBCizGMZKCyhuvQM0iKR/9EiVi0a4v8H5gFSHEpzjk
Z2hG0EsPbacJfwGy0vT8AXt1sa+GcacTdRZljUtWM5HBqxT/G3N3pMYPXCHuyXXJK2Us3RcZTKMg
x9//VeycMrD8LZwSoilsthM2WDVRG8xTejYI9ib2ofHcXyVI/jryUduAqmJVF78mq/EbAbDfdXx5
J5Rvezu4Ojh+xQW7a7+87jLLHBtJB0Md7h2adQdZKGZ6fdFrtLcr5giIMVlaQDcVU9eEoGxK19ko
R1uVU0DByTRQH9FQXOBF3I5J3a7AeuDN0t/GP92Oum04ch69s8nU9zPunqhHkBYMylX4xPcVxAZq
62H/SchVT0M1c3K5u5nH/cEzhFXhUZ0EvlZVTJagHic9yn4r1+ky+LnEUmOrX98Fvw328iqeDO/B
d2FZJ4PvL0Yae5LzP9FV6BAMoG0g+vnQ86IBjkCHe2ftH8P0ESD0800XZTTjTBhyPAs3ZUnZnkyc
13HzM1loajyWAKqFCXUdrkI1Zmbz/MAxafhu9VivkInDYr7tBA3fM3xwdBsftk3qyS988PsVYD5p
1zYUpaZMK+VchHGHwrcXe7AZQ3gIBVvdKbyfd+ODsLqDPHHLBi8RtFRYbSV6rrrN11mQX3qYc7oN
f3oyvxERBJnM38UqqqrxRht00nL1D0Eg1W2dkV9GcKg/Fe6Z7jeBJ0vGWB+73wLLnq9zWNwOd4c3
3GzKb/qPt/f+31BbwhbQFxyj7SInNBdmpPIfTWyOjU7pdFg36KHrlIukMn0B0Uu6U3a/6D6val3e
txKuMqumO5e6n6Jlb9hZQWpHKPLxdXgMQfj0SXD6A8QfTTS4eIxLtCES1BptcveV3USxSV38+/jO
db2qULJImOLklkS/b0OMMUk22RX1y7YH122lEhrWLvoBQhw9N/WgxeMbir5cnzWSIV98gVvtvndc
95Waad0YX8RFjrDyNaIiYs59uKpcgRMpavHTecQ2n2+fEnlABhMVhOxts2VSOXOCeJnHc7V7nlUo
NpKZxzrLKzAK5s6NfX6B66ukrcBmq4EH5m4aMqOtFek8x8sJ2fyF8M5HzFg21NQUAylZBwm/ZX7h
2+2HA/zUV08yXuKMTzZPKYiNcheFTu8KXnzvuxCDLoxx5WO/4UVkTOJySejb5WHmf04nFp9tEmT+
3R2wDJL1zwfsxIgrGz2I/zDgUkp3nqiWvu1+MqFAO+W488AUoSGgax6mcO5WMYiNAVkVWP+LzSfT
wVPVxds0uCkSfpbGGm0FLpbtuYHIkllmK1J0DKApgSDPMAynFR0u7xdyW9fOyF97AzyPRpQ3WkSb
N5TZhWQqpDtMkIM48xJRH4BUNhyBMA1GHgZ39fMuOmboFH+Cskb0YyxLKG3bKXVnG4/uHxkUTw8c
7z+GFZvZux8bKcIjdCgch/l45bFeuZI2TByXbOqBlR0BL2ja+oqH/AaQJZSkV04Rx0Ko3IbJwqng
JHtJVS9gtMcLVKB5MbIAtJF/ySK25gZXrRv6pZ4Ip33Kf9y4CVM8GfrT1mgSiGhnyoiFglB85W0s
Ox/TC+C8s6pMGpGF6EbwiANKPo+ucN40yQiMSInjTJ/oCIDIWjcX4r8RWRQX/TLmxF/sTzFbMgzr
TqMd95EVwtE43PC41zTQXaiYl/fCaRG7jp2TmoQV60wsjcP86q/tLsDbsvxd3ZHIW5P/QFXnx131
sanon3NqB+lByBhSC0zcwryKx+cW0/xPmVHJ3820ugDzvcaHZ3SGk1EnT4WEgWOyuH1x/KBwxlGX
yc1t+JB8KgICVpdXEGll94XOClcwKXqBWch3yyWD+OL4mTehv1/7jH+BMa0PZoXWaQsPDU32yqVy
5Zu9J+1E5+JKLvkBh38LyISMBnUU2Yu0bGncoqXPS9k1M39UVgUhuNcUOnfJJyJ7zOkfjhk0KsBi
ZziYyTAWhugQ6zGYb2u1h1UvERDvMpKd6NQ/v7WMiKI/9agPhum2klBoQBQsEh2ciDYhr5ibiaAh
j1DFSfESSscaKFsaWVDj+ww1fA8AaMQ5nit1Z0uGAavEtU/Z/Aobqz0Zu3LXuQBOD0ta32y7WqgM
aKeixSFyPsCppq9XKn5juLQl7HCaeZ/hP1yN1RK9rv+AT7ZwBDNB+QGUg2EJkF4c2o/GKuRN2eYD
UF5gRS6CJEj6sZnmKuj8OyXmA+lJoRaKRTqQDQ8Sjaf/gKQFvK5ZJoTFyLgxBNG6OwBupXi2nUb1
8u0U5WBB06z5cHjEZgfSA5qikMnYWhdecQ40rsYuIto+cPXP4Ocx8hw+2ltAL7AbZpJgjMjxhpUS
zUZwAP/oJqx9y3TZOn6uLC4Rf3aWrvam5yTBqR+8Lm2ovpI7Su3GtnBIQt8OJq2qYXgoCcYakqQy
O5yqeEo2Vmp/VXPmHBZ1H8VfJHM6TV2BBQnot28VuS49CNVGfO6WyUEKZvxu1QRR1vXxS2WNwdSb
DjEEr9OBTcTPlDv+eOmIfubH2URRGTQJy7KTd4BXDx42xGZWYzAf4Uq2qXVoDwpaPDAYroQbDOPt
j1pVyMSFSXBMmob40xLFDQwZj6w4bTK2qEntIT4i3QgOw+ppxDqXMRLmfJ1/2ybeUmr8mdkA75ae
khcYt6bLIdMJ4g8/c/3gB0UQUYde9uAxjaTRmKRRpqwhbCHR4FH+vuPNcno+EJ/HQMc5v1hDnPGc
piMyJK7eIITSdZXGok2IGnkdUZ+yUUGPhaX2YiMMUpFiPJ3nDxwdwi8LqijaTSjh5lAavMwhwLSG
I/rKTX1pErZPBsO0RgsAZ71y4sor0kCkp7nvtmoTteqIC8DfCWS1C1ZgIdExrJ6AJui8bTAMLzek
/TgmQfPY1OG0n6/p4gwNLTXDZnhYjggWUCiuNre4VIYzPuii+x8q262HiGEklaCw6b2B4GRx53Wn
/8/i1CHGyO/jE4uJ6AfIm6t1ypOO5x3Z9FRUDKypsUOgkoQGoxixYtjC1XKskAGVBVtGdcNLlk6e
07HAVZtjkW06uAFak+i/HmyFQNMaEdKIesJ09SJecXYUqKC2jR+FiHqAspp8N6a1fBZcFyzkwNJL
AdDU/6V9+6uiT72UeQNwXLHL0DMZZDeR9uOmPLW4GRRZEZfky7MloMHrdaastKHk+JfA7IiBDPPM
oOc0pLgH7XlfsEDEg9L42lbZoEs8xeV6PTgyQfNAyIvbBDKCQcP8ZHSdWLkC19GSfa91BDCkC1/w
LH2hE3r0wR+zpqhWNOQ87QgafLwCoT0chZVZ5yOKmJB6lsV5PbyvmRzddInm1Z+0ezcx9/idn8Bj
CJNZxTF8gbcpf3QRHZNm4dwO4Kz+wXiA9Au6vmjAe+MJ3/9SCavoR4B7UbCNkjL1SpnsiV+y7C28
TcnUBVgvloF0F/jJlk9f+1SQrApMXA4TtqIJvZxThi6Ylltzw63QafgyJju3ifedHjeSVuCZGsXg
DTePASA58CXBqbEP55AzIlR6Hw1rk3FUaSuOAgyP+kchs7bgmUknGHDTa1QuFn8Cq7dYTI02HYq0
q6O1fot2QbpEacK+tyS8Ri6FIR2wgv3jkoptCmSWOLmTpN3aLn1NjkDlUPCgnE5KdKBeASN3IkES
u3kzjeqTV+4+X4ftluwg4OqxF7gUyx4JcQL+9zkJYdVVlMqd9DQImKF/Oc5XOwC+Tt5OB2zhO+4M
jL/FvjmSOAY/8E7zhFpebOZ6eGYfjdTfQWO3y7bOPDzY7WF22uZSZdQsYZnU/jVhIa9Q6Vrc8Pye
QpaIuU4l1Ni+3Nye6HQusOCgpC0QrgER1A1xtgFBc2MZXcGdUeKVQXW4U9KCxBUkB8qB/YFi4cBx
AW6pN25YSQLldx49nTWF2Nwn+MYfUtLtIwXvFyHYcY/ji1H0Ysft9qnzKOeGk75y9+10WYF/fg1p
D98Xhokz2TJ7RxEKwuTeJzTtIFcV0CLqU8lGamZsyTCY3RgbV39NYfytU4pmSMQ2l4v2VH5YGqOB
Z9viJ3t89uYNNVV5JHV7d/fap3eBKExJuM3DwbbO/jeG/JSTjbGzKY17/rw+77TN0uWlNHhIvj14
3mud8eeWp4UNDoHEzV1lofdVyvQTH5OkB2AE1Y57w/JiS8Diux2yExU9BQdU3vyVpil1cZA/vCcj
tfRq7d2iwBOpjJk/kXA8U8CbtS9672cKzml4WLNjIbttqI4gZnD2u4vAZloEo6uFKxRaJaxi2y4N
4mInByuZGBW5srLtFdpxgt7tbxjCLfuAxaA6ctoxfy8IkzVhFj3Zjri9W+Kt8O9GSYhSK1ufkM5c
jPdP6HtynpKKXebZZinccfOi7ULN688k4+Ze9AYpxKNb3uctVf+axKb3NEEFJfDXmpx+BCmOK2Fl
VGY4zx7jFB7shRbnnML/uDfuR4/Nu04daSiOjc4Xm5MYyZCOAzBhMP79QIWJMs4JLmkfC1lX5PP6
I+/8iqqpmBjy6rtxh+N85u6Rg5afqoaN1FtIts/Nl3v4D/kJX6PHgP8ei+6kvhr+y65z5kN4Ezv0
cIl0g9kvVAZ8CdTub2RA3qPSqZ2jiQIgBTG5y3c8dtQa89oQNJHBKs1Ukh4Fl0xfFAgoAeeBjsXg
lviVltFFnkTNd8sIx3RRajaNAIokYicT/ExVERtmYoLsHq4rZswRy0YxWs7E+XwB6cqQasd+48tK
nkvDno7Tzlae0xi9ImrMXh3OGg+S9yTkImmCcIi7eeTpl7ZypSgZbA+Xnryvwmspdez/DmvuxEas
idZZcaGR4xU1Nde5L0qFRKhbKlez8NxmH5+2sJmWlIyvQkDQJbXLfE9kCLL29f0s73g2vdDyjkL8
UykQRLAJfAGJKrM/Ta1AY966jmlg22ziqUZD/hW0VlKHech2BxcUsWNxHj+8Kd0Np/W+imbSvs9c
XbtN6Y84gkbr4uTEmokwKhIDHYVoTdlbl/ri4spFhjYAErzQmSbe01ypjzyJr9eBXhgQOd1CqSA6
g1X+yXMZBXvTiKSATcANuUCXgdOUHZiLtozkCF6HKylCFws9h0dH8gqDprmt78DLEJuLi5V4CBmn
sCePG2P47+FH/R6neMmSlh1BNdSqGistzX/mEaADnSc5zgepjO4IFZ6mRi21yejFss4H5v3IuxW/
/bB0oFathA0WkgcJOrZ9VDfhMITMwdLmWOh2qmQJQ79hxrxPZy2VjmIMrIebf+g5FRSOY7L5NCZi
2mNk49zjETnNGgPENhZR4PIcRu5jytO3UDwIshxb0uGSvAYz9RV2D14n4vSBvw/c33UTnR/6N4v8
PCG9MdkBw5i+WPRhbWV5gAj3aNBnmUHP13rYcZ2vj5a4apaDmpFPtYVCgm6XBpW1aw4cjWDWzDZW
ZRfMtgkexiAjjam023hxKVrwXm6lX3CSjDQtY6dD87O46WJZmmZAcl/msG7hkHfEI6DtPQw44UaK
Cly2eX1dchatvSIsy00VWgO3G92+Y8qHdFWvguoBOVpicKCIQfgHQPO1FvavwcxaZiEXEvqkgral
fkIirwV+mJ6YNwibbEanfkN6XwPpfYrSIG89AQYoPlNI/qDA6lNAdm0Y3E27qbi5EQdzcG/0VbPO
HgPruKDB79KTBTRaCubLcX3LGaatVG6eA+m9aZI1WixFmgO6v6ygE03Aal1zjWCIK7EhHaUcxdbS
DkoayyYsN81vP1aV+D5yRGNyMpZlDG00mH1WN/2SWaeZ7m9qKpzBfcMdAnH+Dw0Im2BKoOVlIwQi
RT3x4Rp0GcPQ/JW02JS5ZztetaQWOpmV/oqIzNpybLESrDln+6WQXpUDA4/EMzdfqH45TuLYhKCW
aTg0SI55ZcuQoQxhb++Zyzh1JDcu5z15K6Pq77i62m6lLHlYD8h+Gj0Nt1tftJmFc8QQkAWdfmon
gCj+OsvUG3tyXqTEs4DU7VZHT7Ts/X2ExLl34hnfHVdhWDyD8EVcPr6VIHrmEe7rt5FkFPXIkFQS
2mmNmOmOyEuv05DeSzAs3S4KVT/f4zn8JGiSMS//2zxyBNvgvrI95Y+V8kgLa92TKkw0dQCBTC7W
3iOPM9ETEPyzA0dGo/DHhqwHuRQHv7fDHo9DkRpaYP/jyQnMjCaTIXCxXWI0y9pL+WlGtsf69ro2
pgs039Fhx9yVMoFgjw04kXWP54E8NPvpPXY/c10wc/PGinNhuQu2YjJLuKz0Dxt2RSu9a5nZWLiv
f5EaCPAbldwb6bUlizNsac+gQQXPcBOUYCxmMu3kx4hq+ulCbyZl/bVf+oRyVSg17ks0JiK9lR1X
rjolZKCATYU0aj2vFzgXbiJc15BRwnz9pYuQ6fw6Mv7xgLt29og5hYDivVZvXwP06q/q6AhM/tqg
AUq/WanrUpLtN7lCJX43ghm7RexRSfYHWRVRHMkpVP8cUquL+hvQU8sF20nA+qIHu0PIGr/TU2t9
Y4soXlWQf64/mHXowgAiotoQferGTdelJVgvAnbY2CLV1eSVJAHF4MUp8H7kB6AWXSp9pUWOxJyR
E3Lr0k5dYWz7D7StC5QcOnIvDoqCSkusp2wUfIvS18EB0KT/c/n4QPoaLeHLwqjdLZhL5pzedbPa
i9B0m4cWZAsSHEvDXf6bDlXA+3tKVU8ThjC2+00KS/xvK81vUvOfgyJ+k0X50CqliG3ay5gtOqAc
D+aJ+W/Q50VwVpwCR1+fXV2+OPaC1V269wJ3p0rGIFa6NpVTNHX3nyScTuEgxRvOOSeZrfGVBPfy
LAcE66f/ZAsX28YPYmavDgRkqVsoBGWDCfhH9BG3RYaRSfyO/SJQRY6QYCr+XCu0RANKm7NxEofn
7dKubU1gA/uQNOzp+R9tiukHRsXVIeA9T5xQcqO5uOmr01bFvQYmL8jxP4Od934hQZaIZ7mASTCh
IqBzaLnPK5GC61ANGWdVnuiQA2DUN+9O0WOtQY1eLwv4gc7/QH7aRn1ZdS1WkW+HqrT40xkzyrol
zGC1sRRXvYURxNJ+yhdPe9QFSGeJnBCI+9vgd4iAu8Ga5MNbCqPuXyMPjshTNC2sgS4QDXUU1HB9
chYOPAZMhVyqYJTC0pPAksUCxcUCRX0Zb/psp/+aiuqV+SDIntP7ZQfnIggS9lPXf0Ch/vi9ZoV4
Km8CFLnLGSjg0GQ1gRF8sUmLNHTAX4rNWwm4o0ZMJq3QtEm2jkCivpiujkI71cCImyEnbxGZB71w
ID1vM1gDPEyVG8t57kTe1bIydIvFlwvJiACj4B9EXyfG6TcQsmsTjZ3QBDmT/k3cEqezDxVpIgYp
DDXUxRYuAZ6TsKBBg95cIKhQvjbmgb0tiRFYGEl77D7+CF6RUO7B8K3N/VlUIlDBiQXb2FyLWoR9
vN+pBVHV5WCZRzzuo5wacL9R20KhdO+JQECME5oWeWTIjvEIGRvHqz5vWOrE4oGBlo8Gl8X8HCPj
4IsgW5Eny0t/HkfrKo8842m+z1iuApjZCMYDEpZ1NHrdw+ZKwjmPrriNo9DyVXkUyFTo2Ccd5Jw0
W4IEirG90LhIolEqgbSHJjlZ8g6xX1DRdsqy7jpoSt9b/ZpJnsS+Gtjr0nnv6WVrh76JbQRbaSWe
KHtF6XyZ9GPBlz2kIaCHQ7Wj/gXSnCTOnhfPEbbl3QhQT8c8pjlaTwDCj0nI2uMn2/5C5mBnm5Cl
sSJ4K92ENOfz0xUwZFvdK9Wkn1qPtnqICvZyrDmhY4riBT1CeD0PC05TXfoiOIMvpR6XnTFeq6gx
7/bUZkYWwixxqCDQ2Kfj+uxBMfcPlP8NMT6UcC3zPBty8A6yHy/zKgAbX55yYouuccBcqKcm5DHA
u/NNWSZ4egcpJPtLCzp1jj2WdMkpyHDoVWQ2lIUc3Aczo3k3BjSG6yTCxotPSinyP4ESorn/hk+K
ukUFZFHlmTJt398/yhd3eBcqN0rk9wfsArnEvEBa36vSULDVGYuuY9+tETal8JzeU4eHM+pCM90q
gRz9XTMTMKUiodw88gh6l4vNw+D7L9yfLMMwBZoY4F/7AXBZTMjPg9I7LuBGFiKGATlhfeRSasym
H2ec5nM+4fglOAhIHtEXuNpRV57d2pJTC0ITm9YkeLl3DCDrQRvztWSu7xM7ck2ql21AynsLtSbj
15jafrqmZBgsHWriAxmSncnWjHsqdCX0WQXTxsepkn0DPEkyvubT3nlXxcNt8rs0CuQif2mK2DOu
cUu60QtCsLZb+Y+mfLcnOMGt6E7NJDYTQy6EqAisuDqfQLDu4zW4EDM6zOAI61eAQ/tGpsa682Ni
Kg6at/BGCZexZCC49c3tjCWzZ6j/Sa34CT71HQWAJksDYBNgH/GkibUqwzhy4NtjwxYorg9KE5eT
NZ+J/1GB/WqK1zS/HXH9Rqi+Hs1zC7f5b2+hGQ3Ox4Zfg2JB9FzHch4gpYkMMBUELr4L0WpU/027
nwCZJTZEVke+YGnMW/nvvUyoaXFurMpl4GfhUbjyZYfvl26S3Jb8zxfcUkb2mvlaQrONPB8u12Ig
cMkTBtLQDaL4sWGAoUJ7jlu3irvLDFBRD2pXNv7QvyZGmocGeb1iBUlJeOsEtOh6p2PVii3HYEJz
7vr0eG6zSMScyJpBshaY8Tzp9N4ndi5Zn2OMGaAgt/XxGhDOWZiSch8aChmUDdZvq5JXmm1FPYTK
HDNj+J7N+H6GL0ApKRyiJCkv6xEPlGgLLQg00S2S58bgP8ga2IY3e1tdI583z36i/Uevv/6Dpm0g
yIUwBqrFG55N2lrcuOBEM6wpsMGA5HCrTSxRoqjOXewwEjVsSvfxk70Br7+ev+KwB6C9ngcTJrKw
o58Z6hG+vJgI2+0BBicD9F7iaoUSgBTHKSQb1S8viRe+OjBwaAWw2zdT47J41WCiOB29DwE/LQlG
tNPvdSBQ5cmWmQsRUEWoMceKEN6JkkkpoMfV53BAmjFw4799KPNxjpUWNu5WFkSh674zVpkwD0vT
PNd6CjD61s2/hiGE5+fLt+vSASgzJaLFEDfxyom3FI0OnVS//csdeaF4Sjr3KZVcw4F419sN/0tP
QMYdcRnnJXXderrK+dvClrUom6+VvSvADU/fRjx2XDqaaLgCzq+uMnzDX2GmJovWIraAx6e6jjzB
8v077d1ixWxcw8TD5xg/Y/QpN3hG5zuXd1NEQOXe32JwOEGNRjazuhdaw0kQeVSt3Q2ekRzXeblo
IYxSwS7sG4b98dG36BrtSZqelv8oDOSfW8FRzgii6Ki5Mw94MpLZvhL1n1kpsGZ5g0ITt/ahkqVp
ADPOFezSA6mLVZp9cTOX01YRlNzsrwLKC9Y1tWHQz7tRCxzXlR65MNfVW5cuJFZ26ggaJcQUUzQP
f8mtyhHLzic/WwOPa0TDmCz7dgSk9ZhpIvYCvVbboDihmqCbQxjXyfRlW+1O6Icx9QHqkj1Q/A1l
pYBBvyofi8UGqh1YhGV3tjuJ7qmFRr+YCCcOzKd8JrstdsqoPVC6NMBCXveV9Z/zyDgWWfFBexet
O27lQ42PRVMpDZEooH8cK3HHFUDKgQdgghKwRrCe/2SscfYYTqQtLVF4mo6trYtsYlhV8/1kzHRU
n0jB6bOHYd4y6x7+0NWQEZsLjvChfQbYA2mcpTZreR1UDVJK1Hcb0vdGEzLEreshJVoOkXkXRTy2
D4vMSCszDDtIDRsWHQchu/OLnFjO1tRI9sAlkhqqIanOYetpmaGaPMQEV+YThojodPlrpwyMhtVG
4Ni8BpPdqQgqNw3DNgf2GkkqJRK4mcAyhz86ygmGsPu8eI8wmsuy+p+2O7AT1q6Kdr9aqVA3nnZa
KBBsSaRn1Juk2iS4mcofKjJqjexPsIRlStFN7+o8V4pphugCvriPuUag9akl5r6FxSWKMUTkcwpy
hEHsX8NWnG/PpSfxmdsBuGRpAqdR3WkyzjwCmKBv23EzlBeiTIgQ8hwlzNjJG/JfvM0n8esVR/I6
fnkH+0CX/t6SQiG5czqTll2lZsGqxb0+6gSXcatfjH+LhZxw5j0SY7bFSuQ5h/H6tKY8EM4g5YhO
/mktD1if+aRRmP3oDm6e+mYp12vM+k4b5EFaGni+JzgnNlEu/c68YlVthjKwmF+xQXEyqu8og59C
jNRTHpFKxgf0QlHANz/1X8qrKES50rLrYVlfiZQCPgwacMejuUKtDmsjS1eNcEcwhtTXVO6tNPrb
u4zvF3HlJL0zYrCK9P1feXNN0cx/SH5KflX8bZ8+FwTnSS69tRt6hjKu04lTrzi+ff/Z0HYvAEQA
mlpTQegrZYspvqpcA7dDi5FnZ2v1L5Vs1bQrvooUS5R1cmpoA4YIXi8J1QbleWnT51R6Qc6OLBMW
DA2ZHWiCAgYcQTTtQYdpzyuNb/b8bXiTapaO6HOa/JMH255vIkrikDkQlT/BPm/r2hUc2v+aQ/PR
hQRvnRip9Az98XTK9qQ1eQlK+zzwUg+ifaAY9sh05LZc3pkKroKR338eRCgZhidEawpupDJT6DZI
7muzmW1woDGYMyeRFpm2HwSjEHu0Pq0nYvmxL0uePxDt8+ue5XX3EIYUyhmjGV52qmOjaLZq5hgQ
cK6TwA4cDZSMjvvRM+vJnDv1fS23WeaLRIBeUYtLN1Ds3OlMJW6iinP7et2dqVlHr82Fr0pzB3nt
vPvx9c4TDgmoQ2Y5XfPrfHlszTbITHyrqoYh/AtzSI/4I7wjpdedUqH3Ni9TGpzDSxjUT36IbisJ
thKEZXxY0KhvUrbIQNErIekg6bvQB9lT+JRG8usuGvYHQNTFBeublxzCRC1O/0gijb71qPNPHQjP
blU0607xSGpqWNxLIFeKiELupWs3WTFBZDucWRE501fGSpfudfXILyaTwSqjs56Y+zRPgjTieaWq
tzG4UdBps89bIxiz+zB1xsM/Ay/eztyIC0106Uf64Q1LqsXr34BReDjXtIdXjUsz2TTIn//gG/vT
FjZ+Up81Vr43NhWH1ycthZ0NJL3XB8KvCN+1+BBTfc5TTkLr2DZ/teVJrBGfK1srBVXZ7mRHeFE3
rQJqOR+ZIevDyODJVZqXeijlCHjh6g427yLX6FaAB1zW3kP83Dj2104gwL2kkXFYGuXu2Xx93QKL
TmJY8nv8i09awNHo3OgT02ctEdsf4Q4LMiLZv1WVNjC0scXkfbNJwi6KW0aTU3mQr6q3kgmPkjM/
QwnaKnlhOn0Yqyp1RnEiwiFgA/shc13vpB5xWb/wHWb93R66SKKaLbPcHn80EFLxDSpSJY0tOcoY
kpJqtUgP30zMwfRwbgS3yF0PAFgZhuIgsyOTMfX66qBXDHUbDGI8acpmmPljjMmDLYl440iidJPL
eqj0wvr1ZuceSFmj4NfnCuSp1WM1Z47vVUEmvhUrYTZTsrV491DCvsbDah/1Doace24u1qxi2Awo
4IEZ0UWAEi99/zKDLwV2zNEgmwB8p1omLH5t//9leocwUwPLNCubjWWWTX9vr1iOqqZiUCGF6sAq
D50QpgnJj2vwJWFthPr2v+iV0CH1nMwC+WcF1wFLLbKxDHOiZyEqsEqgxnrcTd3GFoE2hiN4bdMu
P0uBUgNC2DAwvz7lu3TQ2JoNeXKHGd1FOvKQI7xOWt2ty0AakOpcKqmP1of/HdB+dqWoGEyhrj4e
8Ep81VZ/FDp49cUXxtK6CKUywHJbZVpViEWggfpTaEV+c6kagL+K4Yhfq6qHruKn41n7xVi8Vv/U
ZWzwbiINO76tU8Gqv3gtP+nCgzrfPZXmlQh49nnMbFZTu6oPZ0gSuhsA9mPRy9V8wedQMO5fgKAa
+LNUYjvRfJdqGzg0bd7WPN5fCdRpl8gN3u7ZTijTBj+NDUXFivywv7koPcKrMnuGIFAHcQdtIlJZ
MMMcLWO1EHHGGkIYb6scTEbNdHaOE1L9kQbt2xhYAJNa5irMHslpy+w2Z4Pc3PUenvDrU+Qadppw
P/Ks1JsntTlxImhPfJ+uIP6dTQ/WmC373IbXWu2Hv5h4CRXU8alzjXg0npIrj0xB+QCfUc6D6hyP
xmq2ILJgb/0cjzezkuwHJl9qJpguCYAzbdKchITboy0S8Uf5nBt7I9PaLFu98QxsakM3mta1D8Fl
vrPEmhp7TQkXKwqC5n3MDeO/uzdrjloxPikfyZTr0cdsjx2bUWcA+Lm9O4cx+Hv98wWhTiMYymHX
WoC2Tu9k7S8a7LMETVOA4mPPiPb5ydlb/BZFmcfR7gLM5500y00E5SyoFIbXll1trklPjzi6jij0
j8neQbxkF/Y0kwfMfq9MVoxjK7UQ7XBX8WrUgZtQ95IpnzrhezUYNAzni9Hy1FZfl/WKZioT9RDD
tfmjROsUhJCU6eTjqAMTTy+8Fa/n8+3R6BGt3zw2ciuwZN65hsWeHfaltcLbZr6iFB8xcTAHl3p8
9wygVvvX8lupw+y3xb8XI28rvVWdQuEOUldW5dAok6y5SgVxF8PYgsrMLgienTaRpDGXWVUiA0Z/
0rf6Qmg0kwff3zhhUXOBleWovr390iotfh6kbHl1thhyrw0LDthE4XElVAJpBfXuVffZdpDrgxtt
ihnP4z934KVrSkC+zLdVII4+L/CBecY4dLFUOOeqYm8oJWvL1AjE8oR8xEMt7j+SFrq3L0TSsQ1E
DqjY9WJTcjEkFL+zIQPz52Niu/bfjp5GwGVtWx7Pi1VuTkpqGAP/QftldeLaQEqyCnO4gfbapmUS
QIHsYhGr3zxNYkT+FFxkh+aNHDC0n5ZSUZIb+3MgHSJKEY+OYe31KB7pmlMGHylDGWOJ0wJ/9zRu
qZmtuVHUZQ/XXbyI6ZOWPFLz7fHbr6ymkl7yptLuRIjSc0pae8lwWAoXhP6Gn3BEvC6wS7RQ40Dd
Z9u0BDo50Zhx2TjDN/TI+N01gr/19xO4BbVlfP6M37Xk8FHN9UQ6rcppRECa5mxyhfbgRibZnpUs
LRdUzbb5JrK706jiFFV95hI+V8zusvf3oVVQXiu3c4CH0mrGGL6NoQ8+pRBJCt2/AQNzbNAGYgq3
0iLTo0ynwaIjqmRER0DcSyM2HEwYMF9eJ79Y+Ct4LHyOOJyxa7rfWDcnHkU1KRoL8ysyXAaZYgYg
fMc4rR7DSJU0OYwkg/u8+PUogomcIQEy703whlIvhLbViHssJH2D3FU08+HytvJTH3uq2uixUYzV
vzBxOUv3xjHEWcHQcZ65zjmK7MfP2m/ON6bu0C+LUIlxvCTR1th9zlnUIv5QaojAdHNtEwaCpmmo
VB27P/xovG3uSxJZ1fTo1ttR0r2P7h2p/ZHS/ANcVRgd4TxrTmTpi8ke/eOX1sjGbJTlBMFusOCt
x+B8AYM7/d2HRsp0wojROFvBRTmri/8hjuguBX/KkPdNu62U0njfv+v55Y+0GZHAYpG+JmA+thYF
F6QCLxGy3M77lWxpQzMH+x+QudK7fQEup1pzoBI7bcDr1IM+w5AJrL0Fg9IllsxxvNQoVptOcJnW
Cc+FptZ9cQ594sDlbo5fUIsnessu81Ru9olSzUZEMCwJ4vFpM6JP/V7rMZzHrmqWmiBuX8O6qT/j
nfzhrTuM3DjG3E0tkL0egIgEXN8O8XpBaCnFn52mnkvMihsCqD6zT0JQVKTmVxBfCXBEeUiYeM6+
ze3foy2KH9vyuN7duYjE8ZGboLGyM9iZLIWwmziWzRovszUTTQ/HXqxHfpHw28kgPX9LnJyj+0dZ
UmtOo3Q9v7jUcQ6ReCcjRUKS2G70tw2G0gPBmKV2laAjcbC+qFl+GyAISLWp9avrfuWhZtImqLpq
8AN91Ci+1LW1nj5Xdyduk9N+55V8Kxetyf4fdcSDWLGpJMQHPVmFgzoJyUyBMcm65kGskgYe25JZ
dzKkz9Rl0Udu6TxHrs/NJI2TyBFX+OppzuUcAilCBFVyRWjllfsPNLeWC2cis/nKgRG089HBSgOY
p+E37yUICSQGxxmA8RuN/01vSzrtTuLeZxd1sG3hI8krjdO4mIVsgz3ZdbLoUntc68okcpduwR00
Z2vrrhgVrRobWXK79ppEZ+oQBZyLTznQPAK9aAvg/wIoX6ta2LyyG9VVoW+6m1KTzCLSQ5XS+0He
1kOeruIzgr/KhgEsrRbfL+P/msCNw1S8Mnc1Qt4LtmEuHtcR8B7FaEt4wyg+f9qtSPsm9z4AvghF
3/nPgbBU76wV10C/uOihyNDzQPdejVbTWW4u5/0p0sVbEjjQg1To/Gqp7UL/tvW5j9pWDOGUrbkT
3myf1gxR+W3c1Vbsdh1n+kbGRadd5kNdpQIHRFzFWj3L/vaWAsdbpszZa/dupMvs4CysQJARfZNw
sXlCHzpQTuL8HvMBfhgryFJvFpFaWcGkjZ4uC15jfwwm2d1gZ48z2VhLlKs1o9VrmvmKtdkRhGzW
xmgY/j2TqvBs9nRe6LyfjJeDL2nfXZsrRNiAJcd5R382y8mwZYReA7c7XeAO7KHATtwZGIgyBdOm
klFzOVUj4MngO+eL3qZ2t/2CVcoVN4pDL9QNPgPBE0wwQGFt2BvUOuTt2YtQDkyX6scaP2fI1JQl
nLfOf8fVaOnx5rLtKPy+JsAE2djbIXW9BpxEs5hm03dIZ0YwPR/XCnh4PQnUaqv1V0uUxFtvx7/8
N1fDInNtjgejlfU5BZG8D+VZJ54qOFNjOzqPoZxz4vHqxZ/7X4sUS2GYjTFg9BSLIfQtWxaFOHwe
F1s3Q0qOPxgk7ADkyTeyFXoHpQij6ajPATV9m1CgQLGsojyj5ph31MFoSAt2rxJJvUlkxLoNBSmu
tIzv9woL0mivRzai2MeoYmdFmpkB3LjTt31axMnYAG3yASivhlIT9ALdCZBPsS8ulWXM1KkyIktV
SNKIJJVXNpq9FBEkX2uFlm2K5LoEKAfykdkxEnQmSGn3UqsSV9e5JTeJEXmsdMnU21ESnZZp9/KS
R9fc+ZFO+tjYVbtKAA2ulfBQv79zzT3rUZi8fhyHn6ZxfhpH/Ovh1m4nfrvrRLNlgynMT/trzoz5
cq4eDEsAtbD3AslEggxgKYZN5KnWM5QjTar8dzVch9c0hPCmliL/hpY/bMTUtK+uONQ9ulz/klIy
myWcBJb5akZA9y+eleWB3xMWwuH0k6ZYNXwCyRKV95DI5TR4xjsHzcEyXf9dhEBlo1KgcOt+GsfI
7VURPCZi5EWfIR/Yg0FKkLhzRkgshfdVAPF04PJbUp8PK/YqxnhJ8JTxrY/TOfyKfF41KkZx6Bq7
cG/jFWnuqBboaHI89y9wiCIadSM0iZ2eBrJ57qeFLFXRCriy6V3E+qEKpk6s51xwnlLrApMm/rJ2
pLmKiZ7aPlrHSWtlPqIGOIVL2Zb9lZgehwgyE7NoDTEiXmydUYRivZdgFiJ0laDGr5GGXXHRNuyh
N866qSZicQC6k8KctBRZBJZsAcZLj/Rb1gehGeA3vNlwF2+xU4PJHzSFcZNH0TY0AjCO37Vj9D2r
R1SbpZ7kWTf7z7rbRvaFp0KKG9MTRJCPv9YBlXFKqhWrUscaalqpq0AcbQxq4ZnT8/ZYMdzO3xY0
nOM29sx3dFgkvRk3/WubYsC4s48jtD7Yy1mp01DLHcrXdHz4jkPQ77DPyrd4k4194MCdIQAJcldR
MGMG0D0j5d046WKqn9DNTpdCMTvcbYtYf79XO+RsoblIeNpYEVaCvjCPAlQCZOfepp9ez7rkOQ50
mpnQTBW9EphIc/cuzPFnxlVmrXahpa2SSCLCeAz7Eafm+glVQpeugxOm7yQijH7j5wCuFHSywGLK
zFyN8Kv2x8cOsinOivOxKNWgCvbjVUJi7XJtUEx3egmSedVX4EcXfkPa1Jqe2ob/dIMLckLCgNGa
8LgjVUOzKJxcXxTZx72Aa8U7VieL1SvSspWi/94SKCTEtOpN3Nfm1H/1xmwKV7tApQxPt30+pC74
opnQKmJj9ubp1yutDxRLLh9LzrjSc0RvdjgGSWYX+4Tz9t/weP7C/pTueeLaUi/2A3xQV58Ps46p
Z8Rb8PwiANu+hGLyLikQhstbOKATgZmVoM2zEunGQ+Ngsf+DMGE8cp5b/G2cWL/fQmXTgsdf0B4l
SILtke5a/Y8LLGWBE+xpCx7b8ijJIwSTfvqXrL3HcLrXDzOAvr4lZyIXs/DQXk4qNyrI5eGQZko+
Jaa8K2ihPsyvCZhEIDv4Oe0+aJnEu9+31eiid3n6dxJROLwKgHeez7BHH8mC6ZROnsMJcu1+43l1
9HlIiIa99uCZuLKOaDma8PrzvtBcZA/nIQg3xxay8FJ7kTYd9zrqEN1oEKNTJ6XcdFS6GtJiwVPG
2zoYhCgKVCZ0YiPzq4Y+EqdENdeDoNSh1p2JydD2TpwUmABHmuqzKPWArpSUheZRyR+fbOeRTrVk
1OMZbjdy3SHAvs4Ulwc76k9/GDa+MGKJ9VTcScorDEhhg7fXHsJYGRzy8KNK1cnK79wMs6gcZcSi
ciJn0YX67dZ0mqO0OewRRQ1pENCn9R5Q8WLwrt6mRgzSh4ItJ75f5/Fb8QXOLFyHueAUeBiveXwH
CYa19UBUC9lCVGxAUYU/extHgujBCzTcval5iOp1RZLAqHfflyITeNz331JULn+0cbtO9J8W+w0c
D6/y9Tj1aOik12b5IBfWPPFNyh8fEScU058F6oBr7UjIEFR2Ds1uPkL7KOF8d5eW6hOab8h0Xeot
XHPuvOnRljqVNudiqke86ngPKBN5LNqN2TQdP1VYGgzwiGnP7zyZGwhHXBPo4C3kdjAuVZTc/OgQ
Kt0EHfZywzGBnGoM5q36WmiROs0lAKvsb5dp3ZAPGUFxjeXbiiXKEo72CYGOXNnVlAjZYlfe0J3m
bP9gG+ZqwnNqQ0bHqbsdpDEtPynEqDo+pOgsVNXsSQOyaOgaipFPGjgqQBQmLVfDinAtU03ubF8H
+mdMgUzlfGRqjjLfi0I8sVTU2lEmm0NdoqDqMztElHrxRxvloDkeE4wf29As8xuds+Y+6TvO6rKw
JbRd0Qvync0Ij6lN4FdUd20VJ9VgAYHnf57HT0luQsEDzmvccY3w1it+FZV/X94MJaC/VBeOTiG0
GIPTA0fhrLFCkv7P1gCgJpiZNpES8ySxSOhMuTGjkfA0gyztcDWtwEwSUHpE365Mn/ujcLOc+JeX
iMhR+fxgAI5udOSV8C2hqirP3EnGqG6n1xo/9pmdt0s3mLcL6YsTUItDvTKv+ib57E7JtNZXPeBt
C3X5/54cJIhuJplvn+BB1fAdFiItcY2qIgAWkjaCaXRHA4LC5yDYqPiRcC0fL+OSdEZrg2e9vBs0
u0tOMb6UGE52aAY8I036w0+HmZHRy+ZvK1Ru5/pt/+Suxqw8V4MyFpwtVdeKYFKqDIxUIttB74gP
E0CJefbgDvgSbtU/MoufJSi9oCdZwaPDhazlVP/Qvv5gOAiVDsUwgNBpv1C6BeIN5Hel7MQlECM6
n75B8Vy8Mo2Rl5zZAHCcsRA7Rb2gw6VfOXfySx/GsmwRpeYdvMdvtvY2cceNxnECQQz/4qv87G3O
OEanTcP+b031dBy8xoc+VMhnSJsl9VQNoZW+cOueUwc29CC0+FYYhSut/IDlsh753dXCyl79+ERZ
tdqKPjiIPtCNzQXujiL1sFHQU3Z2takAVx5wmJaQLEjIWgG0XJlRqyer9RipDNjrsYBoYkT4Chpp
1nWBi4IBUzaDRDqnntwyuHmiUZStAnsTdgG8LIBPt0c4wpebJzxdzl1DdwZRFCrC/N8j0tF69G8P
8Adb+f0cnlH+44SrMjT1IA1zS5dJgIRuM5J4jHcvqYdjxQSbb7i8UErWl9m3zx6PNT+U2eoRtEQ6
e84CJRP9/K9qdtWMyKoTOvRj7EHDXa7aXWiMw9mvGGfqG6zMRm1u6jwfbZkNUKo5kSMDYEWz05l0
KNbu+V42/jTmT0mJiPgjk7aqvDx4U9lt06j8T1omiEdCP872zE56FpBW1tpsdgr9eRILIBttL0O9
a7Fv8JKyLpQp7n+V0ZQhp9ZF/Sj0gDt+4i3IzUJ6Lp/kgo9AM5T7Q1KenHhV9m3Ea0N0Awg7XY6p
68UaDSdIzM3z+9hpE9ourfrjZfS0vNDnhLbEFf2X2/hvgPXfPUxLW5EtOHkTMNULPPzh885TCmEr
Um7hYMPukw7La3bynP46ro9wy0GK2qF+M/7FBBtyMhxv5MOAShBf4tvUTsHUqYj+AZqPl4wbJv79
Wvk348aJ1+oKRNdMW5XgS4okY1IMApto565wtFT7+he3kBLLqYkYsk8ooUgu25lNVVADeBcjqaQ7
m+WBgcuMxPOlLN1y6sMsx4jS/Nr+hNMhoojBhuO2HKyxzkxyjnutk0PPovpzgBxhiw867x5PVW9W
92ivePtDl2djoNF7sBwXeSiGdsTSc7cjXxsOxVQkLoE4RxYKifiVRAI8EfDSQxSCG6cfKIxHZRGd
K5O6qvsROLPGa6xsc1QprctxA8f0GR603KI1bxt6nN7fQmvU2UYGvYuKzExUMnIhcPVFCUtEXffV
ifJvE8TMGvJnNhvl7jSp+Y/5Hm0IpDxviNLb6+CvTAjaKUNaCU3G1Zu3veu/rc99krBkNfBQKFTf
t9cZvKF76BKgD6+ebXhGapRNJy0r/GBU13lHYeYUTdKJzc4+CjMUOsqdUimTH4PBn6Pf5giaU5Vo
lPMfKUjPy6DwNdBfmGoDCvv+dYQQdcwL0bNFx+KfCyzxSfLKnWcKYKaU/0UQdMUbQUDaAbOu61Hm
xU6DQfkytwdPCM5FP5SNMB5I/E2tRH1qXNJ2Swd4CmN3NsokTzbJ91iW61ZvFdAPG3eUSMCWeBNg
4vg0H9hHvn0R4vc6fugTWEcffk3t0v9zlK904DpYPkDqtOfGdA4Vhf8fq4F8XYfOwAVhAwtTtZDc
x64+8R0mdjQFOA2ywzXMAO9E1Es346ofIhMwisa2A6W6UtmmbzHEqyuNpSOGIjjvL3c+IMMVbk1N
VBterJnT675V3ZmYCN40Vp8wXsZQRvTHgiN1fY/pfJetSTFm6roVA5nas/cM0ttmIdFhVujvYMEE
uSkuiToxfL+wOiZBXizw1EPeyAdoPQ2ZOD0Ds6hMMDAyOQvmzzcnlnslLfgsy6/ZajIo1sniodyw
GR58tyir4kDf/S9mQyG+woo2QPUHql0cBslWQPQckhYfh5NzmNKgjpMxYkYhRSmjZbfdEoxH+AIR
YPONS5/kK30JS9ZMaB/I1I6VTIWmEo2d7yJmrkrWgArGZm2SpniaxUTXRqc0eVziTXWEJmbgmZMv
QrvbxvWr+IugSRs6bAOGdDqImSQZEOwEo2kqbqcedglj/e+J/rfAUh5fjgibjvWpsOeb0aFQNG3w
eQUxykn8Jrine0torSA9EbskPDJHhMs3scgfBcYYppQ2sr8QTWqs/8NVnB8Wj10fZP9QD34Su777
/E0zbKN12WnfbRisQDiz7Y98YwTc5UpWFgkdDKHIuzlenSeE1pGQ0v45IN7bvZsoFHoUMIdkPB+W
k1w1nXO6uhvxR/dhge7ao5Nfrwgr63P40/Vh/MgQoiMjESrllEGXD6g7sZ0a5qz/vjbjRiZrbP6p
3cWJU+Z+KIP+y8gv5JInzwqd820XK09rebgAEuX6B6u7iCGOgsl1XIiNUylQ/NxBeXofuupLYBEw
YbpBf0wTP9CjDICmnZcAiY3fWNZLDpBYHBVb3geaV0RXM6FwT1KODxo3F3u6jZ8KzRwAGL0q9Q3c
GVIceqSmj24ZwVguUK7HrQXyAW2nn16SbCTkLONjid6oNzOVvl4/FK9ff8GsTIFdLKc7U9E/bn0O
m7LOcagMLjziHwk6xA0MmnxhibUC4xNoHDP7RgvnptI+cLzGQUQ8hywPEsRvE3jP5pFTVMv35YiG
p7WcQQsZYpbeg9yM8OtXKFs3/f4fMy+ZKTqpfC5Mgk0nmYeJf5v+P97wXaNC911xbZr8Bgscmr76
k0n9BqjCiKo5nQu6cLeLnn+YD2Y6j96PouCkxduuKtRd6Ob6nY7Lpkz8gkYYApudhAXwC39yDPET
+ZqRxe1E/ZUyCSr90ZLr6qZCUSn2Zr5PB2QvCNazcl2sbKW3EOQu/JvaUCvWTthXBJrZv/+XfDAN
hJ92s0tqASzu8mpjapHALCiMFDKw4P2FBrU5mvVo9/KwH3r+vsOHQ0bCJLTuDXWRnIK8azFkY+M3
I4Wq3AVVRQ/vyiJDK4fT1b4sYxw0BylWEVsk0Z8IaOAPs5gmje7KIaze9x5BISLd7r86D3qomEmq
Ty6rnPoenBKaMjHkZY7BQN13TXbGDunj5b8L7g6IlWuk1UtujXcbPpag/srvuXkNqAFXlJUh5+gj
tvhg2fpzRSUVg92ftv7pmVr9NvX1bnJUK/Cm4A52Mm/Yo3ni6R/FQTjGSXYvvjkC1DCefbWH2G3x
R1V6RWiZo9O/e6iI76Tq0aGRpVygI7f5RVeurdElj3ivqS+sfvGkzZ3+/ycvuwGx9s7Pic7sKGd2
iIZgdXDNbKeYwd1eD5QAGRh4q74+nnRrofwPu/U4l/+/atiwAtqvol6h9AK1F8LTT8LyDiSjXBXF
lPisDFZX/xVlsx1LtUnLvrhPNCpczzDJUgnTZCdHTPESGtKj63kagOLqpElIsjGO4LFWXni/WP+O
KHUsvfXAMTX671zYSUgq/D+vRaO1mDOcFAOQ/lXyEdnIlpRk2PU9Uoji5agg0G8Y/oHbFWNyePMV
94cIkniC65x7HaEtfIytHKNDPSHsOli+7tdgC7agyV08skTRKY8TV2zNhfb4WYXmdY7w2ApWleNa
ao70beaUTAPG1ru5l47kXcCZgarh8/ZJOWxPZKHezlGT6Dug0EGQcJzG6H0cTN4yKYIXw23N+JkD
DqQpPlemN2POZ/in/WypO2VwfKQe5SVxq8mKOXcmlw9W4ECUNefL5tW4uZCaLTt7ymo8DXR704hZ
CPJMhoR/CjZrfqIP2Nw6I9zn/XPxkmVV8Z53AdsTS63CPd+fjD/syLIXl04GmNjuZDF4i2TZybNc
AyZ8xSrrI/urFHzPOOWlVGUwKsyNOxeiRMjJvv3PTbrHryXBkfdKPFL4uOSCNBpVqZl32H4WrJKP
3Gb5SV2LIW9NThGaqf+T3GhfM1rKh7fqmdOCdj7i4if0f4XtmWyJrEq4Ssj9Zbid20Pv6lu6JJcZ
pXmbctxUf6YG9WcTV7pQHODKOj1uaNVBPqk30Io776dlUB/DNHy1nziijnIxjPV2GaLw0tpptYYd
YZVR+vJP3EcW+PFR/lFElAUIJcQOpvmHHrEY90P+5oGsnxbtTtTnQ3YMM0R877pghp3HW1tuLpCG
M4ZjA/3yI3jzZvrDjiqhAA6GrVnJrAWsNB40pvkLtFFWl3yLtvSHjF1o3/DVgJWYQaDDH6Pyx6cO
N4jYv+uHp4L3eM+j0Gi4cAsxk0nAvXf1QeF/JxREBYwfLrcq9PwWAv4V92v7b74fYNKSsTAwvlDy
f7/7KcLgrh4QcFXhWfzOgPlRsye9LRw+EpuROEqHkwxjB6WscS/B0ooH6JQb8olf0sDK9m3D95AM
a42sKZ6bfHeV5JNCn8vALxisfhWzrP+sKlIuyLOmXpQJzKd4TAuLKZHPG26+jqAtAvDgiacKxpbo
GeDorNdGI7rN4eDQeE3D3OLpAa9D1pVA4Z95CEHXq95PF6i/zrUCL6ZVF4erSbHT4LBNGTUtmfVu
AQ4YMxnkWWf+kH0pXtLstzHFTTQ9F0KPk6ywgeJ6g4xpeDguXOyFEGJGlyKMNmdob2s9ZaPLparF
UDjEVpvXQJ2FM2H3Q2wCec/wY1JPgpOyLYKdPzxONlxNL0TZ9dSHqd6C1p8vNw8Qg0N//xoXaO1L
rnKEmiH+1CGvBc7lT3bOK5P6P1jF+cXqJrkOAViFmqQl5Qot/scwAn5eJEMngpGcCSr4ybQimVG/
XKSnf7eE6dj3xtBnB5wAA57cqXsM+IvrnMLds7cHuxMinmc5mgOgpBiNh+NJj0gBhuW5wzokB0Rf
noEgySkmZLxsZGwCRL/MzKKLNVTw33sodoQE6hNlywYSLgMVH2Y/0wBWJuTESj2QtWQwEm8ZC8xr
1AU1RkWSoAmXCDyObt20XmPgpz30V81Y4R3yxx48t53pIzKyUt8pA2M1m/qmw+J4s93zUSuygczY
IfPrXJJ9hl5Lb2QjHlAjVTx0e9P3kjzf5PjL5CHZktGcoQC/1eVMQa/SVKVHM89/m0YwDfJfq7z1
XTvTUg/HRxVCgtacCRYcF4yQhXw1UNMVYBERCxr3ralboj2aejNlrmcJdyD00RCCaIwekkOomF0t
c9+58RrhQ7yw48tOFYmdG24HsfDTARjZ/sZm5zMMkC+Pwup413c3rDcNpyIGmFjW803KWNNMxflj
yj7kLRIOIc1A/pO++Pe9qL/SS2STRtbmQiZFMp/hC6tg/NDLJ0WLFyAidXusAJ5CepsfJm1XqqFx
RJqtW1Fy/eLuEcQuONpT9Hwv21Ad8RdrxtnVo0zJOEuaOSmCFIQXsI+EGN6BvooTSRWiuQwuDF8X
0GeGISq3+RMuDdYZIyR5Rrp00uPI6Cx+hmSH/XMP/7qbegfbGQAv3LelSo5P3LJscd6jhGdYCHhS
dz6SJkhpR50LMAFV1TrA+MsPxj00B18UpdGU0p8X7d17Eab6sY0S+KbHaQYpeR8nOx2I7mwUdeed
uGJSuyLjq8GZu3LQyZzEkFgtukr+Q9Wu7r7qQoEhMXind0BenodtUYUYrZ0VWtyowLJS4KTnrsFq
GkxfaI+UCxE4k78/Uf/HA9jast9hxep+DSbZ+IgQrR1+oqgnL/XCvkSM7ggz9YAVeJH0VJEmvQXQ
6pZ6MAwwgBbH/SKgUza2IcpvsDpCIK62QsCnu5aNpYy7UrOFWrd026fKNH6DwAodeb9L0FFuk93P
SO9mRhiN8hKRXgOOTkaVqYQoD1wnliuLkaxcnrfg2+PjD9nQdeanjsew7npPoOPmw/Dz/ELshUE8
jmwJ0ETJigVpBHVU/TZt+t3gI9EL14dhiNVAqKvuKwELFWdEiYXi8fMoBCLMi1wih/rPrJEDARES
yBYzATUxHVeKw3QRDUXWXSgZIRizh/P0x+t9IyXJWAV2ZumqV4Z/h7yTmhgshDc0cc6RmNPSFNh8
SvsdtJtzk2BEeFKUKZF8hrN8SbqODrOfNOBxWky6XGuXFYVd+//VNRm0qb9NeLl+iwbUyh/hVZcB
DQvvg9dBGJym2zaA1eCQVWw+EuF+PpjOLE5qHmMwds047dO93LOGU1+TWWwRW1OhPzsS6rBnJ3VK
Kr2UI7AE0OhWuhFUq/jr2j8m0CY5L0IGO0f6h1CV4mvYmXQkEpUXme516GM7yRwjWB17HQc/80zd
xPO2J0Y5ecaj38T8x8b3ua/jaUGspg2/GDKOa6bGf3qLzInt6WMfQBYJxFQQpCyPDlKY8jWfQD3B
LL1fhj4kgb3Y8JMd/Ghpt2ZiyUrvcK/Q3ySIXcPV3ijyYypbw4AmDKstiqrBjNxGMiJfQ0MqSQEU
R2ORF7j8d93U340zJ5x+/UWEUx/f6yeOkZTXhNk8H3Ufp2l5GXin9xj2kI8yciVjfN7Sfh1HCSux
wVajWH+AzuuRglG7mSjOjBnb8/P6Lx4nbjJnbGrKb1XNT8OEZF3rVSbXCexs5fkxl0GcCGiLvcpZ
in/DfSdpVf2uO9y08eR7u7NJnKvvUdrwVezlTDhdbjZSnVYw3Kro9Vg3xrav2MvwKpiqhZdGQGy5
6hT1GViA5GmdPBwrHFQa1U1VpgLMfnIQxM5L9tVdpxyJ6/DFuzmBV0GGxPsC0aYiM5ylnZA2stJX
o0jLp+/AP/X/bvuJ7YrEUKoRpklwCO/HFRvVdG8M/u70+6yIh9c3npSt3lM1GiCql4rcR6Ke5Mw4
FkfAgFw2t3unASiuxlSYOC7iUCgPQSi3fSjdJIRDaGdYiIl5elVYYDkOpjx/30+lsAZLezCPPVlW
CFfqZOP/UWFmtsNoiEDvh2w4sLhK3SxY/3ai9bXn3us92VmmuRX5ohIgs5NhK9osZdAo8cKFU/fE
x89KTDMduYK551y8VZ9TX+gcHvcwp7qqbS2ctA0HbTiVkSS9BtwreOLEp1BQ10yvpiCsRFm1iIqM
RWxKWEWyrO3u4fwk5HR3b5r841PyMS0ZJB2MeuZAcj+oXieZvXtwjPCrz7Cbf16BI7XfP9JR/u6L
Epdkfm7d6kmWkOVWbLNDvk6ONoo809PNg9SLPu6A3CAeMX2KCsX60KLQBCURdiKK5vKGFCTtjIFZ
zSFmPIXtkLB9s479FbCE1nAIgojFNcQvXdUM0lFPKLxCelKptUyiLxZZY3DdJP2xvuEZyLAOL+s4
qQWRofbWkvmqq43wvnNYMUqjg/xfUT71lSNihFr1X+WsRN7kE8edZDwgU9+E84FMu78GjR1+tY/Q
SLPyEaEdKwKg2pcG4LAG+OBn28mUtKZIIXq7402CRx/26BpGdzSXad5c/IGVnE3UMzpO6DO8CbkI
uvAOVJVfdpcMnwiEPq9TEbwY4Oun7RSzbKZK/6YbjWyfYFJIwPXAlGt2flm3XcUZpaAHVx9HJ6qu
EbnkIjJNKGj52L1LzC6BMmjzcWYPWUmnWPq8hQPwepzFFHV6ujUgjsKJ8NEa/iGop7JEZ/ll7WI+
70SOqemUimtLW5oR9VxfX0ObnwHXHA/9aVaLMGGv01F3oo4U7g2S3oLyGuB5a9B3r0ZVhwYyyAaE
XhP+iK5JYOIUuhEfqLmkFFEsi2ujE9qD3b3Tcb/P+BjWRqwD51X4dD0LZTyWA9zne8qnhQp+ZNZ1
D4Pv6tDPOXYuE7+B4y9s0uiByIl9xn8gxPUEjys5UcefhfSku63xnXlibKEcGVoqeSn1T4VaN8hz
zFtGrj6LqraUtfdpT6ioOX8e+jVpbRY0YgqgnA3j8OVuQdWMe4U9EnIulPVrOObyWyRnQCkaOfwn
+gVc5N18Mktgl8jUJ/Xq/N5yvvWVhzKK9yS2PtYcRyF5ppeLTk37V71mxdGXx4pbaEwtm6jQeXKu
G6Y6/HS80zNMtgtxVqw5jnuX11a0iB/NB3+4IUDcJyiAyumEwOslimgI1jUXkgEGgzYkLTCrQVtr
N2dUAJ8Lmn4BnhOtjGXOI0xfS+8x98Ag99AwqtmBKc/DEt/z8cD18cvJLkbjy42WCIYHRbWo4hHI
voYCIcc0iWhlW6fBr3q9ke4BR0vzIBIms9URV5DEFE7boTItDm5uu1fOAksjLc+/GcQmcF9uTyqQ
ztUWEhIRxC+0RJXRQyB76ica1fThp6qusmi6jTT644GIhvrtaJKbQ3d5GAHF1oJykY+Z8Z2yZQyj
NY1QeKgNMPU6aWIuJ0Li/cO6LTPwgMiZ63WAXi4W6rXM9X8O3K8B/0GVFZlVs+9ELAn+WFAA3LML
zvnpBh3mSxQE4jCEdLhCO/4IsVDUvDFAuQtPUj65cFCgBSfSfPeh0j+ACGcfcm4I0fd1qmVYGMTt
3dp8pESOdCTHjoXgMSeAfDih8Yk5AFncUijoQHvR++iEt7rbp5G3jQ8uGdOFSnxfiw5uyzNs99R5
n8Nxx+VoDSJnwIrLqY87vUGBiABo0RuGr7V+JAAckQP9CfCebWN+G473U2tvNJWYpxmz7teA3nPa
P0gMDR5KGCSkXaZ0sKsKEEDx49Q4API7ba6PbHBlT8xaf6mEvXOtNHHTwWaItyOJhLtx9UiAzBxH
orG+IZRxf5NPEgjrAV2LTTZOuiev/O6KGSuRoTBUe6AGG4+jZvRxqumldEBtfGccPOQnLQm9GQhh
K2D6927OPfWM1DO5fgKi0TayX8FFXQfT+JxjCPXgKF7VdtXSoqD9P9afhYY+m0fkYL2YT2T7T3N2
zOSL4ec7ictmlnma60+wTqP1goOvJYZOceoYgmV7j6yvzi3MAtzXWYtTOe9VkqwvV5oYKuRXGyKO
fL2Ym4vbFoMfPKdkM/cHwcVdZj+nJK8wgmBxmm4dth8ZgvUXrxxA+mEvxBZGmXjaxhYKZ7lgBAfJ
vJzNbdlKX4+XQsiPwqP9U5KvK1VyGTBkGKvOXxhpdGl9LgMcPErBHMFIcVkNOczjEzsW83yZdLww
dlAxF2A+IvaS6qc/hRV/5CjcYgFAHIZdk+Bw6DeU1dtTK/sRd8lRk1YaaXr89bP02fJWwwnRf/Rn
ai9xdN2xmTLf3iMCedZ5qPoK8TXpQgyvtFjWEa6Ok97F9GiRcvGx+OpUmcsYVMlFJTsFKQntaSZC
ma5hyRRF5CYqSy1J2SBpJkO2E71pJ2OoKo5RPuKCcaT7mUyam67T+2jui/peOXCPxBYtrAX1VeYE
+cXp4Xga32lZ6QuPSqy+02kNz5oBAeyEZ1y38H6xkSAeODyJvUSgIYMvB7XTKsJvXwcLEZd57znw
FHPGrzKk7iIYtoWKZCmbfAf6JxjC9IUxYg9m7LpLbyV0uLD1GT3WlgRYByMsdS1OWunmHnPfg2nl
54Ty6EIhm0ZfiPO6/4ov4hfCs0AOEp61zbyEtqRkNMb9W6PrfXrZBjHCEbWRruhjVMa0/6mFYlDu
QRyKXsZLPGCkhmLXkLvTJY8CrQA2ZXQzBjYi9D+FhTdHRvOZ8F42CoVv6StR+0v8SJHOY0pdwUco
7X11+n1pf9YMx9RkjIM93GLFXMELzQh5Qvgi110wpHyBZuyNYhUB/U6CshYtfwPbgCe3nhBlj7+G
0JDBLPwCJ+GQYNzfYnjkTVFcmdfll/Qo/Nn5WiSzzQ9H5tpwSRN0N2t/YgrrySEU32MWRWmyrr4U
8NGW7mhQEhACMvK6vxSwkjEsIh8TZMqRkcvHYzAC62jl8fXO7RHINzh+lBvq2fBqyYk/xQv2pq01
Cs85UoP4Fbt35hgOO2kh/9gSiDgYP53CbUDPpPXH/3ItZt9dYzkJFQewGovcX1R3TtiSIBBuQV5E
K438L+mt42MY6/V89xvkJEIYtkLTRB54/pN45NsnJBOfNUI/+vDZAQ1LTKjPnt6YbAzWQthFDbUo
ouqMeY1obL4OOQILKJfbbvgnOTpSRckUwiH96bR7QLZ2xFhDWx47gQM0gPfDB6DPO4bzUjt2NXMU
4NNTRQ1owRi/L/HdU5reJJDF0Cs9GoQN5nlwoZ4EYRmd3q5uIrMWMHGaki59SDOZljz2rC1qsnTJ
fTdgF4HkI5iMFGSWHJE7gHy3a9Ur7dMurL/+qRuXCn3noJ1Yf9EU+CTO0dgLBBzMy2mFmEAaYjTa
LMsIabXWm61S2nddRRibXMi0FQMrB6O91cRROl+G2NtNzNAAWYLaopOTY7Dt+HC4TL8RLnxj/aOy
flRLaSQabxnGyQSLwcAK7hlKLymT+tcnqVEocK6+2RlErVXP01ZKEXA96HKsfWQCce46RaZwlOTi
UG+RXM3Ph36Rspjp+s1RQZXae4prmajLbddcRUO/BC1qOzQYQrwDX5PwOJINtvP7y8D1KCUuapfQ
7fvYXPNLry82ToS4eUz7eUmcnEF2c+7No6w9vAH76Jt3yXrbGft7D56I7Z2ZAEzVXiZY+pLVr26W
EiFSLbLAuNMLZOZ+vtIECN1yR3GZfPZ3m1WGzS8nvBTOsq7rC6I/IkLkdYyKfceTsK+ySQSM9llE
eNX9K0eoT2aPsodh2ko8hzhVd9LNkfV5c+GEWLvhDpPslHL62siK7aasju4tLRtuthgdCoCDY+lj
IujIKMG11ymwaoJMjzUOHa0EcgpfYKE9oaDHwifJLdoP9GkaFBhVXdG6TtV4Wyy7WZ1N/vgsKwAY
6W9DmNij8aXY4ib9Va3p5CbpQDU+5ZQf/p6MusbdsuEjgKcMrTtDryTDyzeNJmkNmqf68HbUgNIV
x0mCApHR1rnrKtrMUrnXV7EAhG+R5AWnyxjN6qtBnI8PYznEqzTa8NAJ2EuGbcmuz722lTym1zEu
fMMbO8NjHNXvcVP6Bq4FMkMiVpV17wzVu4PqHj7BPDbKg7u48Nx4oPGMLVx7azZT5m23XU3Uagoe
lnnLlYtJ3h+Lk00l7A1v1a5AL69i72zoRVePTS5H9lGC86taF0iRTxugaI+GYxvDCkIqy5EAT7H5
vY18gB4a3zi6bgNfZwssXB2CmVJgAT9p8JIGDFju2csL5vV5PDHTV6AT+P+99Zh4NKsNvQLW4EqD
V/wVEYMqxALJVbVaBiOKhT1WeyTwkW2vRC0GJO0xD9+HXiFGtzU3vCRQ22RGQIBip71FP4+PvSYk
szyCrLejKshG3tuq+QFeuBTQdCPswzeDiTr7aZCph/bqaoJkjSEibYcSlIbBryHCwM+n1UrzqzNH
34IrHR6A3Cs847EsfJ2KiPWmOz1XQil2tOoJFtLwYFXb5C0rqHwn37YFOiOqeUstdBgYjNqLMi/6
YkzNgfotOype11McisuZI57uIe/FOMVW72/yw5n8L05BG7UTAO8Y1COR2qqsk9mXRLG75vhUzxEk
TE3GTxs2Rk5IOUV1JdIQq9JgCcAULtA5DwBu9sgnwIdsqVvvXRRQ3ex9N7fWCJ8hNz3i/dQRpB9g
UhOBFszmCVRBY+LyhE4u9xY4bo3iAenijC+R0XZr1KQObZ0kZ5RqGbywKCqNYlzlMFxZXRkapyzs
TgVjrFjepYiJtDgFGLzJ2VKV3T9z7qNf6F8FTWkcdn4+i/u2cqO5x2z6TrHlHNLyNvGMnxK3QtR2
KugTEl8InEd4UpTxPoa2zU+scIQlK+LdN+n0rEkPrs5dfmSz2RJsYllqMSvrwb2N61qdf+dSeAjI
xFEUf3wyHwVQdOwsLPlqtUSGC3Tgep2ipNqgfhN7vy+4ed1dz0BUB0fd4zFl2bjvv4LAUe8guFFb
N0/M5oKDU2EKQT7evktDW3fe/WXazkPxqOJk3u8h7GbJXdZ4UDJ10sh9zG69UGD8thzmC30EhCrR
HKa1hLct5HfNln7nGcDO8DJtP3ap5NWvgSQalKiAE/Rs+sjLYUX3Hu9EIDziFa57iDCT91a8hA5l
fOns73aHwJnjhjxB97Q7CGYInKfpUWLHU4MirGO/lV0lMhveRmiGs7yAN1seJpyI8KfxuODZQewE
nXSN+VK/hYybWKqHem/W7xwYUu65wzW7rV2hYfpL9AQ20DnRanFhUw/RJdnomIpMSNMpXTvxokCW
SpAL0AVT80XXDzaqeG8dxwDT7A8yTPzeQcODxvfO4gtFLoHitcDts0xdcniXs3GjeDu+mLDcHinf
w8YZz28SSUAJdLNJNEpC8VG0hSENjX50yy/FQrGy+UMucSq8vaA+vDsC5atwJ3lNbd8TqmvDG1/c
3I+ad7uXkQmvqLdiAqoDI3WAmW4MZ2oJiEaPNEA916JFsTLwgEd/Bu1H6o/fzeR/pU5yejHJZ/jg
uEjg0nvValuPRHgil0wybOk3IBI01N+NSAKfxz4ikI2pVfOttXyn9e4FNpns1O0oRNjRGwnNcUH1
mgB29xZchL5edu6E+Zq0odlu7jrh4wVw46U4bCliI9lBfr3O2bPf3owXu0ndSSI465ra3uGpiGqp
GNtPOoexe1d04KOmen9g8Ee/5pa27jQxuMDnR0/9QBmK5nFnTb1u68e0klKs4wAKEpWIDByzIybE
FXJVDJ3m4ViIPjwma2MG/bgyenKgantK6PsYtiS82+N0IJNJGTpJXTysHfePzon5vFVYAUsYUKv3
GY5lxwH70vTqxTd6KXdsrl7Vt2Y//7zCMkIiXboQFW3ErlVe1A4SqiwNc4i6m/p7CWJ0QmNu9k7s
EH9oRSo/vdNc04hoXzZxZFQWCVJXowdyWMkn8Z2sgdnvRHnKXG9mzaZx41puZuNA6VLU/2fUJwF0
dlZvzrI34YEv0JWrBx6T6kWzwXjSq/ir/Ev2zVeDS4PBgmY6PPvTjFoK/epa7ZjQjlQhiMCdaRLR
jXg7kZ+e/xLaeO+D9iBc7XV4dzga+BySYPLmZEG3W/FlLW4YmTktU/GHukxI5tdLMWRORzKWZqKN
I5FeC0oARzY9ADi2CaFVM9MxvCMsucXPqU11RU7aXg/o24fjrOH3mGttdLa6OXmBCz4Cb+JMpJJc
ig5LyNaKl2mQdikgtxwRWoCsSsU90zrUBXyC6xpjMfH/uuIgKjO7DaouzgcC0mBYwskuayx37bvS
ZRTA1jVjAqhG7LnSAujnoPcMxru6TKYDUNUKMyYWcFbvw4xMjdG1C6ty2j14iWH8VNSBKevlly25
gMfwPW3Z6kpeSq9r2B/nmOlVa4GF5gkyolrjnZfor/kkMWQgaL+b+ehZZxdpaXx5UeLabXadgKzP
h4IvdVLFlqSwaaH85gtQ32Rmk/I3+v4k7e9EONqboJ+9Km0iDOL/Vig1qpBd32ZKdGuSmopuv5A3
zgCEx3cxiZ9iFjuuxEuouwSdIHL25PKr4syr4EGPqXALJMzbRjdwp71kqwBPF5xNsZW7KXF1MILw
0Sw/cehAVBdB+OH9lVD3wslhDkXr6gNR3SvxUm8jO6teSvvrMSZM4g5WrkwpvHXm9kYkj3rfFLHp
jK/lQ73yoBRPpbvKfEu1tqbtKP1ERi6yYobmgiC9RIyJwKMh/HfWdAhdTeyC27WeikVf5jVAd0M7
DMHxMBqwLyjgxgl0kiz8iCfyMuIy/WkvPdUE3wPwtmxbiflmtaJ5qfOA8Tnj8F8jpLNor25B1q8v
3H+DwxedjKjQwBinL2egAwdd2QoYyeFyBTVmi5zr/kaY87IpKfmcjTQt2j8L5JUJZZH5wwqYpRXW
91uOCJowS9ysgMxWc/eqL0nG2UzqiWGb1UU/wDLI/5yd0Xb2fO6kl1QkXkZjIBWu4IJR2QNKHT+u
4Jijhq1Je+h0JMLZmJDb4e+E4E8OHpBO4L+Boc27QI02qAr8AuCulOZnNILEm5Ex7am/SNz+JM2f
x2Scj+JLFKdTmwqgyyf7sWq4v8AVbLUC4wXg7tET9Vz0YM/2EH+n8sYFUu0Vpxipdfjecg8BZigY
Sn7LI0wrkaCOk4xEd7swgtRZJeBxjQFAJjTOXLW2+4rimNPcjngBK3ML8wB8C3T9KctLDuofzI0d
TKskeW7rwOAaRqxBo2OKL6CkWKLR/4QxMJTm/qic72Q3+9AsSBTAqHEo6Aq1LtTOAfpuqqqX25U6
uQdXtZLkDWwyQVBUy+Zr+KG/DH77SC16DAsUuYzk8N6Zo/7dsf18MDlmcxBHUVFDVsYSlRLswULP
kw8mbz2ZlP0vpxu621xTJdIy18mxBAQ8ZP/zn+5Z3IIrYeIMbpeNrwby3i5hvuUZEjo3LJHw9bKE
OmAiWQs018knkKpATGJuJUomI7SLjtN7BVsQPRc3WClZnpAZA3E1PAlLKxq/ZEVcDeAYP84Pem7F
uEEK3gc3cRrOY0NLBlSbrmixHNUOs6p98fhC8c2vgcIO6ralY1viiTvaPlBBZDfAFi0pxQ367zwa
p5ZYZyn3wzsOb9wCem5Mfo+dHVGbOsESgGPUwTFUbKufKEoKMw5fKJDEW7ct7Izy4EK3gykcW48I
WqIr8fp/2ia2zDxO8j1gm2EouxbUrs5FJ4VOqbtsGln5UfshAkiNQ2QwYIJl+3H89J0o5hjjGSh2
s5Mfat0CWeTPhjrkbww4sA0CIeVhADPzWdyg43H65H5b+E4NKKOhAedPuRXjs7MMskfUkGlzyC83
d8Mbvsc984yXUl6qPAikCxJWwYNYgSMCQ8aX35XfIRF43OOxCUPyzVYgcL3f1vgLd9k8r67Vd97v
dJs4REoIkkfxGXyxAbz1qZdcqDqrPWaRZ6N3jW2TwMmAx6OBMu+0LQwmk9+MGzvD9V4Z1/cO5uOO
pqCx1q5rRQMIV9gnYQ+jgONAtseba9P55t7A7yEPFybKTX79ilga6sLXBjS1vlnqehGeoqqroD1Z
PPKNYzMqtiYZ1h1wD9RY/R0yyKC4uAp02aD4O3tJZi/M+LGwILb65xPaRu74hLv63ZlqJzLQSvEq
Z3M90zpHeLV8ahMdKLYcpKJj1PSRCKTO+5gcTA3G5/mNn//1AbtBcAT+L140/DrRhcLZhukC1YZ6
MIiSNKX7iPlLc68hEwe64LHsggbY5+5R842lUqms3zWvTG4+U8Uv+6EtzM6lq13gJmJ0NfYycK7X
pXgql7Ck8Lo6e2bITiM0NB4oQXFeWrwFaDSIFnFlBZ+MElYVVh7yDIl+bKTCRmTG6ftib40lZYbS
YxrDNZ+BWgIsLKzUvAPACdNC3FvUT16KbtQHYlGXHiZNovJr6PSAJKSzHSTjpfkw9wgud3nZKdb4
zsDyu5KFPgO7Ut918DhGSyos9Fm9SGsSFQ1CS12EAEPXoRpJakMZq7I3pHYQ0MRbbfOWn2K9XZvs
JSYF9c9xTzrNCKJOeoPeR7F0UYVoyNqxWD0IeQVp7WM0n63Au4CrBzXhwkI3fBjQIaPvQQLsYCUv
XKhIDTVgaBYbs+tVJHGx3L62FJMCWNLn4wlyOWXaaeXyKtY55V7PD3k5pIyrT8htoyHMm29Hbn8I
g5qL4gjHjQO/eluLusG2C1r4NVWGV+0WyOndyEGKPFj0TnSob9rxHGDAu28L0pcuFlIdLa+bY7Jh
uNgyquMnEXOM6jKyll52USZVQdCPauFazRcLLO+2QI9wC6GX4d9GCpP8TZrxOOxYiC4vN9dFTgqv
aioG7otR5kjw8a1I02ugHR/tpE8JyfPj+GmkSLfIs1eA26w2ZVpeu5qd49Dk8RRT+jJFIyie66bL
SyJT6XqcbL2cjH1O9lH7DsXKANi6pk3MKn+oBYyfk9Xjf/Svjf5274Gp9Jl7p/7FODXJHbvBS4gK
YO7hMBEBw64q7P0nKtWAo7oedwJDYxEA8fWIORwoWPxeJkAA4aLzr9MUvpO9B/xNx7ip0Vi+JFA+
EhS7VTPcj1hBp/dwIyfbE++5AClAdqQWpAZpsjXWUJgeS0ZNralMtoRu6UFQZrSMeYxNwwZglvA7
rYTe2T5EtUNp/ZwAgcVZafwbhNw0xQ7mFvIIUmqm5pYAn7xLQzFcFMcxePeqJyO5JqpOSokz/VvV
H5JRfTBfBzQ13A+HP4OWO2mroKbYHuwktFkLM5JSrJMWz28boWVBNmkyL04BXcwAOOAiMYw+gT5j
kD0AMYEpMsfgb+/LhyEirSHgagCXUOIjBOSnrgLRXrY8U8AQxinIo7HN3mQFcH+M643MlJJq2R+R
947fy4jJmDQAEv2vy8E+qZkRCD571sb96dAuCkvupKnWgkrtATQvv2Aa8+f0g0jLrjJpr4G3y8d8
H9919orOZDckCGO1wWTchKIJaUyKANt/JGJ2+O6FTc0Fb3eIE7bfjbw7jM7e07wKcZFPZ91Mj7Ur
rHS8Mz+2OIv2WFB1bfncLbZJuGZVKWDG5Xes0WaawQP9tPY6MWtA6xHNRws8+0iYOWLNgpVLoEyP
DBLQLbW+LemEnGWyetpQ+p4ltStpXgiL4lyk1eqk0bH4KDUjFw12okqPUglCUL5sWO8GbJQNDeiR
8oFS+hLyfjmbYego4M06zvwtjXaAFUWTbDeJjwmL0gTghYEnNdUdMC7sJJA0KW0l2hsJoBAv+lfA
UBIZnH43V3c7MC14j20vD0OVgzxeHRoRgDuXfk0aK2wo76enHTZMTs0V/C7Tn/vVnICLLRmyyvCP
GRfYjGMvQiSEJJUHlsmW/wLynbwytVdu/rxuHTJCYFALdeGFDthbsKWz2W7lyYNU13jmXH3iOFku
91KYrSxViN1yJ3c9dsyFL0gm6ArmRw0W/TQbrL+l9KO16W6b79VeZQbCD2hvGToqM8ozF4pHOjRq
a80XX4drNHrmqX2FBu3S0pb7okgZGQYYNdcI68WkoHqapoQsvZJa2eyyhNsSIxAoSzfqdmWX2tdN
fyip8ulMlmkVaPnLNoZDV1SBfm7xVyXgV9nu03wEHdTcQHN7P4/lDMTbFMUui13AJtpV+bec8B1z
Kks/D4LDkzMnWMbWyoqi7vvF76GXCKm3MbsZ/seGMZ7Hz4zEe1snJmBF8/svKdKpV5J0Ho2zdIGi
HxIjfv/6q278yQxa4+bx6UwYLJlKXLbYLYv27yO5vENdv7CtCS5o76dzXpYAvsIUbFvt1VE1LPQy
n1XAFomNrn/7cSgcQ4b5Nos8kUNJyjGoUmFPNCnu8o1vy44z8I9MelH3F70rT6VwSIGdQukDnqQF
p7fD8YIYsgTkBCq8mz7fFSqN7GsouOmev8pC/yjBGbYVg8cOgyutMOg8SLRQHiW7qNTuNwVCDs8D
xKbEzVxbrLocbxmNvdvE7UqZx4pjBC9+mzy0qeS/Kh+9uG0WW3ocFxQ9or7XycQkQ6JozUrE3w60
S7UsxXChu/pLB0rOYJEPhI92W6LmVNGO0haPydgPsBvIFoWppS4Z+zhslYMRu5PUhInZU4OkfiUp
kGM3l8p6eGJ6Ul6hAJwEJ9+4ynCgwLa5xb5kMLhCrPOAS9Bh1BABbeHm+SnB9WAgBCDQi6uzpLMg
fqEBWsqNnAq+uoaAWnZoUFrCM4vM5tnOAKQTU/+SuyVhsXEIPXCFNfKgZwOzRWZRmeJVQa/Zl26p
JFf5XCVT5Xf2mf2FoxbdIzEVeueFQF3lzlHXl8IgAoY+TlQegzj3rsNO6ZHfZASgqyL+P/r4asaJ
Yjs5nFowZ2maLuRdWCzeotY4VA8YgHpk+TlNzlpyKWvyZ1KF8xmoBXKE+zDknqaufltBKNSASfSL
IodHwJ4KlVweUHu+9LgEuxlkBzs78Gn3s4Af0WcPqktj2nGA1W6KdHyitJCeMMwsKsdoEWkexpqy
nHXxSuEdDO6jqu3BrkU3UYj2bylkSciZbW+enquSGC9iP4ZBzxEfYDR1LsQzC91miZeWJKIMqLw8
GN1BqaPbJJucZQlyoNtJIOCIQfrm8plp1OjtEt4jVYIvFAUC+nPqeWgR9EWL+rV6zzr+9NagXjcw
vg8VPfbkI+s6g0iZ7GkZBLhu/mWUVWWImvSRmEsmNyqpLh7a5E8HB2qVjuOwBOFPp1+ZYgjakmKb
lyTRqI9TI40/jMqGWPHce9zV2k7wIDhi/TSjbkuOHkpZXGmrqf/FHhYPSGVBGQSaRvDFWERGugnf
cy9YElaXlCC/W8NrgePbPvKVJEJDWa/kLbLe5KHWnEjHbGmElZ/x/O8q7mwp/ng7Uf34Ia80cfb9
DSOHwUzRBe9pHeqSMfmNBsTHGlBkx3+0U1caOnQakIA70+RxbudhQSBRp0lTkdADcug0wdyjIMup
1X9QKszOrBq0zp3Hj8gBfxGFvq5XImsmaLUYqjIsiLYrfOnWCF5/ffrmUCM49iJRoTYOySvPJYbl
sf9wbvv9g2DZkaHtvmVeMs0yQUYks9qu2cvYXfPxe1z0klQ5oWdcOwRveEEhshJYOBjk6d2lzyaH
OioObULLdwjNYhgpGXtoifkfK313x0fpkHMsKDRqmdS2X72dHZV/XydZL1vjf5Lmh5/bwacZeqLo
uxmqssh6QtMACrp06ourrDx9XiRnFbAHZ6aoMulE+HiTdcjLnF8oGb2DfzH+dPmYo4WndBrMqO3T
MV60gY7g8I71OhslYJKhTugpqvXjdpUjxxAZSBZisBSN08+xjHqY01JHZelFyL8mCGKPH769Y/od
pVUv2i6RhSmxEzGi0E0d+m/wOd8nbVW98pgdvZXk7obKxCuBeLaMQX9wM2l8CbQsBLQjuKd4+226
VWUHTSB4UivsZVcJxRUbbVLgMaIraAnV6IUMrUc+XagDfyj+7bgs6o5sNLYGFMbQcGWEN0RkRjso
P2nJsMlquKDIFUjtmDmZ6UwjYFJFI4xAZsPV2ouhBeBXG2qNJvu3Do0LVWRCPmyy0PJ+W1vVeZ6G
pedT1KLj76gdO4G2ZLnz5smXW6/dyuf+NCltpqWqYxg1KFZe49yJwADw0eVA7HwyFVn7KiHz5ys8
TnoCzXd5Yewrzv1Xf1VWl8M/zhkOWOOfGuU0IyUFnvr0C6DitBGIGHD2VJUFhcwJYYA+h//SrXaw
Ssf66ergQXllhjGUpvHPkzB+qXAtO26Mg2cVanSnhiJrxP3wS4W9Vin9xEcR8YfgYmBTlGyi1AKS
jitTGogWP8Gua1wtVsxhtIl2ZOPx5M2rqCeE0bmlg1x5Uv9lndk3H7Eo6iDmHIi0IcFrAvyW8DKa
yOoXt8tnqZwbCE4NPeZE93Y8HKEdM8FsuJdpEP3NARgARqWmAmTo0pj5B7L+f4N125mPuVO3nyCg
X0AB5E0gR8fph1vFGkFepEgkk5OFRK6LNrVz1+IEFV7p0wgmA3taaI3FWtRwkOor4cS4D8dMtTRZ
OlOakx3ipe2jgTJqsIWITbyS8XiUmdmd9lLbarkrQeKRNEAyFOw10i9trzdBXcuUXt8q3RQeDXhK
rM9qBm2iwM8t/QZSPGJJEOwDP7h11pPF3ANgA/HWC647hldVJe8C6G8GqMoSHHzt1/FoXjEw+LB3
fu37LgNhnw6cIDFnsNXd1PQ0h2KdEx1LqdMmHUCD9xZYOsEeg023eo+sp4cuz9dBxXy1M905sivl
dFtFYNQ6UWmnD2f6lND1n/Ia5vPtBcST9XPHVV/qJIvlzM8p7QqomqlaXZSPBKbUaeww83XJQwTA
gWedanaQgKobXwvRswxYSbXhTr/i5SH6deyicYz0Iq+W7gTzcdI2ZAAMRNIX10OeCIFv2sTuqZ9K
N/flHzYNt1478rSFZ7eKrswSGSWo0QuVRTacfqMvNcvqhrpcOWbIuS/l8q7cpd7z642JGCmbqVL0
dJMyLrgdKqGwxnqR6ffX0IP/EaxH6jIGm40lrHADrYa+ach9k/tJeb8VZ15chx63iMwKzJwtSpQc
hmMyNBgDi2hXQYF7/ACosdj8p7cKN0BuSNtXuP7z9I4uawDRazt7Kx9T5qNJ1NRFEQ73pNiZFUuW
pNszvG6n7bs7tT2SrTH7OheRIAfGun3sPTdqtV4DrVsnDl435a8U9PlGgBXDf9fhR0LBtwgybLZZ
9GqGIaKu/h926cGtT0gmIZpgCnDwAljXkuQuKcY8yBdExKmj4I/B8N3iNhux7cQYaQm75Nuq8YPi
DaNUE3uq8RIb919Zx5WclP9jkRiYbPxpzNkWJ5wODgQ26aFMj9IhU1ZGRdvIB+RlUWywYAJBUT0V
4qtZVJ6ZRM2StteUqlajj6Z0+SxtuETbGggQhpRPlOABwnYwpdu7ZVvn18vJfYcaJC8WVQdFZSLO
EnOylXzYmhsfrNGnZjNOAWKsvdUhGsgPIdiEqxCGs5b8ihdPqRgY1Ljo0bw1bBHcYV3NQYGv3ivO
e6tl/DyaBZCpp0s2ketBWJ8oCRgdo+Y9LDja1Ni5/W7fj6NCtv/R0jhbYDLZDmOLK/yz9++ZwRVE
MVfv9mKRQfVJP3c6XBTE7DOVFzjzSkn9/KLtEFtG5CrSfuLMM/95a0mKaMsCtG7ROGR7Op1QiV+f
i9wH+YuWWRs/dIYcVF+FNnTCtZHlM4J6lVU90Zew/LlYVJoMaqHU47hZxIZhmIRTR7/jozltAJ+g
vNX4kGxlLa/1aU6zynzFFK6Du4kAjwgijsHj/TzKVhjvwrOUnXVGcnAGLdA1baZLrhKhg2UmAQbF
Y8HyvCoqXEgmjjsxcVzQNRS0kqVf9VvZZPg15z1q9ofHRnRVY0bzWAL43o6bSBnGw8nvE90FfGV9
2teogZ5+DsUHt55neiBtp4242BXyXuHlz0CFVnhHBNi9PHAqf2clnjVEl7W7tuuUDx0SkhhQndA0
d17RTTjDybEdHWe8wXXFizgWsmX36F9njBl0TayKXt3Supai9nhpKTSe1kl10nBLZLyb+KoDCrw3
7ClezdJ85OrJnhVKBXbL6Jc4yAIejJtBC1UYqNaSIvjqSaarwrSLVoZyuwyWI3guzDXYIC2zQgNo
kbwYq3HsP9wWmG7lzZSeA2Ma69Xm5z8WNk3FAn7DwLXMJqtLUgakDc5KWFvIvKhxTsNqXnpKZky/
xTJuzoA5of3KO3bwAfRPmGVTp8uNvJXsQoT1YROPpW2vZAeXzlgahPUzs/u9GmTYmInyrcao5e8z
34+9vhyHuO+I+QlYO6uKfBTIZJFKHnBN+81xa4eTfdDoMO+D29B1IVCWRygLC9nE0k9Pb0aQk+MV
qMNeRTMzOvOmITUUBEVkXgxtmYPV4+NNR5ZA+doRqUW/ohRKA4hFnK3jfrNfcn52q2PyAXH09xiP
Nb74Kfgz+DkLh76Xu8CWTxJMB4uYORDzHKgSMrvy4EWUJuisDfSwf42DAfpieWAbe9FKrQSB/Fh7
aVF5N6qoJWjIx7BjR/VWyMGhU2kruamJrLscb3p9pBUCze0zEhgg1x9GtCfC+oCux7oJwBgvqmN7
F0zFUAdLYDfAM/kBR7/bZT4KpiHVjajosqJB3huA/nUMTI+k3Xe26ahNQwhdRf+KxJzohxxBpeHy
MPiPWQ+16M+W/uzduAKnxs6L9bY/YBFJSzAbgKNleSa/fxWRpjzph67AkSV8TrUBu8aeLJ8GT9Z2
fl9/ZlUuRtqGupny72cNbuJXtTgtiWjyu9KIAy5dfcTPvMAfhjAR6fsqQsPHyXtPOf21w7MUQMzW
oK7rsBLdY3rSB0Gm2DDHTlmlMR4hiuxAbvb7hp+k3nDqAAn5/UrkiRYr9Rx0z8IFY3RioVonAP2O
xhj+XPQcCtNvxX4uPFhyxQ7Wa9zFyoN29Ag16sJPLQBHsb2+ujOVQeOk7KkReaGHX9IIXPgifOn+
iCB9nzDW1CXjup03AF98L6G4sp9ODgX7hxfLPKVr5Q5288awfiZ6g+G5g1J37zgcHNJEyzhihL9k
pCjfuRwY+Vp3FX/zz+Au9QC+m9qj5J6OPk3Pt+9qVih4m2C8L6pOKHn7/EoVhK+O0yeImTP+Bazx
hrPoqtLVlcsV0pRF1xzqz88+6j2rmKUXMObTWYD3J8Y35oKsSeHpmHQKmMfF4/0rc7Kdyj2hKtE2
gV8/gQ0QEd4ZhTmXqehBfz1bp6u8SgEug60+v4BO6KoxWr+7RaNcJlRc+02PN54W8gjIKPop/fOk
Q2XWS9bA6Vw7ZfNXTG/a/yre0o7F9N7DjrxBlSsi5EIIyvpRRbWfC8WqmPXMgWzMsAT+6q/Q0vG1
7crcdPPCel5gXc/4TNy7NL66SSrxsvvDrHVzEy5CUWfKpH/OZ2VK8jlwe5qbjy7ctmXkyT408ctS
nhI1C7u/v1L8GnScuqPQ/lYMTbX6AS15uk4MrRmgI7sVgdmjD9MYXV/5+7cb8QERIoP7qch1YEMu
4tNS4BcVYtl/5ngAXDLxZwVqNni05oiOo2TsDnvHiVaRNYcSZSK7UC8RXduAfPPXc6qCDwuw9uMc
nn+BjCZ5wVhzFnxLP5lDgfR96OflNWZOt1zBp1cWxW54O59f/nJ7dNbIiy5qhVJsJ9ISdvo/sVeV
YCl25fb0/gIYkLgBymhUSE8TppXTIJ6BImcoIvKxGcONvXSKLntXdc3PS+sjgS+PEB20y0NWmBHl
XKmTlacrk7nolH76Lcz8WsXvWDhvo7vwQHhHBg/yLZ+Vk07l249DIPAbuoFNuTd4/pF0b8TmE1mK
d6s9HJmnS/4vUgve34ze+yNUWlrsHmIBM+2Ign3I72JES6NMLVBaYkpwsiHs3NjgdBkD/u5gjIep
0VROZv2JHIddcVEND0D0qyKtmZNKJ17/Vh6xbgXKT/bBbGeqNBwpQrsoyzn5lvGAxGX5FR5sRWgh
LgII7AmuiQDKftj10gcH9YUELj3owqahcj7+Li8ymCtiuScWSSqgjHjk7BZTmVCKn/Hwbf8jmfLe
++p+8qiO7XcDxFctfyWt6kjusauefCMdwxoOzjQETLj0LDUn/ePw6ymnfXTQpiYBQl2U4kr1+mq5
rASZN0u58a9QrdB41V6weUs4Fy19uLlkFUyJWbxQS9aP6lYcwllLPthmJ17Ja1lIBGoXul1NPLlM
k10+tiSjmJU6kbh88RoALEDRSB/RG3rXlU77iPavYdyU41OESqWpcgW9b/h3C1MTfMqcP8G7ZeGe
oqUEVhZ+MUjBDkDXlrdpTFgZYTUjWPg8FRhKMuGRD+dMyV9N+QLgJDOMAgXrTQpeUyw5SQrKIYZ4
SQEKVEEo7Yv/+fwP5R9Sw1eNwt1F/7f1xbss803Ma3B0Bt1RGGQyazeEl+46Dn3D3b8GvPxSlqDU
+mxQmUsilauEG5Oa5wjeN02sZJVa2Nqc7BBgRFXEZiCA5CZV1F5EUl6WcPgF0TvzZ13/MhCSYJLY
rmrD89di1qHF+tDajWR8UcKHedDEG6jr9lSvft1OycqXZI+1RhgANQIjMYpp0cvsetKBt6JuWU3q
CqOQWrn2MrbCxiE9KxAWENNTKOaWVNyzTWyunHzG4kbP2S+G6pzoRWGtpz95CdAE2sH7m3MkfptY
m/uNKk5LEbzlV47YU08HBWHP6KLJlW8O47KNoE+Xtj1RSabXeepBnHvyyQGnQjDTfGbd5IM2WOJq
aPLagCD6f6rmbnBSeztBFK/IWpl26BZMifq7iSOtgrpg2hUB89OzfuhntfNtJpfF8QnXSyQ1J7oE
auQ5bvlUTGdGCbfNM6R2/Ohc0RHKX5a0S4gb9wtSSjLCBlcn0YbYPAYSUSAriYkeD5+yD4u6F3ll
bcaIylSpenAGUMiCbjZAXKIxihnO6kJPICXLF5aVsZpVGeE82KkxCWuQYwr/+MSayRGOEaho0cJf
7BkqCl6uq0kVBlC4SXb8lSFGgHYQWAj5gGE/TIPiKmRvXJ+wy6H0D9EUUYWhIA6UyhiuLDjP4g0B
gnX1IbLF9+wAa+/8rWSQkFPyu/M4t6rgmX3+kppAOE8OhwGgK3PKqN2arOzomw4j4M1qK5BVJtxl
ZBSEq32omSgz4qXOXpCGo9/LtxR6zIN+ozld+K5vDFZwlblPHeQGx2T4kV9vhbWR6GCOQqTO9IVa
umIE5Trcmbk5qAUfsHMtI127uc6nBf84oTUuWdlKnRspt/pUsxnVCZd2RFlREOoasF003vPWRn2U
8j/q3/TE6sN4bxTeTfdY5As4Y//GJcGmeIhwEbMe1WyRlxQnDrXCyA9iYcp9dcW8T1WWMFQqZpeO
hQ3uyZGWSh3f0oRByToHpd58nK3cjv0tXoaBXSe+gx4GssEb+1WGBNtsWwZn25jARR8J7DCShXIA
EG8EJzVhpS1BtbrO0K167gbIl28CxbggGR3uvOc1OKU/7lCouhtyWp5R1TxmESZac8NuBaQw1ygR
Ok8rhv3sHqW2AMza/TzdETVOP5LoOFWZkoYNcrAxhYnzUSPIFCyNI435Ac4mt50QtLpogvS6zGiC
F5SAwWbPDMuwjUUgmLte4/PM7SfDeg0j32zRfCo2EptjymxvhcTtyvoDytsjS+WHUXa1YSkdSg5A
XnJi/CGrMZ7vfXomsPBKKzGX1s3NoeFXhlii+SKvh6ZG5hvtX0qslmSr4CxSxrrOwyJH8wxsJk62
ZtHDqlc7XfSvQGADVvMLUNstQJF2yQgYSLWXTrWBVXyu8GdbNHMBNu470J1RXHerVOrkuvGUghQZ
VrFG7YBlRvXb+Eoeumpc2pByeb4sB5HfoL8HoYO2+HozfNM91Y+T3DGBjEDgf4a9fy6iUA1aTK2N
rMXZu6WxjARW+4Y2wEQhoSOMMxARJzTrBnCMAe72U7LzSuNMJr7xVYHhieVXMNT9y5VeckfcB34v
w2Wpz1Zlmf3HBWPgdbVGVJrZqXK664gNGnVFpm65RXawDvvOguyiawm8bxN6iCDRYdvwZy3FbrEZ
8vYpb7ZX2gReXGlqFtyPAIDgSY6NeWtvQK55whb8q1RRj/l5xBkBe95EbBpfCLv1+1PNBP7LVOTX
qFs4QI7s4yFVT51X2I7k2T97D1CqcpRXlEgX/mkrqrLN8+2KR8p9CRFceYOrXtVF/X7/Jldc94tP
anzN0bFJJ0BrClGHf5cCbrNTs4dq8+HIkyfqN1AdeFFwlpGNqxsjVTXkRIOMXvvLVmfbc5toVyKs
xekt9zi7z8kAirM9oWhNOO4o5qCW1oYDWEwbuTb4bnxk1bkqoXwCLzAfblMp/ot3AfUVIssiK+GQ
nCzBtYyKQ+JP5XqQ/YNQkBFJzmjWERmGPSXtTGzRBvLX3Q8/R3mJJihGYg4E1Y0hy+tE879jm9dL
s3ONSIzUdWRnqKcjJi3/foHKPZzxM9QmYJpGmrYXjJb9WXMFAf3MGGdxSh4PBipSZTY7sG3tITJq
8BdtaBjKIiWn++L0O9CU6HSL/8C8XS5TMHh40k7gcXLqxK5Gaoqe+1tGOqmOA9SdONzQOACA722N
teGeFL7nbGvuS3QzWrCf9lacW5X6O6g8YVyVhGk4fCjt786k19RFwfVO2nyo/SHRNnbJm/uaZTt4
1Ooekny5IkZ8ygk7XSQb77sDQDMnv3szTf1wLDrWAymbf2dgVlZNyxaCkcSkR1dl/Fmm9deywU+y
oz+taFq1LAolTLkBQ03kcDiKlF4as730V6A5N5dkIeQwHy9qOFxKY0IlqHB8/PrKxYsjoIap0kyB
+XZs54TyBQhmM3LF/o4VTGJWQgo7ZV3Ah8yWts8fuB6yrYozrUfyyBiAiEGvCPFIENQvPpmKS1tK
/p7woB8nQOlEvZCFx0jbCms3JC/yS+df8GR5jG0a+ylJes1o7V1jQo9aC3t/r3yv0WO0UnFEJhIV
RwNtX5CDzSxKA1bpMtQYvR0+kKvwq0MH6t28LcrEagvkkI1Z0/MmIKJzkv8A8LmAeFgMY/ihBuWJ
JghsqQhlSMp8Y4PNTybwbHmi4KGCOwD+l9mKsdCPmb0g+82Nwoxvkt3dAZRJvVIVyzWC4ahMY//3
oC8OwhEuLGEb/3GyF0DfG/V51I5Ykil+OaG4wWRC6aRfTd7binBM8NNJe3snLaLyIPhg+CVHJLEI
RtvBKx4nqnXKM3Ko3FeaWDIrlUWJ1UrN57IjFifATLtrJtyr0VuTextrCzXPdlyD9653Ocu3bHRx
z7UKqVkPtABIRLOdFWSizjgSbXDjSnRoXIlO2OM99D4vCRYQoRLQ+kn4MjsOq2BoCFqEmmT84C32
r9L2lKkfl1Pt05S2V8xopL0CMWy10usDsbFoJvJIkIuFwlcUwA61zWIcGrQeIcTtXc0rkLCEZ5A7
oaO5trtUCyYhYPGsIpVvLk0mET/7wmLSmBTv/bTxqW7MuyXt99IrTxcBxKDnT/BFp2gM9Uu47L2a
k5BGB/bVAMSOgk18pKhIz3zu2uVjAmLEYb7ZzopXXPHyrniOcqU/MiFXyJbQEpExDJz4+8qRZESL
qxQ09cBKHgdqJ/abf1zRmmQgf33wuSB/IwkLv71OrUmVJk8XPR5Q/L0kyoZxFbmL/8G4upYRuGw7
eHY17lpc81FZWNjs7Q5KIb5527hAy6d7pgrZ9Vt6CV5L+qkLmPsqNHDVDbMJDASC1j9bdzErszV+
3rvK6dtfghX84qpRuX2GGY1KuZ1jJZr8OSpmMjc+y8q1J5GizCVHvJ6egBKgpCVcIwdnPAHkaqh8
xaRVvFTrQ00PjPTk/Yo5X78UrE3HqcusC89ADAQwMS3Sf2M+grFXpvkz28DePyuwu6eeYknMl6xc
kq3dwssc98q/Pot7R6tIw99PC46r+GZJneE2HB+zf005n3onudYqhGARZF/m7qLAkA4BqhCuk3rT
SslPHgqYzDuLYI8Yb1h2te2qgYWVIQl7avZ+0l/POgJqJXy2NyxOzUCsUk0plqgkm0yJsiQ7VigM
1nBp4D3SjehUExVgS1rW44NWeG+E0QtMWbcDnIfh05E3eC3DvEZ3fYJmYW3GN5G+I7LnEyOXJmcf
R38qUVTGz3v2zAF7enXBymaS//+AboGmQObhks3behzaGgpjEBuNjUIZKDD5VCWJnRMWSmS74k8z
usC6sA33MnFPzI5kiprY1qMk6fwHju2c7sHXLkFkOaF7IEYnY5NR3KvaZvmFSIaZjFPB7S+LF9Go
xRV9lEBVpipba9Ze5XUhpTvj2dilfKTjaNOrU++Es8RUWcGpdwSiEQRh9Kabgsl56lVsIpRIMWcr
ldctzHekZxxhi1MAm2EPhsyZY9V9RFpYEWDyJTMt7GJuKVYc7aGjKY4Z+EV91M3ELsQtuH+Jc5q0
D5mtUb1Cztoq0+Fep8w3ZbHHaRIo3I+LfzefqAnm4QjMQmP3BsVwM+zALjoPTl1hDt2NJVOfKKrC
EDtVKXPrVbyEsH5cMNYgSJztg4dn7SyKc/FU10+RIWiSC4qTdvUEXM7kJdtu6w9AODLo3TfftOco
df5+BnsB6imjc+XiKHX3XGOqDWPhMpUkX3JLq+4YQUyYv6P3v838lrsteBXxccPEkFrJxIf2ED0r
x5mavRXDjTHRNbcCDmtPClrtkBMdgUEu5/G47o9WP8Ih7gWZ3iNNh0KNd19T8sK2ECIGhvO23DgE
Z5tPBTLKBHtUgfIVWUz+4S08BbwuHYiwhoyzZ/oI/mSFLVHNsQ8NqASe3Y2Ymf7btrH9fhYzR6N5
mO32ZlI2I5PMr12yC0v7eZTjRuuu3y5pM497N0IozmherfCi/p6tx0HDW6pBYFDJOW+ZrtY7G1FU
7Y64D5Ofv+0yfxm8pBAPcm0ABL68tWk1LFFPh5u3m1aLRzB9pR/TkiglY5Ungq4/JVYGhp0Gre9T
qfcDNh5il/IT9bF+gvBzOI7vuf69IBh9YA2Rw75qS7txc+Xtu/879djBVXyGkNUHkLrjCwm68/Os
BtmBs/GMMj+ocCTw/TzyWwB5k9qm1iQFGYFFiPVAl6N0McYh4BZ+r1hiTW4ywrOBv6V47f8lWQDb
NIc1qWn0PW2oiUmqsgqP2iw1Q09Cx9KI/Bzwz5VazK80a6MqMYrJ5yxkocMERxAiA63/2g3J5QaM
Mb874unGhaYZ0CUUs5GT7xnFNp0pF8aq3/1QPEQHxa4+GAa0hyw8qJvJs4HHIwHZLNSPM6EaYnsB
Yrgs6MrArYmZV8EumOSGd07UxGnLFu2mJWAs0tzbt0KfCxvAEogUqDnxW7LjA2TGroMqQgMWPCf0
s3Bn2zqvgOyRtmKbjxvqj+LX3tT7l1JF7DYyGq9r8v4SLY/xTpa/mDqnbIb2a7k5lAsirll4BSHK
JREKisUSvRjgl9OiQFYnsTW45lrfqqfCHOkjfC0OyrMyixW8XlP0KGeh+fp0K2L5KwpmpvKv8Vl5
4iv5XBrNePTKlM2EI+bWLuyqbW9qQk9kNio3rZQYUs/D+SyVh7TVgVancNOdMbW/GX4fT5RAFM6h
pxTZVwgCIc6pzu7AuefAOFN65ZfLgjD2HJZCI8kl6SWDdQHwqCKVMN83zBz3VjZfx8k6wv/B6So8
bE533ulPZXH80jJcGMDM46fcRdy2djdaZrCZAAyTl/paYE6VwxdyIHsC5O0gBhzc3Y4b6FZD1JL3
hLgUWU/vNa+h5Q/HiTA2JKSIIb6joMirgqEwpKGJ06sH9o8wuYF8XeuBdz/adpjWw/nWb+m8H91W
YxO2smj8e6e+XX6vziLDdIeeMm3ajkhwj1o10CDUbBktVb58bujJcxZDF0CFhncn/NeXyhCvpPHg
b48rXCAffy7Chkkbi+DUyGXpSssbMfRaC0gHznKH+r/sy5dski7RQr92OoyCZyRaXTeCJZ0n+19Z
xoYXQH+mwVG56HPgGhvA1TRcTMA2QwIEHnafzmJP4aDM08HY+a1t8SXg2q6MKVaAI0cQQM1M0HXo
mn05RuFdjMtKAW7VK968/JvbmhGDDLhe4JEcKiI5rI0qb4py/JZ/Wzyt58ngRTi3ZvqjOFx1e6EM
EwyuuRMxzMokM13g18ya+kQ8KJFbrjJklalhwUTAMnM869o6V59lD604JGhNB7FlFprHlqnO76OD
2zfhPT5CQQsq2WhRkjB/1A2pnnVcJvqpcX+nQ/ISTsceV3BlJiIN6248zmTICpmmK8Svp1u9PHGh
yAgAUj51GGTPfwoQxiWcq4fxjvGtchNOXCCoqbM3gc6eTSTZH89/jA0t61ROZGSuuVpfEzCiwVbX
ufeYg9N1EvisA3lRpL71uZ37+V1MAgNSY8cXa5ZjpCqVlIm7BZPy85xc5I6J2HUMssYQs4tmo/AX
uXpcev4lOc85Ncpk0JjLNC0hELWmnJiC12eLhJYf3wQkqZemopVXwVDYTH3tzFDLVi6X5GJKzpCc
f7T7SoBpQkuPyI1LeoUycoq6kcIV1iiVtqTDQNVp8vCS1MNhAPJBOcYmbX6t4Bfc5HIFpu4ew8hU
NbXoyeK/MO5tXIVI2fB/7+ldEHBDVTer/K9Z3pYf2p7kTDv90EXXDqMxPkokxE5T72kjmsETSW62
08dSgE04nBjeS7qSAy4UUtxyvLyXIk3//6cNrJ4AOPNBQvh1WG2MGHLq9MEtWdu/MTq+bA5mnJxt
vu4qhr0GoevS3FWpzvTUvcY58DXj9LeM/CXpjJ+PfKh4r3m/0FlTMwLGr5W8mPqyN3UPO1ToyV/D
m8NIUOysw2B/+sMJoXQieibuF7OgzgOJhsldLGxVcTCBpwTQoe8mY3+CVAp6ooPErDoPIgrV/inP
1FrIv8qcjUBPjM5Weuvt3xBKhtxV3JhMGSR86mnXWfgJgafMKoceOUmtICsFdpR9JWI6b/pwweUR
BORgKp7ajc2m2yTkHnyGCXT1tTho9zskWa80U6TIjb10as70HnxcpogW/F2NWNgA9rRSbidlxvkO
iQPtU7z1QQYkQiMBOREp0mrQGj9xXYv6wSmg8nan5rDk3WAbSUo4H9PxbNV1fIP8afGCiy1aU6yh
9tPTxrfs2wcPPLtxjLs/GMUvIaqreol2ybrPose3L+5mZBHdnzAD+UsK9x8FpYH+wyczwZ2mKYnd
B5v+Aw9Pywj8WWdBc5OEx/u+4aTSZSSNNrsA6rjuQIhcjoNrHVG8wrJnvG3sQNRmbcloVJRDSD3P
jl/vM6A3/oiEO8YfBLNpAcx7uz+aqXI9+X8VO2oGqi5SBIDlWP0QpJ4c2H6aDjnDNUBzv2FQznhA
53dc9s5ecoPFR0TX669LF+CwlhSWk24mKC5P+sjV1TNxDTBz1Xd0coP0YKmOQwN1J9VtBnuAS+AA
c1rhrNW8jvd9MWf7eSH81UtUorpP3Iequ/YHn2ZMSIqNBA0Kyn9BwwP7PxHuXE9pyyy9lvG1Y8Bl
zVazBCqKgaYD0lRXwaR16pxMw6/7paU64MYYoG2g7C1qoVRUuym3QI4nvNkdPYI4mIQ1+uusIm0r
zQpyZ6l5eyW4CTUmumS1wTc1RTNctHkrJ1ERK5b1Ve0tPX/ECegVRoGOfjl1dVAduXgopz1B6Moy
d5HnnZI7J9WB51XeUt1NIGmasMTGt6X7g3HxfHQvmdcdaGUngZX0tYK2yx5nbMKOIora2sIlYkvD
V4WvkW9IwU/qikPYDhJV3ikN0nlMNqseNSmS2Yg/qRU3RdZBZLbltSfw2eQAJDreBU3De3LhjtM8
koo7wxJcJ/jzJbKBLqr4FI0Ma/yazSMPWIMKYnlV+gugG48niTQzQSmxNsgcpWMB3R0UmyYQZSWf
TWC6gOKNzy93l79a95jn3a4p7g4cMKQshnSjO8Ljz05S/MKYghclOGACaajiN4izy52w5v7P2hGf
hxHSOCs0Ygd2Kxtzz69Be+Va807damX7CymaKubWCLRaKIN63q4N8FADKa71mbQBYgpaMGJJd+Pb
0DtVMQPEAnxGU4dSfQS+bJu/g2oFAxe9cJUkSghsgkgLKP1MsZWbKm0t216yqc3/4nfbxAPp81sM
9tWI7kKh1ICFlaRwBcCvQa9e2eAt2ThyMZPDSY4q0cxrN4bAuqlKvF60yycwFLXW/mTp5Frqe4U8
yRkkFrirZSQlGRmLawI5Wz1yc+Ozko/SIE9wzhaoqlanRWCTZSQu3SiDZkvsm+tQqrvXWHrmyCmw
jqcYcGU/9eBXSkIkxN8KNean3SYKkrcCpJCNIRJW8WITRPc7b4WrgUKPZ7CW+QGAVlSsobNEQsAs
nLjW+ijqUyjtZu9dmlVJU55b+9Ju5S7k3IpqqGrqXyBv1XKjaYyDUXZg6DPdq+7UTb6CDj+NuNz5
LNuojxlvAj9JnWbsBzaY4K3gS2zMSHvuCnEED+7ucFI7NBsEGMjp8WXzBAJyPumnAhRDoFdT86qA
rye3L6sHSzvodSV1QZZhYPQsxgPM+y3/bPwkfcJE61yere5IeJKgQhrPgKialnkMmrD+ki6Oa2ni
SBWggqjIXiCk0EKkXjxb10Bbq08rtkVURCKkZo79JqYFr1kWQFBIb4wAaKdf9Dkx+5Fe/W6dzNFc
pGRtXq0pWPb96xes69P/XiYTdOf8L57l5+lebKBtxl6cORjCM8Knv9UUAxWPpWiOA7rezeEEC8f/
naa6EgWmDsnOqlFeXNybUNGvlgkJsyrf3mB45gdGAqrjchpKXQuOUCWAgiuEQPdV6gsY2y9vulOn
TAiYICxWsmxGM0Q2L0GooZj5Qz/oEdbglki0DHp2KKFQ2WZadrvJ7urpLF0VjV1fOII3izsl4jgp
AgNcpwbFji/RM744ql9GCQrDBMXFzzMbrZmaTUFafFtQBL1WMQoTR40SGnZhHoNCyn01kDaPRwr1
2NILkqEe2KLs2ZGOyP5p51ON+qFlmTYolUUQDWnyokypZ1yB8awM/i2p758SXADnaYceliaCe3i7
t1CuwuboDJntI/VPO/xcEuaySO+HgLXJ3IS0tJbtrZgjtZzj4J8kehH8MUMmKKVOSHHxNcOJdbo7
AMOL8epSF6G/ZbxvoIDTFToinAz/LTkYqzNn6veusFBMyoBIgG9IVzgpYcRtw/gN/9nVbRf74jiu
UghhydQxlCYJ+8oI/LCV171FXsaZiooX8/ZfD94Q3Ar5xK+0gJgMaLWXcC7WS+oPduTvqTX5s7IO
96n10VPC+lb5pPheVATOSH4JY0YqNK9HhLS0p/1HaPOSxyH7Zvsioz+HBf9KPhZDZpNay0VS4YWd
lxAlqwXiXrdcmYudLgwUXNLNus2nJt3m7dQP8VWM2CKsyD/Yy+2nhWpwz/Tde35kdAle3aoekaEo
29mJDrVnX6TSLPwHswWiEylDzf7E/CmoOvqKxHAgaNEe/+6WSrSlhFSWXo4MEYK/aYmvfB98DWXh
YdXKggc1yEGMMbry5tHgONezvUx+ygrRFdnMoxmyOFVQUpIDiarlDoOyQT3Cc5JKTwmTq0+lNoSw
lrhBoxU9ZdLJ0MzYaRDzXIbxO6M5BI1M6PH2kB8iiYY7DPYOg1HGcVy4lR8UI45xqasOx5AB8fzZ
864cD0qqOjrBYWQHm55VjNHQvdCt3Dc0tvxZigQrR4tsBpsRtYs1ZS0sSjqmT+tNVZDRx9bMZr+P
tDA+43BC2IOoLstpDKTmhhXRFbJdlPtT+pbrib73nDjAiwkcwvqvCWuBlOSWl3UpMIiJZVY6ByJb
BW5UjJiQAvsTSrsAwDbwMBkVchGxUYWAgtOgbAwNFm4hVozpmBMe/YUiEGdCwiobsLywI2+MFXvo
9IpGZYYrG0D2i1fwjPHHPnUj6gUCWe6uonjyOf5o95VH+uEKQCU/l0DeekAM7MxppAkUbyC/qFZ/
jyd1ggq9enxi36rHL4yK/xSPVaE5cRm3FCat41YBzHlwaBgahGD9cbeD2Dh0rivTqff69DADq8LW
/q0cG/s7U/QF6q2X8i1cGZc9FzLG591kx33kwWkD17FjRG9uiSJzzPuRHlZq1fH1EoZEn1vj9PTY
ZwkWvuXyqMpjl1g97N+LrfBJmNNsOv1EUry4qJZiVc0TLB/3DEyfOG1mpNnRQ8qqn1GGhp7nO1Kp
sYfeta1jxexTjsHOTylfUAbF2RNkEvHyOYBJZhNtPA7RLVu7nMqS0rKJixyJTmUhtwJfdcVF3ij7
fsaKWtItD7BaQmjNvdX21d5eGKjxz4XYG+kBFL0l4xmHyTBXEzZBv93cRS8qobt1nphUGHNyODDo
LPE9Elv11Yr1Ra9TJDUjTj2oOlV9EKVobDPKrwviU9eZrIHvG5TSrkViZuYYWGEMKkt2kKip1ifK
wAYxQPiVPWcgswVIC2e7ayxRs+dsCR12h+Yp9dTwVyUbOZlRpSvP+J4JGbEQTrev0eNnOXVRwLI9
eq+txCLjECt6j3e8QacEutclof9JT7f7jinWjOED40BJ96dGn7pQNsQwC7kHr2hCUpmc8/4QkpOI
2qi06FhC5cXgcJc0EMxp20xnDiihbyhXGJOoyooZWqn2H9Vl8KLQr06toVBjDJK5qisVShaCYa/+
iEVFyG5ofvMNc0oidBSQMqzvrY62CCqvIQ9hAeZuk9FXuyFtwNwkq1XsdkkkpB+ausIGy++0ElHi
jTXji2D6XDvjV06hPpqg6AOkSkLgaReeCTg9N+nucpRxpT0dvlR3o1qskfEDNL9TATpcVIvFjyzy
qjOgQfAge5cHawUNeo45glAcjpj4syNnKfYjWAXEafEJ9NDr6/K3B8dMwJYmMpGcvHwZG2d05FpV
ISuzuq9uz0+m5+xRFzDj+Jf0ZQJlWPOB48W3dRXhGlT7iAWP4NUPAJg3RfkOIo0aXI4/x3rwCCh7
tDBo45lHv9lLG9Rj+4tEP5Y7H85czo81hLeWG+hmAM8T284CgeiVuU5BfT27ARJeIUJGp9Gb8to/
HviJOq9cHmn0BKecXXPdYF9/ytr31kSdHK2bD0VkKtafm2fDh6JsRYLhlAm1jb3WfUvgYssqxFrb
AedA7YSDKPT5ExDqsX86+y7Ct3jDaXdzUbyxRX0A6zAM4bqX+GCUb+a+rFId2VHIFMURbh1U5aV+
IDr3ya76JDwafvEz29mJk/UDwWwp5t56FoWXpiGkcUk91GZDsB8tLAdoWG3fFxK8XccaJvrscCcp
70l4mWHSwL5mPF9OgKLV6DYvOE6K6LnUj0+YSOTe39nU6ZGDAmr3wGNiNH4PQjCRHrjds3saGefA
l7LpJGTEOQM5o0JydgWuC1+oDDYSKxfZdNXbq28LCJZPOLSmNnYxuXsXs3lww8eNW2mWry2NN87P
PnB0uUgiMf5lGKtVsp0gP/UnsYbuubbf1aIUxN4L1N2eH9fxSYaZ9Nb1lSZGYY/L4lM/X26ROGbn
2AAA9wAHpauh928mdv05tELeXWu35PD29NObNx4URJb5TSy20M+K/RFEtGxD7qK/cYS3a2DRt9LT
eyeIwlbLbYelJ236g6DbLTQA4FOjitVuIpHgCm+rURkI/4HcROV8CeaDUhXjvRayZubOjo75QuaU
rEpJag8Uc5obUKKI6r2B6MS72wR/OjvZ2Lz+ZQk3Gv25PQBSqwDNqtzhDu/VSbtp4U1U5lz95xMW
yA/vDmsthIYjpqCB8f0dmOqmABr7uHN8rl/T6sC1SBR+l+M5A21M7wXjCcjVEeCtjCwFekmikv1m
yu2RdwL2oaCNNN5fshajn6KTY9P3+pv0MBk5u1H0JyE+RuqrEZ57pCBDChIFu8Tb8709hdCYFK74
g8qb9sFcJT/qsu4ku67DVm0PT6v1LTl7JK20O5kdEUV4S1yr3NxgAdme/nseIni+7b3+RxNKuNA0
pHoklnoDKuAcC1Azr5+dRMuJnrFLDBUHhmORlcqbSUgg+HZX5FOGcr13/eJm7QmnJG3M9rleGmUZ
F0mRyUJJdizhSy++584DpbKmv8bvbk5Scv4F7/pu5vZKQQW3PBsuJsdwhywIykVnA94rR2iu/ZHv
pnwf5Xptha+oLJjH1ihbqbcWaF4QLuY6v3uIC79+IoFqETfbZh6kRcI62JxyG9tbVO5SGF+6BQwa
eyfxVxarAxamk4Z5goIKc6RYHdkH7StDKGkpCA2g25ECIXvuirW94zCzvlgbKJhVkkKIFEpWTP24
O1HeEtC4kviNAR5t4QO2Sz33N+vwkJIohsngbQcO2SCOuhpQA/RQcZ/jna5HOa2FSnx3qVz96tGt
oriy3X4G/PrPiwO//4MlbmkNGUIC2rtQgY3uWwkD4OYIad24qosrXc78m3jUJ6tCVNZ8QTPT4Mhc
bIurCtdpKutwo19r/THOBPB2jlaotYn2E2bh45FWlNhWHuI99xV8lNAbI4EUgLDR9bOsMHrC8an5
LZnRBNdWDly54vj6M5X+CPppVbvhtGBx+XeXMw6HRSXxTU5Wq4LqdbfhMLiKMbog8GuJQntcZJ3k
7TQIOS4coNu3pyiCtpS4w8N8XQ0WMvbAgCtf1iJLyth2R/poEZavH/+D5IdwQYoe33SnL0ZTXcxN
2mXgxf3kTzZjdOjczw3Ag262UfrL53UUubEOeJ6SUOeQ2f3r6LIEKI7X/h+27DzFWe+/c+5TEuq2
2F2Lm9h/hHtWunMuuJ30kVaDBmg+lFEW4V+n9aIzZ5WBqbtRVS1iH+uKwqJOOYaQ2tawvS0ETHsU
P5DIUjJkrMZUeRMUE/65RlP+ye2zXIp3/2nr6od2cwKUM/7aZpMgtFwtxz5RqCl/MRXPKnLz0TmB
zz/ypiXfKLmQap2og6YayePyO8IktCbKVFsw+xI5igjZdCUT5joUzjaHHkGEysgj7qiyT0mzDsvn
NTK0Txy8ff3sWMhlQPC2LNSLgnh7skwD/UlUipVca7fq03Iqml+nzDDI/UGuehjeGZsvgVszEwVC
wLny/3k49jASqY1fE3Lu8RxZYexiVSgkB7su4+miEtqGQazbDJO51kr+JU/gLLPLNsNUB11BfQxt
tKXb/wnucc7Y3AUX9febb0dd9SkVyM/Zv/WJO2foXZdGsMBjW1IGxg7dMPwIiblQWWgjlDA8Pvkf
RBEp2gRXLmPNiMYHFbFT5AP7wQL0yWlSF1tuCT5k0c/SR020iDnTiKzp+WktEg1UaenSt9bg+PkU
Cq1M0De/d0vvbw1znzlHLxvduhTC/jypYZ2EScrwy05hhr0r2fv/U3QSIrU9TxUKITjmFfBSX+EE
GbNUUaYHyAK+FLjrPPDR64wQVtVMUQKYbxT8RFSw339oqa4Lim2880dcIDGLsxCyiDQJ7egCkN1u
mZbtSYgwoifEWtImfyddHW3zq5/3yTO7MByeYrKeJ1HilK+NISCzhA8zoGZhbelVK0O7OUlTMU4l
yR4iPvtwk5nMj7YKSnOxBCfbbDoKfAmYi9bNBykJWopH/41KDz3U9B9ghMSJg3p2Y2P75ulUJnS4
BCH0LYJTtaiHmBbpq1p3al5TFTvrvozdD4/D5ODSA37QiBdi4D2/iqYTSxS88eskgEMoqyNF59/l
fwfLspVbaAReHamOFduOzebS74SCFgX99p/F7gzH/gpWBYX7yMBJdb9tKTSw2FR2ZbUxckn/5S7Q
D9E/rsBCOU/Dp+iddBjBN71Jb/inMDI1ERpF5iRUF6GCtxLy9OpsbTVQ+Nxdvefqigc6NBl3Zvza
KBaogPWsIRdsJRa/z1xIM5ET56s/U2fFQPJS2B/AjE71Mv+fhjVsa1VSEzXbGXyyvSLbQZ+sXg+n
NjB2itwKkjadSwg4mKT4fZVCW+bqCY3YDaKMnO8+FlIrr6ZVt67NRPwYh0qZxs6dd5/66JUBPSz8
PIdZiAcs+ZEwoy2+gXGlwiXlrX+S/TFKrNDYFcVEFbhJzR7R1MRCQ3fROVVb/HoXvX0rcNYKgchU
0jA+0W+3cPW9hyUove2/85tZn4QWut1Pt39UddjIRNdWLC2HvdEv5ryy1NK8XKpF+1d5VB/kzHv3
vBpmM3A5O69++bbpNcZMBCvycfk8IEqeH8W2kdREXcBkDer7jqXmAgnURi/vY9caE8r82i7eI/Qa
MotsVCwkpuDaemSCt1Dpqjg9ypiM6qJ7sDlS/CyGJRxtnoBzMo69SQM/gGnsz7wJXdSld76W00gH
lFx2Ak80c67l48Ay9iLPzMVybMzZLeSEu7G2aBIrbAJQJ6D32vy7RKfxSh4VFwHTps9Q460pd7O3
fHyzuQ+UNHyx4HCLZ1Fyg/d4syFn+t9Szg5ult/Ywv9RrUyo70oaN9oIUJ9uO5dBVVxfLgwTVV+U
8vVbV1l5GJhRA3NsYpLMXFwkfUSeK62VhyPdX046uskRtec/GcVE9METTZUMfxr7SD/dy4D9m/eT
XU8H+cXLt3Kv/dC/LUat/FDTvIMR/N4X/Y0ZbdPM9jhspgNL+aDMqQLibZq9RwAHCA/6jYrRV35C
lzRYziTNOXg9nwFDenduDuCpX7JYhyGb/iSFAGOnbfET+dR5kGVcQ61PsDrFO0Ynm1yilNK/VaYD
UuoMCfktVDEqBZnRY5Ecg1NeklvYWj8PTwq7bqBKWoLj1rXCrqnxc+Fj7bHhLhLNK4Xa+Lbspb2E
ZRGcTIpXYfIyq+fKSJlaiwA8qconwSLbJUha1vGJgWVrxw7xf9+MdfrPwYhnUj/pI4eEPvJuW54R
v+Ir6j8u2/K553YPOvoeEdlvVO6iMe4PyAijGMX837VxHihHh7n0PR5mhSSuekP7dOQX1DJIRMnq
dhkjzkJ6ufoWN05ot4u3hp9bX9TV74uLWf1ThTfAklX8x2dhgeryejiDJCinAgbF7pVfj9Khw+3x
RMJrw68tZ7JguoK6xzIKA0USTGQDfV+UML5egWVYyP3/rpRe9q+e/NWalyUsOPofET+cTjqsFyCZ
r4Keu3EQpJHI+nqNpWvsc7xit0xFTTYONcgL5t3bpWfv+n5Ajj7HyDx+7BicKFkxuW2Hg6IwMjO6
oGi86IyDu45XHmllB/EsSlhBofV8U6OEVmay5DdhCGL4Hlb/S0+/u/dNKmuJNg6q0ve88f5toNDj
ssTu/QCApBJJHSUdVZRDnaBFuuisMI2jG1UjOqGojw/pKdMgvtkMyeu2GvRml+Z0s1lg7uat4Vtv
s90rHfShnvIfi0JbOzW6G4uSoq/p5YRC8Ms8zWSTPiFTqyYReQ1Q7LIjJlqV56l8k4ghgl21ceFL
4t2vsUkgWSi/2xgcmaD7eyDSAqeqsSmoNSdcVq7cpil6Kk6bri9sJg1EIRZukggk+vhf/qyUHqWh
yO44Kmg2sz03Z2eA8rkfrp9tsZTgeZKOqUzElWt+yPVf4bR1hfW9ng3VAluTXqiWugr/iw/Xtqp+
Ya+F+xw3wxvqd4P4Um+Sz9b150AFJTmvHwXUUCi/4uKlh2dE/hiLp5RCx0vNjYve8TlGx4OdaOw7
f2/E+tLp/Vary3A41Wvif4ju6f7p9HJBs6nF1bRPESl+I0n1EaKSk3Y7DXQFR0/T6gZZJY3GSlH4
nH6I4vkMB8OrENRR2arYxx6I/aOOVcy6R/MSlRssydSEPkTcN8H7hU8YJBNzlkyLD/C863qp5h0k
TC9VdjcXlPYDMXWxW6020ULxWOUVwcH0CXNB8l0CqsYKr4fOhZsCmsIgdz8jiC69cG59RMPic0RC
8KlU5Ct+hESZEysXMr8DuDpDTwsDDvm6qPXYHddx6n+l8AamH6Hfp3MVwZUHEYuXDL4I59h7Tkc3
O/68mjLZyeBqqUIev2OjQdkMqQl4gdCKaQ4crIs1XxJxcGj6zKJmN0zc+M1KmlMSMkfFPRW5S0+L
uV7batWBKcao5aqznpYdR1l81dk894SMnt3RGAOZCAG6d/Dp2NocNYaGSkelf8c9f6hd46TL7lQc
jd0eBLqF1JNaVqvM1iQF/PRQBW6tQH5EN8ovwqvzcK7f+MPlVNQIcNr/h83XhcgveQRZqthAExWg
kuGI7RAgznOceh1vXUhhlE32tjqakRuJjMM22smDQJP5pStK3ekh83YljxYaw7n/cOvAgwjSJC7/
rSp0Rjm70cndiku2JoopuodaWeOaa21kHctf+uh9Tnx6gu7fPX5hveNyztMlLafQIHm/jnbd8N4J
9nXC30ynMib1EjYGs29yDXovB4rLlCzw/V0L2l5q4nAEPxIkPMjpvHWRxAbyl2YRzqbUqgdcfoOa
lysNyDUfr3824bjtHqdVjhFKJ7w6DEPNxU02P7DqvB/V8ND7N59NRQdj9ODHL1EnIwk8zx35cxWj
0FsmcKG3DpMoUNFFyKOlQ+ZE32tQ2E6nxr4CwVFeDbrbDP0D1V4ddHd2jmKxPBswBz6+5bcysQqR
Mv8gLmUAarKyquayskFFviE0Dh7h5NuPlBvfBK3EBtjQ0Ids3prDrLc/bOQoPngITcytkaxD6e3T
CE+w7JcKqPZxwrf6aoA03mU5KvUtQxCH1KJ5qFW31L91QaDbSZJm/xpR5ZAjZ6haEUKfYli1V7qG
S7CYkHAm5JRlye0OJ+Waiy5inh0yT88ERAoj71ha5DOeb2ZCNr/NEmSoho+Gxhqi3U3a6/d/991k
THk7EwXONRHauNkxuWgNDeve6qa4R27pDW/DTBLnnumMM57rbtiyASs45wC4V9RKNLB6z/xXWNGb
OscEaRjGMdfhg+JTCAJBdaHt+9XI2dI5M0qjXGr6/ilkz5nGD5ygdqa3UJpn74rF7mu0az9JhoJz
StGXNLK2gwglcnZulpdId7WhpFuYuXXvcqAQ5z8jd73hpxR8BpZw/DUJPPMmTcueoql9K86CzZrd
wpwslfjYIBErrXuyRO+R6b60jVIekYe7aZHihLZNZhzyBmli6MS56PBHioNfBG7CxuckJXHNGG1D
cagRcMGZ2bwCrcUracUm1bVzEIkVI/IsTt0KxNhRUIYPl3XtrXjgy7QGwibLhnl7GG8Gqd3X+4jp
CRApha7MZqEwk7086M0LqFNVrAGcfntJloRaQNkk+ZnxnoAMSI9XOHkW36F3KHY4AxAy9Vca/tPv
N1XQTgdpswWEqhawvymISLXuzUEfkPql94q2niN0HZx+KQsv79xcjV6+dM1LnalayGob3PbRxime
sXAwG6sXj/l1SjjVJyRTforVX+Awr42yV/6KWb/ohBypa4b9KBPkELqjuM6YjuxW7LolGNMHZ1wU
p7PE9pPk8sSGBRm6aLJsuBt64Cs8loFvB94Sdzn089HRDSFhT0q8XFdoZEED/VNkdFTCbUv8/kyG
cchMoi0aJtvR9MRtoC06LQ15NtJjr8KmoeB3xWbzNmyx+Bl5CkYH/8X/gfE5g4Ne3nNl4Ppaq73S
0B+WJEtQqP6J7H34l27IP0fJofknBKRgl4s1u5CwQQ5f9biswdQkjY3VFVttTGUIzMVGtzbMNCNa
1x0QsMD/rSujkeQWUkEpxSGKQ+DRIC5oTbawJ/kVvspj8rysjk3ZZWZoJChz2XBWxsaYQl5P52cN
3JPMw2Vxz+CgG6Cr3u7HXMX8YC5cs8ctPmBVzlJemYimxkgykAf+XNeO1DG6G24TcP5rXyk5lAfS
z1KACmAyaDaxGJ9V767c5trqTBQLQ+vLRNXeTd4OO321TLQwhaavBQL2o38NMltLF/gUWOXU/KuO
HKFoYvhjiH5tgKAeHa6h0x4VQMPq/12lJL8Ou2fiHYqEWGexZ+HZFZq6gzbCwEVLrj2p1xOe876N
X7Ngk2B0KYMQNYza/0cvHddQ7Sgwz9FKf1S19IC8J1wB8iuqHz2sCe2KGzgHLEPe0xifjF3dmMB/
WMtDK2r+TVMa3jZPLm/vPuNUbCfIhVB3iXiGjfxKwEattKXPmJp6klpvvkOcUn90hCSGxfT4QoIj
EQIm4brzlAthuYgIy0enY3omSDJLo3gEn9R9LryjMoUC8Z7M+98zCQoaMATxCv/UGg5OpLh6UZms
BxTc7839P11puVTyWN5qNvUrL0nIIdw/ldGBA94TiT1NNngjHkkNEAbpc4eBM5yyfloTnCZpjFWl
zXf7q7toEZRlH250RmOvCev3uN1l3MlC4l6EH9XhY2tUkMTF+mIgN4L9f1EsDua0ASzj7RE7F2qc
hG4LfB5n7bywyoVUDH/xLqdaR+6+kezXe/4Fnnx4OGmMxHQNeLE3K/D5pw1WA+rmOp7xYtYrFyM2
dbSgSTtcBktfcSev/VXbqe7eeQ3F3yYXqVj8GK81GzLV++L4WFQYYnvgxnKrdAZXqbh/5AQ9y0Uw
myDu1v+6YppGXi/Oo7chXDf4/ssRxxtlcBEkige24CDahiqVeWs17L/4+zJorF+Bxlisj3d3Yc5m
H4LKhUfRC8poPvdDM6ibgwPuXcvFg+w+c9sfZenvItp4NT92sE/iA3dyfK+3zOpvgTBjnT1fiZ5D
TEEycElkZz+z2EkullVyY5q2O+CZpjndV/ByxzUXOqc05UWMHFNOvhpAheusEfPCMGm4VI8piG58
HAPgU2UtGIWoOLh2siWX1uU+q4eHeTRcDkobwxuk5Xz6bKlZ65fNard7YUiRdQGwvCHE/WYSdjsI
ZSPlneTxOpLArSeM81oZHWuzN4Ocf7K0XPagoqUkAY1V2lCxJkOUagwsSrmi9fSizJBKH77uewF7
Y6D7RvlzmeFxQASwpqP6135r58mPYp0ipqtYo4Q/9SyWv8eVfza7bgnBgL6sXCgaQTHgA8BFG8tq
JbvgGV44xcb4hOXhdNDXWWR+7xyOLs6PF6P2T7z9SUrFr2kas0o2sPfuBL8iLMKacY7qJyS/Be3H
VsWaocWG3F1Am9NANDCBB7nCxnCVvPP9q16SyDdjEDZ6qia9/S4K0UOr3CO+jSYMVAWjLMIdGDJQ
bQv0k113cAUXfB0KAyZ3r7KE4ITQO6RV6tnzVCDNmJ32RaOyXn5rk0gYydWXgv5PH7L7/rbioqQy
bDAXb6cb+goGYWSxTowsqeT74doiBhb8yz+npYqm/8kMaWkcFPuOH1GoR+DETy8eWpLHoL/llquL
+/ARxvPMWAQAL6qHJ2yLB376vZMRM/BXNPvq358rk0QbC6qNPc+ELG+OvOYjAC5/Le0AA4sbTZKy
egda/wx3j3oAJ+QYl+dwSXh0qCT95kEsPbQx3PFIT1G3hmHpjypSGTSigeEO9bBQtLc0aaC0bZtW
K2RHm/AivfVXDeJ1YLxPFLjAEA81fbjfrHRs3c5vFiQZD0D2diiVHhpEjjNe8WFWxDat3bdGcWPs
T+ldynKuMRT6UArcFx+3lf4udi0DClvKTGjQyP97Y5E6vuM+fkjv8IVyAAtZxqR9JeTSvLCZ8xWE
MxG04bNmOtElTzOpi8OAzjSwRy1xRdff3OVZpyp4qnmEiJWrnTNSKnAq4Er5OigvnWzfb85sgT/b
CRCpVoUIkIOKTS5G2WZqplPkgqtZvuUTOpkj1Eh1Y6VczZRLGVXbGbNT5AbOH5IpkWMeefMixYVq
DaKRwQGy5X4TEFKO6qa0QkPmUNF/mHnNxJMcir9W3XmBGYJSminQcBBmfdm9wGNuYEDCot69nvQS
htNkpFvmojj9xRSmaMJKf1ieB4G0uoUmAtbvuH+yzGNqp3CqK7p1h9DppAOmZbv682tzL42zm7UB
70DPiTcicxN2psyCFrWUZoc612aYgmvab+tOce3isdkDPG97PoskCPke3lYYoDERfYdX9zeZnQQc
rsJ202d/y/kdkwU19UYp8GEAKjqtZ1qEcHjeoKdJ8JzuLCEsrAZ98f85dPoeBRvYYA6p2fNmH1q4
H7lEY8Fyk+AskP8Rd7w4d1uO5ugapalG55uVEAMh5Md20MIFC1lnuxXB4IqKEC1unvJFyg0G3oCn
FDhdku1zWldClfwm+Q0UUinnxm8ioHqHR1vUse9kgrpDF9qvbwUjx+pSbiaPkleMP1fuRhi9hofi
ErH22+SAQCGRZzKOyvrPj4gWEQccNx9cYDs/vyaEz+xX7gAra7moO1PaXxdx0yN7GdVvpTt8J2Ne
1x680lyv1fLhio/HgzMBW/1JF6u4HnHAmj5/FhGDXPPQg0RJu22QhVS6KVUUTR03anySDM+Y6Cd4
coYgqcC/wrGesHoNzv8tGRgackexlhBaPVBkiz6pTGOkamaWR/TMQTm53ZORVljs0YnLRBptm2+O
V1KsS/XaxeDwXiW/rDlog5TcUR3x0gTNc+BiMJaMNEmP4Wdm0ku/KTFq+GB0Dk6sh48eJhvnp9XP
CmU6/F68qf2P+Celxrf+WlSbbf3IOn7cpB3D92HK8SX/uqSqr7C44wFDtlm/FIT06GrURfKXXYia
GfOO/rqf3yE0/dGFJHCCgybZPAiWCpVnDOiOaPlodanQKguQg63vTPHEWrVDKfjYSnolE/fTTat2
qn3bTlVaT1T0DFHKVGFl/mOjeoO8Owf5NOT8QT7mxuMF6/lgqzOS4ka8zBEsDcvJCHZggYGUPTSu
86I29d7tWjn6LYqqE5PUVAbcQlRRKywY5WRJKlpmwCOtJzMm52Js3nd3POuDsBxUHLz8sYGR31RG
yE7Uheq1ryIx6V7JUTbeqWdnXiF2GqSZzyn5C4wqep1g91bDljl7Cw6Hxidk0aWfahej7UPnfEWk
KMHicfbdYSmYgX5FV2Waik9d+4lwlTeBqQHFShooIZcXS/OTitRj+mkF5Vud24YRUaM96VZmIr8M
+Si8DeO25jeZ+UNtP0gNtXMJCmiGZb8Smg/L90ow2rhlfEKfixcur15/y6gAzWwdVnJqVM41zxln
7f9vVwHuot/3nQSN7hbvtmjI6mFUXQQ8YZe4O8INJaRV+Zzha0/O19qt9ZYjgrw1jqCxT/PvD1qx
pU6NF/KRnlSElrg2ej5L+wWjpTuiZLXQiUmlZy8CuCABC3Oxi8GiO3TJHWHDnW/qTWR0XbMLfQ0m
DuRvzbHVmFX/q2v9U9Re0LZJTi9kLDe6JlkZ1coUsgGWW4aI9xZjOHR4xCrdwseMonQJaUiiFQt2
f8GPdaT+MWUFNqvt+2Nj/75kDjtjZfRNM/x7JtsMR1+mZtUXcK+MYN6I4L6F/LFeUieUrCl8ovjJ
/hnVANcRoNwERP7Yz67b5TCoWm6zBbgU3GcJ22d/LFzIzGJ7i8xTX2TEpg2Pu2JuHJCxbb8yEeZX
SspbvWFDGGH7uvqiwTxuRQ+aOMV8mDMEe5C0H+xqc3J3XKgoac+PzH4IeyJNAJEO0uypcnvGb+il
q9yai3wHm1lWku9Dy+WrVXG13eo6mXla9izYQslvU0tgAsSe9XJ/4b1tC9dUJk4RfwxZ5HBIiNob
3X5iFffF24NiWjhCiDRYf2jw62fcTwd7kWk0RuV2eAInFaHJKlafskcDANT6wjtoTGMB06ej9uqQ
g8KTpDZIyRLP7CNHi3rKief6AIt0tFNQf590pMxDaB1UU7pbmXHqEA2IWvaAyW1XFNWaeX+ubdpE
Nj3/cMl9KHbJQPuaRfc+Avd4Ku4uswctx0Bk//qJC+SCCJ6poOjySoP62dKftOe5P1wK+u9zZrcB
9rAQIOKVkz7l/0m5IlG5F+6mR/Gs6GKGLkj2SM80nvqcoIa5DQhafcVPmpEotUrnG3vRWbsVrMW1
/LyJFTvFTuqmq+KEqxcDLN81RYgfV4D4O6wuUn/hejqp9mVk20aCGtLe5UYu2JMVCYs7YSkIdwzJ
rVn3Mkd02ib6OwayHwsobkhkMaQ4vAFIUOtzmu8FNjcCTaBrZpCFZWgoZVchK00iLmC+CF+IHdda
uVDltGnqggzGiMfj8f5ynSfhzJ5rnN9IFKH8GyQ8PchGfWuUjtgmAtqjS3D4sqYnUaUfF1LI7RHe
ek+JPL2vC3AQ+3+0DJqIEo0feBBc0j0CT7LIrRoPwyzcqULFcH1d+VwC2xFfOoN5dSAGIt8M4/3v
7HvF69qyTvDudcqELKOC9POYu3eu91zZ//1AAS8Uo0N3VYuVlTwK7zU1lWNLgAqA7N6pa1ulTZaj
ltplfeRGW7MJQoIhDxNSCbqRhtDFWioZoOyvhUfFUvp8C+1L7sjKLSypRMESiCXgD9MC+s7rgbBc
cm0DO54846bkCBPQnAlRXSUwrXw/12z3YjK71wedjD+GX191DyGaVeULL63JuBqL2MFTQuMi2qQb
pcfWjLPBkoPOXYwnlPuqazJaFUHS3vgTOAO1wGWmhdqEaMUhub0vJklMix9l+51vPxl8jJE1dVsv
FL54u7AhYcUO3N+r35sU3KDSdM5P62XG0C+LjkwFkPAeMFHTR6Wo8xI66UOZy/telmxXmPUZN57q
Z/2aUVUL0Mmbr7tzI/Z0hHyF3TiMH0g2Ac3s6fw0Q6BCp/VmA/T7im1DKa3Hvi2A5X8wnEQ0v1/P
FW+lAHaVoIEah1dMfx1UOikcysr+GNncCWXkDgy+IhiB0sKLxu9gqxuwOLsLXPCYyMAym6UnxSq9
7uqSx+ACC4pPT306vmV4kBU9xvPxaoHZCRHC3Dw93NkajVv7MIx+P8IywvSjekRyQmkNG8OTFtUg
ndFYVwP6/zfgInoLPuSVzI0QV5EM/4pVknNCQGmuRZjAbxpMg7AenFA11bposDcXcGnHIHuOG/sy
pYZlXdrrZPsi1wgEazCIahdEO7p2lRQJOJ1ON8mS4+oUKpFlecqohCza1sMedvgAKJf7e/07c26e
bt8gdIwurEMGnVhuSQsONpKs1hJZ46vC47bPQdRBHCzEHMlHE4pPS67S1jhkLsnAfEOIy7zKEvIx
W7mYM8K2d6HAhcx0KxD82jKidowVs4QNRtffYFEf0FqTY6NfZorqPX39ZzufjPQRIhQNwzmeoLww
WY5Elw6BVKCsm3l8U0V/MTeVrVk28+IO1xDGW0Kh73Bz7w0NFo+2cAPG7vV1535y1rYK45/ra0/A
glTy+QAczudMAHTzw4xoQldYIoSb76iJhJHGtDqP0OdQYH3lM9EF5zUjPp2IMokeDorqnzgKV8bT
8wMWMEpSRkdrZ27IdazAGtIEncrTK4//Qrq8WXeU8Iun4MHsT62Uu9h03KBuCPviI3bpfMr9j0oa
1aXWcdRRwgt2je8gv87W8OiOPhIcCh1D25ydU7APjrn4FwZgEHjdUGgEut4vwR4mxL8TUG1SvW9E
xDXgfDFtqiGHYRwt0z9F0+kc5FZ5wwZ3DkkEM9CSGOkMZxLPWwOqIMPLdxpI7T7orvtptHWEOqEK
BHUWS3jtc3WfkGgiRE/C49rdSCh6BW4tVBEQ3DBXzi2rJswe1vF9aZtcoI9kKwCc3KKDAB59ODX3
9YS/LRIlRQLiSWmBPZwHcJJzjWub6fgZdunqFjlQ+096/Cl+m/ImtwAnqLyo1rXieJpgSbmBeFl9
ON0v6msoEOskaeT/Rz872vLIPt2DI6FGTrLr3rF2jir+hRrFctFwE3oHUPozDb4bX4vjBcT9km4a
wpTqpZfkzMSuckOl/ZCcjnomvFyWaSeT7erMdchGtmgG8HXFMfj5A71cTForhRJa/sKiUJe6IkV1
a4Qn+94IMk110QEg5dFeJJ2CgtPgFM4KbdEhlKO4anWmbXreDN80Wh6sZetyq49YYogRSpq6Sn8r
yLKFxdw4REL72/O7mX8f1LuaNHZpUskfZcg68lctd/8nt/irjeaLaa1Hevb79YV8IXwRynLGefTP
H6GrkTjKoDUuY7iXLLVAaownDipnaUhLxRkBc6HqsZtLPRDGouTo5FLZn6af5rWJaDTMM8AeMG7v
IRR4DkPBNTa5YaxqIj6JGSRLHyShCtdj2E7iyj1Lj7h7B1//tq7KM5RXmss3IXMIOD5H0TBvEmQx
9icIl1Ejy1Opr/aV/GTxvEI79Vtuzp2/EQgrHFXaMrf106bEQf24lcKQukowSHpySd2tCZ4nfs7o
K8nyGoqftjSlbLYKufL7fipRpVhwrxwN4phh7bJHqWto5iDwTU3e2rhnxYVEdL/InLzfz4Gaa2Sv
XVrHBMgzWMAh3MMRJHYmlhkPyP49YaoSq5JzpI9gqu3ndSEUaxTmns1TsRvGpwjhoaT/t83alHLA
LPvGFOL3DToWXbRm5m9pxQGVMP616uXHQYCB6wpYYnjy7OU2aW7xGYD3eoMpsGTMNuweY/RWWHtT
ssbgx2B3Tkiv1+PIyFnWzamPUDiptuhdpGbZnat/OGuQcsCQifVjNM/jhSSaQPRYg8cBKuAmi15H
wt4sTYYzTTK03JRj8F0nUaGnE99tV+d97a/mvyyY2wvbyL+bfEDtzrYb6XFlpRt+Ig0mXxzRqmTr
SerC2dYATzFXCtmUyUMbNClFqXA943HjMA+0TCuPNoVcuJbB/3oePav1QbNtdqbbTSq40DGzjiRE
hwrYlk7lHZq2Tq1KpOhfsa0W7Nd2mMeC3Ubjb3l/nbZyBVSpxSoxMj68N5J8jqdSrFBkugokievT
IC+QPcv0KT6BWKMop0WtcF5UsEMjqwypBLt5DDPSniSl1nFP+IDU+CFsrOOT+TZSTrxy2/xf/8Gq
6+baxw8tQz3pgiXpFlvK9Afa4mC6lk3WCPgVXIZe6IT4llNjdTOiTv75V5jzodD1nJcFCl5dTz2k
jptLwlQzz5Kc8WADQ88lZjstDabocWbd+cPT6Js9Q7P0woE4DEN7COWUt6c+p5T03wyHT1/45gZs
2viZXxnBEb48Qfko6bHBHP/Z05E20IQrHdad1GYN375ydhpuN7uqBiC4lIkrxNqYcrv2/U0pTuW+
URvB1geHyTXXUEwzZAkB4yA82LkUagiyMoV/ls0GvnjpAXEpdm3QdBLBJNzeKp1DBO18aRqNm19S
uIWjb7A4WzbS/5bMOziCjljmDU9QfHUB0RDehH7bAo0gVas7olf8HvVZX5MedXRGLuEB8alLG9V2
u9D51cmjI8z9y04yKnG+iTIHnwJ/FswtHt64yVLHMhl4RXRAyVaUoSPDe2BPRgm2rYznWIw3bf5T
7rw6wuaoHc/aic6jyQiqjnIJAn4z6/WYekHIf1Tq2Pyg8xs+YsR6eo/YeAWn43vAChkr4vaaJdcO
ko8uS+1LcuIz21nvoNfvzQ83B2Ut7Oa3pq0WnfdPeuwrPMrp/LH+rRdSfF7ucpYlZTOzumBB78IU
OuuSVNLcT2arS7LrW4Rb9h4xmT601ARKrGfwKHMvwBX5E9rEsCpmf51t2DtiuiB5LckF6WpnUFqV
DW67T+ivZjP2C63afu+KyMYa7oZMzRS6WQxPzSsLFk/mJMsBOagjacWdeJqyIrOCDJ2Vkh+nfoIF
mtJ1qE1OrP0Ha4xSxuVj8U7LKr5QlgeO25/GFXyrm66+giM3yZuUsqNYpfWShrSkuLjvSFkapyD7
Zl23YaB2IS3Sk7x+jAwsjMC2XYuCju+pdVB1OZppYOMEQDNYxAazBML5gJ3KvyssbQ9BvGGAg4kZ
Y0BwYPMOwIFwS9+VJtZkgtXiM7UffUU80RlTm19pFOC3aEqZsCW3AT5O9Vvcaxm1OHpUKOwT8abl
gP6yJYjyUW2lSSd7VGxQWbEwJkGY+trP2HszsdHHhBTUyn5sJg+6SxcHXBfn+eRofyNQvHF6WIAJ
zKTZwBn+Q6bnl4uXh4FA3Upsh5vtuM6W8b4JGWviLTTwx3PDm5mXMP7ZE23qgTg5PFPM6qvarIhp
GviF4P56rwcwzuVi/98AKcGBBzV4pxzImvXSLTSAWFph6T7A+wF3CiZQsTIBpmwlV7PDas6gkM0K
o+elUrmQPo3WwTpAplbXHESZtCsGbdG/RKtlsLf/OkOfltg8LYv2XVlvvc9Z08/zpgx8jPcNas1U
71e7HB4CdoR5kdomt3Y2DToQEiLWtvVtkI1cjEAGJ31hR/h7wvrbqheeMxsFuG5bjQfela0PHSYm
RxNcL6wzlwdT1ZMPdCyGn9jGth2pdTSL6gvRSx/gItyrghO1kE01yLB1GtUoIkdOUCLKmvdOptcV
TkH4A+NFzxIpbb0Ae09B6nom+7Z35/8VJnSTCU7CaABZOZ6MyQC3cyDMh12p+7+m8z92KwTGic5e
qGe0WzxEiXA2FPUktBY0+yxsA4lKaBUqZobG9YM6PvJhlFyWX7MgAuvItRwIV8mFBNkKKeFnBHNM
Ycv5VwJSTS/grVDv6nfun5qJEhaPmAhKe491FFaF6tlsC3/W5LdfYKZOiT19ong6mio/iDsLZHkm
oSgOH9cxerGK1/gPTsCKRR8qNg9kl4KfuqL57ZX1IB0vfm+rVphCgfLxywaTaZHwBfuLaOBCtKjj
KfUMy/GXENKE2YDzELhL+QQq1vKqW2Cezk7rh0zEMc3hUOa9nX34MZt/E+hraXNkJ5rn8VMMVncb
272SBSu7gJANZUS2J1YUmLrOzb74fnZ/r1xJdwBGuhBnHbkbSNwxdRlRnnZFFZpwKdT9Ir9UwlKi
K0TIYfdaPQEZJMDm95S3JbzIOHtHOFuwuZ9gMDR+qZYPM2muOpoDzGfXac6u49ZF+eqoOzz780sy
hdWO66hlFXHcqNKPsElabUIVFEQPcovR2s3bfhDP4P+pLQy/snjfK0NoErbHfpyayvM6yy+IJ8B/
7JvQQKIyyIRMEJZ01mVP9h3aRjRwX9IpEF/VabCunmMLgmZLsHNbx7kQBzbj/EobtcsCs5CJ2kbx
eVEtuIvGjhauf+1Fnx6c8cNZL6E+UsW4uJDVLKSIUnBM2gLRdO2eUy6b8eR4tdVB+DNV1xpHV34P
bmCb0Vkww9kTMD1wjcfcJoheIpJkIsdeqAWu7/oZwi7eVN1Z8gfquRefBjG3GKL+uN5+aa7do6R+
z6Lw7fX2oU8HOKNbXoCisG/BfHK+tqTO7uYAuLp+VCdTtOeCXXxF3nDTF1ylwyBrStbkTJ1ipWZx
t5YZzpdWywy1Jzhdzw56ti/14MOWE7wFyNKvGjd6/iBChRBLYOonhaexeSl2MraZL4dvdl7Dv6/H
LIOYAV/NNqp4GJkT882y/pJU5ayMETds+AUlWb0Jl4PBXARLTJiMkMNdzbfoVvZcGlr59Xka0yoR
bKZhvg6JA81c+j4agr3aof0hUjbu9ep3wfXuduRJpfP97JfTTdpO7DXwBPDVkK7q6+mkaxqEINHH
5o7NaHi1eZ6Doy2oD6cT0KFxyqfA1TyiTr03CCavKDxpYyO9dsfra23A71lhuMNJsoOxviF5+QDS
cJSu3URkmtXIxtR/rnNknsanGAiFEigliKfbSlmtVUU6C9PFNPwCJ9AFqgTUEgTMauD96AYcy830
sEHJn6hLittWRIt5aEo2zcgj+OURg4MLmIYQcmoI6Mt8v0vyI0sXgAUFONX/EmojX2O0PyWsbo7/
OUF+NM31qoQymE0mSh6FNMxvpxkRYV0Ei3IYpLOXjPvyeJVL0Xh1EnonsBxjGQDxhJiBzal1KEPk
fH/uMuNDqlfPBTfEVMpqlp58vz0SWNflCpSONhicxAM6aRnn5W14oTBq64PvppKBE//9iYUKXl+w
2sIa3krVpXkFLEwZyWLBeetjGfzvP4RkJwMhuNt6meHONEtM/BgpFmlCWQWejPvPzeJ6wb2bWRPA
2kiKKNeRQx+97HQc+eNu001jM0hFR4/ce0ZqUtqi2QHntzg7rLElggkSSO3mMF7LhbSZy9GZBI08
UNOo6QcvCwiqCzm4s4RiN7bQRinKxpKPKkzP897MtLP/lnK9+EN57SzNyf0/Gs7H36SkODSx3XBu
8wsUZ9hHMoI5vc/2TJHKuiEwtfF2sjspqOXbfj1AdzdmtSDQ88XXljbuTgoK5GmXP3rFqiUpNG6o
38rkwGFTVNpzOiX/Rm1XrGRNtrsaVXmxpnk816UmhHDREWzouybCw1fzwLxIboyyyBa5QVpMtuo2
Ir8qb1nygFaUANkwH/s5BIB1u3FZXGOHDUONnvyeMTa794n9UDUEqtfSDTbkrM8bqccmYf8fds8h
W6M5wnOVVQIOGkX0D8bbn6vg4L38PT1Eaczd1tTSm0OmqYwArnLwl/0PUsL8CqSoS7LlXsQb1RZd
C9zH8mvvatQ8cdL6gyq80HpBORGvUpjU6+vBUG08gk6ZMY4pybaNhtU/wsKWhz+N9J0sqIBBQg5N
TH37xpXr5W5bAvWhGv/nUUn1RmOIKzgj1JaiPvqfEHc7Mp0SLm1XxOKRAenjP/wmybm4IcViiHxa
mqKGgxAbsxIY3JJP9+LJ/1mkn6Vd+4l9Y/C5GwXxTfW5YAXCVHbrFCt7HC1wP0zo/W+bBVThoPTy
2owkStR35nwtTIJLYkWXb5dnR4HXkLTEpU2NmOp2GZes6b9l34qqFCLfWeGeiPwUgcYk2QnUadra
w8BYdhKtt7lLsR0bbY+rQdhBRG9cbxLqTsxUfovJrxs9F3rzJQ7gg3bHfE05umT1UjPiLSfxRDgr
JVOFgNCL6adYsUlC+wiQjV8RE5kGEGL5nIgBd8jsB9fFR5rdixvK+89VHCmnxTJ06qPwW7ghq9pb
oJCtOpqT7QMr19OvR3aPZ/xmOdYV47IpCPRhRlS4td++OrxSfjlN04bZNsKK/fhzZfICUDrRbSIL
jj4EzaO4aI6j+FW26ABvZgbKp3srFtLwm88vLXqNvM/kEhq+EKxaRq588aKnc4TGEn91AlS7PEkq
BjDTW2khrUxNBTwT1Y+XFbhsnpGYC/hvfJvXissIkiy8IpjymCsBDPaoaY9npybFArrO/xw2y9Qp
Pb47apq+Dn9YQ0BwUXFuAF+ui4PO1EnckG15T+SpryfiwD7DYb1uCxkH3ZQb59xcBOoW5BSDSscz
VGbfB5F79ZOn6fLuNZmM7wsPsAib1pktS/1/zPoXH8G/sDVNwfV8y62pzAmSsmd6WKegWV4MHw6o
w1Ba59ErX+S4gDsRqscJ7rJalS2DN1Ty/7xMRIxEa5gucnpO/+H8E3jun4Jram42bio5IndHiLjz
RvUvdAnp2NQQ5e6Y9XPBIXHyBUChX8yKTPFj/qdkcS9ovk08BXThUFjDoi4IV9/8H3t/kHN1GwYX
X/mVycfvXIQDHjU0T/vCE7KqpfxAZoRXFeUy2Kx24pbqpIf0f0P5SjqMmwjAWJHsQV5R32qkWjdg
HUzvA/czqyX45E5cBHWxTFWHPJ1IT+o0Z9RYRVZjiDkpNAEK3q0nDMrN4fl7dBieYTZE1l+da6X0
zHGOEN8eSCd2KrdvO5xs/ExnNsolopDMeHzGgrZazT+dueREl4afDkyonmXdniylD9pMwD3bDNfH
RY4XcGJsFcOJS1KsYOMQhiCVF6OsIRUiopcHkALUfjGtyFvNFolVRTm9kmVb7SrTvJEl75JhJPpq
WOf4KIOZNpKLxXxxOadixgt9A580qtIGZCXjwSqDt2p/fvcJSgP1+bedUlZjCjKfQQTlNtwLiwnB
ZC+4HLMJ1aWc/HJfPR/jSRRVLnSlw5pqJyo73idyPmeBNtKI/sDGEU6QXGuUWu8BaqJW/VB7qFtK
Ub3IwQD67emo9Oa6vR7823ZSf3xASi/MLgkPyRVhjm7zowbgnT3AjRb5dG/FjNFjD0PqvNLEPTDR
/zTRv0kA8hPWrM3mCeDog3TxXREXmzHsoSZQ+Bi1i8xKvESHRXh9pYqrmLoKntGw3kxgSsD+HIs9
sZIREUJ7pNd/P950ICDrstbGYsT59QwbGlCFD+geFq6veR58e5frBa1T8Vc6Tz1pKx6VAribqXgF
+3ABgK7pbQvaIbiZ7QWRqOScCZ3bX7bE5myCETI8qg/Hsbfqyz2l2WD6FRwnMA16W3IkqZ7SP5Zh
DxCRjzOgb92PaIyKbe/yTklrG07iAPzKdkEyzWJYccCVyJ/Y+5uP5wTtIImhY9DqR9nyvmGmqeXP
ow6EcFCMKPfsWMPPNsO5taGEowbyWUMcoi6VL90jvh/olxiugmkNguEdO9rmNEJCgNyfg0xMDRGj
Mg4a3WBo+PO6aZf0/4+tUQwQf5mTZ2/FjeVWAh7aGPJHeAtVtGX5mERGI04JN0waGJfNRhXoSxjP
Zp0xJUW/OOGqFbK/nl1xWlPecUOIjV2gCtAqiz7iMWBY15wKWsyi0K1SIODzbfiXCLbaOYyqdgyP
mfLyx7J28ntwbd1mDD9sLZJmDD1IK5k5K6AR7Kkjkdo1lQvL0hi8/bycbn/vfCPLoUyQNCLzpyya
LzoBub+KNLFQVKOVXvIuvMvGQgxNZ6jcodeI8p6o8NIJEQJ/LtVPni7jFn9D76TJZLtJB9X326Al
5p1lUgDdxaKU67ymvAkCYR3d8jOhkneDwo9LaPMuWzYaB6PbM4iFjKETUtWRIeEYgChVA60fM4Lw
u7C74ZjkNhT+sYCStxpeIFGSPaDgrxT7YjJdjkgvOKaZyw5PNP1ws8KFkmz1h4Map7OC+twmVT2D
NpmO/wTGiy5n9B5Vk5Tx5Yfdwpjwc7BJnWXSROGOz5BF1x3uLsWHutIGw+w9OydpYf0BIFrUL4Ow
xnwJA8ai94B5DOWTSnJmTD7bxoS7E/axCUCKE1RozCy2hqIOR4jSOKCHdZDyb1JMyyrTNaKoNmiR
Y2skVKGa1hIFKWWwAJ6mo7D1dXWhiNV4lDKBL/NQja+/LMV4m/9VhFWheB3FKics7JNzH55oUqBL
ljBqNT/qTyMbzsHv1qmNb0xpHo2erUK+AmQCIN81C847LYTmG8/HKactrCLrusdKbvq7I2Aya81B
ti6MUk/caCsWlMy7rRWDSwSPS24IJLhRxo12kDMtX19/vgvbc3sNcvJRnRf4KNTdd6qtloAGqawx
WsN1s9t1fUa8aw6M6Cx0ULI0Qi6vNikNFtCTLsgBGnWj46DHx6opyKO8C/vVsE1tcPrm/8ogclJh
37+mWQ3wu0xC3ndSoQoknhXMQfudntw4HfnFTXxkjI/PB/SQL6NfFQIWVB7cqUG8Mx/vLRnFiy5Z
zy/p8ci2OgOcXv+Yl1aGdyON6SJQmqoiaGDzzkTxFp0/MpOMJW7uCvzoEcframpgp5BrM6I7SJB1
J+seGj/M0cOh0svptpJ1Dvw5XO2h1zcvhxpNsr+h8o2LLsR90rcipJ3u9gHOWyaBqJMogPBH3vgs
h+xy6b4hb/AiNPXD5T4pGcYd0sDks6R90uQ03v+kPzjMajzAcVszyBIbQ6HQeHLeLTVYvXG3tL8H
GTObtknk+82znpBB4nLPlgYFGWWvKOWhyUDKWu1+5vK2e5TsE18rHXqXLX2uPEBW94OZ9YvG3ieG
kzn42FeIAudglSRapDz3ZpPK6yV+ZlcH6z6/UK6C0iRxqiMCMfuslduvLqxEtGQfKra6u7+4Ccyr
Fgc60bfxkBWFpxOi9F377Fx86ac7wrg5jTWjw5RkmPmB2kt33ddzIyaMiJu/CeAZbCtL3ubUACIl
LrOZefb4xffMduFCisjAfb9qXt+x5Ya38Gr4AZMBC4GPuV8grTamQqbQdcvZF8kDffx3+INDlB2r
e34mubzQIHB3DTGqHzFEl70J2tLKIj5Wu5pKqYnj2bLDaeuqSA/cgCyh1vCJCkggWvIiqGweBQK4
oEfM8uRO6yezNyue9+dFEQmeHyNYZyodVWYRWJ0a8+4cMlFWWjeAAwp8hdrl6/oMA2ENjhkTSFEo
M8XcceEZ1SublRFBryvwQo9w9tERQ+MFyHJUUL6i1R6rFyuiQE6a7HMvgvbFblD4mFTOJX+YK1CO
ZQG3Tyu8JS93Ei9krszg3vZgpuovvV7l8t5pTVpBis/+NmE0I0hKAC4HAwmFzPTA6w6WDfAe8UbJ
uVRTaqlNxKy/dzxAiV47wos8QYlXP5vxpzIdVqnML4SqTZS2y+8lrx7u6tUJvVfiPqXSe2iBFbJI
vGjjeSwtrk+9h0mGF97269FcbHeAlzVUt9jEGRTdDEQ9iihL8RRzdYnb8o86PPAkEMZ6Y+jUV+Yw
P5KA+2Snqv7G63gLJF4FbLm3sqEvDfW/OK2a2VxcyxXQ0GniFHSlNTAro6QZkSZaouA0no+qrdPW
IErwoJqZCRYRr9DQnztmHZuqlbYcfNiuZTk6xiSCIWIoFukRM8ap4W7GgYENOku68GPPWV00rf7L
GC8W1n0QtEtTyZ14gl43ZmTQaM73VEYZzhv7rsBHWancHydo6ogKT5OdU/H9KQWCZcNpz+wm10kI
nbCBAGvViafeZJJntJCeymST4FyQTiGR66FTCuQhMUazgrdoRZM68Aby1oS+Ll2Ci6uSsoTlFgjl
cAnceWAVb0p0NOM3+6q1Lg1UioVInuo3UF5BCRLW1+eryeE4lJYPnzn1LeNoPwri8cERVO63Zdyt
877lbHxbzkmIC1qV+HhfOap/FCz+muFX4NMC2fz8NsEtH8zA9Kp8TSuNQJ1eHggfreRK/OlTHthm
cEpJEgKjtozkaN58EoOxTfUJItroyPCu9xAig+ZELfstrwy+6Q4JqmcemlUVYP1VKgYqaoq/6+st
04fSQMCYJ6gUhjevGPiJ3H6wb05dx6krBWAW7IlNXX+ZvdkEgi+4GfsHTNpZPrMG3hYvG/KSYDRg
pkXcQjAOYaID5P1Qfj7w0nJLvDSGnKuaE5sVXHTl8GEbxnVgvByjP4MfE87ly495af13VapKqpqk
EbXh1sRFd7cMwZIw84Ge2iiUIoBUWJNTi5kK6u8aPsGHIMqkv+NLgWwxTv2rkso5EjbkUPVuKVwR
A3mbnwZ5+HUUJoT5oN2ObsRIzFy81qFsh6mD7b87fD4Q/bIV8gAVOj7mZ9u3trDDXWa/dXWmRD+u
mT9VnKW26/q6SZDM3WscVGBlj0YG7WxhsPnhw/f7ZL3hLv/XIfp46gI+nIyXNp558o/Ktg0z4Bx6
i3fgkqw70U10TkQgAoJjigH/NecmQCA5RkgnychMowBMIezCWtOuPwvZN1Le9sLpPQKyfl10cmXO
XzQlPwaKQTkbb6PhFzFLJB8F7A6GUesSERLyII0pK8ChIqJ2nxVzBDrQNZdbdOTjuQtWPyOsIqnY
ZWcwH5KVtuP1gdqth15FI5hZ8EG+Bk8rQVgZdfzKAtmy8trvRT44Yjr97lEM7dl6r7OCyi9ALXxM
i1fQAI+vNKRMQ2ALx/sPTSbQ12VREXAcxNsEzkk0zLKJAt6Rw5xfNzQ2QEmxU8R+XAftcxt1PWMr
Jnh27OScJTOLxK6mYuHkLxA93OSEQSb6m/65vyDvZPkiWbAqB2nMmYRBZvwQ4fuZGs8uQ+rAEf6v
zcww76aWJTQc4rlM1rlFt6hs0vdAXyo4IkKCxTiH5lv5jeIUvrW8l2Xk3LI8T9wIzz9RQ4d+a9Jj
KLdMJYF1GOFU+Syw4wmkJ8QOYZFPuBZhIZo3cML9hn9DjYnj7aGBHPkMO6g/9CPfgNPF+H4CU+7a
SwH7l+Lawbp0UcDyEd4MYPaRAgt+4BNWKsGYtxqJucBHatYu1nj7Ekt34RrNNvAhT5/LiHDpgb9F
QBl4qBMJmYPfqLtl+ltIOvPrTP6MpAKe0laZTJqI5sPpbbQ80HwktQ1D5OYl4cRS3038jC/5AKTS
oCfbOLVIJbT0AE/8MDgYM7whQEdBb/k5azQghKbUc9Px3IcFaeHA/OEtVLzU4l9nr8Y8/cpwRIVT
AzMQIg60VZEl6+rrXvaBvaXiymcMm1RDIlFEU93SPv6NyBpU272e64Qa4eV3/aVSIQkLU5URJWBC
0rF8HeQdgiTtOKsR/c6houlkVq7M0Qmdh3NLjoE/0R+Hst20395uswej4EK3srIN5AVBhiG5CSHH
2YxPWvXUb7/8u/meszdcF1cYjytuHWNT8j7+S3NVQ65mfmnw+p/qLsLzIARSdUdElukCe5vEcLK4
Gr3xXlJ6SbpnttBP6NK0P2dDI7q8F2eLF+9Z0xBLIVYYYcRVeMKSc8X84HirFXxLz6T0p/8306bf
1mrXzcxIY3yCrfFNlC0XhMi4kXqPtdvmpMmFh/JpDzHh+4IVnKjfhMYlYlE9fxrsO+k3lrDNk1xS
5kw4Bqq1NVudBJ3Y2/KjZw4Y9VPOEDmy39+H9QHeW4/vbzbWYhTzEa1RfdiVSWJZOXOevfoPNnm1
c8Vjje03Zj1RCQOHqXXwbjptgB4yFJ4J6kZVv6KGbRjx2v4MH0STFhGsJduD/u3eBPV8KtTKIycW
OtynvHK/9m29zx6KuEa3Ltiu9V8D4i9nKrDw9oDUTN/yjiypMHiDK/w72lmbz+v6cDEB98/Iqhks
DfF3o4XGYzCmPZzu98gKi9RcsA6m23VJ4qvJFrSBELZ+CGt64JjgBBmxkIFDf9PIG5EHme6mN14f
3rUM58ZKUoGXj/O+6YtjgxgyyIV+2WrixP7i9CI5xx5GbiSolm5fg4E5ZLnhmf3KDFd7GV13W9Nl
7h/78xi8yl9CqsSmOgUXtH+/uLO0nLkiT7yPG4mtncrOh0YBmRRnioUeMfFvW0+KSEDFmK4rNYyw
jIs80+wy1eF4q16Srnqng5ABaGz5Foz/WuFhYUZSmPEiLHwhStXJ2T2OyvkiN4o/fuOtq7Rg0snA
cRjrsk10bNAOiZbO67WL07LZTgI1ryO98+RKd3LzpcIJg0MnT1L+L9PXGmJbLNMHvVnxtfzaXwzk
CUs8OhirTZouXz1cqfqyRw/5qL+GAsuiKW3sn8JkgvSQH8uUjc/nsjlnoXs2b6cvxyqry2doZEEe
WvXR2eYmotho37J9NaUnkrkLJcNeLyn5ftjrnhQvx8LWvBU3s3OG7gpNToqN8eqz5OXVf74+5npg
2Xi5zvncVsd0518aGn4CFfdRqZJwvyk04cVZhyZWWzlnttyELV5P73tvYCRRhq5QQVUAvpAg/7Z6
WguhylYG4RzdYz2v5sxA/I43xRHbBrsPrRi9rOGLk5tFUaVXSmHRypdVIuRI7xaXOZ0IXffKYLd/
It6JcHT61972/quvDOeIEUxJKW+7ClwhSG3GEtqEJ4MZy7vBwC1YG1S3/U9HsAb4N9PIbxLWdzSp
6nSP0q6y84RnDrTjvEYu8n+Upe8c74/BKkgwQorsXmr5w/5lzzRDPv2fg9tRwGDg893+Fpg9K/RS
YFy/UwU+qZ8djX4+e0swNrZnKWcapo1gUDQYK6bpn4MFQA7FPm7Zy1L+/NAhpwlPpg+6MMLFOnHe
iGO9BpBCH58FW68/B3qmNLtyykKzZIcWIYxfU6/D97AUR27elNS5AswLDZ3XEaT80gKjkGaRnHpF
7s0zyaRRrzEd5C/k24mxqt3aCkqlS/Q1HW6YM/kHFs2SYX6K7uk7ny06rl+41a9QPbu4TrfKctB1
uiy4muZevI1jqE5AJ/TsyFpBaQ9t9j4nkjmdX4HZ72XcoI4MlSXDqpHFPFbsKpzvst8n66l9Ts6E
FHmt03BGjzLcLIJiwNd1VHSPzXjD86ngVf3O4K7+pWd5jbISOmxEdoSR1oi9XMY510Va5SN1dE2M
24Wr1go4JFN9mN1BhWOJLhefdyrBXLb8MGQpl4JK6fpSwXlfDnD3H5p5gt/6k43oeQOiKwr//djk
M7ncfFPm2byeDYpZ5w7sh8RMeTTYSoVpg49vaoOCAvqN7CZxF0ya91Erhj1MZCn0skD2N38u6buk
eume4+WoO0PZH7F6sdPD1bMoOb8txORgioNJelTxSzJmFP4smUXWV0PTGYWErqkPziHJsl31uaYd
d8RPd9o9IWHBkRJeKPDrfmUY2Bnm6ZBKw2hFKEEWuIRP5gHQNJtUXl1iMi8Ua36XBIDN69vnxvoI
RtRcStOtEPvtP2y8To11v/PthhZtH280/sNc7eSrOdCDZLZnZI7P5paSSX4ORflCjPZw3jrdURiL
IlBTDI+qs3dGumX5gTkxWPJPhR8/Xh4I5EcZXxYoFvxEUauFbW6+pnl5q8wjFn4zWZtzAK9tCP0Q
J8P5veYyQu/jxSAMCatj1zEnSy1/rFT3nPPuHyHCaX2air0nc9d6gu4dzAQYySxiUyGi0gnPTr+K
7ebgEZ9JSr4R/DyBVFfbPd6h102mKkjK8jlg8SNarhBorP2FrMsE0f0bwD0k3mw7TcmrIIW8TUjq
2o4oiGjHmxAMWOUD4ufFZzCa5y9RXAV1nqcm/a//paTtKuyDiB1dK9X1ZAfHOcI3gCu9u0Yxyo/I
hJLEmZx6PoYDJPuz7nvhR421nnE8t32yKuBCTHRHFHei/XLF+B0Y/CHCvNnYMu4BXTQPa8q7uYmF
HrhVH3M9U2KKqhcSWbsYT2615gX+Ji1i572broPLfuFjwsHSji+ZLvRm7PKy8JmLw3I8eLQ9K+JR
rxKuvgo3XXdPIUGALQjxtuP5AG4bWQOWwRrUKvO+q1LM0qvzoONAL2+nyUro6xBaVdW+oLIuOxB2
zL//AI9fJmbkvw+bwOpsVPhdszD69biKFBWCjPHOBr+WlpOAQwqwW14Wg9FnTsXcG4uMnKmdf43B
pe8314zafoA9xD0DvcSDbEHbdI2e2OiL2PmR6U3caY7POB2dRXBglkV51gmtzsVZzWMpy78QYphr
qyqrcWT4Ythxfa71Dn6haZxjUU9kJoObA+8qaARI/AOUNVDQwWiDn0HAmthrIw3mn9xqDwbNVJSp
IA4mEPeNraIJRhmslxuVJfJYLe13uf/+siRFSwaFA7iW3DA7uVHHmF+jlqAT/e7wgNiH1CajdwgO
FjnDIz/NYAPh3mqTP+W8bRARExGWK1Nu0MESBxklFUx3PRPnBPutjsrJAAvVFUoA7X+9bNRIEwyg
ytrm2qlIlAnWd4eCP+xTfi6AnRyuyYd8mJjyC0e7brAIltcL61MJX5manhltwlR0DPyZFIVL4kVA
4T6IlN18hRycjwhFCI1rkPKFtYUvR7aEWNVngqPL4kNJQNDiXbSdvOZzRu6ZA3qfgNGjJyj2U1UR
ci2bkZbMk4aiei5SaqKnZwELqJ1SCoNsRYNyGlL05F9YaiEcYDmPCU0tlRj4bXhvfhMdFssa7/4r
9UBJssVYMhmjtZ2jvdFaxt66zIe4DrqY65M5rny/M5nQDWOQt1ji8mUKe8dZqu0GXxL2F2Z6Jrz/
g9Tsxsv+YXPHymsErTqtN0RK7iMwrT7aKZUi3NQlAKRZfbM7ANk5umetJP6PoB6E2DukHljmuyve
73bluDRiPp5RCyHtFZCxVjD2yXRlQ2Y681IQUq+aTOmU7w+mjRi3pUpKHPk2QOUF/s4NtD4lhYBt
wljzNyIhkkwwqcfOhmNWXZ7oZ6CNh6MPEiKR5ZKS+FpqGbM/k5OVtVuirow6bp2DoZPluefOwKEr
h6u4+bg74hRjNAqeSfW6v5I3kDdXTZx/fh0xWF2hijyQer+qrNrfqvbomzd3eq2jZL9muFll4bES
pH/rc/wHdRdzRfP/cmXJo8uMM5+NAAbZfFfg+Jd8vo7PSAWuv62fnouaJ1k2tt1sA+BT6PuigDsY
n4jA25DMjkckbeJ4yrEjHfwE5nd38hVpObd/ScLQMZn4qc/Jj1tnugTn7Se4L8UOwbnbnLrA0c8m
pyc8RJbQnulrZndrP7wJwQJ6JTqRDFaf9fIswCzeGD3k2tIosU6WW9N+KybwSTVW+OTZXcPgq3Ps
ZXZTq4wOH4vKXLCRWyqWsl/KJwvfDf6qZGjM/H4GwLS7KokZRtfcma5dIjOOkVVWsvK8yRlfE7RV
MQK6h+ZlxOYODvLkMyYn/ZPzZF1wUnZOvLFmkW6y7GF79iGSEbZehG2iZxFjGC717KkTVlMpDz1G
BwRLd4/FBt71O17JmAo8hJw2fElKnaFxcbtKnDvAM9TFAFMJQkhQmxtbEJYhDuSPbdvGs4yZx0YF
EgIyvAw7/c89HzF+6kFL+w9I2NCiPcoLj/EJlpWVjpdpfiTlcMZUTulo+/6PSj4orOYlYSPES76V
JtPD03eBwHnwxTF5mB/FCtnO8P1DH1WRjWUoPyw/MPT/afakvV/2pKOQPI8a4rbjQeA1O22mdTzH
pnOAyrY30Qh0YUDBv/jQXanKf6HadWas5lEvAFBPflwzLl5RYlM8lXw3waJShWMn9clOn8ort7t2
5HJ6OnLfFJuGOQYBhCJhuewB+GLkdp4jG5+oPV3THzbbfP4vjUVelUMytlt581XpEInwpJRoVmOz
cNlkw4ejmlmhZgUK5OYJ7XHly4j+U7JIHh298x21rpAHuwu3mtSCel9jYikUqur97lD9vWFZyHUK
WUPA0596OqdGstLBogtInkY34FnxbXpQspj0ma+ujtaqHjb/VDIoMTAyQPheHHoDsmxocXp5gXKy
ntvutWqfBDz6hKnaJ1DODu/qgwv9p4UeDnwN77zLmr17ZChzibnPiLPoB4pHFFZUmmNv45NKnmBb
WNbmZjB4VgPZGRTxkJEhOhZ91D7kaQMEDVpG5QmiV5DE3Gv1aA3EB+4UAG99th5xyHCEVwaw6jcR
a3WXsFOkCZn9o5VxgZnYRw/Fefby1r/cwpzVX+UWC2OPsOONFIyjUT2QR6jqRi9phElzyLoEoTeX
jcQgJgNxWbnrduQ3LfMYPvNzk3hzdUBzCRnpz3nbQPheMUzdhJZrGNkW7ugceADw8SmXgtKvroFu
PxxGnY6ky91bTdjwSteNy5Z78m3MvXhismD+di1fQa3vu+Hb1A9emfMR+FbAUA+U+9GhQ9IHTgvO
1BNFjUdoxmvHqtubZUc79OfnDmIARoLaUxy8GpU7Pe47D2ExelCiCCI24GH1Mx7mVP+zXOQ7DgvO
/z1B72OGWVWKFwUqFGMdNHNbj5iZEh7VK1R49qvjb/g4l3uzmBq7mbCZDGgomZ5eAOLvmnkt3hqq
VPsnOLTaQGgtJBpURA98xSEULUwfBYYZdxE6D60nqBNvhPWv+SCWUxlw/cHb7Jp5lAnmrYTNpzJo
sUKPBFald1uJ0/D1BS+vhJqYgtUGWj0m+w/L0kdRRmmE8EpnoIShNoSL8edx+O5rmB66MJXLcL5G
0Lui2g11bzzwz0bn8b/w9vvlP3/XSLli+apYH5vHp5JVNGOYmmH+/ls038weMOfB7uUJQbu9BXcC
fahaiUPgAElPQle1uFMzUmL/IssesXFA4mZfpJcVMwUDgogyy9Zy3Vvf4ofRyvG6+rDzu2f4h//9
8Qnie1GGVPPerC2vUgcB1TXMsQH4F9pEq3TMIRgRrXFWBCEaOmy8RwZ1fzA8f6ylgEgQ9l3SdXfg
CMr0DNk5XbEYYau4VL4hOQ8aD3deqh/sxyeyQIu5mzgRB5UoEwuQLy6ZTwhlQR9GThv/YFdktx6V
tddoHHLaF9DKiD4hfTan1LSRrORYblL2Capig6FFIfooeIDLATWYTJJLP9nY3KDvXzMVPfpWUFZ6
TlV2Vw0rzJwP/6ckSzchvi0KjsyRn6IjLR0ZOjkvb7cP3zF4aP72+VfSloB2C6Y3fM2aIcM/WP6S
jJ4AqZlUwo1oHS+T1l++ucisZVH1pOHVH16dJE/TPF/L9Nv1w+8lj7hePLY892z8ecWYk9uNjzni
TnMXcI5cEGubfjHGzfHGgfMApSsI4XjcX0XzC872IxtKq4lQfrrfdDtanGwEYAz81WOvCOy8Vm+r
I/TVCg1FbPB4YBY0iihzFClPcW7bOXPdSuRqaLukzutn+CaThW3cQLvu7k1lrnS1vOvvyBGGKXld
CiAqt4N+t8NQLJVuUhB0xtYp9NJNXpqmYVG0fWfTFOs19xcfxZaI8IZn6+nXGpqcyDC5dvQOo2UJ
xbXTQzThtKl3MK+GP2hOX/xcZug5QwZ6oX3XeaRSx9QKeZ3Gn7pb12ZHyW+Fyn/6smk2kyvswsHg
8+YiDefaUbDTuFXLzDtSgen5x1mKqwUbSGfHNX+bcYnbHzqV9cjopwbztkKmSLUznPnqOS2ph2z6
iO7vOcF66Hd2jauX/faIa6k6GBTUx7wOJx01+a0DTz50dDLPEWtlyXSQjv7HW8fMqaUmBn575KUS
SZzyWB8OngmXUqQ9OgRBk1aeiiAsV1CrB/u98MszZHMxaEcno7MswENGW6I5amhJVtiT3h7dE+M/
9cMqLNHoYjO3rUsi5tl3SgThMmPQ+3XCfjHpKGqtChNMSqIGAzfbnfsduoF3PYL2ePWGDcOCz2Qr
HHi0wYyEKrC02/nYjGoyiy0SDtipewrGe3Dmf0jkXVawe7yXPGyi18pUVTpvAz0LcrNeP42Tlsgi
O8U+J4ynQovRkdcCPAvw5ZfU+ivM2HbuhDtqm+OwEeJAeByAuIhHYZrFkLnuNVh0LDCkrxJGf8SU
j47w9+WGHa7p6LydyITbVLUuihlHpSSQevG9fVR3+Pdo2l9clpxvzmVfklAiwpW8887kalvNDvqU
4mIZPEbTx00YfWa1QVxv1onOVIV/WQk7EBMjdRKM/za5Ju8nY7RdSQzkE7579dZnmDSvkmL68EpS
OEiTBflxJ9WLuNx4Rr3lHhNns/nT3kuW5Rct2tM38D8Hkz4MGqks7/PKFpPM8F5oWXVWoPIhhwnF
vmS0AxHRAHd8xOSUmQnhp2BzLoV65OWAeF1sfXfWud4WFaN/S3QkWe5SPkATa5IhPKHryLv7xBXh
3/9EZjPvR242bGhzU0sJsl7eetfCwXEwz8vBdTktiIIiuAYvk+jLHDWelff4SEZpZ3ugOIkKFByf
2p5uMRqF1u1Q6Cb/PHNyzVhQph6N0lPmMTx4d/N2xRQbLnVOor/rSzfnbUVJdEI/m7MsbtSuKjC7
6C5jR+QmqqRRjMXKMOvRW7HOE4sZudGzWtpDvKfCWZF4/MxsprYUcByEAfQew49erMlcFxArdraR
ha7cJat1UdD+lq1nEB3awkQ2vW3Eltak5HJ2KGQrNne//7LkmCz1rleL9TGp7NoCmjU6q8OA/MrV
sRemXLQ9XScFTDyXMu2g+ArgBd2nVRrjP0Rec9D1oqfRvatrmu6gGNPeypjnI2dJjQmk4xUf+TJ5
OJz/0z7ZSrO0Tt/J1lKZwbMWZUSU79TD2H+tiwJ9m6gy42VO4YZY6Hfs8CQzOzZV5Y7jz4PPb7hE
YvFfYd4U8Kqv++WRFa0KvWAMKL35m5UpsNNFhB+uUD40CGXS52K9dWug69Ft/N/PxjK1CVk56T3L
mr1j9NV56Hpr+3tRDQbgJDPMnVzZkSQ9EgZQ4KTboij/90IB/91WjgiVdQ5fN353fZtKvmRaobOV
7v4M+WjjXQ9N3JZD/uliTHGhzyWmi2OwoZSP0ZFItRAAY/fSxyjTRCFslqHDTp3O3j8iK6hOn/+k
nYkzFWkFCKbJXn+/1A0fx07NHnJhevQWY+Lme58NV4zi8JiYp7eYY8K5dH+5yUhhDhqMd5r9sHsz
TeR1OBAzLvOpyMkJ2L3R9FIVIlfp/bmckCYZoyzIiKUcuYZwzEGHv2otTvgTe9OUd9sqCNik8FRa
dGWWM4xJCqEx3hzsvfhzhi9N6Z36iSb/mnGNT7a3/968ZI1J8Vvn2SWFQWVmLm2FzBTluHrCqYlD
EMWyLJipNdWsR01LEl7ppf7aX9DTBGP5uZcooTOHL6vOJ7vkXYBUVG+HArNlXlo7+uWKs8WuUQFT
3+X/247tQ3pUdgOouZ6PLNCezDe3/qHowdG1fD9+ZlsmgKCV8lExitWhuZdF2mQs7EZkuQEwEaN/
TJ+Y6Qrej4rK7YK0Rqg5W2oUXEpKULOLhWBBotszte8J3JV9S72S5fdoALZpbpVxFdrXMGn/AZpr
2k3/ebtfHt1CJ2RxJYGa5a5P7q1i37+3BL9W/L1zIZaXVD+oK7xYqw4Xk8lL8gNpiqNhAdf34V7L
CYyamDdEqizVPm3tVzweeu14MNsTLq8BWPZWnUBpcgq6Lj+u2L4UQZ1sJWMx+YGMB1pVLBbZ9dZb
woJxpo0CpAy4+RpPspphiJWGKAgzcKxXXkk2w3DMH6LkWZF6fWJKB/y1j7Dcw7sHQAKG0Kbsl7Eb
jiksx+8F4EEnz9e73w+rSUv2KwHDklLalx+zzeF/+qSSCKLkAqTaZ5qVX6iwiWQ+YEqivY7o3rMP
GotxzfGi/82S2SOfH2Ig9JGPT+6Ir284sxdBMSeHsTjUx7GqdJxEDLEOlIe2oBwNPJKq2e5DRxU+
SeSyXpfnCI2dVAfxwvLh3DSy5DZfwLW2FpxUPD01AQ85gqZmuP+g5g1+T6xIfZjrvZ54u2367bC6
eLEyoaLDBCMcv3RVxgfykXy3/4wXrzrDKsna1EDu9MQT2H4P9NSwsTfgTVx4GCceZTsrwTXfAH+n
Y87ILlra6iRO8OIhTmRwgc8yZt2TiWC8Tw0+H4YnZsKdGjpSxki6zjeaIR5Lt5H5l/dc5881XWi4
a03J8dT9e6IeAyrzzL0CxW2pLzcACGyLqgA/Lw/XmvU3EA/nskoih3UxovkSGXT57pyoAu+UJ/Sr
0GGjJkbVOSU4nNWsMPi27QfXHaNRh/DUXxEfx2PtpXDo4AAgQ2Xksm0rgg/nrkbbMhZ4Km1PD3kp
cTkzWUSofZ5ImPK539G8hDPatfq9ZyqcZiYT9GmdfqVfCHaUuHlfhk/+FWSPRjp89D5IsrjO7Q5D
9Y5to5JG4F3b+KCAXhyZsuZ+hLwZPuBf/56eAhA9aLHE12ZmNGB9EjgWg9LHC8DqsCbHj7f/ZwrG
QezyQjG2SzNbxFIB5+0nDf4UdX8a/G7sBma1Z3az+Jw+eUBVZ+b+6XPp47SiqY2nuYdcKxJFAOOq
VbThalsmoaZCLMVmNcNB3jyTQT14BdxGu79+y1N2ZVei9hGqJr0c03SZWuNnhmIw5JuN10jst+7r
C+YWQEzqUj/7Q5TNm8m/VHLx0HaL11D1wdtoQ4RglgKgtYsVFm0p+MbYmtf8X67KYtldteghCpVG
r6vsfXeQr/wSPhGfGv1gjFjWKM3FTmQWkfqD4F1CD7VKQmXDBM1MqxEErYNvah0RSJW41PSFs3e/
SnGSXh07tTRemeMIMEzQomKof4tDg0K5JjHOmDP+FG9C2a0KONI39r/rVTKfCTppVUDvMjHux7+o
wzgLcTbboYoW+4m9dNjKZZ0SiIriWu4b1XqMW8GTPKuMkT+4/VKXMd3TqH2W/ASxXW2bDeiNht+p
lwx6DveNJphMUfSFt/M2QVmtE2g1RoCYoraQT7XdnaDt2f/bToeSSrkQ6PUa+4XzYY95NI618o8k
z/pe1Jg8S4r5dC2ZWf55t5HCe+xQQVAN8n3HudMFEoSNU8h8WJHG/1pIx7GRj0S/z5IG9fvCU1gd
/Dv1wN7ZjZHSR7c+PvjelvyiZCIO02/PpA1cBKCMJuw8Fi0I2pdykQZVfCCdZ2LxULWWrqQ0So4u
J9l8t44Bg8xFooxuw3xmh9F9YeqOmHwUM9na0L6dT2ELdZFOhHjoFq/ItG6m3Aav0bqQp5RhjVNi
9Gwhh909Sy+dT3E1L5loOMPaIeA229ZdNQBNKxXpv/d35gB+bcWebb1PM2ObvGSvdqPA+wzBC+Sh
2dgF8r+s86BuaR9NN0K6Ht2JNresU+XlLnfOD2+RVZrfOWUG4K1ZfqsE1a42Zwa2fs74ADQawLD9
hzDB2gHeV+si7CSnWgMiN55q01gG9jkqZcfoqhi9W58LvLFjhXDEtCWx9cWWiqpjEe1an2e95N9e
ty0tEUu3+t1MTMLqwCgdwRWOasIGdK14arZ929/cAJg+HS+g0y7c1EFvSZNTsxUjxkLw9jioVUR8
eKDsbF7zoyWlLbairzZ7PfWSaXQ2liJ75H/80XavpGTx0HOStYnxFImwgf561LGt6h5EfoipAlY9
ftYZJmUfDQ2RH6zA4UN6FBFm+1w6zLwBydKU9MX1vU+XZb2wLGL/7fw+YWLYUwvuTf8ZhK0fAU+h
+Rvo9izKlv5COCoGlW/2M98TZo+DL5U6taqwnQp3Wc093Lr7YgngqjhxkELYjvU0+e1TvPpYhjMH
fKrSLgZe9pxxc+I8E6yxT204Ksg6PC7oAGJEY8FmS+O8uAKuoqjJj3PgJ5hQw5TXcIQCC9YIZQlA
zIKiYgSnlrk0Wy8qhSHcduciyp/KKzTlg01fIED+CZkmIkC1LdbH89cUTEhXdehZSTIdChpNxYL9
6yZ1bcaLnvT8Jpy0LVr4iBoGfda5/qQB9N9N1CmAowoa/LkL/8mnIyQ23gFX3VERzjiSQ37JfNmT
DAiqB9ZwxgZGkC+Z69eNgXR442HwWa2UfGo6rS3cXJTlXa0milPRIG9xkiednNRSN1b0Mkbk5/PP
uVIWmjWCfTc5az2cdVxdx78/JlKmYQQvK+x79Kbuoj6KFJ9xit++iLA3zKjSrkic5Gv5s6bHPz5p
w5QAF2nmr/vlckMCyZOhaZNg9k7SKiHyHlnlhvLRfAMbGh3xK8q5f1yATsrXEDeQO3mLkNP/GDhT
onox/J/AavbKrTo+HlPfIVz+DbWXjaUGwAJfQcHuuYJy4gAsJ1UAarYRq6xjtlDKZ4Dt3mxw7fAa
rwNX4hZxjv2QCXQRgFIKlhz2F17Mv1N7ElNVj59bdpPv0cpp+X5hWoQuXtmDF634Mo71SoTxJm73
euwGsHhX36cXbgn5SYxoyOUltLS0SX/V4e5077syoLXC+EXka27CjAf3BijT+o2dzGFEVSLjw63f
Hoj0o5yqbwr7gjqMIX8Q7jfQtc2JahqwzKOksSGg6ULBRn3euVzcN3hRlW7oKAfeztoR7dlOK8/e
LvdBQ5KQY0AgH5tT4NPoZVVDVRDjvH3X3Ww/PO/krHrpSa7w91NB25oaYKxzafhHbsTVeH3rrO3m
zYSxUq3eT/jAfV42YZX+BfRQi1nmvDDA3ctnAliWMDbDu2JMku3pUsZaGHnzSmBuaTo9YN+6g7JK
5mRpzbSNCNj2xlS+Z9oDOhaaEM571J+dM0QDnmATpY/02V8EIVYMcbMjiyXl7lAgcTf83X1JhSFW
GIcgbT8hdfcSx6gQd85UmnR65n/6pujV2fbtEI9ny8nlQkmbdn+ws48MUKVsSOGpHchMv9qvjaXG
mj8JPgCrJFhw3pyh30G+UNKpmXrIo3tJYjiGsr9ebpDXm2K45/odHwmz2e81oEzCeRH8oSGxRU8K
kvj9EvAWBehDYtrPg4Z3ecs1pdXDY1OCx77ZChO1Y5OijTu5wMq3goq0u9i0/DnFST9gOXKWSjJ6
hUka9bfYPB2lpbqLMgHY9rgV5928wAFBWwrJ+5/0cZHgVKLOdeAiUsX50ZWwDd0atxhM0bck4tTy
DtpBlnwh2wiywXoh7Jngo/5zZn8PxEFXKAxDSB1Y6ElV6rLJIz2gbZNFs6NacrzqFdUl6ln9fKFz
QeDDbVz8kt0wGi/SK9k6m9rG0gboeDnBYN7tnD2gq12BKfV5EIi9frwyXBzM+tS9lnBwQ1P+0nHz
3ObWzYeMhZE+KpFG/veAZvr54yMqbZWsvBMV0NjX2UUpY0e0uLpCVxdqAjyWBW8B/mNnSfcL2nf9
1UYCufMIBAfyfDDhMzMFW4C/2JH1//QNs1d3XXbV7pE5edGdxgEi/ILNVn9kGf0R/V2dclSM55uf
SQHjUyyZFkBGgubA9Dy5wjLEhhefLzDQKOyGRQkP5Xcp468AXMBRtizGqJFKl5pTFpi+jkXy24pG
OA1cW5qcLG61NfUuR4qtsFvj5nROv2AXOCYh2DVEPpQlIBDvp1/ddel6i8hfH+mOQpxM3BmXWn+N
SU9PUUslvI8ATmAL4lmWD3dp11jbUO+vDndGIaVdIhc6KHkJUBwZdpzYiX7B8070dK+TfrM/y4z/
6/kGY03zO9KbC1VrK2zFuIl8pqpa4tYS7Xe7oC54ma9uy6Ri/XRV9JmlnEz/50q/47mYYlO9zfFW
SedHHlKKAl/u4gOtXvK9BSN3+NsZytJoihR8XKUxG0/IziOlKLaGgpcq3Sa3RZg3nt+aIkkXhQzN
dmHWftx9dG7tAQDwi62HUeqCaEo7GZO+Fqk49e124cTtaLpnEP7+OcNQFylwerRnY8iAY8wk0niQ
GLUmukmVcfPdaWEAhGF8p8nP8riAv2UxK0/I5tuxRGYe1eEGLWjBkAYS9BNzxIZmPUDmc7+16UN2
hBhC6S6FpknPa5qZshdY5L3DdHfq5QCiSzzegiSgkHx/19MYfiMbHcOLRT6+qFWC82dABQf+/pNH
qjX7Obi+FwBnNy6jGSwS+M5Aw7qk8Hobhjhfh7aPERC6brvTJNrVyx+3wEkvdtP7mQaT0XLo59jm
QkmDkZucjUV2Xa9QpeYu1bV14v+aiFVdO9Qitopo3XTKEQU+DOFB9jvoyXnBRx3v9DaavqsMWKFr
Mt2HiN2R6QYZWDA/e3A3Wp4GKCIc02ePVjNyCwod++pzyO45xlXteyYy45iIk65B7JSo0OZO97v9
aehozXnumGjcKHkJ+I1ddEqioL8T8RgVzoEHDayckuFtBtgnlE6TaHG1kvNp1BPiPYv2ijeRZwAf
NmWOXhpkQ42KdZaI4vYig92crIj4fkCvIgEPyMweot8G/KULAorvVo40YQdOKOJMTftz26ctCymp
wd98dvIL5k0w4QOzVY6qyycjmtz06oksHv9Nm5i6OhpD8Zf1qJXtVyLhLkKf8nXiqLSDzqeVq0Sf
PDU4nOZKVOiOxWHVwQQCvBfAi/V8mgi5CUcWHx3bVb8H+CI+ulwcL9Jf0jLt/aVx2gyvqPE01x+W
tbnauPmqnhDmmmWCJ/JJhD8kaXexiC0DsflU2y546rECRjjoDDjwnmu1wDQ1ZGnINVDlmG9oBlvy
gf2hHDuI52lry+4hj2cUPXH9dh37XwuJAkGqZCM9qW1D/fiinlBbcOrkFr7Q7roeOvbSwDCGg8pn
OvZHSzPMUemoWr/1H28vsnfVnMOTxM27Io/KXV3idhzv8eikRDLblwkvyfVkr2l2pnsrloyngDZu
w9EMHfjxSNxzhqgDCg4J/diTs+R1ESk4l5gqDF7WDuTT2idwlPIf71CQSjpVz8qIz/ZqSNrUFZKZ
Fdq++uw5wKEEzKcLsVEKGHkKV5Bsh/yR0zw9zwTT8DBI9TYCo3Pg4/1vZo15WPtVDbadXNiXAehk
c1EN0sSrxHTysX42qRicQWEJ3OCzXNkXJAue/FIhlTcabHRORj/ICW3thMQjJAylkuZYlIE0yNEX
SELj4iAc9AjfvfS2YeReUdTYz2djPaw//lRmV868kDCKbpHE88IEjbr34pVwInHu4w8iaAezYidz
Xvf42dKb6VDw4vkxeDAnUtLyrd1P28qRFKlbF9lQWmiBulPn7HCgDmtFa0fsL0ZrTsk+N+EcvD7c
cMp4IbXU694ww7HuGeF/6prvD6SL9xCbgusTUblTFlO6FjEb2i/x+Swt71TFSVqtcsS0jqEbJ/Tc
Quvk9+vtuz+oBzC7ZG5qdDQkEuOriJ0X/LOhmJvec4pmk/XwKsDeDlKvK1AEFhijIqzDJ73R+9I3
YBnGEReh8VskJ+HZNeSBox8dGp/JD8f2tdck2Kui/ix3NQ2bREy60YOsNhPvlzj+67lLQDc5MRqk
4Sf9r0qLWrF61Bvbr8b5nCOPx5DI/pmgxE/tt+Wu+iDSVmQyCeWDOYALIa5AyArggM0qRKaLv7Ew
VNGiV97lW5saN/Qj8XHfMd+S89rmbxzIoueG3vTkVYESWNz7sS3GBRo+7UKFsmNIUPR+okMfrqaf
xV1bllV9Rs5VPiRVymoTuHzKD0XOY+gy6KjYx7pbAy4/VYzG9SuRAXj3eO8iFB3+UcAnp24fHlgd
0YcXwxkTIb10nO/eDN1ijPuV3+AMNO6tZiFwqmbYGQrVSQkm4rBxj+t0gHrVydtxH+/rFPtg4hlt
RyQJCPMwpuWY2nl8mED7JgbYlePU2fVFMZo30JvvnV0R4Eov2S+4DExhvLiX5cfeuWjb0Eh3vN7A
B5ut0L8rKf3Jawr3sGDbcR5ZL8rwTr/a/a52sEF+wQSiffbxmtqDHYLpZBENkih+cITo0Uf6Ew+T
4yAPydKfQfirVBmiZtHEhflJfXlZJvFD/Pb25ZDAo/7Av8YjFsHMItkYgwggdc9kfLK2AdDtiS0N
aZ+1pCLVATWRDyggM2GNSU3gVRpHSLo7BuMlNJQ21RILfydyENlBlA8z8aMa6AIDC6MTyY0TMJE/
Zp6FcovkRefEFpjQMffloFQRPQ32rZa3sCcqjJfmUdvqiei3uV4qgEPOmGfw/g4aSP8XoReBsIST
S3FQsZPVvp2hgDmOlLSksIez/b/Hf3i+SBzAbR0B5mkn3vxM1ArTYApTWWv7uZxj8QHPt630EBgt
W2U/nfl/VZrB7csq/Q7jSH7HUl/lGEE3TNDk1rrUhjIbDqfr3SREVylxeVMhyKUEH3X/TMEJg2FL
mo2E2W3tH1fkcoxzlITuvUIjaXyPQ+HgGxQwYafzlr0xNN9IYqk5y8wjpn2Z9YrlrtfWLq3Yw7Y8
yZGXcsY/JJBZe9UlsHA9q67HrfmyvddzHO9nV2s9GFMloDoeEXOq+4lxwj8T4g3uY7zGGyXnOCH0
cc5eoWjn1CSXk9CuYwHbdOtFXTaXTdoxvGgjav4XOoa7UXSqwRNqwDgfZF9MgjNLVak2qIJk+S8o
ytvpHSWMh2v9tohHbxSY39F8IR0XSrz6GJLVGG5QOHof58qXWKqEqGAM+P4Mv1oWFtF3Nz+LK0Q4
MXUIOeAaX+2q6eTFvH54j0m3i85Rnx5gEUVKXqsLfflQ51j988vQvrBqcWb/MOYExBEBGyAOnLSq
vt6hQufwWtnJt7hOym+cCZE1FFmwY74NnqfCifVXUuggxrFJfbQ5p+nNRz7wmuptmDYJIn+vn+Ms
kK47ZpT9YdZJ1JF/4DpqaZ+bFrZrnrugMWv2jhwZEOFb9QRJK1wZ+0FoCP8duOZwWgrQxgckC3MQ
BJ5S1Pdja/f41VXq2Istep+NqRPi1ZPtNeewxe4ynOl5U0FPQ0gsrx0iQnvcy9VRFOsskbaheLTm
CvhHSp+ZDCkCYnBf+OzewpCLTxmh22477gzTlzyAKzf9HPC2xSZEXiUVuNECTIdK06+8isUIrEQG
WDRoN5qzal2gdF7O8JAXXudcW7QxjAz/5kRKxYQSqO+WeGBVgOXuzJ7dUA/PRIthjpLxYsKrlKLx
L1tnM4w0g92gd+CNgZfIgKHUsJMIvX9C5he6O1GnUFUwrXW9i/YvgEQKcq/5hIP6ExFb6H7fRAQN
TyC1geE/OvqAWril5XFqALh9pAW9BN6s7lrgf/Hj9aOV1rxP4y3VcFIvM81L9sHsj19EGFAelf2y
KFbDrfTDUtytVHfuRD99QH3VyX/bgWBknhjUmDDKjesTQwtdV+ymLJMRC0thvt4AeITatt7R7kQi
DScvUs/5GfeTVE+GFiR9sJFnRWovFWzk8OuI3lnGl7E2qDj/lp+EyvGaPksdHLl9jkhD7/G5fK+l
io88Zi7GdyZq437DhTLgua28K401oaKtOPZ3JpXW2rt8DDJ9hLOKiPkNnhhEWNsYEay2OhmbOie7
NTaVdr0Nsn/OdBjDJgh9yCTl8POOxwcTX1LPQBljHa37/Lx61X42La2+OHdNP2S+8M3uqYzLGkbT
iBjcjZt23yzaWmsY6FNa89TVYzax/4oNHn+oR6TfBNdPyaYjPZW/h9ddhRzXcVX/kXuzhu9XWiV0
UhFJw6fCevEmSsMF0XG0QL3kKl7qV0pT5k3qHQMx7bQHSDojtd4ZYy/dR4pe0nK9gfB5iL0J2vyI
24CtC+Zpg/tARaSHDQTjyrlJEIgiHkMNEQwyU7ntHzJTxZrHl5RwoHLQq+wmBi0SOYzoc30jtaP8
svdzMqJS+KYQakdvHIvOGQjppUzZJ2Fz9wxV/aRxnNt3AKBgf7bPx0kaTXi1nCV7zfGoVCMK8kBO
g0dwnNElNWJEK/2VyCyPDld9xA4JCyWCEnvmxZLVNZ6fgF0vH44u60lsxGsTJbs/lbz4KbPDMCm7
x8DhtrNZkf+7WljO7HbOWAYBv448rfV1I3bDugBK+tunDdlaxzFOUvoHrAixroq0R9lJ6pSIuqbF
XgJhHOB3kmRPwVvB5xedWZQj1ABjiIG0OO7RLIjFThgb8Vg/LPjzNcAFYWPTkfzqBobP2EEhwG9W
fP6Wf9diVliq6ROxngxpbWZ1yv+3phbJ4a2pzAPeXXJlPooGLUIqAcZk/P1KKdk3TW5UXVxU2NNt
MN69LSk+NXTAiTcpNdBhV7CnHckamnF7nPXT16zz/JuAI2DgeW9f+7yVW3d8J2rT+grSXSOAXQfO
9J8DL7oeFHk8+D7P1dew0Ri8YLT6WbKMUsrfXYGqDMwYNgD4zuC4Phmpf3ROIl+QB0i/URkhZjcI
JPKCCqUzi1Io5iS7lErRnX8mck2BRqcsRdO6VgVSJQI7URg0ktkF9j3fdQ0fskNqzdcncQkTAslN
nc/ynQ69sbmHom8+vQkyviiWul9sX3TvvB4PkFgDlbG3adBqKF0i4eESwoXs9pOCbmfrj5Xo/N7Z
q/Pwu1NhclTBC3qjbtFv010ao3Ku5oZJgfK5XfTo1QwLPms/9jFse5Pbffb3KshidM1fsIBCS+SH
Uy64PM8qY5rGqVHhSGQ4RUELxwARKlI+AkAmrj30o3Il9jomICH7G2onDPmH0lCZnvV0EN6RG4EM
gtfaGG/+OGXpwreQKqSe4AYYkU1R9h+aAMzK6at+/WJN2WI9jBzYRkPNMxfRIst3fR1E4xaWIwWR
6tTC9hnm9PkRAozAA1jlsjSJ2J/l/rd8GlxQpPMgAN7Z+BCPIYKBADOCxwvEPerVZRVGoQgxEsuR
tr6VVhYJ7E9hKnD29l9F5Zdwt0XYAxqxPFeI0ao/L7PQfR44Dn+HMovZLcEJMio1FYrlMqTHHHBw
ENYAJn0NUhBYuxv9gEzlzIezL0zHhsHleNfg6ZBJ1CU/nCpjOFieLC5a/Y8Gtl7X41ZPjdOhrHQ5
2hNkq8jmPYTzUxz17+moj843KwtePOeOBkXM+Cs6nnhwnBM/LwoKbTIz5iArd9Fc1XJrJTCeXHlD
nyRByftxez7GEysPPDqDcE2yjCIzgsA1aXO+uFD1F1bmTlVx2uUSUSTGBVaY+sWVFq6zL04sTLqj
lP2QZANnTZ0fV7JkF/WCaJ1ko5M1Vs++wEcD0kKwQHNz/OtxY0yl/jvzprfz2wvvsXQkiP7kgmu+
FQFQq8S3m3NBug5zMNr2yjiIR8mNAFQSOUJu9/3TNmhg16Ey5y5XZoxN8zXaWBI8lyv6WMGexqP4
k6InNESy8e0BtNTFbXucqznM83vxlgGrT8CUp7ei6gY/Z5PObBnfLd8ESMcrYGaVIRXqxA+VlxkM
RQLOYjZ8o3XR0u0e25hHE4YnxSLwAPt7L+25GU3T/whOvdpWYyVsDtLvUFfqSiSkKc7UZCLrEEWm
aepm+hfEHOYXS9iM2fCVR7x+3HnqBEd1O5TSY3RSKgRtZJdPRTeNAKtagI8B+rUf8rr/9R7SP4dE
39Hb7VeusKz3w/U299MZKNhzOenceJtNQmoY5Dp6kqsCHSWqqdYjg9+R36Sn20me4L/wt3mOoX4i
Sx1CJ3vTvH6y/bCQ64c2LUEcIkCt4nKjT6FBmofDOGq02DS/Wc3wWdXG9jFdhKJa+hNWF1trL9+e
PQC7VmeliObf3a+RxGwBeHqpe1rmFcZIyacyy2LaCIEzoJVRjEMTjMEVde4dVh6YWUgYW62Hev+F
YhqanGQxesF2fWUhrtwMXRz3fVbcgfHgyyV3H/6blJagkCRXTXZ0zMGOQQxLnmF6bhHQfVuNXdVH
hqYk69BiZ1L1vGGUIFykFUIUAfFLxtBuztGgnlHiC9aDm21L0BDWtSNbxnwZ59nYu/a5F/JlCbLc
pxnpSrBFNh3RQUS34MjJW6czexjyxJp6YYO6RjfZC5NQybp+vh7wdonvxcedW85xpFSMPmTYQTzc
1CkrwiJ+aCc+StgVCKR+3U/2AOhzAo8zkR8uTH0Qat7hs5UEoMZbKEiSRWpboKayn7FhXqdVmUCt
gPXS9wCBvA5jeuiz70d1sOatn06mc1EZYLaugObG8r8XlY+T+GKEbP/+C9TrwqvYeaX+HX2o8ask
SSDBolI5m51elRVXlydYManwLy2EifgGoY347fDj754UI3o9S3zp5+BQIy0bHAcs4mHwgutpVObr
BecQiys6lngjzgONLexKkh9NxpsmYJkkvM6EMp2JQQ5ggRC93d8Jt8OrlK6+AGaTTW/O83zgTlyR
mSkzzOM8pUtIpsoiyS2BSAGNLH5B5UOlzAPFC0evaEww16Np05MbdKmmuGgRbKXy06CpyCLx7SwI
FqO/VAqIv4/3HRQ1u6EpWXjetGh1pdR//+XdUD2jPLHg03pSF9yWKLrpPlp2Sr2+5Rrlx4NFrgVQ
MtCkBUfN22PRoVYXUoraSWkhjElLitzrha2P8QMjGUGu7Sey/UAy0H4hb0zV0POPNa1/iC0E8dCV
gFSW23d0r9egcl9PaRL30RAY8fziD1KCHn3nCTckgWuOOIABEVaMGBwb4PS/1WQIpQFBfjCSiaQ3
iY/4zoT9RgkU1nKUSzFYhoJiq6ULixIdzGa0x0Rm2Ag/9EE3DLQsFpYwPExDpvB2+emaxW382vzl
GFOewHf5TrWhGHgbIBuCj94sUXVv95xdJ9gy+fOEtrZQbKGWSbMo781zwOESt6gipE2FXqjoiyjQ
fjQzTrxhW4HX2OTAiKvsyNCBOrJbTXBN7zM5eS/m862BqILKE0KyYE7TOSWglSxTJPSlcF+tbgxi
WXDmIPyMWtxTuh0Kue8H8mcKneIIEECFbK1JyxUKfh1+BsTXoWlJt5DhoLARhcQvR/CjUoQKR4lv
nx/sh1LpDoRmvxw2hOFLDXfKL9qLt4C6gyNuyrH3RP2+tOJIyRSt90RJD4n6+7mhYL7oEDDstlgu
r5yknYVAPDOvzvii6fBNCjddBwLT6AslxYAgslo61COcAz5Fm+JP9AHMPrD3q2ISmcvF+ioK+BJS
aazvNjMDzzmr5rhtNjP26VzAFUMwVC165tR6GZe5h/zBCxJL1HNz01rmNg/oZcn2awKyS8Jm2/cs
1aDKIk1ZsKAyhby6rG+Im+FvUDF4XEN79X+rrHYdduudJbFZ5yyejg8qJpoUAyXxETOSLYZKXxyN
k23cvecBKokCQ3wwQMt1gpdYKakJh8D6SN6CRmbVdDkYRHGDCum/8tjpcHiekGHOc7pFZ5DOMMel
oFyixlSC0U2pI1IEjtS6J2lurLdvxP/Q6cU6O9OCcYu2VS1M/9zPoI/grnj0YXDyZUtuyIofkUie
GpNixHzJUw9SW9m7wjY9kWBsBt1Zi7QYQdpA/xP6JVKtvwJOIamZ9R3e2+neUxUxUjjo5+g8ckgs
q48ORMEfB/HE3GiPbm8Klkyk0GzwiE/bg5klOy0s+3K/6yA/UNSZ1bT93fpvugjAL3SHuc9vAAXT
YjasjdkTAukIQXjaTUOJUuYRKAKoJovhHGB9rE5fmSc+6GhIYXrepuc0US5dyplPe9hKkZEX5ios
O6kaxSBU3WHcL2Opwz5QCCN1oI3vR3Pwc0VXTS992OIh5T7v694BBabT8wPmp6pSmZLYvDtAk+pH
jO4LToSLZg41srR4RwGQOHRhDd2DK9t0ScjEO6F+tKGjd5PHznNhvmA0rO0mFeFzdtYWFzbBESvZ
W+cNKpUvobITdyWyyHpeLghuoZHxG6Bxdp6DmUoJy3zMb7qsCwmjFZ9aBmtHOb7WjKzNPv3NrRAC
6DRLmFrMDixTHdqM22vUZMUtnDdwC9fji2+fSJshEajz7wO9K7vz7UWPaQw5p7dTC3AV0iOMfjxn
tbKcBtYQlWXWwC11mx0Nj8fnmnu+GCXm+GchTcCDR154wuOzzg0T9s7D7nC6AkGNNsbTBE3tTSOH
h5pS2bKSFUL99vgOkubGBEnPiJS7c3uPYgiTDDHHze389oiechGJEHDmFyhVylcWZosW5Qjinv3u
Y5fMXFSMuZwnux2GDbWCpfmC7x3QK6rynHudR/ARgoVNSJRdJBjgt9Bt3JnMHa2Jd8FBhwufR6xN
RTRmKzyabGoLhjj53iqUqdrbr2m24Ltw0fLGyKsu413xI0TCotuCZtfRXFONqIeaRDoPZ7rjoSN6
jckKOYjXrzbme9x9sl1l14iSLOzKMWPKz79IR5ob4gXdBXhKi7ZqjU7MTeOl1Iw7q/zlxhx2LYa7
gH+saR5Elh7GJnzbJhDFJFViliqP4KOBschrU2d7MVuYynv66IXH2xD4VT2R462Mx3MAZ8wrhGNf
lVc2+HI7ehTb/XXKr3EH1gk05z0YsKo3XZFvT/cVN9/VndBZAETcV1OhYkzcS04A/LZSdGYpPYuN
bZ1TQsxa45EMDsNPv16pGjF/rNo1qQYtB0599SpBtJSds1DsFHILUcfYpxEVPCIjXVCs11PyjYS9
L8d+v76hGPYzH7IgL+qymfU67/BMRLLUFVVKe9gqL7FWOv5QHJn1L1yM+Pd3SARaw3daPLECs0JX
2KTRLxmCWBTDDoeCfZ5Qi+BmfFtKiub6QnnR+HK6Zdkrd3mJwywZRzwGDjUp/53ZNdyVdNP26HRu
BBrt3NRt7d0lJ5aiq3lPDSLQK7FLLU9/F+drUD+7O4qq747T9AODHrJX+9dfc6ds4y5829FijNR6
yxi5okG9PaQXXBFv1brOP9mnFADCV4Rrlal+K0qt4KLwq12jaPuKMy9k6/G6aBa7abuQpEUNHjXW
94obvDsFBvpTbz2SvxQA/i1Q6SUFtg9i3cwP0mZgdNtZ9nVqpN+09Ja69dbzSwb4Rt6kKpfL/dHQ
TzRnrNe9HImNpom4/9XKSco6yLZyK/9P9A9jBYCwQljt15UFIX3HON6KyWr31ddcKrucc8tQBx9s
YxnxCdHSCyWMHR4iNDY0gSDRjpU+svFRAuUGY/xrbWUDOLRj89I0jkdHJkZrVRiUd8CYWAXlnCLs
oJohu7NnKd1PodT04doVhWYCcbt1pFjbtpUdY+dcmW0zo06s2uz/65GQmz6RWxjbNwte4+6pharD
8KIwS8wJjpIVx+I/kQFi122N2028kKq4SJWH4K6wK6UPZ+XIfrqOrR9MbEGQdUz57fpK7gsDC/Id
AbzRpaueGEkw4kohEyfqW2S/cCqoHqH9oBaYnX4Evi7rJEibKtGXVw/u1U0O+DkqdFH4xYcKVS3a
m3SH/swdjsJnLvhGk6mmtA6kjRYzKc2PaKCUkNvqY9MxtuHMRq+Kz+KIrxlhl+eWtI7Xx/n86fSK
bZ6gI8E9M82vVxsdTPdKy100kCTUzEwa1PQYaBhfX2NZsutMCIrMxsJghPhgDKjNGVW2ZPm5cCm6
mNnEI/pk2udgEUfs+kaGs3IJW9fBV/3gAjb+qxujfvXafj2T/1qI8IPaDOSHTvkG1AM5b1K+K9I7
EONVQXRFbCy9kFqx10xNYO6bMDSn7BxatjfJzETFcvt/zImOx1873N4AuJsA+kIdBerI8Xpc4QU0
d6ljmsrhFWopOlwy1J3HsL/lMKogNwgbYyPFK8iL2WogZtJAoL6ls5q9lVI82dwXBvwt0VD4v/Nm
t3xIxWBh2cw/8BciPONV0+ftg3cPEci0RyIm0EKXnruY9FMJHmISoX5ft/ErAxdf83hnzZVDAh7L
UQd/MjSOeVbYr6scZqVJNhE4spu4rIchpEXwvJSeJp1qxf90TcVBltOjWOqfIg78dIxG6pf/IJKc
qnhO546isDXQwPJxGBmvdlote4XOXm27qahuoe6Zo9YSpoh6zIzRnceoiOYwky5xM7yK2HP3+X0r
9k4m5Oyfad2m1EQF7lBUM/7yoH9vUXo38YwmYBtWUQnU0UlyFvmcxvt04VDFAH9sSiEUR33zGYnC
UlvHlaNZ7LWr8DovW+2KyQe1HApyg7tFj2HEXi4nDGNzXvo6ADZYI7mOJ8B+WYxTa3Lqu6mO81BS
be1i1+GTD+4pBkCRyFG+XyzLDWH0Rt7poKVLyPr92qWLRodsYqG8u3romgry69aFLKUzL/LxA+/W
I+ZzEYQcC74fdwF2o8Kz9FswRWKqLCtWkALC8TyVVnI4thBHwtYRW/JPAvbMvQqYEalV+VoOwXM0
pCeLK+e/PaMV4IzXgah2Bo6IpAw9iNKXpV/6WGKP/mEmlbKntxHl0u82NCTYfX7o3cORRYlnFC6s
98iPtQhdbsA7y1vM/9qD2ozUdX1Xatw0vSLjaCUhxnY2TJNeYF9YCUF76BxzKSFnVQDIG0fWTHkY
FefKlYcjtJC8gmksSDX46lsVi0DFWPphAP6zaXfysr6wGLsMTOPbBue0iNpq2F713lZYsOPXIxLX
Jm9EJ+k4aJZr7OLOk8UCtStytmlQwmNpGONsG3F/VF9wJ6CDb8ohdVXAijfxc6hFDiljQXFrC+qQ
0v2o88SvbBxa5IG6udaKLDau9bCUeIqmBaF+XTiTRqIvj05Gx12nYZKFgf19KuIJKuYKurtkQPrL
am5TEgw1BvawEaKSo9PKv58K82ut5xCWiPZiQuxcXDjV6vqO4LNIjJbbPseuVL9Awf7ZMp6YqFy9
Fv9nwClMmNpgev4a4ZjOSvdxAZdSaiNq+LFYM5p56f6wUBgYWhwv0J6dm1/eLvw5mNVIV+ocoea7
kNQzVHfo5er1ltUR6z2OS5LbvBfaOQvMQXzYMWghDQQaCHdzjE+cVApGjPKY5SsyruUiyq6ZsnHW
XpxoJLbPchgvmxuwgkO+7SWPtjLanFDHr0B19uCDJDFlxOnFFo16kMXM/k8iOjcjMoqptnrhft1D
6Q1R1y5q5bg8rguaQid0fdxcLEIXW5lzeYHESRUG1cNlCBkhL6AVRrgtN/fjK2lUR++/LVRPd2gC
b4v360OZVeos4nuNI46aFLyVqFXjcwbrFKlS1BYbETYBMSpM8t3by7rm+4oQUHIA0psm94Qc5trs
XdzbyjqwUqZjt00xY6nPNIQSL49F36JpYyYtWeguD0BobkgysebWKqYnVTfLNC5XVXyHlOxcwanB
FiUmDWU5kG6yLQ+eCd/1n6awCQr09c/zGVUcJarxwI9l+rscTGOzW5HfXB7ReZqcd4jYq8RYnxMA
lmJ4jJWUm/TvkzN3YlxmiA9U80SdBWYGCrR9hsMW3b8HDcIgONqhpf7iZjNcc80uf+duDVwfKSG/
VdbmSi3usDC/fcgooo2OFWM2bPMpvCFWUug/nqn5xTpRfFCWb5VSdeARQBFjczQKzRY7W9eHuMJh
QZTf1JLIlPYW22hS3ThgzBZvkCUevgiQwyCYvGYO1ugD/vGTrhq97QZ7VWY9625MBbXsxi+XRTC0
fiCIEkS9kc4AA9D5hx7jj7vlv16wUdAjRWcYQF1vAhBWNjsbvqDRleYNJWRhz8ENpQKc0bDIcRIj
UGVOLNY2F5vMxESdjB2XwvE3xJa7GQFYVIjcwKsefZVpx+hFMVfqIiN5/9fwS3wIolVH1nSbLcaM
0LwOwjC0KDHi8mnH4INv+rpt1TmlSpbmvefrZ+5gp90Uix8MYqG1PyLDMV4Bo+scqMkQGYbAsbM4
3NERVJjW1rHxNFSp61808yVKOHNCMNhRKMM1Buhl/bqX3j80Zral4IQHzrpT9wdepRb/5NV3CvTB
LNk4A45GxuX0JU71IAr1vYbtOk+qYrMCwiZslBbGIW1UPDQmBFxEPQ+McWTHGQoHtw09a12nzkGb
8VTUE97CgVN8iBjd0yZAjef8BczfKUDI+VNukVoBvVnth07Nfn0Cujw7K/Z1VLhPmaoLiUYldAHp
tXPhfIiPGDijmskvtGeAW6TomezYD0tDvQHdMaBcDdQxYoovTcQPv/pxXNLmS5PdX35bb4zQ4bJg
KnYEzBXC9Va3fKlSBp2pR+wcUfOQ83abRKuGNFdT28QZc7b8WRm3jBNpLrzc+zslGmnpDb5j1Zpu
JpaKAOqGpFhtp7t0qoDrWOAflsU1yvSVO31adFKO28r4fEQTkJvqARjXltpC20dOO/He4YSAavBR
+EpFrLrk/k8E4Tt0PuMDbVBwVi3PlV2ZS8kq+RayPcbRBQp6ZR64qhv2BqP16x0DAwBNv++DO6h9
/+/aovxVb/d/FMwvKnWjUkm3Vg0EMljXPqyo8o5Y5KR1T14KBXwrsPMMgN6mBrhpugTeymIpkuGs
q/qGYdHzZV/mCthRbL5CURZgRuvhiANbYaCcp5S1LraF7b5OqbzkBhJWnt1ZPFs+zjdTujg9OA/n
wF83YI5Wcw2ERBr2ljM0i3me6WIgvkghqsZk0AcU1Xj0p9t7LzCp+fwxIZ69rft5GutLYqWZoOM1
EuPv+Suql/8puUq/dkAZLrkYTsbUkv9Znr29+dbT+p+KzBRwq0dBXgOUdwMGC2G45XWNxrNa4Ikg
tgAlJoez52ws9t4Hqzq9mIPgkrtqkQL1iZkt76LzZ7VQIo4jLQ7CdHPuE+If/l0eI3O8a3PmxY6I
aOflZ8Mp33G27hMpbcvWYlak3PfeW3M6JU9Tb5RxUXM24BtBxMu3j99JPaujZa9lhqKzIc+rdalj
49Ifksa2UmDdrpxX0ZSUnTT+4kbiR9T4cFGy4g8ZlRCSXxvsQxQF9b5ESQ4+XzkGZOk2hFzpMicL
t9SkI+CJKmWEBaAa8N5q/Y9CH2jIS2+Qc2PXREKQbIhu826nipTUP4/FjYaJ9mFN2rdeszzJ9MSz
hxwmNpmq2nbOKqEOEG+Ko00NtipvJEbmnAgZLE0ZhZx0XsQ1wxLyez+TZFrHMmaWZG9IVaB/tNMZ
FT2NJkHBFduguRQbXoIx1hyyyydyHtkbl6LXrYRzV3l40IQ9qwjoPh/MjbYI3/hcbce07URsH5Is
O3cH4S21Lx7aba9JtuFaCfiXYAlE//bZz6qrzMosTQDPpSguhEXQftsjqGjF0Ec96oUIyIKpy9jv
yx6YTU+PIy/1Nhb3DZpiBP3PzYQYXeMQGxFqBfObH1kaW+ecAL8+wGnVApjRxn5cCjcyLRUsr6Kp
WmdbDtKGyBPkbyFI3JIs5JShLa7rG+xNACqJmIxQn9l3T0YVw6AAAkBWaSQF8w9JurIcAsMi3tM0
lYoBI7as57I9f6BtSFeb8fAoG/w+aucFKpPk5fK2B5f9lA/maKxCE0qty5XnnOOhxTPCKg+JAEQJ
4hG0p1FXYJXxjJsHlKZwThvTJrsFa0tn9n2TR98FJsakUW9EVuiBkGDJ8nJBLB2Yi2CBIHcPXptq
lKCbNqlmcfFao1f+VKospEiS7AoR+1ruPCIS4CROil8ptrvV79POypWM91MisjQ07zKNQGft5WVc
v+kqPF1Ws9xc/Q8RFSZ077On0d8pUuWr7e/f/JOsqAPlam4pL9sxZ/umZLk39EoNrtJPG8HT0Xgm
1r2m86YsCZY+3JBEck6gduHCZy7vJYEIL2hymejy5kHZkmXRy6rrnFz990IuZkgN2LE6COW8g1do
sXnuv5QBrQNalJejkeSM+oXxa8F2vkDjl9oHh1DDwa6XccJcsebWMXE+ZkhnpH2aNS1i64Hy1u+B
eb9f1/tL/5De0dphw8vLd3HDFyR+MeSXAx6dYl4ZNCKHdJlxxqM6ZGLAGWNgP8gQkVCUVWSPooXl
ldNRHPbehaUiPrvWnJWMWCObyLKRC4YprsHqlvcaUyPGZIkmq6KhKKTWxCtPeOYSwnt6M8hCr5Gc
2EPjrUdL/98o7o+VD7VbWTsNmKzjKeGs9yEK8FzTdkbf6u8objmhyTNA65V9Y9v0fHH0k8XmU78w
yoKysaD7/tOr9imV/mpSFrLmsopnchezQYYEHGPWW1unP4TkvJOnwUL1BL7Z+wUc9rYbbnVhOEbx
8KgiDLVmSA+TX5kZTSNwAeqLdw33wIIdSHBXGB2poL52li1OQl1WNB/eYP/W6adkCe53YjKAC6g0
9d034cccs9XPq8EMNHXyo5QSijprrYEgCV951CUucDBhfrhsGyqtlKJ4VTBm/qBTov4tMtpTAHJ0
2XmSrbGK8qcdjGB+nZ9qiv9IhQdvcO8PQcAfYbF4Ru8QrMmpvZVvvVcQTnzE7eK4icdY+hlQzFTP
JTNt7pSYFKPI9uOildg8RpdKNIGwcsnxMG5C8edjXPNTv2R+qC/bC7YFQ9TJJcECPrn7ygnLTrpK
FYvd9Pb+l+TJ7wd74fyxKvpG3Y42ewrwrCT77SKjFmlDIf0EK/13TYIVBg2B9FStRN6/k59FzeAq
kMJH3NuRcoHjGssQsyZD5xwBff3M+V0skVQByxi2U5VHBs8tXtzzWDMZzMrdMs7AIlZ3UJpAdfNR
ejmfKxJpRqbBr1h6INeHofcIe9AtJnzHAGQtB+DjGFziYpyFCEb3JOGDvvYUWEw8o5epv4+nsTZE
0SVFlRKrm9zpOW+brFl4CwUJEIetU38Pw3VeOcfrbVyYV2vQnr/WyeKkwGA4DTHCHwzXD1nEzmLc
zySNCP5KoCMu7qKJ2vdh3H/6DkD+RpHJjnR4Ghkx9EusK5yzCSQlt7jO1u8y1R/Ho5FJUxOqpD5Y
z/fBt8+xORYBPRAl/YuogUIuJM4NbzVj7eCyi3/TKffo9yVkMVBXUSttcaXAJuP6xlafoyBsjJYs
PX9zHhjEbgvXHmv5RETd3X6oTg0O8hsv0zQfmgwMr1yzFOkgaglbenWjMN9/Tcfy+uV06xynbCWs
WkiEuPvUQEF7XCA1LigYuQstDbYcr5XvXkwGG1b6gITvsiCNoEf704EeDZoWsuiTWFRFBoQ5nyBP
Y4DbJfhJwywHAQGoRuP7l3rsqCr9LZtL7Ws5/MfmZGp/CfqxnsZBivPuORqWImSB0dYkI/UqCd9i
KmCFpV1C0+JJ06lu9t/8m/umKi8ptAjuZ4uOfWUC7s9UuRJ+eEKL22ZhqcTeaiyj5VfLUeG0EYeC
hT7FxBa2M0NrcaEhDi4+4Ic8lMHRVGIZTGORQ+NEd/Ndg8S8y+vwLZBeZnOnOZ1IVa12roi50kGL
Z0voHUsetORV6XPCEBtSxvhg8EhbeY/FSouNZf+PgI+9m0cARrKRO1b12LXeCtaZU8Spu0sqMO3R
RPbL3PnaIY//qyMff4iqZYgL6TfR5fYHD/KBsLJbNLfIuEeX9JLl9VdiIIn7DZ8WQpccZWvyaQfp
K26yLf3YT01WcpOmqPZkMAYXnWQN6rRkL38yFIzzTBuY84Xhp65H79heLQYlqu5F9Ie5dEnYw+39
rbjoLvY2e9N3eETpyi8FhtzYnZbkDmRXvxkBjxSB5yHzjuPMyAhv7XDPKu28lTNSxwLTjvCMPglo
P/2YCiWfpAXDV+F4BgbK3twsJe1GgltFS93m/8qJ5l95ybbbaOJauSo0CYUJlgHK2Y5VUaoxgJZb
UpUqswYuPShIeFerTszKL5HpQKqFlmMUn3KrWLARiP8OGoY1VumjPTTqZlfLRY3usFCJYOKjtNBM
zp6GbrBLy07CgvEMzruBEDJ+yrr51w7PZ1rF7TAX9TFK1z/3F0Wm2ZpsbzbcFvN/iSvvI+eOxdxl
baFkiOWQP0a4OYrlHm9yPl4Hqccbu0KhUyBfUWx75PsoZQ06UvrHlhp1I8ERFpdYilUEIRdUjKz3
wZOcDFB8/dTEPNaXET20H219qXREmTtk8Lm70Mq8IArhTgWDI2lMvukK6phAiJX/ogH6c0tpRmXl
Zqt6LSb27SMkIvcJVh6fCdF7BW3yHtqw7Z8c/7PkwgjxacNwM8AMgICDN4WS85sLPWgR140uBqOw
eVw+duo8SK3y+W999gdanBNjUHY9H2HrglSmuyvpPDuQuT/Q5tB9hNP2vBsVriAGeSkW/U3LNHbx
zRa240OE9/yaTPfFYjb57cYiO2H7T/mlVdJFpjaKSbb8hBp20poM5ZTnD70YhTzZDs7qgZlVD4bP
S3EHpIGLawK8CyKoSKGR58PTiwooCuHNQj6YNXFcfTV6ab1mviwUT3XTiwzI1mXZ57CX0zloV9lH
ACHLWOM5LvbpYRi/SLCOBHh4laJLL2HdpcP0Bb6kT7NpH5EyDfBEoK+CJb+8CHbuqD3xc+4BKHsp
Qt0RCEKSO6opWZLy1lXElWFp320u9R+HMrnXaXx5eRo5NdLzvoBBwaC56vSGFALx+c5080lS5kID
petf5iK/xqqDqIVXgmICQeW1KplcU2JA9oCFiDM6lMQWi2F/S/1aCqTygddhBPjfOe1mWSx+eGvr
vwPaVs8Yf9rXQRkz3ALgHdIRkr3WV1IaAiSyg876IevP+3yAfZ2V2md95/9zA4/WK25Dek4hJbMp
cv/w5ius5UeKOwHYWKxUm6dPYi63hXWvEUBhHb5xFrF9ZT05tXARO2bSCSbgVgbGjiBawdMXvcOc
6Jt3PulPIy26/2fLvtA/04a2CN7lez/w0KYZgcwHomJS1jwSy6ALZRLhpRYEoxk2lxgerrq4H2E7
yzt5YMqIANJt7SVrrxFCEJ/XT0Zd1k6oCTjfFwvyO980TQQuciqvJuDDavMXZSNH2GXUSW2P5Ry/
cUgFaeCmdMqanKyeG/t5q5LTPXbM1JahfxNvD4QQDpl+C+v82W+6hVfxkp8tI6EDu9L3pJT38itV
xZWGxoX5RV001kjAJNtG/FfXRrhQ89PpY784I7vU5k+6PeePZqqhaFOfNmzqJuCOy9d/0ns0f021
j4tp2NGgQXDyjsrZAdTkag7Q96PyYPvuK0r1sOf4u30u53rRKRbz76AyO/IO7Dhz62yggEUolWjG
G9+RFQrb2QH6CHV6UcvR9u+vhkuPZuxxV04Y+QvG7fbK64ndK96W9BzNq2yuCWF8ieZQbhLuCUwv
vYa8lgEu9S1tStr4tvWdIui8wktlic94zXponAErD9+K9JpB/e12wmbOhgagiwqda90MPtnNE4E5
qklFF5q/yDzmdGWnchJuLTYR92n/4l/0Qn2ErZwPGCexjuDSF9Z4qmTmQqDnO0+k4g4nMsMGfJjY
fuAaBKVGk73BZBKbl2hNhtgNBHBN5SRWt6qkpX6bL4YZHJmcre0NDPl0JY4ZQUiOqMVIl2vaFsbl
EDfUe2Ir2fzU8CkycE/d+l3WiAzbDw53ZYbAvHGWSToRRX2G3HFgfxwH8OuBD/bUJlp4Rp230qn0
Suy3sKMgaCnm+hPNUGzqhCB22Rcp+BYtKYWLQ2vLKdlIcpMuAwmUGgYuBUDFZmms+G/J16JNxokt
qaFT76uTk6f8c+rucJJ0rcI0BwM/r7hI/9sOuy0fIaKyXrokyCYHszZm7SJy2Ikc/E1UbUXuXq2k
7Dpz01GJNDFHgh2JWpSEyEIhXO3fZcqZpss9vhZqjBP/HwFyk9KqYgLI6NNCIyEQBkA63aZ2zSCk
s6NO70LzQpbIQw6qH0gZwt/k0zYf6/OvRnIl3GCT8iy+4HF1gwRdgxhVh9R/ymS0jx8gpBfkhOrJ
7YGfMaKpqEhbthXp2oZozZqeldBmTu2+rzxhO4qinNYXQMPj4tlN/RKEuFlzPmizSVx9m/4gsKg/
RgtXZSBy5RVPX4FQOm2FRsTnmUZRMh61bKZ5Alo8Donoh5nAs3nV1x8hUrD1Si6jALzM5uznOM0r
uJbtS0FaQ3cLbGNh4PSOSloD5H29cQsuT7wF/ebgiKQEm66CopMdhmYLNDOh4nu74YL9PIrK9NXD
LqE0rFvrfLsG7GN7o87OzK3wc7B1B9niTIFJon8qEjCaGVwdvmcuav/nnurpRz/CKxq+EZLWc9Ki
a2RNRM4fMdwgCOOsKBjgDZtKQhrSa29XaRL9DgUMQaXJdz2XeorW2tXad07XXmHw2btSsmhJDRk3
Ak6rn10YuDysgZhgdqXzbZmvf94RY1CBSf5WbWoPmbBu4D4RK/wE0wKmqma83mxBkeFCb3G3AktF
iwMPXsHFbaJnN3Z4lhYBnQ1+be4K5pjzzy/v8yczuqAlV7k5r4LI9Xz5yc6AEiPvPFDTPhe1dcA8
M/+IIknKUOrXO5qpWjVlpijzwD/FVDZ5UD08lo7puZlwbelX4Ms5c9JFlmfI5P4biFyT1wHPPQPN
uVL0sF9C33LqJZT7emuIGeLJEsszkO3KldVb+sZGn7itm7xCBK/uBwiE68w6Wxfs0xmsTcILpraw
KPMbAMMTBN3FHvbjo0R8JsPm9RpA09X0yMPoSA6yiKF9hp9Fcvijg8GqbqpQhGwcwMYX1gvuhyC0
GVf6yZyrieK/QYJxYzXE9k3kZRBcqqnm0BZro0qvtT1JbKDwHI0HuT6xFWJmEXLWVJOhBV4zceWQ
aM5vF02PD2mcqIHegS7s1JGpQdsevccJhoGzVJR18tnFCX88A6eztg//HLvHNbMtiUs0OArKg6Yy
dFdKhgm2o43kRLFytQWR27zrd7T+pptjqLZdLsCs/6pwVCXLbkmsBww0A+G+f3OQ9fqP9ms979Lq
znCWSKZ++n0odtiu4LS6MBeo8Hp7H2CvNhD2HTqMol2hmQyl1D0HByZNAVT/kG7jrm7Vl2WmhFRf
oAADa1Nut1KXDj0b1UuqGCbrV58sNyjQg1tV2MJtgLEHOAE9Tf8o93QijyOBVIHKF+X5RaCAKvXo
yCGucVHtlEruBM4YdXFICSGbuDzA6xtmplDtL4Wt8V/VPsHwYDl46MY2fKc98k8PWoX7rNRgLm0C
cqu9XrC1xAUDXJiEYktUemn4anA/cBHiHOO/+WSLMat6naghswit1xXXMO/5yUPBt56L06s0ulZ1
ZbElfJw4uJYOLZYrLIMnZ02tNELkw7wwFekIYa9kjVJ/itfw2K6ABvdmzJlTjpmWP9WcGteu7MAU
3QBKR25Ft1TTED0/kAQvkpjiobUCd+zjyyUP7eNwNID73wnOBr+VJub4hhhwUY7ui7R6rUIMuE1g
vEr88eyRSNgDKg4qs9YJnFq13HCsgL+OIfFNpXtW7JVDjmJKkYQ5D9p9CS+frzWnVkEq1ftcPRAe
0TH0FgvFTHGba1g8pXywkYFhlpplHLwashLXuvkroQIUTcIZRTGTFadvjftm5NSzgn1OP2QqB/s1
feTH/ms+Bl7XUJUFmw2Sa2DsoIvMHc+s8u2RQ+6S5SqAYVvgCpUv8P9SEGI6qfDOfHuNxFWsNw2z
UGVEAkFWBKIDVqejLKpB0WC4ZR0Eimm6oh+M2VE3vbspOrSMko+aP/g9vB6meFS5TkjBEukDFqhE
xd8rDPvEwg2uzX/ywT8xJF0GGT5YIWAVqy10AlW/+pfQvWEELIx2kFdtGTf5G/WlksVj+XNLuDHf
Axnj/VeuPzgDFLoDiPFjEeZtvzs9+f2yub0SLOrlTh/18PV8y8VbiS4w0cEWJ0DPJHOLhsJbL7nc
2CyQZ+R6UT8LaD19v5Mm1RraXt6McNbXMIz4JZIRg59r4FqR0p8hHh4kMB1DlwLcI5/62TR/3qIC
Wp2AMQnGIeqeZ1+5Q0o8FiRKxUQWP0iyaM00TC6Uk7tFpzdlTy8FnYtg1ZD7vb9uxegKLhD3Qx5t
1/Ycfl0PFAHgW31IfioDkvexkWMBbMaRcFyDZVh/cr/2+sTnG/qECiKz1fqeELvbBhV0fp4W83T+
74b1Y9GsfA4vQ37cvK8P7EaHKxgla94/Sb9oXuqszmqXVWBKvObgX3R9iWhc9k1mvJV63jXjS7Ka
mCDpnq81YzhUyb0gfVza2/gOZEH75tf6PqTx0I/5apPvpEM5iJAcOQDBdDf5L4czuItqsBtE8e7R
9Z1pWBazZJafqCOHrHM3W/GTi6yR74rc4JmkK6N38R9CU/qvQl2id7bZe4D5yBF46qbx8vDw6H1B
yd5ueGusszBUgsr6Q5naKDhac9HwljG85uCbJzfutMs3QpoAUlcnCBcBY7ACgXQVvqE9qVhvryv0
QT5vmpjOFCAAeQxVWqfRlTvNMxpznoKXEfq3HYk9vCoKTe0iggKXo5Dyxpx9gOfutKehxsNPCks2
79Vgg3HPF3NISNLIKeLjkIkrrM0r1vtzPwUwoiPefm1Hme2OBO1fRBjUu2plw8rTzKZ3TjRmVY0y
dAPeVHesCTnxudxPbMkuDShFEDdRgBZ3H8SUHgvq5jxyzk8jABgKnUM1E/NZ2F06RghY41RI9vB4
h0/RL2t571FtXX4uFDmpL07XJeqtuDsjrBV+r76zyEGMiwGjBVAgzDtqSiRk0HPD5viVgIhNo7Gk
qMaIG50D4xLYSd5Lc+44vpb87vXG8Jz1NNJ1BCJjfRq5mYDrUa01sPUr2h+WFRcOOG4kJwprIemO
CxnSYxTxGgECWUHjYlw6xX1CSp3prQ15NIem/jD9Lr8K/Cv/50chMaliFqDWu+ihOl4lkwTt/GwI
a0r4Pdr9a5tcoZ/UWDSDucUcIzg73WVtzaa7p+S3ARlWck7DUqLWxFSyB1kZtZgQWVv/ZFfN2vX6
2qoWkCU6nKTAV3s7gJQn2qP3q8RJMkeYlDfyXcuH1EvRiKCzxVRulnUWGj87+DKLi5TwU18QMaxq
9ecSwu6R6Lldy1Co582+NMi50O+NY3ntZfI5Uf5wSenRsGjh65NBz9MQx9Oc2EIYIfxeaRDskmZr
Vg3iAfhWypfjrB80rj7w71DrtxOC/1ufzD8EtlHYHkZlOn9981iq3IGLneuz4ewtHmn/Gj6X630O
B38k9DI5fH8BxpasvJRucgwX/R+Nsq9M7hqyplr42QDVSrwg9DGUuLOc9l0nj60oUevBaTYSd9Ld
bkNdy+bUmvtP7pVpfS26DNC7s7dokrzmLA4+7wXJ6Ncv1QGHjVln5UOFk9hps1Xi/cr5i0rslmR3
cOElrj3iDkPR2aIoiGWCKqIcVSzsXgXfgyl+mrZs+n6Xs+0CAgMhMexvZnj7BuMbO+Xyox2jukyr
AkUEThubD3jdouZIM3ztnUatpMnRGXorkOD/oLtZwR74IdceIZrG++iilLd3/BjlqBtsOcUhSQ1J
vFBFnO+mr2HXHzEinHiud8atD9J3gUkjqz2vBJgC/gmiEApXyL9GHroUM3Ec9u2XBu213zVI//L8
HCa0Szm+5ASqVzaV5rHYuEiASyRhD2azA8g4WuUPf980b8I4qN9CNv7FCA633zpNzyNiSaxK/7Hk
A/tycwYGYFiuoWgi0HPVqUZX+6BW5eEh4eAvpWJLDdlAoLYfWlqHCsXitUchdRyAGmk0H8tHv2Cz
DiXmh9KTenPA02FcJToihGcLnD8+YJmJgGkX2jPha2I62+KLNMPx3NjO7KpEzmZoMJh4yHCI22I9
j7xQ3wWiet93Q4PSsPrODKnnoj3N4V6PIXIdGmIUdK1u82k2KmVZ/BiPZQbLeM8mCM9QvdegxtO5
sBulkYG8pJQDlW3zUHPH6az+YBkZZUi4JNabnpE6omMKKk6WBpTsTx+89dVEof1SDuNB50XLVvbg
r5OO4zKxao6HVOAA7q2mHzBhBDLs/wQPaLyTDxDgVsamCgclnBkmBqgBVo531Jm4KfctQQeNuGYt
gbr/PEPCYZC0x5nr/5a/gnAwRfaL0MQdrLlIoDwmUIrfGGssciM2QngU1xywsfq3W+niBndNOCoC
UjZ0ZUXp9Jyflh4QJ6FoEmSYYZ0KTvnf0g/7o2BThhEB7JGpHafid9OVs/5Z6V4AdNNgtUSxw1NM
hVBxgom+aH+oXKmrxkCIwclQF5On0Z74aumR/2nc5Bp0tj3pS/gGGHGWAktLuZL8Nf/xoNG3Qu0+
L+xc+So4HRAd6ma3xx3N2uoPRhsM558WPfHLsEk7FAwplU0dxkCys7kqAxC7LPmiQgU1G5f2FOgq
WjYObQALfwzGOB+IrQmXl62087Yn2IVTfhuGqNgTCVvX1Nf94z3g3joTGGonkwtRujQT9GzchQ4t
tPheK0xgqO6fd56XueN3JhQ8/ru5kKHOu7AfLrDGmUSzKBl8IsdP7oRsoRaUe+kMocBB95AoslCO
gm5nH8/t8y+yB+5MvbyMGam98cXZ4vAZOZ0EVfgOqPliezZc6KtcpOGrZUimHdveBw0MAdmJ3Whq
20bzDteCZXnHvycSxxu9i6D2UIjB6vQ7hctm/qcGxIJjNStmce4vU4efAnpi29vYBCS3tgoKbu7W
a3Tdx0XaiNHFToE5MhfPwjrDiPuFJY6X//EV3BDT+4m8VVtuFkXb8ifZZaqWurnbrKRVRLd1svDm
gl9vtE131S0JGnhOe1kKHGnCBnfBQj4LkIU89sPV7cs80D+A9HjUIsuZAyEcid6ilgU7Gcj3WCKP
IHVf8fXI0lAuFex/W0jEP0DAXDiHmKw0ggRYt5ajZwLCDXEmb9VGU8i4StXi04M2FUky7GD1nS6m
qTsDjy4wcRtbZDJwWwq0Nn7U9d27QAilUU52PELgDDBXddB3Vb0w20NMF2T9+3VSTWRH3xdXRmUM
HtkJCQRLCeI3T7mYeH58809gXJhEq1ltZ3SqPZRWaudSn/N35XO7Kyu4/FT3PMK5HMZf1naafY4t
i0If6/WDu/DZeW6djdFzGi3JR1wnxs2FAg24oxObrnbIrFutwF3JEdA7w2J8rZczvN2XnmZde6wU
U/G6+21HcnqQuqFRqwRPJCCszcPizpe5uvlgRwGqdH78+YfdFZn1JonY12FKWt82dUxLwMJScc4/
wncx2tT1ESq81U+iz9wVpF/kURiUAYu5rUIhRLyg1snmO8tG/rPx10lzSDbpVQa87nELovuisdOY
EC6/K5KXX6uRB7KQDpO0svfGS1ETNGZ0oLOccrnY9C82eoXIaO2slu3y1QnCCfZN6eHNnSzHpIai
8NYCQaeqwXSnTi0qKjGm+q18hHdNSNqwYjLHHFEI4S5pCDsfXnNx7YU0Xa6QKW5q+4i2MzGOq2Ri
y4HlRXcEI7Njg21pPBTuj9xngRBGtWbcmzIugNMqU3355IanOnwQ6DVgd+2Xg5rFFhLm9mHMGC4R
ukxWM3LhZdOuTLKAMOQn51H0N3VB2CgI1ZAa25B3z0/Y9KtnQ5YHrv5Nk1UQsITJHWvjW5drdeLz
Tn8tdtQzrpoO8ixSbV8EJick8Was+++kDaJ/F20mMTekSW+EBh62KbGtAfJ8p5xmuRecM2lUBiB7
muM535D4DXhwcC6XpqMjQO9IjB3Llw8K+KZgorYJ+GbYfWjtj+oTBSCzOawBQ5Uuhr+5+1DSKr9a
4XW2ndkyQoT76LvEAfaIOWAdhWxNQ22AJSGHg11XHEhZuWjWDDVVc+ZhU4aHVCPk2JtqjLdkLsfe
2jSUZrVWhL35+PJQTL5NCjrLG4iDpF+ZTPI4gJIH13g7Js6ANmU/rC5nzAcSygBBYW3p72EvvKeu
VAHRzUoPvINwi0E57IH5IY6wrgyYfuIq3EGFNFYr5cagE5uU3RTOe/Owjm7/+YynKt+jf41UJ4HQ
R09hSzDP5gtW1SaiLDFFrFxeQtqH9x6hmdQHrS8Odh9ElrjAuEmMl+O76DiubeTehnRbHJfVAwdP
cMJ6o5NDOqsf8ER0XP4i7jZKCycJd8/fbvRaBTZeseFcSkBctSBBE/LMPSV8+2f4TjimuXRn20g+
m1ZfYxSdb9coyga6qs3j+mDg9Ah8vvOLnkj6W53Ir9HXzRnP1uZLUVaKlIhgodHuu/vjyCIybBrH
qEhQnda3A3K4A3t7mSzUtNxR+gLE+KdRcGxquYhPMwUL4WwNBxcyrbzTJR1VquI2itkMXgrR51Mj
nKPXtGbiGDwqeaP4FJpvvUZq//agMayhmc5LktsCxWAOVfidtSMTRq5m33njnj1W87gNlTuC45+g
o6qTXC1J3Qz+ZfI2kWQk5Xu3Bcb14jXA0Pq3a3V+hlF7XF+Cwjh5lDqYOP/odMFF8e3XfCu25iny
yJbHBLKQzuWVdDr9QwXQ5kW3fS1Rd9Cs5rafA/LjajmKkzVBTfPW8DcZcaPcs1vtOUv/l8KrarJJ
aYC+ywYfzdmYZTdQlmlTt8W1MclXhnm00utf8gOsonPGD58AyUm8A77OAhe81I3akTAQ0e2U2ucH
s0Ll95gwFLWtd+hxjP0Fu/lGryPhf21KuvGMsqWalRPx9KLHv8zvbzz88WDAjliECY0CU91V1ACR
WyHsfi3pI5rkWdynv6HMriPlobO9C9JvmZqcbQ6aAOahdvW0keapDtBcLV3Sx41HD+L6UA7Cb14x
nt6w0yGXlU9BxUHE4IHI6XiBMQA5UFrQgPBJO8Ha5FbsFknDcDpiOoYnw5SRZT/Y8MOo6OobMIr5
iUGLiAvgu2OfZfL6knoG7NJ8RIq9uijf+VIguDEEx3Xme/yh1vyA2T86zBHsNwkSVFd7dzJOTnYf
Om+4BCSie1g/QWCzaYnJcg1jMUWQnR/tza+Wcy9IuZnwE4pF48PapCTeSNFqf+1mTTwn9E1sOB5d
p547adokJ6fiI7owESFKHYKfq914kcg4z3T1V7mDTRyt1cFQxgjIS5CjLWmc4FBg+E73gTVdtlZC
7jfsZMOjI1AkrkTbhJ3dL2pzf7hL0tPBSukz5xbfB5K+ETqRNb8B5ZBr1TSjn8B8BPI2QjOIq9xn
qgZ2ogQYQrIGZEv+IHn46Ne1ymeRN5ADrK3Hn84HT15ipqygGCb3OLUTpkvrBj9yOqczdTZln/Lf
h8xfPbS+GP/CW0saneqPoU32oo6nXhY/kotkkc5J8jQg7V4b/IjAHXzDKz86YF+M1jGPdZQkXhCw
OHLsoN771GSgqKvFf8aeh+VT8FLyjqdyTXMBn1jE+AR6HcJqulmBbnjE0dSQaaT0cviFk1+UnBRw
v8uFJh/rRf8LfbduEbe6P5zktrYgQ1y0ztKigOtT96ICjpUmoSsx5/cyMPvm9CHGzbjqM0SLdaHu
FqSOGW3cYA3mKDT5rLyntWeMjs0Ye9UK45L2BXxv/LLtxFo3/OeWATjttK4/DYaweDlzwpKHTQ9F
Jn3XMP93V9732hbs6d0vt5uGDzWos3YR4pe03aMf3LBHAeo96BySom4vcDbPPS06n1aHj+QQEVcV
l41JVffjkTFwJFtAD/TO/URiWywwf+2VaCUaMW++zIkgC8MPHfID/iuaUiId6Lrbb52RS/klujN2
yGLloe/QxurCnmyey7R+cJOt10F9UNLn+76I+qlSs14vRakUmc4wc/xw5o8r3t4tn18m27sJwsZC
ddH5Y0yuA0iC1QkqxslqUIDTpNcmlT7dIOjEXS4NsU6mT17MvwKShr96F/efnltWhivaZEpZ3OaL
0ZLttuNsI1iaA+M6sovQVQRZ/65qOUeQl6Ds3fCg+OwynpsQLjL2GqtNNzHIR88MZzLDn/LDHLIp
YQ9pFwx4MRVFmfYseMJOY+bygJdBRKXuz4WIFBf1u8V5ptq/EiuTwYM0bMwKrmLcSCbKdoxJ4qIo
GahhAdY1jWlfgnp5oUt1uAjqIDKKSkSr7nH1Cx+okcUtAC6GXA1yXue4PSrvExCD9wbaCEXl0ZYg
h/HPV8HObHjlJp4k3Jik+mD9j0N84cdnWHFr2CU0FTBkL2YdpjsYsxNmda4etGGpJ2KbAuv5yaIs
gMT3TYNvrRSjVCTEnA26qshdxUPW+nCy1EvZlu8Psv5VXbF6JIQ1P/xVzUiyooeMHWFeyBQ+DMbL
lUkmIvBpy4ubOMCb9aPUEoYWboLRFLTOpC3gLZCMnstI6P74mu0xcBiPkOBS1F+hSr/FaL5wQAmJ
s4JoNlSbFDBTXzqGviMLZbVPoEmLXqLglMNvM1BlKzgDoRpXIwRRjIA87RsQhPx96VI0SoFbE+w5
VVVXjI7hEk5kb4uaqoE4XqAhY8MC9uJN38FTN13//gXl/KGvZ2haed8rkncmIzQnYWHXfg2ICfA2
N2r1iOj+cTewidzqGpiBqQ2/Lfp41yTJBCu5RF9txyBekkkQgz8xoQoGyO/HGHBXeT71dJ8DDZaF
AobvDrzsDwTif0PfefLAx+phJd+QiAvMwwuJDQ6JtXwjJcdH/zbkwOcA+GDnzyHF9FQNaUMo79M4
1vqm2f98qQn66ma2tRZJE55n1R6K3XnX3KNDG7PUHQCB4Z8xJmMFv2vs+OERsr2r587iu0EJEX3P
qGQxDN5MmP7hSsfrMvMivlvVrH9vdgCm0ycdL/14jurI0Hgsbihd97pYVuNEI6MY3pBSfCS0+MWY
6VGAWuMdRcz50eEMVrigTkyFJkZhR8KlcEttc5HJKKxhSXrCMkVsDT7h5YAifMAbFyeJUv0FfdJs
d8O4mdaKUfMumG5Q86arVb2Amq5XlDu5xQeQyXUdnSzYXI+661PbkkyKsujRwBUVgeCVf2g4UmPf
EfoRF9J2+m0tRPg1bo0nNXw0oFOpSrzfJAy235n3ex+iWeNgbz3/AiGnTG/gXcGpK7QtfAjhbECH
7BSlARjTz/kfpHUOFuWlbShfo8X0+R2OIVgd3muf8Gz0a7sT1c7Z/WRnP5g8b+hxoc8Mv8aA9YYm
OmENkgUt5C/r8SSnzYlbNI/LoIj6SLugZUiwp2mTx+9W/vta5TbuHHHrQZQOy2PdBjZ87hNlCGm1
mBi8S0/2KMfrY9ygxlvgT8MDZ1U1vHq1jejsOOJhyTzMgmS8w8e0GbzCzEMthi9syvZATcib8pFc
pX03noewV+eBGt+cM7+3HDVjOMhu3CXlNsL7kDfhnZ+bjjW9hfobarlSmHWxD5Bw4/2mJuRd9fVu
dXat5PVoVU6DDu2WmZIxpYpj8RhmWvWlw2PUf5FP1tBtU8GgniX9WM4n6Oj3wOny8zf+QkIJKLJl
w7Qwhg77nIp5QBqdIjadB2uTxylnrmzrvWL0yyLEpgomH/qVzAMMoXM3sPjthRbU/dGG3C14Q0HZ
hsH134ZpWuv3ZrmBx08w5ub04r0jB24CKO5pcgkjgRJrczx5FTRo/R2rYBCDbWwNiSTQYsdVw0XT
Yr92dG0PdDJYOMudqWfbHsr8G8SD1qc/MXQA0Ew/SKFa1eQ6b+ZWhqZQVULLIMY020PAfpVomFuT
B3ah6WSJkck8d8tm0x76X6PmeC3tGHKuQpxxBE2OeKz8wIagAmjPFov8YD0wk+urVGdZrYeDHEoQ
8OUzfYVKJOFzIMirfQKU/XX/TQl1mLDClxp9w0798Pggqm9AhJS1tW6uWl5swU6uG0JskD7YiT6R
jXbl0D6ahRC8f75jpeIw1uLuEzJilMiH9czOtkOz1Ir3XsBMzeKEvyV3bPwT0DQsxhIXmu4gQiBM
8qHVUXDTOgNpT7l2mo062Gr3EQErLhrNyfJu07z8/nCC9rMGGlll4cvSba+muLJCq2z6r9zU9Xft
uzh2AXmSn/P60qu9JI409Q7XMXP8F3IstszAwmE3Jm/oTxKaRWLicWl4IEO/E9PPUO/Q1poIYkLE
QdUemYe3lXB6q00RqnBSMhWDHCPTsM+Gdq6YaNLKaVjXRnCXnl/ov0QFL0NYK1njMp3P4UgF3pB+
2/71gFj9saj1f+MWQPvt0SpL1ipSUO110JYG28gGfN9GWLjrbq+NF4TRIti5dqzQ0dWR7Z9mEGv6
Q8RcaH/zm1DCxbeVNAT0X/JKqpDdXVpGIUzKg7FwQhJX355D2bddtOv+DqwCv7a91CPXDT141e7N
vBCZVo1abNAcu3rXWQcCUXiRsir1RgvYZXFlHm67UjAK7dqVPCW6z388pHwqXaUcQTaw9t3GX+jL
gTdNLDpvLl1rhyv9Eikj3owb1sDkr4jHtTLCDp8KsOmQYaXk0KkcKVWyBrAx/N/5R8+XCJSSV6KL
UVxI9fQj9lnUkMexhS4W2A+IjGo6sq5k458jsaaApwZutZEfrfcRjPQLR4UXGof42jHNzzku7cyz
2NJEZCWUqYly0Crg8YWnS2fYDgYCBkC5ehpY9swYynfF4eWcdwcKDHUdpO1Us4qdN7alRnE9PQab
wSP/FZnOOgWejjAc2ZfORljCV5+nDNV2vYGEFbzIk5YN8lvDDGBgfOi7dpj6bFJjn8m+M7ONyfPd
WYVFmlWWs1edIZR0i2vf6bUa1uAL5fY3Ga0WRNStsqtU0UD9i2ibL4v/fmXdpu8q8Tfrd4g0YdbK
miVK44HTj+ywfuBmydyHwHQVnJIbQXsbGKWHw/efi2CK14+H+qLwQt7KRIB4ki/lFEj9109DkoFI
2J6nC8HN0uue/zeBHcEXRiBMWNPK5St0rqrbVy/5lTdsrTFkvMp7+qVMepD+Jx2dOfbqb9JaCl4H
1oKw6/pNxHAs8bsSFmTuTa5b/oieryeeGXKBJqdNQAbbQL9R+hNgbZeN6itDrrRQS5IXKZwEpZXu
+wt5Wlh+6IT1PQ+W64XndCc0raYXTvJv2kGBLhcC7cbXu2V9pkLLizIcYpQQgPMts0RwZ6OI4t+W
fhXX6OQ+gqzvWrMzxxiTaAD7EAQbal2+vTxC3xLULMH53eQ0n+7uMhlwdLfftYM2VhVAYvajYHJU
zYa8ubnxO466brwA0pxAkirN71xndN1H8G3OiG/bi23zyloRATVm4cyPCY6x7ACdO/lc9skUmJJV
MAVFVbtWHW59DwJoEh1eMkqGSFD0Wy1ni+BUiNT+cUy8+6V2EXoJnzf2WGTB0ekOEG5qeZQj9qvQ
E54al+fpURebkIsjXR3NOao2myBpocc+IGuwxdVBJsRszISbPxAnxCFu61z8uEdeIInhjqLtqgFT
5a6pgvP9UQQwn2meWRGhWq/cglub1Kah9zsQxEpO92jsrcAPjH95Rd+v/ue/eNdYqgqMoaHyVBWp
O17kLkkEUF/ck/1/jzCp9gd0fXStGIy6s18pgyRiZmVhUAP3fXdnCReK2wcAmzZ+xcNU4zJ9mO+/
PDSWgws6UXY2WlNmxDtqM4RSX8+HsDGKv2q1fdPloxhhM1HiOfCUpshp081XPs3WLiVK+yTX0Q2e
lI5eBB07v9jqwOczW/Jcp632SdK5wcKusGDMpYqHF9EEBOKNAbJ7S4J9+RN61iQBuj1Hiw3cqSLC
o1Ywgc219hqgkCn3HPuzdHxKKN9SO+18kQZXLKmXRxgDMs45GmSkV5M86hdLaqV8JiTucZNVJsj0
p30++TQDGdmyUdTdNBtda3AabQ3yVlRNz334dmfA13fZ94SRK3xzkgM8NfvjdmEmxapDApOtjLdi
ITsLtPRDO3S8L3p9j3gL6wSPp1KZiR18cPm5uoDGyrJP1116jnK2TASHX4w4VkcpUNmm/XqeFB+O
Er47cbM0ksJJl+nokM/HB/YIyl3STRvrreX2XGqniy1M9eBy/h1dy7lpbidqE0/I8XyGxtHx+yiq
ktKqdqJ3NQyeLeBzg1CqnX/fxLDFzGLDwTNf5S8B1qA7m2S62WbTlGBn6gugVotA9OBv2MNNbCqa
NtEzQO+K1GZrna+zhzi7yBObq4MsSSzXfUpnopfPd5Q1+ne4DZYEewOu8GeO1bH/Jratp+283AIJ
1boI6cp4bq7dRW6mvy0i/GPLKnYs9vIzxvAWbTVN2bE9li2MaXbpo968B02NrQ5ZtcSQSnd4jMz/
rAwmuJRVVZKjetuEZ/JRBwBndw21zLSCUU2+wFzqGBAh0RDEntPWHUw+GL4nvAt6KlMdGsND7QyT
QIlmmDaFzdmpiBRaOTIJURoGPf9M5TwFL/0K0dyITP3tcDIJ9qlRj0bNmUjsQak5eKhosYUucANS
f4lxgaetrQB07hhsCkAYBxuD4TjR4r6lZOtGRNIkxHM/NVUyJhBQp8fdHoFJ33gZS2/DQmWZFtRK
LXJfo/dgnt7fdNNV47mMwUs/KS2dDhMmFhmoVXDwwnVsVRhYG/xbw7iXMcm3qri8ibMLmbEno78F
2+8InabDq5n5/EfQXiUDsaXhkQSjHcIM1pyhsr+twFcWqE1MKb/r5ud+onvMkZrbBvGKgnu1YZE3
DXYGiRwg1vXghSF6aQA88S39NMvi3TqJJrLxEMqv0oE/GswN8zxJnsyBGIUWl9nXZD8f8Idx7sSe
G+o4ec+WTHPJzY6gGnBodPRD+ekqIZgeBnjMBINKJ9D9grlKUpR38v+AmKSbSXH48rzHrbFfA+qX
wG3VLppQLGNh6/C6BdM3akqUM1GWvWhlZG1nlsFNQZL/0Cs2pPCbajGSrfl1BSG7pqdeH90agXlG
i9wJlTDny0ywjQgCXFhBF8lTfQjjdP4HsDIrwtymn1ydAMpxvrYl78gX9DqGGUhp7g8KtvfMmDV0
qBtT4NuiFHeiJumnEZ6/z09ida1h8T1h0o7GC3MAwL/Y6BFi8TyLxVc4zyiRwuZ7bzicoPnwcOZg
JZKe/Ef4uYRjN3SE2ZyfDUb25JzBr6D8b9CkPGlLOHnNzv7S2uUgo6uY7ijqHklF4v/4NTz/spbc
E+V0MjN4Wzx+sP6Ml+wIThHxZxEGNM9EwyNu3rEwr8z1FdJvo6h8uFKASFCH+qZjk6xstW4slFbY
BfH1VfSsRsZkREl9tr5BAg4Z+Wr7YOGkQj7cLvwiF1sDqKE7PW5b9X82QKygBOLmSTUSPaIz5rKm
D+sJdL7kXmNjQELN5PR9hu4f4SQb2GwFhh9sMEr8xl1ge7jQEjqIXP0rXihltOkYxnNr0DV4gmQM
Z7oCDWHgNNr8XpzX70tnKMvIkclhHuhj8SyGjSS5/PgN8JbS54cdCfoRjRLd2Q5VBc+NSxjMgn6I
nQTy3ycVZfLZjaRlLQxId8t/66gSilyIyoECaQdOCjP+1Uba99rzNgmDRm0a3C4kWZp7TUjsltH3
m78QGY9DFFHCJfRiAUW/jcPtnf1sHmoHQMxOZLMHyts0bLpAJSlR8RqGGBhUNghX0W6guZbki6Yz
GGWJquakGG6ulfB2NiVkdjaoDZfEcrXCP+Yqk5BkXG2rHMJnju08e8YmC+MK6/mji24UsoosZMAC
sWdNzR3W3Ge6lU6Hn+QsfOVcoa1ZWQdV2djUrPy+/fXRGC5KPu41MG80sF5mHl558zfoK51yJbiM
VRJy1GfTAkkktASyVMDhzyMxOTa3uV5ufWwp2go1GjmyT/FAp/dgsr4Mx12s8lTOwHzVzHHVmDbU
eSsfiha9OGjcNDu/jA7R027XHJktwMWSMBrH9MNe1emUhXTeS5HKlT06kAbyIWR7vR6jhRoVgZ61
/YIMwyhOGrr911L5AzDafxVhKErkm/s9podP9LYodKq71QmZdTxzjlRtk2Pc822la7ccH9lnxux7
cVb8b6RTJz5EO4oJIqH4BYQv886GqhhmAJNHWsr3HrV4HwvnHEXx/LDsFic2X8TK2vH7Kx9ZLZL7
yhK+rczg67Z4curUybIhUphZusyEN2J+s5lvl0l5n/HxBFW15fewosBKUozUM2hGNWLBWxcFrRae
dI5nx93qLz1+tAbWnOwt7LH6Odl2L10iq0x/TfpwfUuOtm5GwxxwgVBBkVtPkt3OmPzSwCrUNNcC
xs8l9nqS6nJj44yTjD7hPwZ1H4c4HOfQKDbaZFrYss5tHYpZsPjAd/hP6ViGvc/khaUURPrNT7P1
fVhVhLf0ad6q28pVQZH/j8wYRKMg4uHymWZQC8p5Ub5gs0Ipr1ubQ6tmZLvaNzpgO0j/7Ob3+aoC
JEgk2ugSC+1glyk45XWE3SuE+PqCrd9KTScTXfKoAtHmndi0bKkyKFiEoVfCQK2BTgJqZooHpj1U
cFpA6PzojUSE9nKAJKcR1acZ7ZuIwIO1fAppD9W7EoVC4iDayNlCMeoCSCz81g18mqSUfiTAXSCw
HtDdrISDkwFMRz5ew6uNJ4qWLXPFOlbeVd4wgC4xL3ebVehD5czjBFK5NUagy1JFxBLc6odQvpYX
3X+gWqZJJIFOiiuEGnaWlFEJZnNavCPGutijoy1+eEv3imzOauQPYmB3IWsDzpJgVBLjBtPdx2aA
3tMjh01zxYoWlw4Hd6AJDEjyTADDWCgihrjENjzsJSaFvWqviA3e+PEYkuscx1rTpCozZgdVD4wI
maM3SYVfLRiWS+BIRfP0X9YA34BXVA3CM22sn2IeDCAevW5zkxSrXGidbZ9GzyLvufZMicYWWcMt
JtmIXCvWaveS+yQ/M/fx5KN8KkeYh3qlAeU1ntWpSZAc39Lm1EqDX8yMa3R/n5eY4Rc8pnXgF3Fq
DogpOivfBE3lRTBdTVerMsUsBEFYCyzuWj2LRznr+cFRbaja3bt7xLyS4W2QyjZUi7R3ScAO5ZQY
BkStjIzFRbgg2fmmiaNaGGLkJhCsckglwPrXiC+cFq/+XizPekKHaUxlPyJm85KGCVQ50fmidJji
0wUQNkQn1l9KUsEljvr4bXnbqXs/b78pSaoLqehh2CvEATBOZ3Ua0aAYdbqADke9HmL/6HP4UciO
rlhYnrk8Cw4Vlc7os7crz4PA321hTjBGIRm4PzTQX6jvEsV8EaZ8XQ5HbSZ7qTSGOESjQgbTcz61
gwyFXjZ1nU6l1NqDEA7YLHwVHllSCzwzGWBxLRug/zLZRdjE12w+yAkuNdXg9PNvvqDs8p3EoKVw
6HRdyvwjbtD+wkIVfSJvuwU8OW13HjVjF3ANMOxw4vbLKKEqKiINvBQMQ/1RrQWZy51HHj1MmREs
UveljpPig3AsOKcAqXJ4cf1vIBep7xb0jqMy/tnCtVPmHzev479WXq7dBWhbofrD26kp7tNC/fjx
GocxPJE5HdAP7AaFNlf0IMuPydDj8J4Mw8Q7XQeXKNHAihdjyYyOF8frbd8MVlYrJHZVc61wiBZz
D83lxzMX2EcL2BEbQ5NjhqPECO2gnRvqfl869QEU4IuVKIdRpuyUUfRpsIRtE2HUL3qIgZ8erE6S
KfQpmDRvrIDytFRF+7G6sjQGLrn/BZLlaIvUg6JlrE7uSM7rRfPYXPXtBoNlfi/uLRD6kfmBtzTr
hyo6apHabiht3X9qp0lMrfRdq2KOg4CfxfM29vPj2z1gnnqcXOWDilPsMx/vJwJiDbl6DAm5SLLt
G0j9dodYseEi0CF6D+LEf6bf1VoeGzCcph2EDIZ5kcLzIS9G979ZLb4u3+dLqvFL7NuavQ9wMWoR
UfllgPLFV46NAsiL3jA2cvzsJEBAWP+J2m3aDHlYL9/timZYdWSu3UtXUB7EB9/XPXew/m8BqB60
i+qRKcGrfJ92ia0xQGiaJUu0fU2OgfPQZCAPBKMTZeqi6XZSHaxx2YgPPIOdcg56++f4Mt9cQyNC
6HL+GjSITEgV084gwGNtNr2b9SjJ/XlRNAOWoH5+04svwHmnr//CvjbQDIutiB8Lq8R9aQeTjK51
T8va74Y8hpfYp9uz0YqrnX9cSNJklxz42k4+KaQEOcPLLHYC6kORr4D409eZ42dehCdhGn6LUmrA
bVbCOCtZGNtmP8cE+pfyXOusa9ue543s8Bdu/XbfGR+7QcsStBbl5gcwD/ELCuBeA3T78kiYjnCc
uC2oWjGSF7SaMMzjxrVAUCaoEEdV78Dy1DdhiMmE+hSdYr6ybT73ojgSENKYkye8HNHYb675MoLo
ctAtDROkhrbPK4pPRzpT5Wro6Zi3aepTirmw7wHC89043e55TZf1eCrJW17GUdFdVgdAy/aMOBUX
yl1Nlg3x77W7b7Dg1rcJvXVuFbqLe+yviOtmpxw0lGuGr2SeaGm5KfuLKWGyJhfAByE1o/KHi/Vi
Fx28ngi0PR52atmMUSRSlLatfGvchVwvGquQYdwFcQgAOoQDV0DlFqq4qMqamOtF13s/WtT3ZtwG
JGy9Hp7hL+kciblvA3R5msNaMZNcSS5DumJ8bVZVzP+tZGlFLMKE5FsplAm4XIMEPp0KFwVJEMTZ
AAMlvsoGa0+JjOXs0T53RKqj7gPmcexU2dn6HUXpzR9U7n4+NLPwrNUJUiWwjZncDQ0q1PrOXH5C
T+oEwlsNBoc36rx7rW7pNwqXKIDIanqId/6feCvCaKcMU19M9eQzwj2VjcG5hMc1Crq79o4Wel3G
1UgROvLLLXLEUak0TR5dQYvFyQkfl335ciw/sJSZeqGTPwVJaFPEk2E/VJU1LVAES5bvoKJcrPq1
wNEPN/JL/1AO6C04xGgZ7KD1EWtERQ77ifUuLHtMuJKnGHCtlEBsdQxU6bdDi2IrZHslY6MGrgml
jKLqjIcS5eEaFtP4zDZaRVU/Yw9gHlHWQb6m3EF6ghTNT/0pNS6dSArshIjM712tP1zFP6qzzOki
o+Z6nz5TX2v+P9P9MbCc6MlneUKyrUoxHecG03mgJv+KUKiSiuD7AEADVqF796eTOM/Q31nKV4P2
PvBzEkcvZvM7PXYN/v89/h7LEYFXPk715O5SfUIp6crRBKY2yxX3xTJ430pvqjKGh21evXPcgdr6
nxel79WIHO9EKyUs5cXWUQBT8EnGNPe7UGHhYd5r9+sRGSPmE6IcF/8HtDQcCQDgrw41jjSSoZuC
R7vaoHdmpxJEk5e4wUcqh6sa1Ornp+A6DF/cjI31Ey+ztcYWR1F+Ny+idA1kqdzVhvROzLjTFFYs
MfNTb7T3BqsVKu0Jcd5TPrc73Y0p6NUiWZJXoKkn9tOO58odIzICFJoYDrgzDGJHf3/ZWUrvP3Hj
H57Cc3wvKNwKQ8GIE4Ke57E6SN6ZFR5MJixkVKg8XfvuCO6FMl7uB14qZg5/WDbpYFaHTvMAQ6JO
S1uj4pS7Ehr3UqiS7N9aDcO8bbwCppqfG6gxuFk+P380G8WcUBSUdYIE5mxfsyixwsWB38FX0//F
UbXt62XINj70/YlyYHB43scKbiLBh3EYDNgVsbVDwrcQCrK3RWJ4taKIy24Ibi7khd3db0BKb+tu
N/zotuayGxEUP4DCLvSJEyl0EN/3tg6KMWHpc/GiZ62BGArDqmOOQ6GmvYbo1WbzQvyt2/63M0cB
TneP2ncV00EtsbQBls0OiqtBq7/FQ9MenD8XYsuHkfgDtPzn82iVc80vfnJqDaXjvheZi4KOkOrs
ReMKY3AANsWRyiQGMqrLJprTH0Cz2W84aEeiCbubrV1q2TbS/YEpKlWU+PMJaQO4378HBzoYKCz1
v/7DnDt9e8OaJTnLOKYo34Pr7jNebJYGDDDSrsDhGTe+U/TezTBwiGSWE5neenhYpaEbzv+yJ7lM
pJR+QQd4LItLCzBxRCJS/w+6xtBht80h2pSXMhG3oDVmtTayWpvEaSl08qneD8f2LH2fOLwHz69p
q9dUwDz+92vtk1ev4X7GXdsBO3DBiZRCIZ4sHGwlJbkAvRPJ1RQGw74Hs4GdJRBLdj4PtOWh6o4q
DAbpUcdeSfpXA6EMCzAnokcTAi6RxNUbsZSBHVRtPM1RSGn2ygt1WGF2DE7A6aeKqOdnbG/KuNg1
LdZa8jeEpVWvffp1FG/XrwWliWggHmszFThRTdWD+Ev+3gRQqUJJfk5XaxJufUcCSqfDxVYL1gJi
0PPkjlzqrJPMlINyuZ38M8UC6QPFD0V/7B10Ie97ECapKfg6Tf1KOSoJ+C3QMK4lN4ckslAJiZIT
4J4S5PqiC9OrJPP7RNkiKZX8au8t1zbtSmHTQZpwpdC8xevjGzESns0vC3taynxejoDtncbsE1zC
V2+IsMRmjA8uW2DX9nSfTDx85o3zU48y8aWQyJmk4EntQjymuA0EwUY75RPZpnNvTkp2aP4H02OR
YTHp/+iIVh/2vcM8cPWL6Qa1zpQXXl0N1YXL8TI9Ewfzqvf0TT4/nHQax0U08TU5Yr0HrLyerg+O
WT7dBYK3O+EgWxI7maBW09wZk0fW0/1QnvUQ270MbAk+k+nHKwC52GIDfpZHWPwRqhotvUDInc3O
Tfma+cL3f3KptEDW5iTZzR6lxD12bXkY92Epy/9XU+GCDZS5tTvBPFpNDlO8QKtEEq24dvibDu0w
gevbc4SMcoX12qaWj2L+kTt7dvbWjJ1KH2VCPzNt5RWoIWSdcex1oyolD7WtfQjGk8V7DUOC3ZLc
nQ5vo/H6FjtIqI8ImW/yJX4XJQprwDS5Jr4NDDhMhpknLFdVMLNBTA3yIpY6xv5kLIapgC6/vOe1
mt+MaD2jUf4OUCJXe6GwPas3CysujaxgXNWX1vkZDXQuAZw6ffsLzd+w1BsSh2cJqxaG0hO5Sjyx
Mkg+/BW5au3DO45xylWbOkpkAFHQBvw1J/DHymkoYnb3b2UXc5WyBZPk3yXg0zYUt1QNiaF3tRvb
CWGXtFMrJ/xnBy2rkZx6TM2OoVnl6Q3fkmiMZI/1RyU2WdXdUk8C6sSiQ7LtvWVQHLHg0pN3G40a
5lnlGY0lGVeVhObibiM7SjjHQ0if7TiMZ/C8sRWvC1Db2L/P7bJ1+3kWvcpd6rNHzMFKlqLenfsx
nnvqlyAun3RFMOCvIvuzHqCOTINtLuUtyDJdDNqp4/KB4DyQQ9eNxR1UHpIpkbMlyIgakRZWLC5/
7PazGRGJnCJLybPbtRJqO6bA6Kf4Ej9KSkJidWHD6pMRs6QUGL4H6BxLr07E584eOOyY+866zb79
vMwl14EWDKB/7IPb3sRRwdnV0c/XIvCQW2wN21/aKYrmBWlCLwIaqq0SUFyyXy8CmEcaV+fFyq4D
4/PH9oi65o9e+lFmWcTF6s+bCqOWhihV9gYGhENK2TrEKKRDUmrb8L6nXloD9hwwbvxlegHk5Uq5
goja/nyqt3mycLLsPoiwwFHujQiYn9qO2NgWXY0xoUeycU8r65EgOgV6/cXr3bY6XarTnB7zM3tZ
b4TkKPx897CXL3d9wkdF1LqDuVYKXHNDjQsaI0WTGlVLnTRxQx3K24SpKeR3q8Cq+OSPuEM60X0O
nHbVDR1TWArXNtUuj149+BdyELR4GtFhLWuTzuRz2t61n4mxRDrQRXmLSdlogs7BBwiL8YdXSO8+
SRUscg/SbglsLry7VaF+INV8U36kJatgh0ayRihnuIhHMC4vcwzEZkfVZtHrPWzf0wUyG7a9VfAs
BWpT/e5L9pq1gVquf1FFl/g03kkPoUImy0eNCLWBJIKOsIsambdtbSuLIjVjPrY9oJYW7r/yeTSz
CDHhuhamUkfTU6FqF9ZMIDBqVsgs3rFq/g7d7kqBhKdnUzVngrXZvLWMKj7xYImITh1Bhtxvvfsj
CQbkd46wI9WlKREcf9sLPH+OoOUppl8zHQqzjEb5tzF1N4sa/efNZ4rf1XQqqxnt/6lgb7J0r9Wu
xMuHVLiEqGw3Jm6vA5k8o6KqMg8OoOAyCNo1VJ7yA0q7aOdmguBGEMXBicL99iDvYnJxvyOopbgM
aKsb3qf4exr2/ki+cAvQ36h6aMYmANzcLJCAxaHabC1ZFTzVwUiUeZ50223rDaocxyEIPGuQAdlH
GW0NHAdVxEH8fHI1hmISpvjmeemW7mfBXrjc2qlF441mcQ3es+z/O8dgTB9w/DL62D/E9/S5fiy3
Pm1e/1QsHNzwmyFOVVrZc1X74ZyiPnRUhMAKFsK3PCKGlef7y8fMEdpD4bbPKNvyQ+VDcIX5qjni
XoNhW0t/t981plmT7/xOERE+P2fIstJgHckODWUne/kIQObekcnOlkAx9lqeb320JOUIRhgesqgT
uzFM7C8SfnjVoFzFCTnGrguQrs3EHo9NT5lxOVvAzdQ3ly5V2kdF3XBnNAda048+3TSM2C6EoaRD
aU05mSvIpHxT3Hs+5VfTax9B7O9+BUGa2XJkNls+Oq8d3BmQUm1R1AguxmBm6+DasKN8LamKRawC
k3q/Amhgh+S40eYg5Tymn6To5o8mkEOGVoKXrrIfg5N/XM6tMJZBmLfyC5Dus2Nz7rVLJqmQFUmx
hpbVjzdE16ZSRThePEz9cDJ0ikVxlWCHV36aoGvfTVQJC1Z/ahB1Om3XXBl+8kyvaBG0Hf6uSEwh
2Kb38dTq2dJs34nmtqreY3ZrnCoC8WW2CVJlZUCxx85fRAgfF8s/dnXh9Si6gVrm8GyHV/j57lOV
e2VmTI2TXHcBq4wsDnkoIwVAa9OW/LDKVc4EVrTM7DT7WzBOgW8i8hFWhePpNN4wWKvEUCFxcaps
6f/QHMh8Bu3ba4jjVkEQS13d3IJBN8VsMm57akyieEKrxrbKY1iphRQUo62b4SykuiZPM0YgwwO4
SmX0wfZUjLJcNs3Ne5eW9Dzufftj2QG72imAgGF8AATL/3WfolyAC7rgLzgS9S7QL5/1MJtdNVhc
r1zuVu/sKnNqrLOoHFy5GfQK93CxilFmK2nHLa5zpZkpptOAa7wUW2fmK6cgsd/FCCrFKNICre4E
TCULLg5Xwsv7IWqKWiLpIc/1j/zIQiSDG0ZGogrW/t+3d/9vTbkzp2RSpeQ1wEjnGb8hxIRpUDzP
kIdasAsn/WOkQLLpYky6ip+sjrssaBlfkJ74SH4iRVCAMkRMyLzXXod+KjlgHu5We3caQudY4mnU
wPABxHUuR8TCg+9/ZFxObJG2byfREIBpLEgi64zMCjq6fk27TxoA38Wj/yeUCKq4dv0IYIQDCPQL
DqFk0XCeMCr/v7roSmI+1i5lVzMsVd5tOO32ZkJ65eVz/pVmKyzBJ+Y4ojknqa34+C5aUZuswHk1
hm5USKHYOguVq72DGmln4O9DbNZgVEiQ9CwvZtA6wSLoNdrt+KuQjlkVsBwXhYf2uYzZB1F3VUcY
SfMHW6m7vPfODIS0WP2WG7ePQ1HEf4916Av54LQhALzg8PiZ4664TamWu8Z1ssOSNjTfkz26zJTu
znSvG/s0BbaZu5JMo+BIQCX7SDtWT62hT1ZgHEkxXM4rZD9CD7OAdLgE/F7OUafr01+NkKuzW3K1
chyLpWnERKmeuYHl6jO+SIodysOCEvzyL/B5IRJjGVd3FJHtnPErZ7QxDJXjGor/cBimYkSvmgOR
EjHxyVKM7yyT+z3XBfNVxzzo41luUA96o8qwCtz/7Opm4RK0/Tuv1eAtcRUDdJXtB8LUHEAgRakB
jOrr1ZRniSWglToA+3NTxuLdM0dDjlS8CmjCpBJLHsxej1NhzMYt/bcV76ZZ8Aht4x0pE2t2PgEY
gGEvDX3YBkhRdmrII4900i591lV1z+tGpr6w42xBFdUuVoFj+o5odHzTuNB9D6qu+F1RYPjYdJ1u
fo21Xm02Ktycu0dL4J0Mf1D3x/wcEs15zIcUCEtqzASxdZJK/XXtfd/RGxEVIGIHmzhQCIHCMova
bv7/HMsVFWCSzey3hNnMnrlqkVrBwtpQJZtivG1KjsG6rmI0/44zr+hYHkpUgF50uHARaxOLRFEa
VjnRGfH7X6oDLdiSm3KPGAsiM9zw5SP33xs6FKWpKyNfgCSYSp+P087jesN5E8bwnLwPJJxeIwDJ
nTnyMp9lDGzSem0Z5YxOe71BMzWrPv/BeAaDm520IuVc/Al3K4ud6746/2TuHxwyK6bsHad4KJnq
+EF7YsoMtceVhmtnnCzkTtt83VBN4bAGBxQaH8JQxGmTIoh9VKEVSXsWlJDaF4hDHywyBV6nK573
TofQMbl55Dw0ToJWs+b1bvJIzGL7gY2Xy8DE1Jzik0xi05iL2hFXVkXzHfdUoblAHMgUoR2SvSxr
N9j6mIIGkue8xqixignTk464/4XxGKGncqjNlaLd18toSPNDqPvnwzkVc24adGyE0TxiQ6j7aCOX
+zq2To6Ybw4FuSKH+mE3QniRTQq3fDhXQM6YvHFrQrerNJFec5N4ceXBsWRF2FG2hBeJ48EGIX9J
LbTZXI0+cltdSThoLKvq+wrU3tIxkM5/8oJ4aXehR+qEs7iDXOQwtLFgU/sFXdfkNDFPYk6IrsKR
0RXOQd2pHfYaGaw0SdFdYW/UXBF6Da/ljwSst83e9wdlkOYd27Om46Izdxl9h2/u46FgvwRzlSrl
xzyiYNz6xiBBlgQbpK5wfviTi292Y9IGAoVzCo9N1ktNaZWef5xgRBPY02X13wbt9aXpBJEys5mB
AwzsQFXigRJzBYIkienCBRlAOtSX9xtJrsvJ4MIeliekspXbdairZYbIguE+8t0iZNCJRs1o06vX
idyEoyUu6pvXO3hjMJZLGp10dRN3vNI1rEyKWx9WHv+FyltiEV0bTAexQyyJdEDdgi2JB6JxcM8h
z4thhTHxdq8L1VfbJ6ulK+1jqlIifjAAC8V8YAMjUMbv7tmH7NHX9A/tQadFviCMyz885OUJhjZv
/5R4KaP/DqKFnoA2UJEAIiawaTfQ0Xy4QLuBULsXFUIkdYYZMx4fx+VWbfUhhuD3EUei9KYxtPd9
7qB5We+7bufz2+Ed7WHl80sMHGV43irOraE2zrqzxzjsYGWfq9cs7op/6x4LJ8nnhWOfX2HBsDcd
g9SWEwtGXHYCvhI7sUfmqSXTRyQ78eCLuk1N71FdYNS6jO3Ghs+PXAX+4OZutFpWDjbBnc52CRke
3CiHU+PoneXGupN6SMcKt9J5SzcI0odBeIlhvT/CXNOeRI573lq31Oe2Q5ZlJCUBcvpIP19/m5/4
XddTwuhVMPiRTlKkr3iHcCXPNUuZopBHt7eQu1iALeLMFvvdDIJz2Q/nkzfglSxVIxHZlY5jbf7A
YYb9hkjb9t4lBIIvTHEiPZXjof7KInuESwmxn73bQEBxcfZ/yCshBHnUhbbZXFCb7TPwMseypHb7
I9qONx/BUCE6k+mqLNeZs7UQll7Z8h87vjfUdp0Eb2+pjhY9F9jLO6OUSsAcwHm7XsLd4m1HKxKI
r6qAQPEVe1RESuUkiH1yX/0NUzL1MYfAAWjVn9clNfEL9irCb2MAgtH+l4K721y68xiH6tairZhb
NjKQlncbw44mjiBhXWaQejvFdiVma3tNANOHtTynfBf88BizVGzjcLRplR53Hu5/9iX+JrbCqfff
IH9QueLpD0QoHxNoz3vZ5CWSadPvObVT2+0CpJPFJ1elWTyAy8Y8kZRrmk5YohdPuo3Usue+KNbJ
waZ8n1HYKywaSWpalSNztqssyl15eLfnTmtiOhO6XAYgN9vGTarjw5EiRAgtmdoSCXWhI77Pavsa
b/w7hdHDaO/aNQAtBAJUyWcpkUIQ0PAEWNDIE+JQyQkBLMJQjq1S72M0N7txxRigfHC8RjcZwBfs
GHpVfdWbTJ25zI75hOW+RdhHokliVCNU8qRJLjNhcmYSCKUgd6hSaqIWWggQSsQczYbgDoxFt8VB
cg3VNKrCLgFWtTxSMIY4Vu3RZNyt9LUiM4Pw9pNWvJerPDoaSmGs5pM4u3F352pHPIx+u9ymPSz3
P5pWIyc9Q0/Nr46cDiqBn3FGCw94hwkVrGkmQW/tKv2pPYoDTaJy3UBcFvHW8NqHkxphcELiCgyL
y3lw90imIy79UtYKQ5y54TCDENu5y4CY3sU/1XUfytNw1QJh5NXRDsW6U2v4ct+tMHrmrAvSnlKf
wALvCaxTGPNvmNBGixndhxJJXlL9Y1L8b2TqVMTGZ4yu1G+A2xnrTXCArQFEmtWOjaELWv4ZDAMa
jxH1hRuEKCzvrakt67SAaKrjjj1am54XEWH4Sb60B0x/NeMTTm/m51XHEySgR+OUZD42z05SrsFP
6jvAdjcsTgLyOFTsZg3wA2Ywdv0LckIvM1MvPz+T3i/fgtvcdfSpD9eQEJBOA7DwAsdoB+I5lriw
Uxz7PX3arWhFnpXVgiC+9vC3bJA8bfGkGPHGHNmEt6/xlrGv8tpELXP3C/by6+MymAY8tt/x3KKt
0kGScQoEsqo2T8ibqb0W9uui3iNP4V1URCRsVZa1cGF/P++rNUkrQJ8IySb/hPBMUZfCQKEbRe+H
zZoTCUT5KTeaWTtmqPXH0gJx3OfZa3OezWZtzXomaQRWAe5KisEbzkfITWLqZGRns2EgvuSIlzhQ
hoUpJXt3MEg1Y+L0igVAAMqm0wcz4Ms+aeIsepTWlZ3NcK5tXPwUUlpFX/R1lC3+LEIGeJ+ECgXC
5i+56jZ+U3x2SAFDws+nG2RCwIn1vCY/XVZy+yBHy4P4FMEXHUKK6Zolc1cejrmvNHrKPOoRJfM8
qBkv9iPqQPRGAAjBidGmL/MFoqDRbYj3sbFK9FrO8RogVKGKsdGQ49ooIWBYED/Gy0Qnqdhf3IjV
JcJEHcvhrvZ7Z8aaUfMHt5uwvrjCau6rnz0oZ0RHm4lQSKpMq1I0Z22G+No7xMpK1Sbztejc0aeY
NYbSs3dzeTcT/TlvDcXhu5QDavC9PStJpfcGSfsgXnVysPGhcMMv/C7iKjWxu7X/Sdm7uyQVK4VV
VRrEmM+KWY6oWT7pxDqBVhuN2Ilo+oI9MSVJyHSiJMjaxy8gMwOytpppDp/wFIzXTWoxrlbOkpTh
SjTdot+m6EIeR5VmNQ0418ga5IFbUV/uME65XHHjfA1Gjd77d3E3buiefhBZpKXDyMCRrG6KbUod
pJnYpNUrtsqotUlL5DnSGSh58t9jmOnuCkV4S0GNnEax5U8es15+g/7EbR09T+WcdzMzfr3j2xG6
LImXkiNn38YAjzjSimx3WjLaUH8guC+fAu311PLfdV9M81/DpYZ+sEHBy+bD0NAnexfsstDCQxD+
/Q8kZvBAoPS92rletr2yDTpz8m3cnCDUti/+kyH+ItFBhGRBqQWsC179meM+owvKiiYc2TqaeDe1
GaTk0pW5fodqX2C8arptcsyAvv6Y6xAjENAS3H2fBca2WlWFf+c3PpLMcjp3+1NVe188NorHmWXM
a7+dNho6djdK1sT7FX1Kyf/7DwTkFHID5ymDc+pDJ631FKEvcBIkjMdWjjHGUDIeSKbIKKUplvwZ
inTWVlMxclVzbM74fLqqofG2iMVAKJENtAywG8yEp6o/K7OzOswFjQ6Ch38sCDg6vsRZFdZd2+U0
01NOs+TjpeNDzaeAbDO7PYuurYjY25u9hL58LJ2i17xZ/C93ROX7l0+eTS6ocZ4iH7q5EF+mn9vP
w1qA9DNXmUVJKrpI5WqxCsn/uZZzcKCYhYY1VkTZR3X71IPdbs/Ll8tO8Jsx3A+p4VnHLQOmPVl2
WtQYRRRwBpeL/FvviydL2wyVLxKQu9yLF5TFJRtYRLFUivS1JxO80k+ETRq6g81IJ41IuRVjKyLo
sxy+p1eBFuA0wZwi/F6+RG4V5eaXMGzYVBz6781v75aI3JkbS+5wm+OIdA1Fg2gqfzFyWdutNX0E
1XUAJK+F8MyzgcSxZa7vHHPep0zmddBNSiKM84O66+ycIxTOgk8yuUzJc97M6xlGoglHAJSgJv/D
RifnKQGTNqnaYR/ISqHX0kTq39MlnR4eKqZTTqS5xaGTlrA2+3OP0rM0pGlfDR4dvUV18Hxgupvd
E3n+gNh6lQlgaCrkO3/DGr9z92zYhx7rP2MMBGwNklpggw0VQs3KWsrrEdzwTw28KUC8RctQIkU4
48lMgZ78R7YFkINCqrPVg+pXCMgpmhL+LWsaYc4+HuT80IqLOeW2szW6qjZIEuhzRmCSTnW5c1Hp
GCTmA730H7iBnnZ0J89FyceoR19ipKhSrde8fC09zImzoACcQU9MJCUH9MIxeNifuynPiETrwM8t
04Oug4G0e0jyVYKTkqyKvyVX85Dm77WoxDAS59i1tYL7IbWsDGy6DjNDkxYW+rV7LCI5Hw6DSpNI
SUFP4O1uS6dBa7dPYU0yNiemR1ijDXKyYE5ikM+Y1FW5PANkrzbTmJaG3V73iPL89+7t0g9TJkfc
bkGlKeykpnu2UYNtwFoZWexoChCtwSlpVJmoWV4C4RLEfzmvl6iaYiQIuNZQiAUMHF6YIeM+k0r+
V1przcuHoBVGM40X6Ch8dcEkIXr3X2oJzBOkXCj5dUlPKOH2pwlEbnpsbLDDFQsXjYmdEWAR8wyh
hDTaudwhkyTigcIAp+HvQlKfklZRX+awkqcMUy5LKW98O4FRiV6C2Bwb2pTU1dtkLllTq1wWKG4B
htIKnSpM/rF/jmnYFIeHrYAzSiA0szWlecrwm5kNXMYsGdyxI3aJFOJoFog63Kw0ANAnnH1Jv1zX
mTzqwjMtY82DdbYEayXScr3HDF+Gm4THttZAKuKVaxZX8CpId/cIIoNg6TWWXlhpi5980VKbRDzV
IHQTGJVLEv4Rbl61+3u605LK8AuH0974VjX8erQNJ1GGMirDWPqUBYZZ/OzhnFhiDwqXNSdwGcAd
LvANeJ1Bn6kzd4+GoB0Ks22mvpiQvHS7+0vhjICd9ZfPfSH6wJFwC09hIVMptUtSxtZsiQCsS7LQ
6BnQNa5KoHz0kZ9afYf1nQKk3Scq9RE4ZhzcNep6w1FPrXo8a/wsgfg6dtCSRsLZ8qbzhP7ZVE88
Skeg7zRQhdkEQH2k354moTQ+T7C8itDrbszzKgf1KafwYctfyiFmc3VoXalqF3o7YgM09SO8L9cD
2hm5K743tl4PhJkpoyz/vuSeja/LK5HxpIP0tBtK/cDbeIMWTDW6OkMBy8mLJiws1UFB+ciL6pyQ
PriYF6enrxtYABuwKqGTkb0a2xDwf5NxObqzqCgX87JcKG7R/VSrVosPhTxZwn5fgwcsgfb6Ko3G
xDT6R1T5mKUs+6C+GsdhVX2+Tp1BVl4Q6hbpa0nhN9khDkgfoT1waN5JEuG1eBfSMD9cFNA1oJB/
YRbs7s6o70hwMkZDQxwX/KrSYgr23NtdUAr0/8yZnRhPyEYjKPhbhRN9C3IoxFyNOX+yJicgL9EN
Ir+4lnDReEXyK8dsB9TbgKKSGK4TM9j+41e336wUn9TakRGHOBrKPTdWDUs8pecVxrJ3ORuE9gQ7
5814qeKJ3cph584Fb3WLERKJcohaCazopjHKxMKp1va2zIMB4tQQgkHJkVYZiOCavr1psN/Qm/wX
SszC/A4HXyzAEp89qoQRDrnJdiED+tCc7XkfPkJWaerdKp3fBkLA3J09U05fPfQjhxyWrQboZMty
+wriD7Fa1RCGIzIfeTiRSWNpwl+d5veiLuDoRyI9e0dCyhdWJk6KKk4gap9Hb5y778rveI3JAqcO
AZuir+D0ANzLc3TLFUafBie9qfqtSEkfDCbAdje+1f3LiZdlH4P1NTqQ7upyXzbiFVtBWYaNRHSb
RvmccsaU8VJXBC5LBa7ZGQdYEqhgML64IMVsMFB+UoFODo04RcL67afc/J+vm2OMOYh11kbuLmTF
EYvdYaC5wyuKq9hfctt/7PeOYkI2js0cOs6o4tQw5sbGpQLhintLWcONMDBEf4yUCQ1WgZhOVNeu
sEAp0tt2vQGBMw61ih6ZrBI4hLMTGf5xe0FGC1Z9cEvnRz5MFhDGOfZ4VlYy8XWeP9gA3SlGCgTv
efboAEDchim06XNW+PiGPV2fl4Ob7ZksO1X0OrRS9kqCoM/rrLy+/0D68WBV2VMT0M1eA9D7mFQb
7d+uYeBA0cvPAsUn5MSwak2Rtx0GD2enJAGZhE4GJCf+KFhR/j10DyNqGavKWtHQh3yeZbDFOor6
uuZ4mJ0zKojh2+0UzqWVx+aU0FRDfDDjRTsfH0FYcu0H52dxaPfsp8dVxRbYuaSypTVrEIUKgWEq
yOFhIEgFKaRikVgOuBUkDtzC70FOJz5U83j2rCe5ywz7/BMyPGWtQCUjElxJi5jMNjpyi0n97KVS
U0UIklmxTrSJ1hTx4hZIKdwI8WNRDX9Kwbja86B3y9ESkIQr0/pvTjwTkAcglOtvFIg8R1uI175p
0OtJVyg4N8ISGVM+gyPk7ZAJ5eQpIVmY2Qt1wMgv5rJ3/9tYPnpo7j9ZstLZ0/NHSaASKaa+r28P
Ak2BiAljBJYawFM98gId0JOeZIsnm8MPFNGlxGJndJwJmDzXBN13kd4ZzZSAnJqJnzABAexaCTf5
PYNB+UAlPLCzVq2ICTmJL7W6pLLjHQF+gPKRP6ZX6tG7wHhOxDdBWPKob8He8pxjQWkNSIUoyeQr
Iz3j/tkFxx3SVXn1OeDfRL2NRBMZAQBXwUV8DW0846iz3+wb2OyBzwxlbuWGP17iNWH251MeRMnI
RG+Hdijtfly5uVzr3MLgFRAUfgW0kdBlk2KW2ld0roxk0fcso3FmM1WzbY6q6WSle/5OG06e88VQ
XXDDiVfE7dhsO6tEQQjLzbRnMxrhQg3YLPE7HJfWoLG7raqsd9YdL4jXJ+LOQicpsiHa33NuQJNr
NIBLUCVMTd8FY+UOUpWi8/qjgMAxaoXUsCNr+5VNQMQCOYMEQ0PxMXZt4vgRrNjgjL85UCE+g64q
kuyDXJofcVjaOG/SWI2S9ASRZKTkc89dWEPdqRU2bWFtwNS7yQsBEoQfGPJntCeFWAtLrSyS1GrY
zKMvNJm5/1nksiA3DfpcU/8bOaheO5s/4WbmL1hZ55XtFYFFxySKWjl5cok36yw1MaslYj7/AxNo
lgpaDGWTtaI2NNOLDy2t19KkEqQn5Y+sJlwySIiCmv0HZvztgK6jjTz2Be6oX6+YTAJ58/IQ2L/q
7NMZEP++VcVDZ5rwvuF8EJS7kt1464+30mWuiBuRyBw1hrTDe82fRve0DSA/CrDrH6f4ZPBOQvjD
dzWxay8Fjc8N1IoTdt+gA0bFYSb8nk34pUQf5eBrwHa+8zbTZYZi/fwaTED62oo6i8WlVevgLRYs
MWnH0xwsTFfXVVES/PPJFr0I5Op+vEJOaSpk4jfkoBB4kq+f/E1JFdUvtvWiDhEhoXeO+9VxidjA
HpIYLH0smCrD1ofIG10DqqHOW0zZmPpQM83tYj00UbWvp8vQ7/u3sCWB5ghAOYVYdUcNuPGS60/t
f03mTPHsUQO7L2PeUfDAxiNs/m9KoDMXqTy1cTa6tniq7QHQDSe1d11bCP6+FfpShUkU81T3KOrU
xE/56c67CF6a1ruIN6dvN2tmkk9kPoWimNWej8uU4MXQ+nCf2h0fMXi2KMLOY5ZlxXjBzYgOxx0Z
yF75nrrqQ3fUqahk9eb0ezJV+4C4nfJDaTTFSMMag4vx4/jX8E7jlxp1FD6ebstXxcAGS0gKUOHx
xtY9F+qOo+vkjs8xA5FYWWk01S6DTjFawqEmX1OY9Z6UceuD7nAY+VMWm1PdfzAmpmZtIpWaeP61
A7Y7+YnR/p9Lx9ZW3vkLo8LRrmWfJDsBmCuhL9sj1OIPMmu+9D0nTQppN0Ox9zwitUnED109iu4O
bedobbGA4miCPu0u/f2gsuNTJw1xP1DKnoXVNsQeME/LW/ucjAVoZ0E1XNg4tWU0W13xEHONAQEm
HtxOT7Y7sL6bd7DhnNjcT44z5eo/zA3I51b5UnCKKCuetRjuuKZifHY04K6IlCYV5sFYS//ZNHGL
FYWuWz6qZdoAVi9SLUi31A1kKuCFf1ajH967bdFq45oNGiPBShzIKnPn3qOqgO3k6ztB/sND0zdo
k9nzI3HKHR/hOw5L5SrnlC3HYH4FUxVqgQ7gwV1GDq233TeJvKDTpNwSCmmDEB8M+T8QO4+0Om/o
VJStjaOtpyAO77VNTvleuv6ywH+gOUUjhM9rICYuZwU+JTby3KOYOy0HthbsGT9aLh+EBzqhTwEo
NtI+8h2QYnNXYVnq9IeYq1JbBmw+5a0QXjFLA6GP56hpIiRW7A9sqrj6rUGsjE0MOlLZ3odImSYf
k15OAS/fYzCG1qjnFHALpYKFFYXDp1U2l2K7VEfbrC8MGbsYvEf+KDLYH4TL7vIb7Cf3rSn15Lua
lmaMQvMbFqN4bWwMDcs7byE3iZfni8LOqfUNgCkotQaicoBhNsZzksakUEMN2vTVU0u5zimLpQ6x
WBQzhpSZXF3Y1DFFlZbJyvTwzfQ70KYIq251HwTgcF9um7fExa+W9GR+Gp+OrqnGnbsEx79eaHzc
TMTNWGVPs3MXsHCEfx40zB8RY4BaeyVSJhql9vnWyDt0HCsgFP4+gtJF1xVagMQ+U5/OTX3U9ovV
kZQhge7zXoI7xjYk9AoGjh5fIOGysznJDtfjKVBkWaOWOYnJwxMAjLL7kIWAjx4It3AYcXVsPwDw
0q0k00tvt714NeUOJzfkUja2CqdoYLMlAsumdfX1j/pDwQtbhngVagBIwucZaF2nbG3D1q9oSz75
lDQWhtOT17yfI8DUE+FNP4pzXRr8DWl3gVxpAkLpNfBCGtIagRPIJ9Yaz0mkQUuu9x2ihZdhXNe7
5TK4yAugrDnQclhWZyd2Dg4lK0FBsoE9++bgIw0mRLGV7LR/6rWZBdMfwYk5k05i2XkYtOYBSNIv
v0EmdaGByPRCGWkzKtQCLryy4qTi+Szlv/vuXGWhryX0AGnd6/1ZikQZ54NTLnsc/OY1LNQW/DkR
/U9Dd0unHKWXx5hZYA2G3Pl1mAT6JS5SVuGN6+pT32wPfK9cbYiFVsD+Q1hKCHfAOU8CFbRqKS2c
fRlUVblRBidgLXEPhjbCTPDzBxifDpHOw/bOu0tf2g9t/t9yk675Ll/Qy+4JVC6huxWoi6/jQMtV
HGbagUHSLhrlbg8NZy6JVpRMc4//7GYC2gabptIw3KN012ZK+wwl8vNLKugJdODmhQv//x4dyptQ
JVc/fHrOuJcRORrGQaNZUbYsI/eGjTlbKBmMp1bUgoWFZPOPdcfEgUmpDvul+Zj0BeOsVXCTTASp
dhNyno7ueX8hL6CwjYyDQi5zq5xrIqrDA666IYXZ/HX2bSlUHaTgj9s/sfUUHZh6jYymAEtanXBA
O/WNj7jcbL90ZGvE6NVKF1tnF13fx4WG/LmR/2/JDmlFTXw7lpHIqXgl2LwiOl6sEyPEmrbH4m0U
8BV8S+R3PrltvaOzsXxEtzmW2gMje7TVVz1kOfISCYnSgOeHcVfR7CdzQAF/rchhK2vzeSHOUVzb
+F/8YKEYDOOahQapjPELLoLVED4pzIaqh2qMA7cnkncsyiMSdj1Eg93THlOPkjHHr/cgqtKrMw1F
TQG3YkCq94ZBq3mWVyBjlp39536yLEJWLQ68FML9R8N8XKh9lf+wPvI9i0xzenpgHBlk/Nvb1ANL
6mzZqhF1GphLHSWGwZf4QC8IuZyyhaE8RxFgG7haFVTgBh/EUVyqSNJnM2rS+i8xc4UPy37WlJZc
mmReaX0dKNbOAiph62yGHbLmX3Ys7zP+olkF/jGa4kMGPY/nSKWJKsDqVU2GUBU008xfI/GQSn24
tXl1V5ytE3Aco83S4U5DoCefBhmPhG0kTkGVO/X0q/DZCv97YLD/MdtplD6rd8FHA67X8k8LeGMm
lKh8o+vD5pQsB0LZDu9XF8Ymxfa2SC+tcF2+wf5mZQV0U5mVNmhFvriETpP7IwYanNg773xQeoys
RUcxCtVGW3FCl2at1E9B4QI2FXpuFxV1ZJdYjj1KesyhaeYPVPc3b/JTz6+Nx68V18e8TPHjXSEc
K6QEsFlO6jyTMoDZDQJn1AT+VWf4ICezf1nJ17j1ZfEEP0GqISnyO8AWqmAjAMb2RMJYK6LO6o2Q
n68mhaGv/wfi7aQr55dhuJW94UULn3SL5wUtiS3QYc3II8DmF0j9+3S4fhKED6M7OisCryoQHd8C
SuwndOz24KAFsZjDPaTZUG5wNZxlGoZ0X27YTg1Vw1mCWujz2H3Q93/QaVI1AgRa/owHgvGrhvr7
ONsDq4QKq7NdqMn9UiT1jB7iJTab3ELWyqesu+N+O190uDJZ/2sdbQZVWEnvPtDb3nRVSYB8m5AF
OEahFwgnzwtBBem+TWtlkO+j/qZNcNSfJgYHCD4QHYhd4JrETYwJkA9c36u7S2axr8um4TImdJ73
IlDknmUo8HVaunmRpg0meFto0tbQo3oEDT8d8bJgujzu8nQoPCuNW2IM8sn4/bC4QVGqf2H6qc7Q
n4rlqiVKaWg9HjQ9dotxCecOHAapCs0ON1MyrlJnq27r+cGcoOZksL94nkRftWSbfm8IC5k2eO6C
nissGp5cuhYoSMIMQD82mtk2d0ly/deRfYxj3F6x8va3KdLQb9D8eoY+xVMdcOqoaCWsuvYoPwcg
hLN9DXq6DuZQdppo8IWiDXao2lTE3uhRXe+iqaNajohvM9azs4yiBEsMp1tGbH3JFz7fbWO6QdRy
o4doFycqUWjH3q0/tdy3yRVRCA96nAc4sTLxUARIuxGVs4oR6k9MXEYoGv95sjGQlRbdCP4OAVU5
tCqkDbBwNbsCRTrSsInbhQaORQDgAhoHuy1ANmEGjAZTUhtHw4KuC10tlyc2zzUHfwIdiIE4Cr/s
Z3ogIZEfKcAKU+WFInXZjVBLUamsaq3sXa4YnRN9Irpqyk57m+ez2wBgRERYdKVc5v+VyHCMg+XE
7Vl2v9VZhqg8CGk0TPm72FyqrctAuoP8esPzRTblrZoUIfOEpo0oXw+ouozzcSWAXWy7keOVqWvJ
DqdE912gRjnrFoWkr2OoOSKtIR2yP3cyLDhbVkTkZB8LMVxY/wCLCi2TvxFlEHOQN9yxcbRqeaaZ
HO63hRgRozdTTu/PhihYtWnAiVIWDOB3N6NPrCpZ7THjHyAsENCivIwewjYD557VwboSzUi23MRu
XC0cZVaIKctyDmlRX4+lnLBJWrAJeof4XIfICrRBFJT06PkRWkeJPbbj3SzTbCRhaIx21q+B4W50
ghhRcc/xyvjbiIOlOwM6hp2+NvXE3N/PiMZRaOCBQv9JnUJZy3abRRby4B2PSWTTUdItnnIpubES
F95NIDd3vcf0HfUJ/C5w4rjTPub/EG8BBNgcA6Bk4BoBWY2zhItwi72G218tJBiS8n9VcMwI1MER
psQOx2l37QEE5YngB9EQt/nw/GqD7c1NUckV4yHSYeJrzhPPFHM+98mysenksIQTid1JGyVhGVuD
FTP+Dkn4eOxJddRque913U8MfAy0sKShE8Rp5QxXOAssl8ul2pQRRq1+gaC22TMHPNAsT0vietx1
YVousgRkZtHKZSH/aBeTyiy3vo9eHwrVL24uILRG2OABWT1PiCDfJDPnzZZhRXe6oNHdkPjBoZ8Y
aCIWBj1oFrzn/N2tnRxApZpaJRIclxjWR/zAxqYsaMW9hLtxuK9YLVW9rthiWsRSN1xjSwxU2lro
mZzx7Xt0b/gmNsQ318uSh6b7jb38ThV2dKZq0h6HbcraA+Q/LWkNwiREtGPaLJ78D3Ro6ufnI1mN
Y+8JUJz2CAqXDw7PDrJs6vDZm/SgCSvx4pcwsMPzM5gN2U30ou9karesYiQPLyf8WvGLYXPbnJEz
0tLWNz5HTkincdsj5iK5IkodFzqMYm+disZd7TfM2r6bHR6LP9Ng29r7eOeKhwfMSokq3a+L6l8r
aEYnaklupsfH0OPEM5gG+AdEBbvJ/fTz0nS6TjVMv5N0QzUIJz0/IZgRJy/+Afep/yvNpMlGP7gD
G5+wQvqc0qGprPy7AVJ9Gfk32EZ++OdlBg/G2U52txU3OMsGHv8+L4G6rtwo30l32Kfz78A1lN/a
ky5dxuksbJOt5fHqcKRkWWmfOrH4ihHhz79tVn+xqh7tRcprO/WXY28zOvTzEjJPSgfHI+TpjPHK
U9aJnLJeLzqE6LOX6+CKzB7AiXBkhyAjHrKcynhmW8E75UntEPyTTQ1JwQY8Xv3vFiRUSS47bq9p
NY5k9GeelKDd2jnKoPH+hnZdooJYruhaptfTrcm0WUHexYLxpKUoaXhik8M9DXqg7Gm33Y3gY2RS
sNLP5RT3VrZh6Pzgx5xKSVY/cPKnMRtMu2mCVUSSdmNtZ3NyEk38FQLra/ScYSQaZigBtO170wX7
OfCvAvGGPxLpfwXR2rxsp7wjuMLSDavYEy5XHqXMSiRMiITjxjOcYtpPae/+m8qFYwjEwodUPBNG
AHwRypBkZCEFemttTHA1J1melFR0fqubeIZb9TYb/eduRavoKWcKbH5x7ybuVS+KtdZizDvclxEK
Te11yBEAVmrHla9DyL3J9abjZFJiczvkbXg60bZecM1oG13a5b5gk6WdooKT3RINSRTlxRqyzK50
uBmzYUgCRyI6PViV47AApu0D+6pjqLSI/dwMWHsShkQYW9lzsHvSf8jkDrcPofrRh0UYuVcUeyOI
PIVeGd+BGTWboSSndnVGvZz2T+OgREOMjsrsFAv7uc5lbEmAID/2xdOK5SSIG6LYPL6V5h37E3+5
N15+aKpgNlQYeVoOfSkE0hckeOa4jYLKRBkai7MCWLVf2LqC8ePHIPrvsOBC8sFI3iFSXVa3vMca
cwwcN8ohGbxvpAWOWV8tOF/NJMxH7ZgLxPx1tkUYyXEyoeTrmpM4KxhDkhAzwDwM2bFWeGfUFTDq
qS7KL5FGTj2HItzyGLhFor6FZcD0v259w+MiWwAGSsxinUCf+Mqu+CLN3xjuWQ393AFum2qWRuEn
/kcp+Afnr4UQ8rMgLJGe7/x+1wjQcfDtPSYEz1XxNjox+4FINeh2ksjOs7dhXBk2JZqiakqM8LwQ
6+RYL2Tlnclej76GxxRE4VpbO1DTotoTwRc+OzrleTBaGR+OwuExcHwMcdxiQ4VA3qBSqc8Znn40
SHihf0NDNDvl3mQ6AZRHIsGnziAQIs3xhNHFdQAIj0a2HvXDsh4m0YktDG6ymhOprZhxupzC1AKt
YuVA224/bqQWXLs3+yrSYGUIveDU8JVKXwE7oCPgz51otiZyLOSrX/67ADRxsFKLGHtID5th/sjk
01N2am7Sn8zaA4XPvW1AZViDDFPMakXJvxR5z5NiED/N+f7oFjFwmKW0XYdglSJgaOWfw7awJUHa
dEzwsdHhgXEiRx8kAwQoT8etxSPjArXLI11AEHbAurST2QtinSAft4S264ERzY8W6dJt6Kbj/Qtx
X4tYAGKWTUqlIFQdU88LaD2Kd1YaOKLbZ7j98Av3Mh4udPE0uFQLip/Fk7QI5C+KU1XEqZRLlmc2
BfMaDc74Q9oRImkLYTkEBZXUi0k8NDCt9PkzMmKqpsd8D08VrRCDZJgOx4GH2LfUjqJG45HALlVU
+9aPY34ScFnVme2h6thEpEIHpGYnGF56LCa0mCOLUaAadIXt3fNwMwtU+hY2bAQpBGovDDnYOlqV
0ub8snaM1b2Es41dnOUVM9HIms1Iy6ndyQt+jrHLu/b2zgaWfHd/L24KBPINH+rp7Njgwk4yEUeA
5P70nfTRVAa4utfEKXqHL4uRcQtaLhouXOem2JTtjptQu30OkJizYawEyWH1Z195mCwng+EfMotr
6BetdAms/TUOqqVgf2xJa0T25dpiXKJejV0X9b10g7UZoFl4wYGSGM7x207LECbxkOdzpZkWFAiX
S5zmRwqW1H27hGJiCsRsX/P22SoppqknbWZvIsid51iyOUjsUze2twE1AP3ToLrA9+X/G78nfemh
aWPaqdFnfB8NdRMr97rwznwoUbl4NNrUNoUj3yeazXF5QJN1261wkIiB1z+COhiRnU3JSRhkVVFR
vSGoZmXBfpbqd8P8463m8fGNavpXEVKRp+ERK6NwOQ//yRb7DxFjQbrlcHWp734n3jvRQwQSadVm
6pOTBKQEWij84pEp+1FMkgHMrzOfuUTg3wFXyMulB72oRFJ65xJ6sjZOlydtLy08UDPE3V7s7mpF
vohm8WiIC3y6WrHH1bzudy5bcNzKATqtKynETh3oCjJCwH3E9BFQFLrJ2fVcFOqHShjHYa5AMLEX
vcpdiDvzUzvaag/VIKKBREdApgYF3AHHVwyBEyateuSqF2z3N+rUZZmMwglnZ9PMLHxo924mwTuA
uk5ly1KhwBjh2BLkvzh9lMnjsbhwQ2RyHbKY3ShtmpCKl5nXEq0isv+IAky1KLpulM3murTD+6/K
Jugx6hwKUpObjrWwHFXY7OFzz7zv4II5PD9+6fGQaiASyWR6bMo0aS8y+lyknYAANXA3M3P+0mJl
jn1LAw3/hwrppqWxPkhxLh5XtE/BOV86zxu/EfL3de7K6ggSZFgLspcSC3ch5XHLNnnUiFP5r1YS
m15PHl0zOHz1HJHxnSaq3u2/zNvpkvK7p/EISqLg5uuSKWKTzZYPxB5RCeG2AewhSyBhSNVPGc/w
eFpIpqCLBGM/Cld+bcPMCosnVSPUfj5Sn2xSUDXHoi3Nr+2BCRmG/L7Iqo7HYQx5A3fbr1Gvtydx
nruJyIhlrTRL3m5Iwcu5uUo0dBvRPC3YmXXoSHdL4MSzFOaBQdoyLnXi6IXYCAj2qEH4/KmFhTI3
GYH0U2C1f6AVL3y0MgVvBP8OTLCtUZUqTARIjr/kLXQ4nr3/pf38/7WvFlRKBxxCpd1+izSXaR1V
YelwU/AGpsb76Vzkgt/iNsfS6TfUFayeLv+HdKYjSCJb/rpszkK/e0AGvDUuNBHTcp7MIIyd/oWg
quDHeE3RRSF7LCO81j+zQ5dxgqUF5o0Un4TPdvrfJtf8bBr8UHhJfaPr2Gu4VWXM9xoC144/Xy1S
s/ZX8yUZL4BwZ4yuYjChugnY6+7UA9XbBtgXKNXsDXZqumLidb1gFxjvdmV0FyUM0HkUK+mbIs/b
fP5jhQa/gtHcwOWzqM8jCTphYACJ6r78/8ZHAKB+pythnyWHUrhGH54LXHI1X7M2I+KO2ifEkj6B
mD1YS7kMdwTYsO9Sxz0oIuF4I1rQIFNf+TndFdC+1L82tU5X/dHcXgv6L8lqSplKmdNJBLQc6wA2
b5Xlx8SlvjsJdKrQpWAEKxVa4dA1Wp8GSrDCyHk3ixSTpXHB55y2kFqsEfCumnb9cWYxbrOhwDVb
a3FULGZckhCXs4vNI0z/LSgYcdm1x3FyV1nShJ1u4FtHHsMvtQqb627c0OkPutDUNTdpAFqH4HNP
BS8JR6H3J8g6CAlMpzX1A+IPnzXk9d+fF7pPXIBaOr8sGdGmwXtKFpJgn0GBBrBzihUccLn1Gm6M
hPXf6fp9aIfwjfYzR+mnqtWVteva0v51+SHWa2rcljBrqzImER9R6FOJyi/bG4/dJYoWyH/hJF2r
BnFVDCvC7igcDlkNRRMYKigQr7DUJerslO8JbsqCzBS8adNx74bDa1uWTexJKYL+Ov66ANFHQlwA
r8BVEtu8/MKCs9hf22pbgX5k/Ij9UJwapQBPtkPJmAsrvBu2dVjGh14l7Xrd0bK1lWxSn7VjuTdi
QokuqTHfZK5nryIwwKngCcKOQH71spu2VCZ1VI0aVfIY3FcnTSeETrmkThD4U6rq3a7I8czYnDH5
1aGjzZbEtABDIF6jDpfl9/75xDwL0i96neexBaS6DuwE5j/zpvQZsB1qgGCCqkFOvR3B8EfRQcAC
mNTpp5zWHf+9RTMxwv5mIuzQPAd3QoEO570nsXgP2Ahc7v2baUioyoRa6KimsTNudOG5YHem0cUa
9Pq4eAV+9jP3tkmA871u07X4vc01YpyuczTLWuMhjhnzHaUUKfB5h2JFElunUq7uf9JFMLCwT4Lx
8mzD3wiQdVml9zJ2VASGzga1Rad+5Q0oq081fWsKjY+qCRQ8UEXB8Fd3Jckyaz3GcE/bn8GRbj37
LNaO808Bt4u9k+OVI6OVAZ7ZnbPaQYvtNCUaeHAyQ372XzFP0TJk/3SzhDSN5qaN7zsgi/n9SNg8
9IF/ZwhVZqP/zMGibFkQQQa64xMaURG1aeJIytbYtJlUmWNaUJa4g9qyz4jUdilzCTtFtIbJF8Jq
G0aQrLN8VCRf6u2QXlft8/z1VUfZy5QOYJn7Li73NB4acaxd20mkLKl13bPFA9MkE6drpmaQ9arT
1/oPaRZ0NTX14i2qZ4kBJgRw7flRidWYxqPIgsU0W4xlVCCHsyQi2gmu8iyhjHFjxn5UtbKL89+X
6I1xT144dXNsrMEUGeH1V6+jZL4l7khg3HPkfMjKq/qL9PGkWEm8mfXxbpq5N/P1uVpm5w2mrFoT
e9aEJEFblzdM6/oIB63fwgWLuEzJGr/JBNtIaJz5FjIJwkEb5lswhW/tR6qf2uRoPji6004Vsj/s
70VpSkbZOMuR0FGJC6qco5w8XwIEmahQE8nHZ5tJzi6lk3AjbTh5IHzcHlxOeSErBVw5fQw3xz/Y
QWa7Z6DTsHGYTA5oFMcZkGkd9D9enedV04gIQMazw16E6IB1PQyx5+Hl2yWB4JmiK+o4gXCkz2Vl
TFm+m5ial9tWqiudcrvgg1LxzAzo2hKdEV3yPewry89KLOeyoLR5JvphNTo7ibODkPqvXs5uCZXW
zkAbhH8dVgUFTni3L4aP+bNnfhDfe9srA+rkL3jOPfBXrZMDwBTAcmZac8W+p1gA0crCQHcclxh7
EMx2prAhhoyvPzU17S1yFhGALAR5OKKbc+RCzAKru4uabgZeEf4cIoltTBFt5Rppjqb+Ov0a988i
xvChaOlEFoBeIS4dd5vC6/4UyxnMGDKik/HAy5W7/Zw+1O6zYWRDPzE6rKBMViW7aFoVHPx9zulI
r5mUSo2fgXLiE1fLTLRpoBO5NdKAc0vlskM3MC5rKVl+AG/Ah05EVftsU1Y7hYhlEpccJdhNiark
JopSvjh3kQiMzVu/BAAvI5IiKdV2bB4+rmq16xQgt2K9zf5eI0nPckjWVGaVgEpnOG1F9zFb1Bby
PXqOmeDnP94taOWKcClDRgZ7ieYxghlKMqotekiEHP2GNeMV4W8y7wqVxazkTV/TL0lQdVb42nFj
fra5a+5ISpIi1gZTk82c6iTt/fL7nlfL0hCn8nm7azkIgpWF8c7bDq5HO+ISA11fTe2HRPz2lCVj
D57ZCaBZBzxIkv4gB4OQdl1iLO8qWX08eBXYlM4Oz6AS7rtzw15kxB4aa0wcL8ChYpIMBt/jfY4a
pAYCnay0KEAmh2TXzBT9leH25o6HAJv7XpguBZ+trLltP2027MNdJAIgkWfxbveqhqvh2x7s+VkP
IdciBtXiKSx5kZL/oAhvXiy0zq3j/ENP9BF9Zjxx8SvkAci6V76YE1RX13ozWF1f/w3COuR12P9D
DQCKK1H6aB41mn2hiws8nyhPYl+HoLNJXuksUnl3M4yAPNcXvpPKHnW4hHfyM9FGGiTxot6GUFFb
x3wV0LZlq8C4g/pziMQnR5DspPlaP1ZSAwHqHlWBdAqP7zplWypxrTZqJL9VuO9z+EwlxIsSo49M
3PE0HaB+RmNbBIuLVBx3mKl0u3TFo4PnZkV5JDncWbvntZZes+Dh8A1NxCgDmKZdzyZYO4OdNZfI
9x2wqP1hHkGLZ4ndsDWwQGv7MRrgtCmN2AUxN6byjsvOWccavkjBCg3u3l+R5nY55r9EAaVHE/0D
NCPKY9TgkXQxDGjMQAOfLpCTeEUZGIiCWxxwHgNkN71h8suEkBKYuRxs8Q3bxJELAaaN1RfH3k30
7XISfK0HbdczJseUyXOlfcUJ99+Qo0GrphnmGDS3KPTJvRhergxF4zVi9bhzc5Lca0A0Z6CmDW/3
4AsAn/NZw3olvt11X+4MU5MqHslRrPL81accAmqspdEnnC6qel4/9VHGNnUS7XuhG3c8U96rJ6yX
ElmGFbrE0xddZbaWGtCck9wKxaxjG4ARFJ5t1g9wJPk3Wb/tfd4xguwx0dL3TVPRYKbRq0Fjpx5w
5h0S8AKXSUvAOP3jyY2DL9oqUcbDVbRii46C6uqiy5j6E77ozjpg1akpLXxPDnOHXvLXR2Jisxdg
UZWBMz9VwLrIhOCWoXGa0Md1tIA8tyG/I3XqarJiM9/9MgRoB/Au3C8IKSCn8nZjAiLOcto5cNH7
zUZjQHq8sq4xdjB2gvZTaYtSsWUWuOI/niF1LmYYEZS4LdnPNknV5828jecJEDvjxPaij1jn4rtj
vXvoyv6CEIHutIaZaYCpbXtGEOsbivHzfgBaWtAtthPL73d1iyht/FcDgJdeiO8Ql+dFR9Ov54Jy
VrujQyagHf6xYQjFzwUwuFjdrl+8q2EujT0RN0QXlQU9A2MdkeIKapHUSEutA9hjpNws8eXmxA8F
6BIsiTzzKu/zxyzXdAoWD/7IxMsO/Qj5n2bUVmFGYQhPgpCca6KrXmuK6ZRfoluV2OkEc3LTOmDU
xYvRIYD62RthJVveJiG5/Z1YRfU3MoH+8vR38kJZhQggVCaIWS4W5DoIbpi6Axbqmoj8rZwT4sa8
RQyCuIU7fPENAPn+dHox8Ejeed3FRk+VVS7Hj+jsD8b8EXGC/3Rbap562qWuXgSz1hgruI6z2T3W
mDshB1tlJvdCNXHb7ckRTZ2MdtuXZsHPLgMD1Kxpp0FbHoFK9mLfi6hfcCuZML+sJ2L5Iwx/xHMY
sF4iVk4OZlBtrtGjHkpmL4xvzPZ+7FqqscJYP5yJks5PfJTZj4jH7b+5xeZyXpXlK925ZsSTK5Wx
rrYzrpV/c82fPgfRmJPwE44UQolRDz84fgPpl30r2w8BJxhDo0MLV72OpZZXf6PJX8G/qu4K45f5
ytb1dObF17YMggh6J+zQ1WWSmA8WMJvVwxXHUC1g7aDcGMWC412+7MtennxPJH93BiQ5Vq8YwB5s
7d4ox+KRk4zrZ6tDIkAT+uw1hprk3j+501+JYxwdJli5+lyF//PLWUyCmNHpNzvLtCaeezcb7hOp
Eb24OgN5APCi3BeOchA7yBxIAku3DoesAU6kXCzRjFu0I1axP//oa6K2nAtDe0Fe3Wy38+Tllcsy
+Li+PgkiXyxUSofNgOdgq1bS84q4QvE9fQCPq4aPzA6doVpG84TPBU9ksbvl7hZ/xmDVaHUm1Q0I
ymYE90MEgfdCHDW8Y3EkjD75i0I46EK/H30xU7wcbuRzs7sTQ9TniTMG5Or2jjttXr5rqKIMzt83
NpU5T66CTUY7s5s11K9Qfto+8ODA594tuBzy9GATYj87+3qSkh4d/y9+nfSQRoCUhWj/dzHXJWXW
JytAQxG1aeBS+bxxWeWl4k7ftMLMoyafQqt8uJMuo1hLJxd6OMkC6/Pk4ETLdbbKgqMQtwzit4p+
n4Wa+2qfocFKhfXlgwFIGBZWrzerEJqpHHXLP5x39fP2xXEdAMVB7pRN+ywPI7gRRbmsJMuQ1cco
L+PcExvkFBaFEBbLh1/gq+LFxWGRW7HBpDfI5G5sN04QyW7yjPwH70W5OZ7V/5oLa8AC0YiLlHWk
j+hhPpvEpxgTvLpgZFrZ/BDFhqeDoQAhCEE73r7s0hr6zdeCU03ckScNhH9apJdrOZJV4XHprO6m
VZPL081Yy4l/SGZNioy8lv448rG73Ro1SHbDzLQeGzBDoLkHz+CkhzLjiW+D074tQrvL3EwRjiAy
IfYKUQfMce1/L++dSswyV7rYuqqd3KuVKXTd9uo05EiP01hiM2SxkZL0mal4W7BLXwdFSWuG5TFw
RpDmSRTgtK9aSwJJ8X+0yrFLZBMxu78cXhts7mm+TI7g05vCvgrhUShSM6vL1wHLP+qLU3sC7XM3
85IoQGAiAnnV9v5nJ1/J5WFbffVvBTxpPyYGzrADHNfju6LHY1k7RvyRR6tf2zJUQmQaeKhf87D+
xd3ioJ8YxVonSbGU7zjIu3FZibElY4ahMazH82jlOSDReIJZHs7mCbinXnZ2mFqwH84+DLmp6Je4
VROSYywe3UnOob7L1AAh1TPn+f+RYMIyVi6pH1p7XmO1vMvk2mHfBA1OYXkUlPJPaEpPmyBJOuVR
nHU3E5gTA4yUHER0giwnXHExzxrJNBtauHAwwKi5b67kDVXgb7+8ijQ51C65YPGj+xj7rKtkMHMe
gelvl+3rsu9fVhnLjMvWT/mQXmd9WbfCYH+ue7sVzjDdDu5zDj8CP271oUdbup9HUTLgdFW5jfjt
InrxDe1fSOfuBaN9oANyZ1KiZvOZ7fuiW0Z0jjRKXz/ISIkyT70moGcIQ3vd2cCNIDuO5SYHlna0
1JkQLb66Ro0kTHNuDWQSB1fLPNmAvTzbWxHA/L+toj7/bSaVjzzjDksCnNcBDqbVzKBe+lh0c7Mg
pcyWKJqUWXqNN5NBcjSpAddWjbBb0xCoFS/aU6235glMNCwus8If8PK7siRFWGZNEQd8Bi98L0is
B1PAmtHX4kVWiQyB+LA7l/eviZe4qfAkzot+9PRrWkclxFBoTrSOOFLS1zJn9js8GQtG7EZo8J5k
YSsltt2Ht0Ab6S9NdGXT9xT2evRxZGVP/jnuGeyKEZh3OX8rACMBcMmqsl3SnR2cckvikO+GGUu5
g00r9pg7tr2kJZPAMW5jRDrrmto32W8rf9BX/xbJ6oIPOSSc46j6/YY4sRRi2REuTexbblCaZLlI
rNEtVlbSl5b12zIUWxkIEPSKyoycywZykShefPFnb37Hn5agzAnVOlVNzQbUxu/PTSmjyNdZYXb6
cBeD/6lik2tW6FCIi6lehlOD0u5dEgTNbCpABzxj57pZqDYdWwFDTI1XawBPssM1bI75hNCy4nb9
qlmikdZtrZFlSAglaH0153LZiQ7wrW54H3vmRyEJPdq7FTSrc+n8G5XK7T/Kiq0yHyz2xaZSZ6KB
37ThS/wC70N6YqF8YD1Laj24tmzw2IZ7hQrDm/ZyPGW4FF1w5IK0T/Q8OSMmLn6mhVUc4aj907N5
GDYm0Rmk3FRJq1xvo3W8FylaDWtrGoce53u1Bxuog+PcEr2A8fBdYaqZPRftdxfEuPTuS8NVD69m
N8VPnJvONEV03vQjmfD7EpxGCLF+Qeo9KZPtQfMeBGoovLXcn58Ue7MLkmmuqYa3c+Xpf7cB6SZi
bCRufC0tLQ/WbHze4PI+iaCCNrwGiGt2Xs+pYX44kDW1jZQkCX+S3R/fG5Zfy5MmUXY/nvcKYhpS
pfuoEvvHIBlQQH6Ne5CZwbvURsW9NV6Euh+kTk2p5RDVHs8HAqizaL64BQmOgkbtGQxmDx7xRQxq
HT5hVdl/oOaA5mP7R4cIgpm4pUI4DYKRqbfbfn69oZJ8o9xAesP17VoGIL2tvfHv7Qp6NvneKPej
T0HC6yOxNTDrndaj4MfvwdCTeEIJdxAdBhOzKLlY1BKI4JdJ+WsItEPcwOdn1auuxkwddnqQx0je
0WwRkRB5nahwcbuBYp+6gW1DiQD6XB8e9v2tn6Ni77wRJEavPsjn5rErIKno5ptvjH+P00peGP1j
tYgeYTl+ngaGf+hDZHb4Xhr4R9o9JoMQRHH5n/TgWTbVCuQqHejjvtRXoizB+JHO/XWUNjLMiLfY
ft4FHWe3EbOGSkDoDWGydra8uEwUYQq3l0xBbtbyaYRmKRWqdVWgDnH8MalAXhuYUI12GylTN60W
B6kKUVdgZUvG9TqkT9d3YRZ86Qm3yszsIRHJoXWYg9GpDb3REUdv11p7pazsbtcCWNBdJf48YEom
/v9VuQludWtwcYXDRR8HIXvE9sWp2OPaw7og9hymapQLDN5MQTbpno+gmP0v23oxzGYZZyZfHVx1
IcB2BN8NY4S5pd6QA9LXJjf6gUtKDjJFrvOsuRCuTvqAvqrG4GvZ8RUlk//orN84UOnI/Gj0Cqfl
xuvyHzZPXZmeHOSOxVUIgfepTNXNGdD/WY9zKVTDYOVPw3ZFTgCX7EkmcfEv2FrCMFeGi2aTGXXK
5IE1PdkVtmnR2B9yAMX7te5PF9ptKK17EeSD9q+/sTXqUOR028FEZJnNoJcLSI52m8XYWpHFdosm
Ze1U8Cm5pZbNJv/yggzMva3B7s+r2YswP2BYqY6wI9nYTJN1lm74kyYm0ku8YXAigc/4Pwhr5AKy
Y1LkTHHBOSe/4csc6/u7sHFxlHLUyc8ElVr5twzoYdACRYHYlDAedyhmDTjE/FrxUpnXL5RQsELo
G57zzo3vp7OUi+pGGbkxOJVKqejYWFrr5E4e51PQagke9TctKs+lICrhNJhb5fztiK1/iQUkI+66
6bamKGx2/l/PqXduAxEMjqROnt67ir4dLK5vL7UqWz/VbwnWWFulYsn+Xjjy+gqhtpJyZX/i1lPr
4MhRj0/7Fb9oGRPv+V+nRXW2S8ztMcXZBjDCqNtfF+dgg7fiqFfUK8kySA8eUJoyaIa+r+L9PpB0
lSH5FY4yOuu28OXBl7r6CQlxroVRG94OMmEKbO7rsyWdLPTqUlvpS96gV7lKoTCDcEG8+gC0jAAC
tHrYURzPmiGkPVoTQODKzNtMPc4b+O6HwS5UHzsR6ALJo0+JaGAWq5ighQN1YtZVIwTVIRkUemiM
2Yg2CPMcyzIKqVZHG/uCJvPJaSfIwZtE1vVOXdumZ1rnB5UWc4LTjOdF+2I27ju2ubZToxkmgH1f
j2Nb9wxRNHxHtCvFIKfycFeYqauggkn37dmAzoUlTDjgufGaOyEZ15BxDETiIrUHrjkcHuuM1vOJ
ShDkTN+WR3zhJ0DAWBUEtRzTU76a/ij6dPvgJAWp+nu+qXi6UDbt82bCQrNZ1o2rZBeZ5WyV9HC6
deOgvT4yJCARVIJSL4I0V30QLZNq0nLAKEs4eW/3f1qXKemj0GGl8rJSshxFKKrKePEHbqpI4ZRc
+7e3pv/9REBorTChYS/Bgf5Wf2ytz5D6JSF8WrnnJNLdUHyIJKP4orf0I/KEYM5I/Bhc736733fc
UTwEGKbBvFMjK7UYZ29n9Yu3/TS0ytuXzKcK7h9745PF68B2nWSqBbzkyWD4/i5z/iJ946CM37G/
EGbt2ZrLoL3/nX63i3KfgxapNMZZq4S8P7BKS0ju25zGhzkVGCusRLJBlFkA8+rXhIywIugIM/DP
/7JnujLdeebcUKz8X88UPYrWueCK0CYvbH6fSeD09xApueRlcjn3exTTHFaoMeE2hjuBiadlb7Ey
75OeitWkPLmJwiUH61SojYtYlNtLhZEDgXLme4lLd1hc/55qtrN9ouCNgm0xePHWYk/0w3RWxr08
6enrwOfuKMQtdylu/Lvk1EVPveDSvRoXBqZUHkReb7ehsjcHPv8JYu9bxOqiPOH/aawbaVXgseud
PuXkYeVPxGHBGrCvXFV1UeeZ624Zr9BCyNLdV+/OhnOJ3H7L/MoEKgOe9NjnfbnMF3Vht1povOkS
MHpkdnUPIpG1TWAJ06lNm1/+3lULZNouFvmhiB+rD7HIpCVe/sXg6GihuZfu6vSxnPNppTTBMHs2
eTVrS+JHJLxfTunBoXIIKqhlNZm6OfEP7VzGdI5wuI1FbnMAyAEZEG87q5al3hyKHiacO5vJKUZL
rr6m1Bl9jChTjGobihsohG5nMAfmSFHJeZzL+2/ivA307TJ5XrYhsMdWHsKyVosjF6oo5ClWAIsI
dVev9QmttwWo/6UYQieeiK2AXZicmQOAOdW3FGQvb8rKOCJjcnVYq9NzKOXHyOEoizkD8R1PNgWg
Tbz9G61VDE64+NAS4SIepFM+QrFIHe4EugNs9QGxErd5nySgidJNiagywG4SQKshn4f5q7BEVuGz
7e3f67EraO4tKT+e0PMPkliErMjLZsiSJ31KhHWya/ESBMrZy1Xhkf0HmczXuSDUISUUhWhEFH15
NpnC1R2llXZMgBZw+wsJzu8qwTfEYLM/uzKyTLFcJqBzkK4Vw53xcxL2Yb6ZFkde5WzAdSAccmgk
xcZQpk2anWLVJHtL9fJXjkTxpC0eY+7yn4u34DECKZI7e/DmZSvlfyOlNClbGV9tJoB+imk8i7j/
GCLSUTZN9z7eWaqMlPcdkYgWQyf5/FaS+YMGcrccCqun1Be9/s5KxGzzmMwTjz6IK+bFcG4VvTHK
YKwfEmuHAta46GxxvTV73DG3prp6bVniDtXTD9NeNqQ7z2EouCC4nxbMvf3GzEuaEUFNXH6lRpVW
kQTxuDH6pUSWvT+KyvRRz8rN+c+S9R75lTW5K3PND/U9d3PyFy4Rv62W+iSb1nCpDOFaludeJLVK
kbtygPSSbbVL5pGaAzYtb5ArgHX+ZpjMNlDTgx8jZxyp77AHaA/P/pg2UGU5obFI83Zk7v0MftET
Ruso2sh8HTLoZhrB4tZskfu4yrIYzq5+rVakNS38suSKAC9VOF4za2nh9aEIfcHGr7JAq383ZZSk
G2qP4RBe9qAi/9j9wryiq672qDugg7+CxGc5mU5E7VZQNCi6sk4G0tAqBXieFwfMmjHvoAjcpdK2
eDTNngLhE3VoQ5lnHfnNWAmePSNWyFys+RaSJBy9Cxvq7V/bbiz1tVlE8ZGqVjMJJ/N3L6W5jkDt
Rh7j+1BJF6xy3FBPuNlF7qndN5IzJR+AlcfURiy8ywKFq1tB+gxsaKMocIW1iVT6I/DR/tvd0rLl
mGzkYi3X0ZvBgW5w5HjgXxD9JbLn7mknQ9CYjBOQpmV+NUDL6rB3rIRntBTyuOcOTAF6zgmUaVIJ
+UMTqxQIZ0tGQbrAhLJ7nVlgScY86NlTlb1Df+V6LO+qja7R5n+CRfEKk+1XhjQoZZhl3FSRcI1b
y8SxtoHDqyudqWUrHOrB5vL4nCmYAOGtRN/pUW7tH8vb7rMxr+F0gfXnoDBJ7exuabYPBdc9+5je
oy0XlfUxILOU8tqznV++foUbk2t3oJgt/v5UjVzmP6sA6UK+ygRjKf4tp7jmwrcxSZ8MbqyyG93t
QsU75QyGrRizK7qUNCWPojPuO3RA2De15AhpFpjyOG7R5QoYe48ph2DfVCsN88MTuuJhAEzOaik2
pQURXKW/Ikiseoca4JxsY1hU3k8zXrLLj1S9mqEWPUEZAzGhGQST6uqLD+prosM2/QWwIR/BtJSY
DF+cp/xNrepJ21Zpc6t6GMfZOKJlmBZtEOvxTHIEvRy29pi09l8cdlE9KWz+serVqNy9S6Ot8Btf
9HvPbQrrCBPt0QOI2OXkSetCeVx0V8oLMkEwY/R5cl+dK37pxeo41sRAMGE9OyrD2MMvt6MWe9U7
KkRcKUJ6NScjrILv9aMRJ/L/6zIAP4X69luAsD7iQbk4hoPMYj+/JIhsvA3a+9cNY5GslzMI+emC
rC80H3vKypqei0Vyt9YE7HIf2S2MxTznklc13/YHpHgezJgtCoZbTl2CNb+cxxgi0aa5X9iyR04J
LBz2uopIeku09LA8BhNWRQrw6IgZCwpjBPeGXx3xLf/Ph2oFEkx5ploSiQCvcWFZuYcCs3DHaaOo
0LT1YcJgNwX0WU1SSPrgWPJRcfCbcZ97AiMrk0wXDIuCAG7jX6csv9yiQxiS8y2XMI6i07E/q38V
Bw17W3ZK1LqX9FJqBj8B1xuHUvm7nHJswR9k5yWc+ZSaVckd4NX81XukeRqhYAz6CkMrJ/kC3asW
A8Y65B2QHMM9NrsKn0pk3F6F+9LBGLf3xJR8f3VnyHTtPZ1kARjJsE2PvnjvCyUvGPGWpVxCA88L
5j36/m53BS948EHGKGy59NC/frfBE5zMEcyskKY1RBhoJKozm5QoRncB0EkyG2WiUoR68s0kBeBC
AuZwHvPWr8dLwcKc88kFgUA7TzhUnT8OPgs/iE3RZ3etiU6YLFqyi/jf3/XSU3Z3vRBBJ/xkfbPF
4lq/Uv3KGXlGrnlNMVCKTDbGCUs+4oxok6SjmU8ikqntS2lqjmGSaOwg6yCUbDPRisepDIhT/UFH
g291y5ZEemi8A649rW2Qf3UAYwfc6/EGBylX6maLsWFPcCXY0HgSeCQpx6LWyh2+IozXhODvCU4B
2FKGnOvrcddVICvKPZu0iXYpNHJO6PdEvnn5CbYKXlOfu7Qc5FyR8xALGdpxBr902yq8FmyQfenN
ssMBs+e6mHrb1bmg72jRogwTqshekVs9IYwMA5bbS/HhWNtGUU7Qg4vU8I5AzhvSTqEo33TYg3EZ
esJpqGG975vEACQA/hhRj63pAtAo/Byk7uMqF45jcJwOki+CfvXSlng8PA2gzG2Pbe+fpSs7pz5k
jEhyiQyRuUlOLoZAtfZNpejON3udNsKv9A/Xf18jD0dQbjf17t//TIoiE7M0eEJfBk7qtE5osIsM
fvQA6H44WLv4Is3q4ytFG/YWAsreTcDhfWO1Mypi+L1e2siEgNKGaW+t8V+abVr+GNgzI5lmeE7p
x+y1EbOX8yvz467Qu7K51jjPy1mcfwTPMKPmQHTkp20J8Qt4aEVz2MsDpfGr1TyQGYQ7ikrl1qjA
fQfKwkJ9x6lMHV45de45OG4TYApRQSA68/8EgJEl1Fwpd+Iv/vMbQtw4IDTAoO+kChdrvdaby5u3
aMF0NMRmTigk056aAQ1jpSmxTJaGNqTUcj2nXW3AXMnFBBryplCL2u8azSeiOiMtXPYg3V6xuiBL
RBZjM1BWGMArwVwEO5kH5zC4ANmW/Wa39ntTa5HqRzykGiePVQWds2Jgah4lsElqoG9z64K+CWJ+
9RtdDg6DxA8Wl2tDCEOqNiuw21jTmvuwN3ZsO2yB+94db5iT47DOwaaIo/wLogbGfxDAUxXKdJ1v
bHrZiIX7aACjCAjk8Gwj+nFiWmZ/tftiRfoZdN1OPW5cS27OdF+/l8fg5F1TFLvYXELWvStfxj/9
PiG6uthfu6LmLsk3NJ6sWAXORwtxq0UYer6biLuu+geJPZkQBnmvIKEHF9fL6Mcmlh1SeuirNWKt
C5Ky4/eCGMnQ1UVHvx8O+9gqb0F2mpnSRl07VCXA3o0ugbEbEAJBq0FtnEyRzDyHMwdUBRLaarIX
o1rqJTJTGCI5O227GgE/DpUaGBd0PITdRwblnNUpgWrwFvljAy4uXrWvFDzdgVMzPEgdX9o0M6ji
JbEKsju6oiKUkctnWl2BBpbDZbWHH6DWAPJPvd6XYc8CUHeRMAKlDACeLGCjvURQ5FjRLQlCuW4y
87xmBe6btYolruE/66UYbbUFKIBHDlmcnH6+pgEGqwNsOzap6zXG1aaOUYIqoIyWcddIG6p2RgQf
RRYcx3UEOuyEp8PS/i1RyqkagNbzbFJ/7mGK/8NVccn/5Ngs1vZJLpYHLSJCVncuOtDW8ABnrJtO
As+m42ru5RfFdxURRqfZQsyju/sAuDodlRQWFtc2peHPFXkXC74H22kT/tLLj1Fk5Q+8pi8s9kC9
69MbTcuxAtFgMYEYR8ogJqFcEKadT0rn74Gd9YtoMG7M8BFwcVsaGDemLcDQIA+DbBejxOjg46h0
WEa6/0EUNRJyOVwbCJGUIugszKasQ5xaINdTPO3JsyxTTIukRku9BqAHnE7dsaPUp3ZbYUXDx2Om
Dq1/o4tjobEkFtbrLixDaRhGkL3n10u8sCXaOrao8TIhglmwRflZMMTsUdIppZx0OQsZSwUu/47H
4HZuwuD65SxY0qFGu6JFWcFWm05OeM2M8W5voVvQM0Ku9EzlSInwufzCr1uI/fT7FfJ3Xq4hS543
pjx5VQe6NZ3yWSF/f6Sd6cICVi9XACfwgtyylTzXfhhmal9kGXyhpJCFYu2LQDRdiCVqa0pK+bw5
lTovKWJGYy579Jq8njrFTXh3O74Sz+WASggREqF1VbiWiLNgT42p+xqsJlCcgFeLHSitRv2rZprL
Sp+UdrUYhilYIJu28MOhXGNsvFXVGcuAG/pfeqmUZA77/oBv3J7tJFN/AePMA9gZEiWVEALFtmEF
aoCZzUdxmdSWqw7pYJKo1aMHKdEgFJ2uwc0+j3lIgKTGUX1/eXndSJcVxS/Y8Cc5e0LYlKYilDHg
/eN0xcrZ+WjhxNg/syufwPUy4HXiutBHuo8LSRdYi/kkm7dTSKFFfe3TWAmymp9TvWsMJO5O1qIP
lslJwYlznK6/4hcrzLOBsYpZenfs0bzbQznaz1RoQhKHXUfkPzXau/o+nqTtD070/9asomJTButC
yL83N6CMfCmatPAEs1MhdFK8MZTOITszx+HNOZpCQ+wFp0tExIc89Y0OQtLaCi3BqzmWY62pVOgi
TCMGX0Ohfcfbr18IHv/PZqWHmeH8KbWIYYcDs3xtBtfpv4dMGbiC+hEZ1oLpB9VTwxfJywQE7ZMN
Vt5BIDQ9GGuiWwDQDgRFb7lY+F4UnKIhYX4YO4AErq8Q6ZrU7WJx8HdVcZxTRAVpE8uudQVIqYqE
DSMh6HW4CBjQt8RbKMMSkGmn7kiDTtHw/ZF09nTbGSNsG7uE/jZnwLbAuIKbV+j63XNRvG8vK7Wk
rcRlTCAiVDxLpuF3sBuUd66ieFigMMAwN0YLe3CaBaT09jiQazDh4/kOphWF8LJygjbPc2vWd522
BPf4RdmKh0lp4rAV7+g9i1N8YQ2z/w8wCQ3FKLFkVkAF/7/jeKnNSJNfFeIMqaXLxNAw74NS7Yz6
5E9TqU0ldhy1T/wT2QxeYto2zKmwsQ0lnAzC1kekoCKnhBPrRrTKlwu8fSlu3HgmWCWozzBE3opH
gDqcoo07wfTsf7+6wSsC/Y/QUirH5cZizLZCzZUVe3Xzr43J/wssB8isAfTYiVUyZmmLBW9lILUG
zj8K5X1plMM9zXmkcLPDC9xuMY4X4+lkfFDJfma5vS7I8X9BwOH6aa1Dt2IroHVZx58NhW/287qx
fi9cdKRllKLNwgV5maUFlYIpaWcl8gB2aGzfwtPXdtdpnwgVSGegU/0dwsRBTqu+xZ78Eo1awRGM
whNrCw6BTqbz8Kjzq9lHxs/JvyGaDiVvW+5O5v0R1IhvfEo3OGBOb/v2/kYw1N9eyFPz5tyR4/nK
MjW/e7xkEBHr3qI1PIS85hBbLObbKVQpovn5ctCTvwVo/a99BImhuwOo+gRhAGq5QveAT5h+5gsE
OEyfzAQvWOdB8dNY/pOcnPjLf7yE0Nu9zxXgYy3KIkSifWai+zXugwENi6tyCXoGYOnX7AwSgJpE
y9TDB5Z7VfX8TwbwgKPXHhMOHWYAh9+eCCHXmwar2vWaFZfZCaEHUwf+WtIAndrLdjgIT+gs6p+A
Df/CxnbM1cbSnduOUEka2kfFF3FLfsKU3/rcfxZD5mZlpzQ72RpxD7oBAE63ibAiVlOUB2BAp2wt
S68hapEAHhxuq61w0sQM8DIteZPUrRweGyzNVqKaJM40cCr/ubWrMz3m+D/gzqHZZr/OLBX5U6xp
vMmmX3f+5nz/DETJs2SlsS9OSLJu02B1bJrnLbLgQxnylmVQMgAAWEjafLJXApZpAKZHT8YIpa+Y
5IEod34d0Y2xqTQZVY7Huiy0G0R0BT9VF9BY6xqJrBMPUk4B+a1KgJD/CWhhZEsVUykaUllacfQi
sNQjctLdaM3HgodWLcq6jwGalnCG106t5Hpn/8goaFkW3+SyUoZoEeQB6SWHYIoPqU4Brd9aS6Ux
xNuHp+8641rX86OUe0QiY6x8/d0OF1AS5en4vqZwdg3erwjbGoqKt1V234UznpplG28Y7ziEol4c
FZ+BAzNC31ErtV8bMax8/Fk+bOqSG2u45WMly9EYOWiJKN2cs+aK7du5lf//xQe/KLv6F/REgFhf
xkMOuU15xoEAt7iQ9yh5qR/VfNdzx979RuNEm9i1XbgmQmv6HGId/sRhDlEGBJ0wCj81MgVxIUUp
88VLUU9bKrTYiA7Y0oDJ5ziAp+ytFY41zp3BX9TqWVfe5nl4DD3VJ215KDRXO5YnWFpra86pGQDC
eotJITeEQkIQ8Pov0oPP6DdXNuWyY+l5km8tbJiu7WO/3gRcDM3oh0DcmoHfOApaIzq2ESM0JXLN
Kz9SzJTKeV28uBRDGlGMwY/l9mnmJa7EcmwZ9x8qxX3D90Du7+8BovjrJnOo49ynrzFMoDLF8WOA
x+M9O71VMqtxWe7cmy2Ot//LXPqBJ3xz4ffHM7mgf79TYyVVfzCuDrWb2ob/XqZue/2WUuntAAXH
4yqJ0Erkzk916e+WN9d3Qi8Scr6vU1ji+9HGspf/a3tlLUK1OpMl854kX9tUNODhiddAL+20UYAr
Otyg5krMND8QxP6lBApwsTGLKGb1KWd7SJ69MD7hSSMC1nfKYav3ptZQWB1kswkBanyfftrnTko9
kshII4DZjr3Gp7PwJSXvhoytjzyn7wuLLOhXTOOv3NTBU9FppHpy9VAzPYZvI3XVMdb8YBCZ0dOO
AQy2g16etZ7QSfoI+SM8XKFA60ip/FnEzxkmbbb2ERFK+INePqAKheE2Wuo3eUX0cuqZ8z6ls+CP
tbGx8F4VLTZz5/cvfuDy7HSSPEauBUgFTJKCsDwZbIfEACviJUvY19IvvgYFuCnjazF2K7zs0dWh
0wa9JSpveN8bJKGsx9PM8pR+CZfEJFCGalJDzgLY8IoWmwpQMmSxrp+Y4bNMGszNvutVq/1UckuE
KicfV0rxHhzVSEp+RMkyCB/4Z231wDQGjntWE84+SE38bw9epXKoO/REizAowUtJwQclhXhvKIOb
8W7coAJhjztCudZKKFALfWtXJXuZZsu3aWWGdvx1NpJQWQXcgLwguu85zBTl6YNl9nNvWVlteJsf
UcyckQ3AGF0+1hHXfy6dXkCS1KCk3WNrXRe+FjkS3LU8zEVdF7eTw3RBCnPSmwsifQQ7+7Xl51ug
InBNhhizXRF8xqPvQCqbZry37XTwzNNJNJB9yptRQVO7X6+0+RMQ0iZeOY1+q806mKoIAv4Dw4wP
GsC9lMzObt/FMDHNOkgYxlb7l9F8KIZBlCezMi6h3ubak+wsstC+3T5iNLoTOpWCafM6xsKyw6Fj
mopbixF6LrikXD2dAU24U0uXKM/FOfuavDSARUX8lI2UkYCSJ4TkOVnSaOnI8cYyeTEnI3rQjJa7
xe+kTK9+lLmhwn+rWduC5BxnceloY4YOcuFH1x1unFsIsVZEG1e/oWmxVCTyd7gLk+/WfF5F7lmp
KZrZEBVvW1IQkRyQ37CaZPthqg34seoL1NEKBK2d37lIFVUCcI+eSc1n6LPpKVMq1gmvn6k4KyBO
v4lDrK5I4i/rag7UmOs+v+pleGAwgleL6NNlhDyIGw/YeLSbZOvC6Bk7g4gGD0QYFDWqzC7JX6R8
fmag0cG+i28gbGoYVPzZshkzG4yW+ix0MJysYOLuxur5RUhtnm6QVXser5UdwydbLYUNbKhcnqrq
BNhpT6beRlvDKxDZ39xrgMTb+cZ+9YxEb6+srmRI/c62XG1KZvp5o9Ij3aWi9COGmj1bQAffa+Xt
yAdmSF+kf8y2QA/FMvrSOK3iCSkuX5CmjU6vDGVIeflCgMCVPwBQRCxo0dutU7F+OW5u0/mEpU1L
2RXJz2Stnvm/A3GwvwC/UNx0/RJJZu0OmIDTuc6yLUNHRdUpb0ATM2GStD0c/vLq5Hng5IgHu51I
gnqo3SzIMwCP/tRAttwg70KA0KMb/XY70keFvp62qWj/1y6nn/T6YEkWFk5gMxN9EpoMe4MFddVX
4t0lNJD4tKI89zk+h1kzoo3mRwbaEo0pJWzrDSUZlMYOrLAfzZ06wap7/RS0jk6fWyrq8eANLzH0
8ozU0dvkmAbMRiRc/vsvAoVPwcTWEyT/pHHPfq7LpTe5BIzCB68ojUMrptIQilrOgxyGd6sfom0U
JZn3gRuSV4gKEXRSWd75LCGeCDJE97gECdNEyjndDO7CvGyGOANymLa2B4R7fD/0NodbS0jQjW5Q
HfYFps6+CtrnOolZ8zcXTRJbmNQGlCHYa6584tYtYePUNtBL3ckUHt5UmY10A3NUD37acjQVxLRU
ETIg7b4yx7U8FJ65kNzu9MRekT7iuSju35ySiSR61sVYI1uOJcsb9GeUAn5TJtq0Razyzp4uIepD
ghuea4m2mdPuO4UXra2qeE8LQDbY903kLEbsQ/3WZZSiPT9qau6DivRaKMBgTk4Z6kpSIvEnbSbJ
Tj9hrY5Sd+pql306aWmFEAYY6rfmD9cjmF/meHVhb6EoqpViutxEs4IORFh2XfbTpKSWe/AARKXH
+H9ymeDthrm6eBYKCQQGXGc4pJ6wZG/uFqmibjQ24iPvxhoW+cbiHs+4hamb6+0MK8erfIt3Z1Cm
Km5+ObJjVtLxXCDtVOtBPVM8wEhNZk/FvJkDF59/m6tlGSy4ZxTh83qeLqiSDVXZyBtpPRPWptC8
BDX8ZBcukdnOPoqSGWsxxPLcDUUWdITa9x+PCJRUwt/KKN6NBBgqpJHHUZfQpDh3FLyT5C90bLBk
BnJmh0V4y6lXZckFoenaXrqEacHny5Y/+H4t68858bS/KDe5YqyZAtyiETKNW5s7lZO2GHmFrfsT
qv/z0+Ovj/i6l2F5NcccKc4N5DAwaWeJXYLHJ05aMj2V4gPhHKGj0SgAiY7yr+SCXvTFJmWGGwTE
trLBYlbP+y1AhbMHwRUSCC+3MjwoF3QmJUfv/7C7ECjDHwD2tIhC+VIxk8xB9bPwbX2/2wW256gP
xnGEshST5bQ6yIuFdRdmkSSokavwjwOxH34xWz8JiqEQ4QFkOJvNKbOkg9BkJQ+gUE2cxTXg789F
G1Dw0qifjD3qvHEWcTENzXIJvUlPRRYyCSKl5EKvL/10F0zmmCeP0nSfc3UZMl+mtjTywoo3kMkz
ht6Gz3fHXqWHjkk4O12W/HW3fCWvMaNzoiODFrBEpSN+Ngk4rGSydmZ4UGKyTnd3LoSUwZgtC3fp
ETeoC/vCDKuPx/Yuc3pQkuajtPeQDdp5Pz55JkkeEVUUg1QCqPwAr7JwwlzAK8+W0tBWHX2JhlFy
RCqwPTKR5r7U1BrtEftfnwJ0Gk67hdS9vaUoOVMWJC9RNNJPr4NUZfygfEhL5hjPNFhPveX6gB0y
1FuU6/vefKOzaHz/Ay7v9opOm7b4hEFOpKDTEgps0bbk9A71rz+PlGB0WCX/IYqkeVg/sZYooLgZ
gn5zv8zIcwg3elPv7fECxs6xliQ8fi2rKeDS7jiBiO1G3XC8j3x6h8leTWi87ZGBEHHoKKFUqstS
RKVwKN0v+uhU0KzfTSQkT5h2IIksCO/xaIdUCnX1ZNMvro7LS4yAPuO+V4lszfzG9gLYK2OtmEjf
eR9ZnjpgmJrNWN8QslP8APsPRhCK0gqId0Pl1ykYsIcBnhaM9oxhAleaBdRgftFJsD1/y473DYcW
W1Y2ajkV+VSKzFB9lkFV3oW2TVkm97ZbRpkxlQUALfXIMaH41RzQbBvi7YFZj1w3Mmco4N5eaZIg
Cwnuu/Lg7MsxK/Zq6cHjt6rZGvOtziGaHHX0OPPMnIYbLLPID47p5L9lYZ5/xS2iAuH6469Flchw
FMF29bIyJCWAJqNu/hfRX5D+yPq8dMxX+JOGb7kCKwijhyNNfzusfTPfrIPxi7vTpWkkgA1ZZt4c
eMyTOgvUWPSiO/uyZ+0/ypw6X56XDyJzhwGJK6gl7P8OOGffl9aCwGS/BHflAc/itZW5FWgylzRb
5dNqIBvQCoV4wZ1PB6xgh9DqlEL+L/mJwSij3gB9vdPil+6gFKcxisCFardAVBzzsd+MJzzgdj7V
GXFBqLjLi+167BNdIoWbN6kT+UGzSQpGirQZsHk+fr9eAJ/70y0TkA7QXzh/d81svrno5kawzsop
lSt9BVxWOjNk/AEDNCl4vfzD+P7Ime15i1EReAKz3eJIipl13Q1w9XUeljBaGT+orKZd88kUQUF5
VSqfHiMTBj5B01eaRuedQrWNs6Z2TRJJcuTrssvfaAioY9QnapKcFWw9l/x9eGfD03B5K39c2J6X
3psu/HaZqY3bmvgECJ6aOEmwLRT0blZQyL481WzK8XPPNbAfbOREi23qbQlAl/0NcUdH2Z35AtmP
3QetIJFOtmRCkIm/bzq4wSpoHoMhuarOMDkSH2AMYKk9RzsWA6o8xB1nwie0M4RJ2+8MNr7wKInz
7ol3g1KJmKy6qhaHtxJNTWxjbPo6aC3XcGU+Doz1jMCxFa3rtowjuq2yYLLY6SVV4oNVn9xr1QY9
Ljq9IMGnt8jnzmdEX7x82fFPq9Gn3JfvT+zWcIZFp6Ec7r2FrJtm9nAAd72/UqDjsSpFfMtDFo9o
UVuG18yltxELUTJHWb/25bUc6+P4ZUL7+q/EXnIRjkkLJMBJxNfuIUsu+m1KrsJdcp23ia/A+rzm
iC5dyuR5OctZ1VcN2jtAT1ZJCUUuUKzZHQTvS1DkIjBo0MBcAGdTNlop56GkgnyTKus8ah6N2Wvu
ohc4e6wy0r/MdbEf07JkhENnVSzA3Js+QpSc/gBipT2WiWFKmZGvzDa3pyXhivLTu5ZB4UDd03Do
RObqmw8g+PE5ireQNdBqYo0LrXomYude1N0JtO/cEAxvkIwscUEOuXOy/5NznqAltWQVp0/ovBKc
MhljZuFt1LQwRNZVAHhExarn6BP6w6hyXTus0AbCSBydXPfG6ourDjC5ZBMhpi53vLKh5U0G03jI
zlFXVbBNEZtGo6Iv7nwCA+3C38Ent9pIkLPEDF0OIwWXgoVfOcheGtfo3QoNTc+o8n3B+u/vZWGW
Wo//q7InW3aK5L0p2b7UxIX09TL+Z4TyOBv5zB8dcU+tnGeZdeQXMDTkYulVMnRu6QdL8fra6ApR
K/0FBtKqqc44sjLFbow8wFbAtD14mjsztwiIuV03E2h6TiEHCncSwxS/xbDebZCU+GX/81DndxMc
TWYSyCuE8yHivl7XbU2aII7lyFGf9Ysyld0j0F4xAZaPrNPtYdwaaehVX2XnTWR37qaehke4XBQb
hcr+11Z0CJyq5B8QyOHAW9yj4rSfslV9YRVGEAVPpFNHE5Ox1fyWIlFbyf+BpynvQEYQC9vCQ17F
o2cDAWXdm96GQRGASUddpd5WOuxC+kEFzIjL9d6Fb7PK9wRPb/CY83c+bO8Ojus8jqRJ6T6xja/V
FO7uCTir3ru0V2LrBkOHRmTCnI7fAlKFpdYZuntyhQSxmLKPRHPuFpOLZBfpQzByPTrvPmGc/+1/
d5qI3b5zxrmxuLSeXCfMzq2eWC1dp5x1nqyzPWNbGjW5ZG5BazJYXXYgLZFLzEvk4O2rLDqXPDOB
vnK+38+a+B+Ow9pZoKy0p0DjWjAac1BtFMXzHsrumrWtwPd9ilDxb3UhHh7XjBH3TN+3x1PykBw4
PhWU/cVzoYXgJSlc3FmmMRMejFF+Ljw5oskGiu+aiGTjSiS0Jm8NMqFemsdX+GZWo9a7vnrp5wez
IwNT3iY/4epqq9qb528bgwdlG6QjEIqYz7n41xTOWtO1lyaovxNgCAwXQHuTSLI4n/0ZM4YXZgAV
eO4sdzxZT359hfUuEFva2U4g4pbd2CrdDH/SusxGAgls2kVkgoebnQJVCIsMtAlOPbs6YAWjK5++
tnqHFmTt7xrjWh3ly8H+oxfAXYqNywwdGat9qDlVJflIQQC/kHfc8/fbPtk6Pp78E5N5JiCYDxHl
mBpowT3gr6iBLX+1Xa3seoAi5O3HJIzAoHEVNPGdh34o3cIaYtk1iQHv/Xp/6jNDSF6YHS4gR1nu
1+aWFdzjZcbzVNQ0QoG9mnGWCfCZb2YIKPknHt+HjPUMd3trBjXn0fOTS370rzbltcmcMaZ9tCLg
M5LugmDhpwY/4nZuB2vLK7cTMQrZJhusIdu3E+gXNclco9HR5SqkLQmn09Ap22noTcPlicWdQEwS
gxfq8E+J55vOeztYuy8+12dwkzXrVX1hUo3a3EdmMI8Xo6UkADyEDqtK9B1ese2af5YlVAU/HD2M
rcGNihjhX3EcJymf92XYZ1b0A8/FGaC+dpV7J5fuXVMrV8S1Va2T6qvWscSEvEp+lED1j/gfZlml
ZTGf2pbE5sC4NSBlfAq0/gPhRARINP2SBRR4ewXV09gRbi/iNMRW09JCjpF5oKxjQ2j4okJkAD2x
YHKaJ7aSkKHOzdri3uw7YsSb0dm4mQhzauiESaBpW50ZDxQSAWG1aXwT6snwJ2Nv4L3z9fom+aFz
GL4LnsUQ1K7wOIgOmhAY6OQQpbd32gBprNk4lLoDBHTN7MEDhbDeDuMP8X34yDAeCGMhIeYmhPDJ
/1zfWqwOIeoIg/YdgCdYR0ZlIDFbUjjM9JluKsmMUkCGGRP/Dui6PKfn69M1hfT0Y/qA8DrK246x
QrX+IZ6nd0Jr/rmii3UyD2h9QyW1hntdynpD99FQ1TJzfdBb6ImIylwHfaPLLUjb5CDNs/ScRZ4p
QRN8+hSZvLuRrTf/kUoIBCf4twuEObPldvCLP4eL8+7TCUMw93zZRTN+CLAcyGU6Yx/bUZqqDfmW
6jDr25x9B8Wgw29Rer85VUjVtj41PkqsGJjl4VK2Yq106nL4/qISmAkoo+1l19vMClhfWhsjTv/y
75AYHXfvN5zpepoPMn0AeIt8bgibvwPK8Sa1lcStFgQEdjxdeohAd7BP5lh6clmaxWreiHZGeXLu
zIv5/I/kaoEo76A+mR5mE6Fdxx4Vua1UJZ4fFyadJU8sTK/0gxJqbsIJWvRP+Js1aXa13o0h0HlO
tVFyrOAQZe98eTZdfaOH1caEaU2SunXRNtAq7frK5UDQ/e1zs7VFyALJ5xH/SaBRhSQTrKPslNYE
NMCuEMarihIaAqMcFGQg4ZURbKMArN+Qz1M+YlN8GiM3jQTqnITiA+Ao+bUsQeUTkdLS05S30y1b
jKcAkB9tOh0bEeSkjwuixQgn+MLyKNIcy4gtnVgLJ8JraK6ue/K3ylR0psz20mupro8W1nosAX6D
LJKyyFDc0iRXX9+eeD7EqztZaZZ9xbzYAxiyz6ipSf4BBy+JLbqiw5Dj6zWubume+D67VmL1Yt5H
gMZPVbgHquIt5PmkFfp2BPeQR6oHTokeI2HNHS+FviANF2gzFHJh5iqhZdgBtFTi7MJaKPpUXZnK
GCnVoIqZOiudTfrbhDuY+UWXxQBARQWztUoJntUOKLMNfXVQa1Oa4ZXirm7V0/D4Mw8UdKKkdJMx
btqI2YEwKUIIOYXsZL17R0gcTatUBuRXICt5yK7pGVUvfG3ub4NJEpCmS/fD9NPpW7wwIuan5LsG
rufDwOSk6LoPmDLCGn9SgpX7pBuA+TbjqwUazQt1etYHaAkZPdnf0O2qnFCh1947VYqjjZ2alQ7P
T7RpYYY5ScvXWpZiot+m6fFZS15l0fXS23vjDUdBueYFY/iFslLCL5np++hLU2iPjZxH9SIOIf3/
RHD8/J7Fwkzi8PLqGaXmBmg6tn/QwojPgHZ7q7RiPbsnWkWCNEx0uaUuZqAoD00cibXTwf1zqVP8
SnlGk97cFHd/pqRzlpXZ89LFqnZ7fF1OlulIlQkTVSVRP5Dz4R1e9/Nqa+aNwuresOg4+ZikIBi6
7O9mGCKZHFCuoamrZFvDTOW9nMtpLuvJ7Tzfa8DiFsRGDDUumrmfbOs+BniPhuqxpAkJWnctfFXl
YrzmDFDzHqUfLMmAJigZn8MuE3XKRQg23NUqXnh3WIJ4FJA/hlS4wZJwWEKLKb6I+pWXe0SRj3I+
xPAc8KdncHyoW1cpmkeO1PCYu3sxbAz/fl4eK7BQzG6ZeVTGRHm+2qTyKLb9d04oJQkr9k9ANnB/
XyLbmyoMvgu9yDxy5F8tK9YBad4nqt7/P5dZHJ/JKLingMIw4fqWnLVg+1dTHxT4NsXScHQrDtWf
G1Vc/2wW2BnjcNjgOwuNSxFmLZoT7Aj+YZVeXTTrq8H0dRRjSUS5VEKL6Cn5eMyCD4rEZLRhPdR9
UJiGrjnwVu2fgmY0ZVutHGEzDWBV1xBYHkH4bbNEdPHNLY7pZ0eyaP89yWnsjJdtBfm0s67yqtt/
gqj9OoI1wN2AutWTJVgGinII4FGHfhtWswvm2fiJQUAUNgUIH7ML9RpW3LG7p7jypvDuzMojp6hZ
sGUyw+wgrH9Ps3DvlNgILv4i0+A5RaUFxdSj7V5ko0qFGhPyoTGSPZWr1uTjTGcGpvHUZc5De5Qw
u5Z6NPByohzWfGUyWSdD2slnUQibhwozzQitEg10dQrfXw6x4LToJWi9RTjTw2zgy9F302owh6rf
B+4nhFP2urF4aPQHCnVHMyH74uyN9/H5pxNqTMI/C7FUzzqbS4v9gLgCTqTAoGQ1H+xaQ0QMJgDa
69AAAajJjpGNvri19veYaJTGoOqoNE6QD/oeBxfx1eE8/UDYf9hvxTq5QXw82lKbHPbkwI1+ESBi
+458wjx5ljL/jNOOMHv7Mwvsj/WjIT4at1g9fA8wrsZ/6PhFpYsZl5vmdpv0JKDjbiwxtAGbI2WT
b4/A/ml/T4wXwuu19jfWkEFKBuHm+enmGohPhND8/UuINlVY9xDROnJCn0XcPPsfgZPd1jkbFEXB
6+z+R62H3h4/9Vh0+Bly9SYMFWwtDWeKyVezx5x9/uaqb9Alp8LxCjajXyeInQSFEwZWFoBgqady
ZGklGqgLyT7UIlpkkh/31Wex2R8U2HfBwT/onbyy0W/QdAfPEY+UhSvEG7erDxeM9qJhvwbHMNs8
bcL1zxaJ8sFj6O4jdA+3qph/DSXCS/v54pqGPX4qO2NGK7+hraKAFzxXu9Ipze+h35yGGXJqSeqm
DIjPrzq1orURNuNYJnDA+SkZOfusBN2QbCZ5Gp3Pj7bZsuFIjw8KiuMBkQE/Fks+qhHjXCEpi72m
+znQStF8wkcRFTSLYOcIeyjrDg1MVhRgWI3FCqQzykjLJ0+prA5jVmMqkJJWGLCG7A4fpjOFeT+p
xUTn8IKXrLZ8uPPgUc6W768Z2dVYJNKJhtP7veFF6gKOOj0WYDQ9TYNcXkjkM6lFthZULHwzo/ht
qYnx7ItEBTQb9vgVkugzv3kOvsShf4XJsAC6R3cqY1jxfktwXQ5JgUpMK+XMI4icelZHCeABINdo
akz5ogmUvUQFBwsZaHvg1znmfDt7mU9IEsLqC4k8StZKJibTNgehZ8Xj8XWy/Iss1F83rWjo8LZ+
AVWzw0wBqHMsMZZjFXkcbtJWWV9XpoL8pJTG+zA+aoXzCtGojYab3JvihvjDbKCspIccOf6Txryn
wp/h0Lwxu0gHKNdhtmxUc5kcMx32AqE1PAAVNiHR+KaSIj63mhxOZC7ofZDhAlrUR0xbGP30HjHA
/iPwhYpMlcRJMsspyprmauaD/CzRATBVpOLn0SPCgFqxoavTAK0Ypyy+RKxg1cwjFxM5IYbKFbrn
VjYkz0nSzptzIP4bHauB7ghbTl7k2myn6x1QGhXVrrasKokdPqLGo8c0G40Y7nJUDbDMQUiOTYVY
w+5ovhour9Ii0ZtPj0ksNj2ysBxs/xem60CqsbJ1yXsRCWT48U7wIk8uaXxhSP4dbMG3Tqoi/i/j
tlkzjXuCd6SvSjQck/4CyX9zWW8BmMxOhmLrSzE4kKrgSF+VYzur1lsKAzT1QF8/ryoEMxjaHcS6
K+QZByjTGxu511cT9FST+j8l1qq1/v5IwuvY/g4nfiu2gIuYlcZ7RqwWrrNZQYYk9x9roIib0iM9
7NkjiNseAaFUjf6OWgcqRNRq2mulYbfPUDuJmDZHpO5q8qOLJFEdChizrqHOTOgbgkZIuhGox7GW
IA/AEQdsXBrOgqTkpPj9XyntbnGpNYXNkqBUaYdKtWT3J+U+a9wIck985xAJ7vakSeMs9kOUJc6Y
n9DOh1Zt5rQDYWvMUVI2zCJQDRuQZhx7K/8QfqIk/OX4zf2E05+LODY4Dtn0H9hxnABu1z3zqEtv
McYzxgLa/1h2hOcwZ67lG4ZFcDNsJC64+BDeAxhmAfAQkDqzIqHLXEgS2s5Ry5CmW7XxvtKjMzFe
wtLkjFrj2jazH1bUlVF7sj7tZH8/8hshfkyFHtHpdUoPUGY/b/jbWkv3uQJbDxoR7sfslrB8ZFo+
vt9KxB8kpawmr1FQqCstI9IqTR9uriKI8KfUEqoTq/puEKwCk4pxvqGNxeVDWTqXzCGYMyFjOrp6
DFpyM9ay42EyJslRlnfmNX3JQ/CgWe+nhsr/fETCCGt8BEB7M5d8bVaTqTc1fSHbpbEQbEYBZD7o
xwbqDe6Q3yiyom97mL1GEzgswIBuzTQOMxkLxd7a7kB7ll9mQiOqZFDjjMwotsvND1Q6NJYMhwzg
Byynd3W+1bjA5bH2VaHetZRZex/JAceN318FLfh6vRhf8lVb/hKjFT+eKPW/AstJ5jQfqPLFTqbw
663H/00tSrVwj1xvNFHCpjDQxM5/GUjGkVT1xaXT9w6MMoxZHYXvpLj86S3zy+pr+SLZDNyjheIc
/yeEKfngaFxNs6+MkllYst1czlEbVGMgcDg460IT1jminPtUsx26rgwySfrg/P4fx/yD5711eqIG
JjjXrtcSa/5z3hngxf+FewyXDfcvfpScy1pc/TjKvnvyxz8iMop1tcUszSvjKw4D5JcW04nL5sKf
+DzHReJwlMVXD9f4RsBs0OiUCbNB9b/xlv22H70S/8GN5hoqUA7vD25aLkM6YNxisIBZ6nn5Q1/p
12hiXdRfdjvjdxjsooddC6F943FDQ0RP/qyM5WQGL4KBovM1sKgfXD3D+j98C4sOg5rgpOl5mEMv
s6X7EmIMeY8qZpzjISoiGkN1eTywsUq34HMJf9yupDu6qHY4Xz46y32auvWHhBNIPETBRyjUHd3N
RA838kczhsAQfr8cJxtQYwCkAelusUZAWJB/MYIgzGyOXCZqm1YSh+LD7tVgip7+r5U/MruEMv+W
6TYjwC3vmJNtogRTL4NibBKjqynlosKLU4SGB4rV9/ngb2pJ+pBLkvd4JabEE8Hj8Zdh1CXEngFA
XbHI5Vv+tQQ2yn/EnfwpsLkyjy8qAPOXJJDTs+TiKtx81AKV0HWdhlx+fX9wFvV57s1ZhqUuk2UX
XYjjzqeylEBmc8+vyZtHsCtax7FIlv3sPsqPPIUDSjW9tFO+m2HhBPxm+5vBva2V1Z+XHqJKPP1n
UHCZMvc64pm31cKKds0Hxp5dTDP+gHc9Ap4vGAO/70ON5WfQge8B3578K5j+v5+pCQeIOnipozv3
XSDOBQ5RL4ml7Ac/h6bYM8oDYtnXBlIp2yJE9JVAdyNs62Y6WoN9YlZBkAKqeboqfFU5TYi7A8PH
z+qFrvYP0z66uOQ7ko9HllDqr5GEiGkyCLXXybgYq2noqr0CXYLYkJFpzb2uPdj6RJ4Dk+TDhA/8
Hy2Hk9hLVRSmC3Zbnixx2hIXZTRptaq3Ro+oFDyRGWOypBrKCnqEHWsgU5/MP9nEVIzACalh3mVU
+o02eZbgIhEbjb+kHXwlGFnlDr4ELpglHrvSlKVti85KsPyv+1I96XiA1puW/656lvJjG9Aiu5ZS
hTKHS615JAn5mvJyXKPkZgd3eekumv/4EZKdwkE+l/vOd0Vsu9mmj7wk7omOBS11WIV7KADaK1K0
EnDwQdZnFaRBAllIjUURyDYp/8VVPMcPM7b7hpWL3Xc1sssKVIYty6BSD/0wjD05+GREujH7PgU0
pRxVojQeK9fktosqA/XH/yYGzyFUILlQEhuPZSpCLQFMbTKY7nD0VvHZ4bKGxqtCXA7o6aLGjGj7
iL6rbxEDPi92pHpF/+3cKpAbbfjQZ1Bv130dRCCZinotiArt47V6MSZvdNhUK7ALl6Lk8g7ojjaB
aUMczjOJFixMJq3ym2rkR2yP1JDE3v2CCyqNtjYTxn8b3uVHK/dLLS2dyGndBMfrUH4zPTSDNcVD
+gFm1jenrYxzzioEf/gksCBNW+bfa+qo5awEwyem7Oab992no85y95l9034kx/THXKz8Tcu8Zurm
N+AdSoIGqubxCgIcBfF3bibvYm9aiIYaAXBiQ42aAWUwDT8l477T+8kPkIS85Rk9kKNkpmktNC4+
v01ottuTrkUnnMbUTKLQaImBVIfmiNHIiHTT1SjfFFy2OZl0BDHEtZxedRxY4IuywQqoZZvglsph
gxhnH3SaUn0T+TZQqxTBmMVjYHhVpjrH93HJknbPXgjW5xLahcI+qdZ45nP5cGbrQCq+4P1Si7+h
nEhgdcmnSPdnbt8KxHyYk0B6wcUXO1mYBqga4+GeIRnPy9zgVyTDGMojD5nXjyN7aL37PXLwfNp6
aIvk9chkVFVwqTlMTMzjTUgLdYerU9el/hI1ABplie1k4huaD481DWAL/D3EpHUJnVpM50553EBy
jF9a9vbhbbAHUO270VnFt3V3RvJZeisoRsZggLfzQ94b1CilKAIzHqykXjW6X1YVJBNPvb6MmN4g
9lnpyR74cT2XeIhklxGpAYlbprdENAWVIhBI51fd/ppicyAyo8t3PQ0NfvNBcTPw5J/TyVJXjehs
8EBYIBx3kp53JrWK9uVGHnaRhWuq637iGhrEREyiBlUSOmDeI9ImtcbOgyyRHbav1K8wtsGIqOqy
o6sYV/tEPf49tvKB4MArn60EAH5YsFWpsTrTGcIhXK7Q57vS7LNlIS70BngNBolvzgk2NNZC+nP9
gMWcuNrMpKuxTs7iNzVMZhNJ1A10YtuWiQd6dfmTddYwm9xjL/WR5SjKxgDudG7N4bgzdzJ3bT14
mEXei1HE3H1vS8bTnr+SBu1D4JUiv99XU1ZOrm99fLfdyZLbluCdKmho/FEmlmz6++wcaeZsfXJU
eYNoGpEdB+IH/U49eTJwzmWF6oxyNuPJ+GbFlBi710rxsmSKJ8sbMVVdvcssS9yuyYebjDoMOPyY
d3bWM4tvJKvum5i0DESkYXjy4yrZWqG7eFYfUMGtWcrfzq/jv514TcJ47jQ1XvPqJxcz4n4YJGWG
UCvu3scbNzoemEP+tzM/3CmVNd/9e47mcYDt61VA3Z2rhIMdBFwKpGADRNX2CnEkjf03XLORa0k4
VHaTGtnuwj9+8D1yzLxTUPyCALWJH1/K/RjQLs7HSpWzoCBSMJ1oBZLr4NZnQ23vKSDBmXhV2nda
jk7jBbA+ZaFeY8w5dNrV5tFSCbo/ZDV7h7depzt8XWtuZTw81x/eU4+HSllCkq0HRm5hiJI7lCVu
T7zZLEGP0resxa46mGIWTNRPbEcYvomt6mJren8HtgU5skxi2sVihImQVbkBryere+CTqpbAzknv
TSC3svXBCW4Vef97rmnu9auL5ErLxQALI41N8iV4PT3WrCMJKElOPJgB7zDbQEQ9Ip1YHthwf4w8
Ww5UUyd4ODP7tiP19+6gr1EQI7gmvgbmp5H8oRfn4eyAQub9aSyR4f3Ynot37subC0CPNwoetMR8
aJEYJGg0KOqUYprDPFrjl6A6swJsHXEx3bvCPqurEjTP7EA2J+Y/w7xte092wTEvV7HS9uvcRVwI
yEoZRg5NgYi9u1Giq2s7xDWgwyvMtxtmuYSiuiPLFCjhshVKpf16iDycpUd9hxr+I5xKrQZtKE7J
AoXySc4u4/M5Z8hqsOc9+FG1l4DU/E5UOGWhTQcIKDw2RSBJy/Fa5Iu6LFeYM3ThCmIJ4rqlY4Uq
QhPDovHB7vHVNZEsBBKVw6DU3wi2yegTmLY0CXjXkKivDKhs3PNhWohVS1lt0omrPzDKs5iZHcBd
QST98g+cwp9nyS0oTYfSDp8vMSYeMYYBHVbWL00hmyjsvjMnhxeBHjhUgUU8UTHbB0WFO3JD6GW1
+5KoCGIyUnygI4/UyuliI2+8LT6RAE37x4THMqBVcdtBYG89+K4j/5qpjPaUOiyCyfKVd50Dwpi0
h9bXjaVnEEG++RKXxiYZbIIw+nsj2lifu/l3jZHUGCMU3E8u8TIiQmxNea9INlz15VUAagKdYKKa
bTAaC2l/4WbNa2XTGhHr9n65cRQY3l6Bt6m0SEL/MAX4GY0A9MTLvKxraFPF5OVRR4FoGWlezKRt
OT3ero5bZLNPP4FQy60CS3JVoy2qD5cllGY7pr1CFlP+aqrnGm5336ajUkunFcnXg4CxuHFeEeJH
9QfWBv0cCO73uvbT12CsjZhOfmr3FaB1feUJMVj5f4xIkh0TPQOir60Jnedcmkn9cxXMKc9S1BdY
RIdIsJAuz0hpcN3cmNGE+4XLVoWDEecl9VAUZ2dLgp3gmeQN0aMMp6Erh1wBiowpB/dAvtG/qzYo
y9tJOe+hXmJcRGZN5IqEDSMDiTQ9kuY1IMtUp4V0eoR3mLCbgJdQTMRVlCzemQDdAmc67sh+iQZQ
Nz7Nh4pl5BFLuvnPIhRKFHpBpOSX7rEoph5yMr0g55YwHJQVV3n2UzknDS1LlFUiKdZKYg66gSpp
n1mrA3wYnSk0JaaDOIBFFt2Tk8f7HiJ67xVTO/DLg9VziMv8FuR6C+EODqoqywi7kPyc9/e7xKkn
LZ67FA1jjSNHiQxFI3ymNBc+NUwSoSkinJueCfIg3VQYLbvj1vB4uFvluCZSv+FP3l34kteWzgBh
c+0AQiyL9cAwwLFxNuwH5vFwAivxnRYL2nU/f41s6shfTEewt5WSO24Dv1eOjtXMixkAEmDZXYJj
5yuxPalA3qL6L+4Z5ImJrzGUMyVjV+Fwu/7YUeJIA0NaxpvscKcAT7DCn2iuxrVhlqaEwkSTlWrJ
fc8iWMyVSyMnimhhi1KkqHzYvZgjO/nE3LC2KZask7+7UsKx1NHG+qQT+Ei05yhK8O3qb1f0H7Ry
to6JJcd2hnRdMQ0I2rwKCXMPsiR0lJJzsGGFLBY0loLOmcn2kXZCand7fAAmBC9Jfuo/5FyOA6QD
usLC1pqWMlNG0VPXRxwEHJArGJEkEM1xQx851g2fdJc2yKC3cRdwEwL9zxNwFubNwfI70OiLoJqG
BekAH1NksYVhmlDHnOU/inwW0aGpZz9IxnYNuWwkWHqZcdwU4TFQFCRxsJEy/2fIqEIDza5atm2j
VpfA2fik983lwY93w+veUIgqCbOZn5trAD5vJdotYPRoDTzcow3N7aYT8Zd4Tx16Y2VdPkJZNsUq
W6zCc+kf7muHYakJoC77pLmJ58eop7nNEFvkvsKTD/ubdMnbpdwhN1hzdjEdzC8WvQXshKO9K/Z0
sQGhZTuWH3QaWO4FqF7Jc1ESqcoSK3rTx+LgKtuMBlKmLvSCUC2okiUewhRcHnJEE2zFa/HCVCbd
JgXb4Pzrx7dZmSqxQmzVBMgkU+sPgrJQLTmIo7EAgNxdekvQn+futq46hL7lQvZEPaEuGFSjl1FO
qHQCZtOxepOqq17E3muK1/L9NQ2G28s41X/nao585YZSR15wnU9guACi5I9CUWkcijfIgHCjQ9T1
z3EOmhHYw1Yo18S5WyCPaPYHiKvYhTxQzaWn5e1mogR32oWjvX7D71jmksV7YDJGTPvMpPdI+vai
H76Zq8EaoHVo1PZxVWb05qOx+t35BINzirZZR0ZF2RAMP0mU+Yr4EtkvoMNRZeYnGMSZysSX+6pq
rpy15iFt181YOUCN6NN393gcaJF/R7jdfr0JL0yvABxqb+/XXF4R/O0kjcJQjVHaPKyQN53CNc66
caSXjFauZuXUvxuYYJLlvmiX2HuuDjCRumF+kwEyIwlRA3eZom/95JJdYAswqBT7jYW7QlovIrk/
j7cWgj7TGNdTGMJstBban7TTt3cneRwcaLDMvrWfoXVoudLQI3IPto7QXfWAUdmAAHx45v2UZRtp
zl6XpMd1ffKPUngPpWIWcgpfimhFzBcuzVCBmQvtuVJPQTYh/CqD4YFOOXR3B/00fyZlkcXVJHj9
egTMkCrFL7SxZX/0++LEKk+KA3U5fX+/ihaAbpX9eCyWH8zQDY/LQ2etk88xdZXhw3TqWXWm1l3+
f9tqsoMqB7x1kqfL2bteSYvyrqPrjygYubp/WR1rFzuoKC7TVu9HIfmPaYq7dVptjXmSz9njyUhp
8yYqJAxrYCd1MCkrO9dQdDhBqySmImbBcWYGabEtJkWEdNyeSOeDa9FrjEVMen0XSImD+iTvGWUJ
h+iDEtlE4efBOOmtxWxeJm6VyutpTKLO+ONf84tU1ZlmMNbamMJgq0dckNKCatejltJx/FlhIKd1
4FtweKWmvPdwM0TDI9m+sn1BqIryP7MXxFlbCeCCTnGYEjLSOTylObtsXED61bEf1HNm4M0c+Vi0
qXNvaf2zLKxrGwDfVvmpcvLgeHrLS58r7i2k6R/HcyweHWgqmN7qjJmHPA0iHOf0eujmrXwv93he
LGZKy9Leu6VCX8Vnn2fXdD4LFeYEQZZjgaZGryOfU7B2CXY3N2pcJTRm2rGeygRp3ie/376DPnv7
I1oZwpC6KMxBucJGtj7jS4XwI8bvPqA9CuxRF2mWXkWtIsrNCJc94pscsupx/m6yc21AM14k+1VG
UbJuMOSQw4rQ8dhzd5Mz1/xkhsRD91H63tl6o25ObvJyL1+5dB44zHym4/CSpzPXMY5NrBI47F4x
/00Ciuutx4dHsDJvQazYx1bvaW4t1SsviQr71UGSAoCpcopVJ6yyPgjn0sfvA1yB66AtkQgNDjK2
Jf1WarQdlmhW/1JIW9ouZdB2Ard0hR6ItEsXuJ775603Y2tl8IME50UUHOLuY24+XMMUR/uiUCvo
FvKTOOFxSi+8ubKj8GkiTc90iljQeqsT7hybm/ciWlxSKumK7brr8lySLshMSMtA16a0HCQ96G8z
3L9pfsDaAGBAfQr+DPaiVstuMskaGuMZkMqXz0AfP4MS8nlBOOv8Hp8D8P8gm7vROASbqnqttOSS
0bkHjlywlC1EF9biG7N6MONhV1biuX2KRy4Ro2hHPF7JS2kA6ESs/CKaS58ZsY3bpoAMFZcxqfio
kYCLs3ftDXZYl57motkLbwfg49NtZcUfSBINsRSq/Orc/BtVUiAF81X5hyqjJrqPq84cF9XdIT0A
I01gI0B1/CT28t5BQ9j+24ro4hRe36uPfBz9/NDkRlkt01k+FTvJIMmtQ6GeFPyHzjzSO+8qLljF
dB+DIcb+pzBRw8cCrWXen75OTwfZvec4bwU0kSH971ZgGGh71FROUztht7Hg+P4U7+IvqCQW9ze7
EaC6M57WW00CnXk/plR5U9FJecij/UXJaYvhxIUtR6sLRhaVCyT75UGmNDcr7QY4ICAi50uTZBgC
V1mDGW3+Qx94m/Nz7k1GnAipX+zE+R19zIa0GXfR3IcUxG5zhGUNUTOHer6LO+5OH/cHcoC1WC+0
stMvGYDYrH66zqkk+TI5m+f44T8HTcyLNKPzBf0WI7uZoIw852BBorGcOnEiKankg1/Fb1KTidMP
KGcaJtLhpJKvoTTZuN20xfzu+H3Udw+fWO6NJCv/ePfl6mvqLb2Epsvb8DSp3m2fMFbuY/jsS8Tl
Us5UAsvsFOegR8yGW6IjK75Va+bzRGaYLDmzzfLOlFclIXAghx3BNQ03xuQMVtlFkkJKzwy9KQpU
bwzkcbgSvCV05qGPyIVhaMcpq7irIi9M0KpckqnH30gVZ25BsaDxGsvLBii+hFRQBhR+iqiIej2I
HZu8BJ8KitZ+XgQeyeRaPfMhN6yU1UbOKOJ2pfAH+jDwr+abO9xfYRYjwGtkP+DSq6Sqv+bKh+te
i56zVpYM9m8ny/oGvGr9JWG8dKA+N+CzdfO4clbfcgRoJNN6ENBCKRuSW2jhBAnTkvNs+6hLBgNC
L+tCeCCduTR6ImEqQoHyCzHJjrGiMuJeZ5xfbDzF482GeGVojzBrzReu0Wz9fTTRJIpIx4fIZNcy
BIXpx2prBMMhGQ92ZK+85YYZySCO3RfSgrYcFwJTfyYmYE+43yN7PqVjifKqBQQcmzznArv7JTzP
5bygISYY+ymFKBjtxVNCLcQ+R8c8mlrw2rq2Sox6tfB90mQrB99kYSkOAfD0QLSADGVjtpuon3uR
rYqnz6t9upZbW2XrAcGgkVYT5SzhlUVINe2DbdHejUP0olS3i54Bs5bFr+wq9nqwo8s/6NeKYKKu
Hq3me0nYf9qv0ZPAV3Zd3MLLVInYhEfvUYXFmb9k2CuCSFqt+C8l4aASZfb9HJM9yaUyM0189wWT
Kt654nXXvNEpVWpa3M+eEv+GLEFRCXrIN+BGBlqQ+7JK5u6QwvoSYF/5OrMPZu4nspSTe+rInsTH
FkJvwgE0k9djiJKpqUP5EwQgYtlZCOvHm9bSR/XLrhpiNN4Qcl2CsZP3xy7TYu4nAp0j8Nx/xJTP
h9l4nZOFcjjpmDf7wIgEbtXniRLLsBEuQE7ANOzs068gJHXKOFkiOHPoOVzG9xsJMbhSYLbAozi2
zBPBKpsSKPcn90v6n/WHxmuALPi+0r7uboi3cz9cNpQTq9F17ZzNtllzadREoFbG+EDwFn/dCfa5
/nR7YEgWj5+PA3l0FW4+MW1IijR8SjcoSDA3FI+pIOD4YFJyBypLRSPFJljUdbheTdH8qVY3TWjC
OR5NKVvilWrE5VEi4zqRFVAVrK0TnXmd+kUwZC6VtlGCF4upJSuiG7u5RdgmgYioizbTmourg1M8
is0Y29w/y9eEio4Bm2wr2TDGSaH74sVWuLWRuhK1exx8VlK07KMkEb6LvVcBJ7jwxLZKfUy2J59L
zPAWdwiObSG5q66ZYX29fUOa8eJXqQVVhgWo83icS6YYrNXqdpT+USGFX0eZDYRImBV69+Co2GFf
Xu1eUv1NJEiJtgfiE/3EUwudYAPOIo9IzhY1xmDmCHOA3mAY3hzHehwJnEmTayyTq69KKYwpF2X4
lIJhM09dwJlpyRuxcJaWqVYOPWYfd84FX6c9HSlOZgGKx89nB0jz6aTVU0TL93bG54b7HXVTv1YF
UI6sGNkp6XVuIcH4K+HSwY5R2weL92EtQhOJhbzUqAzAR60ZZCRDhgTyJzj62B55ghXI7rRwmJwX
MuK/n18wiXSGbAyDZLEJ+c0PFFYo3jC85Rurc1yRcSh6mAYLmnVdlRORhsA6ANO/sXkeVSS7nuME
njSzwuXGc167Bm+Qs+55zlsK/uIlAkvPKK0ZPkUjDgGVy2xIv5rpCKOLW1ZH2eEq9qjc9IhvgkYS
JrvCr3rqC9wesjhq6hci0yIiTyxn+qMVY+d7/IzTdB6ccrqV23ULqOjBOgVWDPNHQudDdMbucYaz
YbF+oTFG00VNM8OcH7GU+VAnDzdPfzssjIi9OBh3KDE5wQalsZtbggg4EfTP07G0qTfDgv7Y7NRS
RMhNcABN1Ea1LWqBK0rN3nJsEIMAWDXCbATiVNPwv9EzMM/4qXVuKjv08Rcxx1vSpFfzFi7QKFHl
NjmteOTmDGOigRS4TBKCJyQrw3y9zl+AT1RxLSf3RI3BKeGJZgTnP8zjvhnoToOgWBS1eLD9Rvlz
6ZciCwSEGti4H0YuSp6jdzAOKdBVzj7MJ5g6voL8jJZ5D2ABOUYJpxgwr2UU9XjLzpXrPWD3wq12
NUPFr2gvhKU2TLSsOJ/E5ml/ee1HUTvuz0He1dP3Ncu7UzAWAzZs4bF2XZlQe0wosZEnAWyqGPbh
ulwdLXKZ64lQZluBkmceDtoix9VjDcOQkASBKcuWMSjv4ARF/m6e6Hgn1S1cMMTx1gcKiNaOgAAb
GUra62NUJHxQ1P4tJu7FmhoRcDbkaoCHXh9zHIVgRbK7IyZBnWUw68Nt33DJ+sgtc9rKH8+6ZS4B
h1UQs7uBhRgj2vpaKveMW4FUcymTaP9d2AStMMQSm2G+P8VtnvkwM4QLd4wzDxSGeb02Eaofl6MO
0gJ1AVhafzMrtFCR893zQF/1h6cgWDLDDJzPvBvXbqTxpzQ0EFGljyDiPOhkcq2f/CsT81/PEZf5
WLEb5PoywywdBh8Pu5BZ7ZpssvUShk0mXf6IJ3jStXwF3KyvJdRoF3ifDy/jM1n4WSgKWUWZWdu+
iTeQObYmrboEVV79O41s+iBDKLMrHddkoBE1UvxnF4Himo6twVjJdVzprssrKxV4YNJApJ6Z00Ng
KWbaKE2xDWHWm8KSYoxLvls/QaOd+kQ8ckU9XYYgAq0gM5Qzff5I4nxC/FjL5POZsF8HsO/fAGOt
JX+l5UW+SoNjLzA+JVgQe71SAfNKCM/r9dVqLjmhgvLWvc+r+gxdsxAazGiDqPM0qlZ1IvXBPPAQ
dqF8LVsfJo0/FU8AAwvJ1AQCqVAFA9X4xui6OHg0YoW7t00ZIuA72tfDC/GwhPcnQoyWvsfsXQSh
O+gWLirBrmcxSfcuTfrZ+dZy5mz+cgtqKB2wEueBNwoun+ChDkeu1zK/FQ7MHLq0lUlUdLni52mO
z6sOt+tn/2zBFpMC2kUsUNFoTwJHi5UsHMu9DGVlYfREvspgE+dgJvGybh8NRCzjSAZ+p9d0ubf/
cGmHFErkH+tJUqNH8VwlEKSGaPz/i2o6IyLuqgoZKSwFniMvYb4HqF6UB7KHi7cABX2K8DzDXW1w
5kTC+eVw0jHqew0fh/eI9JmpSGlv2tHqKc1fD9eqdB+DUYHu7t1NuSeaPiyA6CVlx2rCxzbwwd6Z
d1oTcgnFUNVwNsJL3YrnH0PuN+1eJnX4Ne184cpCBnwf1G3pRZYLE/ZidNIa+sS5liS3x2IrK35M
t4LsvjBy2ts0h4CaPXLu2YM7/6E658f0zaboINpDTms+UDinJd2JaL3RKjT6wQ7yT2oCzfBXESs1
yWAN2c3u5G42QsaaxdM5IJNO3BhLAL+PrmanvaRgeQJE8r2t2QHzO5rPy3boKM1Ot5f8IO0hUXhL
79xQIPtrnUgrHJTxnuVKDU1RCwtwa7NSk+wkc8nPsFsBJb6ErmTtGQE4LzkBlBiBeDRnUEBc0YH3
eiXfIjy7ci3NJYCXovoDAe2FPisUvRNGji0lDuAfm2jU0w5xx04rwvco1Kvi+GVfZ5n14UbOAEMu
OfNh0lW0Fuizz2Nw2ANpMmCM0CJszbQrHgxyzhCla8NzfSBPC/TQVybd0XfR1bycqY6f+twXE1ei
iROiPAijA09emT2JszrlwwIN1+MD08FLcSa5HEWfPnBVOuKXbdli+IQwvS2Cx8KglIJePMFUFiLu
OI/VEDwaer7hPjRpLCUb3psCi0l0au/aLG/FdAoZta+DmaC4/g4f8VBUrmv7EIg0WKatRMDzMTXd
PjMmtxeWEWqMaj7+MgAQ/M06SuEn0pZH3cSm9tIdzXnmqWLfEEJs7Niz53q0uHyJ7nzSnoVklRzC
3RJqhnjt7h4KkkKkFh5uf717LP7sMjl1iHEgTpknpvsZ0+tqpSkKPlUasrntBn+rZetXVMYal0Fo
3EQiSVu5CUVuHNUvIsZwSy0u7WIwDBKjI1Z14Pdhrv6PRWh9hZQ27NdvvmjuBu10pQNH0wMhDIDE
ea97KA1QFDWtkSnHkCB9d3lNBKfB8IYd9A/aAlC5L78KjIXbLtmiqG6dV5h5g6jtNOLkLA5Gx640
1+NcEIgudCSb5svrHOVL6AzwoOKxep+QCS6/Svaa14XsbcuoVB1B95RO49P6CWsq+q6GHzXNqzKi
jqBF76LjtDcF8izWGar72pUAL23ShtiPv7Vjx9eX/2h7zi38tu2bv5afGEW7g4LnUXxdDJ0WF68g
fi/4CtB/o3E8kS2pdvnW6S+Eywc/PpM8uU1roivQkg77YIOVTLRAqv6CR0isFphyYWJk+VXGZ03W
HQk62ylpuNzRfq2K72PpbkAfZW9DTEzxqBTlziU691Y+jUokzbVu/ERFsAtxCP/DLxR1BN6jCvr2
cU5FYcs4uvXlOLw7cyU3oMv9B9eKci3m1JzyMdyndtcVvtqYN1Yio6jCS+NApMspPhlplw6JS/9D
CdOGR+3COos0Xh7zBh6DNoRtvBQLJBT5AuE/9MPmjQZqQgsFx/rhEjyegM+bl2sQTKiuP8q6k3Hr
Y0KVx3v16mwNdgYFhHSh+WwKBfppMP21vyv9kzntMrhVYsbzhpXWPNaYh4PAoQF5lRo57ryjvgo6
Ps9xrSHJkRK+s466oyj80/o4Nh8Xvd3yaFPQELQOfpbTEl37VrB9NMT3enr7rn9ltOGcVxBi7Rlm
Bx1CekvEyTPgEKinrUf1rmPafKCXlY50tuEBDSwru5xJ4AO3c+8Iol67fIUeSG/CUbPcZoPjKEa/
4bf2QuIV6AQF3/XRDtx+dNbYcjJo6987MU/aNKQ4c/oEAMVz/C4b7v3+s2FyvouywWBjmYgDAVZb
ivLH8gQLW5T7fbBhoODzJBUsxKFqhw0jheyAVuWfpHOG2dvtEg521X5zmAs/8hpJlxG/eS6MDEdu
EM5ejVv8JU9L2aGzYqh36rOBWpW4vxSOavoyC31vfmSs5agEd2ouof+A+xon8g1eTgKITiM/BK83
EJ3yL8NetKVVObhy/Hj3JE1BR1ADR21IM84SOaohHpRrqFyC5EgcnbUKmdHvZsZHXlxUJOhYuYS/
pnTnMLp5BI7jX51DWP36VCb6UREJpfqA7Jh0xgWikXFBGN26Y++jRanmZwZ1UwysZOQVukzStfgV
b2mH6Z3aIr/8IClw2J1VWdaaJSVCz3CSgergsZ/FyByn3X/NQTqXctBqSdaemGvF37oome67D+Wx
koZAhrgRE3oqZcYakJNRbMnw9K+RWI80JCxeLOMqiTX+g/shXtY5/YjtB+6iKKYbvD02ign3YdiM
85M7NEgkAtynRUTkI8R/gjTC4mYM2Pke9JaeOiUA05eM6Z7aC6BU/SWZnL/CKIbAMMz+czvTi8SD
4TuZhZJH7nrNqfqOAmg/Dyac9MKdmE+1IM2pOUqpQbWdC4C3AHlDZExu6wUnUZNOmwKBQygYYvHJ
ht6c+lLg0d6K8+p2KodLfHXa8fAD784Cu7Ac47v3sn06gQJ9LKOjSUG4+myhsB9GMMYwpX/obgHY
Jway/zO7zyhQy38H3OwQJsGKb2wuJjuJM0W67hWGJx+th76tRjxYjeJ7GuuLANkde7Fr8uCbSVda
gsl9dcGa+dPviR/77GMHTFDOKdBqnWjonRtR2BIZXZOtYV8ukNZ2HkqzNHOrsZCPSY52//jMlHiI
8y0P6mqj/BEWCcq8FhPyWJ+H4Ni4cdsRYyJWyf/m7zC63FADgk7l/PSFM2GvDQyahbXkUctTk0PT
XVLE3YM7CPZ0Sa/s+OGSILuU/GJqyaJw29A7Dj22X1E0GZAFJyz8h6Zeab3L09FaSAqUlHwPOAVg
R9yU6YzVn2H6J+7WC7PZ+sQc1RmRlpKDk4sveXpdsfkNRnOtNUsbolXHlalKnCPXbLikfBNh+kpa
pIJu4BTFZQhiODgLo40gY8rHkCOs6KSMEQIYB3Bmdz1xuGZJttPVt7jSyBc3rZxKzJoW2TlQ5jy6
n7hvSz3nmbYhmiGgt3JXm52d36K6noIIaTQpwGPIEdW+zAX0yEG4+QhpcXbGM/OFptnuWnGF8RNu
IxBMfIMd2EVwO0ILB/hzt2WG/mDfP6JGDVIWMLFGY9Ea6I5K4v8OFezG5IaIHBT4H0q/5gn3X5uy
QdPfY8mgJ1No1xmDE9ok5l6Pzr1fIn3el5y1ZmBHa4n/Eg3WhRRkaW9akkJLkSRZWSsx9Dp/hYXs
Z5hNEVZhZRocsS2S4ot0v4XNYsX/rTKfH7PijOtFN78vyuDLGHcoahC9Dh9KmWMSkpUsC1558Fy9
RAD61ebTzkpKuRSdHTQqjHlnuNr98L5j0N9jRadjXhfjCViSorvfOWBTNFF7+6AAtWdDi2a4jJ7r
3qY2C2psIFHr6FuucKiQTkQkb2fakzULoWLmW802uUroGNjyJ8vlzYdVM+r4r+xcNlqn2sql9WdI
CddYwGYNnTVZkvAnSlGw3+Dnx7AQ+8jc+0MTW7JYE8QvkIr+cmtulUvFFSvD7mPOd3PmmyRywyyF
b0t3WJ4JlmP4u1r0US+Kx1TKC0dqcWzTOSGcomsFkYrRY4DOgVcvoG/pm3cbZa8eYqEirzKKGdMC
bg3ttI8iUPCeFWfIFs5BGxA6YP/nVtJU8UsVguVsM/vrw0UpHRQ3zUXkCM01ySsFY3MFs1APzMG/
HwO/6EH1IM2jD44ucMxzHRf9n2GU5FBqF0bLjBLVipSVwzUdqGAN4frKilaFxt6eYQCS+BWElZ6c
6xMlEUXFc/mxMofISstq6ebo8Bp10afTaxma4GgMp5gvBcIGLBvWD/cEKwtsFDsMGIuiVObhZfuW
LbId1djLVoXFtmMrmLzuEKZN+PA3dUYcvrZ/FjCcP0nLFhqu99s3Bsscn63dkp/tEqINk14NHOj+
6YTN6Khinr7RJxmO7n7UQ5BlyQoSoSRboGZ7wxGJeWFuwR0B2vt7L5iG62wEjYitumiL50fTlrnN
IPkBJhTH7n/FwjIV8kdVG2tES8CoFWQcdKfHx2Lz2NDjhuLlxz2IFmV0s1x0h+AG557qSSz34muN
fLVwSCKTLy4QvPT5nLYN0vINr49ARShaue8quD89SsvNyeWPoe2cptryF905ocuybG0uViRGwTSg
wE8+Jb2DDUsS+wY5kb7dSdUznFpw3y4vl6DqvP2xvcLUMtoefpv8cbcs7laEw0REH2jTTnTKkV4F
Om+K8nhjuu/RPfIrqV+LlaJMtOiOFeFaAl6tWl9Frz8B1wVBtuRjiOAU7dUCLydJqeLhaQ5kuHbI
XvGvY89kteUBXMh9WfCXMtME34YCFNjUrIUyUAAnlSXm5PErqiwgpZ7nWtPZWvX7hj3T20ME6v6i
6ra3vjapSVea0KSUDbQqI5OD25WKyjzWuZGXwa2ov7jNTtLiHs+Tw3h2Ho/Lo2jBvw8cek/7ouAU
XZqrziglnLlXYZ5ieiA+fsRT7r7B+rbA5G6QKIcO8qtws6Sryzs1D67tIjDSXeIk/AfiMVtyWbDv
o285NqeQMltlOJYC23SVCW0tWQfBAO2bnDf2htQbAlMLqSrZWXV0D5YmabB/C9UaDva32s6OaH4R
uQ1ZBlCQzvst/flODdGaqPPn/UqlumEIpTJWHORcdgV0uelzRVpARdGZGrjzdSsBS/KXf8rhqchA
5zBZ8XGVzIQBud4QLV5KxAp5wScZ4IAWmF/xRoIGNGkRclWSokt997cVM7pdkUElD8980XmeFgOP
fGbzqg2YhCD3r5w8Mr44qgH3FbhSOwd/686quoNH39b8KS0OnQni1tnkMTwNIZVIz1WrpByrtBir
7+uoKUfh7e7+LKi1TeffoczPxpPHq2UoPNhIhaNcjexmiZOqrom5RKME6slomAydsmxmv/4koEFT
rWEjinE9cHjflnh2i6lTJKyXhaMjv569aAmEG+OuLFc2+MOK+PQLZCSed9h6D3pVAimy/696Gpte
vs7PQ0Q/e9dK5VGZ6hlfPyuZ+DP90cd99BL6TclHmYqVzr0DCPEY8gNAsLIDjXNlM+g+T/jE0Q3R
52Y/6jTrdYKZX9ELmKfvD/icbQM6bDYjMrsURfR1gzuEm0lQsSNw2jlM+7El8TMxIc4kWhGFgOxt
NkwGx/8BLi3zYQ2AaLDIvrgcp1b4ShRhYD9bHj0xWE6b7347J6FjpnzAdFlr0eFVXlOL3ore8N/O
AU7r743E4Jk7cRiC8m6DLaadPFV4D4oJt8dWaornTCQkdB0dKCVgy2khnkBunhCpaIV/bICsD0nV
/YLpeIfQZGH2kr+7CPcGAa2duq7SfjgshfLO46X8+bVFRzCR8Gb0XTYBB/Hc5T938HGPbAhGsWdP
62hobUIBnA5btKpyPtUX5A9D79ZvtrEsHWbK2tzjvfu+e7bwf/TnExDCkFNfQnwnE0tKSo9qOlZj
ncvg74nlfN6ZVxo+qb2vuKNRViSPVvzPFykXYDDRQOE/U/UOBOh3sFj5cM7cdNExUrtW2bQx4sVG
xJBclQXpmMT4vJa+Ylw8sgKBRrakq913H2X0P12tm72NI3JrU50sVWz+gjga9UbEU3C5g0llkUT2
WtVCZUYdDE2bTgW57n82sJrnLs+wEii3hgIYCJ7pNY3SKGEvLfxzvsEJF41K4mXB68mMuoj+uRtE
Ms92IFK+kNVM4j7OajguC0krX8wGW/gHhD5cBxj5vyWFqt7zUornqfmcN0tXdbaXjJa4nqw43nD6
3Yt4ro2YiYUkqIiGG2WpLCAYbrZkFCVjmx8tlfmO27RaGuHkad91wj4FpRL69/LOth+6uM9+Cog7
NirFxTyot8WRxMUz2dksQpG7lTc8jS8+wwAyrc+h4xPFbmmp6vTRc7FV2H9XuPmXR9GjxnnhEjdz
wpuj7xtBjrlDLMv7/Ie6qk7Zc1ValHndTDQQYEUnEfQXx8foTL8X7b1rdqfMNdF1VWCySZcjw/HF
17PPKmxQD8oyb1yB8FU1unfMZTdSGgjp5FsI5IpEQtjCypFPdggFSkbvq9BU/BWBBjOWstAYpWPF
shd1Am9QZcjeHfHMY1aYjbyVBcMsh9KXZGKp2J8UKi0B8e7yeIBSO8RW11xyShLIld6TvEhbfZo1
Hhpv8gdgDt8jHp1LhnzfMy7CHXW1WEmdEMdiBXtLF0GCD7t7MjMHGX1BjwtOui2TVB4StcTr2nFU
k6KsN10J97Kq6FnYRBeSgc9DiH/SYBfV8DsyRKXC9Mj14OuaevhHMYXIcjCEN/tzCswo4F+LYBOP
vgw9VjXd5/pIH6/lV9UDmJotnHG59bpPf4ca/c+nRuNe0e4mr7fi1POs268suYeNU91gghKmr2cP
+Z52iuVGwFI2nZKKc26LH1YUd5e9ho8QGgejCdYDDu+boLDL6X0ilIz2ymBfEBOW6027mrQGZd0A
rlkwAfYt42wh/HfeFJvwX26vEkx9Og7/9qWUbE21tUmlf8fijPTd/K6xhpTUPjF7r68t0h1nB9ah
nLSajAgrmJN6717jl77IT7oC4+EUIBnK1jbeq29fb4i4uFJ2lj60BJ9pHFkezRKXeiQ5DSj4d4h2
R0SiNaJVQfaTSvEQVe+AW6R7XqaVTQ/7CIr6bzO5xUX6nLgKO3HFCffSgEzyPrKognh1R305+QWk
UjsyG3XoYK0Nduzg6oZ4YCU59b+yaGWdlimRfU/z8fxY7l2QTBfFErkGI67HI3FzTAG/dRlrTKvf
E7IZ4JbUAo/fjyHoooOFoonA2KbElqHXEcVbKJsblYQUJe6FfkPCz+5EyF6+3gYkLX/XBTjXWv8S
guS5Itgsq7zL/DrNtUvWPk242Sre3HMYrw+5qusPoXCwAaGYe8AQDS6KdGwga8EPpB57nONsCVzc
Kg/trkazpx8Npx93tl1BkLRGhpM4SRKc0Rmz45M60F6NMv1JUYDVWGDMOkwHR7lDTB9jWWUjxEGt
grxuvkHBdryFFzoTt1TCZDlGECsycS3+nPTXEQtfHi212kQWursYXX2bYFhfkXZm8p2bgjLLNmpJ
UDtlwcDniz40uaaYStm5o7T1sl9zhR7jBNuVH46sHauMoXXEyWcxFWpxCJodZvttCewEIIWdT5ed
INA7x8y4iz65hmls0N45LLFlp8lDb3m1ZSsQRAnOzjBt3SSFOmYsth7zFfQTpocr/6ud5OM9hJnX
8+jKlCVeWt4eSMXpsuSWnamzjogpudVpoOJ4J6n+iwArv4zQZaJKBhw52JgxcBfJMOeaVmtzjSkl
v5TVRJQF2RdIeMtgEf3EOy7kkkqF1qcy4AHEM4XBSz6b4Q8v7oK2837BWAfG2eBk1bZc6SlyBvXL
vBV4RhIIPUpVPPPmRgUTsjfJwSf/H5Omza3fibgbMBYpzLh24+gkSMrSFi+fxJMKKUZbZkh6nZ+Y
V3cEDZuZDplGY5tq7RSDUOq39bnhuz1F5xo/ms8At0e8aOTzq3pXM2rqNFoYxZ+Xk3sAKF+pDaLG
G2zuhnlDyydYF8dga8WD3scvWENSQmWbu2PUCd4Xbzp7Xpv3xnFNhXUmnDRSktTYKBfp4CtHhAln
EFk7Quzio5DHRFGYodHQmg4gGKDP8uHxUhbLQR0UKs8AE08QtE+S0t0xNAJ3tQkP9Nujezzy8lOr
y4YavP/lpwxF7WSiaIylETe8wNk20CL7yPFcoWD246P7yPkKytVWHSD4yhaaIS87zi81ho/RUILQ
3C0hvx/ZfCDyC2hqsAq3fblU1MKdWNTXTWhz3oPc0ZGMHAdiBC7mi/sKC6NWEDhnq88yVRrd71aw
9WACUhdQyOuAqX0LNVdmIfmqnOW2LuSK8DbmBK/t7zNWwY7NsjLXxjLxJ+gc9LrIKBz5ToibOf3i
APaHduNOmOX5uM/YguNqqztfEYFVu7OhsCUKLNR79LVoqAH3TqQCHp5S36+AJ5u4qNwTn/5KxLAG
EuB/Hq2ky+pehgzBNQnZnSsPMmtf2D3eYHAm30vuuPZZiyebxpU3sHCl1qZwI58n8QsMlHpW4vqR
h3KoqJA/aqpk8EzIUmqKsBhU09fY3+14DbDL9Pir+LMjcBievoqGIhKZYkKYSpNYYWjYFgzPgGEN
QJ5SVuoa3GYK5bia2CFL1agajPtmrs/9MFuRMBd0k4zfQAcht7ovN/bKB53EAK0jmzwFbioI2/dQ
mAazPxdariPuxadQavG65Li9tvfYpzg0V/6V2c2coQe8AqChk/02GHkVuP53x4tejbmSCU5dX2TL
9y7yjkZakgJQVRuEeyn+sSCDPTFT7kIElx2u0H+hoGUtfsfJBVYw+94xnUoDzr3Db88Ic1LLg3LH
rNroj+lGC666gTgtQif9GFUIb5XY3PyAvkUqoiSIF2Lg56GUHnZ7sx1giL8xZzNRJBdxDiUVVL1L
N49lgYcUMY6XsJwuG0H0Jk5qZKJr3b7XxkPnI2sr/Cca+e/vPpPQhJ3z+7MNafta6tAPSDUr4eme
SX1db1NvcSjIjFjJ7EySy6tOYitxTaU0rn+xBIK0H+TJgLMUUOtmqkWi3Ss1Z1lH7HsTzeQq2KSA
DoPubmZgs3j1QUo3DYcEWip5hBEgOVSLMZglFBcK/903CQC+ASrtYNT+4sfaOKLiR/GiIL6iNWaJ
QCZSkK8xhoRTg+6LgE+BB7G7duZfXsnYgLfIfQDESjmDVHICfkRoWRrWC9pgKS/PUDS9ejPfW7ZR
SQ9hbkVWr42le1d1OyUPPoHy7Pk6hutW3oxVVm8b9Kf5X7MTzaha9AKTLoHlqzlfDcIrz9tk6rOM
md8DXzYMo5EAcIDzD+Qa9wdXCeJ/VRtdbqzkB+/RhM3q7ydKRqO9v7pD2lGylrY+5BWewEM485Bc
xNbmt9s7HxTwv3FpfFYyGC2DQla5vnRAd45vuliANewTfFKe/u2DH11PJKh++zMLCS8dzVeaGm6s
GZCe4qhw2xx9vFHghVx9fBG7iaasz4RP+iT23LZAybWOa+7nONsnPOEMVXmIABDayK+crTrGqjyQ
6BdwTPA47hMVbvn3bzRBwq8d7NFF+ld0ikXM5M0Khc7KIgoNGtBcF3LfzTfpD1QW4QHk1tW/Uqwv
HWpVGondaoBCoL07LXtHKcgZReCoMlLv1jZqsjvnln9Wwrds4hsXrB1Z7EbgP1l8IXgfzpIpoYPH
Hor9nJ+LzczWfsxwodyBzef6ZtyjazNkqJ/eLCrhwdQIrCHsQFpvxBQ3ZezTFCcZAZVx8glmkZTu
ELSYloucTN/6A+c0gL8SBJ17KCb9RdpMuO8/pThpSAR7NIzLVRLXOdAzAHwvxpVu5hJxePDeozCY
HhN3dLduJ6AWTU77j00sdye/gvNBQDM4LPKUmcGdwqtnaQETKQCEvpfoNM7AJElrIsHsOCETMECH
MqmKnGDbPbdPOKkVCxPc1/WawS8+mvyNtOv0RgxSkvIFiY9hNLmxCDZ5T3YrZPEWC4I509QQ90qK
eTRrMcbD2VwWfwkPYFo/Lv735fnYIAawZ/xp1wfPz/R6tTHjZDmsn54JWWLCVagiVArpS7hMCEeX
+sxZgrqYk0euRZbh2vKJY/XMALegFrF6QsoX1akqNQTaTP0Q1Mc3/bp3F2+62ge8Jt2ES0p0KqH8
gDcTgS1YmIfDXsOgCR8Dcx17ohE1pWc1TY6FsvXNRkdt9kHN/G9smRnTI1ap99rp9FOTf2idKT2X
sPP/ifdivc7noMXdyGOWB8a5gniQmWC36iss6bXXl17VisDv74mVqpMxx1JcjDWUSCrUIvNjWP+7
zFX0qeq7aCyNg4Ctau8iHbB0vp1GJMLMR0cl/Pldv8pCTniP3efTWVenmB6QqhZEh64P9DEcoqr7
X/yfmOiadslbaBAWnT2T5aAryP5x3qfEB2eX+iQzSwbczY/ldseEIO1t4/6aSTB+rmyiMyARjYwx
OF2qeoRoIUUB9KAT8HbnMUcJvtjlqzgrAnQjr8JH6SRw+t7Lm0ii3yZ8HsDgePi2bI7Ejpx3gr8r
9BZgQW8QSaRYd95PE7L6e1aQTYQubGa6D/ND/jsw4A16gmrv4n/l4OMCKDc55CZevG++iuXW0b1D
DXBWfoCkXtg+IlwQCIfEkxc5PFmWab+lDaWlXGSH4b9kEBn/EnDol9+1lDn/gDKHLV3HT6oNEpqu
O+Kx4rtnXjG1y2EmMZcYAKgthBxYns5wagg8JUXZQOZcwh6fLsp5jP3QDtz1FmvcedEp/zvxT73+
+wzBiao9v7CKZ7m/RHZ0F4Lxgk/fbixMOZ7wfFBPodXMVfP9DiHwZG/YsQNLwszD3ruQAcIGK5f3
Xb27jKxcRjtQQuvsA3AunjlrI18lFN/yIuY30rqfp1woqLETOeKzFj4WoAmaVcTobNXCYdhhxpgT
GgFoxE45Bgzl1PmJ1h5uKDNmX1xLHtRooZHN//nJ41v7wy/vQH6/E0uCS8UdAmISEKc1jk0GZzSS
wkHTif3a2WOWDvb/NJM8nBw7sPK1qThhvWoJwzc8TNyMZvbHJRq0s5a95AnQ7rk1uLnOTVJp1p9B
lI2Dpt+4X8upkf73Q8RVCBDquDbw8zsJv5LfEKLaWvz0zhr8/OkEwTnjQSnI/71o1ZC3vw579M+R
fs98aT8kQvRP28Gpc6V8STJI4oomNj6VjERW82fXUsYNLYOvSBTgh2WvJj8NC8Xi2JhNrSEndPOC
YDvHWm+xkrVxyHtTHUT0q9YygqfOm3rAY96IsGSZCRUDWmU9S9juyv0B37PODIq/4XGD4a0J0MDM
Sl8CRPaEtdJQBZhuMlZZJJhpIw7kTAu2p1bZfbgCtKVEzl5lkYQGMGgse7idAW5Q3zGr1Bm8428d
13dCdmo4JLZf/XK4p4s+BwUa/zdL74SQD8/YAFT8DpUO6Jo/D2ssQgVATZMay8o0N+JOnAuXU3PZ
S+E0eWYFQjTZ1fpK9l85V5VRsOWG9IF24Tue4Xwx7v4v5aXzcTBZF7NzhuW0AlfomPux+d3ff6wr
SVP+jNDkIh8WzeYOz/r1dasfkcNUsl5atdtXoJgSWMUZlnoK51pzQnqz0plsG0urK3kt05TWavyj
yK+BGe6JFZh0qFxdcOQpA5Qar05woDsppwGk8qvM/Zoh9/D8f5mozOFkeq9O6t4wHMQKc4Ri0LuQ
YVXeZ462Ka8+l1l396E7luQzMr5OEDpEtk5HP/QB1VQtcjbNshb5FJB/InPbP+fsGbIW1MuyiqZl
iNHrcNM4lMrZLu3/aabQP4NvBFgqtDxBuZYrlxZAvGaL5pIevSbllp+6w3tABx2Tj2hMNBlKxwnW
9i2f12H2jrOTMKv2nbYGeQlnyvbLVzlD2R3HkCKqbzMFUW91pZciu4oIIhHDW+mRTcXv5yfp4Xm7
ioWJS1nSgJpu1O8z/GmyhKx/QJ+2/JVWV1ZggkEH4dTSgBbWMapn1oO2lwpJKyT/Qj5DMMqXcEkn
S/XKH+gzmPjkQzHZuKA6kQ8AuwZP7q/BhjxVMUx2/fGkKzWJHbt1ET4tdhdni5y6c4omIAP+8cOa
4nYxv5oOxI/1V7uQQRdn7GYAmWw8q8BWKm8oSn6gZi/kW/EtQ8QwxL6ie9NrpBBLoxsgNcQkqZw0
2Q+U1NAlYmRxF9d7+0kCM6suaF5WcrWaS6T3Qx/hcokn7QkJr1+SYzpa8mhGOphfYaITZbHZA8Zq
Q3MmcuBQZ+UnIElt+QlHZ4fm5RvX98CpXoPSSU0beF0LPPdyC4UGounFeXKpzUa0hRdOX5BfBM3h
kXgumdtD/7RD57PXMAVV6EWJpimGS5dtB93sSF8ftZgIW/Usc1T+OBBhOM38890Idw3OS0OtutRk
29V90ZIdONRLmIRJTohXFS6wUQlVTm2pE8xB/YGCTvd3303H4+0uimPKjHB4ZuaVvgMR6M6DC92x
FMohfrvLH9xjL3jZk8RyCjLXhDnqDOT2WSdIRd3AWDBtZEXzXFmbqJ/F5R6+SWM8Hcg2vIQpqGK4
uwe207cSS6l+jKA1UidUwnm/nfoliP1kTBpYbEMKXsxOGbSK3m6CpvlhevamQgfwy5KT4xmHKoow
TuIa6GZWTSKjRXYAtd8TmNHv719x16s60u7fxiGWYLKHZU4RyKVokF7IR6wN38gZllz94tDfmcb9
/8WTuExcuZM/QNs71ljKuYkzG3xuj7N2BlWx7ELPqj5UBmf2CBOc53s8N7JjcDJUmIV4Ljyv+vN8
Xc2XstkbpJYL5y6TznAvTSMSGL6t6I2e5FZpnmfByNF4PAkGGoF7UD/ghw4ODrdcmHR0rVvwtlNk
EBAref+m2z9Le1gqa53XV1uBT1x9sMfGU4dAg3D1Pif0MGq/imcwkG2vc7S1aqaZYaQD9HhLusPG
S5Kpo3LjM4NThM2ranhz/9ZcfCkcy+pf6Dl4jjY/HzpyLqd81rcl6cNw+z/MMXOg1cmtiQvYXxLu
/A9o2aJlykKEMiD35N6s1PyCpsEuxMnYCV2hwJY3O+sKI54B6+JyY5IBWh8WaJqNhvDiU3HM9Zyp
egM9wbLaqF+FFr0KHrC29BdpFuzZhcq46Fne3nDeaLmWz+Hndy95ZtFPNTl/YyuOUaFEIaF4ySGt
r+hBnqLatPF41/tbJxDwGOm6FU3aMuSjqSsFx7VJ4LZON5aCb5jbzaniUUfXZ/xSVATK/Vt8ryYX
crgsg0PBo7iwgAz54k2SEZVH7UvANYt46DuC4eFZkrgl3r69FBJw+SmTErp7BTL3Tfd7E2gVIdRz
xQiKqoKxN+HRvDlBzovQGy9o3ER3dt5IiTpxS2Ue2RSb4XXVaUS5J01kQWVtGhVYGHo456XU+kzt
vES0t2aiksTnnlacLFQWVis5SW29amI3oFQqQkvCa28td+OOLN1DdqbGL9yqkOA3XctrH1kVh6HB
55OIOWflm6auuKzr/K9d+K357/aAk+J+T0HKF2upIEseOiLif0gop7h4PTAFnAtNJApjZPawB789
jRhI5u5f2qT7BKE3eYCWXDI6+atuJQs1wsrAlVz0yynmBIzcErhZwD4gAQd3I0ullyRUzNJHHNCu
vk8NiUuI0SBb16rpkW8rbm+afSJ8yDpfhXj3cLDy2x7ItU1Kbv/liwxwdNM/DiiLJQ8IUPcBDGzC
lfu63vJfzE5Q7imZS7QGXhj+Rf1KNvT2E2+nYUq3Fr08VJpETHMK4FqRSNfGtbRfE0ynP4f84yKL
8G0qeztwuzujh4rGPutE5flFVMiByUF3YAzGF7zH1/W6M1oge1oY1LfHG1kphVj+zKlsWAH0A0aZ
Ot3HR9Z6b1JFve/0pQdfFXivTVQ8iJJQ/bL8KEyjaxEh7hDx7a6CAB+ZGDLMiwC/nRrXjdqGPBTs
jK70iQhOV3ZEEQGT/nKQAhiu5d8r/B9u9Zi+KAA81JvL3ccAa6Q3DSwr+NqFyvNlbIKsQdflsfi9
D5/biT1qLNXHLqRTUJm6K89yLw/HjJ4GPGzD01wqkxLZaGh+wHm50bsxLoeI2QV67ot5IN8PHqCp
4pyaXyXVkpvSbnL8IfRvA1qsW7Hc6A9dJTtg0FmEoWN7r3kdPFteRq3oRJKD51JA0Lho94w7AVQY
GRmj3ifYwwD+9T/OLvsD9Zturoerig6ta5NpeSZhOOV40/xByXpw/2yxgj1ZJCbxJ0aY6/nzHQ6a
i5R7ZywH3bUFyDITHtuLJZD5VCIuqGXTx11EnLXj4GK2fV8/PkY9Fvb8NJXH94BnoZkIjxwkehJl
iU6/i6itRTpbMTk1r+Pq6CyQE9OYYzaFPiP1OuyWSzQicEiJB+SQJMFG4xAU7TlaIT5yc/90DbBe
pB+SKaGtvvdAvajY7pinit1xszFqmIUsQNvC6vN+0bfea2ZiNZ1pvErWCknhrIeDBR/ueyU1BaII
BwLt6nTCk46QAM4fHOE4D2w7n4Q/XshePvsLwYc52ITx4cWL3qPZS0fZv78QdVgGO4bjAypRDo9E
iueXlGoMF2jiocIqKz/aHR4IJf9W8fWjVsYgehLGtnQnN0339wOljrXtQCCkuLB3/URCv3vHa3Ub
vj4U8OOh+zyiQgS/n5dJOKa2xkLlkSXICAnb0JPVUMeJWMQ2/pulrATJVbRMm5NcwqirVuuABo4+
z5f6+7hpWvT3BJt4I7Rv9XHCMHAw8J9inwNM2B5bLLWL45g5AcJZ1Rz8M85XRInF+DgP69qFA8i0
9XL20ZUBMQZ40P5RTT2P7/zGI4Kqx8XHztGJ8UFkIEHIE+LXVmVGzZtADX3xPb+g5ZDIC4CJsTeS
DRDng3I+1LxuhRnd2QHmGDC9xOwEs9VTrXJl51o21Bv5KmqXhtP3fikmZAhFKtUqXES1Wp4ojw3Z
Bj0fGYXaKNscTRHkKa7QTtfJPnxmAlR7fCfADlL4/NQF8vhGDlgGt+UQnL5372HpoqoHnctXVG4+
x072zHM2HW9r+sIeiR/l2oXlCK5vovOueQ+l4AzuAt4dUb/HATIsGSBwbETa4L6h8MJBhJUKz4Yh
LfLNbzvBV8Z9kkZf3/gA9wGMBXElFNrVrgduruPCDlbMzL7eWMFkBeoOdYUeKSgoDoRDxHbFKxg4
0JyzPrCBj2gMZrW9Snz+tDxmGVwwlcxAuXVz4/IhdzClZJH6XeUsBcZZxsfkuI+e5AmDD82JLQIC
5FhDO3BoXeaALdnVObrUWekcRNZsqKGsWN6aPafMUefQHfU7fATQj/H5ZcastJUBnpziEtyoScaB
nl6QtNmwQQra27LOd7eSuaLyiIBGT7LAqq3HN1iKLsIhkjEMLjT/3uTX2/K9kmzQEuN/axtXPkkg
RkwHm9ydTdJtW8lRedaes+jbhbc7BCWdTKQJ7Wi5og7tClpppLl7k3jvRd8Tbgi/QAXKTLA03NvX
nMxYxlT4JD426FR8cRLxoE2lGWHyU24bMf1MlE8j9EYF1YenTyp5hZYBSAfALWBKtQUCUw8htLCE
5oIrOeB41KgsdJ16tchvQI7NMBgcWIUCgQaF91DCO22LZ4vnJs2IxFwYp1Pjhw/Kzzvi229imwxT
APMtoc+FP7P36WZIZjz61MtjxvsBOG9wfZdazKSD5L/hWKe3b/aAPZWalFtjwVZSGP5gIGHUc/BA
26es6estSSx+qa8eZltAW5Ss+B0cL2/6GDWC5JsJq4co5+hlFJNw6HLIFSGqQPqp1RvH14Ilaoon
oyM2og/rz7+4yODk0Bn6OVZnYp3ip/pHWyRvFtKiBlwbaGfSQnoiVZ4VB80rzfo7A//QoNfBWvD7
PMWA0R0MbwmIKxGXV9pyVmkvt/pOl+wNOUHrsyAlhZAjOMYY3wTYe4dblqy69jLYlswm+t6yujhh
IoRtppVlhc8A3/o5hEV9RUImdhWjXWStLxtoXFl7mcYc3z//MsDSPoBIKVubge0G2OJQ98NorArq
s/W7Q/bkFj5qh9CmVOuTdzC9D1GncDBE8h4gWGTO2PipU/NhGEYgCFJ1g1FPIx4RztBpttjTkcy6
aRWKoFWo7HnQ7JpCcmiw8rbXFi93K+Cfn1S0ST8Ve1xuXkBwkM1lbcOW2djjYESI0zu2WejGYza8
+ABuAyn3JUgDJ1aURFgrS0xOQ085BzM4ux+3cnXoJxqowz8Y02hE/a0dNgSCZ+bSWgu/V/3nufrG
kPNeZG7qJr07sfoR/lukqDPDDX3vN5jL6Bk8XdY5naX6KjerSy/GbVzoy/Ogq6cnxSUfHWnU3+5T
4iI43v6tUx9gEX9ErahPZ24GtRSyoW0o7quE8lz6kprTwp/TurCj7NGdX5wO0LaG+XrWTI8fl3xm
YG5jSDQ0RTHhSHzRZn5cZcGPBdfqFDHLDJltLR6m/bJKfD+5qsDg0dITcJEc3vBzxvrN1Q8xJtfH
QwfECGEMn8EjyPHLg6D19Tzt43wj3+edYZPrfg52YUqhFc5mNSY+KFDeAvfA3HrO5pDfIQSjayid
y/IB1080DIEkZMUlUl2lUBYqURwO5FSGR5Pu83Lo7YUcuiwqCxRdn5j9/v2ux85++i3YAABxt0nG
SwENyrpy57dyn4dF/KJJTP++iJrTbsKveEN3+pnLp+jtkns765LI56sAplUaz8I1LyxTsJhphoyV
ESkQUci4bb3N4ayjgUQ2Vn7DLJseziLiQvBpl5EOLccBLPqLkmTDH1F3N8iqwex431BPgDWBECL3
eyhR/HCT+rlIef0L8gItwwZFFwiqRihr1WcHM0p+DsT6RvFvdFnpgGvO586H1l/zSUjKjGQhSjdO
qqciAGO+DEg2AL0rcjn6azkFk9W/UMkBhwyoz+JPA/STBZ5POktX8o5GknGrkcW8WEmN0dV3hyeZ
NlUEv6FK360qJfLkReYflGCrawL6jOK3B+3u+m8tWmsVCEgodu8wdC6JI/Iln6qhCDlCZn7QATVs
Vb6HXNR3eJMz6nAbej0qehtD+vdeeWf0AyGRCRe65/TXNHCBxgd4iF7W82CLF5s3P53NRIqYtI3I
JyUcHR7jRjukqyXNMCiPn7N5Z4tgMMh+sdDYG0CyzaEvIi9laktxGjHI/7hGMekRPKb13PoaURlx
gxnA/GTo2m4c9qwVtJUmAdrMOskmazBNCFwaWc5IqFgfjkwNqtbzW6BPVIo0KIJC4z4cZ5NBgtOm
ofWnBQo2UuYKLXxd3iFMFKCsy868cFyNgptkwj0vStUwOO+ro4DrAe/Q9FlwkrXAIjZdLsY2wABS
Q3RqPEmX5EijNeVhotfGj0NEqmRJnll1aXHxjJxIFIJ5LHSyEhauKSiIODiRU9GTi/NYbk3IqB7R
k2OLprNcoXZEgIZUYM1z4pA2WjWDMZu9Z5AL0sugdlML2q1pgqQU+XIoa7QFVFyoS3Ccj11n/1v2
UkpPvJ9tS41mWaKZMmsLBEHc6qUnx4hcXnRyVQrQMGFXPXYBbU36kid9uOBUQnErob96S3GctpPe
iRyyB3biQIYHWBzLZrB97uqaqXF/g8pIuWa3C+wRQ+bjjMW0LJ1+YNLQJN4kPpweNFqDnTkvd/9q
bAj9b9rvRsVPDiP9Xqf2wm4t6HHR3rp6ZLbsOmbhQM2zEkr271WphF/+C6BJE1EMRhlyPIk5RH6U
IMJ1VQ2buohPlzui5f38NA4QjNFKrMbbexOo2FN8l6wHG43nU0lUllVCqZ+4SmM+T0GP9vk2rWAo
RYtOuKzyDo1cn47WllB/F8HYMBQBoPPlRDfS/Xl5HfPWck/sfITU2FT46rQUk3/Kk7bAbBHYJpnH
redq7dGjy4+NDrH9R/x0ggf33O7hQS9HyTxKsE1IuazDxQR1mP7+x0FPjEb1NEMFfYsE4MMty6HC
RuPR3k8yDCxpalQTrjvPsPtMcoZWrg0vkNNROt1hiYfqjJ7vnYN1+MJy0sJJY9KrBHd5oiLYHtId
KafEkCeGVOhmWsjdi0lwFMnA4VeJ4bOyc5f70H6bx8hvGr9PH3drwKLbwkBJA6S1MH5p9PO2IeBa
jOCgfRLw0n5T712BuHa4Pd+772AyfSv6gRjixqJY8dW6Wq+nbtWoLzKIig6IHbR7cIDa3c3Haiet
RT3ml9bNif2wN2/csY410naxdmlygl5rVMqYq93Ii0RNshdhsotAMfLm/dQCAZ+y621qwFzWCXyP
QtUX5+9WA/4tQrXhcgA4s6K8x2b4LdMrIORXO/2zJlas7qkT+YPU3XOt7DiDzMdKRTR5eMz6negV
PY+F0F7JdPe2AM1WbS7j2UW9h/P7VWG+2Q3gie55jRG4L5+31rD7x/YfqhRMvdFalk+3uJlZS5ki
ld/fgcvDazjcDj9kbAXjAyU2HncVJdkDcH1PHAWcfvtEt2hHkHtNoAYDVrNpeGi39NG97hQIwQrd
aiSeZahAVgplJ0yKGJe88wUhIBE10nEkpPUtGWignboggkiR+LLRAgZaS+599KDHvp3mkkP+UmJy
KSzeybCSTh8mVpIL74yQjzIirO+KXraStw+U30daTMu80raMmTn8MATGzsoLH6w7vK9bOf4fLcj3
lKponXFsgiteoBkZKPnzlOOM3jB3k9lPwo2EWASpjH3c3k/amq7xTozffn7s5sLyZr8BgrtMGsOb
Mpt4jArPVcjHvn92OeWUqgqQCgH6Qo28FCgFSlA7s0RS4cjSz7ZmyI8/+1pbWa1waxDV6nlq+PY/
r3g55CB5hFODB+z0ZEseT7wKeeqDJJejUGCCzU5TNI51fYBkCvLmNaPh7zMdE2WVD4BI0abaFhRS
ZnF54f51dbE/sIOmqsWTfOgP/iL9ZnK9ilMSUTkXftedKuXa/tt4A/eBjYHuBE2X98D91rfh+1td
kieUFkUnLDbZSd67+Cltx0tjLrbL0YCQRgOPZlvJCZGaZimlx74u54Xax2XRg/PJB6RM8eKDseRL
EIpJuD5qSl41Dsp3JZFg9XcI0fZVzDcLVIPsd/lcHrYE91kXVZG0Urc9WmSv4k9WrUZ1soA6qCcY
rmZciZggdDoA2+HyDGuaGJR2rcYzmJjf32sGhfRslYdYPiYCPclC0hul/HlKLa7BtqNJUXYEXAje
ZSbmh8EIkY6MO888gI59rOPoiGN1VkxgkPJ8DSncd9vrB2OG6QSdMlj/LpISM4PXL4qt95OBEOHA
Zvhc/Fnf/GqLl7VhWqDrzKf3dz1sYCrvDUIsRriEQx4qFRimqWbGFHtn0tLgb3BM7FYh8lv2GL7o
qZkLXUPQ5C4yZszdLGIq9DkgCDSJXtg1Dc4eAKtVeZs8H41TH80ErBoWZ6nb83czF1ccwbwAyiqs
lXepXGCNv7dqK/4zVt+D9zFXJlRmNdylTb/glMArvFk3nPndsk51F+Z2d4rqqy35uru8+xLW9OBc
/sopaORdO+TjSRsAZwRY96xvTK1JMTpYxHO1jPXyO1mFvTIH5diuXkpwQK6p1ihgcXLaGH7NG7Uo
46iE+/IgyU8lDupyBmwPHTuBVoN6zA9er6cVFz2WiL5mY2ly3ACHC73hd/A9qZY7ST+GkdfL03fg
voPzsRfsp9DY5vRN4J2uaB//o+OFiIP9bi67e+m/2ag4MTzu0NEYbmwGy1hEs+g0sRN3AnTH8L//
CHlQfH5/y5QEHDW3bi28RLBy0pCFgcywKxEEpUSXNl5t2DO1YYoBVR8DiFdTEd2al/tvy9ZLIc9v
nKttN6KWp+BkjpwCwNv0PKQdFdijjHkXwnpwUYcM9hFg5M8eimNAyo8F6XpTK2asCsyGbSjDRKJ4
DH1I9Ui/jyHdvCruaH5ZBf6SpwndxF/cEkwZ5dh1Vj2C7SjApGXyDHiKQ2gFGzKwKXp33sPh4rsT
4wAB/jMJgv0Y2TZyzLOIzcN5k0C4iYMw83V6Yw/J3rtiDTvPxwirBQUdEkZjvvB6iU9o4tzL7pF4
2ol5uHwKQVZbTvW+u2Vq/7StAQX/H89FAYaJZ+qSkaLP0yReIMJn2kUDtl9ozK/lnddpGmBOrjtd
604ekcNaqGHppQ0pfQfMZn3QuEr5cy7UHtQzMt18gtLfDjkj9f58lLbG3TYiiOf0SWDnP/K17kT8
a4FG1fIc+2hIzd4h80Hghshf3ywPRN0IpEyB7yfkVuu5TKCVKK4M3heNEuUXAJJzWMhIN44pOjw8
b3AcmFPS3upR8Hw9og6tjQLkgISRjxYqsO/TeTDMBscIwRXaoxF77XY/dG/NnGeVLxOsLqWaDg1T
eLvQB3zR2PkPxPurXaPxDZDXQTYC3si7sURevxx3RpTPDp3Gt9Stz6nPCzcHqo44/WKluR8tYCJT
pDAr0ddcCzNN5nGuGvnOVK38Yj82mEQH79OHtUyWGbiFNcvoSYZVa9AgatTqIL3L3nbBqnn2Wc/q
tx1xf0sAFM4YsIMBhooAO9HrpiiNHBSsJeKIZHBXUIoF+bTQs8Lu3d3BKeP23dZvqA/tFHC8vrBX
ynbllLE2jMZNLQ0WuMZuyW81hGA13J43xPLUtuzZG3o6Mzog7TePXkSm6/KCgzoN7PQjOGwlwNAB
Gv2qwl8lcjjnQb9cRIiNuJOwy4ybihsCNEU8gOwSzZw4cYpZUN2Y0cg228E7J/oeeMGVcwYumuOW
gpqIOKBEuvekP/wITWKj/NIao/TGEqqi2JJax6STCCr8TpobQ+Nj6HRZsBShUKJQiNmWox3GVfQs
HuH7DvCGXe6bstrn934UN+Psg1UvG/eF6xjLMoMxbkYLRPmCLOGO47WHHaK9DmRQX5HnSlxIpAOq
IZTP//33M0kH/nSTwhvuKM6UWqRw1IXoGDWkgeYMx0L5pAb71VAZWUyQKVy3+XzE1ZDViAFRo4Wa
0YrZrO8yktbhXuc1Yqe5vmWGzfqdlpIU0Jm25nL6kh1veA82GilRJ9E2j51uEomcNh7/CdW8DDfa
xCxcWkzbdWx/8kmJ9pDvk6ce5eYZEaNnyg23eYW4OPwuPA5xZp1CgLPe3hgk8R3EL9BNVMQev6tB
gzcMStbk9hiaTHcTGvd10DglVNi6dbwzbvMWHjUvVbfB4LPUpXQUQdTXcVOC9EAGPcjmyEDGwyoV
EepJIm+J+T9HGFWww3TGCsislveN5Z6hxcXw+d70BYpT3MvMZRT2v7htSTfn4iGCt5pqrjaOj9Ks
BKfVaD9XfqnroVlcwSYNFC7ks6epR69L1VyorIxudl5NKsPAM3h7kWX7fbY5ZoSTM9SIca7Jeds2
vWfTQZj0L4M55p4ZK/yYsb8DYByKQE2haB2tJMTkSHJNIVXrnC/bdsDzt0vwNFioupkJskRAx02d
AI57V6t31uRtdVvHFYcrPyGy0D0uK2hsSgYApDfFbgGJLg87AY0UEbFvhFqXFWpYsHd7y11F70XS
HzBCBmP8NwJ6AA72+vVhUe33rgtXiAqiz00/Y5CvjDkgehSMrk+/WBtFmLZyi9cZ4iCJXwLeJX3k
tc2xrPVaTYNyxBmWpmJB51LpB1romAlOeATkbM46AOa/WuIbSGAusm2r5F52x68fRs3IUlHAvony
g6+R/ZrjV7ofsbX1+aLtqCEXKRsLEjg/3VLENCpJ0IQZ+6leP2TbXgoQ2BbYhDf1sjKyKP6ZRlu5
B4ZwChBbFqMHexwF8GDffLnalXHPzlex0TBv93wOIggJTdib2s5dtzyaBMGSx1bPCw9jiYtLhzFz
llWTodd++mW/hFV6c4KchmhS0WNtdeVuXveNcoujfYB1LYbfDT/JpQBzDW+kmO8H/RYi9ItDV4Y6
mY1AnS26CUPicjD1gjmkWK41gQjqXVAv7s6T5+qTZkUluy98YVzloEyphor356ZEaqq8SKSlVQPt
GQf1aortK2DneftHA2awFBc1KMCjG437cJJCh708cH06vxiDXn562pL/lcelg99nxLlSCxdxYL5L
+UitVg46wcQRSsAXg23eGpK9Yx7c2S/GQ+dr1lPrwomYn2pxseMNnmRF5Xnz3z9W3PEuit3qxWod
2FI1+l/PvNOdXK9tujHQvbl0Wk+P/voQoQ9g+FpQuSupbEyr4i0YCKF8DFy3WGYTPShuDtWl8tbo
nx9D5aSQB9LFScbtCLefn4X29XkB3IcbUMO6DGyPDExIQcpEtuvFHlHprCgl7r8AoFEf8fh9rotD
Zj6aJmEWWxssS3J84/xvXw7ae7a8tqlnAITP3aW8WR/e1cmE1Vb8dd7upkQalbmheGK2zMt0j5DI
UgQKqS4RBiQ8RyqiJBc7TfAL9kxBKtSkego01YQt2z+DhnBTTaKfWwsK/RFORB8QGm2FRkql77aS
f6g8XdDKkhcIt5qoTMiUAtJSmZUMLoXJzeKPL6SORJNm9Gnl0oqZn8eZjJ1YvZUem+p2raaCAOU5
pEI54GXlzhZCftEGDLXbnUHXyQ+HjLImG7uxEzFF0nPRjcX/mTi4SsPBN+ynxmxTGL/3ONYd/Tby
8zufXvc8cPtzRuye0oTPY5cdhRsZdrFTGkL82k7hZPUjHlhNRSCionDbmytYvUnXynKbQFyL4UfH
jm0c5g2u4mhJxOnc3rsI0dCRBWwSdI+yHDjKkwswcAUSJxILvBI+l4WInNRxvs2wUeUYdNzF0lCV
d4d2+KHdLqbvb2T6zV7ejRMjnCVjYH8d2xQXnrZkYi+l2CJ6DveXsfoRMdTnswY7mxmStz2ZURaz
BYFUOgsqm4eY9Q6TnYbc+JtsFOvV+29Qrt3XwHtP/sfmXHtWvGfgiWC5AzlAwyQO954FQOFloUfd
Hc/IJXnNfONucuSv2lZAed285llItYCeBHg/G7TVNy5eEWcKhks/j5dtWCnc6wserhB3sZoRZzlC
DuxobicLShhx/6ocOfzsMfQaLjf7dlFHLcbYgwkzxljIPGTl/vlnaPrjsemDi+P6l/T1c+KVjr3H
NwZ0y2QOshV8mGnk2f9QbFwuNz/E6XHWpXTWlJUgWWJ03Sz37+RajJExXnB3U6VECMoytegtoz3Z
2Jtf0ZxWupSl5z71NsdhLwhA3K4fHFA8zCWdEzPJ8+lI+YKUSPcett9CSBfEcXCzkwRltiHUJcL+
Wdgo/OLv2clwlW2G0r42tb6FH5YZZh/vui2X/cBE3LffvB5f06D+FK3CPt0uj1SsoyyS1eH76fRG
KlDv/bnsPb+3QjkR7Ea6U/NxavMdUZju8Jvi+xgBEalEQXQ1u8PsH4u6Nt8Xb0s/s1qtfPaoAfk5
2OByUsM0vuI1wd34/3eIsw3xvVRKqT/IYbtO1dyypZDTKngZ7yx+V44la4FmDP6VZwQZ8ZCgZ3u0
8ImhFNZjFz71z5iscWq6zbGVzqF15tnLXLOkfoMUR5RU1KDwTOIjKF7rBjtt49yWN1au1N+2SVGq
cLsYO3nfGBzfE3hwGMnXBZdt/LcylJlz5qcM90lDpBAiVfS7RPmlpM9gvaMqfZIoFDZRC1OxDeiA
+wlp8OhsdKDQ2nyftPJqx7gPjuaEcI+Bc58TbQ2YYYwSN3b6cY1s1cWo+OxHzMql9vCvFNNGFGMN
eayftW0u/Ifn3i3pfaUhsSN5PXiNm/aPqReZAJLHoghu6SUXxB6bxZgpkg3dJf436NZGMpWsmoTE
cK1UJ32BCpLQcbtxntq5KlvNTnHUGnJYO9hW0ECBe1jjUZiBL2A99SmR3SJBOOsstemJeWFMVgE8
fe9UyrYHFgTPwuF58mk+1VtKaZvHeYTgNsGTobVcSQmfTBNZlgeH5Om8fZdyY5soUpi2CxIZ08b4
l8n6FDT8rmk1FW/kDYNMEBO8DGRDtVrJz72Rbls6ylx453LBhswouppK/fZYx+rrjqqJStIixlkt
hM7TlNZegFWCRdRhqSo/Yag2w0TIuoV+G/j6zNV2pxYAqh/+Hnh6PypoSM3Viz4VOdsQYbq2WTh0
haBNAc9+iTjHzIVtAHwuA68ancJrmubfCOfdgHXjXndpsk/hjal2uPqZONQo23ZuM2WWD/CXbf65
OHiEVRqjE1nc5Rf1OlJQ6JSuPD1hjZFI6tRMKWewIRPPI5VLyfzcC+HC4iJhPxCfuZsZACjud+MC
QL6gIlpB/W/Pu+Ufeiv6B7AA73XCWb9vIzG7W+NySoa2tNW80PHnEkAbN4REGEirL9NCi0NdA/ev
i8mhuyRfLXe6gXapTtWA6nmILm3VtxWF+UvoMoSgSs0eLlYQ1LNTSYm/R3ZY/iPSLZ680F6lZoIH
PHbmgTMFk3tBE+rqVbDQ2vtfEUNXwGWeQqe/YkXahbOD2vvLUid+qm/RwdlaT6EZ08SiLyJIjjhU
gBwrUj0Q4iVEWz0c8QPoCO7CcTCUrpk63JBhqWeBJg8do8aEv2PEksuYwZovg9PtLLKHVLq6IHqA
8aQyQFnubsJidXUiLgaBeNAkOvv/mxUc3dYpY/oXJbAxRaqMnfqQYb4qsz62IuX9PJECx1e0GMpm
GObDPdh6sSB6rlq1ioEhmirG7jIQsjeWcLP5CDdm5cPgQMia5GyLKNmrVam/SeC40W3/V+JQZdfD
LPkLDSYOSZPqGBZe5fhTLyN2TpqNI0851/0aM7JdU9rINgMjlTmdkQ/msiPfN5w7X3e1EWAclRWU
/5WXTfYTLGLoMYXjJshjjJozLPXIJ6UEeGYzX/bkNc3hsKrPQ6lMK2Pg0HHrt58MP/sE7mwpXEEj
c55FCfB80rluThSHPLFsoH56FpBrJUGEWaISIWqBMbpTbdbPJKxvBFnFrvOye0hO5e+lHtT9/7fw
4odZ4hNglOGIE9bJBFgbrc94M5fpWz+JRiaAaj+fJyBQJq0zIhj1m7QrIcnxSOhI3kS5+SRUOQTg
16eqs5+kW2ULN60zfCvMkoIeSDiA0L8fl1DoY40tkTANiTQAkE0wASlUlLevcoKJaCFv9dDApm+j
edoiPZ4wqni/BWTj6B7ZjcnlXGWOZLUqRp1idgCtzopapckIHjxOBbHeKJbV1iQDeOASY8n5zPD3
hvYhqjJI+wSnG9G0ohnFYnYac8v+O/yq5yUuP8Jbr2QB4DUToprAd5JZA/YiUKu+0SfbXhOLjOwt
f8VQDjEEBcWmu9Qz6Rx4oWfYVDNrgVOsYrdthoFgKbqucLp0pQkx3Am14LYfEE2U/pmqyphq7xYK
EUJ6HfvWtzsrvweDRp9FfT+6FLI6jXtWhGw88vJ3yNY7PhJAoJ0lHBjW2UcymVYJWWqCZQMFbTPC
JesaCjiPZXKfEEftTY3j2f4aZwnYx97NGCjK5ocbDfZ8Rp6TTwaH1RY2n4rqm8oLCBkScdIaz78C
ywe/k2uRkO+JyeABb/hGKWPXH6b1yySyMENMFqLinB7QbuA4jMr6n8HiAuzEpTTSnB9WuyaaV3XW
TzOg30FB/mlIdP/L2OnfiHo24r8q9VVuYnP0s+XhEAK2OvLdN+AhGNdGdw66FuT8z9chx8b/mI0n
zNNf5Dyxe7GbX3l6TPlQyV4V5EcWMCZz2y1da5DsmlTzY3wCPResN4MLXw3CF9QEHSJsY0BD+hgx
dWQ+B1weF4K98nkyIwztnBL5qmDoWCYjI9O6C5+63PzG0Xe0d/JwwofcO0d65+y0d4+aYX8YBmBu
7Xjw4W79/awAdvgDO7j8Xb89UXzOpHpgnm9qQqOXmGtLbJXEduBfgOP9qEFBJXQ27f+f7pbs2WBI
Nm0eRXkpJ4EKluSgukjvsl5DxRZct+dJpcVdQFlcKLZI3gz66Jiw6IAUoXXMTOmc1QxGw7tbgVZC
hwBiM12bj/gdqwsbkrT9+N9gTGlwiNywU2ScXr+FSZZfjF1CKM+9x7vuvqtMgf12/++kXPnje4gT
takMTvMXdxTdBJLgFoktjU4e8UQjtN0qBPWoWfoN1xoopO2L7OnWfJqiRBLLLCTOYy8u1QcToKsu
bJxKYxd3GPADh5vo4r03TQGw5VnF54JPsv2IaX7/bKxJ7yZ43IOvAStKFOZNKrgn4TV/nI+zvTyQ
ID65NG4G9NkrZvSLhSq7oueompNh1c/6xghbbBgTt2JvPrAHINIPjxheBN3jWlv7XJFdY9ltfdRa
AHuRC+NLvyxIbGngDXjCCQF8TgYAJ1aHhn+fBnVaDbxY39t1TdVTqm3Q6INyDZ0CZLpAsxpRG6wc
kYbSKD/2RoAUJZKq5cbnmvNp39uOwihO2oDWbjTyvH2JCcOnfeWdZHmGLH/X/VhXKSirFh85yVrX
39sruI7IpdAhSkA1EJdWznEMy1Cekf/Pc3vIRPikgYtID0M1VV6MvZaOaACXApg5tNptVnXs++S5
bwU3WTnBR3kYSw3+HD1ul7K3y53jtIPu5ejcG/r9xbpibG/vkiUBZ3g/Vycvv+NEjzIjACl22utN
/h+LCzRpJmxOxNpzsTAv0PIdfnoUbUO6BkCH/B6ifMo9wL0kltedpAiE5MMrBKtXalkyL2GkSkR7
opfVI9UJ0GhNhX/d146YwEn/C3npznH2W7aDNFDtqwQfWZu+EqOsa0kbjxMKECYMcyy5H7Xsw70G
Tf5UEdedV59i8V1vg55GquBwjMZvYZnhyiXsUwbCeq8lfSWufHy8N75UJKeyHlU/38yOqPlaJtHY
+6XjcqktlQ6zeplJXke+ZM6n8r8WwOuDFoPN2RIJylFe3hmqzXRJDPsHwA6BXNXXX0pFd94dl62z
yR3HEDWMFbhBz+yWSezRuNLPQYBlAUZAZqMYYQFnhQ6XRY2UdfvDm4MT9f7ePPlcQmQ321WDP2oq
g0OlhXTxmpF7IUsDOq+2hWnuSjWbQCgtpIV91/nBJqyAc059bFMZ2KbfsAysVSpXkQqyLnUOGumZ
1MzpQG1RMEqks7x9DIAwlFtK2CmgDYyqFl4Yat78K16HfmocRPm1VPNbIB3JbQEm596pp09LoJfT
0OGPjSHI0q+BKWArCfGDHExa4wmGyE8yL6HmGuwBReiCRq/EkJhZNmoAQNX5qrN3C99TbRnMZp6A
1H65dxEliiobZE96995gIGuxtSWe0HCf3AhNovXEdCny0GVx/AI6mflVQrxvUZ2h/R86nACr1Lpu
NW3eziSzeeLOm8mgihDGRcbKbMfRy7PbIGXC3SBoAcS2OrOyC6ZCi9sVQ3CzFKkt62qQObSqQF+Q
y5P+EWFFUER4xu8Cu/ZTQRTfYX0VkFvx7mHgekmskYj8bjtOs5f/VPPRd3qKv/Bc3DRpJloytCM4
r4KiHWWNqWbwr9cllUxXxxND16SeQ7NcL6gC62l4jUSknnXiGfkxwEWryIqjbB+6IBVyjtoFpN9J
sztTl9zBva7qpyZc/Lwk5Ta+S9AgbRA025nS2EdMdz2H04bvOTbTaysWoPLKhm2EIxiHspDNm17/
uuwUUcBLrP7tHtBrkhtw1dGR5tdhAq5MfUUGRlepazT0124MF+ocGDQR4SFfeyoDeFwOdauJCmIE
g0xXD1C3DBnnzc6IJuTj0fcAyO0sIzdvtxqbY5E2JCqfT8ohYTcAdHzpjo0zoIDphaSCEcRofK03
BWyCoaUDZBzPbRAr7SdvLHZPTzUHNCX4pnupKcUtYYo2ogGs+L3Vw2p699e8PYRCD0trpWlcYHL2
BR6b8qIFfKmS57QVKam+ORXwMnaaMJm2ZaWrlRJ8m6lXqXI4Ey1nTiC8pdk7lTECJy0DsGkqOFzW
0zf4ImX1TXOuCqRAfK50eGb7h/uELrAD/ngofP88KqSSMmgT3wiKH7Rr8n8P6Eup3x/x4SprU6x9
Qi7gqZEZNCyyoQDxrTRP5hPFDK4tLVbQr0Z6wFiC046fq5nrvk/v3TyGRsXW2aL+t3aHKsAfFSK/
UqxcZMnLUe/vKYgjxvUT1nOrrxOOFmXVtMbAYK5McukBx/gzNdibdmAAoPx+38R4k4U1Xh4jbpB7
zE4I7gnecgKg/g9lCAbg93CZ8Kj6BPcX38cWA/WbWWzrx8NsN+SzG44pmzA1HyBJyJG9bLaLIZCx
nYx4/22dIgAk5WqaOG74LB8N+ZvzYe+0r87tjLgVoWI/4AF13fmeibDUmNZGXBKrUKEjXBN2GKAz
UO5R+bVpQekExzCf//AA36l+eq7qRMEXYE+hrkfBpLLicPkrml4k1d7MhIPU/g36cULnFnks4lz9
GfWlG0S661DMLO7qBrPlq4p/GAmtf9t9x5liSTc189JzqLXWkMlqKRHpqg0gBM+fXD76EB7rJMUL
9XaNvMsuaL8PsNlNvIb7qnhlj5Yc6w9RqZ6f8fM3q8/QHgS3pLOMZsM2TIIY19RghIKUd7ew1RPq
Z2AhOgs5jeB10MPFAj9zDyqco+LHIZriutFzJS3Dg7P82yTQ5TZq+jx8NnCqG8SurN9TdBmgbqTX
ZMSSIz84dWmBmYeq2X4yClmAuuyExcQ+MP6MNcYWSg0ib1fGSK0hLvTEeRtzkNbRES4qIsMSa6fS
GPDHDf/loAQbNPvor6sMGwa8UIh02QnbqObnmg1Iqh945pUtTChk3WuOQy2H/1E7dVMMKxofFMyI
4ouWtqpT55qMlQkij278LI7rXsrdhviINZ3c/9vlUk3YdnOdKW8jA4/N8buAcRmCFiccsuvTjm5O
OUpBIW59gqZ4OBcMNKo6HQZul64D5OW2pXitkKksM3y9AXsnNH8Yph33B2D0HDWn43pg8wTvNxNB
8dclOcxJSmy3LnpV9zhpWogiSKg/M6q8UpeKQtipUE3Tjjqwbr8k5l/W8I13u56DaI/ZTANGnMR/
2tmgl5Qppv2bbYJ9WbEA992nFuR9jJtZwwPKywhU9MjABjlE0ZXZWIfvfNSO1qsKy5mD5gdx7GZc
5gQ55l+My0kzcwUZd8RVvDEzEzr+6UXqSsaXSMVUvJV9PBeudftSwUJVysOp5Gz375khCvYVntms
6Jxh95ffLxcREpgfWHNtvE3T/NDjRoYY3jxT99eszKUYoPdjmQ9X4zkH2kvT1v2dXmdycEU6QJxO
A1DMAVz9nZgWx4pDJmFTpK8HrtYHaV9dBPX+efxkjJLDGFbKBmFJmn0NHGLM0773dlwyZ62rG+O1
OC6bLrY6gCNhSjtOenCnbvaD0WG7GnYQYI//FXQzG5Hvxr9rAIP5vf0vH1eQinAUKomiXF1cQJyM
zH+HdC/7f1JZEuUsUMWidujBB6F3KDVhA1z326+mU9pwlwIFn4QO+4HjlnDm/q5Gtw07MsIYqFA6
8pJDMuVXJvXscREZM3B/0RtINqM5dRi9OGlAn1r2m5r95jsa9uq8s50DN4qBhlHDxy1+vkSywuYA
13+xYuJK1fe6j5Cp1fXd9hTIG3GJGqALzDqZXD0fxEMNPypxLBvZBSSsMCaql9VQNBuN9MoOt+rS
bhkcvMA84A47HDTf5MN9VwpH7fB46Bv8Og2yi2Cc9NIMUWCgEP7GjEgbrp9Lbvn9+2WZdfLP+cUi
/6UELYZomIskf5kYl4LBvxx+5zmgX5OZD1RKEPxL4OS7gx4kUPeu6iA4DU+qFKCqJTEJ5g0cnNXg
RUVT9aJtda98xUBuGfV7Z16VRssAf9B76ITOr2hNB4jmR7Q43j7PrwKfwTvHljyOEXfl8yUPbKPh
GcCKs/Hv7ZlN3nfwomtk1JZ4eUmNO1H9z7yKFTJPyrunbhwO+GdubSsV6kmxg90EfAbbb4f0Q6dJ
lEYS526+0DVEzmH/aIuLXQVIgo+aqJf+paVetmAT7Q+/a6co9gYid7ob5+xT0RyNNmNgSw8EoO9a
cBHW0xFuHejPuEX3QeeWWIUfLzS5aupXY54MuOGueoVXtXFcE2DqW0b5OBy4gEgKTXn5eR+/nrfI
q/xiMoYEPRYqQaPIhggYPbdMCXo7KBAMvafHT3SIc85ifKo83xKdmFFYSufDqfFdjUfsN/edgdmK
QIdYk6m8LU2TydmSR04JCvN08qs7KMj4T5m+YgV2Lz71oR2r2eQ6l5C8CRKAvfeg9EFsHX2bfe7O
oEtHe+NXlKmnnYQXecsYUXWB7sRrF9pQWL71+xHbXFpTIAWDCxmjvTz3H1Yu4RiThUKkLkGx9ih5
oRRq4RXgqItG/Expk3i7ChWt+U/GOd6IweHJ7PWtoDRejJikd9ddsKe4ej6MCWbtJ+TGcHqp5flG
8swaKj342+Yh34rXaCe7k40TxQVWuGfjm6m8WVQNNQgAO8Hb8nmVNH5GMd5t8N8vUH87WIHPYn82
q0a2Y6/LPN4haJpqNMW1mSy+5KwtNVnTkczJiDf/nbx0tUkbDQLZpSPP5Vs1AVdN8guYKXTTssku
PVVHwfF0JrxxcazHLFPiqrZmMbFsp3W7KyhAu39CpMZSZUAl2LS8lHMNf5YKeLIaAqR6zbpwuQlI
6664tcLfURssxnNAeWqJBNsTJCEFyNoysQbvb+dOjE6cUcissDqkorPeDjxsf+UG6WKgoIk2h333
DGgdtfi4Ivsy7V5W8VxxyRkGvvzu6heaukufRL1DPnA5WWpxfie/0o1rhIE3G+Yb7KhSTTBu2vUO
zYrEko9IdAIOlknQCEbkhtFUdkLCdaEjkIrFXchV6EIARAeENHxI6payMqNvKUzcXjnDz0lBehyd
muk5dfqenzcv1ABGjBP4hSO8Ao+Sv/mpZRbKhSlyCLpPBZLkpi9VdyvDN/QqSU03omDI8+HDR7Kz
Wmy2i+MeFTZZTMMdgh6lPtKneuuZFy7bCBP6TICS3yqe2zxRAr8GZNlTcflKOy+COH/yeiuAE6wB
KI5eS2FWIWkWHuI+BRlFmwdw3+fvDYCTT5T60h9uMvKGx2eIt0uSAuZElQqi8T8wh4y8+Ed0C7w6
qDeha7KRxa5BeazEDpRpEz39B96r0MFF3f8WHmnx2+tkw4RDFz4bxMeN2/ri9Lo2oFzGlrh1zm7t
gLLiPRXIndsmA6VaVQV8FRdBTcftpr2oiI0llmsF9OTBGA9mKiNp3WbMvXYIJBtLJjEQfrtgp9kw
w7z7/WBOZ/NaWCuUCsrznuudjN51nJlIefyHvTduKBCQVoqy+curqn3ZY/N8SJbr0bKLWGxLHemZ
kwYrGdepcBNmbeudHekL5W5VpkEVcz0uj6trCCEK2kTWhHN1CZa4e6obesiVU1wvLL4nYlKlEhda
yuTZ5LsVY5k/qUGbmVJ4y/SInFuFXMwv4oYM/ZHrmWfSThkMnO57A5SPy36+2I0hxUPcgXTpDBX0
LGkgLnA3T8xAFSSTJKXIZmBlnQWhI5DkaoXcXauSP8rkZ4bDJtt3G+k30o178jSOV2llSJCB1lOV
sTvhsjvNPtFnCowE2IZlQOFjUlNJIP48Vx8y8zM2El+gB7uNSRTRlzopdC1LKaO/aCcQaRzBYJDz
jVMExEH+reCLBOXtyPu4ZusuneAyKV9LiDKwbUMpmd9TSxpCO1GeVo/wo+OlyUUMsEOw/urZIzRe
juz9SgD6ydSPlOQ6Ex+flr1i53+RbqM8JHV1nPyuAXbvgdjzYQK290ltWXWHu8VyMBH/IDPiCd8E
qNVZxTlLXU9BuM2oHUlKBsdKtFitPVSEdxBFbDyUS9VUseYoB19IzAPTrrsGo4fdDo0GZih3rTXv
C9Y3wyEtEzUQTYKixS0dm1x5ZWCSqfL3JYYnPb42RKpv1JHECBNYGSsAP8Fbym9KzWQ+3JOUOXFM
aBwq9wWPFr7d1Kz3wBQC9Wh87X1+Kx30C4o+0CGrHrl3mcLXjZ6ftUBZfTLRYS0YAp3TdTOhSg/C
1QG6v8slqlSSTmtZhseFdfCfNL6sUfu2v1Zn7ZlspWbmjM0eT6tTgiUdowFbDLX5zwnkuYtbHa/f
ZrtMDwCRLXSNQ/RIqxVtoMFSZ4E1kHGWMYNw2Y+AnMnb0N0XBX2AO/O/aAK4+I2AOggtzuyK3lFq
PXDI+pZkVObRwu9IuhXgLyr50sNVsxY4SXQcfgkA1OZFD0NhxpDrHLZk2FtWBIAcKjiAqRQt1mAk
RrYsPp/jTjEdzdrjMzHziq93cE3GnV62XAqdUOtHBd0K9KlB8RNp/IwiVT27eHDS8Hs7n4sdLunB
tFQ9izISp7KbRSqqK7aGNMa8W2AsHIY0oL2LTCmMuI2UE/nw3jkUvwSO/uHIzk5m0np2m2t4nNVH
AiUwp2MUKdQd16IgJIAjaMlzQwwx23jaiKyrAL0P5WUDPTqubb81cAVT/kICKrPIew/SPauZoEMD
vOjnF7h5+iHGRoMVUSbuvNPxgutyiUu8d8fuHYNMEynwMGNy2kuOdds2GRBq/0CChgkbmlcT7oL3
Yw/JQEwJc07eHjgOi1xHQjVaSIHKr94yOo3Ie3Ewf53jc9sDXDRXQbmujkavPwISCXv/BWldkWnk
RQgjEx8G1Sc4Wdkk+zh+jTpL/HQdLd1wC9xAzfuQDrIU4kPvp4/rt57TF5SHXE0mOx3fz/PpgXYF
uWlvzK/NlSvAvYmsFvDnlMxkqafaKb6sJ33UHQDXc0J3g6AdPHRmFJZwVvNu3gBc68Gfz0XfRsKH
sivpk6zbjun79pTUaBlxhH0vqzZrnQjSnkOcy+fLtaF8g+4xOjidquUB54BBqBKZMngwOyHGfhsB
SpA+okmBcTIXoXG6DeGlISleW5zW+1OoqFFTIuOwtFCHJ8wBPEwMjJldVsCcUEOcdlgscI3QFWV3
Vk5BDWEp2+bssQrUZ6Hc94jL58W7AIhaUf6IOt4gWc86f8A+vLwmGh9uX5sV1ze4yBkO+dsuymuk
WENZ6vV190ENXnKg33920wIFFprq3HarsIkqMUzq7pXef6o3WKE5AfR1ATYTm4VOiMcJwZuXZPAv
Uy5l/70skEmpwubTPTPaZ/zy80bDmG42NhHwQ7TnM1l+rRPAB89pkEMNADNjwJBc11pU6bP1dUi+
zUT+XmnGhn0XAWKcmwUwTIOBb2ohCMyZ2cwWlqetc8OIeRBgFslcGHuQqCWgKwPMhuWKWGTO+qNG
xAxi9NbA4QA5V/wI6LTnjptnqlLFW6vWOqFs0cV243Ma5LNNrLfc0/tE5+bgn/+H1RrBmQ8kdrWq
+hwI0FKbVilXy5KLzKjXymIXgif2WqErarOORdSzMo/N1eSrPTkKtUhLR4sODe/cUUxDgHY2sKBP
3Yofj9++yJ59d7VnQx7f9yDDZx9I9CLS7lYD0pkThytq29JMccKfZVFN4IV7vlYKT/RcOkVM2dXp
JrYwNEt90ddxNxn/7wy0FMBnqzlrPE8kOr55DjpaIr8wAAVZYtZ02+XOgWPlhca0A01cRZEhqCQY
aOllExVH07p8rkSsnwU2KOsIjI4NsTu9dgZCu/1qELyt9sivRcBYpQ9Ei8bEIbbmwNDuCPc64JNi
Kv8XDmsBzI9KCGDzTwqrohO73lfdxE/l6dMQg5xinUk0QLsXSqxol7TKGV9roMbaC+ZShrlErDtk
dmXvFy5Mrwpcucivev7CisdMx4DEPybAjgnzfVkcPVOHHzxZE+u4UiP9+iVevuYMTYqPQymMnvhF
TOWvSF/hUOEj/4a+/lrlvDKrJwNTqtFm9dmMMK142jQv8S2PQUCEzwG4imN6wBG5hf8E88NOJ8cl
vXiOkq3zLPG3316PjifsJ/ymSEcDu0cHG/4fXDYf1xnn2B28Q17juZQ4QO7qNuHjmzKcFabO0WVT
U0/Me5UeOPBeR59CX+rdX+AtcVkN3syOsIP4sftbPi+fAh0Eus8egyzaLHb9DBepW5YyWFvjCo7y
ce24oPQecum56I/t3Y7Sn5czFwNGg/PR73/hpQwVbOSZl6JnafFJckHdWDxQb49QF96lfNCyWwbp
Knp1KlIajmtZgFCkvuZ1e5XA9XXozFqlVOSkygnK/8a3bsXb5mxpWGhUeqz81nn2wEwWjcCjhi5W
AVm74uc7el2eE18TlX4gTRbqyX7cIsrByLYElrKQH7fHHnKGFNWssJFiH9GEFmQ3Fg8zv5gK7eQO
EfDAjW9battHOO9JKiEUbx/nLxSs5PR2OxoYK9Hhl2ly/ie56D4rv62lF6Cn9ET2apvngWVVaboN
tWNtGcrFij8vndT47ukNvO14KG0e+i2skFzoEv82Q+GXud4Y7Sux64Qm9oXuIDeYnQ3mcbjuYMLx
aLrn7hxblv9Gs6AcQ2SxNcGRS8lOc4P9DzeobB26fZ0zd7YWUbWs98U4NASt+l/Zq4SrAbZImZa7
jEggmK2TDR3nwoUskjHGcOfPY6HB1Eon4EscomnwJFvV4mda71pRJofKZTCwemPbsGbM50kku5nK
wWEu+MXnZUZO3Lpu/upIbmI20PlaOadpjXJW5PpOAwtn2B+LhmbVs1fBycYUdF/9ILt5KQ1stQ7S
gyGohNJrAHDkEO7p2n5CUwtPpjvb44Q9Fdy8GFIw3CmuCuhGH9sj/JkFvNR5x9f+dS3iyWSFOJMw
XdrIz8oN1WN2Jl34pa19pOR1RcnSagW9ZSv9++mlF9IXKcO55cHNIFNKk3NokpXgIXYNMlRulO67
zCHjiqkr8nSFz6qzysE/EQ4teLD79a/Zn14ROyD6EkxDhMPT9SggAe7SHGsqqRqhsWZh5CKR26RJ
669rkOYPa6HaHIexmRhNBOcZDR3SH/glXRJ4Npp/+Kuj2xYYK8brEV0/aJG1+SI/+LSLvA9lpNnW
27l6OdtEr5aKr8d+7HzY2yoANB6+mZjEAGSZ8NIeF3Jc5eO59pXoxxmoUXjMY3g6cjxy0acQ/usy
p3XdwNqvLPPtqBWim9hBlOhmGHsTT8V63MBu7dOCXrASQD/lCqmuUH0uELRpPaoyS7ikHYBucYj8
rICijvActx0tDdxwNonQF1MGIM4ffmt6QxvtMriXco9QscdSYk2Vkd8zeUv58Gepkt5bziguhRMd
gDI+S92BiQ86xfn0Akbd5xPqMxvTFU5zollpbE1O3diB1gSZMBLD2WEbkI1K/ZXwL5gl35Z7DTIT
XtHHrKzZ7G3J6nm+l62xv+lDaEnOt5gnXP+aNc/71kH0Ksbrd90vTk+SB/dcil0++6OSLhw174Ri
vw7+KMfwYebX1M1Vm6QNOKL8r9q8Sm+zp0f+yu7jQsT3VFHfueufCBsvC0PHa/OVfh/ZGXrciN0g
FBHSzKrwcyMj6xEZrwF3Go1ZBQYhBhPJSFEX0yDpa8BZfoQnUkIwxi924jgR3fwrRkuiIc7JAPRs
p9yUr5dD5l21gucZgEL/gXWgEyqH8RuFgv7xeNrdbQl1UxMu97HvIlaJgGTPYYlpo2DeFQmXs76t
JXLlsZR2VjcvZXWuJSRqqWQF5HeTllpKSUG7ss1pSji0/xqiLVut9o3ilCyjunj6YS452rEvOcbp
J8F7xlPWCQr20YGDMJGgVc9vfGJQUKqRin3jEESFXlqg7N4Rb/kk4wM+xDvyCOEretfsQtpJZP3C
povuTtUVhmGrfaLypA2crZ3+Y933H4VZFwOutM4dN5niesRcxlrSvX1CfEP6IAN8jwyu7HaY+YSr
ObmIPnea9PJHZmqwRC+YGjK1EbwvEqRPPP91o7Tj5Y3T0KIXPxvstw1sViskHhxZ289fWRW/Tgkb
4Q9A0L+Qi8+e8FDQeEA8qqOu3/msWILsGIA8zDoo/pKZMNQjlO1X+64ZnSXNabiVjYndQAy3syFL
+P9+xnyHc/QOHGPsDPohl55yCeg1OcgVKgM51xPArFNFpbF8EP2xA6uZYDgeCcfhbAoJvG/FXdxq
/hf8ZlLdaYeLSZwEuZzmdxCukBY0jBjaLcbqfXz568yhEZM7L0eTOvl+Xuks2V5ZzNMLrGGOgw2q
adojCTXfz4xxNScUzn/kBbediJr8f5nw0faYMOsdS7qWNLLOyaMbO/Q12w4Oj1s+6aDHyLmQ1Goa
jcA3NzDQE5WiJ003zA4kj1aAYUy6rInhIygf3EOSbymubWD2jrn5sR9Xo7Ds2WFzhU1bRdNxyDuS
GwJSr/AFnGOJjiBoAQjh9j5UMXAaFIAyOoLy8xTawpKTYTEAAFsaEyNJLXU/rlt1v2vthIKdtBHM
63hgKP9oPjNXBWGVF2XbqvSsvaZOnXNgNwPfzqPwPW1Y7KhGSbOzBPwrjFtyU0II3WUciXJ7WG4n
AawFBU5thUv1d8r6bXHmriJb7T/Ocs8JOupfD0nSlI+8vkbvrYe76EF3rKS5/cEBnFVy36XQTGx6
oS882x3Xw5z9ld0OYw9NzWTeUwUsSXH6vzoJ6KiljNdETh+wI6hnGB54f2VsRm08jX6ufILgL6WT
RxgrnkdP2xsZwv7Zea90C0LqgNh+g8uY0FSu+gfIWmUCxhl2aVswpbNLTMFYJ3B5XU9ALMyGD+nh
DO2hLAAhxK52hXxSVbV3aJgdJwFNYapSlwCw88DlhKrhfV4POvlii4rn6l2uE+fpUQ6vRUkVadY/
iKhXpRIESEM8VY5pWLk+bsNDwE1yF+9bOUA9bh9ZjUGmbljXI5PasbSRDMdtEWoA78Icq9DbZgOQ
lYAPCNI5efs7wXnwCRElXeLwzJszSkUnwdM40FG2/B5CepprXvnGW2uFpvQ3poTZ9kyu7eeij9zq
GUFZTOpJ4A1wCgphHgqD3nw0/kzdZBT+XOQBd7X1+NPHy13awcjOsiAwb/3OiampIguIkd5Joiva
Oq7YnUm8Mf0gXzeut8Vwn+yFHAiCRgJTvvAMt5PHetElc9Fk3ukWMBRWQgy6w/EmB4KpfmsR/iG2
YP8heUHaMzp44lYPXRVS5KE52NeyjhRFLeteCF6yfDKuj4sugQBXtYfljN4zlAZt9OzxFoNyEqd6
YQfdoGqZqjwu8gh5FZM9BZhyzjHwXR07XiKkw/1nnIXZXkvXWf5xb0LxtPv9F++wB2EjkMsC0cDg
budB4eWSmzSxBfz7+sxZ0RFp8MDHpDysAMAidQXzV8uJ5qcYCFXNQd9EPj2bhSg9s2Pw27fNGFsu
/zgA2A78kN7+PrZK3GKHaAMuA8VlTRjDkoI7yXw7cC5V+FT4mA9OLgfxzQCMvh8xxC5AFCJG+cUZ
t10sYQsvyLqFIFMvKz9h83yIPie0ztdrBaEArxKeV6VqaozITlaOdyOV7vLak2r7WNvY+8zyO9Zq
vdLwR2KJ4DR32WZh3wr2vTPy/cszPtiOpi6AwAYyMIEwCPiQPa+O4IZ8P/LBJZzc9CfxnZGBSB0r
6YXCs44vbL47XD6+HBuAWHXBfOKlCzYG7/23AMYCbZcWx3wUxltPPJw1jtAnQv+C6wXy3VZjbnq4
gj57O8C2Q+4lHItQ+lqYZNjINniW7FSslRrIl7yAHoZFH1oxaAdpjRP5MOB77iEqlQLf+nukrsO8
1rKB3+e18LSEkeu8yysq0Ll0JZ1WLtz6GBIC+wsWExFePPP6DVohNIZzqBpgPPXT3CC3n/r5l8We
PmeGf7Es8pim/ip8koitZxksagK2aiZOxwOTG5ofQi9dpkelgjzlYc/letq5FsyGQHiwI67vvXcS
/bcVmE+5xfcoM5CwLxT3r+a1rIsTxjMU2d8sMl2o5/A60ZSqodAHdUSWs3pY/ccjD4MGdsTWQaDx
2bWnwYgVYzZjhSHV/NbcrydxOx4BCKzyo9vkL4gCYVhBfnaE0iOTSmtg8ySQsn9wGjFlDSuslzYm
3DIImYAGmrfawcOrHKQ8B484Je1OY/S5PbPdH2mvmU7h7zc6+b8PqkdsF7xAdd1vDxn9JdGoV+iW
E8i1DPzxifDngcpj+hS+IMeXRcbfqaleeQIBVYEGEBpGNHGcVaozE7CpGlvzaHDV6p4qvQP/8/Xe
tEB1QHwjIngBVRtwlNG3O/8AUXSQLO0Zd/h4tgSQyKORxYh1gF/PSZpjsp2AWeovToLOin3KpMzF
pgjhTeNaaZ1jx3ltTSarq8UYwETGeWtBAk4zxH1/PTV1HrqgHPflMsZa5dc6toUuAk/4yxWHooZg
IGcUfFP1YOU5JJpCT7Li62XP2b7KIi6f58c0736zO+2czSwRrSvnlcgfIoRXixoY+ZchsjNWn/bV
bB+Iqm0iABEw/Ia55/13kndUlWpcWaEt92wnF5jEZtEqdvGFhO3UXro2aaPS0KTC7O0dgpYCro5b
gl7QCsX3/dJlJbKTQJ3xPhWAb9hXHgt+N2dNpEgdJXfyd/qL7wxGLeYHfuX0xN3XDqf+CCMxJ5wz
EyLDDZi+QLaoVtgm+MI0dY5SrlAPnyieWrqmkhmk2ORcDEZ3J2lz8WAtPfWfErPGfncjPUIL9JGB
kpvuKrV3FSZIySShT4JKbrea8lcGf/IRcI6J842zS0A4S8CT4CxwPBLBRZMI6Gj9HbqIzo351yEH
x9Kpb335I07lhKR07MdqO7Y14LJne9oOkKcpZTAwIextG/pNlRoK8rZjdNEne7trbw++8t3BQad6
xAlFCXgjBFDVTITblCVMUWabbb9d/eW/q/bSho/7zHVE8rkkraWjdFvgCwGeTSHsj3DGYtG2Ur+c
NpH2ydu48k6JXsGlSvJAq1WWHgKHfYsjWmZ7qPPxsfgB9PwFViBLK5cehi+tdbF+nzWquSxlV6Jg
iRH98/sshOPuR1V4by8XeISBH03+Xn97bWVoPOmmsujkZ/+bYuXUUanIiyJFGdhKYokKC3LYKiAO
3D0QHbhiAq1giS4Dl4D6sZs0ldKG52UUgvyHgf+cSCLx6NRzTftEU9OFz2tCm85tx5dAyyyF3898
dOdLY7amU9LFqrlH2+aIA4757TkrWMAReQAhQOda+R4qLDv9nuc50KSsKx0FLbxGENhmYiPzgm80
ABbTYL1pX+8ShaNnmJgVittSg6vAnRkDhUXE5UCsbpwcuysXmYwmJf230nMRs2/3xTuCxKrH55Go
MZhRT3hSzUEGHRe0Gkl5OXKC3K/WXePNVCZnRJVXlJRUxLZrKmKYCazkJ1jQhhmTS2bAlIHIq9d/
wGm6fFIhj+qVq6xsq67FNzGCcz/1sTR72Zk/wITH7Qm+J5bGZbBZd414k5O8YvdQ8hUS0S12G9+T
OZ4FoDsUlqUeWUlG18XvgRNK0M3cBCfz7GWOtLzraiRAmgNacNwM+kWB0v12qOzyBjMptXFFFhmV
+1qiQhUj4HD9f9l9duWgAsZKgqEEtQtvJWHPREP6tM8rkJWSPioJdsUXARMqzUQ7T4JNe0jYuu0D
5E2pI0I6xhlcDNXi6njbpkMOaU0LjLRd+eVQ62pWyCbJn7Km0H7c7rGaMMqwuL8L/V8F8lkGwpoy
2InRBoGNE6QpraYZm/Lb/1KSeD5B/6u76cpb/OvRu1j/a9OoG5yJy56Uq/Xn+H634q4ewObxMUVw
tw59pRHKk8FdEC4yxbzMRiW67iGtsTHaPoFf+qjY9Lw9kYKKl2II55jGJSR4aUyLKsESvj124Tyi
7JJ+iV2ZToOZy81HK9NAPiP0kmw7v1RapAL5EXFfV+qYvcZ3eS2ohLgpWbmnR/jDSwOZJwETNaxX
P2VRc18mqrPsGnKc2g1LL6idgPKNj8/u4pdQT4QnVIpNnHNMSqxMVKwoloHBI328Kcyia8p9T6B6
N8KmrvfDBHDkB3l6UFV6pN97+KThcjCB/rakak8/3LAtrNiKcc0pNeONTQc6XFEiKrfTlsuaMRIQ
GOUfMLdKB7GwHxCvoM8IEC7FGbCSXDOySd62iBcjd3h3cwYm1SmiJZWLQJjBcXD4Q0FzfmI+uq3+
yhGAiVCoEDL7G3zrPKTt3plRU9hZ3LQk/I3hu5Eab8I0WJ99fNjzcADzrRsJnb3Sn7T0MiEM10uq
9MvmMygQID7n0h6WMW+gmmq9xLy1xYaUmoovHn3EGacMdONU+8lvkDhEcxfNm/jmnNsjFo1nRadA
I+ZuL1mAhJsxpaFncMPKsV8ak/4ZbpIl9I4G8MGOcPcdtBl2q8FY3pHud7gLZjFG7N74WnEd8K0E
NmdyHvb8Ct4xr7oI3SdA2uwdw6knxwBZQbVEI+LqZuRq1sp8yf8dO8la8Nk/IRzRFHl3AI7iMkrY
qzKnz0xEg3O6/vIVatWFJGUZqwDmCQ2PaOzmmB6HEWCVxWWD1vxlk1pgdLKqCsXztHwZdx6xlGVF
nWizfVlEMr/uUnOqPd9MdRqDYWjHocuMXvkseyaGna/wC+bXatOZIfJtfyhlzVE+PkLb2Q90bfpK
h15KWOZL1prPW04eNWqafy7rbU+KuRY4BXRoPR5Ny+3Tb57PSKt1wgUavuc6DbblqcDtsfS6uHg2
NUoM79eilSwGEKjHq+AjyJEthD8VHOs+jRH5k9gZi5nijR630aC1FdcWK5uUTkcqdhLBwLbhTmjS
1zoiCZyMhaF3Q+r2NbP0unvXE9on2KoYvwz/tGfy2HGJMAXn6CCoAwXXJHDUMcUpCuTyO9oxvz2e
T3/4hD+Mp/g53PEb/RvEFZAvHcycBpqwXW3bxxYeawx6dUzzZSFyIysJTTHFf6XrIER4zRtikpe7
mTNADaEZfJ0KQY6C7LT2v26IxaeNPDW6KynBftBOG3oGEjVmE8+srGYt2cT68tGBoRBYmi493IPH
yRxSDOW8Lcas1a7ufl/e+6XUJGMwTA9zZEHRdclCFWFIFP5cIx9Au1wC5Ua5yiFPDBoG0x9lTOuo
r7SHcjOK/a4kb5Ge1jWx5eZoRvx3PRcA6mGUaFgX1AoTQYyiqlIrGGgs8yl3xFgwNacvge/7wVTq
Vzu3qC4TBsJg4nrtt8G2ilM3gYXUCjhod5ek3aGwMkMNkmR8xkiPDADdPneWSNNTiau3KHhs8MNZ
YUwpY8g+OwDhyoGc7eaf63LKJ+l3saI3mhFomS2lCIcbacSyRGCrHkkX2rFSqhOpmHb8EDOqVfgU
21uHk1TAh7I246ZEOk9Ck4n1+qwjhbJnb4Xt/h2wrFTytMJXpBW2AIbxyy6DFamY/SSpI7x96CKW
uUeGvy2IHSCX1GcdyRYWfDbV42067AaNIdpEmgARIyRwIrYSaYSuihY3geMYlrbE5Nr0wAtfmF27
7jjk2gAvod8XppkdXP0i+NLrtxKx1WGxdratH4Edd9tdefdV6vLlSTCpWgF4+jmGAyjBF8dnOfZH
II/j8+SsfgnxyKrhYOOmVj/74VSlfEgJ+15VYVkASV5Ewi3ML2imN36CuDIsPesaCnbM+2kFRJbp
UUHa6IoC7NOv7cDzYvMv0WqcxlbtvDQTOK7nnkjMKb6ZYliG0Deuce0c5P/lTMTA14bla7u3CfW/
/k3Pz67ERJOWb3Grf9T1g6t1csHOIqqXWRAzI55gxNk6hldZFE7I09nC9eGXqIuUfzOrlcXTX0Op
0jh4oIe9vs4nObi5XtKr3fGZmjb4WlDs/i4zKdaxYr3jkTPcKqM8YaBilgJFd5guaYyhqm7CFNYt
5ciSA1/Xc/2VQbNCFssMvas7w8CRtnXoGH3kKkSHgMts1p8GvnkXAnCLm3QB1ig5qX+bfFaYPUy0
UPjqJonWxKqrx8ptC7++mYrhIW08G/OZN9fVe8D3r4qWVnLbNPoMMDrJOtRHbdYne+8nNXg88HDx
RhRzFfXPixK6Yz0hhbc9hQb1OIXU6l8z50pVAIjavmmaHArKEo2izDUINHlCk3i+OjfvpmnpeyEa
dXFk39Qu3BhXB9LkGFGF27hrfJzj5ztwu2PxOPB+IxxFTnU2VJfZ2SO24ZcDT+1oS6LOuivaMCsN
g/fdLwr9zkXCKYufHLCRLjK7GX17/ImiXdNWE6+3hgHvx/0ucPpmp7uQ0MgvFEfWuCcEtih9vFfd
D/59TVQDYk9tTAdzHFssmqTxEd3Gim50mIqV0TXpU2qX+Iw5SFRaNMdRugSIoabf8Iz7mTd6eMSs
COfM6ya5I6Dvgcwp7s4gWLOXVkkIU9LxYOb/m7YwpWYZjSGMgnqw67VQ+GWq6Cbjvern2siFAijH
wQxyP+vV+b57EB6v6oJPZTtPRJPbTzQBKWK9LzNlzioK2iFGgQhoYgb7Ex/bjRt56R66/WfYZIQh
IU5hMmKzQuGF9wCR/33Qj/xpv6wVbS5BQEMaYVH/evTHf5dg/ynV9hyycQle8PIAwTX59wguhLtj
Oxc34Zsn0zwWXN4Kn23xCk4L5pXwYdAiNFEEq8gZND8cGCcow+iwwWXyGJvmNzjAh9cCdjtfBJ4/
USWiY2Ac+dg8Lw6PV/djT+JZfwQZesJxq8hC/AjbzTRGMTXEWaADRhCNrfyg3tx/wteXpfm8P2+c
x33+cRTwITcyY82V+1zKmldbq80ZE7xuqeEIkRyKRvyMj7H1h+Sybd1NUrsN9jTZhhK3WDn4l/mj
RtqvYqfC9VPck4qYU/vhgKkCGT0pZjTvnKQZK4Ne/gCfyOGvrrPFnB5y9GAazPL2ghUzZyWZBsdY
Yiv2Dq/Suxd7LTOCCkDIIg67wXpXlGNuQHTD9Rvi+zJUMuOD29XE3F+ZvTt4M2lPGebm6X9mIOeW
pvINh3U0cAOj97elLoEmYn+7q3MV6sb9KrN61FBS896nkCYiXnzFeaOYE8oJXzTDKnFiupGpozc5
W34kbYv8hQJv1dWOKg/6+1cJ5jcLLd93xiLkeGUyFHeME4bQypEvC81NDPCYQTovcpCfynaRGZAc
sFuDnlGx9Ov+uTRWnDjtm1W9DBhQWQcaMHSPj4qX7SOFpmZfzlsLSrnD+4wnD3IFOPnWSMKzaap+
MuU2VpFPeGYFrP7tT5Hjc0HNJ32AuG1g11rx93LGz2pP4wt00j6iUGdFdhpcNv+dVCwkD/gnd0Ad
b1lc0ZK6mxuDgalL7PXpZakbGfWw11m3Ly3FNlZUNPlGwbEe4no7usqymcG7CsnLqao7Eqh3zwfd
lS+fuR8Yz3dSrGlKLBgQu54DPtJiLK94UxBbef0P0FT9Zx6KEXnmawu8SxdRhSRCnCx63dx8BKaE
Oxo4sMmBdL4cxO/bWZa6v6mjpWuPWBEw3IBaGK9f8gk2IrZM8+D6xLuJxk1WmezljGe4ZCy8QNW7
xMpo/rFqFdOiJyx609u7NJzT3EJ9ZYPyeqRqK0h7Zc/g26kTxakfQv88jCG2vzTDQxTek/dbOypG
DI0jOQMKwlcfSnZArxyD1FFhejlco1BS58hS0p/e9BrILstlVMwPhoVqzhBcUkpXgUVpuzbrngR0
ecq4zWiDMZvVpevI9exndSXo9NmmdtwNEtB23Sv8UxfJv6i7wZQPELUEws2uLzdX7ZFrRwdWVne8
fsHdTaSDaA9Lh4V2GSMpYaHJdCiAEvCLFmhiFE4qQain85cE8O29uHQWeze1fDPbj2nfLm2ZDYly
ZXBzbYNflXIILNCp8Arzk6Y47RceO0LDfNEn45nMuf9GXxNY8vCCbgH/h6mijfzByQlV/JDAhu6u
nwy7TnA9MfWd4hLrcVH8dnjP+vovJx74SEs/8fs7SddqwMttdOndwTK0eKnZ4LLkc+37/JqetP2y
KBv7KSnwsBvhexfsP0OboxeepdQwHF7gLIVL3OmUDltPK212F4d5ups2NVN8d6wX9bTK0aCDwWpH
xf4IypFOBab37/XeHjNVsGwU+Q0peoAlEwqWmC+oNrylPd+UJJv8ZFEw4FRaMwuTYDHTfyGaQH+C
4NI+GQgYjAlO2nVN+dq07jBImJe4fT4rDlsMQkiAyZ4liVrxx+bx7xpO42HPAidrXd8ojdJlS/MC
3NyuQCgC/wyhhgXSCfztSVX3v1+AnGSvr5qfzsW+VJK2nGGBOPwmaI0l8jBL/oO8X9UNIPYevWDD
VMvYte8fr0j40sKkL9jaiWrf4MY1vFH825oPc4FlUhxVp99Evg7VHGsm4o1129M/8m8wK1RrDJLZ
nBVDE4QHHvcv+FA5PqRM8ZQUa8Gh2xfVB3Xp2RKG+2m3I8tjrg+Q0Zj681U8JtMuSw/YSnMCmiiS
+4xW/LZgxA+7lNb5Zacu6NFGyMZetXXfP3EDoRl1EZ7VMGX+lRPcYs9grBYDgEVI/Zu5Jp49GxUz
unCvoWSZQ+Wg5rYt1p3aeLsnhQTiCXQ+pAGSkX/jSa3OiSyg0BpoPXQevG11bksdP4Ks+pVe2xzN
p4aVrZimg93Ny5vYnGQ1yjR5BBnuoS7uJoMzbd0d8grbOOUQ5TxxVmWxAJfhMufzZyboLA4ZvbPG
a1/fDjwAfoQoON+9GObjlMJJ/M/Z+CoaLR+hIO7In4kLCIaQ6qKRP2zLFRkrRTHXpcz8Tkv2x6S7
any3KLlAxl1p6lxRv4hvM4UDjnX3XQwZaRz03a5VE4WmToFruU0PQDYazxdEdfYfp9w0THytLfvy
X+Zyqqr73UV/+1keCamBy1c1LF4fsij6gNbzvLRstNSNw2+2wW/bfrLNmh6oDpFJN6LSYpg62u1z
o4lGn7aHyAOd24poba2vT8hYQ3dScDcLfkBTLBnwHbe+tEFT80wsRDfWrurglTCe7+JhNt9/J+46
YEmAir6ywRMRYU5OMlukDRMeSIgchW6iI3gByo+L1WN0cjiJ+V9Gi/YJgDRVaJ8r1ecp49/sT7Uf
DnXuJBwLmJzxoh+1tMW14OyLXglKk9qe8y74TdQCX/LTletkSALGiFTuf0JaYX0oLJ+bm7POcjqh
gc9gI6fYanKtVxLUqPcnsNgG6k9JhMny2+Tf2GmJ237wOucnjJ/59PB+3xeIC+ftpytJ6Ygsj36g
KbjhF6VtqGZfnNWeD4pJ/Wh4qVMs8VSeMFcMEYCVOQTXftfyrdQwHPvonlBROySI7cfPHdoLWeMw
Fk7vB6UkJfcvsP7Y+So3XniQ9Bsgeu6FSazt/g9r3CMARZehUsehqbXu0GEDQH7dqWgBsxd3CMIx
CYaJc+snFAJtH2QUaycjj/Y8uoLENXp89khkE/BTisf+wJSIIiP1+afxcSxPrn0EyQq3J9DVo4DJ
fEXv8msHFvYXYpRVPY3pyO71de22CNPTzGZlljwypyiUkF7sqLraLl1zTZ4eElXqjxHbD4B5eoon
DGL/uzb6jEHDPlHPKNkwWpGUytDXuBozH/V5VNagxUBRZKV/evSlWqAemFPP8A9SM+FdBlL8tZZa
VkXVTZS48w3AF8bex93zgVC6opLEP3SuqWK5yRZt6iPoAay1g3EkAQrUEqnjKseKLg22fl6b4Pxf
dvT6jpODlYXu6HxZ00y/3XTTMTM0qVSMFCsYcqR30qrdot1k/cBfL7Uh06oDXitZPf5BX4P+p8px
YArkHF8PsrFWXn1MpgA10mDS0gi3DzAj0fD44TJl5x/XXkk/phKgeSRWAfxRcq1oCm8mWju/G/7y
zxu/sF/B49JTIe2c4qwXAcOHFs3sTIYB6+kF1mkq5vATvOGn1/fuLsuwztF4NjpW2aZxt8upkO0i
7GJfb6nqDJrWwYIEQwjNP+sgtBx7Fr9uWxKO/H3vozWN/eHV6SjIfzxrNlZGFAbjP0RkMdUKgWCV
JVo1wRTJEqgkaPeyqXBQC65XNbFq8swibXQkzFy1fZjOo+mv5N3mYe37eD56tTEgcpEFwplTyzKH
SFUInIItLWaiYiejfTfqR9VqJAUNu+bIhtokkpXW7/a66ARsnVApGODQJ1aHJt2eG1J9AI08HqE3
MWS1AKjJrcI/HAD12IY7He9vRxp1e/nMUbrfnpUgpdbQhag+BrGON5DhRFoT6KCEuPrRpPnQK8JA
/4UZ01cMBD7mxxnh+MTsYL2anlIyIBQtK5/FRYqU7mki9polzfHTvdMlm+msMHoUIwiqvNZgSpoH
6ObxM37S+qbW2U0N5Xj46Tx6rgEA3Mbt67wl17np+xBfZWVMgqH5o9DPvo2jZmorGl0YPTA6lXDn
V/2K5/F9qGIcesFK10feCHFxM6R9rn/eCFZUf4oJOBfADZ+LjBqwnWcE54PYdmJdhiT2keiGMX5P
r+eQcMG+Pm5xdjgRmTSrJ5sxJ/Hws1pv/4KaeJYT9++UAWaMsqRCq7srdznJ0wm0FPuklRUGs7uC
ybTnjkrAWeSGZolnOxpfXE/8Dhh5KT8Idy13CwG6wBUzr3BDrDiUlym3OMzBA0IqmpQe0WQFUs7T
cnwgUZj/+Fq44ft7VfeJV2GaIS44mbsebOk5XhRj9LGD9AEQeh8Otmxpsnb+DE6ilxAdI28IXL7s
KM8Ic9fDvl8j1JnDwtTEhieex/fIysXgvdwUYU2EFt/N3nXkfvZP04v1H43VMELxDxa1Tx/vwT5B
4lyjybm/9YmaKgj2hSuan79i6eOl5HptGLqDiOdNmPWyWIeyzgJcQKzwcQmnYaUEf9ibk7sve112
f4fRe/tzJgDrgNa2nrlFXn3jgXKBSuOEsAVzWAirZ8vpZYwHSoRY+jkpw/1CnU7+zfsXvj7I+mW4
9hm0cy2ZBwYqOkmrZ0eigfQXAx8h0OT1ku16UEQRE5+v5Fu5zCDFixJ6Flgl1xCHjHdZfWzerST1
gF7pdWzwNkS89LlsXWwH9XZ91M0r3AGyQEWCJhA4ud9ZkMR6c34z+lxkqcuHMI7OVJQmxEWvj+T0
3SCB1qVsHKCqSMWwMB+0cDSDLuuK1huZb7mz6XWaqGSmbDol6cmHV7JHs+d0UKKm7MkV9VCOGozL
+Z+QPqUcHmW5p+unzSTZceCKhKv6PvoPHB84N8G2jyBfNagsR+4ZPywihRQ8ooL89QPVw1mq3Pe0
0VRsEuXBfxB6kn8/1vvNbnTG3p8/FWG2ZyrS52lsxLQbR8vbPug6GSRPgQbE0R6yqgbyglzDLNvr
o+m+z2tT6+i1zv4ecHtwkDC3GPUHcLAvOHl7F+H4Z3BRnZjb3y0YA0p52qasLirgmkqAs/7NwTrc
AASplAW3IqA3OlwyO9WgYFzuKk9E9xbEmm3Qcaa06OQw3hM6PEAtcRmwFYzAceqCvLut6DyJA44t
mQdSKwefF0gUUgoPDmpoE2E0V8S0F7Mg90NQJ8+umj/ob0q2liKTE5ZEQKO6IG0ZIZprULSpka19
lHkpZH1H+YrwgxCJDg9bI8Ao+yWh393p8aMMNQtEDAO9MthaYS6L+ShQzr3cg5M6gbZTn0QjsOPV
wa23mOOeaTrJWV45k2DtjUrlmxUeZ7FnHjBUMpB0KxWaJzOJuv1bcc2TXxegsNAcQXl9ixZ6vC9e
9FuBTVaUwrHfo2DLZM6Qsafv5TongZ0pavOXBu9tr3FqBCSEHLRxgT+a+jcqZqSUnTg9f+mC11T0
WG5LdBND8B41XgIk2CKiQHbDiIHHfDaEsV/FduBfQh1jz+UAvsIEkhpYSaWWR0OrypsPsBRJuGyR
fx36DH333jVGjsYAJwp3OFDOg8ji9C4T1yqMQNm/HPrr086enG5N8n005aIwRnH2DQoIv6WAPzlQ
2m/BtnNXHSwS17Sm6daqEx93tRltU1ygZkfl8rNjKlM/J8zbCVwcqFYQe6kfKI2rxBtKUrFB8Bw7
68+qZ8AmTDDCT1t4lZ3oI+bj0KTQ3C8YY3h+M9K7Xm7cPS8lhnshs+Hq0kkWnYBaNCezysMelkqK
iKKAP/DvXzaNcKOsmYWpBTU0bjgkuNRMxRegzjvlLrfHgbK4pRlmlb/NPLLfWjJJ1PeuIarXQM3S
Brfdm12rdS2jkFKVs3DHo7Og+gXOMoOrjUYiivwHTznZM1nQj3ilhsYlZOlJckKcQu8ncs59LMeb
HgeLQEa58Jc/BiiJkOthw4f9LRIlIxx1kXRx/dX61D+Ihhz97vNYpYGmfLo2fr5gLR1DdOg797XC
nL8a6PoLEv66HMA0Ls0+AQ4WNrNTqEXDDOAGph/sLlWoLJih4k2f0814yohtoapqkWdagUU9LVlQ
Oz0er21W5gX17a9AmDkmALDNTEJopuqUgvguuBeEyAlRfzpOY4f/UFX7xzN8d5KZVUNuc6waHw0O
UmpxyMCgklQ2pV/aU8G9jVVD9sawMmNa6fyY7jb0ZQfSrcKXKbxBfAwUwNLYbyJNanW9CGHdgX3y
M/cLOFe/mLrsIcRtK74wInbGETpT8Ezb7/Dam6q+3PnUDqX1es+rTY4iOcd4YyIMsJTXqlZSpGZ6
aQ74c7uqlgI/OoKb67pcczE0IMkXNUvVhQ3VJAI1Fc6yc9qk47pE0livxVkCPvh1cX963gPXjV1b
cdDqdPgh4t5+iKisdJzUywqbH2dTJClNG1bdCq8ylCnl/AaHpmwgfJjY0+LGyJo8U4appwaG2xa2
p6ZooQQCs6l8YRCmG73muh5+OtDspM0MBD1/QCbXBePHRys7E3OPLsyPgQxHy304wmRCxLr9FtpY
7OzXfU2OSXnPjuja7QkoI0BNO+RQNvob2dv4k4vGwCvfCI+R2RX6xICjoJxOHIIK4VnaDq/IoDk0
Rf/3/mwZ1SuvzdFGgnZxUPrv8jPm5vYvVyKPER3azqvZbLKVDfna+fYOQhARSYFyMIP0p3GpF6Rv
tAhEULuuaD4c5ggWk8vHkHXrzdiLuofI1jOfjFJtQqTzn1zqLEaKkfi6Oe8tyXc1DK6KveO26Z20
phIxEWe7yn2WNb/DHy1JC1CN6HA+oCRWF0ei75eDZ/x7PzF4pAiUg4cwRAFP62Bl/FM8kF5Y00fc
EU8mnkvvl/O72zQWds6sgtRVnHHShOng2Kg6Hj1upuJItkasBU8FEWS+fSHg0/4Ta0iz19322o+5
VB4EkM0LjNRqK5EUbdciWPxVKqQ/LBKqXOykuQPnb35gGOIjl4w+k1Ru37pYiHdF377MRcfmU9k1
hL95SBzJ18CwzcK1TDYHw2fdVySRkqhkJ3dLbxS9WuiHYQlo1B50nKHJTnpvHUIlRbQYE9VjuL2l
ncyQkzMfUvXLkOxMR+GhAZ3MSjtIDc95VCAsh2KUJ3SOpLWaVFJsFsM2X3JvSk7tMbI6B8mfYQ/+
LHgSSIz4QMkm4PAdQnvGFeimjeu3rtEF7CiKxCPXi3n6I2KVC1l2QPF2cZUESJktNCT+abgnPIAa
xvmNzHvoRDJ3z9fwwmmAbhcZ56XtshTg1kI2aS98LoY8hcFsi40ezga9NcP6/x4loKC0AV1vN6oO
9D6aodSELKQhb1sTsS9SUw5qnl7KgMQP22EqdFXszpn4nFiiQrE6wiXHYVygjbHK5LWPr8dRtkgV
XXcietdq7jGujdtfD3DQq5M+/SkMKILSfDurHnWAMvvWYdEbD/ifGOMZ2whxqj50JCRre5gw1z/b
SLPMxZbMbpHVtnKbcom9uUrCdXNp9bCuMuvEGbwkDGe79JGHjL2y4GujDXF5Vx7oluHrtdlcyicI
9LXfmD8z+bD96zszyDkywiTMxm0IJY2LgCoP6cB2nbA3aMB1upS+G1g2z7Ld/ixqXGrsO8SQjwZZ
yjwxYBgktpuQb2THlvBG7FskopGAcLmYDSGM1FHvqGjzzrm74LguFedwNa5l0NlOpRxKKKBKp/tk
sLshuywIA9zhK7n+DD3VG6Ul93ZX/FHNsoWay+n3KJHUQZKNT0o8VKkp9nip+AbToLIOzkl3hQ2i
BanoRvLnRtevuV7ZtnKmgj2L2ropcsvm+N6eZeAOt7Mmz0btjf1KodEVP7+Nm4lXsnWpjp7q6juG
QQs5GWUG1Ccw1g0cFT+5VQJoyrD3/dRBjDdAKaIol1Ylp+jmxV4kvfWruBzBx6DKD7/mpFZZnt8i
QC3Xa9zp2uOsE6Zur0xeAmK17sHMSvkWS5JyB4kwf5AAiLWSvTpz4XSFGozx1Ao5IYaHuQFf30/+
5OGxuZyaxZKH3lIfKW9/RgCpOe/5aKMCncstlk7imv+NtJfdBF10ApNKetvDAPqFYjIIBVY4Km4j
TJ0Hf11gkCe+uSLHmKIFS0g22PQwaWxdAUlydKQBbiMSyhCJF2HrfPlCh+BGFInrmEXRUaUA7K5o
KfDl3g/Iva2MaV4iCn8vbsDcZfC7mMVIVNIgywFT1tQzJlSZpMCKgpc24Y4QgLoYUZgn+pKKHA9d
1hd5920c9nzhgCWwdKduljRZ9sbZiSJiy+3nvgXFsvbM4XsArl3pSnzKxhxbmFQLrURcFT9Z5YD1
Teyo5rw42AMwT4fe+9Sd9pORbW8h+56zRWuflGAdIznCd5H23o+rAwvvr/oCpwTMKNnMDpdE/Zxo
XbeZsSSelgPzNBE+fDQYMW0RfLTE3201zAm51xx16i6cEPUQn7of3Kjhst1zEPSWmNe8DBLPZh2u
dk7vJkZCxrJeGO+6xwkoY2gU25UIhc3wfyPBebp+4USQES6q4tFNkqAntbkhuXzNJMLzPmagGY/W
HU/bZ1ODxT6x7mwf4TuTgfEfGbrFqzkaLW4hPnp9/RBlwmqqu/JrAFF+eJ5XvDb3/r/g7SoWJzio
vW416H02/zDJoteneCEK2EFu8DlSZJHT+T/5tmLVfvwM7WVHx8//AuPizK6txsW7feld3Fc5qIVb
nj5LQgar54ntRSVdlztt1XkbGd60GCGlSz9oqxt2VgnwOarU1VKqbTWlElCeuwUOOsg05jDz4iB7
cqOG1wgq3E1ufXeVCLAG5As9kTe88Wcds6lZWvcrWeZLkcGHE2i6DWgts19wjaqW/PFNjO2pfBd2
i/GWHPurj6Uss0er8Yl/j/3SXQPbfV7cIPztIuH8UAyEZkjT7D87stztbQYssdYbviQljuLPzvfw
QmnN3Jovqt9TNiABlUTzG/sanP+VWaEqMoQg1pvvYeMkA1mujm510+UXu/hDExlGp7xz/7OdZgd4
vYI/4o/ZYpKA/QFTjdyaAv2Ydn3HRV1xuiq8aj2jaqeQUq1bSgL8E32LaQpUGUcZFt0cI1d7c/Wp
VFjaFJ897LDNjsQnk26/JcmOWkJooMoqdiURoOu2/MPpXzcmg8g0SRldA41pDJLtl45Oy7V8/JjF
lhtKOrfEYCcTz5s39BMl75dkv81iURkHcU0jNzt+3ktgJ9cDvwsN9FK5BePMGXR2vg6YokUPV7Q2
2rrVMeRu42GSqAWalR+4qG3Cd8jT4vxXtbSeJUK2n5UbftiAmpy/GGJgL7ZYO8Obq2lkh+Dngnaz
hk1muPDuXuIUN7oQB4Y4qs3Pl9BKR0y3Arqezg7+YzGl9Hyj+WlQLha9yWLM8an03JtiIEiekCv/
oXUovCsVh9CPgJ9H2WZZJv7VLM6atJrSzVioqfDb1vwZR2jij+VE/0/Lk4CSfDaILWYkZlsHekEB
FO3nwhUfwpSgkQp+NLzIPzd1rEiB0wBV7Kzq6uJlZ22iNPA9puuCGOfF8Ojr85BcV/Fxmm60sjxi
1gzBlWrJgWbrtOTg8wOTILXYutqRLHhUKCl4PQnR0fanlkdBL/T2tNEsAYVc92xAF6lgQhw2rF0e
gQOFJSDo1NTFLxYNz+957B8syLJIvHEFJbsEMFyHCa6l+vE9WX42mTbNz5DNWvWxt8l0nHt4mCJ2
zSOXfvwM3yTaeJS102ehIPo8Q3vTpTZqyvQ6tLpwCWTIkyWCWx8rY1wwHn5SanZsm1TT/QaDa6WY
NFYfOAI5X+e0o6qPf8gyLNWboDG0uMege3fZaVLaU6j+jS+rTTuN25d4gt7gqaJlui9BBNe8wlGC
bxYXQGfrHFHDmaB86XiyFrv1zdem59h7pE/SEQ7sn0GrBBledWtG8Ttax4+H5qdEBPERccobdviE
Go7eltjq55HU9lzb4UJWm4suy/cfB+3nlJ1kSGKzDmtfd0mItDUFhSXEzPWJ9DHWlvGR7l3LjMZS
WbJW6KvOu+Z37hQbVqakoJcPWIjz2+smWGyzGud+Tq2Vpz7OFLlzP0cC+RBmJpUfenxNHPhAXNIf
IZgdBDF4Nkorqfb8PVMz0vC4NiVci/sfARez8ZuNfx0Rwsw6N2GsEXruPTqzRnrbq5wn7wVON054
kr5QjUDIYiXw4KymeDTlL+vDw7BswbcsCjZMOP+FkIe5ahie8qwoogrq9vgcOLsktXklU/S56EVp
Ij3RYnM8FZ1QpwbCSZ2QJSVZTaGw/lRMqOkbzzSLwjqhsSOBIEumr7um8s+qeEijvNVBzHh2ymKd
lmLyO84tQyaT9B+D+dnU+TRauDbQHo7Dn3548s2JQ4CTTHWVhA+cV2eJEhw+faE3bYkcbk/1KWTd
S0/v4upKp3evR7xMI0SZX9s5OOTw3lPnapbEjVQzYvYG6lPeU0IEnOdmSMneyh0s6hnvrFM/bSH3
CqaVHdI532VlONJllnz9pOI/dreDnRN+l27lRR4KI3i4800z38mg+lIcwo2C2mm96BqRSKjU2oif
AfLsdbFfIgrB38nOMH2/W0OuIQ1LTEqRo0cl1n/33Nh/X+hC+PBriWBhaDePd6ziiZpGOrn8vBGe
D4gW1ehzAKt1pZwBvbCn5QtlwBVgI4bXqhFG0mUouErWpDIiWaG8rN3SVflc3UEJqWDbHWnnA4VH
MRsysU3L8qvpp8qrZyFD5QeDsduQFI6C2qTqL+RDzMNdQHHaArkuAyMLB7ZRPMhhclRVRTORT7ll
4oOA1iD7N4zIwmWwtFHnJtsoZOgAatojlHTwXIjr2Nr/jwaCKzxh3JxpzzntHbMCeyVH8iZMHcSB
LNuDRAQg4tNMapyEYTcKjv1GFa9BtOxPPlaF7PzSIWcvLta7VvZvTNWG4q7A9DS5ZZKEAFAC+2XS
d6kFpkhVOBOVL0BlVvNpMZf3Kvym04OQVOtvif/RGUvDxUtBB8d6qj8rXYeqfgvy9HoKOUB4QvHv
sZPb1iRatMG+AIKxhNUZBTEUsRQqnm+b20rBYWkg0qwSoW0SZih769gSktVchWMuqN82O4nCl8qC
yzTWr/8MRPUM0vOpDgQ4na44KtfdA6oA/14FRnE+U/g4+8CE3dPwoFNbTziMX0cXx/TqMiZL5vZ8
ERtWjWk0btrlnwHoT/ntSOBGkPA1hMXiQrKhJ4vGdY50i0AXFZx83zPVzjiAd1qP/KIRSe5rygxo
lklobB46vuhGHsZ6Bai+H97DmSC0SyMCApZW5b6iv2DcsQOHDMAzC0MX5TgtjsseqnCuD8SVrIRM
VrG99SGcSSE3B643zDX7R9fOdfBsOLrp7ptJZKRmCZU0Pols2OKxSPSkWeL0ElVRLTvWWAcIf4pn
rKSzvuifF4cqs1HWIIitrOmCInwyaKryxYZtDVEpHVJPp8jSfRSU/DWH+5PE22Gki1UO/mDoPxjQ
3iBqyxyMwH3NelaGkanRQ/BCu2KeCLAoF+L8un4etTpt7GINq1RW+51RAVeGAa7XUZs8342osquZ
/20W7Y/srzJQ+iw9pJ7LMwYANF9ZUly6Co/92ooK9yVg4R7VXh+Gr28oniOqfEVld5GNe8A6zEAK
GvTQBo0SOQxi61tf33EbBpRYY2E03vQAsJW4xf5R/sRv5UwV5R36/eSFrY9nRPPcET+LZ0CrdTWT
2fVAU4ETFPPzFCvPxysR3DKDMgmVQUtDlnNNwdDVauDRoUGqGqUci62tskXgb41mTI6rY00iJiKT
lViiPX2Uc9NZmF2wMQjR+bP1JPAPel0ANMwfonx+YKdu17Q6FE7ccENDPiSIjlAX3nT49pYWaNJm
y3vIiNwfvfPA/J5FGIeJRpALbe9d8P3KMcawlhq5ZC/yYtoLWNw3KU8XfmdxcQjYWWLAG8zW3K1+
Nsl7gR1zUpISL56625K41jdWkEc7aPGOixPjQj0Ch8/Mu9vtbcnzuqsz8MqFRn1F2VMNGdEGrCaD
L2PQ5KVD4XSzWpoQu1udV2GWrvzXo56hQPofOwRD45o5A8kcSNXCivzQoNMa/XExcO6Xi+iI6jJJ
U/t9p4lW8u28OIXb4qENGnVKlsESj4T62ohUwroxXsdahku8ZuAsqHWjrlgR9CNTmN1WuUnIk6vt
r1EgqV1YOjY1FW6IpyTLHXaKQvk7cWD6owjGXhlVzQKfIrHuIpiBAKWFNUAB+hUanAxCqFOH30/S
CdmXZZLd241hcBqWwndXoS19Ts42dV0o5OpN5t0QVSqrt+xvkIx4R7kGkozKPfOBYqjE/oAJNZDO
aKihkpnHkIITP/Gr2KUiAh5wY+nZVDs6Cqs18S8MJChEiauWXi00g1jHOnszRyBS1/Lrta8ykbN3
q7LuEqxtZAOJZBejfnwSPUBFrtxHhHobCWdDDLgWGwJQyhPLhnIUgFihUpVDfG90k4ME4sZ6xu9a
ksopw/31AD3yUChc62SrbXcdZrB+LRMuJV/4jkTqi7wtINZhWQkkH5MS2hBIFnyZcd6jzVSbeIo7
iAIQ27EmnTDLEndtEMAlIt1QaUoMGdVwp4XIAxieRiEFQr533cpZ3MTB5muTYm0zd+TjWLORI/j5
N8VOUa6FjVb750YIXQvGHiVMRp9TrLp4rTXXL01WaJPqsUXY8qsWCbCnUzvbM+3HFKIvD8Tj8+qJ
L3oHbbCcHITePj7ujHuYgJiat5X8IcT2PHZYmdpdL1ADd5jlXcrwCT98nSlwVXMEIfSt2hW2utGi
I4LmJYNNu+AHyN5eUIfIpKz7C+FU16MFjC0BWTOwoV88hExqH+oZgY//YC5B1lkGbuDNlYxu3v2F
n8VwJoE2RnIwz61Rm/ePiI+BqeMivoD1uYDSC6YiobvKlGUmg5+C85zeFCAZIv11bJ1xqOFhC3vq
St0EVYf1SYyC1OT8/WwTHhhL142cqE6wYhk156i05hPA2lgn5V7pxhorBQ58rUrdpYdxY9KrHTsF
tFV4hNVUdx444zraxKIXwWUZdftsUQePVqilRpv3QirIVLaL622tepXsKue6h3y1Cmx2RNBgtB0c
AcqHGrHTSgAIwNJWwxugbmM0feexo78CQPWPUtHopVhUSn1Idn7s6g+B4BspegakDj8yWOfibHsN
Na7vZVI0HLVuICdmTV9zrHACihxSPFTDy532+YHOCJTOxylG7MPkiIgi7u7UKNpAFXjJA93TsNTk
K0cTLnAJ5druCgE7FVqQAmAkhW1tNsywr7F/HxBFKzPj3e6p751YZQMXn2b/ARnYaQ5qmC//1DrX
n/C+pat6WD46PhLkML1b59Hg5Qben9eBnTGylFqBQva3dSQXC/nCPwXZD2qTqrhzy9wu4fkmz76w
Ag2GxOP8t6Mis9UiEj75KszwgH4cta7YlkkqIKi5brtp+LWNrRwrR+IwYkoMGOppuqGu3Vzf06oi
GL2CrfshGdv5M+v3v+jfVIrd0OtrB0wo3wEVIMjgBPEoqZO+iQqD0CdiDEUQKYdZzB9TlkIOdd2f
m177zG8INGIyzOvwDRwOpUZLdth4eg9aD1v658c7gClq3UqYj6zZLNYEcOs26Lc3hOH1rn1ab7no
G/EtftkukuEMFnJzrxtlepZnAC+xAi66GIJjlpBZPXjFSN0xQ7RS2R1CZg69/1UA0YHGzDSLF8J8
TnMOAduvgItf3kiDWfZ//L5dWD6QQo4HMSKj4RH4zAnOXI46FCI+W+Y2MqSmNR1Xh9XmGhJlnxkT
hhxfAiDNmaqF3NIKxoc33F9jk//VWgbEmBSkVP+puyfd7gb6mxZW1x0TL5sDX5NoYAuhmR9JzWKy
QbJvg4I7VHE5UW3gT0gXVQUAoUNpkIop2WSKRc2UygpaQS3ES09Stmjevm0ux3GwNIHnzVy2sZWe
+Rppf+ZZHkz3rDWKqXKhnytY9csIwAiRhZpQDv+T6cCqzUqe4WDArWbR2fEOFVhiKiGid5ddrb3t
/xbf/zNnwTuGRnO8AlAI9/SS4/hqD+9R7IYeFjGQxkn+MwsRfbz2J0tmarhnOUMvFpuJExcfolke
CEzq9V+OS2u9iPMlzzN8ZiybHEOVdiOkiusdoaZP2N/xz/05f6QGjjJVCDX5Nir/sk1O8S4gYMcw
8LMQNjFIcdqdqL+82qoXphYA1ym8df+qhWQEQi+1EMRxsBvsDBn4Sd02Cr9dRq4+z7GnLLzn48sF
p4lPJVEgNPea3ARch/a2HjAt+gAFfscncSHRIfkUShZrEshf7kub8tZk+iwrQyVgXleIN7/IRzYD
XKft4Ex+/kGVDmsSKLIeUDHoP/l5ZQFN7+VGvz3CsHLnDe3MlHt14gK5xyVzqK/ZIlYPcpV4eBb8
tDk6ydQRIfWNSef+rK2F7dxc2J+c6vpCeagYl4G/SkXFYDDyE8YvYIg62ZVbLCi0TR748fKg0ySa
QXW2P2HX/mKjg+QZ/C2//HSwQ26F70turTCjiIEefH0rd0+GZjE3+QCpw7+XAKqLqQQyKG8RFtrk
Gr4qSxW19bZlzfg2Ivl6i/VbpWRWsJTHVcmcoehBfb8SQB5ZZf1Mf+4B8XxUuoO8oFoaLthyLtd9
UNKesKipj3vVJxPRATvwbko9/eqvh+8n4obtPVSVoDHU8G+2wgrtdHW0rrzXRqwr6PQFKVKt0i+Z
oM0bi5z5xl7rkjmm92M8bREF2oxP5Hu+XgGShuzLpGU1f4p6zyEBoZ2AAYqgySWct/fbFVqoZ+Ts
adl8fIp0qs6Cl7IUFA2V1vGly6yWR3Ayemez4Lytn80tP1J3B5+Db0Y+q3pzsy/Da2Nj6dL19Fmt
ADegsbdHXpZ+Oiag6MxcGPGWhoC/JUAAoU7zvWXBiE67hJ9DfFTV/Dyk/kfGGN09WdfKk6dVB/ke
fTy90lGaBKwTRq8LC0g2YH5EgAp9aHWJ0LCGaAKWyMhVaOgirjnyzEhSJewhrGjrl6kehRTpquuG
bT5vQ8iG85+7PLls2lF58xR4ckb1wHbcFA0V3kchMtlZye3X+NAjCO8PdMt9Mz6wEr9ksChhyxmz
n38AmTeomvTQ2wQJLbHeXDM7HQVqXtRIIFQ4J1HIeYjpwgxH23BJxX4FkEM7bnc552CW6oJQRqwd
hN9qXN28yPI34taFNcLcOzU/+v6SI6dzyKHnfKyS7Bx+XIyV3e0Cw5zIPANsok67vl1O20/G89Qs
M83s/b5V/QLiJOUGW0FT1/O6W2xRajsbhtoXEUz5cpGI5cZCjlxvqHrIuD04KFQSgf/q8ZYRZ9zI
DgGSGDvQwKLEgOOQ16oTpz7Z0oG8VCVV6TD4UtxAwl7AZDKflZMpSnG3tyW5+k+XiXkSbn4p1F7A
5B7OpivHIShNdRDusw2IdTL18CSw/J8Wc7xf6+BPSTevrEVtP+H105rNOxxaES5j1JrOJNXc4syR
5BJPcn5WlEX+SJHIhaXx8DDcmYK6u2wgAmVEWgTTArLJ4O5+qhrJ6YHlbKGXcUzhIileR6E7Fc+z
0l1AK0bNgwCP2r9jqPXC1/IT/X953BvOj+60vUu5Ze6zgBxUu2Q399Y0t3/EAIsiGCZjXwWKcAII
jfxlro7yno9Zs5A3J5ook8q3qfB2hkj3Ivr4g0gKFRj3ZPnzkT7hRRJGxuszuJMaxkJRUNnsmWrO
Do1dbTVmHmaw+4/5Y1Yu1dhXpjwHs5hyLDDrzgVmofrcNURex2ieJRjpB3h+eY9CDF+CFmKvy/yP
ITaC+3Y/+jSPHLh3OBBYgfxBZowV+XeZo0toL4uKn5ZkWK0XyOt3q56Qd7T914EKIqECavAkNyMN
Rwfun/LN2KSBnCXvx7dL67vg8I5VL7OmpEhdNwxohgctDlLrFJIA3PR1Aqg8lyI7AchBuqsIVuho
h1amE7B5NOOaPtROvKIzv7ykpLQ5W77ey8NC864FoiUNRSTLzJLBKVAwsKg+nQ4rwhmNa/zt+x7r
vmVSQDlwtJAt3mqg5v/9MzBRfWca1BCNvZILVb6XkZCVJTcx8HFdCyFxHnM3H2QzV2fkQoU8tO6H
j6L0I5TTx6qC/SV3kcCql+iKzUE6EubdldCypXtG8U7CYTmGCOVDQ0v7NUYuXXqfS87yZP8zuUGa
O/3T1XQq9zmJbjWaGuKXnGLVa7VClrHvnOmz0yoJhdbkMddsnvTMU0lZ5SCNDys1lq933Bz49XL4
Thp/61KYt4s2rDy71+DJZrD/vuLIcY7Gh8b8ibtRKF3w9RXlvoM6Qqtpk0YAc9TO2UGTCkfLoqzJ
ePjZIi7dUN2BL78JACi1jjNcaR4ffPbuojV6lBoUK9WHzdA3ygOm8NBpm4GKnozqbpG6ldZACpPV
mc2cJD0+Ui4ScfwXYJCaA/1ZWr1Xu5Qa0ALNi9e7OsimT56R81V216EXFkM530y12EikL9jo1+ki
0jSc3866UypYHHo0v7cmkasfwhMK7JDtyehf4Lhzbe1IXNNigbsXUaw//gsRfLJPOTk2bPNCZmWP
n2Z2SiE/2FJOmuBXVGCqiD/owP9wck9B5X7Rfwwltus4UZLqWU/7lMBqcbaymlB/nyLDIZehZ4i0
qNSj8OfbEV4iytm9rhuo7+wXATqeYdnLhKHv5k+JlnzAMYUTVDvd+5VUHfTyQz+JjiwkgFCE7UGg
89y/lJCJJ2LpdzhSX1DxtrL0ZVDB/VgPzXOX6r+5ZwXTlFX62P0vZozdJ+6MFCkUM9I59qbCb69w
3n+lqAGz/y7jIXhBod3bKe/vNckzc5wYyaapUlzvgqWN0vTat0NYlTdIjqFpqtsKOQNPGGxCWt3q
9dqdTw/sVX+W3XyfsvLgdruQheuzIgpWQTMOEwP47ykAAGBuZGJeo67NaBgA/TCwRE09k4gpLa6w
yW0BlRraVgiqqAs7iybTDoRE72VLsTOy+Box0dNBw2NDLN8pBeQHkugMcHQ3KQ8B28PmqDUcwgRn
s0wGS4nXNXeFlQ7VENTKx7RMTwHbtaTz+EqbHiLztSlUznNZVE6CcF8Ey7LyEpxiYM5E7y4T17dS
vubAN2iS34tSFZEqX1U1lYAK/KWHRZSkRsisBIWK9ate/oyIu0aonwfiE/u93t0F2l/9K7kUjv9H
7/S2Y8kVKN0wMCJ0XpjNG/BsCghQpZowx1Ar7NHHI5JM18wLjPMY/5R/zZdvNmtAmhw4uuLWNFEx
MUh/rcd7k663kn6l/1Mr83nC5xuQOYpU9FO+nPPNgKOzsWYEzV2LmACyWcB+iUFpjoct4G+dsyQq
9cysir0/7MGgq7QWHHxWt2LIfjsIdcCQyeDN3HB3JNUVkiZmWg0P7UaRKiN3b2lzQ7fE6y56rQIg
XtEBrLlj7nTT5jME78bknPrOdqD/oIuf9yuUPJKZEXnBWu33rp2tfpcPK9XwsgnqcleoJM2gSeCi
UjPcrcDrECFQSBPjYIWvHPqHK9AEYrFSfP1Iln5NJSLlfbFQpN5Jw8oYyTjzkq4eyZ/CgqaO/N/b
VlpUTBYA1CDSCVLUbbBJQi+RCDzxR8alfMALSmN3I1wi8Y7P5l4RkMEonGnlmWy5NL6cl1A2nxzr
iUG7YB3LR9HyDFehtWMmG9MlgoXivDjzdzC5fQDFS2tjDkBOXUm6oT+L0jLlT/BAxuX2rGgoPrLW
SZ25BIS0ZKakQB+yxo1lmP8WaRLphIZQbRt/0ZX2/feJPyswIrNvjpbDxgYOq2g1LpCNyLjBc3pX
hGjEtbqNjp9KDW/Iid3Hiuj6vu9L0688cq6zZ0qohL0gWObBVmrNzY05yyOS0rxP5yG2E5oOyoqz
sXwZn3fPHti2bHpoXwCMQFsZmAx/N6lYhkw7LrKCRQm12+VPyn4YfcVM7hf47RV2R9ODboCX0euf
thedpDFMQAgqRK3iBjNTYnmTAAybpxyzuUDKrY5jHH00jyjX306YISqxdMaM0OF6yaCGEgrE5TIU
nCwyFwKNU2ZwL1uzKu8fAWU67kl+RKopJrAJGGVeEPHaNcANlWkHvCQvXXQfi/gJxd361bz9c+qg
C7MT+A5uivWHELSpMZh7OFBadE1RFMchzIl4aPlW4UCFiM7iVQwDXSaAYvtU/N61SD11o/LzeekS
p5cty2Du1ua4p0JhaunkyQx57GQYeQTYT5flC1iB1cms3cF/fTKmrYRSfN4mTN/LrjEir7Njv1ru
pt8UYnI9erzvCMFJEqB5uV1g9pt2PP0fdrAyPNgT8aRDfY5yI/v/njgTh4/mmsd0QdVr1rPLGnHr
Op1Ykhi05HoML3szjA2LSyofQ1PP17LAxbof6JkVsdZtJ2EZbiGJC01h87TGKAuuJEzRkWZA60fM
VonUIoCj6rZsHyAmaerAPbTyrmWHPHNCd4+Zg3zIAJvGe7leElwS0fW+/jUHTyGb1H6FVPDz0gn2
4rK9UVlptCuyEfOjjLnsope4EKq31HqlGo3rNJgdzmin31jHYYx15ZvpD+KUAmjgUw2AZOqXWYA0
PcaaN17uHWqsokNmIl00H9Exzh++RIR36GELOQ75WNn22g8L/pMrA3nOHsvlgfTIodLWxwo9UAM1
l2xiwQ7NQvxrzEzOM4qZvgCnMtDL+p6lt2oFuLMSijFrJdT2QXNxBtOx6lbj28d/gSpzCDtAbaNg
VjCEt8U6hotO2EpMiKh8RnMxTwHRCuBdXfcsbDlIba+pto8vqsZ2IOjNicxCXXoZSq0EBCzjh9nM
Nw0p1/GlBM53+84mLy3HO/3e5yX2KsPHI2J99ecocRS5Cep9BDGleaQefavY6jLbOqCnVwc+KxUI
WnH8zNvdeKk1s9eCejhfSmSuG9yBckpxTs59k9b9U0efN2J/qGKVSUGBZSpKMgGlapGgyah9MtqX
OkpQJdgpPRN3AzMnmQ/Evsg3Vr2EFAjujKaUekUc3bh+FLwsZhqbrpCbmbiLfmEsTVz7JO4gcwrQ
HGkujWRGvx7OuiWkmpwqMlSz97ujhFlejopPoCCn6HmkkXyzAhVNhn5fumRJtqOTPe6Jnezioarx
uG3hT01AX83kMOt5hSHoH+yRA2WnRsE2v2cm9AJA3a7UVQY+O2Tx3nKl7xj42L5hQ28TjISB0d7x
VXI4nTU4Z9PPc+bE+SaQzawuWwf1kopDAwB57ATV3HsdymUsiY6jZC4uoEpnK99pLriITxl983vZ
HdQSdnHVdbjxfPfqbiTKXvljBIJXFFtJzcB1aQ+hiYW5QIKCahxuIhwNp1p+cxEEUr2gxeL+WWDd
SUPHgzxNz4VYAcuI4qqmthb8Vc4KP5PtHNIdfnN/U+LfTXtX4ni/MOtaXWrGZth57fhyhS9ZuLa1
aCeLvS/ZWMcx1/nqmgTU0Ro6+t52cQNCPrPaKgJw/eECvcvp9e0JpN4SQmBWDQOaz9vcdSeEBdPe
LKls6AaEJsQNs3vCqtX68sUfj9491QFoJF94oyVkAze9gBjoXIpLJ1IQz3GsAKWbtSifExNtUHoN
ir43BuBNK/OUs0NtR3D0dzUobAg0c3Jw9fr6f014b3IFNFsPBS6gkCG7uWO4zciz8pB0DaOeFrhA
KlT9iRIwi+qjYqvXH3+GJD9As0NUMNRdZCqOJeEwDr53F5vR5cUaC8Ako8vzqzjjGiJVOVliVGwi
RvPG7XfaqPhjPXa7SiZQBBEoqwaKoZbujWuecLebQYwH7neOH94ItlVTvbCaNsGpzN4VdYA7ibhU
7ekMmxTqnXwHf/uj1aV3P/xwAhJ9vphaL8ect+R7AeqTBOXfgqRKZIifwGv7XB6qFW8DVmEmceFp
wj8SdTlLnhJFPhvGpgs2K2wdTabfFqgB5W8Lkn7Q5hKPaJowO5PAYL9Adt3qechI8xubsphMnsmE
cB/JkerWCIBuvUt+dmYMfAxFHCp4M3qa5h8bfpXoc3UqCysSGr5Cr54BjGjQfOlVxR1Ufpm0TV2d
v8Y77DaPU6s4HZdXwK3yqzHaNif+XE6GwhMNyABo903J1iHCSQL+Qw8wEoQykROujhwFq6P3rCc8
CpO8nJXxd00+AkOozlazfWYJ0xoDawWxCXmo6YD0NZ71ZowUJO6aX5aZLZ9XexZvyxVXUpOcjHV5
btqr5oOgL9CI5av4ogysgshgoUDlAIDwV9W4n5dRyCg6wNIfkZovd7/lHyklOaz4SZutbYGSgfDr
jbpUa4641MRn//1Zk4A6Sc5UWKXydxk3tZZwDqdopvJCqUybQuPTSxiWzI5EkEQj8qEnm2vbPMS7
LWi2dd0pFRqRn+viU+iZLAFOUqmWPzDZe/Ms/iL+MyQ1PxvHLgNearplBsQZr2j3ij5n/ocEQyA4
sf6uWBtjmPJkj5GXgf0O63Brvv9FIfVgEVN/VWAB2toTeYvvugBydMMRtijY4uC3oOUluFwRNctu
/8Dq/iwo/PNDWNoqqpMp8n4wUet1HSjNwQBq7X0OB7cJtuox7Gbwi1bvq6ao/CMfB2xPgXXo4Ang
QavxndOhcDFU3u1edQ3mQM6Il6MwcoR+9ZGLQvSFyJ22TYI2inl1q8amEm81ih6KCuAg4+g6LhW+
PXg2XMP1L4L2AY2ZjvfZ8pLTMmbOnVBfh9MjCB5qHRpv/JubHMNjFawFx2XZN1IaV/8XABios+GY
yGrx9RSSScsluAi5nBzUWWmC6me8zuviiiH70TysagdhJRFfPYSi8+j1K6LiI/Qu4KZfpq3k2+CN
Y7jN7rjVbr4ikssxScKmp8aLNbheWuJqclZMhVKh4t84n+M7jlbEuEF3iGZ7MeV1AZHyLagAadIe
xdAScqkJ7vGqF9ic4pUZqWtDtXJjZHvr5621jbgm49dRdCtYxT2H8WEUzVSgouMQBmy6YgfG6vc1
rl/mH+GoQ4onnJOo1hJKPh+lYGlwiaztU8LjFf1sNuQMMEQTB+SV7AitG5POjI8OZrdHtDnPFB2m
MsyGHMdV6DvXMDxOLRD6VUWz5yzldJb3WLs8+DqdN6aTIAOU5B4a0hVKiOe5b55EqlEKq0F+kqTw
oNTny1qmF6puzDQmQmDz5Ial3k12kLA43CDEBP9Vt7LkRpI9y+uXA6KOTH+nBK/xpM1OmBNPNKRG
T7npAaUSFbGbd3t7mw9O9BEQTjnPerbG+8C7jZH6Vit1vH1amjgr3Wfly/AFty7v5UHTni1n1IQy
ySyERR61pK/9bWv5lpFGipmCCqK7yuGu7DPWuFtyn6dy8adowsEhXz7UdxZM5wKEMaNqxtuLc1R3
rrUWWb0o0iMCv8GzB9+tPokOVbNbg2dzexEnGlF9c1hdpOXL4kMnOEQIaQDejQyJmomzUfpLBIgP
N/7MAOyyK2wszfDtBD10E+L6Nq+3BGF4ZKeYeNDyQ7vOGqUNMao90cEcvHTb91KOVBQbmu3uQ5E+
1ze2LW5L08ftHiPXQrVXui5k/1dC0UhTXS/mx7hDs/ktOYU7kPc1oRpi0iPaJNGB5EYp/9dgiZlV
SqvSNmHMct5n2/8A54gVSYVXTkxwk7PKEFT1r4jD4U4FXSpG3xZTJFw2Cy68yAYwmNqJGlrDIDQo
l6hQYb2cRzvSEgRGm6AsjFdrTJeUSZbUIZbT92sHyrN9QZg/RjEp48ae9a5UqAroh+KPcZSiR5Rm
bj+CzyPdbudacqABb56PK6xHybKQVoSY1k6EoIZ5jkmLYPwhK2YFT2aa2UhTE38yiRY3AAFTjpND
7GddHQcfKDq6HXHiXX9Copi+UskX0tH6zNpaYtqJprpkmFy9wSIle3dF6XNpQGx2h5xAwCScCTgw
VS0XZwmQtpXAk1nzrwXg8FM7aep8SqxdYrPn2xKh452xoTX4i33z79JODPcbIVde212VqZrV1xEa
GItx3lgYoicwLSfl3DMUVLEAdqPgL5MfhjEAPrSgYV3IhfFbh34ZIw+NkLqBrH0RP6Y4nSnvGdqN
VtCU9Ofq8Ojf0MKQ0+xTc8aEKjBsqroHGJTCpOCKsBC/aPYwFsw24Qbnba4CiwG1R+1QREdHVLhL
inPAz4Ei/nmS84l31wHTWwgBFTiYib0dXkzO3NFSMVWDHNZ9zLttLMSUZy1NilNBfFiz7fRSZbME
gpzrauHqi9PEEXJYODqg98HJWRtGYdF+xbrZYhczOTaXCkAQ2torp+HaFrbSzwELeyAkzUnnzOOI
DvkJW29XNzn+mkmvKotPzoMk6o887njKCksSZY/2P0beDwhFMNCKKJFejhG9Qo47K/pb7Rx3Htbh
z2cikG/+pRoz7/HWl5TYOBkUJNhXitqUuOBsZoXmxHrlLNc/HM9YQblZpCZKD4yWf+kKDMFWblcY
lrdVCEADfeV7YpuI90rzfawH+CzSX9rQZK2KJ2dzlMKLxbWbFFaK2xQX8qEPzbCKXhSK3caslKMr
e6gm7FmRwt5AYuiuD5uLQrgSJPk8nL14IgHKDps+LliihBq2/gQ+zZHhUElmxTdRJu3HEZQLNFoq
AUJuPBwUBi8v+4kkyokQC4Yc8+FqOSzVnQAZs5cYTRdwK+NKpSd6YgMSLAixnriNBkBgtkFCfBGx
sFn9iayjKy6M5BUn38LPpe+nYIzUy4Ntn3huVHC6TyHQrZFDCVivm0rU1ONNZfL1LQwvfDcYAJy2
W3LSkAfl8JSGuggO46ss+BGkZdyQtlHW1xIpgEhewaKiIFuNJaftxQqlx8abMJctZKc6fjw25cUq
v/hOBl4008Un++f9DiTcUNejU3ev4sTH5h1FilaDRgCrgfYG3yDj9Z3MCF+Cim+wis1ccDIYg20T
7K5FWf3rTc1lEGFcK04JQNDEBPyspJoGn1WQ5dhvW/M5hm10p+mdCW36nHNdiyp3zUUg1k6ywirh
uAMYWazJLZh48DgJiASj4icoygX2VThtXcO/bydqVSSnZuO+JlleRXQ46dJXg/rrY85l1TKUst2x
RgsW4FIFmYDxOTsb4QY302vEgO/XGSiiFs41yFmMYHOohEkmWv3jJeXvat+69W3oprCtpL/7oNZy
X6UqjOhfytZ+Rh+43L9gmloDpT3fn6ascWdUvCCaC/KwBkr6nIogs6zpUZTxzN5BDOL2nDCPrO+5
hk0R0RxLIg5sYvMVUp1C9IZ/u6VnAdVNOorAYCcGNTrMcFcVB3ulJSbftsq0xS2s5pF9Mm1pqwAb
FUtnda13B55WJxueJflbvVMrH5IxCblWjHlYgNy2dS+pLO/y+eu1XSMS1r5YvRfqHi7mG7HUzWGT
GV8BXW7b03tUuxuJ0pnp8tTN0q4m/4mWWHezCVAyd4WOJmspI4zjmJlvd3CzI3N6C5RyEitiFm6g
bfclzk1WKzEwj1lMhFCnJg+upbuzLT0p0MgASxC6KCKN+IOE6i5hcQUVEVrx7n8sjyI21NpqJxrw
vaDHbH1gkEJnaOkW9/o9FBhmAcqIRqewZnlgJbLwtTBJnF+SoBL7tGPIA64GSLRgufAt+ZRYejf3
kwrBHk50Ak/y+HpkzDI5V/hsDShA/tN4ul1clEI+5FwUuQ+gA+BKDLf9mU6mRBTDxq2X38oMWFUK
Kw9XUF/sa98gL7lcJpHcEHtKTcB1nDWUTIt+ipIDTelQgNNxiRtRVYVkjzdEeEYHlwIzCc7+RSh3
W0CS9gZ5EYez/eofkJHTy1GCyxYX0rrxNg9/fjemaXXPuJ8i8c9bLbSOdA2ADq2DlDByFSvVcW6l
Dd316aPQsi7HpmMvgDzXSZmra4cfjvet/RlAjaBiIjKkjpLrXhMfIIQordYfVSlL74W1k2DhvHJb
rP5j9PvcsMSSBc9T4AcbCp6Y3/pyZJvXMsdItxD5+kdnMqx25nu3CTQlyXwG34rzbqMecgZQkaYh
Ngf9HmRiWN3b7ulhKAvlFhQ93k7gWvnvsnjoSgtVRbidB3AOthpDCEICbDoamiZqjfS1dY4ccD8/
zGLTYbcLcp5uo3qTJlfTLKFNILDfSVL88O7pciV0rQUWefF0W0o+nLtZmeubJfoTFGCbFI+gthuj
oSDw8gG8tM8v2OSrw3N2ZeSww4BRGHrwhZgirSQOQGfrgbP9F1G1xwVb83aO6Knslf08nKna2XfZ
baT1uL8AeKsCJUggkuz2VbeBd/rtig02VKAsTJEqHQqVmL44MZ1YmzlaBN0fwxV5p2FCBXj1cIEw
6K2iY4nyis5lnWK9icOL625OUYCjQksh1lqGLM5sW0kM1zm02puCe3m+zdxq+BkHQ4vGSNKIQ093
DTgF8/u2cwJ3H7RPzMr9q9KgT85srnB3DeW6HZWjdPXIbtxT77fA/2NxOSw0TavXuYo1EZ5tVkH5
RSE7i8Yd6WrbCrH0cFddglpP0WKCXoyE/clxIQDjzHTx7M4+gW7F5SlE9MT8BogLRQ1LU6gzua7e
RtPtHoaaV06e/94L0gp5c5O0BAjWymcKENnFJCFItU4EtEwk+PQjJtscZ/XFf45lPQVrdU3/O1DG
5FQSfYBBJda+4uQRVFvnk1bL9eGLRdNy5b1qBtCi5ELGj0zpgQGb8Pua4D/o6RNIrGYoooK0QzmU
godwxKfcVbNsMmdw91PVv3nZwxbiDXWFuO3Yc56zSZw1VeZQnGhH3di6E97hnoPl2rSSU7dBDouU
HhNm8BTt9EHC/HqvgiSdEK0+xc7TjetIGuG+rXZ2F9TM31JtmwJ/7KRKDau8YOdQFOG7HBIfwVt+
wuq8cfvBeob0t9mW4Oa4uTcByo9cLmR20jlGrOi1TUKFJk/HPhNMVeB0yupgNMK5z8txLG3qFQqR
Lb+zvxE6TZU58iJ6uUhXccw8Pb2HWelcHbUJ8RNoFzl4M36YvRmAHAgjy0b9uxgq8QmJJg+nLhnp
P5z6sEaYueL5BptPP/WjIC3LU1praT3YOdAkeNLLfVuazmZV/4kAhbeeJTfRpfZwC8AJPN8ZpA4y
OafYrCln3HbZTafh9ZW5DbNIVafVV8LYPT2EnR/RibsM5Vmz7FVoml1uyQmVl0KewMXlKGz1Eqmk
dT9gpl8+Dq5akbLyEXcrp7R5ZXSJmw3Xg3feuX6dJKUsPhc7Ks2vq4UjEzJWaTQuEFqXebU6KOsx
pcdYml0DWgWVn5dqKl+AMyLWcHR4dv4EtcB33sg70dnVSN2eyksWgwKPge0jM7eymVIBSpwmfALZ
Wnm0KzMRQtCG5dCqeZkB0nb4EPleUgUzFJI/o8gN9Nsq29mrrRp52M0i+bEzzY+kzuiO3P7xoVF3
RJkWNSdmlYIZEHqE5VEDK1jCnbeB/Opxf/Zjh/Ub2nIgfTY/zcT2WpMvsDbQ5k98UmShNlbvQvvW
IvcrACLUkMHZVM8MHN4SV49AP3lrvYW90gWH/K8vJyY7gL63IYtRADdjxGeSF+dwZbMZqYMHKdy0
LzqrifY7/Z9a66hS7p+mi8sJkC6gubRNzUFZ4IGo4jYyDFuqksle3F8wfEdkYxZlehRAWIroxxGc
v77pRWzRArCZRI9BLEMnEjIaQRnHWWv3jt9pDsmN2twWBSj2cHA8ZTvX/GVKNtjrLLIUa5yotITf
vh4OY8CcjhU2egggyt1oAkCQmPwgrLAM7juUACnLodqXilq/YzS4P4bj/hUQbzQ4NnUz9OkH0rHk
uDJ5hpt8NWiRq7GKim3IRtYR9J2XQv5Y3FG/xxOVDQmUl4548Bb4O+WadpmmKdio5Lsny7nau8Y8
V2ce35KwHV68LvoRW4r5H7PF/Pa7QmPocqEeirBT2qG3f7FYXcmnEKzLl2Jmzq8pgri80VADGGLN
QUjLQfXxDn7mKX39LjcAZxl3wM1c2S+kVNZ895csMFl3XtWpj1bl6l/sBTU54t3Od2HdnoBSr15C
i1AXLD3YZ+g7xwfALJ8lHdGkCPYDIg5wp76LhchuAYQd/RpQgjUiYUa7JpY1NvKQSKhv5QNLv/9I
koMzuMN/40QDqiS5v3SGANYAf6NUMggs0wRt9VaM27XlzHqFLizUqAivNbsmyl4xParTjnzHlKrY
5ByYslbjMRJxo0EiWIhTcT00h7CA4pbPLI88TxYRPRI3vVLyh9iaLNb6MoXrFfZLpQWgfkoaxNCM
dst9xjEBNCgBsV/xc1XGIoMUDykTxAT51W/mwGWOT+gnDhMPMmE2PD6wl1Pb6Sd+8rmsM65i3QN4
3LXAlShfKQs9o3jX2BFF8wagze8foilu3K5ehJp4P9bjIQF5/03itmKLvaQgoLiV0h/916yAvPNq
26ruCZh4rWXMFsFlkKgEBk1XE9jYT4a2yPZgKyz7GoQI+7cwPHpEPKp9WMcJXoy9qWOqJ2wu0QPl
2uqDVVRDObC7DEqy0H8TDBTpqj2E30VGVnwvzfHdqlwjWm/uAdUiaB9UdnkKzWCBR0dXkT0AkjkL
YaaCHVe5n12WSr81TdceQjIawFCoX9nsIG42Ht5Gpf+s4GO1lWY9HUcCjtcG88eurGo7MaZ8LqBw
nIlE5EzfBwVu9dDlxhMd+D0WI8gQDFW7EbwSh7oimQCNMx5hBnYK1sfaAyGJSbadSGG+NUTH13O7
Mnkl3OeUllxDdM4vHcitvlKGqDBBMdWT4PRK5Y+V/7g5NIP5f3nKLrohtWR3iLZKZY6XQ+y0He0H
TLWuy2dQ8z+t2QWUtQYgF/F+5twhfugJ07re7JwruIkCaQq4tRe++qYAIHCl9rtBKCArq8eR15hQ
uUOq5gk97x1CmlOEKYVw6fqq1mWYuZOFooy7lMbDhyIO1ny67tGTPDymDu/0A648b/xne24+01ly
DXF16Dd90wh1nHmf5tCpOFuH38iMqGtca7nNSyiLNFwRR50u+xxDboWycq+kZ+6taNb/hB+JPSHY
bQ0TNKrHba09/d30g3BVGcwfnihMIDxtS4emYiHP5thZsV57q0zE+nnn3b3IU7/iXijDGiW3sr2j
KBgwcKH3+OsHut9xoKuRB3J/ehgf1+5VAAcnEVNLEr6hbdt3QKE/ofk1J3cbzq7H+G219ePmelLb
Qo+p7AQBJxr9H/xEWFR36ZqOxiRzaj16jhyVx1lTl4bEip6MyR8jiHYoTJ2UUU4zRTSSdOPa9aV/
1ruaLv0ozgUb/tMPyHhDCbEGrP8a2xCIxfOEzsdAcTsLAa8rulXLe/AyXGcXW7f1gT+XFDknipMF
LHJ67QrbC/HFa7ssxPfgbV/VbtCWGCyPmtiyxrNRm9IjYxzU7t3Dk/ZgZ3oFei8t0RSh1zPJ0gS8
MvFp1L4YURvXdvFN3DRauyses22dxHp2zW1rNyA1lJOe0NItDGzYQ5DO/nrIAARCW0aWYfE17n+Y
cLValm2fv2eRqByQm/RYD+LXDNt3JvB4ydnp8f+LhyCu1lHUnVB/GmnV9uYhKRe1XQLLH/JbYJ64
gSZ8fPf/0cMkKA8TkZ0pn7NHbi9puncX/HK5XX70Fghq2arm9GtIf/PVZPd8N9ly6BzKPxnJ+hL0
vI4IX4C2ozXSJSCTT6n4JefrhufZ3vTPPXKkz/XKMRbqwk9SGfkY2/i88lx33IGkC2yQozpGcZ1T
eAU8EMCpPB9lauYtxjTXV7Fz/Q7POxDmHbKwSGaMAQkwmEI6WflwOtmhEn86QbcS7fO4HEb9vJJF
fUmiiL3NDsD0qqO7aEDFVGn7ZNhL3SYBikezfNWnmleGD85fDhwc1eEsz1inKcJHHPBLzsmTYbj2
WSTNmw5YBjLcHadVzV3g4D4vdCi+f1Ki3OEOth9dl8IOn6e1fbl8IXFFZmr66FIqPcJGZjkFryDE
RhWcinky6Ai73qKpSDaQYEDMXoUQpKrgMu81ouQ4Nyy4JSQ2/DNLYeHP1gUL3sP9/y/khF2AdJES
cBEFt2e4wLjNdpcUBFnW+OUNb8msuUJ2DIWxVhGvJThy7dLsukcDFIaLkKx+DBjUoAKxf+QvMIiF
LrF5QRuNMHQjrIYdverwzt/KAyEy+ts3gOcuKEbUp4v3FBT1QHnkAQhtf41R4D0upkt5U5WYiAg0
w6n/e6Wn63tVz8c7Fm//6cPPLid+HGhVEh8coEl3Qc1k5T6FE1A2u5kOnZeB5+fF8ckK4aJ/ucQ0
EK679pgnVvBdV3l8T+TdEYoB+/XFx6fYVToJ88zbe8xyP3/2irSqhYOSs2VXx9oq9SjwkIyvfGo7
KfiSpv6UsdowCZisyqPe7FPeMvbw/KLdxh0Cwr/COwzLKOpvr88Sn776/9sYsR690V61EkAXsQfe
H8Qo4YSSWBs46ns9HPE/yABK9xD7cEj+iR86oST3jMjTNIC2VR1dBGiBOX+s+HtCLcMIVpvRa5rT
MBmik7g21hRb84Oc4g7GOKZzo2Yp+QzVJ710J/PO0WWGlv9cjO5cOenRWN0km7pqouZBvFPm75Jr
TzfLQIFM6ki7eD+NFOsEdAXnkvBh7bGWg1F3t55eecfONRrrhPVKTGWgGS2xhwrgKzkfTXg656p9
dvOTX8ai/rpVTuSST+KVQN7OuMdzVbkqNgeDXEPc5KA7FwwP7fXUK6GJ5DZmtsbVnBV0QI+LZm3a
fnSlZT5onBbJ298mvgcymNQf24+5Je4wzAi6YNviEdLkUl2ukYPOHq968k9aG7iNgn9kyXFLykih
pge/VhNMXGR0pyyFHcQIJk1rn5oKqg+xLJ2fKnko329pw+skg5SX2Swy2hTrMhSyl+6QszW9VCRn
iNzcSxvROuUe5HuYIsEpxnXMKWBhfHJYQdsah93C3j2fRGwdcNOz6stvFs+76XlDfWGAyIVvcLeY
4uiv6KH8MW+mxpsYYMwTRPTMN0AVgBAazeS8wgzNZBQGYxbzHM4AGb1N8/Zbc2O3dY57J0jnyTB2
OZAW2sSjarvMtxcejc/pZqv3tpRv5mY4tx36XQndE6GqhfbD0qkbqhsD15OfyDnhLZsM3AgDXKAr
86DJMfrtEyYGdXz9s6xEOdZCsTPnd0TEtG6/xiwzsqs2mhifL92ZNSCbUMUXjuCQQl4Xy6MWNHtq
XY/BKD1oAvKiIQOPoFtDxz/vX03I5bO6q4CKdFumNkQpLW4S1ysP5idcXc5KmUb+6xXkCqvuGGdL
u8Dn9AQtAn2HyJPQcG3ZfsG4vyXw1jqL4iT5l2nT1aIHp0hMPSPONOZhFMJI3w0r9SlyKtauavlk
colPV+BePlL6OnBKyg0TZ0fboNCBprPePOk+VruCG3FdhSQXSWNT3EPO2KfMwKHzDgPHk8FLWkuG
puN+W6Znhi4XZR53cRkiTnz0gMbXVRNrH35l8Ufja9wuZLNZYDxox6OJ9TlI7XmbPUQrczMjkuTn
PDm4RpZ9ofWKdrmCynPPFYoXioEqwl6SWaT9euX7YRPawd7eEWs0fITEpJp6WoArYMajlErS1Qvy
RwzikOIBQpw2vkSTWFp0/ooSkkcTIMmJkVudsQmsduZgrl728MlOalhJb6aOtXey6NexLkECpLE6
blKJ0Qo0lBk+Bsq/6Qw7T6pO6WfHtnZtrYjEPUZd6oPRCiCAO3TNG6yjuV+t9m6u/nB6+OgRAdkb
5/MIJpMzpcxyjR48iWjHeioQXKvUDriQQnMqDrhPYFdLsIJCiYtraUyhm6lfBUAxTB+aM1x7WGOG
HRgiDT3GKMxN2b+8d7oQynTZdE50ePg7pa51aQZrVGL/RO/0aqN8KvhOCJFHj9GSOaXo+fhCu5zl
1MvfPhmOvsr+aG4PGUjvFKnffjhF2h8yTv2P7o4BI37z3NOtpW4Eo56cYYwfaIvi8Cd3/DQSYkxu
lAcLzB2VjLwArTykB/BFctx/LvWUuyOlVzypA7nAkeqAZfT/GSR6qwqRQo7+81nRFAhofYiUQz5f
aTg1cKv44ZrnFfsw716bbCdd/Ch6CauRovqPW3RoZkP1luU81ClH7s5g0kPJHFy91tGxYnwpLVo0
0EuPI2w8qaMElGyKP48woyq8uZbMvD7ydIGsAp+39hZJJ9N1xaHz2WrGSh5/KataoyHIEXFjlSSJ
wIOxE3GNzd8/koynQo7BGrwY/8az7dIndOV3WxhbHBP70+vr51L41jVf/C6XA0XVjDlKuH8F6jM2
bjJI/qdKvJcaFEkjjTYcm1ZiLpbT64BgqICtqmeoT5Ch4FxD2xQO+ulSGhBm9wMF6P8Hna/pDO6n
LzHt5eYFlf6X2daNqDY/8WJ4DSUVN3Hxcg0CncDs+2Htfw3iLx2kSnUk5QkWQ10mhaTSEySL+Htx
MNokwvBTwLDGqLr1VEwKSNFbKhq1vfoVSKq48nxKIJz4vgN8IlZcGE1NC0Xf/OCkJn79VhmgTGPU
qbZj4tzQoYQQgL6QMoRLcAXiN/bY1Cfh8QZbmx8DAFuCFdLPbRZ9aURkhLS6wbaS3fKDlRjhYay4
rvS26EWila0rZt80lZ60sVLPaPqxgA4d0eVzjHtx9HkeDRAJmpDlHbyd0LNsHsMLUrgiUbo9dfnP
7N9Sk0YB1rvRz1OzEn0VmQ3FmtD/JyHqJqAB1jOHZ1SrBC1D2XjXdAiGiKmwxfVwH+kbGzQ1EOTH
Xvths9ahjIvI2M9VHI3dbMqMeRdwQaPRmgc4watw4fj/rrU0ocRTr4oxKON/DCEN6nYJso9cDWaK
PzZNHkjsAJMV5cWDhAjIn4HrK8gJSCWXJY9PtuNbZiFantjzR9YDANkPtyItGkWEAPnrVC8t2vow
fCX3rRO9igzT4jR7iMZt79hWK6jLU+zkP+SyWMx5WbgSI7zGSYUv9xAyRPWJinEv7G13P93Fmcsc
SG2wnIzS4foI4CiehdJESw0zIzyquTy8FUZ8Nr/C/fjCGU54x3yvUwCcRl2pMHWTzKX6RWGQE5zU
0TIugin9xTWLVG9ev8cxUXjmLfOwlihKTvnjXqt/S2GDeV+wA7msDoPqOQelEitJoLM8Or9xnXMW
UIRYjoPFaH3ypk3Q4StINxlXJjjUh1ApzaEpeCnUYUrlMK92VsxQ5ZztW3TQA6/RL1fEy0265PyA
wjk/TCNfFXfL5wBsunsmERnUade3VafyNSumznaSMabUoa8j/2tl+4x4xqgqK/qIxw/jaWxo6SCL
DrM7tKLhM35HReDY/WIy1hpYA0AMJVEzKJe+aqVRyyDTps1YCWN36a6DI5MMsl1KTgephuI5NVoy
lVWVNo8LtI+1x9UMK/m2NIcLDrzEAfUfAq3RAbv0ROvG1EqbcCByIpEn2izsUtMtITZdUllq1CYp
WWpyRu6dasnOsDLKrOWEVe1GPAI85dc/Vhb8R0gJ3A4EiIvT/fF8gkRUXhMEwaGAWUHmVhWN8pRD
hXoJP29YjfsLwEqpoVTLRSDsZRnkBBkT6uzYHKmEfXr5hq3FFE20r76iaMH3EFEpH5VdyDUZNrax
qWkapYflEMmqN9dmeoWzu4gYfyWCBxlB+mcpjUemG4aDmTXK88ZIzFlkyJeXVz0/MUxQpr2RRJPE
dYZX3VPQhYBUc+jQWt13534+/dI3KeT6Dy3vPmSHrANgsOhjiXAM7xLEyDCK2zIopg+zL8UykN/G
uifdjSCgfK44uRPpBrRC1KKFtjL6k/iMYgERUhvYC0+XGScD76/XWpU0a+j+B+qniGDPkY9Rs7/t
zB1Bft4dXPMXhlUwvXHUDOcSEwNI7cyWIN+7ZDqdS4tnD6LhNBIzoQ0aVs0h7Vh9U49bhSxYh89j
tn2BNndvAj7dI7quY4bjzykOHddIeFMK+UgSkB48BwIej94tXc3uRXFchhvRFFRs6aTuKwXvT+mF
k+SPAdS/biOzz2XpbHussNrE3U1JD/RLXBur8MG1Yjo7GXGgFvBcHycIefDwrxHAl1OOMAiW6ENx
kITpDGBGcP1Ha3NK5mIqXFdE9r2G9oNwtiPz7z9oLbqzqCWmARlr/Mr7aupJMiKkZ72Af+rtljoH
GGyRxm16jGQd9IF0KwojMp4rMdjYH03eNPVOl6rQkVsEOv7H6IKbkKNYxQ/pn8cVhUmyTsUUpKLa
Yk8C1q/CXmFNrzPiAfA/yQKD9lbK2a22CCc+oFo9CO9WAY9PMDY0Xq2X1eq8q/rV0DCz6hpPdQeK
8nQvE8ZSa7Ul1OY6oddEZTn18/3PNcFezZh+HfFOIYo06uBSEii5SbAg/AkvpOL84YX6tIBSMZ9E
Qu0CMhgzD6te1rTTLXuQCyN6k/hhU4VjHN+SfbaEduQNcc5mSJD6dUuwnrLLxokTH98ZfZQJ6zAH
yZVciYXji4ddNXT+Y4FpORLbC05f7aoMdkp030+uBUTbbgUCWwfvDGNDwXVd3ZmhqQC1ov+cgZ8q
ty+s837sS0MacaUhz0i1xmr0JbklYzGtpvvUic53YzjOLD6CKRzE5969enHwBX43knpJhcCYCjPq
frVBBHHpmZAAWFEYFXxWmOdjUvBEpp9aM+qyC0UWuPoNeFUXm9SW/iltLKM6RJQg0f9U41k7hIP0
NIZauMCIy58Qe242Gc7RMl2oeAa4Jg3GGAXhx1+411+otyGBkqNtB0w3ngFKAGailyRzWk8+SDul
l74xQpCzyPpYd9DCdxdIpTBl+v80XLCQGrnred3MF+ENJ469RboNwvyJSOPJ+nbCetLTDQ1kHKhq
yzlvnh5YsLd1tzAoT/ZLFtn+x0IQJFkP1xVLc7NztfQcgTdPrw20ixdwfkQjW7rfL+fDhU93REGB
AnxpC9OpZtbJsDTzwNXV4PrRnsyxBR6435v7bsxcV9eRJYzlPvMm8Okt3aEplWQdlCsDv/Mod4MQ
UVPsxXtQkwIJle0zymmbIEPMQD13ol6p2t8Nr45XYhh4MgSxZsx3KvkRpKkT8srl9CLYFgQTgNhe
UZX6L0dOdCkJfBp5qOg/OxrHrzTvZVJpA1Iw0hYKnGvwq1K1NupjasWTbXSrLqc7fZx9Z7UQmXbY
/o7KBu7Rgk+CxkftUmse/5PDySF7aMFKy9JBA2r0rdn+QLDbagF3OAV21/scUTV8NKujawLNncRG
hE7+vKEk3lZB3Xdbis+p6lTdMjOIJLMg45nNKSo+hL6w3qTERlDD5EhZOcZgyIUcw7tsqxWhKE4w
4esjc63wa5oSfArfhKmE9GiRHlyPNrAbtBGuzfF75Q4ccZn513kriMGVExhZDAyShPl5Ecnhnmgq
z1gZ8sVYuTNaiLNs1YZfxrmeBpj71GDZ7XcUBlBdZ6d7NZ+QU5M1nfUWW7J7sYi8PFDbGYoa2rEv
9OsM10Xb8LXqHLqNKLpdpQdNHJjWFscZPIHCEYlqIq/gdzhFLSbeJbvEWt5M/2OfjpVumc2zAHH8
GiuQX0wga8jVBgW+Caw2QQHAJrtXRMJ/Xvv96Lpze8F0zkE/T+E/saV26ArXqxx8YwQJ+tbsi9JH
nGjkbxQ4Dynwx1RnBvHvTt0CF+OnUCn22VwMyTrdQI8gRjGxLybyuFGTuROrnB8Cx0CZHr0gi9C/
SBpyqobEtIx0NN5UVMvpYujrd6zCat6jk/diHV9m1kw14I8MpZTTpJkUf30mG6O8LJEDV4RV8oD/
8NRHZTZSGm9cLzJSUg6y7Q3u+if0LjOsMHxhCBBMo57CxLrtaVpJHfT6gP2anMPvmLSeU2gvZvlQ
lFxLjFokQbXccML7xh1oKzL0xXKAoSgXU5g9l6D0XMndIwgXwHcTcE6aVyDMC2I36RYgBtnUWK00
wns5H76UzB2Rj3j2oyP1fSEyErZE9YEgMF2OwNmWiWfmfnBj6IivskJXyKjd9o40iDkFRkx/W5St
eaSTG9gnHCfT4yVaWK5JscffYWgKEOcU7CIgYlA9tUT4fRhEz0WniHoqPIge3hlMCLe2hL0O1X+b
Y51/ZALjvD/5gzjzQtDcP+rf0iIc9kHiSRwNbPchwTxb8cXHacJUhxjFR/NGKw7A5zAaWwLuwPXC
L/3b4jBOkxv1GJFRNCr4x2U8VMbub66oUv95j6xgj2qr+gFuu6M30HNgmq5US4fqka2OZ8BwEb99
moC8Lx0GJQHJv4TfaOzLR2IgfnQwRfpiDkISZJ4CsHqS/HrGqj65HUPeN8vVl8GeJ2xbAM8kiXjJ
2lsSfTRz6DceGIAnEpB2EJThBVs/l38lDfMVEhWgxmlGDC5xKYdkR1299gCVYRTazWSeerqtjY3z
bW4s2kukpxoJtHx9wU7LhlTsFBdIMxyiTB5b2Oh7mVvo4pZ8r4L4AQX8eQ3Vgzfqz/Wgrt8kxxH/
XB2s0htW2zTqdB/bmYwpF+i11kuhkCFiNGaUCvq/X4NBCDRbDyzEBpJnZ9nIyTLjDIJFtQaoCbFG
cMGkcAlrHR/st3Td4CfZnxSrnJDIP40q3OEvAP+LvPrcF+D1fL+JVxKIwB6X8Hifm7DV2vxp/YPq
ffkyIy/D3RWQXnJNeVuMcbuAUgpq1/XbBTgsTm+2oor2N2R03xl1Q7cL5sJS8HCvp9Y2+riVpFWZ
uqsxLX9oqPnHsNkyA0TK7m/dGbvYqd9brE8d3heM5XXANJlbLBThxe8233jiECGVIEVH+G49/73T
T+xH55b170gfaN00KLA/ChmUNVEJHrzTU3MWlUV4hFzS5yMeR0rkojU7M+d7EXZqaf7LZV5cPAIW
9JIYMPIs0j0ahKUcd1iXuLg0vSOk8wrqP4/kuoCP7WZ3OfsPhvkGm71meBhckApd7s8xLRkhBIwB
vrZfcd4BfHWoOrncjz6GskDaSeZOkQ39SzdEN1zi3vNkuHXm+SvVa2Kl80fL3kzXOCRBcXGtRaIi
ecDHSdIGv78nYMu7nSYWJEZXsZNJti9xyLNwoqi2WKjnkVo5SeWCBml4VlnZR5kRLPdXhK9bY2Lx
kVKxUq4Y3Lnp/OKVJdtZASQ9/5GHnZ6uNzW2v6q71DePeaqISU0pHVLc6g3TOumG5C/GRg1KrCOq
IcUwgkIOxbdIBv7bThVzzKSmF95bm6GsMM1peUnmutEe7PsZ4H6qhL194U7BgZ4KwsuonFE13hIN
aTX82JNxAn6w/Kf72LX1XqWOBNVC4yy0Xf+4YritQ06p1jhKO90JTjOjoooqJKdYFJ4JWzFLSLw7
HGfoQDoT4OkO061cPwn+yLiv5NSv38eIokPevZePkT/Y4W4VACjlFhMyB1YQFtAUtgRczByFCZBE
5nVzc5hNfR8DYjDsQXeJ0ak186JCRS1qP5SvK830zHK26dukyI5/tpHrSYBjh8fb4Ps37U43bbdW
4WaqthvWHgWw7ZfccrXWSu3lr70b0IEKUxhCS45cRRp9IssuGPO53kSZ5BJad53fV1Uz05Nut3qa
xZJlSyMQOEFgfyLqR5Y29uIZ/AR9XpQfxbGjnbB1VC8W11luLz+5RrgpUn9Fbd59EZa0xK7CPIEc
BrtXXlKCKqrcoj9e6Vq8hoxrTaY6CnNO6SuPB+xHoTh9r5H3vzfeVyfV9BnrR5HHEtMuEFUJ+HW9
HPYhyo6mPAyw//1Em5N9P3oJoYJEfdQj6UkfAGtjQ0+yzu9QNpLzCOVqln1FiwEjaJz8RcNuoopq
W3gkb3b5UBkYoRi4gg8T8sSW59mVHqeASTUVmgJ/tdtge71yxrMORwqU3meoGiKktAndteJk760j
Ig8tiruwytJnMzkaOWwYqv6hS63TALl9Joj9D31dD9htraEFhqgawcGd9fFRmzU5P7c6fNLrSQ7I
0fqO/eWDEsfHO+WtWfqSD1WDzWkgm30kaehwBJOKv2DB79asSy+YFPzMQZcClW1X1c/8KVx8kSTc
5Yuqe77Z0aqoKYHkEdxtlvNdH1CnQ7Po8iQg+hFDaOOChLKjYiRZofczWTAmI1H8TbiGGUPqc9OY
AVmPS+SeUeK0MECaNXR/1a8Y0N6RVkCCwo1iM09cnGL0OA7mHWZenMnEPEHxidCKDyUBl6ylDvj0
YujsuWrHu/ZmaUnRCRV8ZdASI5haQcA6km6+Uyq8tlf0BRS3Rvc67oSP2ut1r/go+FfyqBueQ5PI
m8AjkAIr5+5kWPgUgrnR8O98lhJOZbt+s/oY9Qom51w0oR6FdW/JDxSGJKwRXFmWOJ2D/mzu7pZJ
hHw9i58YXvpftKrQB3y4OvObrar5afMhN02pDm1unrXbpw/cJBo4oFymoCeM59kCiB/XfoI6PsgI
l7Cozst+nsBV8K4Wt43LY/sHSyCO8pIefysR8er2g4b/Uit2pSC7rasIr1LSqvCf9FIpBKirRvOf
ikrlvRb6Pxk6xmBg01XodFov87JF+2jsOFK/g+WtckwMnLrb647C3kdy+PbDejmyrzRw3iPqJS33
T4KNryVizIdnGn6dJse5ovJEWvtF2wx7EjO1Q+u8Hz4ikzLO4M46SE/Th0jPmV+in83qe5puBmb5
MA1U+R9YX9CLYYDYpmQUhH0ptyHXK5E1uOk8LEvf7Je+r7y9XpD5V4wsBu+6J5ZXDGUfLofH5QDg
J5SfAU4657mlXqlK+xZlDuAFjo4kpPV62QcZMs7b5rNr8Mc5p/CgrYXbe51vZU5b9buFxRYL8xdl
/3D0ZSSkakVOEonxa+migs6orhEuog/S1IJaxyNQpC1BnkXY134fuGbOU8AmprdXZ1Y31z8/POjn
RBKHWc5bBe4A6LPk5R3bjIAhEw72g3HWvba20TVu2UpkdGqO527qLTlw05sniyjIwLrmLMzaOErC
mFrDnZ3iqRJuIPso5yT+f5mnf6SysxYvVpOoX/jJ4DDtTT5T/jHX43tbf+tmAyaHULLbdG4XUxo2
w7AqiK4ggsmgRmroGmU/ae+4gTvKlymaiuCrHpRPVi1AdIV/qb0EpBkC9s8L20Oj0ietH+YfNew6
aTbWwalF07qrXgzG3aR59GA1m47jTs2XqprX2amavHVKXGeFUOe6ax1UA99GeEhIhlBulEfzPj9F
ixel4mv+Gf1ArxYhYIOkUAAX4ZhI5BOV6J41ytYQEEDimB3MHz+8TVHDhDSAxP/thi61igsSf7d6
cMSvdxzt1sUDT4rCVZG572n0hOz2hfEHXRz5UjP3KI1C4isJHhNhCu3kIU4Bz/9VLfJJtWB0lfJ0
svUdq823H7GQqmxdtZpaJ1v/y3xpgTLRGvWV+sMhtevtps9O1+hVGZf95V6HN/QYr2hsIVlkPaCn
hcEedo4TaYYNdAE9GzUig64VwdQo/w1PIwH5TFAwf9wlgiIGT/cYDYjDkCi489OUT47F+7+nlwJX
O+YCCdj0dvXa7pWwJuoP21Z9DnGG+GfdbIHTaHwHGGamZPY8102GihlxWWIXjoPAXKcD98aS/BYe
owLtG9ONeYqwGFFKyQYZUMbGi3r3pnWu8DInzXXjl5JUhyctJyWBAVhj+1+l5o71VD2CiKTXkiFI
AHUt+PtpevXgk4G0EOzVxuyE1Hu1uCBIx0uect+DmH/p1ubpodLz8n7foNcHKDap3yAoqzv0VlTd
iuU1jjcmYIwTDFG80eSvZRHJK+OfvXpwuOkeS6QGVCmkmGMtsEkJVQvELZZaD/8t1Aa1qMLP6gIJ
66ysuRuy9u6Z4bYS8Ku9oPy+OMpDZn/AQg6oQQJiIduWN0se3L22xKHhZ8TBkCiXlBzwmxH1C9Fo
qYo2+ATR46HdumaeFhfockavEaSPL20a1PiqVBwfrzyr5JARw42XFqMn3mpZv7freQ8X95CR0rOf
wPEbtBGoxS+Xb3JgPfh0agM0v47voaKZDgy6jmZau0GjuQX/LKhzEgcgBYnRIzCkPcWgY1+CPt2C
hwxfOW8wWu3kAr9iV9oxEtYJsa9rAJmD0RtcI0FhZYDrVAOLHw4GjtjaQ+uYZdC0jMM13GIoseyq
iLcJXc3m7iraXZ6i17PQ9gqCPVi51BLpjGjiwpf3kAy/AA1QguX6jDw6xEzgCPMWLs0F5IbeKuYB
1mQEH9qVSB14xA4tMS+/Z9CDNyktMKWTaBQ3P65ez9cb+Ks3uqjSRxOmE4F+gd7jjHrOsaYPJc1/
UvPvPmkpy8z1a6R1voq/cuokl5dGBj3a1DIwL2TfgGXwMqz+Wq8qTkfBqiYisl4JftPQ/DJ66U/S
sbrKXsbLdRrQAuECtx33lvucQx1rZMRHXOqTqXpgzETp1QOUGTpeGOA+8SGoUq5UAWZGICXCZUL0
HRaG7GM2AOpvKnxKI3OkQoFLYWjnppDSssrusmBSg6q5XIxFrkhR87c8Mt/OJX+X4/SP5xGdF4Ex
duGbULL+Yr6Y1wkQXbZHaXcPYkAGKpn2MgFBe5R8/bshncOoOIAFEtMRGfhyCRMqycVKAGrQV4CP
dGyMFCcmuq2jnDp6YDM5BiSsHDMD/LR8MXvoH8bm02LpVwe3uVJP+CbSeaFjHiklZpR/MYaEs01P
0PE54loGKiI6fx0H3c6ruf7YjMLsXhfZzGQ6JsPcA0sH7KSbYLxO0wfA0Yju2aSENLmlzH9jnIRC
BTakVERO6hIjjbJsw27xm3LA74nyfOevdG8GHDC8JOEi5TIf02Rb6TtpscJiQHT5ey3+4VSIyDQW
GhIJ8mJqeM1DR7iyLU62wLi9c0TlOs8zoRUTxsDyXQhSCUerAkYty6NnhV/jE9GmxDh4Wr0AEkEZ
xDEyMhsVNS1IQyEe2lrgqvzaf7Mww1eR0DqZC/HE/BOaumGkm8TLDo5nNca/UmECYpMA05YI+C4W
3d/f7yESd1ILC7+kCcRn2JjUV9hzY5xda906DdDgZeGKGuZ1aUl1/rGXictAlSall/Og2+V52qNd
vZi66QYLPTt28WaaNsVwCZwpnR9Cle/n/lJ0bH5alyynKbdbk57BuXAHKv7xUQtf1MDhdkYG8b9T
Q/RyY+F6T3cc67qw+dSD7h7Bacfx/F/WBByDlYgx8FAJGb8NfRY40KS9YVGGVHDWuUZTpt4Qoh/l
ZD5UpRqko97ULe7jkWDrlliozuR1y+IIlyPkemAnu1/YZ8R1GObq0I1Cz5l3ZtdSJcmA+CJv1hkH
758EpyM6I5zVV2USXTk7h1/l6fHG9bZnG+5KjR2CunDNmRFnJG56dCASK4XkarOARpIeY2hjPBdp
2SM7tkleFpw9I4KHl2duvMVuwVwwLNv+iPD77mJRKIyOGKdCYLf3W2Gle9CDCNABY5dmbvS9Ci+7
JCV49REcdcVLEWZfhisP2gm23v+vZKWDy7QPuz4MjJNcNDhmxu96lmMSHd9n4hU2xKMBqRihCnXA
zYfaKR/9lrURh/PVuojK3ngz2nXVTAuNg2vKODBrYYpCetqytyiZtGhxPMQGcM9gjb2WQ+OEZ5pT
fJNp3VBy41xAMmYU6L7lqX9MJK4lRR2hzFpAs9QGX8ZheDSYhBhX4keJPTXsNgBE16IviGwWzTUp
8OYRmYrFX4dR1otQ3kZdSRNt/EkTtU+f++ePpf21bIjcbFUCFrjxZ7Kw2DqWF30yXAmuT7RAzja1
MyhP594MI+RkuTpZzfPTV62v4f5dSmne0IYzOq49LT/zT/mIphfxmfT1jk7kDPET7CkwexzfV9Jp
kQj4s6znMWFU8WcMMWZLSEP2rJ2ClTOpzbwPoea+2vARzIwOeVrB8JufyicPy19iB13fbqrNXSDS
btpMsFkefTdxKA1eVurlr6VNoAD0Co5vYHs+ebv7iV3h2YXc5CNLGLG3to0uXQp/1bkvKpN94eEK
fNitVkfER26RCLKQTlqTRZomyNb7ReRbRgn79cWTAkRva7cLpE9fXOta1Ot/D4YINFe5ikk85AVl
m2v9KO2Vq9qpi/nxMOMpoo9Y+EX5UjGg/By/AjX6792JlY+4aAdqyG70+9wtUdxR/U5p/QNo4AEW
d0xvOINPbiqAI6qM02Jt45NsEQBU9D7wzx89fEz71NeoOTCIMSQOpR+D4QxZ7ZmBlbdfteTNLb5l
UibfJMw5Hq2Bq3jN8auwFPE1GnOIAihZeblS1wASCzQiQ6kSP6pQ5bmRvXH23uS5OYtiiA2a+w+z
7skBdWi8PPC+npc6NFQpWgK4vaGGqKdTuqBP+78gv/vhp0rFerfE0E7jpi5EDKehWnB2cVB1wuDp
FvTEfebUwQUTlCLq9tbC98N7uwtMAR3wrQBhdkm6eTi/amqFVuO4pPEUTQJQOHJDl0Bo/yGoSayC
Qo2LruGhP7Cu4lxVAWe5tiKUgOEkLjtrADZPAOUrERtfy/xQ4kpvjNMRqbvnPuRqrthi5wFQQFdv
BL0pz/tdhwfVHUpRp+8MW8O6HOMEacgEXR4/6497cdUW1cpoVA1u91ONLitKIf8+kMrWqsXvnyGz
pw/VUy2FFcnt7sOIZHg61LDKO3S0Gt6r4Msg9eUxjra2A35TRDGtEFMc4nagJk7X+Y6Y25nYFqld
CRzA8Kjz9WMqxoh9FQMzJaUQtnrzrIaAECUAu8to2CjoAyUb95K/tptuem10l3pclLlEP33Dddc8
cT3aC6m6XzFiGqAh3my4jCwwTnQZmLFHcmbNyXeGPN71CqmvK4ORRHH2EBx7AN8A9AQ9qOkwMNZ4
g2dDXtyhwZK8qyxE3Caz5M/v6A5R2sxp5m4mxeACWSm967cOa8fDSBVfNGucDOPrM0UC6yFSnUxV
CfDZQKmGoRy4iBI2kRKjau7HWGdbdHF7vVup1BfDWyaAy20SE/G5eFQr7UbfJzfVBWSZcgpqfGaY
0hRtfqRas3Cg0PANPuvOaxV5t0Op6yl2IJk1jKR9YUyXIhOEnuLRZM1C2TYcevgj6QRrV0IBH+dY
vNP6V7mhSzlzDWRBqiJ6bbAnqsdLheMNoON3YQGITSOONWYJ9bqXUTi+vinIOI5clEwZBSH2hIwo
58OOb09JzIPow61AOXytlQx+tjrYjQ43rXvCK7iHqYJop+aD8V5urqffQrWhRM99ZMGYkuRPiDTa
/Dt0YBa8TeiWHxYxrE8zskERR72OmLTpkSQmXj1PlVyC9gXouTqWWtDkW0x6wIJTYQ86ST2kq+Um
8PLgPYjhxYXi7oWoN0ZjhtZs7Mfek2i/zrpG+WUO7wLilAAYjOVAVhlXa8emyOAWYxn2AQl4nftN
3t7wmAzHPQ02R09WWzAUGT9aydLCBBY+6QyMJbHeipH1/dJEud9I6Wl2yEF4n7cRtW2qNYrjqYLf
WrpyHHyNXPkIS+kr68RAmjenmaXubRkiUtzh3B8H67pDuJaYzmys72SUKRX84JMttoTvyITNjLFX
Q7Jj2zDPIdcbXktI8CXAowJcE2qnIDQJTCOTQhvBLyyFxSI72qJXTQQ7qpCui10AR1J1Oovq6gd7
bxIzX/SwpMtMzxTY3YTb/Gz7AonKvPHhM3sfh3YL2AX0VCjnQQMApYkLn91p6dTjt+LbaC+NmZDh
3Yp31NvV65uaRS3E6sorBRUuRnZjTpEg+DILXyggwSPiKVDyQUtYoOFO6qO2nBbGxGZhMQuqwxNe
X5d+FeSpl9m54PZeENK1mZr1rK0giWIWYpRkywmw7bBMrDXO8Ck9Qpo9VL5b/oyE71MqCOx/CCo6
YFv+yhYUJMaJMm2BrsjFbIBP6bkdeWh+CohywbSiGh0BFRMxxdXQVVAg41XALkKXTFLYX6aaJP8k
I6sv43VXXXaHJSYhAMVMFSZ+aHzcvMGasajs9ONKIAFkd48H7KGyk39PcckEsiOIqa/9BijNJFm4
ePqrWsnVHPai5ehseekIz+j1qwSsrgeKBm61GadUIfKctme55gkkvw9vK+BvQGGSJLC7tOyzS8NE
3m/cR+9/TRahUBA3dQCRgIcLQfuIgZCROjyAlU+hTOfez958BxJfov7jmElRRKJBmtcQrooFuswa
XeYXnwxFmD6qCdrue1ilrtsTvwnAbayUYAIsFQGioYPFXi765GshUApI9EAq5Sg2bHv9ibW8vj4s
VTHYwa8N9h7WNNebDR7v9tJ8Gor4JUEmRQ2aluYgWp6/xvmXBeYV++1hhv27UEPkGGOECze9kdHp
mQTW2Ua/2Bk3Pl+eVEHEwxI0leSZZKnkaVSWt/4D3B2nW9GBb+2Pm9LA16W2ojWz69xkgMoyLk9f
63tnOkCRv7rKl16C9Wndm5ddn2Tc9Tm+hdlihVX7QlwRg+zWet8Ffbidd5sCbvZDA3aswiSq5sDS
TjNRZjDnVnQRFYmJBr6NiP3ZCsSacf+I2sb6m8IHvR8A1VP65S0tQgZ0XLUcUJ+/H+AJhCusXotn
JQU3We7PrVdEWy+XDR2/bFpLtrqVQUtnKoZwbac1Tn2o8/KQ/fvH1P88FvQcHw+oZnffGUgGGXDT
740sZavQqYG5sK7dPuvKX5Nitqx0VluqVxVildnA9/cDQGaq3MdzjFvMwA/JW+pDsoXYWgUpy4BR
7moFOdYkv+FHSitZV/G6Srcf41T2xDo9ZCCNOE581GJM2+jEE8EbrNSQSSXrNkNZj9HIge5/aDvz
1SDgSr+yPQXGOqE+rdaw5mwMPmqqaeTMv2bFYJZJQurialrq6OLh4E2anjDx99HyQyUMvjyl/jJH
zj+VE3ou7rhWYk+rZcIjmfaLKUXmLYEQ/wAEy67J2xSphD1pmojPJMQM/1WRJMyeMDqLw7fVL7BL
X80Pgnrad76bghRm2gELBMSXl6naVFCUcOWwDYtZ/LlS//Le3f60mPfWoMBS8AcHG8ByNww8pLyg
9XM7lfnSt3J67dS9b69Lmq6uiXuEnjNWSmBEYcyivtWy6RaTaaYAozLN3oDlDM6DBC4at8Qcf/B0
QAtf/BDDnrp4WQgakPSegH4rqfp1QpR2SoTJg1ANUd9NUYil+uZUbDjgesoUMJ7PZ3XFMMnXdp4K
WQAK1CDjR2SPapiIt7zu/biKy+Er2k/7gtS+WxbocZu21XWq3lddrzum+zLBS0bsuPvxpp2ofv/s
qAsmt70ZnXK2sou3Ftw5Tiv1U6FZLXQSrufpTohp9pAYlXBdjvrRbyTKVwCS2xWeXl6oFNTZIeMy
oSD0Uo6SkiFjb6grbiT399r+9vD8G+eiqIal+k2v3vlHd+AmdRfpCjQ1cD6xq3f6lDLyukBLxK0I
9pxore7YuBg6fClYPWF3BVPR2YQDtj4cXYj4O0RisDUFNYjk2ATsSeMgVckot2OY6+5wnQhOP8k+
r7TL/8uqlJMAo1L/MbQZfIN9a3AnWidXOglQAAVioA04wOPp/9DpaQWQQllhSkbOjhDXiqav5ifE
zYGQBsQaUXYHMOboEeEHZfzeR9ydnFMv900nDUwJGRoOGchbh55cMKCJOBON2i2NX63AhUY12eYL
nug0MROowrQyrzb0uiCm5GpeuUwjPAcfBpUg0NQoaTwA7U4dP0H2bSOq9v/s5iqVmvmd8X8styXa
Ve/n0B9gMm2ihvBeCY276vIJWk9WvWbRCuH6Ia44/shZa1rM/7Ajp6e45vSkxMHDnTEE6rMtvzzL
C/zOJ0ewgBrzZE52NKudJhtAsPslsQbCRoc0/R3ZPRhlj0+pBIH+je8m00LRgEL5Gos6tUjlTY4L
nbD3wmhW/Ha6AQ0x4g7GMLBNErE5aM7P8nzXpBLvIq/1RE61sTHywE22WY3xSqPZ370xNr4vEr1w
HxAn1koTVfksF+v/0y7gd5VC1Nq+pfuuLhyt7wFYlrAHZ49TnMDX/faaPYl4BkXeE25kYjX2GI1s
nhVww1QTIhdIfXQRR6MI2Ho+eVb0NF8Tt4tOkJg2puNAGcRw8WxZaYJS4mK3wUXeDkTgHJIYXZtQ
ip4HXfDAYLJDat26++hmpGmzzl+43XZET01HGEVswDPyWD8mE75kolAOv/z8TksRP0AbP5eHio8d
oIHNjhwUbdeGVZeJMQaaPgQAeCCpsTcKZQaI0PTEboQo3PPHzue/e2W1iMafDfKthcb20Q8Rd7xS
ECvesvzARrRDxcnb6MRvEW25gbAzIn2tPqbisyfS3PffjRDvWUlmU6dXU/kFDFk8iOua12SKSRZM
1Q4TOXUs5n1oaoZzNc3Yh8ZqLgNATyqLHUBs8NtWvyKEq5/qjfnLvh8YLqF7FZAXEikOGDTCu6EW
cV/cEWYWuEbEsgWN7a2R1auii+NOvgjyPc+xXFfpgEF+ngFtd8/NVqFBzSwVr8IR9EVc5gyeyiyd
/GmrLq19Il9Rb0HwBkxQx3z6q3p50CesJ5XWSZ9SusjfooLnUL+9wPro/KZ8kWu4B9B6TocMSGdm
5tBFUXT2zOUI3ieMXsKDt0tkeTMGPWKh4osl3R9FSgnRqKCuMAFw7uxz5i7kxlqy38bZlF+Jo7tA
hX/XoayTYo84R3iq55Xj6NcSPizQrp1K/HusndxkdyLYO54rXdAYK0KEsG57oCQr5rkegoJl/OTc
IEQDuhrmlC9IYNmRQkuAH+oBfEMlJFaWwlVvGr4v7na+JVAZ9SLtpn9CXYAZZdkBqxNwmua9OAvl
smntVWZXt3W3QFI9n6++0UmK+uflayn5268a99stAGP7ihjrXj/lE+pLTRp2E3WvthB/vgjIsRQR
VCvh6PvsinUc2IsvFlz3ujrVyVHK7deddRubnC1Zni9YQ07Jyyqs5vbCW5qf0LWzI3mH7iINOsts
AnncfA09as4FuomSSUpCSJ9yfkQsZr0mVueo6SGkqmQOcYLGpKTgGflpmeNEN8whlp54f8HI4mcC
+h4XowWQuA7xD5mjY6PphQ0T3KC8SoVDL+cL5uFVfy6SFgojBIXoqezQQfBKN4jmB/iB2HRj3WLM
kFiWpx7KKWAJznUo+zgLVcMDhpPJloBgOWb0D/yM2CWsOzL/FAHcSKu7pHagXa3fr2JmfAtCLtNE
MB4t4l/A0LCeZduX5dKhVqw+v10UZ2bQdx9971xDlJcLWvBEUdYNSpt87ivoQCbDvP4AzmlcEA4g
YPy8dTTOmHCXA8aMTXEzddY+2xGOg1MJdNttAV8jOcZXre9fSmMHRAjjWc/rNp+7iJz3LX6UHRvs
f4BEJjHlhL7KjiXJiAUFl9rXzZtwlNjVlQfV+q1NlOneqzhbmkmGS/gECto5pFX6J2nt6y+MWAXF
o3zlPzs2bjegjoRFo5yR2IzZ7Ne2YgYXd+omFwRMN5vu2wDBOS7DUzzObCcuypuqWpaWNe9fxTx9
3VZ2yMrnfKQ9B6UooLrzyGCsO5EFn4Kv/yaPpqA3+aBPN7TsiqldMQX/tKM72+p4u9/X6CeHJ3dt
ZxwGLT1H/2BfHsv5q7InucLg+NcuLNtfNbuwCd5bQmHQBMesu4L+q17RQF7t7YhpBfooTk4T7oaB
dLrBM+C45K5qnVLulTdL9IHbVKY5xFlbfd94bFhdLvd7tWY8JzSsJh314lztTEdnplHucvanY1y6
oQgvRrxtjX6ykmqhL++pr9YMGcmMH5K4f/bRbAIDDNjV0zap/Vssh9pN7DjHy6kbJHnYQhBxw1J+
pf59znQZidH/wzRUialtRLnoPAK5xVUxCY6QrpzNe+fZexcNVpRcQZGg77V5aaeaT29Bv6Flxds2
kcKpzAQJOFkQobC3Q56wzkxUaoh5tFUCUFX8I4tQsO+x2sOLFLFicfIWVvmvsOk7lQsw2QZLm1rt
csT+NVkgkfAFscDeUKlOAbS7uJGC11wLfUn2osUO5HuhiW6VkzdCQrgdle9v3FwzLEKrMSDpmMh2
mRJgkTgL13X7lWVV/rfH99HWMhvcQwr2AGdWg+YZ4+2chnYNa8OCYzCcsIdguGmzF4TxVOn5s7qz
bYZEcWsImkYKQnEu+0GBVLTZLK3dMvSWrJSCDjabyKNoub2qUtR7+SOw6sbqGXwlwpHld6MfnMYS
UGEu47bMfNpmpwtRa+l3Jd/rME3KSjdxIhFGvnk4Mf4bBKHmryMyiCui8FYNlzWg0EhQzVhBOYOC
whUKkblmv99/Nho7xmFvBtEW4A3uXn1PtJY8PSNx4aY6eTrqakETBLAzRZ5Tkk/jBh7H93COemrE
8XUut5iuZ2oU/nna+nHeEk3hJ4UbVxQB1C8vtWlJcedsCkPLLwYw5NjdcYS5BrbWluq42vwwjuWr
5FnoVAWrbongsWI4YyZ3bUpxLaFex/FFRQe7CcuF69s+SUlgGPMMmAEO2cG2yaWbAzA120TejxnF
4r4DVjJAd+B+CI9UFQEscWDGM9j6NAcYjnl3g6YpTtMX9KwPawOLz0sqXr/MCHEHeymtXeCQAYtu
49O4bXGcald0XJHRRYV065GcjvrokLC7rx9CLQh6SP61349BTG4GQfR9zWpsgKTWeFLjhjrV5wMD
rzNvVrZ7tI+STA1VPtU1iviclaaEX/b0kJWAaGg0q0KWvfXx48OUsltJxO5kLqQDh27XzDh+/jGe
FZRceMQa4Ni6U1hl8ERHDB0W9Cdqeg5X+zmBFLV1mAvVXKcBM+6GZzjgvASRdOxCLvSNQYAxkTb6
y68/eyE2Mq4L0R4hLyRaBh/U+svoG9C8EtWCY45uv+shtNxBCfDgDHtw8KcbfH0cHHe2efYg3e4o
Rgjj62WRoBHoDSTK6ni41ux16C6sNiPp/GvsPuUqzc43x7r7+ZFwCQpOmyl19i1rhxrm8Ny+qH6P
mWFR0pwadmTMBGfhTGFZxaOK6TitBrrcrjc3T6pSBeOz9GPXoT+NS+ugW1NxmJ7MERVkvO5FUezz
r350d8INpoDv+QI2LruygBL/s3XXFJHwfK1k/oS/m3W+OysSfjm211t5D+UrIExPFxjT4d3pfdh3
i6ureLIMlYV19r+q1DCQMZgCf2qbtiikPJc3zg3/xDlPTrYPUvPBUOoDUjDqQKrLCJeDjc/KNb/N
8Dg9xgcctc4K50KnrdiGMXq6LN/z+k2stc4/TXudf5OEdSPY+t8wfhw6lmH5R4FET+RWbRdgldqF
xg2z7dFs9CVUXoT0gXMG6TkAPB8iOScK9oCB3+ENYmXWKeV5wXYtS38iBrq1nR80LAbVerQOonlA
Cdd4piGMHgLDw4aAMAx40LTJZmvu7SrFdB1vR041z1HAKYKo4ZmpbNfhhh/U7i3gnhdW9DeewFrd
qRAN/5gj5ZQCl83TlWldTbQO504pbxGGvGIO6UOlnF1wNnFxA4hchp4Sd9PVwnnCsctLrztyUXrU
+3r3+FvQ1OIjb6Hlg7s3mWL3453nSzxIXdVQP6XG4jeiqbntUGjyCQC537V7aTqIrRXyUcp+BrBU
dJpE0A1Pq4qg9Ju1wMDfHg1ywbFspHhtCybEJy6NQ1yz0WbjA7VhtXlbJFPiO4HwYKjUvXWuMb4P
Q6Yf5sWZe2UX6e001nZRFgSrIVh7LUVfbpdItsNg4dJZ9u3s44q5JIKiTuW6ztbDNKpg2BLqJ5Sn
x0LMdtIfbJ1iRWDXSPaLiOitGnV64CNyqWGpA2B++Lel0OBJORreiXyA20um/4ouV3U1b9AazMpm
Qi+1y/BWRhu7on5+ogtg2IvfmrgZ6XtasUd/Kf4dgx+qb07zVJRmaH2KYWsjMuAg30Qco4dT+iBe
aHmvGiEy+Nc9XpUFWgH90JcD2fgoPKApwlpRGHLCPRCD5rsJqkTOM9bwHnzJoPi5JeFkogIuAj1c
6yH2L528oUDqQgGbh87fsRhyHSHcHxs2SzbIjHS7If+p44khNN7Ja86ddwNNIx3tvR5OBmCWbNQy
a5fr6RWSpXhSeqdWwbt/oMSViZIdo6qOmf1eTXI01ga7c8JIJksEW1xKN1OKMVFPr8tU/v8ne6Ex
pR1CZ+JhJcIqesMuz1Xh3mJ2hUPRCb8YEsH9NBxZU9UT+tEVdLEyn1kj4QE7ApZJ6XFdL0h8RnzC
MCUmeVmmjHKvY8nmmuTMs4HGJRE9sSqBQAiESXSKEIoN0Qfe44rpCzqKvoiWcalODxcyUev1IM6/
YcloI6uC6aW8hi1qiMqFR5Nzz8/3rPrj608ZXRTEKAAxzh6Xsd/xxdUenRJRpPj0o3+m3Pz8ax+u
/2jnj+AuS0EFf648VzKBFmXd4L15+GFQUxWesKcYlds+gZQ8HbhJS/wfraDRNrCEZVtoBdOEByhA
lsqsDDGWDkajM2dR8s35pbVfG7y2znk5qmyBms3dAzDZeixpCtoxcQBFqDjsXaK6on91VzuNW7PQ
XssobeGfDK6WfPkCS10SdSJPSOBCh9r/j11Ui67P+M1Jk7GsiD4V1AF6CWdwHX7JtbnTvLXYLIJj
9Ukm8WFKaY2Lc8AsK6zIUzhzNJtWGIIbAfN9huN/KTrXoU0nEG/8z6X5DAzfIu/KFJjnLYYCIPdL
19FBKPkJdRAZ1O1aua3AJPutzJ2dnpsojBzfmk5Zx5Fdd9PPGTYEL3l32DFd0xWEJJK2/tZx49Fs
qydkuRZeIIHSZKBarqc5OVr8vVmT9ydT/ly3HWX69qT73vfWoX1dLpXPGy5s0kkB3cJeuVrZM0JD
GrbwdQ/n00Ehymah3moxxMBD2GOSaObHtZh1ByujBQ3socYTAs3L54hlYcvFYNm6G+JidZzs+WE1
I0F1KZJPq8esjtC6s4GCGPBWiOqYAG1q7y5xvly8NV1zjB47qVu1LXJeKZDUnZsSgat+0cfUXgvE
1t7walk06Jpc+lSpLutDj6bQoirAInasy1ERb7Bg27mevV1yxs+OikS0AX58hFkxVCA2qZu6S2Bb
GwlgvaB0DK1Viohtn4oHWSMjenRShNfVobiqeSP7VMauilfbO+pF6IZuSQrlYEh2Mh8+sJBA8PV9
/eBMC0mv+DNqzwSJ0jijVT8k3mJBPdKDTNwACnMnhDm/sllHebnkbYlzSpzJR9Ptu5DfixGdGAGv
KDozCfgmEXvOhN1zyAcjmW5L3oF8LvpX/OY0eaDrLzvQ/YvKd9IKp8vYh881d+uA4V9rZXZUyCY+
Hq1uKkgxfidkv9L5JA653eCjI+apkvAvzEyTDCpOjzmW5NqkB9c+kyU9Iwjqkf95mHUvkJKp/iPM
8NRWf4Iw1egrVvA0GU4+zMnogNArrfIrJpVQ7jpqjyAldAW2rRREvcbYH8XLHx5h40FciB8m5v9F
qcN0mMAlxYFNeMIsLrlhXS8DPo3JfKsqiWjuqVgEbfSkQpBUVQLmEmmmSF7GfkQuevkW6KPZpQnS
Mt2+KL8GKijaKXaYLUbUaVG3ia/0KPGYLZSguqj/r9VMT/RjFo9dFTzQanQ6brd8ya1Y1U2t0F/Z
n3byo2M756St/KZptAAuDObTrS+L2ZLBiYPr4bkl4TJW/7it3TL1GgTCy9adq9QzONRc96HJdOMM
SFeIdsP2ghR+HCdzWNClfPidJiJooFkNvk4a5IJT4yvMkGXi/Ao/4C8JxcGqRgr/P58Neqx4HS+t
XLCkIkxvuhRkQCEg1xOtmnLqkO9vXD6BwPGM6JqvMHfTc+1oj+WcsijhTAi0feDWHvVIiVo3WDsi
rQ3Em5uk4ErLADf4SpLu9r3ZtvKE89FO+Ackuc192HxERucC2XB1mpJZhyKGc8YxxYnuRNCoEEpq
FoIbgkPwcYIZxxQv6tJZFQ5CHbqEic5UB29bGEbu+Dit2jRAM1lB0CdToAv0hq4ZlFebOyu6siAa
TC4g7W0Iuanp08M458YY5WWUsPpUEByHhEniiRzn8YfA3TkRCd8S7ix9lNG1OikAhVhYx0dKkiGw
q/8No9C1ToAlQGYc32ufdSBG7VLDrHWQCswTE4uuWZGV93dB9J9eqBx/pn8W4rS/WW0KmnjhTMBG
ZweERxV6yccRokDmGTKlAZqPMKsWzoOXPmz5j8+Kt1bpjE23i7iNABdgzsW5C2SogF9tynamen2G
QYkTKoP0nNZZWvLc3H83P95Lp+skRsvYqIgrQVORrlIgTMWHWoZgztN+DURrhJVFR2b7H4V3LaZB
Zh2ircoZCqPAufmt4CggyqzP17lwU/+KE5b6UVD6z2JO6tnjsx2LZKZwjYx1/8zE6gzchvYeFyHq
OsRF/7sykV8+gmBpE1+83W4A9PTOAzx8uF9B13FMc5C4vS3PwfDFbZHn0bA/u/pUrKYCeqjWEsqG
yiHNeo9KQxJI3260J6qMfOEcLpdL1Hzr/OmFKAFLvyXCvJuh4SfrdXe/yN+YFDFVQwFvzJRW6d3S
ClytqeuXAr6FtgH5vCF9u5uvzRzoiz7cBfGMxeUXRXKVGyXroJzE//wHCcVr1FD8Io1+epWAzPpz
JjdxYRfZNrOtxCPINoeJ1+DYH370Jg6K0o+N1rjRQ2o0FRZbm3fV0ag+tzsyn9rFI2z3ZndwRzBU
0CUz4jFdcMgWzZwqnw52DVpLlj9xPW6vV1QLAhBfOrnHfrpYLd+3TPLwzcVUquB51KAeHr2Irab8
zQ+1NSVCjRhcBW3fnCK8x0K/oZWXT2/i4X38t8xZLd0ssTrVROdZG/efSygqYjJccvu0b97w7lgV
eMdCml7t2NszZ9pIcRXs9X8R7HyvuvW/aNqDi19l/K8ZLiliK3OVX4XObGRZXHPWxWEa3duhr99q
iHQHe8QjEwDim97cNo/1mj6+3SX14JMisv3mTYTPtga9EdrbaPm+DecWjop0J3EBBmFg517g+eve
JHUXpQRs4mz4vLJ+Ny1dw7iD/BVv18LymM+gEdX5d1HfImoBAu1R8yIxq7mk8G9JtwmM5cR/5WhV
MrSYcdJvXlXiZgYN26dqGHKc9kBnamXWw/+3dpsEGsy9/Rwmxy9JMLYO8B8n1wCqCHNUMfYYfXo8
qB0fi/ut13qrZuNvpfboTjpLpgxfXX747N60EWArtl+J9KoRNwb2JlW7RXvdyafjLgVRjvUNd4Ci
jb2Oe1Rk+rfew0uVz1lsygSiwNJsYWWCRDM8H3FS//8lKg0d7ti0bBPF/PepYcUicehgzWMuoP5w
PX34MS4UpTY+MIxb3EbZMHYN/oI2kDCJJx7TMB8P2CeUctDSddm1xPuS5YWdcY5WDS5JSeA7dZla
ZNyQ+Xp4Rkl7PD9Rs3lhiIQ1Mnu+lIFj4j0YEcE0orbftLA2Idz0pRhbGcTvj4/GK7US87LNECGV
Px0ig8wFsScjvKEHDvrkEsHxD3MEsbRPzS+yaeJISPuueTJyjjF1EaWn6pzfelO/Q4TGZcT5tNpq
3ovN97SFK/fCFlGGsTomyKRHZI9ZNzgFI00q6PrIq8s51kOrBKgTs443qTW9mkb+I+neHfoT16vQ
BqVgOhOGgAxdqdkdtYUTeOgfH9hd+AojLBuKinAz59c1PBZlSLWabtSH9Lcg8VDGj5XhATvmDlWd
1XjhDUjm2t9Uajt6kiGqJR9DL5nBMgYq2vt4BpYasviLZPXMoLb9oZ824B013q5RVCNokh/90095
v4UHFSwYgNvk2hpP93CXZuJgeSXVmNgrtkfXxd45sqeqkvrLcgEAtweQ95UK+HhomB5G//yOiqaY
OIZj/A6StkwZ8Iv9rW2+u4GenZDlKiUiFPOgfXkKHVDf6F3rVF0tC0Zsg+TgWSWny8NUbYcnQrb0
Fm7ORsdlpYiPYEyTw6MG+mZjvph86+Ioy7uI9lyn5rHIRIkrb80P95CY0fLtHEYK+WrC761teaDa
rSqHd1qmCquQaeTnIeeJ3hFyjDf5U2L1y2Uoa8auLejJhidWtwxWRvJ7xJNStzTqu3cq+QZRGH2b
LYTEinpw5JC2OKVvy0+CE69Sf7cxmxqTTHW1yo6DUw6mKeSKjXa+EJfF3lwp1W2/dYV5sovehO10
dLjfBkBES5oh1jzbogMeCfPUIKjJy4OMJWF1wnQxXOEg/IZ+Q8+jcQbW/ra2/nODwk5PEGgf+TgC
vM2zkY2poGIhYwkPK+PuxOqudIN75FuVUKiCJx1oI91YOpHOXYerDapreuZlEPn2voHI9txSEMYN
bXCs9pO4G6TqkDL+ZgHv/h/suyQHX6lKa/os6Q17+p6m/LRBFqIOVJALdN+YknElCv9Fq5Q1M0YN
FJ6CGra+N6JOl9xeraTrfKtaz8vP+P0JHhSfGnyWutOtVY9kO/CEPppiBh7M+i2RHL3cUnxbz1/m
FZ4afd+F0cGS23wrDTUvf1AxOQgpqUn3UIWXb4t/fESayQS2LGOvVznV8w8gsNKTo3hlD2MKLb17
Ahg5qmRlTuIAUYSUOqkZyHFYH0bfEdvr2MSO8doIXAdCO+w3Nhr6/tEH/W38HZ2i35olExg+Ln/y
aucdJclDNW2UqScKmn+1FL5EaTAoab6LLk0qC0dtFjwb3gOqEmn6OBh5f+xuuPpizrwpcULG0dhr
x98DhnlwvepKSdTHHohxWzx+OLIZeLbKM+P/WbcbGQ3LQqwNtWlZnWSDzW5g6cbNpalozgiVTvG0
F3vY9V+KpKYxFls+zCLpXLN0ig7VwSKyhJgu5bKQwh1+0q4rA1SFjoyjq4u9eoLTBj9/h7BrgivJ
ihhyFCQ3ithVNzbRkRiP64p+brFXxw7aQf31Y2BhvWoMFzviZr4vEMe89/Z8rU18amEv2ey5Afwc
QLwwngGXhTHLYsilY7/cG9RLAtwxOYD8QSexh3hAXL/p/XnGDV01dj/TX9ahBt+/rj6WRY3QdKQy
UEym8DfVqXeF20DJyHa/HY3f0dFpEQJZlwPcisoMfs/D4b0DmHsFa68v9MIrURFDlEBqD+M79dv9
SPf8CIdjX1Dom2ZzzYLjinyByrPKMbxhl0kOmYX4joNQK2sML1tvozWBFILnhSfRQmi/gzHglnl4
EnhiU7WVtQ4pduoGlbR2NJrT4GbeL6I+Jih2PZOa5vFJQmAyaXE0kLpnG6EpzlTGwWy8CD9/BbRn
8md2oPxvOZ1a+ThzIxRCoODnMLYtzXCbKrxjnVqKcI/frhcaWg8DbyIr7eRZzf3ZCTo2KBHXeU3I
Ct9f99whx+uW+gztDY9+mCfTqgVYmz7UJQgvXqg5aanlckNVqos7N3KsSyZB/fcR4rhCd5v+3rOF
g5jmLBK5IRU2Jc/pLQDXX6kC9rZx4Uiw5fdFrHa2PhNbLUo9sQUR83mCNwdOHfwqxZVzYyKx56UL
8sdJiOROwdFTJiiR2S/3P0oD4MIfuYgIJ+fr3KwhAasSstSdOjfN34TU0FQsetErp+UtpZZ6n3FI
VkWtfVKBsREy9WU3BSRW0uG57nJ9aCD+3siCSFffPJJtL35rks35FA7selzU0Vk/s9Ug5v8H+YBV
XXECIYtbgCVi7r4QP5QLq1C7/0BNhi35l84Vi+JhQYBw0itCkmpqhgeRKplvTZwRttoEgwqHW+F+
BEdT2ayKiAiGi2v/8LZQ68wVYubnqyiRFpwBI/I18nDOryesAqyD7940DUbZGQ6JxY8qs1PyIKbR
4sAnDdCiX8zZbgC/9CR3gNv21Zz2TY+bSrSA6WNvDFyWQ5yycNT5k5X4FQyrlp9Fx6IpnpBu3K8I
es86bbl8NyzYBZxCpvnLih/dYvFsJRvTUYQbsw6DjqhMqtlhVONtPwP78nO/ecDgPVPOPa0bkpHQ
Op8EgQDhDlM65OMq0TZXORFbivmLJtAhmGJuJNrjy6+osHhGwVGpRPl7e0e3xd29ZFf2Ngpw5qOi
v1y8cTJrnT40iIB1cq1V7nCrYQxc/NHt04WsvI/GBZb+BnEmhIVfyWLcWg6ZFnb55w3FMn4aDdtu
oD5Oola+Ok8rUVhoX/ygiVe+MhFsLhmgyWJinQjIPU1PbiTtULYWYi7ZbPen3fCE0bznuJLztMf7
cCOeLbrWIQfgrWMj98leKfPLW7JZNAFU4wSlXOneImO6bS6dyNpHGdhLAHQhNrCXqxq5OwLlDUtR
33OlLhsZ5HJp+g20HvLRe3M3bHnOLXY6e71t7vs9plPLFGsx6y8kEcNcFJOOLOf4MgRbkEJxP/gp
VyHCM72U++RbLDxWxd5xLb2dnqxkp7Nl8Xt2q/9zGC28A5l9KEc4r19cnY3b8/59MbaiLqL4sBZM
BUs4joRaeqYhDxMfziDngkE4+Nd3+P8oJa7ga/DGGJ78y/ghngRkAi+7HCQTS5eJqctLSW5X28Oz
X5+T6hbsCFtftwvIQD85x2sE+ReHwu3h2atorjmDcldOYZMUSenReczfMX0SbMTMsmGxestXgMdm
SfNiyW9dfDcVtJBfWXaLLXU6WGqUMlx8NLT52VcqtpM93pQy8l4yli5i2P4w6Dnz684/SHBKcdDl
bKBB3il6ssqBIzUi82hVgF7gO5OYCB2YKHRuJt5aVshCPth1MFhCSquBz0w5EB5iC5T1gBl6xoiZ
2M9+eLZuSPqxKDvRu1dVFXczXr+PX24xVB/VfzZp6smWcPe75WiJzKT3C0xC0MfLeoPVeuwBzF1S
b5h9Pw2vygtHoETckEfAgd1PvJV70+PMc0PKEitf8WGxlabqHBK+DD6kG7WDo+cT71UnhZ6D0o1z
P5o/tuykRuMYUgrBhST6duYuHebWaxG24QqP9JfD6DZAzkgr3TBswElMm5K1MtyoRCAwzLKcSHGc
1K2kw/NpfxNlPu1u2wuPek5OVqDwEw16voDb6SPb7denD3l48KT/ZR6PyfD2fvwEWYizn2xRsWWs
o/hCP4xX9QlbAjPKiCaVWxqb5MFbkHhrHFZalLpmP5YAHvR+rO7mXoWtobfuz3DP/uH0gTAIT4gP
YAuky+lN6RGWMTmPN0+Tc2BWh9xbT2pn1zdSDAP0EQonjQj6dT8FVjcoU4WBJUW3J/riG4nf+3RY
QT7czI4V8ZgSH+gFxFATU1BhB1aUoHY6YDjJuIh4TYXwUytWmhh2BsEHCKcXnu4N8EMAPeWk/koJ
AKOF2vPNZ4kNrGnMoJvpt5ZxR547UvZqRFNP5UmuXbKfk7QC04o4zvCrxe3ppXHlAcmA4MJMDRZX
jRnULJDte5zXU0XFiZg+Toe/Ih18aaQ3M+ofKmVR1wOI80RcZTh2ifGiG7bDfEZV8EcIL6SGwzzU
vV0o7jFkqTwT/9avldIeLHqoLRlXQKUVN1Bg6yb+Ikve+a0LbXBRowx7GvucZ3ifABJIf5ZvYAtR
f0B7bq0O7i4GmS3WzUacUp+WqHAMsJpwzbSudolkuiYPLgqZiOqMcfDllBpxbdM8e23k9Q9P36iz
BosyLG4lMzR5CWXZ/MKVAPfOHNyWVUJmOP6dm/2KDH5taoIKFgcZMPlkPUCeuTTjZUPJnRKY6Lv7
mtX3fW8Zl1s6gzT0vLzbVZqI3u1tWISp5+Mic9qUa4vzuzb/i9W6Q46UEVK1UlaSXpJ9o1JvBc/W
NBtYc2U09W07bbyJq0IRVu/oaBvZbremR45RI0IauF3bDwItdYaxNSQsEZSBIj9MyfmwRGJEd7pt
tONxHNgtfmz1EhO60ti8BH2BVxMegjCKWpQbeAqJdLNs9JvY61dk+eLYKqrfcyU30XcHOPj8E2yO
7uRiv5zHVWPQOSKvYlZVMiJR3efh9iIic/OSoA7xWkIp5Bg+xwuXRFD3ZuXmR5JJaBdjDyLn46Wg
7nTaW04aKM7h+jvxH8xXPD0EKNId4N5rptnYv2g3LzuTdwggnuC/n8YvSKERn8F6m+gGD9RR9FaU
N5QxazgvsoiOrB3IvS+COn8tq/SmjyOsbWhQc495j3HZDBLC+ajM9vrJFFIli6VsplBMqqkTsBP7
MWnLvhcMc5Xd6RgJia4DpQPZB7vw0idmcuNemh/dEkIv97NiGQGnOZP6pi5fGnRFokSVAp/ZIOcB
ePODf1ITtoSAjcKhUn2xwfz8G0llrf7U+MA5JBEo42CF80DE8WWfrtXBhh8Xc5vx5rZd2oDnI4cb
+g3P8YBHhKC0Wg4yqn4rLTWUwbWerNIBNI5zhBT7aJdN3BIt12K0YC/c04+J81sqASAnLXljzXCF
kAOougZOAEKdXn9ssmDbCyUfy98Ed0kSPxZkwKFucTvD0umBuaZFF8radFKgmLylSPMSbJ2ymOC7
W8RH1Y1DZ+oLOQoGzmGSZpaRGvCG27pAQcLaf5+oee7eA7gTxVb3Ngw029xfGrWisO5KlxPdVm6b
eTeseg9WlvJ1gUgC90ZK1CtzwLPo9cX93ZWm4CitYzbX4+AtyoR1SMmwfIn42f1mcpi3LdZV8ovi
ThAQlcyN2Zj9M2c5AmDCGi9O78F+PhYyhS3KdqLcvuCEGfeT63wAgJG7jvIH2yK3VHvSXbm66vQy
HKRf/dTPXKthDpSqkxW+qzSZfHce7ujxhL8ycQjMf262LhRq9zmYtq4kPPGWlVQfxwwj/lprmbSP
2slWMbprThqbPvQs99fS0yx3FATe5EL10Cq8l1I7c4kFnJoLxaMgvSSB3QevrrV+Dd5TLLo/64kS
UNQMELx8wMaln3pAkP2bnSHwz4IeAdpK9pyedmpZphBuZRDvKu8U+s0JrOc0EKWCburuYUxGDvK5
ICSAxyaWnlSzbg36XceQF4DVt5UsjVexCRPm/KkdhjfgG/YpgwzJtLpzedVLh/gnlJHGhMmzPWT5
t9JnRWZy3jDgmJy1npiVVXuWb9z413B0daZM8XbO0u9IF7n4a810WxaFJJ0Spr2ICro4cAi+rUgo
pBTvK+bH4W8IuPLlxRMHSo8kbEeluIK92kgijoxVtqx9HIEc+cQbU5v0Q+y6hpxIQNI2lOr/f9Q4
DvDOfs0aaEXwjECa9nVxndRV/iHagMCmKR8MULbGcn117DWUpgvvBoTepCFfeTxy7ejFNXqHupBR
Yvn8S7OTXlwXHv1bMddNBo5tk02eCFby3lvXcz+kd6+if7M82/YV3nDTXNo/CypTM7KpPhdiGvcQ
lhIwK89teyIzHyV6gC24uHw6cCP8noNax4ZRxEceDwR6FdkZmdg8Mx7jJj9cLExUKhBu3LcKJZr1
fUrgzeklJwoECuL6XYMQ5BB8NOfBV9ukJ3zEAsTNAUh6N0KytI01p2W+CMGyrFOvXgSVPCuI19se
VaPGWKAN3/8UFbVpGiK1sOiCwDl17hUxGGI27ihy8mtRmZz8y7+LVSsyA0NzLu48OMefLBHHr0k3
KAC6LmAORzZUZ9mZ4/jHkTkXyk+TmudlUy/m7BfAEMH7zrNWw76/CmAcHvmt3wZyEPzn2NkLYXdZ
S6CjXQ95qUxOy9zQ/6Rl5m5oJRA+Y/xXzQ+SWPkYw6a9FTIOnPnfxXU0b5pacqyLn/4O1SptKYEB
jzkFEwdb85z4hsyHWxvMZfvg1ygWOx6fH4jaOc07p9752qyl1AVrePC8XXnMoODSXs+9DfmN0Utb
9ZxLSdx3FTHWnrQ/9oeeH3g9uqQDGlMqFsDJPvs6oCIBqRtZsJq8fl2vXeqJ7fEF3BZHTjI7kKe1
guWUDwBbGKjEmUjPEXwv/+lWykEKrRPJHz4LTWV19xuN/xLh263znxzLlJ+One+Wii3B6T0maYub
C+mCKcP32KVvPPPB1kOuUlQOrJJZirj9ugjS9cx8D+RzgVIqaOyzQ6o6Ep0cvSCAN0Oumg1y8UNX
qOQ0eRKthbI9Pam0hNjzG3HJ6CM8/SkdJm6yHqbOIBfK3aXLpybvE+Wi+1prceeyAXmdMf9jfuTO
3gUc2zWLRkt23q4KxeLjsC/KhzglJltcIwLj5Jj0EZPdusT0IxY0e0bxWjZ4CzPfgEzvWp+kjJJf
49znZs6kzSuLOPoxgfG79yNWdbkHDzv1OHcYnj8tB9gaEGaRbRkADfePpBZ358Xy7Pfeo3RmWCKg
/3rhXjLUqsUOsuyt60V+rpXu9YObom6nE7uvQwxIZBVynClSznKyy5cWiltbL50NI3S+PUMXRsXY
J4ab02efkdUBloGcJrqwXz3ocwbMn6nlVMKBOIEpC51rWm/REqrfp2LhNqcpNj0q4KbUAEL99dx0
jN9I3nx64JGFr7xTmZBHkjMeXDp+siJd9FPBdhUSam+zuSmnAAXP6GIUZql6qajKeQMBVLd0fi/o
4299axtSMrC0W8wPjWLhTYKyp1u/5ssvSRDFZ6XflDjahBIcuI2n8C9yML/7GV1P1SV1lkUZfrG7
i/YW1SFBvyGq5w7b7CcvHPNiWYAo69zOw4MY8ln76WH7NAqA3YbmT59JYT7LA3eoyOb0ePIa6JQU
F6/d0y2vMqI7DgNxWb4vaKdFW8+ENGarLU6Xj5NyvjBOps7S7XCoqjxKR09YuZIGLmT/E0SW1qDK
/7puHj9P2NIyU9VISx60GUFn+uSqjIrAPR7/xkNyBytb4TYuO7p6U1mXVc1rqv5PBKJzsoyx26jK
rebXmbFvy1NwaAIIiojZ5XWjAMrVBKjCUXSp8tMr9oc6eftDXmKmBC/GSIQuUI2nAIfyErVgbXtR
OFyXsnTSouE68xgVDRtsic+yhh+eS6MJejvupXzdyep7WB6eC8kKbl0WX7VFzQIPRLlKrxibZD0h
B0BPOcQfcVz84TFuoGIGaRloBiJWFjmpirTBTXgdTGD0lXFK5wRzocwK5LAoAy/0F9f3FBXrUzH2
7jF81yFsrd8Q8JDYHlLz1OfkXMstycs3HmywXBtZ+C7ZnH9wrpiC+P4jdOAX6PdUaAEFbXt+KgbE
uhoti5ReF6PROfpZj8DWtk9RbtbasTNDe7fuRd6vpBKf/5n06WC8ea3JldpABzctHhrn/PzBZmtA
JgW72y7K8JPtJPV0row4ji/FG9yRYUuCRRlGkIQEEZOl1pMzNqWt03dsvjEjhHjTY2M/CCVcIkMb
03G4bj6uTfs87lsCTUBbBj4OqpJjrUfOy0wbcntCyVxAqlEPmTjiF2xl0Aea4R2oSzyegRWFTSgk
a4EYA7whLoj32yYWcRY1jOkEqx8iAPMQWEvPqdOfdCuxj+254ORe1KwCWehDrjBG6ubCTg8qigRN
2rYT/EuNO4tRoZRoAbTvV+nJosGOmKGw903mccTmDk5xFOym1etiLUGD4LLOXwHmLpwATIurHCN+
UQj+BsIyH8Q2nVZJgzrDbNqGZ67Ap0iqJ2ZcbXhpIZNssD0Tyfcodv90ur14DjYUB9FDlAT/6rm4
u/kw+Nz0l8TpZdVYSSjjTW/PPanmsfHl/Iub0U+q6C14gWslv0T2qKZJw5pbWdWrtKATlZVmwVwd
pJXqLO0p4j56fCsJTnj+rCheCqHvbqLEyPe9M0jS4/a+b1OLgFKzusMLBPE6ZqxJ6TUKiqiPz3sg
CaGz0qQ5hvnaDOVogp1xk3tc1ZjTF84ggR0BpUuQtFrhsUDp0Ivv0YT3/gixru1kouMBEkk2WWYv
O/8b/fA1Mr3pgvQJjjTVFa76YCUWfDSKa8Tg/hYArzcMd8I6qJwEKvYgl3wHANSlOXCxknT+ON83
hEPDDW19IH0GPwjIagbKxGju2gJkqJg/OiaB7Kq99goaowzxnxEhvxlgdkyNGHE7hQkO8LCAg5rp
JuOJjsUkQaPhnnUE9Fa89xi+Ts7XcRSvDxdwfLuGsvbujLk8UWXJIccQmP7Stt8hINNo1nppQIWg
pE5SN0KTQAtZevWr0LFGMF13IREOoK5woeYT0HyQBti942ndKY2O/Gji3b88NcIoHZdosdhovrid
bPKuVt1BXCOTq4cNsEfNLrwkPZNtZjg1oBoE8m0Fj7mOWOInWSXX05q+nC2yLN2aNKkI8qIcRrpX
PBlJrwDd1+1bIyIsD+qoMGHuElZkWaJMhui6NGSyuR0REIkhhwKjHJScX/sl9f51AMNI1CG+08sU
xpeW7H8uxaRaaGeHE38gfdOYegiSVVTJoMY07s1APxZiOVhVHd3ENRHyMNfgxqony/AY599W5g9x
RAHPN/7VrQXSfSIlGeaRqVY5soR++ah+5vcRbXSikaTflxPfVfKmE8jWLu4llRbfAoabciGxbgZr
Ba59ZP9Mjo40Kxpp9Ws/3mzKM46w0NMhz4XSRGyoIlshSL/noie7m8GUqsEBjGaE/lKKcRb0xgJa
R2D2nSc59+2Lzi1vdpXFROGv7TpeIAgS11BOCb//qereCcjCZctctl1ZrkkBoHYjrgNgHwDZmDYV
0HoBWpFhz0nvsYMNaqZ7gDKBcrPVZWQwW29lkb4qqalljr22ldL3v/O9ZTGgE84ldnhDOlRJBy1H
6QxkGZYaFYdhFhdHc1bNkB3+2eb6lz1MVJq9o8Qrq7juotVrU91GEQz0q84SfblcHGK6lTUqQKx+
ZaKbkJlLMndT0E9X/R9898rJU/gekb5gDBmQ+1yU3sdgrizvEcpxV3QCCOhZ0TtDw0ZASqTBmLg9
pFqePhHTeG7UK5SMRgc5oCtr3q04EK+K5/VJwxG3fl2L0F8t4NWpLbGH+Qk3N/lEMnT6NgSG/M3v
szVY+w4aC9pnC3SmMrycinh00gIbWaSR90ddT+vifIWjM+U01MITiaiivGeVEhNJ+nx9O80B3czs
tBT4f6j8zBnMYBx9symWhFmtHJJAqKeVZGiMJJrmlMRYWGZYAzWunSWyACwGC4XtlPrWvff8bkyb
T/GG1FoRwj0wxiWG0e2Ut3IN8TLNnJjHZqrxRoxvjzpQADS/qevQe67mE3Efk/1zuKTQfHSvhMBz
buJq0Iwenq6Rn7ZlnQw/9EkBQZFuVCguIgrjLQz2Y6kzpxqaP8Pwz53Za/l37SDDBxXPfTvV6C0Z
9+5wjAA0L+DKJZC7H3/PWg7dZZtyJVM2j6zncAvGgul6mMzmX2zDsxlqcEBDicG+Oe/WGcnSzvsR
VJVeTCelZdwEufXAkdM3C80PoUIUK5Kj5nL6zEtQ92jXrhEGcguCLvnep/Dz3e64vmlEkToTEKYg
aTqr8e06K0dQdFgKi14F24rwpHXCaPLaA9/RjxzU4gHbR/rc9GPvIbLFTwv2auVPhqO1+18QPlgS
Qp/7DrD9xdUBth7OA0Y3H4pQT7VSyaadGnbv8clvFmi5UjYNCklFkJf8U2+W9lTSQW1NoS61n0J7
jzFzVSVMy5hga1EHaKjTZYGRvhdigvQDUHVz6UhRuehZh8txXYx6BZLR6FqH3/mUGKarzwuMpsjV
WLrcp4vlvhGuY6meRvvbiz/2dFuCiUUJx/FTjHYu+S6+mW+xfardQM21N7OUWE2kvSCklTQdZ34s
5Lo3MZOG3AOpcg1dVIJDDPBiyZ4hFWnHceNmZhbFL/1T/hCA01alJCu5gBB2S0vqDwc3TYaZ0Wcz
dkub/zUom0dVHGdvQOoemT2ZHU0PNJ3ANnJWcESA7DTwoTBcYDiY0k4mw4HbCvxaan7o+F9lm2kx
cmvU6JwNEysOELNBAmai9lofSkHkJxO3Q6E/nbnTVHHHBcAJ+DNbUHINmRa1ir4OnVRcJmPhAI4C
RtXiMKH6wBX3P2ToyIn5ddz1vRyO5RMJm0kMnmxYzaMiPFBelfIYzWlPV+99ZZrzy0levUA4iUhg
6nSOsG5kggQhubMzPHgUhJKGK8Wii3qKaUBcFf9I2o9jaQJVvJxclvN71iagLu5LA7koNHgL89ms
JAAKiD141vKP02NSMzDyl7Ki0KzurFP0S3OPG3vBf3a0hXg+XNg3cKbouBa6eogP3jbFhk61nq9V
iL+OSLR1vrQEwNYDQoafmMGPfVsCShS8z8BpyrGsG/JEKbPptCxFBYydhH8iTKERg9y59sEzjH5D
VsoUYpbeijw+oqtFZ2S9Zexfk4GsOju1oCgnKBfjLbr4Y9hupHuh02tS8lWag7KHQnnH+q5/v+6C
1J+xl2O/n/ZqElgldzIuEzauk6PAhA+xUCobeg9wLbKvKZ8BP8yhuMBA/5eGd3qioeuOX4LGY+az
cuBK377t3m7yFc/Qa8pCs9ymkfvtdM3ejSHb6wnJffiHD7tkUZ/TvgmPCOSxdYUFTChZwqdh9kgA
EOXezeb/Xx8k0MeljqnT8okbtNwrZYRi/N5K5sU5/5QnXbKnCOdlo+pFF9IwrV/F1BWZ6e924igR
qspEFwxeM0EudP8qLOmC/JXMSS7rKA/J0u0DjU9U/3XDwgQsCIAexJUkgPQ/KAEta6Wn62f9xaqm
IxMYP0J1RMf+yUIW7GFcXJCUb3aflClv3c7st1cvMplGnZqDG+NWjGt2DVKhrU1mblUNBebkF3tb
rVixzyCJcCUXkic7LbSA1KO227nFsVlI+05m64eqlBiqrIOrapoh03nRI72qE8IXfFpbe3oa8ige
y92AxwrNhWvivKJElGPN0b62OhMSGxHPQIjsPTKetTWtvzPG3vhzlD/72hVzGcy0fkNFbU7jF2k7
gFojN86OgqfWBZ/MaErKwizMrUbSWLqorA51lysQD4iN5b0BMQm2qsZNfRYMiXk07CcIrY0f3Lco
+ccsyMB4ptnH6cJcigqle5+YiBjGMEU1kuoctOrgYyjPX8LhB5I8cZRMuBNWvL4/efsQ4ee1jSMU
CpPu3VRcwNblFNAhqwOcIiL2Ov+8Kf3m4kK6bQPcL/5s2duR3+foHDQeKlZ7dbUvmAvFf+5vsBbQ
jqmfUNN2kPm93Scut7YUGkec0jEHFe1HAlwfDqaasHLreXO88ChHLifERoCvY/QIHkbcdlcQdthp
C1fKHK7ms7Gcv8zxPtu0eU9K0ze5E566shndeWLCZwO0djljjVkik6rSjs6Fhsw13IaljQ/ShJ3g
ncm7Vbh39YcBQkNdHvyxLYDAHITuVlcMMP43jURE0ESH5zISkZhYf8XUiQ8ldcJiBI7V81GscIDJ
8Cv4Y879jsVTn5V+JlmXC8abT6qrL+vo3TCUOyTpoy69+BdfmtflyUp5cTjh/WoBG7nicoxIYkaI
1HdxcKFZDSKFuH5Y/OqHe4QQL6H8ZqDIm6x8UaapnvZq5wvcJqli+bEUalrBhis5LLDK6P5Sbtd4
eEwnEuHik4Q+sDPsZq7YnzEUNc2fVTNgo7IPqFcipMQjko8Iusml9KHhoehEe6+to1GsrhSCY7mB
n8nuWxyx8FjyugBaIr2xgN1CGJhGawPOv7UKplZ9/mzbwBMY7Ce2BTEeKzCPUn/bHecEoXPIt9T0
eqNfI+EDF+z2ZvbIVEtOILWVcHX56phdCgFKy38IjDqkF2z+0bVWhsUcdhg/2dNVt2OI0ddyvlFw
496NzRlCToJDHC0OQA9UW26kwlpJMgQERhsc0a5TsusFxgTfkcpOPVPWsDseiPK877+m8jHs+Mn3
mVFq/ztpzyIqClJWafMGlOJDVZD7H/3KHnUC/TIe4eX2aOcKUl0wjAhHNgwNq3z6PLAvU2lOfOLE
YTud4n5/0hr7sQVxEup9USsNwDaH1xEXkb/sDPZTc0lsiar30xaf+iUfG+1hmPHhjxBlPEMKjr4x
ZIvXLznQcvO4QVVvnrt78b+f2jHX0weYSQvkuiS6LPOHCuviZzh/t4JuRFBPqaKFw8cBG36iWWUv
Zc8oK/f15aOnZY827F/5AyOOgVvFh23Uwao0XK8MQ4QQAZeP9bwGE+/mWkRTBbum1Nzvh+xHmXm2
ZFqhJnN//vvB11uy4DTOSzS0Bhp/qgZjKae9s+zEMZAU+GLSil/1jn5yuoeixlQ/Y8SxVDNG6AEw
3/L9JAhwp2lghxhWpAmGU8ZUUkwbbLhow/PQE0FZA0Y/JDVYt5nLspsr4QvgWbKHehJFokE7DolY
Gjo4UKfEAWahhM+hfRQhCe8ycUOeuoPAdIg/B9onxRG3JeuMjXm1PL25RzSZXbcqaz038y9s9tf7
gzPjhVwh6ad7oSkqnt/AlDuK/EsMAc88zlfD95E3T1tZ6Hk+uaz7LYwvmSge8TvWP8jUbJO9bYtP
8E/4bOFHfhMu8Z77YW3PZvwdeq89IIt9Aa7NP6EYhMwTpKJgPHILDv+Yk9lhBX7q0kZCB7a3cTok
zQt1xBcpjhsNukrZG/EMePBD8P7E4kI4DvpAFzTSxJZb9W1d181ckD6UtvfUe/xrku2SmdY8fNrN
0+Zv9PDNN6x9ZKJ299ALglyIcPybRZRHLozrHppiUMNhANHmFIzrJeBk8oImzUdcfglWbktqV0nf
DD5HGXjBWO60dJgzJ+OUSbQrtG/0Bfvo0qZlP8xCfmsJIqKIW8R2GVkLyAITjgw2EaXlCauhHXfR
DMG/9/g1ZMuk0e8vX/vlI6tUX+6j6aVk17eZzoHT/hAm78yYlyUvUAehuw7vhJpRI0iW3kDCNa/d
IHmHBUKo9aBsfuJ9IEx0k57u0b7Cmqyr0PQtdKx1A1xFwUM2RS+zxqS/jcXvF/UMNFN/seMK18P+
yxDWI4Yk6QGytwg1WxEbJIx2AgRZxVE5MRoccUEvBLx9TxQaHWtk7CW4jsR++zrFfaIP8ReJpefK
JnB+RuGw4CaO6D5NyneJmkJva84Z07tT6lAURwD+FnWWMJUWNYQca3AxqovCn8o7WBcZJDklXWEU
Es7B478lgn4WQi3EUA7awpKHl9vNct7vHhgupjyDtqN1eBN2cnCxYKYu7vKE5GYxpQnvPLZOprWP
iuF6eEHaBTlDPKpC56USw4y1fjB7i7Wvt+QJeeG5n83EuBRTUzyguSItHYR0t6v+iQV0zNs6fqNg
siaZrH7KYB2NXei38JiCNg/MAV6gdKeer8qv1eF4PWObeTwKIjREviIVf42ykqmVs7I5soSmXIai
OyLkm7hkldkWjF1wraWLjADSI075ChHSbC5/4YJd7TPOScL9B9ZO+LmxuD6dVNvG38Ut+SAfSs+g
H4fFa8C3mZyzLYaWKa2dgkjQqQq+FGYhqah0Qr1fFKAig0777EPZc6yY8SrUPpBy/a5waqz5J2fA
jcEkNeINQWy0dABHy+Yxz1kI8l78RdM+ECcSzQH/5KmXc1eZKSPE4FRhqJeJ5SOc4FAJe3QAkZ99
hhNtQaoKrhA8V4/hsviJ0mv9TnomjxW/dZKALlq65GBMFAbeqFrk0loPKsGbWxZC+M+ySk87c00s
/TCgT5Ghxp+quxAIPY76SlzSmDxESpybISPKFb8PAPjMtJCvSp7svKiNCus7oEc4Lo6ZOY6wu9rM
FG9OiTMBRBLTOCfsnC8lpe3AdAuDoXezFxsziyxVbtMfhuf9NqbDwm2EwlRmK8P+xQhVgIZF7J7c
nPMAvfH/lGCivG65+Xk1Fi09ui/Ur70OMzGpgAxTn4mT4UoQTP0XtZSBIArH7gfvMVqLY2UACjzT
SESVepUpcJK8K699KWShakKnDGda/FnsrQJ/8Em+iwKMgsm65nJoprUTzdPqzZ8J/jCdspNZqqjp
6qpFJQDWOUuQU+BJcqubHTaDY0ZZCSAus7HTGoLn1WJ9OkhDVdlWMt5ctMYv0jDtHL/aBggvDazY
Zc+CWsQiAblkOfeR6ydUZORElKS4avKu7gQyjL1uxeZvD5XtTsXmklrxWRVWBkQheKQP2Qh6b2i/
ObfoyWBjbLdJJ0FotxaSZH9fkDb0ksbyMZcYL004eZJiHlzOeCOYXScQ6HQUPffUY+FFUyNFbrzR
vO6+5YLh/dKhqWkgRuN0x8KRCi4msaPPWI+Pb1J/zAbkf+mJSjV7ak3+Px7bYwZp1i5tSNdVAOyV
8grIoKgWfNUachzKo/ghJCKTrksXvmiOrbTqnRxzbF96uoJIj5u9e8iQjyNr+fLsOj4yg6/XIjvl
e3HVvngRQIWVw7Zv3FgBVfmIGatoAVz45e+DuTC2w0lOgHq3ljDfA5jZhq5SyX01Z/4C9LvnLzVe
nOb4DzXmoOxxryKGBuo2nvu9X3kys/Z72583qnj7p0xdCdjDk1vsiwpYnyTFt2jvVkBO8AdlgcPN
yvnLlkLU+6b+012RutO+UpPwVtgz5HqZ6XFWXdohIW4lTIkMqEbp/q9etrzT/Bf2Vi53zBOKrdej
mLGpu0jLAsMHaeiPC/eNOtdxZw3UR0GBkoDL9TjCZp57jdcDYxNNJ1WGKUtnVG8ZK+52AvK4HMzH
LrVT//4tX4+DoBHoaDrYYmuxB0iDJhIAqWCsuUlQRt0kTECeVeFOlizr2hj3KLF7N/ziZU3mYD7K
bANNWvEtbQbifPIckUe4QpUY9EAXm4VGxo1eN8iXx5q0yKoMXaqzPUBTGib0Er2hzsaadrYqiYyk
xmjeV/XSb3PujFWSZu6w8UNqKmA6/cLLdv8U69ybPW1GBWogTUM9/lD3wpe0QGNeJDBVoIo5m/Wa
uF/uYxg3wKvteSEhiGXy6Xjp+Uc3vHA/gn3EVtUtZ+0l3gA5POGpnLC+Aa5PAmcu4eqpTzs9TVvM
GYY9gXOK154rb1OgtgqSQDntJ8Q6xtXPZw+uRzvbpn4F7dN//NsRxTN8t484X+OyVnJdwN7pC9cE
AETPm6cIN4Ou4y6Obj6OXMfLj7Iy5p8U2NdKI+caT6zdJnHid6q8HX9YDFD0Dm5MHU1ttbdUKxir
gfytarfgux43CCm1t6fIxrPvZ02Ygc/T5jgA2ab4Xpg9fCdoBhL+GDK8c4sKEGlIj4zmbBM4mA9R
Oc4q9rrCqq/bi/5nQcFXhPejUWP9b7P9DV2fM1dEdQGM0PnvyVwuLbNcrvWsnnRTenBbC1xzIdB/
TWgThmATmnghG2pQ12lcUhy0dy0/wvMhkIBS/xfmfhfDhjJHX+pQN7GflPBuSYYRlJNeyaeZryKS
Dlp6NVqsuBjJg2VFO02duCJvQGub2XvTqaMq+Lwo15sAzO2X4he+pS5nOn+jBsmvQb/+WGDT6hPN
NaDRsBpxi3/X3qoBl+sq3ngRHRYHQ7CtJRdgdmscKHXYLxiS8NwGZL9S4dHZAalVJkdAe974DfFN
eZErG/w7rKj31VHedWG9lwBpJZaPZPHYaIq8jr9XnUfRfrqfAbTNHuYTyB5QfO5ZxHMwwM7Z6jnm
7SluGVPeFBnV+S/Ha58ceIjfQwVaiMazJN+C/j/SR8gaG4F4MyR1cSbVi69P+t81gEMASHy01FGa
+gBigFFngVnObX2WmtsMXmqzNSuXKms2xsXSCMHHmiUK16C/AMSSQADSHbJq3jAniE/6HLi1ZcMi
TNPtZuyBoV4rGVwmWOwxG2nFND51+ZVjgriiUxi8oKmP/04U/TI+iVTHGaR/Y8CILLfe2zKjbIcP
5nUd+fk6dfcHVrT0bx8sre7guqvZYLXDzB9SghgBtLN/o7SsWg+ggEdY1D6p+v1AAFdEPvZ3kBcG
ueWZwdkYIMyQJsG4yXReEmqz0ucooyScsBeo0MGnqezkVIhvFe09xsvuhr3ahSAGMhlKXfgVW0RN
9RS5t1UQPcSDHljcKldyxSqJZ5Eh9unVH6hdRGZBQFY583GRe3I8xYYaMPi73yj8ZwqzpFDEyX8O
Vq/zwXa6S6naXbJBc3a2TIFzf9uWvUXsTmF8ihyYIl5SazSQlp89FjdynNOt8JUHwXmzUiTjVMbm
8Gmg5oE56d7zHLQFELH2ZfkQpe7sp0m8y37y/99e5h+3ShYx43D4Zi9TZIlFjdx1GQ6MCuTLUys7
jF2VQzNpZmD3l/u7pLFODMOFs8+0iN1Q0cWiYkjIIMrR6MgkrS3Pf9AIvGwnEHShLOCJOvbl7cbz
4k0wfriRPCkmej9FH5/wiyLeLWEhk/mfGoGkfMZbSzP4wkikgZgnzU9lX8npFY4FjhWWIvEfqnDK
UvP2ruil4+ieAPWplBhSpib9kyMHnt8cRA2unK824F7c+3PM218CQqFxKg+vUymjZTtaCAj6TWiB
96CUMPAzotKOJxScoGGSpBNIPFrFA16+ESS6lhhLNhd9mIfynlxXZqoRHEoxDsLRodjPJqOtzfWF
D4X49N13p4jL7K7MYel1HPFl3wSWq5IMuPWfXu7+ZkkTBVrdnErF+Iu7h0/wFCXv3WHX7IVi+W/t
j1pHVSNo8cS54drAZ3xjlAkOTDR4Kk/5ccw/8/zRUGCoeTTrFlFfXCAom9TRSUf8dTcF4mj20Vf2
dU/CT0YbDeT4P5Tv+w/zEx//ft7YfnrLYkaLcZ6dLNRVRK1cm7AObcuW5c2otgU4ZxjhVI9dieGr
Cu8/kiFWBcvmS9pm9tfhAFp8/4koagyUtvV60sbv6XJiU/lAm9/nS5SQqUrbHYq1xBWSoJSIV32x
4uh00C7mvv3ZPgNIPSiiiAEIsJ0vhAqVtkdgV/z+BV2zwGvZYMOFJCgSIOvIPLfusQO7CwexV6jm
gjSYvWmXOzIGCfseTx8mqrtEtZnTzAQAD45xd042GwpfpJTSELUsryEl+BBXqulkCs7PT9TGiV/3
hXUiJHxSbk+efG6ncoup/SCQ8/gvcs12Dr+Dzm/+RtivVt4+S4pcaga88LhlRnIbOA5oGdrSFJR9
QyNaZIhVPUrm9rsEjqgOq931ATLfDNhgZgRAnuxTT4Bpbf9E9bHh4wbyHYsituENoujowDWSmY10
Ipt4ejI29uzJEajpzdQc+EA/vcXFmGggBtdKo2GRgUzg1nt0f7jXZGfD/dovg3xQ1wZQQYT/GUDP
7uWmBaDSjaafg7uiOb2+Vwqzl1aPMHYvdxySeKRZjxtH1c0tqva46joe3JTXsGSiapogc4QqUBYd
WU7auBmbvqpkX1zFBVjpbRAoCKpU2cS6xZ5+64L/twWQQBd6jPhrGW3Q8TXa8pHS+Wub3axXO0DA
ogH5f8rnfsqryOgHZYVRZqB7zfQHaiXWkOaMOrmv0CgllvI5KXuyN2WWyuQt3mJslzLmBZfGReBV
SkGtQYva3Es2Q2UQDXFs2SW7O/ydAQPKgeSLrm4in90mgfV7siRZbEPx7FeJhb1NgD3RSS9qrmXy
dsF9/igE0CxR7ZubzJXVs5qfhkw8nmF06K/ttKpXxWKLAxPB8KdpSrllkePns9RDMdmFuUFti2yA
g+yYUTSR4RrfoCzbTIvkqwmuuivrQNZndwUDSPXRwHlsY7V2hifaHug62nTBUNAVun3M53LnZkpU
W8h2bJ9O8iE0JbeaC28ve7JoG+XOLx8MSyi37HboWzPLA9P9IurKHbuxLIDt+jqSbXKvoWUjrGEA
51npQ3sd8QhayBJwi8HDZpxSvC05OXtWcEhlko2ukbIVQnzlaaV2gsHMvXVHW9c70FbqyyTgHfP/
2T7UTjYSLVvfuUPgaOhYCem4S9oDG8/7KmfeOwhlVpwnwRKu4CF6Cs3+HCV2LpSN+ONZd/Bm1hpk
MZ4Oryu9z0eD3P/cY4U0b8Cc/0tfySebOZJweiKQ7sSC02XMt2DVjQCLJt5UZcMZ0AQu8QQmLxFD
lxy0n6dcL88v2GqqlfXtzAPEeC2LTLpeykGHctUmigMgXgAj6QKtE2juqLCLXZZ3swDmr6HItjas
xQrwu7Jbebk24QFuvQVkl8wxmqX/b/ZQuMHC1vOalHO6pFVJ72KfrTquqTuUlvF34cqESa5l+U2l
OBZh8ZNlxwCBOEuwrgMXlAdsU/bjO7r+riKqrTFHJ0tvrABjk/stP26HPkLAqR3dzMPctvGHbD34
jr2eyv2FcCZEHcfpQuZKcPrSlpOAzBf5g7XPWeKsplng247JIiUZ/KPCujJerhdq56thlYmEr/yh
wBphtkVuaQKx205OU/YC7E6TDBimozx2mmfOhQWcO4ueZqNOwHZqjtklJ5SQnj9V+/O0TdBCy+lJ
QKnSBEHEUa6s34DIW4WiVlVIHKg6mvbLhlbd6dk4x22OlGiznQE7q9QgM1to7Qq5oiIUbPFPUlCb
MybC/Ea4uNDYidS1PLxRUQ/dBzZWo17vB8en6pBP+Z5xqABja6+iDwwcebeWPhMwzEjC20YOV509
ZAaUFHew7sIN0FVNcIKRubcAkB9bzqTU0Aw0hiznxagwF27nnMgYz1mnWaLpuRhaII9tHeMXdaSW
tKP+4jVN/0nZL4nY2BSsd0wXNQzv/ovUreGAhehoFc6KqcqdM1KtpSo6pfSYIJwd6uuKMzyd/JwC
tZ+nIfJI+XobqXnwbNMLJbesqmuoSRbMUHJIqC83wB/WPYCJpqHCsQY0cokpuDWfekln87swdTjj
q4IAXpnQ6EJx2okLzf8KL08OrakCriEr3TRPsKLiFMM7+QxbPq/pX8fhE5vFPsEx6LDEad3Yhi6q
uxVYNcnwztU7uF88BHiN06r/l7hcAdzMbKYnj3bEG9aOUoABOyPJmKQqVJJqfNp3Ovw00FWkyspf
8g9n2AUzCg3I85jL5hLt5qu9/J4gyq28ecwiyvqFDFfEcTKgziq2CV/qJohfePX3XaYuazu0O215
GW8LBE6eQZvjW5E+MpVk313mco6dxE8qJF2wcS/Ku5TfAzCcH3l8oTHMWi8HOe+1cCDTq+bTw7Bz
dt3g7XvuSpafTCY//v6bZkJmxZLE8cImUTX/G+DngLMHSG49z+v/UKLke6FLnnt9bS3AvqOya53z
dMayeUa5ibzILhmbDddSqan0VU5GlOO179wJ9O9YUBpK0Y2a1is8upb9mGvly/IrzrrtCf+E9mi9
baPNplY0VIzh1f65PLzFBzMTpNuQa/jqPNr07RRrrZRG54/mRpbxr4yZ/7PAsVVC+jelrFz4VZop
ivHEUEpgo3ooVXIl7JEQEoEBWML2u9U8f4+cY2uzPly86zkC8ETBFfUWVWB2G5iSYdtjtb9t0d2v
GLKDsOJo5NphTejEmFWyqFyP9bxVaK/yi+hnNXPgwlua4KQdUY/GdSJgheInd3sGP0C3yLOH7GFi
SRl3UAMs0TgNFHNdYfOfrbDxfJVUtCHYwfvFmoU70fSbzeDNyelz2d6R4ZIYmbm6kzU6/X4nncgJ
OF2bRdpLi4IGLGm6j+HAfL+YE0L05IADjGmt/fQMw6RB/gRn1UqR5Pbu+vDQij6tnhLnvZLQvO1P
LKxj2cy/X7p63wyRCTiko6+xsxbPnToWZUrUqd7jhuYtZXnOEIZfN3FRr8fyB3eYmO52P21CQVvg
O3jIQaXc2xOTV0si3fbvdxUB4mh6zfR1EalMOXNIx4GPcFz6R74S+nmgTyShLH8OO2e0hGQeMhS0
EvyIR6jBuaACQQPNnLhIvfkoeZ3XSTerQmT+JjVKzsmanyTKcpj7rNUpUXjsIEkvC4ZUnBHtw1c4
Sf1tgRfg1wxLUUm9UaBOS5zt+e4Ub+lI0S1PmvoRHGvNS/TobK5MG2eV27rUAftcUaKrM1QGqpCd
YXieMzboNjVrzJD8IYknSQtaMNhQp2PQjwNsHo++6Th48ob1zbjCu2ZJ2tqcDi9EIykjQNMwprcJ
//cPp0KVSB2A8RBSIDJCir6R0YonqHUzRGVtTzm7K2P03i/nJVK1DzpoF2eehg6lqqkbsQAcKNVB
eL9b3L1YYN4iwu/XVhyfBe5Y3M+aB5UgIksc0l9pjb2eQKGITnI9kOdSBD7U7tF2ME+VQjZqVnLr
xoHNn5s6Z/iU6EqPM6jzOND3CxZXbgGVYDW0sh8ZR45Pl1kFu8JN4SEYlpUecMxMseIyha9oEZ29
w2+1sSCu4Zk0oA1WpKJEjZiSBmMHbjq5ePr/J7L3DvbIujPf6+edbCuISvi8U1yL86Wq+XqI+/6N
UQc913Zpbh9ipUmVL7ZQCAXNP+jr+C8abmd5qvYEx+IM2NEYw22YCCgmfkB0HfG/fE6Ezs6SG6uc
93rr4oJErzeno6OuCWdPuAD33AEGlfoHtGe7WHx5qOn6jowEwEZdXmOULj1WbzckyIjLQIz7jTA/
AOyMrcXgNPRhlabNCrmz2ByMk8bglKd7+SsR9Djw4jhC/16Ghj1Kf0+oiSJB5s00x4HtPRcqDlRg
HQxF11s41PEgpfGm58gCuBwOygIC2caBQy90a4dJlsafGbRuLzqW6GHWv1AHiduuJcdHl3FtRw8s
LitKV16g/Ln4rVH5CqhpoGcLd6BEAElNtgY51oeq7KfwJdNNOt+LRrl3K6uxf2sPrlvFG+l7LPqe
rVhvkx0CTy99NaS9L/rW6yCaZgn1JcNf71oDo0YWVBgUagYU/FL7tO5rUFnzGeGNrdgOcK+6TAjM
GHuntWhj8KT6p3gd3I2qIdkTFu4pw6gHGNbO2B3etqXzkDoVDW6Z/jrA6OfTcqrtgbTJnli1QIc4
qOFGL70JjZJqWDolu5fG1S6kBPQ7jML1vRwfIP4XwfitCC0VjBdXVaq3J8usTqdaitjJ2wlihH0T
QWQrdOLq8VubpWgWVSNr/8/ZdLQDlIKequSpvbgOOH8n21wTbLfA2cK/05Z/pgy9yQX06l2nm9IF
EpSqb2tI4E7YlRojus9NQTK5rXML/jyn4N3FIFfXq2c3pjqJ3SpegViS79xG/Rd5l7pOJFrmCp92
8+fQECmrodv6BC66Egk+e03JKBRyIt1ac96420S7d5+ROKLUIyS4jR9InP5WbQnhvHULy9M7cOtQ
3lj/+PtWwOlzpKSfQnv8BURGQ/UggF2ow2waUV3lhC6tdPL2FVR6YBkn/DcPK1XWu52EaJydh8Gq
CzYHjM0/kWtEVwpPIpbHijzDxFkgvgxv9G/5oL7bPfEbHiZDiTj5vw9P5q90vfo9YERhCyXjrP8u
0Ia8pXzMAhGGz2Kfpjui++OO9yH6XaJ2fGTzlRntpKALnm0DjzyN6duqQo8cYYPs37Ye5bSzlkix
kaNYnfBTQ9ypO/a380/VqQjMuN/pgGIyd0OogN1Ma787mdwWBnprwoCA48fpWfeAcv5mDo+ZPAXl
oQZ+9G0QfX+w1cHiJw5YyEDRvJyV+7WyHvZvaanrx8C0n5nJ6YBCpABpxH2Oa7n6GjkUUT23oWAI
kMkzUwPqvmMt2+WpvWJNJswO53ny310H4qeNssWWoDhcPnXd2TiSTJgn9NdUXCdIVcVG8CxxO0EF
IMnG3r9y56VpWdbE/k9LXZ5tc16YzRh3yrcn505ACyfJU/+P5MfCYFA+a7B9A6FeUdfikgTAF0S2
/RXmtGqEg9/EiKc+uLJVi1ntaRPsp8Ble67ewSUiLD4Do5mvBWgPMyCjFQJpJg+APO+VfRscwk8c
+ZO0df2rdEzpayu9i0Rz4gKUPjO2jWjGidfusuCrFDKt5Jjjs0SuRPd0BzI2nPKP+tGMFOPgfI0R
Rl3RpGiDeNu/9a0FokRBQ+10beb/Q2bje1gKLPyQ78dUBecvS78mBmKTXSP3Nd2KnUOVQLMFDBiJ
TevAgRoJANxdn6zTwXqGqTBjKLTjCXEFegD4/nzYpSOddtCkgO4NyxGXxhRgCLWTlQqraDFdE8Y5
As9MTKipmrRUMTVwFSx5LWLaX370Cg9z5RWbRPN4ggMaeXRwJld9J2Bjant27SPAFFlxOt7LfnAk
ksTAvTxL92+ZtjzMAx/GFjaOvEsf5N9CpXINVxXYBS+lEdiIVbNaL8Ot9Ws71Z9jf1eC0oiqB8wE
+5Rvf/qCnF9IQByrxfEQ746FCfRF4sicC55b0pWRdoOE3clzhi/IS3z/TGAEjIBUJk+KcS/7VdPb
WzDqMRQnBFl3rrb7f6jWoo7FrRqGakIUH6JCR4tky9tJGNGpYA7hQEHIN3V6q0FixqWS/MsJdEW+
HoRk0RV2DJppftS65uduloWytoP8FlNx1E0deoxNLhZuolJMCcA2OGluG1hkXbokQBezTcVgOxB2
ubD6asebiRHe02oftrHRRt75j15Vs0Cyq7WN3/9iA3fIsf8+LqHUplWCZxvFWOgRdXTdbePJA1E0
EBph7lugmkB6I+KS56YNHyT1RvSXlD+byuYfg2Td96xRexyeq/4uRP6pzPree9to9RY3odwdoH7x
HOpH2Pr/qmCgFRX99zT3IDUADP/Y2MCKZvifq1G5Tqx7mEbaEPVzwV5D0WdK7BnfiXVeZdmAnBy2
6cFJ1ojvo9OnTfF8amp8W3PFNl/oNHY/f/JtjbpL8KsP747PajdTZekfIxtgdqVH3TfWcn+9ACC6
wQtTItHttcq3jxQPllfdS4okZQ8EgiOW8u5bhUfxXiRIejtjy2Ax+BUm1oIfDaWsxwj7IccIiyAg
QPECe5mo4hi1VDFnM58pvAAElPEUx5oDUP5cB25mA5AhVB1OHUep/yL9ivtiU3xH0fayGwhyT5Q6
NaZV4egrqy8egELBASkl7KbumHBHKLY1yslMwwipYX/kNoSsI4iV/TVaLNbmFJG2b78WV/VUknJP
MBe1gjPUIBj+Z+RfSWhbvYMiH7vJ90MRCbT6g9CD0j3GaIBKkIhj9TtmE8YwWaml+j36nuEWBAya
vpBPJUw2eKqbWgkLaMcbpoK1OKnP58ClLiIL5m2Srp0hEy15c3sFJBI76pdjMX6gg5DF0oKoVefD
myiKnLFXEnscUVzUVcotH3ASlLouSe68/tTvWtnUfJ6P6QQ2rP/tsLUHvuI+WdXbVy7Y9Ng09pxx
Mnn9BXpiwCUDyRLk1v3AoWItgjPwdDimtLrT1ihbLh+a34mONMpQ8X+iU0TuWnrRxBLEjijUkEN1
dc2Re125c/OCdj4qlzvPvmkoJoVr0ppIP8xglczMChEP2F9AhOoGC1L6dCELo7ZG2gxvGYeB+Jaf
BX90wRx6V19Bg+kmpJR4IZXcUa3PtS68WK396+oZNUt0P5HwgQWd1qJuGNDm0eJuHQtEIeKUXYt6
rEf9ELOUPo/83eWqDZyfmdnrrLimzhypCKBNSlkE5d4pw3Ie3UNcOCAPVlnwi8Vf+XU/eLrtnhBM
UnV9xASexHVI6dVOZnjg0J0OmMC8h6NFMcuX8N45oNWwXw/ZoQ9hws0Jd/NCA/8kPW6Lo4ZxfIpd
1jBhMW3Z/Gl9FicXKj+Kr5ZSpzb7wkfZsNDKWwFSp+LMHuYGMs3IIph1L7OUphRRJTTKUscb2rwq
1t9/XS6N6sFgAzRUOYLfnxmV7RAKgNr2vBM905MThmod4LYa40ViBWPqxRcGQNjZ3Wig/bQ2aMMz
ilvNNjKXsvnIwAwGJGIswK7Z4u5bGHPfdm4ZKbDBuVba2dgiSUnidILIV74GDSdT9TRS3EC3YlL4
/dyur7vnphS+MZUJ7SCC3bkUJBPU0rOJCxrdp+bC/Tgr8ADaGPDc72RYs1V365FQgqgXSDaiJ49a
L12TUvnz1+kiUrfPpJRtn1b6+B9NkzLXjZn01+UySpyCg/H+vNjfRYbpvdzOYbCtIkm21482N/Ov
L3yRZTBNKFsdXB0CR5lwEZlOkkn49wcqSu0OYdwQHoEB7CED+36H1V/WY5xbSUQNRRdzAsWlKvyh
1EprK8AuQ/xr3NoyDZaEalNbPMiOW3F8CwA/AEDMleQoNL7c1gqLAY35pfc2fzjxxjxPvP283u43
PG8kONCKQm5I1MTO5gG2qz2/CblkCBiFylqZ0Oav+Lxppfhuyyct0+VaGc4VO0taUivtz6lMlT5H
06y54CS1//ZbhCaUu7qbzeP1FLvmiiZO95OhZ1nOvd3hQpy4nRCduOI8CQ9JsaaASr187iZ7Oqbl
eOyp+eoF/I/3QU6lAhTPxoGZEAiylOIewyrxtBVCQfd0Xv1e+6HYhF5wHtsCWZjsH5OaXbNlbzD1
OLjg5o8lEA4evt0GgT2HDPYYuLiJ2payGl+34VVx/nXyDpSqA4Q4lpMwjsR0oYQx/CGWlCtF+gA/
/ic/k22jEhn30rU7xUH5O5ih1lDfABAeHKSkKj7iXh7z75Xvv9HYOeLKPZvNQTRLaJ8qAMs6LVsQ
RM7JhCcxCZ77PTiq0IQAW2x5M0Fjn+ypkG+Pj4XW0eUxMu2im02O/Fh8yt4e0pc7KRpmM7ZYP2wY
135Nb+QNLwEaUqHgoghQOHtf6fKr+LqMncIsvGYqLIDjF/W9/2HwhzRRNooiHng+W9lHwqaIh5R2
sGSCDxvWtbZKsiGZajawP1sj8Fyn/1LMtKklelkWC0NetUR+zNBlP6AFexuZqb4VzEHaP52JebSe
e2mO5VemdqhYrJH5+ndjZ7dOwt1g0G9b9x2dS0zpxyFhUKnvrnoxn+m4YzD8w8f7wqF+w/L5n0yw
qo1TYfH8JRGTOC5ZOtlMPkC0UCX2tkgx7ZxZZQQijvTw8B1Qhv859rfAfKFMOPKIxH3kg4/HV/mn
hAoZ/EycJ0ufDglWtfVvjU8FehKuMsuLAYks2z1CCu6Dhb6uDMPR0DDs/EBbOlItI0Sh8mwDOQfw
RhECIar3CopGyqTBakzzgmBkkFv30OAKfLbGQEO9W5I6n+UjY81jZuXM6quM8RrHzSJ53Nhew72J
dmRNJFqbpwfil4EMnJatFedgSuEC3T1/Q8UswWZQTwXDQYE61hMqXSjyZRLnpGIriklzxusFRmKD
kTov1y1rK/szKFoMGjq5lgv4/R64oZuNUi1p9MzIKZ3PvYOf5tZ+2pHLCqTFyUOuqROKOsKHl4zd
LOjHOhFFjI10Ci7SbarWlKNRvntGZKKXThqoKkcpaGeIjOy4tFnKNc2lOzwlmM/v6FqVEVSo2RZw
tH18wf0vqzWWwyJbRFK4cIWGDEdysCzhUXX3Ti5lFvHk9pgXH4E7CJzk+balKz5olFnOwoNGkD5S
o4EnsxzCeD6mlBNYEAFb6PXs+2mwgVl+RWH/l4uj65xWqUVgW4YQVILs7a5v2tg8VY+WtkRy00U0
eraeTF77RYClFklWmxPRpsI/ETlhVLbC5Cc7i73kLHxT1omHjgbuCYTpFLULPlypKZ5tZPGM/0xH
7fwIZcTERQoozWJmprwRtkz7ex+ZiK6ZCDQkIMrAZ89fwb7BBEoFbN2CyDTwzPkPiRKrkorc+fEc
FXQCu9fMj738ijgKX5eB7AYiOglfeVynx7MzIMte0TdUWnv6ElsAwvIUI/h9ZlZT+QFut6fmRov+
M55v+kVIYwBWcGXPACprSCRxssQTl5nDIOwwkTJa7tCyHA6U1w1ir9kZNO+4Av73dONgMTLgktfQ
q/J7VmZ+q94Wwlied/UdyRPPjrzbn1A26nWUcz5CH6kuAvNx8AKxWbJBzSxWHL3+e8N+diU1b6wS
EcxfNCxGWLit1oP+chMJwsvlsbLN76kWlwqRaU7x/g4vude2Xp47qRpfY4ZOuNDSY7VyHesYvwJ8
Mrlp0DTf/wj1nwEuuBwU84fCUly2ouaIOqPI14968TnQfdenaLGVbrbI6eyXjnxuJA0o+HMLVJAi
cwlxbAxpKhpxtgm0LM6rIGnDjbwspcw+7wehm/HM1mq2MJn2h4yvHxriWFHAjFgnPr1j/7wLB505
IK+h7BGrCxuInvxFhNAD6E94ed30w9gHiyVySKJm6e1aOVy8XM9zK56LaAUTmUGAmc75LAb7k9cC
XFFOLTISh+uIMtaM47nfLBsvEnLoZBWrLFDwATf6E5K7u9VHr/L/i7Q2wd5CiTRvd4zgpQiiSls4
DYMN0LC9/474HtfGHdi+/QBQfWo+aOSFqcG9iU8nvvyCLdSFvGLPxCWbIkK5QGQjeNE4NG+dvKo6
C9hxJGDLX0U+8iUBQlgRoi/8oF+JZQCUvoJP7w+8ylHC/VdG/dAlFqG6/OWRYWn/RR1fRtlAQpdY
hkySvvBZ6AWopdR7JUFDVTRIU+Sme5GFxo8Y9RZbEkAILoIE7+4CBHfiaaPIIKBOhjf3Cj1WnbYr
c51y6aNIQjLDPRliHjwYsLrB+VXviEubIWrdk2q0zfsorUjns4S4b53BUX3QLG7e7TLUGQyqIojj
IKktg5qj1sKOmmSCL2ywr4xS1EzTeKmCP8OL+gFV22snVp+o2wHFaUpl2cQT70M7X92/KGwom71P
ZRnQWlw3whxlmEPgM7PL+TZY6rDPjuaYgw7koXLQbgoNiewS7/qM4BEo78HViiTXfTq06+jbuv6l
JBmE7nmbsD5jwkhXQND8aEuN+Wp+JTACHFv7LIqchVtwMbT/L5l8H5Mp+V1KcJw2124/43ebNnVi
HZPoxcQiwWLte6q+I5wUlqpv6tkCJ5TxGxyq+si40MN+tBAFdEhcYoIrY+7zb2GohETzATcRBfK+
W5WRIyecexmXFOJx0uaAc7EUG+VWrOcZVFgjm2eiKbaail92b6R5tKqvsAlUThJbz9+V9YP/cUe/
m5CYdkMrhoJoXkpXs1DBGUPXi36cIFaxMjNQsngHWsHlj72Cj4Xcz1nzsfXi6LaMmdVorg0Yv8Dj
w1F42R633rXblWKwSzHoNa8QPtJwj5CdKkPdt+ChgXf0I0jIgfJQCzcjOOA7/6mHqlBUCbqG095C
8/0uPLP0amuyDJy2vpGrRGmOcgwS2xSjifmcOs6mww6ba+2K86UZYsjPfVxRD1ENvTm3UzrVk8eU
bAWGzz/EsQIuIOayNoK0wNx/wktiUHDeBJ9CBlKjyGmYOL+TQMfoReNqpGpCqcWviyY17mu2ezIO
At45ezRohLNn9Kyg3iZ5VoYuAB8HRbpaKJmmZZdqbekleSu19P4Kk91G1/yJT18FFvSmPRHreBwk
6JktmPzCqvZdlD8mbaWdiuXjkzLyXlIFUmJaMtjyzshEg0iPXBfH1lTOMniJY5y51xzcQ4MKcKve
YxiF3XZlQV3q8Jpk7htXw++tP5daGeg3zz+StVZ9isSn8wu044asw6YVd6Tpv4NctZtwu7VIOvNv
WN4a4kxX1XT3t8MzFDhcTfC5ZQvonSPgw9aaNQ12qulB/2rZPMowqLPmDH/960dT5KhCSuAEFtJT
OyrZnooZ4W8jdqK+GSqIhY3WsSNHBNjQcuNbuXUbsyDiLdyYHmM04U2obPNlCY6taTI5YUKSUd29
+CsWL8TNhRoedkP+ZGSwyPh5jBNc/34PMZdUzfFlmMB/h9gZ0BA+U48H2bGS6bYNgHcFoecry3WB
r8KPEW03pJUCryb/ma+vqOfiyVls1iAJ7toKqH74WhQRHjESXwvTsU8+dnTcwNxdv9MOPz0YtSJf
Njx8pWa/fXPpj3VRnkjI61N7C0xgVNnuKFAhEaa07OvW4FHqnluYijHVyK4xR51Ut9XWrJ+LQaEm
sl1n7RYa2eV8MBbmc2prriMzm4bTfUyDFG7S9aNiho09fh+soY4XiRSvTbGi7hbFT9DxKLY1aEAA
bjpR0GXbIuY7Rt7YlZav3WgfI7Sx7/myVaMG8qQVFQU15lTE6yfwT9R9KE1QENH7ti5co3dIeJJI
BhGtwGSdzxFDMG6YCuCezIP06J+BpYRmPDWo1o86GDZ3ia9DbS4qVQ+r7QX0NCsC/NYhop69ByE2
YpRr3Wa9sdVuKJOlup81B3MmUU78EQqV7a/gKGVUwSGdzjjLUvFPax09o9UA73d6ZxRhyvPZ54hp
YyfiCsZaNffDah8vt/uEhbuUqUrzgnm9x26l/uMA2ppLYnwCEgobxrZ6EGsO3ixLZacPsX9kVOuR
ZQ0OPsYZzMA7nBcvS0Rk26qJ/+VsW8qADkC3oeAenA7I5rAAR91GiOKjpAp2nArXNET298lyx/Y1
lmMx192hkMe5DpS2VG7bIlJ9OA5vKUbVpL78tBj02A8+7SRe41nHn6Hww5TXjHEKOTiS+6x/7+cE
w9nL8Ia4VUU3HM/ncG6oXRfimyf1vA0ivIsnkCl6CZxIzU4tP+xVVnCxmi6CLduNTj6BNWTW8Xwx
XQk91MZnT6HuzCtaZMUtM03j1ct3gfYI71huCiOEy6MXDTmSKYHrANlo3iDCxUrHf2zvfso2ei9J
tYLKj3DL8rjChxUXqi3nMmxzvKZWvtkZRpAcF4Q6USZKOJolhUrN+acPs+os6PBP0leqsu6MNp39
7NZD0NWN71bp//i0lJsZRLgfiY/BuJbJ6VdXWSJkBB50ib9vQmyYDSygNaRKrQiLMjckqjeqMMGu
hepjGxoj4jFXmLE4WiZanXeCQ20EriRBYgpdHJlgEey91KvZL1VXV6i1MI2fC0deZFg/6Y0IC045
OWBpjQ8nAUo0LwUFeFMVRbYBQnABrnnCJh0/RzGedMzxhssEuJWMosS8Wjfpo2yn/2zVmAJ/2cup
urM+ZI8zRLTmbAxKoJJTAH6fosUpsA7Cun4XOV3nsMq481oqRU60iqVHGTqGCjSli4ndjv+pJG30
iLbSfDU/3KTA/l97MNo6ar1tAhlzN2pZch2Pe4BPGxLfb009wLDGRVWgoZqlD+QKH7R4ZkshXN4e
kp2TqmihvYT8751/XpEmr7jl+WjyXGpk4DG437QNMudOQkc0UURVMl9KOOlDJHCiNhZTisOqYO9Z
uANzNLQR1+SQGlfCNXNSYYEw0VVGi/egAPQJbJG6Xsi6yvo4XKklOlXC9wyzUzogUVs6WOEWYj4X
2amHkGSWB5oDlKz/LUjXNOpsDB/AY28dEswgnACRa/wkcCBdt5QzuOHCgCxHqMxF+4KQ7yWy/UO/
XuoAObLpgDvJoSaJu5cUDRMRoEWbZg8zHWJsLpxqE9rCCahxmzorjOH4F0swBtZIapZOOnAWVLI+
IDcYDxYKB6/bGbb3bzhPoK7JwWo/p5MsvsNLWaC5uHwRZnnDdVFS/a5k+2d3KNrferzMH4giisrx
OOI1EteNk3OfbukWkqMnVAvunChEHTQ/3B9tDVAT/u+RackN/BP38wY3bRZ3Znv3pQ7AouyFMhB+
uw35y2G5SEC1lQnoQfAVKzJbuq3srDTwkPH0m/oTkAu+Y9TV/yKXHMTUM9KSDZZRp0oqmjPzQR10
q1x8eAAtbGuExeJC4+hNVfgdq3jL1/LWFFSRyVEOoyvZkNbd/ceXBVtl4Lzk/Y5GrlAQmySofGIH
nYjDScDW3f2CcR04YfHBeAFUmmQWZE2ROQKYPx4mMam+EKvWKSvQYfWuLFdk2MrFjwRmq0Fv1fOy
DorCne2HbYn1c0Eu2G3Fok8E50NrLPgszW9qJ7q/4u0U/OYJw5D/G9QsVit7G0Rh+/z4SermS5JV
90KQ6PxijJfU9NQGOScgKsPuJUQ81Nj8K44e5ln0LGreuATqu5+XewMPpOfRbF8UQ90sly5QXQpj
h3Zw40DXUO+2QWLYzdDhDsl+AOG2Msqc0tXaSKWmfrpFnADhuWL9VhejBOCmN0LsxqC7Mrw+eR1Y
IGZYelDxa/D7f0hbD9XqZvZXeQcxVKQkIUka6Ai5FY3wog2tp+FWE+SJTFz9AjTSPbpUKDYqrRKW
2DpFfpvrvpmLkjqEn8YNDcqRlBXvE4wxSotQIwywUXJL3Yv7EjLc9fYVYIhFgzCH7V0GrqVgPYRI
XBw/c+7UCqTbxGcIMEPv9Gyn3x1XkAvLdIjHI7t5DMGwDKPLYfn4jt+qRzbqRz34ToMkP23iIpk3
rMXWoimx0wvlTzfSG4qPf4/kjCzIwl/FFICsciX/4XjGEGvuN2Y/IwDaqYu8IPGsXAmBbxBd1btJ
XeIYIwGkepd4ewuZwa9UN9+toSfGc0eXAWaK2hoMUUtfBQRRm8IERGEpAKPaQPfxO+Bp9qKw+xUx
Q481hCbZ12v/xDzYwHtBIlTgrOXMScPyG4I40lOC87t55dbnXJwzdUjCjyCNJFGCR2Np5g50PyMk
PiElTUIj4zCcN1P7gURGXyTeEFr3gXgFdn+fT11cMlI/PeI2wHISyeY9pfZG+x1xCJV8eJoyf0I3
vqoVPKIxzjE2c6u2W9wz7NlXuz5CI113Ip7/0obIcXflJl38oU1YgJMhagqk6zBIJEUGzYEI+m0D
268eWEEb67o/xsraRfVXjcnsCDhQlhdMiiZNCIBQ4hj1jergOE5jD2AFbUgVxxTMlRblcH5NaSOR
2rH4L4JFHWo7fhKMxCJ0yIiEuUWIXhdG7MyzHgSDbrcSiiiJ7FBgaOBw1OlEMYIOhi8omu72uklM
7GV975p9nZ1XVtP/X8aF15ZVF2P/NNRKHGjA3Vc0M5BnW40RX1pDvtApjxfSn5KUsCLVkrXj+BkM
WgQbfyZ4hWXrtm8MVUK9dfZarD9cNPMXYwywORbEso7RoqDrlDpdeNwmtuFNhtwZCnFBWYZTWfFo
N/JInqD5vlV56Sp6fMgRqdGgJ1LZo92DsJLVF/I9l727PNQP6HuIPVXD8TMgkKo1bKwQYqRjFDhw
m3zNWGYeC0xleqX0OdugBNk6Et2rbi0wJTkpd/ALzq+iJTyVtRRxqlfnksN30dbHgFW7Br3k+keM
hVGTHJfKMYgg/yjvDezvO+zTErVTHhHu1VUR888KGSAiH0HkBy9MUpG4uGmfT6axR19ulzqxv5BN
Ac952beejCKALgJWHI+yud/VmqP1MZXZof1xAAYjgvMFf2stCz/W5eSZPv88zwTrIAqp+rvywvC2
9FYRpYYGED3yso87U4adPv8EVZ6+iXa0aj0YL5ywwPIrtk6Wty4gGyPQ9/0fVuhj2h7zmTblq5j1
v9TfKm17AAC+miQp5eOoEYdz5bz+Zk8xj4nqUS/p2vzgdqY+XxfZ2X+4QERe0GThjrjHHGXtVgW/
Qpb/i4wBWRhWXJGfqpA+ZHyH3lmzt8Xa+2L1ZokNhoFa0S2O6DH1IA5Ok5Ue0Z8PfwW965TzHq9e
zB7AMUivBJhOr+6fC9u5pHtqYPuTDeKZvguxC29hra5O+sqeLkvs3S/iEVkfFxSCTy/hhXi3s0HW
fXxCoeTxsXKszVSxFdiUnT4qSYN0f4+/j2kTxvx1YCnsgWKnv6sp1+zQbkcMC19tcymLYTEn2iRk
hSLCqV5Pmft/wzDO0/L02h+Pe7VJojkSlgJQh7MYMN/WIGik/LRSwqwAldbi8y91Dx8q4Zcb3VHS
RCmty1wNqYtbHJPMRIW4NqKgeEgmNuRzM7ZVTe9oMKUF8LewMVhMTyCh8AweyDS+7U+3bFMSYOZS
MqvElxJsTgIHsQArxkI47z4MMmQNMxYMz1+ZIG1z6cNpv0dcSaPguDsvgM3bM2wZvYtaYyeMjjOc
WX643jQkM0Q5hYAeYYO53zoRFoVaW26DJphiQe3Rm/VOtTIr+5isHQgZa0m5h2Asu/dPhuowdON3
oneRWHZzVeMIWL/0PGRH4AxAzIH9BGLNTKqRKUkNyBPLtvOoPOHu1KkjNWbBdfyD/MdS8BPuy5N+
e3Bwyen48c076eQbWuiYJMjcs2KIE/tlM3OtnXXqR1uqnX8kwTI5uLCOpz03OS2cAojV8Is/cwJu
y6WGGwgNQ5sjDrsGZ/sf830GISQQ6E355ElRm5ckMpVEY8NKWIC+myXKnqZQcaLf0RkY/3tLRu9x
HNYBT1dDN+ef68ZryAihzPlnYfwaGP9LYr1noNDmK1gbJ6H3hGNRb6Avf6nkhAzo3FmlZTMVK7Bi
UMlzgjOCdz3KHvIf4kQmSFlquG68naqCLh0K6xt4BOEfG3Y0eFmNqmkPUVscHMdJ59e0ZXM7dDdc
QsSn7iXBqB6GgFlC0kTUoiTAD0DAUh9RasIEv7LkdipZFJsKqtNw0WQKGxKtR8yuG549p3KveGCj
iqTnjQqECf5UbKXc4FptnG3GeCHlEZk4EyC77UrbschWxXQd8RrFC2mD88LxOPr5LZxSh2kLzD+j
Kvh+DDiKumk6rIOR9OjYC+HmkxAOCuq2YTmTmEKfxKq37jTsd/FQfc7UKBWxEUCv22YiPxCeherr
tDBPOAgusAXgMy0dHQtv4jJNztMEaiLEbMfSi9Rae+H+2y0ADHK9bJaEmgeXKqZvfKo6LIjXzayB
c39RVVBJJntowPiQDp+gEJGdmH/WLeVvF8YhXg1bC3ffAyTYSxhCUHKHoarFQB9VD8Ou+VCq7CoR
WYCFUOvOV9aWLecweqAHN7uDAsTVK9NKu33157NleXDKn1pxEIwgyGHnTqlY8Iqykyllc7G82fm/
gg5X2c8NdkrjA+Bnf9zuDqdJyyWDQWUfr3Qc63Fg+owf9sIs/H0uw8Q9y0z4AdOasdXZIAEs/an8
hMJVDI4O/aYfMBx7aYN6HBvNWHbW+g50aAs5yb8wVW390mzDoCe9rOv1krY5a+gCw45czX7JL/+l
tnEB9foL/lKT0h8MbTCRJ3/XKjEZV7d6LRTuGn4lSESqSmQfm8Oq1qO8HbPbOO6BKqVYGT8DTfh4
PFxEQf1yelxhJBpkBOBgAeS5koY6r53PpCAfwiutHJmtA0uixp+I29VqxDwLBDN6A/T1sKPGPM/o
i0lsT0QHPqauWhPX8vzxDfaCKjZ/CZcDedAN0YJgmGmGNWy+QEvJtOw4Hh8plzkPHWN1B9CzHZQ/
Ia8pOCwjWro7KGlRHfx/y9vSGC/MKsSPyAU/errwRTKnnWKW+jL5mO1wlIcFk8j6EtlmAvjQFivn
Vzk2ZnIfRcGdajaBO5UR21NvQ6T4cIDz8pYoG/WkArVGp9YR2W0mtAMV95BjgjUl95OHRrMYc12y
3KSmWfW2JDIa37dE9xRTcAifJzAhneF9h5bB3SYSsklimkQDDa3zQ7CZvI8eFmDjaQ6h7516koF2
Ga/o93tkdCcHFgacNTWTxBsagw7aqFycgGdrkLpCLv2uM9f5qOS9lXMyws2rwNeywrS9XXCE9Dzd
hKWTFO1vKQdadLE364hB2NkBXXmgU+006vMZQFAuIm4j2LYlNIJpoLFlyAMsNFiKHLH3EMeTYnml
JO8EjTAZ0pt/2nw49xm7f8reoJD+gJ7aapNtmAI4eadaL/dh89CZCxsH70pn/tioRou3yVaCJjS1
umV9ZxyLPZrJbSVCoB1youL3tv31baV2z9eIk9yPfkcbPI91ONQBwaA5YuFFv2hbPwhGvHoK9nbN
7b5RHRYhNxmxu2oCygvcCqinRwBNJKbdwje/YgD1M1r/Wa2K5ekYqnzSdqd1wXcdxtcKC4B4VljV
+rIW8bM8Iy8yQ9YZWVgXRD6cYAF5yKq5joEOBbGLz4XO9qepjpXcvfRflVkIQGr+WC/PzA+kwqH9
+GnaxJKEcdBiJ1VbDyUrVN94qIGFVM2+xXRM4QmAB0vvQwH2aF6huz1aeNIYL2gX8JbDOCNnzArq
vw1HyqQCFetAdRvVJb/d4wjMWrWw5xIxKB9w1URf+zEljaZiOUazOXvBNIEX226CCBO1c06GSE2R
MVlDgPSgbGxnsR8ziteJIdaiBsyHBz6A0d5hnzFPV0/bxuBtdlVFh4FIlL73sPjYW5aebn592r4R
ffM9TEfNn/ESIBPoVjAeZmyra21BAM0kyExumynvyiUhGfrXUnRkjyZh6ClJPlcjLINCVzn09MXq
1n1eVd/jyTO59Shp63U1BMe2W304l519XjtGBzHJgeNvmvXUPpxbouC65QYwKeBHC+EE6o3zhMDQ
OEmg2UZrkkJ95k0QKSrX0ZYPVxpjJGFtsUrFM4oV7HZo+hsJAgecV5NLkUQt+pVElnmo+aHegRTh
nWMbgkPgshslLBV5yoxFso+716zw2ZBPSkQqnM6RKFkmr6Z7ww3m3jmat58F8ycOEAQ/6tDJfcp8
NHRw55tNaUcva+eDzY5b1EK7zhIhhDstBuTuUXyugBFoel9stp0QBhAdJdA4HZDcLUNlUzOvFg5R
DvaxTGAwfa4J6Xc7ySwgglD1thkxfuDQHpDER/wc0jzasvZgCf4yz2inATZcF0tu0O74V6ke2ZLz
m9Zwv3+7SQxpHZ1D0Kza2dVhZFdeR3jy48WDwZLP9RH2m/w165REQjqp8PeaZfr6o44BGZaZxRqQ
RK4BwJUwWKOxjSkup1gL3yFEsRisCeHia1Tc5w5ZyJWwpfyU7hIKm5gnwXuCzvLWPe5mAo76rQFO
iJgNrp8RkwHMTnB11RpkJoIEBdtHpWCKBs8zm/vFnLMV5zPF/VubaozipOUJqMSGds+ogbAsHlth
wmprbWXqtHAF72BQhX8uHuTH0Tm/YgH4E0shk4sbPxEEoKveBaj2jiAMavV7bJnMolfe6rnPQ4fq
K2/la8YxNX6D2ta59liiVZNiIKWaYeMDluyDWHs3VJJKNYUjuRQQFtYSgcpkBzydKqNKFRoIKqSk
0Jf7TxfIDIhCJJw49DJGVQ+lrNI4WjM0EhoNAcgQcpUNS2KOz7+gIjZZc458MXEFsMOCT7m8X6i2
+RwF+vNRHySY/ra1Zcg6WsMFrRKaS0/Nj+LAW0+sZ3aDt4KR3zAI2MxkmBDc5/dNzYG8SuU6QNBC
K6rJAkUCryKX45rqU5vr9Ehsb2x26zE2xknB6va2rXwwhN9gq6RNJ+7BU3IsTm6y6Y+aB35dqlMC
gg5ykQa7Bn72KRuOf7ETArS+6+9Rjx44+xUYkQaxlgh2qiwAhE//9lv/EIRdbnNfY60weKMlAhr3
4i06bTe7oIpgiKpdH7+otuwz5/40mC7mk6Dl+npq59pp5+pq1HAk/RTaP7F2Q2hUrLL1f6WPy6xL
prky/GmLj+Blvlvzc+hoCrn6pA7ZF4ErG/HN43hFEYT/6rN3q2wWCZ8M1V1CLXBte/O9iFVas9ae
K5+5XUwnn7onDtDoxH9XKpsW8KLSWSneI/BseduheOhXs7oEdpPS4T8LLUl9pK4Pt60VLekLyqzK
yrhY0bhu9yw+NclPXCODV03tktKOP9mWQqNm/Xd7G8OBzSnC5GxS3y4nkWc7M1CmX54bUhqVq9kb
+sMdaKmG1ZIZmCVFZq3MQvmhuYRpqFJ0bNpJxPtARg9zBSlW3Vo6YeYKX8lLhccxcNCJFOr8impC
JptfzId3YsmZNjWoMyHG3weGtu5ibRVdVUF3JPM5bDkpzv9fvArD2F4GyMRvBbAMevQ35wlbnWhQ
ESSofbXqqMXPBE8gGnQ3dzgvrWGQEo0Ab94HSLF0hYDPORi4Z8qcDow86djGvn0A5RFMLzseJPo6
wk79FigWvbZjbBAS1FeTTgeumt2+8iJMeVpIqw6m98fEynau1cP9ZMjqxnwfhZGCH/tMc+DhNn1b
l4VgRkclPA8lWBMLkBtHSVGCrSS9FHlPspKKnW3UQ4CuBR4vF68BD+9ju+K+eHpkigVTO6Pk2+eO
sOXIikf7fuNrxLyHaD2UrrmZtihzNp1szCvZA8eGieH7WdVI4i3EfLP++Qg6MLradP5WfXfS1bPs
O71wBt5zn5ziwmX+BIEzbhEcWJHw26eWAVJQVogehX8RYs0tsdAFr+JTdZLeanIY88onXIsqqLma
vRoCSqtFgR5w0yfJeqFcSFaaYyFOeJ5DcMhE3Kc/DLYspkFj1yq2Xj4LNf0cIZNgjRx4DY5IhWb6
oNPml8e9l/GDmpTuQGJvQJL8FyX7SKBx2ljFleqPoY2sf8EE/Ys2V4rm4sReWKsmuw6E8T9yyLTU
N3PRdJ4tlWYhdUgVvoyx9oSYDgBE403X0cCw8VqDtDVKE76LbF03ZIk8WJjw5Gr1pNBHRIRZHLhr
s6Xw69ahPdwk9P2OH5aVzLcZIh3SlKJ9k76Nsk44awcRjPg+iC+SXG8XIW3rbWaUs65PVpCAEEq9
xdWvQaaGrZQItTpcH4cFGBwXaYyXG9Xgr7XegSkNpBmwWXE+n+K+UtIgazE8uKPEUE9RrQlUr9lR
pcRLNLNGBXXe7O63cLqMZmPKOdYgJSnK4TbiqNpVXWU1OQSKkjIRqmiO8yzL7Zj3qmQS8ucm4Xff
F+lrM+tK9nXvbg5SR3iTs+fzxUONdLxWGV1sp74DOECLgmuJMjv5arrmj1rAU/9G4aWEfXuwRxA5
lF0++Y5mmIZArHr2h97XhfMPX39YDgKGplJXmeKPYAwSU+3Vgh3/tMUj3wBlmcg+136eT3eAhc8N
STpGthl/NjevqPR+tSSqZnd9dzYqdLUkeyawC/fL2eO7GeesC+8n54s6E+k29jigTzynfwhaw8bl
GFFQ8uFsgPk2DFoLeiuSQoxJPcRqk9sKEFC7Zos0IGViKMFjnyKmrdmQaSZ16J3wdBiwn02vNhB0
eAPNnkydmqzW439Jl7AoY5xFs5v07idJr1oDqfmCdDFU2KrpmX/xm4fKmIdkgixNtutON+v3n4L7
KOdvfSte1B31Dj3zMA24bAFGHrtX4yHk1UlzE3Hbvw4DAcW93KufmSkcx4Ho9B8RjngL3Kpdrw/W
JemliGREgoJe2sorQ7RZQmvQpxtm95P+jfTHVQs4Ke+w5OTyIQR5iP+HPyCd6+sCWpXBu1sZwRUb
090cNo2QwGjaVgbxV4WtIINAT1Zeb7LvDFbE1Ehi27uNhbFdr6lR8bww5XhG5+9ZKPRoivvMtkmO
Kq85k21+b0mbYKWrFFwo9uPUdN/qb083UZu3YfCur/Kzt3CyrNbSefJXTUMsLQZ1a4CXM4l1WNCf
njK8CrITInGNN+wKze+fD374G/EjZosdZlOxDVxOSCbKcQFkyc4/DuNi1Owijm728avCSk/7TB12
C/Q1817OuolE6cLisX0Mh3ggrG8d53JO6EZBKX/1EXfEavzLjnj2Cx5U0aVCfBTgekOa4J4kkiqo
Ofq919nPdMrhGUba1CfC4dqnIW6CysZOGhe2iCGG7hFMCv0BxzL5mD0puKxlrs+qu8sfsyi5o7CW
0VMXkiKvCLBs9HpxzMECvZ1PiXbQWAsK3FCLxHrj2Q4BhvqqINq+yKP3T1+dI2WORMV49qWNX/92
DPrj5FF0UOwItPTznxVDxivp3xknkW54+K9+lh9hMBrzb9KffFttyAoK+U4xSKhajS7UZnRLU6fy
i0db5sjXJDWLlBJVwypF9qenkjSB/WNJrhhT8xzo5pzB3oa8Eev7usM9kj6oJfSWdrLW2xTXaDLz
aOvFukV0nFkLrI2jXS3HExyiqTAI4HjYAE782WylSAKWKkJmyDCEerGSst8VMmVVs+bYrT3DPMaa
PPa0+fNIgvrB3uf2smloGG/Jhl9+prJNCYmP+mdNlA476FEPQ4O2SRYvwZZu1laEZTNQmmW89H76
+eUUJK4xbP4q34zE5zWXpR6eLtDaJnjOXcRDXF6Xt4HNWuhnjDF6oWjx+w3IZn2wrn96EyhY9X6o
/rpxGQju2kKHet7gh+nwL4W5RACKTxdPBQzfZqh/y83BraV214bdmz88G7h9APUDXZDx0DSd88o7
FhHy9mtWQQ3M7X1MlCL7vDVhlKS8X9r0yN2UQ72IIuVeLC5mcSZ9t+Mp9a/FioylXclwWdr3CUHa
mcqRCNFGpWDE6LQIkWxsIbmguyxttbHxZ7aqtcrplogjAV4uTrryjkW2Qvb7mugQ1mYH/qX8SACk
RjR9Is8AE3QrYI1kDqrh3M9iuyiOKGLe21dYtLH24kBUyktu9B5mZ+psC3B56S44fXHgS5GCjRnl
0vMvLex1urXMks6/y7KG4AmWjzd7L4kcg8vgK/fuCEKufwdX1KJJvuTnWyG2KaNIgoCn8PR8js2C
YaG/EmIXyf06sfbqsgn2Op1FnfTQ5gCoMSXQN+4IOSZQiVq9UH5zg2q/AcWpNRb7F6RP8v40Vmt0
mbtP8ubdrBvCKyUgPqwVJxKgrjo0BONeDS59Os2r+J6ktLg0+NxTnZvInMmOIH7pamZ1pgOmmBTU
pYTZ6KeqD6PBNZXyY0kuAcTq4UJjVIz5ohB1ddfm8wTIuNq5r9qRNOasePIJCQFX3VnwJ+Ux0pXR
lbtwmvPllmvr8nZ34tSA4thx9wtW6BJiZnR6aW19hnpq9EXcvDy3fED8eQb9vzi+jOLKrrgB7QSF
brmvyU/uRerfaUKwszAnSn6rfJybT9du63vE+2msAXDq//UoZ6BKiYDpCux4srWSjOzBtWBHxrTl
NpvGqkByzTm9ODMJbqHmxuyq70+jikEcsbJ2u7h/iPGWdgjaDX+zdXLifP1u7fv3VfsPLakutO85
Utwv1Xwi3AZ14T/UAsPI8aRj3Zi58IFzs1OM+PD2XPpv6kP+D4gTcKbG//n21ntSGR56RpSIY5ZN
BIHZPP7a2cQQxAoVMsg0GY4KDVR/EZq4+6EvogRNpr9iRt+KTQvGfC0a6yf5Q1gXSqofcspV2LCT
WNRPGu7KYNH9FxMgETvJQly9UWVxYDuh2w6Z04B/Bh3FjnlGICQBjb+2mbfy/nEf/RjLCos+Oa9x
y4qCvmhvaCM1fK/zbxzkN1d+jIEW0mT8SYhoJDB8PEBa5uNk0AcZoE5lWYJnn/L2RCSy/GqvDfOV
AF0Db8y6lF13OWzML6T5u7m1V8iWMM8mVfa6FGyM6HDng7UMEUUcFcxH5IyYQ2J/l4m4k2vQXm3S
i2RZ7TGcG5YIOsKgkVuz3DxbbeFxIpN5mu1qlql80tGdUNG5dpBNzkdwBGVxDPSyXkCiFOu9a4Aq
saYLhPs6zq/YcGz1tdyqVQVSTULQm2imrhI6KARBfmJsHEpiMz0efnL8mRqj4KZKjvwgs8+53SUt
mhYC3dNnDmicro/iEOluoEfZb5OUoYX08/meTBUgytw8OWRpqeuHH+OvIAMLdbTiqUMxgv22rldp
YB+zNcybKojvrzEkKoL3rCZrQBXzPA+TuVv+rt0FfH7qCy5Ci2Vd+zN2Pl2hPobt6lAnxuKsYYMX
k5kct2HdWORMDOCXUH7FCd0OoVSqegIoNIBtpcVlHjKTbr6e2/OST405lkOoX6WLiJzuSaoqRUyc
isUB+zNbb8U5n21L/jZJJfNht0YnCL7pi5UtxodLGCt0BYGsdvuVUj60TTw1iV2l8mFWd18jwRWw
/rHz1lrAey5qD6EjA4C6fqEBJbSm4wQxq7bPWroF09euWyUAw4GsIGsOwADtKzi0Y8twqO8StRz6
AK0CZ3d2INHdNmesvUjSHUzjiqTkbPMDV48c0w/QS/TL1mUWPExeZy5IUPwE8tN1khLcog8xh93O
/KrMFr36JRFqrQYEMRLnnN4zQFK5A3a37Uverie923GEy4lNqbdJ/p7yFY3hykp2T1JIJQMKqmcj
vfQjfaemasl5zVABYSqqtDK77vgdnV1UXs3FVWl017awVzweQWGXTgLzs7/v1qHkDa7d5Dghhiei
H/GXDQs44XtEjlxBqUG51dw7KJDt5OHqQOoh3bnEl/tsY2QZhO3HA3llb2kTkO3FQVNJYpDaf/rF
avuQ4qsJ9EPLBiRG7U5xtF/UnB7kYyu6LDPre+3GYQMQQLYVv90PRyrFl1RSKEp2dcvIYrIfggEm
AMXxW8/GDDNsIgTL1z9mgenMI4/iOBBsNJ3jFG+KtYLfmedijye0eyPiOnZnqO0bxwFswoZchURZ
tBsQBufJqM361M6YmDC3zZYw1hdzD0+0WTNzJwK1LMraCSdKSDZuWATSbZeFgt9jMpkxbocCAFJj
kQEI8+uLOscM9mERbjGepXCg+hEARl4f1pi/V7H9WyiCCmctuT5Zlvzi0Q8hmQlCKjp5smEt3bsf
w/Mnd7wTtk2f6UGaNBgjXnsY6WXBNXpO1mrBxZzIiZnYKLGCqjmunzn4Od926bVrRqxUnglew2Lx
eNI8GcCRztH1IDXNbH52S5CsqEL06SO9BHh1Ztmk31Axe/zSek9POWH6MIs3datuGqN5/djRqFrj
d3SB0r2k7HkuIePGmEHvCLjXE/1hRRBx09Xg87wDzwzNQevA96gY5vn1ybjNwfWqWCgxZ6mm+wDa
NGB330Rt71q1dhMw45VmNvHWlTzf3oxhZRBmgHHS1Z+CnLLJUxlvUXkaJ9IKvGU/BpMX3jDx9+va
iynhgsc0s6F83rI6c9c4xa/MUq9T9QJ+mytQ9evcIm0Ft+1jYmMIG3TNmtB0pl9Krp7rU2rTdu9A
ORPlA3SLDsSYyO7WREUtIhx3Rx1zGsRewf+UuK4wesLzKf4h6UZbEjkqsYtsr6zd0Umv5HDzEvKK
ojoxy0rjSYamumFvZWWdODmy3VnbpghBLqN6IsAFTnpaxkfx1wnV/EPcyMF1jIBhyXXAtBRllKPr
JZclPOeeAXdbkEe6aY3/JJ5VId9pipIYqk4d3S317lw0t/X/ZXoE4Ocp7gFldXN4nF6jR4fveV6b
xsWI67ApzDoLRvx/vZsmY6SN9cflky5TDrtEZ7HMcy7sC47RrzrsUQjdekugVBwfDzxMytDPfkVg
kliia9fRBdbQFshuZpy0DPVm44SEVZV0JBY1JxVQKyxGWs7S56c0gKAnjkBgQbDnKr/kddRPuRaH
ON7DyaTZMnCteOyL20wabGrCaXvxcZ6YuTW0tuprLsl2FQsGa/xPVHt4oH/ehnebtVp1aJaAKCdG
izAevA/+E2vKKDPSd5Ks++AkFkRYF5LhBHyMLqzte22CAkJvyCU5mnwh91hwdFlq3Ldc94QHoIKA
B4ccqs5/KDOkPyeQHs+oLogHwOw30TauVBS9tDnaumPeDY5Plear+FyzLGjb8cmuT5ZrJFkAKz8N
pM3YSKGepNWHDbdyrgg47x7d3a+9EBBjKIB4lux9hDA2sS9i/QKQI1vVZ/W3HJHo9t4Vl7ZqGdkA
XfSC4wPUnwfseVDYV+TUjAn61nvOTajZ3uSzQK7ajDhLgIUt8Rqn4TqvmvBJmOo1orsFcMpoaEL2
P43wp0hbqumEjhUss7nZwtNqCRvca3PfuNhPMSic7urw5jkElKByp1wDjdPyk9+ZHiKjRz/3Wu5M
gQTdU/ZBdj6ZtXWo1cAkf2hDoHNzZPB41XlTk6Taum8aMe4IkVIveoYAv5AuiAbmkyKmjQB6YxSW
+bMYhmedaLgBahk7M9X0xJEVJn7J0LndqTQDTiTn6EPi4ilWiUKP75MwYILYKfdIp/3ofKpklGVd
9AbXtZjSI7ejOGIn0k17jBQJWcVKRdVKg/QvECy3FhpXJ0gXLcfSH+Ixwx1VGtKhMMnBdl70gvVL
/vKPWnIzayn2X/eVGLyOj4CCMK+cGQiYqzVwPo3yX8pHi3QO7WUngGsImJq7Xo1eeD6lGgbhHsd6
EazJO11b+3stffefHG8hxoCoD0hXRWrsbf9QglplFAi+nlxhc/UiifDpLHTAOD8gfMbWcbbKX8bc
0SuXUiorFmpxlJX1hlpB892ECXtdD5QHtzE+zGTOWmeSe1f6Qush1Kwel9WLzmPbaXzPtprkGt64
g08oBcDVb+bxMdE5v/pS6bz+kIhbmYCunVZDEh3lRCFCFeL8E3abr1lpqY9MA+JrEEn9jii5ycEI
nwLbkOEFAN9cOAlqaDKs5ENMEw4fWyfirbXyPgo/Z1o5HR05rqGyh7kCae3LpktUnGrF8L/FuOvG
9yftn827gdhdW70vTRqtvpVpQBVQLR8yZ8MSV7d3peIw920FFvsxGHoQZ3fMprcT03txMlXnWI0R
MQtHK572Yky1PtCgKhOyl4Xli6MnvDRlXeMMfesrxkoxAxQrHGIv5Y0/I/mS0lt55EWMtDvCBdvI
v9d+jjF4mE+9J8iljjpI0Lt7MaWUiTzJ5LQTA0FSzaTXIhCKp4HQ76MtKUEU6WdXD7qCwcAHpLWI
S3Jldb+qKstSmDikWdV397hUD31h52ERkRDfnz93NUK/t1DOtyJf2AOLEK7PBxtEWVm3NW3eh3O3
VAQBCZ5Ql/Z/H567wIVxOcQQgA7LuDd/0ojiJqEArKk3uyJTjTVhfakinDOvxJrd2egxQ8ZpBucT
P+IK8OENUP5MTWL8EJEmXUiNIWeWsHRYSSgkRzVETzIdNTXavehsdEbTJBvH8lHabM4dJ0DRrt4o
t2o8kFPydUMShClrLtnIueIc9enXlezdYJmiC7FANpnD9OuR4pR7YDPRDHcAk+Hgow6dkps5Bybv
67Wg3y50pXAJGfQRigDTdmMaZlhEoRfhpZj4Stm2YJ2FM0rc/NcNdhbBryDR9Sbl8c58d5tQVMR+
miOHB4sUkxFoVXxW4U7BAuvDeVk9ouzvHNLHTk/jYo2V1dpLSgpry3zlUsiaShRiLTWBjspIHNL9
PD/1MMoYDdRxzm+5aJ7v751XYwDBGmNN2xsmGuXIHXO2fMNX8e0+PgZynAMPFHbdBGaDwjG8/MUD
ClIQxf4LFR1hJjqyawzWD7rU4z4D9YJsOGXllR4U+AXlqqrjQ1pwkxlVfUtDS4GBD+/i26Jf22tB
1pO3tislECp2Bvvai1iRL9BXohxDzU/Asmaed/DdjR6VdBsvtRB6TAfVNJmO0A4JO8kH0O4VVEj+
GL9M055w091amAHci1Z5YlPa8/kiYdNI9glwiObondH8Cb2hNQa4m2Dcik7ZCjrFUwVbUQ0YZiw4
ZFsumXN0sMXGLurZui4XWoDVc2Vuer1wKpgVy3lPOEkvVpibjJwBAuaYNNee2KdGkGp/qJ/pXFO4
cVGjaV+6dQXOzvuEyOjZGw9oEesKkkg2Y2JEi+MJ6Sbca7V+CLoFt0Ne15LD6XJAkEm76P/zg8Om
bbHUgngBaXF3biqYhkHkfkPmSH/AUQd86vS2sl+2O6AL+H5+lb6BwqERS9ax+kuzh0Tn/6v3EW2I
KqiLsnzxMK+XMzVCOudQowuXoYklyhSy2JLyooAOQNHJaOpE9C7IRX+cKS2FIzpyLde10TIUNXJy
UM8NanqPbWN/hcp34rROSKnt7/ZvHVfOEGT8tUMfMkEXI9zZnAnIVByIrBs9te6ebBx6zfqARvuh
U53MFtuIapWU4+I0pkJAeBSJSgFRN1UDHURzEt5U9GfOiO3NmxlPSsd9KkrzvID2uKExcmL9gxFO
5kpKCoJwFdOw7beS4fq4b2n3wSfnkvFinaN5GyDIycdfi+/zRkVnhSBXTk15a1D6kA1A5owGsnXU
zcP5qHZvrpxECEUzrmZpp4O5fvJEqhtQ3BXyGHz1fNNJjVIotfRVLobi5TikcjK+NmtHnWFp+zMj
VcjZStiOOR9IfU+Rs+sOUp9fPCV2F7/012NQ1Bli107LXjhLCNpDA/ReYx7Zj6y2F61E1QFP92cR
FNxR9DOER8Cvnp34lOfboI2nTQw/bqJ04G/6lzBIsPnW1tqI4hsNsm+xzcqJwNSZhSEgPocfylFw
MWfd+MiwjJEuKvw0NOtPuERJbWyvaTjlXyMtfDjmmJPWwBoc9zGLSRixEdC/ij1SBWKRLCI6paLZ
93JYASzbbUUobS/pBXam+/OyL1e65LjQ9xTV6tQVvCb82yzFN4qn6a6vt+DNffrf51bs29YLEG3i
eJNuCtVRMlMckpgAM0QvuF0fCCA//euVUtTgrcJCPsLXrtEZQsZIbYjxuSJXI5L54+7lwkFaA7qW
ErqFxcyuudqbOY8iNamkuM75o6N3ocjQHDeyuD23oblmtGn3CfskoerPdZUS9j3uw24aR7a1tQcY
JVOMy/Sr930nzLiCfZglVebCSLrE1zP+8rcJ5dLa8Hv1ZyMS+nbTYkC08uaWubgOEgtyUqk5Fmvy
ZEJxdb796QF7UfqS1ukPxq+wLUYkez5YzRZRrIFZMq58T1qeAX29lOOJOVpnxsEF9hclFOPqmAN4
6MXrlliIE2GIfPZ9wKcyH0fnyhYpGXIlITn0vgLC1JmCSFnuUA7EWHXS545/95vbCVYKazsKWfNy
/jrvRFOaPyrUg/J0tlUsOrt3GH8eQr9KZ27khDcAjGkWcpuuG1esMaZVTsApZpHXlfO1FQSVlaHb
sl9K6YpiWWFc9Tp8dFA94Vgxcvny0CsWG5AUgoilTntnuuxOgO6w7YWc/54b14aHk6Pc4ons66MJ
+gikzrhdHvW9EHC5NH1edc2HkabAi/hDxpovRGHRbUMSiOLJC2JKzmNNvxQjDEit+eFmmEhXd6j9
cypy3U9FhOU1hPK58qZ4Jaead9MYa3JNRbGh4qB/wMc7Q+R7Nj6lzIJgwDZFUz4e/DgFncVPPYjz
M1TuMiGBQOCtZK11lqSxP3Y/WQU7bqqhwJAGokEIFkaIZaGuJQ5DtA0LPQzbDd1H0fX71BIp4EFl
+cCT1qjzpaVciZhREcDIeJEFz3514g3j9x9s5fMhrui1tKr2WQ/15uplgcQ2JYONwtjjb23bkqHQ
ynQ1FQ2GmzrlzUQ4xWuFcfKEG8zi6TwU8YwMbTZnIJNqDRWGKfr+4lamP5s5AuiARdAezMAy1Ft6
cq3QOV+KKNxcLAINrX0aE6jX414AP1vBPWcCsuDu4eDBOQWGc1Un5hL3k1IHTuxdLuIxFkX/A7YB
bC6rO/xWcZk/GMXEMxz072jY0rwq/1i3DOBmECAAoDdgr/NyIOL+X13qxPGEGf2/9usqDL+G8bhp
fds+hZH2Ibgunltgpq79naknHsINwvXlWRR2ZCqFKlUCO8WSyCGxfA6CPuH9DzRCaHMB5OQ8z5tN
a9Zkj17LSjV7z7MHpkAZFEKnFIQW1JVK57JpBe4sS/E79/1EGO9mhkDYw2A19/6qq2sV72pAnIhl
Ha82ZcM1JuETKWOv9ZBVpVEeweIFL0R1e6FbBtBE5bzHOHuAl15W+JUkEocA6yskvs1j8EGU1K7u
s8D/lWGeqHd+2MhTb4uMGpAsJ1LirG2WJaab6Tf0fEFGFJrtghekChbuxR+WCprj09k7q9EtkgQD
zlWW+g6N6QgqA5fAA+PpHgyzH9auXcd2Ay57jF99whZ9I3VJ6fdSh3/ErsLmSY/tb59BInTTfNly
wYJ3Km822eOSe5X8/3MYOAdTJO5hnm4fTvoZ71EkD81kOWKnNtdOn+sVxBiYWRpiw7g/sK77Kmz0
rL2+pQJMIf0r9M8kc9npbZUYLDIvvcNmwnqjsb2Zd9YcxEgvMY64cY7aQ5rT4VaxFumaMroZF/ts
2SiKw2X/6urW3QsZDFDi42fen+R1rWl+AeRID2yq8W7+9zPUtFvlMpAfd4bj/YhsU7I1RgrhFr1y
ggPZtnlx7lRTL5aL5L+KC0Gc20JGUzqGuBOlBBdEnPOrzJ6iW4UiLFM1XvfF6gQgVgV7wMhZGx9x
vGz9RFDsMr51OT2o4I8rxlULuUtntMO4sOrlbhN1ht+1NcRNFuJpWpeCrG7cL4JZnoqrh8GAGyzo
H2JSIsezw7uYPR3pgcZxhl0YMeBW4yM+jIIFNbg8TDQ+EGtudjr+XxQS4uBTESG0IYCqw9CRRva/
oxt1dae58MIEmGrrgrMCXd4FLaJA0DA8QyU0Rc8dWhrUCk4GTRaPa3C2e7cGuR6IBSSENtXiDxaW
ZmAmnTY3WTtQ2JCU0r9FOcJRIDD4CYekSFffmnp2/p8JiJvUNF9M5IdybaMeL+jahSrU/RyIvf4Y
fklapsRnPa/RRpvF801i/h1RzRlAHmaMbjKuH4vi2AF+/a3ZgDzz88BsdtsLzI6ZvLJA2qokrM3v
RwVaW1ag63YaQXhJt+AZb7ytOf787jAOWRiBAE7gyLhryttplo1Yk6WdDDacmTSZnrDmRy13dXpN
vGR68EijYeyNTmo9PWno85CYSTT8TCGQdDxs1IhzmOoyUMd3tzDhYeqTetylPPLt+571pFL05EPS
sTWdJJ7mZ8gz3wTfMrsylwRMgloqx7AUpmo8mNCKm1sUw/cx8urhcapXkdF/WTveXB0Mm6/FI8Cn
m9Lql+L3pR3POLvpVp+hMtnFPVux+CcEgpbOhxjZTZHtSsajbvYedP2sfZ5hZpI7ukmFIIASdQRS
0otjBra56wgujREAPqUHHnY96Of+jYKKs9WYswapUSO+QTnFs1wQ9IQFvEk7soSEHddr09mOGd7y
f/UhZ255GHmdj9RolRbZz4fxLEtIrG2SOjt1OEqTF4iFMOe1NBH1kqabBV9MsWZXaOekMFnKHoGS
T8A60Ldn9IrqHFDMY7QOwkUG7WWqQhu5pe1PLYoewM0P5i/siU+PYWXbHM9+eV3Oq2h/DXhuFnQO
N4mVgkgkLLsBFuy5FPppIzFQqNFTFBEPagMyU1MRdclongjYJPfq1g/6LmIDv+Gb+ZUztyzU1Xir
2Sm311GPHxH7EuKQrh3ykLF8wXDFovmqvOpos0OHA/WVCNoHDG6OUA5YguliHs1WQ6eSGyxh1jDz
gjn4AdpCLoPeFS1wqRQBxHjowqaVIjEr6V57ccj0NeWEF6nRmytNCaAEPtsWf7OwMHggVMdYygHC
/tu2mKdKGqk7ISj8TBKiCt9ocf57gMJyRoRn3nuaVZRyEgEa1G6H9OsU9OIGh+Hn+mwK0Nuev7r0
cBCufZOI5Dq5Txtm8KW16hug/CxA9n+s490jis+J10S6yY5DcNimZTzw2vgQf7g+kXuISA+XrHNy
4qF6/BRcxpNrne2u6ZGbGG2Kw0NhtHG287t5N1CfVz7NwUo0mUVh60kGzm6f1YfTsfPoa8U5R3az
VoC7+lpOBdqTGlZMyNrOlPZPKIW9dszmVyIlFIrWhZzv+1lgOrrGV19oJVxMV7otvzINp8xdK1rv
Akcvlc15nbLXD14uI2h+frVWRDz8zBo6LbTqWDPnlWyjcgVzHvH6SQJe5EUSWAcLO8vnPZ6OzgH3
MoennVNsmd+dTBpvyC2Pw9HGEQTCySopaCo8fKhfdV5xQ0yXUlz8OeB9BBrGV17S+zpsZ41R6tmv
SktrpcpxQNeClJEtQC0b+H4x2WyWdBUVQr811U+48RTnlgvGDEFIE8KBydVKVQuiM22QWDm6R5+E
OdGFGmyB8+EE5pSWekH4bRfO3OrASs1YwnOS8U0Dqhc8IBteyJg3rY44AXC8l4IfQJq4OLxb0EKL
fauRE4M4TvAVZxMw4yYqDSh6mH9hkTzpkB+2Ub0lv5oL7HFWpYqnIV8RUrt2idlLYwCiE4Gsm4iQ
Md+D//MUSrPfusx4QPr97aV9Aulx3VchmZxyg5asQdD92diqDVoicTTTBoN//ip4FrmGgIHzUQGc
ORTa0uozSFDBKFsva9WPK78OroEjQ6n94PgaJwEPjBAQrasgzJ4sQ7MCBbrYfbJAfCTLhQV/EIEk
wGv8PzsJY1Fqo11k38+MNmIy7RZxexqew0+bgjpAOKnxj3k+3jsItLDP3PUCMnYB5ZyiS6NFYYDw
xkBLQ5PwmTI9SU37Fl/ERZ0lcw86jH37+CxB4FGU3TYILpCjFwXGJrH8oGWlebKNPWhA/g6sIOQ6
xeZFFPlefiJIeCncvTBqdNgVFec5zrMLiEHXn1pIyMiBeHA/nMokKfc292siw2g7UqnSIlcX/jJM
jaRsUsIKMYA3pvH/jEBYbIctRy19lZfm5Ks+EdZuiMx0kyZrT8PYtaTRW3B+szjJOf/KXJzDkxM8
lZ6wQd1cRyOXr7oQ/IMvfWP3Id+8pvcDAfYlsNq6Xwk1WQ+XATNJHIAMkXNnI0O5hXAKwXfUJjfh
LviOgSQLmEWQjVzaYPV8WfVYuxn2c33GGfb0bNXtYojYTmRnq2n8J/eoYNbHaVTWC52SZTp+4pte
hpvEwe2eIjPbmm6zA7N2WbsIzL7GCGuCUbDCiS+aViEMnhexD9AvA60acp91XsPSaKNLF/qOmJiY
4EllBOGQQS3JkRM9FNnJrY7qJr+UTzqJob3WZWTv7+Z9nSgN/c7m59+dpMBovtm5kRjUMtma6unN
MgH6S9fHsXcwQbnjqqMrC4juhr4TAmY8zW7SYYRKd8/CmyXx/hJOy5sTZH6g9UzzTAkz/siFCn4g
oMX4GX1R8lEf2mm22z1nyk1gqhF9uAno8Qwk5do5vY3KKOSDNjuN170Feq4bHJfYIN9s6nsIgCM3
xjOajRMzKXsm7hCA4G1hPgr+5DUXFufbfWXF5BIUdScEi4rZ8MmzFOMXifYAG1tqzB74NPnIgP8r
ufUsFgk8gDvh6a8K+mAEqf+EyOSzi3qec9qZyIx0E0h5WvmsQMNlT2QL9sVKZv/4BbFqT4YhgXOc
vvUsjkiByPxKpg7nvANbeDjQJphWDrCZFMEFpXac4rAfJ8dklNcb/1muYi5wLPRJvg7eQmzPZaMS
/36BK2XvXstp/fiNWSVFY7EQS9he+gKSw4p8BVKcKdOK8xiK1TBzY/5paIr9+VmBi/ckhpxdbPru
11kV9jNgdVAU0Jkrg0w8dap1tOycg6p2aPS3Af+TRbqm3u71fsoS5w5goXwiqsjvB4YtpHU3qzQm
+RM1jnJ6ahSWQ+xITjvUgg9FVYWnMwPuMCijkPWcdGS9mZ7ZzfbbBcpUQwxEtocWoOic+QXljHN6
AQw52f6Ex9tGXQ4JPMzcGbetp5fhzMmc+YrJdsHP9gxHAHQ5dRx0PqsZvSp0PdQ8U7ROV/P67OBp
gsbhxkwBW5fkSw9GuBFup3FOsf2uhLsDbuDJK5Iat7DTG0uqJcORWsk0HLFos8MwuO0NdS3TcO8D
YUEOIWW7veI1Qz3/I84poE4K1UVIgmmA+73mOxTwDxIetAeXvLzSYJ7JlENfPEnzI3+C3GCHpM9a
wqO/nCLCp04Qeezuf5VkXSs3KLtUXTnEwuIVgXZ/VhqzTe2+gVU6mmXZFyqxFwt2GzrHfiFoEbLl
EIhBT4KHLZ/OBLDWUcBtgzkPALYnFKcHmfhJhmrmZrWYnnZw5yjWVgvj5k2ZFof+2komhIxfahd+
TpxDy6XgiFeOwWuLFJDNg2Ev8Sg1taQtE7uU6kGPbrt4FPpll+D2u1Geu+GuUHGWFX/g0JhYIean
ZS62q8R/5bZucaPBFASS/BN6SwUQfV0v0tvx7EjQyVNns2If2TZqhinoDSuP7HrXtvR+wjVGbi6Y
SqHkcxlizufHl24n/pBXXAC76WuqX8IrdpKxIgXjVCpRZt7y4n3/T03dNc55vl5Ln7Ro5jHMsSyr
2GTenrzmaLNr4KThq/wwMFWKXaHHG7CNE/WKQ2/Utc5lcXLO9A63qXkiHp23A7zgVqPi6nKLdmP1
hiSbx5fVoLZLMN6iMxdkAC3CR3Gfvioa9mOK3fQqvvtthrSDvFS3Mtlw8nx5r0Y+lULu+i8TkBfX
k6YsYXLyeIAhFyRbQq3eHoNmgjTIanOYsyN0L2SX8cSQWwPLR8Ee7uWV7unk4+t9LCaUIbLfX0GA
E7+uTe1HNKXFWzfxDTk4eENRJ1DlQWt/1L6neDqhsdXHh7X5aoSuRWn4Db63H4xjQpyeohw4T+US
xbmk+cyAKtYNBhammOIsoLaDXHVzPjegJRf6uHX7PlGQO8X+HtdDWZvVCHrmxhx21RbUQN/aCGEr
qqe1anrUDr7zJbBFyilPJrXXqSaBlur1xU1Tc9qbVOVKN9DpWH57WsnPybj2UTmqioNGXRjw6tC3
XYVcBXlPHBNQI3hakXiE2VICSsBnsbHwfBcMXdL4hh1/Caf/OFkV1Bjnx+I5z/uc+EYpe4HJBpcq
PwuyRg24dhGgRRgGuZz7VkmMwkHuEsT2uZryKldx43WpPg7sexEMsDiLcWhP1BYijrCk6ZSP5Nht
fN1IQo8TNJDwpcjRN7SG4sw9a8zovaP7wz8Zk8mMo9HfmT+h55HeyvZ3WznEWIQ78Ro21dWN6T5s
/DFLVUPpjuvFIVTVHMQxIiY+bybfgweK7ZXWgyaaGfJTPXWkns6kNmQbxVL2cr9MmbGQDL1EqWag
eRgNBDudbGCN/OneAKH85BwLkhDP2cZnAuziu8TKgoJSMQ2Hpu+db41fP+bSO9EXV7eslUfpQsTH
1OMF362oE4flFS0BMKgEOlUDG7BM7aM6zyfs9+CM0VmOMcik6XhdQxHJX+4Qoqkv+iTF5IQMgppJ
dkul8/efghuaDtFYkCnq/d7qO0KEdBoHfJiJK5/iSl7fZVub9BYg4xvstWzryp2H43/5pMNtRzEg
usJpPX4ZmqIdgmjdy8JFiG9kVn6XmKAOfIIECK0qmXTYqXs6JmnrOGUhYnqso7HEB7BFXB8YYXHF
2UuDPQaMi6eU6pQ0pRdr3xPEvz+xfmtM32VtpCR3Sp+bmKfUiayWiL/CE3q6PqhYnEH9GLP1l/9o
EufU45Pl/l99F6rPy9btVj/2wPSmN5FPsX/z7WOBT93oppivOA70ffw442n4wNhz+zxtjmdQT/ec
9CPV/qPlafC2GUYZwM4YRG9VjvgYypvQsZ4uZwC2o4uq6Hy2axkkxShIGyHwvFXSpM7C0fbLEMky
A1kXVD9KFOL/Xpfq1kvPQYj1C7YMIVuz/KzSeydE6B3Ds0qZ5ifUUxozoYmvHaPJdnLtWfgJXjH7
qo5jXl9OUWlacR7kWjTgoQqtFpp/JywAYzWGTC52yshEMiTkM5yRMQCkqu1Nn+HQs9ACfdYuT8Cz
Qd8UXx63YFuTGF+NtRpe2qhQjhKbN1J2FE1/KRNHOfTna8jWWNMfFYLJ9xd4rzFiFbtdnAqlXuCi
xenLRQnatPFwtXeGs3eFtweT7GXf5TnpMwsfMOaNgHMTzt2a/aL2PA3ktn+XEi0k6vtQxkHo6A9N
NuQ2RRckDJLXsn8BWJ7VM6swBER3rE8PJWJydOfLTGAqF37d4cRwbyefn7O+69haIPMoUvp4528/
z7sM6olGP9wkq6YsJwHPY6KhwQM6doMzx4RqikXtFMLXUnRZrVOZBHFkHQn2Ppjzgs1PDYQnbnci
sOAzXpD2mgPQVl/HbitcH63m3LKvYbtCF+lB/M++bGt/XqVqjJYzj6aUkvQjs3Lz4sY1nxlYpmpA
3CAMURYcIFRHbTMJDVGTQw4pOSVlVVSakcmMPssqo/ydE+8eVBA8pU264QlSP8zyn369HyKD3Ggm
AQOuMZSv2c75H0jYuz9Qv2l8cjAFgNhUpHy2BY3/wm50NgFyHjUba4ifVck08hT3GU3zJv2ZUsJ5
HOePNat9kLK+HrGjY61G98/W0h7wigABqelsbxN/dq5pDap/N12/8w5ySeCqQ3F3mxPHXiyyx7Fj
PLVpxQ4kF2jtNWdo9c2wrCrNEyE5sbQlaEZtEVjlRLOu+0qAYYGtteC/qx5L/FbDaKyGqRAev9lb
qAWSTv4q71ZG+Y2kTP7uONpOvXuqUeuGNezg6L+cymZc7X/Tf0JGJbMjHP9iRIPycjP/vC4mC0O6
/Kf5uW8tZNA3TV3J3S8BtIV13qIFCwr/J2Tiwz3JaSD13Hv0fUN2zYmRI89EKlZ3BLjFUG0c9F2b
LNgU5zBpxZsjTCwEOtaOxQHDOS588Al6OJ/2nT6yabdYK7aw+Vz7g158aaGPfc5M4Jn2vW6XxIYj
N1Rsq8wipeI5poVGJtrT/iJI+vgdH4rDfJsVy2tuOwycqJKVY0ttWgMGF23PZS+miwegelSH+n7N
vmjPQqkbLNTG9Jsqfpu8vIcLY0G2axnzu/Ah9T/BddRf52t3D8RJ7oSP63VJXm3uNufstLfZwu/m
+DwkAe7jd/MktidT43LW0VVxyKWo/qw2u1OmsEEGsV8AsT3yKm2Pog0pmY6Ez795l4mHF1HPrYhi
LLHWbtPgDHo69aOJ5471ov+SUdngNQtWWS2KzKr6nyN+45UCNBddfQHxSzSDCMIscR9HrL0X7xUn
K82qcd+Vthv1RcFkcabEgs2DC0atwcQugmmszkYkS0EfXnpTr78uyYlxURoJoSt/R/ruJcIr996O
se9iji72D4xizW9vu/beeJ+kf+YuHevxiIWCm51kDCYfnqJah0OqvfVG64JE367HAmI2ehHEC40R
bQc43sX62vsVEaEppRU/JAvl6PUEJLrJEepg1RA/ddMGWALZ/XmER26jCIpr90HmrBXiIHo046J3
3TwRLdOQVueF8YZ4jrbxuzuHQjnq+QCQYFsEE9PMXZVssqTppa3muG6FWDLkjWZlvon1ewOnCtqS
WWqBhQb5W10++1wOFxuM4V1+0zJWKL7WG4gjv2amyDcKW33e2gCjgoc7a61bJyzNW8GgmE5rvPpS
n1f7Tyz6GmroTaZ8mKxdEqBmlQPP70gwDgXyu2MByuEP9HFOcHOmBghGxltsvMXaw035KzhkJleI
vuc73atE7TP3HOeB69jilzfYl6aY6H9jZLNTTT5FmSrS6tikwmwkIU+QjxUYukNXLi3kIygstTj7
uZvBN3tQr5TcK9I4gx3xUQ5DIfvDH13RbNROae4Ughfk5IGyFjEHMaFd7THRNvN7znzAs83EUNZf
AV6+JId8oQLC8Upsu15TxU69wMQENrP8LKo5Z+5lN+TOfibBpJWw391T1lHLUjdfzRaC9ox1fQjW
uPCyGXNZa/SM+U5IkUhOB3zIZNi+xfCG1JUohEsAoy6EbS7eUNH6shbIy/SZUIxgFTNR76MQ8MPz
TwFOu7Yzbon/S7rAIznRfou3qONbx94P19dK06xNSt/YANA49QLXsFgbNfgyY+cgaS6WdP+00DRT
Ctnopyabm/dHC6vHCpJH2vvcH50SCbwnx1LlaLL/uLIU8hxamhXjGIkTszVAee9Zz1hYpujkOGpf
AiLUKc8zbqb+GZ3H1Upue73ndgB6ij2En9F4nvuKjn8yGcwzPFNg2w+h3RHIwh0BBUFDo+ZePHti
fw9rNK3IzjJWgSK285zLHWpzICscjuDw1dI+XDFP1llu+yW+BDxIiBGLaLOHvjKQ0mSQwV1Ob2eR
VrW059mEaSeB6d6lJuoYHhRlu03e67ybToNmAjoO/ENFbFNw84cSJ2sqhSONmjM5MLRElu0ddIa4
qHiOPM/SQPJyE/rAop/vFuZezyBvi70Tq6XIDyzN6rkTMsER/x0rXV3FhtneBd+HsDEfQkxxrDDZ
UpQR7RPPOUSjVZeYMIUpk4EwCgeV3u4vFapSJ72SZ90QRWcuZpDrvAHU4jdFfUtKQNJgLe2bLyN2
efQAKaUT/9ixffKo0jXbdj5bBFj6lLAtR8XIvb1EZD7rd+t47u6DiAohyAPaodrF9pHtPfnndKVx
Heiezh9pwJ7A3ZrpPg1Q/aFKsMTRY3dwrDpfFwOWNhGytJBEKk9ocySucrkaOKP1ErT1NM6PElME
3vUCZGWcIfpvG4cLtMCuimlWPaVAwXOgs6f8OPTopsvMAFtVZtlVsahP2VXJ53y7/L0jDsz6fqFg
T6aolKZYanNTlL9XdIhHD62kGhNGBi7bOUPs87ybuqh5Xtc1bjwVLj98dJZ5bfIat2pD74PxVWCj
tzOM55ihmtTZRX2p7M787ocrFKy/HSDt8fDM22vfJbxwXJEFig5OYg8sHImGRC3AlnpgLHViIGru
ovYBImECkO/fT0MhrKqmHZtuOh/98x3aLHiUXNVG208VLPErOjkrpLqADVZBqWRTMbnohNGpGQZv
jO9NHzNIsRjc4RsSwvMCssUtAFpPalc3SMTExRPsJwYp+W0ZQZqkVcuvZehIQoeZ3jRRVF6+eG0r
s8JKfqzevdPSr13AveRj87K42hiIlfZqgRenIHOIsNuDTxF735us4ecnPcuMgqfuD5kcufeFhX4R
dyYrjooAGkqDnMK33fGfM0YsJ2ioudRou8m9kgegl2EYHQ9Y7HVil/8SMD3xZlfgEQ9VFhlHmBFf
f1GeQCNuVjmBjSQnpw0qv0hALr2yWxG3rwpSJLO0yJeJSfMtTntb4+iuOL1z2YAOr9JAoDVkj2Ml
JaSAD/k4j5f8xq4IKcNeXABtRn3f0w6pFkEjLihHFWdVbyEQRpJoEkavgEsnU+Zk4ezgJBkD8C6j
Kw16BRXyjipyHYsd4Mc8aqA4wOv8Y23vzajlf6ZcE9Q+m+gHkWIGDE8WMXvUQ9c4+gQly5lmt/SR
Ne2tMnSJpMMObq2JvzDl+N4gD6VTcvHx0u+MOeWU7LmzHXglZahy3daTbhENYuOw0hVseR03vv4k
Z9FPleR6FCzJpjE4LG9XZMKzocDMIQKLtXMxAMm4ZkVMY8jfHx5vc5VM5dCzvOvhVkDamSOpvaDD
Pa4bMr5o+e/yT4KNZLiCSUCAw5nCZ1Fg1ke0630aJggXp8n2BQLLRatppwlj5lYk7oZ+W+mFnYyz
bsiSLFXdsEWuKqTZ1mXnbw0nqfAuJY+acHUWhsM/hEAEGS/kOW2QAoZJeDdCO2pfbsmHH3XPSvXE
9VLpRkc77Q6VII3PJ5KJbknxlIxdvujUjMUxmHVwAFCrKadIGaBTkcZkAHcp9MZMMCPNLJfry2ru
a9gvsxjW03azj2Z04zE5bnYQ/KWPBvA8MB8nsPG/K8gfuUVVO9kH3arwE4BAxog6O/AhuB98BCXY
sMiIS8op++ErMb+lM+ebde5OfqBgsnh0jgtEm/KHybK5CluBymaBO8B05RhJElMY9fCxvN/TZMHx
g/oXpl6c1YOX4tPpuk/jbE1Plwq1IlKW0umCuiVaVQER1TtSrBxRWxmv1rETK1cyuDa1NnJJtXsq
V5OluAjUSbMY04oCNiB3cqbC/hCFOvluT4mFH+6e3aA06dlbtRTzPT9qFoHqQscjuwhDHK1NT8kW
Kt+azItsPfeyq3v0EKuyGgDKSQO8EGw5Iwr51NbRy/Lv1j4SSVrNP19JCRD6SfVGKbDK7VVVthu+
8Lo7F9ZFkjGLevObge9heZj1y7OYIoA+K0etl7zRe2XaX5hOlfQh0LfM6MOTPWBC/auR4GRMNeD0
VU8DQPeAvAC6wucQKr9rx6q5x71MvL3jMLokng9cwJ7FDgifupXsaR+eL+5DpHxGpgtNx48EaqSk
LD1VN2UebpINg/IxZPPqR1jRF6lUKYKOhk1azUF4UXMq+rJwEQCr3KcG/S+Wr3QQy1nIYuO8pzyx
Mg19sLY/bjBjTQa3gd1ntDX0iiZmu/pOyfvqrmMftaFRZ1M9zKE4Xq9H5fq7XKA4h/cjckzpcopO
NtFjE7oIdj9FfSYXArWHVWeiDr9vpZi9SjtvomyfyGs3firQ95rjZnS/XJZLBrxWF/NhYmwJo4th
cp+Stxm/oqM/WeyJb3QopsVNWVJhrj/dBkPT+DdNf45OHo9r3V03Z6YzqfLEYqyZMpJ08NeyDzHo
qjxaA4d0O23owrMV00QIfvKPwN7TeLogAawYyK2UDMjEwIzR/JfzuUpim7GZx+HENy8HXX/3nHRn
biZGCIRdMh2JAVQvgwHnmLm6XrbphkW3WZr2mU6e5Z/gKoJKeOZAwcMfYHSZKP1TtKwRCLqIFBgK
RCXyuoeCsVSvWLNr1y6g0r8ASU4TdKmXRXNBdgtSY8LwmlZlGapCXYYZHy6b059KOGDuA73M4UOB
6PliLjxSSCcm/HsvULYBLpVwoIvi+dwTSlO/fIWJwmvGGQj+20wIvplaUVoO1JoHC068fg9/HKX+
egcDHv2Z/mBw5g4TIglntZ+q0wQ6xj1x67Asv6rEGjENL/Tab0Bw2Cj45zr7PeWfejOXFuCgU5L1
ssc8xbLZ8ytHBexgtRzjr1qZ6YCzDMx3l9ryYBxMeNvB0zLy3Y3jLxwt3Pd74vi45Ur1EM0PU0Br
cGeyTPvx1Up/Sh/VywmK6UioC+sErCAKEjlt8oJEgWfdjq0Z2qvUpvHq16bIsl0igNsdXis/NCJW
E+lsDLFlzJlWH2ZWlZeOhS7zH4dVpfgdKBFEUFkfD08DK4sJemmle6XYORwcsuFB93t++PXuW5Kp
AfGXX2lAbOv+PrsxxbOcYLYruOhCevKbe1t3pNjVF9mIuHPXJTcZZ/OOKNynkCkJJvKz46TzoXqm
tfu5WRQ8+YQSlIS+JIhVSQ9UvOGV0jpsoJT/4pJqyQDcmZQIgnhz/iivS2vtp1mfXRDosvKIFJF7
Y68ef2DAist0dFj5+0xOP3VD1r6S7z8qOpJwdsAWCR54QjR2Wv6Vw9m/idmW2QIN8ad6ic8ihlJI
cHQfg/cjHiHLzIWaxP9Hz+mEvTdhJY+jkrlVlcJ4Kscg92UTk7g6qB9HLj3/0s6+Npz5PmvkhrxU
fryE8OZql/QpXIcONxPyvWWFZ1liSbvQPjflnngiWKoZkEIlBLZv1Ap30fy/2DGtgC8dqOqJ+FkY
FVxbpIMrMHfUATSjA7C7sDdJH+YwH1T879kP3JAX2l/Kd7bd8bBcnz2wvZU/VRaHiwOjPOOUOkRP
/3U0llsZ2lpL6pBBQRh4XZ/T2cAL1UvLhvYpa4oYPndQkzQ0yudKySde0BFoYOtlXZzD6EAUKQjA
H44Up1fErdEuNbjh3CU0MPon/HExOiyfASUFdQXvozaZ9mpDKo0w/NVHzIeqh0VZeSVIIxkn/bsL
TfpsDFArSIeHdLjMPd8XpbH02HLYVq6sMm26hLWs5+f49oFG7loI+Wgbk8SjFYDDF04Pv4qQDtJT
PlhlVaZI88/hWY39Nfvzb7mc7a3YQv2k7+bQYscmTO20VypUXEMxE2y9wYWoYE2Z5VqANCtr6tQG
yAjMoq/mNlr0/k8GKP0UbtW/ev1M3c4l+amh7pMHCmDCeFvtDkHKJK65OBOZ7rKh9HepVbixMbDl
EANmsOBCfqRrYuuGL/r9HjR0mYVB/JoH910/eJRZHg6lz3acy4Hng5WOlRbTTgV4cVzRvguOL7hU
UMO1MSAnucc3VOPn67ijpuMZZjBLadkYW4x6DhbJSVbwuh7r7GdOe81KOXV++UTa1rVxveG165My
hJcdvB6vdq9bmMAy3OnHOBM6JFvoYsO42LHhZ5S+m1yLS8frxe95InU0mOAlYZkyqZMxyt31BGDQ
3ouEn97ke6X/Z/2VpKu1UCcwiregS2xWTehoV1cXJZ2mO3YvA2S4m5XlWLzUvcVEMsOD96aAIuvT
nRWQ9vLYuR2WNPJ0ucOAm9qL19D+lIP6NxXm30OBGRepKtTtLL7apKTQOrQVWcRNPypE6r6SEKkW
wVZSBGi0kgD40ACG7KGwGO3mXtye+9yRoD76tgI7Cwqk6RkSyYLWPpU9NaAszaJyF6Y5M/M2Jwgz
i0ugsUYYbIS4LD2iDm9GpVxIL5HwlLDT3Psrv/77xxrPLqo3FQAB3b2STnRPOZI+2lzKyUJrTtWl
UgJPktJtMp2WhJI5Bwh9iyLHYiwEvGKm1XyYTgTMSVUaO4wcWtysBfdvzTI8lb+Pm+DaCblRaP1n
vsH8cjvRe8fD1pyk7GatxdeTKfPdgshi5xnCzKQUPy5g++VHfEyjhpJWK/+wPqaJMPJ1KRK7BclU
dgrHHwodFxKSnSEqhjuT3CnelZbHuDzf61vPC/sdHUAFibfCqEtILakSjaZE1OuQfY+T9EvqcgwY
78WbGAVcimbuV2ErQE9Nj+nf9pVCfJtr+qE/N9eMzw45R9FG0JoqQOEpnw3VhyvVRoIbUUoUDEoE
nU8aeNUu1vyT0CUHaLdJvAwq6ZA1AhBYMPcXmSKiMY6ftbrksZQoiHp0N3945yMyrVeC1NVty7Ww
AzqFPjCV3PfTXESJlzMMaDsCZeoGonhwlUeuuAx0mRFFbeNJlhCG315DZ5ilOOa9RNphQdWCuLa9
FhPNAs7xQvZgJfRCNJyCD/ICfRoGLH7tf+iv7MCegMrNNnXWou2Vk2XJltPkOc5ejQIQMow4sYaW
T1MdsBG26zO5HMbnEt7FMIWN36EJQoYc+ys9huq+uAP9+LV1R32uhfU6jBjEjm8okKsOMRL4oqeS
H6lOroBVjf7jcPTki53W8UA1t3L2DwdB9rsljLv+i0BvswWm/gT6jlWIE7ipb4c2kd3g2qFVjrQq
GXUbQp7DcCzwkLuWckhwJy3Yra8jddWpNelSet+6bBIYmUkqUvZYnaZrKx1w4W84euaP6ysrK6me
WGHCynFZyIwCXN+l+jO9XWqcpz1PIWoLbqGRQtTStea9r8fIBFmvGXmvRjOO4iXMEG67fCAs02TH
K40096B8jU8ae6nUI00yZvGWDChZWIn51WoUsA7ShY5LAubK+e11wxEPlTUu3PdBdH0xpWl+iQKB
Mfv7TXUXV6Nkp5r4sR/WsZqzO3xYsPv9pcNtQ/kKpNl8kBw+IwqaoENdgvJgzV42Gc4iy4RODdFi
AfeDW2zE830LI+tlXh4O6MvrYm5Hu0zqy5xAgNBzNNlWEyiDkT4pkdgGas+6pdLYaFuM0Xqzptcu
Jm4hFrE9hp3e9KRDHx4lWVBBUP7YOwIQlyMAfh1DRjE8NUS+GBXWFhXMaltJVY0aUjZsSwXGdHXE
dEsXrs7LItfNt+FBaxhcptuPquwRB/lfhcwMd7imsdLPgD0EXVZpSHW6IQOH8UbStzYGZC7q7Le4
CB9aPMugXkSuO3tz6Y6TPPTDl+YjsxZEy1DD9ZTt04ql+1402t1jcE1xA2dSGkZToHJgzKAQkcQs
p1LpLsJk7dYSkWRBnasTSFiotycyTd0Z/0sv03nmdGMCt17mpOKyR0fVV8HtKsZm4xYvPN6Y+N5y
hPlDaevfPE9WHbsuYaXXwAO+zlComUxP1VguApySK3jDXa+rrfR3RX7HYMSkwJ8ei+mQjeWNbmKR
QfYOJF7X6FpK0lkJ58aRCioJA9ovmIadN2Wjtlqk3DU4NdRjRafa7LTroL6vawua6T1KOHFEeldR
kJUMpYtaEkcSeC6JgOQS9VcAc5sUP4XLz9OLK4iUnA4+9dWiTrrSoodrfna/vEATo4Psk3Sz6tuB
pNeu5V4o3quBrzppxCFR8WGHB6dGZ+6r6GBkAyFntt+XWdRIQKgGs1Mlpa/ugHEzeIYP4KjcY8Pl
yZuZwOz/QSlsNn7LCSU5qpcVLGnAvmCj0uDEVz953xq2w13kuudmuCqDIlqWqp6Afk7mNcDLZp8S
IKC1S9BRmhhRcZSH6dEJTETPvW5TgsyThmABOPtkECaebvFRbJaqmdNrIqd1pZEMTcUKxeuebTbM
tGyBiu0jsEw+RKXPBS6TtbEL4t3chR3Bag+D31dHnAcyYMjj+A4lRAW4vedxJ7XcIdj4hJpB+9mZ
8z8nkoTvjWrMVDcIrYh+lqqPOYdhyXdqGEk+OX4jUEw4kbK/1LjwiGhrCmqdjcFIFbftfnQ6vGwW
uO37RYlorLgi8Bo1rSrx0BhIrhJu7Wjtd4bx74DL+ZYLbfjZ4WzRaUJtSAtnNHNdDhgYQIwSog8c
y/Sy6mv1CiJa31DIB2STwcaNNftMvV8xk/ad3k/2+sZos/mqrpRSkTdVUcjSUCitccl0nQDWJJQ6
tC2GWxP/1Nk1UJ+1t9kFh1PNQC8+GrnO4+Sxv6c344lU1KQvBaddS3LjkLpE7045TrU6WbPsYFvb
VrWduaWZYD2bBqLX+6cFgjMKhHpslD4A5Eym6M2E/613hHR0H8qzCtgG7jxqJE83aX4MFeFcR2Qv
W9QyYPBADZqjNLpQtU+fMctgDDMs/xdHnOhcy6J66iOUe2ejXxVrm/rm6o9hrbJSXrzJssNby9Kh
mLD7hThUGk+fyGRXFVK7DZgwrxkYYyK30XyzcdOGbRrQ6aTYk1fl2mC35CO+t3mR2D7lYUpjdJsX
CJi2tKUhZptCKB7FJRfnY898kuVv/zF0H3xzsSfNF9j5/Ng6oOYq265gKfcN/VaQV7M4eockwXPO
qQ12IIjaMEPxX1vuax6jXT6AjV1BVZmcBb+w/N5ozOzr8SWEarkN5+MunZiZfoOnN0OEiWx+loTX
iBe3Jew457uJY+xhcyF9BYe9RaTlsM8sReI3SEceke96pC6f44XbBUG1HL0AUo22HEA29lkL+DbH
s4zWQladX/AC4yTzw/xT8+oy6g64MxRbL4juI5h9sphwJFtJFqBVxneti7J0+qc9TN/qgZOMGQTh
TuhCC84ge66RHzI8BXy3/bcpzbJ6F7eH5DXqjUEn5uuhszlhCkqvWTSwQHrv82cFZB7mfPqw80/C
ya/lQZVy7VZm+FXGnztbyD8r/vp/P3gcwzG9vFoCEFSWhPXnbT6I12l416MrIhYQNo3mLqrFxxwJ
C8UN8JxByIy5YPvJVmk+PNuiXgoknj0/eefv0VzU/zqvtr+rObTMhKxtB0EB64txYk+nzDpSNVuW
84ea7ni46bvj+IjpsdNtEl6cJW7V7RoPPRTOZ7ZAsagVxG47oClIIcwyL3nBS/d2G9s5PviO/Skz
xEk3We2nC7QSoTGpX/HRlGR/E1oEy+BGSNOt64na1Csx+RrTEQCCXBlIb6ChPv8/xJoCYjANIxAN
2z5ZK+X22MXuCponktggiPJl7NxqP4iRV/S04+TjNZtlZORURueQg5Zortjtz+eMDu95zEEYMojz
5rDPgVYvlwyCMVetKroWUjJ0QebJ/RbC0lCLskJRH0k/bqMXfPReaL+JDYqLkrAyuNEKjVjZlrnt
QbGqC9gyPCURe+aXQ/Y60vjOTg8AF/hxBVCivultadGccInAPcqK0fIZzRYJdnMymGwJdcyGxt4J
4WHsMAO1pBLzGPZrxWPOCRe9LIphZoNfmIOf429Je6SoYiskRIoxlsAeHt0KegScm8KnXJcltfGs
ydyriyztTqWmMqv73x07VVUXUTYs3dfJbvx77hS/tWy54ohh8cYIv5d0UsUiC52ALa/8HFwC2e/V
kngL6Okg2CPXSFJS0YA4nOVnhOtMZDZ5PlaH4FVR4ao2G1r8LgDcMxpcUORsX+nIKLTEKK8i2+0+
2WOOpd6o0lbm86RkfHE6ddYZW71eWP9e2eRi2bF6/S7pVuqROxD3BcXztlJf8vKJTAEsMNdHplPJ
xSgozG0vQHqlB9zSekckxLC8r9GBN/AjHHop1JV60iUrOaE2G6I/xOKRAKFQWguR2oXZwYEhaFWB
uIUDasgBqujuAz0ppwRjLGO1cHz3lp6JMMsksCH7siW2bF5AtatmQKjprQZFt9y/Skm86gyVxpr5
ElzYy2ENMbE0rHVj7JRDm7y90xn8IL68ypNn3u0G2enEbWTn6oU19GZ9b2SKih8OQoNpi8hzjZrF
yuCZ9B139ZHGplnqgkjrnz9MZsYIbZE/W3yewaA+exUZkJyC5fi0K7yIArAcdqvL5bOQ9K1xDgsT
QZykJQS2xpK8S132i2K10V69G6piVMxhFzyy+cP1x8ATdRTokaUP1v8LpFKGpln7hEsaeuw7kvgJ
+M2ExpaxcbGnr71hzWJyQH7e5BdrjpVuFnDGjPVTcnminZ+PklyQlbZd+V/NSZqeAyFNjvZwNCW0
fl3vdj6mDwk9X+oDu1fMyXuVHTgblaliINjAYMTy4+QLmT8fR767y9QHbEkPIvoPFYzAWmUM50mY
pp40+rqVxvtdItH6R9flpM/3ZXAEr81UKOtEdybu1nnRhKjtIwqLZ+1ZHSTNcJeFzFldcIkgPo5V
lH1rftiFrq1RfMVoCiKaLSTkq/EdAlLZ+vVTN+nxwR5pxOmoAyAVdgq9Nc7H+IL75Nk2qNUsr1aT
zVcf/A6LOvj+xHVxSFdk3lfkS+Cs1irJui3HnE/wj9Up1kCvu1mkmyksu1ex90qoAvB+icmHk0cy
9rcEqR6a7X0hJSKluLU6aMqUBLwupxLV19B/pHXXs+z8s5k3NLse80pIcmftyRHqeNapPrwT03JD
l6dQramqEHKu01bk20ehsH+SuAMmVAgwgVAS19EDcKpt5IEOkCpUL9UNTnibpZMmj8PrMmLVHpIM
F1P8re38M97HyQC13rgTA0xgbiGqcdh1BDiEFi7r933sJWwGzamHSYmU9fDgnSZOC/uWzB6VNvo2
vQnlJRwLWkndszDpSR1TQdEXWwzrk/eCdJqn498BQSl6CTVwQXT5Osp/Se30aIS4nIkPddQKa46u
cD3HMPgVaxXjvYXXtxARhKrh2Yj4ZDnxMBRlDMT82ascd83CiEIyWsM27mWshhtOVLuiLtLEk2bF
sXbOzCEG7uIBN5+NjeqWBDn6/4GXFa2/zlWtG53Yqq1tifU74g36AYTFDQ6QDmQxV0VKB+zqdTY4
xxE6gqXElCVzqzcoogdupKzFXoDnhPjWVCJDPyoYvZpovgGgJJn3/CYBa6RtbKlrwUh+N2oGnROC
ZqkINr6xPBTfsLMBiBZmQzQnaIonPM+CcSJ686+8VlQNqjqGRJnjzJP2C5kfyhT6BVrOBhZJTFjY
L1ygOJTfwalFOSUS20UOWzS16QjK5lcbgPbrD6xl+Nn7/dYDB7AU00/4+9vDzy3u5y8SDPCxzU+B
u6yFFpkEVfkhW2e+TQyJAnySkzfVhCuSQVCbHJ5r+kLz3fP8nze2hZ+OmLafi/mZATEYL2kCDdQf
YW4D87zsAk2bX0afxKz3RSRpCkMMo4gI1cJ+cSpArJGS4VVAzMdxjC01sEg1bldBn8Qyq5+nGXxv
9qeMDEpekOleVOhsmnlhFaVX9CrPjelsn57aMyl+ozzSeWZIbixhGm78wEKxb4CX6mk9/CGlg2RM
Us+ZBcN+z86vEsSFEY3FOAPXu8hsyk0yz99akWRU+iOfn0pYc+2KncToWvNLSEG1RmCoPpjTCZsq
Fc1JIdg7L0FyczQSydWvtn7EdmHb1USFwBv5NGa3F7+j7AynDO2EXnTRRlgEx99MyY/YX146pdmu
hi/zX4ZG6/ScezisC+HJv/Ypiq5tUpZVKxkJ5EJzYYqOGs7i8RaQUQ/ezZqfDHZm0Su/6pgyEl21
62NyVcuHUw0LCEDvjpxcDSZfTC5sU55thugfZMi1hj5UWn2Yh3wsiylHA9poM6ZHsGYdxDAF4Asa
rX7MRjhUZilVlwsd7R0PzF/Xr1AlGDgUYIlZOUclDUOTG2UHvPQBtMX2W2c/DasEtGKxt3rGK5mE
dM6A6f3jVLPAaqR8WORw9Eg4+Loi/VXvnXGoB5YaMPAvzmY/8JgVOXbXhLP3FyU2WPlE0hO5KgBm
GXZXrXI38YA1wxcOk5AOihVjILTCBr6sQHXPIxZJ27CguV9Z4ShSDNG3/1gLIrIvkbzCaracZwsc
TkHkuN6YsaFJ9qfmgq4rczpxQEDT4Y0MGsNSUx5TJVv9pfFJIclTbH3DQXG6QH6OcwHAAhwJTo6p
/hQQNGM3L7Aqud4BOQKQ8k9jKdQSxJgSL2zQ8cWv6FvlnoeqSfbzyJmmMEhzm1tJhbgjrCxUd2pq
By2by9IJ7T2tZImPNpOIQC3j053yl8f10KRPmjFXA8g1CLwTzj9bHMeCYT5Q98bkUQsPp+AvfYIF
RahUqEheywDbUzCrkp4BTlCvJxjmm1bZw+1S/zIqoaPbMgIgVb8x1z2GZOkjmX2ypsGYyxuTqimr
4AjIVX6UPOwASuaLUeSGMIqF2CxrXmoEJxiEKilKLvI2UqAq590Fg1wWFomNhNBc3b15cA9Scc0J
gYkX//0OB/vd3hnJx6BWFhd4HTLFSZAMMjzZLoeb0Zp3nqy6iREjaZYiqoKmx+mw6lRZgBIiu1Bp
NoZC7zcU7DQlPwkCt8Gl0GbdE9pJl6FsBhTPZ/8f0IBOT7jbSBmwyd92MwgAIhcwZp5bmfdLez+q
mUoQ+VxSNOt1t0NTt9A9bRpJnRAQ1ox9oRHrRmDR7Z0EJTZu01AONNvyiMlgfXyoXh9uz3/qlsB4
4n0OvjY7qn1pe7Ej8uPWFo4wz6Gu45KAWub1gSQ42Iaf8Yt69A7hdHY1E8oquCa1p6LVj4H6T60b
qp1cYt5iNJ69swohqXig7ssAzUwnpzjBfhnJsFgWjnapxx5fkbPVLin2AUx6CXtf81aTx7ECXW57
yrZjjG2pcg/j5y4BnhP+21tkuWoIyyOvNM8aNCocj5voRH617/7nMlF63Ey0WRiIvsphO6kAVZMr
eSRScH3a0nEE7uA3eRCG1+KlFgW8acHF+2iE+qgGe2rtrtgLBlqqjet+WdeLktv/t41Vw92ey+Kx
zkeYFsxUE3Og+bEKsDobICYgODseC3laubfUUfz4vL9ry4Es/xlme91MTn7sloh4j+UQQEUVQgAo
wZpnuqP9D1lEpyXVbYU9Pii9pUecLRom6KiMEYqCLTswPHkf1aaXilkYLOkL3DYaRUpX2NcYYAKX
6VvXa1KrPoVM4cDgr/9XmbI2OF/QNHwGgFthycBJTh0iEdqLLBUPTutBiYnDf5G4n3vzsKQ4U1wB
mKfvTO37hJQTk/3dsHH+0IY2ytOJsyEt6Ce8PIWi7qZf6aLODwcCwdO9azJx8VQIUgSOTRCoA8N6
WZfZOi3BKZNJVAK/UtWBKi7tg32BK0pR4A3DzL/pxVEFhEDYXOU+Su5fXjGmxqYeDY4d0aW2JR33
LreHvFn2LVe7m5AdF7akPI4SSjg+WWrsBihxJ1jdJu9Nl7pPFT+sqe6SD748Y4z/88OKexb1fu9Z
qC69olR5JyA/4+OEq0AluS5HkQ3COOBmQ5EC6BZaQUPmh6gK9ivs7hz9SVXW1Ab8CEZVaisUXXSW
xwWw/61lqCwoHS+pGECS1nfYRap91bIW5BuRj1xGaEwqFBUI/uBviUuH6ur1jpcYzPAmS4FHqW66
WqrSRxM9/liQwu005Yuf3GgFzHHfCnXcnm3/AEFdeaonzNSho36uQASnU/XYPL+AOuyeFtuBU1j+
6oakt82bkh+yGA8FGuRSpKRnpLABwJaHL6hC1wKRj0cwsOpfpsO83A2iEm0CXNgerdFj6wdav7vB
GkKlOgsdWDvSgblI/Pz0CG4BL+4YsNE8KTWhSd4J2hgCyLLzpw7hjow3ieAys2pgaTYfSpvu58i7
JbiVL7xXcek27XIxRtXmuxa5JwzPuN+yHVnfx3kSdqrT0c3F1ZfJwe/zSPTZGz+/8M6BTPCWZ5KS
kZKf4oF4kS+NfFRZhcJqfGkLcOTOHHHJNUdWOs78z+AsT9LqwYNHfB6U++LbQyCjWIwy4uBhb4HJ
+gR+rUDn9770aTZwm5mN3lb+dv/OpSUB5QRPZ/4dqRcdgbTNy2QaZXknXa4FH2TH5WMjjObnbgNZ
0bgHBfrNsSdO5OTfzhXkfEqgmiTP3+DJOeWIjjoYXyDxfr5/aGS6x4Jm+g4ifhHAfzw4ZRtAo0ui
2rCF5374YfiwgleKthJfRS4cdIUgthbi4uvoqaGt72ta7gjAcD8HEP7vd9Yep6dpKBubxXGUZwLu
5hPUIwZtGkkc+Oh7FA/KJRIEf7UHTScsQ2bHI5nS5PDJ/hvW+qboPib/R2U88IvMky03y2aEoUoi
DQnVxC+vr0Mtjo5I5x0O5dmjYjGFT/1TK/vJTNXuAnRDa4GN5R6E5EUowhCU6CFk9F6hBhy43Hl1
LZpIk5g/UOEZEh7uDyVNXddLW8zfIIOde5ZRqrv5xcwTJqdGKmlKHaABnPxCaCa7Z9sVKb68ZBzV
2cjDrw4ZTbhR/ZUapXL0bLQ4q9rnNuKMJ+uG+/f+BpXU8QTu5a0RZ8gAU0FFNX13BblF6MLYCYJU
+7xETdMTczQyGzQ/2l6AGEuip/vID1rgEgD7sPVGFwTO+xvtSuVl9TJoma8j6dJ4iwywf/sipQ4j
vu7xTL5bxfMMnLi3SFpYinkDaFRHsz0nLgpxANoscgy4+hEYt5Lvl21EXq6qVv7cR4DHbSytaHbZ
0CYvShJKV5tuFYT5IXbPMbg8t7Wi8o22MgSaTAnNQNDrla9bmQiuLMdifFzsBYd2oqFpDzj08bJ0
3M25xxab+MtH4C1Dj7FRyiPjulV2ppp5i5LgXPmkqNY0Dx67W/w7F6DGSuUvEufbbtqSm1FHHqCv
GqVb8/VyULiTPJtUgbTsfp+E4k2wol8aHQvWD32UJ+bsHtChRysuDVLTrGvsLkKw4DNMNR22H7vC
kp3epqGBs1BhWA/LNB3fultbK44UndcV5Jn7p1+v0XKqO78640an9dZ9Y5LECxUvKfGRn/M8KJgW
vb5bOx+OkVz7Ynthn4F6oqgbL3ZjjdyjYn7AcDPMiRNb5uDLHxlzxFKrd9VsqR5lEkQ9yyd5SZw6
QlAIF2xsntayxg0aP4I7RI7cCMmQgT3PfkLlu5YgFs1tikPruyyNr16Aj+LgXf8oxWbX6G7c9nkO
I/eXSIaCsW2h+qEmvg+WezEGRaYId/gasT5XzXz+rThL6Jbe9Utti9J2x0dBeQ0fCqSid71iUJDQ
fNndHxDCNbZSVccxKKg0nQGH58Ky3OwC5Cs9Opi68mMIwIwiAzsSNLKCk8MfGlaWlBYdRzOnolrT
aBLmLLooRzHCL1Z/vBcQv0jKmpl1QXIZjlp7HeFV8AMrxo2eTYLiFOvZwyIjO7JAYKH9NXQpfkKh
lRR3fBrqEeK8ejRsNMGy6Wg8UGXKS7NsLU7DlHT8YUAa/+KkJDaLUErG+xT+R6zs8CDpkdeQzogk
akvWQ59sRPhEw/jLhnh1vas8wV6ChrFj6RAzJEUaRDSSFOq8aN5GLDgyHytUZOAlAL5+HiSrtamB
TjjA9VQsKHxsQiioWEh5v4D14DuxZdjosnTSSWwbK6mpi/zFHidOdHxDGt4TjArz/fcLyHapklAm
czN1EWeEse1cBndnAx/al3hqXAxzNuVe3k3PjjXIopsExxY9NLRKL95D+SFRrdMhZag66CXt4XtR
NWipLqMzXj2Bj6aNAvuGOa74SjpK85RM6Ijb4sKbVd1u1FT7DKwDdTsVMuxJoyZ1QMI0Tnr6fa9V
jK6v6+eeFYiUxs/40mEo0Jf1h0rfB6Cgg4Z+N30BaRAIm62uah3m8fxR+NQUtr2WNDGTCLS5rJco
LXlSnBNMWh7DDq8ABUC5xSFWdKz1PqoKGNDjtlJkSIB9ea0mj+BipfgcWueGDUJjzfwPSBszpd7g
Z4g8C1Y34SqxRsEY0C1I47tcyfbKS4YhFpRMcPatlizxuim/AF5gH38qdPtQWFf7E06yhICE3818
h9/5JWJghkfahLUYmNGm4+MPK9q3jFrgDNkbQaAzH45PnXJQtqesz8BLXxUjQhZkn7kAYJcRyZ4T
D1t/r1pkrCh3RIFnF58fBuq6vv7V09oAfu8sVkLQZOVpLV43BqzN6kAAI5ryktbKXgLW2SmuOWl4
iaeqlW/RNlbEKVb/JZoGskLqyq5Rqz1dz7cXXFKOfOqM8XBOjoq1lMJDBjkwR/lZ+MCEQK6oNEKz
DPwehAuLad8TvPMMXn/QBLVq4CiJKcrYIOdLqgzzfIXWZpbzolK+jK+t//uyGbkntv4vx9a6KMkV
OG8qwDquCSCaVHZFbz7Z9B7FgMMdMFUeLHfq3Xo5l60t/H567J01tPufLHIEh3lcv6YdlyBFH8+m
asI/Y8tx2ZZ5gfgNEnrJVYSP2VTisdRp/DGs9XBEoX2RvBncNeCU1BtGE2XP5OaPhmkJ83XVi7up
mBgszCf+fYEYs7wlgPEluAMSrWK56ECAK3Uhe7NzAx+2z5gUCX6DDg9Owl8tDgo3HV8WuPN9PnWW
6BXXtooJHMAoF1vt+oQ60G2gFNYkI94ZY8KYgU0i9w4j/DfEbJauYmtn9y03hWphe35P4o56OXQ9
elPilYLM3R50mobKbocSiZuwZZ9o0c94rH/WcMMeRK+lJORnqaS5A7fLnmOnXF2PkIax2q5E/CuA
XM++04dDbmIM6494Rj110+pfjNc4eOoBHW78/vtDG3JNlVmkJUgct4S903xEy5o5rs8zFfJfxRgi
qudnwiLnfjrfnJYKrnAbP4kFIhqiWk7Fi4HdIOKPKg3eAnazqtDaB5n/t3LJwsY0gDUThiGyC1Nu
PCl7ViMDAPIrebBx57DJRRpxkK8iWxxJodFelUVK7YR4IB874vGOMN/3Cf6K0lcJRGQVzEVoLmOJ
Jvt+OOUhdS9biagdk8uBGUG5zUSx86mf7KUichZVddvl+MkPGkVZryxsQXgkhJ+dyEhOQEMP8igA
3av2nnPEemR13h/lk5vefAs/cUq2+pasl0TEkss6G32OP3toI5Ko5/aEGhhIvlJWcnCcGtG4/kLo
ji6m48ATesKjaCIeYSXaOZ85LogkXy4u5Xr5k8q+dyxOTvEuEI+mEJy4qmenhe5OGhiSeilTcUhT
TekszJCNNuMRuA2EDtib1TtAB4ySAZ8VKFEwE/ydEuTX60yn3rtmPaVxiTmwaTXTgyScPTnhzFIq
ATv0bvz/in0nJ5OCJeTu/swh0PvnIxGuI29yQOu5zheuktmZu/dXGq31L4XSjo3SbHxzVz+yYqM4
+9jpSfOpEZtmJKq/Z1XvtqgzeSA7kJi1B5jTXNYBFTEMRs0GGJd356I1rI9xFbn5N1ISquJXYNpo
3lOtMO/bW+7oZbXUUK/OuoT0+WPkaQfOlpPTbf16ai0T64jWuHQIOFBEHS+tU3JLq/tiFNaA3cN3
gQYYnkyjeAdJkEdDW6CEv2SVkx8xagvRFQB/8NMf4tiydJq2U9MjmICGiuWiksfCbT5KScLwsFSD
Mk1OKFK48Wg/99lDXyDswi+eXEoZ3X8LqXlU3twZKibeHrJBv+vipt4x4FpYyMU0/I2hyX4lCIBi
KJygo/1MhLZ7sfDNDkeWOEMUbzbNfbdvljfYyl1MGsB4WHNVRBii0xGnkZKlmdyEr2HXGiOOifW1
hgZMIFmRV5abqhFvVlK1BTF7IfFB+lGf1vgACCdQ1wUp5EqrIL8mgLiC84OoRM2Qo7nf6hcRp3Py
VHj9WPyx/WgU01GUjuabMt/mfoZmINFu2lnavZs4QP7MWDKzn+gxDrR9M8OyzVUYkRH5XfC3KTqC
CzCE2lYlppbzGuWgrca4YfqDXfjPYtcaBzsFgZlnUGp5fMGYFKjeiB/r/e4bUFvMlYP1gFCrqaFO
idLEr3by6/Mo+6mwr2b1y61uD4Zy7dGNzb2N7HeIVa3xzjjre/mnSPrPrhMpd8E98usRHk7XdUoh
P0EuUBboRmU/q+lXPNvGX35QhRgEtp4EH3uC38aQz9yfc1PPhArxtZM82Iv9MY9yWjbMGa85kbMS
0NSo9zmrNX+NeUV1iOTTa/7YZtRB62yB14gzwF51M5r1R2n99SHhqrvM8+QHqgKqSvJyHhVomk8s
0v83VJItJvFUrZpnYv48gB0gKUKUkO4AWMqU83bj12Ay22DxzN+Agew9pR4+SDusA/I/5ktU8LiK
SbRI2c5O4xxgNQDr/gztgSP5tx7tlkk7Ye52f7XcpSH+G4eUczQ/LFi/h+CquwVf3WuMs8Eex/ga
rLr4jkLDIln7alqdfcsmGoiAdOj6dzBZCU0hCu5Ne8oYiUmEUGr+67H9USRyasYnwuaLsBcnq2pZ
N013suyfqTKzotWWy7X/t0ksCZmnyaGgmjKE0P/tYeyyug2HLYPMo1wOA1jUnNIVFBwnHZOkzGb7
mYPoC1JqY+Qrg/eMRqSMLgAuxxJXdOFU8Ou7IWq287Z3nDve/aDIaUAXBPhpgBnfgBVtT+F/Eg0Q
otUD9KMTjFo8ZMNPdgsuSS2BuNyr5Nk54XSGjkrdDnE8P1HBH3qmDJpsv/Ri8q1KxHMpVLgD/xA6
RvrJVjsc/rI8JA/up3jz4y6R2UU2aHgM6SeuTTnQhWS/MPOTx57nHjptGFGGEcobuC2JBLhm9boL
tCcvI4Q3JQ0o6PltKPvqmp1TkSsWSRbeHtNYEYxZiGXyMY2fdbS45VXUkpk8Des+FPTnpFAyt75V
9klhZ42z/aUc1NS2EKb5Ql2/MbNgyLcDUWxmPGvvZNKhuD4vA5qBHH0s5SijXcJq+ohjkdiZFatR
TeaUJIMB45DPkzV351d30o+/VL3iiDnGujGWQkbS9h3fkwPOXsRGZKXdC8AH+EsTnl0d/qHdqhew
peN0iwby5zZcKWx06jg9QPYGncap8SyLxzexOfYHFi4I07sGnlMnFKmzphAoPbabUv4Oh9opbm+t
tggJ2FeeVGvcGSSF67YXLlsu0fEZf8ZunImmfltuvgu5Y65+yvkCbvjux34pI7hqBT7vmQufWxb0
E7nkPSvYFWqj4ZLN/NF0ad8FccV7SJnuD7ZgsmtC3sa1s4q3hEwEQqUedDmX8l8TbrlND4YWwpeP
spVMeSA8L/0XYH/TyWSLYfKC6RL0h88srDis0lIXXJegAxeNI0OgA5aH88Cd52Ehid3HTuB2WxYe
7hWkEP5TcllhIoY09gvlyBcWu/N4dB76G7zzVIH1/TTxSA1R+v5Op6OdstDdS0B0oigrAGEMDOmk
rbq3xcar13cpyvHW8tm21zP5rz0YSEWDDhgyYS1oA+bweJN9L7qtFz3IRcKH5+ssIZKk0mS7yBV4
7pVzxUDwLyr6/jXHEvyctx35qQ9Q/+YskgCby8X641KmcejZ0MbMszA2U9N14+pMzKVwN9RCEZlc
AfhJeDyePcK3TjHu2TMZuP2DXj4CadEPP/C6JW+ygcJhnqcmSygL9xuSnPf0IiB7tIbQoJ6B2Gu/
X1PhxzhHhCAcnvv8IIEKMCGHygZo+iwJ8vDhOo1CLK7A/tY1yCUYVKqVqye2rnai3cqj0nbtKwRK
KRQzpQGhy9LP5585s5swUOTUh1yZubH/RVko+93aVO7Iomph6zFHcrLLSvx0ve9mAhzsgNP17JwI
D17g5DsEH1of0+k/FWdaFsSgNkzsGmLnf2SPzCKYX4lJBwR7cKhsqNj9hVYzyLBYTazBWDmFqs2c
57Y273c/gmvI5oQwv+hu632s8usPzGlcDT6ANW7yTKVepvRm7tcD9Z3BX/LmPL7BpLaBpvK68XOL
EMnMhF2sXlO/hBwNZHkoRa3lrTgFDK6CBeqAgsqIuqIrbFWK6wW+yqqWf5ofJ/vW+SCOUNoPW474
6PdNDHIMCuVxfNR4hSoF7thB5n2YIqyV+u7BcVAZ8VAvuvlemtZlJIER36v1I9amN/lFOpw8vAzB
lVn0IPgmA8bQIdYyTWNcjk68NkbJzLX4lttFSFJZND/psFTwUFFJhxvEYaGW//JsIUd8hcL/rCqp
AR+Nslc9lOVydSgPgmXR4HhjbmsPuUPszJhWl0kSCcAVambz11u8VEzvywV6E7PTncdkBxRbZ+MM
2KOKwn5Vy5vl/qpeiypVgQ99mU/uEsYDT5sbmE/DxnNJwQHZHGLzs7PMduHdLEosh4vbIZOvbBRp
62Vxn0DWRuTFsc8UsWsRpylIsx6s5wRUt1f8N8tSZsgprYNyf2uddUylVx3WvE0WDqSD6IOqm7qq
TTlkS6Ps6vapr94u7LInDZvJiBZBmDcATjssvxNBcbeKKVeQWbSmt0wJ5W8lyOZT/RKMa7ONVfDc
BKvgetCoAtalEJhsWKiZ5sd8XfRaJkf1PGxwhuDrRA+PETk3TgucScqTs7ud2Mmk0quKH2zpJ3Du
BdKipf+MeAVc7mMfdeSkXj7EJbv98cCclZepFNk9SKfhURvCtm/TgHBMDojCiZ3epSW4FigxbJwt
6lVH3EOkt7pXVbdPjdWvl88TBcG6iC/4YEipkWNmtyNUTffcDuTo5pMRulpCnVLqH198PwPZN+Vr
d/6OluQG9kzSooKSOKU/n+wo5xoSOgJkIpR1A/zRde6MXc6LJiHsJBWomb0WPsmn2PDT3zDC6afb
WuvtrsMjK3hsmA695Moyd4h8KWsMUdaZBojX9DZ6hQMbzd1xQxpTGrOmpYDZhNmf9olxasGBGmVp
D0lNZS6Yxt2INpcVuR8QJIhxwLYeOujPaYRx4sLe2nxdBVviKOEf9z1IszklB1GmxIznw3lSYXmB
E202N69zn/zjuyJKS8c/rELTilvefAw8MjvkxStmagForxPXERMPD+6BXDNkhjqf6yYKQJFS//nO
8td3bJRXjgbppdyxI/vIEgawjrk2u8KSPcx5rDBLL7Qsir1uk91vJCxpfVGpMF4HaNjUHRV7AiYc
pvQKC1EmTyPHKCw/cATcsoDjK0wsCqINtB78IT5SX2gpXTUUnRW5YF/n3AUsG4/IMKu+vWKExoRb
FgpKjq+ADAH695VKirmXvzuAKUzxpD7/v5itqC+c3X+ymk3EX4RF8BP0NgBQ1QEd0F7yUkOz3ZVr
GqozQKPt2nArC5GZQbXV9ZHtpf+O0JJv9/SgveL/5relNEPmrIuYzjMzOXn7JFP23PuC/t4PSzh2
2jXCIFQTgaxkfB98i9GDkC8rzy+c3+0+iperq183/xOhCBBh9p5KoHbv3NZzl5MypbYlvm8/W8NW
jKAcWhjhAWt+jbuuJVZl9ZKRFe83dPMgCjXb1MumnUy9F499Itbxu6DbyryPbTdctpYAgxFtzcTR
uE7M3I4BK7RjmrZWxz7NeOeahSz6xKgX0k9vNhkdSRCOHNCIj4zca7MGu5OSHtxjt2t7RTbnxz26
rDAAsRog4YjruDmh9ha+QoJGWiz7NGAMYcudAOWIsqpGpkc0kpfR4IizMtFN1CJ4rM5etlkG0wQv
6pQWCqB5Dlb+5SozguiAlTJGPWCYsWhYZ4o4NTK4gnlaau7zjZaG4X8zZ0BMaCjNFsqhd9RjKphB
K5GzNjiREUfVBlHCmpFWXs5V4ayzgDcmvooYSVpN1HcRoumIAJEhg/nI0T/94jQf4NfaK1x8ZCOk
laClCyodOCtpDVDDiHQAfBYywWGdSg7i0JAQbu8FC0hwe0RtDCv47GcQ+MXTgiW1Bk3TwlmYU2LL
/utAgqW10dtpui5We6e8KZ1lAJhDL5SAh10w8F7/+QdMlXZHoXyoe2BYlYZlQXR7p17OpPpTgPxY
n05gOS1kLNmGWudzHdrNpSuFrJtUrXe/jXq796ovKjiQ7+//l6iWIpxWYQZP+LO5Kc+TbZLamdNe
ABkPPlDX5GF/hfv3B6f221jVqKSPrJGeJZ3s8L7RgxFYa7T0GP9Lz4lGUkF9u2OXf/+rfruaxCVY
v9XM8f5Dn4BYTJ++9oYEANKyJ9bRdJI3Re1OtjL3zC9G1X9/B0Lh/vCIqW6HAMS0PVMDIDh+wPjl
CfwCdL8S0M4ZRgkGQOWr8ewcE6SwuI4aFMayTZTofMxZo+ZMJ81kj15RkV+5DoAF5iGXdi/k8c4D
MIPG4UecorEIebpkEsuMOxXgVnVW4uaX2zWMLIIHpi+8UIpN23HtP6xsH6z8cUu2F6yWheVeCqpQ
LZ9Y9D+C++bOOkNv9u50IQSG1pjcQht8TOksTsy1cvBqgo4uZTTIfJNlftBZ4Zwf3EYqw5ifHm2A
yPTGYAadETelz824RJo0hnSGJvuX4Au+peaWAfZDTlJA38Pn56HOZ6UqgsF+Pny4vzJI2vS7HXkF
8J3LrU9JQOZ+NLLIMd8G80jJKALw3cMRa7qN6ZXTeTt9IPMbTO5vzClb4+lmdDw3hquipv+IKUxc
W616BxVQ2CzpzcSpVCzPF/VeWxM2oCoVPDhFcGZDj3+IYVTGdMOKwJsERM99r5s5lGR+FwOiOD+C
Nx8XKx8ZR+POej4IGhuojqyvdN6BS0ivGsi2DK+MVZIIJXZa0JonrP6ieMgEAVD1x86W0YqswoAP
db5NCXmpvj//OYUurWPuhUOcCqXFyra14ZUQADrUcFPv9/TxqWXE6/eZWeWA3nVw3hEd5aY7GJw3
X7pFSsHCxSUW6ilwi2LIK1qclvQczLOshkPvyudooEOi5MESEAi6PxnLywWvUKr9Ao3YSh68ARON
vm/e3E4eYBelVCjrH3vOR3JJJYM4wcodja4u9jviYey4ckejM0Bc0W/0xyB/nY0M8eRvGdc3223E
f2bhRf8N+2V1fCZoUE6S6CGFHYZV5hwWrjUpAPfmUUfbDHFsRiZlP3hKWHjopLPxgaM3G/9rtfIS
KRexQdUmZg3EloTt76mXHCDww4aAeH690/MUNGuUzR3v/gKhAwY3p+9JhlHq/2sPPvwq0b5wgWSU
NIt4GvUQjM6pxlXbUhkGx+MDLrCMGJH745jpuCJix3azdYyW0URQ78w0KhHQ5gX3jQca3sUG7Q2e
71XhlPkkkDv4fYwrTJIjx9Qx4Bf2pvVfg0ICCTLGbPmd/O5fGJuLKKhi4UPjrcsqr9Nox7Ztj/fv
t26q0bT5v808Q2c8oLOMST3Tl9eXDJgQ7GxpDRp5AKcRrRl7q1jflXQrG4oqx1lbv5glKRMFiof2
2sRGANB4O2ZJ8d815JQE9zrejH3lSUxBsqd/KttDtQzD9nb4MaGdIPlNdVpbHwyttyvnTehnzzsm
bhR2b1ygfwes/PaxTMQGNfbYWP4mcUzj4UM6tigUYzBepTzHWxPHp6sznfjnfFtE6EWpBKNBg0u6
Elmth+kU8FFlduqEj3OPik2hKqLUNGK7ar9Yit5Dw39ql9kOeUM+dtrZ42vNareeeUi+K/20ttI9
WCgQqgeTWhxo6DN7Zn7wx3955lXQQBlchRlX1EPJ332hFkgkyyWwWF37o7DMho8Ssa795XbiVCC8
2FZD+67wFFlA5b3+STcHs2ShG2X8v3ZgArQ3ZWU7tTEuA+a9Od7hwujYT1nGzwCvmNZ6k2AXF/5e
OtMda61wTvX8ZF6r77Ya83lzGMRJm1WOwtJonmahw5use3Q4ZMqt/cI6uvZ5hOLW58Tfh1/HHH0w
H/Lb8R9kzznlSmrIBFgLEDx1GVM/iW3yRRzx+zsADvv6PyDf+kS91rMyo4AYqiesXpO+8+ytQMwM
euA4BVGkmaHre4UbYnMnoJmXb974RgIHbQDtC+qKgSam/4pQXgvej4nwOXrPdgXPeHc5HII6R3Lh
/sAqeOi48APPSboRKpUjeSUnuhTDX4omVaTq5G39w1gU6QbZHvB/wBqODOPAKqOwmhQWru8VLfbz
HL+g4hUcFB/rLZgIyzAmrSIrGQWQXiqb3b4XJJs0gJN9SyW6Z5RCZfCEg1KcMnnY15Ksdm+1iJGM
wvCGbBckf1ina7mQBDfyDPeDK2UUOeg6OCmzWyumZxgsb8ZSOs8aZIwEWZ2P4SOjfZXOOu4QZd7b
MKLiKNuBXsiVTT7Rnd0ANUFVD/mHmqUmxyO8zMNA3Ib+Flia/ZV9TWpx2dS2JHnQN62Yx00nGByi
vHdnFd8rafNPFtv4LTwu/WpLDw4WJ8tzJkTODIGXx9qkzo5yisiuwDij9BpXyfNh+Bce5u9QpwQs
pjjTqa1BXQDmhZyhjBn3CWT9z7YXwTa1xaQKMTK1prxdhy2unC95ypSStDz1LehPHiujQVxdfiPK
LWeBdvjHr3wJJT12cq9Hy1hIvOy7jYZpRf9BOyuZ+72WnK+a6f64KtMhhyn1tvtvE61T4+WACy5O
fdsTchgs0j+AK3/lb6A31Mit3MeET9o3wzGqJsqzS38PrXNkQA6d3qex2mxnsO/HsE7o+vaT6nHk
KmhmFbYzQe+eFVBY8yUAzOPTl6KlZJW6YxSv1sEVAEj6jg8G5w1jAszlgzY1t5LQlYuUcqmutcji
lq82NIK07i6xwCxRxWZVnqwRn+dgYCI4/F8BL/tfdAXjBxWYFnW06o+8ObUXJySX74z3Hv8zgY4c
HcKNvlSuqROAg69tD+wX6g27LPLAeGLhlXWzOWA+3lFDPHpBTknFyUdVNHMazqsd4juKZb5m6Mqx
E+AuFLJsmaIFjBnCQ1SjWCZnUMKo1KJpTwvAB/rT6SwSvEa8BuQ3jTgm3Xwkm09rGH9XWrY3dc57
PtJegqzpQ9h9L4KKeN61s1rXx/SNIOkQYpZiXeL2XT9bGU8kEppNA/FtQatnCjqO+AtQwoscBZ40
yDxXOrOlHY3gEXoipOeAr65y0jjHOroLXlcoQw0ZlgsXKeMgrHQcx3U95nuxYSr5LdwyumyhuTh+
bA+dhI7rfq0OKgAX9hdmyCz2Kx1Lc1Jvg2SFjkvaHhhcBwD4f0brWK1HhMx7jOgH6a262/L7ELNB
EkXOmpiOhEqLPXerCtZQTgq9rmYwYBX+lg9+tk6msXU8XIDgiduzqmmjioWNzaQtvmrIme5h5RSr
DqZ1M/dFFVEmNIybIeRGTX0IoHOzrjr13+O4QxjelJR9walOO06U296vINfzDlwronX/FkevE3dP
uFW0/rArAzEro8yNt0L3gMerKOS/0/bZ3EBDFk4wnnJQaUXSsSvY6aGwpIY1lJ7EM1Uk3wnUTIzP
Up0iANHb/fWaUgx/SdW3aDSHblnPggmG8ylA8bOvf5U2UaBnzJ1XMTtOhnBoK+GNB7UEki6VAX+B
V2ZhwAGDf+sbx3OmPS+FgTeMnxoIqnr9zWaMQPdRAjQmW2tss4hT282xbGZMwaVqSOWl4OFkiZX5
W3S9VyJLj+WbphIMQyP8Ddi5inAPWKS35FGvZG8+2xe190j41wMKVH68EyRG+px6EWDWwQ2KnF+S
/A4Dx3eRuOaNBQf8ZgVw4eLawyDzfYY/sZolAoTkV9j5JdxzvJLZ5RDunWDi2MX1eQ4e5RjVis7U
nrL/1hMgkLIU7fqGYD6nFvUZFjii4ZA+0wnLFe1HkNlWqp7w4pLLgZpXJTHXAWrUzSXeloyhQid0
VGeJk/wPxmYq43/vYxbqK9N2wMTJpiCPFqjdBcjqtV928cm3holbyuMiLCc1esJz4SxN7liCjPcw
5U6esNUIfIr+fxXL2Hs8p9ruyGdMD+yUxZXEOxW5Ttc3iZno4VzeuozCMik3tBzHbqPOn9V/c62V
IK1fX6+m8JnVLzSZwHrg4Jxr+Ucb9CEe9hi2jOYi8tM+GGo/94nSaLyq7rCKvfwtDKRejDLkKgxM
Xs5/OABnXL8UtTqkr+F1rSVZCFEuUvv3WGpAQcySl1YpBLj1lQ3hi20bpz1G3jeSlzPEANChSBoC
wibJJUYY1H6rvAyiNMT1V9bkzQdasHAIsmp078B0yFMyAjEJO10w4OHsmy4AyPDw4Q5LXA1TZj+Q
b+jjNQGrvazTvaa74F8bnRh2hCpOAnYey5lZrnRydbn7P8IEIxDxljROuKLzQZpKPEGD+YowkXyP
JRnNaYhVMnIaoLJV+7U8AAUXK+iAeETMi+uBd0mwHFpYKVPO8GVzFHpGt/yuLsYScyCYTh3gYMjQ
u8yF1zFcpOwAGtvvSmjhp7EzA/6BILmDjLs+kFx9oCsQ+HOJrJtFZeqZq5ASGaJVm/TwbJnm2hVU
xgbACg0qDwGoy3wwydYnLOkF4mG/ApwUKkVM65cKNqqov9CFdovqZvz8BcBynoH7RS+l9FljAwf7
MzGzsTDeM0t7vb4acblW80G4Vmuxfj2vNhU7XVZBMku9FHqKnsJUEx/VCtUEoq43FqpQ2V0dZFiq
OrsnYbRv3YHkRqG8UszkkxpFm3mxVtPfXsn9+wPllOHiZpvNU16SofPO8evNzqqtmFljT1vnHYro
j0t6Uu48sMnnA+WrBmOMFlO1/gIGkz57Gqh7dipdqnibqlvjm7Aejv/SB94etGQgfnbEIlh5M1Re
8h7c0T0VBlChLnBfRRbrgPf8zHd6FZJsyl4HBx3kKm6+KocFcs6/VZ4MZ0XCVCj0y6IfmkeMzuRi
Uump9F07q5vK0Z6j46gMu58soxS+g52Ywl0VMsJ/vxuHO9dj5FIH6nIZoQNNNU+WLdtpbJyi/kZj
KopHuYUeqAhQHws+soEuKNmFxhy4ECnl0N9uX6mS+OOVfSD67iBjc7qEOZMploKQkGZC5uL3Q4RL
TLHiFJY9TdnE9JPNJ+xDHqIUYngm8m+eVSoPC0b7d02/ot52J0OT4ZkWmeFKJ2HiD/xi/CB+VdJO
hb/bxDAnLqmG//Em7Wrmq0E/IVsZyNNIlJlmDbhC9++NEhdUkeLDah5vtxDOPdEu0nA10Xe7fx1O
8rn1Saod10uQhKs/e6tNwMaz7Dpd8ANyppTFRYkq9YVW+5wlLGwqglPp7Zu9N27Ydq7umJbywJGR
wtpBJtRMnFXZ6awY5ZGJJhb7zWy4Fs3ey31hvnhtS4AOCj9k9UsDGIqr2bfb2YjiCkKo63NNO1EH
Vi7QiMJfoUqRnFp5bVuwaplMsNQYA9IB39ZelQ4J8ObVojnIwKKM/sC/18TA0FRYi39EdM3dxNtw
RbXPbQdTUhVPCpS7EeTIi0v+kjwDU3hlsWQcMoAroSovwLy91TJEt6UD+GxuKWcZTgfEWWwvpWhR
ZPfmmKieVZfh78cZRUAsud+0OyMMJDpcWpP9j89y45r3TP5HeZ/k2J9YJ41wj5h9CdbSd2F9h6uE
/5mzUm4UM4yR9GAA6uz3/g8/tqrHnKM5hjIufnT6iD+VypctiDHGyZ27M/GZT4V+j/yyGt8Sh/0l
MP34UYg8fFBMyK59Y267YYIXShMAMAnd3c3y9K4NCVAUBEY+foIUM/FVRSrxXYL+fgTa0G3VunWJ
9LtypFzY0OtuuaTpJkr95lsJr/V8ZPZhPJ646CNNBbVItKcThS3rfEeSLzw9xfY24908UEvvWPVI
V4r5M/2nor1H7m+TZwD3q8n0Iu3UCH3Qy1dC964T0af2xgqwwi/kje1MvJmPwcIOoHw0qrErfgnq
xrVcEZbSxnUF2hYeTiTayQP+vqyKD3FlxaZ+UaGFYub6bpjfP3umuPsadqe1gSd0xNoTvE4Jq98X
TfvBta9wEjn/xU9wP7CyBaBNavF7NfIW97MP+krnXL0zdlJU7tpv+rcV9LGI6otGolkb60HRJzKt
A3vwVDIobBAzwfHTaEHKFEB4F/jIR7IP+TuevNR9HtchTkl3dp8ib0N51im5LK6VFrqM/iQnziNf
0/6oeAB7KRAb4kY+9rdBxkQdjAb5dERX+aDsccT7tc+VIe8tRtJ6zMaTkmxLd2PjvEdmo7h2aLiF
bY3pW1XOz9Q1tcUWUbqWPSkPOz2yqkWD/ESWuIE32gWeL8G8R+3/M8wktk05AZWnllpN9ScjkvAw
Qyp8BnxxcDx7ljpktHQa1A1F2HhMxI9ibN1fV9zR3OJ9TODxIThrXwW2TwIHtboY3JwdBvj6MbjL
aJ22tcFryFVLVk4sF0iwweG+jEMBQC4pFVCz+T0FZnkcsQrCG+ZInEeyimNrbExo1kZeN2hSxj+G
IliVGPif4mHE18saFNoswfwsqj4ggAzAMfnpRTj04N8ibUAoPl8U7LntIS7MQ/TvgqRCCrJcioY1
pX33pDrds447XWs+qa7ob2dlqibh0widhbKjl9a0rAoVAwLY3xvBMLkZpEKT2QtDXLT8MrOIu7+v
FtidsPrIxF755OR42XRbv6UOMRs9+G9TR7IfdaA5OcsulhjSyD2hE71HWQnI85OC4LmcKd5+Ug/+
GRrkwBX+gPo6SAn3ajmam63OC6B2u3d00Tu8mWs3yVJqRUgGYPgakfh373OURlwBv6bvb/SQMMzz
Bk9O0Rb6O2RiEAOtIqyJs8LpmpW6XNjJL6EXlb9dC2A4ibil4CA7HPTMO01zmTr+jc2N78Q4WoT9
NS5LPQVxDeiypgvVxC7gIxnamGw6xvor3hpg2dig3h4v+zCGckxRm51I9oFnjl4T8DudWzEw84Xm
w3xw06BX7hKXRmfKI2Wt4PB+6sN93AZM4qGSnH0tZF9YIDkBSAFMNoPvZp/YP7nnQN7Bi+LwuDvN
O9IxU92b8DuEm4QdF/wosVryySdB3Jbaa7i5Ric+/DB5dVxjlXMVFE6K8LDBhMEScAjXPAMJb/AN
myGVMvE3FpbqsSExrcHl/SLMkyiF1y2uEpdg7+BkTp4gK51a3aXnloI3bZz4KsbPNFo1DdGSHED8
ArbMHEZtUg0GsdZnOV8HVrRBGsUIRlwi8CitWidGCtsFB87DByFiMUVkBGc+iPL/eLMGNZoiyclo
o8tOJNy/iS4BJX5q7ggOZbHjJUHkoMDZRzJ48lC5F5IGiRP4TwbOzgu2Py7pQ84oKKUEfFqH1nND
auQFaRO796x+yFcQxRDacH4eMU4G3T+ul9yXroy5kE2p7LSRoVTaYT8Vts4Sh46u5fEZTZjZ4+z3
gEl+gPJgJ6pl98YJcmqzKPlo6EZesU0ptOos8GyWk5wxQqssRCX63rMB6vS6EM35sVVuCRyaoLrn
LvYLd+2QKQjQKeWCOdQJOFsiUEw/B8WTl+S7Q8g/NoUs/h7rgCeeJpLfYo3ePy2q0gjc9ldMmNlm
iUKBZdqbNz2rthWZ+6BeKXW4JPclYeGRRxoPgFKDROIRtu7iHYumNNDnohVU2FVfehyYEE0OZKKw
XsmG1Z2Uny2299Lb6fEW/n28NJlZ5ryMvLyxZWOcqmZEP7etz7xzzFyM2MaMu62hJqHJA7ANG+QK
AEZMsxDiCXv7jyNWiZzptVmXslqOLA1AKL30qwq7fKm8nqz2bBxC3Oe/riZGs0ry1TuJvginNJn8
6kuzTJWPknU2W7cqRhbDr+XwSzPwQtEhrhxbgB7hVxWveOum3Kh14LE0qmr1Y55tI/BGfL52LiIW
ELHJhWOvTHib+cjf3vbMrzWLbvQ9Uu5+/RHHwapQymDGRo6TGdLvlSwzxZq7NUtu9BPxWuoI9qvi
rY+BRQLXXeAdAXfCdDsyC4ldHtcvZ8fNyl+VvxNbJSEqLKNR/IG7cfgx/P+vMbJqhlT6g6zmNZGZ
9zQvXdHYB5IoH4M5qZz0gA3BPoqarkQMJLQqO3GsoxD0rInlnpOs7WRyzsmBA3j+l6G99CMxUfIV
BMmc6OA4TyZM7MaXV/A2U86xArUGdCNtXCnDKntOhvFSnASC8lBo/dKVV6aohYkZmE+eD8Rc7j5r
AO901ktmbDXaczaY8mRwfcmBxa/0VCrAgsPSMkNPAlKyQpg6rG0TwutJrXa5u8PBPp1b6XNY21D6
QNzVef+IhEYERm1zFmyJqeDIDwP5ATlhHg7O6qiRZuiiwf4+jZNgGVdIcu6ADZMwfcF4Gl+ZTZr/
z2yvZkguZXnt4ctBv8PbO1S/UG3GaYow8cnYhR+03ZHYtpqLrXQT89rWDVHR1htgAbziJNfZEPnH
Z+XiKTsqskStQgmUzwLADbagLks3RJWVNugHDpOpEUpErA0NZEhMunEzmL6N7GGSFrO0YbaGGMk7
e5k1rqaKuIGCRtlqchKzoGC8/H8H370oHXkQV/PKnBhYMFs0PHpT7eB6QokMtN39Z7shxVIRP3ZN
vBp7rUaWUPtq96iuZtqkgmbRWxRi4Hw5ixYItl0Ko2SmgZHy2TcVXl1gmqe1XBiEwzZcBkZvMrAs
eYCPhfUiIQn23OZYfmGwJfFWQ8+FRdoFYdM4vQme6EqfVeEp1vUSc49/F/sfp6AgLLU+a8yZTL3j
CY7AFn5iKQsWwVJ0lsyGm1ChguUK/agtTNyft86/x68lkhWm+M+scBOi5TM1NqumN1ElbyStr+Rg
5E59PI2B6p8YeqKIZ+/ES1aRi8OAF3a+8FWJpxSQZQFcSPNUc8T16ENVumjjbNnbrdV+tlV2qWzM
NGXRrsAIAUnyRlMjQOn5VnxbpV1EyLlMbfZNf9cvlU/emnV0f5u6aDjc6Wy+DqPHvxbgzReOQpI6
6Az/EHHbHmb+ktmZAGsGF9zz8IsiKD9BZh2DeZgMjHhC55par+mE3RowcrVw5QRybwkxjviHRfes
4qAvz08BLD1/eYmxnCSbXEOOPj2U+46L/nVU3YGDoLC751d1RerbaxdfxjLDtq/hN2Yo1g4VkUeD
0fneIDvYeot9ftAfVQnB/AllHuLrmexwG3Qz79Egxk7Uow7k+mKES5ATfnxMZuUaxHV9E7iC0WS8
gKd/LYMZPTwOfc9iJHfdkRiIRqT/ULb1Cqa7kgJB0xsq8bUmc3i8fECS+wGY72LqjApctz4hUl/U
pRUVITLYxvQkwPMC/uWfgxuYY59gO1YodvGhlv3TM8LTyJ8ktbHcMBg5Roh6eJYAjrLmA/rLw6Vr
IoRqCihb0PLMqoRrLtPTl3MUNsgIEFm9A4xUPwZO5nDZkTuD+Pc8wVUvXGNcBtSgzmIlIMtTZ8Pj
+E7uG4jxUOA+uYWRUwxQ96oZZVTB3NhaqwFAnW4xrLCOL0VExbqivHFpCqd+y/z4q8by/ZkKjd1W
WGPl8QIZhkZnXaOUC0X3SVXDY0DqKmp1/4KcMPQqcHYhuIOxRNRMtA7qv6m53JttGq9QFjtDXcEn
8Kwtw+ZIzrvo79td5jbjxwdSwIVHNpVoNi6Ost0373brg4jvG+Y1mjT7wn8QULu9ICqRCNE8fk+S
bk2tzQsSz57V0Cj33Z7heBFDriZqXOhvW4+RspL7GjQEhuGvV9hmbSjjMOuI9RBKGwAfn5XyGCOu
bjukX7qsYCdIyAPj9IEm1z1oyDaAQOmdNPWbrfqrPr3S1Dq41jTm8BHNQdQTLwPh33x9+CWVd3LR
P7ZsPvgNcc9Ib5KfyRyoArsIkYS01AuRJtWkawvLIm5E+h3lQqNn1EySwC7+xIbQGpu1fRxQwgv2
FILgwMm8jSgTicnRcvm21+ppgvPql2SX91eycV6052tB2GJvU/8BXBU/7QMMeDyIYmqZMZTl8MzX
Ihv/h84oIAjfLkwUTmjHFH5pHVCksF97SFgxup+twC+N+7izv9OF6m1VixhVLHvUmfc3RVhzZI0t
vDbEmId8X0+puUpXnOqaqf33IqQndCygp6nqyYnwwR4CibjB2sgnZ47HhstQxqyHEM+Xz5krORd8
xNEfNlCpM0Qyy8LUUxBp8mvFtibC8fZkNpaGl7YstqvIf9alzR3LLkez0lco3w03diXi5wi6kt/e
bbXJpsAxW6AFcXzkvXMacho+Qx1aC81auaq3SUdweRSHVsiiL17tvAd1qAf/e5nCWjOqk+ecGaEQ
e2T9+qQYDRSB0qaRN+adby+NgBdoI22oFjneyPTQDSLbkMwKvvA/fGJLeJWg48rIBOpaJieSQw7v
/mh57+WzpCxQCN26Z56QWkjALXToVCSqe8+GGGS1qXV8h5muzt/SZ5TlvgGiyp8Nmkamlzxn7pmX
uT8YwoVKsZ++a6LSkGs27iVS4c8Ly3t+VNo454P4Pv108iU72kbD3c9ls64W7Q31hA/mGedK58Mh
KceChWilL8Y53uWg1QciKUtZNcqExo2oDqcpPsPQfcDt37qL8dKSi+tcuyF2ksSoxei6L+8I2jCG
r13SThfjUwOtVlVQOTPNiFgGoknOxnjqjHOgDs7xzQNLog5RxSgVG28jPW3ag9QUDs/OcJu8+xK4
SethKWv8sgGGSRT0AL4O13BOcKrQkQsB8RjQ9hKRhzIDRPAS+gcUClvmQGRahj60bWMRxcQ7ZA/G
ItooXuzqBPz+YCthyf14mYUpGQAwhfiVZEJ8tH/YcV42td7bdMjyg3MayQ6vJrfcsXCnifYvU5lV
nZjFEhdkGDpQUztTqljxz4df1/4FNOgUu+P2I4uiet/8a2BEGQ0+YX/Wdx0Bmo0TcDrAECl1IE/Q
zvEvEmp5HDBVTPS9pHP4sjv5K6m2C/UkEzoyTTUbuoU1FtIUAu+XhXwr4KR+FdHYsXTDY6JeYQdc
R8kI04nbyk13QPaHwt4BkWFh6JunQK+sdm9ezzH7jMAcX8EXXCZL1kfkL7qrT0TzvzYyAlK5iGIc
rrO0vc51UMLM23JApaTiB5Y+Kwek/zj765x55KoK6gsQ/HLw4aEoxuay0Exv7GgNtrVCvCQkAjna
fsgBSvdHjOBMpSoo7nNAFSXixTfI5pTE1wpKsj9uMDJLblHegsjczmZe7GSvAcdr64msZLsi05zK
H1kfYLqNAPK1oSYYh8lFPVoDjH9JJHOqaeUNgwvcjuRuBXNkgjOr6DkgSiqx16yH2d193e4JhpYT
zcpEp2HMnXYvhPwa9E6+fJA3KuC5xe+qHOw1Fzi33/SNK0jPlcIgWWJ0ghaR7SRIZfvcXa+KzSj+
ipqwz6uvgei261OY5MwOQ930QkhbXVCFxUpzZvjF3HBUf6qbhKYXW/kNcmo7JyT7UXkl4cm+f17r
fL3QhaUbpj/iqcJHkDGPflNIIqylgfD4z6H2ET+DcrONyGhsjOMoJKoa8IHiQxoU6/QCEUG5ciAU
DmSD6Tab7++7v4yzXgzcGYpAYDejWookd38sZlLPFhweXafLnT/h9Q2XHT+Mg9mW07CF0k+GDtKN
TCkjT+Fc9DyswVQ/riUULWteFzCVbdLhSBxtw5hbK4n6GtTEgNqakQvwGk9nLsgIQE6Y3RvDQXyY
wG9JAzrisjedhhimeON/0CSpqBcb6p0WBej9984es7zmNtrO2mC6Cn5LEJzclo7Fj6iNAYEdIAPa
CjJrd2cQwFRADRGLnivdQwlVCMg+60Lwzhx1l9mHUAnn8lp14/sNXupA3BlKWDcrXfAbVWtzjRNV
Skob4AudSQTEeAV0IAHJXBdHGWF4oa39PGT3AWZSkYWbMDtakxgFbDgYxn2hb5mRwn5PmOLz7x6Q
HM6sozYz3EtzF/KHsGcQppXzJzvMp39+RMxH/HsDlETGbPybhdmuxjHGPkvKzlKS4icUc+rEyu7G
yX7Z6veTCpiiqGVjaNFsW7IhTbUgpJBeUpfuETn56BFgEdc14AaReBcHMolZ4GR05yTQ/kDpkbTY
lEKx4goXasqV4cYaFISLygpvygA4e6flEp2RnvGXUKNkROqyxK6Y3ZSioJd/F5IBRiGEKbQLiZmG
5vPb3Gi1f9sEKaSVIKs2+I0RkUS5O4IGE8X0zQJcU85ESqK2woNDKWUvWjBrRv0bIDWWAdd0WqLT
Evuxoi+XdXOU1YE0gcBU3i4f3wmLAqYw4cLRxXZPSsVFurEKXTTrwUCICk8Hw29P+aWRM5KUAbP1
SyRMxFpkVrT6uSG/eLSZ4p4yALETwgJu/sW5rPz+4WYLlbDNQXOPfsGG7K5ZhqlSgLXJDxB2KX9L
//uKWxld/Kw+rpTcPAITbI4hTskPm/xB9eMbk8iEeP5IwkAfqEmpDbU61CFdHuE/NWlD7frDadmE
9EVrKPzo7ccbID6+ofOorrMSkSUWFGHqy+yas47c/DbQE9P48jpnzOwjDCiHHyDpaW8XEM0MxE8F
AfVPPTLxV7MlMbiqAyZx+I4FsMHpxkENrjXBEc7nWeqoSog942+8g5z7Paj3+ptg0dhMyptqttol
/NCfvTFsJt6d2tDS3txZB5E3/FEcDkWojcmTgox1HuZvcOsAtM22cx5mGb2GmCwno/ejb1vSgX9J
LXr+9E0P+JBrMDz7PMzgixa7WALqtsKpD9JQQ6X/MVDanqeSmbxuWlAnIinVbwoVFn2m8frb7OHz
vNQDrVKd+aRejQlw6gwIXCEtLZNnfVRU4+2sHpWKteMailfYh1f0R5p1DLQCL6pNzRXV0I9iIPAH
VAKe+fKFofUrnTZjagnnlXg1AQ4evrkXNJaMiuJjPC8qcTXijf9z28vMLVzv9gEPjxD+BZsn4VHf
9G8H6DPc8Z8jF02UD2DQPZi1MB+9kJuSIZ5xCOulFd79dZVaFTZl84OocZVUIHS3mf8t0IMV0fpT
/Y6sFYbss6Ah8EykZrtjtE/g8wVYzQyDjbAgco6lwBcOF3XEnrGA2YutwRu65sZlhW5MVfTO+LwZ
fG3mWyjms+EKwQt58PBsB2LY5MvX8pLVwEMBpaUidCHA0ycgpB67IqP83kUorntFZVAQa4TvQIOF
eGzxAWl0ZnbdiO7odhVicyG7Kl2eK2NKJx2Hg3Az2f8sn5mkKevdefwh0oEJfNt7GqmanAqWn+2R
+FcJTRZymgIxbdxWRqUtlyC1f6molv8W/S/nj9qbi5XWhBsuXHN8VDVW+UYpsIR48c/zbOgSrJ1P
dZqiyCArMQ0w7YY/reF4gqEOYo9v9ZrEVPrxpcoVCqoScNFLyLmta7eF7QkUNJoCnazFwVfJBedn
iCHxBkbkqFRAJwfal2Uft+4aXicEj8GWyF5e4NKNnqvJzXAHcBYn/Wac1K4yveKLYAP+FkD2LBg3
H441bAllQnDcYTYKB70nMI7bIIM6abk4INbXFVY1Brp5I8Ut/GX/vpyMjyk9ogVowfvCCHMaeL1y
ynkt5+99gqsSE1Uv3bDAwMTtf5ZIrB1+FExiquM7zlbr7O/f44/6PbO9HU+Po1W7nRcVq2Emv+CH
r4ci0/fGQk9qkJYD8L2Zj36KnYQ2xDqwuWbIKN6e7w/hHJkH7V72T8Pw3LXhb7NOZ9M9fjrYnBKU
Mdg6Gv8U3ZFOds/7/bGz075fyAPgYdNE7VcQZJP+03h7M2p54EnV3XCKB680qgIVtpMXXCbDLJRU
Bl1jOiYPiXdhcWF7x5G0jXWBQ21P5+s3zEUVJNxPQgDidrsouBgJvTBmX0PPggVBYzFdD/KJ7DNH
wvBe8Rmn/Fexh9GcxcBKYv08dTihO45YJ3RcTfcUxrHQfdwdBrjfJR9pGChY/3dsPtiRKqIYwG6a
CtUaC6NdC8oNRphXRV9m4LOdZsYJ/D+4jvOtvhZUBPtWqsrl4ogPjBmIUdUs1HYTIaiRQngxFhZV
4IDqSlIuMTVaHsdiDl5ZqL7jHVrvM15dK3Gzsb8qETBTRArHOtZgDHkU5VnXfV9kBCy3ZbALrm58
XrgBzqbnFTBVW8JZFtXkdrEgF6UsmVHhT6RaxtnJNYC+j2cKeIQiXCAgFADtxy9MBqtsjNZL+iDx
XDyiI+3PZWDRE3rwXAViQfAl4+UmQxQt8r6RTbiG/n/kNd6StgDtoG+dl3WF5LU9Ur7rF1KBpSAN
RLj4DR3XyZMjk7PuT9sLJarSoAYaz4YWd9mjvR4kI8L1qJGHNKmxFkhJIi1+FJljUQryBf6OoA8S
BpQa3zGT8ctxTVrS8C6HVqTmuTeLfoqkQD3J/jcbSt/IpChLurOQzEg8Rv2Y4pS8C4+pKeklhCjc
Mgtq6xVtGHO7A3wsIynhOTwj3UrVDpyESsgDIsHblNCHjOkVv0Xg6FqdBaz80noIQf1triRuvqda
fkKDos+F8m53tgxmOTC5hF1gY9Nw0G4ckKtsaOitAw9HbSVfkQGcioiQQf1LKtQCpL09mCPri4Vl
5sV7WankHSHKqchqln/RstTp+uGFIIjep/Ypl6xV14FAYTgSdqdXvsyYJ1qBB65KWMPlTDZudIDD
lP38UyhOT6hftUyClb9+RCVF4p5o0sjEBHe/pC325hBjuOI+SEHh/dvvW5BWUJLA9a+dTmpvpz+z
TZlJu02OOP9fOGl5NayB4Dw/PqTJE7nYOiZiuKp8wIOXVCvRfwAljUoAJy3yZr20BAU2ctXa6UJq
ULOGHsDZNMal4PmW/E5H33jY4KAcDVx+ebSaMtfoKkGJ+n6vEPpls6XtsSjqVBN4StHadWq5CahH
K5MxBED+ms+mCA/s/KXs+eI4eXOsLAhcgKPC1iZH6ryTnrBe9U9rFmIIdqexh+24PptJcY1fjYZe
3Ei9/Gry6d4Lv3luqQk/790hQWQH033VtOiQiQyjim9W+7Gh8jIiKu4cJMM4cPzE3YaMHSGi4W0c
wWve/+ld3ulMY6TT+ezCbMFIcwgjs3KpBttyDl61744LXgh0zhT/JT8jDj2RNyDAtBwcrnZTYfdc
rL9+Rqr3bLLBDveNAmRdiWoh2+HCTWz3G3udDnMGQ/SJNKPsZxJMv2FEF38ZTpHLNKQPHOO+Ddat
M537zAxUAPiTMjgY+9A9DCEmlDIBREu/BVjv6n8flk4vZwaaN3ECbwVUYWsj3yxx1w/WwTS1sZ6y
rOINN2KCOi8MzSFstQf7gO5P5P87kOh2fNy4hMqagtjUm3nS8z5RxgfkCSr38d3B31J1u4E0YrCi
sH/433aDAArKJfTJypgcZ5m6JYNnU7FguWXHLVTSSfLuq9RPMIdzQLLe8zKhCoh/zWnMZzUrubPV
0W0VDn7GBaZpXU3LRnqCBsu6QvjaUbDSjQa81poAw7utgghttdHrtbENS434/zSlLRORV2GYpG/H
ZMP9+yWNWY2ikDdjtU5/4onzUcmqV+zNwLKjge1IEQMuqLn9TVp9Q/zFDAH34jUpEeyfYlkdFNfj
9NGLj7UlTjMbpzNi6oCgIUy61XqqRzUpRuRi3rWZPkN/yyOCz0wa0/tG3zAlNdXxhil6H8rIFn0y
48wDFvbuSAul7Robz0LBELXGR5zgNpHhYtsxQBZbSy3Vo7jr+YZmeaS/0GqNg9nX0hZ+gyOC+Zjs
ZmsrvHO9FVzRcT38vPJR6rk5fdp5owQvGQIvrTxa5MmMC9toPbtsy/S0+W5d3TwHcWBIj3IJnsGt
AjtZfg6rkEhvXpD22JFsK/XrksSN6Dy7PmffYOVJ4EzEM2qjJ2HpOnimOD4vDI9wXcyw54W1poxR
tu6CBxhEHVT9PO4k5X/aYlPbOllqxXsYyYJIOoTy9LRHTswW+JQbnu6XyPgXeYr/Mvc+V76P3RNT
8i8LgKgWt7FxjbBMyZTHcJj2Ygpn6vmBlce5CyfiXKVYlCP9UcQpErknTYqwDpKyi3MLrVIJM4Jh
K2oNeXUhr0FLARd9ZRobmO6rcIQJBO1SUI4yuMxqaCet1g3IsXDvcoK5nXx833nkWWEsaRxjDv/p
P5AFeXnUSBKU6g/STfhKcl9mcbqKrrlSAFr53CGlbXbN37QFVkpN3OBartYfFv05JbSvT6gerwGS
T6bcR2WPwduKaowX+/DZVPCJSQ9dTGtgtL59KYTTdsLm0BqzB9v6AmPyoR+WgdUqMNASr+Jvguac
rnLNCtANNC9c5F30N+w8z64cr+oKgBxD72h6ZH1cURn7WWynCdUx2zB1Oj3dwDEoZbFOKiPDQLyP
cMSMWv8QXGMzXW7EOgE2xGR52kXewQV+F59QFjhWZBCrl5hVZUJa+gWmR8eAATg/wxa0ojApdtHq
KUW7s/lQnJw+PkpmNHAMfNZ62NKHm/heY3WhGbFyAhzL2hzhC6sfC9s6L0xtMzcgC5zwo6lvQGMG
mf6EMeLMvhf91nRhjirhxBWN6C3uh3sXqDFWuQ1IyEMoCz16TbWHN/X06KejliGBo//PPraqQaDr
HZrsbDVlejcuoPJ5B7U8WfG7HOtJhALxAYQvmIX809QL0ED/vWLNkaLNnI137+CvM1LXvER1mzOS
HaOsJES5iKcoYHn6bucSymx6LEfb0562zEoxGruwkYNzoEaGVeuDXJpyEjeuAIe9F7wS1Eg1KQbm
6g0hk1LyMdcf9RBXkozuvehT7ZBcONDCB5wyKEHAFJwAcY9foyYH6FdQ7qc7UPTSrQ2aygIZ6RP6
sjeiBTpiZqXXqWgEejaxg9e+s1AeRt+0FkcCge2P7UuWL56r03Y25pOO34zbVS+8Sft/Fj3QKtGv
xNUHodNpZ4RO8zwT8Dvua5eUsgECCufN4hnR5BDSLHMW2D3F5qPeOgqlcbQ7Ounbxh0YIkTXC1KY
d3ZTfUVqw5oJpEW6mcJJJgqqqmPeLOPv93n5VBNVIXbgnkjX8T4Ap+HyEcVf3BaHZq24Ui3N/Pei
BDHCNf6IWFJVGjBHJnw5Wz1DpDV39BnuDOFyZeGG5X1ix220R9FhYblUIWL/PiA3LRW5WXaaImgM
ZI7ZDyVSjFivHU8AvZnWWLlpMdyKfw9mgsrmqIsAxwtosXeb7VbJ80BUWUOi3HBkpWhzQsr+9Qwc
Z+Q/YjQaBTB6TwtkUnL8JWA8oqOO7aQxLmlkaz6ULlXBd9hqb1fvLBLRQ5GDQe0KENQXBMBLJO8h
bUzVCNYw7T1grm5MWRmHStbMBDC4dVTHCf0wcoiquao8kd64i++CI4W3gbTz6km9DdRtM2PaGQty
ZIAB8x389DkXJkEfAgG2diMFF5tzuucTckeCBeeBdrQeUiOur6oj8Ng5utWjtWkey/ildp34xF2l
jSXg+lLF9WRYlURZza7v25y2Mj5kyIgw6PZjjou9uGDwfbRn9x/9iyc4FZjCWamovSjs6YmUdq8q
03QOAC79YoORvIEDdZDMyKtWnn1eCSuronHI2bDGg/XXm/BesB2LWvCwpqvD0fceGg/gDkXyFaHq
QKDT6YrIsK4XK++tmoIAKvAcV7dgTMtnoK5hMpu2UbSaYqOQB6V6WcvQ3C/zI1EZQH0PGguN4DBR
gTJRcLgketDhZjdJgPiNtQjiY2R5HVjOyPRRHvaHkLIzUwStwSkNlieimMp9pvM40CpjYjLwJ9RW
WITCZmgql5I2cYt46Lv77E66htCfPBLPt3nKVjtOtHlicDTcRrKl6JmOTe5yTTOBP3OKA/W5B7x6
9IGjsWoIxmZw4iU5M06n1y2Je8LpgmzFMl8imSoGRcEq/aFvhixldIQM9DCXt+qyNtkjqlbs1HMX
hwXM9Jp1iRGrVB9njU561ksm9xlVJ2w+ascpFw3nV6OJPsAyVrKPChmqbTWUw0nLgbM9bXZxUH9N
FqfJ9x8Fi+gyqD9UUM9qwXRNGYWBZRkkfKm6ZgFUASw9tUtBBx7eKWUmJbvTQV9zeYn35ZbcI3/2
P43fsdaaF8DKKjrPDjFQD32vkDMHfgaQcOSIoNrtSPmL4soGxB20eSr3BOv4gWAynLd2ykBk+hi0
IRMjQ/5P4xu8MNCkYcx4ly6VI4CReYdfbc6H9cnq2WclMJh35+aPqRULbw1xEdlOhKT/AxbJWxGr
lF0yRkqQotcMtv52E6wdM15i7rEggrKHlGfcS29EDbzyyC3p3CTEj/cdgraA9mbjfXM7VPnu6MD1
IMtQGgic+wkEXQeerumYAO01LSzDFJVdm6qGdOfgOra79kbfx/Ipfy/YqAdFXyMquyN9d2Pbma48
5aXQOiIgmtb7NyIQ/STt9s+QnAZgz5XsGzOxxuzuyjnRNC+JTfLLuAqq8wBTo/FC03+C0z06l9i7
u+DTHPMpTobwqBvgND5MnkUB4EegGjRwkwDNax+f7Jypo3g3wRO/QOJMAAB/HkFkPJhc0uXUFWau
mrrF+AC7xa9bRWrx+GgLx+vunJTL7x8DZG8Kdf5SHs4eXhIzoNmeJxOwmgr4bkIJyB3SKzlUlBhB
Cujj+kv65x9kDMZv0YHq9hWoJjUr7bfuN3AmA4nzizV0+ONRfRy7dnWYzFaeZt1z45YaqWFvnG0V
HuKeAJiuh23nXSHFM6cjY00KytC20Bvsxhgo494PWPgGWEgQcfta9YBG0TUMBi1C6PAzsbUGHPCN
B0AdwGCcfGMxS2a8YWmL0N8EXbS2H7137nUvowKhY1C7fGmCI2j/BC8RIwrKpgaMvvarA3mzS9as
0iUyaquXWIOFjORwkAWe46xNgMrzAarH1r9ua2X4p/SCR/NFUyw278sJkGH2/h4P2Yrlw9oGAu0E
/40UPglAI1OKk+UI5b7D6fMTJvKAyknbrIqyx9QPepQkWnd+olaKks6aa26AGn8IK8xlvUUfx+eZ
A1mYG3UjUwnaU8R44Rh9t3RVayjUqnbcklv0NEavlFQIQ/n7LYbNPTUwd+a8araFBBJAaREipNtc
MM6ErqYFFNvNO49xf974ZulTR8FHNsvvCpyh+EvA7hQo37dXDfY9ZcHQ0yA6hyRQFBkCsDJuBRwG
jH53P9/az+T4FNB8H/Y5Ruw+XFGd+TGYmceB8yxfVZN/+dV/gQ6iE/DdXeIy1xA8V7sRRNfWqeut
DuRlz9yWt63/w+30TKm+bdrqw9YG4q1dLpvs6gEuQ/J/ti2F9Ds/g1gXQYtjBrdN6bbkjHJ2mtiJ
KuKt4lKWjMQCmNUDoQzfBzrUDS9rkvtFGYRBGDG2CBUon0Xl6VtrEe/sK26ziwiqOxUP5XBockfg
k/IblXKW7CjnX3JHV8sAjK+g6/3shR5FlFw6jcYAL8ng/AP9oEtBtuw/Crbq1xDipwto/NEHnLOk
gmfddMbEdtFiiVnbC5jZLvY/WGFhcinAoTGBWTv/yA5vK0xH8rQDg81TaJmuSrp6tlVjBAzMpbba
fpVYK+IDbiWBU2hVi5ysjWHxlKuuE9zmQxe2sdAQsShAzy9Jzoh+0uSl83T7cbq0bFASPg+umvXK
MMaYHZZ3Nz7ajK+65oYH5e3Wvdd7L99AJrovttYCBmjFsskk4ZPHf0EdhigazMjYcD/YWQa8naZ6
t3neukBz9nJUDnsiQKZUA5WuOHwcSReoEjWpPFM7PE1xZt1p6mSsKBNFGscVDmYl2RJqySrBXRj2
yGVDh3ZjWBSQzvCe7/pQU7Me4WtlePA8G1BmDz7YIkQBiqvI1d5v8EVMYl0kwtKjTNMcAelcxhjY
GtGJ99tazVedQr1pgEwiM2dYk/vaGi+HlkIeh1fXyRXbbOvMFvlcUkde3h/cg1il4kxeh6rHtgfd
l09Cyrtw+BW3ZoqY5qqLX8+duLhHuLnQMa2w5FqQzf5suplmhoSmopDZplUdmOh11LtZ+93mlXrr
2obHbLVbTVgAgZI346JYzkcbJMlcXCzswA2DzXdsdqewALBU1Y8ajq3ofyaE7ejqokdGUX1SwaNL
ToImXZuEupCJZRvXcJq9VpTl9zYC9WJwzKGFblbu2zy0axB38V9g6yza+PCToZKzxFTHkyFT+7ua
MFUebRwuf2zsMFFqSOoADuePTn7gRsKAMhhcj5g1Uq/MMPfi9/hzY4Mea4fYJDOpPrw1ak1Q9Io2
21RQhj4SvKDLYoQ7WvGnbxuQ+CwJlLEMvtX2hgdUrdJsBKQdq4/tSIBFz0qIGSutA/3/GCCeT7ho
fxzwQdhlfBfdDcg4Agpsd28lbuRgcWVX51TZimnkRioYWXjeJnkhMW8fobeM5r9dtK3pe6BzgzNr
YtZKSCNtHTBw0Ean3u2IYcksZ1vuMA3/E2OB5c9mZ0PjvBmANwEcGSwjvFcIhANfh5zN4dA5gvq2
wNeK8Kq1YtBahuGZct05N0wksnRxnd0uCa1HbR2ea++4byDkBXKbjyNCp7UxETZ+8m+TfIZQJTE6
LLUIxyd6jIEQjLil7vBt/UiiLTwKlTfgGS5DQ+9xSKkaDC97C4ZS6YZgoCQ5UvPKdFfOilq88jIf
a63k25ItjiwR5psGBmite2/4lILOdw+uAcd/HJtZaTXTJAhXYbhb24xi9tt/whXpGb4xiQn/sAoT
8BPqxxTtSRVfkRiywBbj4W6AkBcZQ23QVjlnGQvnd/cJhUm2syyoImYwB941Y9oCjQY8w4QrzxrP
zZuoSn+qb27cdgFWRNotqZVnEwbUtDK4v7SEg+Ct+kDAoDTH/Ik/GgwBO9ABDfp7iy+I3sLL5aJT
/xAJqC0V1LX61ofRlZw054SkY4W+paApKjx2ce26bG4NvdIeeZSaPdBljmEDpA06pkgqLZaoyIg8
paeFL0tcR/rUyC8rFjZdHZ7DiSa+pgdYXOfcJ6Xq4DqxFSFMyziG/uq1dyBuO7Lamb/YJoc5Cbdb
xWD5rvTA0Lurbu/KJmHCylN3/oXyFmJGb3vzLasJavly1hofxQ+KgbJ+Do3JQHYF5mnoXnJT1JgP
Xq4QDsREGR7r0DO4WSwivEAmD5EpBb8IUDnbVx9d4rgKkAm7ZAwHFGxfWMrL0HiiKXDjzKAeubB4
RmjhtT4ACWIH1U6+OZLSsdLoihwFQvDLgHoEBNGeyDBBV5UPNx6BxttojzyXNLNkFv7Unc12u5LO
BwdcMfMe+JU1hUJ44PiakBnH8OgavcsQw4VAdS2792ymc8Mil9A9fuAaChFhZ+Y9I6TQpJ+jr7Wh
9/hSmobs95v6dC9dLnGtTbozE6vDCzdqRo7BS1XjSTby6fw6d4Tr2GrnaZ5WFGYLAY0AsSTB6Uo4
5BtYcZQtXiswXKGR+W5sAWGwolOuQgFuL2vTn+Ht8Utob01giV2HWEUuatSZJV0CARDbmOEp8sGa
qU3WuaIY2AXF/76qLah+0cmOXfSIE/oZDMUeKZI6FfxHGAnTj1KdJl5GI4u8O6LXZJwQjnVOs8RI
aIx3LdVEM0nYit4StqBbwgSuYRcjO2+zltVzmR7hJ+S/XyJE879WpF8trJKzI2Uf4v/UgSX35l6L
BcAtHgDJwUkLdTPJpOWe2e+3J4yd2x9dUwaYYzROt8qudqBuoaKnHpxHildMtc0orQllPmLDGR+g
eU1mPpmWMXrgpwgCZb5AB9+W2yndyO9WI55x4TCmrv5tHKnKIINzbpQOekhpAEKV9MZCHJuj4uWy
9PXCuBeX+SeDtk/TrlmSJOV3YT07D3YSexYbSRbX6TNUQzPtm+rlnST+cr79L1cPdJ3ra0OghgBv
dMhP/00wHzI+Kxo1plN43H9KxDdPRvDP5VwlCB5RBIdUO855RVoC6wozSbrAI06GGzIxNHHKqKEY
pqnbX8/6TF2sGwFTjhvyla8ALmQd8f0XUX+QPpqsBI428snEoyyGWUgqhODmPFfAgD+rLhpiwAJL
hogRDwVqMEjBEAlHOQkWDIQ4hFMHw/km/jXgiit7Dbi/jP7/bcQkNcCiggaej2UU+bafXnQXebkh
hEnw3GDMGVWp6a9mmHT35RpP1r7ibPZKBhkJUGMR9OA3Lm9qdlWNsKMkvC4XSOoHT/kjAVxSqLuN
IMTpKO4ruYdoD/Sb1CrZj2LwMtP5oFpdYqnsmPj6b7DL+FCt0E/Npme8sQUSiQRV0F6UcoDPdyiN
BwkGtT8jdXdqg1AvKLNssjCm7kYnzyTvLsjbjip6f1RIH0LoSoQ6guoIA4oE7tebg9FdMe2XGmDx
vE6uoRKNketurHKpmYK/acziuaFuGaC7B0m6eOdarZAEWGVeMWAVJEIhTxBt8MdSn+eK8mKHFa+G
9AqsPEst9xqEgAnV7hqIWxOhiJDmaQt2W6L3R4I9AmuoXWGTwQzFAiX6omTZRaX1qfSvVKNnsUN+
82qIOlZWHUteTsH+A9PntQxrmnf28ptYQUVEaDUfgB1Ee8SHWsLl4djAwsVWVg+vwtiGkbP+9aqs
9T80PjpgzW34TIF3f2BE7vSyH/WaJcPZWOZRF9Sez88p5ninIbziCdMdohuOwRUuTn5Hj9r3QQPF
0quvdTsZf/Se3zOFIplcj0tJkmWhu4Mlv2hFa78sKSUFQBPoukySFmowHOrrZr0fpMzlXEOdE/aV
u7JxPQG5El/AM40NUbXuaoPrySwIWbwZ2z0/RSv4a/VCZVEOPuj5e0R5YAXLE4pctRDlfnnA8Hvy
SwHTZ6VKUVWiPY86Ejc3DJ6ihwWWP/ARPt4n0Cs5bkANYOhsLxDECRDbMZaTCNKYXRtmnOieGLQg
/rNuX1FVQwFdrI33Gs/7mWHiXf+AFrYDwZpC1OctY5Ahc4HS79+1GJOz17G2ymCB4UZM7WQZyXmK
/GfNDCS45Cw956INRdsS0o6TUzvQPUEGsqpooV6l7blaKbPfuF1tjB0hqG6mYFQwekH4mNnW2iS8
+LE71ALs3/3wqqTNh7wbgDEI97oacyyltlMgsS96fwKFa6KrjCGu5ni942Iz2+LChngbBSzRKc/K
Hgu/3BUhCZTG5C4HfQRdSUN6iGxMfEdORn7bas5YFZ+ZwHuz/mGBZ44g9f5aDzMFIanMMBhAIBE8
oOMvJ0xjKTse1beJj3e5lJfXIb1uL72AQjMCJQmI9kHzKK+YcISXvns7f+RQVFbXjpnuUrIZQKwD
krgeHWOfhK5s43ZlUJVynE5vyYM6Sxc8eoqRTY5HMsGukW6sD2QZW+4W/GKn0nxYDIFgyfU2/7ss
6FrmqWkz5XestOSrf6bD6yu7dmYEaHrpGa8NOOpMtHo+nqLA17n4OT8X9nTjczvpe7ZARULIG2Rd
ZcR+k+dx6XFe3NJCBxWmEY2uMBlyJgJyJhhjvs2STViXoFmof5oNO/GTg6W4IlVKEAxa131Th4lU
OZTTpaM+ifVbALUFOWRw93REMYqGwNkrwG/M+vMpMuV5aKZA3NlPbO6+04edAMK/8I/71HKUJe3H
wGpZ3bRQyVGu5jYiDIP0+2DFh7sPntAQyoi9BjBVT2qN8BOHMeTKZ6pR/jp+HAZvv7jynM8rPNLS
/qfRJAeERW1R/Tl1KqCTRl17F7Y2jUVreOqrldEXAjBpt8oiGhkhmM1a5hcuyZ/v/uLqnxNol1LU
YWCtm8O5EXN0GH16gwIBxaDgsNu+JwbttnuqXFtUVDMAAUHz7CMq5jRLLo9X7uPav2c5gGt7ETtp
jE2VJ0UKwxEGXJr33x6+c76CuTtUDjd00VjvUUGL3nRtujYsZnmeKbSkp1T3zqpji+AEz0cxOzW5
KHF7YzfQF9tFxnl1qd3Mx0bkXa0Lvb2LPp7WmiXs9176vPjDES+zkVVVAIxIgJM4kUId+fm1hZcC
ifQfArqNSMqME+PUd9oJ8qDMGqxUR4C9IaRa4fHIb4c7ICJ4TDSiO1NI+9GrtOzhIIrWhVqNIH0K
Hf+FgktwQHC730gQTjXqkEnAwP6FXpPMzcVFIcWRBmNzlZ/f7DJSqnu0bZRYLhowVPbTSikjfxhW
P6tzN1rHeKE3/Orx9XGEJ8xfkJi6gL9mEOj/AydxAifYvoarh95BIH9hpUHOp5BBuz9io/IugxOE
O/CiF+o5HMdgq0SspVmSXfwnxoXKA7rah2L7jChC/HFMRip4ufx4zhSU7doqAMIL2hK3QDhHFuXl
kSdc5sEKMfz+9p9Ko+MIKoezPBf7JjLFZUVixHbxzv9q75LnChoNYLOR9X6Dtp3taS9cxnb8h3Ze
B2oq3UpZ8gJgcH85noVqEg9lmfUEalRyTTGUhFXIMBHs3SLoRI/mcx2DhqcQ1ahsq3GF7ZEwj/rg
tclbLSxN0RdUKlnVkTNIza5nyCBZYlw2HyouYDrCIU98zkz1Yb41AIYXDkmTYmmzmY5jOdqj0DEm
adG7G10iIBtnGx32gMLNEP2LKOswLSotFMMdatR83Ltm7LeC1st3kMS2vmGqd2M5uKIYkocSgm7g
1VER4JGNR5fSAYeFaEa3ydz6djgpUFcbd55rMKxkfckU6PkeP/tmgTEPwGAeHSUOPgEDAPPZC1cZ
YncYMwWgOnhg2TnxmG/s6Vf1xsAjCPHIWCAP/yRMrl7rksqkDIzUKEyUNDix5xN+NbYvui56LSKm
Ho7efx+W8JJ61qLWcQwZc0Ue4AO3Qz/mP1E1+mWNOOyavCs4VFF1w2QAV/CHDHBarhc2D9Yhyonv
qNiebYodheYmqPyWiDc9AjZsKvYUHWxoMref2za4vgsTAK8TRxCuGjdPQC9NDUvVeeLDIf5DXdu0
fngwy9aWpbQjyMB4Y/v9Omsut78cKxbrUwta/1MVQIHI/my7GaXsEC7dWQmM7BIuXNLmFQmTMClY
bAM8YnN13NS2XMC/hIGoR0bVT9RT4wJOWCB0CzkiN2tzCGuvGvImkWjj3EpjzO11wX2MWwolb9/h
X6KLjWuhj8qxDb3R2+wwJHPp0O0enZMVgvYRiuJpnnXrSiKhR8hzHbRBby7DAvN3yh5gNazO3xJl
qlJYKAF5qhXiOmPThdAOLnsK2ZOTlxFXOYQzcIbnZqanWBQ/U5tDOQhA3BYQiOMGQ0i1qnqPIuF7
KOzMWebGpvaLMQeO8htyoxKIPbBsqO5PYLMRqbiaf5IWI/SVIRhWPlfMyXwWr0pWYlF5ae2cCnPp
RXpc62AnRGmPUraBIo/VLVzQZDWXQyyNc3PkVHux+4Ci+5Aajw9LDRYPYJueFv3vTAtF4BIkio1d
xpl2pWMedM12PVrRc0iJHoPkT4dqQvu2I0VNiecktd/Euvo8W03f9i1/vwhYPF994hDHGVzYQhPb
Gd1tKXB7tohfuhsKmKxOTlCtpdcD9lVrwoPDAglTLSfYJseP9A7E5nEjcvhYbbiLCqqRS/N45m8/
ip5d9YPxPVKkChfZMLvV4rF8aJOJQA6HGyvL4LWRt/Uh0laMlblm9arvbdCroQGk/HO48R1BqNqg
soIBbxKnD2Ltxi/7Rg1wrVuYBsBCvgihCGsa9eV3BPuGlQrtdlSP2+OLFzrivZIqqthIw8zl+ZgJ
/Zx2BWC4AN50j2oZnY5FF+FVD1olJzqNFtr0iDTC6cnFZQd46YJCkFhVMHa9xp10OJSMv4vxzpFs
7jU3oReKBv0A7uPZrxc2gbyS5RfOnnhBLXaL7GXqokEnLO5fulJkFDoUrhmOWAYvCZJpVh5obkGA
WbWoz1Aecf31XUivlohYZ4ws9fZM9Oki/x910KNgQBWql3i2MHeVzGcoKuanhJWtrC8vJmh2P//5
Lhf8BKu7uVLpjUf18mYIHJf4oireLNJQUfC+P9EHYj+rbIsmeXrHT08uxLDP0pKI44I68V1ZFMia
rNXcZUcGKYIjzfgUWRtoTo7RXKUdI7L0yrD6Nc9VFBohWo49pdEJ/N4pobMU+0/3L24GqWDzQf0K
hqfS4QWZ87GpVw7jBSU/FbI2sE+ttQKCF79A766wmBI+JmWQV7s5K3k5F7fFgYW+KMyhtN0hkp/w
4sqE8IYANQkkqUiX53qSiBrntlHeOWsMwMIvSwEZ+wHZjOmWLtAVsUkTl9qxiAwrnQGXMleAKlfU
DZYV+MptEsVG0ne6P1Q8OjMDlQzsaTp6rDcIth8HmX7iU4cW3h5633iRodjMQYHmkTFxU7aZ3+aq
KTi+qjizEQpApT3bTPXc7Qays6vKdDqJRoZMi40ttealZBWPGSP/5A3DmfoMDqIbamWVfI7TwBPm
kSmKxe35S3uPimwbNKT9qJLK3izVY563H7awoI4eTJhf+n53EbP/e4s1RiGileXLgLKUCLcSTaCs
cE37E1zfc/a5OMkSzbZdYdSOxGRMmPnte6CypZJdRbWwj575yrU0oWxy/qVqtRt5iGYgifMeZaXQ
xNgnGRi9oL5/GcW11geMCax87HTvAXIg0pTPfJOLm+Mq6OjPkGfLZimwL5M1BQ8jWl9gveaQ8kZi
TxZtUom3bLmBYyfJepV+CgHvrD0gRoRntLWbzAuHBdZmXIEQKUR9MamKfD0pILpgxk2CXqyur4Cn
khcINEOLf1d8WJpRXE4bkJIcEosaKL1/pKrq3NFE9aE/FRCbVh+WsyuuaR2r2Of16k1Rn/mnRzVl
P10WRS+KDfklNPdu8ObhEUrrNfZAOUnqy/eXpsWIkeDw7Q5baPd7mgme2JqZ8MQk6maU35fO70zI
djq8LydXnXBETDh5OX9irHUEKfTQN6Phu7hTP8x9H/1FhxMOjZ4B9o7cvOXZc7+c6RVCffZdwSCP
m+8AmeJaBwkZssRoXOlOTXNSf3CqjgB3gB/eo8UKP7NL9nst6BUf8smGLCSZVOwwTCCguwFWuJKe
d27x55HHK2cQme46KqGSTFasMwoCkC71Uf9Lt+/X49Omx2u9zxr1wRQMi+WOCIRvp/AxHm7o+asn
TXljejrnU+7n0yp8pOw1/JWaInxiLKb9uc/R5UcNKNCKo+pnZTtkRMDQfCYcBLU5cpYs9ZVcfW2j
iIY/uap7qX9bLTp1RwZNLvEW1t0lHc0ZaaL/eRJdd+vy4gfinjqYPv/9IBn8bZ4CCgsKWpBS3gvm
EHqiC7MvPyPHV6lTz6104gl25ATMPtL6xK7K97+bHhqD5uuWqN1opneRGFy/6Rgs2RQOjGzYFU0B
8vjZ/DQFxE0kD94J1AGPwT1Okh6N/FKiACaFytEejqQ55sOcer4CwvXXAHfJ0HXgcBr/EmbzJ/eK
+XMdWAb8wyhUNzRzkiaUMTBdXtr+DiA9E+DFZybNlPA+w4rjBMtNfKHzfSKe9T0onAwnjVMa5Y0d
WVmXj373/YEKDhn2E14hoZWkNfycetCKpmjMKDn6OGTKt9VIc4ftfgWAl2T8nGcOlDAOxihtAyYU
K+GorWT7Xwsk1nGH5GJZVHwVcI+foMsfLIddN1tw3v2xa48VNYA3zxX1XHhiao9+L6hOhl+PLm4J
FwAGJEQtIrcPll/WWsJ4sdpZAS1Ml7i27MZqCb+5WZ9aR+QsegD824sRGqIF1tLeXE8GvP1qdybj
1iLkWCOCZRPlEVE2RWAODdBYZ72LTC7REqKXDXURY5zLlSgARkN5wVuLF8DWqRVEGsxBkwK8tjua
aVsK5PGd+Mw/9vUrIGdHZkdJDpcqRvrSRNVCbd5Uoi9rCCc2UyLiIAcXvBar3p48KEYC9Qhz7Sfm
g1SN6Frw7H/Tn5A/k2LHrv3MZC6URutnCEwom2rxqVPtaBi7SAEWRJe5PtEwhuryy+diFRRuIaAF
xa22d67JfkhvrZ9IvetanU4yVGcPZ0kw1KtxRW6QQWRkFqr0zMD+Z/Ycvrvvya4dSLXB7vr0aRMd
yl2uWlEEvdvRQrV2m6+aKpRiTqpgdw8VPivLiBF+iC5MLyGH/aUR2PpIGPlWgrNNAM8BQqc586jS
Fk9xHcUui+qrbRdS4VnSTP3xXoVyj5q9F/lJCJ9zS95GkU2E3MSBAdOsVQFKcv4xy1kvZ/X1jxpI
JDSlbrf4TpZ9Sx9VrPoFfWnpG0n/PWDs9a0tiH3JXunGS2Sd7re4QSlD4UeTW4nmwt7SDjqAI4vJ
2IvDEFa4dCVbd2eRgWwEV+V9ezAhw8px1Gw9C1j0mX/OG1dk0EcOhh6BAFey0YRQICx8Pc69iUvn
HiZQxwN4RWfR4io7TdAkAJyiveRvs5y7ooWwlWT1weN0bzbGTkJYcQ1EFUYj2zMode4JuFiPJXGW
p8kcXHyyQncjtlWOIVo7AHdiUZebRxQWTsp5BOz9+1bEXVr/8B3eIO196H039gh47NxSFjVf76mE
0w3uxY2g4ofJL8Nl8raWG0ueEaIXvxW1c19alp3yrSXZ2wNha3QcUPDu78PaBBGHwaRo4ttdk/B1
wWNPlStDXwymoQu7/kSt8EAEIpsd95/bw5cuVO+KNsr8ZzESASwN8g53+1paExXE62dWGypa2bjX
1BlKPv1K4dH4UGlG7Zn+cely2/qx+ZRifFbuY4rhOj5C/BxOMmqiUZxLMFqe6e5KUfW+mZQJpYQQ
qAkudAyKYKxkZZSVF6n3FZmJcCrQT7PjB849CKxzgfKg74btL/ogvXRb6fzWxKaO7Enc2fAWh5Hw
r8nFTWW1KLOx9jOnlN2C0nCWjacyba5ZeI6NifVbs+T+Nl06Lpopfu6IfN08mzFNsJvu+VcirXOJ
XlqHAKGScVO4aCS1HZ+rtHhY6LXpeNmOmqtemLOg5NpuMXp3Tj5wUbUKYed++x//bP/CAADCVxJl
7aelyKosZsHErWWCWEzQ/cDdHiSX2MALDDpGXegLXH2Fbz5bnYIdrBlRdeTLSAnAi8z8+QZaEAfP
SRWHVNHaEGnczKtCxH0cF9II/shY+WDBlRfLo9/G9FYfO7lwiR3p+ThKgg8qjXhhzJUn0T+oNAaW
a9BeBKgc2yuq/TwdSsDDqZQuSkTjEvRMhGdwkn6d6veBhj+AHoTnJQp2w+F9c0bxBOP0X5ouG2Zv
Z7FKtc8GD8Ld4YJkZwzkK9O3FbmHgJ6tR+lxgnwe4Q4U0sfeokkvg6DYJ78kpBDAmvDncPcKGTq2
6i/UEA/u2D1ORXZj2iUUVPtjnOHBAronk44uUaHIVluAVic18Cq5gbPMEG/kAcmSH2cijhxeKcLU
8vMVrmtw/HhMa3JzcNlIatd62mTJ5eVaKc+ls3ExElhwakT3YiInJEmXdQztb3nUpkEoNBj7zQyk
SSBGllKRo6Kn2mdsBCq2YdChlLLWonZMeWcNiAA88qseA172i0CmZInSTYUIgc/43skVCATjXp/K
3jVaAZI/FktWFq/oFuB8xw2VlpFrmZy3WjHqIN3TBGsF6fvdl6xjdnCC5d23L1NxGS+cYKIGT/Jv
QMOEa6xg7FnT2NTuW5T9AHyRLsza0D0m3BF7omTDNkiL/BDTXUOazjMKx7Oc3T/AHMjfAB+CLGKL
msEUleZqEdz/MkQVcgA9jJJo/ckp3hLwuqVTlXwycWg8ULC1YPviy5WzREDvWnOn5ML2XUf948Mk
ndgW81EHot+UvEN/kME/73gyNU+AaeVIeTgeUZwixoJG2ZrpDDLn5hyGFPJUBVm1tsfwQCBBPHVj
bH/pwdACJgyzkY2HqUp/4IMBTM0rfGPexFTnAqbdPg4nk385OzJaKEVeu/+WdsceGcXaayYu2s4X
6D/zO7mNp2WlCFPnjCADdoZC2EY02h3qibGdTneBhLWgXW08Mjc2v2oK/yiS+HT7tQFmC+ZWf6Hf
7Wnb43Ifl24BXu9W1JdRpbqusUPI9gWhgpkkeF0pHCCiM/aYT8FjuvaiMpGcR6ewdIn8LRjnOjKz
fG/atr8dBhi1NiNZuQrYKqeuWoBgDT+eNHRMAwC5moCIRxpQybI8Da1wbr40cnLGHPbphPSAwIE9
4zkVBosF/uZIvQMnW8iSGcZPtRCEPCPIwzMSYxyfKzNw+1cyE3A1f59Gduak/ID40xYgKDj9Br3n
eEgJV9ANm01O/zkqM3oWj4IFRe3Mqfo0LOfPxJwLchGqj5sWwUnJ0XOjOhHmvyjqSWkRpqUGC3Zi
G01bLa/E2NxXhn50IVgaHbCvM9YcOsj3ddGbiiiicnbOJZxAp0scwk1CpctRs/fMhnI0eCYMVmDE
Pmhcy96MWn0RT5pd3bXQrNTIiYDmcVi7a8iRdXvLnQb5PolX+CtAqloG5VTvN9oKqT/acMfwtTXo
IGSqK7ddmpkLrRQ87ryJJEKz9bHKmKEsqP8Ygk1XtQXZJeqVFiGF0QP+YRJWdkljoJlWqATppNJU
ZgpWVeYnCFxV2knoh8UZYPYQVnXwSYGfsi3+ZoggiBknp6h6tzepcuwWoU/F/eTyWjRSJPMqrXy5
Piqb1T8vpAHimkbRlcb2nXtRwZ7Yy3058GQceeQ0VBnl61t1y5TyJg4kf9j3213UtEFi6efv9HXU
pTTxda+LQCav6rUm1C1pc3/ZIEoyutjFejwnZRKWXsbUtbX5c9olXjT+hGC+8PwEecDRbo8aRi81
MrUq64hFp+Dt44BY7DHf0L5NZCzM8T/g3YouP//4nQvCVH4QbU5cKa+pUeMr4Lci+GrprQ44XtIO
l0/sImLq6qyikPNPSg3wl1KEkX04z/hz71UU+EFI1kxYAHw1WlvtYVipqFUbi7AIs1ww6J3eQZYS
OudSLq6+tRrOTBbySbXaHtwIzqaazBh9bNIHa5u1eMtu2Cq7296uAYrVy8nrt6UyOdxq+GJri65r
Nesow4yU2cpLnPNxuESpPywHd0NvM++OQ59P/Fnp6l37W6fcabWgRiYd1QQV6woLXe3CuqglLhjI
G56PrsrFbB6PvfjR5uYWvFtjIa88g8m7K9RA4D7aJojZBHVCt3mWJSpDqzyvRbaIM1XQ/4QTawxT
oInQ+MdkNwLuC7ElXJ3fxoX3OIJJbURaxiGhA3fewCV7vwKBlKGJX1MO1cV8SILSUsM52qesI1Vd
YoG/WT17IRDgSU49fDBZdyIv8XHTl7yZqaRz7PtKbNZnVF27AEVIXLrJKON7MiwOrenkZMfK1Du5
wTmVdFO0BJjJYZtIyOceYyAzLGlP0QDNUCZmlgXk8UgowJoUsIxR6i1UzdLEG8dBd70lIsk5oUXU
d9WrQyuvaQQr5DDUkM6OEfKyU29Ht35d9+mq1a2KQzdP2TQybhNpTn7ilmQLUiDA4nTZ9KzSxnA9
WP0yokMKDyBFBfOf4XPdAnEZyev3WH9QYIuA2PIUIRSe+OCMjcnqKXuvkbEzJ816oFy3EWZy6AYp
LVpb0NIG1qsErWmUOYAURqEi/SIy3aG3INh5KNWuliu67SdJXmtc2arwKBvRDabsk6ZPxA2yDDgh
ALk+0gPTyNdeb0Qe7urhR+tV2K0stUkFuqNKY/N0zDvLuxMbuW6djYgo0Zj8Q54HePy+iwLj8QUF
GPuP3U3u2T+avCzmO79KLjStGUC7RZu6RuP5fc/0LSJRCWmFRiT32mP9d9oOJiAyPJd+k7uEF0u+
X9VotUpIBOnawm3SLVHm70j1JxzJ0a7S9vVNfeIAqya9bQIj/FQnGZx5UELz+M+9gfKIc33Zd7m5
9L84W5+4zKCiYKxoMpMbooKEXoEF2/901ptUOhIM80+fDQbKdtRPbpk6oPM26rfud203/XnZC5tz
FnDgnlz5ThRzWF6Ac9FMaB92Gmj1IpbGtj1f/iUG5mzbIPVpW/7w/ohG5pvLt1m4AdxLrGjbwqvz
yBQjJBXGTmBymkZ7ON61201WLws1CAI+Fd4XH2cxw3D7ljEoZgsPhPv1gNJn01Eeu1dxZOOsl2HO
U+AlK8VP1R3oK/MRKnPw/0vCIxdte7XdSnkn0M2a2IOA2Qjl+L8wW5Z30M9CkXVjUkKxZX3kOcYb
ajKhDl6QQtTgRQm4TMzbgGFyzc8KckOViOqhm5OcdWasHqZ5jTUGT9OcArew5bUquCJjeUInVR6b
hFEnqzHPOpAiyFifIs72bmNIYL7k8DPdSRtMOC+Su6BTVm5k75DY1nix4i4R4jDRthLKqGuO6VbR
5rur6CsHf9vzIv8CR7Hqun8FEPz/PETKRkDnrrTKD52ezmjxkGQFxN1l6m8jnk3UDTeDYsmZMFJh
ofr8XXQxz4T6eYimBFnRfY8sj6gTJy6PVys0YFjm/yv2+V7mW49BPidmn4JY3k1zQDVZ1eCdZ20Y
Vzgvp+YhEvPLzpy63NAGE+HOnsi0WUs30OTQ7BFTHsDlwN0yoNjtKsflEsq/wkU6hyM2BhDphCXQ
wxFnTViRoaVTDAhECZQ4DIo0ShyAy9J+QfHIDmzOje3JDm+HDpaFXtQKX+HtgAqFbgaP1HQVNh2z
00eqdYb0/3N8Dx4B1gNSiGgl9Afcx6qA54t87C36Ymz1SnY43Eb53aG8LoZf3DkoK8unlATiC+Tj
i2Aqkgno4E8Xz44XZmK8iNd8uHtv/HVPIXPt7D/XujvOxHnHmyySykndNp0XoeHAhgzwwi/Eh8Vt
cSBaf71gBer1XBHT3/Y8nQfwOoKI1tM8yu9aNMeHa4R9zbOYbdY9Y52O8HBAfNOGT5Er41wWQ0qV
x3fR/VZ+J0zryImgYPrPO5Z0WQKQChvfrcKdmxxRUWK8VL2Nao5V7uLm/ziivgwucKZRUAfcokBf
UGxs+4BhE3HzPSizRzKKw9Fh86WAEnLR2xmdULJvIDxlZYbHwXLg7lzXfS+9sCbrSc78HdEzbWa2
TFJ2n2IajHD9Efa4x/P4u2jYkxt7NJRj7S1dEvyxNlC0UsPfCSbxaarjJy90bHFavf9j1Bwd+eLs
4lULuHKPh38kQW3LEGBz+A6lkBfJQW8kWmNq49kWdldSmiZwwC8RTeQ1dJSqH6rQpdSyKUO/2LhZ
ihu7fzR85ngkiWDkMuwsK7/Jc1NjUXPE9odbRq6H/00wz9RVcg/u37KkvZAjSE9JM/mi8iBKAZFk
sQPiP6VBEw1Dfw2Pt7HTBlowVY9kxXI6j7LeTjJ4YAEQoKltj8fAAjZ/E6zIqELFJokd+Bfj+RFE
Fm0Dh8dau2LK4ikL9/i2vHZqJqYDwCyrzwu3wtjwFhjwKyHNOM9YeRt9xPlB2lm8HzbL4Hlvvity
LDxhTT++d6AtvCOShl/cdQkoDRNcqrkVP6Ng34Gay5Py+u2tBwxFeaRWpQw1V0JODetjiGtR5HlJ
qQ6iRyqPaJWcpk6Xww97JAOump9narrY88M9UwzQawBtaUG/bdhqi1ZLVG4jdk3wP8wxtfjEdQR8
B3QLaNLJy6kpbm6f36+Rvwctg16Hk8+8vgxV5wPgtLFPZS35E1nVSePf4dTPgCE6QkPf6E1AzWpD
ROidwiiZhNe1y1374egPK2/t+AwAcogSmNRUwMENlVYdII+0bBfYjT1Cvz0Pf0ys1VNYVGOzBN2i
QgQASdQdJgfW/FDB2ccSWHCQ2cNXtVKCVEdwKRE0+Bs/dcjl8BQVSoKQ4OuhiTlbUtI0X8hHSn6z
4jOSjQ4hjogeCbyHi09gy2Pe/dp1bhxrDPT1xzuv/H8R3k7JTiLBKyEaG3hw5R2/rZ6h9Ni04Y0m
vV/q+45bIaM7czhVg7OMOwYlAQx0e8LXpq1lI9gzPEY7akNAdvc4lf+L6wga3QcBIqKc9/9u6rhV
s6ZhxayfAlaTgezPK4OyDO3RIRUCcYV3bqkTDkIKiS/2MqQurI7MTdac9+E8ec3ZwwLHL4D+5zyV
lW7B1eNAdiZAAolLNmKvB/thkRzIhPLoThBxB7qEWuvQ1yO8hcI9+MAeNivJmGctpS4iYMrLNeB8
pBvqTP5GWXW4iqagbILPesItvH5W37j9CbhESaYfQ4wdOX3/Frj204+zxYcNibPyYHB9qxnR8eSY
RHbfx5Nn6KP6LTru+s0byw9DoKokWRxuqgwx1m19qOfa1kMCeP3vCOqDnU4KAxungAz/551yMmcZ
q/0wqFv06IsFfSkzXXvN64nE2b5YwosKOeyih5aW9ig9vO4ppmkg6sGX71Ov3Abr4w660IotWyxU
wW8r1Rgv7kSsiQVV8U8fCYEGP4mJVQZgRaQUQDs+abJ19PexbwvhFJxO6QcSVmvanBa8rnyPw59H
TjOebuZn5tZlf+ddYfLdW9+n4WAIcn5ygSXVLdXDYBbEj1SYMHN534FmcP5wespQ4XUAEenmpm/P
kLiuTUNtTDapr8q/Uj7CppKnZU3YiO0GXdIvzzxXfwdCyGU6n+8N7xRurxQ8GJIrISEcyQjpzS/T
9FC0adLCA4bxgI5iTf+2nuRC6fpsJJ/zSG3fusC5/ggyD5GhCJqzYjWZmCl+lJ41ylWUP6iT0DBL
YM8cWvha7sDf+n0ojLFX7kuy1ypaMZ1HR0f59wbAhn3yNgrHjJtFm8LMdqs1H8zWlkIl/dQHabtX
2gRl7u2Mqjskv4vjWW5U8pMJ4/huwJ+xQWY3EvdwGMQHd2VNzgoVGqCX2oat0K+CPSZ4IYaTfgW3
x2r1iBMZgGBlWOk0hBd8FzXdM6tP69Nj5j4y67BbVj5ngeviZy1hFhWThrS19dG+Wu8XqtP2jwWZ
VcsEC4Z2BIsVD9+ZNZTgcjC+Q9vjDFCdBbO1Klfoqj3gr1TEkOrOGiIXDpf4n6BZ4ykFMcslHZGV
lw3LJP/MhBOpD88MFE3LrMaRkdwQgqwOAX8/pCmxKl1ZWidb/EJrjYF5rNfFZyP0EP5L/W9o9gIN
H/VnRbZQWKewSqlwcWnT89YfJC8mWCRK0D0XDOytwm1Srq4gsCGTbsW/SecpsV06xP97Lh9dLrOI
OIwLc3wznX22dL/0ckiyJF4PjdwP6FQLQp3a7UrHXbAYbAd6eh5dYasutLOUG8FtKYkJP7bD6Gf9
yqz/V7q20g2tLxAutQnX1TkVsTDx6xNXpCqxQKPmIpqTf7ukGgHgsjPbAHDW0XXRU6auE/OyspYZ
G55aWOqxKwvqqzYFHXjmQ2skzXyLPAzEd5ne2Kp0fEj3rw9nlC31kubD88FhyrSuAfRL0EEIQU+5
6eM214ibhb5S4W9tIFeWjVZxDH6tC1/3ccNIHRhKluSnD8DBdbg5hkPDZSCD4PzkBFh3B6CIGjoF
euiOOYWDqniXl37g2iGano3ut7lRkX7gMAZWTeg2pofxC+ttVawI91QyC4qTGSBRLB6JEaeI0Kq2
mgS6U8uwfj8HdGwtHAHa3beWSiPXGoFFldNFohhu00MH0av6viHobpGA4EJR5y76+CyXgXNm5JSd
FwiOB5nrH4VUXg+GqrPuFj/oJIp779CDKYSs189KWD1RM77/QYCOvoeedeBeWdgt4ulDjVQWZ/7J
DIhB3rOx5OOo8yN+WJu6pvdnNljQR8/pKM6ATjhTdrpVsEONvLg3+lNWRnYg7ORPK+xGv0TdPDSv
TayFZbVlcH/M5MbEixXahCLHINVdUpjzojvKEZ0MoKUz9UWhMzjvuA61GWO70saTnJGmaI98KOoj
KcJpEB7VlAw81GnAt02xWttA8bXyZ12IqxCcFNnUu0qX/sZgv2R2VEx4OxPNVUwdo7Pp5Ac3Vzut
etBRzrgkMaH0uLEMqon7aPSLemiqPukaM1Ed+6z4BfuWf27L44VhqeLcvHtlFctw3TtJBGIknkpM
aMDfHb/lzvXbBLkSvDd/iAwMxQ5LRXSBMvXxU6CyBY+CBeRsvAbYbrLFAPl1WHT1fflKI5vme5eR
+2PUCCQHG5v1JlcJmuBUsQXgMu/M7DYrUa09PwYLBgF9WzwypTgIMttrJPgeLYrtjQN/PMK822QO
58rKCA9jNgAvV0z23jxngvRuvMuo0SxWcp7cEhbACe1mJUBYke0tBwpLe2pu+pVUvf9oYuNvBd08
4v+IQJQQVahSLfVu2MRn3NT29rhEdZwrUXUNYYjqyVx/N7VJQxOOCDev3vSeBi98ttwAGUZqLetr
M4MjLSC+JTfZbXyrNfaw1852kGQ6mlygiGr2RCD5g1d2o3o2ZfClHJN/u9qDGVe636AzGqNMEfPF
68UEaTRSNRwwTNo7dH9j9NVR45+9icANLCShWCAsEm6cq+Gt9yspKR1wnvpIxWui+KMRg9jaNSCy
PwBTSCnjYtM5snphiaAz1+m4ZdE5M86QiSqHIlv9nHYjQLXCgqs9+LikV5mGvqCtF4+Xyh0lGzkO
7CyyWXtFm/9gVVpFuBlAi1XlZw+Yz5Uqn26lvqbjg2kIrNUgUN1Rt1cHoggfVDJvHyLdCy8pxEL3
ffGe8uOXLhukG+FjYSk3JK3LW/1qNXoU4M2gDRH/FLOgGB/WdL2sEuBXhk+0drDyujEzeuVKb0Ri
nV/UqzgdZF9WS7orZvpn7BZzZuS34qoTYL50pJmoNMpG1I51MA74TUt6Xoefhft3nVB3Ll5u/usD
kBPkTDX8wxtLvbK2rhvQijxfmKRPFJtte6OprqNnLbg7P58WHu26j6vzJoBEqO3JboGYME3IYuOn
sOLH1uZJkmNRVi21C6Nd+r+28YzqKiWbIQ0RMaG1/+a79clSZmaJZ6n3D5ihF2xQWVS/TGg5P1Mx
JLsmAO0yLGdyOpEgCMkcb6ZE+tagwJpLDRJBVUx3N3eqd/D3B29L4zzeQLqGpHXN3jpe92RulMDy
1Vy9p8naMkRnuPxlLyLcJutqCshwvPPoRndrxd9AEiNbzGgnRlPNiyrXubo22lT7JhUK3UN4HQNY
FGgus5i6fP2AwwJTDn4jrYiXS4FeiLqZOFACfwx2XErwgTu0o2c7rDc6amPK2rkx62sqcc3CzuKH
kh1cZg4UmbSvz0SNkgZwq++2inYZtq2dT30/Vdt68BPgqaUZVtsrVyUMv5Vu+XCKr1Zz6bC8ydY/
KxXYlSnzm2+zkEMUFI8hPccft2kLbMAHQzvBjj9giwcEfDl+/ugapap9y/uncEmRMvK6NV+zh/vR
NYygBFn/qJaw7PNcIUwAKRaGWVgGfJ3z+fZ8IE77//21u+n6vbwJwPcAAkPTNBoeN0PCUL3fSbW9
8qQUL2pIHdf4fN/2K9q5GcnjGVQqdf+qR/lBRx+eYXBU4RxALLzLoXZxb1NPMXKZIsX6vP5sQg8s
LVirKUzh3U+nSQQs201xei4/whkxJv1Z33i0YSdZbKkpesJ338XbNEQ+7IgLDdlYQ6ka3hQL/RWW
MDzNMqnC270I2yI9bWHaH/B1235/psAlmuCC5hVrK6bzDF8r1c17eHkF337LjkNLyaglvgWn9KK/
oL0V3A412XTEhtrLqtenhYkErypph12gigPz9qEqwJiBt4JBXzkWtqPw+tsIMOCDlAXdREIwH1Xl
BzMU9zNLjtTwbt2z8pOl8b5yLV0H6NE7pVtLRhluKpPwxcGE3CdKTgYKVYfu5QdBhA1kTZe/7JtI
UtQoJ1BorDfkLxsHCA2aC4rIqIjpiiqhg5Evb8fJDlc2NSjaD3eNoonobd3YXk+QwFDCd3VI/G19
TZK3oL5NqOJik6fILe7sENNg4i2JN4HurihG65Znkq38gMCyUVTiihZYBe91SiyDeLf5/IZ6bfv3
hxTidix7YMiN8j4JkiroA4L4tmTikLcIu/LjTbazr0FNx0AYRuRa9oZ/vogJp2OMgu9BU6E16Qed
BaE+50fM5iItoZgGaQhjRRV90rVi3wQWO5ZW6grK4S5L7D7h/bC8mnGmXZCKal9N+kFTuUqyF8lh
28Zf3R1r0CSuDZh2ryvBQxP8PiQ3guKwpwosjK0pGa90DKCG+XlgolMTYg4rn+EMXLcd0qZzRuZw
SLYkllrWlI8IQV3CpdwC6K3e0uDdatqOTBOEwD7l1j0XBtu9b1UYMNInE90yNXnFQU8CohL+sNGW
R/OzX3PGX4MsOfpuwSG1K7anbf/O1y5H0Gh5yzlBJqmNMNtzqD4B1FHgOY8K2Y/1MLnQXSrsNXLh
dGxtgpQBL+OinYDt/Pel2n4vanJlaUDGCl1+liV2eAFa/tV321JoZznEbxxsFfrCtERacHRUn54M
dXwsDxfbknnv11ESIAxL78/knAx8bhsZ97bE6/XoKBqGPbguzHjTHfSPMO/FZIDvVhyDVs9335vo
tg1tu488KfeXbVchuyfBsxLhL856gPhRh5JeVehusltk6JeWbXSKqTWYFs3iTknv5WZSvKxCVJF6
Tc7nTiYDpr+XMTM2J7HlDIXKDLAxNA7xaaJPzxL4uSo2pvZRpT2iXvQMtgrP1KpWUO0Yo7WlvBU0
C6IF+gsf2xWwEl5vvZAdgwRhlLXGh2xgjouId6lAydI1KsosB6akpcpgCubrA/SP3XO55e7lOcO5
9A6shdwPv8I+T9SdiVU6q8d2CUm8Hz8V5vI8QULiVlNcKqmY7bL7GsQ8+bQ7U9QvQtX/WE6LgRbS
6yIbRhZKa21tic0yONbEQ6V9vToiWIE0PsWHFTlHPP9WHJ3AuvIy8g5st4CvPlJWcwtub2lEJRfI
bcCcikZNW7t1Fli4MmSqUHQg8Ma6fby5UkS0waeLoKbzFhri1CvAoJOF8H4cAS4vz27iEWOMdouR
NxWsau+Wsxj8A4BwvlrKcpZlJ+Tu0RJ62twqSrmorg3aukq9C5LUt5volbgPY4EAzFyPWXnJxTpi
puW7/DP33UtUa5mmqYoUDIoepM+AJmRDg7YKAL0P5tYpegyKuR9KcsFP7732R8Aso4r783bLoA0A
QW8Tejvi4gVNvBcr17iHeE6fH1sPluvgYqNQsenlWDHnXf09piCc7T3CpvUkSr7/nWVlSHpm+631
wOtJMEEUfFpuLpJN6130VsxnJeIyZ0FV3BpKdUIphfzMdwPAh3bcyLrq9l8Z7KoCzsXIkoE+HUmP
yRvgpKfxru5NCuo6F5k0tc97xS06W8zH9Ey8YmREevBqZoors0WLhV/TahMAGfod6O3EylTvkNyD
OqgyobzCRbRR6Pl/Ml0hTNgU+kgyNNAQVfX1k2bA69IOWPDbNveetOjXlrrrLhZF5Y66BI4lYqWE
/nBsQ0wG7E5a6SA4WeL8uuYUIlmu65iTx+HJU1L9seiKWEAFVXzT5iVuo4SPN2g6Y+eduSfTU0K0
7ll/qBEch/Vxylr5g4jOKn+ypawhFOMX9B11r/m9BPJIBHdcZwszKbHtFlMKJBWk+gaosdLcahgl
X1NmrKSZFH1lT0cZm05eNHo/sJGXr/Xu91UunXEMKBKzia7iH824kyFXJMhr7UgrqtV3Gj9TOXcj
0XquuukmKdkpCXZG4q4JpE5a/9oaThYOm6t/hDi/YjgqnCrkYe4A6GiPuwXGPMEXKyOjpScLMqTG
vSsTm4h0CFU4EM/4B24PtutIVyNtgm5/3v3fQL7nKFIP44YP95r+5y9QAoD5E468BVOtcWSficCe
1Q7DENxcQLRXdCmnyjZvxCxzlI+RKWl3fMELfhkka98d/XR+kftD4FOGwybvOHafkuXGK3PCdmC8
mCXnbfq1KEfqGIdoni5/eGm6hrO7p4umJ698GbiiYbrIgn7fS1gV00GgMbJ2vizZeI+KO4N5ltK7
oo33wHQqtdI4sZPv/yDoPhGtEXPIyT06+w3pYoLHAs39nEfUR+hncn9rfXsOXOZV6npx1cF9FfwK
5zj6WuXZZ7Gm5F8eu0/g4JKdpD5mOIK/clZpcTr3AIe0fyFVTOVNlOufotEwzZZImDQ4PucXEqxh
MF54LJ9wby7WAdqUBOrxP82iancxYZ2QQrd8Yr6+97F5sYAps9imomwBla3a5azlwmCaNtXNxGI4
MUXvImiS4IYNk36kPBmLENpWUV3Znlxoncg136lKBydq5YKxYqD03iazJBy1rprkk8y8z4BJbRng
tGVLkzL+iPuXz45xcZgEGkqWSbzU8PntDqkSN6UXpJs5W3H5cPqBspoiPnTa74MKdGM70OtGNMCf
REut6VP4TOlk67ceauEgKPiTiCy3RhqPQKTdmg6n67dYu1diLjxMpXFYfGhKzd0BNDBECAwowgK4
YSRkp822WQ1K6hRJQpzCYpgOsrGsZaV4i6wV90udD428E2tadaqS6MJgidgh4JPiw09DaalSN551
mXBDYHvD+nUQ6Q7GQ3D1NnkdbFZjoTfF6+4UgyagULJEMuPc0eiCIOoGBZniRPLeO/ADvdssIFDx
zmwBGdN2eT8N02CrqjB7C13D0XPyTKZJGIeTloQd/aIg2RMwTTJX0XrLaKjvnKpQRTIuI3yxcnUc
4wI6k52DpSCTEh6nlK+N/skgQVzZjsvgR5u5cpSfW+BRTqc+q76aK3tguF8Cq4ckyWJfWhuKiXMx
ohQl/1gifJxUvkjdZApcQ2JTau03VypdTwhU8smDCBW6sycyHCU31N64TBzmE+7IDEKVTmhs5cVs
spBVk8rW3L9Dm6paK2MVxJwW3h7in5DbPXHTO+MQPCryj8dRxFx34hTcUdDzvaKEyzxiDZnwaEoF
Iww9h9KMueSf30E5c3lUtJ5dE54Ro6U4of0MZocsMlXNncJ3BS5rjobljr8paX0mns3Gb6pwk7ZA
VrHwUWJR4COkS2O6iEYV8LGkrYgdkI50o7b446NAHmN8eRhKbp8vKOlleWg7VJ2r3WHH1yi50wN6
ztaTHrvTm+u+AH03dTWGg0eQ7WSl53WVMCIdPDKxPM8IUfIoN8dAwmwpxBKgLS0k/ZITjyrUEJBi
ViAMFVf2un8PTAWl3jI1THCZQJs1gVm7zEh0Vpy5pgeKSXWMyeRkgu9pE4kvUbgPPvdHojL5EnOT
JBxdZ4/qj2oX15uMgehvirbJKz2WQk4rFYYCKzuWsZ2nj/D8QGXfvSy6d/Ba8Q5kAGpS4p7N54x0
tRCe3qreEvc/ADA7UJcv3kfw6OQWIyE6Oxro3g1YT29DvZw6Rh+YCgc4+567HoAYp2353B0j+36S
cY/fjGrC7xxELnUMO3KwP1kKx3DqJXSkBz1wBWFZPO/sT22S6UbD/QDSxu5vYl1s2GeYvsW5B07K
k2UkIvGumrVK7LQgsQ3fU9Gk7Mk/ag3/5B5rjkFBmf+3qX2w+4wmI9NYFb3dP09kDrS1tftIuMiC
nmDuyRl+9qz7pccWWato6wyaPwqxyNjn8IKdrUCJyHNQAesxUY8tHl/qOSgr624duhIi3XtE6AaG
2bsQZGzyFFhWu0k8V0gvGPTFdxBzgwbB0H2gBqNNKLKVuO7IB6qrWA1NH27iegLpTNiACeeOsgVK
bR5LN61NCMESPPg4R89BaEeaBjKvu9WNsH3KJqnoxZsc08sjqZXUZDTBByNWZZLmf8AOHAka3Xd+
C6ZFj0vpN+Vq+NTDwbjqAGtMLodM1wQN8Qax6flSkQEJ1HQcojs/erv83Ce36R7XukkVgZo3M4Dm
2OFd8hR15VWwYpMka5fOsl2MEBXqjrRE3rQS5a8BOgTXeDD6pv6LDEIacUVDBO/mBFZZBj0UE8WA
+qQcVu8duvJ71jBhgppsFyfcu9x8MRVXNllsFGTF32GFoS3S+jAMKB1Pk5tEB0cNtINVnw81N8lO
Yc37H26WIg1eA7MwbstU+fTIpXcBVeHXV3guGwibyYbEcIh0A4iZtPlPrHLrNef3icX2qORp/WAJ
3/XnmWO1+pywnKcgVWN0328SVscFnuodPd2HQA/wev326PNbtC6MpOVVlDAjJ2FrmDnFoW7PGyCb
XUC40s4Yf0o6YsDjK5M8+sxcEtOULuqR0/YRfk6G/4ux4gS3zMy7utniz/2lCSqXXQJLrwBF8Em6
4MY33Znu/5CX7FuoHQgapjx3wkY+Yhs86sRGxnkPVGssHQGKE3B5IV0ACKexRizW/vdQ+M4FTjZv
PB6XZiOJnVMjG7ngcYUfXe8Lxb4fXYti+K7WAC4HBD3xNhfh7q0P1KfKkF3tZqi/w8+afgJkkwmA
/5UhIx4YIfBJO1NFOcck759BYgvtOPyvhmHnAt/VXXzucUcr0Ls/MmP+S7n1SPflZnZLiltt4JI5
6zZ0j3B2Cv3KNBBK0vCdly+yqPRgxeGyFU+dqyu1I6sI/ymqC1VkoWU0sI8E5NWIHYYgV+iWYcSh
CQgmjNQObz9Yhi1TK2oTiXaxMjse0+5XxtGxh7CKVzA6e/H2GQHfvYdtSuUH/louUBbHJrWGENbe
Jkt7TIq7J15tCvZjgxoVBTEz6jPUdcba63KO3CFtJmk9vGNUjmjf9xvai6wWXzsya67lnQWoGHdT
fJVGy7vFI7ttvwpv3FMaEDcpOvDfJnNVYUBAi839IscNHJSqJF08tu74q3OAtM8sIaT6Ua5T7/Bk
9MvO9xNuEqVn/dBfQ4kRJcHNA4TkQUWPWUvG5m+shIsZqr8GWVEjIyLyUtpiX64WBliliZx81TaJ
avImSeEwJSRyfQI7jzai3w/77fJB9WdlamJ3zeFyXLJ0FdTFOSELwahY31/6Xt42DSjFb4S2fAH5
4uNIEuzU7I2Eyo3sU0PRCtz3F7BnlIheiM7ngOvXuXnFb8c8+jCp+TBnyUix4Nh1MMTubSQAoLKp
/URRVx3Ly/AFeoT4Qq8++0C4ngNnGZhzztZ1XdGLgEHa6xh/9WXCYnzCkGSAl6psx+/755mzeDj3
DwMvMpiMNhMhk/z2r6Bk4MVpvW6tatVQ/lTqAWQ1XMf8HESuziL9nHq4ejtr53l4ldmh6egsD0xS
rpl5Yc4s8GBH1T6Rw8i2kxlBjhqv3XfTQlhCB/nRPsH1v5ISVmQn/EZPFvHjLObWM71L9pezC7jF
piA4E6SGdGH/Lo3XIHQF0m3fT8vKPoAVlKRwX3/TZdIqBdZov8ILAssa/WPp0xxcK2K1oDjdne4w
byCBVcLGrxQMeHjqV4n1FlYEiGzzX5jteWzKox0A6zb5Si6q+RV3SSqx3dJS/B6OmHvsnnto7g80
Rcde1tBvKDtcTYsUO+99YtV7vbZanC2o4TurgUPY5XRePHSFWZtzkpIBjv1hY/WwdP/6isznLbjT
7aOZksrIzUeINPsNwqi6By0DFgmdGdOyNGbvxc4qtULZhS6blGXexyUBFDnoZeAbYcII9EdGQA/6
UIecDwSSKC0SHU/lmkF3f1qrHf7Xtj/APjZkrOTn+ojOln/l4UGsW5vVQ/1LTl7ayAYbo+cnU7i7
OJFSmCrZvTTfmGTcsDwGBAHHrYxl56Ko47EVU7sr3GSHYli3BUGlbVcxjNxWw6rPBTcASVCWztPQ
9MHvJd2b3y2oAQPemWHkpvcYdZkf/RE6pqsBMSq5wWJ4YC6WeU8OdxmoxNETGXBOYwmZPXZFgC2f
gQOUnOCIzo2gGbMFpq7wF9//7+HZs/mwA++yYZSjqYAMZbssPRfD+itMu3c6yVr/W7vwe2dOAEiQ
JJkASxOidaPASOYHzW8AIyR1x0C6EZmqcdsPF7GLuDUyjCgvaN6SXPEKZbYIHsYV9TWZ9UhN040M
VUP0kIq4xxME9i14ENuECONDu50RXZ85CitExVyxVUObau/UZ5QrWsJroF8Q+ZQjHSvxw4z2kUg3
vys1dK9CD9MS7+ESo8oKkItWFm4VpK6ta/AbnAAoNxs84rc7/nGWmrsz95iYFrUX6CzdoZxlhgKh
Ml4QPAL0g1R1+my055muscfjHGibOKztiJCWlIQejJyDyJzqLyicXNAMwvrCFhBAK3gKfVuGukm8
LGs2prNaJzQbQtm3srmMDPkyC0sY8OHj30vbS2xO8y5ihwyjPCaOA2aZzwTqlsEbU4nzxZhOTjC0
pauSYr1reXR7LaJ8/vDL7NsrXrJY/XC67O6f+oG3Sfhe3uGd0yaQM7cYCD15nnHDGUPh02X3AGvW
HYudK0175H+YlD7gSNur92TITuWP0CvBnAm6iazt6xa1HFo3wEVXybCTDmRclbBiWPvv6miKBvsS
7Csfejrinn4LY3YV0nFcBAtMsr3zEdgNikbGMTXcJVYWKHJ60fJazWWfthAfHQyc9Prf9T4sYSJu
lvJzjIR/IlpL1TXZgepBe1UVYIDPYsaoAHEFFw17m7r72DkyzLxepBfdciFRD2SzSCiUAUgRp/ey
3CyugJ2/bF4JP3y6Bl/mbbrtgeroVx+ZHgecMNDT56Q7aQSvnsmcOMxCWftJaUz25Wy7Cv4BqIX4
Bd63wKugtUTo5v4XHxVTQtjkLvM/l2l6Zv6AodkB1FgnwXsjrg9AaNbv1RwpXCw73rZ5SRok5UFt
sbCnNPEsQdBH/eGAHYR3HQqcUp4zj6cgBIuD9FOSaT8ZefhERY8tMgMhgBJbcd/tOXg5d/38CNzH
sDofLGItyeYWIef3vhjGx00X5abxc7Idoiw+juTckhPA5wmnUh4jDSbD4YfFMfOhXgKV8tCwDw60
vpOJ4UlkuzIPd5nadzZcI/VJ27RxX777p/FK/sVPNkc3l15ydsaDaSQsr4gaQ+36jlP+knqfv/de
EqhKMaUkGDYpFfbsQF9gcxeanV7FP9mDwhA4OY7bOSDwL7Wc5oZ3C9wK7ud12qv3oFFrBU0VeAbL
olUErxsjwZjt2o/jpMS+cJoovN/UWFaWEhm7BJNkHGEM+Z5W2fl/iq3iz7Ooz81K17CQOjS1pv+Q
JZ5srMxYk2zXdOwZRqYHZZP0SwfpV0IKitedhnoBkzGYOSnumhHCQp/LTSgBEULgwovEyeFSRUzI
kytxm3hrPgeOWqjs61AXQF6WuI+WhvCLeerQ+E72QNboZyFhQ0b7NjmfL+jhhGEktnLaFbcUt9mX
Jc6aomeTi45x4u1e7dAE0jSNKTnafMRpF7m9bcBf6fH2NIg8FSrbrElRz8fp99GABGM8e2YJQV/C
Dni9gPHnQS/Ax45dKzB3B0JL0KYOp2RBVkjEWEwMaizNKTRRqIaS30uzqyNYhUE4tGeAIbHQdKev
+8TPTyvUSPEa869J2Ehi0CrUaeyw0RWX3pKCBTkqtRWn/57zUxFRVOCqpxRTdCCu2T0nfSwe1Cf/
69Zrq72zUN6ccpLMd605l5WvjmG3czUMGuDl6lzJnSa6+wNPTpPDgWqmGIvlG5rZmqGL+gkyoXzd
zDkd3T6wOdPu1p8uTlB2nTv6CjQbQHAl3pYeoziB9qe9txPxKMp7cU1ka9fv03COlmGobGkqWhow
jPB4eQy1Mjwk/tJGY2JGq89qwkni4Ty7b5L6QxPwsEfcDvsz9yxD9AkXrCU/u/QgZSi95EBSVk9E
7CWPX499xApLKtRVqhynGcMxYxJt04pp7Zet/yQ0x+nhTFxBIhi8c0Vbqr62i913VFfLvtgNWDtp
hW+Ai5ZcpgL61XMrMN9EQKDhrCLCfWSBNuGockOnPJZmBJHdVwot0ty/O7ESZLHqOLcSXVchlUF6
iAF0IKLL3CHf3CaglGtgiZUrWnnISjGPHdgBBaCHtPRVA0w9sLWcbzjMIRIiS40nNG9mrPbrX4Ci
Vb+3XkEcl7OpXsQ7E98jdHQCtkhUSjdrAZxA2WmkasI2G4Aoyu2K32lLn8Zka0naue1pJRRIZOBt
jxcpzOSSpPak/tpge4j39VqX+NcmYwTJybfd3JJ3rG2jHf7Ll1MsL8HpUlhs2Wwyaarp2DZXLFTc
9Y68mWVDf1N6AkWFFYIFic2Wg1nCfTtvf3J4yGJnq1uizYgLoC3V9TokJMGJi1vRs/bAxnm9ijo+
EHyKMm52GIQMX9Q+rIhecIkUr20qNp+sjj2wjMHStVCWYCY/O99kYbH4/ETmS5xox9/BJu0yFP9A
49XWo0Ja0yKUTws8aNtvdgD471nupDLgHtb0IHe5BeX0qWHs9fdBBTXP+aYPcYTqC9ZAKSwQ2nWa
CCWOUZZ6QhBKxg0aX7t1CeqABmCVfIiMv9oSBj3mWi7sK8oW78seyU2zWKfodgKVunYo3EmGNWhL
x11l2iMvk84sfXcysHoduqs6s+NBEYZdkC7joBToRIBFeIH4bRq5+Dh5lsgPQakPj/waPHbRBbCC
tRTWxpObWrr6IxqVSmn7zb9Qmo0COxfo17zgb0e6C+dYiHmPflhHNPOZdSOjekaptjPkE8DQCW68
P5Z8+ToTLIP8WwxRmdom2jKXU3DoAHXVPOJdKJz2/SpKWtmWioirTSyhUJ5R0HXh6b4gd06vDnP7
XYzE0/d9y3NUWXsfbYzQgv6uwEaZXPGB3fp4i5TQ/yQl1ldohP3XXnhU9zPQpJB35UsflVmZkuHt
XnkOtX//rm7SWK4tgxiKJGri5F711l3zaU0rTgGgf2L586bdSsQ2adyUkqfm/H9HYqo4GAcCU6Ol
TY4CReP5wQWRYPxFRDsymkyLYeOCgfI+5m+XjAOaB60+vCE1y2P7Hgzhm9/dL+RfqiaBQJiy9Qcz
aEl2PjaQACkb8YLqN651DxDM4JA3mBkx7X7C4NSw8UE8TfRO5p7TXDXtXpA0do4iTUhcLkbaKpYa
0z/A/RwDKPSn3FT08OT1rMagI8DrSUPQDqzxL4LuiAKqY9uj7sUSYi7OnVTdPFBOkhl52zWuQjDZ
rhiUZ5Zz7BQXIYb8+TWcr98c8btl6E64NfeHwHOiqVlQZCbFD47dGhoCQK74Exd8TtouAsHAUEPg
p13c5t/fH+zrc0QV6jZPrIPm5lM9Ko1f1O/I4s3pyxOZFR6ulOM3AFWGYyselN+kCuwM4oiAp4qp
WUNntQtcLYchUpDjCvG3Bs0Wv4Ju0IASaQNkxZAVQloBHOjhf1DeJMNqAEV4dg5Y3ibzyaZryOX8
Wt+9VE9c2MfpQl81DsjPYiMQO/csZuecMxUNg65Lmvnisc4dKBY8Hr3l5VtczyqCpCsfLsB5RzfV
KCRzkt/le0yVWaTfQVbWIgE4+tCqGUDS1hsc94LX0RD/nDAZOYy5kOntxwm/GKVNOK1bW4Kcrvpf
PhZ/p+kWJcKSbgexATtiNkpWupTJj1sXzkS53R4Ct8IIEA6hXtnEWfhkU4sFAeGN0GKEXTeIdRDR
ay9XcTW0cFtgNxsRiMfMMr6Lrh3R3COL194FF4ohJ/3hw8xAl1DGVsNbn7W1By4PocFlrKKJso6/
ql24mDsZqiqhzxJvvS0DUET8JH/19FYs4x6wf8Vcpz2ImAwvGxGSCrzY/03JW1uE1T955CqCnb9q
9r+euDhDiQL5MYYjAEI0yvz9068bg9vyyCI+podkmbCVaL8pQaIXmXZv7enIkJVvIYb7QvsUwrZF
QXBFG6ZI4gWwtaPOxgHfb6ycVDw4OsqVnWGYPuxAFo8eywblLPcS8JGOTr/c4rXDGeZRkwx4Hmqn
T9Zy/fXvI9Is+NXEqoXR2gW5VvZ5Z2dWvPAO6B1S+jt/CoaOyUO+/rGxcD+mNxSO5DAjwc6VIZON
ZGXZxK0oCwhcJaxy8tlQvZzZDG/p96VjCT844X20seq3etnDhh6990znUt5tzm/xFFMZVLqCWkoH
tTcjF5Spwq/XSNuOwVJTusMA2bHqAGX3B9Ez616/BOojvEJSVbwBaKT8I3gaCnGRux5KF/DKkYZH
8K9C+K/FlCZDoJcLh2gKr/8sxLbJqF787AnsPV2bRAkWikQbC+mZZS3Su51tZA5SGQs683K0YWHn
h89HuTf/PvKvLKE7y4Jg+zW59l69/hcLhdNQIQGYaHfpu+uyl9b4389anxhnGOhTalWB+/mCymYC
TmuGy6SvgQA12sSJMlJUOhqTq+LIIkIuZpoCZNGM5YD+n4uZeWtsPltzZfdAvUww/r20G78vnV04
JIXS+rAUKT+7KTYmopkJojaO1zPaBHS9tS6adGQovEx/75qbfXZTfXD2fUqMFL411Oov67ftzY6V
wgsXd2eBR06ccBOFnfIJHMaenOS/guBUEmz5YXuNtkFe2afi0kaNSwzdXoaZOjfkxNMEMwxeyVpf
yGQFIMF+/1fl40ipYbcaIFDhD2Mo5Y6izzKp9PNwvmZ66E/7pJYsupvEX3OA+0EVTlLGp1v9Euxx
MoicQZLJjwWzSagr9IpFYjSuZPqIWh+z9Gw0y3nmli7LJ9jdx2evHA1pGzqzcjCjBZQqao9PMTY6
rB6Yac/YweCDHzLGTWn/2+uLlso8DYObshh7r9rdAfw6l4ZyZqmwFPyQYWiaz1kZQLlyfsa3iT9t
aWKXShS5cINGoDXgYwJLAaQcLJRXXSyrv3/o8MnzMn/LlFA6rZSKjSoz76RI0gb1aSTwxfGiD1SW
Go+sVObSn5wXA7DD3LGdWnre6910w12KM/j78rxI+vpYcpk+9gGJajku8/m4zcefYW3zmip3A/ZC
i85PfJTeoAcrw/nwDm6Uq//o6MDLgqR+BqdFYA3vgUBBsFSISGU/DRcH3xTIGesMxYzJzrYs9t+W
5EjCJ35fxXS4JnFBlaTMEwJlQkFPLcNbeVmfsLBJ4nhlpbNG+i0YYUw4sEa08X23PoeUmYUIZH2A
vV8p1EsTs+DF6K2aGvINpKhjSLmeMe4aS4cPDDtXd01oQS3DfBuNHH1X9gnUFbUn8oJjWFV5h+mS
QgXBwUF6S5Sdaozd/SYXiZ9n1FnO/KOlgReZbSLt6IOiOujoKlwpEuN9z4IuHlj83oEqFz07Ists
WUkozm7ZZnUY/s5quGuBhW/JM99XEsC8s4eBLGJF3pyBlBle9GtBYEKhUUSTUp85HBzRaJCVPc6c
056HYisIOiTPK4+b2onHHP5KGkJqkPNwQ5SyEnw4SQsf1OIBvq45h3ME1b3IS419haFzSIuRZd7h
4fiVAc8qOT7QzBMk1SZllIVrtsNa0h1I3j7FQ5nVpzZadpol/sQQjN7z6RV6+nRl7eOl5lAoNuol
0cInR24RwVtNbdSuMsWWPA/tLnJNBImy2iXoWxZRQqhQtgEKqZwAVrGb94gpJPES+76FAXDQo4NS
Sr9GpdntcAc80bhVCszQbYs3ifMvAIgYGwOeSwO5Wky+V10ZTcfLCotrsh4N93WHoVj0iB540lFc
waVZBwpS1gGirv0ng1twKvHgf4RwvBjKB4jhw746mu6Ka6ITY8U5JDs+USqm/mussBltCYYGjD80
wZcfjRaPbTK1cl/X5n+2pU9u7ou2Rhi/cvU5myd1DDLy9NwaytFVxNjS9xh4Fgr/Zw8c6PqUYN+8
haHPAKFQ+BQWHBD3UfjJvu2Wz38FFpk3wGgqu1lw2Ln5whzo42nRFD3BaQ33Mkc8Vt7y9ASpxZK2
pDzgl2WtqMaplNqGMSWU3G2T6ul2bOXLFl0m/pTRMHVKJG/9VwuEUaKm1x1BwNMut1o/PECVZZV3
Ei/+0oHLmLg9t/AmxLqgWFDrhz1M3zkIr/k2JFM7WICe3txAOuAszhKrEoWxrC5ARBathAKLBqWu
R3jBTPsaXWvRgibhZsfyinzqjU0NRqdktStmjduVdbt4SRng/nKEA7Zs6q92a4i1ZReivlwhlUnz
ldLn+xbYN2cGCF4I40GiSrmJ3RZ6kpfVt8CfaiNs8H4vItdFfjgVXrut0c6iAAalfae3vHTx6xT/
APhqb3+a4NitSQFhwahulsJsx8apX1YYOjDArIgJjSOW8/C9Fbfi+d834AaypIzG+V3Nen4NmJpG
zdQtxjKfJTXyK5fXOgXENJjljB6mN2Mhg0lLTD6YGU92LltKKqL/tP7lE//e4WOTEF6SR2iN9tUm
0pPIBx2UZyV/Hmbp1Gs9EBclHdfRLdbiEIHuL89FZEjRw1Np5lokGRJRi0FpiOMRHByHxneRJFpI
Nwhcj5Toopc4AYh3qgt50eERegaNh0Dc+k2DRP2OXUnBaQBaLjA4TW1TehVnwWcZY44bYLF13pny
7xX71m7nU801lUR04mkzxIIzp4apdPehtUFAP7dezIW75Dp65En3hIdIVL1IqXAZgwrl7zRn/D16
jHmsolos2bk7QJmkEQvGdbY+9voo3gpTBSp+SwYPahTKq70/rY0zApzIydSOQbSMzwT0S0HmTdQW
7ISVyJdf6e/JvObMd7Eb/JmzuONQv0g/G6ypHsCJxqGsAG2zrgl8to96Zpv+yiOQT3CipGGlkw28
k8fCLKXdBMjGAvIvGt8eU6es0W0u5/5fi9WFbEf9pwk+jEuIjhBHfhdak5AEiZmePlk+s8LQM+t8
iWB67TD9djRKVtgpUQHEgl1W7+AL2WCD3IlqieCaG3EfxCae3FqSTmmFmAINMoNGcMXBjKZrP5Gf
u1UHydZVBIvnkk7m7g1bFSr68vyP+HPp0SDYVzn/ziCtWoi97BPQjRNo/mHjIaM1q7qNjR+MKU1m
P+7W/0G0qNtGJo+HnTXhR6k7R6Lszrw2yR4rAkHuREj/PQ09CGtyYP9Ox2ldaVZWaxfvJbt8wxsP
woYaEbTYh1wPlXsOWwGUnz5vOffnZ2gFP9pxxh9EwcSnjtnjK8KJbsmM1WSC5/6ae2/rGF7GM2in
T6ZuJyjm+Vj8I17/8+Yim6/XCuj5w73G2ppOEU/RJIXJool19JkTOcEWYhazOg9brjaxzadXvPqm
NRxjRHvmrKr9N5rOKWLV3ehBXeyp+89Wml9ra1JumhNUyAOm7zfPcjP99c9duLUscXXwzTsmzvHb
Mqrx1DRfKgoL51jIoyPke/AmnqaE2oKHrXM8yzlqwnZI1dsnzTE3S7mVYlyjJwlbwz2RvdTQklKu
WYoEpFLcH/NiYDq9gyIG76479rDQExyNCvsdBcRLSWG0/UopK2rpazO/EkCjbNQNs8pxVQ0rknIV
0B2+PBLLqz6eEAHTV0Sf9gNL+rdmFIF5MTHW0PSVVNXK6Gkyx6gwdTArr85mBAp9pfTWFHolrPuH
1BuSWum5UrvG5uAFqhih3xmgqSrc/gK1x01Nlj9qJjuIIoPiy3dzKw1kAOqlPLh7h1VDmzXI3q9V
nJUmtZUPnVo7ijb5HOmiN7go8Zrjnq8KniLQ2XAapftI/96cT1U7l2I8JPDehps1L0Bj38nOIHAj
IwvpAYZbTSkFOhuLeS9Z+PUONky+7Ei4AK8brUCIEOCN5OXzlRlDFM5d/FyOEewefovGZBGMNcON
0Gc4MrTArFAKNvKkKwE4YySlUJnTUcfFQPqOws/az32cHRHCAEzAmMaUS4h4gsXIGrWCmzW2RhCL
4LlHWRgYkttHLjzuPj0gHsvg+5NJvu6Upl6RoeEVeUWsFErSeiNQbbVKhhz4KKUCKDWNMBqLWIDc
Ownc7HCt/CnEiILWEM+J9UzHUzZwV6UeakYBTVePlFAefcHC09/aCvmvUggimHFS2o7I8Y2P3Qx/
h4AQYZUtZxPLS5bKJjNAhV7tUM75uMKf2tbzUo7iHkJnbUX56YIFWKLdz8aIkRzW3YOQhiOTiEDn
2Fxg33H94G2Jhe8kJXoDN/eRkr53tNfGnu10fs4H0zodoKrsWsA/jx9O8aK560Gkp3pk6vX0TbAG
sbcWF3ednfzARaAJ1EG6b1iE/0yyQ4/KbrX6gt/Wc9lHAgE7fTGTAokgeMSzgNUp1Vpt3GSgBOE3
E+KJJPEeUD80xRxYDfzj/Lrp/0B7HsILu26s5X2p/vNuJIwjXBXFXkCvMhRZuQZDzfnY5bq7EPWA
uDXAV+qZ6iVG16l2CpGC2NLBw79GO31h/s8iX8TKhp+E09KegxmdFwRz4xnzcJ0Ab9BHY7VOX806
h0Jc4/dZ4W4rOyigF3Vl+T5K3/B4a1R+HmLYS9R9u+ADUb07B4LafL4sPE7n9kOKNJ0FoiZiNl63
VOBtNxKXhLsBuemlhN8iD+XY7l40kRuRnRIbDSHlFbszeoyW5hnNCeyXsThSBD6kG9qIK6g+IIxg
YSTNQK3hdsl1/UNDCn9E9t/XJmdnCAay5/IFIQpLD2uJwLrwggz4WZGju7n086RFfb2BtxW1XcBE
WstHzlKLspiioF70o3+L0MfZgOsqZPvqSCRx1NrCKzKbw6lyEKkVqBjJcYBqpKQNfjPE4PrqW9lJ
pi5OvGGRGhsjeOSid1IZy/GdzFExArbrSHMIV6ZdlAAZoBro+GJIoqc8H7mpJhd5ZyjneEbE4WTu
10zk3RQFSSNdq403Qncg1agFAXeCQPzdS90oJ/jpob0Op4Knpf3N5I+JQ2bOednSpX0MfwhU/ejE
n2koVCP25k4Cz5yxwQqEEC1GUnS1DE+ZZLrYmeWvGocGaoar13xUY7vWaX2rvCy65AnWmv3R0jVR
E2j0JYsO/U4N3zRJws+M6yyejPUfGTEgIFDq4bXaJL2LXoZLAEVo5iZZShiXLMh1pNSJhj+ccChz
DL9Hx8JuFWUGwa2iUS0QnQHx0jmhLlke79Ib4NuTpEesUdsdlcUSdADifSOyXl2j8Ov6wPQqHyxF
NyUkXEWEHZ7NNnT1hH2T/in872P1L34D6PZ4HUPLPVhx+UowhfF+mhtzZBuaJzaWLQ6OjE01/lDO
FADYkT0V7iML4Mnp3Sdxnk+n//kM8/5guEy/hYrrvlr4XclfpKR7WzgcvbEZMgPbXe88/xBFfqSq
/QF+xkXTkqC9uF5YIGj4+l1a9vZ9HdT4ZOp3Bz9dPAwhmOHfX5XqBXUvqK6XdQNkmnpDkaajotoY
HOPCruGq3Z8ygKtAfweILi2AKdQf8IY0nJzLKoz2hqUYdYNFNTR1fh4WouctsGnXqgOntThOsxJv
YPbfs1nurAKDLCuzwZ+dTv3+0vko07g3mWJV06XOW/AWodDkcWNgRfZKNwlheuFS5YWYdrEvZdWM
CLSFoE0dIZmDZc4zU+D6R7HHl7FWc39ZRwqJ5y1iSOUERzxh9RYO7+K457FEQrxoUv2N4PdoYla/
enaUFRdbbvn5z22veNRZ5Tqxe3KcA50iA4aFyrcgP5D4TaDWnxzrbdEjrJuQ/U3mPcOs0Hi7vHRa
2Gv8nKIB48yzzie5v92qn6i6Qh2xna1VEoxu4DR563vMMH2EvKzlnankLaCOL9LtrE5dKRHe7fWP
piMUc+PAROQqQ54I73DIJu+B1LUTjFp0lkF/Bwc7jImEWH/N0rUAFe36v0ZmBMyjORitzGCLB+dc
bIU2PHNJ++N4up2JyHrYJlBOIZ5FW2ALZbKecSF7lgj0YszniRPTdfs2KOjbi5kvddxp0r0yfskp
IMSpZtWjvcclZT4zy5BMNqMsqN9TGWhMmcR6NqGktmxOTSqlXCvFscSXJum07ZIMEXNzo6CBuXNo
V+wOvSz8bG2Zz25GkVWu70jw1Hj1fO9aBLAcm2IO6FTgGuDgnIVyx0ia6Eq8W4x08gWuHYCXWb4y
gWftwQyQgaoJbUUub/kB+mgxCM+svALDubvmlK+kaZ5Mhb6gTm6TshNvC7HVyBiIWwVoMstCMyWA
xlHpZm4T6QKzxZJ0BIqV985iJJQxU4l5OxmeTRat3hEpyas0xxPgK8jLo/F87LEriOVBc+NHmSWS
adwjrB8xkN9YiQofh2yjrHshtb7KoedfnMfB7VtfrtzShvFKUROF3j/++YrVtOBBQvdD8RQ98YPJ
07dnIasOr25iiXkbILbILpjWeXKIbUa2S6WHKt91z4U/zP15PLXjB+GB8HAFJAlnShNfayjn67lI
g5W0/dZ7qjQ2JUuvDOqhovp6QH7v8v/o8ETZtltKBJWgEr9aPHk/bk8At+svxqACA8/cS6C+rvSj
NoUcFVQuP3QWqsE6qBDMjOmnU5c71UkAqIx+P0nOKDl6wJQqx0cRgdxpCB39Y8/uwWfL/SEhYTrx
gHyPa+CB68hTkmQzgP79BhfB7C7XvqdCZHg9wiQOLLy3e95j5o93xPBv5xAIeqPye//tvda7ezeo
Ri1ZJr+PhuGvoYSLPb34gpdA4QZHUtnWt/RofhZfgOUF7vehYcPdv1v+I8kWdOi7Qw3feOS1CFh9
AmZV2xRkxcJ0VqjbLWsxmE84WvWZD4R1c2D1LjZbReJKnECiHRQetQHO5DdC5u20U+2cqKlJkSPj
8VQFxeOmXg2Z753fB8svcdH4Jm0FaFEihJSNlvrg8HyuKmmlXSd3c9rzHlVobACFGmOomvphCtbk
5hhgGwGsHCFbj67jreAhSMrSCBV0a3dRUWnK+vnACYpTEQmvhe9I6U/9nnE2zAR+03Z7VefyFDfM
3gkp6EC2g7r1VOL0o4n7o3zBisZf2CS/xrvw/QaI421cgd6vATwXEgsQXHjHp11eZ39UWQ2rmxsF
QuS3oBQAY3OwWMWplneN+T6OOfXDlHM9BSCfSgFzPX0EBbMrrSpPD6ITBQPT9YZ5QD27jugqJK7z
SWVcM+Mf/exreXfYe/valdK0/CxiPkf5P6JbEQxYydzkRpVVZajIKSOrsY4yscXjnNEo/evDmWfL
lOcR4fXgp7oz4fDMSd/Z+xs8qocT36f3IesjkDf6YFMMPlD3OeLAvPmQ3CM3PKZd4o0BN5hf1zhu
p6zaaWWrkxCsEFdYu7fiw5x9lk8UZkUCXIitBqW1kORk3+2khj1JUO/Gt7HjLwblMbsiy6IWfTKz
SHLTR1rw1cyL+RxhEmqfdLgwsh8bpx/rjGEkJrTXF0pKu2bKA7p4ILUtjJ9LQOOnPD3yRcWtqUYt
fGBbRYiub800Xx7yMLX8DsKHqJILjwQ2E/gKdPneRukRmFlF6na0NOBYGzgEccDcYsJ9Wgvrk3nf
5UrSUsuHrTKeivbYZqWXnu1HKjm8MMSFUHekEj8kzcphkCgVmADvfpBRcKMuCB4q0grl9MJlRq01
gdilXkdlSQONxo45HGkq+zZWKJfbyl72bNF2wLtKGDFuHgKNue3npgyCVB5Xado99dhZS1dKNdrr
qAXcsZaA2tJ/nW7zpvtVp4QoyJR4m2Kld5ITi5OYPay5NGZv1vgqvZgUjUz4oRXnjVI8Q0Z+L4pd
zgy9q845e3uB4ACLQErbgUOEsqKr2B8YpyZW3/oDiqafUWo7lenwpSzMB4KcfviKNViok9p1Skwb
yWBL1ZW19Ee5Uss57Tale+YPsvpaeI01aVg/xnkU4o8JxqW0f4HJzDo7BqMIZl1RzNv4YaTdI4Z1
Muy0jr2AGywMjXEr90T1CY9yN8TZEq8yKqvN8eq6lo9rfkkDGtGBhaqrmG9CMFh++4JahbL2lHyt
iRT0j8Vwat7TXzA/cVBOjtnKGgHymFojEDKOB0IYDljOPj0l8U+71HbfSCJbWIAaxNDBE+Xu4H59
X9vER64ACAZnygYV6LwMRhr/OONCsUFSF8M4paIuKWW3GZMdCL0E4dKylTeR5twTZqHLEnPaGuo6
dFVu0k6WTBXM4Nw2tg0JfV/q4JIQlZ21ZgwsieZ9vePmmvoxl/t6x44dTfoJWeFFSY0/hgTwg5Z5
qwSSuN5DZt2LGFa7RWl9chm0lTYqWKo2uYf+2D9yKbeEdrIonwtmTL3yOHcPJlnp6vgeVAubutJn
nuBqnD6LXDuShyPOJFBN4sscMc51SwihaFw0lfGIt4sQsuEm0u+ByDOWkQEsSe7Ov0hKkWgumZep
PHzrrGgkcso8SJriP4/lPzySgPazk3Av+DRnsxhXBfK6SJ4MWc2m3yz3xYYDYwIPOh9SZME7u9Dv
Wobdvp9ofHB4eJYfCyE7Q98+SkCWdQVUlUpZEpjQpjzpN5AE8qmFBokXXfaFB7biVJRilQoKdNWP
+gVsylGGCf/32158/h12cOvl94c6HcrLUzFUOpVyJMMkKZ9OHsO4F8L+BnDExZxNkr/mdHA+1X6h
sDJK5D4/iVPmpk4kcf2jGo1GGV76QAXdVzhDDIJvi+aIoTG1JWkgotFOuaxsUMnb68qY4g6mN2D8
9FBRVK00wnLHNDv+Eb+g9eSmQ8Pes0F6QiZOZRIl1GXbzNvFnc28I0NHu3i79nHAWU86w8+1VOlR
nCF+NAhHSVek4zUyYPtLuQVBM1CkyCIBKMzLNSyv0ND+3LMJ4xT74wg/FSZ/AoKPF1EHCFuB/6S6
2wtGCR+dSzQlZupSbLKsOqB/2r+zCvmfLi1ssRROAAsdLT2o4PZuecL+UYk3xJY8fcH3dJBdPyA1
HculgUXe14Dz1pK1l+y72fWFEzlKHucfnaifk3kdoEf3OggezfWediJbMfGNAVcVIiU++42jp0SA
hU6Z6rloCunHtoP0dzq11XTmvul7iM73GmCR7XnpZf00IJGvYJjneHTcbBtf2ffuC1qEcbif7KTf
tdoEeSa0jEtQDqOiHIjovXX3H6UrvHm4k4tZEJDAhQokb3s0VRU6yuyqqoQL/mlLGfQ0eL1phGVS
1FmUoXKRBmUSJLdCqzj5V8XSkcvflGKJ26JG5J5+mxPhhMs27xVxNnXmde5p0+8V4nbMe5eK3rES
YRAG/SD9RWNg9wyOy/NvQFd6vs6hXoE9OeqH5cAbOKZmq9k/mgMdBsxduYHbz4wHEJyJF5IYI7p5
z+QSOym8H3SGBeljkvj7rd1LfdFoy5bfLN5x89q42wuBqoCqVgK4JJqw52dmrsh0j7A+7uXG27dx
jtfx5ZsuqxoLYUFKLEG9tMEtr4KJo8L6caDcdLbjUwdTLptRxU0SVIZGlkV2N+HPloBEQMeVJuda
078F0NZ3r3wev63BVJgm7tSoTTZx6MN36rwJaRDO8qCAUEupTQTF53+Zks0wSjfhIFYB5ntdPNIp
UWbMbC4aDvPzrJW6j+nvhJywCc8biMFn/lrEDzk0104JugT/cCLKqiJUOKosv9Lr+UpeCb6c3oxQ
vRN80QduaPBO9hmRbCk/gU3b0Dd0JtjS/Y3ayxlslosg6sRGharLsfIA/OA9Fdtiyb7oz+a67z6W
U7GPv7MG6tWmRVtU3f2bB6XVpBq74izZslADTVMY8UozjdTd0Zv84lN2nhC9KNyWPCq9yxTE2YXk
OEyl/HP+e4Zm0L5KgmLhbYdYDIaoP9SnEnQlUF9m5i5Nd9BGPZGRmrbwLS962yq1P3WcgEqLrDMx
dmpq2Vy8UDmkuE1vw0P/HIxETDd3OINdSagL63Y0zkEgmXMUm49rVZ8am6U2RuJ+wAeZSRpnw1nV
rzX3FnzeR4hVlYDzi8xQnp1V/vWy/uznMad2EvfbpmoOp4j4KwikNLARz82iJM/7DgIIQ0Pvgccs
+f8P7egEpAfkPoQpTBrn/lxbUMuLf6VTJvsk3VaHr8PQX1U657rNIqxKhPmRM5kJ6zp2sjuYL8Is
45BBS5YKbjX/EPXEcWWi5CLk7hTiEgYjpds4gvq6ygvuzbQpO8MhwN/ypmoKjjC93TNVjHKeV1pj
lIXgWzsdUYlL2Jlpiu/HZr9GF8gBkU9GtN401fH6FmsISkviTctohmXK4a9SlzDeCaN1iYM5XIc7
IeEqausZe4f4UMrpnxQ9YlSz2NnTfZWjnF96xjPydRRv8hTWSpHaj2de18w9lXe37XfLjW1V1GQF
NEHQ8QQ50dEqNnsti3TaH3uiYqngIb9pEkgghby8uLL3AAn9ydmprYPNBnwbiMkAYJ0ebmeWWDqv
25EfdsP/k2dXccMtSMrPIVSfSN9AFibMMgo51IRkkVyEa9ktpSqLZf3KmA0vH9FOJqb2gkpcCkns
iIRd582LNK2s1s07n6p6EsMfFNuGMgOtR8BDpTHXhNhn7KEsUedOpxzq74OoNTvF/LluJrO2n5sO
dNkpsJE0InoE22H+I6ezL14DBT3Bh47SJ3GoPTXph/oyk4CPw/RIsV8TQ5r3sO7qmIGhFX8YKZdj
V/0x8R9+S1/5VTUiGtp82GfCZIfHjuYXK/D+0F1Wic1m694PVCWJaGAcEA9caTNWb1Z5wtKFwu7t
qilN1wks11miWDiTES0R4BqPOqzlzvFmWWx/tvGc4WF75VMPRhJIXOx/AfY+hPMHuByzNK3GRhV5
XWKqYQBjwYAa4ZqNILBHrpOxPJuvAWe2PwKm2HOIjSci6Yb7bYwBWYE8PrLT3mkDxqhTBk3LHMtW
ozkvKvZJcqqlRR6cFTvTugWigFU+BwsOBnVv414SWVj5e2fXNIRxqxh+Ti8uBsXenrqzj3OZx7DO
eiQsbEzwttWYdXoJIXK43QZ4SKOHwqCt44Ro/tWSiPE3iNsh9LVzwwG1YaeLh4koedyPnIcwf2oO
4LEj3uaBacl+soWKTXb8u/tF8Oqy55HjG/QGnmNSqTEFa0rtqEjlpXZicem6n3PL+WbUIV61fIOR
05RgzCOfSVmeydh5kBRPo8/QZDwySMLYf5HHlAYaEtZxvOwQ59sxdVBltVsh0W61U8eZYR+mBN4B
sqb9lJM65cZ6Y1dtT/QEWsiki1rj5r+AruTD4J+f9PL2uMAaGCTs06P1swOJmrGTj1KL9FmY10T7
0EOa2dIHAppKDseUKIiOMbOIRqbycvZAAS5r8YuhGX46N+C/dZO6s+R+orYyd9wg9QHhnXXj218Q
ODtfqUQrcDvo9FJ53l+5IMlbm9763mxa9OWjYklxBQrA1aqZpmDRavG+wwzuFpGwSCgN1b759CJw
0iWTABaJuB0e/Kb3ceB+6YDUMK5nHAoDQ2C6v7RLRk2h+WQkCxu4JVqNzU9NdqlIFszuZeuMXQuD
xearuozYkDZLF8ZIu9Fb6oOh4RfkqWdIE/hZ0xTOT7Ow4Mpjdqn+qBpmwGMD4GKC7o/qfMwG8MJt
+cFYZi01DJAs0VYR/KEa6tAf+TuAkc3CJw62dgjkHOZGOH4s3GKr+ePoaqnVaYnpdVbMt8MeMqT6
15SXHCEiR9+klO34er4BxoGEY4vtF5lE0M+V7FJjxPl2krgvzdRwfkQ2iBBayF7jZ2kcLLaqP13Q
A6OHPR6GkA36kjHqdaIchHAM1Uto6da9e96VByuHq5U1NefE9Rtfxvuj62clxUUrZsy+lHoGd7om
BguE4tOKl1uySVnEMubXH3f0K+IABc8gmMKb3Y4O53DajRM5yTU/VKESanz/p9SyBAp8kA0Y2Isb
WrkqodS6scEPalLznSeTuhl2EJeGaOOsBuylB9isj5nnM//EekLyDI/QJqCMQ42CZ9IPGxqGvirf
CQjh9R4NrTKolhvb2QL2TaSwr9NIs7xdR0I2oLHzM3c6SZnmvtZ4MLCkW7ECUb+WmHrNUnCf32x6
9a5R48vpAs/via/6JDdd2a6yZfcnHK0bXGp0M2/wFIbaKWcaYYL6fNyB35svfE13iTbjIj/nwS9A
4Fnz8HsQvktfASt1pVipObqhA9lF9IxTNVNIYEuM7EdXrRyxN4h6OyWQfPGJU+8/nEtRnAIYEJW3
+lVafW/+efr5UuRfCcOPHsVY7TBY+okLktXk/YegN6TbdGfQ+wy1tQaRBspu33CP99X0POntSRo7
PHr2qcWiXKZslKXfBqkeCIZVlcPm3HSPyk72fmBbU39uKmBsIF0ITvcrE4ylHxJTzF9rh14F5pvj
2dQQqgDBsfxpqInaOL+bT16A5xcdUyqJ6ZdfBeFy3nji1yplqU4c+jfw0BKr2pCkxQpOZYllTzPQ
djVYz0o7SxJYWZP4qj+UitUOLwmrt9DeRw2bINhVvxoFBqoyUaC/Fv7tMxU8iyByj1G6buTfrV0u
qMyw/mJLySi5zmrRooi2KLkCl0BLd60/0CgPWNT20P5ho55pyBW69GHgStdLEu5Zcl03CsgxVKzF
qCHW6l0eKLZ1Q1vXvG4S4ih6cPT2L5zgDnSrE9gZyboU6LdyPRA/otXgGUPeK5yRJduDkGiMF4rX
SAX0+2nJZsWjwBAzh6iJV/SNZUrwmUKJr+O7a6bTGVJkYNsj61uulHjqMFG++I9KVPuWfk5P5DBq
PBL5qbcFsHAV7+vOWjRCwM94DIcDt3TuaivLaxvzQzreB8+E7mOM8Z6j1/ZPZ54ESz4nFYNWc3my
Ms6cCutpl3m/mC3jzXLyw5VgDpNJqn2mWdCcM/evzckBJ0G/e7bZqFoaa+JIWKuiUvX0ck9edNsy
RPi8v07KPs7AEAx+f9IXNSrhVPEJ4nHRK9o2E8N4unXN3ZW5QqC9hyy22e3Kq770bAe/WKcJTqnc
iQyo2nxjA2AvF9vTPoZk7eT7U28NLQ1t3puy/W4YUNmNFJdriZsWi81OfUv8wYbyVr0jp+cpOwfa
PPVl+mBLuf3VIt/XtL2wgt3tlZ9Ed4TPhKvLjXXNKq4PYF8I9H7wjskI9JXUGZZtWR+M/yc3+qSM
XPv2eJ/+o+LND/iUG/i/GtQMU/NVggkJd3rYK1psHQwCMfnEQNTrW0xDqcSHuR+mOofHgyYCxFRJ
ty4Is6Bq5wuIOgcscXzeX4rP3z+1ioBTASpOYxoP/9pZ7wSQWqcEFlYvTCFJMBnRSLmoM+ivNfLf
1/OYRszjj/HHslOxZKyGr4Yyt8FPGtVEaWqAJsBYAQosw1Wr5j8rmSnP0VCac+TktnfOiwrsw8uY
bPJl33pCXSMq9J4PM2+63ArubQvEfa71YsFOSbvlapqBByJXZSZb2UjjjLNr2IAD0SScBzA9Md9K
+BRyEJ2Tbdj8Bmnir/+Q8aDUZ0KjJn2f6y1Rx3D/9vdckgfAYamLDyDYwAeQjkPskauJwxVrEYcj
9W9iJM01/VrZqwgABpE6MFl0WRtcDJt874MBDXrBUyW6U128lx8YukVb9darkt6np4QjmjtBxg1f
SnF4VByM5iQrwU3muWQHvLOPgsO2IWRgOySbQqP44+poWzhY0NcHkN5CQv+vIzI7Wym4uGQ6W1r0
ADj/wm6KRMmVQ2VJia8lR44VHm7xRkQJeLo9J0al7dUdmGg6ZuqTIh8722LMqXQtjQ38shDu/gPO
t5je8AhdD4+sOaKnD75zl6WnQFx0AymS/p2/1cFfLSvXEnto803P2odyulAJ9a7GlpXuMmO3Ckj2
yYna/OsM9m28O3j308pCxJLumexjNZBqlC96jxQVi+P8B24FpCSZCQq2oqQxvz2RaPrnTo4U/BiA
JDKJW+KsBBr3EKPpnP3P3yt35v+smMpg/O3gDoFujatSSS4zXdhM22mafMyeZt/iTuyWb+MakrLl
DkjfkyfJZTMkUgqN4y7DiE3gAIQvFODThCMMxXNkpXcrVbNeq8ZO10jmgURApPLdLP/8tdFLijJ9
AT/qWrwCEcTte3MdZKapXwwq917iOFX9Y9XMFj609GoxfT0SHf8yNy//EOvTxuI+sKjXD/4+gBoB
QLhNGDtkLuXnOmYiiLXzQpesTV2Z07dCEcg1p3nVxpHTVVrDuGznRRfJCpqgQOS3YPqg/wHX7I9m
6n3uuTTbHIucrF8+fZgsgb5289MJkIHL5kpLHJzPCCNf0CiqUGo/ZicO0Kzx8pSwUDM/tuOZGS7v
9Hk/PDKS0KcnmZdTCq+Vtfd8pokEm2uheUpJ7s4Y7A5Oxy/zLwYE9NcHuqsTbaYDuUN+ekRtlnx7
njyq9LNLnmowhZH2DX56ALl+HccbLaqLVzj5lftzwJdNFGREpPlCq1orDQbKeTYIVaq6J8tdI1B5
5y172vyhXVlrwMwBR96AOi0Nj5uXx+dagSaZZMjSWqzWVdaFaqBGfk19lDIhm2LHhxh4lUbRU+oB
JZsUT8A2ATW3HTV7VdQmGLcnqZuFRe4jhU4kfrByp1plzDjIXmAnRc4eAgoezhgwC8ApvWjfQSc9
sT2VWeJ6sY5ApoOI8ydBFVZXjjJcBw38XdngpF061VU0s1TV4BwIQhY2ue1fZynZV7dlLen9cAe4
KEaBvUA7dkN9Yo5Ki1mg9j1PRdDvvKZ3SOeqAYCPrn3diHrwIZYeoYJToctQ/ZKQdVsA2B3XgQZw
YEGKxpo4Hsv1D1C9kJx09iUExiixOSGAAfDa4+NGtz/T0Q1MJs+r6ILaOMXlQ/1Ybvn2IcHCkARk
X8nhtsKfOcIHaOhFJ8ZBL+fQFF7z07HtTqZnAHOTVhpqOuH0euYxgya8Chm4zUEaASqToK2EsiZS
cY1a6MQlkluabC66ENUWic7BnpOw1AGneUFBCB9bdF9p70UE+mcBnQLYQaNmWSqS9L9NG+ItUdIQ
mmxcJHaUGuY036oC54yCddHwcmcb+jFV3T92GFagtlyssqqojCDKxVgsRWtpfTYOb+YLveJmtZoo
NFHgXEXtSh/Xnqmxqp8vzyBF/lfRFJ9K4qDP2WGiB9yuOkxngR5O55DiRe2xoH0MLx6dm/srY4HO
TD0QYdskAlDs62iUf5OZDW0mS8pa6beBJ8nXI7C6XNFVbkzVR3Bn3wFdbXV8Sz3VzX/iDtO3xp/H
acm3YkUTxFCGkvWa2Bqau9sQ+vVulqS9OpbbNDUp09EfFZDqd+13RTlZ7Si0vYJYONVENnKDIzOf
8J1FlkpAH/BCHXYH/RvfHxAYPB6ReN6BxyWj7gLOo0ABCazQ/XgsVbBX9YPG2MbGebLUJhr7Vtn0
LyMW36h685PBIzDVfJ8RpqYLqCDR7CYcaeBtIDFoR48WomcR7Il84A05kT9ez0FmmelbMWToPmAJ
QFk1NYDYoPaoECmqR+XNLFVNvYdyWc5Oo5zFFrBieLBlgwDHpF5BEraY/P6u5OZiNM3Vmvff0y34
kolzmQZIee7w6lWr3A/SY6y3D05l9v4yjdRV8nsK9Cm6SITAWrKq3lzE2aEeP/jBgybj5FSiQH2C
dsAEJ9BYAwqQfsqywLZCTK8EqiBwLAriDmlrBFHTeBoY8vZF6AYuDz1nYiSo9Clc442H67LgXKoj
7CkEcr13MVzpnKngbz3Y7oIvMoVtQ8yfwLk3pkef5bBhVkKZIsqKrX8swG/YruLiaHWRlMV6lZBZ
0gQXutMNe1EFfwJv9d2d8u7qhnt9r+h4OqfKIddQxKtCWruqyeQTTbNhIEsHXq8Ufr++JPoAptAh
oi7MAkh87wkpyuHfTEV3JgGfDouU/Oxtu0HEnoitImTSEdE6tjMiBxzKyrZc93KWq31ip9zuuIqP
MqfgKazvk0hjQUXPLofFqYau83nUl71wvzEaH4JUJe99ps7cRWgT2z56rEQiH4SQLDl7hGT3frT8
AtfBFdSnyGdEY+BxPxbPZGPUmQrx6hnzBJLNpUwrxXHZ/5Y22LmAcdBXzdcAAFbyOSyO3vwt85NW
Vdidh+WCKRNPoR7OhHYuh1R4JD/xaDPri4DyKep3H00klI42veX/E9/EFWahGzAol8DvulMaePDh
DEecZiRGN0krup6cYwBasMeNLCKCJmfI2mxPKnEtxRmPD+NfkMaye8xr2VShGUEhkqL2byFpeiqV
wd3j8fS9GHxjF6s3mpspSudMppZROjiV41H9f984BqM9sJmxqJ0U1P/YaFyq64gToYHGjloOaKH4
3u88DBmG4TckznUDBtSID/XNzfH6fM374ytkFsEsMlC6/CmJffiUbAo83/WeuwFpTk00Bjgf8Krx
c/jXcx3QgWqutvV12u7Zo6V7jXhW1OSG01f2Dh4JDn7fQGV6nTCUncR1KnNxYDwCCsM7VFx91j6B
MD1ShdL/K2aG6hUBKbFTweQ4iZh+/xv+aey/rVuxuMIQv+RUpxmcFaeQ+FQlAl2zfXts/ZGvekX6
JJ7XJAbQMbpZqPjolaASQQ3mLObn1VYjl2nMchd2C7DdxqAMk1mhJlqjzujqnkiTQrHsU8/Z8aZB
6QjJyzkH/rQWYlGOeMlDwFM7s7Kk7e62MbuLGa276hqzBA/rl5mnS++BKvK+QNkT2e/Mb3XCot3f
7YQUQg1V/oAb/0H6n0RNtBJB80eoDC52asjz4y0qaysRsY9AweRaqO337TS6zs/cAySKmjnuRmH4
+pabsVqyEayR6CzEZZQmXDpxVT998mnrAYKAH7Oe2WvsNovbkPjvuWKYtJwKJwPk0J0uSQlVgg3k
5o74X8vnEGCDi35uBIM2gNv3k+S2xMEx10D82/aPcOaqQm/3qfuojTIycAy2t12NJIbH/Y/v5g9e
S1V2S2jb7FnR4spEheFazyeeHiBuN+74j6eiGn0oSPDamIXBkcUclkbN/QdFQhddI2K+qLdDb1gf
7Uxa8kMUn8KATLrkA67poq9oOaflRKQIh8LW7MrXWU870vf/wCu6J/BSyvONF3jrbRJQbfFAKHoe
RQuggRyDpJcPZjHnTtzFyrJP9GlD58904FebLuA9VVzg3JyGgV/vcRLYp2kdVBv/5eJJBohbBJES
O7hUiZcNOujk0XIbcOT7kKbLGEQ5N1CwthxvUMERAOinFGwleHa74+7CYxsF4gcgqm96Q0S9kb4M
/7AHNIV5tHjpQFezjNqlgKva0iPGJgxt/lW0qjEHLGUIijOpA2AGZbyYS80JiDRqkvGpas9nCwp4
y6lsL3NGQBzHAU8w0T4YaxlWvcPuRNNIb6UPZ5iFfwdQe/6snQewKz4ofMxLidwcX07lYycfmSyI
K0K2R5i5BiPvcGyr8cW7fpsRJUJNMjuuOpmbqgzfSdCeJgD4nB6gxrB801SCQ4/H0yu3x2anYmou
6pEsFlmoavsitstMbtHm055Xoc5kMn3bMGmyWM1xOVEA275mNE56JCbNg0Eahwk0PIZUMNB33jKC
Zgiisf4kRsz5HuC4746VJ36IcxnlKHrfBCIF82kOJ8R+7tBXw2DDxUpM1iy8w/gabBPlh+FIWHSL
pOYN2wdijgWCPyLraFzRjDy5jxsYklLeVqmem3Kai96UzRpUyHiLSLUiBahCM+u126WVxzCiL+hP
fgGKosnt2sKiDc7jfmdJbzg6C2oOkILWZ5yZKoVFWHudqymmABIWo6drM+ltcEW4KQYLIlKLZJeE
P/Y8+KUF5GTyyCrXkwpYZ4hk+KiJ/kYGod8vpDoY569KARcT4iPe+pNHVRDsIgQn8B8OqB4RRKgA
zZiNfBr/6mNx2dlBWuLjrQFHFU0kiBOPZdiyHY2TNcmm5ENhLdC1F8GnFEjgZ+kXH6DNBG1g5EsK
olRCJrx+c436L2b3lHgsVNmGjq2dGySoN/Wn/eIUqjyAItliUtZx8zQzdn/nLaVUB8pVWCtwBnI1
imflxnJ/RJOZBtjkj3Fn35wA+cw4L1id6eJ/r0rCfx99Iadu8PjecLlWrIM6mrWNelwSJBZsljaN
Qh3xqzFHnBm2KceN4NgeLwLbh3KGfToax9dqmmBhOolmdht0nW+ZR/HKhqyNTF3svq40UqFstV6e
iUOAGIipNP9/IM+3xrRqMhdURdWuz2TTzIqUpu2fR7evXVMopxHg9Yn/Arns5vIlZH6p8TL1MtlB
cMGHtRCXKIfO0TBwyodGHcfI6PUk/hPfcmHX+NG4YXdwHYfAP34EQbo0P99cTK3lok/qcbFPdvL5
3ukau/2ZEdoCRWwQX3UyjWbvWdGJWPxVYL4fO3kuJNUVOs3+CP4rdUKOOU1FX+6egopWsUjoDa8R
PNfEi4sWb4rm4NWoEUvXsOaZvFJ+oG5G5h3HcmSeX156zLdydLWImHqQhmdUmtvu6X8IKeKZQoFU
ur/9G+bF8GaD0stJlDxrEnFSN5vxwDchwMICRpDq32CnU9ypxF5cH4+Gl7JsMkjrxf+nHYkHr9D/
U1k0x4Gda3aUW7S1BCSINcwNRxu/RjKjh85YJQfkpS0PGEGwjuIMsTuE8GBbzXvc/H76vCIJGZkr
W7AE6MMkKItwyzusXXQ0PicB08nGZGzbwl7k/bZcVF9eUJ87eV3VJpKHQ3H7vESZDm4n/MilR6X9
aUfGIwUrMZuk9Xhp3e+zPkEl4Z+JwyueSMZ67qa/eQ0F8W4qvYsm29TetU6euSUNvcVf8IMyA8te
7cvTEz3nOtp+PFxMh+lm+xDEF/VRu/fdLm3hPO1K71+kXBHZFNze7deNjlcWTQB738qU2Q8ZqTgV
6Q/L6v43p68r+kfW+w7jELKFMHdUzUmYb9dUWjXXuHof9LKISD0CTeCB3WwL603zMrDE0CmxC9hz
GrlZx1jixVsHJhyJpuCthxtsSeM5KTYKcWV3x9u97XqkkaSt5f5j1V8E3nyeLFIQIiTuos42XfTv
9B/iW3iroBWOz6RMXRX3POGUIHJrKBp3Gteis4sRvT0Wp0gcBkKrYU/c9HyoTjTsR4qid0L/BTT3
lmvd1aA/Hfv0TDOUNIo0Qic2mZm5ckXIrpZic7nFsz/6ik0WFdvWDyAWf3UXPjLZIpgynpntiq3T
V+QXPaB7KaQ9dGBAKbCKZeA/1FHuGm0g8zX+o2cOsdWviV+Zo5x+M0iAVdV1OhNfmipulK/ygrVW
lYRctFhVDxgOWOqQZOcYoZjS8Nm1pDQAF0N25zH7uV2gfc1dMcp6yjzTMMLxa+hvqS4/NI0iRiiZ
RGIOGugBK8rYRvLYBfVc5YzEr/cr0K/Z14TdWmPFe1MDZUioPYd/OUeBDP1yCZiXuDo0tlrDhqhL
caJOF9VS239fLgqOG7Qd79QvuyeE6FniuvALxn1oMeV99A8iENFn1cn2VCyKvvqzvZQzEEehRlFe
PW+iWFuHrFP14/JWomlOaHGYwoIw+/iZvfz3DDT40c6jCgVzEUSD4bZz9oikLR2nAI77ZnXfU98w
y1X3No7cU1nb34P5M2NSWKADKBZyFiqUnPkBJmZmaEkB3rS0idvavIDIZRrNoXGhmIXurCZi1YQj
On/BdeRHHOZ4XagHLQgZ86A3p0LvLKGNxk8i1YklFVfwl0lfGotcvA/mtJv7eokd6bi3rV4fj7kz
TNprJfplHZg+gj+0HlHBMBo7ibXPAepq0wdc/ddxs9MuyJOVaQY/7cCIlm3CSL/SGzqDj1PjdwmJ
6sDtWG+CNuRpLbReQuborMBugHHCH+SHwGkrvZEzW7BS7fW0oWyOIMKUJX/VuPpcnG2SazRHv5az
heAsUBDxzpI2LNcfGhnC3bCwuE+3QuOfC8APXTMxLjSgJjBU+7VYP9VJIrWJHwUCbJkACW0wh9JQ
aoQSPOPcx7b6tM8Nk1I4adN9qA0idixpZmF+Trw5decAsHAOIhS4OU38JaAQU+FGvDZTghVdcslx
bMFPbDSQx42HmR4qFlG+yMUy0oRE6nY3KK3n+3S7Uw7iWnekBu7/b5cX10A5e81znC/6G85tXjaV
fMPk4FmkcgmNgSdRSNPrxy4MFt/+ahBDA/QV1e3D/40lSrFORe/kKTCnc6a1zWo+GXEM4tyCT5V1
UN2yr5h/xSZh8FFaPJGymSuHFHEPWxReMQTSDRnJElfjbakrZgOjIQ4AL6y/bniqH/FlgjjR1R7O
koI+RtqfO5i51fZzpD+PsJI+HeDrcAujZ11FaHsl+qnH0GfkZDnhzgdworoeI8b9uJzn96MNPbZ4
z/1NCOD2C/e29rdYvmnSAAJS6G4UoN5mmYIWx26bs9lXK/L9s9YXuDaXipwflWIsPy6nQXSCW/+0
hZRE6U/smdUuHdHnAP3bmyIRlMlaO8592q9t97aOBAe3uPZEcgSYodwP6D3lZVWTCGp2RnO8pXS2
hFJkkOrSC+1E7v+bQSgIAN6pFTYsEus9CPnCkVE4hP1d/Wo5EL82DSw5uRDNWFc1aSJpIxaTVezZ
A3976xdBjLr79hGVbgMn054cN1CnOEfAgndcdPHIIze7OWdFF5UfTAXz9k2ZZcGOsUYkfHJvcLDM
1/tPcBILQLzK2bni0RcYX6iP7bihJy0G3PGOr3gthfQWpBvB79euiwRZlMCbF7xckfZucSMjALxC
0Z9g0jaZ5oLp4WjYDvau+xb3C4eiczlcElvNxvflv0GpY9WI5PbwkgZv6yJG1C6AHsiZQwlb2rmP
wiWQbDnW5KQiXyNRwgRIIjFv63pjkk7sml+VUQGzfMWw43bZbLYbCzgyzpjJzK5/09NXKmP9ObX9
XqcRFFSJ4zrJWxkI9iMpgSGEQSgxQmnbYc7DoPZfWZ+fdH0CkodT9Ft44jeDdcYmId+VJtawC64j
ep0VBSoT8heDgsVer0Hamdyt45rOz6t71Xl9Ap9ujUJv5dzzS7gNBQP0cl/h7asG/Te+6S9fT5t2
4/6qW0WJ5SRdDWtSbAIvOJj5DazG2HiLsRoV9dCUutToGWBQXLtXGHpjMu3RvkqSgnLvlpp/N65E
bXH0gp9tbNmVai7FKtyAvf4W81i5HyjyIWw5636xnZjckEKFIkBB4rmbRHrmzLsoQop3zDF9vjVV
jHF3ciRAYM9mmeDYBPTZSNVQNvjFJyE/qj5QQw16LiVznUwSvsyqkzBYJSaWmW6l5cjUSRtz86Yu
ikM8Y0XkGuXZpcN5nHd8w4JJFl6lKPLcivON+qqPp6g7CXqY7j0z2qkv3Pbhn2Ny5Xc1aRd6AIoY
OCAvEJemDiIPSnkj3kTxZX0rXHTa0IhHfKaoh9BTrZjGO2G7VwtXM+BJUI1XzHMhJ7v6iDtJBKvw
dDE24bGVVMcPegoft89FhSlrOTvjw7uTe3ME2bm7G4P7E0R5TVPBFwEEjAIe4MFHn1PMnrEqlTFx
TD/47VSSgII4TAsPwkWOgBcqPQaF5gISDZp9LU+l7T0f02Q8yTV+RsDnVdz2hjiyw1vj7NiRTF7J
oaR6w4LMNGldlRfr7pbsEQI/Crk4kle3qMrzA+THHXP1VVSI2c3IRcsjPxUls/E65GMDOtPC7LAl
v6tKZpY2Kxf7rnP4tQvJ9CE+FzwvfT5Ed+TAkvwA7BVhVIk0hc1JoKjlSm4LRMWlh0URUMcrIk9c
aUN8kG4JU3yT7GIKmAfmlzCW+nNCPLRLbW7Mnkg0RI0ffUNQIwBtVm9wjQi8WNPXH/FUQCX7tLh3
cf4U3BVQkT88I7xlozkXVdwvQbx/bxDou8KeP3zZAsEZSVL8ZztDSkUIsDDXgHhgnk8PYvCngwBX
xGNGiQ9QstirtSAmnQO7VpIpOj+P+w+oUu9LPqIWy/xof6qXPSL4Dz1tgbNHdgk2/uiSS10Dkj9h
q2/L0m2ESI65rkd6005smizhuNcfuxWzhc7PUIHf1nD64GTU1JZ0IV5ceM7OSjOYCpbKdqA8YHYW
kDNjVstqCB5PY0dFjVAuLcE9NVeM2hjVszIN77fTCEw9iIFw7mmoGORv5Bfq1UW0eCUzVP3v07Uw
kAJ3iPLA7LdG3GWEesVzhT9ckDr+iejfoQwvXWDqiPgHLXpRFsUjb2iqulUZIwUG9F8QvjBI5S4m
Jo94rkZ34yTFAIv9EzZqJyFZ97Ni/Po7a1zUKr7IAiNqeyabWZ/B/ept5Urx/XCjyxPYwl0Lywlo
w6uLIToiMAuObFtnjIykrafU2WgpoUVB1fpi+CTD97VIIqdo1fMQqvnT6uW3kge9Z7hZbhLG0hhJ
6XFbrcwZuXImJ586bg6BlIFhieL668IlUkjWn7E5iiBL3wv5SlKL5r4NiU87G7kvxmOm+7EO67cJ
5yQyLACeU0vEx7dTHaQSC+ckd3DYquFhkjJyhFBiSTmtk8EgbAJq4y3dweshwu5wZYF+Fd4yRPNf
nv8RR867VNFfkhdh5kyj+eENnalGgRmx3xY8NpW757zCiHuqOSZ0rvmAqQInFRmUPF5uq0jMY/vB
ToQcRWQjidwpJ50V/9fqQYufoLjVz9tm0+sgi9h3t10I6WHUj66y6SId0NZMkG+JzfmQB7g3qCZ4
ZOQH4cd2aiUlHWb1cpLWiO4r9v+KOL1z+3Rn0+pt2P9LneYKpkAAu1IXmjAF4/TU8J7dwgtg5DeA
FdBesYmON1jHs+jv0D2CLUawVSvMJOHbv44tCCEnXDk9DvD4rdbUUIJZCacTYGHrycS1uicmUq5R
kdphegH8ITrHywNnnNagc3lM0j0PE3u9sOKZo89DPJti+Egrh0PK2iGEt5OfdtX1u7EBkMbcyTEN
3bUBdr74Zm1pmm1XDuxaMkOxhxabZpj8odVT/WKQFfPa+JHWDHXNzGwts+ZtRAs0/UR3zRfn5w9d
gwGoSJZuF91F5/oXs5KmxE7A0HeTuNbUS3GE8AXDviPvvvwuA8Wdv64GfK6zsuONzogN05wvbtbz
pJIaWNZtXMP9CEOtjSpllx8mebtV0B5CJk2HUn04JcZLH3emyxG7jRTETkWgyvddDObyI2CDpdW7
p1G+ndUIAnrKCJlecsTm9IeSFSeFpzNTDUFuYX48ofd3T3fAvDq0wucluoU3hWvkor9qffBRESaF
iV8SIwO/mIqUbCzpbk9vZlHO7i19Iggr+un0m38acIHNRiLuzXuavz1Rp/LLczGbvw82rmjcQ8C1
zoE3WyYg66SzKivVjS81e3dif5+XoaD898JZ/XbgwN/VwFagGUBLLs9coK3cmBLLqBfXkGG8ExON
+srgi0dob/M7zBwkgeq/ps9xz87TIRtAyFNuOCCtiF00vJG17ZrXxHn7SUGWpZgPVUHKnofr6nwn
szm4F/5C6XkHNSBIrN1eKugWmU0pVJH7LMbQRW0Pdxj3r5jeC70Sw0GtR3oE1r5EuCidEEt6rI5N
6o56kwz0mK8AL65rnljOr2Qcc9t8TPz1KvQ3WxhUK3SFfGHlbGoxlflbXhKdJ4fQxT3cvizxf8f/
I7OVRpbiiHH8CLm89t1jrhhycSsIvdayDHBX9YHhkmN57fsHG+fnKwpBYWXWw6KWQKH6C/ZmYmDT
ljoDAaoOUS36jQGG7arLP9JPvvW0n9b7Yf+4oIkHa651+5CNAvhFALc+x7eSgpbB8P3cEJWY2qa9
bbgQMDkOc3JfODJC90vqw23M3IoSaMFxa2WrQQuMcOCVCqo57sYjhXpaNtw+OeM9LFDbBRWllccJ
NETeCHaluNojgZKGYeshBD5eoJS1tWX8N4Iw8UgqIlTQnWzgfRcJJCYk6ig6G3dxRdp1r1aGnhJ9
ImA0ZfiHgyEJxVOXXMIz0+ZGp+ROWFgF+25+6iwtsz4hw1AYA8sD1UJAev87d4Cp59pvWXB2ZscU
0kwESlluXF8HqmS965HQcpH0sKEEHjM9D7GW0hFpd4xv0RndqBzwvd4o4kZFmIobK6SgGUzZjDYS
Z+W2S5TzWwTTCw34bcnNGotQTNL96tbg4iDLxgd8ocpXS5QJyaDqkOMVcBoX77Z5MQEGs31HH/CU
S93B1rIdM4jVPubUduOkuzsKiF0DOb3tA1exbkmY/tpjsYsa0IlzEthGHPl5Ml6K6Ve4Fc0mIRvB
324PszmA3G0tAsM8jnXxYo0iplvISUlMAZXCdjzNn89Dok7Dr4mDHn9c4kbmy0+y6WmaQmuI8rMe
xc20IQtuPGN4pynS7LzvYhBMTx/qSzQMEOyWbLpvIIRS6AEzyL2h4+D3gFH8AtUQqEtwIdpE1dSZ
fenoPc47KLjDMUZ1ZTX8GUb2aNh+cUvYhFNN2CS/arjDBh2IS4sIeDc2S2PrYmsLtpu2Jd036bVf
+vD17ZlkVO+YK2ZRCfZQTiqfWbZd7KwrUJIm3QR8qHnXbmHm9MlMCEfLmRkfcSu5h7n88FPCPNFf
ifZWeYeIk6U28VluRToKhxxNuvkFerJAMH9OjCLcJTVFnM01/VY7lG/nVjl59HsAC0pm+D9jWElg
TyzFBssEHYpnjQk9eI696xCsW6TqMF7TsWx5WNPR+Cpobj1Thg+nLOyzAB2kiumXwE2Xc41ZcD+r
FeoOECP9eHmaaBohoKCa1SvLjPfISELUztm4ap64YeWyeyhGySLA0pVpkV9C3BLYL3QLxEY75ju2
qKZ/JedaqqUdKem7UzoAgW1G7q/d5/0HzGrFKGYvZzYQzuuuKhxVAcHvzM9W6iJt0LWVh55Y0lRd
h2YCJYeMAg50Itq3L4JB5U0SuQYks36QNVBWmCkLGwfvP7msRnCbBlfyoZwr0OuQPYVKniyLlrwX
xuS9zLyT3NjXgsZ7m5ExRyOoR+iD+3//OypDochYQMhcfrpK9HVPnkcRCF/dMlUIntNqeoLzAVcn
xiSzjR3+4qHR8p9rO0d063tQ5rtY4PqK+b0CkNnHiokaHbDC1c/oC7FKF8hgGduSZOW75AjDDPbs
VJCHPHzdXA8W12aPg1cnzSSzWo+696/Kp3Bz5oPjoiWcaqvJLmwCfBJIP78keAzu1/KhXplqNEBM
pnKxRmumL0R4QvX95J3OEu4BrkKNBDDoQO/Mc9SgTn3Fl19iQ4km9MPegOV7QrEsfO9gh0LeH2tp
jiWT8rpJExUDw8nSEPLddE20CQ22qFepZHvxhbZh0fyvZKwKdT4UtL1I4N5RRhl1vDAZfTpATeka
3Lmrdu2C8WETfRSrrL/X5sNIwEyqoVDPMNTRTno4GU1pmixS5ltxKEI6MBi5dZoCZis7G+ttBPZb
5+2yhPbwcmGxFPD3Or8abqHTJ9GrEljaljUHgBjuCvT9y4MF6G01C99q7ztCnSfEQT4n2J4U5mYj
IIyy23p5S5C1sCL0F2hPIDN6V2k+wgFoR3lOf3Hdx4te+Kt5PLaUMzbgJ1pB3szXxEE3dO3B3Uef
jX6nrs4nPMQGRM9nF/eFPTb10wj8HOAOTemxTVCvU7L1cNYz5Jnds+bugebu1qtbcn8Lj6RGXMBo
m/ct9r4qeS21ipqZIjV0yRVuQg1wi6IxB12QMnwkMoU0EZFfBOmdeR1ZX8RHfdB6Wz1Qrx9KwKyn
2yTcI/SIQHU1WY42BAEJEWg6ITUBnWkEv3bt1WAn2RvgQgdSmSTj9lNXxHU0mlB2F74/CEOFfvRA
FpkB/uWbCRt/K6Lqkkde8P9EBgUGU+hFKdzKLbUVuBbRPM8+AWh4/Eazw/fugbnJrqhHU5xQT5j2
CWfB8qhtKUaZFUlENVFizXhKWcVTxNSBdCR7o/RQo9bLhuan2qRWtiWub76ZhDnsRPlBQ/AUkgOJ
TbvUmaFxC6iioYXPrKLPNhFyi64PIYyKAd/UIE7ca5/mYBN8fRJrslzCB3Iz2FdfQwOlObclFLuN
lciQSrpz/yK+j/1x71mzEWGFIlL6C5DfYssUX7c8e55RXHRvYM83N4qlmuu0vZ/4W5h7NtmmQCfG
wrWLJVeg6xIWazkibGzW9p74W0czycG6ISBLfRX8K7FEoDhPTZQtNYCfmBglOGKcUz6/WKlWTXsu
2f5zsz/tTSo2jzo/6ppbJfEn1kLcm6eNXO89UjiNpq9kJdVDk4jJX8jnKWikSsuLI+SyjPx2eUzQ
Fo8s/wv4Tam0SgG+F/E4nJshWXiFlqxwt7uxg+1/UTJHv4c43sR60eKlhzkfCswd2RBhr2MKNQQ9
eOktU9LpuoP+Uw2OYIr4SxwbaTeSAGdYXRcd48eQCU/Sc1WE1Met/Y9BjL2K54/K+LaKviz+apoK
EYja5CIL7twRcpbT3BOYjgj6TuUMU3pQsmByPc5XVNxof0ikcOf/eQqaAODCVijF4uOfy93Ngail
8E1slXQjdytkCRFgxZYUPA8lSP0PlwnQXBFGrYw9dk0UagGwIyL3kNZ8oMvKhDilgTINK7E6b27/
XxZ7ZhBNia+VZm78kwGbmACyelvmFaxXec3I2RF11tmalyYFuIko1f0OMfzNnH3Dxna22vu3Io/Q
7M3FQKcpOn/pE1+Rq7yjnKpmDjf0IVZ+33zD19AU27obOdrUn10JbUpedz89Qif4YaORWtxDqSLb
x6ppVSBxtMShMU4usdnMKWmRrrUTO2swHOayxHFTCIMrdG9VOppnt8m0tSU+g3BJ4efRhEsPDHHq
/xZ0MfNPGdsLKAhEBC9lQL+8O0g2TVFOrkMUKuGJt81D4KuOTaiaVJ0HksZczVlNS0PY0Dq98gMw
SLY2gmiyfk+f2drWdhiUBJKLHKmlguuWWd2rhY0u5alq5QZ1+tsc90fQ+2UJAMpOVLHCorj/66ww
0feEUW5ABPam6E/9FZ0ADLDY70epyP05DG18McDkh5/iArI7H/8qreu7MBhfgPMJgURPrdqWHJgE
eusHe7c9Ro1DSCqx2vaf7K8hlj2b7ILh1uhrxz8b8kKuB6M7FMhpr1PPMk+ROkAblANEHlLBPHcE
Ep9OVt8Q9jNxIY978nSZM/OPbM3AJntYUuo8iRpwsS4dAsPDE6/vOhHpdxMrazWz5w3EnCq3NKcD
nYRjxXPVWPQFJiZz/4S2sSkx97Pshq/quTrh6Wt+okpEk2Zb2MqO4Y439MyzIXgoMoOaMuIL1qmB
8aPmp7N75joSAn0XLw2iqUf749VWjCTX5N12WHUoplTop2xrUFJ70LgZxUI449aaoNeOn/FucYcV
tIHhJDoj/+19sUzT1Ugb0dn9GMjlFvfrUw+HIUOxwjiDj2inzsj3NGR2qQKJca8NPX1NGWIiAHzU
yay/4ojNWXIMhfTLVGq3ij79GuhQCK8uDgcoTC5Xc2xt/QGPVXaxlmATUeXFoMrfnwJYzc4diSbd
tKsSu92QzdVlB84RhbZpFKOSbA8BXUPdpYLu+IrEzUYSeuXA24eFAnXirokHFCijwVSUxLJAM3qO
tVAkQo+1vZCDPYpxG9juW3uD6I+jKgEZt8GmvI6ho0bMTvfjCmJdZ3lIyM3j9GaPnGYTriLDYDJj
PWiqNTa3anh5Po8XeFXzNxZHNEIzIQEak0KPL2/LKAw7K4spq3VJkoaJOL1gOczZwLjSRbi4kE1g
swNnvwJesl4aAwl6wkGyIEq39eG4jZD+aQ9NDYxXtOICkTFsoe0uGPCfJ9L3gLVR1QWT/zKvyRqp
Jhjk5QIT+8J9KR8S1kzCcRtcu/hVXCvcrDs146RodOhRUL89+NxRgqSl+FcTcR+OSJBD2iBiAZ5x
uH02YdlCDbxS9Ty1G7zTE0IzzvjwOW1JL3lXmcMV7VfYw4/8LDeY1rWHxyaL2fhRs7D9FaI5N8nr
6CMR9kcqMZPrORWGgwT3gvg66bzulMJ0B/27w9eHoOzWpGHfp3o7tA2ZHycZyIvZAJCpTDaX0jPE
LU4kFWZ//yeixsyiV1A9BSsM/ucFz4WO6XkNkeieGvr9WnZQQG/sPM4Jjextw/A8c0m9r80RFAbF
EkLsaZna4+/6SvBdqcW42PA2sHRRC34xpORT5Szxe4zlsveAo0KUqJDrfPKjx6dIO5lZGRNVeW1o
pJkunaBPbthv9Gxd1dgFfo29zGbgeI+CHX+gH7lpLYiZKQbXBIpRcCxB210oJhlmsPjBBlKlj2rS
JBhgEibnvbxtVSttkpUfgdvnYPfb6QRam2gR/RhVwAl37er+eYgB2VIcTJ5Q++Jlctl1zKpU7GhV
LCM526aW226fo8hnV68r+fusJS5yBgACWU2gGTJF/WJ2OA4+9kwLIVkxbcu8SseS2HzsZJbSTDQf
KvTODuXMyc3kw9h6kNWvsjg4V5w22zvR2aD6T4uuR5JjREZLTNgGOXxeG2CiwCKkpXkN3hJrotRA
sKErhHU9TyLYF62YRL14yUit9orh3ynSKO4rksW1O/9S9QRFPFQdTMl2/lCjFT8heLArlrp10kFw
xUyYu/bVrFL0AjcEnZkFd4YwjoPZGQ5X30Y54n4ATgCLrawaXtRJLfZHEI4lOIDOL0jK3guaBjE1
+AqgYkBX/v1mELdTb0lUn+A7AOwCkip1ktbVBDWrGn1cJsfJVn1HQdVPlHae8fJwS1Le4hqnnUfD
uX52O+9hnRxuiZpqTk/hywv5TL8jIgmBlYG1Bw3ANeP2fKEfYlMhyVdb8Z1On+2GfgOOobC+IKuk
ItzZAeuVH8v5tON/9R96vA7eW7nkYjleLt30dR2TQBsRYijYc4WTU2nvkdaOmZYtL31mBawdTAtr
unceoOKa1nSNWHpZEJrXactImunZKSL+7qU5Il47jTAzZMXjsQKcmQIL5sncu4cIZEMcpoIQe/eX
KDnu0KkLwwUDKbjVD749WgET37avpMd3aw0j4iq894kw4Va1RTU24KAM5Mpcaq9ZhrLaRL9pj8Ph
0uRN0M337pgFj2fcWu2wH/d5LlBpxZ+0OYN4SrfIo4sTgt9c20gZWGiqHtlxiuqlBwtipCIw+jVB
2ATn6V0TbyAKdH8epRW8vNfuQOaAB/H45x3hLYLWu/0M+ukCCbg2qVAJBpouDExgr0CtTogwcNFP
w7+0+Id0FnkqCnY1XKaLoB8mDCFpHxHG/8EyXxg99fE8WHmCC09jhpYykX/3ihdyLsTx5ksSd2de
HzrhM9OZKbZeSWRtwPnGjRVvOo/i1ql1ziWcT3e3/MzeorVkRpmTHc2J1UZ0aFL/Cc3W89lCoF4J
cnFl/dUg9K89fVCRcu5XXtCNGfaDylNnAGu0PQldUTzg9Ejh0oaYFESEeq9Exsff0v/LnJXr6D3I
tcbL9aBOy5qhnjUGPcSgy+W4/2GO9t6e8sSr3cJbwc1XmSGr4Zwo/r4ryckAygo/Z4/ShPhL+bYe
9Q+kV/Rr2apr7E/oXWIAVuHgS0OAlKG5qSTtY/d7Nt5ndbfWvYu3nFN4E/Fq+SJK3AkgeAXn5jBp
gg6ddRwYXsaZAfYfkCCP/5VPnVZJu0fmCk2EjWuKy+k0SOypcIkH5ytjQj58ls2y3FyDJbkF0I8e
DyMGPso5ZhgTD1TwLzLE7DLw+GFEQBe2nY/UK4KRZLqUDmhjlPvnjNwAcJU4g3eLQMI30QKrjo43
w+Uoqi+gSYWbjijuR7d/R9Pm/BLkMoSB8AsMaU+zj5QQmfaqHLFzYzlBnhpfRBwcuW8yZm3gntB/
4qyRqxnaKSSHkA6Ol7jWlBBUPe81+vUWBPAuOPZElPOOO4gvjxR2Ixir0kdqitaWQprvJIi8A4j4
tRxhxJt4W31v9FfSYB/PWFVn51+24zObKK6rvYE4YABk8ec8zfDIY6l/MkUsB2PykTuhH3+8Kqn8
ALfLHp7Q+NwGIEaEl1YJFrDThSXshv0JIMfdwdhbm4G+GC2XJWEaw4z/k5WVOVc7fks0sI4oNiN0
HWsdMl0HCsyNCYeEm825s9e8x4xhd2GFvTO0mgwZaRRzZEpt60FeBgPY8yLs82C4xNP4qdzeQfh0
2Zhi157j87sp2TBgT4RkY9WrYnLjhwG27RCRknEVvg0ElQaJdhm7WqPqBQSKoFkgUcFgr/MQ5eSm
VDQ+OFL+RBOfVeod9DCkBqHRtsCtEZNZ697lZn+rjHMXUxq5vKnvJRUd+I/2USWvRbZ4zuqeNkJF
UltqI6x2v3YEMEtupDSO+DF9n2laxGTqf1o0M1Txoz1zXSMRj+qRLN8H3QUSIcVQ8/QqsOUm02CL
dYE1JoOK3kbdJKGvqocsywLUJTvPUk3/ollqcC3k4Y8aLtrkNTwRF7oQ906XBNYucihXnOOPkGPJ
MjJhR2wgbGUUpyqUcuQ5k4Rlbb3cEg7fvELCD2Ir7aVxQaV3BWhoUOas3vfeWFEs/NHCpa/JctQz
GjjsYDRpbcLcLEw5NdmdZFG7aApCgA9eBVtyoUuL+MRcgNdSUhf7LYESmtls0UAa6RxXrO0oWkdJ
pdeYhcynA9Rk6hVJ2jjRNeXM7bgN2Buue/V8oYtWASyKYpLkzHcaI8p5aaB25kNwJeWHD7ISMx9T
HwnQHpf/gmBt2yaxfYPrA7qCdD8QHyjNjTcW9ZUlxdHb8uYRECQSx3JFafa9QnAdSunEp2m6cDdJ
H5AuNFuCf0Hk5sXXiDpFFhgWkFuv43qEFGcGphr1UgtiWvuXQLRMB6m7J17Kps7ecu/eIsxvDgvz
zh7yo4iiYjyqeyRI8KILRs1rW2LcmJ5lmjY+TZ6EiHAZZ7N/h0TyhG7iHHHw+qBSi8FasjDZvnim
3s1A78uCPOtk5cN8Mz6kL4Wn9UERI6G6OKH+2gb4TmC9jDHUEtzcrt+7bi6Qz1msC/1qCxgasKmO
uXPJCFCLkJo8FTrFCYTFfSUKVisR9npLkpN2KW3uPYhWhbT8mtTGUqOjTwv5dUTzMWHR0LoE18ud
2TiDm1Q6+r5XpO3BJhjmDgUFTlAzyJjMWYMvg+dlGrkYcGTf9YWkYacYwubzy4fDVTdJHOHSRj11
RNqABwjts4IGid4rmDX0rdwVN5fNahMQmzO0B0HJiNth/YqSbHce0rNVTpPVKCGmVq0yRDo7Pi04
Qlvqjy5dqlpi6/iLOgDymky9KwKJBr5oAVZvmo59uH7SsBQP7W9IXaV5Jeu1cBNwrRtaut1wNaU6
CRvQdWKPaUze3nRTApFTYj9ocoOvhut8qxfLnJclmI2kIelQHmDIYxRpjZbR7/wnKCmoK9hX8M40
9Z0DJ3iRsY8WgDQoVgWpRvc1zaHfMHH19o+reWiTSDokLej7/PHQh6nom24Dr+dgpIiSr9rutKkt
24y0Rlliv8nafnRXNMu3bUhmC9CuveXdi42xsP5F9f2cnXdEnLH33FPJDU0PfdgvJfUulAGS5tV7
yTFvd5i3WtBZgItBZyKZVSdRxByi7t2RK45j9AyXrjhPqreJcFJP0ZXGF0UKnFjvuEUlsmMznfFt
24V7CPI7U6z6P0D9EO8BWOUKWp1F55qxqqUOytgdzF0YYOmF81ecGiaXXCGW5wG1yHSk3av5xRmt
+vToSxe/TGRrT/nOG1+nVMyn1IXplGue4JDuP4DJKYLfzUJtkGDfDRIoAQQFWOS36cMNiiooCkog
/Zjsv/foCeFF2CUkYrBYP8rjXJJFQES4/Dzpn+Ua+1hTw/pF2m9AGZYam9eRRht/tQXMVEErL2IH
pjhsuxrgSJGW3Bm8LKllMqa1biZ8Mq8Tuo8wUbXKR8GG/K8FZ8B53eQz04EOKWyzYptiC/yISJf3
8MQUxVn75qzlSH6RNAwd1cox2t5rJlBJ0s47tgA9LcOJTdHP/mQMIo6U58UEmfBEu7FijRHBazYA
9uIlBzpiFaLg2FTAftd3fFs/sLVGuAZM8M67w3urNo+dGsdZGwqwr1VoQY/6lmWrGQtc1JlSHvvw
+vtUW1Ut8fQbnwXnxLUsF33lF26boEt4NNLKHvWydiVQXiy0/fYTREP6L/zXNm/PmW7L00OED6vr
mW01uKdQ2iZfHvto8Ed/6XSGLKJrYj2eRpXthYRnJKF6Dwvzmt1351jDBo6RGkqhHl/MQh7DYxvG
4j+B/sPK0WGULPSuiTGkwCgyQ06nV9Y5mBENSZEs2vPw05SQMOSOlaBYyMjKHN/AU/L3TKAPKDMo
fOtPC+ybilRvOCO32D4Dvrb7WjjCdZKUHIj4c9+ynXMht/zkY4bXw2uAx2LY5FxYYM23oqX7jZBC
5l+6al755gHYJXm6rBPVbZkB4CSF54K5+alN6VH7AszDWsIOfxFueZsQOtcRMZ4xcehJ4mE+H4//
cDpFhFatVMg6mlA/yGnnIDvDGTmOY1y2ZfXTwkjg+SwXH7oHcbf69VBTeV7XiqH6wFPCO/Yhe+/m
uOZW2sT+wpHPA/920ZrsyM07A2YkHHNFwvRxL8qUODg4jJXF6QoiSoxHRdxzMYeKAFAkJp/RV8Uw
i/zxwFzResZ3u5oIPLkNVsOAKzJcvnmUUekonhNjp45fnfq6Ns1/uduc0tId6JZVdQ6Z+3g8/MrZ
bZgb8xBYSQGyzMMqf68Ntg438hitDWMekc/zXCe4O536p7xqNAEpZxdL10KB9pAt+3jFyfrEq32w
GnsnYXUU3t0wndTjlxcnAh2ech9D4B7vBBa7S9SR3uP3jRNGj3G4xygoZ/JIlKhXTevkuUaxKwpZ
5GMls+w+riWTQeqQplAI7/+TtUOtT4+ApwAzED3sgSBcLJHrPGKR408GM1DKV+zv3po/rJaSCTTY
S5GrM90k6vbZWaO04X3QJFq8x8svTRNX6qgc7tAfVN5hwXDAOQVUZF2Xj+6+UHpCkDuW7Sl742Ve
7rGt2U5KHhgvVJcjshNmX2UmnSS4uXEkmZj4pFbDsMDKOUErwcnhxJg+F0xp/ZB7sZ+eI0WUZK2U
BvvihvC+yjijfhyCtOMaUWigeONNuF5TVaiylYHM0jm5Ri7+JG9LC4k5Fkkb5cGPmMCQTDu2Yc1m
KT1WqIcwi+a6rxUDny8Q3le1sQTtSSfm4eszI21D7Ia49qBcLDR9pkcU42l83zePHROfNl5NIMG0
py1j17m+oWEEAOum2OZZ4BsanI0q8K0L9l6RxzBJlH3s4Ckmp4cgmNL2wF3tim/6X0XGmnl5cSHu
k8TzkjdnlwqFo+qFm2o5emDVxJh7dLbyXCAzeJxxVwnhEmJedUdTpvLvVoPsoYm2tLZUNytROYkj
1k90Y6V5xEU/vxBndfs9oK9+VSlit63ic0lRLs8ITRezuXd04ME6FcbZ3YXaaULXFFprydmtsRCe
OGl9UPXsqOYYXB3CKXYinQwCmBdmhRpMhqGI4HKkA0xTVnE/lfqHO3PcCAdd6RgsCLLrdlr0Llut
HJkhmNvRsvHiyaSN+u+Fgwi+aSi5aZh66osfWISzPq/STX+OsKeXmUXeQkk6Cszb3KJ4j+XtSZSY
qDnlCtVmQgFqSZvyD/2YOqAGtHFhHYVx2DLTqqi4nokJfg71CPkxt4ZOn15NhujLR6uMfDWb+9vc
oh3Vd+jubiUvlu6da2UbfHxmf8iv98ICGejwU0A6FJN7SGWk4tHZwzRXpcCxmOcZKCpTepSosbEz
+h3pgDc+itkRmSa8qqx8UsfSv4qeE5yuqIlMLAP62lJ7oMLAGQZIu/nmsgszhZJiB9nwn5vmsp3P
6hHUKd9TJpO44vOrhmoa8tp3jq825iuhSjxXLV9kJZBxR50T7e+Qr1qY8dDftmMlYeSq1ahPlPJt
Roa3WjU0i6zklvLzpHJ3jgDQ/G/rUsMpSZYtJ8o5vvxaAaHOJdH9+U5Wz91/JmwovkDegIy7+GXF
yiQQblkUjFECw2xi7Tmwr8I6e8+2Vsj3aHl9B3nyw42mQor8buCjq5FiM+y8Dr4fPHTO0bQkhqbw
k/V6dMLfS4ZmsfN6VSYmXCF4of67s4Vpkjplad2PRa47NeMV2WdKcp5bGMSgg8EHjwjOY51obUH7
5Za0IUl9YrkrItVHmzTjDzvgTGA888lBZnrpuL39dwUwfkDKBR+19dBU3Jx9Ub8qHrHUfXfWSFRA
e+Y1nw8WZRhVgyDgj+dip38601vV3gRQqUPvvPRnJWutuSSYZjThX9Nu6PyqUOAkKisBaG1hOf2j
ednk2zq3dd1afeNa+Ciec6/IeWDbowdS6a1PTzE6q9KKqiXE+yw2ksCjcrWB0bQmYnRMWjt0uVuY
iZTaVJlt2K6hINaNSaF0wAlXY2iLKODqfJCKbCki8/Kkx5WUbAYKfgVMOzxLWtlVyMdZTRehuxsw
KVgDa3EEMPrB1hk3CV8QnsOn3qhUitn8nxj4qZMP2TJi4R1vHWkIweg4nwAyrUJDgXgXOJrfedie
WSTHuYT1dplr+6WTn5hNrIRPWPRodQ9Q1HTFV0SM+EJ5TwYtRbh1XO7HQxmlYReanlx6qAnQJSKP
rJggxMGEt2G3Hkb+uhK4GCrxMhq1QtHejdoPIn3OFt7jsmfbWlqYzxuF59UvbPCGz2wVyhsQ61f9
GmPmyYtAXq52siVx95J1LFIoLo8SckusvmKzzTZ55QIvElIclU+HFpUDGT42lGQXVNak7CEv0KHQ
4MWjIIKaeqV0GJEqVhrrFm7EzwUlM1LP078eCfykVOql4z5h8JFSQznFMI28kjnnmdQPbUy0PXxN
U4jFig+OiHTsC/PMyBt5H4D+z2Pt30O/ldocxugy1a+9eEg3YtMmNu37fMH4Y4dSwGbccVVlde/n
z0Kj/13OYkKKydK6BiOkUeAhct/41CilhiWrvj911h4Hx9dzwnVrelHl+iZuyl6VOhbIJXaHq1CE
TqTw5giq97qVc1Ca/RC0gCvspc6x9YsMduDyxf6VEGOY8a50/G7CZAMeWvub7oD/FEsy3XIwdE4O
gz2HODTH+G8FtrOYCaTMmm5cyJWmZ8JyiKGxEwzzSjy0N1YhZl703ZI2Z1Wj/CC0OPj8bDlum6is
XDAbzbO7AexIVrvEIra27q2uVoKdZUQOB6LRCISf/Ev3Oco88Pinw8BxlaDq5P1pUUiwILcFVL1L
cV96ll8u5MXaX50Bt+BX32SlKqy7Rfgl/xWo1MvISYxEqctR5vS0oh6MseJ9tUesluwRR70s+lt0
nZjcWE/XiArUzhhH22ZMmWOIgwouLo2bzY+62+vNm2CRLmAEAfB0CbLKzenWg7E0bmfntfi3GRZU
BlDt3eoPSNbhtVvZvAiZQkCLZ9MDltKFBtHBf4uBEjoRWiSKM9vSGMHC6wDHDEDF6fwMCPGcRcEK
96pGwdhkTFPj9fkbjopBCpCYc8j9+50agsbheuGCAI0PuzUP05ltNUrh3HCemQQ3JWmfCwV6wKet
TitEcx3XsidjgqV/sPKKMOSLo/PTEZIpUGImIH5eMVs0d0xoF4u8Whe9vGwF7MHO42iCpKBG6wIQ
2A4Bd3Mv6rNYo7JW3E55VdGc3BJ7c2uiLvS8LsM1ssr59JhRXWI6khRcGhdMtk9t1YBb69kTBll+
LtEp44WF/H1DrJiWIDftfti1vwKjVqwnAwghkYVK257PvGxP3dEjcJVIcr/fShGWfg0mq7byY0mu
WhMTxbNn4QBqYTrfz4QPaDky/vTXs6g5khJtRZTKnE0FjuJC/iZdnvu5oZq37v1CtXsnk1vhfnAX
DTESGwWPPOrQODP45SeBI81eCerE+OY6F8ell1X/6TkEsDOPheojJmlppITJTGYcvanzkE87MfS4
ZlMNTNpqJOn5cWu5VbqFnEA7B77kkS+IgSPKc/cfRgLpytmZgcyaKzRuKmJHqCBJUzXOIZeFnqf5
HduhYq8KUwUTNTBWyPIHhle88XNcdJTykr4TL/P9dkAZ+CHRMX2DWj+BFzblTELNPNYtXbefmfkE
dSXVVNxbkkZ4m4XgLuFuhb1OoQbZoub7g5b5QkvqwDY/s2xL3pOUofMpDfbXcbpDl7F1cWxVrJOI
DCt4NbIdYKRmIpdSMfOT1Cp5P4oYDAvNasraWVt4TZ6GFAwbFgWh+lRqSukZJ4Es+ja5KVOoYDd2
1K0t/I9JZ6svD8ZicvB9w4wFx4aiRwMSY1jU0VU6/GmD77NY9GYCanhA6fe3tbUa8os6QCW19N3o
8tFpEkpxxoPnNgvYwH7r6DO41sauMUKtC9MJ6S2BCx3rlh1VURya7SeXNtapRgSHA/4KmH5yHDQ+
MXkvrU3Rtk4MdyrWGOKZu8ympAFgDNFZeuTDgvgFQt7zR2NtQsTG84A9060EhsZbCQpn/eQ1OONY
2cg4byNbTzaNNqIOLKagET653TDO1VmmKQdrHhcoDjelpcxpL576WxBcUVbbtC7cBuVz++snvwES
bFVMOd+ja9uUeVeWDQCIIbDTycMI13ysL0niwBSEuFYOCno5MGlJaWWSp3tdrNFDPjWUWfVEzGPf
Xbooy1OJT9m3E7WFjbveMb1GdiB6KpRnTftgwakfWFbqScKVYc4RNQWHYl3fOPbl8m93TEwAzbPQ
26CWSac52Jq9vMW7qpkLLa/IgiZARqyJMQlUPTY6QMuWrgsHud4ugUeUI7FH5oXB5hVQbiQDNPbs
ZetW3nPxU6fgdYKZEq7J/fit2pH4swx2ezLXuZvYP6GAk0jl7hGYF2bQSUy6C1z6qQrG34k8X3v4
SGhnvYwg48CJCB9q2iC9KdyXIt6qxiyxBu6pOklG9kc/9wa/XVu6V1n/4O8GEd/3yQOOfSsL77Ih
4aJtxopfnkYzioiLjSPKKmEOBiR8/9bf6ZmYLTmr+bR14lGmM6pdN4HDhp03ZWU22g9mIAVdcSMx
yLahkuduf3gXnravldNY7w4STVDvlEWowJKpcwJj28gB0g0TLfMCUZC+SQjN18Snyg9Qn/vkr/3C
rGHK1slNel8yyqc8Gqvg6ADMIc28zmOfSwog/lnbegxNtHJSX5iI+E6yUEypWaefYTtL+URXmqX6
mQYqpqX65thFcuM0JZqTXn6crxf55U2LXUhQO4q/WTI3x76KHL2yjgac/J0HKEvtgAl90KjpCiH7
AgufsvIPgRwg8eB646kFWjrz9ScpHIUkqO6+cR+wei0R5VNVuFEIsy0i+aX0Ly8uLHCM9Q3UotgF
GHYHlfuP/9r0aN8SyJ5P81+m2Um6GvtvfyrWNfyCLuiwnW22D2ObQf31FnsCH/aXRT/jvQAmwVEM
HskjCjSWKjYTmfxUbwutzhdK0hyj+oOX4D775IF2+3kT5G7nAwcQX2wOcTNR8NLlOadkIvghlajM
4DclL+eFSvuu278mo0dVknZpkufDDnjx9abMPlw2OmGy3aJ58kBk9AAb/xdpcCwjGylAzbsXop8U
/MQB3/SLqPZt2NRoJfW5Rl9k9u4dp3LDWNG6EKovEz60mIhBxcd49fFdqB+Y7CxfBxjEus/KyMbV
H8mxdv0rynvmT7OVUVdjQa53FrBCkr17ILv3S+e9vTQTHH+p+DTWM+WtqJrqmvy4G97X5DKD16D0
vLgnJQBE6D9hLnxbS8cVZioBTSjr+6blu/24Qny3t7uPhwxQQLQvYQQF41RnFNb5shfiodIDV8f+
FdHPGj3HcalPc7J8r+ITRnFtT+axwNTV/OTEfOfPE4kvrKrqY3089LF0VTGYyW+rNMANw13BwUEo
mqmBIN7tFDkLinZjhTSSKyRZygrqYWO2nsK7QA1E9i9pRwfIoR1ypLj1GNO2dvAdU9x13vRWfnRk
MDGsmzqnGBzB+IUrOXE3H35xyo+8gQV+YiwkGulNVSy/Yb5Z33V/KKGa5oplyJW0TouDFLBDA2kv
pesBJTZZ0ET85/oGaZHy6W8O76UIu9wRZhWvrPhfFSuaQSbUu48imf9/w7zqy73s5FREyRWsRYPD
Nxt/2UdddzRefbwlfKAd2hqleGfChsB4gxfOLXuTy7pblLFiQ1/etvJw/3yaNwIgyV7cLWr3p0JP
jH15cFs4VWdAN0GPgPh655vNtDy9Z1akuOILp1Bi2SeNUtPBN3KPiSLeZHRhZEEBis0AvdWt9PkM
pUMoKCHtCkcPOef5F7YMS/5OQC7Yuxh2P66C0KsXxMsFMnZHX/Q146opv/sY17iUjd/jCnIsxLaH
SjNfbzPnKQvV79Cft5vvNgAy1vEhyQPi5L7h/E4NcknA+LLyS+lKl/FD0DSNBpgYpWQQs6ZUkOhP
sNFZb7mef0LnotRblAIwsxUvTxa7xVoT8E7NweC1FbUsrBloB94Y/pxAKAci85EC0oZml+VnLXuw
kjTCs+ynP+cELCTnOiNK3Q3jvVRzmiX9xyLsG5sGL3lkaCJPamWJ8AaJ8AetkuBRY7hiudFGuIJ/
AmYub2oNmi41y54KU17VNLHstSH0h2YMDCrRJbMZFu+2JiFbT5pFW5G5iYgkZCiQje3W0rFi8dkD
BdM5VhMw+Atb08nDTbl1GhUQaBbO/xMp5FeGoAY0nJYVyavwDtbA3Gdv1GyoqrC22b0ztgjhKt3u
ptRAgLWvqX+/W3cUBxfd9DFJuMkvO8wnWwwwnwFQP2rKz51ydVn4YrIWaGKsIbqmtq6YT//HxG1i
RHiczmHp4+EbXj9Tj0EcUpBRd96sGigjZSZOLWFAASryx7yQGw1KyVbkVd6PsCcHuihECAF6FdZQ
F8Stg4sn2YzknV5QQk3oJOMXo5T1R0m8+uEEbvcAuJLgh90Kqb3Jw3Z28axTMnXb7dE9RVrK6qjN
MwZrWgu0c7erg6YtFY40XdZa9NYv5BXBqzXj2SO4OPIfj1kz3oIxy3vIYAOfpLaR2EiyK0/9aDA3
/eWPDe3oNKMy0jq0J0XoNOJDZf67RTBzxgX8aEewWJUAkmh3mVxxsSm/EdVVbn4F7OJyDA/QicvR
QAji7P1RU5nVRCTOkJRwvN29MJ22xhGGqm5IuerGI94fqbp+AvsHSv699xjWAXdr2DgIFgvNQ5AA
BXYl4GgdeSzykIpZq+vkFGjtoz2HMuDUurUmclSCsZnc50s3/FxwGOF27xJpUduPyokLXkmYCOnA
DovVSzrTd/Zkbt1+4u4kkgAK3MCk4sgll5K19vtw6ao53O6WLV8d3L9GEeRxVezFT6qMfxDglOsi
yHa7loOrYiLI5UPAp46V5xDYotDpaakHnxpPvrb1Gw6S83xuP2lXSFmqF9l34GNqhdeFq+vMhaBl
vrhnC0hO6Y+H2X5T7jS0ROwhrka2QalVS7oA+a3Fosy4xVsJ8k/abSPoRjQ3Jx0gEUSbJmPlXKoJ
BK0Bmr/kCi2p100SSVLaIpXWkUYkyKEy+zyYmW6SwEcxJc9FnxRc0KvU7FFYIbA3IczkSlpuqYMD
n4s34mlUHfp75V5Y9Sb9LgxMxe+AhhDWvWujEKptQui0dvQox53CL9o4V0tHSY3w+eNUjms8r8IJ
u5TthKi+WuVrL0WWeuCGodswLgpqzS8o9Ro46sT38yGC5b5SXi0vx39KXkZ/037Rp8iYBMiW6gv4
rCBRPJi+Txk/V8i15Z7AZkMlJxEEqu2d1kIhq7zXW79CE8SK+GS9zPGxDV6IZLwo2IbXZEV3gWBm
gm7LVX26dNt38HYohPhv4jvppjUY3b6MxOCYyHwwY5WcJJzMDefO649gspAS5JOR6+N/8a5kr4WH
sJ/PUaVd/4Rxb7RuoNKF+cFTsskSr/rn4s6xMHOho8gaFuQeB9MwoyS+NI2PGYwm1VXE31ikZfjW
lWmkB8hNVqUbY81gQzGgA4rPp7JjXsZEDKWqFJo8glPap5S+m+i5FUWJtr8oCEI/0aoty2XK7MfQ
8/EYyad8fIePbmoYFXif52vPISWNzGJH7hgL5Kg7d+GahpEp6eId2XPzHW+W8j+VHKhk056U/OmK
ExW0laxErEdmkD65jIwc/C3EyQZrOz5/cbzIYKMmovPOEWgi99VnY7eTFl90n0sP4cfx8iwD2msw
Xjq1N8qs76/PVqe8ldveO9LcwCN1kvumlcMlPS/pthYEb2J/rWg1TBgu6s8+CaD+BkxPMExMrLnj
Wr94DorgFlALalS48ToVUzrKBvc/i8CVPNkmBorKI7mFp2qF7nx2v87DMzfY0qHlP2v8T/VFPSUb
L/ltobIhhMNrMz8MykXK8dZGbK0J0CGihzqJWd0K029awr2dYxhECHD64VGElqDqvhHrgHAY1Xnd
zLO2jbmuS9pp+5iUrNAvfu6hHRi/5AhHzWRtShqrUhCojpamekZCBthrMD5qb9yY/ggZvKXUrMt6
Xeu8Xe+uPB1lF3qmzTlbLknQtk2x6XRtDvoHH8c0gLKebS6+JXdfYCzsErHBOWISQrHruG1EZ+TT
NliyQGV4yHFouN+wXDNRStEnjbX5HKJILn61M5beIUd8EXVMvbkoh9Ea8p4AfSL0d6FwnIkBADwz
sZP4Z46VOeiTiTP+kyJU5WUYrDYkeDwxckxhJ0vn/MRTeRBfy+eZBXoXP5ptI9+lLSNnfcHKXBg/
XmOr7YoHz5TaXuq5K2Fq/NNDvrn1RRM8uvXz+Xe2nSX2fxCrkjpuyDtqVE4DjFC6/A6GpQID3gas
Dmd7jTvxfYW+KRZiI2I8X5bJNLIFoxBLak5Glazdn3hAt2kmG7U37c/slFejvrXo00cDkQ+lm61N
UpD0vsCVHk8BVnsG1F65d4nyOuWiYsjJQxJfFHl3qGbuiA9HVwzNLJz92Wf24IOKzhSA63uRHKrj
4ebZJjNNT0gl2yJXrAA+0lfQ34ix2UwKX58Sw/HLjjqWU5leJMPC6oM3AsHbnlTEK7F7EYYOZ4Kh
roTrP1T9wtN0YeATXDoDeSdO+FiUzF96ThJ6BANMBjFiNbLs+L8qbcI8wEuPjsOjROiz3RWpF3GK
l6+H7vxLaFfaQJeSAudHqRIvg3QEl6gvXqoJ/z/cxb6RP70OJYrCSMp/xavojcuKrcvvsj1mxg91
Za8FhH9hgj8mMnSMwiD/WQqZoRNv9IOhnlfpU+7seSJLWQQLW8ZYhM4Ylcb9hTeKUep/u0ndxNDx
Q32pcCiwGdmRxiWETtZz94pM0nKPimzjhJUqsdJ4auqghWcF1wrMqEu3PgrNrR42NMn4KfihJ49L
V5Y02RYxN2FhIzKuZ/SYVPlDsZqDnLlrCFZ2nv69x/T3ArC16/QYc1Y6JYT6tBgLCh5YbeIjCBYz
aZmlel9EQ4i+5dZFs2lx5g3XzY2Qr2gaLEsYWyGcvfMDOvrezuXD7a+j2bD+1UpG6MFBaYH+MYxL
GLwfz3R5acmACsij3TSMZMh0RGV6ez+GEgZLsMGTaFC7ZLzElPi7R6P8A+W3tSSAq3qR3Gk/bb8r
Inv6RT3GEkz6Q7Im+cP6mSvAdpQTf4tCOLhleIJ+8343xEWM5ALkbrFDg7j97RsPy9GQnsPbjAc1
GhUhOm/sn+mX4nF9JQM0kK9tos5alDVcr3XsiDV6yDEXeyWcH1vKwZSpTDu6b66sjP3GCeVbE2iH
2xK9IXVZmE8k9MLU4C8WNaqJ8MCt/8WfnjSbqwejiI9TcwwLWZZ1+AE3k3EtLNnEr/78JHqqHOXR
cNgm3leEa+6/8Hiu18LsKLH8U6rEuQvuzm77Tlr2qeoI87GcqKiN1M7DV5qkak2Q6fvOio22u4ta
A2XFQnNadkZmeH1u43ujuxf9M9snuPKqAytll+J8uBigDPoLuAtNNMk6IHDeXTNK348+dis2n/g5
G3hrUultzv5DO+yU+qekOtKmrsGURJD+iLR59fKfmLhSJYdKUcAvmfKbErTFmj4gAOQXVRSRwOgE
ipkkNVv6o8vrOT1iY/KKslTG6fN4LzptBK7Vaw9AnvG5+S4GXlmGVKRn2zZnxMKGWeq9MWR4iP8o
py4W8vucYnhwcmYxHV4DjToiB+Aihw4c2kHE8IDQCaj+zyneIXvB2d4wZwoASlk2PQLiohJi1t5e
GiheaK7Q91nZv7RoqujoVWMTUyO1hQjniyXcROuHB2aUIzTbbDYYk/2Ll1d+d99KWw9BmihB6zJv
8QoyslT6u2ilSOoLYd9cD+IVym9IRuAzpPKBMsyxtdgOxa6Ng7IDjGwX09OYbMfOPYNv59S2Z7bn
taOqfMis8TzjrpqKUkut3Y7s5HikkX+SNoY8VF8tkD3vkacnS2ZvruJQgD2t/Jy/dJYQn8UMducT
hLCAwYQUbeWpHi/a+5CMLSkGu/Nk4WwgHqNir9eFF/hPh9nwdrT82IeYLNWbuwil2xRPhRN1pRb2
ITvJgVp8eJ6w1VgU4UmaH+fNeAXmwpb+qSpXmYlMdVstG+wTBuP+LjR9ka23gN8xKhi47PEHqu+V
o68jQ7laIKzQLIMSJvlrW/EW9s01/RGEkSnPV+PT1z2HR155a+kJ095o9ru5Daz04iH9bvPQxrQr
ghetxbGLYp8qiYQZldLTAQd7GDHX+oovUcBtgxSZOV4sDXRx2LVeDbA2JzIG7erjRca0P3gmNNsJ
CDXumHm8qc/08JzONlcWxYtO95RcCUy4bem8289+ybz/26ovwYJAeyW7DgKYWNDch0bbANJ2ErUZ
UdOJSjAwPvrgPkzKM95s7eGRfvEKq1IUgFRAyFbE7E0C27uSOVWLQe4sRQtSY5f8m6ksAcNMOSdM
9qIror+qBM94OiuL8y7bGJA6zBW3LVGNrrToIq2JLijZOnpuEhui502eT9BVl13pLf5w9wndlkx8
s+4ohQhK/EShs2/F1hYJp4gUM/TWmteQ3S+9PI4FrZPVl4LS8OWDCcnYmjzSeEeeNAQANMT1rBgH
gWPW90BW5wUYxJ6zIfWLrBENOdc26wXN9PwW0gkmaG286It6ncbv5MeCEt53IYfzWFCfeu+WSu8y
A70LZ3r2JxHt8tcVij80E69W1YJrwih+rVgi0/D6be4Gw9LKKDkmu758ShcBV0KF1wNO8EHMnGBj
Nh1crnTzJhThjmv1QewkQISxh/ujdvhBJ6MKc5QDAOSUwRrvbI20O8MTuA3f4/xTCpgoLqrx6SXP
dCuB9av496iiCjJirgAyN5T0ZYDwT5Ca2GZdZgIDrRFla1VPN6FdNyS7B1oWXBIdcjdpHjxySted
zTvFggcUv9ezn21dkto6o41Q9F6ZEnUXPmMu0CwHhaI+IsC/WX4Hj41zwYI5+nu/uQcDRGdV4KsE
NjexHk0C+hKTltjTXd5DyY7db2GzOFUmCy3o+W2G3/+nzeg+1V4UnVNTp34LO5+HCrqop3sz5GW/
1LDXq1bovXFjfLa7gO6PGrbzVRHKRqwLf5jfVK+e6WA9vC0Ph1kI4Lo0ZJNAS/Xae0P+CsviSDsz
7pmCgLzhrRE8i5wFEQ++AX7ZNsKtiol/H7faGqo/VEBC2Ujf37WIhCbg4k+yqeEdwsvW8l74x/uv
nmVnR9+SXcxOf77ikUFPgH3/5C6p/lIEOGT+yix2e76hrJJxwqTcddUisceyazJspunLqPtgWf4G
S58yWCVEWzYMeR8koDSiY7X7fiKFaHkod6hn/OYOUpj9FLD4P6nvclpQ2VNdSgP+WUg17NWy8g/b
6+4nHrMyE34B8wVF16jUZg1x9r1A5puDvVblb5Q4/2RvXnJ3OoWHTWrEj4jImljFcp/NLfDLRyAe
64e7/TCjI4corE9M9DPkxgugiZxuXbMjFxHt6Ay0Tx82MlQ2GsdPWhsMVjkx+r/Iwh6h1YIAy7Bg
lVflANOZ7k68eIckeT1A7klhe/T6iEPi0mowNlPcqXGJLnybRMM9RwfcfCYHYzc0iGlp6jczKfhH
Ozu5Xh2KeK9fJ8zS1lzMmE5ZOBmmqVQJKLmP/KKhSj4Sps8uAncUdc/H1nT3eY4pV4bv9Vmpw294
gKR2Sjo2RuWZFaPEGdbVJfq1LqnW1KDsa0uscUrhQ7voctTxY51DzIGjXmVmsANvaA2VdaPL0EDl
PKAbDxNMnk82PF78ORE5yZ8VBsgEApmdw6FSTFNObEkcQLzU3IAjDMve8mRuMXFSe1tjZYNC3l+A
w4tJqyaZ0hUlbb8XUAk5wsxR+CGI+2BiExM277RO8dUBnL6Dqu93CPew9hfc8I/Wwp7hMjIIrmpB
YmdBBm1uHLvhlL7VnaaGWwdoAGqBtl/ZcB2Dly71k5VOccVoujs/yRRnF8ksGaECsJhIm3NsLsuj
v82Z+5Kd1OvqiaFcPO5zLo9rOQU07M51/iOHPjnkOJkdQgePA5eEzSQh6rU1Bm1/jxoBlD8sKQgW
OcVlRfy32r+3A34I74qsbxkKGet2s6QqYH0K1upbcn++O/sm8KrLFG5Y61h8fRYlJU3TAtiRZq3I
XAv5NZo116i0ppOc3gLkwsl5yghAFc9AFEa+W13hmz4/Ey0pneagWBqoCgMHb7kQAzVkdHMWFtCW
6rwifhvzX49HhHuTfWJC+0X83Bwuhz9LCvpFNoxA0VOeC3ePoP2tVHHEH3ptHcmj0XTkCoaJ5s/x
JY1+SwNXJRHS8N51DpJV7Rv7GOc+qSrbQhAMkLsWSUUubP6UWQwGwDqMCjcpUuUVZhK+KBANT/Aj
k30mhdy4ihDjDzgaCOlPrPhnspvrV+5hjDazhig0GGbLtqqE3tTDwz7BESFbReBlvlaxqplUds77
tQeiKTUz+5PxXGfc3OQXg0lRG60+zNSINy3K4JyrTbnr9EDu5N6s68JCWVSg1BhIEqQ4V5UVrbpz
G2sf+4qgWZQohtKhngNcFwGebAthPtLzNv+S0Z5xwq5VTa6RNV1fBWKEOThyZEuwzOxq7l4LTmik
opupW3zcymGu+1giDb8lkn/zNQp9lAmAe7ruduXyRZz2h5L7J18RFP+FNY1J6i+cZi1EQe19+D4/
1k8tpUZCTJDwO0YnkhQaQr3v7/h/uuTnlVhWnUbfKk9fBWoWV9twJKBdQVbm0SRp58o9DlyJ7gSq
nyB56qmJLK5kz692BFecd3eMdfGe/xYE8j0/dJUEmZY61J2PGEjuW4SitaQg68mKMc0bZu1vBqq+
tEyBZelAnnPIs/Q2QRNCrLyjpNv0Q11I8UjJcNgST2tHx4NeYIg37iE/zCvA6kMFlbIW46tBEgYT
1tZDlGsKDb5yTx4y7D4oylAvPooEhkxhPuMowfHl/lYdqq8K6xXpYQ0sruOggvhVcJaYcN5OSTWV
A8zmqDgYDuo++3QcozZe6HAjWPpZzO1aeyRJHEugjaMeTxOs89dzZlG14Uy3zKONfNn6EoKZi5S9
YxrXbjnxD6uYwkGqdxs1lFabAQl7+kkzQtxReYL4Gv/qy9XI0TBN5BSydOymqx5moMHWKnbRVlqm
MoaJSeOp+RpJ2QQzMj0uH/+nTkDURrdLUXQv+IxWNrkFyUkRQCrJgybvMJ688plDcpCJIGdY+slZ
zigoaaWc9J0PAY2jkcktNJQ2Zk1mnqcExz2+LnBogp6i1cPOo4UnLZ/95WNni/VJK9f0SWKGcPka
aip4aCJvoyyl7CP84JV2iQmtoo6t1wVVKcn9mr9fGp724Yvh0TQqD/GpDJEoPEtaIGSUGve84U7p
3udLENLCHPUHvfW8LOC4gPpJufJaA9DfI4yC4GI/K5vCSkiqALKhB5JPRwNM/w8DXBjEcs6O+Lfl
LzA85BX/PSocvYNqg2QG1PTEd0npXLkL07/Y43YNulUqqAvsdglR9Ch+5QLocu5Aqh3/zqQKGa8l
rH4yQZaCCiD20Djil/+jtbGbgICY4ieCG4w5YSc1skn9l8hakoWHwyRNJidt+oCLtPcUykkR1BW8
Xy+YghVk7+cPETe9UmCrD8j/GuP11kXXyAFSGo7zFYcrZFjPLvb5REcYlh98LDeGFTcqPYTRy4Km
KPGPaOTEKyK0+0foZeqKFkgfrNnrO6gYoc0PZP87a9k3IDyUkRztSLeDXEYFmwiAoC8qoxXcswce
M5FDVMOFTsdV+TSM5WGH44Nv9i9MZF3sgUywPr1qDSnAA+kxNjvXLJsfhnHFgUb7T6Ul85rtkxUR
YsA5z9S4lhG7CRMFmYVFvMaok5q3N3uB44i3GoumCpeMrtZEblQNkeYyQ+I4XuU+vtdPWAM07b5B
a26UZLlkC/VZXdIYcEgoq6rNACIYwU9sBB5NubIDrrVmG8b7JXT8Yv3JG3g6RTrVBx2gDc89N+sJ
hwhvt/1OV4I5c2rlDpnctv1eNGboH2T1496EBhUBOF5PkEjJ/omF+hrbepQsgp8D+RCSv/fDqDrM
rKbY+d9QB+oR4WsUtlMEiTnIDQXKOc5xIP+gxbEhSqgl12pg4SdNrEpPen1nvpnCBihGUyOxSkGv
at0veQPkE9jEzOyPBOw4IFpyCug1jCusLqucmofwVFbiN79KvmaAQzVn3pfK1BGkpZHD4YpX870g
egOn5JMHO0hfawM56zKiizV435DmDBUz2u03t1GHxD54GecAt+EhSXexSX2pu6HKe1rC3vP3iHit
LwkqqUMUeI2tisyDiGU9qqnV5PYXMsqRFbB6XjYr6tFfgEpJ+EalbeZmBlC1oaKdJ9GKTdkz7GzW
q/uo6VSln5PJgWUdyEU84fnM4R52xwosug6w0Yax9aCEXs1HcnslqWhkzkJNKKhqHh0TwIeqY2Z8
fNNhc549Jt3ArQIUuD9bSKCsbWqtq3kGu63de5WQUx5AKnjRXtdH1spkldes3GBxHN+58kr5iq1d
veDDrqR7aAkukFhA6o/dJrxAEObfT7HeJ57QsLUN0C1iuZn0XtqwaO4tJQi/C/2oNUsr3tiTuiRj
Q1SpLIkyQRPlQ5mkRGM+dhBvyJiIrYP0KSkFO6gf14PajAPeAX6I5OekobT03SQtWAn9FQA5Tl/z
TtxZoocdznhoaUqkldjPr5F9AsiRk9X9s5O6ri5d+obEAxWlK+Kqkf2IY7lFBbxmj6fI2BuFvL0M
5toOIsViOxdI0z/tX8A5TBd2+PJxfPzgrQVIM8Y3mnLGuNb84D0LsgXw3zgstj6TMFc+iHOPgCqG
mYihCUz+FqPb67LkPvvpEZysUDLFoHMfDft+1vG5XDz1SuZH7ZGX0UEp4Xh3WDSbzy7Hp/fc9Qow
XCMsylxiOlJv34ewMfT6UTDkQzeMij0oVpC4r9dSlnE95gohnAzZ76MK8xdALHve64IDZT//TE4R
pWUsnzQ4CY51JW+Uaat0kJfBryKwdkvoBv2SmWWEZ12GOG5LhRmI+YtYDkoD4vAKbi5vDC4uGb9R
DQza+ldr58HN52fA4THb1wILtotV+v6OKkm8EuK/DU9h+t/1FTjmq1ml5z1K6rDuS56Vqg1BsgRs
IFYwKxAY+rZLzTPu8MIuY172qE+5xmmg3iEfgO/wWjhSY2+nyrXHUOrawaANcBxB/NYddE/veqMF
QK/JUFO0w+GnTHHQv4uNwdj+fPPT53oIBZlaFDelcmCZN4N9nURdrHjK5KmvEkRx0kh8iJqJh4ev
QKRBt1OrIdPrlarKcKi+3+IIElCSw81uxMmqyzRipXzVUbUJnsdlqjD81NsmdqJ7oylo3YxsIUju
a+HO+coDFsPaBUfzBNCQDhkdk+zDO3WwdteMvdEvZbOxSdripuZQu4TlXGYK9fG1b0Wa91OBfbXF
/YA4rMSuuwLwl+TSCpm0B00ojoQDKNRvjx70Qx+b5eqjEIo86sM7hXzSCUiC+ZKw/jRw/4MgQrTt
tFlQw5RiVQZcaP5SV7aw6z+lNPTL5JwM3vgI0zaMgw/Nin7SH96RRmytfv0AJSuxKpY+mjRa/Cpx
wwwWCgmJtQP+KAh5knWgsPGN4nCumgqnvVFo4J+V1zgzYFyO1a6c0R+Zbfdf58Q+5UXApNcbUplw
LnWQU7967tlqyhDfgVsGo8PpPpiifr0wBTCh4Ts6f7I50hNdoT9wc3ziAWoT+7duKgDuO9ut396g
SXJ8cMzGmXZYu3uvDNnHfvoHFU4xyoQtCAfh2V8J8u5VdCT5f+oitirf1B1vNbOSrKRUAqk0F2K+
X/ls9w0hoHFv8igI16UXZINhrfNQJ1qTOzpjEe5PxnG8WRIovecvgHOFf5dzepk5uUkUGFdL6L6Y
l6V9Faq3UbINmNKZTe6d9zTAfbbDCNtP3KnOtZ63a1Y83EtpBTXYt3vQbIm1LqDFrlt+ukd9DWVL
QL4Mg9nPIIPi7ziikAxzIaErcw0sIqrMg3URVP2isdgJw5cUqYzcxolL+z5Yr6mDg5IRNvzWFf/l
mDbaQl17edXsCBY7dH1QKhW8Mxtric/iTmuxm9EXfuJOUASoWdMJV8INpLLmwWo3D+jCRBdTW41j
Fi9MVmWHCasYlMhLkB2RJXIqX+ENOgkShVqahPUl50u7IRPH7Nh7MuX36z1p06xXakIM8nBpmynJ
9lEuPf0XkNJWFJ8TuNCC9TdU1G4sS5Fm2mY+4kmXmqavy9KKBOW9O2IqCDZ2pzGUD8RpgAzm3lNX
vAWHysHbSv/5ypQ01i394eDWnkSno/HCF6r6mPedx0f8mtQiO7bg+qRFSeMvblWX110JlYrZej+C
yAnxAvkiF1lGfsZZsykar9rBfDC4vWE42bOLd1SM6kR4V7L2fQPRfN3nLpkVdp3ft4i/eDJ1Ipws
cCtNaf94ovkDy/tSr71la6S7XCosoHExJjW8gGrJ+xnuV++29V+NPmV44EOo22DrxRHLwABP60Iq
ysbFM1vPREZNEOYW7EgtiTnK42QMLPFI1QVhWMWpG3LIu2ZwbXHKcaXrLizqPixZ5A57EC20ZfRy
Wtax2vCbiOVG80tYZhwNSIR/UoJqa4/xBrhaFZUaYABD2j2SCK3J2FyOZ9ugHX3+irKe1kvPfdGK
gIWuZi2HzgXwJS5KliguVwJu4DthLP7FOkzEYGfZbdNWCODmHulzP7pFnZNIuPf3OfyKQ3liPmgT
pF+Amb0HVxDv/oKg6pfs6qRPVLn1JP2G9vgcgRXhNBSmb6ZY0NvQmAzEfNF86yUHkqLHQK6Ccyy4
IlMlbXHqy488dS9Tsyl7dkEoOdXGDTX4yc6y2o4m5J1HU83uVYoVfPGd1TS/dYwda/kIfksvLLJ7
leLjVtHpAFf6vS6k3V7lY9oFnG4fCM1d4NuPODfOzgz+j/TFONnYPduNJrQIesuIwksvBlfUpwsg
ocUUsAI3Vf9s1ORLmuDNMEGE0N3BmfA3t7hEv/sI+50bWn/09ZLwohRsGod0ChEEv0LDkanPIeCd
ZsZ1WEl7LlJzU6JkU1g4xzu9qC6R12qMk4tpTBVA2xw5t+rYQ63pd0vuMzNnGUXeZ/eSODJU+5lb
DJlteBsjZ7XrWp2rjyUR69556k7FdFWM5KgIqFjfeeFIuAMWtIOiLZ26x2l4Xc9qRsj47b+9Jm2t
nQxtHnIx6K8ODBHPzO8lpgrURx5UQFjdK4GX7p0ePS3AxrDwqk3t/g2/XE9iBqltovPl/lae3ui4
6xUL8e6yx1kGqPP3eCS7FUb8lyboFffZfQNDCsMNKoU0FTE+MSDu/nWHLXEZOm17YIEqByhshIYf
qxL6s4zV9q6MXO1BryzJn6oObT/zAoJYCFgUMApTPDOnPfjC6tobY0oeqY5XdS694MnRsl5CTVkf
SNWyKwXpZzcoljwHHQOoFXerzX9gGyipBBE+avt3VUD5gysZVYOZt7h2dhzMi/GLKkbsxjl/xsjK
vzKHNxPX7jwdvdGnxrutxLbY1PNTJzIsa/9kEVY2ZFS4wtL/eLy5eg7clpyRLtW5bjwveXhFaiQX
dFkOW2K3BB8tE3JTAPOSmuJRS4JKwOgjzTX/nXmF45RI9s2bnChPYMCV7x9c9AlH+8xQOfBGGXdM
dY/0SgHk2sqVF9/EqdjVc8AwX7tIJFQLFnaHqFuSaEKhAV/JvvtquE1Wz1RmNzca9iHqvy0u10U5
ogJSkq2nROav0AE2PLkEK8xVDOB0f89mPVlNUxv0Gd3KpDqCTIuKmQzeC93PZ8CdMBsL4uYQoPGO
1ap6TMvmNn42bGuC7OoRmaAjF22eqi9ilFFff5Qn+q55E0i0s9A0vYV8YPdcX5F3DcL3A3gXO+Mg
zvCHzzu8zfffIwGOwui1DVqGwDR9VPuGrdnVhpBM97MfDxO8tb1rlbTw5IyDVojWxamx8x4AuE2o
W/9T2WH42U/z51ZOAYwB0PlwmEPhxeQWSakmgEzDrnmdy0V3OhZWaMlBjLIkKeY2i+AjvItEaPqI
YGrBeDuyoKSxuejGrXB1ariIg91vG/WflZAuJrMBN76y0K9C6k2UzosMfF0JLKTLUkVw2h6oE2em
rIFe7c0wIwgLxUpvX+a8hax4ZCRx6nDS2vjnlFSG5Qxzk7Gu1XjnO7WU93KhNkNo5AXJmL54WtDu
6TJQbELTFdBN4xeugImA1WeFz16Cwe7GmjAN4tLFclWeJ6cMhXmaltpQnxLnIZ40UAIufmDOQwoR
ARk+/tLKCtncF+Xekx3M3WLFOK99xQfLPj9Q0BgTl0hzBNcZ60YP8tnDlNUdIcqJkDLnvECgMg/p
hJzFP52qRKFfRANNRqQYEyz+27APg2jHocd4ATvnswwupvZvQHBZepvX5S2/z9VU92bfBbypUDsw
UwhurnBYtWOpJIpvJIrGrjj1tDcIR9IWgHnsG/XDVA5pvbfjdwg7yP1Yvj+DNCxRE8/T+Krdkfr3
N/IxVsKf9epeDykA/pv+njlCfKKbpdBrSCGau4KjkQKOvoC2rVPQVPAMn0c9AiiSrEiiL0uKVn8C
ly8BdVd9jEdQx/7Umb1Dgje+QmBHvho26B/CGQh0U3/6Bl/jc6m2bM/d0WehqR6NrUH3smb1U5g2
TbQbz/zY0e7q7i0O/cWqL4klC4y54gWslDhUYVrXmWfLwVgYydc3TCjzGOrvrjTEpCUdlD4y6pjl
RQ50oYnWkOeoSd3RkBlvsN65v/6cuVq0M/drpMJXfAR5v5/upCfTyWG/1wrp5HDEXSY6qpjMAtSl
G3Rr+Nhoqb/PAEipA0LBEvvZCvkJYV4VeJtvDpJz4gP3Q8PrCR+4faV2GUD9Nz8EVTo6WRSGD1xq
U9Aagu5/VKWs/d7rKSoMHfgbwW2PWjlRe4Qn81nmJ3bBZkg85ntT4KNkYT5oiBYopUr/kcH6TRJZ
h+IU6L3FqHGHbuJ5GqgwTIWLM0+Iy7Cjp8mKTpN4WtQiS0aFv2lIMhEYBDx0fsRnsLxfGG1MqebA
vo/KFhxo6n1nexHpovBvSJJ8ab1YEjRZP7rSKtfMhh2nG8dp1MkMDVCq8WkareD7OLi3K+NkBfwP
kl4GPyPK7bxCL4CqUYMpzJq2i+UqVikX1UH+CpC4AAVU5H2X6G/Z5k2WxMp1Mj4XVxNOLug+wPL8
3ourJUtZjWT1UThiynhoSbpCS39zid3Bq9vzE+eoaprvfpbp37oweHkWpTUvltrShqdS2dMmInqC
ocL2iw0wMGMtYKjAmwE5v5AEDxe542uwNxqjBpfVJKtUj6w9N6DRAiSKijoL6Qx1C/HWzxEr3CAg
qrRTmIaNiIYmdSXGf2+PYvNevkvfuxiZ7en9Q8r8LtsegHwj+aMIp4QLyrOk3bEFgjipn95YSy+L
T9HxFYltBelhm6+EqsSauPBQJhilri7k6A3EU99m7OBtPFMHEzkZo4c+UH0cp4wbfgGb7+tO+wrL
nPZiLM8O5mlCyZIp7WkdJ4h2LJWsPWAg3dbJhIQJk09Do2dtEVrwdPVWYcD2NzGbYf/XenJPBKHE
yjs6tMMx+lupdrn8F2LLBfeTRhdF0wyvelTeEviFUVVMiKBhE7ywgC3M1kpk0xMc6YOQeeEqeYiH
rheyXOYkwwyCaySkfBgWV+RERg6eyfO+9KNLHi3KR2La7diUd52uCaqTTbMuT+o8wzBRWSHPCml+
wqankqB+SwbQ5Z/gvqgndKLyjhGtEMM+gtCO1CS3+Qxj1mkeH1zcIUMUzcIerf8RXGmK1d2nXmOj
qxL1ltOHBkczqcFHsdqTagPSu0zUMw9wrcpTDWzexTtbP3O7ux4YjOCbob/LP1Hl6euZZrfYchz0
oS/XCglG8qrkuZkd6Y1wcc3L45N/I0+B0WUNXgu4/y6+DaYYecSuwW82esQHbE0y14JW7PWLIozA
KInJqiG1uNz73bxy5zJc/sm55lJv7+4TyF0311lUZ2U5ikAs3EGg9Ojn+HWYQflh3BplEa1DnLaH
ojaudU5V74m3fk5VXof7xl6UdbTiLIeAVVrNvYkH4ufM+4ob5GH9n0L8lT0Hcs7OtZWh5BrmjgRK
l+BAGN79KvPAkbhbeiU7DjNYa439gapOhppJ8iUAHjh+CJezur/cloxoLldEQ6ko4VNeN6/NmUss
w9e5BPYKBJLBEGV944G1zPKkT4rSM2/jZbII84mFPkMbjnGAl7QD3ogeyFRQKn/0xLUvLBW8JwE1
yiQBjvLDxYFBEQxwRGrNnOx6keuLYIzYI+Dleo3ry05BIgW2kwJiSqjsm0KaOgN8E/sktgFzGJWS
0NmPmMyLGmRMnfD4LgK6iSxStu+ozkpcy9sAFa7u7amSVkPG63bYS0yZw17f6/7GVzx4qkiIap0l
yo5tqOdOvVkhi+UUCRWbHtHlNJCt2XWL+ArDeoRFYgHaOqKuouvNPlNqEkwjWXPd2jV6zdlPUt7L
WIhbWIw5QrC/a5Vzj34DrGK0evKxYBdbfvhdr18FKJ80MMAd3Y8s5zNoxNZY2K84JCBxp4Qr3npB
KRxw9ERwn4xJ4Wdc+q8iAbLPKWy0kt77oIP3XpdqYK/MI2KGOoiQgvgLakrqEF3Gmb2QzJapl4mA
ybAGQbC1Quc7hDPVi40zE9NTnv0SZ/XjpuDp5mzN8/ZgKjvxM4SwyIfAa69KT7iDxGFCby5A+okr
uFajO7qFZwwoD5CcSvMoBsaSLU/z+QjbObBeuZGA+GvS2LEuTs/Vki+FvFDJbc1IcbTlZJtwnBd/
vtuBcaZ1C0Kso9/JGX4k4OuOnDWcWMyMyViSD0IjULky3we12KHhoXV25MPMg1mTYlaVOOqcBFDN
FbIMVrF7UarZKLUB9/TrpZ8bErdNIyHnFL9A2HYCna/+0g+AKjFcVqGNoK5qBG6/ihPxJ3tytwOp
fAQ5taiVoZqyv6Rm3HwlAWwKtCXEnjMECQox895cMzoUqcxIPThh1G/LaKcKZQZz6GrmsNUT8qpC
RfcW53SaXSCMZEiTNKcdTj1lps4Vwspv+gzqNGYiziS0dKOtirWrZip/hbjmNfjrB9ndDBJ/Bwtp
flA5htv+hevJkPB86FRcAqltlHniVsn8hq7qf7yy3GC26slCwdJ2Yr527UzsqwAmK0CvdJ//DWaD
fhmTDRcDwqGCkhGXYqimLQPI5x/WK1yvLYE4iDpQWMaSnejBeS1y1rBXGdm3GMLTecu0O7vSwuWN
DkNivW5ddAWy0EwV54olru83ZePTejJM4mbqnHOERdy1DFCM8RzHd3HuOVbwTvnpIquuoqD3vzx2
eYwO+cB0Osd8cpwALHu8itGtGnz1n0pU1D1cl9mMNqo6E9v1idXIKOsRZ848kPBjTRrzl1y3kfZ9
uH6hIhxrlKOdG6tAuL41Pih6mjvL7Cdl7pwiV9hsXPq3KnvfbOWvP73VkkpAR61N1XpwK7LREuac
i0AlJwxLItmlRz9dq28DAhyLHthoZ3Mdbq0yxqa7PKKP/xFusOtvUNTudVcnx4v3NdCh4mYjd6gl
p45OD+wUmrSDk1S+F+RMR+lmGxm12kB9X0QBXVww888psPh3l5uKc/k+NUQdWP+x8XDv7HgXzCrn
3Yk0TFynMh+eaypN2sLzjqxqdbEBvs8Hpa1pr3QK5jnFPf04ms3uHV3hG96V1JMDr1jt2yVSc8pG
AOamDX27u+3bTj4PuWUbwW3KAJjeA1nl9GGv1ksbN8x2SC3+cu0VRtgYufRjdMWlgLsfRRRyyOo0
cXS3reeyARuBm1WjhFSpkboku4e5rIrZL8kNUGT4N/ovm1ZoI/YZPgWU2oCT8e2S9IQlPwoDyKjG
GENBERX/8PtM4r9E+B7WnhGDOUE4YLCNV58bpdqHb93FNo2T7s6YWPV0kSoOdR8Vv+OTd4VFkyTX
gR2Hbm143+dlADpQGUNSbyeIJCo0SR5svGZovoFz66OKdNxczP3XOO4lc4mVKQtl2QaSPr+Rbgb0
KU3KPDRzZ3g/fNpR/6WvSd2Wzb7rojGL6oKBD0JsHYq+SytYs1Hm0vZCTmR1Y7Q0KoeYl3bAyBP6
ETQojmgUPlDX7BCQ2d658Qi3XhlAZrXIBk0DdeXLJ0MZtv/zF+iAaRtSmyliIJqEiw2HsfAlNrr/
DAkYVZRAoEspkQ48Xif/tM7eMvgl3c0eYcFf1QDOiy5sptJ5O+bbHNSWOvjwrYzLmmmc39jPfy9D
V7TgAqTjIA6nJMf41v17Mi9xeOU1I0d8nWF+skQZ0jE8wkyM3InAHUi5l7ffgUuYd5aIvVWp+QgQ
Loy9mh63EST/hdSeks9GDgFk/O8S8Ze4uyqHhCQUUK1Roh/ck10LHsiAFZKfGb2ux6OKep9h+ztx
JI2AZn0nBmD36x1CkuFh3YFVsvjVb8OdlNBYhAZWffBpEeEjRj56IbcKGhjwPqTisz2uE3IWwKkk
/Jw33gTgONv/vMLpDEgLn4bKdBMVy7fv/T50EbhLdw2HqeIlOm+f8nhOKpB5k16iVviT/miT3Iu8
yTzQc1cptd+0rl4KpMPSlBRhd+dlubrwni2bWx6RFRYE4nRzpaHmTqlrWN7F72muaYN0kGD7SvMF
XjEQ+kXXYKgwe2Hsm3RNqHLmHf7y5qgYTiiynjnY19ANNyeoD6OATu22enHIgu+G6wh+jIsoVHP8
3MvGVPtrxsBrH3QvuPkM2W7OIgPLQ72TUvhwFNmY1gnF/Id2gMTlJ76WOEG67GhfCuWz7P10Dj9V
I+pd3XMb+2sBxvkHynlQDLuthwVvASeGtTs681lSWUnPmIWShzzwW2lYU3+Pz6Bdyps2uj+j8X7U
UJSSCwSm+3kYiIuH+YjJvG/vAo3FWguWRfBBmsCLNBG3mpMJ3A9kC6r7ng4QTIdYsv7GesiW9Es0
ZntpvkESdSya01XgzBu/tzPSizyU3yaWMUJkx7Q9OxleEarZZCFk+x96NYLJrrbnnJIQdL9tbWpp
W7maGK6JybQCtwCWDam2uWYRJN6+g2+nPKr5OVeaA3g0lJchlftNXgs1OBMJnZAlWJ5x83aLzu9B
UOpep45H8stci+pCZwPBEx0g/BAmCsciKr1bFSVUWXRrQaW9X0Yc8857/xywVMBdulY/D3E+a7TH
Eu5wA/zRDHqFKApXlEDMA6xVAD9bZq/wT1OeW0qJ7FYbfwE2iS0L9xMd3PYKpJnAzTh2aDFZJKsD
lWtHUp8OxTXJcIqA/MTPlwACg6Smqbtf9cy9SNqQP7++GjFk0p46qh//48NXb1gRCmsn331B8PPD
VCC1Lzw6KHT6dKspQs/9ngV643iq/ygSmyvp1ZmLIpXEytQ025FInsJ7ACTfSZ4Uzt1xSvFSkctm
+VYMjYdkF5/sIrFF1ZJAc5ioxN6vqTml0eAYE2zIJDPMxEIMh8eWPmivh5DbLY1UeEAEAzkq92uw
4uxNL8MPsHusL/XeN4vJ+RTcDGM4xvacy7ARt4Akz069Ykk8CIoUubtZMcFNwHpN0k05xR4Gay8U
ieDkJvYnWIbvml2CJSBBFWzVRZ4eJgPMQoCKJHu/TKMA7majIDmL/BVVtxnDHATvvFxRNRbh8o8/
j6dbUKDi03ziT5gyzd8Cq+r0mB+wkVxd7vQhe++uNjQkUfgTPaBjT5BMYgodZ9n6kMP6TyUMs5wb
W9DfdNX70ewsrqTULJb1WxdqXu8E0LEIoELvLIVhf7K35M3Z9BSfgztJxXtmHsMfnxSyRrqdKM0u
cIbl0UYrfZF46tfOZaBYYStC08T+q29BsSAZhs/PwxT+z1kNcMp4VTfwcyu9MzdOu3Xpfozm8ydw
gDuWJyr2MRKMSMdh1Ek9wp6mp4pbHFsHlmjHIOSd16DmexDRAwtXkrr544PFKYZlzQwuyviTb5kv
XCRJUSgCYFrvSD737zKzlLk/utbCY40KVrNKFrakMB9Ddyfinb8bnEttKYs9f58XuZy60lTHfOyY
p9xfhqbPJlAbweUzGOxrj/bTM5Kvch+Huj1GjhC1M1taPkD/ynpyCYIle1aBNqE6Bn20bAOCQEHW
eU9zcU6MqWkEBoZ1JTZ0SqFdyK6obB/884q1VodrmbHKKtFTWRXjjAcqVsgtpFetOmmqdzn3f3Eb
c0BhiuaoE/xBmphZxphuP2vgixmUqUbZt90+icsRiaHzX553UAKqeUUtRIlHjDYSKxQgsnwkh2AJ
hze0BBIO8XrhQC5eO1h9DQS7M0T8OEzPGZQr6X5Xqb+xSm1e6wJXzg07qobpfm9oSdUP+Pe2w75t
bZMMmPAmSofAtuSQLd7HBNY8eqfWWaBF7g/6iH55fXaoyqO3lJaxDDyXiu2G48AHN2zyqCzFI10S
8udRfENKYVdw0Cft7DRbUtige2zamnxCP5XJjKPbr4703lpYeBQR0nrCtlmMMbgyhKJThmvEQVHA
tRhrmXKk20kqpLycL/I7uDx8ToWjWX42EJN9oqG65lc7OiOt/0sa5/W6VNEoIEyKOLigbcscmxO+
khm1CKqqc9YlxziLxa4pd4VLAy/hw+3lGxQ8ZqurjSg1oyfk61QuJXC5BlOslRG1iF6JsCf3+sCs
Y/6ldIldg/FuGVqiI8QEjPQXnVGJQ/1s6QcbJc1W/eCD4FGlUdIgHG44GgZgMM0is+xr864jRl3Y
Ufeni3Xy/K6mELDrw3snrU0k9yKu4jE1aNt/dAk5J8TTWJCKfkl7issgdf/c3RPdJpfkHlc7O7L9
CJYwU39A7QTLCiUHxkui+wHDWIPTxaTOrcAMJTa4fi/h0umG1pvtYTzdXJIkW8EkgQcdicmWkpdr
nA7rA7EIm5J11883qRl4+wApYywkRUCze5DXI8qpdVvST9KH1WUVHpmEX3Rtx52BeOV6eO2XBjnt
CQfNZo15JU5J+31HUvAhLOHVFEtP4T51YiCFkNMeXY96J7HZYP0oahAiMluSSinlpsgX3CyDNJ4p
hVa05vhVAPwwXx6GZarirCGmxU5zEFQLkeZEM82Jq1ibUl9tWNu5HrO7Jns3wYFDSGc4toPTzOLc
wZmMv8gr3yqtjSftdJJYJFvrv0VfeLZYU/sSN9AAiXqaqfbbgmfVRjNWVJfTkJ/rt4/6NLhyPItO
GQFpsJhFtQD+a9P3uxBhP+gDBp7+fhLzsrmURn5RrXl7Lo1LuLtDwS+06eB5LIu4bw0AE+UCotNF
xrFJgOGpHWaZ6GuMSUT18qcabSOVxqWrewijopzWXBtCeLjDl0+XONNVSVvO6HSZnglyeI5l4xEH
J58Z7+f9apF533dQJ3u+otjuRnv9dk1uH09eln2E0B6h0JJSMJl7FjOkLcj0fjCs3L4pQFal5NnH
MtsrSZWfmAegQVezaK3nLh19mIALZZi1lSywGBEoFvyg17b6YbljkeZ23PIMQ3DsWqokKq4h6m5K
IOdOwaaWaxHzScjB7/to4fka69T+j6HbaIgmChRLIAd6+RhAn/hrHGFcDag4Hghit4kCNNcARCkQ
RxdXtdBPv4E7shiC6pRXa3RU/sARt0JLUMoa5l2Y2I+ktf0PapgP1Ussfu+nW8gXT+VhBRPqKRAK
XeXkHZVUiDqcGldIALEfK8y///Fi+gW3TEnRzVh5c16FIgDqeQRGuIfh4jd06sG7GGMV6GLbPsWl
8g2XPrTKJlcigp1jGQ3ZEN8Ktl/1Y53VlIRZbInOXBumaV5UcfaVXx0zjVctTZix0H2wZyRUo+L4
smkCh+1qC70UPKM2PqdHnYq+u5bF64PELoQmMqMN7F7cm/8XzvQqC+xOjhjCGXk5p/HnNLDD8OKl
qDHto0gh9jdet6RCuynVf7yn+sCkNmlQsqmFvrFY1NmVs/UcRanT6eFh+hHKpbyY//USBqRP9GKo
XmH+GZ11z+qgWXdRyRo+XU4rRuh3eatmcWEWcLpf0CT4YuhvFrD4OJ+WWCMyLH8WSHLbZ6jmIkCt
iajTW16jWzgCbcB/SABLTcZ9Z2rA6Zr26tmGcQIB3SjRTZyi0xV1CN1JybwC5Xpgv8J1sNw+Sf7C
hQd3t/1PT955PUcuQsS8aygnpLuwRwWrmVxyVrCcrqK+hTBsQ9R/NHA6vCFNecVH1P05Djuni/kv
TYWmSssefwX2+JJcXu2hbMIKA/F3KWAvRxP14oGcb1OjVYmeMCO2oWNjlu1V8KoH/+jdiKmGEHpx
AtRT7ZAH8zYFzMzQtQcPJoFiaoN4pK6rOpz47nqx6ghnIDI0RSbb9XMSHGX/Wnha3wSPxq6FJMwf
62Ga5t2ys41M4Rq+fW2EwTVoJM3w5o3pjCUPfwRn3LgtqIiGoYZ7vVdlFbpFPqhVi1lw9Ny6QlV3
hZ0nSc2T+4u7tDDkC+2jZn2ClKCf3ygoaRVsiZCGC3AnIs9XKBOSbU/7l5z9lpBmpkSA51WK0Fk6
9f/x0cOe7MGV3gj0kB3klY0B46VM/IziUulVRdM81qtuBuOnQNg0V+1s6VsnEkH++qj3J8BSNuft
z9eu0dHVeBY/m3jvIGO4TB4wgG14JNtQgStH0ccNTN86Y2nLuF+DC49WDn8ptAYfOkwrKpsPzMuQ
tmFuzrQowKlpOlo/vpQ/6jMJa2PNZCCJZ29PDSi4DLDsRE1Drb0Dt6jgPShN6oNRPqIS3goTshX3
Pd/T1a8wIsmWNpWI2GMoqgnMX3UKE/FNzdkr6SbaH2E25rMkrPr8PPmyDRJvPhMpE0QPfb4XQ2hO
I7nRQOhKKrQavDJ38Hute1NVfHP/kjr57h65ek5jp0h+jTyTS0stwAZbcMUnpyLBD07nCHttk1rX
Wv5xhfZSNNakwA8IuSM+3uTKBhFyFzC/qtXP7AfUeWFUzlow49u6FK3EbmHuTprMDnwPXMBq1JTI
UZUcv99y56wS9bnkY8XcMxrlIqtJnhaEQGWhocSqSaTx6KARat3lBS/mr6yB78UyvG+XTk3Cp2Bd
W6AY3cfRjYbZOi3cPmwGslqmg7H4iViIZJ9PmIsNcHRiHOAPR8i7t9rDxRJ0iS5PmD/uY8O1VrA0
+dFk+19e7HIgSF6VdX8UwMBIWJEXmaiA/XgYOD2zOnBD98tRIINr4kSIPs7jCVvPPGM/UAgTu/qn
T+t0o+fubm54NhjTlBnp3YjnboBNtA5Y0LTGCDpBIS5JCrL6vBYa+Y3ox2K5yrAfEpfr3teIydUS
l2o0f0wc+e8GO/RQrh2G7SBoneTkNGbw4BOoZiip1Lu/h/E9nseMFJzO5k4gkKAZgDpq5Sqlcc/y
OU6aHSUz4J4Q5yh+aFrYlMHtBUaK60Epwg30LseeZQpvOM4YHd1OJKm8WIF1T9IW7E1vd0X4sdJh
r74pEo+78l+KPwb8Wbyt5ze6Tl7skOOalyFrcX5GLh7khTjhOkdP9lg27Sfp2O8R2v23U73c3q3M
D5Qtpnjp3vVmZYFtZTdfXIgykLw4AcciiHjv1MiGtK7tRW5xjahvAU4HDR/Kcq/2KPP8SwZh1HZ5
PyiAUaR08wseZZRmSynlSd8XgeamIhq/oayYNo7Os2vZesX6ccZr8fPfzuWnDRmOL+PeDPVXA+Vk
/c9g6OCHg3HK4G0Hap8pF3BH2NnpKAhOQtTvFfIr4r81TJ10oWNvAPLieL3F9i73E/dJUVsnud20
9hwdLzKSv4Y25uAw8sSnu3a9wssw0DB5KBL1UbKKrkkFkRIzVUM/D3llW6xRrW6N4a8V+ZbgOjWM
0SVjvGzD7MoPLEvwBjDFXDve/+j5MTq3bQcfovPjfxCCFEfohOsaoLazRx5JD6E96aP3JxXvXZu6
v/mUKOzBmmaXfHmbYdHtbbkrbIWCmi8guro9L71PxZeVFgGSQFGLrNhvMofwGHkiKmjO2qWSopnp
eomkIPwW2RPUseE8H/lPYCtlSznphXxqYdfX4zJTVzIYOgzAGRmldaA9KkP2UevnkkwVPa/P+gHB
QoGLXJ8JUcsS1zxrsyW5C1BwXgPzQmYdbrLXrAVJDIJoflmTxf7pN6UfC+RtGSjGyQamiBTgC2+E
Zd6eBwnsAn5Kaj5OXIXC19CBtMMzB+wZwE8VPE0U5legyjCVii5U1NjnOme/T07Ekw4H/cfCqy58
6Oc6zpjE8kwBrqei5vCJjIDLj+ZLmlpII6YHKO67BlkHcmGDmwszgM7JraSWMSGl66hiMWO1mbS/
XgMPqB9CqQfWB9He1aZ5TX1Rp207BQ37G+16ST1sAUO9oxQlOXNOWgDkK6jcnbY9xQnM417MPlfK
zb2U7cJ3CwdT3ffBiI/aNUI73BjxLcJE3ORHabxTFn4D4pDvmbduRO9Hy6gfeQupHtnkDyRGAJ7b
qv4evEo6rQYr+SrWcQ4Ulrw+L1pKQfkTI0TCfRsvuB7x3ESBeyQzQML8kdIv98LWksM1FFo1zlvD
6O8tW4C52O1LVk2LQhfTeckRA8jEzAY7cyQQvJyIh8CwtWOKap0m7uaIdskAnQvWdhQe4QzQsR3j
oXf7iYpZgwDuvrbx2e3hgWlMJx3bhxgBlNsuYeor6ce7p+L/bA3Pwm/PEUIMViJa461V3THEsv3P
NPP3+PR73sA822SBWNNLffQP0J/U5Tb669Oe0Nszuh2o5rnKoQ2YkESDv8wXC276oXvDIUWKhSJN
pec7OaREn5c0HKkUB6PpEq2zVvhMu2WX3QUli3rTWfB0KBDzljmJ+6UOnv6YhDPIfQQ61Ng7oySC
7bI49DT685mD+jNfHMLCy3o2RaYoRcvnpVZwWttPxqcu4g7MA/jNEifcaHUOs1AsEPKe4MpDZDiF
ZlRW/Ug5aG/VK6DFHM9MoeebfcQyU14Np8/uS6RI3RBYp/sBxaacJbUwKnixkCh81e5Rzw5Bpd5z
S6wZU2A0R648n2lQ63SJpoNDZ46c0x48I1EFjBRg7U7/UTGSLPbY35/UlJN2nY40aJgIy6+80DBX
CJTlbdyaHw1XG9Ox/3fBBErxVxZSt+ABZHH1Bh70D3JNC4P3HmgDfvLSDrzBpnp+gebDcMMn/e4u
ThAFqs9rzeHAi3VLkIlKCRJXg2uPJ11fQWFENOccpKgKzwfF/ZNTH3msYUQiGedgYF6MLbK1Ci/6
YURZr4hMIrfCZ8J38SpOF7n4MUIa2Z9tet6HcOkmAtoOQl/c8DKK3Pyl/b2WIHAV12kXFpOejPdP
M4IlPbcO4bcN8yPvxi3ztIYqfLdRriW0szCYd/SOIEVnukqb1Boz+WMMxj/xy3zDBOh51VUydtjA
n9oOsGgDH5Ev5U2OPVT56PoBYfFzRZai3N3pnmYDnc31IO9B4rdmj2d5eXCUTTihG6264CzeDc+5
w7fOGuAQzEbMoaDG6+el0Hfj7gqxWh3dbfUrKpEho5XI4ye+VX9Z8inmHzxHtotABIpnByXQxdp4
0Q0U071ULTNrGnI8IAkvW1/pVotZLBfYmUkTvBRZ4YzMmIpu7SEGiUEVgCftqulTLJHzW8xcds8+
eEXLLA6xFlWxZUu9lreORts2/pMUFHMV1lJIi6Z08nUP2rVBL122Taf6Gq7W8bODjUCqnifI6YmJ
WaAFBUySDBKHgIvDubS6Z5fKnXiYpT/2LS13DrlktZ60lZVuIVo8fp6ScX+2wQY8ZFGkAnK1P2a2
/+0E5/GZSXxnmxXxkIfq+DlfknUkpIh+Zmk9GdcYEilGudoyVC5tbBKzuMA1uGis5vWffN/Lxni6
gJbPe6uz77vGFcagDjEw64kSJtsx4Ia9WvM40Zh1vV//Zno9blesJpPOqngIOr4X/E9r7m7mmJkm
J7AlYfaphcHtEkDU/OTrnyhhSmG6G2oFgg0WY86EvWHqhWq/hVGv76T8jbbBxgonT8+wr4FFHy9N
dO1D09cMsjUFc7HnNmtHBEtgU05PaTMjhgE0aBqxnSKFSItMaR/i5wpqZBFCv4r6chQxYtFME/3Q
R64ggzfb25QO8vUcd7CvDct+lVVV1i1KaUsXVqFmXhKOz3oEtjERPESfOClZ114ADGce0zQGprfc
2uCLeLoYswF3Ld0phE56Slcdaz1P/GfB7jaoIBwRsWtrVyVhZWacfo+MbIZKisqaJiEkiyRLiSPP
FuYI3ABsSKCUbG7q19ZvJNapTk+QQycO0StJ5kqGmV9pWL7OtZQKowEsj+cKCapzOFIiPs8Zo3cn
89YeUh583opYQk5n0EaaoGw+8EqBzyBHS92gC3+BvCT/ZwR36fKHVMjMFXl2EdwIacVozG3oC1UJ
4D/5fJbRb+npT/S5zg2nwWMfxBFgBiMFIaukzsbUqLyC2AoGEBX84KNdqOD3yTME/jUO0E5jPtcq
st8KNyXaae1HPPDLGNwsn4TlZmdfXr3p0fnYJSpsUqx5qbILVf0i7RvIsR1CX7DywZBegBsDHG00
o2ruffJyjmW/uu8buKWzNlUo/vqZ/enwwsQeYAwVyCn6pFRv6psFiWTzibIqR9VjPQmSQdboufDq
I9+YYa2XZMYDsVSsUHfFVNviyZr9K/XM+TE0Buet+dm9xn+bndA5Rhw13ToniAvhTkJcerKBOfmo
V5BxXLFgdffHK/B+ROFhbsWKDeg1e0FA9nQAvxSUGW9B0dfhPKKDfjh1aTKmk0ZywUnhGGkfNekh
aCbQKNdNqZHOQP1UUBztYQNR/3CgkAd1sObh0UOR0/Zgt5awi8DSxdHfmmJCfXmZ+JHGgrOhDMJW
XaQvekPA2IDSw9uWOkqdAKH2bTw4P+cimf1M/9YVH2ktg2tygMOsd/GeTIL1bauEQI+9JeaixFwx
fY0MY3XxxSobhWeJNQZlopDPgbEcr891wy56R7jKnsoJEUbLYRTUe1DznSkEZzIAK5tZHqR2wga6
lodEX+yMiHXwOc4uPNN+Ar5LWyz6ooUfJkEheFOqAh7dIn3+M6QqRK6f9J2Y3060K2lUAhrHIrqv
qHFzrQHayRrM5UIEJAUIlk4Kp7fTjXOZw5495KtuJkmQAvuSQ87y6QPkh5MNLgOmzIot6Hup0mip
g/CJN4+djTcvNppW/RYOsh+AkwN0iHe83ODKldLQ3cZDA2P5wShnyqKic81zGESfQBc9ydfOZqBl
PMN9oyHqvpBuZLFxVHui7n/c/gmfZg0FDuufiZOlJAL+heIAymO+OuSKFqcmh/RP2bUXXLNXjBZc
6yUQqlLB2qnXbJdZpc7BZafcSOAbQa/YqZJdpq2kKr37BLq2lkbwJjelkn7H5xbFebuHhSxx40Lm
IF2IRR/47X8Q1viLE9f9r+XBVWacoJIHphgCeZOnDDjabRLvf7fvYSS6RGnH5L69acfjfgvU+fMr
bxbGo+NRS9lXydRDz1TK9pf3oCL7DuAOI2SfYjQoFGwigw7PCC1e1yOeNEczvL+pBWsntp8km5So
T5G17NFH6wjW9ZguSIUMJkS5mQkHM2Jv3cocu3UCrII19+yHTMtvnuP3lsU1bvkMUIWfRWtQrtnW
6omIXEj6fXmYSppC2k2ysVhnxXlNqb9fR9QzeNpgSGPgOUiaqKfCmG++nUqO9izOKpcHyPQ93JHA
FId9YxbLX5etTCLc+qs5nRSm8JwNzTprhi2f5tFLvNAMe0M8A04WI9R4OzaZBxwX4Y3lZZygSJoa
LYfk/CeCOTGULMy8J9+nzgaNarCDlCF3bL4LqDpv0iyrmBXQcoLrX44cwLByBmKnG+vWf+AH1+mp
SHekWRTl/Mf4nzG/XJoppvZ06g/VKDb3ywvLI1s/j7KArx6SO0tbdiiMHCWkpx+1DminNmII/en/
Cqu03q+nWoCcVrCInaKBaNYVuRm47njzZLulajIf2hVSPDz6mh1sCKeekiu+MchQ0P+kEmu/gZZ6
r5TCA4fy0tj802IYCUA0YHBFxn1DQmBfizro6sl/bDuvl8dbcdtdtScHclc307jOkjWgPz1qFtaS
fNp1UhDubh0zLHGFNdTGl1/YKNS95zhsZgB9eWHVglwjJGvo576rxNp6D0UEOwrAbCTlow6riQ/B
LjzoygkDeFDEcrlk802O0Wk9a4qHIypyx4UKUE63NWCfYpuuw3MnuPXWGZsnMkIRPUeJsmD5Xg7t
BKF66si+Zq3z6zQNlWX4DsbZkwnQVsMNO8EdMcyY/O2t+bLAKQzDocaKQNxgGfZbDfP5ZhW4tg2g
zhYmYaDmGemMm28LdnACwVw5MgwC9Y0Ccnz+/2FWv70NpCr6UBR6gJbjwPrhkGP0geCe8xZ/BcKY
6w+kx0GDSCUZEJRuFowbEbKMQXdRMBEs3hEoAQMijeAmc4FSkcK6Svcs1J1WY6af/AvTU/sf9Ne7
EaXq4tIWfb0bUxwmXuc+o7Ite8mF6iOar+WV5DHkpakzjMdRuGEKYi7qdcJFrMHqkijdACxAPGxY
yxNtGrsIvsDN+KSXs/XAqbzp3n+hANBCV9qfv0069qxuvPTQ2r5fkJgWAKvqvd15nBSOdpd/MSui
F9Y/YrXRhgjqhqVPfGdGBSsR+OAGqPL5JVl/SRi+KqGeRzFV7jWyTkYAXQbC2QA60M6Eiq9KiW73
rho8LxcHl96OgOKIFag4PcRPT/zHfBpJP6ItTS42btDJSNy8f8x6/E4noy3HMuR1cweFriqAmUqL
6iwXFE+axpXBxlHQwOSJTimhK6MXT0g2xJ+R02sn0vQLSxLNzTovQUFQhcnCQlurD63/n7roNT/r
+ZXTspUTclFqBLou4pWrSGNwsgcmD1Bwj2Or2Wc738Mt/mxyWI60nzJMMbLmMUfmYNvXU+EaTFWk
IYpA+bQkICyqsLfXzJ/9EARGMVUFrdGN67mdRYLIBnPjo/3hlBgYBTpbJtYJbbJTVKmx7EVpHF+I
dBrweQqpERzPaGmvryJAWz3IcX5qm+SOFcUOZWKXJnXuL+dSTsuevCh6ERiIj5/SwFlUticvI36D
gJfiQ95/smYawd5W1donAWjIGtmcgQ7yEleZ12ZE10juJ6EwiURn2lvdBAI9Kqyfv56HmNpSAS1Z
0hfV6Rw3E1tP4pCJkjAMhFsRYiv62WrS3uxTOPtd0WEgX+FM1DeLj5/dg2eB2tu7pcSI/kHbYnfF
AtO9nbePiBIdF8Zq4zB3yeFFtqgUM/kDOBmjRX5eSX2SaSMoz2Wi+43pLe80CJ5RwzDUp1DlkG32
LcyMYnLvuVv8nfyin4HAwG+nmxn5WjmptxaXnc7wFZX1LOwoV5Dpydma6G3gIxJAjSLwxgm+OWa2
PEot6NvqOcRNNq/+HlrRRxitQo1M0s+2m3NEf7AHzhUCPkCml9RwYRmx/AcFY6zLzDyFbIdp94tC
hoPF0pOSEYOUChZpAgBCUJOc+vnM+2N1GHECkJOeb+tcxYEc9kYFODs1MDNGTCNvp6l6cF/41IAG
IdGU/1hTUisYQWyFek2iHDSAuAGTpKtBgpTPQE2gGqHefxZ536DTGQ0azbd7rp49ir2E/aLv/iR7
a2UZI5/gXgo+iZoyyFwFX+tnLuekkMES+WCgUhZ+o/SOZdsHEeDodMM6f6eQGZKWvxIhiJZYsvFV
Ql/MiTvoyp/FxnqgF9ZBBb3MlVQssy6lcSiout7lXM6kqAYZ6bPvP8wVtXB0mjGxXN8HbJAoQudr
EDtXIJJAMT9LCjF1c0miM9kgOlF1Z9q7j15ctsRNtgFcAY36CZ0L+pqTMSro1YXf155DDSGuWteK
OIzFE7GQTtlDWUnJkT2NBOrYuy77lqEDq0PtJ1NaEEMfkoFYeBwWXj4W6D5BIw9ydzHsEFTU5V8w
5x1p1Gq8AqEEVtzKOWkiQLGzFwKmgt0HM04qxyzhorY5Evqa9C+R/2wKQMcGbzDGi14AEVxDpiCk
9SU8TdHxWtDs95a/aIJmmK48MJ2JRKc7oe0wHphE9WtgQmull3d4Jh5QSSaWyFNvwZprFPwA97WR
Vclan9QcOIPYR8UI87nyadf2EfL5cBj8iqfYa9vQPgSXLUsQ0rsTspBLLq+g9QRTovm93iX+4fKS
TWjUu7dV5ZrIyaIHxdVCp15lrpF6Kgzs8faSTN3Wo7/mC4dI3F17upNAWrpZZnMX0XgoHTOLvPGM
DSXNr7ygcg+BhSkCm1AAWoMqH+M0BxI4LVha+iEWayqBgDo0R4YQNeMuUnKxg2pcJ6Ajq6I7vV8s
qLMQG3C1QsIcTGl7tH4yNZX6z166E3er+Z8Kn7cKp7wg14RjdF+qki05gigk+oL9A58KNSx77xvl
778KZ+SV8vsovFnZLawQ5q/iCg/V/6L6DA6e8wS8fyXajAm+9ZvJSMTPCnHs2/Bhukj253mLLdYQ
pnEi/Bxdze23J+n5fQRFmISVQnyvE72zC4aQqZbJDOzih8kxmE9SkCrbC2wtbqmuAMKjqm8WgaYB
QDMLbXMjenDFPxDhHKcHDEnW4xD1DILbRYph6VD2/c/OvtujKJ3ZOT9v/TuFdnc/k/tZ19H93cT3
c5FWflXj9Ehfh5Rhas0+OjFWSLlNtz86V2uLjI2+tkfO7ida/gbNdZZvQbyCbkSyBwj6/qYcoMS/
EzGuUboMMS2mvvFvW0ouv0ClKBkOJ/JtzUch10dhjUwAT2YwbmqR3M0pwb1QIRVSGq8sOZIyT+nI
0Epgl9EFcwp6C806QqUyiF1nvVWPYo+dLAXI4koojYloWpw3ov6rd5J8lrm9S+K6hxhE3MnQedDs
IveTDUTKUNcemFPoER3f2YC7mRVwkuYYZkuawD8f3s6xJgag1F61RnqMkV54GJVBT+ESPdlHPc8/
Wo4hR8a1TB4hkmpgkVXV01hzjQX7omhjpfyUA+QdPRYUXs0jRCIt6SVw4wETBb//SIlWkkYQNHaj
h4Cf6Jw6zjnktAkVugsMXfLGjd46hvlKUMimF8rE99dPBdtSNdlvpYkO4MT6mds7slbQgIPwbkQg
A7h0Jo3tcqFCBJ6jJF7KG2SJFT9TRBXMQx8Pt0ljFUsXfPzLJTrNuNiZh4J0Zv/c4KDEJfSGLkza
7NaE5cGL12DayOLh9T9I27UcpbAZ1Ye9ZBYXVo2hbZPPtLfkbk/NLTAFUsERCRqBRpw/Kv9eB4Fi
y1c7S+G3GZUDtf8J5cWgskEUdsNrOhZpTzUTGis8ePNyU1VezHXuseTVkPcEvnR1PTTalaqSQfBR
WzcW0g/FB8xMT6dAjHj8ysjDK/J6Q2kGyyp3gWZbOttQ4XP7h+4vujRfT144BDgJ02b8ltKDWEJz
DbFlnviNrkyJAE0gY7nKt/2Az4A1obGeUPjmjs3FIGPYNbiljy5UipGVGt9OgRPp6KCUPK0zi+bx
b7LzpzD+msA0N5NDcLSROdu1dx732AESAU7YvXEByDmYqDcym/C2cgXDZVRUWlZzg+l7wWZ31Le7
Gos5dxpClrIhAQHAjGFGuTGfoJJTdZC34cQunRj+crBJc7DSxu7v40UsNbtcIvy9kmOH42XERIPD
+zJFYeb5kIAH8C7XF2zXexhHDJeonTRhhCkHkc1qBp8ulkY9gtg6UPZnctkKeY5F9HjrL3RTmojN
YFujfmqyq3IMWKjCiYUpTvGza/vpaWRHw3+cnIKqKWfBOEqH+kPFS3922RVhv3FHFPDJWPOj21dN
BrIhLnNAGgwYKtT8CintsC/Z4irn9Ily6gZA9OfDgJl+oGS4cXciWSVgeEqmms+2JmNPM1BFQxXv
lF6o59eVY8qxPyC22iqeKyAgp4iWTr79i3MES6jDFluWeze4cDmSt1mVZ0nYBFpielgfVqaF7poz
qtgHVyf3yMJASYsYAFThIxIEeydtrc3jj7TMfYV4YGyeVzFlrAfWNyxU+dPmMuHhR6f2GcmqTou1
QC8YVvyshpVItNtnn/sk1O9gioA+ToesHz0BPciVtVu8nyQ7Pn5gYmZH1FyEwVd2E4VAWNCqa01/
YOpE99UgtuQVPLCgfPG/t69lfZC8Iqqpamc89PEMGxG1qcmwrFtBc1zZNqky+tob+/Liama7hKLF
o/dWX+SBmr92I7X3XDmOi1wp0wuqgMW1Lg2QPLh/1S62eugdbvuCWrqIvCvmYPv34WtwaRhT7Zic
PHpkZzga8m2B8xKCbnjS7WUVhzbX0wtOiFcVthqxmxurfHjY+SWJqtLbdwF2Q3qdbvbdTUQFhDyw
Zs5/lpGN081HRY7g02MREBkOz8Fu341QSh8p6XrgS8bvzxRrdJolLLEfMGrtnNTKtOP/xQeJRsuV
gqpRcYoUP/IC5/M+dCrbhJKuQNRZh49cCQSTtjQLfbLEGFZNRrI9x1DUGFs++KrRowA/C5q2ilG9
mTiZgO+OkBD9pHGXalUJhhcsDOSIbZVa0vq4+aQeP7loFlxuPwFZP21t7K/gDeP/drEmbyhbmQNn
xY1mahv6ShQJIC2aRscCVZu5mEY27cCUjO5uAFiMkCRFAwtnaF8VYBY92XeJqVN1f3Us+RRpXphl
BCOSAvoNsbnbls5wvhJEY5i1DYDjfoJayiNS856e3HCMarboMiuF2tvSVnCyQfKh8QAeuwCewgWv
/v2L1kphpMjCS6LjFv/9JvX0//LIs1KgZjXWkOpQ0a/9stdrl6oMZltLLfEqyOlrdACtV7j/OC+z
KpjFUv/eJkq5YlWIwNlaq6eSv9winjgsjtCJaJff+HTzsnu406LvG9CwGyVRE6L0vSCxcpNXEWo1
Pa7IVTZTU8IKb0uCC3g3MWbvvM72ex/VoarEf5i4MIvv9HzJFHlDQ33glNVHag2DfT5Tl398HaZe
gmotYj1n/F5OYUsUQLR3GvE87tInxB1ND8PyA44nMelhsP6EEJ37efvivKDrtKfU4pVvIoDuxVSz
vVFHdjwSe4NjW44wHp7HVEa78LOpFAEQDIO0BXtF5hBnQn0mPWb4P4KVzfLnq4v+wxdCmNT/4JiZ
v0IY2RAID+uBHzpqRUGE8rb8Tv65dod1tUumq+BVU9RdJlFTBK4Fx+IZFwdqChZMc7KxVchyt3NO
wBOWYY/ymvxS7VPyw1AgRgJYPyWIXdTWYD5A2OLnAmj6DMLNrgi9WYt3chUs8V5OH//ebKCd5fXK
KnxqsrN/dYcYA24ZvLpN3qGLOA7bJ46MMxKEum5/A6abHL4a9R+4crznyi0LBZ3u9vNNkekwN6zk
zvmMQHE9oN3a4Ctqs4vfYwIYUJPOarNX9PcE9z/DRmx5TbwHFnyZ6O4mHj3MRdin2pKB8dQXbWtj
i9hVwZukZAfdukDoT9PK8McZrpPkU6MmQ+hjKeiy1wIUOqcdhYIelprP/0mMMgNK6KpVunIfpUj+
au20PDsZaYWxaJccvCKUDDQCk3hydEnpCE6y6767K3pjquX50MAphIJc5tko30K3QkNocZaQVxJ9
0Zth4nIaHIPYjYR14NXTkPgC/dN3tDW46R/fwAkNxf708dCSY0Uj/1d238orvwj9DG9P7AR82jL0
0GUf0y4f4045QCrqwItLJEsFStMkWlStGt9QHlRAqdyc+vhNVljQbrmRg3HTyVpxa+2EWalWNI2T
bWOpvfzgltEAnMNL54mk1LMpyoYqQiNKImoP24ISEGPJ81i1gz1mg9pgiXObTHtejVTl2KscBCBK
RmfoUunYmeC5b2AaalaHZB5AB0VXGuIJNXS/4DFTl5uWsqfFVBK2OKbajx48uR2lInrPbhB9KR0U
W3LrPkp2giHYLL3WXUECqP9BKghGoK06xL4eLwhl9x5CozlSOlFTuXZrTfmDx8WlajdpYqnc1QBj
OcJWuoeLoq+M0SpCcWahFUER3AvICVQrOSEDkRuHby8n4EmuIN64huRxp0PLZb4vOq9oqVjrDl74
rtm4Xmnwzdspbcg2NQDTuEEuQX9qtYK4nVfn70IeM1qwoEzFxLibkCeZBHy8D5s2f02ewl8Vf48x
XQR/4CgWwsfnHr6aD0SeVA7KtebZBxyvnHut19Ca5yupZOkZfywGuQ7UK6Wsah8VOuCUjzMtjM02
xYM6pgVcIr9O1sPcBcEk0iwotoP2OG6Il5gBEg9QVQXUAUIntKVFl65KtEahWicGKdnSGWME0XNh
f3vdpsribtI4ieCo0MwqQRc+hzTX14ZKIXyfDbwffMiYKZJgEUBfyT65qNudaCgyKlQilTE2swVO
d7Jfq3kGzCnZe6MOwx9CRDhljo2WO8NtkcuppeWPFnFAQnJPHUiEU4rLxgoXmFOv7kfWzXBNgbS3
NnqFx6+esfmeL96+B/2zYPBKkEvpwL7XamrA50aLCeqYwg8NBmpHQNHRokp++RjDthPfEG+bIlJq
jvazQ5rodO31NCeKhjthKUnmkul6mJMRQeG8M503HaIcXZxJPTqvB4jZGSeF1yI/kZahx3wYrKD2
QhIKJtxoyG6rRDI8YXTVbaDlcljPpmnEjLtEdqGe8j0EavKl4XZQH4eqsBTP6G08jXB3L+u4YcFK
J3puSmNLq737wcIoGaOksqD89G+AnpfkpcsZihPqQ+mdGBYPCIMw+pFH+gSCgDP8PGmL60MGnqHp
SidACnaq2Dzg/igQuYIvRTl3FPladgzCa1w5KkiJM1jTvqj68FbCFX5Qexatouw5UhJIpe+Ez7p/
GeJ1bYBx/y1A5KLeZu3n8rztnpu5Y4jZ2kgg1Ebtd88W54KK3jCWs/5hInfEK5DTet2rigwV6VnD
Q7CHYciqW2p7B/sjWVHLONypBQqVCuwGXCmsaQdNxlq6J6O9+q7HyzBa20pHNiv+t+vZlviWei94
PjvY5ENb8OGiHhCHPy9A0OarOxWuD9e4PNboeWJYT0RQlheNyrMKvr/jEX9Ux/b5/zw5gZuiCZXj
NNeopv9X9EgU8unGtPErFpLt9RIl+mN4Y0YND05BtBygxOUv/71r704WvZAcwJ7lbjkOlZV42Mk9
zn1SE5w6nyztWssbgYuugXIgKFA55RI3t/qRUK8PVMYxmIQtwNxH7jCEvHYW6f/KcONmoS5rvxxM
b1XsPLfuy79nuO2HKjYe5PGxJPmZ7W1hi/K/wT0NAG4oCa+g2PCO4CB0mUFGOre5Rpxm5z+24HY5
ADOlIFgEJTK/3GFT8S67AT8VDMHEorFdJ7baP2KhNDYBTipeitZD+48P0e/KerOmfNW+ESJQXfs+
E8FBaH9L22Q92e6kzOw3RsdVSjbDltRk9NR8EBc9HVDfm7a5mC0FsmY1YLajb2ZKWLf0C3Ksl0/2
X8YHps+yhC7SfY5lYtXK3g1FERlpuoTZf8ZaWxlxme9avGTfWP4llU7EJL0jzTJlSEoKW4Uq7A5z
EoePnny8Gb6TcHrShI5dR2le6pL+YSRcF4b/qZh8GqMfjKsgbXQ465ODqN8ymmbGIPuaZw+WmZS3
/Q0QXw74lecaqKpUGq+n2FZSfdhXRb8THjygCXThlchm9fCKyVomx2ou8XWPpnm4FhsscuovHaSg
zGgwFlJvxVrUxrqMRTx9fxiGzXy7cFzv0aTIAeIvq3s+QMRKz8zOFzuVW16mqzos14se7FHXuPQz
BL7O4iPGCzqIvKDLwcDf7DYfB1aenXjhj/SWoppLc03tr3Yq5aHqUjc7npynDcD46GKUhSgdlYR6
7YWqXZXykfcpOjbQ3EcaTKj8VVKh4+ktFfTgz05I2KYi5qzCDHQZYr8uUDQNgJ687Zk4+QP/+ngv
6pEkq2WC5TGuZ5nB6anlYeoNUVtwGQ9Y30gQtEp8bLbkCqtVg4wWksZ8/jZUeN0MiM9sPtNg4qeU
iVhVPVy0/0/VStSpgvHjjSGCBKqVe/2rCgWSxmcV87+L7MIgo+OmRNaRKK2mH8Hpab5czdg7+8uO
sW+628kaqD/IsxQgo27eYW0gNlOL068aspLulqVx2nDfRRAurdS+fnR1NiTtDrOzqV+m3In6/jv/
ie17JQQgspysktuEf9ctUy0BHLokt7SoXAtf6rJK0V/sX+mNoAKIS+6tsWRTxoeXplI2GqgTkytM
oBHFcFIksSTzKP9siiM+fpPlGcH49Y2FxcIgPgcpNMM+LuavOEoWlvKjptfVhLt2KXAU9OYjb2AD
bbXnYJqCTpKdpazrWx50m4JUjvnSSPwaGJ2oEZXEUjSwEcdEVR9HpQpuCJBFrOEuZEAHeLAbag52
t8b15Kwm20eVD/xPOYMSZnfl/P2NVekIm3d+YkoU9JneKWaVCYgoRmH1j3a6xUq6oXeEtURIiTbp
mOS/I/siaLb1YgsL6Xi4F2rcsb11wKSosoDZXA/jz29uxp4uSqhfZWmRwATC+decUVvXaPC3V6Ir
6djP8zwXLz8o147Dvk1vbrSwuQF2c1muZm87++4YjMFmR3AbxGlQCQxsczQ9fhAEFeYBUOVoQChE
RWdni7GeNP+93CTf7/yOoSQ/YCNzvZ2r344W3w5f0e63AgzXzIGTuTKPZ6/7MjgrhqNR7osaG1yT
CpBqF2d6ZPf2VimRFys5ag1i1Vr9rDsOP9yH8nTnkpmJyDBDfzpkA2kLaZWdYG7L/M0lk3t/lIHU
2MutyqsllfmicrWnTqFjIYlkacvoQecX9qjdW/vQZQ/1ThlXq0PJEXsD5pkypMnJam/cgsweQqd9
8A/zYF2OQP2zna7eYlsGvSv2htz8BDysSc6aCgxjtslLHKZ5F632Kr6SoamHTCYso2B6cfTEexdA
f2XBJNb05ev4f5aiBPfrnhFa9FmsELkyR+1houYxQ6G0EThYKrbCgxaFQlSPuDvrgn867AaPJikG
xZcRAhKU/cB2FJqKcldKzltO68tYxgdQOMkbssrMLRRX6bjQTmNgmJSqQ0D0OC2W99/J47qw43aN
4/+ysQDV8Gem/9dqwd5TtiwWimPoVJmuTE2Ry7qduMVtCKAdaC4HY18Z9qdm9hMtmB3opMHBNAyM
761tlHMl0DxPSj9Sif/69bQn+8Bl7E4e7ki1/v0VER+dA4LGOyIMiCinoCN7mi6z4hguon4toeD2
n4PCpqrTfwAtGsnma5G4uPTJjXBJ2te4PPBsZG6tEwjwkO/xyH13JQE1X2VJIiwP9eTja6M8pqiR
7zx8qml3Tt+9WoFm5mQoQvXOHfZ6bih0XbdhgEMkIGfAxbRtlvLZRxO138JG8yEptmQvWlXkPMvZ
w5j2bAo1FqKqkr2RqdobcgBrhjmYIfT8Mw95f2MSau8+1vdcVJaSKXbri0fAqLMIMAkSKppJTs2P
XgCbIJbeAbyhm8FOxttQVvfWpuqpnS5E+syG4b5AVnXnof0t9FLet5nxVx6+Mv77yh0pK3yaw1S5
oQn1A1naZ8eRjRFVt4ZRcxQ/tWLEKadpGHEkpwZyBtLLUeEIbYnBlPXYgw6Dgle+fhonkdLjbKwJ
RRmY/2Tp+vD9HM/J9stlZdIDjZERn9fQ8p0z4bYgg8s4JykHilJTkLYF1eTYD0d3WkdBmkaiLse6
SnCzeRC9NeAJLuo7No80+ymEzFgNuNp16Bq0HANyFUK7ETMGMRm1Yh0t0+ifbhG3HZhtNbwCBUSW
KqkhxYty4EeYn7pjTTDPCN/rzAlOk0V5YU6gcs7PspYDkcgGnyCPaBdIHTankL+G2PgM8j4Cno0G
P8fqpMF6cqk41F+RhjUjLq8qLDpL2+WOPdgjkI1OydxBj8M4CQ0TqLnCqkML0aZMW09yrNLOLp+7
XjnwDWNRRjwvg5lYKSfC9/yXjSDyt25q/YX0xMxXmHTxMokRuoHkTDcN113+HiiA3vx2i0BzNgZ4
B7Fqlob8ju8eTsT/ALrEueVGs6l94IbT1qJLSX1QJEEay+GyN/meLI4AeHWCT6KRkU4Jh+ybHi+2
pcB/livhnLyqx0+qxMFKn3HP0D7vd5BSzj3qmSfTusQ3wcxS6HzSp8YNOXu7YGv5HmcHu3btWNv2
Hm3G5DyvO1S+sKjGXWZGvrMfssQv12x32CMuNTiTyCA1HnZew+/Gz+5RPnEwNEkhgDV2blrJihv+
2xEja0s/3/+CrorG/rpK28wnmNi17x1RaxH05BNLOZqQ+ZcjxejhjYi/fjyEeXUvbAQpqRXn168e
1POrivmtwR/kROFqWHkumR6DKJT0QUXnMGCAiA1nsKEea6sf7CzEi2xFf7M0ZMA6KC/ZY81iwr9P
VmK2Qt4gIg8vdz3YQDFnsHWmoDgHyZW7RNwy8QOB3hIP936+S4Yfkfoh8YP69UuHfgDEqyykKOK2
LrxETmM1nk/IoaWtS8W9nGqqmOrjLrwqL5YYW9X6/5UtKR6boNlvW0TU7XIPOCsIYFox2BNlOiGb
JpYB9Q4mgc5AodwOGc5068cCTRj6l0hBmxIwxhJ1g4iVI1m6evPlZXEzqe1jux/4QAcn+BWxvdwr
OMwSkFANrQO6ec9m79XaFND1JlzT5F2wBBbwFLiFYCFOYSrGGo4TyhXmZjBVCmRTe5ZcLPLlF8U8
frCnG2WJkqXV5FmcRLplNA3qp3jvdtf6hzwYZKrxepG0amIMx+azT4swChNx8Z42JfJFfIqgO2OP
DHpVrBN2JB+Lib5RgDfS9Zl8lgcdnZMFNtOTTIWSgyHW2SoFJDmX9i7FjdTE+N4oAh/qdJCFUU1t
1AByfiEa7l7dYqtwob16SDwsWT3uYNxyD6RxU5tUjSRSNspRjIOA8VdrHEXBHF+5xPSJIKKJMVtZ
4T2nHE4pbfXcm1sCRjYj9HlZZ+zyQXaJVzbnFxEcuuCSckoL0IEiBa+2qZv0RPK2Gfyj8oBkk6qN
FD/iFtezxKrZWp7ajuMnwlI2D1n93ch9o8Q4uq1+TU8mYjlKRFynuByImpBvyHklkVC7Pz9y5RFF
rIw13tUHP1vLCe9d92I0yhOg7JpGjQBaDEIxLMdpqu48o8pCz3gsSIR+c8QVkuph/wEpIphN0PkS
KPZ8SH5v0/T4hU+/3C9Avr8GjVc7RdB+q1W+mhReCgSwTgtHcQA7GOz18fTkp0ECjyEzL2JVu/wk
2UNaO7Kxk/+LjBEJ8A4pRlwpCQCjfBOT13JFNswEUDNkPnW67NJSxp17kf3zD+xu8HLRRnPjdYaD
y0c+7htWWFNj85AUetYzta6RZmAkE3/r5mEVDkTnFxPooh8cAffF6yPaTxu+YjpL5S/2WhIPEMW/
7REsZSYFoObjn7Ua7Hp9+E9iphrBz1XUKobnsSc35cbXhXF+++wYy3AGeTWOGsRtKmXdZ5dSL213
FC/VsPE5mgtdrJEUfIM0oNDwXJRHqknBIJP+vvKgTfEgLB1hGD9HeLSWSJjZw4x6uVdTSJUARqiI
ntneOuAkVygScw55w3MJIUrax433AThjqL8Y2g6eLtdY9Rq0SXRbh6H9AnnfO5wJen3Vj1j2vZCY
PmbhWSUPnsKf9LlZPKvAHR8HIcedWw3Bvgg4vq8kCOxWVu0b6sezQw0BGA2mOJWnGssllTG1WVvT
8AH6sYSDXc6uKh98NOB3xV7eYXCC7qRy9heB8QJQ9I8GHH4jrVGzfI1hiROG/Pd0kP3ZhmWw1rZ2
NLskN8aH0cmtRsN2JxdwjdEQqVXOAk4rQf+5eCHS5Tw81Xid9bLRAbJ//gutMKSKZlirbKrQo56M
w1xhdWSI0Fp4nUzjAFuPW3PjzxS336Tdk+HoPVgHW3SufUJlxT92KnuPcCCxfPA3F4KOyRrtpD/Y
UC7KHalzTPPIGNKGaumv596cW0iRdw+PU0shbjNvgtrRtKPp6hTm+4pCP0wiHz1bwW+oW+I2vKyE
o0rf3jNgc/eiTFude+IE1DSLaWtc3sCJRT1nZB7efatbgomKRRBAkoo7wzMHwgYQd4pcMregxHKX
nWVUYzGMv/drtem5qFyn9yku1+kXgJulzIlyIfeiK+zxHzJXCOuI1ZT8tgEcERkS8Q4yaS8Pp9m/
dYEXlkStFuERAqTR5zMhbepdEGDN8w7GjQ4iUVpJI2L7bU4t9Vi8GObOAwG2BnB0Yie6OkT+vkaL
qDm23ySKlYOX/VEtu7j0IWt8L8enmaKjwEfchDeKWNoMkTx2puZvYeTxALUeCqTh/hfkjV87KCbv
sEgxp4yG14ucychDYVV97ery/RLX6I5yLuiJN8Itc/80s/E7nbhN2iSA3FPkoS3iQbwnAYRqhRWe
F/irSN8SFKI7LbnFQHsWqRVlmk42W3ne8OIrdfg0zDgIpwXjZf1NoGRR3i8AVlo1rajE/dOhhd/t
sh5kmN1vf6yFM2S8o10APLsnsQnb3m8TTHN6YFm6uN2qmKIeT+zN1jPcZENvPxvW7Z/Giw6EvOm1
ySuCM/3QEj8u7/dQ8Ij+O2DY+/tg2qBzNoHkyivyuoHJoWFktS/cJWqdyvkQMK/G3uMotwJVM/NE
Pq0yIorkBhwbqo33CaSrLSYZpN+aGLin+giTf9tvykCudgigPqG5G8pZDHsMHPZjpI7JriShMMPB
Su3LSzJWjGEUCyyNcOm0KstJvIrRBfxPnaJn14Zdxi+MG650N7TCXbejP+bQfz48+bAK4W7zDU/7
NdevsN03t6hGmYrp8oVD+AnRF3f4datSsjf5EuTzqYvIKTlc+CnFRZCD1f9I7awTvoA/YoK23fNl
Cp/bbVvdFrHfKiqi/2Fp9cLO728vkdo7A+cr3bJc0jbEj8tylf6s9am6BtjI9X7RcTC78RR/OJw0
WUbhZVyN6TSr8mqqTtUcXZH8CX9SzPmIEHZqJhuGU9Y/2Wk4ci/Jkxt53ebrxWWpgalcPEtbaS+K
d2QPocbNw7AlYWZ+KCx2zhGBQUFIW7v+sRqHjWkCx3jyIiLMNnRdPRYVt0LjB5hoPGrEVHvBs7i1
aXCZSfY24ShHiQFcgmGnBOOYsunrxGNajbcUJcvESeqWUsvy7/uzelQHJzyj4kbRYv/1KC/lDQXJ
bSTAQVOE344c9QPFhoj10I74tKes/PBkTUQ65cKKbc2JDFC9ek7e65nP7Fv9sIYdakT+T+Y/pm5A
qSbHdveq0HYHYqZxdYNd1eVqqF4sbT1bJ+eewLWok9MuSD0B0XNwIH2blNwazAEVWfpX0p+9ghFp
4k0VksYF8taj1hlPCX/ICzw3mwuJZD7KhN1pbxmCyUUUlGZhTqkyLnxvD4yc7eGY9ImG+N1NKdch
nTea4n1OAviLJBSVqNM3RU9F0/QqEoZYbGpP1ZUscbYva9QS7K5QIzzOYakr9hRHzu45RshVfVpD
0lgUVSGEKw8sEGglWAYli9dUr2F1++aziAvsRjR5z8OqSyWzks/o/vUE2bNeO8R4W58yCvRT+IJK
o7Vkyq2qboWpMffRympzQFwXmmMDrBBBAQA5S7uKbd1U81y8g7RRH8T05NTAHjM0n8lkrydjP9Ns
tezn0b0qqmH5A+lG0pXgWXrY4ChKda5UVxxjaQYU7vTbGIUIXAREVSk3KkAMgtv6xz2tjx0yAsN/
wQHiCv5AoqXifogCDdbxmdAgopo6fngaZ2EtnN4qzqy4nzTJDEDv0pVxm5e7C7jqioqn6WsF1lh8
sFAWVn9xDg6yWTrIjbS+/ztcjU2tnye/NcjKHekXzpoXiKYWVDzwOFZ3DWaoyl8XO/2S2tWf3eKl
2/zEnYth99xaWHr0QPGzZSNa+XG6W3ow1vWlwG2TW6UXxmDB0fMUVyaz727HSGYzPuU3ypSXV/Gx
o21ES9OW9rP3PU6uJazZBBDds6t1JXj/TgzsXGdkQM4jWmjzuO95tFSkJEn3igZZOyM4C8nKwh+Q
naLCBROuhV/az9N1BJfA2b1S41sjR5j8ExxSI4U7n013Kg/eZPgAygUGGEnsY7NtxFV71vuu37Bw
7o3/kGEgHmmMa+qxLUeJ2P58s63rP0XOpHE3fJBew+oTz66ke6ajr5x0YyWAJa302VIo19Vd2OGX
LblemuAV5JRvSh74VVSK0yiQIrrlCYWk6ZaAp2d70rl17YPS+wFW7vfXWI1mcdGXQb+uRfhaW0Z8
zO+JIShYWv7CiVvjlWm67tpEcVrqvCpbHV5GRFbC1lLf+h0+ug7pKzWuuOf4L3Q3iEywmAEzwEyJ
E7ZwtDTa00k4E/nL58j73j4OSdOu/CR6OUyUrQVPixZhY8Th2Pmg7hjTvZF+s0wpUL9OGScDk7sG
H8B1eGcC50sF7s4abNecLvXbfQewzKQdj/cjlT2C86p1pVpu+4h1khwLQD51qoZ3797ApaHDvkiZ
tZtJ67MV3CnbR8L9fBctkzPGySbbJBtLVRY0LLqi0IfcRo61DjEqPyJU937m25A21nYmMn21sYGl
FzGdV4k2L9iJIPnCxodcNYuUKDA9/rqe7clHVtiCGqauGLSMYvZiW/LWU0zSKNIM8uaWj9moBzkd
W6377O5UOjwwHqDRgU5YwnSLBpgoS2uXGk7pDNyTv57LCVfr4YGETLqIAcRDZ+3j2DCaJyenDaUo
dKdIcGCG1E9vzj/k+SevaAc/A/WQVW2qu1V4ZYSeuY2WvZnF7dbNeu5VD7VaRytFi70Ev3lLO3lW
OMnvytqEZiDI0L5DUW3ZiKhvBe58dZtuQUFlGMy7Cf/zwz6tFTqr9LTfb0UTCWu6QECY9IxT1jfI
+DcuxVpaPJOjoWQx73mNkbKU+DgonCsiE/7S/Xom32srj5G+c79cGqoii5nO/O0Dh95LppLTJDkt
ScjdB92Zj4ngOpkeaToMHXju66b0OR7BOhE4/iPVai1R0m9iBYBSf+Yvgr9lJ6Vyrbzau4bXdgWH
QiLsElk2EIgkZpasdFTNu2lHYvk7nedGADcmyryxjNJR3vTJcPc1wFDR/OEEVuhLbYg2gJdgk7qG
hKO9ugdh1/Ncg0tBw428OUJrR3QhEh1e8Nu0nv7kXERRrsgI9Wpqh9HlE8eaMU+esx6pOxf8x/aA
qHDZFCXA1IP4c/r00ZzxaIgFZPkbLrSJn5ukbDnVeN6HL6x8uuh78nJpd3kwds2HsIW40BvUuH4M
LCA2FGWoT5HM861n3q9DAVU3GonFSGZH2bLfG/iz22IiyZtRwVRpSwWdNL5VGO0PeVuqzL3yB/dA
6yg+qSjLtN9PEG6BDSc8Rw2CTEppP0RGykCmxBjSS4vzXgF7GvNTQtyHXPtkQNUDiNu8jsHibvgM
RR1OjihKTIkBr3p7YDVtkcN9oa1ALeA/RGa+y/8wdqxWHiVST4kbj+l0xtKROayfGQDKSO99VrWa
2HfOXZmVKdqpNBXnVXBeY7numDasdWfa3S1kcZJSkNgOjeL+WeXxRP561Q3sQL/nBQouR/mIfPd9
dtr1Q7EpJ08MFUv8HQYzj3xMnV5ncWSnKzc8AmaAQ65U1LXkqgygnOkaJgghVPiIyjNW3SuZRGYs
jZJKfhxry+dUIQK/mlk4GHLx8ROYn1BLxypssTiAPyjmqzLgRO9XV9p6Hro7GKdJgr/6U1TiUQR3
WOm3U2rK9HAWNQwByb15K/ZTTZ2JpUmfycFJAOyiES3EJcSyFPKXnXEhg7CciYUXlsdM22Bc7Yuj
TmjoEwdl3MRjic18KQOsSr6cOqgijlx6K5lTHNq4VKWCqUIXL/d46qtDos/79H2J5aFdAqjvzIGn
PvwOZ2cktUbjXm+UqvbZ/mXLvdWN1YFS2j9lzg9+ElEqQJJFdLksrsfEl6PTIevvh0sE2HNQF6DO
h/KiDg+/xwtrmP6W2dF9Br3IZ0UnbXEj38LL24NGetr6wvTQhYYK/GZfoDbx3S19llPGbd8QS5m3
dmAbcsBDZhut1eDBarKMptvDsQC9xsknOYtzucHClkAv+S2QPV3VVlT0XxDQBi6Md2SLyV8GsK4j
OdUJb+LP+vkM/0cZs0ow+DEzGk3xmnBZJgA9tvlO2II5UUVdFqeUBXqfsaXhZo3HaKvzUBuYKTDQ
2eoRl5ihOgQbbXoDTTo8YGwFzNK8TJ91xemgLshP2+UmOphbDhi/oSHtvcgq68tdI5RwRgtQWqYQ
Z/b8XEqfJ6IXPSyEIutgqGFLLJsUecTF8ToZ0gULdSWStrjgyIzEDFlyffIPd1ScuGSqC3gouaCU
JJuSSINVXbaiLKcKefH8v0ipEMEDZ91V95FhEzaZLzyvYogqm+ujAVzwt/hlb4e+/CFPt9N14k+Y
p1Lb4yaYdMq6ccVBCAYjSPhrZ/o/BDE+tAts9LwiVOLo6e6uMxXxscvCU4etX+FXBOfhMGtyVTBz
8pXSZggMGKqzvGpUzyXME6slnMuVjO9EHYzDyVou9CtD3WZHvVNAzskqgUX09JGO0gUVeS9DUQsf
goDvDDrLQUTu16PKpvvXVzVRdhGKerPgu/XW0c9sDlijf+hssAAsqoxWZBRwwmooCucq8tmSveXN
jIDjTWVCcxwEsOnDhfrSWh0kd2hY2rjLfmLiOXxHuSB5LwXbDv9/FQ3DnuTaJDvPiOwUT3ChCw26
eXWuuAcL5EBz2+Ry4nwGbbE17xP/jSaiVi7fGlK6yOXQUpRrUhMg3xCkadMOfKM7tWyPmoIOsl/E
elc2JTUT2DAqhix0oQijn7dqi0qWBsevsKukrgH9Seqb4i9zv3ncZgvHKbip2IDD5gBPvlGeMiK8
RcYJ/MA38sAO+FpxoiCdIA/XA4b9I0r9deOR5YL7PbHL+kk84xSmKirAH3ldcgMR+W+vbxqWiKsT
3tuMqrG/fEeS9Ee3Otr1Z6T50Fupg2fA6y1zjvhuvSwfkpUxMRez4FxYGOhVNFEC79bWJ8fhudUI
7YllbRhXtLM/ddX+DwgfJhQ7oRG82oF5O032Hl7jM1fGZMLaPZ46ZS5bkHMS6uohA8J71tl/np/4
WfkZv/iY/Rjd7Yd6M4Kxe+Tj5rWRi3fKNL1DyvaL+wwXfHAnCP+84go+RLWu5axqawhiqaHxb8Hx
nRYYUg040RQ7FpdWfRtKl+/yCJ7GmSRKsiH43EaspKDa1Q0ycc6yZdjblRtwPWJd/HTltQBHHPDf
BJ1yJW6TPffy+jAgUm2An9ODiBIdCpVNdDSCwoK+rekigZaM9QCZatfWG4NgUnNZt2vGMjWF+anC
igDxGuB/989giMPzau5ac5WlpckBvi66HKW5W3Kg7BeedmYJgEm8ACpFSl7h2/f2JGINh+75svZu
PQFZ+D5Jcw5LysTDOkpCne86gib8LZV8BKEFVhueATRC78PKMvO3mKI93dXDJ4wsssR3R6xzcPA3
gbzVfuaZgtC5gbOszdpdigNVOhAZbgghcTx11QEjMNVqmUmEoEv+XjLuWR0H8oT6/5nad4U2uCHl
TzCdB07s9nPFpIqDoxJzWRgS+pkhf6us6KTFJcp4bKMaKjrtsVQQlWc46xmAFKcF34c7DiwVcjWh
CM+vPIvoxWzN3uswd0hwDXsr3ZaQ0CEt+YjvDHB+hpamfuzr1sJ34s+ZyzcBmwTjOF6sG54fzTex
qwjObXR7BaydkseB/9JyBFrqM36kvjhFOn4WuKHwMB+g/ygUnTNbs090WM/Pm23fH2e12KziTXvK
TpJurgwqd4J4e1ZHCQuWIukYPyelh/UymyKiovVK4krc461E+Qre4W5uWQ/ZiWZD8/ePIZysSlub
YO9QShdivfQdN40dMlccQjg1IAZitP4YMs5LYch7lc3oFC19kjp5bqYNy5Nc5PKJBZS0R1uOS+bx
UT9U2RumSZXpo8j8OEq+2qh0fK4zPKMX+0jxqbOCC9KJ5wdKJlYvVnGfm5lOoqaixo+oDMSRMWvc
894uupl0hb+Fro+l1Y4L4WPgALKliVBXLFLaXkU1Zm/C8VRMiZJR6rVYaXDhdPZ1FKMYcqRoXmMC
UyCncioOK/iw+k6m+DoSXonLIRtPemTKrG6dz+KPqMARkXjOkNuTU/ivo5z87ZChOg2g36bVzlh7
lzFW3pkH9HD8iqWScopAaJqZ3Ww9i9eXXixNEzkncJPwG0q3fVt2ISk5vkmxdNk8aTaytSybopQI
y4Oo+ZrNfYh7LCUnJaoo0wILGGZvqdOrHvaSqFg7aoem5fci0X2jPLtkyZ8Se/RVPDvVG25E5JDX
TCgbXgOrCvIPtnbQ5OHSb+y9GgCs+FLpka/hQenUmQSqVXMntCknydYk6GKM4VH6q4SYgE737CZl
dA7Y1J/q/9hVV2D28ySdXX4FTQd5Q6PEZCUo0GGPMfofYXNb9RT8tFFgTKdKcbrStEFHN8pA+kre
NSzsFqjSyzGBe/TNQIkXgMzKA6tlE7XuWCi0l1uB5AC5RT/dh7R9rLhqEH5LTK4NP3x/Xf6I2Ge9
YHrKcnr9jfTyp5fU33K3jbL0XB2/ZrtmWsKOeCQCG2KJTq2gzgsBxpq7vyFFN8HC861PedIj3Ca6
1MNXHoWa3gHD/tgy1AoLIveSv5fj9/rk+Zb2N0dncG1rs+QB05EKFEqXKvG6oKuNcjf9ShI8olCu
d7pKA2B2e5NDByJBjPV/F1QiEEX2JVQI6n2n9LqZS7nQL5jUejxupD3Fq0R+paZgzjFi1Vt4wpZk
z/d8WXEew0Sj7iYqQ/o1WVWQe+/gbzGSbR7Vof+dz2rz/R11pUR+jfN24uNBsEpibfxXnQ6uLhka
pdSa3B+400T59MfwsRKqUqOrNPQdJ7WB3rwpMUxBqtGxX3mirRz++hIYlWAnYEI7TLLSKe7/Dr3T
zcZ3EuqnR1TrnvefH/NNU3DV/B+EH11seD0zO8tSySACphOhazDV/rXCAU9qbIp1QLo+uCLckfIA
LPrMzEUDTBhQr30WsB1ohT7JYrQHr/uiIOIvBN6ii+gCxmq95fzY7bAHcqxbUO66Pn8RaqfSvxET
OpRxEvq3OVb2XNpZDLQOD+woUqvt8fLEjnmXpghKnR40EqbgGzqImpCBNWI0vnIMajqBnRCKOMO1
EEZtPo0D1CizGn7QzAipcNQyVMnpMlV+7rLNMKNLCDlKk6BXTPftrOP67X5ObIieVfSIgRBBEkNU
i13m2HoKWE1CQrFKuCKGKwksIVqtMG+jxegiKawMIMVgpE+SsEIgaK8BeNqyNrVkH6vEoIUf3i1m
Xme8Tj68yRjXaSSDYhyk7uTcEy0SLivLDwUiHjkqVQW1GZP7rxXPi1Fz2iO6vXx/KyqeaqmnS2bY
55zs1lpB3Shu/URM5snUIpEJYaPprlKy5dk46etF8PFbBxq/ILd7ZHkjQK9AArerztBLEQiLfbvU
EloMEfd3UwfDpu3DoDlrbnuBKTmr59XNrIY84ouMGoiZM8onDHxc2CfY3MUxAzwDhPqY+OvOtQlC
YDk43EhEzt7gyBAXDKUnDQ/3G2ouYdsgEe46BL+eTBSDXgXgJhttW214RK2OrLg44luTi22HjDSd
vJcL39LIZiF2LVXlf4HNBf6L445eZBlXTj/LvIGQDKNc/YH41PJnbOcPuMEL2nUynO5rknBj1ylp
d3Y5vQgxl6nnueCTNgQAdQ6Qonqm/hj0shPWBcEzG+O6E+UbVkihti65WV3CdiK7QI2lohiw5UKt
0j13dO6YCtxCd+MS832YAo02O8Negxd7EmXtOiMpTx49zNKsOfqGJj+0/8k8WsDs+64ZwkkzdrZu
EjzmFZcrvEe2TGREd2vyGkBsrRXFKSxzq7UK9obemQzH/bmJnOnWmt7Z1syFTzNSeoLr1OniwR9S
c44L5a55iExTFRB/Q2fGVfIkCnvn83Pjvckytu195yxUFtVWAd6rMDV+qGWfR5LxJsz/mjmw/087
FtuamEGawXLj704IPmwERGblPe54eaVeb7x9wzd0uhsRXLmErfa+H5mg8edwsTLaMVdCJ1dzJi9q
ZTgLrUEkLsttsRVJzFsIoLUxZlvsln+aQ7S0wIlVmYZLW2kP5jwtPDI8eLvKBlWje4DL4ZuP1mI2
zueTJDTMLpUQN+RRq7LbPdN0JKzqDluUuIVtYGFLFZZGSfgyxbs3PIv+CVpCbpOFp8eohqH5HptF
7SkNNTijCbT2xYCaGKVzugjzxuqJZLiuugh2nLD7uENAnR9e0xeIF6ggjEJQeoAIqNPIIvwkDf8Q
lUW7nirIssWwXrYKp6717KPnQ1IARY4yUJ2jP/NmEzYjKO1Z9LPo3X47gR05um1Mt1J2lUdZt5cK
UKa2AGC3mQoQ4GBWR7ViSJOsdmLPC19WLlcRzuYuWUdKfyRhlVCfPHN81ByHNcXK7ZnsJEUGa+Cg
NBWCZvCkI5ImEM8iVnhjQEQZmNOgXCiaG8mZeSSbH4UUan025O6F7dzrTVr/DTs0h+gSWMq2x/4g
9LMqBemzugNfrPvbAzo8G3skyKBSedbXs91Vr56bpl/6XgP8f+mvuMstgAhmdHG9g1aeo6dWnxbt
V6R4eWgBl7elOcDGpg+DtDaxGkNtSMv8eWfwjlbqztyn34LEHsJq6pZ/jfANSLb+U4A1ol34iFPz
qU+/ii3mNt9XCopzuSf1h2p0M5nCPNIqnVzDNukmBkk9dS6rrD27JUXKDE3Ps3YJmgkLdeS5ZeE0
An7vIdr9pa9yLCsP2VSoBM7MnT1rhnUNtEknC3aH8wXoPX2+ZhXL/Q2KHwxvjdykbNNQ/tnwr3nF
4AFvNC5YJrrDSBjubKNKe9Ojih8ARW2OCyud0LxLLY6ONitWs8MSHDYowfFNDU3VbQGYGG19gyKO
PZkEJ5RnhFkjwvuQFpDZ7px2Wi5zAiLIQu/dq/eFcYADw4Yniy/hdHlRB5RkDKnN/ji77I9mCONq
m1LI+Beh36tUg+bc3WmBkDAhHuzOFwYlIRp2JdnBYoSzpAWKHgFqWbAtZhH9tpZDS3eBeEDhxSRk
6RP5K4AfC+aoz7ucY4dMDqAOfoSCoBc5oFiudjDXaszsHDC5Gdi3PySPtrmjgmKNA5hNhJ2gGgMU
9VFIXxEOzJwRyOeymXVaOpUc4JFRlu+O0N0wnisRu21nc9i2kyi4j935BgzW224a2AVQbiUX+s3a
/dJQPKSMnzxRBlrQ9pllTlFdJsWvTb2dwQgv5ISxbSYjSHWrcB+ZHrjTLClyBHoj6WgDD8VJbKHy
P9DmLWuIGmkIcOfczaUG0L4JTUfuelfMgvhfjNfWI87mz6zRn0TEn3CLEc7aKc3wB42KtMClsvcF
Lk/xHVs6OynUHcArEZ4MKa1slo4XLWhBW3wWe6SQ6nbv6HQk3KxOPHR/W991BB8sQ+kh3PTxb/vX
teH+EJVDfyKjpeTLVZn9Q5rRXQg4jGbtcYXY8mqDs1IYqUJZzf9og7hcpU3X4GszBwS7iBYFEfOX
wOY+y2RPbz6LpwPfJHU5iZ17N/L6zYBm3YZQ4+Y7IyH0W+nNuyYOGyYlPBcPHAYzRB+pxAY6f+ak
JiPnvmejHZwZNU8iZ8ptwq6HR+T8UGsRs2vaURResvJzxp3/JhghQMRXjbBoFSJsVv303oo6N4mc
MYo5SGLoYGTZXQ/ds0ncJz+JqZ6/Ob5o+dk6r4Q7fq6bEF+LlvXJoMe+cQgYqFU7YiDgnpeNG6l0
EYvbsuoKC8AjLT6hLwIk0AvUdsP4GzSiR9v/x3NPatGLbQrBGo2NUb4/qj2PPxq1rutj8VVgc52x
dG7Gt804QW1aDb5tG+F9U8pvmpSxklI9Z6HHIuaRe5ap8rtW1B8Zjoim8IS16JKz4d8MqNxHlI+R
g0f9AJ6YZ/oliSTIbgHHpBSVqo/YgMud/0OzrwBhLXfWaGElhpsGETsvIVk0NFgMwyiYeIyowX6n
lgsnq0qzX2h7kJsbH5MuZYd4hCvP5Vb5dDyV/fYjWD5V7xcjycIPNO7PDcQkaKt3sEvOFjW82OhQ
70KFKpSWCP4gQyj6BFGbut6tnMg+erN1hU4DGfA42A/Q12C6T5VAPdycx2cxke1y4N6LGpRFzXSs
ncSKeiwmDp/OS/7aLbB2CFX1PXYTGJstsw6bFEz0+2OX6djzV8cXpNbRrfaEoquuxrbJBq65Help
IXxNe+hSSH1p1HehXTNmTPOil2gd4zWMiHR6fPhNS79PFkrzWtmpug4GtNX7jEojGGYdGcw5kJhI
pO4VmsIqq5vO1KIHLrNXGjf537BQhcvp9al8Iqvy9zrJcMZ8hJpEv0Bk/6M0cdQZgqfNjNZWFzQX
pqkTnmqMX4j08ZdoKxnB9WHMiWyGWOcWh/0B+LOXw43mk546y6CEJd5qlkkxzAGsODiQ73OAiGE4
hpN+t8bSMEX+qvw0aPLsZdoitVR2uKM9kROFRpjr7C8TRh9HMssOh152QIEZoKoLllNJMeVeV0wB
PJTHDtnihrnu7vb3Rh8KaKu1r9jvuYPDyqdazKMibjKHMZ2aBCkXCQL8wWvbCNTjr94Cn37ck+J2
Jq3RGkILQ+1p/P0jNmbn7HGxyWGPt9NClJjVk08xuPPhjd3jJDzF0BBgrjyEBgHyiJh0mQ9xNqva
6t0bC+oTfSETgBh6k41Q/yk6K6kgnNZRTpqTOroxbrbTdTjZ0WRaHDpAL4k3hiF6oOGmG36YOHIM
Io53mQ31ss5n9MIj0dcYdkTjkaPZtUFqr1JqYOYziBpiJyFNnX+lInDTH2npbz/+ASE4dd3EJe61
GOGzgQgOEiIJNFn05PhXU3svvnhryhRytTX7k/OQrCosKQlN4scBqt3Krl7x3+Hbn3BtL2K9Hte1
sCP+QESIwSKTZJvJKHJJa167ZIqAYo9zhwvJ5Dlr93Wucxyh89VujfrNHlw7We1X2u2WOmYEa97B
CBy56AcqBE4oNaq/vhTyPjkvGzu3DFXlimju3de/L5O4S4sj48bnwtvCOMdORrAugKdVDudWGhXY
jHHEHG2lRCzomNP3CL9i4mrjYlRwroB67LL3310XflDf65vpgSjtv34KRg8rko524UoY2n63CDQQ
EBWNGGWTh7k5k8EVEb5s/8oLUSSErF1K8eoCX/NaNvLPVwkhBu7hQXVpdfpCn/GsLUGRNzi0P13X
eyMzxYGfuaeUY0pgaGauisHeefeFjIAjhaSVFxMi5wBHy3pWwOgmJXpi+OZUC06fL4kUWpAogjJQ
8daQ4TTOptDV4KwBdNxlDq40VLmyy5mexsRGCxXTpV8CA7ZJssvhwDfAUQaQzNxTGOms9DkuTOfP
7YGzaBN6ckb4QYNMAFpPkiIn47SqajpwRdlS1aimx6KXCH4viEu64tYiV5wuaqHBrr43yTpB3lq9
uYx4vX4m2mz/xYfZj1JUdO2s1rYxzfZUipsVOKIPsvBDTKmysfIPj91PC0ubUMwiK1fxQa3fNlbN
xyISJIjHaw+vHWbJtnEiIQlnhW4VKlUY7RvIJPL2QPrJq4WiTdKXTJ8bwLbIjEIAdBVqpD1nQliI
s0Cuc1jpdkb6mgWlXEo8bMcKwOojNEKqJFSc0mJcZLBvtQhZzcb2dlE2Y2nvHpICwnxeh7veDtJu
YKgqV+YPjvBcaFQbu4UMRhgwlJo4rVOFrssGLVW1uIj8aZ52/2rItncxHZS53ZV/9hTl4Jjusala
WZ8SXgXsV1XPuGKixOf83ks5MGxM6k2VJrpcwOTFT670nouEwfT33LfPUfMJmItXoEHD0waWf/rd
KyNvFdXqz8apBot+sGwJZwz7Pf+NogDYTZaY+7pbTRTxby6T91LtJ4xdiwBZS6wAhv08tn0k42ML
R5Uu+Uqcj3L3MMTEZlAJvJ0xQl1Ed6VHjAM0gYGS4QYGs1N1jDpsPrPCkhbw0meDuLBvt49BsZJK
5JE4X/pZmuxS+Megu0CWhrtgI0bwCtSPAjcWXtdjQ1wDsupCYsV6tRS3KFE1WOq5jLjaNwRZm9v+
A+7y3XjXQSpyFHOZarx8zGQyp9j2Zt403zNPBHQp9Z1I7Lcr+paK3CcUGe0nOZZwuXIBp6T3bVqF
7PFphMAiuNT8JC61K193H5rZkOMWNybtViKZd3lDzVWxZnl2AXtA0KTfP3OGqqnnmBgZzduEVEBE
6zp3RJ+nQ4/OQp2SSAyEYvDOuHIx6t1PO/ogIMNbNhsUTPCa64dYA4dq9+woWRAXE6zk+F1Tm8CZ
9VU2pqMTjq33zlDyFG2subQpLAjVsJr7q6r7HvF/Sq4Xjt0Aoftmu5OFdvo17ljeX0PngCOx8UUI
ZiA74XMYWc79ACTC5YYlCNdh96HjCGudiDcvvripKgrWfeVcmW6Mt2579F18QgEGWkCEZ/RkDTRr
JFZyKZasR5vCr75uKZs5Qq02eCYY7GeRSid06HSd4DOTeMOilgx5Pu3jU2aaBhvD4K+oVk+GteAK
B50fQ7os9DcWh5SWSo1yaWSJmiFQZk87CpMVoWZz4r/UAC78Nd+1UZDjAIrVB/Y3AWU+CP0C6Fyc
nUz9qCV8OHaCu8KdIua/vMyHOu7ZJ/R/YCvyMaaaLE1mU7XY+1QLbx1eLwzc4R+NeHD19Yqx8LZ/
h+2zf+NNSQwPvEWu0MwqPpMgp2y3VmSxKi39bsR9enbi4qPdYIPcAEsMGoCaHvshd6dZFwzT/chJ
pxHFEkquUshQIxW+4R7goVyT6AHHogNx42RFdK8yEBWnM/TP1Vg0Jz4SqnxfNT66NBq69LyZq+8q
PqsRTPZ5a4JJrz0FVOxLloDrbheB6SwihbNP8b8d6dn/gzp1xT92Mtmde7gOIWeQ0S+lXsGUj/Bg
SckeDuE+0oZYTt8d5efNE+KJP76B7ktD/xrZ8sk3UVA2gxot8swZ+vXXCpjq2PjvdkgZae+zOzC1
X+pLfvXr9q3O8AdSIqi2H3h1iCBQ7wZfQ0Ts3waSHLf2ojwLmoGGvISMiR7jIn7D0/rRX1gWdNMF
Ux446FfiMoXUol213FCkjPt05F9U8Z9IbWk9F2JSuot40cLvSR+aA7JeIjYgslcH3eNx5TGlU1HQ
odf2eI9GQdkoL6J2ScS0L7a36Lnx9vbZSixMnOHvKLTKV7uerIZGVH5+B7hIRhSu/IxXWiWOJt0b
NXdWuC2Q/e7rP9Ag/QisMGt91WXyzToF6lkcHlCeLMkjH2wi90GHzVJSWjfcrDhVzlECBomwtLED
EeDBI8VB9vSJ5PXRzUKd5hQjUkqOmwXGTYWwODvgMQcQ3VwVzbB/LvXyVmC9q+1gy2aRnoGwvO/p
wCOYFRviRD2VoFmHYmXQk8n+zXyTf+JNNfbgdktxwHI7LrNgEm0r28CDJrAVd6g7hbiHHgDfoS7T
evuEQyu3eFPqVVcwTDqwaVnKi3j5hN1ASV3VIfB7jblUoVabjZ4zTJHC9WDdoY985gXj+N02ZqIW
bMJNBqVkNPxT1qxYy2C72Uv0IHIrDtFejDv3gvdyErf4ath+pXJGSIXHvuJaHEdBd1XU9adr/T3L
UJ9/cu7PszQGyrpPm/tl+AVHUQqwL9yfbVkx71wo0o0aMgYM8MUrMmzgZK0+WKm9K9wcCxRKHVL+
HxGMXYSl3MtnDfkdVfcJIUmFwokn4BRq8coljgiymi6zJ61X7CMFqk9Bq5wXbXFFklPE9Yn7boPJ
j3+PcKtHiXXcvoTX4weTTH9mKp135KQAng9Gn/PMvJij2JAaHgA1K1xJ+oRICul2xziYDsPsR4AY
ct0RPvJgZTt4ztMf4yxB7h0rOrb/zKExC6uQ7cqmGe/GWbbCKvu3awNK7las3g3JXhqP7XSFC6vf
nvtV37a/z5sYI0kiXWQze1Zl5RS3THpsawGxKj2+IB5SvCZ5nBnH+53TBxj0g2JHMPLNcRJalEt6
eKNrskNlW1q8hol7YYLWslkYx/FrJ2tsrZcnXaK/f1ozBpODoqa8JM787H6LWXPPbpFwvvD8AvZg
K0jPqcqsoXJXU3Vuo8LiNoQ4WLuhIVQGd55dLnKxjwGsOiXkqqIqn0/VhfGbscCgo5Q4pBld06Dl
jHidfKLqhun21pn5xxUspTbKokS2B413xZR4mdL3NkIm4dEIh0JUUzWexkz64UN/dt4Nw8rVG/kT
rOdfO2mHSpOl9ALRNMnEbE4OwzDFvZaecJc18d/0D81T197/NVKw9LrVpw+Hp/ZsWf+dN3n6kPNE
iDWDX2W5m8uVlc8xaQQ5JfW4CPpy8bWRs8Xf0+71bE0vpYpu61AnKJN8szcQ8s7yIXfgDm9aNvae
talSRCaU1dCPkjHkWE9c9e7+qCxA+BoDJef4i2pyER+nTRdMDf4Iv4zzLnkQGVk2y/z3E26mf6HU
c/Ci4c6QJwPFcMAcQDkTtI4aSPLvLG3f7QOZ5ry0IwLG4ycWL2RqcMKn82RhhNV2M/Rl0avGcSBE
GLD3+pHW0JvEJTmXf4X+pRzpmuFR+dKAB/UfEvR1owbppq2QWojXzlXPfxI2b7i6suAo+l0xrZVl
1JuvuwELmqATQSkD47Db3/YwvLy6BjUhLLEAzO7NRAA9dRnx4ETehbgNPj8nWHqvOv7zUEtV3uHb
o1If0Qjea8OPGtVZDdAaDDXZSjqr7p1Wsm9mUSJ6I3zO794XlX1qCVJK1RGRcJtaOlVc/wEacR4c
m9gz/o7jD+H+YYwiS2s3Rf4NCqrCWiWTAuY4sYzNeZfaJvp5lNLUcJ3LeKd0yB4zDAA2Bg+IDO/i
Fvu7OzoCP031SCbUtZmJU38hYqzE4CORGGoEK8tMI1PBlV2OMSKQ1bec2KEc9hJfSMjSUJqe9nvx
HtUusOYSEwbNJmePRSsp9R6dhYml4LM23SexfCf+QloU+2ZQ3Pcq3PEI//nKlIFqWThrfTeOqwSw
Hf07fJ77BjLWGa5etTTT8mCvhYwhZpOY24QLW++mtToUC6mHxxKERlBrvnzDibsm9HdvR9OxAhDe
KgvU4xLuT0FxmMdSuCejuBZbk1FC+U1RXe9GT6akA3SPCo2UHy0juxt8kQmwnHp1D27k26w+Bb+H
DHBr/TiqKJ5rIan207L4rNTZBBfz8KrwKjZB1camVuizIG0m1/xsaHBsW4RgeeY+XINx05KikV3k
poqueVpAcjcHIjV0iQy2ZCrevpcg6CHa9qRtAkI1YOKGjt/+CbWQQXz9tmNR/f56M50rtbp4utWW
fm4CjNGjT5jKc2VxAVwZoGKtcpXjfRazm7BGceVC46ht8f7fnTw6pDpWG4XPVtkzzD+YkztYerBq
4Tbxo+82w43MN+LDY//Jb4wdZ6Sh5SnjTwd2KU/YDCg8a6Qb1myWcLEc9lXzCfTnbIkYNwZD6laz
4Ikm+6UuwVjcYIQ5a4pfgtdRVuwvDoYFIsSi7i/dfAO6/4RNx67fgVa1aJ4T4MVR4HMT9763Sgk0
CFxAUUmMtm/CP34MqCJjoeu8cv/JAPc1S8hZvRQrV6yAJJI53OPWTUOC8/51IWCg8izlsxhxTjrE
1mBZ3XrXnl0ns6zkZ8sPRNZ/eN6+tCXMDHSuODvlmNEJ9Adac7KHQgkCDMrBM7TyCw3+oJPjXOvC
LQ1Xbo3jW3lvYd31f+fKlsXHuoqZZWZwAVfJA3isBZJm4D7tXJw7wFQcWcTUDFMCglBuKM4Kr/wI
gIBFungU6BY06cQIXtCXznKAm0mdGd8qfVBdnF4wYGQKDGGYwAG5hC4RMNp4uFH/feAlP46O766x
5iVedu/4OmVithSwzZqZuK5XTTnvOKL5/AKnyuWAK7yPIg65y3ACzGcx4oU59tPx6nbo0lnHCY39
NXAjY/uOcd5dv2STqKkD77rP8/tiX6UYcMOxQ5WAtlrwOiS6UzsiFOkf0C10cVres2xX2TcbBVSv
gRJhx8slB02702S4neMSIHrCQ+BGRx7IOH0bgnod64cMWBb2wLJqkATKkEKRhTDFuZjnqtCIqXUI
LFxzm18sEhQMKs8yvzfD56EEzK7iXsc1H4xWw2AFwik/exp/lnsMPWI05IQMva152HG/ysLpDpI7
8eV0bDo7HQr/mDLME7OXHPSpOTeJ3inIp/CcRRxw+rHs4MoyHsMOx2QZtyGHg6k5rZaEA4scpsqN
ZHTStPNEiMYGIxk3t7ylthrORnRW26KyX6VExwAIoeOKUqZemaZtE/lS57w0TuYzZgNnX5A1zWgi
1T/zoNTdsMgz5z6R8TLmxv8wn+rOUEEQXDwqGoXUP8sjNPG7dwUNN/Wq+Ih7PqJ9bNDAH58fRkvb
o1WceYO2h86Q3R7p746Qs2/vxeii+x/yYCwh8CwZ6Q5uukisgN9r45lvPVQ1HKTOcAmyELqfyNOk
lE0eXMcPLNy3Eu6VbF1sp5BjODJI3503sr/MMRueU0pO5YoUts6XrJPfJh2hJQbx49eHgKPJKqww
f8mnMz89Gczykn/Uoki/XYKY5gbhpojyHNt+3dFh2lLS/2KxRL2srK1UsVJ68SkwISc3a9NRNpYp
73JVh0V+O1GjADQFGa1EHf2x77lKsLNabNFfHcf65JtcsS9Sq8Q/aoICia0rAnig4lNc7KokiXjK
ENHEFaa1fBGh0zhw+uVxODDSrCUUsgQ21JQriHeJXjkqXSSax8QMGohNt+f5C6Ql/sF68B8A99HP
FJLBSZhmE891as3j+5FemPIE08AvbrnUXSW3qC/VISUeiGjYHXkZ3vn6dkn9H2bq9J4Gf/EdLDBj
4DOkIOHe35WLc4Nj4gXsTvL/f/jVfHAIGRTE+5m5twyKIyzJUCHABeYBGRy92tI6niIf4RcNO5Ym
KGIg6+LaBcf5L2Q6/Dk5W7jYZGyEA3uUr6IfdYKC6WycZ2d4XKB5E21Ru+/W/wNXM4wsGqG4Daft
T4Ui8BTntV9+VcNWOaie0+MaSMvPJgWketLdQaVQkv4GlX2s0qQ4shm7m/+MYTcVmhxSwxQS2Dn6
fLGsbxQULnSx4G4vnIGs9vfT9+wyjrmKjRa5g2E9o8MXK7sQ+Szz5ELorEdsmp+zjuw8KLKw1IvI
gFRG7tWT8sQlmAKRk5geTXSzNE6slevrpPN7xARRF9eRcIAi3WiUo75HMKrN3UbUI9BTHqQZDN/z
vfL850r9jRdGPzAPANShT5q+PJXra1WahVOvp7bzsEOmNmDf+FFYRhBWKb9Qu1p6MhUzTDrmI0Tf
r57cFIfHYbvMxrnMouQ1AlU0AFI+iLA85y7gXH3qhlNlDMBbz35C452mLo0YCgeDns8IjOMyBkZT
4lqJFVUORh03xKA24dfPMiFomkuGXJbrD0KKmh3umTNmYT9KoSH9411ABK5Yw1CYEO/9y+CRZjSR
NzSe5t87UYOsBgj/qzCTkfGwCuGTBnE2YNMiDKhyF34iHu2p+5yrlG0Qrfl4LeS8SGd1gKFiYHhr
1sj7arrjQ/lELpoXi1RieNcWHayGzw7+Y2aBAnpej8NYL1A6Fhtfgkv3eXx6t30f+MTnrWyEUX64
lYZyZZ0H+MUOdZ76DvhEdFqnD6VmitROpfGVxouG3TH2IB+2IXbxGLGXEgYUeGY1X6LTkX6Mf9oM
kOuzaHUZwiCPOa8qkf029X+zc5mOqXis3fWx1qyFLbsL6KEXXyfsuHbSVXKa3gP5JuNFOquZ/EVV
AbbnZUb623IKhnTFz96Eql0T8Q0Qk41+qPicxaewP9oMaCHek6wmvZgkybmc19PWe2cu1+HNH8dQ
ulxtTioKSnIY7ggBsFhHR9CXtmzfGYOQAV89+VII6m4bVpisVRShLWSerQG9OKK8xEq/mjknCaUV
aCBH4+xoFbDAq1WrWO7nzx8ugk+EMWK71iCeEavTDQhxzDIEmMytpEhrMg4Xw+WQQtiMzpDJ6zCJ
c48qMQ9iHtQieXYlxoDRIEmbX18XghfDwoDPhGvgY/gS5kigkmRypr3NqKQ706JIrb5W0q4fa64Q
Ul+mGqJKPlJ9su9DQB8rrNFa+QZFcdG2pcp+meV4jLTPOP9rKja7ajG0SqQBW2ln8SwL92fd/Qn+
/Zekgzwavy7fluydKn5QcMZHUpTH7S96U/BL8CvSp96sIFxodWsXS3ZfjYUoRmzdTNSeA/R2hbcn
IyPneWf0u5YUvXLR6QgmSQkIdXamfEvvfeECqkChSYc/hX0b7hujLTFfe4YI1/7n+0Rjy5BMhPWK
p/YJMfqrOhuHAjw8I2aNLLA1gIUjdCRRl83q6gJyDt6CSlCpbrYLPF7i3Vb6zDb52YWsRNy/rNyO
9JObxNUglTupIZ7taazTR/KzuWstDi6kXLePPmv74IR9vuaP1LWbfMi7yDu/WpiBivDQkvJsr3yX
Cw+kYyhKzRSkVZLybbLiXriR1+3b0f2HW6K1DgSbPZ1aBY0LBNu4yR20mOkakZulxPCErpd61ia4
8R//8zNv19K8GrYZQGcC9Cji1bQcseoCEbsJGhSeByfz4yx8dGaoGINGDQUDzokCrefyGfvI70Ki
uaiQQUTcE8MD8sM/IsqlbFaDBrddMkzEcuNY+ei3DIPm7uT8lc//r/mbqPZRIfRtJx3es/c8rE9f
YBEFXV+BJVcWXescfGiLlmZfFH9BuHGzk4etGjQDNvcD+25HbpwPCBRccLzJT7pMAM4tr+ON148i
8jGmcovXRp7IfV6h1HbbgeWXZkUqvyasLfE4TWyLY9xehkxd9lm9EuItSbFN9N2m3lJc1uNcEbR3
avcYGkEB3FtK6HEOFzngBCwly/0c16QRkgji/1TyY89mtEzmls+aGBoEtIj1B+MsVrTfKVLXuCM+
EaDjiBGlVEDbwxCO3dPX5UyEQg2bqTuoUehB9bAw5n9UnV3ZuBKdXpxUeCoxv+9tgLekob0KMIQN
lqQRgwCG/+XaN81QVIXf5QaP6pNAYgfB46CMbhH3zplxFCQ6MceSmJHxcTXOBrJTuDdXi2XfdZCL
dfU1a59xXJKMlW20M8gv2bvtLeCKXkRdWED0qcPEO/BkR4vPMXnWl369Ssr/yRcB3phNxxrXKz6O
o0wvxJEOoRBapwDTcdD8ruFuxC6StKhPAtAukzsnxVZtwoc+Vl9NcQmNUBxi+XhDyRyulWx5D82/
QFcv+trIDPJc3G+S0fDSNGnTCdp2iJ/DE9oiGpwtxBw1p7Damn9tH/qrzcbNKGH9YKLcjw70gwfM
XRR/qnMC3dkeQajUsCum7a1w49168kT8Ko0UGyE94SxwwAdwqZxNMWyxw8Gmt8lg91w8Qw3N1psP
xfjJkwTk/eZMH3VWXgstdAzgr3r20GZ7S03f77ujAzfFN+0tbxCgxd2BpuuvZ6J/3GdgNkWhlTuK
B83Y5M3q/IDilLQbfNcgf593HLfePbOiLiBSk1+Hk98Rsabykr5W4VfAavmp8JPnCTXItLgIVUue
feaAt78NBuorQw2FMwzoPNAO3jigsJ7sHHlZg90qUxlNeyJ3pQHST1F/aeOJyilmBI5zfQdpZ923
Y3R+yLB+J9NDa5qLqAyBSTLWCb10BMg/ZnAKt0tH/zE+wccTnaeFKDMw9cnI7NXxYFuSvusEKFqP
t5uLCqF+SmtxXJ6KnMhs4sRjXUwk0UIzBLtYRHrQdAOcxBPNfJPX2WMvlHN+DFrSQaS+8Hxzsbvp
1P41lNh6FF1/riThn30F0lyWllayOaNbHAoEFJULOmlVcFKJV3Pm+tFQA9T/Utwd0ZtMavzqgCId
nQqERZHaMWbV59V8lhM7jaLjPEO1shDBamdGcYzWR4bbptZAKlDweBWEVja0Fmbr982FVWdd33BV
ID96dkpeb2Me75QS24DNj/eh+BYtO4uJfsJz305QMgV9v+OZxbfKTKuaov6ISTMybaDs97wuBC2D
E7BPxNHCptYGyNY2RGzG4xVJwgJ+6Az2dSxjvcT7oPFWdzy+zjN0cBGfxySo1dZNe5mvexzI20wX
/NPtP4P7Vc+WAJfXbEPAhPt9v/kvh4SyaQpz04uCK1shPnyNrWaZzSwVBcxL9kzXQG5rk+x+ouOf
gfcmKswFiQxcB7J8AljmsjYUw6u9ns2E1tcRtYu9Id8b6nq+cu86OO8JbJW3YDE8as8MXksYhkyV
RhiWZten4sOqufGpiyuCGB4FIQQXbYXq64hXLKkGi4OOce03Pxrmyi+2zNVqmGZsgn35CSmngK2z
6Yn6JvG/vR14eTg/77oH+hYW+muceY/miZUk8DyjGvJzN8et6OGte4+q918bGtTnVEyEZxcxN/pY
+/RhacfYsNmX8IWr7QAU5eoE7gnB0cOS3sEQXgcmTRcOLQQz7PZH3l7wU3dkTfb9UdlEeSjqSc38
wb2r9Ya6Z8okqy/Zz5Eq0XnePHHEAI0jdgI5Z593upvufwtWEmOtL71d6cSkJ8712DvYLwHpSF0Y
1a4c63O/Wj5YUFPaoXe8mk5MhvfpjvHn0P+7nBqh/E39qpzYRWD7n+mnw6mKKlIQ7y7cUdIoL2cB
iDZ9M0CjplJugKdK+PJGbbcs2kn7bD4SbcDTt4/KmH3u/8EQXn7HBtxjnfrs9PHz7qXB57adnWob
62OaeriwJcZXupqiZA8hdo3O2lVhJPcuPaWTAv3qbk66bF/o5nlyb6qjmov/yxfFjtZEkZ9USdul
eNCbQlFsrVxxRwvRbiYNk2YXRGJi1cDpEFiRgLbCu1NAYmmDUHGS9wxgfosRU/C7vUp0Hn6qfzKJ
8U6ss4tmUD3vTGEsSkkI5pQNV5w5EQ8UJ2ujvr59h98MKK/Em1mwV20SC6AGL0+w8HbjPQE7nqzx
XSN3kVHwP9nDVbjgiKldap6qxZiTWikn1dXWGMHJg34CY7pePPQ3pc1Ksn7j9ZRaI4kHpn8TKHAd
JfCYTY7XubeOblY9txCGNR50CqAI3pkxf3u+cy8IjrZ1vtXdS+83d6nCAgkkw7uhNJqcSARep4+B
t+jXVBMTuLOhtXh8EqRn8TUpzx2NlMAgdnMULIjVkr4TuOvbg5oetMF1ElDvpqLgVTjceidNdHsR
EQlsoqlsCx9T2pVRC5iX3G41fUzLb9mrBJuvkjGfwySzy0MQDdMO4Z/X4UmqujCUWTixjErl6hP7
XwJmzkUPHtPu+bFD00WXW7XS4MaMg9ELS64UgaT1kXC2xGLXC9jpDy2mryRZRWRYabMnWIxE2ANu
3sEwZkewBW7nPFPy7pTO5rVRTCdCLMhm3wTLBaNF7fZPIILnv46isH3zjiDpXYgn3qe2/3Sur1dx
Iabc83Mf7T1gXPo/lVRHmTT0ojr5muq4+A2sMjK6nYFZrqKGvsvingR8HaE8eJ9Ga+dChRT5BU/X
MFyNeI+UJZu+BFMCBq+KBeXBkk/xUyIRy6EUWPmLOoHL9v037qlVwMCBgNLjLN0gpTOwD8OS8Ru8
AUFYJA0yeCOyxjZoNumpjYCrBzDpQyc373rKLZPxcfrJCMYE6iOBMsI/P1yX4GBuZoydX5efNaH0
wb17XsFnHFvGIhWkorJ2jI0lFQQV5XfqMr2B7KX4oZKil0jT5hvBW8RMJ3EJfWV3jajWvxvZrAPm
1WEsYkVIx8PhJw2s7gUcdjerUncdqRIN9fcH1t0miwgSVVAdsw1U3N7pJtKuejmQdNPngxwa/pzm
BmbootBPw++GuPUp5wytpEYIXPLu/5tlB6cHmBVii0MfBlmP4MuXgy5nF+icH3FVmxNsMFoUo3KA
Wr3U20v+GenbbBmHOncLTD9V3USpF0LJ/5pYx3Geu426onLFU2vfHEG25zFtUve/chIOIGCvvZVM
/eNy/A6bMz18YXz0U55yao/fpvEwdwaXTImc9pl39ChpS7F+/YnLee0Rv0WOcrojj0ZmnroLKdOS
Z81m1VDQQeyghTaiEZDhMdX8s0Cs0Tq3eoLGKFS4CD6arSaaDT2zjzI3ToCKhwdz83qbqHteCovf
d2ovEZPNUg0qNqyPgW7j9VtuE/nb1A1lAL5M7H/BYoKL0lZHvHX2vNLhFLaeFigMmEZngQkA8gE4
xNzzPxFOBDtrWvabMOYqoS2HK65+Y9WbbRLUKBxK8keHu5OkP+ch958+15WAmBfvazPXqgj2ZCmR
7l21yxUjvz8SO1nYqa3ZkTke5S4Hi+aIaeqYRODUEXCBT1ZTsYU1Nuvt9kKx7yUzfyuWzregTwCf
LI9cxEgPFHqV4alAa2/aQ0LSw81ZfA+Q7osQn+AvIa6CpDyughlLCzxTwkdU1Q+s+ZS1k2d4DSy5
+axXNXkzQqVoCIoWKyDxO9Qlc3z/2QChimil1N4FJff77MyjlPytvSJJ8yZeUoyoAX84K8UsTF46
8lXjGhyheVKONNp6K8sWLAeVrso5V/B/+1sy/x/Ps7TPx7d1cBMPbV98dLM2BP0O9C4dHTEKZVcM
sc17b+DIGGvCUHhEpVWvUo2QTaS7Ex0MHgTwREnmCKSqGdR1Z42ydMcdZqUDcKorsR26eNYQfZC/
UjOYquStaI69YBH+456OIeO3NHJNOnKzrLMfneA+Zu7zDM1mxA61bjhMlN3vhBD52sOF6qiwOIGp
nzDtwSbyWpM2ZRf116VMcrESRt+iOmZqlwDb9CPgAjQI4WeeEnqOut8HfigNdQa5oGdLMpihQJmn
6ayKC7Su4UllXlEK1WMSxVVnC4dRAFE+eZdQWT3Cvq2dCFrv9M6Hl0EUTg+kVKyd9RtQxCsBnviU
9j1Yg2YaB22iymuD4YWTcE4NkG4O5cVeRq/g6lj1ugo+JQl5lJIawYfDvTTC9cZ3Hcb2CZOcdMQx
+y8R+O6YsjKvi5tR1nN/EHhIScvuWuDQzS8Mf12YbP5ZhU0bb/t8ZDk1lCEOflEDAzYs6brXVJKA
U200SIpzoBtC/nfR/P7na3Ef8lJ7a0wULGDXoGapKZy0jMV4057tZH+EMJaraELXYvyL99cW+zbd
fmG9FIDIy3pjAyLbEo+eGRzd/debl242wx6oU9myKDzXgUasl7UCrFSyhcZwR8bn03NlleMeBu2b
4Y2SJdWMGX/TnGsM+KHYWWL5fLxM9+cBgklGe5l3aTSaLxWUtIE/KYSJQ3nl9Zh/yCGR2Kv+/ejc
4qiVDDE10aWqjKOdv1ZJPtepHSwusA9tkqBno3AI8JI/JA8les8EYdxMGYyoRNGsghsQYrQbMzDv
G03+Ag3OjmG2X+JgybVqvyDML/vU9raMa/nuvZvOx6OfST216D4cpIwKVxZ8Sg9fNj4GxMNYUWOP
hy77HuApX1TCw3auQ2g1W/GDcMpoyslnzQPYryDNV6rFG08fD45QLsMK0GZyJYOBhZbzFdoSbqUL
Z6kNS17wvNkmgvd9t1stTg6sTghuNdvC1ojj2uzVaOMc1SHxnTbFJ7aqJlsWccSByzONpX0VAwUN
sBy7S8FJhNCL+7tJ9N9+ISUUnEtmT3reYRnn9Du3YXufsknlPuOY6oN+BMBsmP6OqCCRAGoBtK/c
gMH+JrWbcjAQr6BnhSD/mwLspWMZTrXHBL07K1YaJrRIWCmltKGzzm6nmrQfDa/G5ecP7X2PNSvO
/SdSNKIEQkel/vU4dAldIjR5x889fjTXb2j4GeRW15E8pRfO9QwAqPPvbQPl+nVVGq4NcgabqQ19
/pUx96ESyvLBM1bcuLv24c16Mqmm0tSkjN14IWHR7OkN3v0U5WT+1U5xm5wUSLdPF2hsE+abikQP
vYchUxI/S7i+v+rvGNlQmWdk5nYrAKZmX+owduX32IXeGl8p1ombJTNkBSqWMbhXo6ytKmUulHAH
udHUMhgnE+/KPDErUog3rQkzLUeAed4Wj6PHMZdwWDwmmePDurWzi9OPSmsQT/jATJFVXVURxpaq
nG/9a/xQm1giSc3c+9/HVBMCMeHkCdYn4hEQ9JYYY1vWWAbIj1/PwiqXU3Nzmi2LNzF+imj+imJ6
JnWU0Sp/aQEu00dnIdjrrKhrulRHr6hUz48/ViC5vMetscpqS8ngMzc5XQ/UbbLGhFyY42eQsyzV
fRpLm9rPtts/ioVzFhvYHaVO9L+XpND3cpQbzx5TUgxWqgObwioDHjWhSnpzzMQMOxwfHspQCt59
VVlpjcR+dTIEVV+kc504EkNreFNr7WS6zLRv8parKVtnUnqOACgogAT44NMOMGYfGuKbISNgT3R5
cvbKOrHOvHfYufcg/6BLyB4KEPywqAfXD2FQGAwsVeShYyPFDg1G/saTqq/NPkmqNcYxZhsYZnuB
Vuc2QssNuQXh++RlVrEncp8u2iXX85P3aRh9FvhvhNtv8muBrFKxt6lrf8o7F7fl2jgC3T4ANw/r
9c7FqeJhL3+AjMNZjufDb6h1rI+PT9o4J1bi5SzS1mbtZ5Id1WkT1YRwRnXw81RzMPVFyLxJ2xx/
fcSPPUbeDfQx6d88lMlcrGc6VoBfbCa7JBVOdKd9Jy9jU+BLefYjb9oNo3Uh/ekLG3PieUyR/7+X
psKckc9o9WVAcE9QVbTMqCfEMuwRygUsRgBhcnHrHEI6cQKz87tFgyXz9lmQLOCHITD0AJsurP9x
0LAjrR1pf1Hj0qD6Xuy2BvWF9Eq1HpH4mFIXhCgPNdDo6yyNGrFWPcmNqP+oElttmtMw2BLyWmE4
R1PqL94Dtte5lU880e0DHc20//kMlVP1oZn2ojwLIiW0QgiTzI3y65KosCfJstjgqSXkdglpMK+e
O3jKPGSP83H/54NHndI+z+3kZ+VuVFI2bG+xuGBZsX9vrHscJT0aZbPwzRAd8Ykwv/+0IZSdJDoN
xuPgnMpIAjwhdJ5xqeBuu5AnK+hnpGtzYs7f/W05ZG6ncEkZVZZeTJt2K69xXSJ31FXLHX8cT04t
hGR+G11cCAC8qJlh3hzc3jWEuBOXURIhPKWNNYqiI8B5aaLnmY3s9OxRTigfQdI7iwOiyrHC2DEC
+q8kvVeNXgpWwv71hm9x1dCVQnsanPQk7T2IyS4fv4IKn+JGeYPZKpGXsFGEp/t2BTOAk3BYIEDA
3kN1g8cMsEBRp/2r/FoWGj0Z9ZSu4HGxsAFs84YWHvo+iF3Q3TkHyxOMUG1kUrLTQtgf/UNeiDkF
C+aT9tT7Z2kCcemkivToTvMcfXRPL3ftvBoqBaAVXmYHH6XpNOcooLlw2MdN5id8VepLneqzEzIv
oGT/O5xSPKoL9IN1S+hr3VGyYsuACvJ113g2/hYW9+Mba5vHNcV5zEUCXEtdpt5k82f879A0XOfm
CWwE7Z0EsEuuN2brO0GcMDMoD20rwqToUN8m7Ih9IWWzoVWp9vRkf2d92AVVoVA+AUuRSHvMg5aG
60YEptecgCMKYRGYPW0ZAxyBumUfpaOFp7nePltseG7sszb3c6nh72lVlza07vGGXYjL6vJLHzyE
in6X/LbzJAj27gjw7pdYW/Ix/NQWjOMkiuVWYwyeumCnADKUecOBxmlwxtSWmzdUEvxSOjcq2djI
C4y5sksoIfyMHXwsh4YhjDko2jfaNYUa1exMLO/KlEiaxiIV7z1Fha1oQ79EtHVzBRVxagOcCFXH
wrCgA8spSw96i63Iph0tjMTfuTrXbFjWGxsZzPrQGN4AhrxwYpSEULoioi6+0IX6fduu7LrVbUPg
J9qmUTnLNtDRldlivoyQj/wmowAWUDyAt/b/eDXvjIeMEtytPFz7tYj2ml19c31qNtYE9if9uzT2
P9G25JD5GTwNAlAXJwRMJxCDbu1/MpiA6hrC5iJXda/wDK3RbjO2punbnTdkpzNiElHGqKWWM0Np
hga32fSP9N+/9ZSUXA59tWtqaSjA2gVjEXFImJlLoZL5z4VzMqGXkr0wx0Tr9pcCYDmxo7AepyZ9
TDN5rYUSSKY6ICK+BAk2ZiJkFH5lejk5u1k3yI531Lu75AeCUui7o4ncKx2UsAfMwB0mYRLzaMAk
MQnyfaCdC9HXHTm96GHSe3qu0pRKQmqvgYb6YdjbjRzf/887rTWZGoKD0TdZ2ZHBMCM/LVxHgF4V
oylMz9frn2TxESZKvb+tEsznbzrt6X+gpEBIu/KL52NUnUIgXCy3XUn0wVcpgHcKIgLGFlmQ6Ihr
yNt+7YtBhpVqN4GfYLHcKbjTKetkkkcsO0eYcPIeBV2rzA5r3G2wJkNVZ0aKGtiUN4qFCpwvZ6Lm
8QQ+/eSkCuGNofYUqYqSf5k53mBVPB6elaEUmOuaIFtxU08czmSv8efSkXN5TMY/0MpHE04pkenb
liIZuPD+2sC9Ai0/OrifGrHcdmJlIeNsVAAv1n7vHED7Hwm9ZYerrvjDwr+58fu4i/zGeszNngkW
d2ZqqHBDJqaI78mdVPofZ5OLSdNKiju9qPvj1HbdHzpfg7Wb1ET8qaNPXoQKseimYZHJ9jaRuamA
4NQzpSvhGnbLaQQh6mqHhIeziXREmyVX7jSbqVeg3KVGoiKdqzCzIP5vBwzuCjngae8+QgbXCG3O
18R4WfQtctIlw2q72/VS5xCeOKXVzbypxCWZUvv7ajk2VNRlykUMBb52HOTgsavqyBgwPRDzeBO4
WpCD8hYrUiXC9Pw1HkVtBxid2emjkros9kge6oXHyCoZKOXsybmgK1nbUqqgeWA/uGdv4WlLqexa
2d/0233XGpjCucliPgvbrfKW8XgE21LVkDCnx2RUnSz9gElDIZsq5d5kRoXuN8D1/xKuxr36C2Fk
gZpI1qAqPxy0Q5pQsTyBADh+IxFSGD+/7sP907S+kIO5huVZGJuCEuSgllrpiEn5g060OOSDHWLX
L0Jlp5IB4s5sbCNXjys8uzmJLytKrP54ti2CTSw+06K/qIrNGAgq+DnhE5lyepDVIQwpwmfMDMC8
5ou53BKeDjsxgyMkpRWYj+eZA819/zyXWwlxFvgt0eWcsfu0GD2w30H7StCt0nL/+bcbAMVFrUtb
El0eRUWEJ1THlfISxvwm1jrKUWrhBpsi9kUDKsxtNBg+b/EQDK0JWzrWHYrbzN1bWRwD2iwnG6Fq
xlIyrHQvTxMyVVvFR9wUq1GkUoVK/wLHaVMGO6RALz/+TsoQE4x/eTCaoUxz8orzb3MNgUFdvi1S
VW+YS3szirxrKTzosj5YPgzvatCKfeKQQNsDevVftquB0+0vsp/t5ekoYtZtXQkMa/SDYrrX8mwj
M1vFVbwL1Z4ECHU3KT7/XEoOt7VVhkL2XGJyr/9HDPufl/WyHMy+JxGEdVAPz4N79dNTqXT+cMTJ
tU2SF5TE6QN/50/INQxptw0znr63kCcjdBOvtXWMyNBC8jFyrjkCzJIX3XNuAIJmeOfq6C0f7loQ
jSddRi+21S3lpGWlount8X5EnZBtob9wf/xF9cDl3ph4Mqf/5bb8tBAPGssrBQEd+52lHth4xBc9
1BaCsOdKRZFS82r03n1WGQoXC95Oo5bpQr5avXlXLuC1r5ETF88zS8QGsXZ7HwoM2qZGRWqQ8S2w
D+cJuaMtT3LBYfwO37R9k+sHCRqoCkvPVqxWMLtIiG8J8RY+5Ouw6DJP3JDGDEfnYF+d6R6BRaAH
Rq3FQRuc2isac821aHXapD8d8Yo2W1xDHyavnO5ZXCt4DvC4i/i3Sbk+gXHtL53JFmnEli8W8i4J
iVxNGMOXhNn8JBCzR1H6Szanr+8gh/QMq+ZPXzSNyprvzEaCpmf46+ocfWzIWia7oTOcUkq+QkL4
q6DLRkGbMTsbrmCOHX+ZSZqOBG2UmEWB3yipJs2c97MMPqLJBXRKv7WOAlTaCXczMtO1yvk5Ydoj
/sbqX395YGmB5xAKFav/RLWJv36aGm8oHZYFszeBIhXUJ/u9ckL6PHefeOD0JfKEagVtT+Q9jZcd
f+kej1TCCKPeqzSfoB2laKihzPSTFt79VHt+wuOtij1lxW1aSXmBiDX6X/gdqQGIz/VfoE9zqEF9
KZDcH/m5P3bF0WFZL8gqj8xKLXjdmvl/QKi320w0G+GMxjX3cDzTf8sMMTZYv/4OY9sDjQE3pfHj
L3DT9R2tSTygCGF83I5QgeDQtAMaHdM1a2G43BN8lFIQOaTtNReprFfsRiG+FUYqbRjPQNLS1xDP
3VcrrZW+foEm1olXTgGl2me3SPa3SFKbyytnCI3n4gOG8lRn5iCHiZc6DyXt3byPXCNd3EU+Ube5
LyL8FtZMpM5YdHZvLagVDxO0vfdxBFlEGKzuvBoVxClV/eYn3m5TSEmggfgnqxR+VRRuc58fUyV5
zRJtCpMAF1gApqQpLz7oODQbt4cPlFQvhqHk4HUUqMn3b7LT4yKVdTX8I/lxI5zdD/gptW3GKE+5
H2H6flauIuuQTjoLILpDnm3igTTkJiOM2+e/vD3TtZoR7l4M3ENztGR2aHKFnd3LhXhPFILZH/4b
pQoEj2gDGbmHFtD9P9kfrn59PUN0yy6FQHslXkyaKz6wvD4f5wxc2iRBa7nLPUiWgERYRRXD7URx
vOE90TsWTgLknA0MivAkQzgvD40q9BhJySIFWOwP/cmdtODHmhnjHt/GOcrIngYwCK7QrULgXaPO
eij2fjpjamypPVs6/5KD8WlEaxTyYOJ7J6EZ02WEtDc5TnNPP+pxLPSMdSIqczFs5EHTscz8kxaB
uBjkttyS+GCPGeED9kzEh/idYMZAzqF3kcBjXvPzUehDiBNaogYnnatJQb16cnnBWYuMIja/KfvS
Cz73JwbdmRZUDsHg6R0adicnno0eq+as59G9h7rCSARaPzsx0M4nK7L9bg+GTRCIa1FEKu3PSkR+
qrL3vV8ZZmFvV7hIPHucOd3azP/gz0sKSbAnVSNYNN/du4IyjrpYwrcrgIDX+u1/gJyDEp4Eyx1W
wVQLBE24ZnVwNa/RRhJM3tE992ugK9nGLluA4tXwQY4f6HxJxV04EmoTRG70XBLzx2IK6lbkFiFg
xK+FT3QIepkOFWT0BpparFlXhxPpopOC+2yFpF0WjVOxhGqFYmoThmhAXYT9dpaqeskkNgvjfMPs
1YcpkjLR+V1jvK1Svh43rWivlR/qmXz7+JqG9OiJ4+ONhct4X2sFlQcWN++WE83weAO/cRrFK02d
UuXf4nXXSR7IHlaz/kRttSz6S34FekzatWecXTGzdW4R4/kYLV7AJjtyHstaXADI0ZYVvH7ePstf
HUhIruGlP983J1M6n+r3b6kouf79zBiGMdXE/jAoZzCQVbGwzH6GsZD6GF/gEfvClwv8UX6ytTkt
e+gfP9KaUiMbhj7g168xBCLCJWwvESZAUW+6gIoWU1EYu5FZJzjPu15ZpjxWIpzwx+cGO9J7Pzp+
hBU0wqXrhkzPicGOPxopWUFCYY/6pNOIqYgIeQkv01aKiL8/AiC2v/nm2b4ABqOFoWakYMz2qMfL
E56LVQ+R/cWioM+ZhqZuOld16XVbgml+Y1ZjSVyoYFrmf0HuepI9XRAQj1OOoQxKlFzj50KaF4cZ
CNn7luRwl6K5GEHN4Wyw7n3DuvYItzOMCpDp4UMvYuGKIxbz3Bn/ydvXDToicrFpqLHDPaBiLGGt
6ywroGnH6UYo2/sr5yxgfqPDMALCZeHwYcqeSWojBegcrQd6/8II5w4l29X3Nt2KSXdkFiPIIuOH
XI2MrYJ0Kf3sYRuPJA/jl6MSAYkxyoUYVrl55WcubhhezQNNrLrYsb3ShXAZJ/aL9w48f8RGrYAM
R8CFASd8qLwVqNFVcq/VPUFvObfw4czygBBwhFeDMztqewjlYUFSddL9LB831n9L/XSfsYAdfLH1
HkxDU8QBxRsRzqRjWnExksGD2ZKbiqfhXkrT6JqgNkZfpN4FWGYB9ZeWHbBCS4rKHQsd7YdpERmU
X7hcDCrbjDpj41SrUKChMDM/PXHfBJytgCsf5frbzwyKpP1AnrAtyzwbHkjA67AxhX6KAyElk9KW
Rzi0I+d+OOFg17nY0SNEzV6v8SVgMpvNWiNknEkRyWFggCw+tBFMLNVryQyDf/6/f8ds9zfZ+UUX
+xYyUjmelm3F3Wd9vovHeEi7x/Devz7vqCo9Ryn+i8UkL53+QDzPjxgbuoVBB4Qh4/58xmpUAFkx
j7B+yHRGWFoYt+gwFpAmzOQHyretE1IVaR3QZZqsKcvdyetVFSJaxvsmQLD0LAevsiiulRLw3dWQ
Qq6QDnRhcgHT7/k+vHchqX6ZsMvirCzjU90RuuIZNe5a2aRvNvXB+nzD+slehvxM6FfbAhEPEuI7
//Dle9fryVhX6uyZOsA684NTM6ygqiV27x8jQsWqpD6gG6zoL41/4Oj9KOTr0ES9s8QTht1k04KC
yG/F2/4KD1VYr+KeiIJ0VXOZQKbwHt6jLA8phjN6zMZy4OSjSAnlZvWxlEn1+vO4nbjaRwOOBXlC
sYEgaXOc6Q+etGDNLE2f6W+PKdGBL3HJxqLuAOclS+gYuK0Kn53YWlCBk1OOwCFzxd9hpO/IkGte
/uIS4OQMfYwQ5uwTY+0cpWE5ny1UmY7l5jb3qocB3CVfsifIdWGxyP52wuzkyvbHOLo4mjWG8wPM
cidNnHozs4g80TAYPyiyX000MOCOqcCzVDm8g5M1obAVKoU4Pw4hEAkw2YHs5yzcupFgsLnrwCgz
LSf5VRLlfGx3MlcfdrdG5X0RCTeNhy5Wdk2rJRbJfV4a8yMagFHYwtUvw9LdpOQGTz+hyKZbqUK8
0NRUjBEOAxFH9q/G4m31KxWmaag3kPi33mgeJx6/1oBluY5B5oqJLjimLS4xyYkgXJqqB4rq6WYP
5X01r5xwpeLSx2egK490EKoer0T1qX/TwytfNxyEFoGo6cbcQOQ8cNP7fPdWoT8c/hrx0mSG/WR3
q5wPGRbE0iDEk0Dmo/1glymyJY6GTKeXLWi66BIRD+PzwzlBp+r+K9MIVjHMyrOWKHlwa8x7QRYt
f16CWvE78DhbimDtgKz8ya+B10go8gkISL+5L1XhtQXk0zYgodnJBUmRGr4A43qDuBAEDzExckDi
jN35vWTlwFF/XDFw9lI6apfNIAu8zl/dzQyimM1bc3AocVGr81oLr+Mbt87R1IgQ2KIzme3rk1Ok
i4rpTmQW1JCFqjVIQ9/kgZkWtcB4TXq915L9RT7Vc936GTNemzN6nee4ZLhQY2fbienSmmXvpkiP
6hTVBR9hzR/+sp1Ess6pTty3OYyY465aSkh45cpT5Ll9bSHDvMqij63UxOB+8WDqnRHXAGQQbRrF
F8dW3d4ul/LJbnYA6APbHHeKDLwB3tbjGPKMaPict8asTmW7qazprr8yBuY2X+1Jg0euyyaHa8+d
A1WQQT8yB+nD/7agGWPns4kG0pSQhiYgFmXBCptWj/1dCIgrHCSQ/fTwSfe7gjvu36P4wOQjeIud
9gQZ1SF1qqQ+JtmDKYDeEvZ10bSJ6/fDL2W2cOtBcpdjLYbyYwI1PlNKVJdBDR9m8zNbcHdph6SC
GvoEaz+TIw7KYE2ODQb36Y+MlI9xhLox/+uF4IMkRL0lKpbtb8TuRTS6iOIIWSDCdRjavh9LVPd8
YmRirb1SCQpyW1U17FZSf2w7BJsRMgaQdl6jBoB7MBNKyNj9CBKXgMx+fHOJVLHHTqgvbw7DMcUJ
CGxVHF9kN6lgEEfS7NqZJ1wKlnttrJj3QHvFXGVyaTjGqPE4NzATOYhHptLRr7hnt+qaQv4iybCe
bxHOZSkD/Mb5arKdLlrA6u8kQFtWQYD7bi1Z3QhVaRnQgcdT+Eu4fQXYJTWVUnXqXZEMFpbmKlSx
L46FZzooJYb1YbnDXSHtk8EDjAdEC1/ITaP3nPFc7jNoHzAAHt83qWRD83zFy5jMQ+Mlwa61c93h
cDlkzD7OiEir10QHMMxY9S8hXUfST+8K4uvEQO//QYAcL78I411a6F3kaTOmBIZMSqN+D9eU5p+J
TH7OU7pQ8C9T9B2ycngWp/rYveBXZiHU4m0yIEZlEQ68pLT02Sxowni1/TOCnIgvjvYT139iEo8I
8UOchpJTjLyBZjO7qT/QKairWkxwxIIy8HGm26KXCWaiYMcwdQXdoAXf/4HGDnJEfb0qhzvGJEe4
wZOgi0TklAS4exOMJFykyuF3XSk/er2RoqsoJ12SrALhGK7Jau3EiEP4VTQfEGqJulP+b+Nbm3Ks
Oz9U0EB5FDuWyCqoDpw+VwcIQ+KcDwYLqUH9E2JQn13KfEwmfnLkfZEPS1Cw+ipIOSko/lT5Ilpi
qfbFDWR5vXSKt4YhdudeX2PkCqXzxvEloeKQOdL2Hx2DgaDB27c0YYPlDTjYcaZJqC4rvbu1zbrC
2IIwy1jWXPJRafKAq9xqTqaj17ZtyeAKGC9UCiRH1rELKMUgwPulbJH8x5ASAsN3iLU6dq/BCmgy
m8So3aeo7782bCypF/cVGa1DP0uO9UKfidmgUpLmFVt6Dne0vN4mpRfgbBO519mM/vwO0uqgClQJ
Tnjr+jzthuixaD89ZXcuyzakYkQ2gvkud6jAF2YhCV/PZiRLM6634Xzix6B7m51TBspCLRZD+gIG
x+gnI2bJDR8DvPLFFL7rXiHZm32PP7zxDWoSXjiG77Rqd4Zd10lVV/2yhBRZGnoadm5fNqOJPshP
gE52Knj04JuwGks5Hgp9bNbpBfeNAZyddNFUNMhGx8cbnP9M4kwrQcABvaixaC8C2ohvxtW8heUn
4P7QDPMrRqXhX4FRhrHF44v7mDQXFq4aXD5MWo5quiLl2sWKu65tdWn2cMrdg4hDtn1Nl5nauv8Q
i+iDXlbTPxBfZ8oftXw9ItjZu3dwHOprYhOgjSKmySNflRJrSmtIBwKQ++9iQL9rGP8Mneliq41G
Ppi/ySd/sEFDI5AnqgLTmaO2VphlRKlGb/YjCiiF8lNjc/uD5KWCqUYM9D2oXG85uiIz/Db+dkyS
MEotlVzqDwv5BQuH8pUgeLvP/riYpPOahsmxdcrJatgNkgEBa3lZpxmXycGm/2ZXfKX41DX1WFV2
ExQmNVigdwQ8dvASaePpzD7qtAg63zaAqbDnYthySSHgb3i9CJfXKrW8N7hsuhisGFJVHOf4E9D3
BSM7CACqAsFz8r2Z5t9cMplF2IDRNRHIWEniYNfNjHC1m2inXG73i+WdJaqkq2rjJMGR5ymQXRAe
DJEhu/xTCU9sH9uEO1KPuEoT+cuvUg9j6pRyFbd2MsHaKQUOLQ554p0vu2yrccZADXmH0VnBejus
DTFhoa9U2JNVvJmGv72pqOp6LLHA8ywDuKDeSRTlF0geCGbJAvTR4IHc27uD+U7BnqGJ617kXV+U
PC0YHX5QDhHhWTM3/3RWzyA3oWJ6K5WiHOyDBFAtItt/MznJYTjGOIkyQ+UqVDzICP9BCM2W2g1U
JwWpr12HBJCKk7sJsjmLo56b7pZMBl6bjHWKFv0RwZHGyilBH82KHSudU9GyXhp6YeVn+F2K0iLD
yMR6z9mrb/v/L/TvLDy8I8iGuXu/R2Y+6iwGCRnTawwfA9SYXNE2rGeel8CK4pPUOLleuGkEX7TM
rC5zYnU/TZD0aZvv6/diKBQo/ULhagfLxDfRzVzsBQDpKXNUtpEecZ3OxSa/InlIjYJP+m7KqPO8
AGlZDKpbk7bRXUqPToh01Iyd60/c1aWKMExFuZkaNa40eHvKc1gZ/7FXDVfJEVrl3Ag1nUSRTT9y
5v9n7oXP/usyKI3EqvQLH2awEjOOjH/lvdUl4qtBJU63nnPa5bs14GWCMAZrmhqq7UGRIWBkuRCx
DnD+ffs/1ZoNJeP0XXZce1UdQ5LjFOzIobZv4553YMkgNksEDwGl6pL2C2g0KEXtgeYE3hxvxI4X
QcOs/onJEGwL2QXgmjZgg16TRLeI9QGaCtI2AH6xvbTS78IOAGgrgvIOfAbi1rqeYo5fXWrO57no
9FryULe+L17JiXsjDyKLk4wZ2T1/gBq3lWa+BW52sm1DY9dqmhmuyOz/JOE0bzB82lsC5L8dKRqB
uj6Mg3kHwMkaTJADvz33FWOVu8i9gWGEbgF66WNdtuy10ZZt2pkwIySUW+JoxxCl+YFBG0Tvru0r
cHjD5+LYb9X4UIzXtXaZDPDKYGMdSeVl8E1cRFm7EmUvnAvjKexO02I51nsu5aALvRv0CLUozlMF
MUTvJ197gJYCo3Ue6NlrcyORrCwLOgo1H1rSVYomKjd4LbdNhBd5i//likweOiABE90SxA9LJVPJ
5VVBgca/UWP8+DXzmILsxWwbHxV5PU5ZnCup/7NfhC57HMJL2FKMORzvAFnsAQ3doW/mTLIGWKzR
x5GWAuxr0LUi5IUvS7/2oKkhNL4QJd5hrgKMjIRoWH9vOGBNTde+H7+MfL2DU/H2wlA2/bZ2cHFe
lHzPOg2nmc6ZikDNCrWgcwpyH3jHFNRotjQJiNDWeV+2xv8Oly8c4NV4qXUpPzZ1sZi0ZTatTCP5
j/bReQ9LGMSHDymU9Oq8JEyStrG7EJCT1qOzQSPy/W+kD1sgITVcDMfYw0wb+Ku8mRvRFOYCbI7P
F/QL0piOepUKlTDvzP7hHV1cp4Gigwbw4HI6jWrcaNG++XqhrXiz4InRUna0eZJPKFp3/AsHD/Sx
cggjr3o9undPVgeoXuJovUvs3+8OjYOttBOjpMlRfT3W04BvTGos7FO84YZ0rNXXc1zFAPGhfUeN
zkbS/BCnhRslela1lupCuvuyTOUWCM/sy6C4qrrUnt0IAXRomtgSsRdBCbA1jtJs8heSkbmAYsYn
RwBFi0I1QznaPQEUB7SRTIpikvdEpi3lkqI5VqNKzcpmcAh54A/TFe5afbpkFVJlXfaj6ZAis58+
j3c1BK6nkJufrbh9qH8SymaACVvqxjnsaJl1VTFfPzy5dkh0nZYgSXSnH8vasUJK/k+CRI6VHc+2
5vL5mq5/O8yVLSTRo+YMjEKF5FZxTm4/YUWOmzup4veu2a7LQY2+K9WxTjlCHp+tI+3IoglDWtWe
5txj8g1gEnAO8eaJiVYpxden6k5W8qv/jqocRqbgWnnZr9GvKRPOqVtTBF9d4MJj9wwmbGcHdDWc
yUhFKamvfhB7AUSj4xder79hGcaY2nwTM0lqcEhejoFbGxKvZljkJIZZhB7Up+XyhWuTPp6qyTwe
Ipmp3SOrMXY20i0UxkAfCMn8WL6cAImrRzuNUvi/TzDZhkl9ilzvkaHuByO5D9kzV+koGSZPUfc1
96HSS/gvbTxG0zg4LcpHYR1d+E5fvnYLI9fAq9VCnaloOnAgE2rdoOG/+ziLcdTjkx5+he/vP1pK
d3oUtJyvFhFykffmmvNzs46G9yIOphv8cXQ7CNquVCNlhGjdv5lwcb4nw6jWKGlvEZA8Xy57aCUy
WkL96ywnkYbkB6a+Z1sppRig5dl2roWJJ7EsawzfewRywDLxON1DWwlWaJiC7vg3zKcGsOFwZKv9
glQAYHdQp8cLT/gheVB8zdBrlJOXjO5a5hXhtzz6ltPus1b3JxxceCgsCjoLcW9blCpEXDoFZ0it
CZLrbhxPSe8c8qGOZxwVpzEmxZOszVoLImH4LJ6SHCV5RvuTav+MVu9Q+PYdtNwz7XcKAExWdAeN
wGxVj1cM8hEf1aYEtgf8oMffQP2IZvRIOjWg+TAJ8JlYtgux++c/6Tma9rtj0Bxee8uewlfCuHeP
Oz43SgfqFMDKslc3RNUexR2ZO99iBVvpmAHEjhNg+xVslZeUf3CPOJnJJjPNCF+ABGr3svmj/3vO
TaU1imOyX/AFaJv735rOJy25PWEoZCALC9T4HGJsT/WExevjTn4D/JjgF9dsCUdMJjXHdAdyozke
8PvN2EjStTS8tCulpEBCimjfomySi333GkScu2Fey52Si2Xw+eSf8OAkBj8z0mJmWx2GQKjpYD+G
HpLYLjZhIY/oa1YBZ898t1X+OpsF1/rt/Sq0sHW/cn0H6cSslJpFoZQAvTcHXmcPYDRLa9P8XZBy
6hD5QQJYFtep2oMz83reUlyqUwoNfkTuSFBCIeGCGHoGPVRae7MEicrOSTJzlVvRLOmjWwNyvczW
BWyQunjC0DW52AyJUB0k/dWAM5DMvl4V0RGUevZVHF5cs9uB8d3fsFBAECFkxuY+PcGhbEaiVtGr
uAZIJtfqwgkGLU8/woi8tH0Bi0xf6SP3CwjBRo03kTSy16VoGZv/EYVEAo6b+36cQhf8W7EdBdmU
i9nYP16zJaEuewOM8bpva9tnNiMnu1fsLQZNA2YtABydMhB30/s5qBJeD2IYDw1OU+LmGqdtNJVT
Xwo8LtGKdccmmRG6ntzXbi492y5EgI6ljFfeHTEKn8qip5cxjidNSYf1fDF3QhWzu769IYIhFR/F
v2Rpck+ScEOkcO6hSWyRcP3906sot/XSygYXsJAzQEkx7l96mG78/u65DKppYeCXwp5ggL45IaQ5
3MUkc2zq/PM0NtHVatw21iWctmlkXDRu6uxh7H7AHNURjK1CohrsrSvxw/uqVG+Ge3tcaafBEERo
oIylnrCBpCSG864p86RaLBgfxBOjr6Kd4RDWpkqPw+ObyZL8EL456zeo5zp598dhLxelO25m5VOD
XHnoRgjA68oWwFOZhmQmBUzDto7AolMixfDC0O5uWhaUTZhEM04a9XxygjcCpdaaWHlpLN1RT0GV
EaLCI0htVzQPqjvwgTc3MKAZb3dDXC9gN95Mw165TZGzCfW1fLaj3r0jnV0nrvxR5iZZKjpYlIj5
26a8K4XIo+WiUcJNxhax9ex2U/Fg7+2ExIPBDjmn7QlQEzWePs7vk9j+kdmC2siZnjTvZZnwdUQX
+yaKrw/Wei8MtR9M1xjaDPNAmT5ymV8YU3K3T0XyYUkH3xYKdbUcTfVGd4VZnCiHjgaq0apDQSq4
/jevQGr22r5OXqV0h/pwvpbDv8wQ3PAIPCxUiQcAfbf2MJXwwtlD40JaKGI5sl0kxJ/ufeSQ4zml
XCqUz88vtgbemXZrwY2Ad94mmdu7Oh7Nih6mX1m6CpyvwoOsXJ6mpsBvZo1U3Bk1fBauMafVmLln
YTC/LOEQq1pKRGO99qiQgZFPc9j/fkkzmfvaxco8F151/HXyM8MI+t9MhHafcG/bLv4zPP0bV8uo
ZVBHrz5qNCVv8YEFKVj5Rj7GDy6AO9UsU6sVvQk6AO9rSldytvRe2quEpJgl5om6A9kQQUjEhb96
SIuMiBfqGtwRULRkNsR3Y6TUEA5IhUePvubKB2NdUdwxuZFgQsB6RYTp0WRTyLNuHv9wUTPh2zH7
9p8XOTp9tHY4d5oRrSE3wHcGphimQzxPyUtl1188HlPAJ1dJjIZmjFats26hX7zl2pmZFc+RqMFk
BCgbra0YrP9kS+RulbVB9rP2Iix/9FftSe1O7F98b1+nRTMZStGpL/k/dRmYqO10PCJ6Fg9O3Mdn
QUjGpHkfTE7U/dd9Gke1yzq/yZSzS7VLNv2EGeJ95HmadegRIvY9RC4LKhkxqOLFcCunXBZTBUGg
O8AvE3tgA3Z1ZwvGv6hmNK54aH5r6yfj/49ppvmqGTboxNPxnqPaiv9Y/i1rzNHIuj5Xjh00nz8M
jCFzbSjwk+ExN5Xpn5XEwOOylZUnbkurGmpCdWo/6NeKxwYX95YqZvsmLONLxFIqnbmh25Vk4zEj
4XW1q6Bf7pdpVbHmkJfJSKaYlhtRF2bkAgkYOQDb3ffjzozUWRNF/ybHLsiu9agAyyf4rNwr8a/s
9/hBOKl6lheM4AF331VuDG8fyRwntaDKEBxrkO7quYAj/AOgwaapMSZGyI9aU4hCKc1SrMOkP1x+
JaQ655dEmdRrAaWgBM2nuzO1rgQOMGIUJkErLB69LCGwxCzdb9xHq5f/IHx2P0w42iQ3RzUpd54c
pMpwxJQMDIIeTVy4y/3X6Wr7sMe+/5L5CFHWejjGngq6NW2mykgpFNQ29G6N9qaawSa6j5JOLOJ0
Rtf1Vrza3sOJ5wJdq+WuzMmO1WPJSn02zUedbPPtY5scVuZxkEy2VKxnwBFThZxcjV2/n2V62GSq
iViLhovHYP8RIUtZpnG1+MbKjIHmSVAjAANCqqxO6p914EWbhLIcz4qaaPSbZDG+jcPbYdjxSbDc
WqtgJ+nY/YZUxzUqQZSC3lg2tMlegm/nnCGRoNQekZ4D3s66oXwpWw84RzoM2ZKhtpEmXWBXLcsF
u3YkBiLXDv0IpZIMyPOD/nP0B4qviPvt+3xn8fzRIajcOQ3gWGex6DcPCiDpLTxXuOu3yXnUUCt7
p3gxlPljdiL0vRJ7Qc8IcG0h1ljUg83GO/phqotMT/0sZCOmSWcNaBh5Awxf4jHNf3HkZNsS/lCW
vrgzN+KvDqvgCivIzRDaC7dBOwLCXSLa27K/LUY+gzEffAEyEelrih1iQJSWHQ81lk2d/X+AxbXK
DXSQZmfK434snhx/zDt+ITfLfz118706C2rgiFjx2b7x4ULGLDB8/pRFwcO4UQRYwGhh2dEwDxkH
EZSNcyg3IYEr2OiKFqEcU11f6X36q40WaGPA+IwZxzLiI9GEngjISkXNNOGUKis295JZAYGAkJHb
AvKDYi1H5wI/lgHnsfNQqoaoHDrhlRcYvDK9J7G0M0p+GtdjjZNTDzRMHVjOStRnVmKGsiO0lFsA
yV8mNbdJmlVUANXm1WAR0XDEacx5EiycFxiK9SwmQbN3NzBkFmF43nuPoSxVahCAAOxvBT49/sSj
hDLqLa5ucouYdAgMjLOrmxuPfMW2HtSciSHKEfFRlDhLGRiUHrBGh2sr2E0av33WrR0q5ULF74CN
TcFEor6uBAwPwPibgSHv9UzdtLIbTkKPzry4S+zu0xO5XMWyBfhsfobDZXLXHRRVNjW3E4wDh77O
KvoqlDVohvWnljNBGyiErWMIOrCnWSQRu/I7KfDwntQMVhK7QWItz1kX92KgLNkgAnF+PK70zIKj
7P5GMkCcd1SgvY5B913MGHOuPK3jJnvV8bZh0qywhSSh4ZLS2rCX3ounco+iVPj6/6F1NDXPr9rF
vq0R/v+EyGw3hlE5I5vjxjp9J5JJF2KeuL/EM2UaCOi1WdibNEP960/SxUqkPAWgFSxSvD+RgMHt
UeYjCybZQoPoS86mEtJhKsbpkHgmfnffQUzIwaS7bB2yE720D6xKKLtnEvruicqsVPRK+JLLL9Q1
S+rKQQJDIcUOfrtMVChKjN/EjWC1JHWhSzSd1mdfl3JK9b3CMvqTRh8E0eLNHGUnJcmy9EVxT4ya
CeUP4e+ePnYqAFn+f/ZFcFE3U9eAEss7VOb3YAWllHWQjxeyBoFojZ8rAgDoXwiizQTiqUYcp6vI
e3gwaEz+NurUMcM1KvJW4ta2sISuWY/kEMijZi5W02QlW1E1bU6SLIt5ZB0vG8axyLCPDpECpAo/
ed8odAn6kCewGeSek/kWd7eUB3cc8jBvcXgYMZyB4kawridxRfWAEkmWUuI/PLcbyVvGc2Q/6qHE
9XpGW+Dzquuzw5NQsIJqaecGZK+zlRWIcCbksDQD7zyZQVgDbdChCYqXRtinebjdBpY5NG4dxUqG
rbRvLW+v16nRgQTNvrHJsogxNzVFUs0IMM7JhZI3G8L/t5svV4u6Zp2lEDtGp2OkniDhzbcTqojD
d0wEKw4gk4h2io+p1HKoQDQMgMbUoquXkmWpcOkQhq0vOwWJgMmoGjhFk5Gtm8rD7wJMKL/u8MqL
KW6BI7N8nbfPLbiZ/oxmc7VAwlF6uA1COn/AsVZ/gNJDxq0EZ2NLhNFJp33zAuDsqzUYYXn7CA9z
e3gaulQLF67Qz3OQ3FxQY5WHArNClGOoLTdvgI7VdJvJ8daLUUpoYVrYvpQoAq7QlMwiXfTn9xd7
UGbnnHAMKI6VXGllPlftl94pSJyT9rsLg3mQrQb9Dl2M4xaUeX0N7U702U9cdoQ6/iwskrXl7g1z
wr2EnIj5owKVe/hukzxfYVcte1oF0CQTGSoa4D/UDTNC5n0kcU56UmFTk6E3PePPl8YwRwTgJcvW
aMJfUJ1eezCPtI9EI1TcbPV/GagUdWVapMmctJFo996d5RwtxKBBiYUdU3Zts0IJ7EpC4zsNx8Ez
MEqM/V45/epIbJ7kkxRdPfz3IZBitaLrwkGJ7rzF78qi0F+oNiimYeuDSDpHrkFy1sCV7Ey3tl8d
X7H+djiQ5ry9P2ysSUztwndukdtABl3mMtOa2XvRleSfR+iEu0c7iUWxPJzh4z3BEQ574TfLLaqH
TiHoaWprKzINEUoB+0pIaqEN/gAWRthxzua91GhmXqMkbbBpLFf478k5+IKKMYy4lO/u0aim78OJ
utRIbqpVz3nAQEbzlfufc3gWTeZuOTvkGcuOL3/QHq38JUBO8Zp0pxUeGD4JXa43kjmDc6lWVj+j
6B+czJSqTEHeA2nyV+ogyCRQoIN23xezCwrxDzMuClJjTSdUpYmr5xcjn5LiB3SqxF7fXqE2gwaV
me/WjnN0Q2pQIjCW07fiIxhomMRNSauEifTJJ3y+RZG69B4wvQ45a2MTVOpuUOpORfYGBMJJ58iZ
1wzJkAvnhj+X2HBXTzJCG6GF38SMnChq1EtS1jEa5aW+jeEn9y1tfKnS7KlFUTUaU1RJ9WW0TX3K
/uE8wZhy98OMZuWuS8ckA5KiyeXeJkNE0SviK35Xuva/De12G8vC+Zql6etT7JRJQ9r6mEj4sv8A
QXp6VGdKSupw9KclAZ4Yb7jvfSeCjycz+oji0taxEGuc84VrvG0AjX/TECCbdMvheCKcBgJDcKjK
WAImShnqeVSoyDWVt7/Frr0DYpzQV+C6qlIO/1WcqkANozNR135EPDIsANkqkBPIxjC7j+ZFh9G5
GdKSNidDJQNxhiOTKumx4vTK2zxr6fzIipe0Nkc81dulWz3VadAfJfEswdqdGGH0Mtj2scudkbnV
0Et8Xbwe6AlAmQaCgbcfD5sVcF2lsf+1dGfntFCBFwFjXztwLb8H4zHxBS6A5YxJOVHXhFKkeFnL
Y95VeaQ5V5k6chlDiyofXnlyrHwu+2nUpbPbEuZopYtwSVYhmPrdTSbsJe7Zq6q0BGmg5ajDy+oX
Opnt1eNkJeTkF16ycrCZVVSPeSMiKWSkHhYHIZtSl00YwsDNBqOFquyasFrn9zCQvhsRHJdjDOPq
Werp0aHUrpSSE+tq/zSdSyRjoyXLMhBTjRCv2HyyxkBdkYAlFCvGReg0okG4TVonmnjSQRsTd3P1
yi75PPaSwPsP8zUmq0mwDu7yXCWcFK4hX0pDuGPRrQRa7WEW104QecJTYl9kNeqiL3C6RDxd240v
zOrpvfwI+MdZy5+Mw+RpALPi20VCTyHIplOXxaxoU+w60niXkifnwzORGwVA09+Z0uuyNimd1fc/
qus6xPVAvHPD6MI5MhSz1GFGMTpaqLIgkg1fQEvvS3ZMqnXeEWvFCZWWnAWlyzejBK20mP8iCAeX
6qYagArglj5zGo0xZnWj/tCTMKQfcmJeRaGHxPvg5MQmFrWZeabltNTHtm1GRBn+cpJTvybs3ya9
sZAbMm24AbguufzCr7su/HnUkZ1FYkFE6VRD/Yu9FT9YF3PkfxW8xEZf8SWq7GhLHCRlyAV+5xEs
4z2DiaJMp/CjfJU7ngdH5jZxY2KZCzbSb1vUoJniZd8/cunHOg8ILZ5I2jb2o9QgMH8IhSxtGZKL
PDOqTJfo7Uzu/jIAig+BQdZrZBeH/Tev9RWsgFRs6PHRr+7/T1cH8oniKxUrc/t6w36jHKzyXM48
bHwaQ+QqhN+/YrX1+f29ZW+jIbvBUHtU/rDKqFaA79HfhyqcLqctxk4gIHzsj4rhmhD9R8Rp0Ozg
im9tOcGC6TBnTILufKG/mRIvQbkML57bN283c1GxwQShR8GP0KsvGZVii35bIpybDZS5uh5BZ6iw
P8CWCM74h/ibdUMOuvFLS4yz7YEAktVxCkqYwNJDHMVNXahh9JbkrT5yVbtA5LX9xcvvTcAjqpXL
fWnUMmiHU1HmHboNncp0mHwTtYM890PKyTdzmKFvfDFbTrMYIT0oXQVWRN7/n2Y8NAZzsyVeI3zy
lB92pvs5+XUVJt1quI2O4l1+iN3pIyAccXF9Z+9jzQMDWvjHbGNZmbrOxcqH6a8lZZ/awxNU38rD
ZIm+fYy+1og07zfTPiTODS8uG/+imdColtaEsAvuKJp/I9lyQ1d0k1SDk5+RnA6ea5iLdCmZzy/r
KOdoDr5Mxj7br2SyCrwX6NoZTLuRcp6yLkWubqXC2VmknGGrhX6j4mm2k/KbhAXgQUmIbQSsD5Gi
+/6TA7JpQnlOuuGzIj7cCG6Kc4rQ6XloUmVJ2yseSYDufY7618srngcb5Vtszw6QTNBgtLHqMaaK
0cPnKSzNzTOiLch3KqSjhSAnvuGWdU/zkVhChSlKaXR3cMIsjWEUyEjws/JWdqObEaDqE8boWzND
S5i8j9cxLdLqyxHHDW02abizSiaGAwJM59ONglrxGJT73qdCEBJ+sCsIs7jIjvgb0tmUf5R4mOFf
/Ne0MiCNKEAId4H5KK4DoVqi3yNu8Zff9YJeq8qzBIdgUhW05hGD9ZbAPzfITiVo1uc45BU9vk/w
hL/cmIrqqrk64oe8eGO+MUQ0ozU0Nrc2ul75at2JGlrGB60AY+Z4DID46cZI4fxBOAlyqatw+4jq
uCIilu71a6pYcXEKqmZ2ShEJ3koOLz8vp2vECfhLuhJz+M4aQDX22tPKMSLHk0s0wjN21hJvX+gf
NnHFgMfE2Zbql8XvVABd1rISuoLLwGG3BCMW0VEboVISyHtqET7mYLMuadqr+TpNfF4uSP8LvZH6
f0BgojRLP+gdcWX0WO9zUxDRKIY62l5vwyOPv4DBOklvlih3FhPydRdLbgip61qy5Jjh6L2gaeDv
V/hDmpEkev0LgZ8pHtxXM8A0TsFgRi8V1SLeu6FN5pz69L1ZrVE5EjtzkIlo4xmwvEl6M+1XvtkX
ZaQ6SyrYS8EnZVtMYuoQ9A9UMqG348kgBKQrgOYLii/8WxqbYvz6YboRGi5qxiSUtNkguPiGe3gi
qe3bs104F5KrvedQcxL7toJZlw6V6SPS4fwyLhiUkjeov3eT01fFJbW93HMov8rZuS0bin0OU8th
UUIS+vOAcxDoxEoSzzB4nIQBoGWTyuRc20tE1ZixsIitJ/osVYPD0X8lmn/XimzipNxdw7snubka
WhMnbRSPoRqurohbo0w5K/igWSZkUMpoioHmohnESKzFy29n0ybRKJyiBdpmAMoL7Eq2ss8Go2Bi
PBVIgZA82DIhThoG+jbYKj8hSJcj+I37vL06gL26KANaGbEIRdiCiNuN85/an1Yh/JB/R5drJDv8
k8tjfK4slA+/JhsjG83Q7zfwWOcbIBo/QZ780FTkYZNDPFsLZiSDlY1m8e1F7K8reAb97+kJuwAD
GPlRmXbgVBsIV1E/QTeGVrcxN+8lF5fFE8jWRXMsiUMzZza34a7Z8ZsMwmI6ye7Tdfih7o4CHfxG
2xso1hwqPqb4DwwZlo8KCRrpqr7rhOzkkzZNfpIcKgANc2RgsLfHPqe5IAphOPBDJKMIJJ5iT3VX
0B4nGCJD5CKejWhNsacHrVu6biMIFobHX3Wd2oiFlOdl1ZJ6vL42uJcLkcF0ozGHFycrmwsz6No7
a6I2rUADv6VxiAyKLAYquGnISD/pHVP8sS1X6X5I7pcRLL5eUhIXzNXnHWKpra+FRpPFRdqkdO4B
oeAAN1313r/d8Ob5/q2vekXgaRI/WB5JthJi1IkATcFtB/C/PY73i8bDegrPtF7TyxLnX/Sh7/wi
YuqJDJFaeopfCh3wWiUb9vr/AtYgWdlWZy05R6C3pxS0UOYeHmS2+3GnSEz0/alLFUtElHXF1OXH
IGn9rR2OH/hPZyWAHnqW+8qe2tieVxF+fLtuFibHPpAfW6GT4xmfRZxMhDecH8vUgUcO9g55cYDw
XfiI7WJLNcSML9L3TMGyKFiBOXpWSWEqiMU+ANIdL7m9SFHbrXkTCpfmOPksLS08hIB+F2TYBy0H
E+jbHEmFki3ndqxDPSVa7RRR1azEFE6kvs7QVO8zGgx79lJXSnwqe9wPMLMgJNPPQunH4rl+lMEu
+FXQ3HaaEfzbfHOic2ZK8KMFEm1YdR/R6PRUO+3W8uCH666SdupUMyUPMzp+TSR7pHY6mzXJBQWM
8zHMlMwWOgL8526xL0bUoNNtN/3sUnT8J7aSNSIgm99yfv3IHn+esGXEEABjPewE0cYxTsIZ2dTO
Kj2NGRMHOoBpR2JMPUZxHXCkH+c9Y/N0c0sWJAiAcnTxVqWeYtu9jv7qFZ2luiYI3bT1lGEANkHu
GoDV4on7JHQf6YKyE7PdwOPFX/4o9kzCcEZ/o4PQoGfbKdZc65bxPkKvGu0VI18aLx5jppEzno3r
9R9pKnXjJ4786hmcvm4qwfBDbbjX3g8oNgve7gycTSN+haD+shj7OEaxIIXZViYk+ce5QZPnnkJZ
3uhzCDqcLtV/5DYUJhQcvzrPWc0UATlfP1ZP+HItYvhJ//FRYO36MB6A992KXNR0cL1zmETzpmqj
2ODXtuMpZbj8dEFynTFM9MwmSiakmcaBi6S0w5pVcAoNwQ/ENXdkOz3s19Pd79KW2cXvjlkuIQxj
DyYkgoILBt2TUFjLgsO0Dqgyo551M953FkdR4/bkCGnRANfelW72rCLsSlxGinj+t49DpP5XNGsV
l1yjMd2afnk4Gdo2FHnAJYWcrc1Q2KCHYK7RfX9Y90VvgijcOsq9TC7MQivJO6yFM+9zMlWVOJIc
YGoiYz2L0s5pJDRFkCSoHt0GuWA/vHZL65f7sqxAcR4yp05PgdD1Nm7g6+Jylp/7f0xoKMtVXYbL
8U+hVBSsYtljXRmZKeRRSrWVzLoEoQmeq7G3Y+prtn8yLdrwZL8A02PVg6G5E8IhLYOL2VGnwE0M
oehF394Gkl0zIc24G9HqJHGMCLJc4CQ9DcUx1gP+T9D4oih8hxY4F22fyw6J5gXomG1HcRIkJrVE
tbnsys2u7+XlrAxY1LBCW2W8gL2GEFAzjr/7pwjsqO9uUNx7LtPA/2hZRvWFRKXYtHeBv/BWrssp
EwtCbg40msKNCga1KAwkFHXuW6s+RH3PzHXA+vNeFi+lj96DmgtsNUWbikeBij4pQyEGSWUelXpu
WCwu5nyJtxJ81xoNW8v1t9YuA5jGRkeA7NN8FQjdw1lHOmXwr572ZGwcw8i52xEHwnCQxm94aLbc
VPf3q8hYS82NMGMFRoP6xmf51eZufYYAGg6sJuG3QjNSJdnbVpfL1TReqLLPIjRBp/PkBbMpjD0o
yjLwG8K9vmlpsZghYZHBigP/JuowQwiTiIBElu6rZ4ASyhDJC+zOJ9GxgfFoKyMXC6lpBjTCZkPc
f0jKTX8zm9k+xOoZis4t0c3LtBJEUwj4nuFZaNYZHEfOrmphdZNICdFPp1IAwHeWFmZJY3qoo3Fa
Ihkr4u+kusMYpGz6f/bPcx2tIeAyQRiJt6K4WuSITIc44cry1s9xgz8P72cysdIZiY62L9r6ei88
WXfM9OaKR1BdAzk0SHI1iNpCbcQEy/38a8K0oTkcfNfx50/kupWFoKNTVzkJ4mXTyPKL0yAi9Z0s
s95clfHYaJyiIAXIfvCP5Nmk/GS1TzYjThIM/hUbYQwW0Oqm2tko+7eyx+rGtEMY1UFyHLrA1QDc
0Ed4wWfzt+hjC/TD9Z0izr1eLVD8MEFod33qgpXXYKNSJHJqWvggHqhKyLDDkZmYTk4CD3pewctR
1uDKRCI5UHDJ4ul8vxZOYa6yP5cFBLMzBNfQavoc+4GV8UNs98QULpVXOYR4d+La9k3A2SOr98i9
KZUEOK1+XT6WN1MurGoDDCNcCRYvfCdrHwcMS11nsiRPe99sf4hQ6bBxNLbdrLaWs0mDqoHYpdkB
CfP2C5bDuE426jXVo6iV7l8pipTzHl8jDCQe1H0M+WOo0aB8ceWG4+BJWu7uVDg5VIyMmK8edpXg
2OJfU4I7C1iEsRebKayw+XS0MqufjfjVdk5Z6i+gBzorm0HW2bDOpSHUImTSfqxbybRDbxTfO37R
WrrAqhEy/U3gcUP54x8rECo6BAAlMdRNRh6gIcyaVtYtRaW3XDEpdzUqrrgUUylzOWmvqODM4usy
QA2SFGcgnXRxl56Xsl64MczYvzrKeTNmX6fcqRYRRnW1aF8USYNlPpCGbPgZSF1ReWtO9xWJH7i4
rCGy7dfXiS0mTMB4O2znK0iJy3bNClAL31UqfT60WEpBiUUfCPtEWEnJnjuX5edRFs1ihALJmEGi
YVw3ZS1arUvkcc0BzXnrZPG6SA9wY8cbRnFvB8pesYhMWbUJ5wLfrI4VJvyCJfexCcO237N1MY6s
CBMCRgf6qjAuv0CfA4BW8pVTBWVwo8aycvf15URF3zMKZBKNFgIr76+z+nHwvIU+k6UCniaCf1sb
9Q9zDWukw2ZoCiDcH366LIQ64hWB4aV44XQ+/ZtdBrfvVlRY+Ytbw+L3JEPYlmc87LvMEuSh6a1+
aIpTCwbHRhBNMdlaCDQHe3uA2mRfDPehJektY+mffks6D6nQMxdNzfZPuj9wcCPnkWmr9keU5eoR
TOuchtk1EBS4EdWKcM373WiXgxqZkLcmf1QZnpLwQdiJ3qldZfzxOMVIv1UezhOpUG7WE0I/CmAJ
fa+JddbmnMTCZ+78qPxzgBV8FLrE/ifSxpLZJ1nD6N226AtghDN9kCOoUfu2wszNYMak31NVNFrH
16aSClUVYkc/bsDA5zv6X9YPwtntq4s3a9TFfNkZcc85VTgyG/eihFLYe0q9F5Inv4JPSbWWZHwg
2PxibMgcuAY1D1UUwyJ3T6GrejNmZkzOWtDHr1Bj2G7eB4goEhD0mxH2LpaU57XmVwErd8q9RGm6
YNBDw8chBI+07AVRBn6Z8OjXjOCh3v7Xxbv7NaiR3t9Yp27RXb63eRj+Ie85WQPprOEjtzH+tTcF
UYqPQZy+SOkw9b1XL6eMTyYT0zMEL6Wc7CFV+w4TdKqLPgitGB/PWXf7OloywlQFS9EBr2mwjWAm
DX9SigQnRnGt+XdHNe2NyCh1ln3pM94NBWGu3S8ycjPowSgG4asM62qVPxN9/hJZk6tNaEV8ueS+
H0ey1TuThkVMMK/Ip9niVlRke2v7mghYzU99urhC4Hf9Si9NyOuFlDLSCpSJ0jTTzHYnVKAaMUUx
5K6fXMHqv2XN6gLMnaPMabwKzoJjD+FKxMuNwk2/180lNCWclMk2x2mBK6oKOp9eP9CoG6JaUzeY
wgZIMWmMTNd8IMRybsbYU+Rw7xMbDlIuITxDY5/VBkVYHM44hQdpLJ/vx03zj7mmS1pid6YfX40o
QADbCxuLtIUGmUVTSeqF15KMPdHBZmGt18C1sL48Q66gjpY30Od4QleulwOQ3WA8eVZjLG/+pNMg
3jgLehY3tbGgvnBuQXQ9Xf8qhkWb/MS1TTe059ru48o+GGlvqTItG55sUxJ3tkxzBjzg4zBgbUUP
Xr1A8/JyoaqIPhokn90iqPfU56BP0Z7SdbdOT+Lp8H7d2iNPtimqRCdW1quJ5Z3EGKB8Lus+n4dS
ELUOEU3gF3E+XtghzFvFoFfTRv/EqT1D15YCoUJ/xKhtSTADeEYSokO1XflNNCw2ENRLWEWa5Utj
UMj+JKlKVMhSsY2Sm3p5jbmlaGgLomA38WRI6wDtu6R97Cv5dkibHSpNaP1iq2yvrtpwdpRAG+m1
Z3btok4NQYLCNqRqEfLj8w9xjMHWRlMvsAVoCu6IfJwmRMB7+ZEQff/2tysnSq6FS+7YZQ77yQyY
4tvFPrBW+nQAhLAJlwfn1sDZ+fc3gluh8WJ+aY+FSmyVmEJN8O/gwg3IJ5YEm4HFOeoDB+X56c0s
VSjuk+vLmShB23ot6EhUglylXJXHy3vjVTwym+qZ6vm6Jl5SRkVsq6TXDbtTYfqNmpczFjz7c9Cf
xbcKMCXnXZ0qq+2ueaHPF7ZsiNu8RdL6w1iZ1igdUUMkM6Tia+lSpQQflDrGyjsbV52OmIkCjYUS
+PheDsTuNKCCQ4ufN65XKCjBcH3JPol0GZHfofkVU2VyKha65vmPGoecxJzDjGDKMxjVD3NtPjyz
stOWdGnSmx02teMivFlG6kJKxaU3VbRg0bqYVm8TSOefBlTDWLWPV0fBv5vqryV6lEDIAB2DZwxX
WZ/38vnt65Uevn5y42f4YkUPl5UeQ1HqiMDsyQN9w/ifFtNzzzlnR/3+9odH1fqEsJ8C5yWz/REd
f/AmO+PL21zUwjZMuEmJtwpH21EFIcinQXhZZudwPhE3gH3LU8B4oKZBWBYhDV9Tv0tBoPMsy9/A
bXgY53W3IEsfTKu95L697nCKwklYwdvpqyjOxh1K5s2PEaAGhZGbJIDgdyc60+JOqOjBj2QScj9s
swc+Ov+HRFu7rgyHA0di/zVtD60HdWyZ7yeQMYdo9Y6pzImYO6xLdWnD1cVpZBvE0HvYsjMIx0iy
NTmTReR1WK3QbmW9cdWTw5HQA/jlq55VKAx3NUyrZn3p2v7C/h2uYWOmfPOb/QLnT+OusL/NjNuZ
Pug/ZZKUmYOeAxmvCMxvCEaANf8GMBFaRNkwrLQQE7Yon00jYYtyTZ9e7k4hEp5wluOqT4iS/SJE
rV1cwxj9WSQWCNpRrNF+eaBMQbYM46EkvsUpGS4AjQ6n6g24d6wabGMgahzmdXHNbUVvZCtFfgOq
A4sCfPGVoOYnsoOnauK0sGKAdFjM6MOnKGSICXT77qz7K6TtnCZlo8SPKaj2RL3EsvAkMYeRNa4M
zy/2gPl6yPEXq6E69Sla1mZTU4pWQO5B+x7hujs8LZIxnXtHmYl30bNJ8OuOJocv6uJo6xFGTdQ8
wIJhh5LbADuV/oM9I5o30ubwSZllTtVJMZ1uqriM7tdKzroYBLJtPgNcfBSuUDJwJRbStzPxa5l5
1jMPoSktL/2bXtK7N67wXLjwjcCeBA6Aczb+YnsmIEV7/rvvpuRhWl/7V4le/H1XEuRB35QpeJlE
edpx7E96rHAsHaM/od8BftEWxCAezShliCE+tM8Dcmfs7sLgV5FJsFtgVpAo9WAkiQK14PpZDM+T
virUJ0NoOWAOOg73KpTpepBIUhqYrcZdNFC+HaooKmTJ0LmwvDTRoOXHIJF5B5g0Duds0YtcFGZA
LuYhEB7Xpi+4dpFbZKgMzMxSuzt5a1JDjU4NV7x7T5G2gIi1VjiejNG/YShlongDUhx1/SkkN0IJ
HO/GnS8Za/kxH8VuLveZp3EjCeaBpUhB1AZb3CIoZZ/mgUKIV2Bt+gvSrCZb1u+th9pJmyAFh+13
cGZ1bW8DIGou+aWfzvRSdad65+aPLXZP5WA6cOcIVX+s8DIU4Fp6f/c6wfikKM8M3a57bnwMBgNg
9WeZEbWyX8TTernRO6q+AxuruizBE5qCzHOrNB8nz6Hz6KfIjyj7qIQo2nrEbJ+2xL5wN5FuL7Y1
PXIkB9QT6xSOn6A/7hYih7v5QH+v9iWSjBuTO1Wg3BpyZYF5YTUqhRUE9JJr2fhWmK/bBX0DVT5c
rj61ReuQu8SFDhbZBvzVLpR9/qjBqWPBTGuTJ0pwW5biisU52L/cDtX5dJLnrTnxj8pihr2swzaW
pQCALqOju7IrjKm3oIyPhKu0hv6qrY2aLpiOKnF5peXTj/7I9CVF3tlrz1PPGgCo6/aXW18MGKOR
ciiatf5N1uSS/yF+B91AXovP50jmqvNV3cPEuP2tT/d/uTuLcPIXHP2FlJ2LPgDioY2JGIBN5iUJ
m9LZg9LqaxgdMmv+orQrWOO5zQGK0rMeNsFGz9rKFuEKTYdOSHmXVOPgk1Jfmz6XzWk8xcylDObJ
+Ca5kaJa+GA3OAAdPY4lDK3Ejtwcj4C94o2KeilnNX1U23TLwHM8SeqaK0voN09R21FHjGdLe3rD
9gKWOtY9d45Q8cbnPybAiyf8h2cvVPmnr/26QB0CF4hBqD48H7WDRRyT5VcsfRYss7dOMJPQDYeP
aohnSu8UtvbdPEda6/Sjc3EkdDFNMZuSOjvDtdtraqMSWHQp55qdup2VtKxzT4wyZIKjaMvSZ2SM
03HbNhUGJoVOObsyA0Y/qoruxErJHqSR681U38Mq0o0kW/F4ieW6YKLD+wGHPSR84TZSok3uRV1p
XRdMCJYrw8pWmqv5Jw1Kxim8p2SCEkUE0sMHMsEVPORnvfBG0zec4o+3veDkDisvVom6Op+3tLP8
UVaqXGKCoqL3uY/d7DYQ8iz7QUTWZECvxDHdau+MHqNxupc4L0VcHc7cM5EVWF3xulnTq3tbbG51
Z9F09B59p98/JLIlDvWV9W4SNuRbDnonSkfVmkEGaneEJY5Sm/6ErxGZwTvMBKNDkZf8t8chzbkn
4xhUheKD9xm6h4Gv21Dzxlr95YxAYcEWa9a/BDhIk4+k2CRomv7ohgVQM34ozto6u5ft2NymVyoT
jbuYN34A8nUt+QxTTM+PPVRJA/3CRZUdR99/R4HECsFQhvZmZX0OBYSo6tbAwvTGvZufCJU69eNt
3Hf/SjPaO8DTPlGqxLqZr062xby/lIH1yLV9/ISaJqLDyYGXl2q0k4/lUmZYUeAybIyrO2P/ue83
lA3TeuIoVqwY71je9+DQMF0OIbzpm6hR49cmtQz6tx6wx7dkbAszp3lyTdwy0DuU/CvqitH5GH7k
IwMe316f8VhdG26N6BrUlZTSlB+XlWjekN+5DwyQX8fZvYhhs06HZnCjZfygTWdn4mH1kARsvqS4
ToAlv+tpmY/wWymp78om+RmNqoH9hXdnUhkN0OtLLBAKXE8Q3vv6i3icocfolwhGvUXKKcsTk06O
hYNVS8j0fy0epAOJD76L5F+odITyWH1hSc7IRg/vfE08wqNbzzbnht/mrti+JWRvD8QK6kalepg1
L+Qc81SjFCwY0JUApoykvJCYi3S9HsqQ1Q2egZlUHYhkYFOfjVb1Zcji4XoWaUhpxGkew/rcABF0
LIoFN3qZg/VAJ+piFmbh1w0PComnAf8dKJvANLWM5HIbyF7Zf3xrkzYX4UcGsUM4kzUpPg6zr9HM
XEtk1VfgiUDP8A+iPraiSq/u20yBa67n5cRMnYDtnbggGQBOz9Rll2GkO1IrxcpWWPToWa3euLhj
kJAhkniOWSaMhKtBhubnUITZ8Wzf/ByzaG1utn8TNC8ukY852YkC+MWwlZYuQUyprZ1XBw+5jsse
+x/9zaeHbkUY528Vp5BLpKKBylHxy6evvlNyqly9NyUwy5DesHEXyfkBTZgZaqQV/6ojahkWOPE4
hj8z4f56xzp3uPAOnObFrxOhhodcftrFAqBDXXmX1UpBgbr5SNXE/FizKnJ933HoaxCnjlmGXZJG
tZ8rjVWg2DSpoXW9wgaE0J2UX8tehmqGA65uRKTgM/HJwfVKZLGk1HlzXC6AuixLJgXkA0DIhoA+
z6OUrslvDaxDqNIzABd4b0EniSV9TKmpIRyLYnzN3R5+VwEeUabnooCE5W1tzM9tbK73/X3am02H
NTpBQk9axZwyv+oxZQjKg89R3TVmsnhHpaiG+edIhVbrCgljnOnrBMEldR5UmPnjmjPtLJHS2Qb8
7538W6gkHOSZaC2WbjyT6Np0vi9SkzKEmV8j1PMb0e+zPjJ3MW91Q1KcLGiYBbO94S29A9OjPgfm
RQvvs7Lzo4nA5BjL62aiSN0Kw9Q1SZDwRf547hr0Q7OMMcQEEbqh6ExTnqru8CRhEAwiX6MRzJCw
7gSmfOp1s9XPP//BbJGHsAHj6NvCuDh45UUpshFkLd3SrESh6loi98jsC4VCg8IAWdvGxxZRNBAQ
2AEMT80quRL0X9+Z+6pgEf3O68F7iM+elHvv1RayNIMTbV7HUfEzyaNyoGpqw4CQMhgCeX0vmszZ
92qAfN9c0TW+atwZVNiDLPhbHlJV6JusOQtZ+msQMOjutj8JczoGLiHie1bnYLljdS38syw7nazj
vCt9NOFg+vP3FTJXlEcpzbH0a5Tf+YQdZzBHREpjeeLdaB5BUutNnFoOa/FpD2wQDEIa3ePFau0/
khOFGmmQlV7m1TfZ0pccsoxu6yHDcymNxbC8ftSCG8T5moUYXOS6+Ws4VhWriAdzsvILe6fzc/oh
p8nMreT3DK+ihk0aiREdbmm12XVtkq4jeK5Ith45iV+bpGQeQLyhLgKo/+CGHOuUPJHuHdab868G
ysgaSa1bgdsQHPOU0jKuvspz4YF4B3PXszqNB3PGuDOWEbKALFdDko5fzLNqPCzkFv/hkVh2OtSE
iFZG7/O9XF63/1GygXW3V27YPIr79enYkKiEQcjGgfJikCascF+CFpIv5xiJiWp0zL2f8ImZQ3vO
6uhGRLr3XwwiA4XJwmwMx3ZeUetO7qhK8dXWzuiEs9eBu/xCvPjPI/3JYjaK/3+toJsMdOF4eH1u
IxAmon98U9z8+UZUmagWmK5UDL+a5oBbmnLSZ+GXl+0dHPrJMq31+EvY892KSmCut8k9m2xQnmCm
co5qEJjea6z1zlWHOUDUqo+H296u/ThbSqYJg2vfFr9s6j7iP/7fMi8RtbvRg8tiqWdIX9R4KLLj
NpSL/Dtn2zhXC1A/YtXf4moc4zLimFpyYtVeMphKi7z1iLlx2deDm+tx8JLmIDoW074Lf79qMHFr
692RDv2WUvTNjJftO7+GYrjFXoKI2Fj+yq226DriYDngUxEt/YznrHrix0ZMO7BOqJ47z0m7MdVa
rVx9LW1ogsd+iMD2TxkEGpKaPw8RJhQJ9JYUJmv359BE9QHFfasRVC/MpLAOtL+4gJE1Pyh93GBL
AzbNBAuvGqn7wAU7WYzaRcPRXx6ESzz2KTgPSLxEKpdFxe6m+vHErwK3KFJ1E7mPB6GuPvwuBYNr
NxOXYiAChwPm2eqGtxEHgI6rQR73RLPHvzlYLaRLocKn+ikzxh4b8FAUDK7G6bTVk0/27aLPVGhq
Gjy5U0PQlC5NlhgcWk6j7e1X3fRi0RNvUFKbTu3RlbfwDCE+WdgioNT8sayyhkS+4PmnQMIUHlsa
uERT2az00NtO1pUXcdVn9LvDRY66hd2yeQBLWtZDGgJwSjkVGPY0EV63kkXUVDp6yMdYQNqaYFXC
2wCnQI/tiJmr0cQW6L74J4TRLDT2Gkvy4GpFGpGw+cKI9VY5+nj39ttkwb9Gqy8rZvjVnA218FD7
ESxtdk2KqIAJ3uPBfPCopg8mgd2fCXrzcoryKj/5OTS+gHTpBKBsuSb+S+L8GJ2lMlRBsLx7YDAZ
Kqkey39LTbrUWouLcfPXiHui5I/LL4pu648hRAA6gteqsK+UXVtA9zwu8tZQMHWNDIWIIbN2m3GY
tPm8/TqkfWBVeQfyGjDUKBpzHZm+SzFMOWLleFnc9/UDhnb+8e/e37bFVZclqTQiz7pttsAVaMis
OO6edqeWCc6HOTBJxwzgsTtLds6ybVxn6+wUsadTenVOiham5kLpz4IeoRwIWV2GboL43FSAt6k8
lHJPXn98VhPea54Injhtk/QthEbJOQB+VfVq+I3QyQe/foFdINjnjO2dj5att6JwHWZ0CQ6neD01
R63EI0N9WiANHFDlV4ysZ1KK84h37rKniniLW8OPfA+pIvgkHQlOsu5tkfHruq5byTri/W9zQhEB
I/cdCsDphliSPgMszkXOkJFLPysX3unjZuEA6qWUUix3MeBzI1JJWhmjHfKIuRVQ42FDgvWv+/uU
YObtfYq0ry65pv5/9Fbhhv7vOlDknyymswFSxUA6zixigy3kLHXRhNvbSTsSkGJa6p9i8yqjL2bI
y04zbU7RyNgfHMw4blMth+yLljsvH9caYKQH73xiAe0GZWwPKK+KcTe6Ol8eGn7d6OUxfyZxOcM1
beKzbHlZwWXukW3Eof4uk2Bibqs3Z3/vELbmcf5jO6jJtj587XSV2FgFquGOKc+Pk4UtJ+jBmdfY
zJmA7PIn/B29UP6wJJRe8Qenm3yTI7KErM+/2pbM6PSn+s5jRxh4bR4LmrqptVHKRkKT6Sfa9vWr
p97bBscOaR4JS5tcxWwaVxU22WeocNmBkBlyurUbkeqMZooc3RYWVyvOWxTjxGncUw2KpbbNIAFN
kg/tdZ1CidH8H36Ey92F+cHpjen7s5wfSa/0Hhn1JXP+x2yH6Q3A/2aBtyJqy9BXk70z6aIQmQew
9LdP9JL5P0aWROwY7/CmFrO50N97VrEpCHBCojdtaKZ5iLue8wP9jHKYwc7zYbIdRfQDy9RTy0jS
jvbTLhCCrUmDoBNNrH4BDG3DpUmDaUtz1FtrdJ+mFANtXl9zNRCW0NdCaAJFFK86y2U4zyFwOVBL
PqvjPUF/XTQqvGWYysHDoDF1oMOMxjECbHl6+V2MqmQ55PWmbX+9+MrTBoaC8Pc00Zop0maR+p53
8zMNv3gBEuaSOX2mGFDovNrULjWXdjdd9R8703PKoGfWXUnUkexGRThu7f9UAQ/qegVDON76sc5O
foQBJmuBYsmUqtV+e3ws2+nZF1HasWxpQsCi8QYoRUZJ2XbDPWOTiW4jsmoZo394NCzDKYRUs7hn
7JfaCwVhnetny/+AgJG5I0ZOYC6O6pJpCKL29L51inz6Y607ydDbOjMfZ9NPh/aPqzCiBZvTOpNu
NEawM8ji/RWO4S/dtosZv4AqnJJnzbE1TtsMjH/ZLEbL/eY6yrdzBaD852z+rYpvqzzcxNCeZYHD
usdhaEr0ZHVVJe9cqVEcA96eAgR1cZXfGs34Hxkb7I5dAYzsSo2orFDBegvWhiiwYZfFiDL6X0tD
9aYRIvw83vsonpsQha1NJaDC+Gz6IHnKNqSygp+Ayc1RtEKtOzYMQrKZ38ieogVlRm/DdtmWx9JA
qWsclWcHli6prbBSME2thzw8FO2R+HygSJ+SpgtDNOgNxdrDixbYxmrO/TPQ91vRymETqZ3g9ySn
Q+ycSRKuIenEWE+gPhEZlSRoOYL4pbe1iSE4v2jE7tuxcNxTSAan2tUxbtFo3rB37/ckpXluUlN0
Hef8ipDdxBYHFFgSnxyqySgL67zAdl3LoiODBQx+Iq3S0NszgsGFqeGtcamLvxUAex/WejwuB7ua
rlwsSFcQlkppL1bKw7RongxpnNPoTv3OcnmUW2zHv9/taThZ3US4dweu9wa2eggeVv9LPDF9ZkrD
BWboymhqd9nUlkGO8hZeEOFsxiMIJtnvkucdqHDCtCtEdVz6xnZhu8mrRspGRhC3McGWkTGy+LkT
yUgnYZmst69GSoYpP7Tv3/SNQaNvYuvXQJ+sYC7xubg9pumB02TRr4w7O8bswIswKghhhiEn4TA2
HFl+L8JHnP7GLcUDGzqlZGAWQlKHVG18lc3GwLiLQ3qD0dmB9dpMUw/tqrAOMG9nofPJ89/dL3Z2
rfmpFnHxH1uuwygcKvL14W0/wZDBICqw4eTC3P53PX2ssm90ysm+5IUuZnzIEReBVXrhIOhEV/SS
IsE1INTsPeMkt8aLVz/7Lbi8vY0r2OLedT99v6RIK2kQ48srbjwTelElICqwsFs8fsMEw3plez2C
bKjNUbWh1k6ZavnYlS82xAZrSCy6ewSC8fN7x+/s9ZGe9WY/ba646miKYGVn+Yxk2eTopB2LlrJy
GiBFrMpsXUSm5dYej02RGcjNuJnU3W2/VxSevMw9V1bu1kXSErs+htjghlxSmb46PvwHVhIAb6M8
PEcl6KG7L2jldm4YaLZErCfuw4U1COar9Z1qk37OuNYLHMnBknKD3L8SvkBVILaCj1i4REMJMS0k
MExyCaCDHPWHoxDsCfswuUKYw0elL1gY4wuGp+H8BxRUxVCepqMCjRY4TuDmFVc4beToWzWeA2Qm
/5xFV1NwLA4Zkq3UeYHNDpGog2GfRz2qM2eHHMLenO42yYjdQBNs7+wVzWSomS2+0ZpGL9wMGgn5
fmcJnqBU1FOOdoANgRnZ0TVktTWSzbFB8ah7+jHKtb3W2C2sB6S8ikK0CMRp6nsNPd2FnfWbPy4v
1xuTKymZAm6zrl/R4kgy/CzvkATgIavDXixTMhbX0Ty1cwELiSkYgk7PmSa+C1acXETUfjHofCW2
P7Qt2dVbfvtYlLZBsIvnyiBCvSmVfBp4LzfBC4/rR5M9+nz8oPGhrIQb7BnTjYxTlx/ORozEixyc
rUzUTQupv2rXWLmpAkhxpnVeDXdWpBv1TZOvQ6LVl4g16bZqXO+faBCaCdlyMbcEIYwP2grlsptx
PeC7CiYLF09OREsS0qtxBMwbDlD/zpzfVE/M3SuUgyrpCTueaLUkKr4A4gMesrodirE1JxjelHaY
cr8+UPDcGhFWtg1qBctOLsugP3PPhxLFQJoVLzqjRBscJ6GtzFEhgqwTK5IskzQyPonylMNgz/f/
Rkbe7FCkNYGPJFbV6CcHr5l+cQRz5Begf3P7K2riUw/3NW4ZwzLfulApD2/rHiB/g2/mU/nmEHUy
fvrc7ZnhgrtSw7i/n1tJ68ycpakEPHIOzlQ4+4AST5LUT/y8/0X5sSLg35buAyQ2NiazsAPANHsB
/GrdL+s7Hkt1/excDBD45XE1v9w7+4lOusJCiP5sGmnpnbAgRbMp/Uc8YqijSvsKbwHmlS9i4qNk
o+Z6YhlPxxZz7OTsgRGPSYZH0KnlCFTyRl/MzCg03PT7DR8g4TKSn5bht1bh5Gi4b/6XBrNu23A1
8/+FwXhtSMdhAqrPCoTGfO6oG3/HzzbiuVCG0/KT6pVvUGU3WsSPu5FTUxq2144atxVpz8j6koLm
qlAaDl2zGzokhbwrt+qoorOc1qq4BDYELC2WS5iViRGAnxMkUffV1SRo8/YuQ3eGV3AO+s5Uh2+1
tBd+vWnCY4mHxbVSrJy5Gotxbs8lV8rv5eySnCd4h4nS/S/kxkWVZr+GUniXZiwo/5DNOuls2jZM
5OEHH08UF/kp/AU7SFT/GGlLvabYvErbTNFw0d35w5OrdSEFctWaNjcZGF+SYRIEAGNPAS3FJYMR
HfOLRvp5wNlod+nvETWDkfIjSlV7Po50oF5ArUWtFgFEc93AG6pTLfmrLo04BfvFXl5t1+gANHmk
iXW67e9PEmrVjfKqShxYDfgLQ4ZYc7VyfUt6KZKSZTyoUlHJT/5RRqiD9yUQSpuOAQs3bOFJtvpn
Q6iuzDT1RKyfW9ZQsBWlL/bTtgduPE4JoYRmHVBWZtiRVvN/J39zog/0JgMSH5lmEwqOnXCa0nNv
w02Df98ijEiUKqBQU+grdlAYP584qNgBHqvE6R3r4MEQnWWa/N1kf0zfFh4yp3Iqulwkxj6HOkG3
2i6OHIzohRciEZ/UAWDBuaz++vXIxWitPRwCu1oM5ypuYqH2Z1631O3EcEkGtqL9BsFndmfdYLdf
zThsl5qQ6XKiwaB7wxtqLwry7FFgYI9ESvVfvAUO/82ccNUw2SlZX7wGP7OEu4vtoI+8ItpfHPRD
TE9n+ICN0yqng7PgaaMKtV4fZh0FNMjdp0rIFLot1HdGAhwQWmCUsItQn6UGwEyRt9lpDtgqVHoQ
yykoJG0ZEN2HfSBj4bN201gjdS0loKtA5lSH34BIPZTFlA+KxS51Qs7SR/blUWTA4RnRdB85qtfh
IFba2bme15Q+mC6PWzjhTL82C6378ra4t6QnByOohg67sQLYWAmKas0FNFL1rkrcrXqaeprQRUh+
aSXXNq+68hVMvMRQmFuYfcRzY5Lq7zR8As/A0xM/UcvgcLDFS95ZtaxUrQw+LtnJEd9po4ZiwrY/
i1JSWHvnnttUtIpdQVd5qmiaEGhjf5FQxDMlUBpHOTSI0JAW+zfWOjv06Jussmz4F1xXqiPUMFMv
uvlsSv6LU4mNmUUwS2ksx4j6k7KYrjw7pJouw4fe1rM4OwUJVNosv1LgtBOWfnOH/r/Hb+wnbCva
iMokXhO65qMMZ5svVhpv0DqidDM/KskfhxMJihIbhckfKS5OvMduv6PA2qHLbvqUbyFnq/KB6nIn
w/lBExZZFZ63nF5bQPDJt9ukAR+jKqBJEiIQY6OwKEj7t93RDoW7Ry7X3MZc8cgyB/WIlvScSBSV
YcryEEPvjC5vt8k3cU4AQHAqKjWYUJbgMM/Nebmh+PKyztYnzulP4/o5aqp6yjOT9cBrVvd043AC
aTJWJDvkfUIN7lC6KlHTffofmfdhQ1Ywy0YT04LnExn3VozSA42VMuhpoa7O9xtx4lfGQMnY+ARi
U0slonkUbGe1UjPM7GHzZ5g5inn+gMzGkQcaLhEY2RJBHH5CD+NInt8PSbRSm+PtDS/AlvZP8RiL
qz1Ooea3qIUzVTuWO4F+1XV4XNaA1T8P4BNxmttroZ+AB5aLVhZtyR26yY5LCvp29kr+6sZGTo2T
0axxbv0NAiifLv5AfrTzrcFwMe3uOUkv3uSdzEutygyoT3E9M+3Jq2yJ7s/5ps2cVpTKpSaG62sc
pCU40V2fiQfF5n52Q/ARqVCGU2iDsKHst2fvKaTq/gy2WmyAZzNN/xnyPMa0rPwJ/5l2k2kuGTe5
xuXkBgWWcUei1gkvRfWEgPuD9Re3lPVI/CbgDAlR9CcHhdbMU3YnLbyxAix2zQthQ1+3doeaCxnE
CW8DAl93dcRu1vP8YI1IvDUNnyNn0GyEEAaAXj7DhjpTY4DmXhd0KxjkhhHXh8V+v/Y/r7OO+Lnr
NloqnqyuzVCUsCC4vcgAseg9VXCDyhqTkOHjNJeb5huNkv7xmHjyK3gL3e5+82HOFZ8AEi0OxCnj
ZZieMS+lhVJmvq42BW1rOSx3cf8qK/KxE1+0EVbu5OfGH0e2gDvPf6tNYVXIh/mSUfyTwU3MTQ8n
xuvQ9iJz8VRaYiu+tWe5Gg0yIRIKPQqiLZDSsmuk3+lsxBvu7Pa2JyJZJAK1G006HgkMJa72ptam
jMED41I6oA5KAUNdLfyhqDIw7IyXrYsn5EGhtHo7jvplvaNYNptt3XfUbzL3ZdJfHcW2kog2Yt/7
Mp8jPglZ9xzA1TLzCsUiEm+48Mv7RpjDILLvWBseUxSiJPR1mX/KjZTD8+a8YIDP+05JQJXxSdUL
e2rNcY95KtKpiWA+nHvpUOdfscqS1dyGtRj2PQd7L4ajpEujgOsxModoWJcqDrOnVC+1VfXHpS7F
834bIXjJMKQ840ygaEe2n3p2J4Pzi+FOiAPePdbG5YsYfs03X/330Vnu1jaxnO/rdArNXvFyVGrU
3rL1hHLWaM3HMR55+ifhjB8tMhcrGmhtYSU2/octD5uj41sn2NrfgHfiLUwEdiCwIJXj9cBcUDuE
aTlv2r55QI/rBpaFkRMG4XH5qaVmPeK6RUDqrk1u352/C1CM0355kUS2s9q1rgmWFbZZYya0Km/6
t42SXINbt7t5uRxDd1dPFAmCRS6OZrW4H1zS/SNWugyBRU6JWoufw7Rg6Whr98ke9vm9rptnXRz5
QGKPo1Ea/xZREEfxOd5Fjgw5hJ8vvfhKwNhWf/0m0WMg7+ZKBF9NBdatBLhFEDvukQtw6eOcQpe+
uDw4TOpymkFisS7enX4Q+UN2m5vEpv7zmUiaOuUaHfyhlnV1/oO2KXdpWPkxQedpdgqexziHc+DG
mLvtsgNA0Q4MNVsHKwbw3Bb/swgDwfQ+MsgWwH9MVxRDbFTbd3HUwKfMGuu+kLVxm15KTOikxTDx
GAqZt7uOSLIzLf7XtPbfeynboHVGdP9SAAPactjbcqh5Dsz3mJEHh0IHXwp5v2pYrvZV3Hoq5y5i
RbVmkSrr3Cuz80wDNMkiGRspcq8r+0yCL52bfKO1c/AFgGQoWCPgmsCv8S9rIWIE/bR/J5q6uj8z
aJqZkOIzvQNEGjNXpv0Ox8oE+T8PhQejbBi1PvcWOkObvQVEK0YwCsxmPCRqlr3ucUtxRwVQVQPN
dzUObnAg35UXr20ad9rpG6TDZi/lK1pTwvynJDOmZvstrLRgkC/u6q5NZw16fFhvJzG5cb1wG1oK
HaiSfCs73FD9W/2T2yL4UQ01x2PZDWlqQComvCzEiK03VA6+Zk/hf36c2cckVZp7HYxa8+Zf23gG
1tIw4OVNPHqmZh5fyNr5QVPcapIJXJnhq8QZgpBiitZFhuta7UFIuQ8Haja0fypZjwVgaYFjBJMn
zQQJ1fniYKhn6adtrnsFwoLbP5WMpoFlgZWJWRYbKl/GFTGZrhDaB/4JhhWwVCMUNlzn/MfVP2Xp
skmcyaNSp4MrexJlxrSJTsegDWR7EAOt2fF4S6l7Iry940iZRka0T5nIG0dyvD1LLULAHydaqngJ
Oq0b2Vo0w3uqI2113GBEL4VQHRQCLEgdQbRlNdMkf2QW5x3ofHOFMw0f2YBQu+vHf/fWGgF1js/l
hTWn/ik4GfdSDwaPyj3+HtV1cos7Zwr+CLHlK9/Ru8B4TcGXb+rxDsJ665FcpWcOha1LgNuUXCoD
5j6oFYJGJ8BOM4jVZ8wnTh+euC9wTHmserRVtMewdsq9T1xc3VDVP9RK1NaH0agOVILuezj3I3Q6
VcpXOBsqnrn5V1uUSYPof0dBayBGUGSSI90cjWG4+zXmTz8u2zzRGaGBANCGn3aA/BLAUJDNtzez
dYK6mU6v18zDPu6Prm9H7PXK/bf28aeWtA/AYYeLsyuO88OqZ9wGIxsbIfug7RyKAGUWkLwdn06t
7pcW3btOUPMGEKEf7+9TCgMUH9Lbk8Td4SXypaniR71ep8dvS7bEppFlwZIWqDZuhKfzPXtiTjRR
QRUcTUlrqi0dUpqJPFaJRUE6ODxQcnaFamgbGL5FI62i0Kqj5zxokO5pZW70xKyhiEDLLbJiUSqC
7k3BwzEP9JM4vv4LaWq3ypXTROgx6vniusV5bAR0rGijE6xsYLxmOPQzpLNA4pAkF9boXE5toFJj
L70zQXknykGf6Dz++QDVoS9MOf+dRxcyN0X79uaYNg0Xo/q6/CYNl+5BO3TFc1a+QkyUEeVrrtfp
VArOfvdBGJ4yLe0JF5/mlYrlkSQ703r1sVhuzcc9WAAeBDYXBMY45loFWTryL4QZwVGLTGd2rH8B
uyddQ6qrb09vW2UIVCnmrFuXjiV4MLu/3b7vDHv9ct76WscO7z1YO+A6lrvwa6FRauAj7nKTKUtG
qASKyglUJHuy+WArVOQUB1gKIAsVrpoPeLwJ+CPMDac3X45v7O+qE0w6iClOrJRiye79yw+cT/wo
tfhz6ewLUxn+nqxrXXwjxpzlLuL0sVA096Jm80XIGxnE7M7etqu6jsnnV66zaLq+iZE2i86nlwPp
yuJSoUIfZt4nMCStfwtpn68A/43kBQbIis+q7+F99LfSQ9U79OINyX1n/cUHeAKu66sU3az65hd6
ZYolA990wzBJl6h+/mAjm5aAgxblkykBhONzOU58WteXtsqAa1KwUq+FHiP86m6DHiKaQl3XO3zr
IlV5qhEd0ylOheRH/SKsXbxC93PjRPYL5mpLmtrtJmbnScQ02HSEYXxwkZjD9OQnWYnGAtAt6eZn
c6vjyRVq7aNWnsUbrgFvjToYGdMG480Z9DwuTJxs+n/ZMFP/vhq50dZTT/+hieyPAq+cFh8l2mYZ
qIjUVotdCw4qsZ9W5fh+5jxsX+lTLSeGXODBVgNaW7tlb4MY/oXlln8cR+Tmz02YhNpVzs2rIRgl
+IEHSwmN/smmNRp+dRZ4r7VXLSTu17gLMuvEYDhbEqz/Op24AK2JNF+1EN9Iz+iR8DC4D7Y9Lzjf
Wz3QPcSW98Uv5N/Sde6SPEWDlgmxqZfrYHW6mFph5qqiVUyhtfZdooI6a/ZEmVfxF10Hpjf7/sVV
nTsyhlW9Pn4GbKIr/3rKMU0zhTjpBxLBuGPRHgIV37U7O6OJKIvUbqWuZwlSvpAGPeJzRLyG1LS6
KFJWXvD5+lnEsblifvk5uQYtAbQr1pijK3aa7QPYo3iZ9KU4mO7RMrOYmD0FbtAqGcm95MUOSQVn
OmFC+4OFlRSTkyBv5qZl3tQ1QCF8D9Rh+x52jz55DGSJS4WSBeUNxnr1iSOZnKEDRrfkIoID3uHW
qhQBoY0Ps7EMG8Ir+CI6TimOH9e3ESnHTUeV8rsSgpreTSd5YGWu6MjrMnToHG8AO7Nuqn9uQK9g
imF8nOxssvmNVvIuswjBZEvTqSfADUg8vRa8PD/e1VF13Hq0pSOOUdjVfNj1IaUR8UyPtRAWnuIW
0qIfQko8jftpKi+e8T7pGGeujxRQ+a8FKvUqjuyHsb2zm7/VYqfOVPQQ6j4KXl1nrpqRL5+7nbmh
omAS7qeKQKa/ghoF4QmjTbjVfs5z2ahyri8JaxmvXk8x9Rkc5b8sN51QajbHJIiiacQfHlIPl3zG
49POmfJjjku6sXPUk7y+zTUTsX+RyhJwvkXF0TAQaHoZw2xDoXi/hq/HAjNeKv2+mjlnfLQ8/ZLY
twdPohSOMxKPf96NNarWGSWt6E2s1S7C/CLYX4lufoh/+1CQi0dsuKkye7X+dHkW3bTbNmMxA/9T
oKzelK0PDupo7/uoKYMboGHRdUl3G/pjCfgXk5QcJ+mbA99Z/zq3mqrQ/AX1AE9GQq1RqVWhEpUY
AHe1mmsc037MyWqG+NG6Wn48SmAn61bFt3TXhffjj2fIsnkROAxgbn/Fe2DKilUxN6O8Y1jlfbUB
Q/T2nwmtRJeS2zC5bueVqyR191IVKKm8E9FVTksKXBGPqIyu+aW4FEJ53ViT44j7oiAMifLH8WJq
vVPSBIS5wapcgBOqffW6XQW+SEM58stnfgLnhwbnTuwcHJ6HzW+9S67JdNVhOIIkqRQ8+dkMov33
nOnPgY+SRt4jiO3wqsKKgVFwFZMWMZ6enLZZ/V2MsDHgckyqPs8PKAsymJ7SCxiLh6Za1zzAtq+7
7WgWVbNLo2u9TyulpvQqLR5p4N87vgueiCszuVgz5FCrGbhmcuTQdpgR7870o22n3w3gVljI+gbZ
/HvU5gR0A69kO8OM3ksVJr/5241zMY6++m0QUqhtwCu5v8GsHawkSkQy3CFu6aFbMB/+woOaGUJq
Rzd7bvKlvmgw1wlEodTmnkoLscEQyhl6LNKdsz4UvgMtgVxOVI/s8Cm7EunFbGfNhRCKm5XJneRy
yRYX7qHLIchbc9j2FrWnV7C0LqMrhlJS/oqpcSm36BvyxKy4wibrlFBIl3U3/u9c5Y+2fz8DcJa8
I64mbECjd4p0N6sd1nZXPvj1UyuYRNLI9ibUxJFMkqILJ4Rb6vXGoT6spkJ8D+ZX35bCiT2HVjKn
iOcibO6Y7wsm+ZEXSLybcOpbBSAMgY1aETmHBzUCvwP+Iv2DlCfFX3hKllJxQ7nn5pMeMn/NVA4r
LervBFYN9SQpyQOsIurkNxCwOZ1ahfXirNNPJOJIXKHdnjCzzawZWk0xzn0aWOvI8sF6+9KusKv/
WH9fe5a6gowPo0KaV+QzSMjzIEXdI49yBwiCr/8hTtEm2ttLQbFaQMygeWTqk55MxsmekbX18OPx
UIkxTR4/ttv7xfGLUX2W6onZhcjunLIRDyj+Pakn0JdTczF112QVjJ/uJqsy61HGK+EuGBp/9XJ9
Ev59Ew87hLNVEXBQ4kQOAa5dLvDj+6PG0DryQKT30OSpH5apNRNAgl5RdaVGEv4Fe8h6i3jieTgr
1U+uRok7LnB2FoF0nlX354naOV1nCa59+EBc3Q3jhFexTM6OJXzGOSJdU+0MZvXJrydcbxacDlq8
erpHrwGPpYIb0Bxrntv4n28a6ycpZRgy33QojEySe9nMEOAFlYs0jylufsB/EBuDa5A/zLxIk3mi
hywleKFBEdFxrIO/cAWFXejSKvK6zoiHZA/gaZNP1X7aBoX4bAH0s6jBTXaYONqbEMflrBvKix4l
zQ+KYMDBU1yMkrUSy7pcEkrwbFeRtn1oP22j9vk4KhNEetWWzRS6SwtzMdbI37B5uqxoMnilJWZa
ewI8x+Mk009yUoXeLoZO3LENFrXJ92LosObOL061Y7J2dt7hA9uCmeXybGLFo8BuERRj2a3A/68d
3PrPToySj/zwwfHggt6BY3nLJrymdYBrTahEtzGfztatea69cpz2OL/KODvkyDstIQs4q8v4wbSl
3tsDHHRsnGAZrI0/ZuOD3Bs9Rao6oLCwz/cTSk9WJ5im2BB/CSFSe2M4Ia3U998ArbekAMdem/xZ
hwq3/AiLYnIaCuleRdF7fxlp+lOuwz621g56y2QTBxBgGmjmas7HFv5HQsSHTm33h82rsI/oTtVJ
7cyP2yT2tWsbrUVY8yH/ZHkD+333bU0DgPXKZhSYuqZN6n2f66/QEIHa7MFRmkqWpMpd6khayLkv
QIKiFyTRzpDjz4nSGasABJey9OrTATwEN2HHTIBWW7og8u+koNoJ7ow6iEybjWyUyny9gXRCOvx6
wgzMvhygOrHCWoh3Ct8MP0RWYMZFWh+U2gdHXsAfzgtUkM09YOeDUmqnsPhZQYwHtBiCFWnuz6Dm
t/3isYN0jx8EbOZ7Odos4+puD9MXZStQSzsi1GD67NgwdJdl8+BvIZSUgbPFYLmS0ZkfZhMAXXO9
8BTxGLH8NdrJX0EDXEVaS3wOcSBeCGpqWbiWLz9m5YPy4rA+caz8+IqyiKExp3Gy4mCSaCr5u2WZ
QWbnQmOI6/FYig0tWzLabm4K3bdI+fhjkF1naIFfOmeebAk6cim1qLABB8X7VmWrvvralN6hFd60
1O+7Zpp1/KdJorXU2lfpcmO4vIQsa+cRm/H/aCdJ5xYWvYYUyPsZIMy+tvjgRLpxTjZJQXaR74g/
++enZA/3ymFPVz6fGeh/WGB6yuxMg0NPkoM8Oj/ixOjc3cdlhL77jMlA3S3ZJHcrdYLWamRmqIAl
HSsJRyPHji1xhX72N7vTzU3BtrYTbqpAf9XFYQW+5Lq4xKTkXL/u0XHlbVWxAB6or7051cdgHTTM
2gIyH/kEntHsvyo1wfvVfebw65c99YXDz1DSdqksIwcBi4G6sYSt91EWFumHsQHLbk0Po8jcQjdq
oj45O2Wiv/0aHRhs/JinPQzGc/wf28yXzVCS2WK20A3BjX7idaBnJ1CtaR/jPiK4MTfCNW8RQikM
KZl8KGVtP8vyx11JSBOqlK/l8okmCxzgMeWPaph3+LwvBvtUUHYkbu5SMuP/rIY9BL4iMlQeZeJV
pcDjyVzvMR3LXEoyqtZxf34KLMUfCa/tz8GKG/eYvUwAAze6npBRmfmRrLwLe2fOW0dR8kNxSWNM
RZYAhfEqJMctD2lXH7Ad8tUFKzz3F2uUuTbPY1/r1WkcgrCVnaXIPVmvKshI3uU1knxq2I+A5ANo
mgBZdXhevQ8zzrLTePnHlsdXl6uMFD57qe6DACeV1Cmv35+7CzvB0EaVGkCzihOHw9DzhxkECPm1
2Zv8mOD2NtGDhBGcutrZ2GfphKMWfztXDWND21LHBzc+diaVQbuwVSXot70uEkwtwh7bgqKLZe8+
t8lf9Fq7/5a2ZqH9XOCZKzIvoptdh9owDlZgCNDRu8DAZ9zV2H/nFP26nprj7aMiGoDUJCMV1fwA
IZr/Z7k6G4B4UCe2XAsFhFtrtoCz2BlcvhIOhWxjn+5R6j7drcXdwzFlaw61WcCf0SHcOrkUVGje
VJb3Wz5RHkvJp4gtBgVJLppWuPV22jCyDr+fcJSctJlTrTZsohSwWHln4ZeaN0mhIXwoqtlCqmmE
4RgppNEAE67d7a47MxRbgyp2PxnOvW9IKo+mxdgcPqXfm1SQlctXhZ2sjfZ67pRDOyaBTHyzcKqq
f6MDYXL/G3EaXU+zwlyChz2V//gwIz0f87b7f1hXHXKoqskoybQwl35RkO6Tb2enFRTv2HcGaI5h
vy+FUB6vZYIVvcOatcOejjG089M16okPio7pD4HdbawQRti3T2mCHYJg+VN/VWfa+Ae7XaqpQ8Kg
qOFKGPTpCmmuk0bfpjr4RO/MYVs8THjeeyRSrwGQ5Yf4x5E51RNW9z8ezKHL1RA47v1RB6uQMf/L
AH9H4brygqPLbam7aZs6qidLYy+ht6P4lRqoj6kYJ7pZKCtVOai14WexDV2q6lacAeC7jlnzoAkh
BNv2f1XhMqPJCvyw1Maih5hxmVCirR6eFHr26hGKwt2QVgmoxt4W8ItJ2W+k2uia+/ViEYBAQM9A
ODEdxU8LG3CNPl4wKUz3OpZEPnzaJUt8akuiH0cMSM4+kWnW+VKShn+fbXOBZvC7DNKtV0XqPDJb
sgfFdMezTvpjuuKmoRJYG6cSCw/4+JkMHDd/vA7vKOLMKEbzx6Phx8Z49Ja0klDyfv9gr3EKL7+0
kt/a2SwY2lK/0tNNrF+FYbB5OZrFDOQ75QJT//lhIPT0DguenE6emZHjWfIk4hWHCbtJsyx7/pKP
2RUfpnGmZB7lJeRSDlV3JgsDlK8tF2aHFnaiueE5GKJbsSmGE46XQ5hXZJXlXsJ6Y7miP9GRLcYX
Rrdl1JWXG0AFInVxmHcNYACJtuQyW3bzEndkKfYyu/M3BK3fpeFtkZfzq6AdoqeiLrDa+TyNqCNm
A4pXnmK3hvp7qDvqDw4+4kX3YB51wMSIHv3zq4tz9d25Tejek8rOUvFjgxl1TE5nvV9x1z7Us7+j
r5IM9KtBDI46kcfukadelG325svHjPZaSWeL5ruGG38BYSpsxODLRbDG2zfaE2VRPWWR+NE2bo09
AzXDRCv9UB6aOL+9AAtS8rDElt+F1eo872kgpWypkDQymmxDhFTZ8kO9H5tr8MyN7Gg0bB770ElD
TdxL5K5FYjUaFVEi7Z7RvFWur6mjhtZbMsejoGQ3dOgrQqqlSPegWaeloDP9uzulVSF8/YK+PeNJ
veWgA/OXxPkhxOCfKmYiwmmmp9w4ICa4sMCpiLRNHrWkWa6IQPFKoHNkU5voUwxMNgN2KQA2+/jr
WrMXxnKRH2DlUd4jwh+Ve0545gFBiOfYzOrmYsrTZpda26voDWQFNqKWJ1h22d0q2VO0G0/85+BI
RJhfdVYoTfTzByaWWOIAtSikfBn0Kwg4VSIaBPSKv7pZ3gcDsJD/gfLUaW8qByJnSrMlDKk3yLNs
w1RhpbW4jvSpsOtmgZqU6BPP2+OCLosdI5mAcuK6t281Yt9ga6yxfU3375fusnq+XDmWbzPeTh1C
5xYIF0OYez7kQ+Qv9DXbVFCnKgk+8869fpZoMs9bALK+5iwlVjGPeqJj3/nL9kT7aM68FefK8Xtc
MQy4iHkehKaJbCWyozv1A6S/zMl5RVSdAbm/GbpxSDzGBlUwpDlYAKeaENnWKRYe+0UfIDBPy3ez
Z7Ra43aX/FVrfTFPHm+5oZFgtnjWE1ZzF7ehcv2Bc0m1OfGLvLUzoyFy+aWXFMojZG+sIfd+qqAR
3Z3FlylYoGl2SIrLpVmLChABhlkw8ePNLOWO1r6SYqMbyBfC8iQZ/NAjHYOqZ088t/dvzf56iFkY
NkGNJaTEz2Dw9CcOp6TrQLxMBLt0mf2MnPf/oOuW9MDdXc5bW3k1vQNjYnyUnI6HvP2q8ci+BCAU
f5HyJYwvWazqWxgtbOUvtVvpiUhcaRNpXk4hxU+iZGXuJlm0WIwx1aEmIOOtpG3duOahEeRqKY95
EOGgMWR73/hNoXoOV+J0h38j/OahZEYbhSi/L1c7JEaxJ37hR0p3xH6zGnszJCT2HGnfAvrzEskC
5hQZmxu8SobHQA/cW+q/CZ9D4HJcqU9amX0q4q0Y0wtmg2t+2nkBs1hXvCWd2RORFdBMIJRARGis
xMEVyoo2faJDyblkrh082m1uqP48BFMOQJlopv882BCtsPDAwtocvI/WxU3wZ14nHufIgCzOM9pA
7ouo9DIr6IWOCYHuzqyg8Jvxty6/K0sTFZk3UtOuGjhk+740R8Nnh6nyELOkOlp/5mAxsXeB8eeW
OwBNmwJoW0sLx1YT1bldvd/HFnFKjNouw4WOlCVv3llVFOFa5KPa8HuSrAaovGgD4ZSbAwq58I3l
lLhHD1BnugmHJv/gOhk1r7wQlAFimD+ZERG6e5ABGZ8ktO5+2XW3o/ZVDPtLdNpGrFKHIxB53+ZA
1IsZO9c5malz1gZCKqNkhe7lKydLAO6r+vIkFKOvwe8IBKCiQUC5kZJGXkSHcbQ0RJCfGU2abySQ
zrkQNctGwTZoYb70QZpWsulLQQzGWLc8Mx+YT/f0GUcgB+YaH0ZiQYyAoBrfafhd48kRSWw+qkSM
08Fl7m9cDQLNC33QZOp4eZNzWtEEr+3a1Dl+c+DZoMqw9txHCTwA164u/bBZ+oK3JfEQGUZVQX5e
fgx33paKsM2jkqPDv6uE3Ha++gC3/wOZSXi6MvQTfCF/3s82CDLMLh6ZE4Gi55Zn9Qlz7ixI2a6E
2buWsOdpcCNYjvTkqSwMXmm44QqORzpVhTF5WQaRvDGejTYhkY9INL+C/V51XlYNNbFdUZD+GuYi
z+Lk7l4cQVS9D39PV2AdEeKQm8unD2BUYXYrgQEkbr4O6hYcQQVrMQPQh/gQ72GyaQbyrCPciF+d
pc311coTWoaEeXWsGj8D2s2RANgEwtLAh1aAzo5+J+JW+QvbpFZogfIkgJG4AGlFHTOGWlgiT+/m
jIxGkAUmkGdlFzp+UlYePoB4x1l1PqaWgPL6buNjT/kt3tgZJL6Ryyz7rOG3ogr3zsqyiyeL87ad
dFeLNXh398LNdwbrsnzwuDFX/gVItNZ8qlELCohS+PXad/dbZdhOimn8feSLNC68OPHxB5iEI+NR
+Z7Vj9g6czN41f8APiFYOnZObC1QZf65DuJtGgYlKNcmAPNQFPBTK5XnIYJm/zsOirdnUlQGVoxb
AskvWfBhY74/13dl/4+Z4c3Sw8OKLBnE5Jw9iz3XxVZbbcc3xdhOONeYFqO5XYdUe+gHjsqs51KY
apCZDGMgJgn/OBzFmkQ6OOSlekMKRGqMtDZKSlguxujLDXf4vdnon9deoLOG0QZA4jLqVrvBVEgc
hpRl+pHH6UwBJO2vG1k3ApKF4GLt+mVhyvSAZxFNwuX+Q4EBLuNjB4D6XI6B6uYgx9JCB1zyRnc5
nYH9Y9rmK2PTnEZZ7xd6E8FsJ3rc+MnIMFkeNZeJ5AUamSVCcTB39z631XUomrlEU8Ycea8YoakK
3HgnrdIFNsU33/Bbo7HfqZqh3ahurRhnSvOL0Wfnq7lGfFWJuHvWbQ0jQPQ6Gm5/+R1xPAi8LrOX
Xt8hgSF6zi1VRGS2Xf8BJtG0wHE2Ysjj39n1nzeuRRT0usDEVdt/mCDfsdhbu/93DYEgF4A0hPsi
wZ6ZYo8MULJZdCkwLwQMy8Km8sDFfBx/3qHXtsyw9gJVLhHJ14/UUygBIdGVjC9Wyu+zXhfbvcFB
f8CwQx+qpNDkKGAKNOpBPckiCASZsCZPrkovII6EnqKcRJqqbonT2cGlludRpq9lf7BRbWGcNff+
YnWvlj5oSl7W9GujXmO4b1QDvZ53kBJC8PK6BlAm4E/B4zdn7z08OXh4q5A07efKvyl2FbfI8KsG
86Ygpipv3E2/dOz9Ji2qfaMq9UXulCBqgv0KfUvLTyIIQNiWJ3TgmFkWOcsTKkdF6QKzzUjTAADW
xmEZgCpdpDnBTIxHKadAjhsQDEN2YlI5XWKF8jWZxhX3gmVq8wv5+XjIKBdsGj1ciEVW259N/r5p
vbr8OsOfjaVS5XRJrYillzyPK1U4rWcE08wYMk20tRZGZtmrJHeeWttkBbbguhuuU6LJkAZN2puk
yMrfnxZOGBwf7dLZbtdvs4nFIOQ3/sEYYrG9aVwxYARaUd1E3fLTJqBtF5L9SCGD0wSZhYkL9gR4
olZBoqeMP/tbe2REjJNwXeXqJSD+CZnRpGh7UsfaFH1HjcL26w+A1HDM5ouw3VDVTrS0xSrOhdHh
MW3OZOmzL6dPybt9vJBjla9yNXB7St3HCkBGHkmqZh1j8VAmC7mvijuzxyCxYCQato2KGPZuTzEI
2P58+ebAmx3R5KljD30cxmsXDqOk/Uj6522HVU0eFQgS+EEl2ypK9xE7Ht0UUcsKSLNjwYy4VD5O
T5wyAzyYLcIg6ashgu4t7wzBVb1YTgd0hXSy6QTmYS//4bhRh3bWJG0+xW6w7XOtM3NtNrEA2Ddb
1eZoVNTOHhtzbLPa023kgqrBThq+3LVNibqqytT5hYcgfRbOJEXE0jCCEPRyWFG/rr9B+/oApRLs
rCJXLnu4iiP0uabAQBnIbc+pecTYp00Lh4H+3x++ROnbHS+tC9KDr/3kvY5zL4cm7qlYw/ssIDI5
YV0nYLGLOXs/e2izfTfdW9CYwpqHCzfUVFnXOslrlP1nSUDk3TWo0xQ3F1aEq5jQmOTPcKlM2qf9
RWCckrv1dv5g3fHrI41jzjzAgyagw0c0EVrsjwSLN6We0sHwmPyz1yWiT5q9wjBVl8vs+bv85x/8
9NLDqh4xwke/ZvkJZa4cBk5Fx6m5z+VYSJ/uDbwyESISbRv8+l2fdhvtHG6wmH1tDqLJ1q87a0kL
+jJlAqhga9E9VjVvy3+5IGiehAIuykfDNWFbID3GA2boj20xUjjVgNY6KMUkYKSCul6bWx529hXG
0IieetGkc9NCY77rycs6NzeBOiPmE37PMypVybbaFfitAb8ytLpjSsPqT75/2XKPieGPWrh9wLZY
gAuIMN9TI1ksnGIEnuvx4P6gxcn4eZGyMcsKlnyKqEa3GkbPEHAdWW29E10NbPX8StyIotvfrl8M
VRFnWt+zSxgrbG5eZNmnWNxEbRTP1SClHuqqeHhfc+y9Bq/tCPxVIlGYKJjTYHrvqPGLitjHc7k0
d4hp/C34HxbwdigbpLPItIfT4VntwkR68anlQjbZ3Urbfg/x02ITym8JqsMD3u46O4WjperYWJWc
mo57+LrhX0C9pasMfeO8xFHsDUsBtOVZ2f5EHnI7ePFDGmlTSZAbgiJbBTgOCpt8ubhUbFEEPRxv
t7We3t1/wEBaOm7Wlndk9ViDWEfAY0OhqnavhkFW1dDaKzakxFjwowD7AbRQlL3QsWkD+u2f1A0d
DzGWeipEO1F0zvBYx4FNH74YhHGJjVxxLuymmztL4+9mvff9spiz5f1x3zBmeXb9LD4zFQFKzdyn
7k81qAGHDYuytjrg/idsq4hZDCQje/BhBm3o9qfhIrNBzkvXr3kPPhdeESQEdLo4SVF2in1hMQhO
+T3qSjKFUhVuOGZ0UEtbSTNu0ooogRPVEFRP0Rq55pMoTq8/HZToe4pyKhdYDrtwMxUpO283cdcx
DJg9GRlmmrcGbR2yMHfv9jBGs8P7dBNiGxHZ0rOEiCPe585AWs4HrSfmrpP/LrE8T5s/k5W+Hc2G
O78Alz1WS6VcigO8gQqdl25rEdwvuxXclS6rM+ANy5msu4jYElA2SWOIH7z1+3K2NHnbvf8yyuK0
DHE3nLfCM/YO+Qf1lClTHdWMO0L3C57gmXtZK/BDkGMfAIyxKzbxGQox22T3QwRYoJ2F9nRFnhtv
K2kHbeLYsg3856ZVNwAwUNukIdNlb4yjotOA3JFCng1x56yI/bkcZRjV1LEkDA4h/kp//OxOZZ7s
WW5hFbBjwKf6b/jXochf8YSFJU8lQ0AUTobXSlkBKIxkauKAKW8KfT+oVil2Api2Vjl81xZ5mMS9
pSSPKrffiWbM20DGQZxdP9bYfaRvPOxQhgxbFZVPoeyg/tJKnlNTuo770Lr8IlPNAdpENhf7i8Js
mmdyFPxh9N5VlOS/voE6livu+pwOowCy9ce5uHhd/xIqf8tNcn8iuySM3fTg5aFaueh+tOyOJ6NT
PpWvgIsCrlc5Z7NPBhgUT+NO0TfRfuPY2Ef6H4EC2sllI43tcjRUINS/svPVDZ91g9jkX94NzhFK
WwKVBehuU2W80uWIUurZrI13SqvVEd+LB6TZouoNFXxVD4W3Yl5W1DqM2qidwZdE4HUpvHNhpqIt
iv18EdwYRUL76SmDEiHtvqE4hEhSTcOqcz3Op5Ws0AuXeZFEy7GQh4OyrBrlU+knI/dv/ZzjT32G
5yoZDiDOVOg+VoWOIw1gl0FqtUZc3JeXrwqlOvu4cHIzDk81Av8TwWtBxAo5NXh+/Y2pdyIHtyZO
DfxM46JiIPIPpWDl9CLIIjOGrtBMRF1I+lhYt/7u7phLzRUUBPlAwTQT1OTLGA0vfr2HATMQOg6w
+tDOOGySTx/grg1G/aB0Uqfy2GTYHtHDahFwWSWqJVAymWotCAaY4ooFtcCAHt3nLVYKofGNUv7m
L6oh2/5ZLX6fISexowVpw0q0dcfHnAIjINt9mjV52ACysRM5MFYEL+y8Rl6VjROxIzlcsVDySB3a
GoQV5EObRSOPvgpecrFnwoaOoTCFPG/pDz/fljT3yTufuuvdTHDstDgIsdtYKMoGJlmPW77bCuu5
7HM/NtRhcNYcWJKTwcscbdZz1CU+eUKWUMRfpeC8n3qMtAryMBb7NZVvm/uXiD6QIOYyMZUBzSKD
5pJBS01FXjBTK6ylYWPNPKmMcz3uLvWomrgjFAMuP7CDxwBX7i1LVDmAaw2JkkjCjuYQd3lQGw53
llzJv28TH7We/xVSPHpa3GBpjFsKF8jinV5tMLhDeuORL2ZC5ijYDOZ0grhVNBySr37rPYc+wSPd
8Lb/Tm0TxR1R7wRF6R0LSEBSQeQfY9dHGnHT/IURwjRRRZi3Mz6WnXWWt8SO3t1hq6MDRN2uxm8Z
YbBwSWsbAnQaz0YibD0SsLcda+eUhdyT6TNMN3kEfNsO2iJjHOmerdUAKs23YsS3G+Kt14WB5Tpg
SgNjxGd7Y8b9iENGxV+8mLFTCzPDMXLf/0ocTP6/93zV/lwuxFA1WgAADZav8mWxH61YdqPOrM1A
QvqaAFZPg+y3ll31hKaoQmRpud+dGAbmHeVv5t7djF8ohS0iUcUomn1EZPcBBz7XhDoPaRu8EzgI
tcLT8dFyNtEE7X9k3hm1aAFaFZK+Lg0eBrl666ha3Qo7MGqREO5+BPCDp+ILN1iFTR60UTI1TSyn
ma+AwFVhz1t8xA7IwFo/coYh9RZqyWwGN1njR+eVFGq3Y/YwREUkVo/cJO8Jph2V2bNYUlcu3Hm4
aeVxwf06Y/MbNi+wUnzqnmQHMiWbiu5oYDNNTACq4lAzzEF0GpcG9tv7+6YB6ufVmfAS/n8moWmt
IIGvgVkd4tdXQnjIrojrea/QaA9HmBSj/CbtZ6uYgMBqhxTKqV9aqZxq3frH0vLwcSLdbm2jxzWZ
ut8H5ccE0V7g7QdAffvr5qs2uZsPQrZan8Ch2WTd9piiI8gYoa40f3PTOqDZr7a1snirs/w3xgfv
vHuSwAVDsQrfnEQr9JHUfd96icyvL6oRKedKCsuu96MOooJrzfCB2ALcbqaUAiwhim8+GvdA4h46
tyY4hh3WfT4Vxmo3qIuwBhDUuPyWIFSaVAD2x3U3mx4Ab7bUNxxkkRXvI4KXM9rJAkWhV4z8Pqfe
0Nts0MqtywQ4jbg+O//RYa4qHGdz2M8zxZyWxrsyertADNmiU5KeKLr7jjBz19oCXyLnPSUtEbMo
qHI00EZ8ZHoN8EjOx0mazQ+uJhw/XJmFBwIFXws7Y7vLI2C/Twz8j9KpzdKnc17Xl98dvHkD87N7
1tyWTJZm8QDQWyxakap9GkOV8LMutY+0Ofi8Ftd/YziVhPfcXSSde+bvjKQitLemZBLfubU+2kWC
A6kjoQtYWNMCBDYkXiYwYjC/nZxb22EBEbImMlYYUeFgyTMCNGHsVsNj7ONLKhhcvOT7vY6LZ/ix
CZr+kDL4LWlKaY4M7W6Pa/ZdqIDaQ//7p4QhTUFcjq1Pbx3/z9UY4HKLLJ9m9pc3eV4bMd8p54K3
9uPBXb0/vW3BHlDkgJxC+uAtVrlaEbhvqU8nK5js3TtsmyMW5ZwvkCjhXn+QR8IxW9SQBvRiAIYE
OTl40QWLMoK3kb2BSj6BX1WHrO44umG0n6q5dXmhomlsttaV0Erafdwv81PNqCOc/4IW6gWQYWpc
DsaTP7DFTgHiRnOmuxL/WldrIT9hm/5uDR/NrYqiW3ne/3DNos1q9xnsclROnQUGbJKUWAGK5p1E
TZu6b3sR8/tCrA8TAktcksg7KPzqvPSKx+Fbks9Q0XLTor3hVPwBGoiZ4NTKTAIGvNClKUrytiM3
4w7ZjKhdZKw0Y3xbGco8qpZryN0+G/jYc91kgdYZFOERblYY09DOfiEZ1/6EFJEnf2iu/U0dQqgi
UZ1FTQPg0oFGI0Vyo4EfnCb8NBxGm7MgDg90IyijxdvmkhhUUwnv3nEk+2fs63baz5tHCXitGOqA
x/W7wnpWPsk+spQbKRfGiFRYF/3+7BJ+lbnAy3vTWVAzUydSMf82YRp2rmCSEmRaaJtMXp4rJW3t
C0NXVS2f3qGCJpxrxiJOpg7mj+dXByr3acd10RWr+7GLXsxE75FT8IBDDe1clKsLsC5dgqPoOCm7
/xtADfaC3ts94N6AgdrSzQkt+UrWYpCDeYnu+U25rDjO8hrv2NIMOV7eyUw/Ys9XPsp8kyfhMqSY
gGlYQFqWNGg5hr2jgG79NXjiT9pBV0uH4l2V7ubh8m6/6Z2YPbnnzjTLX/AK/d1r2xFoHfIOXi0v
UuZDb1TdB81aj3JZg9RH5NHQvPchI+niz4Vb/GgLWM2UTgLDiLpVARVdqSt9FfJCqoCVAbxD6ugb
dB+iXiL+qXKNcWOm9wfPupchMzKStzIlpnH7MJrbrGrYq3KnXcyiNmYshEbyTEOUuIAmSQuth6aw
akYYIidHdcGP5JXq7o7ztu9P/EqWh+wT8kn6kQOEMbwJBBuoNwDP3kxFslWcY8wlmSdCxGv3ma8H
xlA7r1+/qNlgr1Bg1YKDYUYYMjcEVy6aKgBXmipl8XalCkuDYCLmn11s6ARwEs7aZmOLH6sul2gZ
eHWl+wR7Y8TQGj7P7dXPH36kTbaVJ7j/1Zd/bPqIP7vz/WaHkVDcNNk/daqcjZIK7zshDPqMUDAL
V2JGOnrKbK/9EX5uM3ieYNCX9B+u5XOFTfULTOq0337Ut3DRWlWdVqw4fvXQS5oFqAbu7V5LiIlC
0kMUMvOTnLg+AC0/cFDw68vxJ/5/OGwk7GnL0QeXD+VxlVHI4dz2iO0s4cGe/yvbGex44i9NvV91
RSHdCN0JHVS0mmV3fXxTZAedOuOdUAfu6UL4Pl6kXRU24TCriMV2tAQ7JCboHN7CVSTdgW4oMGsw
D5r+reJ++a0oOh41+d5733B4Mm8fiN+F2WI28vFfwcJW1CGHtGc41EdjVAB7OwPlVkxzkmgpqI1H
stowlsdKp4KTNE7Vv70M+dD4RY7XWyqEkX0RbZkNM2n1e4GPSn9ml7SIJzBoaN2w4nXcN7hOcPqZ
SAhZf1muah3DLtKdjOdnSLs8N+g+w16o7FgAxsUeAKR45o8QLD+wti+UqapqTMM3VZwM4/uEc6r/
IFqpx3K2ZwP0jGSa2XXFY5MSa2l7T+FWT+baStQMlb3/CNDRvflsnvFqIjrGpJZdGiNwLi1SgIrc
9IKwZc6eupRG46VObfkhoCqRGZoXWASh7L9RuolpVNI52W9rYXoylNtuOfCtPHZxEnvjEfzGsRaJ
SBtzXJ9d3FJXtHR8WCohyVLN6ejsDCSLriyc96j4t/Va9z1eNW0mz0H0rdHL59vRUeNI8whSzI+C
H4vx2hsXPfWSOJWuXVIx5fs03g21/YlPSPCbT5nbbjzp/sDualgccBOIazbO7yQubO1vuu2aFbwC
QzNP6sC4oJAc6q9uSGF/hSLkvTWcwhvLu4Gv8LSWiOV79ql+nYBNFrj9g3FF3097pC5d40Foe5gB
KRcQpsDWzva0JwQmQpYj3ghi9cTXlAPhTH5vYut5SeRBgosAdZqXaklUW0IqiqTncaogl2VaHwRe
lEKYMkZo2ktrOcN5FXFT27rJvu3SHsLZpg6wmHfa/IW9PZsq2mgMMYG/m75z9p3RddSwN3tDdgfn
WaDsl3zxLHnNmQ+Forjr+xnvmtzyL+XaUK6Id1M7GimVNKHZgBAKUc0nWzwbyoNvAKVsIX2BHMIL
qBqRuFYWRB9Q3WZegtAk0SabaBOuKSlfmUpRdzvgIBDcMIy8wh0qwegFwVP57J0eRbsrikOgYGcx
5Z7ucLUDBrLDyNlGRr6FtS6b3mCBJuD/UB/0YeXtvl9OGQ6yNLX2R3FF2TIdYG3zLUCZAeMle5AQ
PuKtDadnHHqu/bsmcZ62Fp9NqZfHfVMgpxjNlMRVUOCJu4A8LIf3N5O3JCjTn5fmdoCWYvAgF3Hq
yVpkm/iZ0zjBnmEGINxoCNb/yTq4nlFznn8Cz7l6jyEZ/zqMrqzyxFgyPIGeyif4GkYVGBM/D7Nt
I+XyzV2IHrAZ0OzDG7oCcLe3NzQN3zFjsHs1bP/5Rf35l+CpSFIqB9aMrohILgwrCjjaCopq24Ph
YJ3XJgV3L9qLCiQRokw0bdjNKcJN1hiI64NJQ/x214BsTWbe0fe06TzPVyuDeA00jdPeLKnlTMoz
mPq16+WVxOdeS1PPWt21uFFp+IzGjXi55NLKpjeUh01pFz3hAYdZoZ8JPpWVHsx4WL6YokKe/9NU
+sbsMA0eP1M98ryLpnMc0BHs7Z+nUcjpoZfethKKSQqTWtmuNtKoKEiWmpUgNB1QWjN6QEnIrdoZ
q0qvNtNya4i7BRqgvp3G59LxC/7NASCTSbMoKcOayX9w80Djn5lWwFVFPhAC7q+zeiW7RyzJqisJ
2njzffTOF7ukxMLpBpYimRbL0eY+UsJ7o+U72Yo4houDMrN1fLoOgwmbZdhTCpUvsaKAJkygaB0z
09klFntbGAfQR69lEicb6NH56vDZTHCp7Ipykn40wVCP8QZ+Pq1L0/3+MiZXGqOI7BFwDvvT3XPK
n74a8cLXJDtrXeiT/dwcDW+0CbxODtuyUfrxML4mXQwnfM5O0W41uOIX3gGqVXUGYbuK4K12ilBD
KU/BPwpMHE9J2G9NJbVuCbKlkoOi7/X7kuAgeWVvw9E+z/axiClNYBvhbOy9RVbwLZHsfLCO8+Wd
t3dulVH+cE8Vw/efyzQZoF0ArjyqbgT52wOIjAwgR5wR9us6SuwVP9xsCaay+2g9QY8342CFvS04
6pfdgIkV7AcnDud7c6YM/QR0N33Q5VuV2Ks0kIk1BEU3jn1G2AEFRIj9iNqwNyNUkW9wDnBfFqYZ
zOwyfGdw/KpZZMXviA/84EExQjR1KHBtFmztqlRQ2Aa6OUIsNlz/oFiXqX3n54VRWYzpoSPpTNpQ
mi9/EPH6T5D6/obDSrWN00zOZhqNho/xvDLZMWnR3BCtgJImPjilGVzSEWdQLUB1neGvKnJ8XCXN
ssAu55y79HO/qprYMWYLLzY46A2Ff336+jZwf1o6YkpVuECyf1Hnhsz3rnDNPxql/7lVW2HPAOrC
mrAZmaJRE12/RTjkztShSYQGf0FCSo/Ar8NKSscdTWCn/SKzdlc+hCXA+IFlHJDEaexf723Jpjq/
Hv6lg4XBFOuyUb5lwh490c/AvrZLNQslToXBVJv7cpMnVohHmR/dZYhRy3zmuLzYqjfiFJWTBkPB
RZ6lg3ysQKVq27SGhxjh0YFv3zm6bSnbDjHf9e3hAXOiyPyHPvozDM7n9u8FwNieZJzzonSQoMA9
UEl7p6tTCh1jn/r8RyAh053PRSRf76dtWShD1QD2jVoxDd1GsNrRUcIBGZpk+jRyvJNi+4gHbeu2
aQANjEGhJI5pwTd+Q+WVFUdAhkglpG4P6AjateMR1oYDHr6nqia+oO7CNMPY/7Q/pvB+4C+ExTuz
M4QGki3wf++fcEWIJJ0Hi+Dy+ALwT+Lltq9UL06QDWEmTG/E3KEXXhtR6ajwHwdLEfTDAHi3YDmY
qLiUwdHETkg/mWxpXdbnbC5BPPCScccXTrYOkuT00sQ0dCZ1REAfyy+XF4L6noSdswEx9GdfZJ2H
a3mOk0NgTq+y3tGEdwRiJkMo+UrX8WepCyfNZfI5oJjy4S01Ex4jdWiNvONHgZqWYTu0HKZevY79
VZOlBIlJRHWHW+fW8ndnt3nsPZ+mOteiFe0Oh7f6K8TtKLV9k8qgUjaTt8+AKjnNNpWg41hCCniU
1D3LhoKG3f/ZMeDJJD/+s474Hg3SEnioGu512rMsu+DFXOo/gkbEkBMES0leiJCnQZ+4pJygxrY+
YWfW7/cTQNQ2RQWj2OxZrCIRgXsG53aA4Sf7pinWOuvo2qu+XGGh/IsyVj2k8TTSVjezrkmM5dj4
YuhzUzMDEa4HXdJPQt48ybtBj92V5G2OfWZEJb+Ct9Hg8mA85LkSm4meRpp5wyfc9brq91G/ybXh
M70MZY++WXpY8a5FrgrLvOvXUTmyYVlnNZXILC3RsTrnIMMXLu1bDW6U133mZfXI9bjWqRDY22ZH
GEM5lGGVV2A8xfg+GS+RLudniGr1fSapgOUar7hL05l1P1tiSD28rHvt1zzk5KPqWR7YPxtIqk5C
JRTqHaKIlSzw3ZDNBo2b/zdLFbT4qOBeluoh/NvvJ+y6AaBLydCh8ZJez/B0riachs6//4N/gLYw
L6BlafQmj8e4gVJo7AVFV53Jqt/Cd7mdiC1oMvstxc4O7DvI7ekELGt3DgkiFSxNFSpQLoTcr1/q
nYek1kKsshp1CHSc5AXBMpC27/LBOvouI43CXh4K2D3BhQdKgVF7ieYh/WaplBX1ic5Ty2pB4gE4
6TOVRdExJRIbnnQkIM2ijR9nsd3Kx/s/oyqQpn2cncYr7quAxIG6qpO1eBMuWzYyyK4leQfQiukU
DKU0uXRpYhkiWNFPHYUBbInoANeq3mfuFgOSf0dE7q7wWlOC3enGlsNwFpRB3XEFpnJMBnzDI8Qk
G/o6LG5cDv7oxPea857cYBwAjRkGFc01q8nuLLx3BfTpnEBqn04VJTKvzB4rzBTQERpXQ86oMHrm
UQxSwTpfmlpYLx3HVbPOC44g0lk5RcAAlO97hMCpV8mMuYMegE7DdpScKIzvvZVa0Nj92FA2FhVT
6ayPBruDnkPG3pZu/A8FDVP525gZipiq7bxOdch5UcBtfu48K1IV8uCr7rjyE36Q8swIBTnAk6fH
bSdNM+MIy/xbN+OIyZ/ApcO8WpC7rLjRhjQuKJSWAum4xZJ+upWtyeXYshuo/20khlOEuXFmRCgV
sFGjsLSwNeWJWWe2qiOQkcmSCTCjthFwwYdPAA6gyRWEUhkEB9g0iYm8wca8aL3u30yqoc1eCwi5
ybyWycX7Di6T6kWAmzMBXTPPNhzjJRN62s1/OTkZMuFZS348fK15Q1owUitfLTHO92yVmGwUe4uS
76RCRWe/WxeBHyVct9LqqAHwyzn+CPPNeShG2JkGLWaOK4s3m1NTjbRIKwYjRvkkhT5J8APk7wYk
XPy3yrJsf0TwHH7k6keLNSgLvyEmVxPgelQ8AHduSLr5P2OrNTMmZYI3T2ZAagusBnyt4DP55aNm
8iBQX1k5RL+OwB/DyNwhVnzfMX55pTr5tDeDbMVMo41H1UdPqo28hZk3ONPBFGmFnzIKT3VjbXFl
0lkhO3EJSzSN0BNmfrDwX5mH228kaWWrqua88Ol6jNrZz8K0lkZMX7VdL8tmygTSiEDBlc4GHQZ4
fujrvcQrC5bzpBURDbdh2Q2mcb0i7EiTiNdKyh5+bADRo+4a7wU6zJYiNiKGdaoDwzXx0Zw9JlL5
vber94yGqSUxWKQTD4NMa1qaShZlED93CrubNreGLxbf7WolLI8H1zKs714oNoNZZaoio7d8W5/d
/Vd/4YyJKNosqRlNYsiTGIOitVjr0DV+4P51qHWTfRGY7sDImBL92KuMw+PoExn8ZKH8+L3ZGV8m
zrpTIoRU81PztetHIfD3ToArRgbswi+hyuHsClk4pzmW21FVe17BhlrE+xKzTiYn7rZf0qi8u1bW
hwsc5Okzb6hBbXJ7bYlxJvj/MVce/xgDRnRip7zTU85jDR3Y2lnkT78HqlAAr6qWAVA7BqUryQDi
tabodJ5KwqHcZERSR+OqYjXPWj8b5dbic4fUcth49kOimhMdQ3MVM1X/xXQIjI8pPe7Kh/DO0CMP
zDhoVFNfhof/lJ7BbMsUrP+97WCM6y6KU+yDc6u7L1vUy70x4x/FP0QCBLLrT6D4k+lW+hX9ydco
/nsOomdVfFrZ9nqmu22JAZU1WVCH0cWlhqo9RvdQEb5Nqw33x9bD3guILFP4ypT4VPDBkM8Z/E1i
qXySydAs93XPvTzL/GdnX68Fn3/FExeeQnVkuscdigL1kHN5Tm+UlKQ5YmWp8GexaWGQmFxHPXsg
xsLwrMjQvqA5Z1tlubQ/fl5T6waOjuh+7Q46FzwVap2hIVqIlWBfpCrMBZoRAsqIu+IpVDZd4pq1
GpO1ScN4sEP6t57kEVMHZgDkmIJMy++kYmKedUQ0XiW0NgNwWtwDGNjasyYYIUzHN2kIekUuvFwQ
1jbPLadfN7eqe3hZ+XkcHmwtzVrDzd0zUbQa4lL2gAm8YQl5dKCqGlumbstaEH1tFWCN3entr+Z9
V/QjbwQj3eGVmx7z0V9pl9Tr2/tAh81ewUGhTN/yA7EnboHRhEvKcnRctSLn+xEehKQg9z2nEjBm
yueBnzWvtDczKX8k2k6FqlKtsKZZeovY6w8GXzYP1NkVPPumth1/9+30aBgiPXIUfszaMgI/59/d
/ALAxS7fdn11xfOWMSZQq9Gc1M/2mIdYXYLOVMoJzpxTckpFYidKasnR1o4yKJ4vH/JDXj55gCPQ
8m6txtlMf/5MJQ7pxAdKDdDHZZl6P9WQI3HPTqxwk/8qEuuEyt26zy9BNKgr2XtsvxMPKDAgHKiz
hTp15woCXwTdZ7Q7Lgig2Vq+bceyXqbZ5mQJn5XWNhMu2MU/h9Er7OlqJ6kADztjuaH1ny6YcXIu
ChchlRgkxhsMJsr9+EVaAsWpF5D6vmw7n3b5fptXQwopT6902XIOPQ+oAEbnKLbCnqKB7LcKZ9GY
XbHPCOyO9NmqaCgOnLPS/wknDrhkS1LcY/GegQoOfHct7cTE6hxWWOqBwlRoaiLrbKM3kWcpET80
GXTNCXUf5bJu11v0Jb0YayWlDlENJ5krck18UQIgJjD2cGY8kGElIS0mB5yCBDvVEwgupT7P7X8f
3KCI/bjzQToW9vwJZhLyVEZ0fU6ir3vvg6Z9LZ03c/qDwyvFCgMA5R7Y0yI9Cl7P/WshhI2jP/dY
v4J4/7adEV+4ktIl2uZBOLhppF8waun4mauoPPajv014tLgtujq7cUxfqt8Hrn0Noy4jztoqremQ
v3xN/YwsBCUwFvJw/3bYypnR3GaSNBywxwhAfU/sHReZNGrnlkucuEIDE6ge6LPqYQIoJbXzwyCv
j6VhnnB0auEyQjTHkRgThNrcg0daeVbs3XRaG97bruO8om/0Ty/qX6KfDS/dr36SRzWsQSoPdKeW
rXue2RW1L1CfuRdgBctnA2ZFvE2suGzXmRP2Oj8XWP8XtTRzHfTDCR4l9PqacOImLXpiIDUdeyVR
6rC5SaQqNiHM1CyQUND4ZCuTpQyYIhCMLGJqRYC/gbL7az/d0zRfwnUlevGiQcuO0eXu3wp8EmKB
76Ayp+jiNa3rw/K+HXceqHQruXu/vkxJOb+/yvh/6wb9C5V3UeNXMaaxZNh7tc2mjSuNwxjuF9bu
v60VOwQZ04jHfxJQoGdzluTm0GN3nH3b/Hw1E98cEuKNy4g6ApC38tiDzlvtNvEn+BP0rgrJWv3S
PCo2eU3iSnEpo7qjAQeM0p8b7YoVjklGdwOa2fff7gm5vKt9IOCqCIo9B2NcKzzqzKegWpEc2qeh
sm0qEzz/ZiY2x0FCZplp/tNdh4ui4r7ZmFxuGY1pjt26r+kQV/z5UgVwrSVROiw8JyKwP86xkpta
sDrJnAY9FSXF4YYUxMrK2DfEhGqI4GOpo6AAcWyMmSWiBp2JQjj7UamEm179BbrGahph1IhrNruu
NfVaHcglAFSyuY1TdcKM0Tl8ZVso0DtOknZjPf0ovvNagORnG1n1vQBwv84wwGQpN5ykoFXQK4yX
VAj5RRsSPOWX6wQtgzXaJiNORvdwiwkZMb8kcsBaKgoyyco3IACbeAmBKqZFjGxYHmGX8oq+uRE9
Q/amGJHL4HeGcQ7R9BefQnFh/vOFsnNoF3d1Op5dhF96yh0PwbidWkI3VsZWJepPl5pahzp01nnw
HtF09v0xw7I2NeRTsbDZ09rhAmt1ckbR7sVQAkVyja5Vkox1VpC6xboglqDIKiURYPqOTc3sFcrC
yfm7012KTdp1Lxv9UTdBt5gyqNdfyWM8lrMPLsV/qx9cWC+aiUxQfQzR3HK/IXKWPKmpvhnc3y1k
MWFeDCEmYE90yjQNLTvtat6Bn9rJfs8zGv6Q6d1nr8hGqyDPoIH++dhtjzJlTOQv+5IOzhKJH1Sx
HIkg8IcHomep0BpmEInzQ7U7z714aIoE7nK8Uyqvxlxfh4a+6GM2NDu8C6KkZZgqoTX5Hokkdm3k
vqCyKsoZxqY+z3BjTfk3vbckfwpFJw4N5kbEVTZyqB4jVtDJnQT3LVjFDMYifRTe1OfgAY7WHk9m
1TqHtStfKrKN8LZ2ctsIjlltn3eUxkdES19FkaJArZqaoRHZZucBigUuPF8BgSGTk1eM2Le3w4rN
cdmE+sVHRvWMFlRqTYOPYXdZ9GpT3PzU1Bjj0lvYvGuTsYIntJLTF2ZOkJzf26sn/ytYX68tYWQI
/spDggisxgCDgGBwtGYa9LjlesNREttR6dLY04Xzq5geBIq/oM8XcM/VZuBaQaw2OcN4kC4YF7YE
fYehcZNXsG6SJecCDoNdpqKfcepOCkirWwytCfttgfAPwa4scytAtp59DfeozMyr4J7aL8w+oNUx
FdTr7lxttFkCAs+0AGbUEzkAPi0Kze8HARk4pxyvQNs8PF+bLAmihN8OVKv2sd6eKrN7B1goRQCc
5baQ8nrZwsqPMdiwz6kuv0BuWsdeBDUaIGDy1SQKcEpe/dZkrGlAJ6Rg0pKJYit3uRxsc1Zi7qXS
UbEVWMwDy51OxNeeI9/DZUVJG2uAIhcFhdZeqsEx5Dxjr8CjzyIQ5T+ZEwp9V6/+da5GX+aoXalr
wrUZN5VEGL1t02hscOdkImJF7RbBXdyZ5EPxPKVNeODUMxHZJweQxYLqZAX3w/N0pzVbBdAyU0BT
ZuKR0S99xDNiVXJeqCLWv/9SzKFJ9kabCERArkQUyrSGnV7XFXpHu7HPZN+Ph+qhdq2j+lFfASon
ui+wwEi9tn/GsbAu8qnNQZ0dzTQ3OefFQJQennH3b/Wap5Lo20UAbJZEfnv8/2LdisLJP2jaSOyf
ZN15JX/7O0crteA1bYkOtkRKWO6SLM4SWRISYE4FBh2Dmep++lPL5arIjCLg8Umsm9wb2oNbWsGb
S2UEG0O5kIiXrXV4Kp2iSRRBaUPgvS2MmyB+XDxnHbOp1rsOxis5wkNgf9NzLljysDFzz7KEwPbC
tKHDwDMIGXewDR5S7DI2TLxO+WWBpqEag66Qv+Zg4kBnFT0X91UxQaAEXznfEilZhdT4JQ+CMxhB
9ismO8QkeI5FDym7vCL9KvtrItpnNqLCuttqtDHVkaHYrtue8AhVGZIRzeVRPw9VKM7LUNYdcXzw
qlJUInZVXX6Gq812lHlybWPdOIt9N+Bh17SK0CrN2gI3t7qS1lHUNeV3QytY7XE5uhbTLOTxDVuT
vh6i7FxQRfD81TN+Rf/jA66iX4QyXbBoZVpAMmRu1mbqkqOfI1o1stAcOxSMeRb5iSuDfaeG+Dp6
RNAsvzi7svxa21fqlNMw4sY8P8oabeVtJN0Pp+7Xrs0egg2cQ5aFPShR10TI8p8yUBp+xP1RXgtF
4vLc8aQUMW9VQkZVg22B9dqlJJmSj97NEeqUPqPWMdfiIr0VPxV1cWpzzIq5e/CCfE7jC3medzJs
usSjSO0T18w06oW9qT3aYC5lC1amN5G0uyCa4q/cm2JQY4PET+ADZP4KfwHeMAaTE9qDDQlbl2+i
VRPLKNvHFRRUgTNZm7F+1FuOESEPNrLiAaPJq87itTl2B5aBKVZJWoc1LZMnelHxhCIVZ2rwoS6L
QbxJTn7ej9dE+2L3DB3VYqwbAjL+I8jzKX+wMgOjpDuLGRCByW2JmPSwsng//ZRTjXQ4noJ+wnm4
Sw0I0W5dKYbOwm6OlR7CW60fWsIkO3uS2ZNJMs2HPEnUM3amnhQ2BPannRUisl7KNs1ocyyezL7k
87HwxEpm73GtVqmS3HcODr4p80YEVCix75lOY3lZ5JpEJvou6nqAeasTLCxLkPXZIXKBFUPi7R9m
HfMs8VLdnB0HNSCwMpX3QoQ8clcMOPvU2x2Pt82LGclXYU4QIj3ai+xskc0ktPH4zFwl0EDhlSd8
ku0KNk8k3AUinFcURjQv19l4TDoHCWql3LtghkzjTYWwWJSaVKY44mPsDnpiApZxDvPTdGt6SoMq
tj7AR5B+HFAauRd0+jfFlni8AqurMTXva1KQNA6uId8bnhLAPV0+OP+H4LGSGAU6sJum8NKpffmZ
2zzT2yEnb8fFxIkPUlryjYujLpvyQNmKEFUxGPzcv+jOZXSFqje5dzesuvODenTOvAFw6Ydhyr+F
+oCGcHd9/RlPdHOX/QaXSG+4GXpAzkiCVAvMdRDET81PFerfwB7x7SkfncgDSwyJI6IJi/ZPImYR
IelmwXgztmuIrHMsnomL7RlIBEtAgpAvbKs1xyvoTNmsA87Bfngxz2gEyvVndKuPlOGKuOn9ok9l
J/sEttL6M2ZDCrhQHTxbS4cTSVIJuQdLRhjFfmzSSYppFQN0KJWovTc51VHQYEvHltZLyYiTF2f0
4qqVqm9K9Ch1D6Q7kNtk34gTkGEPLNyfE673MLl0Ifm3/F5S7wEfYcxZlW15tnHF4L1exWg6Rze0
IQK7B+pD9ut9xJSx8SbpyILWv+G7B9aI0s3iDHDtx/J1aJa5PZuu2+wocVtnB/LENQtWgdopYW4j
yYP+BBDxnBouOXCB+fQeDT5RVSS+eUH7jeEgIiF1AbgWvHSs5M0hiFdQGDrgTJkf2JyYrm67AEvn
r7m2o4DwM/5xGd6F1q+dSteWeXR6q0WHHhOKNFFATbkd/cu/X+8gkaZvjTuo6Vy3MVNJeNTItLPA
8HjRe+Y6UTfQn1OQxi8UigLQ/sDv67EPxvRVjaH9onIg4T8hHhzl20VgztdSwzonzbS8uozgyOsn
UmL0t4QYW8OaFRpVJOEgddzNeuFXRplBp5aEajUJanvoJ30113y5cvj8429M71lIrKfk9EVXfsi3
emWszg/TfGKIV0VwUJHAtJeT9zEHNK83zDLq4/m+XmneXwsTvfY0TQfsvNQsvcDvz4OnHb3ILHex
6T9CFIJvW36hMfUTcPuz7+VnL3Degrghw/qhimmkJT2xoICLAHwfVxey/ojNhUhomqyfFMfyI4Xm
TxsGG5MlyYINlRq3yZSaGhzAXfsvZwVAIQJ2Dc2G94UYc+Q4Lq8/CJ7Ein2CXsNxaWM2X9k8gUeU
KA1wl96ods+PqM2OHZdjWLYhY1PF5Mi8sGPJQAgpiyubOqE+hIp2k4Ilya6SYxdI58mYn5hEwl2U
etivpGcbEYXG0pIS1YwulZmJyyZHGhSdispronro+2dpG8jCooZcJDcN0KVNbLTBnESR/hmM1k05
b2IQ8WDBeC0XmAuCCg6gTOO7Im5ulznF4tdNvEBYXjKrzaIXUTbqqxV8tXSUGi8/cdz2qbcyTKDK
n0lkrj4GklazKxIj1D7XvYeTG8eB0rKorcLyMmMeXyIhbveSwwRa7oyMRPSaziKKfgP2a+dH3plg
eSWtE8/MP+6MHZnaLjepoEmodAR+aEVSlNpFyHyMo+bWxtfKwJi4VKY1EF1UR/nFvZkYeG90+wmL
52QIaqTiJ44ETKEd8y0lS3Jro995/O8K5cZsCf34ou20fs6P6DUWwMplGtS/xeS4OoOAfdv6M4Di
fz5FCw4ATUm8NR4SKU4PQc+iES3dNmMTkVB5J2qDd6jqxm6hgy+YT3URduX0Kn7LvcBYBBFHQ7td
DnolEWixvH5fHxKxGgtdHZetoAFAJ4ZSHI6De3WcQiHayUKVQPn0DxyHZRRKr6DQZ1dhDPH7/D6O
CkIz5qMNesWe+z1JtuEAGcfHKE/SUOUUHyNZv34W4gMpzK/9L2mJQDpOem0K+qDZsAOaVkoNwxEB
lOOW/lt8OhPwojpDMZaTfniuqpoE+FJs+f6EuVXQp/ZZwwUSyxlXCB386+tdjTAh7aCkCVum3h5P
yTrTh4SwR3QtiMuQ2He1vtePaNs37O25+mlV3HURDWRq32kIdI1Vr4TTltXGwXoDWTw+64IEF+cA
biiYnCKq37cLIeKWCsq1Jb4fB4YKfhdg1gcBraLpfRP04hUf3/pNEelFn4o2TJlYVFBEnxEqxIFD
g++ZadRHmAFDkIDBAyeHLiGs/G2gYpCBY6XOPPG9dVJO2gDCZ9EuPs5FGF5MDG4CtzJpYD7oIDNR
8hMCKsQ23TT+AK9xsEAxhe7YKHwZCVmEXIze4FHuzH2XTaFm6dlTvtSRYd4H8N9jCve4jntazsuq
41F72+o1HZhRssizfPw4lX7PNcdvtcIpwf9JtNGiG3V5YBZj+lCYf5kB3yIZrHb0dcG+ImyTwHVK
FMU5DO9JLCv2nQ7dhzE7pNOhI8+7d0eo6o0uocPbLa+Lel8O+RlLrj31g6YwDq+AgiAC26VYyndz
Aw+m3QlE8IxrgOJXRvtqLGhxgeqZFq7vGsELH+y9wHzq1eOtjSVjBZtYPqCF/Hr9U0yl3JydPQYQ
C+IFv9b+AucN6++IzhXsdVCuuqHa0V2OJLHJtha2cZ8eYZoMiQ3Zyu3LWwlhxsSGdTCaAV6Qf60r
CS5Srpb9rMmPWOhcwwTtBmWN+/SELCS0ImX1rgJ4fMVEa1qTjTcslElGWwr6lvWeoLKqCW+39+q9
6tZVyJUp3bG44fN4/v8gquEgS+Qp+PfsfSsQeLM0vo6dIeaP7lNvwA1PLQQntgUxFM6GiCLHGpGM
1DrFH54cjc1Xd6CIG1sNl44s267/HIovh0TbJZK3Fh6VEKurOyUDF/clPAPwxiy96boLlTgcG+6L
kf1XTf6R6Rrwgn0HQXo0dqg8JLxdcwNqapFriLaOUuB9I4uQZtyI+RKAXj9NDpKRWUHW++BRp+0X
Gd900xxo1d3CG3/6bieVPdEwXbkTNuitEecR/NrrJ6GBP1BitUU78KyyG9elZ4udWAs7T9WKE8aY
UU9pS1WGFLNLrmEo22wAVOl7M095+hiasHABFsSxxqS7paKSEzyr/dL2sSqtNbJsPQ2JjgcNkLuY
csKnooeLmmqhb6KazEHV5kg4JPtDU9y0X47kJhQO2pvZo5ItXq48S27FzBpzdbXLJSZbVJ+smpfs
buzN1sc7Q/i9HaJlSTpz+PTCkk3SHm9aSz1NlGZNjToPRL9iGJtTliCNOnxrvs548yJL6KBqldAF
3LiK1sJl4RwEQ+vrcC+gH9hN3783hfHpNikI9K34UlnN9HBUm/0a+VUcPHo2umrHLButrYICToAg
rYFI9tuWmjxEQkq6D3al60tOgxRRynLrqTa81Up10VmYw0Mqeeqdd2JCtv654Xh4oEpbuyWaRUov
n0kGlZsE6HIy34FaAMTnnA1gq7uEgyESeWLlBCmmihgVfcAJ/Ayk9ZFdopYPmcPcmnJXr+Y0WjU/
DuFBbXlTfo83cz4qsF5016c+nqOJcaSYrw0p6EDOv3h2m3WbKVHUfVvVu9R8yC7aGerM6LcOIIs5
SkJFGXuumnQmytMtPT+zNrn5v42cV4K4677d11ADLdFDeS9d4us6ytn63yBCQw5b/cKlfXuIOsrd
wjqYTl0bwFKczTyKjkNCcEHICbIWj+NkBclji8epX81ZpvPm2EQrXM/v3/F59ZNDwNTdOKlYT2Qc
GUBAC2HHmddGC2wz+iDJYxWmzOdqIQ5En3IdHK8xAkMLx0UDO1KMHLRnLfi2RnOGm3a6aZJFQp/b
kHER8qjnzYlKahqrKNDtbzpnz9257N+hT7o3vGDudNzX8gBAVjn1aXlCdkWRQQI/9WBftES/P07l
305aH9ZJtqZy37MnhFDb7xMBgBDOUVXXQut9tPE7TKeP/vsIyyy5t6PumqDpUzBh8ToH05YrupnX
ruY5ULd80qmJVORr99IDu9Hk6U5gGaFIMNJVqGzt+spOnyMsIhGX7Img5u7PYjy25AoyKWf2+e6c
iQqUlU6vO4ps6vliIYnZEPdDrNAfQdfUzIQ1LPI55pOxFju7nPykA6lll7o6zhA+XOPz6N/tKEUK
tME2/T8fPxzibuypJs8umVv0KkgUNRh/IBmOt5uqqPyJZCri00JnKi/SHgifRAAZtCWoNlnY6Dar
9Jr0EkSs7kkKSEOgqD90iObEOJyY40tyXq3LWL+miekDG8kRSQHCh/ihVM8/H+kThuRycBJe6Z9E
ugu6FW/kdD7Y+dFmlvHz5r6GB2S6NxjDKfcu+OrmNLHahyEy0tMY6YVUieqZIXf7jB4Ki5QKX/uc
6/OiT9+qx7QAjg3rt+VpeNWGjw3mxpcijLLc4PxYwKgJibn49aGuSiDdTfOi7JkgmckVaU9JFJGy
uTvwQ7OfxMhLSTEHyhD2Wv/+CvHKmJ+KvUcP+1yJUci3jJR0nziGwwqziWCipfE2tIsZbUafiw6+
517Ub4VhrDiCjIejxXsUWIiR8puPuNeA1DgSkNKUZqXt3m5q7/l0cpG7wqt8flQqlYAJCwYNt2IZ
aIVhjhhl65IjQ4SJ/ToMwqAaIUeAaYKsit6xU2nItVnvJby8nG+ThT/7W6F3jHkQk/Awr3H1i782
mV9rDIl4Grk2dOUIiWqWLqu79O2+LeseVLn+c1CvGEURoWHFT0DXWzA0fVSmzQ6nPnxmq680wg9g
u+fbm+4TEcRHu4hvMEAJqHxpN+L5yb6VOVld6RORC0wBFIybta2410R9r+prERZVNmGEPXASEtOd
DG8OKRex2Ki+mdIz5iI7+ZHzO+vKsNdeYk8AiSKmuAGG4I+h8olxJf7gcOHw7RzXAbP+xy4Wci6Y
xTpQ5d5kKBToG+m0rtl3vGmQs7nZCEov+mb1N0csX2CAsvR7S7+xQeBm56p2IVG8npygnmxW466d
OLd3RQ+yfJwoqiWSmCuh3O488+KwNa5qxQIEaMFAuOGdlVfw/Ao1Jjp32XXMNmVtwvFGBHF0w4Uh
jb1+7W2hKxjtPKzmRMM/gKHUnUW9Ik3p8aKaEpeQ5Z8LiNcTiTISv78aAhyQ1/L6ZHKBAjfb0zSq
TGpixsfVziNsJ+q+D8MfWextIEnV6YPdOXKk0tqj1lU5SnqRChBgcL3O80o/3Mix1a8bikUS8Yn+
43NrgFiSGngpm/4vgdH0lJHjAPm4Hbd3hTye9agzp7mf2b6H6WrzQ4ZbhyYnDrzAJMaZ2mqI4ZS/
/dcYTtlykHNj9Rb9Aw9V9eD5Y3k5R4djOi0W4Ul/P9hy1HTfYbhq7kknZfwrm53aWbOqS6iiJIIf
dMrRa8c5eOLWIuEzc/lKECH3Hq0e7CkQ0OZHKqziGMSbF/HPi1eh663YQaWCujKUhm4LBcv6df4m
x7iMEHSgoBap0S8rms40jAPEtE+GhbPeqgyZLLgidKuPS/u2byz3wP+Vul5YOhimQRKqi+Exe/f4
zhG/OE66St6C0zW050ylGtX28WoDdouISSaxJooh9txrsBCz9DFhaqGBOnLlbs0lmiFW+1Qemjom
moxM1wCOUn7lmEinUCYwfhjA7Bas8mRqRvsuVhVHh6L1XkvPwFs/LFurI8d+ObnWkSMwdJGJKGSI
7MwYai9K1UNvjjQJirq4jRczBnSgafTwlxOt09j1acJ8Wx83vGLJdB56pn6sixTWyMUS55203hBX
RJcVtC0VCdIpuj+1Vhoi/UN20Oa6KtFZJ3WQAWhBDcFCzMpqxSbkAo1EHM5HKEwRCzh6UACEKaEF
QUsFEvevbvq19A0UD+X4vapOXnt6SgF9j+HFu7HNZ10DVi917FlwEi20IpzkQKIAz0vQrEqEvfz/
Vn5eIyZb1xIsWVH7nAb2iU1T1d2dY0q+tei4VGZ+zfO4TgelmL/4LS9hO5G+qELyr7AUMcovmxWa
f1U9LnhUUH71uLWrBQFOvmJ2I0v7dNE8/8Wxfks7KdpkZGbb3pRPgbv5/yxudHPkDlCuop7H5wk+
hw9qeU2rsPVonz+m1wNNiXwshzR3wXxtTRYWxzoMKKXYqdbuDY7WRRoL04J8F1uhgQSw2r6lcHtE
kkrP63A0UG823ZTDABXi6BkEmZTkg/pWbJ0lvKxGSmtyK81CbVnRcDkBpQ413YWe3YpdAnziLrr+
WnDydGq6buoavk0f3koq7aP5j8W0NfXwQlHw8FKAFGYqBFduUeByLGf9P3Ury2uzNQsyitMj4uSh
BUJkQF8wQrpZaDaf0EOOdGvrTHG1q+O3KI7XjuqSc/VKMRf87qjp0+c0WwjgJTENVUNXmYYwoqkk
KVepJLOOQpBpWDdux7FG55wsx4WyqjCvgafrz9TVgMcw907bDzD8cG0IBX284455qQCSAAamJVSW
hSWXjOC8X4tZi2jBZ5qTrARU/eVD2+irnMmPeWTxWZGiOfG8cefN8D5NFemi6tXpaRwB1V29Sn/s
xosJlBOvkyzjfsv7hzVes0YxQZ5rUrKNexFrUq9/eObaTQVoOS2uaY1G7gycWb2xeeVVDxGXQELl
k6Hpc46SyDFPgumfc403BYDKU1IUiHq7d+8erqPbFLeZivo2JIL1H8sP61QaX+n8ZFxpvXYkYLDS
8Lm1/u1v2ZkmxuAkvlNhU7rt50TN/XGf5Ea1mxNbwU3qsRIUiJB7N9bJJpbPl1rlZLmhdBDs+jr3
WBBJLznTZ+MgEqDTVKOS+3IhQmg67HQ01vr4sv8es/SM/rPYPtkEkC5C7bUtLhyUvyhJNaBkXtEn
GdSenbquinQzKX7ziE+cNmticvZ4q9efay/ufbioQVi/pX1sZR8JPhzJJ3rhNl1HxrILRgFRWgRs
byGpsgdzy2MEIx6YiedqbffMaefQp2lYrhNYSfjN34qrcxPadM419AVJAEQ2KypoDVEqVPookxNJ
evLZXSsMDhzCUOfJCT7GngBO6kqoIjRUoS0t5rpnMsFJkbErTn/vIzZoz3E+ayPYkgyG5TdO0j48
98NUaQNDwWBgfRm+RYa9QnFGCmI9L36CNYT5JmSqLVJGxVORUxQkzZSQQ6Yt2BS8LBMWrqCebiSA
17DMaqRvKqFnRirv4N9zcvpWMnlynlsMl/RZhMG3ue6WtOdxLxmv5kJpnrKL1gBRSvXz6JAlDiYT
WifLmiMX+maQVNaARdlheZz1Ha+7/uuO2uNoVWYQYYdXIwOltABefemRqPF7You1VQUY7eHxxO6n
oHQeZ/2G0IxRSB057NCVpaIPmR9qZnI6U4Oh4VuqcNTdND7jEWt/2P1c5dkQB/hw/rLRN2IfuXNX
mFvyoX9FVzw4oqPKRbJn0NG3HMzHmpBvznCJnbZGJwnjqTcUTWOX7eIa9bJd7t0sJhu+1SPTeVgZ
vrXVpR+JzTrANfxJK2q9CADymSPvZsTufLukvYO//HDaOW7REPtRJBKw0jtsF3Hs2HLh0C+Uga96
KNB2Mx9MfmwJIbEVdh20Ido9Eb9XzgdZiTho4xMqsDzCSE2HbrZ3v7HXwbCx/QT/AQTzeYNybov5
Jp5cv3tmd2e8e3KXpPIhlWqOmZUU2F/ZtgsZ0oN67AXc5ZX9h+EjvVslZnbNtwPncbwvrjNpx7Tz
QyxCTyNUoUpcmhkVSMVfZ8jd5Q3O2kaGZMnfbQZ+09Qk3fiJ1S+cWKtMQTcD6O8tKXkIZMyDYSOG
YJASJNOVe+uMfp+1wEKjKU+H8vNUNgV8+Sdga9K2Pet1BBDNxEyP5hus4yMdqDcwsj1P917iyIGU
K6LhLlSwAZCJTQwYPJGkYLRvYL1vmX3KaGtN0lfxzWaeZhVRwGMydyl5/lqTe6sYsvpHaLuTnWaw
KYA4XKCrSkH8XCEMEGFGaRFU0Bc3D7oYWLoFIB9DvijtuESsac2lcehRHUNK0taiDCWcM7bMTrdi
XOnAqcRmv7UgseoERQQTuLPDpvmrAC6KtzSFxhpRlvKCFRvpv4E/fe+8L275AJIotyTAWCzw2tTd
dU86fO6mzzR4H8WBoeJkPeCJvbehYmZ+lpaI4Py3PxTADw8Q3v1PmuvAiaBeBACj1yCodvA1jObn
3zi1JAZXM0BEyVH8dn5hmQWRDC6pwO5fxWJPEp2f+yepBm+gj4noyIqgY5uIx81eeYa+ctp6jxzV
IGByZSeKs8kDjZL48DxSLrEcyEeaaoivkkz6fLAKt49m8eEPRq47tWhs5O0e0WG9dFYMHzXCFrsE
qKqfYbHrv/t/QmACkylql6AGJ146UgowbjeSAnc1v5Jbgz4eKeyK6MdslkAa7UiPLEKAotP7n6cN
+zekKOunK6cZP7yQevFACpZqg7c5tguotZwCoIQqq9jTACJo77Lv28/kwAX/QlXFZZSPLwwHw326
HN4jQ09x9dMITEw2yPtUHZoTFmqyym5X3F+2slpgktFx/flJHIcwfW3Yq4dOmo9Ue/o8uhZr+zzx
7rvWdC+l9eTHecsS9o+ffnbOj+094vBnSh9VgBXw+vI3g4qG2tcxhD+ScWFigOqsIDyR1DCfKkIs
G+QA5322FN7k17TZN0RXIbKdnON75U03UIeu1C5a5oXc/UbXa+/cyLqvNHwpQ7xXhDTEmg70fw22
GL2wYHfATU2W/3dp+n7rmXldZllDuF+Q3hrmLtJFGy/Lq/jvIBYip1sIK1mSdNV1V6cwhRHWC8wT
jEhE65BtpXTg5vNNLC2YmhIqx31P4PDf6WeDlv4x7F8/VN+rqqk2KvQftR+30vdC/XlGnnVougGI
Aei73tSQ3K4fo6nQSEmSkEaMhald5bA358fEraLELjkPupSVSWnYIOghZKTcizRORS6fXgoLEEqx
ZDo7RWyvgwHxaezpS1wHeeDgduurXGHV6zf0yERxJx17ins6Mra2aw27pne6YbsrcoBRBwYLfcEk
vaLgBES6Pj+Vm3xY8PxrBtWR8/iXteOApT/kOpBoNhTVV8y+qGvVsrkgcx9QyiqYMQi6yNpRb2o6
baLQisg4lykxao2rxtn4TqhRiCBx6Vp1SLAdWODgTPas4auQjC6WZlb6rAkELM+fCg6oAr+gBuoI
8Zt+pnq6AcJa+PgxlxdEha2SqwAvtW/HOf8gSxjbeoT3AF2ENi286ZmUW2Xe/K2c2N8edVLcJwzD
sezpObJ1uAKL9a2vqJ1+n6Nhh047PJdjpRjAzl/rq+QMMB+sMBAhSIHNMLjyofQJbWIHc4ELeWsB
w7n+itfEtV0OUU0zrJwqT4iG9MpLkb1lCCZNfswh6IJ4srq5Hz9gEhkDGBE6yDFCZWr4/o55kUrb
v+UCeCC9jPb19JhNjeuVN2GkabtKei/2nWHGCi5ZroR6WKlr955ec8Jk075kWFMMQuNL9cndy+En
JRouFmxuudiZDQUPVk9U40EU9boMMaHwq6Dg6I2bEvJQODVc4zciqy3oIed0x+SAj21XwvBWcri+
5d50eL3BW705DcyLfNHP9nnsG11NK7rVeVsgiACBLRy/oHouWZdul5utUfcHArSPdgM8MVgzUqqj
fLYmPW76Poj7xafKvC6ALhvHAT26n5LVYTCLs42CP6J0Om+SnWvJ1T1VSI09A1FA2pTATtNEa+PC
iG0EEnpkbp3xTu9UxZYcFrlLCowpMNFJJXNiPjD5aZ+TuwXjrjUbgCO/xQ7jnnXe9BnqdOY8u0BM
6EAAgJqzOES8yQUrjEob0PdBlV/jWdRASaOX4einUYGVvEDMWhUg3SKoWk/niuDI9EeGcfM6/z5X
hMm2Xk8kCU/l9R1keNZmM1cekM2c0oWPzQec0nl99MSdRBH5j2BpXt6450B/pRSfzY9V0Y92HNp5
Ao8OVwI0zW2EA1BfQvfrHly7klGYipAfiw2LRJBt6oHxR7xOSXGfBVZ4KT3OHdom9BHwG6qoIH37
j45A7MMPxk8H3wZzjMPn0GRZv31uE6tsvz17/1pbmZqkStXi99WloC0BUi6neEyegRg631IzPsIx
aikqT6QdvQrd02qPLhEz9GnP6rKkOOlYvl4+bPE6j+a10IW1TpZKDaaoJA2hTw+HxXqvS12dwO+1
zjMYUMeu3b/JhflcRoQQu9sJYq2K63usE0mFWs2yvCgAUlWM1RajA6KekqZ6DNOp89+/3AcK5W/+
vP6LYbFYIpO/kOodMSI6Uo9HlEuRqN638/RygsRXzAxOGTTZiQZfcRyuxNHlTtfRcyekNcUS6UVE
JV1muXydII+WsKbmV5yUzhDO/trm8OkLIBP+sLQGMq/uYMSm5aHZRme7yBiy/BZW/YZlyGand9pC
8ZPxgX9dqGpBZDQfL/rkERBndIENrSLVdSW1EQMHLiB+KRxjye+3k75fziVUgQwHNaeV6xsoqd0Z
ic2Ttx/77BKG15OZ7qYNqbrgrcYRLR8vFoM8rwA++ZuGU1eTyh2TmfiphUWyoi4dfTw6eP4aiCqa
jzRM3hHJW0ucfhOd9Enk3tbofVQ3xUZAimWn5z5AZ3c3wsS2xNqYIcVr/2wUpkCorPJ7YX9XSiwv
ny6FToG40/hkVUpnvS4NFNqmQEFK+1KnpeQy/gLVELBAxHJDOUXknIrvsEEjfeATl4DB4aDAIApQ
rSGg/DGtKC9/Zv4y7LlO9nvUWFdcD2WrwGm1i9S1Uay3ycO3w3YDmb6BeiJwNTQRYiAS9+zS6ZPH
o52HW3e41gDgz7KAEo6plFAIdfQXTaTxrF5IM+Rki1NtCl5/RqYqmo7x9RK/D9fg9VWRQoAZNgnM
rfQ9DZ2TPyX0rvKxWNGRUQ1gZ+BcvO0iQ2DpBDPxNnkYDBpKTIBCRN3mdi7BisZ6gX7553YA74Kr
yfTPtH9f1IjNODTGvpjVW/yGjcO3pqH1LKZyZ2VmzzdjefKQOVBfUOTCEPsVUfTZiOFDKNCvZqMa
cnQricnPDWKDK5rmjPJji0s3l1Ifv58BDQ1LBUJA34v/upAQ9PbhRnjGd2Ef41BEfsumMouYkRPr
HQl57RRaSpwp/78sZiv+P2AKtZ/tqq2Ve9mQ+i3b1CIFu/X+ZIblNGJQcpHtimPGlN9Cp14tCUSe
gKbTTFVQEsDRO5NthPhlYJuARliTujnlOkNMgR5MCMEAkRZNYPbBnneaumDvbWFDBJqipvDQvt+Y
chr4Pa8qftemMnjdxOjK1Im2Vbusb1DLtAQSILYpPdTnFtn0/Hs0IBtqbXKAlRmRCF5i3t08WAnT
NOFCpJFFlUpFjCkHgLDHs3pTLi+e70JKcFwW+JzhnzS6eUheYdtmiDCmE/SE19FfJPfl7lQ0CCwa
9+WwuXEDogPmTFWfvhJRqB2oV+PjS3mIS6g/4uwol4IUgRiMVF0eOddfbBXJyWKA3mgU3dQAyrkV
X9x41Y2XlOT4tLIF/Y5EpgFNeHDe2baSzc3sVfTWIsGtS4oPuy9LtIdwn+0XKzWv7hYrwrC1UIG1
StOGocFudgnEmdvRFULdFUhzTTXxDOH5I8EbhEUH+cd4xj0AD12nmNE4Ocu0/m1P6EnrphvFrR6M
WAocwodyEeKj+4TDhjE5cmRYOqrjCQU1ZZbj20Vl/zLYJsf/VWbAiejN758UR1aqlvcqLuDixZTE
/SM0Vsfc8y8jE1aQGzLYc+l1Q0g3ZYGI9yTd/Tsch7KQHdJEzZP6SQIpaUKenmMrS8NPH9/Ngu0x
cZN1cufCd+zSG/xK4fTDMZM4tLfpDu9ktQ6IoodsStoxQWf/918zLkCdvHbfB5NuWY7XXQ5UGtbZ
o/gjlFTqfoj35Y/zWUGOhZ/f30+2n1B33tCGMrmzAPNskpGP/roTJMppd+54fXOHyBkE43fBQ12J
YQTU7CUVc5GhtwL1glOML9fgdlkR+7T8WAHUTq2BIu8lnxIaOKADPysHl+/CLybJtPH0xa6IOrkn
bCjn8Jrs7gvzzRj+IrSEWs/mtZtdHDSpyFr8wU9Okjgx32Wm6eHDTuJFJzpmO6sSDHpj4nFRQ9tt
SK2HFTyEcM2oT9bDt1GYwdnB/4JynJc1HWKJa72acLkLf9ieqH8Ql4/iiMabZa8A7G0PZaQQEBlT
ACPn7Wclnx2xKn1KrE47WFHDA0iNsxVqjGhdf1e5079bW7j/xicpMwOsnEv2aAFBzEgvVV9FQ8qx
KbgJONm9HpOUWvICK6raGfQ+hUHfRSVV6yz2Kc2DadOOGv7aflqk6WN4SkvKWyXt0qcaYz9+kAxq
WVPv/UNRGJIFPvN6xUJxwIYh/187GlG6Hv2cavoRloUd1ud0GTa9sLORPrBXGRWmIWqOS7F27P3u
ARi3umlm+JwG83BB4tLMJV2bj+thSuI2DBAeGF26iCDZAqc974UpFdbB9khqZonCWZwxEtq6ij06
OkLdk11p/IxUjoYmODmjLbiPh5c5qRsp/E27j4cPlCTQ4tSb6mMkvCYj5l+OP7ubsPARjcsUPoZt
JlKgIP0ortZVsTF0vR0UTxTCAtsYQPB7KWg3DCKtOdFFDb5W3C2NCV0nZKByx5AlsTKdsP659jDY
F8/3tBQvnHpepeo8T+qN45r/Y2Z6sUxvhmXB5UTtE+eqQUmYBpLm2Q0ORL6yOcnDBkPKqHt0S9sx
bLihpDqkpL+mX+omuG1Qs1ugn7wr7spAq5B7TnLOHXLvbnT3ZepVKk1OpIzIGY6QhJcO9ulfBAWG
f6clWvK6kGI6WGhOhpCYYQBmKFHUvpbp9KggYiLVdJ08ZeXVSzAFTVwJ1InDV/BBcz1VNZgKC+Ra
3PDU1lKxScmOAYaIUWbZqv70UIU4pdKk2IZO/C7SqPdhV7JrXq+1oCgAxvbtRbD4JIR/Z3FEoWim
+5EcEv0hpSvmmNnkh0js6qE5GxsJZjHp+E3/M74XVNrwos3TzShpe39mKtKXHc6Pl6ZGp1a+IyDd
5Moedt2A8LT2HQxhTMvdT9dFFVnJ+WvZx/+tvM/s9/5w+6z72U1RblM1136Do/PyQLSprP3VIMSl
q0elHbClj4RBD1NzkkVb40/qXKotAi9E0bXhM4z82iuiL6u0QbElh4QtRk7X6mP9DajTVA4Wh782
gLanKzZb7jRO77dhyMrzbPLGfZCLaV3kT53BLb4Q148OPpF/0pr5leyM2+5+rdNFiY66Uarr/ZIq
a3am2yJD3cU0IGnt/I/yXaxy+WUP1MvoqZQ24hUli14ICToQVwkeQfp9BWdxjLJssngNfq7chISD
lA4WwauE8WJZ4MUTlOgftti2js4lkpdstWVOzcr1hGQYtf37i2CF8hWtwQg+5MoOL8LisIdq9w8x
F3FFsig3vMzbcGG6nrHF0A8rNHyqc3peIKivQDuO9mcPyeF0Hcf7ua8Bb3sdgdP4fqHHjIuGiwdB
8JpXX/2QCnnC7Za6C2mPY1bZdEHXK8ay5THqNbdpI5L71AD0bHgfxN5UQWlUOFiXcSW0Rac6dc0m
HOkaXh5tUeboSmkKynjWBKVc3nk9mxkHZupKcy28E4OrgzXrFU7mJAW5wRnGiGvmfWnDyyHMie+s
scZY0xQKm1kxlveqPBadJqhuopDn7qfsvBgCVjqZ+sywxJVYwGYLKl9qUdYWRPorspuTBsKVNXDb
lr9P1Ll5LpA2MQHldY6zzwQPGqx0nz1OwV1gWoG7007b/1az7uOsIpdRXeo2viuO/a0vtRUWQNl4
ov61gnhO+NzbeIN7/qYuUlrYE2O5fCZU9A6hgs0Is6JiO/yrDrTZ4VrCGq4n7Fhkg4emqmFxkBzH
PwEwRlWJQHxfwFl+CFR3oLbRtsrA95eJ70fBPOAnrxlOnPZ6d9FZB9ibZ5kQ7fpL/XLHMSf0hTtc
OKlcKOCIvZwso20hh7OtKyPls8aCdo+/21p8odmTBISr1zE4P5kSSQLGGOsoECm6KYhBAtVB6hak
JQ7gMkBWFsYx4z/gOuJ0WVGpnrCJE1qmF7EGvgxWXtjIUwfobLK9lhfID9UPcadyvU8kIYqCcIZW
21Z6aiJVFICqzj2GVYWxPxy2J3iqqietjE77azgJ/RLuGvS9fWL6aP0Z8nj8rLGTw9Yuc6rs8CdJ
aWAWPc4PfEq+k7Z0wCAYQHaxjMGoVuFizofJDTWh71sfA44P34x3e7CY1yQ4jyUAJik2uS2SWBYU
b8B2gHbbkA0Cuu0auWcs0UnZY6au9YjhsCOFkYEj2zBqz9Z8i+77kR5lFlI8ZAtLjgNRssLwjOZl
Ne6u74Pb9mwaDL/XdKPK17JSc28GrUpnoyO+psiHcZ+K7lwaJA1eT+5LZXU6JEwcH+5U2ECRBRMB
IJnflVDKFSzONwCnirKs4uh1AUOZ6+OcMQq+9tQWzKmoPusaFMbQ/JlQ1LfcWc7wyfSfjbZpQMOx
I9GLN/Z1mTOFuB5UCk4PjJxQJM7lYyaYj+xGf0hn76RBEvnBIHTEET+jrO8f0gGHYrvVr7sYguIS
hFvKWN4U3Hc+pZIKZlW/MnxAPpYk7pM8d0ExLXbezMjSifNgrlJoDBfhTEw1CfBk3DbvqZbz1EQh
kyolHF9GJ0Ei4VkKvHr6QHzuN+8dzVwJx62dRSxwe5aj1XeqUz7sekeGNw52yt6nNS0mHnCOWfdX
QghGDqd7PWFdcfPiGs/Rs5ULBy3TBXxjGrL/OZUZedJcp3uOfDqTQDG34KNjde5xKaQdUF2gTQND
JnEpfi+xXyrhT79Q1py4D5SmjEbd3bigl5ix+FqmKpRrJv20udV6Od5T5xKmhYt8XYlLx3vqB4+L
dtsab7eUTzIOt/3oK6pJkzxHQhPg3Cq19Sl0fNJ3jGdU3Tnxl/oLlRWBpw6r8Hlwv05Ti1mTQOgC
cj2TyYHNIw2LQ3yhSIPzfvCCkjd8DEYFf1NLA6IEGNuBY3XehVYbOQcS1bYGGaLANwc67HYvqvR9
533ecK09nTSxGPOYT8pQMwgdLNUCuFoI/Rsv9ScAUZswX6dG5y33ivypIKzM8+OZpbm5cbVy6xrT
pGakA8DJJGZN7v5jEnywQulRlScriS+DmUH2wuNl56s+DMKwByFiBBZs9k4yD61kEcOK+8wXVLl6
n9D2isjrUTLj6neMtkRUbSVQi3hdXecsItY5lXSA30OD7fYzV/l+rpRkfJFZNdtzPbYdyx31QtoX
1FtuR7hz9msI6ZBgYJXMaAElMp0JHfCOF8gg+uEZM4N17QSmXASC1RwFoFS3SS2nA2cN/99p4Prb
Yt3j5EmCRqRpgNvbS+igBipM9HEzW0kpD0jUlBvyR5iRDGD1ByTk8ovXCJBK9RfNwjWYUCZys2Ik
2oJzRj3hVwdTh3RXvHwsyNgYlUSI130f7XvLF1cwmhAD7tJ09Ci1YkNkA5nSRJuPVQuh8J8jU7/1
DDF6loK4Xd1f2seLLUspNob8MXfAF0Bugb5dGwzBV7YilmRTRE1ClAih3yjmA0LUX5hVn3SB09Mx
W4nryq01PPAidu1ambH7a+TqF90rpk4e4Dl038ygNf3cMcJynory5mxhEMDq2XTi4CtkacQtgs7i
K2pk0J05errxhzeuP1+2J/S4OOSbZLHY/58z0llHxbw41cX9UqEaAF/QxPbXmvpY6JbAjJZO606F
mReb9KpmMgC+mXblofmMeZblC7BTGYhYbijLp3vE7p4MOcYahbam3Dcxq9eZnfQJpcXM6FUvFXKV
zA4yZ4MnDEDUPGuLDsfhHSW7GgwbRwDjsNNKcC22DlXZLJHTmRD3NWdw9aRGSl4vjhykelY5cBcf
FJUlrhrwHm6gP7k3JWgiV9NdP9YCBWAuwOXwuI2PIoCW+QGeGeQghijSO4dB10HqLQ9u/+3aQVEp
dgDrpFTzJ3KL6Ig6YctQwCxvhWHqoNBVhIoI2OoooF38vWSvhx8niRvNSne+PCpewIaYBzB82dUw
Y6TzVd5g3pFFFN1BGSHE9hhJhj5iNOQmjXSv0VOdA2D0tQBolK3c3tjny8Hp8hmGu3dUKiV7sas/
VVfVkfLquT7JwEjd4uyWjZ45LnflyinGVK5TQ1Y0aOE/R6YPhF3BbIhcUOnOrVnXel3zSspFojK9
Hfc2z+/DL9V2ws8QZzijPeFPinKUU40Fl5glqV2uUkBLffVgEp3SMW8YeIIdkZoJCEmMLMDXodkR
1JoNPtpy5AdXoOvgALE0dGdBO4eosq6G6kR1vPQKzeo0l6FoRTk+ufDH6e1Mnp+7BZXFqN32QxXU
zpIpLoczKDaAc+bIDWHfa3x1SAFy6zRS0jYJM66xOyw5R7NXVEHeOF/x17SbU0tM/ugbIbu32POB
g59cYd0retiEE6chucBzUAU6QQ2ESd1dM7Y4OJOSrFl+cMxURoqU0F3NWCmnYnQwGjLF1etm5GV3
qrkymQihuSqnFHKlL9zzNy68cOW0XUgm8xoWn5n8m52wZ2uK6ZkSXHgvTEoBWyrwEWxJmq1qpYfR
mPHJf15K5pqpgFOyaeHuyG0OZMM3ooF0AKsKktYo+0xmiDGRLycOhPSeLbB57pGlP0AKdM97F6e5
LuT/sqvugiRGHJ7A9Q5EofVb2tMx/4u40s6QzYcdWgTEMtegsUC08QnQrmN8oiaeczLApiT9nFMu
JVKTJDlm3/AJy/DDTrihf+ai6lhK9nv3EwGDR3Mfds8Rmx02/74slRMKN4BqbmSF873c7KqYyH8n
GcwTW2yHE6aMUIDEhuiwJJDTM+vhvXCkSXB9PN4nhZGC0IGHFJ7uqQKkkNdMBZqdoKjQRaGSZVua
T1O/TYzlLa75Gj8wlICaUh5gLJyncR4p4gBS0+rmNYnjQuoFipNeXrzUPCOg3zTSxA8okRFprJPB
mdORAxgeVuXOQOCKcIeN9dus50YDW6cxNox9Cf+A4AolEOogrqBp215JLR/TYSxs6MGEVYiZVJxS
MKa1fwuoufH4vJdr+w5AjbqO+65qM2v4UUHTKA1VYXbEYzHJOePeNrrHyzqiH+jeH7B6IPtc3rRI
tpSrYT5oC2nmYSkAIPiB2oa2NPErMTMMKab1szajTprFIyAAEoRwmI6l0n/gBHOCR4SgOuJOgp0J
+SjXQT6CmeJYLjqybO1mLMM3LCr1eCIgnxcg6QnGDKlWWXkant3pePELOc3aj8pkOpp707cT5lv2
K5EyS78wz6gSEuiI0Kxe+SqlAcM7IzT+hgyGLqQflqq+Vj3YYxc1bwx10ahUBLBRHtrwIzj3Et/4
qabmAJw8Yxa6yYvtQo3mzXmgI2+Ne3uaK5LA5Ba+lsA0ivZfoQeWuiliVWZ16F308Z5hBXZZm3GE
7acZY/H8UYXnU1oWdnJLXhoVTOpY+pgBIH1fq0Bpp2bFn5gB3tM2xAS+b0+Ua1aWaEwtqF+j1tNr
1oQ6gB5lfhHBUQN6oljvFJi26djmXpn4uCxPg5uoIJhjUMOTKlGyx3ue7A6OSyH0DjVumi0UkNV6
vXyYL6nu9Ff2yPsP8t15wfG8DptvfKFVBaYCVbl3INoV5XEaIxEDs7nSdY7NACMJ62OgODgh+MC8
iFFaiPICd3SGSOCwNOCYPwQSu8ee8EtX4bi0HSM1ef6DsxvrreMDeEdZJZ/zbacUxQPBQNksOtzP
Yruw1WEzNliV8ll0ZjmysLYFWyp+Q3KYJVsYI183jWz7CnRTLa29FDY7X6k0bY67HFZpCQR9sj6l
HWsXEQvVAM5PzncmLGVHIRm6NUZiJNzk4NCd2V68T1yCDrqyy2ubqRf6kKSxz2XIn1kbARgotzlw
Q+5ZfUHXil1D/XD2Ry8q+HAEjjTyb7QI08p6HAh8jZKIbLsUb2zj/4TH9KZIiUeWplyOAv0t5tE+
eGnPlxOp0poDJOPDZznGdEDpY+T1pS9vfbUSbn58fOKzmKcpd1iZJfWG+yHwoBlyY+hVX3HaDwpu
eZVkVppwCe+byp0GBdWJ/cTKyrrNW+CKMTDklFBNV90BqBtJhE1ZQpCvOCDw+GKbbzQ3mkOrjSOd
HU5UVm8anxgIE9xrbviojx/Yu58qojayiwhnQzvPndaYoQdXQUKooOw7CB+g//89Njq3xhn8e3Td
49xGXNgXQzMoaoPXk2UU6tjcoTvSl4BE33ItwVLAoIH84BCzMgoy9WcVsYxl1/rlfYmDvWQogfc4
EA37PQguwMDwyjMAMBJxysE1w38oCF8xHZW0dGWu4ezk5VKPnhKwTfAZi8TI0Quaw7O4gG8ID2Qh
HoQ5FBZlvTMDFhqrnu2JFZBm7XV7/A/duQSYlFyK+ORTIbR5bmxr6E4Vp/ey7Uhl8dSKiws5x//M
BdgSoj4SJsZR0GnNpWJzLwmB4Ii4594nknhoCH0Mz3aOVX6n4h7sRXgefXUULuY12G0z0uwwQu8/
F/dynKp2iUGzIbx4kn+JZbj579M+ySme2JfEfFWQ00BlMYu9vichDHLk/O5Ie93zeLxElQKlC091
5W3VQedk3SRPe069i0bJMrbHh3kvX3hDb2DmnQVvqRlTgStS1i45G7oGgATL1Mgl4o9KjnAWzCfi
GMDnM0xT27ivvYWspThDNVghI17aVlpf0jhGY7CGeRggDdeXdVxn6BMe2a5h7HjbvZLpuDnWTbeO
B6nqcF0deOOmi55SyrxXUPNLakmoTIG4fkYcyY0sDLuj+i6mMkAwxgLQ7aeuMuqzxfcH+6BaQkNp
WqdvNIHpg2cQqGVjBs4YuZKAk1VfUP92F5vMBgSvUybKqz7+oHPAJFx5lPwQ3AAZaw+4tA8kNRi0
/2Wgb0qR6mvUFwLa7YfYeR0doyUhIVw6/4pBy8Wxx2fWy6AgPdU4MuyVmqg0FyxpjWvbm9EC5dar
ac7of6opxZjqnF1C/bz86zA7QIUR6EX//rUbMyDWYmKjYiHpVBG6PESBjtPKofSd05yR7Lkhsnr8
dR6VDyL62jwabDSiyo+FXaFlPgyjcez59gEBApFIdEMOiNQWpidBAndGjeQIA6uGQZO5UI0NC2FJ
b+Kok+KNKpzyI8FjkhQ7xA5JNDLC49x2xwMSrw9LSR6Qm7g2QJ621C/eFMuYGtqXBWuyOCW30rhY
iR9DwW00cNrLNvq0obz32OCTKtnUbJTuh8SdmwHDgVhW9+WyvwcgMiaqpI0n7TMIvmrkw5KuHUsT
Mq+o/0B/ktxJJTi4pa7s/o5zt3pm9vBNIGOV5JeObXI67xU84ItbkUmbvxbe5BZc25cg9eTN71hD
cnqC5IqI61ltozD+QNUTPn8LPN0TBA/tw8bM8pXAqLlCei3T2QW3ovM0NyAc31cxbHzIc3KGZdSe
p0V8oxwHlL7kWO7sGZhbvHls4eVTR2q2gTGVOZxlvVm6CoB6SNhwsjkJsR/rgsREiRQTdNpVsaV0
RWSlfRb58Ec3LpMmoZQj63CKT0VznADpB4J+/VFRwOsWLpPTPgDODoV6Qo8Bhe2uqdqn3wZ34mje
Q8Mg2Rl7fJ7VYROw0+3BhbQFWvvhqFbjasPca/i2upO+x5p7jE/mDkOGxPdNTzFHH59xbuhTyT0r
jKl39ME8vgYFsbBOXPrk8hphfTL/UbsjhkdvUgHEJlT0w3PO7epA1LyrGJal0gv1waYSbdZcEO/s
IPM0GNC3xkmRzegTNrbreINR8dZjFnNHy5i6ObPbGyL+QIU88rXORO3h+4JslovdjrGHwKHrnh8U
5qVNXuVYAbPP5N5IE3QSp6q06Z3bYP15LHL8NRvADoHqTfCeMpWv0wdUiJOdqIdyWms4kspqyfkS
xmhq9fzcXaR54rCTVZSSn+4dRVAHtQxbgBxvMcTQw5DV8cV6yWO8bcmivPGFLFNKFh/Jsr6WH6RO
/NyPwxoQnXPlX8zFCSlyTJ2ZgvHSfEJSRattj0K60YcyLnVm12khOUpRaAgL8jXxePBUaq3Z4Fdl
mc1/Lvtrt/FiTXtEzZopqT2H75plHaBI0w4ELNOx5hKeLXUn62aRi+65dPWPFN8t7jOjv9xm2ZuS
FvUEp4VOjg3Su8EcBzIKPMoiygucrVPQNxi3o/HgfioLNQ5ISeM43bVHvyiH5nz+5cGsozoxjeA/
Z6W9wWNkHgMUo/gLSN+J6Mt3DpO0XRxIyTyF/O5fNHLjePa+NaO39Bbj0Gfw4uiW+XR+oARCaseI
J79ILfnTYUWJrPvsyj5x/MvfyRi5co2AGJkuymFC950XAnTEW/Hv0RLY4AqJ6x04Fbdafvw3a/m3
f8u5B4mJsmtE2O0YFDRvZK4j+hn80FOrsKIVneNuTmOhHAx+sQVR2yrP/vbew2nZpqTY3XM0qQHo
GeX0SKn2OS/11HmguZK603bBOxO2IH7nHM3W3hbCTjeeY7egTeV6mjFgdF8tFt3NyEZkcBAgiFvm
v/rAtU9Vg3+RfAogDYZu1YbhPeWaPszDUjqGJ2Ot9xctdRNjc1sQzdnJDdyhuFYBekBcECgUCqhR
v1qo0hq3SYLGECHzA80Lg5ZmjA5hdd4feZsmOBZPUIIdDDa+YRFqTRbk2Isix/2E3bdQHIGTngF3
nYOmSBToW4XbwbGdv5ETkZRbPWaVtaE5DTi9JLV6V1z8rPoxco6L8yE2haaHmrUk3iTshqh4VoMX
IWgtp/X2+GaYFG5iuN7dVp42yMU9xg6TR96bGbmMfu5oMYI9kmc13RoAHL7FMsytL86/+16vhzyF
nW/jMF9BWY5LrGms+SExyuvwWpGVdggaZNNRaE8iCt8dm3Qwu2J7tKyHUQ29ASYt480m7TKb24hV
J28/ByfVSw/QDCXYKPr6sW1FMWDaueCtdhwkT4uCiZDJT3hoS0T8z19ASxN/qmdgSNfILr6qd1b5
LLbQX0n7YMNmpFfDGvBSbJ0LxiOgflsRcSNX6RqEgjzDYa307y0D53YzGTh2ZU/9jUoqrIIRsfZ8
wTdmpG9zXmN17y6QZuW7WvmKGV8z1UMDWZyRc0/8gSi0s0JYwmwsljWRe2qJawXzeImBHt7nWU5Y
dQtgq3vFYdV2YpPln56qMcN3MZdlIVqzZtAREHL/0nCscD9JzXR+l2vmSSfKBSLcjqDspT1ar4ao
kerE/nYMxQeadhXUSgdhPgPWL16J8pKgOO6xDdlhRezOhWWh/N6+d9umcs0zYmlWNaxLrKIhznv5
7qO35HPqnWjnTNeIhokg8y4H4rLIgLzQwNUIjLf8NX4f3ujmxs+Gm996eZS6KqzGTVXMvZv7inKp
6Bnt11nIctFAHJJlcOz0MK0Oj7b6pmRL42sLBNHGJEJ2LNVRFx3wxs0Qd10Ntb0//Mt8cKNyTedr
p/mwuaw+w69UJSlZUeIgDhFNS0s4VoQpRqf+b+lfYRQ20MLLqjhza9QEdtGJxyqbDa1CA4BuEASR
/O+CrI2xkno6ler3yoPr8Wsmm+1RxA/Tuubbkho7WV/wwD0Png5PbLTDTT2Y/dYtrMhTiDqgT6eE
kIjZ78jE+3+2K0hW3HYYAmDZziDeH4LYW1vCU50oKjj0I2VqmDZqOo1ddixNbQZ4/wFd5h5q2U4w
GXDFVn1Gti6h3lDrUMxc4gtc8QaEdLVc19I4h5aM7ZNyZ4QthPIiLMrHMHZ5F3vJrq0jdrKvQSuh
ZM+R6qsImhF4Pkg5ri6k8UGq+nixX+ScA7szZG1fCbBysGKFQ/a1qXqMW64vyQkdG9TUugzsH4O5
gaMX4jzGxpVKslnQ8zzwk7Z+fr3uVreON3TZbbCv2wE7i8E9L9KCdiqCN4zIusuUDjRddz4IA2F5
/Vf9tgYg3Hgk6gIod5TBsTpeVDCQJp+v8cZR6TVJgnDBc5QPJO2S3Uv9xr6GsUja1Xa7lvCW0BQh
NjB2NoWN4Tu6v/9vU5VSoWI1OXSG6Df3kZWBmDSNshP5lHG6+5Jk9HcqvK5O4gvbM09fCj/TjEYG
BC7S3y59JMIiq2y4cpCUiSJJjq6B4nd/aAI3aAzjZhV0IQmTKAwW5sHRBbNptFzL6wpjW/PMv8d4
EFFz/eDVoLVGqM5FJ/0R3Wc7NGSoaCfZhXD0GTJYEQyeJ55Xp+/3dnDNm9RTy6GDWDlpI2V4yKrZ
H5gritAeqUdfOFAxfWvkr2rU4Qpi3NqhRfsb8GhVjXZumDMG8xQR03rlu3j43nHf1FM7qcU/goT0
m8lH6DYUpA8f/oeS3sZwN9qLBsprYnJL2aistvgbwEXPT2a+DkOiQ8oHMIgaDiABtqOHypFgkrq+
kYU+w5yytCwpqVl6oHYtAl8uA2tjURUVrYoriZZk9W2fMD1EcFe5ryFPawcuOlESe8LzER+IkS+u
3I692nYiZYvXjtsV5F/i7TogMY6o320uhVJMgc6sjkjtS9yFn3Xx1Uq2/moAmgj6I1rOZKq7BF92
4XZUgoWBRDa6S4APZ1LjiIcVq8AMSs2/vruYrwB749Y7W3SMV5SNoZwg+bWa5rTxP1fkgVYOSRec
1HVGrWFJrIpWMp2Z4w3gIbvqElHsOhJ8P79ov5UEvijP5wKiu1Z36mBpn9jmpGAwcg6jM1s70rvY
F2iqdeJfSxdju8YO5AKHvTWkOhXJRFkqE/efV+FOovJJaM/hFJ5Z/aUXgdZldINE92QJZdJanUTY
xDtdLnHRf5wa8hs/B0UJQLVcKiLnKs6bA+886zDLFzt3tCHyJOVkoZZnWe5CY8w3y1S61kR83fQX
3zPls1TsWAjAC5ZuJN/Mxxllz9evIyxvYFSpSFQcIBltIzyDIPcoyk+PY+k7amWXt8j6c6ZI2Gsn
GKpFAqVaaJT3VLmrz3zJSkva/lKTnbC+wdoOIdXecxjTCowcjCkltXQ9iMuvD2ZiMiVDeSPtn9cI
SrayYeeqKktEH6MpsS7BeE7eR1zPpCbyypHaeWWfmwByYp4NRI60I6kFm5J+Dm2C4TOgIOPwuHpt
UUgQ2ujcwPuASl48h+x+HAJZwVWdu/k1HXwAh/OnTLavlkVbZAIuFqb8TFAd/awHfRZv57E4VIZk
Ijnc7BnfvyUfXMC/wDY/M89r1phrYzc22iuZQaCtK07FIm/NVWuBnvlzem5wIi7ZiAS2nz8vR45c
azOk5+cuOM8m85smMee3rPafNxJy70y7Aec094owc7cyfy0zkItyEwtdZ91pPYkmRZXNOyM8TamX
udUf5gXK+9MGNhfdo7TCG31CIyo0R9ev9OsJWCYW2P2TcPfAzOY60Maz6Cqj3bgT2o1qELLuCVIn
NjxjBQvVWQCrUUzCWMaLuR7f94zPcvDawAt7vorF0omhW0SMQR9mvGOj+ZlA0k8P1WWtCyjYCJ6r
NjBxXACJNdm5kEQnRdzZ8zvEkmmoId/la7sY7Wo1XZQO8s4lwFMG/eE6k7I+9CvmQcC9ppO/g4Hy
imLrzUXmMs5HNaCBIHe1TssxgbBC244hpVwGWL42jw1VkI7xuvcOwDM2oMV7w/xHX1hYV2zNoVn+
/jS3CUx1rlwovFnOYrLWCcwRoCyTWeVuSRPrPgUBHwy+TPQEKJaZtQ9dblBw4fvabqBeZKUcid5p
p4wRD61wLbDKTGjL/g9qkblOg4GrTMMV2FS+jgPURY21g2lmE+hPf8gIDYZzvGK5l5gxUMM6wfaP
B7Mncjpcn/JZ8ZKZcfsEXUEeWIwwdUIOnPwLLo5voSELiqcr0bJHLFC96vaWQWkno+p3pACULSyx
RREn/MKfb54n7XXGb4eJ2k7LJF9TwhW4+OPVbx3Y9NqB08pt/lyH0Fl0EfSlYKYxrSLsXM3fDM+E
MUhdWYenhHQ9FIMvqKo3ts5gHMQhnB1jIUGYS+uW820KLuXCZxWZkaRab+e8nbzji3S9DHW/Eoh9
n9lWq630EY0AWwmI1UJRxAh4u0ixadqYbcQQ4FUUSN8YBCxA9q0T+pyXn8KeD7RTXBDo4FsNl4J7
V6ucwoeoLUtlREU8jEAJ1fwTsJUUqxNR47VTmUeuLnOPrJXCfMyds7ffTdxKXvOfcEKsduHi42K6
RGXKa8YeiBfpFGvMu3q/krT4n/ZNCjhsaIGd+BCGjdrJsJKPjtl+EIF6A9a/MTbrz4LATo5KaT2k
tji759c/poyurSOmVULgWCzKWSpGpP0TcJkab9BOexseinfqAwyc0E/xhl0P4AN70//gUiLd6pvi
gwdkTH3H2aqAAfi/gYWipL8Orysr8U572GnQVigOtD5UOjQv9YP40JesJo2ooH3CvmBOocChn9Vs
mNe7skzenTlRq7R6IAhV0PYsEeqr3Io7u56MXujXw2BBcE4U7TntsoohW9N1vjMe2EoyepFEWUVj
ksOudfaRK8tBduyf3BhnTSb77PNQ1cylj9V8lVM3f73Uxw2qxqaEmnu0Xb77tcWT4O7vZM0rFjrj
l6xVcKwSUQN+fwPGP0/U9TUSsz96q8wQ8qOCAsbhvfQxiyTz8zkTKRbBlH9VzGCWT7W9+mdaH5AW
OsjMPxEniwxMxr66Yz7BrwnSb6CowWRB6G9mdTXdrulj1F2sEUj1Hw2BLw5hODuFsQKwmu5U/YI/
jCIdqG9v57aRnWa9xGMUUGMrlhg9WSpBEDuuqEZbt3fzGDzJUo5FqB7LDZFiu5Oirk7CByaZ50Sz
qYvzwJOP0bcoQ9AKbpTBXlfcPSllxRcwW2q+1tMsBZgm3XCCzttRE3cUT450H/3L8LRLS0+wELKc
NguCB5SLJpvIvW3puCcm0kpYiOEVwdflr4tIlg5bKvG1da9tjbEcMe8oFIUsrD9V0ijZGRjKW2ly
FWiE/sPmFLWxaIWL4tC54pKWTWzvkjh/Xe9oKI/8d10p3fF+p1Akz4kJw7xY2t/UDJ8mDe/5mw8b
NSoyEZIUhvN1zj87x51cieIWKiVi7nOuzf0KZJzkJ5ZaNDaoIseIHS6/fKpNgp0IVYGTqX/u38FK
DZ5tooterNLRcpG06r0TfgsrhvwGUv0jjhNkr/kkNSizzgpf+vXSoHE+rbMF3EXb3b/2wkQGtgg8
OdJOx5hm36WCN25efZCyCzZRqzXN8EBuj6zACByQgPoWF0tQjnMmjlPZ7eC9deH10b/KRXijGTCB
DGla6xUYf8/dhj4MfNxUc+iKs0Bl6R/jUkGQgVanDWx7AkKVmGvU426HbDPBR7nX78VjFx76L/Fw
/T/NVQilRXTBGYmIvKW0tiOShg7yEwe/MV5EoiHxaZ5viya1FvuDeh9fl4/yqEjJbCJXrjeV2H3i
I9f5Y6ZkNcWI2O6Ml1u66APwqO1QcIhleyYo2GxP0wSdPO5pEqC8FNm69q8/1R0v9M8EER7nJ8CM
1pzfV/vIMSB5xgWQmi8VdzkC9zUeVvUkyAeSUouVFnbk5vqBj8UV1F/VfBtXAIgAz8ldAeA2Ur7W
gOQt0CZgmoyJiR/PnnsxmHBs9S0AoeDlGUWAkt7hkCbeBeOZW391MD+yeIJd7yQUfkwWl+UiK0m/
tGRBQO2deQZp2Aa5cOB3OArqObraeT6vxAKSRB3IHnM+kaNyaKC6INZ9IFrLeiDlXm2VjEiVx6Gu
x5lnPNS8lsizkrg8AIO+/v4HNlZMvWK22xuv9TURDyWup4Gof9Ry23LOE2061JyqbN9o47/9b7Cn
stAJDjDpuGtyn6BPeUL2f/NbFy7x/7uh7T8pbHiAG4C0zH2F49twKSQKLzGgvgnFYTAZjCAE47zt
ODFEgx1PcGWDcmrM37Q7aaevYW+ZPlEOCjBIFJGUAz74C8PHB2vlJnNXCbyDebEPBqX71kjW6PwB
UXsvUxoQvDmlzaI3F+hFa0vykhHgvWLJO+ku/jJ54uVZVue5CZOWCkiEK6HCV/WXuEtWzsmkmBhd
Mhu49HT/ZPjQ49afpBnZmv9UBHeBc1bMVhcX+1NpvtS5Q3F9uMTKAF1C1MBgEKllRqc2vjz0E5lX
JucC+Io6yy4yipViEPMT2Lo0oj1v5YOjI+5uD68uTPbMW1B++KfX4CPhKXm8UWCQxiRhzanX/z+G
54iu68/dhaWo3sLJ2VXVipew7FQl5F01evDlexlAI2GeFwM7wVE/xly4X/pvMRmvB7MsutOp8KaB
urzshPwt7Dey+VvIfMUV0C33RLNO0PPNgAaA7cACzn+mEZx8T6JEmJkXo3J0kXT/G2htgsSmRUhd
JXoSWekgINS6dK4LQ35w76zroHAnUMD4tKb4iXWVjsdUBBBUKC2Cpp7UwP2pmu63EJAXptKLt7aJ
lQjDCpq3+j2a500cSWZaO7dS96G+bYJG67NLnGTXjeAur2QALOLeHytAeXEFg8meyUpqO4oXxaly
hzQPRqO686IA16lhIVwmNEf2+lbfVhgrldVbRp3ssx1IovxLcvllxQaeeBt8z1u9ZIUSrMXARE4P
PT8+GKksyhFnK1ohtnzYtjVAbHKnzU4vN3tiXyY932/PiOv310hzkpo1wyc8J+QIN3Rh5L+hdF3s
qWUwsgPM0qfYaSGphRTKeahMvXxaAdaf16EUs++eaLI7r5aIS1kfmIaEa+2uddfSat9oUC+apsF8
H5sp2HyB+WMd5/3bv3WVIlot4jBla7i/jvdKuk/Pbozs1EWR7X/7tsAcN/qi9t0DLv5+IRYWHP/B
NZwP7iTdFeAH5gntGkOeDexuFHe+mo7O4VIu2op+hLaiJXtSIQaAe08VCpFsAlzaMa74wzC3O6pq
19BbOhru3YFn/0utk3wsG4/sf3CrSO1Ed1Ptaz3fdnaYVtsBPaVM6HzuoStqKUtzHPF0pVzyGutF
ouvg5V1G7DDW9bRjybPDQausg86olAPt5aJ03H5uiED9YAPI25VtOTPIkb6urwm0BwHvQzFUWxrg
E6iFaArJXvAsog9HWkGnmEqtGbOoyk7l03RTN9bpFpmGH7fmYBRVYqHexiF4KrlsNE2lPXcSY0V2
N+PBeqi5K7wi7srk53qTw8p6Q0ht5rfahMQbR9vq1kn/XDvxK/lo29LgCWxeArsrJpq2xFwKaaDe
Eg3zEMss40u7qOcHt2zkN5IcV0D/LN+wVgnK3qCz3kbSAgtNheZnplefumLmsTr5XfpmEgAyhsuY
Jj959Q1eYkMN2RHpPF6rQh67rXWPBmBp5wHCPQRSXF8yPo+EFQ96nT8yCPQ72Cz26PV1yFaE7bI0
MgvRu8zATKbg/FCy2TlhUyEzeAttTkkf1iNg9rHBmW6+v4E8ApGIdiLwLyCN4QbiPPy/9hHiXdqA
LhP7/DpviSqa0ludMy+UC2YK6aAJ7l2t/kezkVA6G5uIeeswaWRCJQmgMg8pp9e4lPaNqBmYYCAd
nkKhr4xXuOmI0UMKo9Hs/vKOd39eyGwdlZ7sDeyrmWnRa+ri+vYasGBWBPMoQBFUySmhpDBlpL1W
/Ws1rcHFhpb2LMpGjPQ4gj4yaFNpFgnDJTzPD7ebmp1t7bihrk7kwbyf2/nceyAn48sjMjkpj08y
4IBf88qpcEvm2UEjiOrlL574DquyUEIeBflGsdzvbkp/yh1axWmZrt6ihgkhb7l4VDQEjro51mlq
TgEF6UjSaAIl89PQ6ofCsmu5D2U2ROMiW4Lf3oMCkUFioR02oDP45IaZQDD4Qwcj4Imp+97gp34N
KaKIPr/xTardT7tqXhMEoA05p+yJ2vAj5UDVVIz+hi6MtH8lukK6HvS4i/TkodylWhe4OW9fFmYV
yK28B5KWjg0sNiBiEO8j6TZm4YOxxHAEorHLBIfOcwAObNaratHp6Q6WHW25TkOZY+w/tBqn0GvP
zPQi5Wx4gmQlCaREI3xgdEA9f/OP6I6Ad9e4xs8ZUjAM2wiGqYRoJF/llYLGCKKY5wZ0KvGjwvVH
ms3Qq/Rb6jujXyqVcqGrgzopp5Q2MBiydhj0SRWQLEOeZiEr68pM86Mk6MKL9VIXrKqJjhSgFUN8
4ccH/J9wN7pe5waXBegUmDBT93wY4g4IQp0ddQBmMm3Z2ZskcsBUhrHVTMAotUXfhSpdafRIDdzt
cj4a24PUHoTTbEAOslqeTxFzcO3cvzMiGXYuMl0M6AL6qCRC1M3DD3JeEvAtHCOsAyRw9UGpPX1u
BOBaFSvBi4m0OLvtawHd4Z74Zvf9VvHO0+8GYRJKDenAZKoysFvxLPlEn/vWo5ZUNRz6O4riEZBt
EgRd4ocmkIehoByv9ZInlnThLUqD2C0hwBOD7Xy2KCLIrdSQsT/Vpq1g7BP2VBRKukbXna0VldOS
L4nw8Y/zVE/BAEYRAzm3GY335d0DrIcO7KuqXk9mLZIwIiASauiP2oGcjZF21XC/k9WI8wQuW2pP
NofJPAldW7k3HPSWW9e71+SrGECGnCOQrSduRdm3A5PaEhRZtDi/IcqMTrJFRliVrftE33AJQBhq
MfF+gMk1X2/jZhDgNscczWzj4dYdmZMmt4bvEa1kDQBZhtgobagrSHUUiPqhzHSQ2F8PY2ANq1Ne
jm5/Jag1/uz9kTzMWHEuF6aqUkN8XQ9RkqcAqgUAw3/sXKGrYLi8bpXLebrVoGQwRLm/TqfCpNFP
k9x6wLfEN4IyEJC07EEyxrfWpSmlnTQY+mL/jOoLDhxI11sz2+gGGxLDW1PMemVIFsCekkZVHv2M
hYebK/hVMU5KRLKPn2milI23gR9L1EQGxi/fhK1xhpU4yfxq1R+ld56GIW52I5HXVA1gdT1yV127
5csY/B8M5/yFDTY+TLt4piJUzqKhR2sfkJJzDhryWQOVZZmB6q8E1QWwe/2/4r+UbSZ7Z6pefUQA
svjl2t/0Gl3h/AMZExa4xm3Iydlqm7jqG4Mg1PMDYDyovlZ2r+o5ILa47d3D/T6Rp1UX+oAB7C8b
e/If16uYEmr9L+w28LLOSY7UkpKlUkX36Gl3MX9tC083v6EdJRoDOhZTmpCXYbDLqSCm3Mes+sCw
vM0Kx5sNuJ9dLIdMrxtuLnBf3ZMFHCxZ5oj4MhoUcpvjvsVfdYNCXEsKQ9EadV5+7GJiKCPaDxXX
1L3huA1wjmvTSE30kLiYLfKcbWNq/NO3+b6SVNnc8CJbco8k/nF8a42doF4qHtdHw32w7oujsKIB
KbW2NZuGuWMygwHN9dhrwKjkB4JDLckE4XLD7wsFUZosFDtf4JmPFpDebhn09UG+U0jWOMfhT4YN
gFL1I7X9FpPLzln+XCUEKLo5lLTB2Ha+DOL3KnIaWVuf9CKd8/wTUZcJzP9P/GYy5QWnvujAxboN
WCd7rLxifGve2ttaeKwl3/Ux537C/dyPcyXfqdwnoXJdBRiZjbHX/AIHeZPB8aE+jf1EDpooub4R
jqvGcZRsdGs6wMdJUbn/kAml0aqUoOxamxH6zellij/XhLPNb2btuh7jaV0saS8E03G2yWmYNijw
wyc/StRLh693zZ2aO6Ela31HFVOXQNGDiTzjEGCwFqobUWTTaSIDsRXSj4dG8/GpQTMlQUpPFVDw
qUP6l3uOHP2rXZ3DQfvuh+hbZH2x5jutL8JHgE5l97Kv8XK4+5Gne1KfVMIfwD2EKHF1oIojP1Sj
BhddTOs5nKGu/13ZWFw/OiTgNtFlRTIivCngUi6VkbO3aVcdiuS9xgyl0JKN2xfkWFa4mwXoxV3M
enypomuLdYfMxuu/6jfHEchsgwWBlRu7UiRpuNA0lyCbOoKlCmmm+r1qs25QyLCzzQVKwwLLcmdO
rCvYepIYchNzdC1MRrKWELLV1SaOMWSx9rKi7w8yBhdmC0eHuGLDb8qKbnCJ+8FswTv/eQ0wVszz
fHzNqYqy7RsWr82OiNZ+qmg2XL+CbWK6659NoJ92hMsKu6tr9OWPZKsapn8XWSXwcRUaHRZX9nl6
C9IzyzDt0F7w2edzxSbI5aMSfaEfwsIKirvHjAqjw+QpnK5LOfBe2X/byN3setAWGeKTiKT9eDbI
dWvqsly4owRbmS1Wq67e60uSSI/MNyAlmBrKjLkyubiGHgCBL+ZZwZql3tlEsT4uAj4rGNQ2YwRG
l3DyHKupBVGnpi7sqIpoPn0kw/PUBefigTJm7zXzOgFgsnXehZVuWYhG83l7Hkdukfs6DHiKxPl0
kuBdUlBfjZSNil6LUp8W18b+9hGBariMoVKTUwDCNnoIRrf+032B2DlfspgSVY9lhkHv3abmpaWB
FwQ/Xgpgec9bYRoiy0NJgtvNkmHTVdU/U5eA0fILpoxsokGU5D1aMqy7Bn1THcEf2KclJ1H/9eX7
S+UU/+xXD6vQFldCpDezOTtld41fKs7/FAfou3Fh9uZeAAMGt/7TgVt/QEJxbCtAMCNSXoH8OVo4
bxQBXdPmVskD60Y3k8+XNnzofSvGw+sagwHzxjbRUpTrgomvFrHXDn9VLWyQhIKAUsUuMGEhslMN
9KV6RErBxXjRrsv/EN+tvcs5GRsLGa+H2la2OS1crum855vFpfP+6ebk0YvCRlTPNyskrXnBaPAA
0rLAJNjywrMq+V/BsTupSVsVWyDE5PPbNH/bJOVDghUld1Ok5t3rjcu3MQ5Khd3BJtplHQDfGoiZ
lM2q+jJ4D7Zr/iSIkISxRCpakY0gmnbJr1uvSHlkjseoRZgM1PBZd2GzNSffSLRgRHR5mUFN3/Lt
gOXOwaLBYu9Hb1bAVwvzCeBTENoAh2Uwi/tUOGu08qc7+AijpbWa1oG7nMV7+l933WJ82WWni5lr
MSPoD5/AnJw9IQr2svVc53jun65ghIPM9NSQX8Ie+eVaEbZ398iuCyjnMmlhUKt9ky8fFYEzTXpr
x0VFTaBPZrKVcpmqquc7rWq/ZmnpE+JoN1uavlOVUwTXyShfXXTun2eGx9EwFLojlEuqvZGM4Zx4
N7g1MNuCLi1xzkSOLaFJ9O+WYpFNYfE3S7DGUC2BVH8DaBHJvWaGM7CXlPyMEsQnRhC8QOdGF1rD
im1/F9xvIH67h4vKTRn7Ti0wSmK1b5Io8bHW3otqIzUSetLjL2PNUJt5RjwFM7JbMOWBw3xc4lVA
SXceqcLMFxrsdHuzBcPp6gwR8yxDeoPFUfPyo0VaDHX5mSl0M/5WwVXXvv8s67JKelr/FKFcrddJ
DevQNDwtsR40z4/IB9kKuzQCp05rwldwNkr3YHr7nh8bHctnFuiBDG/vI5yWxoVt8EC79tTQ4Hty
t84ltbWX9h803M7NG5XJ8BHIvUrd1+oKfEro2CSFzqJGSYlFhaC3BaZf+pvwedUYZMZIl8c9GObp
9ZkO0PCIFZdTzFw/SQfZqtdmfTTyXS+ZhUuFs1ygKsO6knGpHfDX5p+jjq3GpaUrs4iYj3o/Vh6F
LhFcyyQ9iow1/NFmVB6EZ423PMuISTUBr41Gqpt0ft0Qg3viwPdLTNq3WQoGR1M4KJe/MyUsZbbl
7olyJpfn9L9+UigLRedTHQbomcEWMA/+nCmpmHFj+d7z2C/RNSzUCvGFS4vXaV/NaDeIknm4G8Ui
dosA+AyvNMzwwau994X70OyMjkxu5Kp9qLTRxXamgk7MiPavygAQ6if8ZRuqNyc1/qQVVqQSvUs/
j6CIGp9Hm1nr3qR956BUMb2gIQ/qNaMMirbFzd8Ifnb+lRyG6XfK5+LHId3x/LeMIhrmFg/FyGFe
Acj2ma32PfOYkb9k9u8rMUHrOIKlDlCAsrGJlBlOlEARPjsVDEZEY+FSMmPyv68BHCl+hu0wN9U+
pkCzzJo3qMCb4C6wcwMlnx2M94clbF1S2pCmuy0ii4CsQ0/zo3Kdldepjm2McKxml592zAN96JNE
a6BmgGAePkdBMbi4uH9+/Vl9UK/FnnrI5WKY+maDfMZ2ci06ctQG0ZxsVBoHJzr8WBQBx2RwlIme
hHURX94+rbrfZqYpXqQByFb8jvyvj1824P/ElujMZBWuOGSGQ111+hlG3AiZWsUeAHkzN9bum/2U
9iY6Q5fHE31xJ0nTzh4tIRfUb/LWg3fxUEfN+BZmOXX5evuIuipWlQnRxyzS9LEYGkAYFGCUleRd
PdWHJQOJzGFxCHFYCedk87M3tfCVaWv5M8B+zU9LOg5C/AQ2jLW7Csw1/gDT208rTT036cIakrP9
JOZQ3gZFGhkKTqAu4N4MUsTB5brYmGaME2TmZWIIzxbhkbGGl50GVSQqnTL6yeiVqdqCz8bxCBd4
+ECgXn+l1cHwUXCGe9sOUZzmWB4NjTACZUVs9CWzgfzYyj09qmkGtfPTkJHjjLxHFg89oNqzwAsW
Ll2R0k9dQX/+cT2QXzEph8j/DNyD0Jvqpw2ZO7a8Q1b6/+5TgVrgtz/hs7XO5TGdMFC7s8RdR5WF
9JDOyEH9k22+vpDD2WlYIDBvVbj1qakgmZrzcEuRoq2FEpCxkd4ydje5LwU0EIzcah7oVUuwxOxJ
JpUqnkmBYKt3ktMfdYjMvxksHV0ttuqbaietWoIH/qEv8NzWeaynIH0bMWfsWa5lsjrhO3bJz5HC
VunBH4Wp3aJtiQoycsU5IH4HcnyL8YflbieuPAh95KG2q11ok89d7fZoLArkRy26qej0GyTDrLn+
abvovolriiqg/QE7ZsYlp1GJW7WX4SCMvlwPz61keJ3wvqD1S5ePf8kLcf1sQoHhCLzWCvFL1y99
QDYljTj+xCDvUJEhmMkaB3QXmarwn875LqRfB15ddUjwGwV5w7YD0+mXxDNB135W9Q9baW0GPe+5
mX5ZL9qKjqmh637geNn5YMPHli/BEQVwaY7i+K3oj85SNiM7H+BKhNkb86/kI2a39tbLFtgOlF70
SyOfPZsoC2CAnW5F2Q9A2vOON8h/2pu9DBlrrOlIHUJkryXnCcwKDvEapKap2c39CIv0+EO4wyPX
arJM/iJmmQ1x2MhIrwI3w2TGJDlh6O+Pgu2dVH1l/dCvo1bFyd5hTtXXmqUSCnm1ZJNIr9MF8pbI
P9v7/25lmzr9zFUUMxOiZ0GopXUUHcTr/UMbOV1mwp0at7LaufKEzZ0HToBlCYxZQPco/W0/lnRA
DJOoTW5PyenQCFZBQRnb3UjLuJhk1aUO4xRu94dimatPZWNgCjaNo/y3D7Zid9YSeq0hAq+Ajm/G
HoqznsGyXa51enNKslVa01p2p+EtX+x5NFTErbVf4uE4Q3LgZzt/ljrNGcVxbJ9fr2snKdNUJhWr
VxOYOzUkwegVi4YJ1VOVmNaddZF2mJDQtCQVWcKuY/yaF9mn6W45gzrX6/MMpHEwjs83YIdqZtx7
xcqT/TPxWeADwU1cyu5PIs6+BZRgf8Zd89HgJfr4LgY2wos25KUYx06BKduQ16V0ap6/HljOW4Sv
9utY990/Pp3bALIdeWPX4DKr99basj+i4Q4TSJ6dm1rYwEQeBiapsnNz66sNSgT+xs0Q/RZteYqL
OItng+np04BGCzTLXb1dXKtpkG1rSoB9SkV+wzJxROpfCSVJLamqcszi8Id1HKakgOk9yJoC6h41
/d24+dTOPqahq3t6ShKadM/nduoAncht6Vghwh4rpBUdCzYnPGYAKBL3FbqQ/8DsLL8QBgXNWlp5
sCwkV8rOvvbDIe/HRftFie+Ak/BPYqWe6C0emJKeFkXb2zHmcYXRwAV3jWTvkmZCWqsZIAzceGe/
HF9OFU80GmIFzjwoZMtcSqFiDx1vKxrSsA40wiFWqnEshdF007yGoNjHweMVSy3ulPe7EpT2AMgE
Dvayk9khA/s9pfngeX7MRY/hIFgzdkmCm6J9Gm9UrjPS1y24v+aSzPC9rMh+/4h7t68prqh8B5QL
NHpaM5T6mNMdSqrj+vp335Vzego7etZVVzj14vtnIJRrGpJAr+nunbADHaJZTo5m8SX4PvcudgJz
+r7kuBWs93A70fKdHr64+5XP81U0qUazgsDxr9BPzTeB9dsLTSayS0gnoEhbsXs/R3nA6lMYs9wB
QR2vk0fkz7xhgqfmWnF14dmlAcSW6KXVAdhTwGTDjE7/DgdwCs4prarMHD/N0Zbjknc/mo2s0O3k
dbB9eeEY+BD71ob+iVsiGAwoZ/jc0YQke1PMNWB0yWF6MR9Cqbnknpl/ri9BecJ04njz8GUsQY7C
DdHUaFtn9X4jaGhmIIr9ZPjdsKKiZ7kmpfntVkIjer7W5FlL3+jbtG0iCsUtZADNn5jQvSE09m7+
Jz61838amqv5yLbRouAOTgv6r2BNX/jvz6TF+rF4j2RMzyqLWv/s4yhsuFLhBqNVY+POo3P2CQqf
6s6Gn/ziVokxhc8uTaiGiu6rYcgkEHLs+RDujyvIP7FPnMl3F2mUPHuha0Y+uMHmRraOM5uEdvjQ
bE0JyMD+bVGMOrF9MhJR2ngBROlVSNcOrjRLt6o2cVHzQppRVBWwRpf/v8p76JY92yuCJaFB3aNt
eqxvYw/wQVg7kmtn9vYin5z630hcsX8ZFMwOosbiJzs6f2JFIpyAtQ/4Urt3mlPmhuXrcHzA7GDK
KLcOixJqBBIcJZzl43JaR1TiKQvnod8+cjehUjQxm6HTqxT8JDiaSYGuL7HAbWadx+3Ih1jirJcp
einm+u1hSStkYqShvANKe3MCiyCJU+Eb4iRfXnGa/xAh9/Edb2hxfl2ZWF2FZMBeAOin69FGlt0/
Hg9MU68jq4dkgZrcrBWGs46GADoHbnWJykcPQnVBXEmNgem7i6e9rEBdDKDVZHHRN3Z/Q0be4MK1
ez0yCY2n14Ig+GG4Z48nqyv4Mf30Ijw8/Ke9r19m2Qz9c7HaM1MeIcZsX9DPnH1odZp4WyPYrPVI
awStYgKRVFSsEtcdi5HSh7rn4htU3h0furWTMMtVbBxSxehoC3Cr7CHpBDv2lgXiqVyhegkhIHts
BNZVkTTt0liSY6EmW1S23V1CuasmCOEI+mNlwZzTVvLW5Y3gWk+HHrDVnb869t2QVTA6GJDq+ebJ
O4btq3fNQh8diuTnAylpuEloGeFdyte9xiL+vIOUD3KDOhBD8Tl9BBFGpiCaC8qV0yoH4kQKIJqp
o2gAaseU57XpaQKNbqt7QgWm4VggdzYQYf+O9T4Sv93Zhx8EMBFllyiqkgLCrHpkWDZ03HNUh0+B
8OQ27mSs3wlOP58QtMDm7xu9HMELvBJ8ZaqkwbWLiBno349tRtUljXWY5XUiiQlaZ0Bu28KQVnog
S90/iwgPp3gQx0vnMrU1Ll9mGzIPKnVBzsW2kaoCmpMC9eKPU0Ny0R1w9/5+ttLM74j4sOVyhYMz
wwBTrWtajxDWKnWolPQg/oZzVQL9hlFno8FK0j6Y2FbYbIFslOXrWKVCXEn9QlQvQBfvZkppTz+t
hUz1gsq6rglkw2tXkUa+sxFgX2svrUzCZj3BTcrzLYzt7TXxPKN2v19LTrJj84Ib+/gEEr5T6slq
+x7oZnirsUeodH2VvBU4IL/B3SFXdIoMMfToz+IQ/KeumRAoTbkL6L+jHDA/l5BmZgDjZrIiygnD
iD4YrYQlKdFsuiCppZCmRRiF66dRgz/HLMde8YrpB9xePrEigXQVWEWvtc/2Az4al6G3kom58g7+
XkqYZUZ0AJ3FWMLLC4OJMv1dhQNsuhQsazZd87pw5Z7ZAueWuQX3aN3BifNVxlk57RZeMd/obQL/
6KoG4ZGt+ZcW0VS5HL2tB103WS8S4uDOSU0N63B8Iamjvzaxr9V+vbMNGUjlcL+7nGt804n7JjGH
R03YeQ+FKO/K+O5J68TZApBhiMZxsrHKkNCDVKlxz8H7rpnR2slx/6gB1/sRtCBaUwPaznv3XAdO
H8A+TJtOT+FiwM2tCbrhjYGl25tgip0YGXk1tRqJUqFT4dwKo2p7nLqdhuWZXL7BS5Dj80uNAQXj
4T0BWDV/Qj2hLQY6XaQFEQEDeUpZqU59EvkhXnDtWICQl8nJX5axEk7KO52tEEvqypEDH7Nm5zzm
5704v4KYjIO5KHLMlRRgNokmlkg3UeBqZGhDnlvHowkiNU14TvFD18+bYR7s6tEARgnFwED8vVLS
Y8vdZnhrYeliGlZt2YrZL9c3/ToFX4cTl9ogp6FjNxLcwTOiB5CwtVqs7z1YCLg9dvoUYNZkMrXR
OPkzEry0oEkrl5zva32H5xsnIxIVG+4VFKOEHPQIE6zbbEBn/dGFb4pGlDsEw7OrsQDasQeQrFdA
GQcusOBD5ase3K5LESJA2YrTWE2m7B8LAa1sR5IDuYGwh4QVTFeyY6mFuVH3i6hBaJxAI1c2oDL1
+TXPxU62edhQ5wcafZ2wi7BdueEFQ6deTwAUi8babAg5iVY98fn/+m9erB2CwBLEjNxLZc/5eF7o
6zqhjrScrzRnnrowrttvM0/qzJgQ5olKTOJXFIvpyZuMs09fY3cAlnHCgHUk/9Fd8bXWhlYr9o9O
7SwRzHWi64dzkNWYTY802XUdcsjow341suW3yDlZmjg3jemHKZIYOltZlERF7TiEF4YJK/sUN48f
NeviI8H9zBzhAhZ3kBHyNP1eUeriiqrVDwK0nvqRB7MgVK+cn755Yd4ggno07y1N0EYjKC74FmQe
+Qu+1fy3dp1fcgT46JghP2+Waz0yrusJ3nxaNvSZ8v3BxMPqzFOnqSNlXkrYJj3AZNEd3AXlOf0P
b28sPIZcRoRZgxf/Bye8/GfSLePjNtdsMef2MCpLldvAQ91ouzwtMnajxDeizXvnqNbtLScaM00i
GwMRG0c+sEmvykJoJVRFvL9ZgX7X6jrIKx8NtZCmvALr9YbPW4NMky+wJZZV7m0ODf+5urr8i506
TKNExwapzTEyubeGsAItsfx2xGsshIBQOUFjPnGD+kvgYOgrYTJQyVIsQm9LqrKn23Vj3j37wFUL
l/Seov/AsxYhrIt/UxrkVrncYUD7cBwo3mmvBi9YnhJWp8yVJiPw4+DJeWijB2fJmZKc4dYUWdbE
pERbOCVwUf4cYkdgWEgU+h9tRhVXAnXCESO5MolqEkRnqlZR8+ADDldgOUR9D4vPrjoC+cyeeThW
C2HzsjpaT3CIie1OLfR2PiHusfP+FrRa8sK5oH92TBUPZuUpytPR4ocEPVWQDusKqMYjnUxJ1U1g
Q//krssdjMP1FaYW8YdqeEDxr2cbEDEgZ74pvju0rS8e5AxToV/WClr64ulj8f0N656WJJPVu+7d
Xa6JRPo7ZOlrIUXi3DiCQLCbZiUCen+Srb8MdMqColyt0AeF9B9nN2BIz4WxwDDkoZUQ6IX7/K2Z
0VJes4o7NzbEoGhbrwIIGUNsVoaVpC2lUJvHob1vbUO47a3EKqXPJBK0CQ/qQ+2rufdu3E9TufsJ
SSxLiJ/Fjz/bwvz7SW1LauzXR/TIiBewadIvKf8/J7eeb3SAfBjyGeHm7WMXpLXtMqSJFJ+h6EAK
gxumaM/CUMn9UHhAEAocalgKGDAFqLKwUw0AFEbYNQcvQpWoVAMxOgViBJatqZAZu+HalC+RErQ0
3A8D4c/+mam3X/jkQFVEChK8k/kyMqjpZnIYh+whcD18x4ciZiRT2b2OxspewSPoNFljqO41CKke
dviaCVoDVKj9Fwl6K5WTvEbI3WXvLr4l4PNn8G9weW0CVN+lmz9wCLy686QDOMnxZpXAramCxuyM
S6hZCtIvLUeSxs4DUJ+YxXauDMyhoeQ31958f94VBtHxtZsNzpWAZw1MhlvXX4fd1OHP41ZjKWa1
wRzh7dm/7IjE4dKDeu96Eey1ks1TTom5fhJm6mLh/s4SeEZTocX/diXj98woo3mQGqDbQmzHNrN3
DNQnbj51rnY0arRV80v6wGiMz8dtQfaU/zejMRTMO8VKwJnqHYCVJCzVhmGERIKbtP6e3i+ccecV
/oPFkS86uAvU9clrrAJPtZwwX9vs78cyZsFMy/xbVhrDOT8oRgh6Kf7Ah9qw2+5vIsGpqoF8+UCq
jYvI2Ox3tREJmd2on5hLYWVWF5k/IqZwR37Fuw5LAa74hrWujNK51/7fwy1wTHENXd5OPnUh+zvu
507Ub9teVTcOJDIGSjWtY21GaxcVq6GmGBFdjehOjaN0li+MnQI/VQeCtC4mxbS1Ne97BvlzpD4o
emwlMQodzGCjvzfh12gsj3GjFmfvvCyqq4ZyeeLbvoM6XqnTrqVN/L0NyXlhPa1/IjLtA1ueAQlo
PXj3MiWSmnX4RCRAe1Qdsl5EMaLl8EpzlAXneKciZ1w4P0GGxI/C0T31VlhrYXaT/XsqjAkXOaxI
LKRsqxgzdc46Wxvg4nmNMXW72Bwr9WsMB50+VMxMjJAKZHBS/qx9d9Xvh45VwKcAahObx8JQTjJT
2U46Fd4683Zuzndjb0iJ4p3BbThTqFbHs7xIK1QVH67lgtH3WJwSxKgD5gJOrG16mHJZcnI65O0+
RGDcd8h2sWhgy78p8vkcWY3/T/nPupvtNNtAZo5yKjat7Q8A1AwzzQFq9ctDakAuGAdVCJmHThA/
RDQGemgan0pu5l6Vv8j4xUX6KPpt6C9bxjgRoFIv1uAIpNO+wUIQiqdrHlf4dCn9301P9p62gCso
WoOYrBYvc4WAzH2x8lPcSeo+W1Ex0NLHVfSFy3N4d7BBbqAfZWw86j4kfoDG5ymG7Qaws2R6d5F4
A/rLVkzVclPD5Ois54149sv/Kgi1A86aeLRsjPqlxJeRGAhc4qW281qC4TNol4IuQ4lxLqTiLnbM
Kie4L4EtlR4UQJPdm07fEAeU9D4ZiQca0s3u5wKlOzCxDJW4vMuFRK3E5F9FgJMgklWzTPnnF8Kf
i8xlZa77hADRixLl21RoPn4n9kBvlSny/mdpq37ORp0sYeW9aXyMr7eRjm51hUjmQ5v1Cs/hvRdn
cleGC4Y6TmHbidYzq2kWyzP/bjVvqFIXa/xvIORg3lONjXKHmmZ2QiFVF/dWbUhLKTDHYezJEDhO
acJ8UjC2OJUvYQ5m/qCxn2q0uR/mQeftat3EPL2y+RRCYXfxWZfelf+VrJIhlEvPk9hayzIMvnhH
1xe9h3ut/z+BHB6OgYjjAieeyt2lgUF2rpvEBfqCd2QHJUOebipDbJ9wv5F9NGKIr5cy9wxTs2Y/
kB6hR4EkI3rygEs9iurZxwn2+cn1Pi0UxPO6lUanFRth79ZOnx45i3PrOl5fnViDnw5bjSnd+Tv6
9dECa3mgbpIyfy7t9ORbMMjT4mUN9BYaeWx2nHtAurtfi4evnByfXrVR9FAQIz2GX5z/sZ5Oqffq
S06v1x+YdPpLe5vK/XRLMCgANuaEHhmYaVxMJ0ylc4d+SQYg946xj0qkk24KsfmHLH+9ewx4YAGW
CA87aexV7VdOcrH16Kn/M0M2wM6MyKMhFcxi+Bd61vH5o+8D4h59PGGHE++oAp0WN5uRZwGrBzd5
5QWK1V5qMoqthBhMHJpPq0aLHZ0cXVwVTOLUkhrmymPWI5uByoQrJfiisaLIdTa+yYU+941K+E85
MpzMuH9keziHx6N3bXAsXC1e6kLa/RPOrI9oPGQcpU16QwznJGL4WbKqktHqgJUyCGZ1ynHwHNKj
sVfmoQz2rSp4/CxHRZkh2TEPD6uMDdklLggpW2E5Yvnm67qJyLwQWlmrdb4wKISmisX7/+Zcgq70
9vz9PYonGIlYdWiMPsyrTdeYJVNimHXOv8eR6l2wtGeM0Rmhx3+smGonSCmvv4vTCrPP47jNzKBV
CDJBfmuwJxmDciA2dmz11akoIb+2tF32hHHHx9x7y/TixyRskrjfBF/Ke/6N91zttlvxAaoHsbgJ
8/AERK8yk5h4aqQHmJUI1oQfoCGtbCHfNDFth6j90kQUB/kDMTcQB7M9eSCJknL2WgxbV787w50x
cagcDR4fHNR+CtU2Zx54rbEZzG3pCzJsf66YCFl1m37h6hgeJHTjVr6u/QrlhdhTQe3Q2hUZQQyK
r0HZbrB9mDC8wEMlECFTPwxuQcFoz/s4Bw+afNQZBx7HYtRSK7a8ZfNDLKYWtBXp9bkMdxRXKYrS
fiMUTmuZkLVEtxh0m0NL+uOZEx6jzFh5dtYhfkA2iDB2wm8z9TlCph9+4ChuFbnLuiTQzrgmXEO1
1B3aXVjvNbSKAMgOMseJwlOqaCscdsz5NFM7vspj5VzZ6coRyr3o3n1remEYsuSOpFhH5NZmjpou
StpIXywkKmHDEiEdY6yWQgxT93QYNWx3dchdhTzvSw//QXRPwqvXRWF2t2lnXxYvKEe9tfzri59z
T864ijF+K8ifvG++IIimjploVt5kU/N0FZYxxlqv5y2kmyYR/4Vhp8frYZyUmBEpsmxQ5OR56+Uq
BDu0oAuALFxtnb0tOepcrS1fJTaJZATjTeJl4SEWGLXQjO+NqSK/mOzBN79+t9GtxpJUgR5KGGEH
xmGWOatQD52BrtTfLtuX9PwXVX92N5Y1GPXyumCTi9hEYfaAHsCxqPOOd/07jzCA7WEEnnXk1cXy
6CyClrHnu6fK7W6NYm8d0IpAwmpUvVQSoCA2oucG94bvVY2VSkfk9cZeeWojZBC0tH0PRgKz4YmN
o71HQyE/eJViePLo/Wc+Qd/fUKoago/tFvAmLZ+WyhS4VnHaHVF3++aH8lqlbQwNvG93g0rE6tbx
jOq7Xgi+AmURMRpIr7oMz4ao5GGSZUS0auAapKvfDzZtM8AeOCDBVyH88nwbMe5YUGaUMKVaUgue
1SBd9S2t19Lh1F7sEJxmer0X5IGJ9REL0Q17m0rcVm6iKw4F3SQ5OgLbprTAkvpUnumKL4W9kjct
30mkh911UejJSOikETjKm/FqoGP6qwnkvBlwfpoQRFTohhCm9YGOG8gu5cGeW5bN2Mfe5GdLLCHx
tndK8eXME8GAAKeHA/6OJTWXpGO1pmfhTYJKCAhIQ0SauO9H+5w3/e8Xx+yIelC4jDli5Xbu5iM6
jqIuSLIGfapM2Uy49+ohzITxu75kI/LZuSFuT2FjZES2C7Krk/KnVjjlzhZTFA3/bCl5gRcw7GO6
yxLGqdWgUWFFp3Sx3HmEhPXRP+T3wlIdPSgVSKBMnBqCnPToQBCiPqQ58bgeOYgJrdT1Kta/Q4Hn
rbfAajOe2pUDNWORk9cSeddAfKTU2iMRUxqCu/eNGVBFdE6UYlDxbW7KWHlGoyGyRvx3/E8IWWxg
nsobtF12JDdE66IY9xy4NzeqF5dC3+WcJXeq7/Br4feniy4BnFiboZElZcD2eoDGjCAfXmOGAqpe
53ADhI747fyL2KiUXBjAcakOe2JMrp0NzckCROa8UPXU7opoEVhGy3Mwa1ZSfDpJ1RregKio0l4P
WPZhSR8wztKfvE6ly83UlV5ZatmiiL2Jy/apAxmbXmMfDCJaJOnbhQ18UF5EGYmYDK9y4pnoUMGX
OFMZlotI0KYHw5KTnEAuY1MWJ7d1ab2SoX63gcfW5YRHJFzBdXRC0LWXM7kUPLxG351S91yrCO7t
RL891yHHq5ep4F+qAt1yMtiJ6+RJ1+UZmMQohxuuiTeuIJHNGEGKczNy4iobnUsU2fYHBTc1Dw1y
P4Yh0q0oigx85H3FOR3kKDxvaC/Ciyxb+pHL67uZ9f8WLWpoVwYfUPSUPW3voIwJNQUlRxHmQ784
rynd3GN6R16I9Gwfb1I8ApqeJxkDRqcRa6DgQ2muJPfSjsLEyUUqCdEDWqvF2YxNC4u8NNqRTlRR
AF0tB19oEUsCfn9Ucz8Lan/LLXb2+24d4JMpg5gCJAM884ImDHXzBvK/9ZHGmkhkfA0snHDwO8du
D0FcyM4WxGTeM0ccJjVT0gxZPLKoC+xRmeRgY3AzoaSTKuzsl+KVRy3p5BNBUXfPYioVhtBr+o9m
ulbdyoIXFIpKnfmDvD9A29p4sned8auTs75h5blK71TcjBj2NoKeaUU7WI8+zo382BYAtusPUOY6
Q3F/W5eXEskZUo/l973O3UigjD5v5L69QFxdi2U5q+zI2NPhO9NauGlS5OQMyuFdOCuc8KcvFXki
7f97uGi6+5gcAICGwtgQCP4dc7EsiGNtbdabF+zYLeQmfC4QXm8Hbx777dMv8LbUjNyN9/M8euVB
ftLYoG942lHXP2VWp9ycU2klngTXejaK7hA/Jn2WqKxlPBXpJPO8Oy7+MbsqliKkWC/IZlGUhLeM
BdTpyaOUaDwkOt2mLNRH8u3Fm3Y2L+eWt9JrbNpQcmTGkBa/XsGaMx8KAC5J+zmhHPdhk3iAnJ8Z
idXb8dCPYZuD/Itkqpd2nZgLvuN8pze08QHY6wNkI7dRvm/3WO7g2FAqOCiKHbeJEUrASaHAkjq+
j2RigqiFkD6XA6RrIc+c6OBCxZMepwZrsMdxk5XwdXlLTq42vetGFUunMEaN6rBC2I8wgsRSxPtQ
sZYn76eHTswsDHN72FCtl866VwZgbh+Pbzooy8FF5G+RKGs/qZCceBdDk0NP7mMQc2r063RIJoKg
Yqdf1PiH/JehNdOs6k/KpM0iN5c3H5a9Muisk4w4sXKGomtAj7I/TrUi3iBByczvyYbej+TNxF6I
KEc4B6W9RUwrunmIUUXCiuEwLfis5O4LzmwSYVAyrKrNsIU3snZMc/QDn62lXMRLUJIwuNfwOtPb
KIiq7k+4AvuSMyelQSRWa5yo04wtXN0T+y+oO2qAj+nnxYCnccjn4MbqN3KdAfSQP7WO+Q4RnIKp
0lUzrDp7V+2gc0TP7pDHbSP3JUYqODhjojKbzsizoIrK4hbMabglZ/Q7fg76JuBXQtmdpwYpAts6
uB0d5P1bKf/Phoet4TLEHCmJmFzeyfla0UVDSaxRyQJ/onRLGFYZ9hSrk2Xvg5zbrmh3+SG3S4vO
MDnBBmd3j+tJ/eBaX/E68pNJgtYyFwVri3I3Ojx/S9XxJKTmYIZ+gHOzCOa82e08OetA7kIz8bFe
hd22Cwigs1G3FjSjNqsTp1qEYhWPhNwm1jSJRjbcroDb3MbGVV4HmSFP6hjI2y0brV7FbQDbysdN
pqxFGSIKZpzXZU2IIzwDOpYn/4s7V2n2TfywHNoL9M1UKHewMMHiq9A7wQa47R5McSXQmyuugeSR
kpCMpurTIEXtRWQJv+haF0SJ7rz2qs957HO6D/Sr/JbdxxX31XnKutmLCQfn+YB1lqHqFsy9BoQa
QQLeE63a88BIfkIOVujennkD0qx1i+6ENmZ2PmPn+YRxyocOInjRN8MKE8XkTcizqI45Z3joNut0
hKxt2EpEjQayIjgGgs7RsRGzcmQM5FibG5nMAEY+lHnEFylK2nLJMtHWa4AxHGw9x+vLlGCwzk8v
cIVYIfvzCsvgiea0HEwfT5kmrlat5CwalxfDJG8CDdG/38BTOV9hkBzQjA0hIj/Y14lj7Nzc/46b
UfOyni1pzP1RHQ8Zcsm/cIZtxQTsSGjTGhbRecmwsq3nRs3PPLxn0jyiE86lM1W126rw2WZcIDD3
3MU/C4HtyGbzzYw95qsFr2+velubOgRh3Ek/nyhQBc0rrvYVpH0GGMZDWlC/49eOZanheYd3tgsO
chKpyqauC0zoZfpLpkbbRi2nH3hgqoSdgZeKVducYYSxjaRxTivzfxd63IsjiQapzug5c4M5LZrL
1dg+WdQiy/QN3TJsTy8Bj7ckhyiErC0L3tn+1PG5VUN6zyMtP1trQvIHyRcUqPZeVoMsFYXY/9hl
Sbab8gnXOm24tZ+y3D3I46lRF9gPRBPOBGRymQ7W78mjT6MW4+Gb69YPmk204CiNBulwJVedJJwG
oFzCP+mHQIl+wmtuQueUf0lh2+YXJ0/kagiomBCAVeh34qG6G1l+0H3yl5YnM8rqDaIKslC6ZRId
g9ASTiE9Rn3giu6UgbtkHZ6YH6FRAY0FLUHQnkkHVVwtq4NwAIsJ3Oqn8rNwpG0LqkxnYj27u33W
Dy+QblapZ0B+hhFRZnBXfwJR238TthK2Bz/bitsHlhxDS8L9n17X6A71VpNzH1W6A7vdbDhCIKeD
vo6213tWE4PleqMCGTX488retOiqOmA+ttaUSrntoHP0taV9y2NLCxTW1r7DQxHGFQNW3Fs2Wna9
xUGdb03qxtCylgR1OE5kk+K/mz6jB76CqLen5UUIikGzlysd7Q+fY5FjVDjUmjzQ6NPIge4z6T1l
2nx/ZIOK22lQrKhsvM44jVtMVFrc2rG+fLTeeyTW6iXZb0/e7w1/rp1UowcsfCIIzvGEw9r1ZN6J
ztZLMcIJBgJ2arBAl8yM9D9QDizXbQa5Yi67MhcpUmuS0MokEW8M1WQG+NZr1SCBbuCHVVTNCX8Y
r+WGznCvOIHrZxlLUFGVVUGm6hTPzT9wWpCj9ncv05znW2FcN1OUWxVTXwwhi5S4ZhSToHIDs6LW
M7AkbnKJxpylICWjNY4f70/AYvbcCYD7DWTD9GH2LJbpc60rgEQ1sVfDH9oKbfltv7NGpKjoOemy
Dsuwcw3gUeWGaFBIhhWbnEgOMUHqJ16hspbUc7mtUmkJVpTBoaTvRB8QO39+72Uy0aj53CrDfg1L
z4XE5IuKHbDvinOrvoZQE/KV89G9tHkyfI+tisXoX4cLzupNaqbq0Susuj9sTG8ORTxP1Rzd5BAR
oaCDp9BH22Jk8xdQvuIEWmPpzdoEWWrmMiswXMCAxmB9IQtZA2r01QVz2qtrXeJo2Fc6JIpviBZI
8scwtU+OT9Y++zaxW6sSjJHzVWojoFAgcKZVuNK6s93FAe6IW/BRAOZZNu0iwyXGKD5bck7+xFmT
1gtVMrA5nagL8Yf7h5P31QPjaXEmRmmZpR4i/qrCp7rXZQYPfbcF2JXUqUVyCsSHG/4BAZ3dN9E1
dvW8H3EohcjcddnyGhFmK3GbZdpbWaxtO1Hq73i6uW10h8w5OYd1G007BLMVBn/s0jgNM8kpZtSx
bqshQb4Taa8kMQRyarjcMQMH5XAMmrm8NhvH+g+7Aqr9PKsMKboY9aPNU1UGQ3jaS8D61APT5O5z
gQmSbWkBXka1pB2aiw/XGeGsy3Rbj21TUcTINjpLKs17AcHXKbWDYI4JzAXccw1gyvWTbKbD7dVa
nj3aA7By6bwh9T+fR4swJOXF1JY/csTKkTejZxI9z/xTVRkEnZkavjGz/6p/jfC1Z9hrPfNMZdjR
hcTBfEYGb6yLZy0mLhfT3oYEkefIUBCMnXZksftK3mV57qnrwSwN2lT8b4WD1Il4ryacaEDItYsh
pGYV1ue4AU0z4gAFb7j5oA2WaB7cL36S5KrHjrLiYIFfmiJ083+osIHoFuvsl26n3cv77XWe4vmb
pkl7rJruU1oqiL8wrBTLV+yiSjLKT/Hrk5tfx/NzgwSPW/BZ/Lwv1ywnUGiAkL53L82oWJo6TCEy
G1xnlS23N734uOWi4SfL8MMRu4gNvKns4FHoYYtDPH6sGH1+HU6bD7jiUO/NGQx4pW5KVH4CwnuJ
xXmZWV7pi33OVPeKfbPdmV89+L850oLsN/IaAJmzwS5rswaAfmHhLCx1DvUqZY+UdCxQqY3KsxR/
OnXgF4T9XhqWGcCNzB1Mzv26YQHfTj3YiUKBwN49bGV9k0QFdluQCnaApYCtUXa8J57h6MrwZ/7D
GDGd4LOFiDi10jdsGgf9DVN3nWpqi4SAuRrpfze09X27uj0i9dygSGE1FAIO38hnmc4ATAElFSMG
rDzsGIUQptF3BxmabPxWeKhllECQ/PCFajZLKiLm7GhM2ulKh/qAKKo+JZ9fRhZCV8tGvHzUPXLn
/ijd9yCq8SinLi+tH6Av7s7FBF6Bw4BqXEtbuGcs1Iesok3CNoi9rQP3stoEYjd0PNDFOBpgP8l1
ZBALIxI284E7M5Zce/AO9WVbv/Cq594tRCBirHX5jsAZGowTSE9ejJcmDaio8GVBV4dPEkOk6Uo3
ZGMNkTqhVPF4OehNoACdC7QgY4IsmP1ksLjD6/P+AsgMmD4GRIBppG893s31sXYcrH48NKzNe2Hh
Am6dmepN0xCVtKqvOH1umLj9KAdSlNOe7xgKaReh89MguaxasZeUh+N09AULv5gqJKZDekAcXZ7w
nPR/RSCQBbOU5Oog+BcrUPhL4y+C0SmvLjjijn9STsWja7SdQzkxkA+YVsaT6STKPMbc9ZT2UfAR
nAyuZoaGO7P98s6lgsncvVauZSnt4NBbAnHqNRuCWxYZ2FDlRLxgK2rCxBVlxbruKy8dDNQpKpbK
es/Qp6tv2EV8ExNuEu4j8900fmHB/6alinpMlwp4+rUJuxDthXCDRA68G1QeMH5eHo2yF68vwXha
Z+86oYAdZtoCRORejv0ICyVJHDCiniUmVQ/Mmv4g7ZwEtrwPZMsEA1a1wqvcR7e9jEVNm3uM2B68
OyjTy6EeCOv7C/3tnrobVZd7PgIkVssPlU2zji3KwX4J+X/qX6/0LkFEytAX9sZxMBgB/Vs4l769
M1FNicsf+g6ljxIColmB/gZQebFdpOaxgSG5/tigNwcH68+171VrnIkdLg31SCEVz+bWVtq5FaVb
2ptQuiWDym51qZSeDPQINs7Pzx6MWNYQBdAWRlNC/uZxYsK41ceMP2QHEKpZV2fI8HlFcCrQ952I
ikGL9UqxV/g9XgssmsliaSuU3a6KWi/tUOFEqY7H8ELIn/v07t1ehLMQr/wT/1YqDaIDEOIThbU9
+fd2UP1WjW7hY88Fn32NlFt70PXq7MbGy5pcOAm3XcyL0EFCYJ2Jj9klvGd6w/Oq4+Zou7ZBRb1G
04Od82MDogJ+GqT2WVslYW239Oz4YP0NnTbGMNOmu5jDdkN10EVFdrUqIGZ02vpUCVLWjlpMGqbP
p7zQa4OraHKSsj1FqGM1GeMHgLdR4uXP0nQTWb1wK211AJudi6J8YStnqh12gnCloHvdjsQnMxBb
LaWD4r++cWpUSdiWKw+7jnRLra9Tc5jNeWC9mFL4GreyKP8ifLi8Q8oCkeWBSDb5q4R5LKoLx4Vd
sxDVD30YPfBP5dtnXZPZhpvEEN8UEmeKKiEK7NiNBIrpsJ/6jcfLGl4YHZ4MaxDlvhvoKE7w9SrQ
HLEjyi5SEf7RJkHSSQyqgH8zjwGg8nzGRY7U7FfMGlb6rA7Z0Vi5aa85eiO4wOOKditQH2oAUZoc
RLYZTz1IC26jhV51QgaJgNdQSxYWz7ustQRxjuxt0M+EOIAU61Ej3Tj/oM4JkPXQxfs/JsrlFzao
c946vyF+DZoJgHK2m+jj9FB3GKNYiqvkBI3s+VxpSnKSBNn+KJ8bBY4FRYubVc1m6620oXEuUy6a
Fr6CjBaFZnLjnQ2GtVr84Z6ls/W5cZclWXK+s+nWb16vRDT6VnWNzvMr4eDw2JDUHkiICVfVbkP5
fmq4j/GvSG6AjInys4mx42pd+d5oHLe204fe2mKbKQ5qV7mEcky2kqpZmi5EO5owUs/raUO+pY+5
hFDgrk3Jc/eICdcpo9+XyucFhFeYXdP/QQEBqDrOdwe5IiICWmL9OEgyPiRqEft1iUVoMX10lwAB
aLfJNu4x4ahiLjHmoCvruOJZRnDksr2mDKPU+QS056z+zyu/oJdib+6pHAImxrAQKmGzJXA4fTGw
6P/0QNKv7rQ6gBNn8DxnPP1Ky2L03XD9tPuj7C2B9lI8NuiyV/iTzA5DC87Z6CmBLTVAXMOqNS97
GHYaogQMAbZkMDzR0O0Z5/iMNWjFsju6hieUoPGgItYwK89J15Ls16EU0a9mH8XfIMwRRMn1GUxv
yg9h5ve9eogEkGbjoWP9TRWcQbL0YNEzhWqGDqk63IjuYttCIujTe4+Uc88vN9tVJik3VzdmwbKF
s853MbzpvP/s+43tnLYurpWOj1cxEGP9kRsS+W80VRB0QBDDaEHIUB26SUVbzJh8AKbZSe7p6f+8
yaEWPGL+RdY2oVRM1mDUJ+PkL9Jw203ZkT8BGirksS/m/Ho2irXH2S3+XPMy8SkIBYkpreiE3wOo
bUmAjMfnvPyPpfh4SKI4njuHbOBz69SF7KEOnbbu/e2dW1/RIfn3gEyA1IP5P2k/mpT3fN+zc3dh
+7wYYoCcld4fye1cHyoKnkTgjyVAMAlv4vl/bUrSEdAnBzF8ZFNFPX3FuCVw6TjX9TwmTAYXBLbe
dgcDhYLm0qGORlAc9pL9LZykkjfDiY5WznTCdJkrPT3IWixosoy2ZIntGsUghEclakeunkFBDUZE
YU1v6cskYR7NWcLZKOVM8XquXsqlUi2wdbC1rdNB4tw2RB4C+qYSmwr05P36RgYX8OAbW57HnOzA
bOhEXgYWG4nd4rDNgjSCIlt+LRV+/AuO4yG163JtQHHBPBavuM06P/jPESn4XOH6Gb/i0yxCW5ZL
9zu25AALFQQLuWB0PAC+pvZvrUPsMZbFO/TJ/1Wl31zjxvfJkMA4Jk1wiAQJ2BAv1S+SSDR9rAB+
ozUFNe69+EFYOrRrGrPZsFKp8d5NmSq9DQPv1LTc0jnVo8eRll8ne1ThhbzgcbG6EXzTAzlGyjDZ
FLzp+et6ND3QNIreggtU8JBeqLLBjhOn+SJ61bky40RzG+kyPe231bqq7h7lasAFgxT5BQgesL0J
zR4JLW6tpZL5x/v8meFrApk+RFnd+70XZPCKGlNbtgSeXMS14KHreMIcqVLs4RUenAvAULqCgAus
9XWWqoRe8pmVEwYTnwNnEUTRzvF7elWDfgcWFvCXjLFedoB51zVca5aAKBOf9RztRU0ubYRXVoJz
9hGmR6DulMwkT8Nkc8+8q5Z12QkRZu1Iu5OwtfnUOxjHc2Bty0JxZuvBr/tNaXZJnrD/l+JrijEe
KyED6CBGQtONH/aqNmQvv4zvNXsWN4oJKXGrQQNxHwpqUimcj7TLk0ds4Wznx5kFKO1gtX3aKP5o
16cGhg0Fzg23AfAfq9dt4KNo3WcABHU1Irj0wJLdAfUVLiKUEv+fp/VOYgY32a4qDiBa5mAOiqPk
WqfD/5McR8WoACOMgd8OZvnKPNGRneKRwROybD4XgCN3ZF8p/qXYnyqHAw8+Hw2JpnR9n/iZ9C5F
DqQ0XNshk2oW6rU08i7VGs5KjNTYz7pXEM55aJWrubpwKa4l8+9iB1uPKkPnN80cVnd5TE/rePEb
u0DQl5Y8su/9baiOugqnkovAuBfMvbrlX+QDA8S9+f8nPQT7KooR0S8Sb+oMfvGuluQ9NGEPzqe+
19Saxn2VG6DbgjAUxZ0ShL5aZOBHcZhwMuBra2h04pIQNIvS91iYa/mg+Q2idNPY9jJO3dINN321
81+n9QbaNiI/vb+d4DMXC1nWA6R8BdxdM8fm2PoYaTKzbSYEgRd2Rnv6TgjaUiL3cxLhqMTNws9I
XUPCjx7/5PPqBp0pIts9AMvKLKoHuko+WcszzmXbQT3uD5vjRPWKP8QLAOVgpTQSKtUCC/YCuzY4
SAYXKK6cPeYkve17kdCwVfsVfD4WTQYl1xf1efK4L+pMqOqxdGWxXlrhP4+S22wNYU61aKE3Q18p
etXigZfbyzBOdHTFEHbEVrMZKVsNiwiqLg+a1CGgWviTU0vc5H8xJWKe9DCDNjoWinEezp0NR74+
gdUP0gHzULo/OagXrzck04NtjWp+ZhqzFB7hC797eAHR+UIho/R9HyE8tvtSDOwAzcJwBGr9igLL
VpHgVmirrRtiaaLuhJF8Pz+uG1+p0amCqv7Z4+2KdEBEu0Q+8pyHzAKJY8JgnKo0w2xdOn4+oQyp
m4m9lP5MM6YmwrrMBcXdtH9sWPpQM8vSsWvH4FhTYwFRJ8VTmkLGTJiXM3+BmutZ93Ogj3oUBoT7
zlnYYPV2YSvk3ji46tfAPAvKErV0VFVmg1/LOLgd5UHBteA8Kr6Aw0G75IjH1pvbz3Mr/ZXGuAci
733h546ZMmhuccCjY3qSqAW2dx90lmWNviDbQ1jwgC/jadAKUCd9W4gz3dZ81/0U9t2l3kk9kFfe
03UcEmz6bGTyouwO5X7Oi+dJzk8O6LZFxyvaD/+kSPb11I0eN3ExbFlWuwCCriCnXEYWw/XDE5uo
igmZW9IBoMgfBvjs2VBaDi/7aizr5EhfE6ct6P6WRPoJAFjBMJ3Czt0f7j6002AcZCleqoynMVgu
xWZ3JpScgBui5ZFacuWctWzt4tP3RQN4MBMnHbHL68sxOEPRIJ4zuQ9QHqoFSdDZoAFlVhCpR9Ef
8dlvLfxnd9mbqj2fEKzS78hWs8CiyKKOhpraGHGyOZL9kRyy2z1H8+9fwUuu68ZJhDaxhMEcXw2w
AoSEPrHXX/JyHLbAxZ5KH2gJW2YklhGQnFrgrC/ZEE+R/0q5ExI6BRs/9eLdhkcnbPW0w6D2ZX38
OIcidymfwTnbWMN/upB6HXM30fLt/XtZlyRGpid/IgCfc2N3nNTAh5toW0mJqzYy8aRh6MnlLkIZ
AptNoa6FC+z/YgL7B+fkufQQRD8c5OGte9imD6mF4WzYbLtFHe0N5k5yPsPQT6Q9jhFPeFmw/A8s
VkWXxkWnXpyY3RBKHgNki2iANSIPbz1rx55N5NoliQiUwFVdQd5OvL+tLBhQU/BU8v2glWM6OkkZ
bKbiFnRDYCJzPcnWgWvFP1D564s/7IopDzqwTTDEolUKDi92vpO9sMfqdYhgqutu8pYEFZJH5EFZ
NrEiJ7uIKg0iNsGcQ2DTpCiviI6Vidk6QgkKuL4J1e3tQYQ9K6g17FaYIzgVUsYhKv0zn9qlFNZy
PA0UGecR2m9+0l+FtFkjhvxkbEeoKL2BgevqOqZFc9p0DHhmux8g1qrPm7jd48av/LJm2YeHO3su
HhDI0uIWV08RGIF2kghOaR2cU4pqDfumgq8Uc/oT35cfIhmKcHZ56cNnS9tEmOdXeFAVBCPf0KqX
bvCHUWWjOO02bJZx1buK+8RUdlSa0amOOhC1Ld9VmVJJ9XasTWerWSk1sWGtv01c1uB26NBRqlv/
H+WHNg47+w7HZLq1tDhKYSx4CQWgrYrrgsEQd+3Cum2H+KGoF0PHFzq83auJFLj6C5YL4MXFhEw0
g2Bl7yLTIiGygYzdwKdcAcnJhqa8/E9hhyp7NiXxVGchLSsmBnW0MhIxlD1XuCAy8/lojlZjEzB6
fG8g8F0Zp08EG9ODBQn3LA1WQuSPjzqGDswHsXU988FSXOJnm1EzWn70/o/+kCtOSGEE2DYT9VuU
m1Y2neTN+Mok9kYAeCZCZGgpUTRYzurTHvsp+pMiiiuBJgAiU8TtmdtXYW3aFLVlBgu9d6Og4p60
C6qm4s24hAOSZCdzug65D04SNZavHXQUSpI4MmQnE8Fjpupi1UDaX7599lPPllgasoKwI/bVKa5n
w6dDaUzV6zrHykX0S24jM/TmDDl48cR3Sn+dYfVVWnPqj0aYKm6wV8J4RG3NiClWoUfLwc/oWcoX
XPQ9RLICTncrnmVJZORjLb2lQw9rGvwa/jWYPu68w2ZS9XUhmyGkrTYdf/2UURyNkESiZtmihRvZ
wmfABBAHxBRuGS/i7YQ780q93UYimhzMpzcSaX8BiikFimaQPXS33G+J4ic5fT/rjitd1PMnkwf5
yAw/rLVMb/Dg5f+X9YveVTy/Vt4pQmGOsCmcYK5g5hL3M5ffJIeySQ3fJeKWpbeHZ6rIS+1qzGbY
yNSXtLvlQXfcdf1iEG5lzmVzzn2z7tetLK6NuMLqG7Ngl/V+GT3JqlLempEHMoSaVj9B/SZrNK6j
u/ypufhyj4LvMX4M2e5Lyru0hrm41H9pgW2uIPrcOS9v8uouJjIO+H7sxO62y3u3maVJ2AzjQRMG
yIgNpxPMLojy02rqlkn55IQnEiBqHQJS0MLBvFlfAT+mT3oDBvBy/SGZeGnRy7b7VDd/pY00r4ll
rRXxwdNXMGT2uU+ss8IhmW9bkbz8nHKznWpbl4nZNdFKJMkp9HOQm30nwMihYfIXr4DCViUmtFtD
QfSuimHTeziZ3/nQQSbhSjd6hYoEjqazfPBQNqcMxDV7/rDLMi0+4/ehVclImzvAhloiYiXR6DYR
8LRNqlYaBIL6Z6PF/0cNUfQsdKQfLlB615ZdpA5nfnHtG85S/Ze0w/8XJO8USNNVen/VugPMI7KV
bcyBkzZv0ZX/3MZQPYJN8syMIMF9cGladHfAYmhf5V79ObnNJNl+XXaPlf08ns3Ah1E6BqSXxXUt
BMSWFdyuqcHqWVedV2CfRROoi3pcHQ3KnAl2AqYIe1iU3DYDVhrGhNfd6nrUTgoxA530A2/WwphO
bgXBRsvh8xTEUoIAr2RJHHt+4yUGpXUl00M6J/495s6RglC1lPRPNgwm8x1vUe4tvqOrMvbYu5eb
ALX4SwSBCYnvDTfIPl4ciKZcYzafEt7E+n3CmODeO+XCHNK3HJP050Sfbl6iaubESzmOA96xdHZ0
oAu4u0tx9Uvf4qaUdazpi+F/aMuhL1j3Y8YHg1nrPifK6dYTu/GgI8ASwQZ4pdQwW7nAo9aggr1/
6hb9rfSjtc4wD93YLdmamfo6sCxybCnKJOoZvuvAUGmqetjxSYcSqKDFHxnM6PiinXf3Jy0R1IRr
PzHPMriMZ1EMpBjbJk3h1Rmg0vaSjBA2zkQ/6A3jz5JKB5KDP3EPqbkCms22oh4Uf3FUUQl0Htvv
/NsTTE8FwWSwFnAwmggmidwzGvXERI8HhZyD/CZ+HABwdPOS7GmpLcgEeJg3Nl7ofEOYUHAnPbKW
F67xAuUNHzututeOQ14oMI7mZiSfx0nJDXlb2NJfrs107K30Mp0yMXA8Uk8O72rJjdDwBuVkB6W8
PEk2QC/nJkUru9pJQRK+pKlCp8sCyQm4Ztm17Dw9utK4i9S0o+ZWDmOyKLiFcQwfGO1VCWIWa/Wn
+EyFDJ39iHtiIMmVleMyeVXRXMJE8IP54DwZPSwOOhMlRTPSRBrCqbDy2IhmQBPpsAa3t43ZId00
EQQ9AmMrhxlbFSdOC/ieYmeUuuzwzNQf9ehF7xOceMDEYjANM/KyiY5MzZAoeJIqWpuJRWlNLGgo
bKbTI9NEd8r9JtNwDZTBOecrkzyeiSe3rosuHfFyLdY0VqOKICyeuTl6413/EG1uPXVlcJfo8TDq
eBgKVZLg2RftubeRWmkXETZC2HkLvGpZ8OrrWZbrsuumWEyMvl6DuH6smS85jZVWx7kgVMLLrjs0
1N4M7IdqtPCtEtbUkpLkubwP4X69kvQ6lLS2qbm9ww1+Uel0KGIn9D3Giy+I+SmSxmLRrXXlZyVC
BfOmsYBwqN8Gn/RGV1+64jqYCZMb5DHU32o9C4fxkleFBuvzVP0w9rJJIQuJbwZt5P7d9vJEXgs9
EAJcvzeE4YVzNO6mWXwsg4o5lqCjhqGXJ9jwWOZi/1TpZM/EbJg2ZKBKQrsB4XQOfQGDhcQ4ewL3
lwm64Q+TSJfOlaU3zRaIlrcXuUAOlS7363DNa/yQn4Y926AxpW4bq8+CgWRQyxff+CKxD30oLO6V
JHVEFZWLhMOxxsYRNH2to0OZqv8ZWHFwShPsR0oQMj/LkM3XtSCv7c1ZVcyeiH9T4WNFE0Nww3BX
JTnNNXMKSNOZxMg7OGDBHxmYdvjWI2n/sg8VNdgwq3wIanFsUpnjpXN7QnHLkxJ/fmMoGFE3JRbb
B67IbgZZ2dh7K/TRnjqGBH52puh2ehgOsVVu52bIzIcxOtjRnRprK6T8WNTjkSdlXvkVXKqFG7LX
+Tb16MZzu6Y3eg4HimO9SK4BxKHL8/53IsvbY7TAUZsW6au70Mmy7E3iogmXFhkNBPLTHgEVLDPM
MURUxuw18OmQGgabcSaUluh9MBR3HLa1pLFnNS2k9ppY66NcPbDe4mc5bPFSaYA2pM8AmBDk+YVK
DA05Xi1uuwvGrB1D3AT3W9wJ6Z8Kfu93Sf/iD6vu69oNETkcA4Dghr3jRB9ChmQ4q1A5YDL7C02c
TXuK6r6eyQA0sw8wLbJiAp0hOx53C5w3dEA68g7yNCBJYt2OUUcyjGYO+3F0+H1t0r5nN17XUqPN
NROASD8Xv5XyRbacwRurrJ4qrEIIC/+jaxjhy80i9BMJE9Xx32hncQoPMnHJA58zBZRmpJF2XJ8f
oGWMUeQ9zcahqAxmnBvyh4dEyTmLqUYtTyqx5LTDm5MohcpX9CvLWY/02yedBlLSuNmvurD61kml
QjstztgSuSisUdNdMIDUgHQRTpYPzie/t3lvXD+BFgzl9U8Tur9btaf9Fi6NbgKI4XrWoHntaOeG
rUN7XhziXCBLkAMZJMHcTBc3wetYAKDgE4qmlifCLrC3yioR1SKDijFgvkT1jzbbiORLfR35acHc
mwNfBsK1uO3NDMsoUdzdrgL5zXDYVveR+nxG4rrqd+LEgENnWOU8x7sLChUxb8ohqgaBQVZK1ANG
l98NBVGRBck4VYl8l1DWCCVt7wwMbt17kylxZVtMrvU40MiuZbljwEJJVMKRZk5CLQnoqA9EHFJS
620SJOPsQiw/JhUl/LI+inORu3zLygt3Jgt33+L3xpD1hZKAl8yKcExYM7lx8Y04VmxaxMd5mct2
XaFZv6L6KecavNK1DE+RL15iMJ1qx5KrgFQHYAfjLcmOXZ8b/aE49unHJMH0J01MY0xfkdSQyy9n
R/xsmgs8G1GQ1BOTVYljNaYA3zJ+cKSbn+ri4UQKTNnL0ciwyZOZJf8XWf2GUdcvjTCyrg1+HvBX
8QqpnAUtyaOp8O7jAskD/warI1zVR7/XK/n4np6drLCuLmYJRzKWAHcZc/xbQbXUgRfXBZJ3r+yk
WGDxISw37ovcG9X+MnoCYoe9RryS8xxOKXM3Ju056IRCirYKvJnNNkGCWYZkpDhlWLo6bcqf1XmR
TydrZZbpnxlWP/uEnrTu6HdcG8aRwDzjkROcmjlDoL6wEMIMX7ZEfkF0cidYaD+4PZd0cP6fciDn
ZObWZTeA3BWnKPM+fIlx687bvIUpxt8qUl0dGajVi+A6y8XO7p+6SdHW3ZF+f246JJMMkpUrbCg0
5+OzqRVc5kxvFS+rILPWyXDfj/Pvmga+O4TWcIYY25JwyxzmVei/WEn7HokFNltfuWzKokzeEcfR
11DLe84+norIll0yTK6c5LClWC1fj4MgLh2QDdNLS3I/jp8XTEYeXamQhXkmVFhnuqCy7ocIxsOE
fnP/rcq3kiFjThSV1nn7zBy75n8Ip6KEFlVOl90Ee7ntdpymMQXFBI3esFMbgHPd0NmvxVkTAW5f
cpKIT9bbOvS1JUwBc3jhtr2qarKOQnNKfRThaZ/9u4nrIiNYcJ0fXXEnSHpqJDc9Qv2o1fkDwHs/
EXJqo9ODXW0gv7pzQwUjLbs9A9c+FYoLQ/N1lHzs1evBzfGUBuEyqC/6HxWulFJ2fqby7Iv7ah8M
vJNdh8NalLbEDMt4CosgBaOdAE2V8wvy1VMQDO2xgWDXx8rPwZRXHaTunIDzzAEq/9UXbnK65s9b
qpjwaOKO+tLbHvQd54HQD88PMEimCztWUGQeamkfhEssaaiE2koJkEyR+ww7gX2qbSWPWOFk1xYG
uaGvNyDoZZP4Z244wcgJYQi5AOZHwy8V+vYoXoekk6FIMehbHCoTgS0ZsXRh5c6NtbW8lY9BT3XJ
0P1l3UsPIx6pzrBucQvc+Yn1Cx9/9vfjUJGs9Oj0KJUCGr7azbKO0I6pfLtLA4EwUchhds24RoyX
23mDMdBxBptdj/Mnn0dRlaLZGlXsurs1zm9MAq+wp/qCB/o0c9Mt5ATmG2lELezLELBv4hkMqIVL
Tb1AjM8y2QOFOQ4CQoS866kXqfccI3tctncl4WGIwFFPrLqWeTi9TyIcxrSU/exVUw1Eul9Wa8kS
IAmSqPJt1fIsoPK+qR5xpG/iKzUkMNMXw3wuYCKW4WqaDTG/84JwVs3e1UrCSSV1pmSRmXhFeXhx
RIGA9aBlQkQKKtX0nKKr4yO09BnsaXwd4MLZWAbWAtfq2qHxPDpNe0QXauaYSyQB3yap55Pgwkhe
m04ExJyjESr7G6Xk++T9vprHFLlHYNNnTItWurqB6Rvd9cF52J+wdwTyk2XvUWZDWlef16idBpoD
lY8+YBYUEMBcQuJi55HWgHi3HlW63KRjG903oufXmsyFZVOjGI6zxrWw5WEVoFHYDugAhUNSoSMb
drSqLkEjHyky0n1kYwvDhhAmrchSMPZzzX+fooPnhIgYjlGDvEiTQM9ixCPjiI9sjGG+B5IaIPkN
xx6K04r52vxUNoYLUan3EUOH9j42D7LjNeFBXXPU77uBXVCNkT1ZqyYI7NVMHKJzcaRwtuYjOd+M
wNEwOBSPluBeng2hP+AZM0H0bKeGUIkyoQiVqA02RsvyMoJG4urdhhNN382ooheic/xbamL5yENF
MMWQbsTW/yi1ocBlB6vODH3H18AlIuucNORSGf4qiHq7AqlsvzBUggh8njOMDH3GC7RzUflzGD/B
zTrc56EV4ri5s/a2SxORYrPaNEDYm4oYFj4UwtPRwzuPrm9vD7Aa8tDNYOEmVPbc30Qc7HSlWz4h
RSHnDUi7f9TVFw540imvXlxWGwnHdBPf7KStM7zxU9QK79H5eQK1/pFGmcND1ftc8j2T4UNwK/zd
40qFAive8+vhfvj2GSqPBl7epjraS6YoCQNx/ik3lnh1kbocn9JGlC4Gylb81L3qHdSKMYBWvZWC
k8QMTwMMBN3zL4sAmMvL5ivwKeaDR/rlNhFXOb0fo4epXTAHkVVWYhMguIL3ofJlUpgUi+jX3SjY
VqRILlC2JOGpzcvbm4aqP2ometSozWRchtdCwDZBVFwDYRMJD4QJ7cDn1rWdIRNJhSwWWchNmosK
RBx9Zb5UJ/O0TAKaPO1IR3FmKem0KokXWw7kyXelc73eqJvmst6YOH/CxURVi605CsTxD19P4rrD
yowYmsyJAc+MQHVGHvtDToNZHKuw2X3YWACcx1QRd6gAw39Q8SKGmekhcD2WvisRzp685VILPvGr
GNO1jna6U2mhm+sfG9867Cpx3taFlBuByrTmdevk9aF9NnN2OMsy7ApoBkVKDAJUVrpP61RD0lQR
nFpIXEZeAcnKtLSy1YCO1GuftKxbU3MI2FL3dsw4YEvZbsF2QMR+Xluq7vkAXvBEeJm6LygCgYTk
3FsHBKkKpdEd0MLJO8Q7B0ONPR/Kck/X9mmBmoDUw0rJePx6AIFonbKEgXq1m9TbWA1S/HQXMG1f
J2VqdPn1ga1cJwPsgQWyYrWQH7BII9G908RXKLlamwwmse8y+TVok0pyZlTPlCeJmR74vtZ+PVUJ
bLEFfp2yzwQaKFwMSESPLghfyZFJOaKwNe4sK1135NF0OsJuS0Wm3YDGRrxQTBpQ7EAjqvtyn17Z
iOebVK9rovQ1URlVfcJAi/oYBCRWVAqbgGfSXfmeRRnQJvlMYOUv0CwPpdJNcNcFaICtbjk2glZ5
Am4YPRdNvCEnsGj6tEoYnH5g2ZbtcRb5vfDxZatdFHShHarLy7FCMTrjXrIaMF6Vy8VwCDPJ1wv9
zhiYINKjllygBiqrB+uzgayerHmIJC1ihc3z6caiLiJ6XggdNpaZG9nyyMk2aBo3mOjlj5AOWBpl
6axoB/QArf00Bnu09jFXSWjLQRvWM8jgQNYIOoIsFmWB0GvsYAgxvLzGrbKBPl2Nm6kLiVY23S9w
xNA/XpwpLwgZhoff6c9nBJx2H0mJbuUMhMSGulpN9a2npG9riipPPW8CGm+OcRXe62CQj8aA+mQl
0yd932Z0gTCPat2TyFSRK9EjRgjsErgymlfPo5FFp7AnWsOD96qO2dDqS9HGyoDhkHjQz8yz/Gaw
zX4+HWvbdsLcru6jDLtaziF13UTzuGxN3d//x3eyxuGCEVeGuyME2P85iaPhBicsGZntvptVyXtd
iri2L1WRR5i8VaVcEv07l4UUP039eLYUaIWry+6BL7C7ZSWE4CbijSyWsd9fWn1kgfLqVK3p8wqK
ms6p8CHNgRuyhZpnbwExe1hgLGu+EXjE8wAGu4r/u+aic71RoNLVN/RV1W9wf0hcSFiGzMVuZE2/
pRJByKETYHRpOLWHpNMKH2Gkr6124PKmPwwaX0gOMqY7S8lpM4uPf/FXFUOo1eC6pMr0SRwc/kO3
xxgofmJQ0Hl6+iwR386/7uwhDoIgjfN9HuFdiAscWaIECYDnyUoza9q6O9jR0/fR7aIo0LH40xqg
N8kDET7Kvq/yamJsY9STShx4TL1HSsZxq/a0sYVE4vuikOKHCPrgHRfX9AvXgQp8qkH9OQ1lQAjA
WUCXFgEIr/EQE/dKuJs6JJ6XkBlJnZpNsdaU18NDMAW+i0G6FkvBG7ibY5EXGEtLjyYyT2FasTHi
musDsb60747yNLWU1YoDnqOvFkAu/VK5PID74JQC3IJNy9SlgYdP2XQ8iyyoT2SYc3FWw8FemIuH
toqVPHQuE8YMkCQfo12qj1Y8ukwRHcZlCihb/K8BnnQ3KIXThkD7ICduhVInjQOiQMCCyEWOxizB
U/80dOLujDQuYoNv9yun7A6czBGAEu7xE0rzeerfvGB5kj21uVryU5AkZPSaXI+teLNljCCX7fBO
G+A6M2pA9cNL22yPkb/2K+yud+IKxd4KS+glXuDQmALvRAlGWNj/XpWE9gZiLQfC19SKTF4HMMXa
jjzLFAWsD5x4UecCCIBTI7c1ZjOcWWqzoZno3nmzsXUed+aaL+g5tJRj4LLR7zQdNDWD9LbuA7Id
Z+NJoa/oDoZyO+err37PJmNpzZvYEv/2ajPNJ/JJs57SY3OBTdIPfCIGyNoRtLeIgGG+rqxHON9p
OIRwVW4JtUoAcCTamhBHKlzMc0BoivjzbbMhN69TirHTgwMs75ZX7O4PFPpEkz0i2N/oMjex08MM
AtQVi7iu8zAeLZoPDkpIGawnkocPdWyNQKcYNyhHgH2+e8Nah9sbO9okl9nTwFdbN0NrQ/ONF3IR
iF8ttA2qIRHbarI/VAQxjJV9HVOhLVp5GaWdMS2Zku8GJXNM6fn0VnqMqgUT3Ic5poLAZNJMMaYV
NnrLfvAWT2omGdPcO1VvB1jQPk0dUXgopneYq2SVZr2JVMu3Nx5lpF/EGh9fUqgrFI7XNMioGof3
SLXAxsG4JSm9QlB0j/eYgl/Ftldg9er2OILd7OlLERsZ7s61lfEl2ANBFH9I0leJCmDo2evnX7Gu
1V8WDZdpDwu9ntqVoCv7Gs90jVbTX+H5rlgJKXqSMoEQJ9urj1M0mW+Z5SgOdAHJkCb/OtkCpTsB
3HEXmxhJs1uo01cLNGARr8h/Ze9Lixg8g/Uj+A27JQW8ZwGQIJXz+rqcw3tOVsZTMleVae5iGHbZ
UAeWkbNzpntt0XrLtO4CQS4AiIl7S+4eFm43PuYOgoBpXYwgOBNjMgu63EtPfRjO2jCITOASiEaY
o8G0oTd/xfNll7KPpqLljWRkZ+pPfo3IzIxg6IpXPctHWxA1kHbGfq4V3j3yMMBg94VpF/SXuSn7
t1FUsFPtv1YpROysg9UvtvNUEoxQkVc5/R6ZplYr/MCntK8A50XotheRI6LOfaPAK0A1EPx7mz4q
yK1JMYhW53RyK7LKbbQiqK4vAZKB7QfA3Mg3PMuVVx5FJ7z0DS/7dCq2mTOYI4/wJnMbVDnEQU1A
SWHCWRKOhgRwKhtwOQCVd9uba/H8jxvoSaWDdITlg5sj+HpxjCiYMMPuaISzBVw3jEyA7W21kGpA
1xh3jbLUSH3/1EITCt6AeQZG2BpjMAEV8iKMPS9gDUiBQLOLRzPFF4OYi8D/E+IML7fn8k8ZBx9M
LN5l/6wufUfBvTtHrlbdXYSQWAGsrG7i3xi/3WgCIyshCmoiGRFkrbxoJ1H9hTqSAehuLJtaqLNC
frpFcTfWYg5wC2H6wl5O7cosW4BUWsHVRN6tRr6Hr2Ej8mO5aGU3piSkg7mCPm90u4Ior200pGbB
MgRxlfYkwA6zuP/RnPLEOzxmZbKCYE7Cz9t7jRbpM37/1M/10f0JG3FUZj7FoOtilaTp3DpU6OBp
lhtlgFwNsUeMI++G95MSdHy5AocIgCqnBoIQTk1WmiDTr91wuvTZatoHki/7zvt0fxEwBDUqyV0h
gQVYx60LP5MRb913aM7RYXCvRJbTaqLwggyQhvU2VIYMOxGMc0iZWn8K05WQ2YC/jjaQru4VfJeU
qQOBW+kJ0jNAvl0Yya0HMmueVG+atXAmwl3NV2V6XjkAp/RnWFc/v7ncmnd1G+C1b4PvJLuvuEZF
mAL/+JsQ5GiyjIM4UcQz+VKt2MA1IqpiaBh9gEiFCuDGhwyY3gqv5k9b4+oLm+ipcDKHgpVagqR+
jomaJeT+fHxpnPU8/wCJfZu9BHk0Rdy9Yb+XXRaustFoSqHA9eLJGvu5tL+Ke+ssK9oWNzUBnCZG
KxrhC7I00/NBeCfFRYGkYsk8lr2sPTSx8IWBf9dwfRlcZfQjzyKSqz4VUV43P1nOEfoDRXDszR6O
46X+ga9xjO6tnXz4sInJclxYcO7FaxiomlaW58Me5S0J7iIVGEUsPU25/3tqcRnwdE9qaqbHOnba
0cmg/SNVlH0ULLo9YEomBWtYfQRpBP2UWtaZMym97yKIaqkfZTxvIOA8O3mocW0ZvoE9QSUHRDe/
Rhkf/Taoh4I+0cyoY5j6LeTxwU8Pz/t/t6JVj7OGeF05deRc8DMAAZDyGpQEePEXfzEd4KCxbp7T
W01INUTi6uJbtVhy0cHTmAQ8UDEI0JYJJ2mt1LetbjypDL1EpbZQ4hCiSdZ1tzNNOfF3Bvu0sVE2
LReWmEgsPEpua1PRGHgrcZfAFpchtt7XZIxf3TB7TeAwVUighMVqeljaOdq1gajx2bwuaUqjxSOn
MYd+ppfmNUNzCy+XezqCpUcR4/bTfzxZdrvNjkas9KpbOf7/VkuVvgE//iaxe+8iwQKVkQV3gii0
KUPC+bliON2aRVXOvyiHhsO3bt6BTJttTouadZNWyWxGj2LW8Zh8vtp9LLzMs89AeKiuKjxkl3Nk
3zMRMnF0bu4ufQsbVkjw8ZmNUJeSegE1KItI8KDsmX8gUFBk9NlySZEw095rFf71hCfp8aZTlDFK
4JfW/Br8QTZkIRHyNQsN+u7tyRjJH8CAvmBe6ji+WwSHLy/oHMYLpFNxGQPi//NkOmyPeyoluDwu
4rCN439qhvGp8OuO0g+P4pFVPctrGC+XNa6ltiQwKK6VTJUrXV5Ja7j0Ta5uMcIYCBbkI7wZqg7J
tyibPhjh7aStb5qs629y3mKvFEEcCsqQgJSl447uf/Q0cLzdg0/0AV6iqxrlw3caxMC+u50mpPzF
UkG3VZ/Oqhi2s+qN3oeHvGkoTm5X7t6mpF3usx0eU8v8x/fJ0Qop0hymfIAMpUSVBVX5NEdWbiYT
/ZBYnWjHmFsuO1eq9XKxf2bBm/OKYfDTw7/m347HGOyHFwP9QU5T1RQRmL0QwBDTFtaNc576jj+M
0H7UjGI2XvdsBkUyjCbO3oYEdSFYAc4XU8D7g+qsV9rNZ2j/Wo9aNKh6bBlxDn4SI/0oInhgZW+M
arKMduwFbJOqAKEZw3YHVOutK4sVUC5dqjg3qvyq3p2Lk4UjbbnZuR/xLTPLlT4QI4Yesi8cCgOl
2euFgCNg7BLBQvlZYz7iDI7V8Mg5l1vcuEfOAbSFA2BtlYIbgq951hoF6K8Thpu0UUVyylAJwT3X
XSBojI99e1xwXTAre0X9M4rdXJRCMgIgmNnBf8w7vrDaXYpYuXHGRCQpZsqC3UIv8DbX+O9rhfwF
bwF0af5fB2Qioyoty6eNEyFSbcq9XiwbO+rux+v/IvK/AVNQNTSCgQFJ36J0YhEuzA902AlA63QH
+8GwZx0d5C8oFFhSH8cmWBQrhQJxEkNn8srK3BlfX1uomCuwtbYFTn5IVenYDGThXrqWbJFwmIg3
4RyiAwUL+WgqydK15b9w76aq5d4XGGbKjDcxQS93k1R0Zt2pV9LGTq0WGGI5KVHwbkqoDYrNgaPY
iLao+JSVevVL6i5XwP08y0n1oAx7Mwq9WtF5kjYN2GUMqXd/vI7P0klAdNt6vEBBSl2pEZeM7MuQ
ec+TNflje4dCpUTJ7O7kjbvNHva6aTTGCUfG8lF+hxvc/W8SOTBRtPdpDi8Yq5tyUSpuyEJLE9MB
ai9zztn57t/gtmc9aSfgekXHkPKz4UFFzEIgNobu8iaFyvDgmg6920g/0SPEZbA0KoRYIjgfAugg
pgrcAuqitmVS/1X1C9eiFxMVmF6Nn+/Js+h9tfHEhZoqXltDdec2aJdgouuirusPK1qCSvd4Jn9j
MVb4mfQtB7LryWGDybiC4KfXsE+Kc+BTL7Injfr60k/5ZcVSSM4TmNCNuqA5+zWvAXDhQT/nyydG
etwzm6eBBBfBv4t3VQL/W4OLowBr60azwXsCKdDztw32X9pM5AW8vAzAovTVeRoKdWeBgK+WBDKQ
qqbbusriTZK7v5RlgM2GSwKyA42YuJdAOeHgnR6A6n67BbQWQMGb134JMVNhfn7/7YJfzCz2G11b
VnvHD4rZvfdmTGv9dYmetusa/Nx4agMmzEElsvfcO4lf7NwK6dmFvE4132+ufkXbIbeNDyrGVGCl
gNlX8JFxu6cRZvijLl5CmcbbUW5NwdIpuM8Gbrag9n7u8VcbTB+XaGdxIQrBFU9M+Im6ZZJ80AdP
KQr/53nB69EyEQiSNefVl+KHoPneRRoW4ZzloQNEmhJ51uUMJHxHCINsprcydUgEFSMcuV9POglV
cJMNtAY6TiSDK7z+emt4pojvcmMN6vQYkw17S8eG4dzSUWindT7+/PNoJI3krFyMhWlEfsSe+I/o
hAUXTonu5xYmkPjf2gphKiwmMDE+CUt19PRPIj65qq68heo7oT0/UkjDRSrxNWJ6JImZM0tf2FAd
Tp5LCNNr/NeZFULmfjKQEoxpxqB83oEPSt/S/feFOsoUKa6n9NIMVfgCBZqeIS6oFs2BsNbvV4zJ
hMPrFYY8QYJS7R4+ihqS3Lh0L46SS6I9EAHG8A15z6YPBled5v72KtxsytAmtzk39OTGSB6GJgs3
URXOH7ystwALQ3QM8oqska0PXj7lrP0pKpL7fjvvNimSE+jimDNIQ5oh8pXB+TVrUbfl2RJ1oK0R
VEh7/5DzMV0LUwiF7cydqnbva44xy1BIZM0Pd+INLRpzjRvf/9yk2rFSi59mp+Fkz5Cu21LW4aGv
beW6CAGrzI/wFBZaVpQqG7FMWncCUDQRw4UO7gjhAofSuegJZxgg2kupgFj4sQkPjsWqmU6lCDIH
TVekswqEWV9YDEdczKGb/AdElV64awF2v1b4RgYFYh2KGGW2pRgwyeG3sw+y+S5Tea8McCX0GoRB
RGXPWCDJp9FqHs1FTDlGnaFxJbu4Kh5a4kjAAWgcVaEYUu+QBAcDdAicPBz2WnPTveMPBsw32gip
81dw/dbIAXN/CwwggzfLD6jm6WoE91e+5ZBevDu1YbxtcDFnAQx1wrZenMkF/nwFdW8NxI56gaFz
fQ/OTEsCxAW6/yCfK9IuaKi+OQ1YHERtuj3D5A3JTJdLZOpcJe7LRQdg09YaILsvCeZj82O+2gXI
5JEcUwbG0EGVD9IZ9ZQS4SNrC11sC5bDKmjyQnByf6TjZUERBwVCypk4iFcT1jnf7HjpLtt2Ukgi
rjpTBiLzYI8DoZ5wHvs9l/KJno3tDmGDLbGZSVLMJsEW8YT+vgwsdS9S38dfMeyLasmHk2PIubOj
fD9IwfR8sdfIf03zPdCURwY0vfAEUXpAbxyyFfsJKJq/O2rpixoXmL1eEVmtm0CZElAlZNa3gPkI
uTweyCDWfdjV/ICUXO2kgGOrl8c3wKE6ge0KwosF91gJKFmx3KdJxEs6FwQel23580qa3RqyFYHs
P+oXZaLZhoj+0oY//HTWhdtHu7A/XI9beWom2jokonCgw2x7W4ES0DeY+uVgFd9Y7xlWLecEXh9y
I8E3Nkhe/ncizMYznmuDeZe9Sez/rcTcJ/W0SNFF72DFc8PLcbUa7zdHb/Z+T7GL5sd9opf0ls2X
Tee6m9tYe7rwegRlAddb2s3jeCW7Yw+qsOecn5MpdHMP1TktHaPPOUCQuQS7mynhqqSDRe+hBE2R
JuRC2rXl53wjuO2ByoHJDYAhfWtl6FYT84s5HBAcCKmrQGwWNWodQvKL368xNRGSCitudVQaIf6c
ju6pCY3VENvTkF6o1hvdyyjjcCjZMZMAU21+wlYrjnO7En54urP/Lr06YS53mhWS/ekAtSEqYSQr
BD/vuR2XvaubZUTpIZixRloMWwEVnMAsCITWVhtEMnunkkZkFO/j7cmbyRPzj7ir6bn+mtgrL3ka
G0HgVKYAenCzbUTWvMxbi/kXuUXk7jJ3g6mUrRLIqTGmKmtf772J5cgNsYfPsRAKKk936zCfLPr1
jneZK3argD99VuU4+CHAKkmlMICzH6cMxjaLvJUDdVrFEZdpBrQLH9sd71/3G9YD/Y2pFzNOBkpz
OmtfnBOHzyCKumAnsd7FmZaxpMM8SJfb6nBCazuVo8KRlTHrg20m01BtS/cdhFwj9FYz0DxHWFJu
/l1+A8ggvfg2SZjNmTIaoSm1PGWV/pQcT1Un8Om0kk6KzrLtPpc2tnACRUtuamdEeb787j1SG3v4
aGpF0kiYOTf8waCoK/tFnJPOUzyROVH8XKhtt9Nxnxp6p1P0P0KsK2tYRpjcB6ViYrbhIIcSKRf3
9iQksPYJlIO7D2yOdsBdnm7AFUDTfsu1/iY6o5Fn1BAIjXFinaAAiYxkdjTDZfHh2ihysKiLKpUg
5dOQWe5mno0nDCI1Q5dsG6PvduHwdjHHbJtmzJ4jBe4ItuIDsheiQDutrembqh1X4jBX5ape0aKo
p5dxQGworwHnhVLj+hSFlqwC3+gSdpZRFWhuMyTlNIYqht/H/4sVOBI9+WMj/0AvrD1CLyFsDTPj
pjpTDfuz7wFvcN+hEukUkKhqm0xzXsoyJ55WC0QJOgvWch5Z7oB7blcbgWBxO2CzWNCAwp8YpaEI
jj/fYBjYs2b7QTFs6X/1cXTzTw12samdrYkEb5rDlLtGiXxDTA7IfuOqyR91GP3/SjdCEcpH4DJ7
xGi7d2JFY58HpHWc1Kx69qJeCZvYsos0tyPic4XwT2S/KleQnzpOZ2BbC2JwjcGteKE79vQFmy2y
fQxP8y+CK5rAL2RPkTpM87CHRmd4JQhZwbMVhJavMGULaAV8XPe9Gmk3wAahx+XGJ56bbznO8bfL
xSyGl89XpqCekQYCnVRdYc++Y/oxV3wSzVoUlcTa0iETKSZUjgn5rnoZrTE2QPM1MQl7w2q3LInl
TAZcYwaXBtY6lsB8btPbPOsuKEEf6QaA9pmE96w6gMvuqaNywD+H2vPX00r7H405KqyYbErQBnTH
yJqBnDJbeITuC4fL5dOqebww8RxhSOUit371aSa/3Va2ljV3UAD15bBXl7Gdwz+ZXijaJijsxbdV
jBQt05IoS/aFDqwSzGFzz9xrpqUZqNHiDZSpQENlfxAYlWUBK/OVRDse62YHmD+CPP0mgLhkFVNY
u2mTHrNGRR9OR3CzgvDJ6fSecmjUTyHjTX2HEAZvle3cT0WCAgRvz5NjGGi0ipyCcZcrX5LCNEDS
WKHT4RK7OPOd+UCeWArPTlDjqIZog/3u7NpIqv3Q0Q7iT9Slckc1xBviFynZUvnsw3gLun9ydKXH
1NXrCwXBl/PM0WnOhp+fBSQlV0iLafpJh5khh+wJ4AHkxr6FNBKlTTPMh0o7v4GD5NiFiX9pmVQN
D15WeH7DkKxMkC8HSovyYl8JB3c82MHTIXVklgNfHR6w8stFeXQplbZemEqr15viBQZzl4ljH5pc
FLvcUo75dMLmW6SNQj085dhvwyihoXn0nXj+sjljJZiwRstXEj9EcUNMgaaZq8JCSgvBAj4/SySH
j+AsGAwGB7n4VeQom32ZcmT7JUXAJEwviqO5u56ma6Tu841kCHtpyTcnj123waOCYLZ50M69/hbH
wztVhgmGSSEJH7VQPMMJveqREWG7Q/QLsGmRPbKDCz2l397E6b9uK4j/RagnlNXPuxvtA29Wmamw
TwhfWGIx5SkbJnBlx2KKfJHq0ud461/zLAMSgNEP1hJ45RsAmsmqFSISaFkWuajFiEgsY5x3GJ68
6PfFKq9U3MYHAbYs0mtanY7MDCTX2lcvDseywBh9qX1Cmks5WExlbGHhDWDQxBJxkZlQs8tNrHH0
CKkzzRSjZGo3MM4jivmmsB+92U8bYdXZWBm+f87q0gql6Ga95g5ndC2eNrHsyAlHnJ8OjIpQb0Cp
lYygcTT5yxlYU3CAC62WxLqnAd0Kdu3NpSZFtVRrBexdkNFGhXzeEApHdWcu0T8S9cxlip4+f1Um
XpMTPjDAyFJqz93VskNOAYHeKe0o+8moYs9w2Msl6I9P8D4fp+qjvZTujQoWTyYlw2wS2IoA6uLP
BVYdnUDrVUT5tfrjl4TCodF/z56f4aBNIPv+ID4XhDOKY57vFfHok55UZ5ZRU74921sGvd2zGkZD
/+jlSQlem1DAeL68x19dbFCpzsRCO/xLlAPVwwWRuIy4h3bB9CJHAkjWUpl+To6656PFeaWkGrRm
H4uyZ/WCPT3Hs8oGR0Qz3Gq3bn9IiwkRxm2nLgJRkgd33VimC3rFS8gUuM/aeNKHdW/FBUsLneqo
yGFEpaaplkxufwdpdHvIRdQozrukQN2+o3tDuhBwk8cKWpDRb7aZ7mqreEoToS0H3sq+lQskapwi
yzhxZoEzWyTWMz5rS1+JQ/OXQuGePWnTdKdUar6fB2fz0/dCDYeMOfYggbAjL71SQW/ab6kMcSyy
8W3jyGcTC+TF3cLBES0hpG6iyO2iSCA/q6LiaQ86sNSYyVFq/+z12wZW6zgLNgXXFjTb9zkjOM1a
pSPcoZNKrSEPco81tnvYvH/mOApxDT+tjgY9X3aMxznF459l4dx76irEP+1/sji2Cd4u/sEUOC3o
tc3dlA7Nkgp1JK9US1lqfPi5W4Bo4d5bw4xQCIXFBkOuLepPx3ob+65Ovedzs16CjWRC/UF7GZQS
M5ko7y16M/r271Wx3zouBbUbkFQ5BaVia8aGeYIiUSmPZH3tVvgbbbNV05GwmDhQv/pdunySQUFz
T3u4y+6Z+DW6Fc2nNMI21KtoRPP7zIl4RQeSoTNzJ4LklupTwD/ubaGFSuGCHBkJEc1re70HPQcv
/rSNzblmfjnSHC/sLUB9211MYUwBiflzjeQvSIwa6h2Vd5L1Lc0qHRXTgJaHwRSoNIE3OfE8m78A
AGKObDb05l/RcnjRSs+guPumY3UTbjLRjjrrzztmRgSppofdbhBgE8q3SYV4SHvlJKSmEY+wSoKo
17YJg38694kUeNrpYwB33S6ln730PzgPTqeKL54oJVR/9bN9v+JYjmEsbB0a1MXtzJ+A23WhOlqv
ZlSew7yQD6DuaGlB11YJAMN8K371h4g+9iWV+ZzvSJkXZOUfADQjZ9wg0Ko6Yx/nY7dqcowiYFOL
wuK9vk1KvPC6OVlOERhf50C9rodyrnAS5Pf1OymdaHFvwOkxSxqczfBqP9a8YR6btMOoxGe87Zzc
VQLvmh0QfKN2DNHRBwQG+EnhReBciKYKDX2XFy2cp3wYxgxOvbzmeyXJGakVMVi55zH7nHkAwvCa
56Uj7qCSqBsZxAeXNZFTQDRMKE/6p1ujUsO2qbfTvRKtdknIh5ObcnUUydgFs4ZD4gP9P0xSZEO0
cbJmx39vWeqUNTBWAZLUTC9etE1w9dtp4AlCdmNk8ARD1+yzz8BXGjiLPPOyIpsOubYon4vf5bck
4YWBypv6p/IZX3oK8UuWozeMVhPrCnxwSbjlXvog/iX55G2s2ikWQe0lRQPtOYHsYCV0jKChu5IA
dzqnudtHGtmB1yb8ljcnO6X43yaCWgX4fdeGgr2m1Hoa/WfZa/cLOTta4EmTdfGmO5SShgVvq/cY
crMKJ6A0MRvClHM6owas0e1hwrsyeBJjJFEI1LOPb3h+wMV17aqRW4ys/I7cE3gvzJ0U5MqwiXNN
WT8qWszOkL0mfd4dpyVsliqiaj7vXtdPOYXW6FrwzZIPhLxQoJLLNfdi+3BenTksLsABSWYdW8nO
ryGEA7IaFOw0LK0PlA24tQedjfsJziEqtvpEou8BXy3QH8EonyDKOuqDiQGn92569BiVBD7sP5a/
XxcwSW9zNojt2HBpboNoEYKRt3N8NJYOHj3qIRhkrBdlE6iuc5VyLWiPYiKAIA42eggFOWyOh9bW
jopMZEaBb0heCX/8dy6vR0rtO/CgMQI96+0lE5MpVFPw9pHphNMvzDqwopCs3DEuLqynLcesO4Ep
2nEoM82sDlPuy7dpYTREjg+UQYNazQPQeNo6C2pHVaKWQ7eL/hv5YEx1mZqJZXJA6NSDFrehx2Y2
+wQh9906Wl5A4sSWD7iwC+1U385f+zOYFrF85KQKIN2G/iPMMAH0lLVAtKHsSaVYGxiUpdxN63Xn
LpElf+2esoZeARM2XdskS8rOoE7pW8ijAwOw9I0Jr+evCD/bysgndNY8ux9B9ruDU2i2L7Q+LDLf
AlMZLXJvQBGUYyCbly3JGyd1LWS9GA7H122IvAmt06VrxBiT3x27xCkw+SozwBn5s+F/sz+OlMcf
NTY7lvzu/Nrq/r0czrTgFNLw/W3PjT+dmvyUBl8hQI0iYolrqbzZTwXRBNYx284HaaM+oxPLhd9a
15Bj8PML3Yun81N8RIxIM+4yw832Xz7Vec3ew7IacF+vNl6SFlb5/VuUiiE5D5WIINCAJSV6jpQA
UEiXSYMbS94pyGXoU1kghPTViHtFKAPLkeXgLJwUh9VpuQhP2rXzWVN1Vv5ZlOfy46Pl+6psegQj
IlrHujYa5tl4ChbT7Ragi6PRXzgfUubsFs2bhgeuL88hQUNv5RPrv4TmLU1gveBkZYq8MjgIIkx9
OmYI1NVtG5coxRT0feIYTArQabeYuOQgUNkY9Xa5PzOm7DBHZsmlUB+PYN2bg6nybHksrLHU5lfu
lrfX1AZf5dDtTFpBxfPQnjbboAieCnFpjoqCgrEMw1yDmjyBbyo9IzZBQVLJSfVmtwcQzn2PnsaM
U9vIsB6IwpQWagdEkQk4UAoQM4xq9hRdyOMXlknV6F3vs5bRrhLfgxkZJmpXHqI0iAP5VOY6DLfZ
MRCKMeAEFig9a7NXfoBYT+GtuDYPIgCNRa1Clr979hqTgO2E+GHogTvCSUSEtQ8XhSATu8LgmbT5
4n2CB6duhOUVLqiHIjAjLUImDlqyrAmbakSFwzipKqYuSrDl/F+yh2Ym3KXvGa3McAWJPn3xuAQR
aAynhOjE5rQnwsgJZkxUzcKJ/oA9AM2/y1A+JAFRnlOKWEQWGp0igVjpxLRwa72G1GS3WkBQDCvh
y49lwIzHOoVpd3MgmwP8GMuK7Fk5jzDYF3VjMz8WQVpc8XYlnGtYBgJRdI6WlU4CN8YADLrvEEEo
MJNMwzKtozSP69eZMQbgVHO9tM9iDyi1qRGqktBdeUgh7PjNKunXZbWQbGWI+i4HJyPro8oCnETc
Md/mtpndoNPGHWqFWpAFpUV7A3VJOUOnXhMSOeppHgRU+6PtlAXUBiErRnEP6Tkhc2tmUqGQiHMu
05x4WGpzp3wlfY82NgdPnvMy0kJULHBgR2y7Ve2GrTDKwISJKGkWNgP/grOMdp2vYo4sjGEcwmhI
joAn5x7pgeyG9w2zgSDce/zKIGIdLwHP/bbUkVk5I/R5KfdAXAhYIGpPm+ib2NLjTNikGrd6N0oO
CnvkNKmaSfirSk7mhEEAmCTK6KVdIJgkfG0SjWD7slJI1j3UG2rDNyXzq+IG5vPzMl8PVstBtV3p
jIXWCWdEJU1ZIwGw/Nq53RDgNy4mQ/zIt3wzYHUo/J7zx2YQ9A4wyKBC79sOsMhVx3jctDtB5DJZ
wd0+s5b8qW+LIunobgFuW67YIwSWUdwp92ayZ1tQFA3qSRiiDVHaBCUtdDniK/tgRwOv07V9/RJl
lU0hwL3WwVRDHnYXukX4IS6apwn+7SGY/fjG8f2I34ii+jAb8ZrvMXcfFLIn0cvran6/fLuFEVt1
F5cbCx+0cx8pLBuKpSuKGmcqw4pjt/jeV4Fma4ukrMsqONCHfiewhdMuAgQJbucw1tE02d6F50Lf
sJOCvv2rEDJ7f4APUyqLsJu1Ze4yUnrRIkYYETrTlVmKKspQlT8yWAc7LWo68TX6bI9c9/4fGcr/
O6BAz+CcjdnT46R3cMhDZpZMNI6Df+vV18Z5MjkrGA2GgpOjwrCHG+L6Sho/252u7QXSFxOydJVG
C13HNwu+XU8EA5K1jYCi9CARuZQLvKv9YwhplPON4DA5I52aVPl8wfRQUvEiOXZa8jnKbtoIVpFG
7cN08PR6hl1jWdpwawa/UHYfIPIA5Rr/iuIKPvmVauTMNEFp/gq2emRw+2Su7TPY6o7u3ZqGFk7f
kmg9jwpxPvLVbXMXbaZxzPQdJEX3N1M2vHqk3dErzGeNv3Yge39ayrSbI9u+fIaHSitkyhd2r2NE
sTbtECD0y6tm0DG8zcoMtOmolSeCx71+x+DpXhaYx2rHgdvjTxRa1HVmq/EJDmW9iQ0Lxl3oZikZ
1pSn7L87rl43HD0YyAt54UIjhAplvo0OwWf4WKHZZK1HnLj89XSpfVws9lUS/VYSkBVicNkdFODP
YnF7Zill38sCl7ThJByd7hDxH2nOCQf7Oc7CEFzvdG5nB/tUojrfkUVQlnrrWTPqv0nJnEY2+uwx
5EJKHYaEYaXOge4b7zYgIkr7Paxn+ZbdSTda6hivJDTb+TjrzYHD3PC3uLPbS2Oc3Isg28v5qmUw
1ELklmUO44UcIV0n/FHRdYZvNa6JmlScxl4ntED53+jKUEv/bqPhJJjGHfG0HO26E292PdiA7HAX
FDxdBwk7yXVUuxx4lAuq8qTqR50wUaeVFByxkQJGnyk18NMJUqMQ0rLXHojbFhYDWvUVtXIS8SpH
0Nr9xsPux1FgUNAFa+LptmFNkh7kqI5fN4VdfkE/gKNfA2yu7QffHn+o16DzJZtF3uOnIohUoRbs
yYvJojcItB05vqsLmUrqV90na0az58QOltM03MroFSfg7IGB3U2OBHi1TemCK2vTS42BtCEBaDFp
uAOwh5auV87ZGlY1w01Cjho+aWSAVtTd8sONY7YXnm+F1zQs7MqOV/sbqQ+2SH73JRTNDjLuQLxK
3EpL12kX0ycAv68VQLGDKPyezKwO3lJiNAKr42/TCoy/T6dP9jexFdAtzjRwCiUmxTq8ysYWt+d+
3HwvA9yWT2mumQkfH0I8KIiskQuEiVDfbDHQiqz7lavsDKQfAzFaR3m0oyDWqKFeUhMGLVsv922d
GCYdIov3V8HcduCn7Z9ToD9jzhAc0Hhu/fVK8zh6+7nXfDVib4MXkcl1dVpfQeC5OG2NHMyXaOQY
jgGz7FO0gf9eJfQR4PJH30u/1YJH5jafLWQGqpdYOTeiHoCU6yTfVzKtcpbuuLCbjYnwG/5fQ4gT
d/+9Ymki7w3OYScrP8+0WR4xxavIHcYOG9rCj7SoDIz8FCGRsxsvSXUppkB7jBHDXAsKFy6hZxnh
S2ObxoeYZke7OOOlivsjNGe04TGpxZaZsBJS4PCes5V/XRYR01raSe5G5PhVxh34VWYq39WIV1a/
ElxZMdHbaeydjGObyqHowZHftR+cGrQsxsoq3JAnTPYpZWWQ2RoPdZbuUVSJoXArTzDGwHwPgIyE
zgO9oLty6H37wOIjiMCglpr2mraY38trzaq0tH8QkqPljt9gSKHf1SL9iDrQQcRsetwQLoIuwJyC
lCUcOyEG+UUsHwAUJAinPLSuB1pFGbyhwfpmETWwEqeCC3Not3/pU2DWo6t1wDlmwtKd4wmwOoou
SCmSxDtLsZ1KtQDh48etr/0u8IAW1r7tqjsIHQKOilCyzk6Wxlx06sVUBY0oaveQOT5V07ns/YgQ
RbF2pZucICpDtIaCe5vGvzIoL+iyo3BmWCRE2LP54OAVfIGVXP63MeBNLvHEAEMHE/KT+Do6p9Xm
QpVMrbGD68NYaEp4OOEY7779cuZCKUa9jRVmw348ZLm301Fvuf+ki9Xw4UujmYlKf31CneM1cZ1o
0G0hIRi3AL6+CqPWd6PQ42IAqlgrJkTUYU2s/+EjQ/XdinQATKiyxreFKOyVMKC0g+yJVfGZByob
IbCQh1HDEHhpCswLWbg1tP8i6drD75yf8Rk6zT2/xjVOUNZZNGwIFOpO4iaIvAKu3xVVYs4nF8KW
QZsOtGHRhyheDGSRDSMdzwrtVxl8JXmotwXVVGQeTZ/tolNf8n3f5ZXBmk8BALe1RiCQ5pdn1khF
7+ugHKo8KWt657TOs7fZRzeC/vlp3SjzYOMYDNR063WYM/w1MNwAFGOrgBsibkvYlS/h7eRpSlsK
RZFtf1+cBMyVULzyyFhmZi9EKUjR9fnhL3WZ0NGDeTTnp52fYZMdK7jXaKYz/1F26BaJST8d9M0+
VcOb4foMuXUmGrqPEhFLtiNWkmrjS9LAJrNh2fVUGm0hl/wdTHNNqbkCJ5W9kGCKgjcU7bygBwqS
M9QE6beATBy60jqkN5WcJ9c6Uo8CkN6jVVoy+LOEHYXbYp3nqWw3qbKtpawBuz7yGllO2kBB4Tl+
ABlKCbQo0zZZSV5C+cHwNH5N4LFnULznaYpEqGBKy+tbbS5AQ6YOpelg2y1BcvaoAByWvZ2UtL+B
IG+U+1PuM5WMK5CWLfeHHIgYCETuTGosmTAgLDicA/enyG/JbFqr7EUPW9xdKLxrAHBUfUTn2ZiO
o8fqmYtNomBfCu0QpS9IY3vW+5p6acUPbUmeILP4zQo5KTePQiayxkjrj0M3pTfQ1B4JMwPMwUGd
N71bhPQxr8HopLLMpj2lmFcOCEniOky6I6rJgfrqYTvgMOGW5Vmj5jxqC/LXcEAMaRya8SBDz59F
9M9nubkrR9Sj2cW7lH7Dy6mL5iei+u4YhgjRFLau1ucDpFQbngSNnJeqw9mM+RsN+WkAQMnBQpO0
5b5lRESOo7+hnHEURsOL8nAYVN8Ed9sp2D4b344RnsaLIy5TCO8l7VCH1hz7k7ude0GzqDh+07i7
T8GkAqVjlq+YGieVJRjkTDEem6vTfNKUP0W6G/qXyzkE1djRt2eVdb9QlyoVLzFG2ytiuNtagjWR
XVOQacRwSs0nHyhcWpUCzpFH8+UqSXa1PiCUuNk6QMtHnybu6NQrCQUz8zG2+0ieSl2FRW/UnBFI
ZN4lZ1EXqPLinIXZuPDk+vugl1hfFI6c5IcEqQQqNrey2Gb/GrVxxrtd1ImuiQfxQp1bsnuhJroV
yuy81FB0fbw/1f2B96GSE3oEG0iOKZrdqiWaYXCO4MvsqKK9geuqRAXkNmJvfwJlYiVEPLawVsWq
h2fJ7VUvfzFIyGyp12O1+iHES9ge49tr8bXgbzBBUXBSy9/G1Xgi7Xr+pBe8spDm/TzG+esuKpFO
EVJM5Lg7NKLZsfdSgESWrUzSz9xpYDLhuw8h9YpZ+tu8kNiIJhnleF1weCxu66oZ+SqwkgHaoYkz
E/5iai7ejT7vFE3Kk+b5j4YS0GmbUDluvHKBLP1WvIZrgmVtvjkWKSB+gCsiNiJT/KATeOKTz9hO
47QQL+2JRM80Bzm2Ws/9qoYxpe1g0Xt5HxH1MY5EgaKQfiwtllaScxMDgtE922DYGwLxbqRtb0ql
L2XXw7hhdQRTO5hfObtePob+MlIJkP+IpOjzqCUQpeoh2B8XKEtcWh650Vp0w+BIIHtPG5QQ0SLJ
qFHlWj/i4JPKeR4k6feBU9RQ+IS5IwUtXFhQFtYx1VX7/cSt5KJoV2vLmYzvQ6N4dxWXHbzn1FHN
WpSW5vtQHevMGaTH69OOJrAZ7NzwCcy/I4dnVcThn/WSOgbcXBT3Ryes1tcqLvM7Pb8F/QloqSol
4h7MKrQY9WYeCxQ6UkQ9YEGmMZGXWTnz2YvENmC/Zo94II0ZRWJiFtvoLDj+hW4EI+wSv/LAcSWE
FzIkTmQarBazZNABin21OGrKgnwlTaadnFXveg16RMSf2ZZPOIZldwPvc+UUMQTQJ3uNfe6s0orA
vbofPBjgw7OKGKr/DIWZGVHDtvO3pPvcTtT5J5W86uM6Q3OtXDBCg1XT8OkStkXrXC2PBO7Gtk2x
weuhWV3optnPTcoNTzFHcSKyiEiFMGyfjueDrfgy66zDCKGfP1k2kXgqIJ9vZIy+b5iGY9r6Yel3
qz25FrNOArQ3FKVgxBlYAweeZxd2TvCy7G2EaIMq8TRwF8YzQQ0K9rj+a6ieRFeF5iem2x1j5b2y
k4LttjlD+/4R7yb/vs8xABYBdXk+dsfA2np1PLCTRVFqmPujdhch0UF8/2Bd7WXRzONPzgHyxEsY
3HKYe9tcpbgp8QBurTNAoLM7U8JoJwUyb1h8l0NC2bC6OPk71gpJIS5ZpG1FO2EfZYCYvU4bOpgv
OknhPpnNN0wCEtKLvlPm7LFXgl9z1s+qWX7v6hVttOuNNSzaVqaCNurCD6vo4Ugs308modF8DG5c
iEc9T0lJbMkPsRNEB+O6QwF5H3nKs4YNtnOi9IOAceuXBTAp8bA2zaBkV8BjjkYUwOSKmditbmQj
/wSb3zTf1pM7TrHwCqR1gYwPuQbIgNgJa++RgkrGs3+A7MqqKM9T/SrRaOwcghkBy+akEL8Ag90y
+oWAxWx32fc8Ovi5Tc2rNkx3W0zWDhs6tEg7WdMi7RuzOHkuQqUNz6BZOwxIRGq+unWXwaGmn7el
hfpLMXAbdEWRztZlEWiPhScXHxM+Yh7sCU7KtTRxrH9Knt/ex+9Kwe4/diJQoUc/SFziL2iBm9fU
zPcs0ItrKjx+GubgVlnECpq6LbGBvDKOCqSbZyIP0n8R997mSdyzI/Py4qWzgGRrRkTbhy/fQo8d
Aup+FYuN+Yw1guky4wrsQWNKRqrNhKEZWPgUho91EzlWqYox3FuA+wDqJKSRhtEW2AHje+WJzoA8
FOL+I2GSN7rv7uPi4BTY9UXkaEPUefH0jgdllPWvf/qZ+tt8JFEmcyCBe0Psu2N/dV5+WsWWLXZf
FzM1vSXKnLbkZsMnRvw3wJRYgtO1XyJhELUWA5XvvXKzdx6zTdOInro0FF36OMLYLlUGYBZWFt65
ry4O87RTcA2dWubQ6zJlU6PsAq5aW6AMteJq38aBBgVt4uvbRi2mZYDwzdk7zI2b4BWRXLGND8t3
4HIQdpqsnL7XcT1BJaJpnDyKYNGWJh6N/zTCKx9IHktWPA/7ejjQ77DJNNODg/qmg/vF0dt7kuWJ
HI/OfgCSoyv6S9by5KPAJ0m6sOi0824maCo544hdup3GaKS6eBjX29x4qC6FhHlEgBUWz0a0ozKq
VizPvnd9I8X+8yoqAQBIEyQacp6bmlRZrioqydNVQum5WvXd8JAIscbkrhfvZiRv3YCqjpPJN6T2
Sj4gIKhd1nXv1KX5VCBYaQ3JBuePyh+mjRcwmF6MiRza1ce8QoxabWEBiQfIkVXW6AQtE+96WZ1F
B/x5A7q3i8y1LDREWRfvJDbDgtvI0+Z7B34Y6SlVhley3wpODdKKdkBgQ8ryn+XCfox5qoJupYKP
ok/fz8yWH4NiiccH3AnFyM6dMNdqXieSiypV5sVzHCHzoj79TeuH0mmUaZWMwgDQzDwenqtXvglX
QnhxpyZhO91VFYjIkDh4/qvAgJwltO0sz+pnDqks6P246Htz552mz3FmWK0FvLVuGXgGBJlp9dL6
cCc9pHB5H5Y/3P28KgiOZbP/Qdn0V9d+fncAOQW+qBhMxaBAJDnF/+UuqTnURtBEriyIzrIvgQz5
9KudCvHxVpSTDPoFt2+PttoKVfjdu2XCDIuxzTUnWJTS+SXffkm9MvS+E8naw4cGebqiuw0AX36O
4E/jUCL6cJ7zqkCeOXR7OW4Ynueqn95qEZOVXsCeEtVfNzUv5FSmZdJQlIl/0vHZL7Hp1XgHLm+o
AR4+7rIeNIzZ+6TFYBCYnrWinlyv2dBPtVndX5qTawVg48dNXifjHDofYNe9JtHO9syU3ncAXtWM
Lzvk1G2ccW/OLtfAL/X7RNZNMoWCBJKTjWurptHBew6B8tqdf+OC0wWbq/hvwNcjgYY4rSsr1d1r
UF5oTs6PpCIYbRQQ8V+XrXQjOGDnsgCEl/u9hfbMN2mH+g4VMVA6V2okRII6d7YTVnNId9iHCXXc
OWZdyxv9OP1gmGB1n8xe89tGBCt4bS2nIEr1Xy+cHCnw4gNS01IlWJL5inIdVvw0+0ZOiye45lFO
5DcnEK7ZXSbcrCqPE557UYJsExWMcikqU88Lt9pakawgDQGhUt3UX7XFJu+8AniOsDYK/QSs0ir/
kGjk7K8e6FxA2NzHogxA3ZBe/S2bj3VwuUn9JtLZxsqZj96LxMz8BXdJBlRd9y9DQm81WUPygySv
9+JbjBKTSUL2hLluC76u8OKh09Fs4tEG8qtRY7OY5FKW9NJdfzoJJKtoJY/Ezht8L1H/hhi31qeK
EDG9wECT+eWcqMPqi7Uc2X/mYKyQAnIT5wRT8SI/ucd6av3RedDjDkf1CzFu5DXgX9heIH8oo99q
L0fOzuJR4jP1D8d00kyZM2CZN3hW1G3uzNxSH4vXdaC86fBh+kKb9ec4BDfvAWaGraVE+/3Uo2PW
UaMMfIuKkDhAgWYshxDbXMaGLtXo0xRqC947AWsHqJ+24kDBfPF92dxkBQxhgtbf5de0p0JXUd0X
PWYbbtS0Be+Job+DDf5TrY9k42OAB1uOZjvWCAVykkdcQE+n30lNlWh6bwxWYl6KNiqitdwNpeZt
ZN+D09Bbksz8Fqb10WH/HA8VeF+0XSd/BY6PV3/FdX6StRSCUdCZktjSm/yKBw3jk7rItw15OMtO
8VQtNld+K3IpykTELNsxhasZq7wnzfigM8a0QNRK3flsYew3Gi01M38r2ZgDCNjiuGJyreqjl7x8
uwxMhm6Tt3zHLOgeFKQJ9pamZNlLqZ/Hj9i1sNUHTfCnH0/BddhATb6ZBM2T+X5IYt2aVN2FWXPz
yWRhbezkRh2a+R+uKPEHcR4vi1EEnnv4Wu8DKoeg9tDRMzH5pFHH7zpFgxUtlBiP/6EZ32iI4s1M
hF/Cq2408UzljCpwVuaMRB6kHCi3UKuzIZzkBCXY4WKLzAux/b/v9IzoqfqYLP4nfvt1w0K8l7oB
jZFoPsiJ9Kf0xt2/+Rb6ofvuAg4mFRHpp/LyFTYtG1xgatcpvlTpSF4yCUR1h+RA2qk7MEVHDhUp
z6EXq7hVEAr+VBMrEzEa5W61O+lbcRG4HdRTsOCQz3BIn721cSvchtEqrn+sqId2rvm9VsumwfC3
j51v8s1q1skqwTPq+ArifgKgpdff5RLetomE4zy3zFhGxYglrujYf7uUMqhJV26chhTU8M1U1Htu
vEFrRf21exhskpZ+9q6OOoHFYePpYxr5NJQhlrIKSuYJlBumvALdRqsqGGRTHTYytSaa8EcMIvS1
tD7/INvzkfQ6Ixfmil1KcQxFMUZ2x9m894fIeWwIkbPLwRZgRPp3vTAazEyNxW94lr6tS08GEBtR
/TbU5ErSKj37L6+uE33m4DwBpaAZ7nTRQ/OlIqzIk2c1eIAQWQFyg2BmoZzWpEn8q6tjbIbuIyi1
ldBDhBkacFxkcOvkXDf0yOtKnIqRM2FQf9OKpw9IT2HaJMFwBUrVkm+l6AQ/ki6rLax0wXrm9+CE
JKx51VTt/3ziPdn7ff7Kq3M3QI12krUA64xv6YGGY/DshWklX/apx+UEzlmwUyPdxU8qmxkYCa7i
q9/C/RM6sPryTHk/u2lYwTuh+rLTJkMOz72UcpcFXs5+AKXXm16oJNFaDoiNU9kD7KUcI13mv36p
B7YtTB+TyQK6Bf192dBpb+sd0A6BfG547cRrM/OEowP1zT1tN/JT8uDwEJdr9KRTJU9pTwgMm+Nm
YrOafyi+OKp9DNYCMEs/PmRmXUO76zy7UbHLdjUuvel3A3GT14j3qjkHd88Re7AxMGrXRSMEZLmN
R87U9Gc4+9L2N+m/Zah+2S23tTM9b8xoT2ojSUzECXX5DcAzOAXkJkGoixHVvEKKQs7pG8Dwa2tb
q6O5/WHkJrAXJYlxsnYzw+eAZy5lCStAJDA5VKqsTG1XE82y90C0NDj9eGt4FEC/d6oTb81CgJy/
nNS7uzwswc49POInYmKIIQhd+5Z/C8J0qyCml+iuHaA7NxdUZiyMSbFdYOLgkZOwzz4AxR7Vf2/u
6acyok3tj8BkVOv7cSRyshyDIibNoNMaUkSdHQCj3RWieMELWCbJVs7+fBei4k+CZDX8LfzWP3eN
wxYa1P21NKZG8wJqOzulv3emACuGYFDQaF/I/zMTPCNqRs+Lg3vziyCYrTXT9gXM0eWhdpUKkvn/
McWNSuW9/BBHf00MFUh6uS5IIpBPJiLmlywbvzC0ivF4a78+BF16dLcKQ69N7G69azCzznSpwjdx
c7d5n80c2/WmAWKs2bPY3/4gMAzw/B0OTP7wAQb7lrzIl5cTTpk8CWG1yRq5VdMarWn9uCYsVzp7
l1pWnYJGU+NeqD9LvxhCzY7/gKXjNbkBrDL8p87k3nJ+byQWugLymQvgSXrmitmxFkmnAK0v6Kab
NkhYPtqHq4BbfU1Z4OHGBIbhnVX13iSHPXWGAEB3eGZfPdOGu392/PejLrMpvo38YnLc6V6Z2cXu
n3qjWwOMDxgFEDPHQxZ2DydaKCur1nfhsun7xIrE8TH2PCXFz8Ei68VxovpaZTuQYkqMK2q9d675
XEBAX0EHLNShcSPnIisBk460JHgwHBfeztoB2WIh3HTLNdIcnvV2NAJsOvfiDUqqqPpRZVGmNVV2
hbfLJlt3xnRKllM1LHflbgjxWCTc6vS1dGwlHe/UMAm8vC/TRx8ck6dJ29DXhwXao7UvwFSp95VX
xB8wWKmyY/0CJx6zHwlEpyYMzp66kAQQa/QMYClMUwaJoC1NcwseGZOsajEo6g/k+w+OWVj69GAB
m0G808cpz06iyrndjQxNwoqpn24Xgm8jlBzoo+WdoI+lQiOVC9T9CyoYTDuwOxwiFq/gto4FDOks
aCgkBnPZKm/pq6lKY9pDbUVbDNMlw2uhf6PnbpSZEy8FDIKjCHiOlgPgPhfTontvPNmKfLry/C97
rxDGuL7ao7WUU4wl2bcRgoYLpZ4nCWHCvJ9YOgWTiDYg1YAm6q5Rz8AcWP/A9FTh3LFJt8kI+XWH
5l8C3MYCvuJy7kMEJRt6CjEA9vJweLjW5lIhFgLTndcRVd0pmClYiSNSHKfHd2vBKnXG6yj1Rt5n
ZJG31W4W9Dc1TikSfSd+9LZ6672G78AxhzmUcK61V67bPNVEGc1I3YW8TPR75ODOId/FDJ7UNpMV
JzMdOA0Ikc1WHyIPhq1zUj5h8RZIiHt5WJGtXD4eePoFKO+FnufJbYkhwXmWG7w2NarKymUstQVK
i1eCmGzsUrnkRNbfDTRiwKFxFG/ILx/Nkbo1McK5ZgIdPWr9xJZA07HbVwgAu5bYrD6orPSiVG67
cu+7LroaAVfCykjlwiCUvtqP++D2ScV5CX35tW59EH+wBdgM6Igy6+PhigKJIUMkNx117YcvSR8k
voicVqe3fmHjMhkjhCLf1ZWdkUTCB8kddkWu5FJkv8cXe01UCX8JLUA2A9ccsJg4SJOSmDwXM+ax
M+ADh0cpvsQkZrTIjJdT7m/99Vljo8YoO0b7oDIZvLenCB6zIn0a6qaIz4mldRLjNE2Z6XhAtUs5
gmokEEwRfSfSqSGZV1Ktis8r5KbeRF69Cyiiuz0P79nyd+8c956shH2PXVGelJYAAg4022hjjSbA
qGpLl4iFwD/uSFzeWbIo7bAZeeey68CjmFgkI8i2tRFNCA3mON2xHGOqNEVq+DP4qyIU+cEMRFCu
b8cSgXJVhY1ZtYxkAGenF7Kjz7sk6QVNaSrUcc8mJC3jzGSaXDgDF6RYQQoCiFfKnLlhxbm+sbzG
rnJcfAlNm9u6IIiL1QlJolzbc1XzJh6X617Lnyxz+QM00Ygp8cRYD0CjEPCMugTVYfJN5znezn8t
qsO8zHDjyeUruPP2U+TnfJ1cR838s7z11BJZdd/f8I9HMIN4Keg7Akoo6/t6rk30S0GdBZcQ+c+V
HiuW3BASWDOfy+b+xvMNIxpCTNPnRtmhvKnymXzt45qZHAH5qAvfU0e2dWiOwRQxfAwTOQtVbj2c
hLZoF/koRzQxcyaOABt5CjgcVKQfh/KZGuo4zjUqMeHKGVJ72HYUGuF99gCKT9z8jz+BRdw2kDmY
T7/f+o32pWPW1PER1f+KcjVu3vja/AwSPoqCJ5IOPiqIgRSAuL+jqebFKP1rwOBB45qKnbWYKtM5
N6frCedMy02BosgjbdV2twRdMY9nbFFFqeiK+hh5iyn4m7XsYcXrYjd6Kf9Bv8XbPqoEsWiHH5kt
ZD984q4Am2l2bR/1LRMuSQDzGCvZ4Rzu7H5tM0Up4T08BfSSUfTOLOqKwwGvjw1Vat26YU8OC14/
XcYsS0x1rUaQ9/164SV+JQUpX9sssgH+EBeNJVkvCceq89M/n+ODqlD4JCdiZMgmBJxY9W2/qkan
RJ7GrwCljriU/iUIKi6XzaS2VxW0XQ63yewJkaR9Lb1WL4VrOSmD/Iy3X6Jdd/AfTX96Xt64ONwd
Y1EgfJCGL+gJKwD7Iv57e7NNexD28Olex/bwu24W/XOlFvGQ6SbO/4NBVn80mZOirGfQiQ1BrBRA
jZmYcX3S5gJxy3C0PwiWGlyGQ5YVd49oK8XbJd/FE5ZbdX6cZHhLaEbyrwdusEcH7awkXBwvZBDv
zKdi10kEGDodX+zd0RxyM5MUJ7+j7aWikaFHw3kurm4+pyT0tvQ2S7ZAapcPKFFY2d9Vh807+vuJ
sz5nXbcJDeiQMR025Xk/pk2zT0yymzdRDS/oL3Rh1oSJS/KjiEUL+7AExj80ZrF4Az7nApPRCnaV
rCRx9FwInMFf73CsITOwzl2gY2uSrYSEb2N42si417QLBFlHNMU959dUvgBvoMsXfvHHsgzQozg/
uScE+ZQZYfnUJg1crAfyC9wg3lcHVgLLOccQi5aD3abvYOrX+wAWPzXP/ko9trYIjszQzUroflAB
8tHy7fGmJFyrmuD7dc4mApXOADU1ayY556hiZFMlYc5QD35eHxzymMSh9YIZm+WzVh4/HvU3G2qX
CmSGlV4pNFggBdPO2lZUR+B/mMhqHpIYRJe6E6Lvqr1a6inkXKP13J8UP4OelBAP+ud3ubeuJv6u
puOFouVrFItHSUuYCvfBI/hLjYpgI0FzcLM/7okhcb399kH08NH1jgqWPXo2L6Sc7EIRA4dT7lNC
6Vj0V7b2lb2lnLYEA1M2OssoldXXI1T0alsqkW88l5QQoUjmUVzq1S//QYG3NCl5ATnpOYGiJhaa
hERyKlqg2N/JMjXq0myig+3V9v91VSyftY+8u7HLXNHY/ePnf7HFABx4oRH1EM0PsUGsyThZ6u39
ApIEsvE21IKljqRrwAWZOPnUO+qx5bCXUNPXnWE2ZwxKOxUEl4yzcE8kncsW0/exteUU1cJCwu8D
8OJMB2K5dSun0QGRhPzvuAWxOApIDxFldHJ+n9dNtw0lpeJkCILDWmgqVy3KgieKO6J6eZMF2+P9
PaVb24Jr1PDrXFTMALVq5XMR5V28EHwQAI9lKxGxgA89KLHCGzBj6FTQqljf267Y3svOJ1+anRTf
o+A+SaXv+w+gwZwQeycb6TRCqKAIgXprNhQtINyEM+ot+6Cl7gRWYwLV8zEkGwmB5vOuuVKwCkB/
I/kIAFCWIq371QdJ36eqr7hrvWALBygZpVz02TAaTGu78GQHeP83OEQJ3+miZa81no0XS7gy20Ok
FVEwBqAqbfPMJw22zYnqwshHYQA+7y7oBv2veNbwVHHiGJjjOT1jaLLHykPFevsM7Lu1RqY2I7kg
gV5eqHVDtgOAhU/bujIHKt89+Hr8qXJ6tbgDvXtMNfDMNsG5zt6DJfO3vN4jwnW7yjhIvGSGSohQ
cKL0VVS1JwkNLu2Zkdx/SLDfbiUTbPbsR+VVZ+aCh/tDcSSO3iCPlBCRCamAmPrEzRrxS7noSguz
ydwZRUMw1vGkWBs3i1z2YJaKLlGLvPnVwO1RDw58svD0PrngYxLiqNiQ5VQ3HxpdttCiSIHh59xf
8W41tYVV8NLSntxof/FP66hlGkOW608BinaSIiZIvpHX9Wspz0hjt/Gg3YTE5qd1RsHP/Ni8iqwF
Qnx4kJ1+q8stgPFikau67yZCox1bZ4f7lh3HPNKaiicu1LcM5z5PQJ3jrrxLkFj1Yl/MO0ewZN1A
z5l7WA+GghaPNgUvW6nOSlnOEq2yfr2Huzs1CLAtEbyF9UISNOlCgWTisa6ZxXFQ9pLi9lBZDRGs
mvdVmeczrU6Sr58IRnuAO9xzfJTER15xZjEPki++4aWTbjN5/V9SCb98skgYqSG1UrBPIyH9XAHx
RmZ5VxtrsVU/g0Cr2m4vrD0fwlebWKpiinPyVFMSE9o0bq517HPFWfmdgT//wQyGjI9emMLunmJ2
uTtPsDbo/zsYW0XTn6ERyQr757XQHfUv3+2r8UOFA9N3s5aeLBJ9u1XpJXv62ep5I2rNXLjmwaLR
qZu9JgS04lWM/t1S6dNzfTQq2X4TU/rCfBsdZZ+5EK7BScbcu9YbFc9l/vTmdWbLg7WD0Cnu79di
U0ey3ATlG47/37w8oICfjONGwOneiwmv1+faZXXgL+CF6NDgPqdM/zB/mNcC99XwHmCaBROM8klB
BfGuWNBWt7qv4PAMBnE+feKVJnaWkewAJel7Ev7Ms3aPDNrz22fUEvHwC9ivzEPFirZhPXQDQ5HJ
9NlTx68U3XvLJLOSMPxaE7nRR6krHu1ebc2JjHSwbs+WP1KPumNwBBSz/mH8matn0rV66QwS5dkS
pjATwPanhZWRwmf0gUHVRsNMP3zeU3mZGCqpkscWtD2Ggig77jp9SFPOWHAcc6moXwKYEHurMMx3
XOjwEco6WhtWsGnDB9AahLw8Espk2gyYtrPCNcoRLNyE7zXIOm3iFf/JV+6/pY5QsvjraZaj3yMV
BfCImHQKCZM8W3huNHe5j3hTNwMLbOheS0fAkY7GYKpVvUs+lRCJ8AdiRfS9WsaQ7ff/2qetyAb+
plgZAP+mLhMfZaEFBgWJIpsxsBTdN3e9N0EIYU7Xlz9polCxcijOKa3C+ttCBWT1uP1V1jhOFxwq
P6GgYDztCvHwV09uy1qC0rsdFGUoF2Qj4PqQ7w07XOmYyIO2AklLLEUaeNQsrylImcmaZ734hq0a
39UbMdITXKO3MVaxglzpI8xHe+K40YIwjXiOg7lDJ50lCR2tIqMCY9sKklCWbSSoIweDMHncoLqZ
bYYlzrGV5ITvAtGPRD3cVQPT6rHbJu47VX23/HP0m3yGqvPV06ftuTmk/FNO+CoWCFUtPVpBb0sS
VwnYlW2eU7qjCyWtgKZglTvrlyyJ31gD0sAXsCLRo/ZLscBbTl757XuzcmIDY+M0bcI8BgEbPCOr
jlRfz9OQgUjodUXcdrRsWlEt65Fyj4tShsj0qxEy9TXAb9ro+L6+3+O+pPkZ6dSUpTrla/chLj4I
2QuZXrl4/4NBwVWgwN8A7QGJ6Jmn5dPj8MNGnyXruifuhoGmxEnXeHPUB7xLiuBfIrc5+qFu6WN7
D9yIEZRhyRUtc3HNE22h29Q/HzpqoY2+rNnbCHjrbtX5zTAPuRMl51/SyJC6ozZRbgB7B42FtZx7
6HGKqeKCUEwavlXI5r5EmISfcF2CYgHm3Pn71UqYfD5sffe2ugrahh/Lmf7roHqnPyheYyEdKUID
UJIHGRLKwWFWrjnEI7yjMAloDGThWRJkmvckiedA0mmhn1U1auMBJnYqsLe223PEkyFK0/311rGn
rF2/Eau4AgNyCO20ZPe+7fsPy7EYiPxppnKz326LeKIvBEoEM1wpjH2QjCJokWt7fY9OXSz60C4Z
KlVBSW+5H7ZVgGlRHF0HXPoEaWALzWpVk8v7dlwcPngkoEwqUXGJOrXI4S41NZoUTC+hKuYxM4+s
oxeQ37UsI5d8vTc0EE1n4rgGU6Z+w4Tyngn5ayje020sNs2gsLjFEBOjpe9TP4JneEUBLaE4OBUO
CHOHuhw76L2ux0abpUNZnM/8cftjLjnEKmHkQJCdqXbOxUkQIXSOvUDCRYHhBQnRaySt+5MOR9hH
VNnqEphReZAZZ9djjpRtkujtL7RU+C3FbJPinsAc37Hrrhp/hJg7f8cQk5EQHLKMFIGEHPqyJRwT
H494sfkfRkFE+0qK4kQRmP7CIP5Wm4J2vfjB0ut1om5h2ArbXnyCZqd437z02DAQIqVO9tyNxlBj
e0nV0UedH0C+23bS+YPE9E95BjPOnHzypzhVY7k4hP6oiL4/65NE9EDO58ZCr+Tn6DsCU5S53uJO
ei1SizdwsfHDZQZbUMGuP91hwkclO1K9tOiOnNvcqYhI67eSVHcv4cjNv+uAaU6+NE5VRc+0sVo2
Yyzj0qiu36TCVX8zO+jHPMbI2TkLc29ELPqVK00WsXyKwl/uN3pTMckfZ6PDKnqS3lpjYGqQdCnv
glQobpEOIBihvBzoS4ca96FLyv/gTCz8Jkk1E2CfVq6GUfbi+6hRNVcznhnrXlxlFCE/g/KsJLjC
1Y905nY1lF3zPbLWNGXSV6pb8YihgZzThbi5csO1HjmN41jlpOHnltkODcZP2ZNeVt5eOTMDhDgb
svrPSfCofxb2YYLtJPSNwkaPGJ/2RhlsRqijYi5atnQUy1DhJ1GnZOe++Z36ilLRMsxKy7+Ec/CI
vKFKNFQ7MncF4iSc2gr60OoxulfHaAYHdY8k26LeoNmklDMxIQmRLRRg7fUHdUGgfDlqCDLx7t3A
MByirYZ99r/o58sn3AybQ2QiG/oaB3yvKi3DmTs4UkpGSh0W9EjjfDx0Jud6b3lB0tz0gZ9UMN79
oot49LpIscS61NL45aE80EZY9Y6vM30/lyPrLhr+s+14ezJsm4RWKwmZKcU/bE7hXVhbG/kpuGPk
PbrjP2ZIHcYsYqL8bRnQ52K/4Fx58DK8tUhHJ0Ik0XMZLWb09Iq+qKPbZI3FdHZCffIDFOQ0cJU7
hJ5qDATkSpdrmBQ2tH7CnKhEfuMVRp4IhTYrKfkt3t57j32H7+1b1Widzm5X/be6sOKg8ESeyoRF
Z+9s/sAvolWq8jUBKMS4vpXQi6mNV2moMUB53NXCTrIKCbguOwcAP4OnSqi1ZQUsnkPztwFPs0tk
Z4RpZVf0F+NbuNH7OveDz9rd0+hRyFtODTT9x0ROfuDX6Sg8wbSFagmFchKvVRs9Znumetsy9yNO
7QiTVVEShOjppD6g83UDOkJcEcGvjaJMX7LDWwMl7kxxglpWk0MO2Zsk0a/L3ZQ7SU9OcNMtJQRE
8UcV97PINrUXZFTIAihx5VxqQIotowASCE6bC8SJ155O5OX84ju22n07CLvhd9TS9APv7I/otL0P
1+95jQ+0OZflEiVS33xoqpGuHaiCUatCbaO5MnjcBI4TF912anHejySDcMXfw8sa8ODCdbw0v1aV
QBkWRNmJXRMiNBKkFwhZkzQxqbQW4APJihOGW67t02EsZSTt9VyYqE48sUpjhT4xs5MEhuvNEkgN
ik+Rj5ayS2Po+Wh3pDUq75nY3AYwR6blus+AtPC7kk2e6+cd8d220lgHF7o7NySyIKtX66RWm9n/
g2u/MM2D0PfsJZTuni5qD3xmCEF7aWO7aOwCjHxMywAhoit9IosdcfiyiGGT5kvKHQIHA7hAcKyT
xrjxmwpwF9fOz4a58Vg9skoED8PvR3h377gIaacsOqrU7aTpe+jFBeuk4z8S7K+Bv8HLkPoTWYll
y4ydkehoqYyTl/qzdFkkZdlg81M/l79mRz6gzbABIe2spFZxAP077Rj4nMOOFEQRqNzUdU8/H25v
wC4aLvFHsfwSiRT94ZN/8FChVdmKBppfTP9S6n1YkUYDflRwrz+ztAXBbfpkhBg0o7g9d8MFZXj+
6+ndD+qTVUeWg4Nisf2bKpaWIGae5n7zfWQoXYQN7fn4BcJA46kcifUEQPuy/Xmv/ZlkXxsOGZ3M
XZzv8l4emMNQKdconfWByUXa1jg1EvNT2OWdO5RFj7c8wzBEcuiv1A6txEuKrKxxu442O4SIPY1v
Gu8Zp91Tbm7Dejlyue0lhaFLF8g+Af3E8osW6JIbBCzVNayaOUESa44t0I+G/DZgk2fesAx3TG+z
Jw/FiVGdR7Q+bFpaBpbTiNxySBQtKlfRa0tsnIgek1UDEyXoBt9v+9nwN44iQ+BnLoIuhh3Tz8DX
JyhElv2Ru1HVIhDP9DppBXCIVk8L35WXZFW6xgdfSAAgCXMuBXSYnbDPAkDA66wE/mxOPYRMJUM2
ie0uA6udmllyY79QaJXsFYc48f4k9kXNgcGDM+dEqwT0+0YPcQAt/AMnzoZtv/MYZnLD06TKklxu
VNLpY8Gkd90cz1l4vufyQmFgcm4an18x8sypit4HmG0U/pDQqhGZDEUzFaSAVsMPQ4eFOynhlOWr
TO9afWeULYD7mdfD82SQovcBl74ECmJnfQUAKyTrWLrA3ns2SsUcsQVnTeNOnAdoEtXmTABFJuY9
RuoutQjfy3y7VLcErj/AoAJ6lqCFID75PGZhz+8jxKDhH4crtWEhua3hXM9WHFl1lme1NE4tRh8O
voPW83mXYG2hOgN3wcov4PyDurqHS1FvKGqb2y/DxVDKQ6rgjkpVgkSxflL+vg6JM7PxPoWXNL4X
MuBPbS4dU9A4McMrcojVyftkMafKz4WvPP3OsZXJZLnHBlX7E8TboMMvmydonHL4r+Kh2sysC4YX
dDCJNAoBUQppC395j2l1mswKVWpel84eXlcHV4T91aIiU8QEuv/Ozt9ecOfHz6ZCcedH1X1Cf9Rz
MeGznTxq13+B2CdRovkDP9VxMP5UmpsG1CroV89tu9wQImKa0z0Ws+sM6NqWCHNj2bDVcXPjgqu5
07OBqB2oKNPno98EHZhuzY/7XwsvOu3FttTuz7DhBRL71WFGxywssJz1EkDAT4Kvg0/j04bv9FKi
SSJ9w44rylnNCz6Gx4YHVeTexNiGCQGrYRkafBpZtTevSOE8rO9tKY42ZVTpFgyh0KOc7Y8wMvcH
R9zGCzTHJ3XEM0L22fXGm9joyPF50us+dmB57oLACJiJdJJQohlnnWvKHh6vbfYBG7XjMI30M2Lk
VXQtwTSYyt0zKN97VWxr3AZly7cSbso1/tPelMgdRuBQls6jpjW51VMS5UStp/kodv2Ya4FAht6f
e2Jh27pw10PGiojTwN1oDIfAC3Q7kbxS021FldqWR0THnUk7a8kdQAk0iiBWwqfANlf1ff+9VRYp
kONM2mnPO7b47JrkNrjYWtXVTTowaNQ4/ZUcS6a2wDJBO/qiEH6dJTiaYW5A46EdKN6XNbN+sVe5
iFVSDrz4ibMINsWdNs0qck1qC0kFYWeZT+XoDyVe7tKu3iWydNxgmmp+9sjdzib59DyJknuGeVIm
9JPi/WoNVkF+pP4HdQ6Aov2dveMPLliQLyZGbird0WvyGHjfsYvLtNXtT8pWtTFbIpeBivtGmgs0
0xCqF2Mi+eKSrDs72eIRRTGYwzvP5RysOZ9dh33dc2Vx145M6T80liyMFtyBnPtGZRdPL5Hbooh5
nKA0LSQDliJadVK3HJVXb0/sUiW2dgO92VOH4WeYWJNUPzL1z4dMz242qPok7ZckTiFHT9xHh/Tk
juoZPp4Ca1MJesfd3qMt8VDVQnqKzk4QCy4YuqiGd7lhtZ3eeehri0izJsxsR++AF7X/4d8MAvi9
SgFvDQQ92r9dBC/9i0ReDQ+i55srmSYyPyHHzz+uIWNS5mH1qN9Dg1XMFBvO1MWQ6IFDio+iQOOc
1Lc72XfqHJBB1ik+ym37DcWlBfMTgUfvEr+euuUjK5GHhPWVWTph3Oz7bp11rcZLuES1NidF3VL5
uH1Lvl//Kg1urihQ/SHm6VuFK0IhQ92E9UhvRxOhaSXIiBnzNbf25zHD5yUYJhEZATosXj/8fxEN
TwvWoWaN4CjQjau1c8OiqKRDVlFg/a1tgE+r45eA1WW0X2WGo3duIGfTtdHA3i6I1ehusYEMjRDc
ehFlWj/0i0YEdkfPwH5ryiCctdzd7aubGPM5dCD8H7ZOGzneMaK2neoN4Zhsz/aL5aeM9wWu6ij6
G+LahfNr9/3I0f6AMXwWZ/D2xPJHhoKb71NEmunTurYWVXgfcza5F88B0F9gIhq8YUb75B0NxFFz
R9UTpsOKLQGFC/LyiEv7K2h/W2UDQMrO2mMekRvMCxNyrdPWCY6oFAuiqBAMnXs4u0koimm2r7q2
/Kjp86gS9Y7zo1mNnaP32WSJ2XmuBpDL4cAFxssX7PsB4ktTDdg0uI4CGHbIoWAH33jGHEJZmeb8
CmCQLMsbnWM8Wi20BXg2YMMkmgJGHahTQnLhE7bgLdmKYl+mTZxG62/6OJNzUYHXwEDIGYHd89H0
7XhPUCyGB2zE57BM8eBb0gHwgPll88DFI/lcEJuW1HKgI1ADTKM1JZna4qJ763wDmLDsnXUOmjLY
UQp1oougSKTO4rjzkVlxnVLwNzliG2P1Vmf0XdIT5oRrGlypTPJnzf1AavThrfLfdB9tNG+QBEJI
rkwTYeYq23Eo1TsbVvNW48SXDkRjIE7ZDZouE0K6lLV/77VKytNv2UKPd7V0J3ePdySL0m1hmU5T
av4uPyAfDd7ySFsstTW+eXcVeVZu/HLWdn0v5Slh59g+yBxooqc7vBs6T+aFtlwu2ckQGQU3aaBa
K9ulkhl+QVzDw/NQyyfmNZLsmH28mwg2Gn2fyuaJqhXrdh4JeQvenSymBP/OkEVlv+hCLIwrNGwx
VSOeKcesGM6jc+c6A7Be54oUkXstscf7dF6yX2ASTaPgjhJqJZLIOqhngWqr7JW2dkxDAyRAwUkD
WUATF6iMDWbZ3T8ecA218iR6G5P5lStkUhv8wcnggaqWWD50+xvj5EJi6wLHMuHq4KuPw0E22jOz
B8dPAG1DOkCIHqbFfqYnZLC1jR3AL0zwCplTC/FfdHkx2kIOs/yStLylM6n/i6Val3hrHz/u4pt1
LFqhHCTh8/pJrQB8yDxENNcyFbZe8V64Lxc86ihDe28LVs0H1KzexohuTbRtcRcJp8WfwueY5YIG
nLwmoDLbn8xUtT9SWl5btTHaqa97kHRe7dl2YL51GaaGN10ccVAZuh5RmpZmMii36TIvtATIovD3
ee4wloFVFuM++h1fWErFNAZTyjOwJsgjlSGq5zvDOi8YrIeS1c+QmU1gnEBq7cY6Znm26NkMhniQ
0/eefDGeKrxIMcxQvbNg1I+uPJlNm3nT6DSb77lXCEOduLdVJChh/+lbsfLgvQ2eyrqk9HxDC/Wb
o1Z3K9Jm5kkjhAf0oHssU/bKvUO47tCmkqphmrc6niPIHJXC+XebBHgRZgyBxLZufRn2w66iNVCA
z8gh0m8O+j3GzoU1cwG0So+rYLU85JElUgTRABCPWVJ2BOou2LSpIh7crt1KYSX0IWK6C6EWoShO
zGbM3RuCb7I71Vfaw8hgH+Fkw0Gyy/MFX77uknn//Qn0SKIEPJ5/b0LTVZ6OF2zmQN7XDDR2Yq6/
d2ENUZFg210jMgYZhlqF4m4A0sAAUEKeGXGhVcDIqwRtILVCcHa0V0MpAIy+TInX7RLuTe3RClyi
5YoBmQc0A7jaX1S2/mMoZupIyv4SLkxeN3A+T0gHA5uaNKYd+0dmjrhsX2HGmrdJb0UwhMDGsXPq
cWfbtXCItb2H/5aD5KlFfV8ek0zLeh+fLtOK/WFW0x0zxc7qzIVbmBRJev64nLzIp1jvMmDr+m6L
jDz8i4ffcP6aQWvL9q9WubS+zzUUSf9zEKwfi2sbh0ngax/ej1CrP8WlEPMT96mYuawVObVGkZuL
pBtPOCtu/jcVwPXij5vXVt+6PmZIrKBLl4jSMP3A0DH7ElOaYdfgAsZosb93vLj/ZVSPB5u8GSCq
LjHOLWaCxfYawPaZjTV9MqBjOmQa988Awcs+ZnW5ho8pc3CmU2sCOfRbghI8HV51JLRwiBNw4x/2
nbNRSa49tDVT6jgxSj42fAja3/UUbOpZcjI3YSwvop6GRCbjBcGL8EbjMLgglkBHCbnumJGC2h4t
CBHrj2is+vmX23JwZTRj3IhJpQmDks8q5eUjVzB6Zqs0j9dY7+2aMH7IEZ+nVtnhRpLKrXNbyqQ4
Uw8jaTN/bIiwmuCTdh1RVTZfe0T7aGtIulcTRLragLac0d9J5obV29Gh0dtnuGYQgdeRIT506O61
ZdWd/EvxYwbwzFYpIatg03XvZgtanwgZZi/rifzrvTzP1nEv8HbgLXqfsLGfLoFHsgOWCXbfroey
jtOxXmUeKh++USEUreLj71XOi1s1oi7+6CFpQTVqu+Z+xVmE9QpOgyYN4ry53MNaktQVYhmjfN7L
VHq0M8h4WNAifzHAE+qeRC1B79BqwdWNgicP9SslqmzZkbLm+/tqw7U9NWNZDw1Hb0txOPmZUcxx
kghOYt7SImktWNCCzyYI2e9Ip6eClCOds+0bFLSJpnrurYbF/B+uIX+idYwYgnUXS/V+brB110HP
WpKmZ8jliSS6gQonWVjmcR4keJiwlY8oWTDi0/pTwqa3k3npdGuHqpiWmSH2UWgiJeQg+AvjgK4Y
bcLIVk/nWfvcyOw5lrH0QS1OnCoZhumx085IaJMqXQuJOMEsN+3HsejBTGNfyvTAM+/OvZmH5Azh
6ysjDeTRgscO+OBZA8z7JCirPHbpnMu8jm45a+380ltdUpTOtBPeNccQZnY7OeTTnZNxnj3L5KvH
6iVjWKac82i0hA1doOkz1JQTYTZveVLplnoPPncqLqwCPtWYSndWKN63IvCpshoRA5x9N+0GEOKS
NX2lMbW9qsHH1pnB6GOSYOx5f/djBP7eT8YqjDtR3sh5nzNcgP4/CPe9NeW5Nl1fDWC+UYs3B3bC
DiPjwt9KvPsOTBjJVwK70V96mtQreQi4v4vlBGqbl/owaqMAJw0y8GfbruN9hZ7bnucE06ge1wSW
tupPHjc62Toz22x+upS7Mj7Ikdp9PoFfyaqt0CoWPpzuLozotpHHZsaufDn7eGrHeQltfy8pDCQl
ew9i8Yk4EfFv8rlcF1bD3EnTLRYSELZAuWdAsg6gbdKqYJW9AxL/xN10FFTJZB5gRFo6gvtQseH0
QfiO/1lMnoGvMtBWlnerzgsdLeNpKpV8czNo9ygsU/pW0FGbfgwwkzPa9gmE6S2k8FUQ1oi8Miu3
UE4lr4V8rg5nDSydxWX7rHR/N6D3czwRRHRZ3jRKrnrrS28Wb9D892aIfvBJ6Ixhu2GnXZqTkm9X
nzLpyIUrmFCABqMZD4JOfXPoCY6g/w8T9FLq3a0v+a4fDO9R6QxNEv6gXtEHO3HF8vB9dvPFWhrN
vZwifC7zQ7Vl3tzA2bJ7hsYGW0CJlY767nAlxb55jnCUZhw+9/BPuL+qNEnYXVUIcxKz7wD4jnVA
JafU3ddmoxOyvrcTPTD9j+4X8C18SChQh4MarQVFXDIOsZOpSxS5g0OZrKgGwG6/W0fBfoTGZoDA
Jk7PxhMU7dpz/Xy8Da8CfRG3GiGD6TtqNXQoV//k2Gjf1kYt1KV7dvdbw6D+fG/MT0/yPHrL6vSV
kr+Y7kaF/Dumewe2RgQVBf5efYIaLvpcS/UkfC1EawpeRH7Lsz88duqauWYGCufKpNroZRf6DvcW
Ou/U9Tha9bwYBEqFBiN+6RbabB/hG3Kk4G4kJO3Coob5rrJHgeROS/4jMFHgSELGHYeYMK6Nvze8
q+/b+DCvL5yNdApF0kg1omafpSBgEz5aJ1bevvmMMEPCJaO77o+dltERmnDhZwD1aPiAAJlhIbg2
/dCGKBJ6hsmA5MdPj1KIjfFPTyV81w70LWWjCtzQ51pwpdxrEW+yPafCLOuFdJwRz2KDZtk2DJss
OpGL2Qj7FUnNwu6uHzoXKxQo8wNUKm3HmHpPx/X5suPf6iJqCTZSvsqjoVDgsqV94WKfQn+JIdbX
2WzR15PSoxpImDyHPW5WpjU/QvONSC0T0CcFH9VVCiVK5srgV9pKNNnRO5c6WnsIkfOO3pHE8c+W
kFUeU04IfM46qY6B7L6r7EjALkbzm8kJIkpjl+2bSw7D7tS/P9tX8KmthAUGskt98SvnNBNXZJMA
UAOPLw/2QYXrxfNXHtnLgdgJdy20xquA/ob0OMoMOAkSbME4k6ipvy6eRuWRtbdmjkqPHIg/vlNY
K7zV7q4JN3wvAvemI+VHpZBtrT+1jOLO5s4tpEIHhn9MnCECt75kziCpp2mAnd5RmdcF7k8p7ava
yQ0LUPERxdgGmBNbF7HkNGtHAGzYfLghRPJEF7nEBM1dGIIaFbGHe1xTjqNOTyZckiNd1C6aXR1M
GCsLKbAuYXth86aKi2fGm1ChdW6UuKFqKWy8E4C25Gc0iL+izvPOpRaIy3mRwFnEPxn0Lz4DesAD
zwgbyX1QSw2WQLoKntIwUCZbtlgZ1AsH6ekAZaPbsL88WYmMknUcncV4rr9NL2qDMRlhacLUZnlR
674tFMMSCpomrUFsGBVG3LvR9x0xQ45Wv4v/Xq67igW03yLz80OGfxUb8VljPNFpD+80ENbwwL9v
h6dvdbUbuAiPGffneVvcecbW7Zr2FpjI80BaXq/TTSixVIPKeiGMvNAKCetFWRax/7HQoswZGXD9
f0gbeQoX22AE5tqh8cmrYmFzV7AiGsJV0Rp6X3Wi83fZF4k72zG7cJbdDx9V+IDnMdgLrjeV2XAw
uLiI4+BzEuN33DBA9X3fRjowLA2mcxH1p50RLf6xGnEnBR71QVISsbR9FwGQpISpNlNpWSuOMk/W
SUrWDX9i/yJhKHcCOEZaXZYNRPBm+QQ2nPitPt4YlWTGYDdLiT88AqZqL35C8uWlJ3eLQZfz8YM2
hQBIgtW/g5EUJEVG5C80/KIbgAmywPwg2owxJ0KEjW/nARdJnxDzeuAQXna5sycX118go+UUxBkH
qAJ+Wae1YLCSsmGEy0VN7qnUAEZwbI2onMo/QaLdSKuN0Qf2Tb5kk/7U5GZE+U/XPLelUTuh4MQO
OaormKIFhmPAi6qm2ZeCk2TXPU5mTJ4OOWTKTqC6C4RxSbcRUrT/shVG/VoJxuMfqwFpGGqeRjYk
217wXyfsMF6G2x4Z/WLGhKeuszBL3x2KvxdU/Q1evAzK6k9wNomhEnsZRBVAPS5wbZdSk+c33/5l
A4G7d2e8KuTF22rS6pJUTBZD7JTFYQ85O5zZxEFFFeBtX3XIfF07+LpxsXItQSrLGP0Edp7Xf76q
fy2qJfSr+hwvQmGdUJ4t2OR0v0MghrcEfgZn6LdicZlD10E9wHG+rmG65DF7yOGr/X+H84wJSCzA
2PgbpTiAcZmJRY3zPnW76GJIbDoR84LTx6NjREtzOJunJ51KLAB3JgDXtqquMYKBYC1KC1TYMXWR
IikeoStMD9JLgFmmlftNlegfJypHbyFYPRrCPrZS9vmntjh0O7vPgmSsFGgaCwPGzZfTLfZdNlS1
BU92X4R4D13nsT1dF06DiS0aEnuIEc79yY0sRrfnhlAzbeDG2vqxLhNTm8DmRfJLquul8J75sn9v
Q7xuvaophsTLU579zzSLzevUW5wU+dkSBIkSXRCHtR8CSc/H5OL2CR0B0KavhQwDmBETGHkszSsU
Zdyy/eLysBimOgO2vSNzcd8L881IoyiYxaWYtiiEr3CaCl8jM2zBr6cC2xkL16w3lKMlRHWVxLaG
Xp5S+fowc1UWh7PCeqJK35WndSgDG3D1/lfPrSH2QELkVXv0TBsHSE1DGZMkgwwRtd+MqKjfwMcz
mxVn8Vxo6k7YazsxYqFjSn3NOYIsR06ehbUya4HBHmcAbX1sOHnJvvvqaTkf6mdilsuv9RnNyYzg
vYPv/wlOCD0niVD6/lbjuQ1M8bkEtp9QrKLxomy+uEyUfArHBsAYzGPgqVLpL3S5KfYz5DdVGWhw
g4q4xIMGad6yWRgYt5T2C2RVgRVAgDa7Bl1v3ldaIHsUFigDXdbL6BzBjQR9/FASWwSUxZ2cSm4a
NQOQP3vZHFJkPHf6gDVdRX5URXamEHjynTnpOpE/da5EUsU2QX+xR2swVhX6FCjRjznE6Qs3OrSO
bRxZEsp5tSCXGlpSE2w4AyFChKEHi9RmS+BNYE+vzDP1fwVxpjGMZQeexm9tbq4EAWUXWmWffCk6
4sZio9OWmFukpSX2xLFb5GQQvjcUWy1kZzGPwg9WSOY5xuRfSAGCKyTfgWBtb/daOo78LJVcFC5u
k5H8CwWyUwbWhn2sGsuFIs1chs7/R+LXSZrR27ctJ62jl2x7LxBPb3Hj40Eq5e7nJAQ9JrRFb65o
IWLmpzCaejB1+QRLoHDeAAt9RK7lL9+oVBqqgpq7oTzcapepoxLvZ5g+OibGnGGHt4+fqSaLmH71
glpM0zuEUhAcmeOV5APqNLq+KXGHuAQTRzRbj287HYp4VK5RbabxUVlDnRbr104/3STdoX8Uf7JS
zNZz1owpXc9Kh3wFxtHFeBKn3NgFC65QnODW9Mb9cLIjjeGucUYzag1Enf6cCfZo38GbcMH+mDO9
YSFjZornmsat4Sn3N9qwMxAYg4zrFeadAj7ssYoZWeeqQ7VRF1wMocslom1E4c0rHzg3tk87qWdC
KVhLke7WYj0UalJbuftV7902L574njHkbueY0u69Y3jSd7gDfQxOSoyJPUmwYluetIvvUx7O2ltE
gzXNcnrf2fvHywVdDotCZZONfSaiAJGE0ETppGjV4DmPo6IWp382ZxFNa+89+oG6aelSR955n0Bh
D/mJkCAzP4cl0AiRCnFXGERLUGip15lXBuLa5fsseAo7aGJpTXl5X7owkmunG2sg6Ylu7lq7GoOc
z0AYffRsSMPlSCmatRZzy2e9RQGzkWGRFqajeQ41NjZ/GhaU8QISQMefdElzsg7PxKKsjJrR7vmq
5oMMO+RAJfk+VY37ES9CwAETdYrh8qphB+vUBtGajY1cyhWBrHg/hELqXpTjxXFHu5C16C81kei6
8tm6kJk5/O1HGljJipA1dzB0CROnazqeyYVmcL/rnuI1CHA8tW47MAc8h5fE6DpiJxYfF7V4OdHu
JzlgaFz7nvooA6YoMxgkKWBn/V2QfEpnXb80BlcBPN2uBvBqbAmabB1+lQX06mZwsDmBHJtCKbuA
ZTxuK+3mdTlzXf1sN1i5SZO0tOLEQQS9qbJvRXII1nIji3kqFkmDAHvknNKmz3rxT/DJOBSjeDHq
NN+3G1bu3bUUkmAgrGZlaCn1G1duPK2VgX8PzdYvR5MXy6C/mJaCG3PUhoY1GKfurp7GRdZdq7vR
jvzVnodbWHFQ7pJZ53aut06BrMBSKvp/m8Jakx5ni1mU+0KE03J37yfXnwihVBO1yeqzMPj0ijQP
6JXenudJDBCJYhb10VWNGz9mtgpOHyiljqt1sZb0+2zppRORxxMOZdzr7uxXnAIPV8vMMbHBBzSG
bm4xFYV68Sj2g6N/777bNtjebKk6qVrEwttiH+eVMAUN47XqiQ8McEnYuP76TViqeMk+pff1Jl6Y
H45R3HXdFvLU1WUNWukhVb4f9DeWXzVaAB8hq+B32y5AFh7SjaBODVfF7Cku43Rl4TPz3LYc3NB0
Wnxe2oCm3xzdk5wuejSdWu4AcaUzI/cimqiZ9/QJWHMZ94rl0jfm4CivYO7ai1k8Ux2ZKK43+fcf
GnX1mrpKDQ0xpYTqrH9t0Y9dkK5IMN3TivT8zDbYTFK54huvqYo376Ro+gM6qvZYrmrhPUaTO3Rd
w4vphWKT3+jomoknO3x1j692N03jrx8NDCq6gTU8IDvbyrmuBeaOot6/yto5pfwi9gAKm1bPGHE5
NwnWWhqYGnyHuJPmWCKu29oZ8tc53VZUl1fi358DSlRLgPSIBmoByW9bfa2/lJuQ5gOYC3hteExs
nNZOflbfm1WgkdPhQnmQW1UQrhm3pHLlwCQcL0Xfc3slq7SFXCLvvc4IkKfP4jl6dLEffwnp3dNL
nGCUSRxJoSk2aT3XvnWRoViYZ+aPWfVxkj4b7oZFjled/pj7JlDdUFUOpkfaKkqAS2EYox5stjaD
JTRMZpKhsCfmsmVFA3U/u3WuXmRI9xZdCCQMbdw6T/V5ibT5J6jIhmTgAF/eMn6CJMtkkn1KJqWV
5qJ9ysoq8bedOkpElrMr7YhnpuSp0q1tFg2AB2Ypod+ftiZj1hHr43UsBJDrbUV+vcSBVPG4+lPb
nTAxdAesh81Ym12lM9tt4iWEZuNVwMQK+nZOErXvJYzA6b/pFE5DUI4gvxLUpi4OM8EtV1SkF60g
7x8YDs4ucXRxThjER41me2BEFIzI+CQ6yX9F2nw+egnK6rqvpEbcttD9DvU/w9oU0/gdmSv18n29
izz8ASufyuWXmmVCeMj0D/DdQvnuaSHLeKqakuYNwccfl3IuUebYSv+BYiD9ga0hB9OOJjjwQD81
TVXU59ZeSKk/70pHbQHQFde3X1y45BFcbAueypWXTRzVK7WwB7FOWnyY4TjIuloP82emSXzBZkQU
OTotTdMS4BhfdG792ekkhumd4skeDlJYK5T839euTyvKgftfACitcfAnHfw+ulEjxkZ1lp1kdRRW
MdhaOeBakvksHZHfODZaJpR5YFKLQvwi7oT6ZdUMWYA+YQh2itKwnart/m1V14wAe0DUh1RtkaRr
yVbfmFlUJIvGjJn3Qtmd99n+pF9/GN63RsVBcB7A1xR88vHtmSwHNN2H+nhHmHchMzuMbzuehEz+
DacaV4c1NHZtBZxVbkvEBU7n3OEI9UtgsoNUI0b/40307hlUkbRNOkf7Mw10S0iUjlffw+3J7jzj
VpvbszO6LA4G1SXgAQnr91N34RZ7ftyfSdM/1qAtZ4gpbcKK3WZZLfYROTLA9OaF6NlwE+D6rnq8
PdE9sxPggnKa9O7FNeqlaUQsdU5VcPv77SGF3ahm8uitZUk2igPTIsyvsZlbCMFxeci907g3tHGn
24n8kNuTl0VXJsBDIgSCdW7Fosq0TZFlkg/urxF94Ft+JhCBOsFAIzjrmH+EV3RgNHJF9HRlnexC
3e0nMAyoTm+aChEt3wSEWYKYQGnarRAebDfk+hmgwJKdGhidkDDvu0sUHTw9nlCmQLQdxoaJgGg6
ZILJhcPS5HWFcuDP7Hu1ie8pP6TWJEekn/xhYWHzbfpbsccy86jsK5mrZE91LboEAMFQDPXHoFc5
PChVvg4X7sDzOYjVseGYC7qfKceByCKHLJsXOyezRVdrtOS8VHTrwRc2A3NLSqRK6cY7jzbX2g6M
K4eIYEmb2C4wHXjzwIAsdcUa0Pe9RTOViZWA3bvPw6ZCaIe71EP0Engej2VZg4BgSExEQfaVkvbC
m+9syO8Ym0toNiEeGm8BjiS4ict6jPApmMpSk+dTRpODJsyt/sV5fipUAmy2YGXrm4ohPOCJw4gh
dkQRnhaiCOdIe0u6JHjcfsPTDgceMC/7w5ox+3Yh8PFHHisS0FkpBlKGK1mzQ2gY2C67lhFpm08p
gZuhGwoITwQEcTFeDVhUeeyWlYIbqopN9CHumZ8mAT5lcpxID6O1/OQuuQk+W7rkLFrJG0Hp+TOS
BxearD5ACXvOFDpatId3F/IAff8eANFG4wDz8b9JzONfoAGxytN0l8MFR5qKaSW1w2cKaf7rtI9U
q/22etn7OWdR+D7FZTv6OQarzrMmYaq0q2xuwz127JrqpuwcPzUC2dG/MJU/CGH7LfCYOMUfI0jA
jyKOJREDD28v4IJHriMRpJ0tiFtM67Ahy/VFTl/pC8hhbgY++8flC/DaBm3dMQwSVfSzMHiDcz/y
LweTV8UtjJLoEnXAJQjPd+B8Z0EXzzwWCaAY6SvwTn9U+86lbUNizKZFNsPA9120uCIVKoM3n2mH
liHLifur0EB1GOsgiy42Fq0eVHPp5efkzfG5/NveRnjW61oCUY1qv6i/m1AnbecO1hZFXYIOq9i8
2Ngn1kNwEhbZB8gOpuh3JVlijItkmYCxqB7zBPux9a1v+vBt04puaeAaw2yZR9M4cH6S5HWZfkTp
BXRB7cT2C0bjJT1zmuI6Vsai/jt4lMHVLY9n7tbeeaeGCAkgr+WJiFSmbL+MlqJh9sKi8TiG2e9l
U5LtacZ8tKMQGO9UkaQnJl5yaBMz0jhJBs+tcOqr9RevGAR4IZ/iYE4sKKytx30qNP9JsJ0vPdE6
KzPrCD4Q4rNmhx0pKvz+kSZE695kccQN9RB71cGU0J0ALVDeJyn1hQxkpBp5XfJHHCTjkq/RxQCH
KXHKcYrIHhekXluKAaArX0j0D7HMxsVr+NTU6dJ4oMLlX6X08siZaJUk9KYJlurANk7KINc+ZCqo
0PygkqSfE2syc1XXssqv1d8ingQss5MVW14E/NsLsL6v//zCDRP1u5FWvsvQ7fQXUI8eLitBZpsj
k0XwAC3fBwpjrruhoOtIGuWruFhgnHTL544rWAF3Gxd/JUB+5YNbBlE/D4kgXEJXK3cv4k8KirY4
nXM8WAy8xb7VdrxIPQ+PN9/r+UDJ2ZWBtk56P3MFHQxc+otlq3h5RTYo5AII3360CpgIXsPNMmI2
8L8K55f33fqL06M0zQzqICMJTVg/tAEeSZtSxlG5pjuI3pblzBmKQVO5XV3FUiSkJPYL4aQF9EkT
TL7qCYPdHXF/3QH0dTMVD3GZoYgSIKUxyV2ibb7THnKHdYyeaGzBBcyRNRBBX/F6zMfmFnzh3aH0
9PsbnQVFlAfGYpHvFRpimdJ6g0I5ZPUakS+U67v6xOIVOmKn6YLguGOwWtRFm0o2QwdDMBOMFB3a
ibj1o33h6Q8LNTNhjADhA+QuSThdxSUNiFvvXQ2LjqJ36921Aj0U127e/uUAE/+u0ytt6lbTQfkI
Yq5dpKsMU5YWzZPq60s4dG2Z0bIPDsWLgeK/+QmwjMMd4S+4w/JD/eKZ2wWW+BJxsBSdIb4f6k+2
pmbZ9G6RxN24NQW9Ei7NXpcMi90N29qCBwcbsWjfjUsiy9Y3xH5GHB0tiWTHy9KPA5g9EpgvlJll
o37AyEQxs4VWBZWzLZPMwP577hZsO6EcELVZnTS/bSnYngv4CMfVJLs9TDLE2liXVAicbIgsgH5V
rSFqvnOP4krueH22rYxnE+J9+Ybn1FY+17iBzx5O4NVaOtDHsgZ3U1HdH+CLDGnTXb1QDsBCignt
wTM08alH4p5xnZtePmVOgwPn6XUuxpRQnaWDjUPIhz8jAM+gToeX7d3H3z6osfw3s1VFH7Ydtm0q
gzLIZRAsM2PGWTWzsHNBrn3Ai8xkgF0/IgoA5xZRhz39t4h1sLJR+iaWIQxWe5WXYDRSQj0/Ie9h
MTl81J1g7eu6zcHz4pkOeAU8wJdb26/pLVI62hodAOLgnS42PJ0qGbpqSviYtXj6Cki+nnOD2K2O
b3UigON4pMl/cIfjEIv4Xg0UHsUI69Sq7oClusp2m+RtATG7hMajN5PG5Hc3GVrnMwCLeCYgel35
mCrThJtH6RL9KvJVUStjQRv1tWK1J+SIHDgCbyLbD4+gIrG6gMgkBrZBPWo+YbDAZ4FNPDsivM3T
ohNiJLo9EhNG3GGPCWJgUo9klGEu3VVZK5tghyq+YSZOqSBmX9LaCTjcCfJPnAkhns3h0iug9H78
3ZB7c2sTlwbGo8EcwIcQ+TDN3Umx6LzRzbS5YZJ65EqRiM/a/5pOh8kn+P9HTy+Bd32Wvr6Nikgt
gSt4M90IpwaByxQMeu0urSnJo/IoZmDrBu1VZisnqcyVHSkbSGapUfaTT7f4JCw4n/T5Ez9tCj3e
rcWNspBTE2wWt84sJglXFL0Du11KO/QSw24E/t8Gv2tw6iHDjG0R5H7UyvSTE8tHZinFLcexTQxj
l7wGihSgvVgTp+9L9njAW2I4bH1TU6rDAa6tsKHkTkYl1jPAxhtKVk8+u7BIh2PWaoswr1HHJ8Bs
Q1Bjm7cvqt5PDx/J5t2tMkh1oaIuSb3ONTkYVXrfsYsPzfg4o7UocRn0IT8o+ur/pFG/XVh0MrFM
86/yO3C/LER0dpZdVHmIi0J1RGdio++1LtIl7XRgoW9bBy+t1NRwh/J1A9Xb6bwmte9DuSMBhK0g
dtP0PJV60khAKag3HgnvGDXZv1hoBW4pIJKS4cffFMEc0hcKzyVm1s2FIbD+tSfkxPn/dMPQhtZi
ITc7y1Z3rN/eH8xaPvVQa3z6k7Xp6xFAw+kBXWbH69zvqjyD/+pcyBO3z0vlahoW5DR1EWdvyTaN
jgbnq6tNCi23F3T31QLoAeZZSZM2OnIrQwf/2902iT3ME+NfdVE2txFBCpcJueNgMdewBe1Y18Nv
WQCuYyrmTjDvErcHsqzY2bAfLmOltwI3jb6hbGtWG2MkALYP6ka7LplTp622ZoN3fMMWxX9Vrx6D
XNCoVCxvAJ27EtP9LlywR6IBWbcXt8P33kHxv70voItXmifGey5ozXJZYcfxVHpvxUD3mcsZaYa8
WV0UUo8sPg2mUejTvoJmcDqKGBJj018BlpSlgrG8Mr9D3Uqtp7K56cEb1gdqi2Lhno0kBmwq+sdP
bTXUkswM0DxtI+Z5XfISZUbFh/sB0TLoJjOZdh6Oz6lU4UUnkbVmbAy1tW6I8yPBMW3DsT719tyB
u0u/hR6BokodHGs0EEgw6qyWEDbpdr+HDMauMtgKg6kt7ibdUDlKd0Dk0o5S+rZjP/NFPiIL9nzp
b1m46UilF6LgN/vG0d2He1YAo4C2HrdlNacRstM9w9RW9KkUNRvEdBPF1zf8NJhqUFejEfJ1o9V0
qG9PgdGWbMIbVncnQLK37ZH9X9tzsaa6aYuOh/L7EK2jEUDEO0DXlb49LmFBZHfsOlJzgL3FfhJf
2tWELjmcAKyhCCDihRRgY4Q94oFUlc3PU4uiSOKm0o4UYXYZasQ6O5StosAEukmePLQhQ87hlUdN
Fq9KvC+8CccGyYPZP9zLkHNz8qx93Cytq33brDQnRJaUbo79Lo1CMRSPcA2QkRmbJPeoYCvZNpeg
afHBGhSTDjEDvghyLpfb3Etg9ECE9/gQVWwmt44dniJIkD4sau/ySD8FoI4XxMg5/4W8pasZJiu0
fJ0KdlVMT1oGIhdrDhzAyCTChfaA/glrQ+4EZksJRraVApPNiQXBD6avM9leCKbLvniJYioAT+wv
1PlnOJih1VG1e5uDmPHniq/mJXQECW8aUTm6TmeW0zYyvA2kWnI2OkrujPdSK6herggUXR450CmU
7OIv5mXsbU6c9o3NGsG8jMQH2747vgwijm0usJ2+FAU/8s270TGMUrFARoBRWg++CMPSIufdENUp
TBwZYFSCgF+gcl8SzWDYqXFDm3mUn7vTQ1gVn3eI7cFmwyVTS47aZAq0v5PmPegaOyJhwBB5zJBp
KYgGne3+PclkfHFAWSewBT0fJACGB+8WsXJgv1pVkNMxQ0JfGlehOlS2K/zfS4DuRT8FOw32LAV2
tt8V7ibVuggVzsno5+Z4CyC+pLA8Vu59KMRGvj9EyxcAZdLahkbXa+cny79eX8obDv2KQZeuPcbw
T3V3XyerblBz1ZWtHqh5yfwgEutTk6BidDlZ9StaMogOMOzHgeXmFQdqBq9Epxbb9VI3pnlXFR2q
s8x9JL8qNvmxdgZV/60d7iWcoIpgYGRHSNOUPKIzes0DUbXbKYWu5VqxuyiB/brE4B7l/2E4TyWX
FO8YWEAD7GlUXlHfWWRR7/n97T1F/CwIjYEaRLYz8t2y+DwrKgDoU6pt8Z5RNPuk+SviXPeHqDsR
r0NiBwReR1mPeSNRq+F5SDQt5+YPZajMvtsIDIakDqZ0Px6zOKnEPw9SkXPgfL8h1aZE5qsIEbJb
GT5J977lqr8JCBV2rsmeApLiYJ7nWdVvKG14VFo23JeR+Y9P/4bHicIJwaP54vkmMRmfzSsUJjZT
qIjt3IFDm3taplWlJQp1ibanZ4qANOSsuqp7YNzJmP737rOcXwuVdsLZDQTy6ZEM9zFcDVpcpjBz
feE4cI2ZbSx1heR1WCGHiCkxfJgZc729yoy2aQZdJnNfo3xoQ/fDhzoJR0AreiA/zKNdDtcZOfgU
jj+ry5/Dpvhky6XCH09rPmfkTjcBL8nRN7BliO0HmdMvjNqQquHO/ovzrTxIPI+V/VReq1mBoJAu
aNHIy3Oy/PsdwAfqlgT3EdupKegPc/7TJ3204QPN08pRSs80w6/pIKKv6OQ7NTKlcGAv4UsKRX1F
HRnqUV48C87mN10Fqdypo8TbV/tpPmOp84I+X3M67HbmbR5MskygdZZ3femEl03E62e4mFut9ggI
Ots6x0kSmKhpyvbEd8J5KWVy3mIoBrpbI4ZVHYgmkyVqrd986fXBATXnUvq7RmTi1dMElOGoYvUg
k6ktPqDj1siTMxsNIYU0AWWwrgq/ik9MAqQZc7IU42cJb/xFr5+iyMsBWGHbIdIurT5eAkrZnJZS
W9721uO8JvofMynRNxx7pGLh9GSGVsYaGFceSINXktqKuUbpZXPwZKYiMMUF4z5+ktT8swpHUjng
lY2B0WiWBfr0Kq1jtMRc0uP9JFDr8eaPPAz+b49OoAh/+LUZsAOxVwe77iOlnvOHv20NwOYXowfG
OxHTwWt2y8sMn/andGCPsiadq8jTXVbKPmTExd6B4ibTJSyW840z0fzR4cEwTG0ej55w0jCl9J/h
yPBYajNHxCGTqnyg397g1QWhwLrL1MuORmyLB9Q3S93fXEPOtYaRwsdiZKH5FdqWOKal4mNCdSQg
mV6o6gvqUnUouZm1gEZfJECr7Ybh9iGDPTWEvfTKeNZWtgq2dBqBUSZyYaUvvJTIpmvXmJdxPxf0
J9K7MruD0UHdDT2Ke/oanXv9bgKT0ZB8f+zT5n8PT4+FF6CqTeJ1rMQ7CNtOXPlKCIB1jicVrhOZ
FHsj4oYRa6yBa7UriyKMDH7+3P7mp/O2IlEtJBYhqbxMifW9xlf/Wt4bDKCpO7Je2oP3cC7KOjVR
Y4w6/9XNJ7y944C82iMjUocexNPPn4/fMZ1rhRgN7Uwig56JHD/m+AJHwj/aK1riQH4sM3NtULvU
kAseCSAa3xHGv/qyna15OioUokjvhMX7wgNhEht77F+LXu1K5lAVvOD0tkp28pHSXtSNYTy1MYhQ
rPXxUFe4GDVnN8S9tPpvQVv7zSzz4iEwi7AtV8AgJLkFutBxg7oNsogTekVJIMub3GFCAY3Ly102
t50t5SImmst/A/IVGjif2bawi4+Dr8dbNqRmiTd6HtlVTLOEbUmFbC5GvjTafzaRntn7Ut+fuUNV
bhilUiLjMmbnNsi7CeHTy90NLVtAIhuWFSb/wkHkoZnyVjWC9uqad/bFglG3qmQakdiWab+mSfn7
40/M3QqItVmIxeLEhwVRqIYRb15jgM9Yhaa74OhOlH3HL8SIXKWfeG/7x3tV54Qxe7CecK9OqPGP
Nh378yFIkjvQQVuMJXHPwdd6hyDtFWvFZlb/KqrVu9vuiLZ+aQaMTa4IbICbK1I88aA9evDhg/y6
E+8xcwDlZWy1RAXOktWoz07aS88YF0c+WVg6CiVdSNOfCS54RwnFXHj1MSz2F12473F0hJkThpQb
HGc7aAEThFiTagleqcrntouGrGDwIjTZHuqbcLJnAIFlLc3zSjLVJIt4Llrz3mvnZ3WBSCjdzXmU
ChhclgPCgQAE+otiFTep5hgaUHk2MYMXdMdAcEU8wuKrqxZL1otoR19LhHiwZVt3hu0kDZPMvuJM
EvU+1ALcmPEVkzCBef/JTzSag3FHDPAF5N88ZdtXsXkhz6dM8KzPADS12NYwsJBxvZqmH8WnLwOs
RYUw48CHyBghbP2JzNu97QVHxvBzZhiOsRx/qZCmEfgKjG+uIsKv8yspymg5Bx8SkDzTFY5FQx+M
rQwxQRfl/fPrUt7oURN/ho2DsWaGus7JDI+ROn/nklcFpG7KzL2zijhv4MA/IUtyj255wYuM1qoy
PwbikE01U3wBZfx4PyfjHb1jsyi+2Tp6Z+NGXoouFb6pChC/iIRdS+fsXT17iy/P4ZpppL6iDzSr
n2aSzlbEzClnPjfaxwu79OojM3iy+JGdbrTUXb2vckMEqIe5qpbxB3hdEIoJYuKkek0VlV75ygOR
9RHrL7gmt4SMeytCYpW/5lWmQfEHvM0IRS+C1Sj89HDGh5Adz+aMB1rw9brL7IFxE8hJwYCDKywr
3zfZ61zWTpDKy+dhX5Wv3txifdVwHfz8/CKIvEjPjPYRZCvUdYpx73AYZNv4IxgcTEbCdL2HuqY2
Xyyc7HAANV5MRFKAVtbXdZPIzmYUlWP1Pf8hxVT2SjZw8A4N1hH4mEo29cdJ8xoYOm2TpguoUPYw
GJwVEIxySnakYeXgSFUlDe+R9IV9b1Jys4OJ96dHQKffaa4/aHbO8Cv11sE4wPGw8/L7RyxZXwnf
tuNN56P7T5ym11HaC/RxL0tapN7j+v0LU0BZ7m3nsFertoU0L9Lqe0SDmzlIUqQNAV4N8ZImo/Ro
g/Bj7zyE3jc0Nixr3YoLYp9U/wKUYztFD3G+VANs8VJHJisdHEGKTwhk1SiEQWfvr8YovRlqc6cD
pg+g+JVOtjir5dpHAL4zCw7Pnu67S+pJb3AL8D7N5dAdb2/0hLMcP8lmqTtARWjzqhJTe46cbs1n
hlq7l312n8C01qleWswKDJjPHWdrOAzRFl3MK1tkSgp4QTpz7US+TYQcridQZzDAq5NJxbhatAeO
5EwOiu/WlbTJJtfpqOuv2By4XOyJViqJXE4OnRMjXMEpD544fFn5ZGXbsuEuTpQ5XGLO2tBfaTL9
mTi5O2EsnPt31uRfYBdAP2z3qV1OoA99QuDrZs8HJnynGR01lna49kQJ7ebY1bFtfgbqmGI+TG1h
aA8AZfRg2LlK0zJ0oKZfTXhFdJMghEj+e5SmOTv7VPt1oTqQ/oDVNmmlb9gorvk9on/x8buu0cB0
ibsPaJuzLJlk2YYQnni4rp3uwJaXsTX+ujlUAMiCSoszI50qzrOl13/IxbuYLx4JdRk/WQY69u4X
LYrGCHT5pukSAPlzSBAbTFk31luHZwZ9gdH/2jnxofLcZmFcGm9FGa3B8QIpH1ufd+hpoRPWLD2k
Z3rLoTmq21uSNwfwir0mt9ECJ7Hxm6fKN5hc4J1AFvBUvzSDvpZ8KD7q0ZgZI3lNZnLSyl+TeMgA
MBobEoeRzdl6bH1YY6pow3/dTbC0aYXnCpf0RzzKCjMXcjPD6XajdbIQ/yh5Az2AR5nDz1/LEAEQ
ysW3EXnx2FwPJf2e7/PdsfEG8O9bnvDmn02XeE/x91Gd/dW6cBfH8pEjgyUPrPl8q//uhjifb83n
WPNw0pDVI29IuI8trxiBRN6jOwATAKlIDbcULnjLyvYcHNp0Rhqwv7AtCTXYpnrJqA1RbIgxJ8yl
K9OydFIOwHSPXLzBTxtzhqzgmMn8epaf+LRso5M+OWiDA4dtZ9HD6nxa7VBtLivoIxyyKmevqbPe
v0NO2v79TnJ3QOsgCmxPV5KQwLve2wvOrAAfBiOxfg/R1K02Z59uGEyRb4uhSzBEpk+kQmenwoMD
lPiPzvGxz7NtTkUbsUGj8MtIOZ1Gixp7nHiVdMTRjizC1Nvstf+WFJCu2I418oIwNzMaYov9iZo2
njX40M01yqg5wt8lYAPk5ynliXGRZkkitLiUyGz86eHuXe4HSz/W/mbmMxoAcZBNvPnPwy7zq08d
iyPZXWL10zHXWsSqvmKrpiKLajfuJYWadTD3Xfn5RBiDI4rqfPhNDFGht31ooJorcbLq/52KIUKk
076Y7217tcL0103F0FaHXmPMGrV3pKShS3AHJGPtkv4XFjDdug4cyYDPAudVvCN0Csr3or4mh7PW
jo2NTcmafXPAIUsVjQpUSSfBS3jBHn/npcRET2FFtLh6b7sS8mhxlgtMXnioHA+lMBc1h/bliKGb
0Jte03jDCRtJNDxKRoGW55Livt7vf37AYVMci80UODO8/5XSJ1WX6yGpZ1vaS+jenY/YZQ5c0ctK
1Ei9l4+U9qD9gl+mUdMaSCZ6O5zula3rPKYCVsoWUzgB+N4FcX8HELcJYCzeM00+6uvShUGiz6sQ
Mq7K/bl6NNik8UHQLZ4L1Aj/uMcGMGbnU7dz4dUhV79ZVUASlI6eRB7cbqkQQEf4qlbcUI93sL1x
A/3oJ+wjh3e6H9ByP5/S/5p1GS27Z3t0/V/DDiFVm+oKnMrm5F/0MkQKvJNkneSglTAxapcJIPfn
KVRSKxwG4hMOo0s9FXuwMidqOy6D2RptW8bSG1hcPeWv/wtJO3YWe55TC3M5rJ2pBtsrC+Znc9qo
1OgWRXAk5vU+4pJ5deq8CSpbLScrZt8Mznr5W6pgUFRHj4Y+41G/9KXcXF0+vCRr6ejGlaKy9jXI
xsU5hBlZru/yi6WrWf3DtcoPUMFl3B4Qx4NR9xDmO7EwSNUUh9fXst8EXrwD59AjZkfWhp6yY2F3
gFJJrOcAdgfVnCZ8515/crC0/c4nAo1PUryYNGKoWPFbb0PsInYLghPEbQj6AcOyGwnfV1g1DCte
7WjQ+zHpneVO8cTqZjedXNJERYCDMqb7NHqLkNOcbbUb9MJAgm8hai9KoTF7VbcDSEK3IteY7D5D
t7c2hrWs2kUBGC1uSR9ZGcwbK/bfAFUqJELyd6JgYZa4fL2vpBm82iDzH9S4Xtqxz8CEQs6UqAZ/
EBHCQ5Km1VXi0A4Sad7BOfc1mOCxPJUJWyVh1MJK4N+65bLBhAPxyI6w1xCVSVLO0bz7ZKSzOoAZ
AgcoaChNmeaorkZ+blcmsx2clGAXOqw/lkFITpjRI1HPqLHzAVWOF0JQJtnDzS7bLGa2z1El17eK
6swWMzX1vPC+Tiw2ZeYs7t+qtLi9enreT3zwkO7bREgM1tOLsOLPdHgO6nVxh7JLUT9L5XU3bUCa
sp+WDADJHgm2SGgwMubnlWhRkS70dliqYEqdkResy/t7dO6YE29EJnI6tVd7Xrv6Eky6iWvElgtz
PWgpPAAcCjo0QRuWiSTxvhuq8GNgfwJErBDSQcKWFRQCFEMEyBW9PsUs4zXlMTZoOHNi8HylP/Bk
rSNykwYV3QqNB7COsbf7NNoHqekDsG0pOLuWSM9zup+5EQKkiGrNM7IgtCu9fA2D5lw8IIdqTqSK
+mbTeXXKsLUty9jg2C9zmZpJ3V7R3IrRAVebAxC0NYRGzZ3jmNo6pguMdTRmPSdB00tpQGejndej
KSjc4vFzLpNxxNKK3m68Y40VFyPF5GvSGa775jOx1IFzA+WT5Plo43prx7ElChTYwukmV1dQjcaC
O25+N2jRvTCDk0df3tJoegQhCW81WUBejP97xWc6M0J4Z53iTHjoIEx3gS+HDHkO+M+5xXhSYJUn
9DgX6opUXFxpRO6FmYJm6xI+wH1azfHQ2gM1yo688+GQuvw519pVyaCjWzhdRUXmtzHA33eVE7gp
ok5ocTRPESWsRcIAhNC68nQTF6zPPHWqiH8Qi0+25hgObYYO4gl3ucAgbVjlkEAu3JBE/pf5T/5l
xT4OictGQ8P+Fy2qPt271ckerXT08gyWAs0BMs+zXUViQiVqUqIhFdp7dLiecHpP36iojMQS1KZn
rT0A1piR8o7kl+yXFCpzh+dTG0GUNU2KFgkmjWHIU7EmddBo37j1ykgImla+5qLVYZNDKpzevw8u
rVaSlaYXyKWZICj3HpAp0TjSB0eM7gADRXKsW0SVn3Zp0jsywcpLP45uSABaYAPb+482n18zrKe4
bRVQi/bfsZH8uZ/tawmFaVaWYtKl6rKIC8FW920xxDgtffPQzMugNqtivKkNNPXY6iRv6+hqA22q
7luCYQF6xqrP/EauuhGGGXyC4r5Gg1hNSzsiYnhiBLWMAm7vOaRxXwp9PfuiJKGAZYYdkbLRe8HK
FgPNrHlQkeKLVa9igOMAfSfBM9SzOFwFlZzPJbjzT54//F1DiAcKFi08GeGw+HTW3ML2HHKrGGP5
KQmsvqLq61Tc4hnC+DW4d4MtsRGcxZPyNkZf42wrK8DdDY9yGLaAWrV7ozQn3cTf1pk+36eEFPWA
qoivIHmk2dyu8PsYQjqeLkGF+ccFrpChluRHSLxvZoF/UeS+wlVQwTBsrZXvlvIQ7BndQV9wLnON
tKHhF7vC/AI8hTWS4VFP/8bjvjflG1mAWWSlbqkp2F14zmqgsC88haZyhs5JrL/P5K6axrscMTlA
46GnnCZfyrHReYnHbDA4BxSnbDaINJ2oy2b0L2j0eO+2LCEUvJ8yovdiMDFPxcgujJOweUVntSW2
gEKW12s4g13va7drT6AmhE3Id+nVIJmSvM3obg5j/BUaRoMa205xQS/bjW4qfIQpEhKrLXZru3xv
0lU8TTRujaLg8Aq6MEtyBppdcX86dxEEH2qhITTKA0JO/mrIfg8jM3tW5iIQWc/1hNp2t688/lti
bg7JsGWHz8/3aPX8s+mSBi8abq8ZXObBa6K1R9QZfPo+3N5SXdbxsVwijWK388KbBoZVaFqqvE9J
vfmGJTjzalwLoTX86vn1gb6ZHu9gecgoF4hVyjIaPsKKiHb9pkmOSyvTjHfBK98XhSJk817OxInw
K74/BEpsVQHYxN4mqlKXh/AtT/QRJX9CoQDUiWcTSc4vabpUQn32sKjpRqC8yaRSly61mS7X9XP7
YR1JXCwyr2eShnzbKhJaSvV/O5w5zJ8qwItfd7mNqU3HDvoqYpLfWxsgDuUsjrbtmHv7Uc6AP8nt
trNTYB8RcFMntTvY8OCjJ4kUCjRyNMOFVe6pTQVEXuIz4i2jn/pgVo/fdRi1iCcqDDd6sAxXdtvy
3NMy+QeOYuUtV70HVq8AamRsGU4MTBebLOLmpMK2eP2XHcEyd+aQwDnIr+BEguQFiDti4xvct8G0
REZZljUIKdzZdMC10tx8P4NuKWKitBUUaIkPHL3P5lkD+hZlEB1wVJA2Ln/c1jo/weBsDpV0ki1x
1IUrRqt5mI5ojnRrdlOu/9SdzDeTWFdVauyqxwDSDSaODISGK8QEZBfsPC5HLgKQ2+G2TubkdLsI
k8i7jabVUmj+rylikjvYVOhPlPQO4cYWDUMACJxyRbEupUJUJfDXy5Xk86ZIgjocV58oVLK6A28B
MKnQ+I+r4Te8eIsbwLKv+VabWzLkS5nBUMswXean3zRxA7QO4kgsxLEJCCqSwNSo7zSJ9BBXZyTN
6jXeRJ6yJVxzzOzBFhVqibqtKJHD9vw+Ggr1KdyHE5UlqOjphprbYbVb7S/5JLXoTYFoS3/0I7yg
bzlm8BTOn7AeiKphY99H8glJU8pnuIIChNU/houqJP/j/Sz+EQLewP+EIkNwXPuxLvcl0KxxLHsa
8FBYOYzhRzZlFTm74LoBAYznrkvCSS0U2/MUbrE0uia0F/d9QqHvrJ2ZF1jtATQD2Oe+KvolutwS
NQd1uSc/5BzcgYNrZ5t4wd5XdYfFYrmynIv2Wkp40fprUHYSji0RryZSRv2/uTIE3EttK9GFEYxL
FLulSXLE0oI9lYSYIqM/SvMhPBzBpoLRtFe3rFQTJdiy4SxXQ5KADKJqjU9GaaxKlydKF+Y349Zp
gbKnOgRPBuR4OLb2vE8FRr9sGlgFZ9qHfST75OoXTxqCYGljasbhe87z9CRz1xbks/DjESfH7bHX
+ZpJ6jUC9s5uSUey1y2eswwCXZckpM4oezh+nQARoj5UY+1lrZg9xRCCvPgQuRzV4XaJNJOnrFtB
1dEs01sndHE7WDh7EFAJ9k/jiJ1k2VH3GzQ7c/gogjdyga4GNGHk2FsSPgNGg/9I0jshHwKRpExm
zD7UJA1AEYtCkwYgpqWsISKtHeWkglDD0hoKsfyB09hZ3tgl0V18A1Wj/bM92xMKXhJCPscn+Rjk
6mjIXTi4UzoEkPqP/1yfu6cjMVx17YII9k9YUgv/xT6lbZYGFWowMrR8eeMJOUvAF+8ka/ONhSTy
1eBjHTuXEaVUlTqKLTbkIwKu1hQJoMMCbReK+CvD9VT4375EpRxF8WgvnL7nA2Fg0+9PA9C9qYDk
ttPtooZkz2RKB1FR3602xQFmRl9W/QmJQjw4P/VOJSYLSNShU9hWgP1nW4fxyK2nZvriDWGyeKjc
F7qsol0IUAdx8m3w09z88EhiPALoln2HgBKPZJ7ppP1XC4ETCKoQ3CXNPBjKaGuPyRn1fnLMFqQD
ctU+0Buhh/xEDylJp2SnGXe3ke1wDrnkBHm2gA2OS5kqeHOGj61XsT1ujj4eq0ZXbHNp6jGFucrn
LZ/kBSE79x8Xpc1bYwOd9BL7dk6TAdg0dVfcz24980d12+i8P8OXT8hzQaGCq6QO68vsC2h7esug
KjsydFFCkYjtJfUUOTSUbSsSMkHcT2P30i6Z3u5+kpQGb53U4qI/jRRrQfZAkbYiV+F3rbadMwk8
wTCRMHJ52u7ns26NoqHHHYc10B5x31FFrlwB1pH1iiW+E/XEcBAs9GMK95tYSRvF//+2UkO2sMOZ
HccGwgiMTNggWd0kAxLnipuCDPQwBErY0bsze4868J3Koo1qNN7XFuN5pYwQKJixLuSEYmdUgnw1
5F1FMXcQVh7IkFp3YAwf4181AJkuOn6U2leyP/D1ig/zP/cWBEt9bho2x2mymUp0dzO+1kAVgOyi
53eJJguaV0+eC570CeFUksYSnfQfCyAnUZepem5lHItkGnu6RhyqGZ28tJu7O1fJ9D3gcJ3r69Gw
vEnvhnpybRSNlJOisJ/GsPnX7syzaFMsJphWwUroHLkDpahnHfAN/40QRZG2nyUrvxcGRrI79ij8
lGINEWru+8sCb8BojYEB0eXRjckyQ+wtCabYXrZMPONUI0FoRREIAk25R7bLwEPOJSPKaRWQYgZ4
6k/9qOY50NCqq+qmJUv2PwZakv4xnBjU0xN6Pqo/MQkdWhQWb4mqCimipJytK68truWJQ5/UihqJ
P6n7UAwLxnxYyv2nNrGSAOOuelT3l+sJdj+WYeGMVFCZ3f0rmms3ujguOUIUGFLcNrFgHG1Rfhes
HZibOKatDxNZooYKcjXIWxkZHR1bXdUzwBIKUigbbh0Y10sKd9tZM4NS5ldUuvHnlBAg15QIiLQe
J/X0osbw7bEhsBTwzq3AAnwKKBRPDHupIcnfbI6bs5V+H8+U6WCLs6zazlaxKd6ohH04Me1SSpkX
ckO5OAdyWbMcICPAk8UgANUSeXEwYsONUmY65S3O5QCGmrL/ZXil0PN4xxtEKByGzmK9EDeNMDIR
DcpH8uElnEDuHaxxUYrW9aCSKXB6aoFIdgMDJOOPQnSSB+2p0oyCYuWWl8NvfCzpYIqykjBvBZpj
/qTCqzRQPMAPCwy3widmm23bOiunf3zt9PAYi4yYtmsbD2NsJNUZ3xS0bHb/pGwno6f3HIGNACUd
dgoog2nI3JQRNufwu6e1e9T44Eg2vdjONxssd1SNQPQATJ3tNDZInHMfVJUCRJCwvdb3Khy2VXFS
KN+lAPrEhQJ+oXWZnyJrKpebhfW6UC9x8d+/XMaVOk2exOjfK6LH47mzYrhKELUbqeSBModkfIjh
lphH0A5uA7rs7C9qZCdBHeWLcYCcu0Cuj9FfpR6NGgtV8UBME62wOq9J7VMrhlJQ+r74Dz4cYSra
cJPmW/0JWIVQ1h7AShm9SHlr8SPWbiyye+3VLMqlhfLmMcxFLsOEy76zEoA5MfRrbzO/I4Fe+oqc
omEhXUmU1PCwkVAqyx8Uuy+XNWvhfUkqJBeffNdtUksIhhdVegMsvs0UnBcc49pEWTRHLVzehB6q
eEO9XndQM2MWK90lcqqvFVQQadJBfOmhgAhJqiuzcGVTUcYtc2dplPD2+9jC0+CcbglNFdRa20S0
Td5PXiaxAFUags8eFnW6pjeVE/HwOKBdu6GlfinAzTXzmkdQzoGjQp4BVBSq6Ml//GdA9OuJwzkg
GkP98x0e5NQ1Nyr0+X6J/FtWM6zpdnpc0yb3jHxFqsPVgx57eOREar6HBhutW6nkZ4TOW9nB/Amb
qUBEAn93nP5dW6FGqQxtfvkTpmIiazI+OoOYlJb3BoyGDGozO9K7HMsUgaDsGZ3eIvGW45wUySVG
Xoj/F+CsU/ZuChDMRzdMQd8zvD36Co27taVblK4uXwivlz3NQAQU17zs94jWuxeheWQTsEK95kHv
uSN8RbxnpB45K3/h2G6ykLzMcRe/lsL9uuzjFPFVPAMH6znZ5TY0pVYt4gmsk7PoRvNV8jkZCJKH
GC5GbAN/99y2x6f6dSiQnYZ0xc5itmfhW+5q5KXkPjBktxyIETvXYxxpww6TvAC01u8CmlJl2JNd
44iN2GyqIFwrpyvWpsvvkVudKiPkI0TSh6qljbrEUG9EUXDqTy9Xt+urRSO9oFaV/KuMy0KH1Zw2
rje0gEYau5P0xyZnCubfZXBlzGU14VHS9O3z6qo8cwFziwJF/0KugTvXgcEjA4p20wrV20IXAABY
ls7UajAjv8VT+bS9H++daeWj7RSilw1KfaXF0/x/UOvKIxAiFUtkD3HvweX8jD3J0prUZIuTCNNT
ul3uBofi/nlsR2xbZqCNe7GpHIBL0pQNBiCdxhWS5apEbzPjhNrM0WGHMnEM1LM91ORausZK4FgS
U4A/lX2XT79V814+27N6MtW2e8+Pp4c0T7Jpj3SKCwwFwK+7AZgnrmMMB8tgFAFuMgZXt4jg2qAR
8dH53vudPnDfiLLqIhT9Smi5wJJONjVrBfC3YQuxUc/wI95NNN1TF8doeaguc1z9WNdPSPx7LD4R
Pkr9xbe5s/MLKquvNRCr875gadTrQXPhdEVELbBQErffsD35wKj47qcVYgxALc/Zi1er0boTLfoO
PiR8zhpmbfG0OMQbjqbaZ7O9g85p+pWDA01qJbbXqvcu/40vh6rUfU97LoWuzosJRZibnHZhDoYu
jM6KW+izduIqha/dtDG1rd8H/Pes4PiofA/An8jXti1Z+dvDnhFJ3ZSqemPghzOLUeIRscZthayU
04Iiwy3u7l+vgtd5WWxP9fy98FxRmks/XUMarXSv7orL9whSsLvmitmvYj4gtHvYTaTYQbucxZUB
flIfL7ViU/202DjhOepIJDDvW3K1Z4EXNFYUj6+7AilFH6HyAmSXbER8ofbaRw12+NM8r3w1/aiz
lYzHX4XyqidePqzi+CoWJgY0g0sbkYXPte5JYJJPxO8e+d3q0y/NkNy90qnR2vhD0QIypLIMfDna
9f5z774ASKFwCp0piR6aOJxc8Xa8FiW/VGFQlKQLKjXJyLEVvonEleemMUhzDgePzGCITQ2SVUOD
zKY97Cekxh6O13u6Bq8fMvtSmWtMYuEVzGmO53EgIaCxP3MWyenk+789C4/sTH8hzWGC75M5o6We
j7x7BKkx7TfiUq4nLOJn1/UqoQefkHXnFqKFqc50lseT+c2yUREPpQ9a+rTaCEQ0q9u/T1kqa6oH
3ZNor0r8Ke6UbuKxtrR6fRm0kTeB8pdKt7Yipxco3gJ6PdNz4DbcsapFVQPTGhniWAzsFAOxXQEX
1AZgmaAyjcqT4v7ZppIL29wLi/mZW3KzyJqGQ8xjTXIo9/iruVMe9tBOU1ZL2ZGCc/xH2vnlRBhH
vbU5aGiOoUDWKnT//ZWwpGXl/V9PP8Qpvj2XJNNcKxzNZPN6NRfrZLJlQ2VyRY9eCRKelsF3GO7N
xhQDHMI8iXJoYd8MY5WpfyJJNteaZ4SmOEjumNsb/SEI190DTPEx8gUjFPcKTQ0MYCDwZJkeNp5f
1cnKpfn5Vr4vlkzDvXz/qqDVPEWZl0fJUGVDDPEbI3/MMGMNv99uIbz6VmsWLar4xe9mq5GGSmVG
LnEu4hPUIzlvulhBbbHsjosC8rL8OzaeRTrv6qWeoCmV8Bu+a9wJ9dZR2FfpCOSgX29x3nzsAotw
F5f/d+P1P8HBgNQ9TIVv3JarDV7EXzjfeC9PwrTDLPEOekPKAkWfPSRKD9j6911gNO3jy3W2q6OD
ppYlGZTMBAVwTk0Va2EjQFkz1LSzYJ8Xcgosn7jWvK9r9EBXrwyyy9kUuTDWGb6rXfCFnrLzUnKK
H8HiU8KOJ/y7n0eSrTWt8xKDUy5ECAoGp/0dXIIhBYYV4wutHvSX+jVct2JXZfx8OQE1lUbsz/Hv
U1XddC70z6ZwPUqk/DxypsJf+y98WkZ4HHHnIfgaD8BiIeg9RnJLI/DHb2j7NAFzCAWlSWTZFGu9
FuZd56i4TkWvVV+FOPKkvOinzrI9eeg34kHWbQDR8qtke4rIldgig1Gvh6KWgxRI/5FZMr2QCic4
jwaSisHg34zEl410W5lR0OhHo7UeG7DNw0QSfLxjH/TJRPz2mG2NTfuwDDtjgdtpBhbrBOBPccIu
KI9nLO6q4nxAqjrQT4+mqsyFXjLwlYlhb7M1wii8NS5RI3FoKdov3nAaLrN58u5bMznyKsU9Ard4
NeJHy3bgaZtjc0k1EXa4rRAzo5MaYlI1nF9jYUIeLRgbmd/Xm+bsAuIGNLvE4t0YOo9luSalTsoj
siaF0IASkzZFZfCH1NOuIB1gHRYtN0rhWOzAs/8O/7pcFb9NaATafBWqkrkG5TjARWv6qKL4L68n
ZJG5L7rrNn7LaW4dYvPyyT4oid0we2WEXO3Ts7nqz4KbAxoKE6JV7Yfhjg+VQj6Od0ylYGPQit0F
QFSLmIM2OSK5xjqiXJvcSSM4XvncxMcKE/RzWAnELP2lExWQKJvRQPpLmKWRpnc9V40B52cqscNJ
2Gi7QO4l8BRXZCtU3i6n328vZKMjfdlK77xXvfmwM95qp0Kmvsnld2LhOPopxyHUJ5xG1bXBXIjM
1h1Ru8SE5UkfwCtuZgIhE1V3u2pyGlBPz+fEPn6j5UkNaW7HcJ05YXjiU8kNI+VAU6AooJ4Bh2QZ
6gLd9fHaCnMEg7A+i8Vi7Rz//1cfj/SZnpeU1+IUXF1JvHmhTUHSX9fr/qLE9+cd+BrTbQ9w+ESy
AtuDsqXXmGoF5sKZQXf1SElCZofHnpEXu4YhLZmNKg/tr0MBCuAL86SPpixfkAKrwmAJMjOkH5mt
/6kq2mbmR336B7OS7bC4wloyP7vQbs45zvKYJEnF5oQbhnk1eWDfwioTh3u0edr9nh9tpznoGYuo
AuEOASx593au/28DhCZoRjNEMrf3IcIk9PFsRfMwtC/PhWD4MaAolo7eWYdtgaLR2GXqVAGZbcSy
/zY/ePQFxMdGdJZV/s4hUPXiRS7Rinugd2Z+IZV6vG2ZjB1ltuqNQSbjd7hnoNsj5r4jSmDft0jv
DaQxS4eu+wH8BYPpnWh19aXFk1+BTzZACNz0S6FKGn0LpaCwx0/coEomi6GttMdY22t370vb7m7r
29wS3I8JvYCK1o9AjweXw0I4ByeKdxCV9HqSwaY/6z+vWYJp7J4vmy4h0tc2GVHlNUCrIjzVdYqv
l3FO5KUK/bdPqQgyOItdqjaD2iZKuoztCj39GW+QDdD1lDfHF9Kv5r8vuNfcMKEWK8BxMMBhYAXk
c09KqBIv3qYq0KOoCbgHfh91jxymziqSApNfUc+WiLOH3XRwUZ9olRv79Tig6FDZY8TV8/06HkGl
5MZOZO11u9WIObesCi0oURAMlM2ILCOn11+ZM8YKmMZGsSwPFtIpLfBBkjq5WZjZ2kTzaWe/Af0b
0Tm1avP156ZfLmPPQZwm4t4ZEAtpE897YY0BktNVH/x72saKVyvlY5MufwgTbUyS/B7b6dzj6lZ/
eUp9XHiZ0vcpu5plfBcworeFlgIGz6qayDaMXWXNPxJ2ODCvh3UNPw8CfyecPDriEqPJIdeBpSUQ
5j3jM8jYeyISFpJHMP2abFfi3oyfqjDr/rk3QSTkIxtEO1/BphqqdGwY+k8sy8hyM9VHfBU5cSWY
e3ljZ/IDa4TsWNZbeJgYgkv0Sv0mY7derFaiN+unfQytc26GsC8iYU17aTa+3zDrHyalxKWliEjT
V8BPSsk2vbE8PpK413/nVZ18LKF4u5CuT5piouXKBEqqtNdgunVEqvg4Cik/FKMnnQB5EGt7TiZV
AbUGmE/CC5ee9WQxW50Ai57Ye4Xnb41Rs170wzWTj7uotJbb0DRDiDaTQNO1j37LtO1Er75mqUSq
qB0F0G/HnzdA46SjpYtw1oO91rjGvA4tmL7eFltf2BLhOsLPGMbJdPs4+0wwPm1MMjVjVMzUeByc
/PdEoJfcTCaQTSmERfZs/XTcPqnJEj9MnVhgMHid5iU3zL4p6yJPDbSeykzXxtXNAsadDCLMpWFV
gv6jDO4su2CWYV2H+GmJBTlhP++9bLRhhPRetDjhOc+Gi+BaX2ZhsdJ09iZCXU80DdDMIDIA7x2F
s7waIb6PmGRP2WMuGIiFKX81UXfqrQVc7H9SnePOGK9XwEbEiHwVFi6oqu4AcL/6gvF7foupaY5l
I6TA/TYrmLbJudWzFAj59e9LM17kIRq/BpUdBjhD/z3vMcG5Ony1LmHW1jc8anOnv0ZKbD5P4+ox
MZ6n0zK2VrH9NWgwYt6oL9w/uQYJf/XkrOprlInKnvbqzUaGdnNTZXRoBjfBuv6b5E3wEm1AhcVI
iNmIeFEUNhrqhAAch/pCSEcwtf02cJO7Lfmm+9H7xtSdM8NwkigA5AdH6W0d7B/CUTb9bgwGxYVR
DvnX1AQuvVZ4qalnOoi/1DwuzgO6jsCh8Sb+m9urL00/Fmu+c7o+TTKSKfAKavxMH6R1hMbui76A
EWzEyV+proiaYc0p+ZEqCVHOM135B90c5oiG5siZ/PwdzqSLyRsswA7Cotjgv9jG71e6VSwFRBD5
00KPxMzNsErwrZgvfFYUfUJQmjE1VwVPmb+Va6oaS+7DMPT4X8FX2aHsOdV5VANWH9AZNroBtMuE
KWSI7/cdKaAudhqklLkrtZNdEWq/tiym+AUXACL5dWEjeLU9YGevYSV4lQq2BkrLqRDWWxQ128PY
rO2lkjNC2KV+lSCHPGpqSGQ9ehcN5iS8YBeSix3LjMZCbkU3c4b7m/aY3K5BCRf5rFp75+4ca6F6
Y4vClWE3HZABHwnBPVfuzZjKQC7SWE37AWuk3j/CbPyxj/3ZfboIuA7sYjNII15FxkHtL8InIDts
QIGd97zV42RgrpnySknydxL2uyypk2PUtiRLR1+4+b5vkyIJ3RXzhwFDRtS/uHZb5485gnOJ/fRK
hWbzgQ0dt+vg5ItIFMIf0+FUFR6IbZ5krCEulb27Z0g+D4hFUcDIJSaHJYr56GDmzapE6UM40LQZ
rK9BUq8Vkpi6nhf04808a4uUWuyJZeoFm5LBrzvE8lyKAVYwSyommaHKXHEdT5nkzFfNU1pAIIgn
RfCkldPoqwICL3NFVImtxfrrQOIts1HUET0N7/SgFoQmsT5q2qI2QSBO/2Koa7aEhROrSbV+0UHD
Jxf4i23+VLrd54XPf/ks4Jh3eCKdSv2rSaF1ScPZkXPqRWsciF7yZnYn+5qC8G9p58H/klrhO0uV
jJG9UCI4fKbo5hWXmjlS1jpCEftt8nPd6qMAp+nwbJYd9EKqdHzenkltJQVFzWYsmE573paFarS0
4ZNw1cagBlVU1ARvZvmjm7/5tPt2J9LArVwwLjI0zTnCSahJgLFprzpQce9X0EkWJLYqwADJgBMn
dPpW4j2rnKuQ2MKdfASkhc6erhUokQDRl3t4Y6sKmqjr736jlmCWBknqS/O7D3JRnmu0FkhbYkUh
pnuVM1700uooxv7xujbBq9wZ3qF/I5G5pDKHq9DBF2d3KsBLg8dNUNDZ0hAUZ+bpcskcO17n0Yh9
g5/Zu8k9O7z0ZGjXXXD0XxEZtuNFazW+2hPbeHlu0iSPyFyIlE8aZ6EOKu6RNqimjAic5BaB3CIu
XS5HmOSlnuFu898H6eG02SlDYCSAFfYXlCoR/rdaF/SHNdBOCo3zJ6SMsuEzfqW4AkCa7Lxar3lv
1sygYFrxGLx03sAw4gxArOQOCauTN0SfEV8ENoNgNEc55vtU/wBcoMRB/HFDJrPWAzNeWF/Z9Vbm
/Q8h7oOeUd4kAkAJmGNgIaUJsPMWgJdjmFMhEPJurf8lpaR72X3dKT+T4tT7iMbIVBug1xo/7qSI
43Gmzdg0GCm3g2zxTrsT2Wu8E7IyqT0NuFWOyGNyTK1vIyK/qpc69F+jlStm1zlCtm8vK2EgEHZ9
2PzuwBIZB7+nTS50iRKNn9wa82yZD4AywErPTFRHt+/oKcURv14ECPQIP9JPR8Ugpom5yQzpkhtH
kwtUiePRt1t5n7Lv8l3vUI9tiTvx2qKSr/H2UkGbBZydAYfUGcPpb4xUJ0wFEL46wN53JcTuRU2l
EYmWz0gBaSAdztSZoeFg9AJRWOy3clN2RZCydtYMH8ruUySyb1jT8c7nh+mHTwIlrP7hpQ5s8Ekd
/ZkqBnGXqNnYmClUcnAexEnNo1UpAILCvJOfayOFCB3sba+r6moLjSkW0Tg6E9Wly+u4Q9w+rSHE
7ak7z+MaGLriwDHRYLgp6hZ6qSUgdTSFzm6HvCNOoVbS59Hzzj1sYtfP/SO8bZ2i0QXnEnSNd3RR
MVC9J4g+UC4eDSHTbTabygKvhNjoC7lhAo/AekhzFLm76lK1F49AIP/U5HOkaAlok8fKc9otd9+M
WAr2YhJBcdfmzR/btzHbnVVWbrQKGyiAQeFi53jMcBjs/UPp9zMKrx3BTEW+tWhIRYB01V/fLkLg
6mcYKdStDuMFIUJZp602KXIY2B3TGC0Sz3PslsG46I+0lcbm3Jxe9q30sCPCB5rYEfpQ+0yhugEz
60sYA8C3UWHJMNGA4+akpRkBcNbON2/syBQaEQ0EvQhKVNELNVVcgGA1Z81S5VK69YuvLw9iVM6d
VK3zkCKG0mLh26CXXWljHVwgzKuwk8CW1PTMJfMvDUsa6PDv/7ob8s1BRM/L4IJigbVYnQgnS7u3
mWNbZwp04TOUxSKPzL0w+/tIQ2ryw3R9qhOC+gKCja7KAE71InA+zC+SLuevRAgounUBWBAjyOgV
4BiVBsgcU4CrlhNTmde5GGYFY6jp2/UlngP4WQz13kWIJhiilDSkknMUFaUPeD7gE35iTRTnG/3l
Enh0UOmcidTW87DpnJampJxyOUr1oyYmjPAW/Y3KnSLIXGydBwN4zjzAbm99eXoY1O9ecJBi9R2H
IG377/oEuiYhLucCqJJ+tchbUP2bCvwohtJ1Dg+zv8lmzub6hx02tQDEBFBBGghRyNS3KEIAuaaN
YR+2/pH8VLAyQnxjBnQwUdf0NT4++9MgM8MPo2c7Iq2KuoLYy+iAmI+R9X9DjPSTXKI8zFdC/WL1
Hi/s+ZuXjyTlBg9ciAXwg6eJx3u19rpqfa2aLzF6ik9lqKKeGHD8+810vYhTVv36GOkqNQmLphGv
stAr05Qc1DwnFOpuScLfy9w0ZgBiYmL8eXaVF8NgF1piT+I6if+W/MZPf2QWBGJTZG69diicE4PV
sccHtHb+SgTKTNXCF3b8cQuzprlT/qU+DqVTzvS+1Po3hBKRslHQwZeLhEb4bp/WUyRKK/5YwLYp
5mPwguX5Eyc+tIrXtwFpllr/g9hFpC+HmaTwQ8WPtDlH7hsXuG1H0T3Q8B4EYsTvPUjd5YaScHLn
9rSroyUGmW+EK0ODKJaSDFX6ZExTg7UCF0K0HzsA6ERa6wQj6q6aqVWJa+oZExwfOszhm/E2o3AM
F6/W1mPZmMHbx5Z6YXMyOoMoIz6B4HaHevfwyHDsa/Hlwq5FpUh0Ud7XRIqmnrI9VkAVW/04YaoP
Yxmdw4V29qYw+3aTI3YRctJwyGBFlVSJ5pKBQ1xD8Dr0KKHz9bv82jTRDk+Sd/cvEYzmWbr5bjh4
HrzqaNrN9XKcyAwxefYQOZoMT5m8p7kcGdoF7R/Sn40ECr8Wz0P9W3tszPCnHJUcEDLDVATQFuaf
pjCLITL/kTVMCL0FMZXAS2aNRTPKqCkKaHwhvArfFs8w8IybJQgzwDICRfLcZx82W8mm+3NtCVam
Pff/iQu0FdCR26xZ9X+3qYQqVjl8FSTVELcpZXky1WUbQEYJCeEPYmSwTOkriX7NgJHByB8vCoR+
Em6eJ/PuHlLvYxDbO59ujc2uBg513Y+qRPSHDwdSlTiXhigY6+trxvQLnK0bnd7BUdRoYqjdv2sS
bRqavmqKFY7Nl1wvLIyY+otoBKqLWCtV5mVjiG1vJrC3qIxTbX8tDR9JbsZc5jF2B/dI8ldd5DC3
AJ99lq4pHoXJPv/meaQJ9v4sWHmDU2wMyIffTw2XLuJ+GInCKNjc04CS2PzjaDCMdzBI8hxSemtE
EmCF7I16nXb18N9TiFuFbJZmh5uMkHSJ1X3JZpvUd4grcgELc/Cce7X6L/3ocpmcttLetJyIDGCX
ZccnFKT90R2mKX9s/ZtOhB5OOSGNu9qX6CV8pSXQhLhqUq0ILc0GcPypI8tskE0322f+0kP+Rr3d
Ospe0914Z3kuAHODseei4zXRJgrFoJl1Tyzy6XdlENJSIo2MYFgdCg89XoXPNySHmoCJSeP16Q5R
9lYaDC7kBRXuN0cwg+rtja0giWpdivOTEzb/okyv45NTOpDZRbWC9dYU4BQTY6m5eCYsUYFFQ1Fv
1F/KUWd5hymdyQryAfc9DlGF/MDS7/qslrb5qRz6FMWw4PMXOXhWOm/+IZ3BP2u03exzW8XarK0h
AqNfCWpIuSFRUmaSAful+HmYLQ/Qp0V8vrX3oMVtxuZH66w0/TlE/tId17yQnVkzCk32EUV5mx5g
yQMwlunhNQKhXN5pWiIxT4zccO32hiSsLgKGrPJHXH5URIH7NPNEl4xqcdqNkpgHB6LsIJxWiMEW
TMKgks5A94kbosrza7V8hpOvnifTvZIvO/nNBNrtHG9PeW/BEExm2B3iBFONmrm68ZeTpnUR3OR8
9KNpGEFCE8kaFAg3RAieOHOno1rSaU7X8wUC8Gd1FGD1bpooPexkdI9wtveuYXR/ygIv5EVUeHM4
pn8Dy3FgO2HIhgRKGkblfRMVQ48Mw+ZSsp6Fbcqd/chNbglbEioZpW6nNUFI50oGxtwckM1xGjUL
hDRNoc56I/7+9gZFb4qamPu1M/yQaG3fzRio2Ip6MT0JiOoxtvAncPgAHri/lfZSddttVQoraVAv
xm+b+Tc/WB9FBMbzceQ8wTLm+0LYxAnOLeT47jC3JOVnY/ncZnCg14XPKJoVY0jxZQkLVvM8QXC3
m5itjsX6AYF9uAvSqcCDEjGwc3dH6a7QVzkvuG1FSHjYiomTylPM5zpC1B5rf5dh8zUFIEHcx1Hh
9qeZdu3rIrsajncrgd+INJ7QwTQSlHZUOidrnsDb31JFTkT4lM4Ej8ztKI0xP1dpQXYKYn9NeTfx
dJpM7ZUJMvCT2t8XiauoPOnz9a5RM+r4OgXLgSbUuogO+8tc5QJ1S1Pd3Br1IUB+tQGmU9BjHfbO
yaE87Kk7Xoch+GikrQg5cp0JuSjFHhwAwhpF1FkHAr9b5Qr6ZCe9aHptukIBfzgsrmABvNzc6tGG
NKIYxBokI6XqCDgDQ3pU8RBLezTzmiqztoupWmm54Q+m6eoOS1dqgXrkK63YWwqABqxXxuEE0U3n
Ud2w6+RdPGy3/CaGCtCCK2Pr7eF2+DN6aGmtS0Wlj8G2/dW+c51l5Qq3yA7ueNUkiU+kxu1k1EsS
YOOSOth9USj0MQ3Ig4u7O75SHNaXtUYoUhn+xVIZfO8U7jX6/dGnqsWthq50LJfHfa9XCHyTUOVw
8mQBSCgqGa4Tvrc0MD+ezpukxMfWj4fUCjJfpVpMlYTHPSTEaO+BIsY0raEuEB18XGXJqY1aZidt
hf4i+aGzuVwij2kogNYNAE0uK7jZNVKZdKofZznMOWX7anz3hZGobHHXw3ha8F21iGb1W7SHIT4m
LoG8EIhTJM8NL9fzSkluGZktGr/LlLlOR+3Z2AwAjJDf/aijSpyR4Kenuzmvt6PFMXaJbTN6q36l
YO/cWEFbkmCv25mdAdVj1mq7LYcWOhQYXhPvufqXhkKcuzmr82XbcnfgTnUIUPSEoCmnKS+dPSzy
pbqRjE2k29XFrPXHCihSlvQNbFtMCL+VZOz5aOvTfZnpWoT9hO9APwSx5wfb9nyPkpM7K0K4fdqd
16csJ0rY8vhWnE/vKHAQibIvBNo4hSpyIedT5IlOO65ulwALc6uipznbNuhF2NlVglJ3dhG8URPb
oFUVEzKfA7MJb2MWHhL/4NWak3YBuUDV5GKwy9hw5J5UbGtyyzSYVszBHTjJNavF/8mma8JD2h+B
v5oa8F6DrXznWyCZRZ2mZJrPlw2Kr7Sry8e+kT8yEjWD8meV3JkufCThKuLvjUlHKyX5pyD34xVt
zC57B5xVN0bnkTmNETno73XZ0rHydTur6BQQpSaDAe24y4HfbocJKqYb7pU+7mgnJiO0duaal7hB
FSfg8ojdGrFe5Kk6BQ0P7WpaTS5bfM8dbhaH9K5TK0hvWJmekJjknqZp//1tsYgnP0tfDWwcNQrH
pa/VgRF+doa0lJ6u96fUC4oyR1lF4Dsz0chcU8S7LxJVMmCfLq5Kzy+S4QFbYed48fBlizuA6RVK
IhyfPf/b3i4cWPvz8JA5mBZskAs45LLO+WpE+TEmW4JjlcUO+gTIWYa3DpogW+Y5xEDE11Fj/hOV
9Rr+qlQ8nJhsZrLqJ4SJbS4HB4GaWXNsENA6cU+IeejJn1dMmGu0MCx3eLwan4dpIvbuD4naJjyv
JQKnTB7MKhRZLd4m98e5EYGhbnu2aXGrQVepK9tnWDYTQsu30ky/RS6342SgDkooUkYBTfh+tVqO
03iaES2xp9jiFh+rDrq55ppBURhKviTw1BZarcEDwZKty2C7blUE/K+0P1vI9ZEr18WmzmRpVsHJ
KHEtPj9FKGU91ioVeWQ0mXpzdFdVoW5uGoQrEmZKISEVVdvuAeyzrBvVFZFqYQf4eOA55+xf5DkN
dsc2LByCayZ5ox6J9IcrxNIHDtDJe++Znifu1Zsja54zjI0BeZ/aBHbQGVL6H2e1bC59YO61Ht0x
Kteb9n8he2gMhcYVsigmI23mxpZ8NRpOB1q2ViAy7Ec4oj87LvnXAkaSyMIHvDrOI00xDQuC5Quh
tV43UtXgTGmIrejK04xVRP22f6N3xdxeg8qbFukd43N1MxpeZqVHhf2E/GkA6bighIqHl4rczcrk
Due6H4BrtGT3ruQeqN/wC4vg6LwDPxO3l1oKtKVXr4dwV7jJBPVZvtPrPyWwriiOBw8ruonLC29g
0PuOGBR8p9UZI+la8OJXrrFtAGlFgkJbLnlLvGLREAUTjzEe8y+OgHvLeGJlEZ5mvI26Yw+nyDfV
NGng0/rRg6LVC4JfbVsON6JLyuW+6efg8OhXPoy6S6/Y2tnHIGnZSo0u5p82RAl8FO64Y0Ozruc0
Je1cmsMm0ECxu45zrLrIqF5VvLeSxfVHzUW1/SyNrxLoWjh2Qc/TmlikP4Z0dCEueZp9vhR3nh1x
OiiVlqHeg+A/P+4Fiy7XZMjEUbCtNOXtuxFAt7AYxYXWJ+E02kCrekSCApstdVLhBYBvX0sEO381
XXeHKILkfA1QDRYRcw+LZEFZ4Hd/6ru7q8F4s044X7wctxHBig+I+07/k64GPvg+MfC84SpEdlYh
W1duVE6of2QKKZI7NaHtiGJFnM/ZHoKpZ1xRtJA/QYjU8CnTbmrFcI68jZp8JbffjtP6XnVEJ+7N
93GkvykUTkOxpyvVdiKD3BIDz4YIfwRg1FXlf5oW8R1D3cPRbNJOiUivMcqOEJWLd4ItlMTLCgDS
u9Jfl64z/bqPuvY7RWvNCp6kHiMBEHWuI07j31u6KMoW9x7hUfPtGm8NSJHICafp+gAQ0mCVkFhU
dwxI3bdYbIm6A7KHWupDw5bbp6CUxb15c9LAZSsOtSekD+6D5P+nDK5VYzFJ6yxdDwZU/9TPHCMi
giQBcyMDFEc3qKYYfRxbQTDpVBb6uz6T/iGVwaM8Bt/+1WsQwkwilHlLEX5vUgiVisNJYKRd+Hmj
qVnYVTZDrn+cCX9sAPSTropjQ3sAJYvMd2U9J7RJeac8dX8k0Xmaiuko1TT4BkaygZid8LScjK3P
XsikKINbsn8B0bzKscFTYkJqa8Iy281BU4By9mO2I8krsD4+wqGFscHvBm2zmjzpG8/BEZ/AGaWG
Nheod4FUWYiL5yKzWetMBDkq5YihdYhUs+nWSoo7jDOxJoE50LSZuKfGY4pkpXr8OfJ5qxTu/Mgd
EscqZ5HH8KuWg9Tj1xu9HRU5NPFqCjdRxiqx+rmg8RUaqjeyOlmTMXl8UbiCwPpl7QReWvQrMJSK
Q3wIR+c7i1ibhbH7k+Y1agEhNcXQPJj8LVRB+Frhv33QpwCuPCUvZFJDnqqayHoOQ6CKLXd9HPbb
n+pq0pZ/x/0+0J2KiTlZZEkC1/9q9CG7I3BoqlxUmA4go7gxKrMWs4msnFYI2NBMqJquJ/ofLo/P
m2tVZyrG/w9yGdDXT+CiV0xX29TbVFb4WBiRtzvCu6qn3fRN/fHeW0eQc/FQoXcyIaVPwUhunJFT
bEI3W3EEBWiQMvk5SJp2/050uYdSn4GK/lGyeOCKhr8Ez3bKqsi8mVMvFI8/2845fOxPk2LCjdOX
bNcg5cwR4/LiZ5Xyc+S0fLNVvOyQ9rjHxaFawuqOAzhrD77Ad1r4N+WivhgjH6oNIbHV3xa29FFJ
+zBjBv7iLy2vsoYs8DpE3gVIEj39DrxO4Pz4jW/V3QJCXy5Gyk1ByhXW3xjX7YTxadrTctal4oMS
wXoZnQJlcFcQc5eCzBSVBqtItI602znCQUQmobMa4X39LHkVcjPshMXLQ0SseBkHzDn+1lWCHG3I
oylFC0ZgWS3jdy/djqNtvmCZ32oOFSnjb6KW9GRW+TABkdZPEYnYB1N/SMgDPwVMEK8WFtq5RxpV
ggxLG04iBoUQsxzm+P1BPJY3lnFV6pL+Fw86dLISxTtLFSaZ8McWFyJwj01iyd0ykRTMe8keWsSR
2mietmzPkrP5XZ/dHvTEtIih3mBMqqYNsGKPs+quQ5r6OfTWwBXBhbkMPobjKMF0Wlm3GC7NuuEd
8sVkSL9Gv9C6r+0/R8r6OH9Ohp9zo0Z1qdTI5fVUlN/80QfM8MmmTKSUhRrE9fkn2UvfFH9cVu/N
X5iVs3MJyAPKkDHKyNEpKi/YN0wDl64JkvMAmq2mDIH+AgFhcDvBKrEyRPxm3bINUjCL69XU7nQh
hy2UvQ0olJsF6FH0yI7bZzyytrfScAbcPDfmkjKgoJzL0fhzLmvbJsaCehuTiDzyaHOp2xTs7Ivd
sfXMscZSee728YtPSV0AKW6lqKyTuehWmGmJDm+BeyU95dbHHS1baUAO3pRim2AvIJihRdsRzMnM
V9lRPrl6zxqWERlUtnIfRA+l3kcXBfRwUv++Ermqnf/OUWXOkwiDqXOPry0OqFEv2B8Fb873zyAZ
CJHlRgJnCnEFTZVKkZXEZ+9uli3zCRDqrkCy1ihFfLwI7NXEP4WZ56y7B9acMaKvyOSpjU99265Y
nXhP2xTSjZ/zDCGCeiNu/LMKJvtEMvD8jufYLye+WkJDeqLk7u90YQ3N0V2eB7RTJU412n++/Sw7
vj9fUbBYEIMFUDQyj9N345KgInV9GcfzWUMijYqzqy2xFFhe2ZomqxUzj5P8D6xA2kszqJeuFD9q
H2EZU3JEp0foIMxFLExcXa9pgw7d5gNvWdCUrPKJSNc53bBVgsjEtV8uzEuvZrG1J5OTA4PFyswR
9BVUGdnBHMsODv1dCuEP1w5z6qkHWB74JTiuka4M5uQhtacW/miTIiNKU/mxbLOHvIZDY87Qp0e0
qzpYTNYCYhv+EEpFuZCZbgnVqTbMkUAFEf305Z7r8Zf8bxgYsBtHoeXp662iRKbQ6z7+p+jy8ZGT
UibW0z710WOil8pEVAPnDAS6/6ECbij8g8ggOn23ay4Hei52BMomuE1l/4bBoNGa+a3bnoYBjo7Q
2hD5k22pDckz7QJeZAbHFxelEy52sw4rwSzRrrUk51debVfvocH7ix1Dm28e+/UmhaadrbMfYW8f
APJiLkk0UBBSWC2ym4uFP+Z3trZ7JhO9HTLNo1fSDz7BwWwquCnhI3TFvdCOY/3fEmmZBXrZnCqS
1sLS0oGXe2v7ea1sINga/qdl5UNy7LpWpanggl6PRprOaNeNVwzPdJSGqJwhBYGWjIT3nIMfQbBn
RwwxEU/Ae4yU2EekO6A7D4U3eCYh8fhIcRIRXAdzKXxOh02PCaY7zejuJP5RX7uhJo3/YNVJ6WKn
NjJBt53MJUn+FpnDd1jlVyT2jZZsfFsWADsO4WYaiElvf9DH4ABWGpcfhn32vrje8fVgHBygqcYq
N/4Rt5zvOU9U7xIIshXadKy/MyDPxMxKf9P1NeIFuXACoe1UwLi3YRDAK9PneCC/qRlrGbC2UVNq
EYkZqqxB6gXK2YvyZsQB4YaXQj23PtZJS0+mSyNbieGASPVGrxTOYj846gLEbWMzTin4g3cy75hd
xD5ohSWAJC3xcBM5uaFNJ+wWnyOMN/1rIjz3Y25Lq7JojVIP81m9deAi2c6se+DjnzIFTlucF4u7
S7BPoOZLnFuP0iaMw3Fkx1H8pP7ZOoVPGafV2e4de664u1YSkZAJYSSJvJAFQIb7wC8FfdaEJxdK
hq8oHFQPmLVFmuS3OiNQ6hjtvreZxkkmbn3mLK/CoJdahR4j59czmRjmzFr62+pSDP043uHdDoY7
HpBLfrPkUWnY5ZUSoZH2Fntv2+h7XqxzWHqXGPxyAY7wiupqsErGnbhrlIDFGTqaMF11DIuRGKYs
gBC1mA5y4xFzufFbjv8MNrYBJbls1C/CCr9RCAC2a5Z7vZds/7renBAnwfiGhO7wTI9x0cxMALHC
uvUj/0qQa9/kxe7i7xDW799ZXHmJzYpwxJF2UAhZl71fju7Eih3CzY7n8+yDlw8qNY/r/+yYcUCF
L6Ydw7vGxMVWdEFTgBqp5HBA2EyhijnYyaAZEEvGZNuxKtJhIJj6K/j2fNbvyNi9louZtmAYnHUV
nKSbVX7ax2Ng5v6WzdtcZAuYnegPVgFuzjxh/GKQ7UGudH/G7d+jbMPI9BO0Ni66IBPform2njRv
Tuu+MW/RupNB0GnsVuX4eWFuNpd+ub8wyFFnNJ2pskzviRly9aN4vXT3JReIEZVXl0qUM++uMzxb
mr3niGGRHjNmPuUbxge9xE4DtGpJuQ2AFiwJZyBerCRaKeYydwhxYfNKFjK1U5fDatL+L8bb7Lqo
DDqelZxeYgzqaYiPhw/Z5Y6v/t7ydbalpkvkGwIQO4s0JfKdWOUu7ZrjmRC81dUC+WCBOnfnbD7R
V6u2hfyZRXEBSOFypKGsK1Z2oMQijBa7J0pKzxy8DF5hX0PowtgffOZZTjxdeVMMsBhGQeLYuRlj
CVTdP0UMBkiyfG+xTRSE00OS1tilzJgKVJNjKbDY/NENdp/U5qeDM9I+zPi6jJJvCIm5vQI7lzvR
o1PlXQq63muhBBkSB4hXpTlaCd3j9/fnLUk2ia2fOrdlT3ibMmkMLdi4V6lLZGZ9Bhk30gz/z/lM
uotbPzibwEKwqW0dO7WxHgO+6QPuU6AfbPxN1PxWkDzzHa6ik5AGznq7KR3f1Q1Sjx5N3WFIikMw
fy0OQv47fbeH1f00VuUdnhg18+fCwQuuCECOy0MGbLAQnrHR4VTp7dVTydCgPt0FHUdR/XvNXySg
3MnqRCl4i5KfzIHQS/YBEb1DWX3xoXPo25ZKm/a2ec12TS5LvthU60V2kgGbyUfgGKO8kvrQqRR7
kUxgtfUrF+c6Lfr525NVpZ4BL78LWebKCJ1lWPgmE713EbndsjuIj+1O33GEABHMs7Eds7fAlLHk
1yFtVn8TwwN4bruSzU3HSgjpoqz7jKY/j50B6224qXZbrEXOotvfA1P2egVPGKRHAgOP0hJwLkl2
qxp/eYJrk61ggcU12/OUV3/SnTuPXU1OmPXz4X37TDx2jKnzaL0Dh299CEs3iGmsrQYcj2XBlfw4
850JRgQhxiTyijj1Kw7J9/pXirEjr14yMxav6wIYPcAL9wiKGF3lefTFWZwqN+U2TIRZ/45u9cVF
6cdffBzTb9eej1B0/in3n95HRWzD+BglsgRn77zDLHosVhZcwix+TCP8ITzaUjKxkstoGg5m361D
m7q9LlvOQGvdgzLPZJvYf4/Yv6550VVDFKS0YjNOZtih/2qbUgP8PkjLIQjHWN6Omh2j+hRuIfPO
H09wU2dIiZeWhKvmuh6YPaud2Sz4bu/AFUKE/9wcuRMnYJqKFIEZAZuHk+wbmd06tFjkSpBmfNRB
a8whNmgpJzRCCe4JSCrAmV5j7QpMrUWbHF+fSdjnDE38/Ns4RY8L0MdIX5MSqo29ZEcrhGOKmlUc
gRQxUswSdv6eChoYfXu7WdazaOWkv7EmwQk+XMqJQgTlL5LaYiTxHR7MrRNG6AqEKbRB1R6/DwHY
oDccNs6J1uDDJitm9c9rPqS+ksxgF4O8oAe7IMy8kEzdbKTu+FlNzHKp3xFL9RZPNcQkXWpitw3B
Ly7C2S6v60iWLIWbMAwVWQpg842uaW12H6a7VSrG3cgJFr58KRsurEXCBFYGwkEBeinMj8Zmq5A+
m0D1RmgAeH9DOia5YpSFjOrI8h3Zb/rfyEkYdphJK6Flg+F74ny0SL5HCgbp+GrN0fVekdMZ8+Ub
mvHeVH38PTYhrnF2dpuCydblmjs/VEJQal7Aokg+9i2xhfVpT4/qSQIUqpZDFZ/uphqkjE9EpH6/
wZJyAuRi8j4LdEiSRU7Xk8eISnQpudrgXs47IwzfewiFpY7M+gPCyv6NXUAJtHfavMTzrN5WukNt
GacyH//Pfjsv5udcjzBv+u984bpCXDyNUSIC2T+YEUro8zS1D8BK6NlKRU7/TnBeOAlg60IEqy30
dSKEyFeqf0KMwGHfA7qpWTsB1Q4TsVoDzsWnoz/orRDI8G/2khviaLh5BHtcRCoBzgi9UpXbHxSY
YzEbXawfjoX0CG3nuWvp6fvEpe4Y/xdqY0DqzJhhw/yHqAZAP/EMpAs7c7RC7ShSvI2z3Sv3/IXN
MO7QNWtmjlzP+5kbzFBVOQMjVkZRHIiIHDuyxnDfY15ozMNr5s5Kqhy6mK9CR5lAOhXvgMUojiQ7
wwa7njHWq+sUUP2innn+WCht7PKRYTp8nDoidhbEk/qipPwZFm6iiaptHHHL8gGm+ExTPIprF9ho
nC4d+ekaONU+/PULFnA6OlbiWVBn6rzMpRG89VV+bb6l1sV0ckW/BSRRiVKB1a2mUhcdsABDltW2
NkmYg0PmNZ+2s+tJ05jwft75RsYxePWeHh7goJy69+arXvGfoSgqNdDI+SpiLwC9W0FK1qCXEBRC
H1dcucg4PjtEqZkQm77cPm7vM0XHPS6j+NykNInA7WI7101JKNQO9jpiCx72xzQHdPZiDE/TzeVx
f2jYBk00J0Y/3vwUf7BdCbFMi/XH0k5c6h6SoOw2+ykbgzjjpxi0zVCmkDs4ITwCpqmNJ+Ym0G+B
BWj7Sj0oSX1VaN9p+ug+2Mqb9S5eVyYZsTO4l87G5YGMgcqSNwJgIolD4yQEvKNRvVEz87xvbFK/
mgyx3IFla01/hN92rqKQhVAjkzzqdIRCEgnIcjGSAnf2mqnInPboXC6agkUJwJYKRATpZg97JxCc
8fhCMgrglpN61/OQ9mHYrB+LKPb3KSIw/m8HugJrRtgmbC6D29E8gjQjEJqYmYwcsqoi8Hyzg65C
MBbOJ2qvtFMhf3xwjflqXIJdIsg3b0iGDb020PNqzDuYelnsWyei02Vsv6ihqwsoCBM4YmiPAy2a
d4PRTIy+Qnb4FYnBWbGS0k+xl0amgRQk/lXMTxv4eNnpAZpL+kuxveqMZhlzQ7F11gcHdraioaoB
gUVAmsM0UrVUc1o9UgrFgts2vRGb22DE4uxmmgwyS+GA+Mcxha+iSnXowc2pu+KWG0U5KhDRK+kx
DKzMSi1N2Im5bkEzE2jGHQVh/PbwGRwQkJqz+3emI8W6uQUOp+6mYlHjirMevsmE5Ksimps67FCO
WWcs3fJ6YRPjdjIULr9vCxiGgTdPwPnsBXiqbjgSS2LjbRiJj6xnXHDOihhz2jMwKC0xnUZxDkTF
oLslWGb/54OTS1vMs3Yx/mHnFSvladWKKtmC6ZbeL9ySlItBrfSN4X3MD1aF7MIJ2VxspxJPEJJn
hpl/eoUeffV07J52xrW3lJZdz3ghHCJjHSN8QOAXao2UeCL+XFATBXAB4Uo+rfjAeXAW1stE4no1
K12Wd5w5wK6F7B2YxOpNc7B2X7LNob47gJUWOMRP6mPLCthAgJrob9Xm5p6M+vplv5+2eqY5FfDU
lQzrldlichdgTQTnS7meE82dYLN7Zc12effZqaNLrRkVeJgTXdWr0OBdMHfspbk2h/VW2K+DStIa
oa1O4MaJTvWYK1N/08yePNPBihox1P9bONfw1xtKSOPTGi+eT7y9a0AWS8RzZvhgr7fVemli4poy
ACpPU/aLUFI3BUo3ISZmS6owrqIombN2IPqz1RT/PPv30epgWxMy0Srg6oloemVheQa8jvLz84mu
55jYJryJ3/t/xzQu7KCWu8fYhMklZXCg1OjwPeNUqdUFRhM46Kjpi5Do8fv0NZRhkNcpM5czZPZS
YFp2AxafyuyjZNio1TRV3Bcr2QDz+6qtci8MEtU4kl5hJhp6CHz+vvw2mv1C/LzsHM8+TZMzHvd5
cvEUNk7zxG3Es1CMfUZolLQMpA/ipdfdlwINe3hWxmXdx1Gk2g6Yihl43I+wMxUUzYDnblS7mDyN
psWSRfgqujQudCpS0wPszDXFpmirk4JCWlM+VeH1dv/SPHNyRpolcJvKX9RvDTFrNO6VbN6tBT8C
fRQ3b82DFwvmq6ZU+fCobziMpS0B6paUWXoXng41L7DjmHKnc7kHeZ9P5NOSxqzsfou5odgvmLpe
IL5kQXqbGIwUrWvbbw6a0hWMOITvlwNCl3kElUCAqlbh1YjqspXSTwVBN5Ea9mVUqvlDKuOgYBKV
ITr9MLokSKKkPbslMN/1gO8m378TT7yHHZWTmrYljVgsk7IiM2yFfTeulZ6alkjUOyzH/AqDw93j
vEsQva4+3SG9XDPhSXee60xGXdQtjj9x2PqXco3+atEGacK3dn5WSeELOAyAVYZY7K5/+ARKWquQ
GDxC6Z/JALOw8/GRssM0aXbngmr83HaZZbDAkTpDaeqfl8it7DzkjzZ1Qlvo8WwYwIDwnu70ElhH
Z5wgXtoBJRJgWEcQgKq4Qz0WQr2ySA/HGPVseAZMB7CYG6fO1xhl3oFb23i3VYAoWU82nuTYp7XQ
VM551tkt1zM1iQGzDzRZ9JARdLtPecUzNTPxMTYrvYZWxLt7zRzRN2DAcRXqqRQp/sY6B/OK9KxR
+ORQ4ebCM4D4th/YPZAB629YId+BBblyk5zQLuzi20cmvRJ/Wa/6NP6+KgeI5+wuJVpiheLX45Zy
Q07JlgV8bkxKse0QqU+1oyzQqx3nrE2oAvrwsNN67yWlgTqEXcQXFpWs5riviCT1Vlls6n04OXUK
0YAbYB4U8Fbb9JgBoHs/xj8J+KZWdPhQpmYOHwI0ddxLyy7kM9O2RFLRTq8T/IaUE5CgwBxVQdgi
cCZeYaQDFuVzztuEskUyj0iNGXgQKT2/WPi2V0PEpTxuAX23QLOB8JY4Mwk5CB59u10mP807OCsI
38LihhIsO3eKk1NmP2v+1w6zqbMY6kosuKIRxILmQ/no5XrVBcl0KgTjIgVfiI/oRKFPXWyXxGVL
xJxZLHMGpTlTipi1mwYGIzLNqH10w/G1fs4vQsDg8d0P7Nx//Y63hQI279X8k927Y0tagIih+Lqv
eFpd/WeY9u5wPVZCHIsZS+dpHycT0bEbe5AGJjHLpH1eOkCg8DlgIpa8b0+GRnRkj0oHuwzTV2Tf
OGcCriVUjEihtPp0UPAWPpPeSat5HLnZbRU/XLBGclV8rl1jRWnxrkduElUAubqJpv4TpW+1mTup
lWTdAimosIBP0I6JB1y8l17vFcRYizwIvaZKj8gUzMFTm4v1u3CJePc79pQtDTATwbZWfjMmhjyw
KSzuo0zL5NSNBUB7sgQ3imkbrCpPJXT6QiYD55QH1ZPTJkxWDUa9usRiqS+iw8jFLpuJ/IMAVcSM
OLYlM3b5ZoLLiENiQ9Cqj0AVmjTQmpLPZAKeEbVWad16nu63IxEfqDHJ0Bxbq0uZ7SnuFPx+Pkxp
tRBMMIJKxK6A5WO6pCNIpTPkti23hao8D9irRys7K/EXB4XwPpobfNMh6xIjftfmSqRWeTb2gOVL
HtWTk/xbl6TWEGSO2b5dXv8CW30W+XQkPCqmsetsButwYKIRR6D+L0J7gJknST/PuP7bjELdjcV1
JJciksbkqul57LzW4++gtoQ6HgxORnnC/h6S1Y+uJbnj6U9ev5qV0kieGMucP4+jkUBopGcSsQtj
Y0ybxzqUbkGLsjqwb6ZeG6+l/E5bm5FJej5idAiIFrVUMXMuwq6j0a3dy9WdN+3Ykunahc8OFme+
h8UFBsVHwb9u/DGjRocoU1/6gMaj1Y7e2q1zKXhBm9qpDrD7ngCUVr4WaufhRFizZOP/889lsga9
Jj6UrXAtZa3SRLE5HPOZ7bXfvoYOy68ASLtU9slXOlI2n+QhPi2zUAHPiTZl7BDAZ0TPsYNpAWaD
yBN4yePKz4YW/mpBRRaLIVgdC/hZ00SXm+TzI96p0DgOwk0SsgTtc55xKPOuD8Q1LfGycmqUfl/g
Hk/xSK+TUibAudNDjolpHrGWSi4TlfH7WrNNYQazdgzv7gqCrvyabDGb2qD+vGbvt6Tmc/p0E25w
01YtoY2RQL09MyI82bLu/pLo+grKpYgGDA+OWpF1Z99dXieo+oJ2rh1p8HY4oin8vGZv4I0jH13g
48GBCvO3JOhWeHiCmtEqI0hGcI/opXntSTk0S4ORH/yus3npjLcbz+m+QtJTgTJk4napyEl8JvoU
QTN71jc11eKxn/SWqb98rCccziVPX/a9/BEvQK+SBR73K0/GSBVV5ZGhL/eRaw1rGzh/HlLrGdCD
eN0G09VPXLC+k7zald5asrEV/plULkL7KGhLEf5RUR4nciUG4ue5rFwlMZxSxD+6j+2rz7tSwTGZ
AOM2dVY1slPlTr2iG0lQs0j/fhN81KtE/2+ufCfQzESP79vMDF86xT/uMF9Ya6scASzGsBRwAQBn
TzL9sj/GCPx9MAmsjwOso4hcTEheeZ6lsnWan91XmjZRhpqMzxnAmma1s7QWLh1LlGKv7MfUvS0P
wSVxsahlYINWMh8hFjgpHkXTMUnD+GzSWVGEEeMTDj4O0DqsCdUa3B+IlWp2H0NlkkoxRrJxQH1i
rZt60+O5kSf5S9k/zMlr89Sguvd9orkimt1ON7M9LjlKXCwn4Ivipdt4qDgWJNZOG2N+NORMvpFD
cnuywJg/SEPP5XhMJ7JP0SoMg5NHn2YqBJLx0dxsXhL+gYNAWNdaD9QULcFZnc7Gzal/VJOQWNwN
oqWc+3nQwrviwy06RsFGz8QoXSC/AD8X4cXes9zUZaEJaS0NPlY7pUbpeRHCnRjIzZL8v/B5VWpv
E0PEMGzgTSTyDIIAU3FeJuwllmp5mSjAcqJF01j3M7CIIOy+PMqssMxwnsmvfZz4GRsWqCEXa1WI
XItN4ILdgCTDlxu2AjQ240hI1zdwMeMFLLMKRhgge5y0G6l10l2c+dPIb70rWRTleDF5wM5/AT1a
b1+yb8oJm80CERvSe7QClQjyZEJvFauJmF1TG1BAEzij4T+aDlh3AvF3gVQe/r/EdK8ue9BSFLIi
t2IiFzioFp7B0+LNWV44qGgotdKV12cRMfH+nA4bddI8sUJuTPOf2cmT3XItYuCwYHr/eImEC6b0
bTS6i9ZRfsLRyZGTCN1yyy7UQSWIkOmSvvWQYJMdNvVKL3RQ0GcyjqLohrjU6L634ZeK4Twobs2F
V7/zxkfVhFlt8VN+Lbp17hshePiooxT4qRsrjHLmXhD53WarxL8+TJgISSj3yHpVPknipjuZH3ka
jR1lDK1xvEsdIBp9fHiIc+Yiu9Nb6kOP4pjCd4Fb8k+vc4h4IZkMqRq1qFfDWlqg6u/XfHA+aNkd
kNVV6tXO65oEdPgXeSLPyINNjs9CH7macBU0mxvyWkpZgV8RYvA67uVHtuE4oR8yeTxmi6qlfHet
mwyuwAUxoU2heUqOAPQwzWiMyeCE5vONGg1IYXQkSlBDTGwytfPhmwvykD9iNLFzpqWDRCx3YFRB
75e8andC2Q/IkluY+ENOsFUsc0P5ksNAh0Xoo5/68hAD/hTlFt2sQH8LRZYLA5A22Sp/ZvcBSlo8
aJFkZyP1Iw99exHCTLwzZoOYxgRCl5n8wyE0Sk4IW9SbLEtoukDkT9vi1c975zaxHqq+JTtrNWCt
aDYupXEoyojTE2vKbDyTE49mOh6HaDtsFs3nWDvWbq2Q7O1T4D/yf7GuFW1HREaWleAJvurZpLq3
PKZ5b8p1Psz2Tl/wqUcGHOds2LrCsjl3sNWRiZQvv6XVa4tKscwEeHM8rqw88BJPJ3FFZDfnoNyP
x6EcOAerUCrriV08KSlsOtwqBa8P0LIChVyzjZKCzkaFWCpetgsWacPUfb2N4zbv72FTcc6ftSra
1QmQ0hxEeQwAo1682GZcbLzNRgebIU2xihv0AI1XldrwbmgpB+zWqJnixdkRa6zmSYPxVtnWjRZI
dKLb1Z31Zr0KFxxgeeLHvs1eNr4V1tLwmJ2i4Li41BAT7apC6YFlN9iuatfuEpWAqPlCPnh8uH+b
H1SQnIDHg48JZ+nrFBg6WI7QRAcJoW4FqmhkKxV55kpaAZd9aEXWWPgFHWKFecV8mZChG9XAyN7Q
LC+VlHaEx8bQYg33a/r5s0F67XCzGqM9WLj36PJ1fgMM9FvlA2xX40v44btaBiOMpF30mtL88jmd
wvu8xS80ahUovx42A6Vvoug74QEmEH/3DbXxrpO5tUyO471GLMVgCwB51LyTK7ygoLynLEPhhB/D
WtkXwP/RLkPGCwwAF2S3bjzJV+ENYWtVEXstDIsgoinOM7kknkTVi9dllBGQB8odlMghNf7O3Tjf
QIzHUDiFyHSXnN2OlcqHHF48EDPW61ZecpnTPGS4MS3AAjzpO1lu3WmkexcT5Gjf0lImNfvDhmkF
2KYcgYO1KF8XgoMR1i5SS/rOHFwxIr80iK3CYdoSqSh+92f1nGWezkhZhDmvVb1LfbLN0EW6Z8by
nNRl6dXa71nulxFSW/2ai3SNCcohfArKYXPZLk1fTNICfGVUdlv08LTKRboDosR87uPxic5daY3R
+fN/UKNjm6XwmI3gANsVshwYJh7fyJL5GEvFEdgyagfGvfo8o0gWIlw5ocQ0rK0mhfgPRyR6qrgT
fNaU2cjYZC6/FGIsWB6863BCQNQfJr9tbFzUo2EKql1wrdpwUYJMcXK0u1pKBWEIeYPNVfjZEkwY
icbVpfkVvhPPdbnVkDj5PLtv4c2hBMVD+9Lf4ISBUEPX3WyA40Vg3nDEuBy0dzuGlvw3DpD8cV9G
oCMLCmzht+5WuTd3RAWO37UVABb+lrM9ekpzV0Fy/hlkW3mjDl2V49FO4hUJxuzk+TIPIh6Ippuo
/my/YlaIXdpKbeHcTh4AexkkobS8D/6GbK6L2ZUoqDDyFfeaiQo8NHfw1a2mxfG2wzhdENTDh2oV
cxB9EB9zcXL8PQEd3x4e9qo+2b7nsxM2lEJqUoZIdT/ZxMuIJmqRFoQ1kZueW9QIEyhKXRqQsIMY
RfXKa5jPjrk9oMAa8vgRywRU4ur/GMrTmWgJjBw5HEQdVtpTdNwBmrde01P6L9LscbFsypW1eT1I
g1BqNcieCUhhxpt+8fsvosygjt1h5rSqxaEjRaos223TqaTLwCXVvxroacP5BL55hFs5C3BPyaL0
qf+nj3X2jN5WN898Nk5G+ecNnfdhE9OIYsO5VCa6CWDYZyOKHMnm1xyXL56VjHkAR4Dq9/15A83/
j/ixBNYyjaJ7XGml8ZjsQl54Os5FlVBhK9gA0GpZREFELkBRrPX7vWPRWxxuY5KeNK5Srr4oNvjy
DwLqzKAP1eN7CtgYMvOtXKSNXJF+lQs4A1T03w/b3wTCZYHOapg2kdZaGGUta+zf+U5cAGfnoS4J
/J9m+D/Z2yd3Qs7yilzl6PaYTRwqGr3q4eVc3XWb+IQZTN/d2cg+MR3sfTLumczZqyLhDRpI2bKb
HUPHQOVFXbyeIbPXVt9ONf1c1nTPdnP0D92kAvThQosne1+C7LdvvNAihw6Obv9xaSD3rshR7j0a
+zw21E21/zE+H9VovHBwlBImTRoLilX/J4xEk3p2ps9gGFzlhTWi+Vd/YNZjg0ZmanCu6ceQeig2
tYVez3KcYrAhsksP7cz17exByfm4HLxbnv6Alz2vBMne1Wo5NmVzt20NcrG4PY8njHOgxgVgUjCJ
8Efcvyoqum+IWYdB4dppZOcLoNpjiF2XtRpSlupdYGUm2hWnl7Z+WYUxuJaCfcBRPFwMjLk8vsF0
/7xWbqbqWaZFJoq/dB2OZPQGl+Q3vZPUEX1MLMtjT8n+kJZvEkS0dJr3bIqpXiG2gdONYOcJdWi+
Y8pYOWZ11Mk/rbRbuLRJl31RDcXwcg0U0eTKQXlzDEUVak0QSBMGLpcrRzIJSTFT7zQ6SoT5/CCM
H0laKO5VaOLugpzlQnaw8O3FKcW1uz4QOsyEzOPaBVz6FF1e0i28wB2FrSlW86kziE2tzPgY4h8B
tq5hI/9Y9qaTmH87v3rWTIjYE0Lwy1LTyGinaYVs9LQKdYLr53oSMMaeyHBea1FSgd8Ebj2ky8Nw
3VauGtqj1a1w7rrRZYhPFMsIA66eTAXL+fo4KBjSv8RF6iIN0lzCF6EMIkj7uqW0UBBRmdBZM+CR
c0YFcDTOC0X7AW+rr8yhHLVSeTkuGUptOM9r2avmj+KJXWeHWV5CdKcraSPJbQbVsNqSPBgz7g7D
NtiNYfUu/206dUotB5WJUx1Jri6J6nA97oUNt53K/F10Or6u2XxAlS41YJYoQnnd66SNYm7F2oE7
gnhwpO0ppDfW5S1tMv0Rq7X/yEWitSgno2FDsNMGWqCuyhubYDHXzt6qgZQ1mQn2gvGp/4bcOT4p
9PzE+rRgrFaa7g63ABG/puNyihD62twRo/M8fbsR1w9G7yatiKoH5+MH0R+U/3BpES1pV3+qWq9P
Ab0BNbmxiGN9CZiH3ObIUgFm+sPiVs5zw7SkFxcfiGhZZAJYJhG+AU940SAcPfJ/7ZWbXR4RuLdM
DFRJiKQImVHh99gle5QdnznDFTF7J1iySjueNkPw/iN+5FzG750RhnLjHYfgPWz9rHKK/8s38SD1
c3gkugZT8Sh29tA8wKrIZtdsv4L4qMDflGNujDMG092ZpRoK2udGSijPpQvcGfk6Ozcjq4yVaqPj
rDu/xyHAm7JE74RYkkvm177WasHlDshvbTDVURN0nUfvs5dxIA+8wL66/4oYl75WBcrDkpTmgwAF
x1idZnJrcB4Ly07mfOXFj4DTOU5Japix0OCDL0itZpt6U9BWDUCHqmkC2TRegjzGi9VSaavj/oHV
7aOIPF+XC5jc/KpRt0BoQYsYPcV2ZR36swW2/Wfgjdyf5P4WK4Gq7ONLpNiYp/QXfW3TKGvSrE/g
pjCf7iWUZLKsgndG54zxaTNFR0X0nPnZQWFT2+ABWif60CF51eQROqwIKOO5uOuXqQ1zXR0Nie/B
qw0DEaboysLaYORKcbf2dhayIOc+VqcQTb1OS6pK8/l6uTeX/7qHPaGuWiA4SMdOHQZRorxhHYg2
V7EJfuMU8sv+DngAlWMFpy7T14nNrKSf5Mzat4+azErmpK9muTZjZiA7Qxz6ygMWryzSXJ/Zoyzg
tFd8htHqFZ2TkOtCj1p8yxl3BL/ulwxw+WjetoE448qPxZJwsGVJMqlHL8WKKOCgXPNqNNJr7feD
6vw91pgOjhJPKa+YYKfOjqRUf3LeJcCVdoEMQrczO80N9ExSOe054OMh1RWGg44jLAoaz0FWc4ay
uxKHEAqaXWfs8fTH6tvokIQZ6u0lDEfGcxkwgk9NBzIxeY2thjSTnxhb/t7Y3n0pIqXV/PAKZ9TQ
DJermra9zGaj4tWs5cNENlfrNS0N5whCtaJslVhPnWBwIjywz4+fVh3zXOrDckJU4FsdwB6PLxv5
x3ImVKJHHoTYlRG88ib1O88cqxoOtlrRqr7ZSCwcd0V83/HOXMBnunY7LW90dXHzTmLCjuodKd7v
TKzoPQOS4/NCGLiUPvNp3NGlKvxMJWfPuJywPb8727RFNUo57VXy+l0WFHFlZ1iRnEoccvabe6xc
wbb0WK0F0BeJuIoksMNCcCdx0O7VVj2OqtcyjIPaK6UfJF9vNMsXKHNcPeOuwKHt6F3/DXPmOa/V
14DmHj6nyM3tUGeJUD4cA41scs+l6fPAIy3DEkeIKyAXdhulC29LkUajyYrGHGvtGUj/N1B6jp9S
D5clLt5BAdPWuG2nF5ep4tDXiL7fytuOiGhBCvPoUl4ND4xMS0GJEukXdLV9Yj2oAqx72+5fLzmj
S2C4NDIn6o1yMkYawpDwSm55XeI4jc8FbJAdta1r8VIc3XJ1NBgVurKW0k1dfgqPEpnOB90doH5N
Q2I2P+o3hXe56vDHah3w9elIXMUmIzeGV+bBJQ4S6rM7PXJcFgWaNXjpCPPmlws3i1GldFmeFeve
4mVEc6Og5IsQU4QDp9vyN/bj/e/qBH1NIJBhYLzivaXFyE4JPOYljGGRi44VGP/62EiX+5F5w76P
snBX+tn/ES9paiRJ1yNAruS5VYjd3RAa287R7vV+UJz9mGH/59h3cNe3W3HNetSrsNg/B9Sz9snZ
8eMRS/oCN4XJi7yZcOlTa/VdvbQ3rTy2rLe7IPu5mfP0FpfAYLuV4nbGFIiNSk1LsNq276wogLGm
RO6HifZ4HIg1ll4gNyfJlg9ZrJSkJvUmXqAyzebqDJr5TUdWE+7HqVRL0aLPNQK1mv0rn1QyF3lq
g3cHyabxAnvfE+GimvvmeJCngspysrpKDhv6O3T/A7vyLTnmGP1rGKOjjbZbAIwxklLa4Rsfl3Zn
kqA8oHhPX9ZO2hlkIXzMLMDF/eQhZXgOvjWymk2lZpCun4xMmCTRqEVpX60G5Su2SpKxjKp8AD86
qjtWLy97NFNJGj+qdXJFznkr4VYiOifXq3Mn09TdsmJEK1gb5DweBLvYcFG1jdfUMWtKnKIKijxe
k2p/WrUMo54Ipmng81Ib2kUMxU7JOmLczD/L3H18aPQaZypN0oDQWYIELgIpe9Q7Tgpiy1uONMbi
K0avin1q58/w0/tAsltndSm2uIPMTs2ndyhvNzq2E8uJQis66Z1gqBhsRvw5dwMn28hbJkxSNIs4
fmmsItUTMqaJTCXFg3pK5SqFRyjVcEwL5itzyfAc5EVFCQCdZR91g7SrhleECiYDZQSVslPYIh5W
vksFEm+wOjzcltLrh0bcQtBAVCd6SYU9sqkMzzNhfSFFov8mMWxwwYc9Nzn5qTz/4cx6qIScThCy
ydF8AJfEi+p/0v85Vs0jTsnd2f5e867lLIjQRSvHTdiICIahM1gfjJyXFf5ClffB5OX5hRdUp9Mg
YZtAxIzI9KrPYDrAmp45aV4k8WfPIKHTNbkRgo7T2Bt5eJ6iiFZBTAtQOmtiFPe6czhWEZy5upWy
dIPEkY3kSjuG+tUvszLUqHpKrcrt4b/e716Ld0J1tio/2D3torjAzVLsjfuS0D6Utj9BjHRY6YmX
ytTqPyXHfyjdlOUVUBqL9DUiMzsOwRB2ZsyGPqxoDlfCX9Pp1k2lOuay/tzRPP8QYuqEz4+ZOWzH
yLz5oR6OSndwD2gpujUHBnKOXzGloc+iW9bike4UU2pqPgkDRzyqR8EeNNX+KlKJixU3M/fPq/uw
jeRgtFVU47RC7oD7iJXlahlNSpjROMj+kfLJzIPqN3p++0SuwH3legu4uL9ccwmC/xazRP1fS5H8
O1jmU+TGyEBx+zZUU5RqMKy6G1HFeP5mc7QJwLB1L4pxJFsQhd4zo97vUn2CmhoTRKiQ6XyN4dvK
oJqZGKPyhDUbsOnO7stOtTeXMH/osSaPrJxMt21HFpGusFYXcNvP0MUXdh8mIWGTPxnkBEhrLK1e
e0PF2eJmHaV8TTB2ucHoS39VwV8OFwZzKygihNbkpEO4B+D75Lyg3vpgn/hLzwZGknDYoL6z5wJw
XlD6dssQ35OSUZJO5U1dOamCX8fc/kby0VYWnHcZjU/3rVxIlnj3+GbIkjjSCZZUdHia2uIabVcb
GOtOqDbQtxYpkxvrT4MRAWLBrhUPUqqufFJAkg9JQQ1laxPAzymgmtnmz2TVn2eIuLKLCR8VMYNq
xdnmYKm+1OQYCgYddWenwHjpLda5w1YKQWFNsayHjlcvqMLe1NPGhdw5ZK72jXtyEzfiH3uQfPds
e6Is9Hlgr0W8+p/j+ZsbI8Q+VyAdFNrxYxykjnVxXnHm4rnNt+JxgvDWq/Nhd7l2bnUQOwvKhjNI
8o0pYcbSDdSP7/xBSqqsNycaKnlB6FoiQI8EVf3VOJitx8J0BaybSVqQ2/pRpoHK2cz1ydaHKfKp
hYkufoeQiXx50BAlfKwV9d4SCypXUsbOcBGJA9uT9nJ3SKIOAdTYn0bMFF5bXwnnKVUraELkwQt8
FyS8/x+tErTsiB+p7o5bSinho4SLlcLPPrOfpE6iZREcszpg14atMEe561CzRGJPHeWnApbwP+P4
JMwaH5EhctQBwpRlEo26ujY5V4weEZtT6nCAvy7dxrd8XFhp2bt63+BLLXaQ8hKyVLWRSycASO6S
f2s+v/CbyVJbcZcqzX6+DbQHYwTHl4Yv2E5KCJtbIl9MDnvjIm6/+Wp7aKfs4OU0RssjeiWL24xC
SUvZf9iCEb0f8NK7QTKY2iMF0n/Wpzx0ihlf8iZsV1sDWM/h17kbwgweckiKqiLtXCpXHV4BQH4v
e9NeMBUzQaa26bJy0slEgvtdmzEfdQ4yqDQx3DyaDhlpQCUW4iVWsQK5kd4PbNVNq2lUMRhoNCC9
PUytXctSuVWCVcLGuZBzsJNrbokzlJkeELrQKMB1tx5dy+JGk7a8iDo3KmkB7diU8M65ja7CIGSK
ZGcvErhlfLsa1cA6JJJT6Yz7SF/77/Sh7YfFOJgfwtESdaNoO2a9PWR0JdeMHAwE+/dmBd+khyow
FND6554cPmHMc84qAbBPUFPutDAbTIKUGw2MxRbYYRFP/6L3FL5nuQxPSOqW4qlo5442unrIXb5c
/XHXASXHq/tmWi9npMEj0+Bvl9MzDs/wTdNtcYomjLk9Bud6X7l2TwwxG8HMe7AwkVizqbLz9TCG
PNvqY3Lv77UYhTS71F3scKKiyEeb7FyXGhOaoNub0ME4HL+0wg1xBGdbCJzFClWfb0d9N9nkzN47
YJTNtQRauGBamcbbuLuw/a3D4XgZoZrIa9DPapiE/fNWTnpAVboUjt+q84JvrDCSq81xN9Ko8YOA
B3JYgk7QnfYilqo5dOXJu8TsrT4407j1Beznc6BJNuwGeF9KUG+Be/ha3aS7NeVqE1z8pVw27EJY
wIFqMf8H0CSv5QRuBniA0iiSY08QsGuw09zZRKnWl+OOCFeyhrKiBdJALof1QN0EtnEp6C7ZEVVA
lEkQa0oXj59eGCPVT8f3aR8NV5sbCTGFS9ZLTqf1nj1pzc0oaB6IJe3BhlHnx1nZ/It8NPTlxAw1
w8qni5+Xgv3gdkxd8ht/VbEFWJM3EjL+A/vUzGYf8iS5UpOgMIyvA6YM8LKUTwKqEp58Zj9ACDyB
EI3955gZWVNxmvS7tGe1/DXwEC6uXK6P4I0zwY4wTAXMiZQ48MP5/ZZnQiFM+EvIzyXf7fyW0TaP
MntsZkTWrDjmY7SnNkRnQtb+IHCydIjm6TXwqKI8y98MUMyAA0Gs5YPhWsJsAadkL2Ld1bIPbEFq
Dy/rjySScnsg4YO4Ab+46V+NiaC+IboKJQoR7PBOxfiNXcqOsqUU/4ICU0VlDAs10ZdEbcZiWlBy
0QTIUkIXt/OyDgHWfJCbLAazdUyL3sJMWJJ2h50F5w6roaSgW7z1nkfmb2qN6AeYtxA9JkiBmN0l
yRR7Jl1RFE2R2//Wpnkuz2+NBp2Ob9ycQj4EG4IrRwt7nnvAzDsgZicuoLWJ8ccX1nlqQ0UfN8bh
AwcyTewYNqWgDsfCTrBeVDwYQEPJRd800NsKo5t9uVljXSHmwAIPGcTjMxfiJZXJmQy7Fm/2C2nk
/xyZDcupfwt2J0JjIuLUQ3sB3s405QssIel+MpmH9kNEYPf6TNSCXsRjsVj4BD6/pEiDEkgfgwYo
sE0EBGG2/y/Utibj1cF3Jo4akL1DKYdz3qoCCiW9QwFgWR88P/TrD5mHoVS5XXyjuH8zQ/wRfGKb
wa5D3wNfoUEW5YmaTFAPP50sVwSeP+0oDetEYQiesuaxTfoM6ttEZd3uh7Buy1+vPN+Qoy8pqsFL
0ylkOdTA6Qu9K5leKtXwmlngT/gMDeniUxAqB25YbqYwQ6d1UwmtjBIctTWI0QS5zfS5QNK7wC+h
qZAACgoBYUPQONJ2zSziHtGfZqvvarSwGOnAQ2v79CMZHM2PsaE+uB7SIN4UJksxriCZ33oUR+OO
JKlf/VfwEj76qpYMTfXJLBo0zLjdSevaSct7knxMZnwVE5WxJba2j3r5eilQgf/Olr+I2yVALOEW
U5CSBNgfzoYu5tiu83B0af1FOgnXgi2O5XbO4I5sqR7Eo2ooYwuHl21rPIF34kJM/QS+AhgNziaY
gqUTUxIhIGdzQlvPwRimRAkyR+MMt+bPjuDEJPKGDZh9bBvvwm7y8KMbVsjLE0Q9SIqn8Pu8zQHF
tWIWrYnaspxch+7aby218KO/3x47ODBly+ao4qJ5O98RsqcDWxFEHmer0Z75kaQMa4t42L8xaQUS
ZN8Wp6iCCoWtzQPasgyzSOK1eZgYwqI+Qu5Xw5TFkQdAFsL7jDySELqjFCSEOC2Xq01mXCooTm3A
21aivRF80d+p7J6uv9jNKLZ6m+5pGGbgkleeBOR+YuG/wvllgQ6Sc/lR42iDi9LElTlWIp6bZa8g
MDQIww+Wa8eJaeC1B+0porx5Ls5OZLn0kSdKEhCINmMXDL1NIJUthOc4VZEASNpuzDalgGLFygLi
hQfDgc6Hl+50LdzspywYa3OaRHhMtj8kiJ7iil3ks2RLzxbZUwv3E897EZQefUstlMb5TaSb67K2
XBlY+X5+XItdQ+bCZQGz/Pol1Xh/TX5c6Vc2tJnPcKuoLIlbtB1H+GVpOmpIfDDgCXTZZPL8cdTF
0RvearK3KdC59oxwrv4BGMIQhgXQ+Uvjrabv+qHlUQUIHUbg+iPMKmjgt2OCOudXd0iokEsW42zH
2WSoLY50xQkp4SQFZNF4CtFwnYrWILLWCIhMVx8TrEIr6660uGr0H24MviXzypdANQTiCZtFXBGk
qaoF/Bjg5mG2K1eycss94PSCtGpk6Y8IAIKKDRCeruP8pVFziqTq102YDblyJCTv7+O+4JvzJP4v
glzPHP9R5zMw4iG1QMyXRewUd1P0L7Gtr4kzZJkSxOGBLD4SDLkxn9Tyo01/CB2v5HFGQUTs8So+
66hFBj7fkkgim2fH88jgLOxnC304e7d+1q26FXdoXpWGL6YlI98RUtoYy9XbOoeii0HFvoYNR8j7
iKY4FYl/fizVs5SMYzPd7v5NKh7DtW7YQ8h3q0+Dw2dnS7NMGkJoZhN/DaIsHbju3VzWztqc0C0g
Onq7vM/DAhTWyMNsEGHXhc2bYiLaWrzLUH6F2HiOfRaKPXEzJ+qPEP8jR7fl4Hz3KjO6hrbxf/Re
rtuEN8wb5t6dwWfiSgO+FoFCiRo1OiwY7ZeV76KZmb3Gtd7bXVbHj2+sPzh88HoiX8PMxfE6rGWb
6tYyFny2HX5vZVJ2UrD9UoCtjCa/Rn0RjOxcwzfdP4EgPv1q0pjZ+AZorhV1YucfXAa7HGTfnJng
DNwf/OFfnHdWAVgMZD1pfkmKWJPxbyAA1M1ChQkruJDMchwF1Ym9Ie2qI59+VJVn0dHlN76XIQDx
x62x+9tyRYjS1TIoh8bEiBt+pTHZf9ueejKXU4KjCLpZGBcecxCvmm2YQaBAP6FWSiVUWTzuZMnL
WEAnkCtKDylGxlca2UHNhf8kBuHSpZ0eJLyTNTOHmvf0Jz0PjboPYHEIt4+PLIqTeVPJczSc86hS
tiTLlW/P+adb+ixOkmhy4UUIec83yVc9FI2GIBRnUtDPkgh3uEc9kDw1FMO35kfXv2NaOxdsi/kJ
4PwVoEFuMwddYm1TBMzh1zwEJSHEsM4pBb5+cyYfWHIrloYUU6hlERTAErnKyS9dTkOaTdNIpbQe
JrUXh258/lPpgPksv89JFvkvKAP+00T8zsNM5hrofTIDx1QjN+N06Qt+muCgB+WwOYOexk0TzrXU
Grkh6W5MWKTDOQPLydjT0kvKQztRF79rKbU5Amgkfc3xQfkm3PY7eVzN8RVz66jQe6VNeFTIerLo
plBK9iFFW1pRvm8aYsyxAA1vSfo8tZvC+PJjNay83VvXPosCS7NPbIzRu6Ofid/dWW0wlRuryoIC
6ZAFl6m6gxS6R6mG8Y+zgahcSorGZGa1ntPuNzLqDSwTyorowcjhzFNUJTmlhXIXXfwTEtSIeVx8
Bnnczu0dIQOkEqEExk9kJc6ej/H/bpGK+uAqCb1EIuagcPmUw7whm3CRm05S2z+CrCfIU2fTo7s/
3shYCfJNiRiwiexudfiiwdYPR61abFp5o2KSGQo/tXTknNMP7P312gE7BFEdBtIiao+bRmq0unzF
PiqxI4YtT9RzIoxrhS9tF70HyIbfbNlukBxvMNwfw8Anx5Bp69MMEzjIiUrWEECvL3he6vF55cij
TFBrv2sxvxsgfxRBtqHgs5Z9B3NfsA/n+QSrBdZlyvDjd46bj4zC8/J/SkqJaP7gFriWnyf1EuBW
VzMSsnpZkpFCWbTyUTERvskrP9ejqGZ4SnM3fKPJae9KK7Y/D7gBP27a2EYSB+ujTibHRI0Swis3
lmqTOnswHop6xLEyDNsvNokaZIASSy3wPjnIQMmwX8NNwFp7uvPLFUqJlZJit7Kcuub5f+kW5GFh
ju8WTswE8iqlZrnzFHxitcYgSy8VkhObOUyOMn68IaUuYSl1vo8lMIOgoy0mgRWPNIE6o3IS5Yuu
X4As3ZLVR0Q1MT5hCDSfZMUOupOI+jXdZqOVD2DmQivmx+flMGrTBkSTY5u4RaVtP9VILlqCp53E
OpxtMklqq0G3F3T5OmuYPQvlnBERuioSaThGGYnjVLQcVBACvFmehHqV5Q3RaQGnF8SaknYXUUS7
BDxdJfw7wg2xMKXhVBK0MGDedl2OxkhTDiDIg9Wa0qzMHYsol7a/fN6jE+0mtK6mK44jp+3FrWFM
rmjPbpEp+n1z6gm9JSbHF0WYA7uAEyCYI0+tWDdW1nJyk0RiYbQypqMNYU+d7vVijYjnqjj2bWVp
+fqQPoS2ISAakAYzwOzpm3A82IlhLuvYgUhD1Cm0xsy1CPJpPkQ1PTZuGOlJLZHWngKc0xGFrB7j
+kuFeI2U7LmRqWdX11adwiiGVw41seYnVxArtrfNL3C84+F3LXWEp6ww/fXU7IMbe4Rva0VUIxO3
OkyPcjTbuYcz7uW0UzRmBkwSxyo/KQPn0V/CCSsC1NRKBWmk8i1EBX3o6GVLg5scYYcHyTcd+5gk
ap8H3GBkru6GMEyPXY9PrN54iWTQ8Xq1twh7Id3bufzB+qSnztA78IkubXpeOb9qCAqzwu+BQtZ8
kldq1evwDZ0oGCgKYV4L0Zhk8Eel5b8SEkn5q/8Kjtc4NYRJCN5X5FL5/cQ/sjI5gAsLYRFWhBhC
FiVzSj050mLmuPhilJG9JL7qUf89cfPK+2Dv02rTsiJ8EK0tlA4vMggUkjVKwkDoANmkl0Wpk9aE
XfYOwP2sgid0u2E4X19/wqb5FA8CeZkR73E9kUboCxTB4+BQRKLKNI8pd5ctH5nBSxM+Tjt5m3Mg
QMedllFuh9eWVEi9aGrUa1zpY0A1auBxI6LWfXd9uO6uv3pT4I9G718eyuaaCk9l4J+4ju9brr2B
6ayHNo71wkE5F2ZzF0ie3zH54OzFgZBmLks2B2VWcjtLUOZGbom15VEwTOOZI+fjpF+ex+V+AsCL
jCM0liqrdw8QeSmLkAcDh3W+3rJfcTw88LCuTp8Ol6FMN/VogR0RJAijjH8ZxjUoQSRisEbrUWjY
s7DxjoOy3sMhhJbwrEIcNfe/+xVudnZj5LfN360yBXAn7U6oTSuZMeNRCMRcHuJiT+WrF6/nAe7J
dzz2Zd2iVgQT6alqbCMeyHFQZZVw4EC9PrATIDJCcjsyhTQLJUbtv3HCjpIXw2XR2/EtiLdRHDTL
8OfKxZU1imPf7yFTmSqTYy+/qHNVI0AyehPFg+rS2Y6oMNkKob/KNVPKxCHXkUZx6hF+ZE0Ii/dD
8ojM3+/jHFch2rp8OFXERyJHKa4m8av+3HnTYoCKrHSWqg0jhbRGRRX8nWKUY0Uqdd238GiuCEoK
z/SGeq8xxyNIIJW1wSkSXeSBgylpt3c9PjLChT9XH0lNST9UlQeRrjrpWNHzDeOZL9ymlUTYezDj
hCR3cikh63+UfnyJ1RFspbZ+aMWjJKNp9+gxPqK9b5IUs2DW8QooqCncl6KzBhF7oOEVKaCwJVG0
NQxgFQ11Y8qmE0sBPGn09XoS0fXYmeZupO8t/XyIVTqsMJIEGUILbP7iCpBIVKKsp6ZjVgSvJu6P
WRFIXQVTJWwhKH0/kMJR9mrH+4tjfztWHfE3bi8VTw8ysRlnG1LQBsVnTnQRmM5sioeP2Ey6qqOI
nqLq+Ea0wix/lRu4d+oLbI+zDhxh2IJ85fGabe5yLxCQwYCe59nVEjGlI+pPxycvthcRr9i07niu
nkW62NTdZQXNZMlLBFEUh+xwsbhOKMTSHq2cBF1/IgHNMlwAmvn2+Ub4fih21CRyuWNmVl+IwSZu
G+p7xfSbftGukYcxqsbBRlrzaTeHS103Wi6CKTTjIbce6niZ6JzDUVBXZod5Rb9E6Vq1ZB7vItTH
71GXH+OXhZCi6wSKlTH74Rf0Fip3b+OoEjnxOp/Oqyk2TBXwVnPA5Jm43VG5gmP6zK56zk2cGyyG
kToCKDvjyqWw6i6EBdFgL/xFiKkXPWJtUk6tD1FbLph7LPBcjghRB/0pLxjAv66TKlayMbah6vwy
Muehysy8yJaTcs6Wn1bSdH9jPusp/LsIZiTEyxYkIW66ksY10OFvNBiv+MoARwoJck3foUBCIJf1
BpUqamPiaESG8YpJ0Ty7hCXvYckcFeTYXlEKJLOhFf49xPbp9WgKEvnyKGCCiUPAlbbW/LJURdtB
uwbo4J0mp50/yKC0JQydSJCiJ5pliRViJnBhpR1J/fH1h3LiS1wjczdf4/1p01s+U2YzYqt2q6OI
V7g6xUtVtdayAJsEMySS8LweGWdWRZptxPeM6pqcq5zkd/0FCY1RMfDpGyUXbtsHWPXNGRr1mw3W
nYI7eFKsfalbXL46V2ZL+7t8BGWSYDEUlUzsh3gdCZ2bRXrYYwO8oDi3kWptJ3CLyraF3mDThhxQ
T7SvyJNslQF8dL/FhNGxj64hwqCkKu6Mvh7MFy1C0+MJvME7DP4+xwKBRJjr0ekkMORrKV9CMB4w
EdZ+6JekM7vEqiGdSejZvXbZdQkG4tj44SEP0/U0tSbkBAEIKsIs8g4nRR1CvY1y9xBWeJCJ+alP
esyn7dOCME72cSff+EguFi3BGOoacvRSSUpO7pWlqwxs9REj9jBExy6eK5HV6HjHRSsa+wSHiQf8
brj3YffoWl+BT8FrchpK89U9FZsQsR/dRwXaJDVi5k/pmaF26YQxNzYq+W6FjD2RHx5hPgFoY1ul
GjhMgSychmvhRV076f6pi+F6mHIo3P2zWDJyTnjlgkK26HbY7ZCKEFpPF7OfmkuVdnw+G2Mp0X5O
fscVdqGvs60N0BmOKLTf1I1vhV2lHt31QalcXUnYlQtJno1RU42zIhYf5bT4qj252z2ZznpRBaV6
/4CyMfgLPNWBsv1KIyCSG6cJgrO2GpUfDVpgS/sy3SqWjEz3ZHI+wcRx7nui94aaZ6tuBMNb1Mrg
vgWW5rbGncXsf5uNrvR6WtIVp877+WUCS61oNLpt3QXHSrxBLG/KDC4c5hitbwVisvJwabsO0qpP
1XbP503KdVDl6+FyQaWs8OXkwvt09d3x8PNNOziGudfdeLAMIVaC6vYJ94ps3ucGBl4nZ7SMYIFt
Dhv6k+6b95oQ0QlzX2nlvezuez+04oqnSE22OIvyuyTUFi7E2DMJ5uWaOa6y4kOQNqiwDF6YHY+R
9Kt6ocJ9XgnGkt+0E8eJsdLiRUwF1vxBJ9blIBg5a2MZPLKiQDnScOkGZpyz672mBCUXBk322GoY
2/VOeZIgr2wRUVGXn97sOjitn9bnsYaODsH/S6QzK059xw7mJhzYdpVod2myUOpTb7jARLQ7YPOb
1xgDr7hZ+WDjpz89gmzbsjLLhiUrsrja86eE6NrEHgXuTswGwFz5RuiP22Hnpf90HyzFYhgYO9ED
lffcVclv6d5s3gkmBAT0Rz1qNxNZnX3ylqLYcHpJHaBdXvTmXTNDaqFb6Y1sbIO1NrpuBEwYAk+X
ihkkSBVvqQ7M4kA5seDbMYMx9pwjbT7gnmiLR7CbtIOp1+1VXClh0VE8Pg7Fe9uJvGt9fhcW/AL9
d3NJByjLAASFvvhlm4MlZfMjRYh/kPYRT/pCtPWMmB3M75ag+8vjwwaDJI78YTaeS4yIDTEg/95w
R42To2+wyKoPoPVuJfoBtyemRNZrKI8Ty5QwnmBgnXun4LV94RxTR+RMD/BeSkf7SrrluDVd3wyW
oZ+Y7e7HPaKEdSxXbziTFQD/6lwhjFV6TtIaJuErha/MaiE4s6hC0hhA9iwQ2oRrgpn1ho89G0WH
6hdXEEIsR5m2NYA9mtcXxOSbuQmg+IfYtZGNw4W9BDXLJlDveE5DV7StL+9bXOpAQ/8iYBVq5yXA
gsHJuNZ5CxxuLIwWEzoVTS9N60CzyXwpnREQ5Vs0Pioc2WHacByE91UDsMpbFwp4a5uqbjLCuedT
8DVwAmIwbFreJTT9mNkz8QdAEFJw2aPUsnG8gPT5S5qaTUdHLSkJZ/KFPI1uzs2mnMvRo7qYVTpb
+lLB/wZ9nuCYNMBvIinQ+WMsiLcpHCkSJ1ifTCN30X/26i8uWN/SQr4dGfgV06IR1IobWSbiA+Hc
xFcDtX5pY+rOa4J/5f+uZCMmnPYn8lPrFPtkrUlGE5lAzQL+pB2NYRcC2R2m1J7vJQXARC4mpO11
YFMuW/Vc3VqrwXZVymMy6FxENAnImUb4MoPRHQYkNxt+HD9MkOF2a1sor0RTOT74ukyRl+e6Lr7g
JBd7D7/KWuXXqgGJNASdANj/thFZjqVdvSANzkd+DzZRAlO8JZDNW6cvi8L4vUXOXkAeGJE7b0+a
yy/+Q/I426gG4JWU5/JNnNuNAoiuoGbxJhv9N7Cjls5Umt6NcCu3IpF+J6cNfOZY4Po4kdLniwGi
BSAuZbgBNjO/2aXavVb8v/Sk1xsIjlM1ed8WEDkQSVJFSq7j3QlePQUM06v+bAdXdB7KJj3Vla/2
YqlDW9fyZeqMBO0KNQrylEiOaOU7qBCrISLbF3Jgbznyw1t9/5Yg2w3afX3Guajpxfi56Ir2BTnl
M5KXTHUxVGfAInWMWZi7tcBC7/IZE4FauhMDSqMFHB6NSsF5jkp7lxNp66rWefuo/az2ep+7fwD2
EChip4E8paoZwV9rtq6hz/5a6Fb0y5V+7Mpg9azJXPVPtRGSjKHn/WHm0AvA86pwnL4/nDODWQ9D
vU97/SBN2gfk2RFdGkpy9KJvEOAOvyqfRqP0hzNtwuoi9bRG1pPyEj5bxacvX8ccyxgEOy3Imp0u
vXjDJDfrchl/nsuADT9b/UyzEHDuM5hc4WippuYaXO8rgxf414ERGVKwMS7aVi4NrhcRdFVxzvVb
O38GPfXTYcvHmQ8aWzWQCIYsr4WGoicCOWRoeeaB2JuaPvugET0sK2mmj8VjaN5ady4Ad8pg7DiP
AdeBglzVIK55p/kvI1Q4k81ovKmeGYJJ75jfAwGDbbEEZ3XI4P6kGk4Q6mJnWjYRK6QWVPKi5zg6
uz4PNCuuiUspzyY5UpoPQG67Qn1E6AP//eniavcWfhg4u94jZ0Trs9+ayWv30WTkukFN87ajIf6O
tDGVMVPolvYMYpp6W6H5kS1oQkj4wmuf5j3boDofr+Pg8aVm9MU5uZdOk3DDlWJ634JabJaEmMA1
ZuD+m64AueJ0qz4JwEb4Jgac1zjdf4A5edzpWWhmuIXctKoXHWJFNK0uCmoG2HMzbupGGU9Tje/O
qF6WZ4QZ0shCT512DSdf1qZbdzKTiZO4Mawtpv+HbU6DsJ9u/+/zcb4QIea4pnKpLPhtmRLpXAX3
DGvO7koAi5RQXkX4G1hsCZzAQGqmS5aPDIvWpXvLqzdwKWK4Jvqv6q6pVRbBtNxiUi4ZJdLKk90l
yM2g0DBQDRIIQUN8lK1TlA/O0c9JOrOUPCcP6eEh1PO/S8rIyLpUz8A44ZdMStpcZrEDGluUbfAM
sl6Xdk3jOiPqzcsPI7j3OpS83w8hmzlgGzSCNNZFawDEUMgIKIAaooz07ZTMCXS5MiZKgPvqgOj4
79MxZRInPA+fAeNHeXLfuTxLyWEMUsoM9Q2//eDZNnHAxpGSUaQaBMuSMsRJTk/Wr8l5vKeMXwxZ
1QgSx8X4Vtstoa1qgF23/XWd85wybTWO2GDxLHl0O5l26LJaZwL4nV+d0RX75+aOgkU73rfZCUhz
WD1SHSbJJdg5P9ezllJWQRFuiPOHauf8K/SUgfDYo6Y0ts/nDET9cpdoJccaw5KWrMmd+VhgTQsL
KsdUauRbjAqmG0qmVFGzdpiH8yItfxTsiyn3LL2Otbw/YfG8z3Urgou7tCrz2TFAnT6t56xKMi41
vxwG7S5EwkCpKW7qVOZjSyYUT/NENV454vXSQw7XZgkEybQ/jTAo8agHlGcJ2zsy5B8/KqPHbDc1
0chvPinSXGcYGOMVCBPdwgaUzbYRaEwN9eUKLadDNQVyobyAxLyQuUisiRnklPkH4XiOr4SA69LX
Zy715xjE9ou6uSDaRz+T3/fTkjLgqMUxxkApVFknnylVRLO6/i+qmLnyIYrwq93jR3pCPPf7QmcI
n/feV9w3tKgkQPguZtIBCD913K1imbXuWOBSGSYtN1M6MCoC7+wHmfQRCmhkrjOeD84b//um2xAq
y5sKcZQ9P2D+1V//SueYxZ3wwCqkuJSyvB1j0Xxjq5H37sb66IJ9aGOjfrv/Pwbw6uU449kT3vjU
z1gvJxCFT5IMOrZ3fZMQ4NmFzUOq8ycLgWv6aueezs61GZO+FgtyrNTTOTnD2afO3jbbPMZCYxj4
6LxYNQpx3hqRGdFElp03P+lqHZYlJMZfCWIxgiRwbxbXU3MeW66H5ShYWOxdk0ZQ7uNd9WnAK4vk
dm42plDMrzW6wC49TpBcEmmxHU7kAUP0HQNevMwIHbmE/Wj2H+U4+z8hhNU7mByJRzLGnBYcAZeM
7TxfrJ6r6+nlW8TscHPJ/e2a2huCkPbIwxv1oskZH5vIexaSb8aztk/rXWsQLWsSp1X44dSp1vRv
GGRLCO7NrgAq7hzm1Fth3HO/Lq+7qQQtPumBkaaDVp/004FdDFHQbDZt1Fsyw8szWMjSKSoaZiKB
5hiSZ37GDpXKm6t9I0InM5UGg/6XyeEZELCFZcJZ00IKfODWBBw2N77LEsB0bvjX3Xcmg7F0SVuc
WjE2pTIo3IcCLGd1RamQkYW+1+svVMBK6H2B/FY0r55i1e80z/4AS7tu8eZiYKQPNVI6atQmc/pJ
mV67ZxAbbB3Yh5fnA1YdDccRlZHtbQpC9Nv2yPjX4EuAXeKI+tSWB4WoPFwO/xOKRxxS/ri2070G
DEj6mn8kVCDWTlgZitS0rfCAXKBqIb9qQvaV2DhJf9ucQPEYKEOHmcQk8ZvYSsft+cB1DnKsX90b
uZ+LIO9CqY178EMvMLCVn0H2qSuMOXEdf42rUMDH4uZnPR6LTaFFv1ACQZv5c9cDQd+jfPmek+N5
GE92C5YmgUNrCwhcOCgrSXbPn70U6zXToe1ExssMzKK5KRiHyHf8NnKVV/+zIr72Snv1qqn+BGLu
QoSc/HiS35dMLinnG+OfbGUR3EioKhuPdGbgnq9+R3aUpYF7pba6B0AUP9ncbEKEIaGvqB9bk45v
gKIoI/xzU1gFdMwaC99+mZEQ2ssa032ogduFlY7yLQBPkaRlOCsNKEkddPBgXJ7aEJX6NhrvHAlr
/rjQL9gJeIkuCSVgLOQ5nCra4LEqQyAhBaluSO8F5aZzQXHRTNwH828EgV+zue/+rX3Jp2O09Jig
pPGv3s1ynG1n5tZXRsh9LIxBQH+JsubQwapv5XvXvJSDtwU+rVUMvWJdRZZMITTOWN0vWanh/MLt
4WuKyMQsO/07NeUitkzRtjDjPe8nJOaGq1zwuzDP+Btw7uT92qoH3ACZbHjme4oclFb/dyqHQt27
s7MaiU0K3/szUVKvX2NB8xVm+6df8IWwfRQGjZToAopPmcFsuj1sqXvjc4/BzooQAZXhxNYMDMn3
AII6jqNodaXPWKK1BlxCjNmcZ48vGtWuHtBBGMChmwOG2jlB5UT0GFd6ULCWqiJmv9Vc3Z9n21o5
4k74bxAmgQY8TncwDWrCBIpSyg9fXcsjls+yrBql2+UhLH0eTmCFIe+W/2UnipDToHA2M03AqpsX
Tw/X1I5fxEjPBtkcJmC0rxYBt6Ss9n12lcX1OpxVgL/3ssuWhTMioWq5DHxBqGLh19GbDMekX7RI
IQujqWj+0T1ROsDokm169OobUr1X90RjZ7oUxXbYPqr6yyrU2DDyyAfZIBFSmfBx3XQ2mhlkdPa/
jhm8uQiYD62MqZgoibYd/MyKPkTSsnotpeN+iFmYyMYDiSkKjaehoYcqBp+G5ubBDqbXvBv8aiE2
Uh61DJoi/uCaZdPcBso9gu4nhYNyfhZf/uJC/BFkt0fUiQ+6fGd+PIpC9eexRL+HtsfWCDNTHDwm
ab4I62lnkX1Xyxhz8+kD9DqIlt6tXvmGa5vEPlzB1BL85joblj6Ube1bYu1dXpOEdskaM7yEg6gg
Gln99HK5IBXt1KRkZAU9aFhAzehhHY6GDo3Z+9Upp7aASZS4Ix0erq6IOzBNcI1mgctOqorOaZ0M
Zek0qf26pUdIdzgDC5wmKMC78moQkXzU/jfcMxY765xSiePfZXotc4pYLUY8Q1eracMv2z+z7RHK
lWTgOrQwFr75LgN6e+OQhHBXCxnGNMf46Es78JtxyWWB0819c8DgRqKuOo/TQEvt1kZ4TlQI7uux
/LToEzNMHBD6TbL/oIroit4xrGpZwNqGFrT2z/cgdyWJNxMP6BTgpHutn2wB1EE9vmOMTt20dEZA
sVX9FbvvqmyUa2J0wEMuRiI6wSPPKzC0aOnjuM0hIMdJh6bwtCTYFcI9ns7jkxR7yHVZeAnAclAj
IfZI4hrrWNvWsya7sfpmd/RPGwk/PAnq8LFW3t40AayM8DeXi0aDpW/RCUailf+UAglDZ43ORBub
JNqMn4d2aOkTTs78qy1XoL1aiah98+Twr3xu7VnJFEph9Qs3s08cQFc7XqCDB5YyTIJVJufr3iMA
qf/UEzK1cTuOPm8JA4MVHxltN2P5N95njKNd6By8eo5ia4dXNSTiMGt4wFUvH1KDrsgfVeCsaNLd
urLyrFqmWBPOA1auOluvw5d0fqS8LaN2QhXEC6FvzDjLyNjY2rM7bLV+nKlpMiOlQ7FwMerJ5jBP
ZoovodGNq2sq8o+fjzzw3QLgLzKCXdt8siaXxx6Hib7be0krbvMxXv/msU8wzkqs0LqdEvxNwlHA
ecOfQaKb01A0MnW9g0pZwnGPjnHmVCzUdarYr6JecHJW+OhHiOMw7pe9brXGwAL2dQmm4c7h/TSO
ns6kw7AnOOY907yC4jiglc5JxTy/Rl7+imsT/kKz1aEESGDhy7MymgCqKegeDS5LHlUYbxTQLjhr
kEA7u9O6xSezEsKu0CzguUPznbmMMPa1/bLy0QRG9qCotFxVSh6xuGg5WJulvjJ8saPjmptcgI7V
hkshH20E0EAi4Ea4tt2FDNLz8sfIsrLfYXOM9XEexUwTTuoEZM1A6zFTfJmbg4QRiAAfpXH7Kn7g
FNqGar8rdu46bqgHTiL0UHA27NJyWxsZjVXn5f44AUtJdKB5erzKBSTOnegukxV2ApbFVZ/e6L+q
BPWoefvhAnnrbUKR672m0JunTKxaMOwNXd7pYcTBT4xlrXIa8sPpHQPas7gmDuXWJZyxhsn4TQYq
YUAyJ6XIjUekPYiE19lhtVsIUjOTRdYjQ/B5QGT4dTMuHFVIxCldjrHrd1CMKGJjcpi5tn77kWG0
f4Lc6k2WkLmDZE/KCFb0mFG+wErl+29fI0iYdnYwNwuysctUmMmJcxEQIZFa7imMB6xDwIGjLj4T
28ty/a5n6yDHR6QZHsR5wDfn6W01eWwfwYhlZ+nbQOz07jEAbdmGXw7CO0WxC2J8dRbh9amwZ2ud
cD0isrThKiSiSgkvtzJv7G7PCXNgkS0B+UAg3dZqDn826SufKHHkG/Zpcj2bSSlJclcGMuC86O18
WPE6M3LEftqOo4ZICo5RXfY378yLFZImfkN4bKOrXvC/ZJYrKfLoe27BnF/wgqThSkWNkAx0OTfq
CUEKQkOB66ZdTkqLJVG5SufI4NAqxL6PlKBl7oaCBLz2ykDJ2D9UvGvtcFAyd+u96ff5A9h/vSuw
DAAIaSU4JmV1uFiSKXk3loAh4dEr4uJY+FPCW9m1GcKerP4kdUsHhC4JZofFf6pLhJrKz4u/NjcG
TiOtDUwuPNLo6ueLCTfIYdGddNUCdYYswOLGpwb3+0Awtv5kjNayNUXhEUZSznasBx+1pQABLAtE
Vo2WAsrbDfOlsB2NfdY3+O/vUvyP4oDhdbdMEvOur/qin1aieyn9r0l3FVahALXAeEZoRfOrKXko
4Z8bgWeWfBFJBpCWx56pO8weNK/nH/sVQfnCW/JrGt2ClE9Nsd/nbHDRII/WllWoHDmO8wCUiH6i
qScEYd2q2PQQX93/dL1R0PG7k5OIK1rQNYXL6i77r3SAvXa9lJ0ErhYOP1P/y3UAxyUssn8beYVe
tv0Gr4I5g3X/YGRxluXUDqo6B085QEjryp1wRURcOBunKWKrhv3lSilSpYuMB/i74Jb472DyOEiP
0R8YXA6N5j2arO6nRyYVsGVo8TeiT3+rhm54cCYfsEaTpdzRNE230xKp/FN6wwL7oAaEaEB58SWH
lVQJ9qrOcIPlBo7CpLt0qZ9r9wFd9ZJsm6pWkhlPGTy20RdCTqA8JZogsBxMtK1MziiTUEJHxi6G
jdC+XtkZrR95kGWXqjrIqqWwkoS5rCozmWufLcvJ+qn1o/W1j9JRteIG8JyCz5QIyWVt4T/YPpIh
ovgGUWhE+vV3Kgz0f8ShAw8PsrSX8mYRxNyZxCa6K1lXPDYsrkIetLd+Pu9rhvB4+8nFvjenWNaB
GlzE1Xx5ArdSHE+RilYrrvvBQ+25uoWm/MBZVHEUH2ye0XA9vZtXWc/60naRoBPV+xAaFoVK60FV
FMc0ISyDmyfiHSMq0Gxu4kNJKWquj51QPiFNzdl/uRA74DyWpHejUJtiZfFtZAM4BqG48pe78q7D
/BkzuW9B6QScb2gHvUv/9tug6UjLpdYIdHAmS50h27WN0B89j4kz/Lr4uW38V2j80K0k6shaomb3
2Fbcog/MSXyFPetems/BCBXuSRJC1/p6ZorT3dM+ikx6bPrGIs/fFXdHjajNBDVoOMc5Frmbwt1+
bu/bTvCvqmVThyxmxURDvWePMzmoQ59qs4Sh4sJFjWT+XKTKvEgasxWES6iqPTSO6ljdy+opYYB7
X/QHOXv6nY/dxhM+zhkrPtK7V31eiglkLJ2gKSuwIt8PMa2SfeS2tmUEo9NAqKctBw5TGuGF82v3
46+tDyX9Pjir/gsHOqPBs686OyzXryvnrXs5SayDAnM0A1c1AKcr9l1yDB1E9HdtUZfXeQkp4cEj
UWoFc9PoeC/TtPhQtvUPGaPQTDECMcDFB26NGyJy1Gy7cDM0kwhqfSQF7L019OihH3WtNb/SI30z
d3GhFw3mVwmU2GEGLq0qeFKRdJrg413hMPS1YFQ37IIjwhg5hchkwgUW08LVZJxgcI4b3UqCSlJg
Cul0nAOdsTU6kD1W27zrTKIC/hy6hT/Pf6VAGFGlhGpiVfOo+4IyFeGpl19qVsvN9SA941qxe2fv
QUM+FOIA5Uzc6HqNz1YmvTmfu7+0uN8lC+G7NJbVKJE08dHveHCBYtlgS18E6S8T9CCBQuCqOMRL
OvypOquLw7diX/DMDOpFS5ufcYNJtNvOAxwno4ZdKApyed0Hy+hyp6odzgp5WARJb2CMs1ifXhRp
YFeNBBl5MPlzBy1qyiN4ymULdo4qfkI9klqYVChvCJIqmI1uTXDZwN5NSxJxAHzZpAT/hkV/F31H
dxyKc/h4K0PcitGb1oo95WM+ZaG7fSGOpHjx8GOYT3qjwzlp6s9Le2fxwkcAb3KW3BvTPBLSj/6O
PnbSramLGcSO7QggS41Y4ZVBRicm+ykHQw6iDIafc4PAlYJwggApppgk2YwAi0aYGAjjV2rRdy3l
y0sCOTWzMVgxA7zxiOZbh3BPHbOLOjdnnD7Wxbps0ShN/JhkyjGZy4SgbqO3q1R40Xcw6mVuXwm5
um6n88QQ4Hg9cO5ALWslDN+nYZ1est6oNmAVtdx6MfCEfdhklkHD+nbO5JD590Wus42ser8MC4De
TbVnGHQTT9HXf4zoHLyEDBfGZ0Wr9FmEcg5ZCKgvNWelDXEhBoBDWy/FrGpas13zdYRas5DqwZel
2bQ1A+xIOsd5cM1abcX+EXHTavSVw8k729GW26u/cMLi/dDx7BH1oriY9FpctH4p+/0ykdJKC0df
JXsox/OqYsN+LKCV56EUhnndnjyvdpMT9+ovwRJWSEZ4u50x8paErUjRXLAG4NmaEkLFmdwvjYFS
pdVw6jD9GxLwdTcYcEVtdvVyggHVa4TWqe6/+hg3lLeho2p2uND4VPvXtRFBYmUhbRpt0X1f9gga
OE3URYUHeXCrc31ABa/kw/bUb0Qpj7nELFDAC3d3cQ4y2cLD8ePIUyLnaAN/NKW2GFPFBClchbPS
dLpbYr+EFze5iMiAQMQ3jZWyAXAdLk7OzpQAzKaukY2j4Sl4TU+qiiQ+9mVfMmPROJki0sYQXegy
6Eoc7dchJK8dy3j9Ij26xWNYgCWcyZyYVh1e4wGUBmP0XftfAN2BuRBydBghHpqUrKXzgWyFE+yz
d5p31tcYCVv0v13785mvLZ0T1C7Zztm5bYTmyjUl2CMKGlL/156pGrZfdeqmgepzSMKSZMHHkmuJ
xnTEws3Lmai/fCAUOuU9VxawTzx1GCDho8D8t0gStwGlKm5llm6Hk9M2pL+AXW+p8Sm+CRBDI7EZ
pHIwUBBwZsL9c4q8ED3c0YLSJoQcMlIbD6pl2JRDiCTExyVamJ5fMCUNdpenwu9JWBPFdJ0IUQ1P
8kowuDisJAnrWraYGTDaf7U5Yp7Jr1z+b9QHklQ2MVFIyPRfFBw/GXlFCC54PiUqaHpCLfRqtCcC
MHYtwgWqrq8SaSj0frQnxztU3XlHeQTCLQ0KS2rqlCPRE2WUw+vMdX+Q7dYOdf25vBZ8RWzsmcWi
VqLTTY9/P7GgAc3fN7FODqeofKmeY1gS30KYwi+u+U4IPzMUPplSnIeuBLc/8iz3fdyuCZQAAI9X
ZX+cQ2Kzbnt1PG2p121CldiIQx2RUbAI6gl44M/Q+ANCjQR8mtii4R9NOnImX41fuo1HJbwcyJZ9
gcF68Oq+LIOPDj+mO6f3Yd0BL8XobJsT902iRxuQf8zIybkYuvEx//CgrZSgvNhsa67P6wU5gsDi
BjiT9maG5xUE2JCkSDDYf8RYeeuF/p3l5Uv5CYULqCRxZj81ORuEdi5gmmcPjfzEc+frLt9s5+Gi
zAof2+dWb939f0RU5wEpsWfOtMnmKzB2i2qn1vgV+MhSm7rRK5WcqunsAMfF0a800cMpmt04gWIE
3yKGPtd6ebfNq5uIyvfKgnmBE7VjlzhTwMLcvEP9zQ2eLmVu2PgXOsY6QBDHNMsr9Ew6GyofOzDZ
2xGgr7qKM4OjH3pOM2QJ4EagGv37u4UOF8Qal79FXItz+lP0gCaTOotP649ogD6SLq64Ay1DWjfA
8F40uXJ1NDgNrJHQA7APvpW74V1z7tlOIliPZchOOgwcZzUhYZL+hoh84giT6i/LapMsGXkX8Pbu
TB6JL7iPFwyxPcjKhiTKv2msRRx17Chv8qwpnWFIARVTVzv5YA5iEB98JCfTvLC3p/OM5SXbctkW
vtrR+vkzDDS6WG4Z/ZQ0PmOadTSp+dax1V8mrwfQPzaECnOLxN24/0uczf+eIWLUQ0ML2PRpJzvI
38eKt5uXxTgMsumjWWhArZjifkE/nnru/AXufd8zttu/D2xYu+x5eQG1EcXEp0LhF6LpFJaUzZ+6
ZThyNfRObgygoY1L9MTrEvnQqwAnKvB0U+CK9Q63+n2gqGvF3Sjh1Ee+rJtLK93QjRAAdC/eLYSD
nlOn/Oo53WZqF0tNoMY8erSo7cYrQ98s3x67cbpTOZ/jysapHWhGo3jPcBtx7X7qKM6Is9cD1UVE
Fet2cRYUvmhgUGfFKZdl/s2XqP1bDl5EgAWydm5WpaBrn8BnzexPoXqlsZ491w3im9tlDevK12WR
vLv1QOdH/hSsk6fNOXn55I2+s02QOVVPg27IGG8xQTmAzul9V+QjHy81sL9SsOA/YLZYOxLw6hLd
fkyfTJoSiEwbnnOfWShHlif7Lx6RVPz8fWnXM6NLwSGwCsnBIS9Trfo3mfnTd82ejvlzVPpfBsjw
kKEdPUIoFwnVTWr0oB/hG+c3Jz8oh34miWS60xIzZtFBNbkB8tp4EwL0cGMniX3IULqJ32gw8ylI
0DB+ypO5KIrLhjTG61+lWlFq25WA8jd5WA8p9we1dLG/6qonUHzexq4USMnTK58tyhlgLCNYq6Y4
v2PfPBh2G2l5f84oyoogzSijKT6Ay+Dz/8vObxeGvblwzqevyVSNHzhirx4nnvQNw/9vA01q1/kO
/qRfZKL+5ym3Gv8Cp74Zi+5zD27B1j2tibicV9uZjlNcWdgtObk74fQy1M2xFPhY8FgiZHYrkm8Z
APaZpMWnq+X3SoqHUdRvu7FmdNAHxidrb+k5ju/wAqCYHAam7btlM5g8tDo9fcah0vTbZHBonNbE
QCZzeYKRiG4uWvrDfZiHjTbF9sLcYhb/40azEJWtj1BvmNbtpAzIJOQGMKZjGhZCE5WGFdWs9Fi0
DoOsprRm0/SSLjE1tL6vTmUVwouPrMzdcEVddeq4kVH32crIlUuH66IgPJbvnED7pHjlZxgy9U2m
VDzWgwAMAUYlCGbSe9gKByNiRikfHsEBWXnz5vLme+2vn+KetfQRFTNoJ56vMdlpBdWMzS7q7+7N
K1mT67fxcTA36I/Cieg5r3etNBrwX62R5GW/Ny4rkpDNDW/BILmr+Ft8jpiEsDaAHWiVelIROG5k
XSgrpGSZSM/40o96HisBoMK/Ri3+NG9Kj/1d5CoN07xG9hKfv1WTXCyhDsOIRdVSN2ZFRepKqmhD
Q3CWqeGYK3Ki0uNehTsc21MzU4GsD2TtJ+i9P2f4J2YebWbZJ7U5gLTqWLRsuxQjZqILk1yFM/Qg
vpLpe3QqXv2lG8BZBI9JuBbbx/ve4lYo9Gs42Vjv5s3hYo1j2FgNcUeL854MlVcAN8FV0NpMCW5n
wPcbjJB7svuKR6BWnY+F4ZmOe95yvauy6meYa7PrQ/+hOTsU1+ZplsJXxcP0NsMifm1UukwSzvRB
SfsXvp1zzCQCsbaaJhQrTa8kEfnVeDCWJUl+WkWE60KxOqpjmn9By4+07vBeJQ/kRDEWsYPlcEBw
xMcyr+7pl8CfM0Q7BRTtAEazcVzFJxZRbXyIORAlMK+qsSRv6CwDNy1kU43mUO5KGauWvI5srJhK
9tPXkICOvZuD8iYup1MEgy7+0cYtYRbp5aju64akMXbuNFqEaJqkv3eYN9ZwHHo68E8rIgUGAEf0
NQ1wW/Nwl+j0nkAAaZtHIZGsNE4Du/CKl0nNsn6Y1pMWaVGz6rW45lgp88Bj/+FdVryaPYltIg1B
ajAoD1M7Waase6OQ36qjsxPQvJyvJ7XsAvUcstq0LAK0ILGAS8es2i5dJG3OZrmbsB7AajEcJRQz
8R/A4Ly3va4Oedwx22R88uOdKoTa9v4JPNHxRBqB6Zo9M55U+SLTtfZGLr+W9Yite1erPXngenid
yGxXLDT8TloM/RHW5dFeWSgVOFZPV6l/Mp1Qvo3qaM8w+oOE1tw1wknXUsllmxWKt1YPiluX22Ry
SJ2zsibOqPKJX7bhGX9cNzr/Cw3i4NIvaN5PlLaPn0wCVEYds9VCtmAm/r+o497h3WuwN9Na/a/0
pfLtSQUe79cs928tUjyfFpW3W3VORLjThHULsbNuBvvdypS2Z+ZoUfII/1aKPdSxnAaxVHQRPRZb
d22/l9Ta+T1lzYzHuAvWf9mSrmzz5T4GkUTa7kr2fiA1tbAGDY4Mvb7NzuuBAN4EP9jzSKFPc7pN
sy7WcuM+PCt/w7xYhkT5q+zhKu8I7kePY5rh4laX4Xlh7kyirkbtXyLeWgklnYK8V4dU+gquXgpq
+r8oif4fpv5bw+VkrE1AWPMHF1pBx3Xgqo4ZbRf/pdzPvkXT+Lh1/27xBpnb6DqDXoAWdGo2fj/A
ypcm+U3C3YJS/YCvxgxocbtp7lfYHjamkASeGKL0+gJFLYQLPuXWL3qrNg8OwxXapvkq+xd6+6NN
AMO5CF81XldkYNgECA8yzXACihp8Rqk4jhQiodyCibWQ4GZl7RLRIRM9J7g0pWFv41LlLBdStJii
oPo4CsYe1TdZQz92/NfKK1LHpiMdYPQral6ssX2nmFpY1uj87yAMLAeovty3F43TtXKauGjJ1sk0
jD2NZ+bOzVfrS1VQGrr3NmZb9vNmRyY1U125K9qciB69W47mwjXYp5wcwsdLNWTrN+IyBDhlTxbC
B7MkiKyPmARonhqm2goL5ai139dwtMyGdA+R5tmzEBF7YcCSlj4wxIxIWvWZPe2YI59iENHd4UyY
C87HW8FssyWxvpkqNNAmyM5Lw77Lfnp2U+qyh54rto5nXWmM5PGBY2nZQGRz5EM0WLCyqLfeCqgC
Bhx6cPG1T3KCAmgQBAOkkw3texz9Ejy8n1VsGcG7915b+HLuQvpvwRH3pFw5tcGoT+uWe8HrpnnU
NIkiQLSJE3gcWurPhVu0FYLeEdNAxy2VTgpxXOwb53bEQN+wH2WdViW2E3SH5m5EPkL829QzWZbC
wD6USxpwUgPW9YZLdYGeNiRD46deWsI1/bfZDlE1DXIwZLo5Viv3OxIk50ONZvSnaPI8P8WUFHUM
0m9cufI02z4MBVk42bvNJTEz513esEFJiIdtkj22liq9oxgp7YL/oxAxWErb+geRMqPF8F0G3jPR
lJJ8YXysZStyWy63nadGjG8GdCTNLATLmWHx19DusGhwoPjPag/jg1nBLbhIaVqrXYL4qLhfUM7F
w1gFJ14VapytZ4kbw6Llwtq/NALZX6Y9J8n22nu0gJ0ntGZg02LaxG31gTBBETrmF/8srwqwuEXr
54ukm/N4pV6dou33cJgTM4VO0xmG1LB+i5ROLeL+XKvx7EsQe6Z089C8WKxWLPF26ckZZETJNsA3
Wn4o51BN2q5XQ0X5nGuCJQQxV+efqeuM03AfayqXejCJkXrniRR2vcFgAfsoCFuMtdrOnqrCkBvA
7aKihuNIvtsgdTkjOh6oxC2pYqIZMGrhrCoHYgTK2UK3r4dTDJ9lu0x9EAJCdA20EZGGjmYczSZF
uqmEZ79GFpxnbvVMrH5TPd3L+FhiXsv2Ob+JgCEzhtpNRAdgmRJXbChJp43rg5qPA37091cXu2UP
vcVttTB7BxJ+35ipj8jKVEpPqFnyUR+wmxYdeT/o5p0/LtqR6tLvc5euFssxDxiOSxsFaIsrSPFg
28PsE5tU+fOFVTgHe45HYAEQ1csqK7B70+CK5F190BCLo7HJnFNCypQdZw7bpo+qqpJH6stt8aN1
VrQ75PCBP7q/3X2h4LqL7ffoOb3t5jTA6cFAwGE7bC3gARMAuzjkqdUYizAv5zBkWEd+vJhA1q4N
khEQD9VCKVSh3VCgVOc5YLc6nbfIcaD2AQawlw0bnFxzx02WgLpdH3uTON8cnwd05z5vlY91nAK6
K47LxYqczwHU1HpvB+xJ+aNjg4lvSkgIupT2dHaAjCtZ0jTCEJKxfCaHKLNhL18y0krMUr62icV5
IPaAA/hELxzxsBVrZXOHsrdV2CvArOZMjXpfoQ4VdDqRScSbyPvxNa9VERB3nQpMkEvPcPko/HbV
4gY0myq1YjYvXptKwT0wKKQTJfDE7xNvpf6u4oQwYvXydpjHGPC5HkW3KZGB8K8sqPyi5KhjL4ra
YAKGAHZ5IG/TlsDbd4OHBUp6Mx5vRjm+IE5/9tT75myX5Yhq1E4Po9wgy2SuZe77mXPRpb2fA6fq
MOQV/DG42qJcAMkfh+/VTA6lZiOTqGN86NB34ESXMqLQDVl1FaSislvcSiRtBis3zgpfX41c+/L1
teQ6aXtMPADLyMQkT4zZqzONKF6RyyWw+zhPOzJAp9girazw7cNKno9pIUAB+XDZK715pIERjbHy
r1Zv5CPNNNLBGTQCjkLh82OutNoCwPPNdIqB7Vwcp3uj/n9ZPQ85We77pdITw+JPxfiYhodtyVNc
83fLc+N3Dv9qRNjQqUgL0KGY205AkLSg0gjjCISb8E3W6PmucpBya+B8wStkKkoQL/6Racvy8FjF
IfNeoFEkfrmO/ibZkBG6F2bk61yWEZzWWUkistWLZTRYgOWdsx+YCJexGLsocFNCtNDKjZm6QkQZ
L6zGfGxfKpDGtKMfTvIE57loug7pZibdTwvu19Mi9ZlBTSwIC4jWX+ffYh+KwAMhaJM1KwJHblmQ
N+z6sVamBbR32Nm7ZSWMEtKt1KmJNSX6es0qLFuBgVus7L/kxo64jJHIz8b4uoGuYoZGgD9f2Pdr
/mdCIIrkWoNKBIsfAQAZiGmhMPJB4rCJY74a6HPJttFiFHhUssZJOX/e40O8RQHgHQsx8AchnTVN
IINa4fK3+GlXFkQTB8EUkW0g8Ch9iKOIxNJmldIoZmcPLVcFWTAflTW6UUvcfhDp2Sf3f35z0j1H
bnweG1l8332Y2pTCvFUSqqWKzZzzxtnN9IwIALl8/YXujcIyiWDKaQ9NKDMtj0TDD7Y37SAVtRdx
A49li10Le6zI1BD7QZkBiP+WjmSLByASVXGvq67Q/aRZcT0IROwdyOQorSAbX6tL+CP9gvB4TlJU
2hxPwdLtbxI6w9xCe9816fu78vmLaxnAo2dv/VQcKbXByenTDf8rrp9HXXpk02F/iHYQZ5L0+9vq
0FQQ1Ir0Gr6UTUSL/kI61j7a6MjYzt7/RsvnsfKVDYaC39VxdrelBH1o2Qw13vsibfuVYRsllddt
xXoJwwivMIFgLXYT6o8QnqCAXL93zD+2crUiJmfF4WlUt3s7CYce1fRNxeGMtFqOS9xzSnMkgQwv
NwnxBH/bNQ4iTqSS+DtoL9sA1BqUSacgXKXpG8jCo3947LJbmWc7wFJ1jTRLHbwiOBhzI8Q/GwfY
AnRaX9e0kvIztt7n4K1eWt/95aA7c5+0yKd8QvJk4YstWHrc0NEYTFMkYTMpfMk3s/RyyXA6X9vz
oLnNHZPeTzhBpO1/YEmjK/bP/dqxFCfadbbI2QF0sQ/4XdWK7fYYhGPsKHOWs1G/D9zlUp1Ww7e/
vs8bULb/biQ1WEDcTIoFBok3T8qSK9Sn4m4E3B6VhmwXDLcF1fOAG0LP3KBR3VwPneQ+WR0V2mAP
V5lknDYL6Q16dm7/k0hl+v3mNev7RaKipcVpmVYHCjFBPZITV7OyKPxYOfoWLGKWp5EPxw3nq6wR
7YsU8rHKTSQeEZhtlikXGxs2x/HWCbF+U2DzbLgtzuiVbkIOjXPpjJPgrQkRDgU36+H/vfFsTFYC
OgvJVaGM49PopZBi4OzP6xswceRhz9Bi4EA2vZrw5r0v8cCrqER5fHJO99imj0sUjXyqQlhH9zVP
MrJte/XI2VvRNzNV792qQbtKP9eRV/f3nJTHVXUEl7HepNG+2X7+cNavBmJcfzDw8INT8EcL7ElL
UtwvEHJaZIYnUZstJgFMES08aJq91LniXnoMPeHOkUiLmaEM+NpYEyL65q+MyWd89jpV9JiBkqQQ
6o+IxXuQqlfMYLhkWt8uy8vIpzwAPMFg1i7EpQ9MP4y9VDn6zvdjeENB7WBPdJ0zs0iAKKsdUyuz
Qb3r5+vvRRtkzt9KzEcMHhwX+VQZQ7RWxpgm/WAqs3qvs2T/LKDRcALIhZecyFhiAHYoqMT80rHY
u2f+1yVId/YrnRgtM/ASyy4sup4gK2f0V3q+rJJHsM80IYizmoDnB0EyGSHqR5w1J0vzJF9Ri8lT
sDtqwETrg+49Vj1123akBTpG+o4rvGml50HQKivSN+M7Z68qTM43Gzbk70GXaOu1MEx9s+/NLFhi
g430vCYIplnLOTja2JRzpinbZzwbB1W83u2YnvCMlVvJ3FsUPGXQeVJRpgbXoAJi0DoBz3t1Qz7G
dO2SaSn4qNDIXyZ/xWcJ0r0Zi5JfUKw+RNPGq2O9faP3h/hVFT+XfkOev9p0hUoXFbu2XrrjAyfs
ngxvdUhoNK6nB/ghwWmgb4LT2L1p7eEk6bkmjacOO0RKTl+LOQMK53ES24fFZfFF09TSj3lIW+E8
SS0bojk+6VKEUYXR8ZV9QyHUyjbOaIFCJJb+VWnfZ5IeGL6KmCdl9VzN44OHS07LGXWVH6tY12c1
/jPy/E4Kw5no0Eae/7kHf7bXicJzKE2wlIKbDGx/UHTlAymmPP9fRQ26jsWgC2acNMc7hxtsg0PB
28DvH5DAPpeljkTixWuUkeZX12t06Rw3JZvdeOjKAZcMJGc3ahnzuMd/t4zX+X3OdAMU+fhW02Au
lmz7ZSeIfrhJLk/z8sMhQETCE0aBcEUaAEPitP/knTYUiT3fRXDmalNEzywny6QLgBGbnGrgSoh2
YpkAJV9FtfCrown36F01ay0GHzK31L9PrSwo7/L51mt6z1pkUGxwV/9CpKyRxq8vQlg2wZ/xZvPj
XMJxKGGEVAqiCvMJpkEPvN5pCyMzS1rkBbZS0mXcEcb9wpJIEWgR9fyh9nReND1sRoTGcjJw6UiS
eS9mKgc5vBjexEvpzgp+3QSOSfRT+Zw8YS1aOrdFhgu1vjCHyU/sioLqJ0nwJpYy49h6YOqcFC/S
I3atGrSEfGvtUxq1AR2v6bQuDTPYXArewqUwWOgglWpujqH34N6g/klOVR9XksYMP0OScOyxg+/u
SQS+e37v2/pBEkn52VXwGLCGvuQyVcZSMiaEGopQr32oHzSRkwcCR6/q6Duxd034bFo6TJrLcURt
VtljCLbufSRFGkwAXWdGbBWEjN7LlflxDysgFzBMB6dPf9zzjE3b9HZr3fyFXenQD+k6bTTSb/oV
9sd0tYskqSkTlCEIo54/dZ9rjmKnmk3/itHpUD2oZZVLYi7QKHaWd+znVn+BoQAnsmqfUnvYqcif
5bf0IBRjaO4tIuDCGbGSWa/m52fJ++sf/LVrhhyBtqh7GqGbvmQXthLriHzmdo6rN2y5jyQysRNw
TbWYaxgqWIRIgw5GcuzvpRDoU4/R6B/bo4KEA2quVgKynjovaIuG0eJjIFjSTnpPj+vA3cjrv1w5
OcM8MO1AvOmoa3JDN6kHgUVWXkN2TFKIffbFp7ejwsoWNQUhylr+IZIlFQnKZFA2V+DPTRMoZJyB
CHwOYieGs7aNcKrXuXrEwDUi7iudGy4buFy+8PyIOHBO8110rXIeQn9Gtnz+5Kpd2R6+Pe1a2zHd
BQGpw09RS3GRnw9wvoEI/QZc6I9p2BudABf3YfJPx6oD+8RLEgCjCltS9IwSn/DEFM/rX5c8hB3o
+maJ1dAdwwvE78CZ+ahH1Dr2dQqpPOly0/WjwVER/knAVNjeBBJqtPc+uF5gUUYFPw29Jsks3I5+
6GxwDaWMQJINmlcxHbC4KmOiYMEzS6yfFxNJSEFa0zEIv2XtbFpxN+IahPeO1fX5I/W/pqCWbDq8
6u74Dfa5gwvDpDYyub/v4ZFuAj5cuUf1jtrBe4Hjo3Aiq5ukf50CqskPssqQOmqCP7IC18Mk6KKc
34NMz/0Yv7OK5DQgqmzgRg51+PRbk9WXYijyB08ZMgliuORdY1Rkk2Y9Jkt5j94/8W+AbPANWO4l
nspag5zqSHT/C3+/4+lPn6P4brp4jOtA6OLv7oqlCsQmf8pYd/mqYZ61J95hj4nXlDtjRAQWKlRN
CJy/IuhY/bB0vKAU5nFNJvaBO6FCEOYKUeueOq2/qNIMlIu0rjP8snQObymPpBeh0YM8lHvJohCY
ykcUiNl7Hoj/7ywwCFiPsA+jaPJARyAgpTBXVdwxmJK0J8+OBKYZOg6qETBtdQkI/v5JS6q2JbAd
oJw/HzAamY6CXW5Mc3xcrK/kHX5czI9Nmtp/dtC3aV2hwVYt3X3ehrKzRYsriPsMtUIXR/N+9Xyx
pLnJsG/FEsnhEI217fsjpQmWYcf2OOBEu9ip7r3q7tEJdZn2UQR20ZcPjkOHZXQf0b5rTHBQpmEO
H5qaDpBXgZS6WF/nNsgDD1clhBtKzJya8Xa9NjpFIC4/VMX915DhhRrtxztovr6bXwzOqZbz/E3v
lKZbK0QUFwurXWeg/aL6To5duzPQ7LdwYuBneQ9h/Q1sZ/brRzXCgOujjSYXv/qDKplRk/Gtv+K5
xc38OK+AIs2tzlKB1tA3VGmg0xtT0LR9z56w59B698irse0zDVjvp8AFYQFBdOJeTVHsY4ZFVAp7
88FoCw7jqWSnA8OgDedM5ahC1Pjm3qVi06Fm9pxqumCHJ/SMUQqAnbaeJffld8fs48W5VeJz0j0b
spHYi5SW14FKA81l/ETImKFEv1K25TUSfGoyt4l7fnqfl6gJtQfPv4lw69fTyOzMwfXrcb6Vs9WS
C9YgzPCNhBUBrNC+j29oV5z2uZGV3+kPmyfzgg2ojXGCnR9yUM8+CoH2Jbpi4LhBF+vxE+qTXZrz
/JGoW+lrreD7PQcyoMjP73GApx74OJnNKaZRny1S8jXHYuXUW36TDzrJVCmtGQnSqVrBCyUqrW/4
G4SW3+c4i33w+lL8YMYwRCPbcuLJUqFs4JdaxlEB3X13alc7acDy1M1P0pcextjZsQAPfytsOTJ9
lFbvAqbVF7JKsz2NOmMdFd/Z27nGaO1ygDf6jA5EWcjd62DmCwtkYqbtyzPDki5kk3hCdsUe1pdR
m1A61qB/ysdP6L0astq4jNw9oOsgbI6L3qpZlZB99nAPbcyAL3Acgq4jbHFE86ZJ0nh5TS3NrOBK
Ot57U4x9Ibm0YLiO/vek73DJKHEFOMqGCrq1bfhRlkX0N1EQoQ1/i1ewyH5CoSUY7JTWAvUUWZ4b
g+nbUuQEMpthYOZNMlEZqvumL06B2FwdaKrs4Z+d+vx8mzo2OQwHWW2MTg4AOEAEC030FTjVaVW9
EvMk1hE8QLI0IgcfTh0KU+dPYTSmLQAAJM8MxsQ1z3ecNVeMb2P+D5Qz41GFr6hsVQcJS8slSpEI
UrqHW70RV/4tMkNklZIV07Qu3EewJ8Rf1llyE7lSf6leZ7eLlu/D9A1S/WsCqZjhjBrhbLRDP+HA
lbpq0xJ+tTZi1B7AoOZ19TcOcYvZ9KjDOM6Y5gfTVQybUcN1N7MvRY0+0j3d7awJCPg8hgGGlUow
VGDJnB6P81N4TaIwgvUWNIyz+l2tgE28e7H/NFjUDK9QRAgg4m2YB8+sLVpR+gAwxinW9/U7REg7
qNut6c788hB6MYfPCHhYv1oNGXz5s0GTacUm5RL9V/mM1NYeldqUqQzcVh34VbNi/0gycSoFj3CY
JXVSC6RFTphyA9y1bjkeHlH2LB9tkCYs90hMvbJvrx0MUY8E4HArfMR4lzRmbewSf2+6hz9SyrkA
GA2K8f0Vhjg3wVarGPmpQzHPZ7C4yjonCpn2VY3ka2npdIMNNnzKWQkVYK6By9Ihu26NJ6SWzOTB
79oiX7wRrhQkChlI+JGpPjofQH+pYZWJXAE1bbN2F9LqQQauMFRX8X3wn+KNWFxqsHVE6EOlwYm0
OIeJGTmkDnQa1m0A6uSGlBKp1MFDM7bfKZq10L+MfuTj7dXFctORnsJ6uIXF9US2YiXKtCBZoByc
sG9EiZN1mYR4lL3lqUmxXQQRHUAHHNF25QoyKAtnj775mBxLuj6UEQP6NIVeheCKMx6NhBpRXU6M
udtyqFM45dM5euYL+Cq6C3hVMh9qUVxtrEBsCUjUQtTWQB1O8o1kHt4kUPbLjAMMQRvJM/JHQ4QA
ecjdsPTSDmwaD/+mqtgIe2R3E+s4HT6jh3cMCsQieHMy0MtYfg4gsr8VtW8xj5/6C8HfrIrqUipB
QQA41T+ZUA/eNfIk0Oy/WKk7iaskgqJNJ/wjAgCRXhVDBGnQ7hQF72XLngHuJysX4c68SVrLPbig
kBc/EKKwA2jo5LgBRM2jUgYmETx9YbxN71GTcetPZiPYG8wp06bWV9L3V7wp2/HPgQRPOEd7q3a7
ZbsZKX9FJg2puYWv4iVsWc03zDXcFRs/wCdyOaWs1f5Vub2af+opg3w+0kHpIwJYasX/kHWokakB
Vs2fKfs/Grr9J8kaYP5d4PxGYNU7MssxjLmlA5Hoe/NWuJAixEEL9iEuv8ybA/VvpBX5L84DbP5v
cDn/cg2IvU4cNSF11l12iXqtGTDrvM55noBMvxiLdzm99GaKvjjCERrPqUZos+c7sfQyZCJCltAQ
XPSH19pj9jtSkjuHX3DmIagEJmav3+zCBg1JQ91jvsuIm6Uo169Z7GmLhIORmS2I0mYviMr0/jTN
HjqzbDJtAWmMUOz4xNjAaDVwRDKWWFlDhfZXqB94mXaxbIDAKPc/c31Qc0Q9MuptezMaBOldMhPa
DL+4Ix1gJOTubBPLsYf+Yhg3H0EnULv6ur+YiXa73tdwceDnknAsGoHHzdJg0ruhfZfqm5p2PMiu
HURBfwllHclVsCbCchROFA23oIjYv76GGUQHILGWMVb7OJLgwPCRqYxCEDgWsIZuT0S1riMFnk6l
0srr+z5fIGfbRp400Xlse9cQ7wGJ/CLo1S7GroUPDE/icL7Q4aFvHShZOozJrt+kGYdDV3z4rDJb
Ue5GM8uZgJCgRtjIz8rVWFRLk9BCzOXMO1XeNNyByJUpMBnAeRyy1RMcDmoEesvoZMRJDutclpqX
m3QWnjMeoMRGO/XqYdWPQItBHw6QzUEu3Rk7ok6jvLt4MXDlahRVqG+nlRM2AsxkSlgmOA4vHqGG
LN7fEm0cygHWCe2ARF4VSqBeSoheXWUOKZL4hU1LuzcKUIbqZx/zUBElxA6ZrRK/zIt7zjjchShE
9wvn5m6VgBd8akWu6VVDemKExFM0rmA7qFmkEk5dg1drKbRhPSosrUuBNBooCqPjPvGu2QbV0UD9
zds1W9oX3ZeQ6/AhgZgOovD/roHa+BST6jkk2/vjKqbLaC45zJ/+muHnyrzL8BBLq4TyVwYYerFt
6Gys7fYkEQ4XyRzcdrZodVa2XklaMB/vv+NnCI150ikTYByms43SWiv+OfoUwmiUF83mWxcJ75cU
NYzkAPfXyP43ASrrfpV5r+Fan1kmm4ud9ipyRBc62OWNpkt4AtuYKfy36Wg/PmOLK+eyPZFKFAYg
+Upd5o0dMhETZbQkBREhvyUVvcS5HNvaHQlaiwmKEhvhJvx39dwLSAB/ZK0CyK/AZomgG+/XcLsX
jwvWIbSawsCVViusdj7r/IQS/aZmVk6FUlvYIaRHZaPN3ywerUDyROjs+7DBT8Ucl9PAhpWlNYTS
y0Vwq0fOzj1I9RwZZGkWYLSnK9jPV+7geCm36KimW0/rBeJlt3l+7dVVWJzulbOjq0ixMlZKaLRQ
M7NHOSH50LyvXY90bKP5gIusB/ED4ja0JkqTIB7P8GNvz4KaN9AzGCoOySFm0OU3UL39/y9VbY/3
60QwFU81a9Nv8vq/AXyw5Ff3lsk6C/sRdBqCGvkES7J1kytdejpKSos4gX9hsJoxiOBpGVrMywjY
jPbycZNyKGVa44+0qs0hUiGdW6OvcGtyKwSXJvw1riImHEtR6FOO6hOZEZLejU0SiN4qlyyqIMul
+8TMthp0+dYhWUdFnrO4PxbgcOduTY/5cqAtiVGmZ4GMqNt/TArebGwtiW+zgJ+yf+TvwnHd73ge
rE/TkSatSorZoWkx7a8gSFg4bv4/z/Fk76ga3+9D+u/HLjql3MilNEsSbOQBwltFTfS237ZcUFhm
PfgiSA8CwtMHvknrmdNIBRxwZjBa0vXrusFLoiOcOwdyBl6vTNULM8I1CZY1nyYKaiFlxqUx6y9b
huZtAdWJF0N0d98vRVe/fF5TmP7xgylVdpnsVOjvssgI3uZfEekTAKWGXZ30r92bSliB2Z9GXUVJ
OqRNL1Rp0y+kAPEsVm+pHatjuQUVNdF0eAyUGeEnd8S/kTies2+IUsO5TkW0bTI2pB3+sfoBEGqW
vPv/wzLPXn2JlhbJ+EjLzxnlgTjuF0+iAreKGzY7h8N5CGHhSnaikLFYc3cdceZBer3kAwHtordU
TfKBKbmR9WtycpvQGX7ygZxK4CWO6K5S61uNrV0PNa0vileHU5CYear552w/Q5C8i3brx1WO4CjV
QWrNOhL25hp7X3cOMbOBOna/J/okZnDQH5U2X1a0d58/31kOoZ0HKpFMzCZ6ddmNNNJ/L77fyvpM
T9TpYs6iapT6ZwsM88J9LCwBIj7mp37x0dvxWiJAnNrw/f0rsJsaJlHVKUqkoKRXN5tI2A5fGiPH
JdN37gLZNHehvrOkRqgpBvjXMm6yfgbXVmF1YPY7Ca5nU8jwfQnfwUKOk4UQPKyx0eelmmDOLx6e
gtIy9mvCQe7g1bcR6vDP5SuVt3QJfFFfSZ/hL1D1l9WWZ13l9fZE39qLOASnDm5/OGSAwcFHNM/w
xLxrwQRhivnE9aEI3Em9KaDSrOXlomOY8R1EVIbmF5/qYMcRjv/fD93xw+IqmJe6bWjgvZgs6+cD
COWR/jditmK7pPVNJmrILwnWaJYHf81qenvYbHUJPcYYtEWZso9VuSbm7Wv5EnjAb2GZHWmRjDkn
kx6q+VdulnjuWBaViZSMB6QpCTu3IUpyTkSney+VVrVXXpFRSPaTpmS+6xQOGy7DM2g3DooOW/Hk
7Xn1Ehm1QmPtxTacG1Q8pFd8JBZm4rVpWUIzspbct5/bcTScy3ZZ+Cx1C53mFiQF0N6ZffPiqYOm
pbnS3ic0GVpdqjJS1PWhXlJcBtIBh6IQBGy3Rb8fJ9vQypDwOZiRGVvzi15ZK0dMGkW2u09UPD8Z
Fy2yaRre1Aklhb8qLH8rOCC89s8fpXid1S6KiIuOfftzunY6dvcF4cM8/pQarwKUzpYVlgCMlW38
ruoiWsp+FiFdDxDuzoRV4HoPnykGFkSiRew/ZndipsWwVf86mEjOMI4NCf3bA8eqkiaVwT6NQTZ8
n5774o4PF69DhWUoGCzNRwSLwhuGJnr81jwQhAYthgl7IrEJ7HyawavVoD4cglA2W5klVqf7UgDI
QqaysOZ2xqZw8xbD59IXCEGT6KVoNpO4tnyLn0+dbzs0TYai96esOl745cOUeQQkDtDVvdFDtw2n
0FcFZ4slschOGwgnh63tFsNJ6OdCzFglgy88jw5pQPeGTZ4RbtxUhS5EGP3+iaodABFCkSBdljQ9
xXb51nM3ty13fcI3I4C4YhchPLL1qmWXuiVWBAvIh7sAJXU3EWcdeiiPVs+TCm6LVui5rYHnr6V6
iJuQdNcv87yfkEbQ9VF1bC0RObe3loRdGYkQYmB7ieqlR9SKfm3yr9D3vkuxid2HbEIO6x74GADB
26fnZk0fjCHsHVrmjENAcJhoxAA30OLSNKbuCqySGLIVZrz95KWX3QvvFuV2ag3qlpfEb9QkdogD
ghng4XXY9c6p5At9YdHgCMlkQal62Ebt4elJrv8wp3bIqvX/GtMtoxCKgvriUSZv0AdEBtbpOjwI
8xhzoSnIBLd1lCuYKFQYLujDH1Jf2EE36qPfQFnvuP7no/vYV4XoO0Tn3XRwJ+ZyuN/cRA0/dWPb
ydOW/YLouDTj30PDu3D+qX1uh1CiRqgwzpAs9rkJLjs93/HyyTcw/aVAaB+Amj89SLof/fSFKxag
auikpqjWA7Vaoi6p93uFB7+Rd5jB54+b27u4EATEgUM7ZquBLifq0O1uagUhKdgi8ewIXlckJnQ/
E8cp2dS9SVR4cqxg7dRX9uElTeWLRo6PjsjHJJ3VaAMXU5wMyumpleStC+69Umv/47h5skBc8e88
/uGHxl3DLk5KL0byhkQBdQyOYIdrgRaEX/lvO6SSrQG5tsbUFtaJfsije11gZv2FEok3bJq15fAw
pInKzD0Bc0YkVRg/vhL/dEUUW7otSndTgmtTISWX2GhCn5rgwcyruFcbREH+LstSn89Iv7vAXH36
yP9dkXqFs27k8QaGNnPs2aMfpEJ4aDAp+zdZpihuH0shFv5451UfGwchFfS8781sWuiT67ioV+/+
uYQ+oQJCJkDYmRBPwKcb+mYTILFiRIYVo7kwPDK/LO+6/yQN/xUq2aKLNqR56rKE13lVlRAvX/ad
XtqRsRRd8HjX6oaUOhsC6ZoSFsCr1yxjaaye3MXxqCs99KI4pQAUBsSiPFBIUbYvpys8JP0enpb0
zzic6my1PT1rGaEWG5lVRJ4GzLbUyfX3+a6glqRme4Vpkx6AsmZbQlZ7rt0NzSv9pSNj50Ry6UOP
YQc87uImYyW8I2aX2Mqu5/Dy7r1IL7UyaQ/yB6NvV8OyGiVdgWS2PEW+AgqNGogIN7ZkzimZP+FA
fNpbx09Ol1iOAa5JGE2vgl3cK4jRqNV0q/d5ZfS01b27qrj5ZKiS7u5qRR4artol/4JRcNlQYLYl
1LLjeJmgP+CIA1uWayDtGZXtSbhwCkDq6fwWu3E2x97mB4h6HSmaAYw65G4YSKf3+tn4usGRqvra
Tbql2J/fF/b1sciYFEVUnRhtBcqHlXQr4BrBXTE40UGMuCAjKu4BH7p+7l3n/fT0nI/+T7514r7Z
nwCFz50JQc1jWPkHO2VVbWFvuNuFu3u6Kj8NvWbsnmiOGxj7BwQfVcZPGdEPjvwGPg6FBGkD5Ona
LfYBC16HHp47h39UswAtxAPV5tejU4xbCJk2s7isefXVqiznFwYhQEM2C3fKwuiC7MA8Nfdd95pP
GvH+z+qcb53moc/jNsy4o3IIqyH5hzFEzMVhdoP3FJz51RhsWHl1I8Trb52VH7QgXNpnx2Ij9y7A
u70EpALqrYPnXTR0KusczpjjSvzBJkUmjJXcx+GKmEdJWz+KwJPqvgepGG89DlP0mO9xkaOQC8V+
4vMBm8soLL3RXLAsOrLAmSyLLn+F2ndga7ruOTe7Ixiz/WPvpSD0XddZfVjbQx3s/9zY1kZ6Ovcm
PPsh4hl/fOwK9YlVLvUtutA29YQaHYwSs2SJbPo6t/9cKz/cky5OAXfwcJHDQBPjGR8LXkKS6bkH
jkDTvlhKXSX6eTJb+HRA5O0uYF0+ulp0KY44HJ+KCoOeA9Vw97CE5wI1ZQ7Z/Czn8k3CFXZdqkTy
oHWRDR0MNH/wXyXJ0rwlZkxc7Ri5yGDwWnb5KX688cVC7VzzAS8UaYqj6WXV7Iu2HAXpQJ+RiEIm
a4JXWrVyz4slME2R7McBP4OAQk3ICg+yuv/2oVfzYaFPLK8vAfOHWULaO9Db7TeqqurUMpDASJOB
OhmvwTaVDoYPDCZPNhQzl5OEV7zxeH4tMg7NRDA3KASa+XvH4EgEgaJd3+IsdB0UKg3wD50hEANM
nutG08eKbwlOvljknJ8HkvdES/inXfgTD5+ChSQnTVNhzER5UzU0Xc/8Gr6oSpnwdYASPw/EjGXc
4nwe88aZ45+0XJEc35Wi8Yu8w8B8JhYXnown7luv5uXN8GUyqW4FRdjWaiGPoNSWHnKgsir5G/7J
WetmaFRumLxwPY74E0E2ipO84xxA8SauVUNqwSl3WZgWOv2GmqAxMTbIs8IfP5WvQ071r5qolhgc
SZvsZbTHTtpqy8IJCxKJcWzLVR+paD9SL16n8QDjLA0AxY3GZo5fWbik87KAfhKbdXx68gyqfonj
gYP1wpOunvNdlXtjSSYuAA6Vd8nMykvD0unkrasveFMXswbt4/ktR29lOqybJrJOO/cH80po3vzB
SCidpV+vG2njwkomBVq4t1BnIeYyzJ+TQ+doWcX0X5H6DNDVbF0+/ai092arDRSFztwLq4XNiFX3
TPDMitBnC5hBZd/sOqkelP9whXzWR7x24HCycXkey1LqyY1DRUy8C3XtTfh/2807TnFKmJZaUKxH
8lh11i+6hUcabOCD3i0Sit2ltnlCX5dtdMy28WmM+taCx/Gvz3HW04TtAKIRS36mtVU4jYvua9N6
9artaFMiQ0OFA8G7L5nONOokYwyXPGu3pvoYz2T0HlV1SK16/uPDt4FtEQQPiiXh47zoFvChGLEd
NnF7OAYG3Pz00oC5oSo6I4A9JoqlXGC47i4pqajTukFj0qluPcbGdNkhDjQoDcZEcHsgFVOXGhlw
MPo7wTY81tNn2eJjRZBwEJmQmhil4CbfbmsGdWu2IQ21FH3xLfbxadGPjckr8BX0O22yh7+C4oK+
hsw6mYYmB1i7wxAzvAAcqFYTWVOEmSDBdP1/urQ62q67n7BxKIKbgsDMMzoyyxdB4W2zJEUHDXcz
oElLpm7vLg2XSl6Unr3ciz2uqge3+fDGSgyMbW9T41YncqfABEcEI2dSXWaPxCJkrBTdKS9aZanN
aa4rj877tiO+/J5XihAXlRwmMBtqZaFkt6FOp+mKu/pgyJCC9/nrWk8s71jIBStSgAjKePUiZzTa
EkOK80H2VZocTbVD18widyQxC1LRq18U9bjwx5Gp70bWRNW3FBjeqj1NwsOLOWaO1xtttsfrZ/rp
GtMoWTXfzsJeyZQhcx6OxXitUDW/1rVAUAfz+ZhqLNuFPjLwhzH5+0qQ+uI21WFh27HLxawWJBof
KgS9MyEWZANbCIR+YDg2HiZdL+K58JZKqFmi1MoSyfkOHA2UjX2NLmHWp9eS2F+XPrj5hZThNOWr
s3DYAyyaADI4ghrLOddRn3TJXmZ6F3Xcu2ZVcPaLtsxRUdugtMJCNL0RIu27MFYUXyK+H95J5oay
bk5EoJn5QYR35zGbQQhDstdkx9ouZBupkVRdFDzHpPsVB4pHZGgq7qka+OmqCPjxyhfe2cPvFnPs
xtwM+bsQu6/Cyt0TCFPduc2pEl7KKoHuae11gfqPl/0Yb9ouYLSAVVYACOBrF1nmZq3helo31UK3
jeEvRdljXxFG4nsurnlvIQQB7mKSohiJWifiwhYlbY6onQ/SYyl4r6fs0mi8677qdqYlx2nKykyM
Mzg79pSHMIX5UCs7O9FIsOq8Cpf0uVKS54xcqPakxh8za1T8cEnkGvGKAq0si+WkkiO9gSF77h4X
r0FvoNBPLd67Htsb7ftAzdyqKp+galFVmao5FLOnlilkUcJs/vaSRnzSMOu1XfZjLopbVq5eHT7h
18ENES9k/Cl/DniwBJbt9tz9JksY11ohPL9pPtChfE/B/ilqWtyNBj7FU5iMba7kDtbxPk19MaQR
bHVRCDRF+vO9qrPFBKbjVp/L8AWAt+yA28aNheG21VLgLSt4U932Znjj7U3lNKt1cfSu/6bCoimV
VuWaJZ4ExzWYICaqKXNPpf0DaHOZ2NinC0C2MHlzKYtnGtiSztxyNXPpnDxDP6PCG0SoTkfSdZK7
U3FwKSypjscWyaQGBwQ5TEz71O5IpufMqrKSlJBmpxjvpS73a+hOEzC8fZOjVDyGwP2DhB5A9I8h
FC+5Qr1t3kUIAElK1+L9zYrjdk55S1H5f0Az5bcPX5jI3A9x/3pDtmG0Tr2IKH3mxb1FWNFxBQcO
5DYh9EGmj3sWTcRadIGd7T08SiV1VwQBPGK6gEximEMsOV4hIaiBb1dVzQ3TCAYqsmRkssdntNa0
vPemz2fN75Yr8mvnR2XVkNHQEU1XIJerE2NDVS8KMHyHCT9/OXI85DdmdR6YLKMqC/cHDL3Eknbg
GvZUw8ztxKPZIC4PlD/JULePOtIPPY5w5/f1/TXx60Sx3Tfq6QEWOIjKxF7P4i8Se9jGwAwdGpry
hy3E0fuw8S+MkS2nmJbYYbaqAWebnEBM+6PK51TXdNHF7FXeZzRZ3QXt7Cx97Ku9sAQNYr221iSJ
uZ/vXQspeZ4MSsU4nSn4C3bLQoio/HJDuZxGHsXJ8/7AHVu/hrSwdYdLMTbphoHfdgoBoVoiMYvx
LXnuybzH4nqte5Vm3BUcxdKojV/uI80uTkhO/ZjTFRGmacsewbMq/JMuGa4QGM9Gp7FNpirGyZuS
rJX9wlXyD99BkMCofC7vRNSbKr1Zp9arKQZBQaYCz87DPyB+Lq9I2CerzfcV/IScpHpURf81S00w
XSKI5Zzn7nfO/xxYDvbV9ufFWA4t3S+5frvax8hx9FmhWnMBWxuH+Tdxcao3zbjudec5SIapbnBT
6lHwoc3QA9NzmMust4khcRD+IVsf67z+r/LNZ2B2D5MiwQ3xaByw1ssWMFHzGNkUldxnUNujDeVk
X8gbeCsvhqNCWNkKO1Z1H5nPoR7n+CdZ4nm2STi8YhT+bACSUxaKD0NqjMQ3vi4AcjKgIUmXJ2x5
JrUyz6GEiwdNZAFugNoYBn+D0pg4m3hrAouZeQNh+SCWY45bcZsrH4EDhLnHgKc2whkTjEf7J5OW
dz7zC1HHgVBYhD01/M/KDeYrKIUlDtRxfyREGkrjjbBAH8QMTATuM117pr4DSSMsXyWZeeciW+IL
lcE+8dlYO2tumR9LN3TzgmgX/B5E0JGOWjEYfeydrwEKpEOtenuhgQW7VxtOjpcTOgZNK5k77IT3
Tjf0c/WHqRnYh4PQF+zJ/89Ho/qWmMIkdNZN4VWqiC9m5GJ2QojvgHP1Zbz7ARRPQDaqZvVYyv5U
DPiFeA+KtFv9+p07DM9JE5dex7ByQXYw3ZjD4HBkxh6KCIbKy2KyL1L2U8b4FVb2ojIdvznK324y
mcBH5+Tes2ifcJqjwq8geeE9ZO1gs+EVxwJ2/XWD1/bI2qtekrxuCnp2sIZKAgZvVaKysx636tP5
Eg5+mXpX2NxvUixYhRfFFjjeL3Sbu+39jqc0lZVnoBuDh2KsTl04j9oLbr/CmcA/E95HCWA6Jodh
B3pg+CIR4R6ybsnuEdsM02pEMSUPR2WkJgFttm19HDf1UqKSzFi4A/jBWNCRb+M8swa1GUWdFn+/
QBOa3Hshp0LDUYomS+pnJ90D129BGupbodcssxOo8EB1lR0XmJjGpyNv3mPzScvv4conXGlH1/es
wr904vUf9UdvJctaMVZu2SmDNPUpN0NwUiSFaGPSKzntGmsXNCoNj5OZd1pZXwdLoddm6djvOUSE
XExAwQSM6//2NgWLP/FEJjQLp/YGlKXc/QxzMLudaazBURatIa5nDQf79wYzApttORZ2wz921BxI
fvoFzjNrnqyRyHLJHia1/cikdW/TfIprd7coDAgtX6Ix7D6i/AbfsBgRbT8eP7xWJ3HwSxZo2u05
Xs80m2l8PxrmZ1pu7D5SkM2ZGQ+c0pY/HXYp0kqyrW12Nis4N1bPS4sdy2yHl7Gv6IVdUr0VhxU3
55Wf4/vORN6hjIaUjm4iym5VOH+EyCYSI4TeKGTpVKz8QIu01Dh/fI8f5UkG91K9USlkJWXTUpSG
enFd9cKQYpzEuFiXoyx9QyD+4Iv3iw0R7/QSzbC/4+4SsjTSlZiNXTyG4HrG4yC372IH2GCfKNjL
YwUlDnkv41X3D8cK2/xZxjZgI6y0Yc77ZwE/LwYSzOiRH0O8p1Mj/mByiyDaU3QC1nOTL0plS5y/
JJ+qb4JmUT51vuMrh2d7QcrQcPpddutK/h9qlyzSmeg/2w8L1W60VlfGyuaeT5R7G9rzvBpeXK9x
mzqlqV5ffnPAwlhLelSyNRlJ5dMwhcYxRUs1sMTXXl4V0dzrZQNpZ+xw5WnysV0dRUcPePmjhk+D
94U4TnQU8ee0kZaBpkWI4idxMO+U03eqfyznY4JViwHTsTq/GtbtvAQlV9IAsdQmCbptPJgCgQaA
nUYQdtUbSSums3araGfdOyp0mlYCZKqKJtRQFjzCNrW2K2y+OHGsqkXdRNaYgdqniuvjrcLCWrI+
8wSV4SRlYmOAxtb8v5MF5rvKWOdIQFySYAtkld48MW3Xn5O+Rri0T8/SB9lvNIu9vQ9QYmzVcHC9
F9wCqH3cQ19BYQ6A+xZCBUlpB6PtG6v/EyetEdHFOzJ1+03V8EMC33wbu9k8yV2K+gu7nYYsMB33
ROdCi02LoXfJ3etOkHt2KVYWTff9BsBEgkLFgKsky9KIc2mwGGHt+pSJxXtvmMLDC/PUwGnwBwXY
x/mXDobMEiPfVHLBq4PRSslRomUCkB+pV9RMFnjWG5vvXH6WoMUnYUKKrx52nQfaDpd4iCAoYb0C
XbVVRm5xhV3q3TSl2E3KndikCuXpgCOw0p/2fw7v8PW3RL5YAbpy2u8pf2QZ8xGACyw6W9SEt3ms
k+pHgSCvae3gR5CmnjTRVxwUEy/BNoWfhtrXvKZeabd/ZeZmDLhn82wSUTdjsNBBNy8DXk+XRFTL
TRTVK0HhODmfLZfIVlvbI1oHC+vLjjE7ZxqZJy3dbyPdsBLo7mz7iEx/zZVgvesb13sEHOVVrffe
afXWK6vcOfV4NbBg04PNZiXyjFYboW0RXSE37xKhJXoViQwjUKQzYCdO7g8VyXkEu1BrMxC1jkw+
IRxOafwUfOtq/sIikeJHX8AJRG58rgQ6f8lvbNxVd+mWnBoR+FK/wvMRRiJbA7LsSEyNVIljvpZy
Pk5LSDUA+IwIuuSl3g/bXL6aG5MCcx4bKGYqvuOmTsqcCJBHM/uQCt6znZ6jZbZchuAGLAqVGZfy
CZiiwYSRLq+gBYhIkSYf4ueJ9E1n+EjXx+fMo3lxEUrHsU3u3tmmchERFJryIhN2IJJ2WNSM6ImB
mEKoGrZ/Ex4bE2DNDqUsYQl2a2Q02GUwHAZmZm9GJaYoCH/1rXjGtgE0j+af5Dtvbld/2KSO9A1l
42jSpzqqvXVHB6Qh2vUIQHvHFT08n8E61wsdGTQ78tWXDa6pvC0R7vFxUIigQZrxTf1G1gmBIiDJ
hfG6d0ctuyzJh93xS+ru3wPRjv9+j2tTVbFSGSR6/SYiJpcT0/c+qLhFl4cgBKcq0W99VlCHoqsg
7u9LtvH1mkViDsTQlC/L0h21JYOh6d1zqOCo23mWu7oVNpxzkJGmEiURZ8MuJlUVCgaj5FewoCQw
VwQq4Cl5khYR5jw9cwWT6Dicm1WqRQCJsEjKTRQstyVhn+P/FCHH5Xds03NDGFTuYm1A5h1L2IpK
oRe0D1YGOIhzjjDtZiinmxASaXumB0M7AEY9yUU995XJ9rKX8lfAlkhcpjcREQTpR0GGjLW25VaS
dtLWfmTH3ELg5inMViOI+VtUV95FY93wfFiemKJDhPW8s6a3CZ2HD1WlDA532R5xf+QLAl91qdSR
VTFtu9am07FssZwNkTtgQo2x214sIWTOoTp26n8eXCIRogTvMWX4SGwkQTBZ+C/TKG+Eo1arqc6q
mGIeenbTTwNf0abELz/0cY+YcOZcdMM+jA972Sm/ME6Pb20e4Gg5WGA7vRhmrXEUHZGDQ03gHKcT
DzF5zy6jYnlXxrhXzwrnGwFgrbrCAD3/StUl/64V92gwY8D21Ew1aoXPQ1NYExCeZCHtwPtY772W
H/XepTf37rp0DetsgCmK8CRJl4Kf1NMnbAodymCBq+8pOTLZEWTkYNRBBIK+gjGGiRM6FDZP3Q+R
xanmhqmVAD6Uqd4s6mXwtj09dp6IhvZE+cj5G58G1/vcLP8tf9fGgvfIJI0mS8n7txnkY+EHd84q
XLJGvCQ2lS83TbkViqpoyZgcZnD4fJcmvXhUmgKv3ymcLaoNFLGquEYNO4m49mvsxXKlJ17RT4D7
dkqec6peSabDwiLy+cOOKcXta+UV3KdgZbVdztcL0av6CQc7+Eb0sfa6R4CEopgzz6z48WJxbpxs
yfxATmrLPFlLYOONERsf45buWSETs/2KbsSGKAbbtdKxi2b1qlMx5GrYDCcBMqQvTlIUu5AqYsoL
QaYMC74GLhXCVW2bTGOD6ZPbjx0fEy0X1j9GeXXIuMDskH6u5Upf0PKZIxfwHiyMfjrbqT1ouYxS
9zdf6x3DHClcdCfQu5Z0n6oWJ424UU1tDA0+SHIubRclQ8IGZHBM9QI6Go3Qyea4xNgPy8bLSOYe
p64QScG89XHcHIQ/Rh4gbECETCfDeWrfjiLkSqhE3D0UnCrUmWzVSHE5w4xC1pyOpx47T7Sba5U/
mr99UeNDH4QiruiBdQy65P9fhU2jfVN9/jxFdr6hykWUzWnY0+Nin5+z1VoquXeDSPBxVSUWSW3s
CBe87ONKTvnd44IhDpGFziCgOG1y0rGywYZ1jN8C+WaLe8dgi6EHcDbSi4YVsCVY1FcQGX5j+QhP
UX3B/d1NN1S9lT8xNbWAgrtQvayyZmF/H0Owql7VBwYNkCoZIcIIBd1JI9dFHI1OEypLDRcBiusr
cuNGrJ3HKW1wkjL5+IoWibEeC4QlDqk9JhvVr9G+v8XQKR00VxEwz5/DB0GFOV9xjk/tmdFAT59G
9D0sDhEgkWAg9eEU+TCnLuNBi4Vit9k2ninXLYyBNj/MPFAlxEhzxurd1PNhyEvUAoLRbSheMqgb
4fKr2TVff6VH07Ad1DoM8chR1E04G3acT1i1nYzlSktyG4x+yUfdcRw6e9mQsIaHUhNq6vnhOQUd
CseQjOVOyW24xLMUYVSsMdKbXDOuyCltXoBZIo8xXeZ2AOsq4W8Kjxn/h3lkw9BeQ2jme2R9c+GX
sjhReVsnX8orxSDbzALDT3V4I7zKVvDOwjsoi+ciSIIor42KnpKYRMWW7aY8Z6wqEX4iw9QJ7Bg5
X9oS7r8rMoLgckCUDiOW8gfZHK0narkLLZ9aNil/Bxc1FfLVqALwzR3qemdbVWWkFpHUTqVaKReO
9LiTf0jGYcOBQntMNy1dr1pePCt7jDTRsR5yo3keBhXC2C7piIjkkC7Bpv0POcOr4kqcT61N5Qke
7lAnR8vmHn0BrL/jN/WHOJNP51RBYZFJ2dh9JtmJ4zrQmDNtQtrAe6k0+i/3QYzNBDfQUWMVQB/I
VlxUzlTpcsF5dvnzxDjYlUxHP4tUrRbAYuRoTAB8+i3KoQCR2BVLRebFNmBDwB9jXkWbqCPlzTtW
C7+T+qeeQ+q/tBGgEW6+oC6IbC5uh9XQ8MM5m54hCMCNZjhJO+VIhDPlOOo+8CZk6UiWIBkYpG+4
z/GqcpjZL2zrGyoRuf2+9bqgIZzr+otG5lxfAM+kWab/daq0SSzBu5CoDHJHfsWhZPK/2JGzUxtN
8MMm54o01kbC7QoqEkBxMATzwwhYVzE/fW4bj1ZtOD3qK5M8tJ1rrJOCFC+nk1qlSBvmPodR/v5b
Eag4PRk3K8p7mn8FIcmH/2FVBn0NdMG2lKhLKHfG2X+8ZacyTNj0P7CyN6zN8vnlNWaww5g8303C
K11dyPBfBLJI4zUfZuGSWwqSuoUxN2f8ehE08VCEpnP3SxOihZwhuv1sMSd8uhO+E7Eqp2Sw6JG2
8/+8xly+dufw6oolChFAymJXinGdyIsg6ejmkEiubYLWN3DUu/NcNXm+baXaRMG1DXNweL4jixga
eQyYTjhw7fWb7vINOs2KABQ2+iORuoJkmBr//OVqRlwC5sKW+iYM0OOZoP+1VYPATAuzf/nDUwUZ
82hcvT7P6H/MkOYtwGYm2G3CSUzgBt0LHlRljMdJAbf355MPCa83Y/fN6Nsjo0b14CH+VKutNKx/
F7yDleQCKNU0SCQU0xAdsKQBPpuYf1tc3KepmIfCuSIlR3YNFulYdOBb1pRjlCdsnecE7K2j7HDA
vuVCftHV+Ei9YSJQZ1YsG08AwupdXni6v+hUDIMgJu5Jw48pI972ow62+daPTe7WUwB7QBl8kBlT
6UAfGB6ibUWIOqjFXmv+LrUQEWvrGh/lD9rPRWglK8sOkSHX8Y87B7BVime9jdIVcdZ8s4iiDbYG
kL4F2qeWXPpW9N2Q8Y05GKnpkUfZlQJZLQ27OEEurg+GQkZPb4o9JkllMuhkqDI4BLpIBPhR+0Qy
EllZBkt3yTfElbAxBTNfH1bQs5AXe8yD9dK/X+Er6e2FjZkjK+wZPRiDTSRaUylM4uQgJnFv0sIE
mdv0abhK2of2fIA7C9iQGsFRwQ3IUHuDZKRRbjKagU6d0axaShHWjdzVSH95JcAP/Ws8hbETKsvD
zK2gQP+0uQ8ywJhapdtEhvJj4X8dHhS5PLIejCv3qcolI5+tWl4cGCYqOcmaPsfi0Q4KxOdYee4Q
oopaXR9+sOFk51iREPNXt+2EaymsZuy6ZglHd+tLChB0WHVjkA5wohM5yS5ZLP6yAUtWwnB5woon
b6e+V2mMP2fOiDydK0Q6MQPCOyocLZr9m6Mzm1Y2J++KSPTOUSgvPEVR2GKJ+7A/fm8s3twPJM0J
/L99Nl4QrRKqsh6yx14Z85r4moPCHP3ZgpFMNqMTjn1H3EZHBrpZE7NVv5k3V6edExxTXHCFB9E2
aldp9k+vjJ71a3yEhKgadoecNNkSvtLEDhH26QO35lcwEgAS+xAUaglVFRvcdxPgTTXgzlsDY9rA
zZYjDd1InV4A6YjBDChI+G6KGS8ATYUUDFMQc4AXCm7O1SrQFxfUoj5+Yg+ro74xWTBz8mIMJLYw
gbSVQHXwH+6vT4HYLX72h3Cr8h4n2s81mBYaYVzyLBbhaClGTvuXck/BoUqov740d0NmP9bGoOB+
89O2yR9+gKCYa18jE0+GdPAWP0yEYaQP1QqkmiLzh6oJxLxx4pYlAOJBdL/HMnp8zzAY5UZ9wTou
3yhsb6E+jkIBSJRNhy2MZi0WH5lWZeZ9QzS4Z9pt4x0SCIx845IEcIQKB9Ee8k8ET3PSc9FQPlJn
tr4aPED+ephkil8NQhuCI7bpnNzs1hXdsbu7C/8kYl57xu+Cg3xa4jhbNF3RWDKR0x9i/OnCfCF2
9J1hZwDm5wdODoAQBS57R2x3GT9SsI9A7BdmHzksVTJuId5oHudPjonwkSPrr6m3Xoix6hSARFCw
bhx2H5MDbAq0DQO1WE1NP3iHvLm3pjcHnPg+DoF8THPbaAC7KwKhCVpVjdnLpOF9t/a4A+3Loalw
HH5ZZfXxQgTyDNsdcjGH0RsIi91DL2R2mcojF0xsZuM2qqzoqvKGn2nDg36Z03mTQPQpDB1gNXCN
wHUVgCppE1++5jgsGS+nrVNKrb/VaqyLgBkBBa1TVfF7tnBTL1CMwVxsKcwGuKNTS7c6tjKVvYnf
zrl/yRvjAwywpBy3TX8yZz5R+uON90dwZmOaiD79K7jqmykDaYfCmAvg7vtIp8yxcxuw+HE83kRx
NBTF0SA/uVRDqkfg1Kv/pJ/jvDZpIOQ/iB8sNLjhuA9tH0z7kNMOxPFtaKYc5YsRlEdSL7Momkfh
22qCbFHfxjemovfzbGG8TLy4QfJ93kZX0FHSBixu0aTes71vgLTOBAerPAJqYtwXwnvW0XFRJKja
1WM04574E729v84elmRP7fAoyBzT6KYCdyenpSrP+/WX7XOcuRS5oLOJDm0mWQGfEWLf2WR4nETZ
ZgUfMZkTcysLKWesLlilEyTWS4ROTCxw7t7xTBrUIiWPN7X7WfIElXYoMeptQf6uawX7lBw/CT2J
xY81SiuCuXEzTjWZjM5CJIO5nFGHtYn1FhUxqQ8B6XV7aImSTcYuYwwQXARjuNLc0KKNc4PPjDrQ
2ROYOOgPQvfnJ8Y7KLTVFdBMWQUcAabg7puluchfsJxyIl7SHdmHd/AMsrAjZ9XGLl5zccJkCeTT
5E2mRcNPgrLlfZQ2RnghCN8nOJwHfjc2se2Yu7v8qBdgxYlv233D0KloGmOwhvLpmmYEqJ+HVoSx
5xN52YBt/6BGkzwJAZTtWv1urQjqYYsrbh/mp25bpIkOiR32L9KmV5NcejUe6TOhnqS1nYC/hXGz
JwrEANl1SzGXWOpFt029Z1WPcMu4YsB3j2nbpVlwTzG0zaFKmdOgXRqiU2L1aNoBT6RmItF0HRTN
yTGucS2MQ1zibhM93XQgW7dS+V8beqXqQNBGTgr3drdkJVQQbL/Sef9eclzckXSAAu73rLZpTKbm
fhsFhL7fuuAeaU3+nXuUxHxNMaSeQOUnZUXOoXGiU1llgX3HfBlYwvIWSiiJWd1gs3o8Qg3v3czp
nD4dzqZqSaIkDWrto5KLI7B4iBIy+yfMeGCrx6vOlOjAgiPT5ON2T1N7vcwjvQHJIGOyzQVo7sb/
ddSpdNz/uEVU6u6RtVVsRoS26glWtmre5kqcYs27IOg/jSPiJggT/kOa9coKN/IYsPFc6QPlbX6J
KBQ/lsYPXAUH59cBnTV0cFegItILYv2VYGqiUZsAQMuZqKGxsZOZ/fia03YnZUfPvZvdTcrnwdsm
7Bb+wq8SPTH1yojIV1Jn1oaYur0NsGQ+baiG3qhRItLt1x8ZzZf4dkh27kEcsW9T1DvuaTjL1LmJ
NJ3rKU22vP4/m6zF5miYw1AJ2T1O4E1iRcH6L1OKwRCBijYT676296DS8JnQoHU79p2iT6N0i0a9
K/MQqsmu/1ZCd3oqPSWqrqVnm8ok9pQPXi2zFGXOciKHEDYPGCDz33QkslJ/+z/5hYGurDhKokMp
t3hBNOZUmPQmnPw2XdIouQ8Ff4URL1lD0sTgLhTO2ulNczczg3Fj/PfGzjGbhuR/3Kak4/WsCgOB
W6c+451mQQWjaiNPB6aLIFUFScPryrCX+2SE681rp67LJyjVNSZFbpul7OmCntYMvTniD/jKV/Rv
qhD9BkToB33FwILPqFQW9d2T9c5KeYiAO/iWdEwQpwzvU/0HbZysQfoHKfviPmGuIwfAVeNmXT2M
3jtZ/M5TXQJXWOvUUhNU4wFSMLz9SDiYgQ40WZ6OVBbMXrnDrERqMgAKaFh/LCVwl8Z60pP+OZAS
uNmIcllON10Owfv6q72H9tVzFCRk6/1ruhhAmn0ivyBtTuN2ESZdMb4DodvEL3/aqE3KDPTLxmwS
Lzirzb8lJ9XAavLVjF7hyFoqICttrujGgkk13rT8AiFTryakZdFch/Er/e0f6oeZ9hRr0Gsrhizb
INjuQVHlX02pZgKSuWzs67Ulv1ZPjxjdr3p7gQ4EeMgOve3GejVRxH1EHsSuuBvFvCmL6TQY08e4
cIBuNhssdghCpedEslPnF3ZcWQHvvRJMRpQGv2NUbVgE69+Z7XG+/U6rj2NIaq6Jv5tQ7GjVLvwA
+qIqK+5P4cVEsEQ/3Ez6FyrtWNVpwwzYCRgWUXz1LKGnckA9/B5rqgcc9OeVjYk365amWkMiOp1k
H/kql7XL5l1ZvlEgLic+6xacj9jA3J9Jbe4rqdlmG8BK0mXx8rP1A7C2nPpFi92lcB+tWY4YX5G/
B4u2dBixsFkmOonfUTv7Oj8WWohdNjEeRKlmOYluF+Eo5Z84SpsTqgUXXxD61fjgZs9EHkBOr+PE
4kVyeH27RrBR5TEkp5jBNMges0bajLd9ZWnqAselaJvzzK1935Ao2aWrw/puaybdqg5He95rDcs5
Q5j/7FsAwNliB3VizE8pGc50g6uYNmNJfZHY5TnLlbzWkXWL8Ur9HAZpxdcbJi+dSgaLqN78a2hr
NxCaE9seBNqsYkTeQZVHdpAWcO6kqoZXSBVNyy2nltZnQ6fmvgc7U5c6xul6gAza5oZkeAvq7z4X
kgKdF8HdtmGlmxP/OfFRvsbhLPrTE4pkWWFCtbpyLDvVk+2wQ0y2zbUrSk+sWWg9lQg8++87IWhM
+ETaMZglwKSZRD4x2CY/B8pm2LLuhEXXEueeXISF47O/VyXzl+KM7a2KUd+czG7bia8z3vn5+n7J
8YJn+7TJgsHEVTyJX1gJvbOR/1kE+Kl1KsjjMFHjaaVS7ACOo/MB/SVz0nwJr6hcTpMNhuDyjmWu
sU+JlB0IMuMVjBzNV/7zAZ2DHX7+zQfL2uXR9oG8P/9y3xToKuBN7x0c2hCwWW3SmUU3vDL2k+vx
IQ88u372D2pd081OORP/pucRhHm+fFHBB4F1KGn3v+fNHbMx2w5f3s0IIf4w6pcKJ06XZptLzZpj
gaX/BDTT2ZX4PuMdb0Pf9XCE/F6jVfAfE/1QkXob5S/KkDHE/zxiBKBSjZJ4c9FhoHD6q8YwYkX3
5iuMzriTqES/yQc0vUTkofSeYqvgq9dJeLCIp+hXkPinylqmaiUDsyZaN/fIw2SuZaKor8QT4py/
cCTPPqOXcew95gfaoaVxY8dmLdyOy/y0l4lk68SKWA7mZrkpw7ncfYAm77Vv/8c5R3pO2Ympgknt
OXdGw/MULixXyuk5SM8OzHFUCe/ojmvYD8/rm8ToA2a9pMPjcnJ7atkUaSQuaPtgFWA4bJI8le36
WnW8tbsvTWkeUJTxuMiZJLLe5JcnNHdtePMCUHv2PRvzdWOGWsckbzNGZXDzJVP1goHsbX8M861h
QxFgENJX+r6AfWNseBcun/oqnCg92L6jdHkFF0zIz9M+ci0Y0q5yMFs9W/Y/LDPRoZ1OfRclI3CY
FfE/A3IZaDjFcrc4gfMw1NVhs/OcnH1Q9tYNYlsI1lLJOOnUM9xM03P7fUkMo352BHfHep+y1nhS
csZL8dMrFYw838V7p+WpZHbsHZRFBYMvomIO1hhs3dUPAYx0yH7oYKEYHZDCECLDEoxQ7f+n7tTv
/eTDKTbv0INaFKJuKH8JBB8t8v+E1TPq4PinC+eMV9E6Q0penr03yKkP9hRkGTCVeufMI/xjZrIE
RdNarZO/Mvy69vuAkJy+TpHNfSTkavA2VpuPlJvDokOW/Zk8t1x3zlT57P0BrLtJTHfMTd9zIoQi
wBY+gE25IATyHUxdTlM3PztOjCB0l0UslEHoRlrXDJUtvgb4NVG2wWQZANLAcwwY+7dAIpHUkUHa
QoOjZ7fvh63UxdgOpbgPIYuOtgCZ65iEZ1WU8JSCuYw8NDHJR2TDkwZTi/t4aU3tm8jbBZ85EKCD
YS5sr4D6RqwcpFvkdaj5tAwmZzfQvMucMgUK1UcB+lMlpyocmk8lEgZ/rRnNBziwwMHNNQ2pkyyQ
nKtKar7OifTl0JbTfrd7KciYtl3N6T9k6Qz+AThk0O8OYvNlGw6WSWBwXHmRvfVYYNC4N6pvu9wf
sZzRoV9IzzpeODtaSzASH4vUo0Gavjr2or5RtTPwiZGVKf0lYowIW2rkIiWH/dEDjkdk1nKkuz5u
2rvogpqdeckatUt/1m7KC1DA0/zkzykEzVmoDJOvlXoMbRb5iWh35a8QH1LPqo/fifvtXlSAqe91
KENwKS2TD16DvVJTMWbT/LUS5y8SZ1Q8S9U0jGQz8QsUgvYmDb2rocCAtA16WbzmtVRG5PZm2ib/
SQxLVTMgcyMbYtTjCVqNuB/6ddkZdNEcXwoHCS0WED9SA7a81U3FbW6vbmCrdPWDmQUIWVbe9D0S
67FpYZvGGXhLQDOxA0aHm5hcYl1AUI4p0RHbP4cfgBSl8pG6nyvNsM7XaRk/ojaaTPECEdPTsRae
ftBBAw8+tI/hyuakgtWOvyFNl2sV69501coiZ01XV54JFQjEv3naDq/qlYiMKyEvy6Sn+SFNNfeM
KmdLc22XNN6t1a7kM+VeIPl70JDK5VsLGtTUPrLnBGyWg8XTytS+2ImzwzsgJa+jv2wbVZMFxUOt
Vclyul3AJtJ1FqIGExO8IP7M3lsa5NuMGJmxzEHUx/Yq/mo4d4FRkTL18w6cL0vE41flwIj6zLLA
gf5ZmRrSHfTgskgexQUzdI1Z6tQi0Agkjwuf/xM0IT7LwZYTpm32u2N4aYWMlC6kRQPmpZsLfZUe
qHpi/0YffrP765HQ/vHmakc+/XpH35Jg1dGe/UFSlWW8sNcm165ciIX/4tOb4sYr+wuHtjO5F6IT
ryluqLRJ2r6ztrCWcFj+Hx4WR5ErrFyFKn/ZSdunnhN/C5CdNOlnysLbtGcd4JgOaY4BOub8OZIG
gXOJu8TphQTMWVHS3huJWDHBcspMWIC+wBSEwqhDbOpVcPFJM5kWIBDNSouXf6pvR99X8KRPZmut
lPN06lHjMPWLt6YP/PTJE3zb03tq2DH9PprMZCfOf9DFwBs4YDjM5Qv0kmFiVU6ayOZDRMEIiE4R
N9ZfT1EMBlWY/0SuF3Mp6pt9yQRTA3NDHbYrNrRa3LwFGYiUjyPOZLLiJua6j2jFntABzYgYajs5
1offlpgtukIeSEQPXZ58oNMu6VYbrsjcSKtId3VV2T1aTWdX5HYm+0GLGt4HdJ24zd84FaPzRVSx
mCpcF5spT+JHYcGFeeUD/bdsRPCdBdI6DKPe5gPbdK3ETlpwlWx6Hek6OtXeZuZXd/pt8wSgY3hM
HVEwF0JQHQSmJoYbccPYETyaV1uUJXCHIsv9/y0G0TvvK71h0RtFDkyhkdZ36TmjcMLm6eieyEYt
e+k3lBBoDaz+1Nbqxcm5owpdPPa4EVt4Qzaox3zU6PKCY+qEAMUrHf+9ez54pxfU4Xg2k9qrHhH2
5tophxkuK118Wj/69TCjA5+1SJAWcljUnXAgEEzCJGcsIdnsVFRdnidbF9CtNp6Sdi0lKexthjUp
m9CN/A8uRCQLw/HnE7oT44FLI4s9qNFU76E5zjeX/yuxMprvVD0EPkGao0fQAB85aDJxYDdCOnn5
Gs3aayykJs/4kB5UpezBcsFt9bWyQJ34sZhj3qqmOhnwUkbZDlOdf4IknVTuUPatt5hRKGxTDTV9
CZcd3DyIymg1qgNYbYhgjDqEbKWVFaP82qGyQE42MK/d2WtwcR/Y+jXT1JsvzBSl/XEjE8+9aoyf
6iCqa4FwJ3eL+bi4NSsrUW74y83xQBQEscrqI0uqu/4AcItrGV1eOJ96k5TRfYAvW1mZ7lxL/RVO
BUzFqT8S5WQgc5cjG40qWb6Wwc6QGGN9sl457mFT3z0f7rmbSGY93Sz69VGgtkY3OaaStvcbe4eb
GxQu8ul3ealoTN7+2nV4wKHU2CKrlh9q9fy59BazqXZGGHZBzXa685NwWSgRv+oQOcMgO6lA1Ia2
E4yhmmDdr0aIHaoad9pml6fZLEDsqGGCR8mj+OetJDn4IqcuHANA2lbsJcgLeyetsMEoeI6+nBrS
IBwviThQZhKPU0z3gB+yFM5KtMImtat6+WtrTfcqeGGGx9Q38BqW7BjZp63gT/8dTIcvnmBxU4N1
SwjBudbb8kon0y4Hd2+boNkV/t2T/YiRt30+YBNl5v/CsDkKYcDLysnuzAsfz5d+dsB2ReKCXAf2
U9aueKpZUn/RCbrXQcYlZub8SwlIqYujJO/5coPuTLJMVcZeJCeDLs0EM+zCmuYLSlepLilqQKhh
HDb12pg0YIPxalRm+iUw5LndrYQy+B81uXOvocEnDNceAvAaoPOsdwC0YtrqGRSqiB2s10NJikYD
Adc9rclu5R9DM8KRP2LdgMU1HcpBm3ScFgXo66gOQyn3XXYA2aYyED4b67l6OQ6iG6HoF5UKuxqk
sgqO1s8uyRI+oEl8lLQ98KuAHLZMGHkryNS+uOaqUIsfm1mCPyJG8tvIxqvGQEHo7H0lDY7r1omb
sxpC+TzyAyoVp9nECoUGGmSh37NuIIF3Bc8Sk8PZzqPb5VmXcTUVp6UJ4E3RNm30z65n4vEDoX/d
/7WjbxuZ+t4Nm9htx4rqL/6722rtQPTJEBS5Ito3SHybjxV4gzctOesQUcQCSFZ5b4b+f/6hj2zI
0do/5yWudfaEayYtBtV/Bry7lyPN4sHS76QqSeXxRjrb5Ss8CgariRtawjWx2ouAE2yCSM9e+s6J
aKdEdbBs0ImmY5/0HolMoLSvMYVU/DlgNyj28jphPKnrZ5f+MNpeyA5u6of5uH2HU8KcuwRMKkAY
viqqDqbAd/XLxVnGxCY9XefEZkt3NmCRyzVJVY0uWc4FcmI8c09SnLM+B4qeibEg3/flBGrSYvIX
2c96Cc6SCW3ixWNb0MS8vSU7lPWcm2s5c8YsjQTrM4NBtdQEwAMAEBswBGFFNn01BiwugKj0MIXf
jV1LCc3D9JPj04YXQpT7GiO1CZHEEzA9YsH4XvFx643QglE0CAC+TWmhc3Qc1cvfBnhg2q83ZY6B
A4jgRkJScJfj+OiLwB6p+NNBdg4K0fcl/xmskSY89xN/tyo9OR/wc3ne0AtpefqpDUFINHGBWF3Y
6bntjqQGIobbC+iJWxwr9Vc7J0BCyec6FJMqDEMVLQ5zx61Kq6ynGaiE+zKAFh+3FXZ9mdvNTU7I
zPrePynWh1taJ3c7Qs9rsqXKe6lEv34gHVdrRzRRQRoHa19oH/rM426a2GoXf2hIJ3/Sh/FKvA1f
+8MKZ8V1noa0yhEisiHjLOCDzRhEgFs5KdhuHhVBv2RmgGEdIqCS4ptRir68JRTKDSoTjHmZuXrz
klk/9/expDMJVtL747DkMHCSsqxDwsRkML7GAfeQKXP7MbajpxH4n06UJNP9NPFRQM9Bh6LPYJo/
75+j/lM93Y9tF+Sxrg2Hobx8OfO0zcDlNR4nPm7n+TH6hKBpSwhcjZcmCRdvt7aRev+JITjCHbmJ
VnTJb9wef8tFXui0I6CJ6dnXvQi9Bpk+kex845Y6ktSJ0WvWM2l3jhVzQms6p8hBTsKHMAGGx0Qd
OPuEXyLsd0CjP0EI9mROA9XPAZBVXk+hOb/Qb7k6oATFLwzmtNy9w9scTUJqn9Xfz4Y+H7prLaaI
HNpbIrWrmpxh7F75o4k4lKYl3FhtZAXouw+53nxaFzU0TKuLkf+EhHXDNm/HPorGY0CuFq/ztY6U
Vv5ElmUT0GFE93uZ8NfAnMW3j5OEN5XJSwDEp/yyLGHOjAodTVWbplLTThDlpVT4/v13ocmFhTsr
IZ/LLLkzzwOYEhG9+EMSeVmIB7gUj7m+SGwTP1Lae2Id79dpiikkV4r127TQKVZ20kFtKTIKrftR
ADQxGOfFBs1SOWQ+9ryU/8kWpxl/IVBW6ykPRdOr8H3FOKIHqGqJqJ+J9MCpv+T9Gq6ZeDelj53X
Zz76nAkxilK3nUxrvD4GlCv+SliSRENpXbTLgvdBP5jlCl7pFvkJbvFa02Ncn2z2hXojtY+VAwFE
yWgIo0Snu4YQzmDz8NtL6sfoMqzzSfQbv/tFqeArD/nRxktyq13p71n5jrmwVqtQ43lPsPUrSCyI
KpdnGfbr9L3+uqFYFRySFCQU5ZvhB3yGEmb1gcDyQKqoWSU4iCH0Y5/VRzMo/7YMzdqqUCrHMcCw
V+XYEBKvvML8LRSAOYBuXOlL0i4NFwQsjbfQYLhDUXcoDJWBKNBLxfMXhz2gzakEgvyHlva0bU1E
DpuWvpO5VbSY3fhn8jsNth1D2y7xCoTmbs0KEhJ+XUYmPsKf9+yZx0RmOYy8gI062dpGkDrZUIwS
kpvkwgW+2dexG1FKorDn6lMKxvWl9rlWg4p6uMOSl/cDETyXfaXGikPYI5yghM8wvAwQ2x8Q4Rx3
ET28aeKdNjxpXDQdscUGpyPHPvGE9dMNJEJYpnV6e+A8po2p1pH0b3+rvR+FzqkD91BlwBqnzV+N
v4TcjHkeTi0J7PFZ3Y7DeN/TmiQ+AhgyIB4ffY5WpaG5nQlIsOiE9++kl7/G1U+IgsB1l9VvpcKi
AgdiRyYphIbWWoDDspJLu06X/FqMF9TdQKQyZI5eS6bD46U/a/M+rN6GAa0ZI9Tj5odi2FlJ8Sdv
m3eg94U8Jupd5ZquXtI4VbQ/+Rd9o8ZCuSpBYWmUKvpwc3p8UV+pGnZXZ8DApbYJW2PhKL+31/qQ
cRDWdYdzvrbaimqXMCKJJJKWhvtG7NQAPxLo0eMXdlP2rrIpNbPOwqbChpUJ1bRYaDTCTryxy0hF
aEmByZOnI5r5e7aWZ8vZD+y2YUaLw1/I8Ubmc/ZQiJKrgx9zRL+4V3Xx+IIZFbIp6f/+aHO+hBvT
fVJLWPpL3eRaf280ufjryRTulXuJEFTcQR/2MyLf9yUEvRi++hP9B+8XsN6Oq9Y1208un/SvhXsg
MKdR05vuQ4+b0Bq4HNlKGuTocjvnIfDGShGRz2hblG6G2znE/AeIJZ+FUKhWIWqJeur9OOGL30Q+
DcgmVV7WfHLgxPsUdnabypinEXEq1kNlmAn+7g08K0GrjMJ+3BwvRlOVkY13M3cChnQuqVaNh1Yb
EXxDjPWlOFz+/W11W5IlmD0mhjddtBZFm4LRve9Nh7YwyEg/L+Nh9PTJdO5FNznNE3legADNllYX
kcVX+g+85UwfTxsuTdi64BWH/NYfF17Vzoj2bBnp8DDllsyodjNVgHcp73uUoqivVpVy7oLmkrp0
8DeSRzFbXhF4OM2EMclCBNcHpHI6z07yGqRO6zRNw8TVCOg+kJMcazx7O794SQpyTPiMe8kjWt7O
Y5ad+/BPeabnOySq1bXHixglMAwAqnrIMzqMrNV7BQw/3n0lncvZvmyl5/aVaQlXpTLYTLRFhGgu
o/PlBR6jpinTZr1Lylsk++Bb7HF+dRDz5fYecXf+y1TcanPWabKKoXdvQ8Ru/jFw79byKnxzFUfT
mbXlGMP7scGMYaRwYsSj+zTc8XciLSTV3tdg/EnILuBFryMbf6UKUF3Gsg+0CszUwAKsSGsAJqtt
JqZr6HQG7O6Pf9erOJVflJddxVu9wYC9i/h+uS/EBFS48AsOZd5xbiHskrCzzMKHoE9NhX/AJpvI
Y426i6fx2PEEjBJpAKlUjPp6X0ESlxDQAgFA1zdb2aRw9uv6+7W/TiJO8gef3VGYWwDoFrRcblFq
tTJx7qLMWzGqgc+oZsojPWaMGiWjb+vVINcimq6HHOr9YPp1f4c5da44CrdGEKwoZubrl3R3JpIP
mHbIg7yUVbfikeXZ+8gm/tlG+J5PUEigQjGkDBYzoYYhhVCjOnI2WN3sZ+4m4iSbQI8seQfjb9K9
wbmw++GNZpBEsDK3EGxtV/bbLDaf4wuOO41gNY//iQux+qWtQ7mFkWfDsu5/ty7jkWBBbvDNIoeH
XV7ze5BnbsO+pGhFki0ioi4L7AM5WF3+mQkjVeJ3aEfBDeq62o+y/dEn8XH+ptGAwobbx1yjBbe9
0axkPsDxupjZEVyPR33w7DqiEx6f634djBajIg3GYgIO5HZ8+ltsHJtCG6TZeS9TyCSf3ComVPmI
vwpIypb6f0sfsBjN/9GhMd8QbqUlVdzHUAIjw6issecVzAa1oMy3c1Max+kCnKDfgG2E5/p3Ed7S
1NpXLlOm7AZj+CF8P7TEMeFJbHqnr22bnmYGWJK89PsFlQ/d0OxjQc4+Tfb1GJt6JO8hYXExEEtl
EcVizcd7Dqz8i7D04rcoUPUu6gVr0VFpLy21vURLKIXxtmPBwbl1ImoZzrI2HZmKy5nV5Hge00bb
KVOYELgjOyAKkDAL2Ggx+Ss45S9X6F+E0kt5R81O2BnSnGF4TgFQ9pLJJFEF24tqqdPTDatzPZZP
oHJ2ZHjC9Z+yYn8ZZz2tv3QPEvyoWU+XUHzyHURG63kC7RUP7bBxaWhaa+Zc4btgbQMpr8ZJq2D7
bNqBMiBjh5c0LlbAHc9FlGTgBUh0AOJsAzJq8yEX5D8PvP4tqYqSW+xyPd/ycZPyir9g58jtLEU2
O0JDs/G2ZPqinl/aSOnmzBgZBjp+SNHM7QnGiRaFR7UHo5HtVrYLqdiO+UJbpbuOJPqJf0zMmb+N
WeBYu9IRQAuA0c1gDLxYVYoNaAgeNcKyna9bvco3s+8PvTtwHYqmry3JAQM6fj+ci0jZm0CpiPQJ
RHIDx0dzIOvWNGqX2gbX2ttejt9YJMN72lckC35Zg9LdaLfij7Rwozk+Q0nbYXHP1DNxtEJKEGc6
FGfFeyxWUEP9iyzNUVC16daiYBamaNibgIbl8xfraBpxBusfXSS48BcSyuCqz53c6R5QkNMhraRs
LC5HP6NDePocPX3lx76Tah2f96QU5/vB1MXcbLk+qQNspJXPNwGs8DDvGg+YyQ91E+Lkd/LElUOv
ijsQ4zHd8XHyBZ91x/xXGbugBIhSjCut4A5pk0D8EBf9hg8leeLIwDboWSsMfe26R7jzV7JiuHXU
pQNbKbBOET6bDtu5V7k6JqGN7e9OtZUCjTebzW3H/FocvF7wPpAJD7Uy0ZrKTzEjsHMsbcs+RyvZ
T+jeX5OxKbYylDo+ADigfnctuWQ+VTu0Rx/RlLEWFVANFkRhDG1pN4JxsxLDK0Efh8XQ6KXq6SU6
jcAwLm+ls4DPKOa/Q6KCs3Z8PCv4lM+sPEN0N+AGjEVSnGDNC8ZLXfqBuCr8i/aezW555BsMFz3i
LQLDTjnqqYWq+m6hs5uHhF2kabt8SmcC/LyYVqYPlaagvdVIP7or9clknl4uuzBqZM9/mCzP9w5S
KGzYKtOa67rabu5G7j8LQfNTHvsvvyIVlObu4Rp0QXmu5+e9RGw9Cv5FR2IRSaOMGHcGp47Yttny
+C8H8IDDfCC37IfSJHp83l3DfM5mvEAjnM3h4/j87W+D6ELcaPUrlaJMxolU9kl4MymKOSrWbrqA
DEJzxJ+Zrpz2z0Nf3r4lpYWOIcMVd97rP2MclLq8felH1HpRJo5i549OPF+p2knIjVbQNEGzK+Qa
e+47hlLj0jZ5vvbTQQsV7n4hYjcr83W53DZM0x7ctElp2P0C4PGoTrWhLaK4RQBXCZcpi8ncSs6D
NE/Jq4FZNtU14eNr9ME6zwmFMr0DQ7U0C9C6pK5iksucLfxWJ46GA5S7jwOIMrWkRiehF/j2P8I7
+3oS/hAhkQO+FRp4zVAfrHNOJ0J1MwQGP3MPwisWPBCGhE9TOqmHQcv04ArX0s9KTSz0gvh99HrJ
fIE9hOrTtErwQjokP5W05p30ftQFa4xgILhxodS5WgnCrOlcVn5Ayicvo/HTl04DGoTx9vIbcBNS
qDurlqolZnN+i0OXmJaqqyUuuLNY8hR7TPfG30r6WGwJg3RVutgSGZfI+BKJP52VujB1s1MoFEFg
NrBLuuy13UXBcAEASNlRK5ZIcZkN6lwBy3qHejRBu9vkCQGsvK3XHspTL3BcYidkCVMeRz2yqns1
XFxveWDapzviuAPRjVVB2Gu40V8EDEo1IlVamlgrCofbjFw+FTAubVIKqdLsDiA/qAf0HQasa8Pm
X+h8nHuq9dTANJna691nnjwmmhUIjefIS659UROjn6hlVd5x5vQZuUH/uLAevCTqsuopEIoh81qV
Scs9aOGC/vYgDzEE/kE7rRXNHNgKFhOK9090qc0sTzrNi1hr3I+EKfP2l3BwOoHSSH6dqmiZZe+D
DBh8xDWkOVPF4ie/1DBLvP/MdWXQn/8vlWE7ymiXnZeaLak7WUgr17YHLoR4Snmyc/WKkRzjZjeh
iwmsZ3DOtfwTcbsuA/WzF0CT8UosmzfFrDjU+fGMcc2lvHRMeAHAdaZUJIWTt/0KRtfFFHr2ySxl
Ik2tDKMc9WOz3dw0IAC6VnBorAgGI5xsMouCepcQaLFi2pr/D2kPjJ2wFuoIgYoyQoLL3hOCad4r
eSwfPrKPPhGazBmQn29hH3H+xwRmfmWTfwBSTPkreZWS2UetCBjpOvZckFzauNUoiC6ak0IyURni
nm8gfOeGSfsIeDzptrAnRl03YyFeLTkXyfbsrvLX4wr3fOslu4Sk8gLNIvZYS964Pd7U7eaaRHCL
z6s5S6s/ZhR7dCIQo7fnXJCh8v6Nmm8OtCpX7u/g8Y5SpwOPc23rTNlfu5+a1/uJ6pp+mrsWpnDD
flOvWd32gXIKmofDgzk05x0m9WB/wkm+J/ck9C6IuNRasjG7HPco0ePYJhIRmT9GhS+zXLizqKkp
SnxoyOBALN/DF8u84t+0g/M2sboH37RpViJ2ktZOdErOdboMI1AILJiIj7pLih4iu0f/hPMcllkZ
PPNrNT4/7ot2lMCigQeQ4+h/CJDGaM2E6xx12oIuqIFVsWRa0Y090MpzH0NSFv5+8xZ1i7cwe4b8
sISVNqJpkGpKsr3LXQL5ZSYKrQB5mUEdeM1YUorBSxl1qCWcmblu/PbcLZKO/cu22khMjviVpr6z
i94RApEH8wgzKn0Nj+o1K/Qh8opb79HuWBNSmMzOoREb3oTcWZdyG9i1OtX0aAVxI/t9ia8iaX4Q
Zm2wjtGun+2G8oR0MDWPYaxPr+xjEGgIVHX3TqbU4IqQ458w93tyswwmp+B3L8z3J2MWhmswye1r
po0hqnfcjZJ4RZiHRw4yw+4DpFuvEGR48tklVPRLpwjjc1gTciSGXYjULUxdx1vYAQiW8cj5BIg9
pARyqumPwdgJHqY9sTJCNtS2ibjm0VmeZEhpMtdm4sXQLEWGZ3J9Cl6aSB/1aGdS7aqKpc8Hvh/8
ZlvVes2rj6rEaMWUJgLre2iFBkcWlOBwFpscwhSv165//d85NU53VAVTm9yydPgSNOfvi1ZRBB/x
qXfasPWntsrgXcctEQZjjoDrc00V+T3yY7f7IQ4rCzl21Q53t4FCoxtlYwX5xI5jSeskruTtO+x1
NpJC8qAaTuyiade3z/OIg/JjPQ6hni+e0DcHZjsFX1OUDB7DNJGoOaGNwBdXz6lFANoF6q91c/E4
xc2Oqj+u4i2y09gT8vKJ/qU9ztyMAaDv3lL4k0l0iO5oAsT2SonhZCJdUkAScjDroCrXmDLXXjXJ
jg7hMX7MHjzgKN/JkUYqeE+W4dM2cUnsgzs+EqkwLZnGzr2LMVM5h5U8A8cNCpbwfNU5hJtgoHYB
5ieLyy7yLjoyOn6JCaCcuswqEI/vN6hyePKrmuURkJD6XMHzH49uTks1rhclCUHQk+1l1tIzxXXk
neInIxmjBxzgloXCnIq80vjSQyhvMlh+5NAOUygDKBB1Sb7zvODqe1AQEOnFiRVtROI4xdv+kv7k
7CTI5Hisbcl3gTq/BXZKMn4aZTyrYX7tgLkP6s+7M0BGa9tJqbR6PtAO6Q66iivLaTLLUheofJXj
MpbC8qPJxLt34Z9mZivCS60guLbpjgcsDa/+yURsrTpQDcQNnPHO3Ibb2pdaqOvO6z3AlelM5q7O
UgPjaBCUzWdq0MVe1wF7GLEfrzheXHGcUN7mH5cRlBjWHZxSFLGg29Fg6YS76Q6OwyBd27xvP9Ag
H5umzfZbTE6wiCzJCqaVHKZmtmyLJce2AvULuId7Lp/939VuiBygDk+9wq+fOSYhCf376M2e13Ua
2KZ9IwxxnfUpUT+3hXLnNGr7tAk5iccREZMe3btKtNQN0zpVZDO8HtNKyOd7ARve2weCWpn3LEjr
peEqu90w+A+JR0DJhWEiBUZ5QT/UkKfS8MS6I/oSrBipmgWcMQODoqVOQROQcQQuFczvCdL9Apps
eguZYUWMvUiYu1QID/pq0O+ycYcMDJUZfKzMyS98jWs8NUMIwpau/8Uonzvk+qWA53MYMSBPKF7/
CZq0Xbzxomh6p3xvmQ6TNpTGnt1jbMJGkro5JngJ+pTt8zT1py7BQ/dKaR8+/ukd5k8kRrsdurZn
/mBG+hVF2Ow/gIdsPdvYRwRsrp4Opv2ltvzDhT6Zp/3tLm3WlFO/5R7K5BBlHqerDT6BA8PCeUba
ax7Viuc+pZ7XR67uacukW8wVXiXygiE1PnaDPVUapXsddUVmZ5NQSplSEXUrjHKEP1BTUq0wF1yY
RaXm9IPIrEPzB0ROoZs7erc0o5XfSn88H9GZEeGP71PHjAx2TSjMrHxXS7iKssfWPYtxT2sGhOm9
Goc62WNyIvES+Sck14TT+bjCYzcZ6FLcCFL+fpr5ViIdBX7jdVm0Lf3mW3PQHbZy+sZU4ZLYkRjs
Ss4iGqUUyglJrdCEc+QQibGjYRicWPW7uMtVqLultQ/zHTfePer9mVmymDhQqTSNJgiVHMHdSSov
Q1uKA1djYPY3wUOqfVDjn5kRusXQFbfhwr4Xzm+37BMMB7hSDi2efiYazMaJe5avJ3SPd3AgCaIj
pNWesOTYllUUVFhYQI/QWaZWtZe0SCHTlpv+mcm3OiKP6ZjlvgLOSmHfwl1kTZlRCaVxD6JCEt8P
MYjT5YiVO3l2gcH9z09bBNexoV2YQwR8NDMHY3OgGSRo+NdzrBp/anc4o9QKUEygNnLXY0ly55U3
K62HAF8SxKJSyy5o/nfzB3PQK9pbDunwb58XSTAqIxLkX6L/IfaTU+Wx5Efr6dKgXnksXkXOoQlC
xVNo13OxnNb01lsajIKDXfmy/SWFNoc/qsBdyXCtxYFpQoxffZqh62ZY8hVodvJHAJOXlfUv8D+A
+dCBjptMEQdbZSOBkMyMlWtphNU4aYgDvA8WcWfwudtPtckIsMrpN6kvH34dHy8Hbwd3eVkyKiAZ
86U7W52vy3ZTeAS96qV05kjGl+NYmeAhLPrq1wQ3llTx01a6EcG+YDE9UJBRJ1Z6ULRZA8m+ZADg
ATabMDZhUb/8eFyeMnsfYxNQhcrj1uEyl0uK/c89GKuP8rVJgsNDUIbtnkFxQSjW9a4l5ZLoQ+qB
LFEPKuf/nfjFKrfqpq877ZyDcvEZopFOJjIwgJzJ3VVfbiSOOPV4yezwclGwP+Xywa+U1rZ/YiBh
HzIMDmJ3PLlUkN83Y4iss5iNsSoz7vVr88fiLs1ZBF+eTAQ6qWD5bcSo5/rcI4kczEc73klQN9oL
qmcCBdPHSfTy7JjQdXPfwFbwXLg+TxWFAqTO8r303lIuBbrnmtxsdL/oFOG8tHv8/pdYtkXjxhLS
fClUtpvixH8MYCv6R+hEE6sPUn+uE12LkLvEUgVdcMHqiB43DCT9lMULYXx/W+dD2cGa3C/uf7YU
SqiTdZNwut4hsmp6LjLWDqPQfpbsLAiQGhHU5b9Q4C6RHxt2adfca20v8rPPwWlyzfVBCJAA7o2t
Hjt7lPImJVA3Q9USjkOvBtJu210ArdQmajkxjnPXRfC0+s0S3YHSWxZsvXyl37j2Q+hlyRvZQTeX
GAvnozfIBFFLDt8BmUGv8H51ArAOCDAwOuMdySjArHTy4OFgUZ/YY5wxMZM3L6uj8T8Y9awB3/Hi
uzyfhDHkf1Ep3VGq3+KTW/vBXkQkxiPcpdjjcRRJaobvcfLuhKRC+HREN3eHKTF/4tSOxSAoTfRz
X19pGOUYgkCvQxNw05fRC1Jf4qRqsvS1M8TZzjeQrl0ccuAqodZQdhgGp3IoK7adBNYGq1ilgQKz
25qquAw7qrvTJjRAwiH4Ob9Sy15HCxPcWDL1AM0t3Cx46g40DlL3k1udf2xgYZC54KR0xwjfxJ0K
B/4OlQfcluz28i/FzW7TX3qsdFbuAas9fqSsYI56kTYkTNN7FkC5G2v71bUgjOOTZVJIBEQ3BjKQ
Sp41rxTrWXRypXDn6GRY0RGLUfcfmpt87MSOeLig1Kqer/Nod9rRCwyC13Sr6bMyl1MsgrkUBuYS
9wsiCykeIt1/OrMWbt/dXudLPGx/73qmqFkGnUwVDPvKsIAzC44eO+jNZPsQ22MoCKQrnDNWzwtt
/A+tzn4B9MISW2egLOUy/ks5CEwXSWYYbZVsftFb4aihNGBBr+lSUVD9kRcXXLlR+0ukvfNnH9WV
wYvs1UGHNGAnYGlpMTQcylsFrM4xML71/kdvtqZsniBMwNOgvBnLXLdYFOX2JT0a3nESHPwRXmc3
xXazEWqBBpgSGKl6ozu+eBIQoBOqpQ860ZWKmOQ5EtFbysLOqDClXfbAosviwuqQl+c74ff5SLhf
fUeA3oaDgV4UXZmC/R/Qst8NYjXoSMr3Ii3/lFI4XTdtu1AWxmhjTebMFpt9NPb/3Cd5kOtVNcB9
fQ9fU04DrsUtMYxuR8Qa6s//yN/WnlZAJ01pwXRYnFh83GqL/Q39tEwNxOy/jmLisPmT7NpJYnIC
KUnz5MASMqRDcvB8e7gulavQk+M57tEAlWSGSuMpBl7bs348N77FtLieKefbpZYp+UY4eYQa+GrQ
dGeB68LD1Tf+3mJ/h6BzlBXLwdEiM83pcQoto6BUIM1Nh/ss2MbA6dsjTA4Fuhg5zZg9Vzz3SZC/
AOGs0T1OBVH7dA/9We5xWID+BkH5hwpOPUMRTMFUFnx9LslXPq58pgIicp+sHy77WAjj+6v8urAO
7adfesjyo9slPyTgKnM5MNgOL63fhru0PggEVr6aZR4cuZrPlPTI81SXSadFpO2gUUf86f2acYgo
hxGY4ZXFEHaRwfT+o8r+ra2jZi3z4IQTxNsJ3z37ZIUKuNmbFimbANa1msNA9YPHEmd1F65wpVFq
zvwEhe4+/vSweS1n6qnKj2sGA0yS0uV7fFd527qOZTDBETe/jXiSXl/mfS9aj19yKrdlwb85+0g1
lucj/Gg0BA6P2sd095SdrKHOJaic5TLcnfodfRu02FZs01UwjROh2fqv8GiAzudOyhNqa45itX58
9kkjNPIk6cKeLJn/s710GHjbD2ARs33Z3vaO5gZ/0qyFeuoEqHa88NkTlxOJaGieygtWRusFTFl/
Qm2SfuJIEUER7LEAWNCUrSY4LlfUu+8ExGxVi18+YbEmZFUxHKWulk79qyVBvfXWJePLk0A9vUnX
2V6i1r2uQmj+3IH/8mfk3LsEWbRyPwy8APOl6nB8sfyN44zO3XIX5pR8u5Ttyutx/ppYvLJYgkp2
h8rRx4Mh0pZsYFUGQq9e4Ty96R56wCSYkLlWgXvA6ECChLPq45ct0lpCHBntBOK6bBXw8ntVT5ib
J4OCdr0AlkJZ5PwUIj3sP45PP89pFpvvnYoXRgeZkh0reMV8F5//3OWdQWOIlj+y1Z+6pw8Vd46E
HwZXaKG+5/75GOKT/4n14IgEqK5AIrLXz0GW01xv924bmF/+Cw5TFP5nt395TIDJC6yBGUv3i8SJ
D276OIwMLeP7IR00Wztxi9KCHCdv/7V/lPycbxW0OuLLcjwXDuXLZVrsV0T5yNdCXqAM181C2vMT
PrZMzEytOyo/z2GYrlO/5E+sJec8kVSS8JV/QfjpgF0BbkwcM5DJb3gi5RW+XjHRYG3tK9mP3B0M
sRd95EYY2zCoCeIjxhzY9us2VBImhLjR3BPHKWZwuNbwTlnLllMiNNhDKgxYfIiPblnZ2E353Yef
Ek6FfmlDA6P+sPdnXwewWi0selq25MxUFbi5v1pLhbAY/APtesmqaTf04bmerdxajduUcum7MyP3
5A5e/c+6/ggXStIM9e/EeL4AQhvWFWFOrr+3DAY1/hGQVmsLrxpmGOAeFBeZ+ZcOh0LQNSSv0WJr
GoCL8CYCCzkqiXVmnJKkJOSHjikIqJQ8vDlozgaRpK5TvNxVvmZdSHXZ/Z4cFdqDrUUZ/ur8ngLO
4tXPwpZwyqQNxRo+LR6Dgq9U7OoBzkRPQ8F/3bYXWud8UPpTrswiMGAGft05wpDkC2shiG7KYpSe
OPoF3yf7GgGAsRyt5YzQ8exK/dRNfIYixWVftgbZ864qL+Mn7Nl+XfkZVhMVstkwnzjBxcWZjIqI
JTQ2IDxAnTf8/nNigBJQfNN2NBT7I0siqctf8MV6Ao9aAzYLtnteXDtebF6FBQcVBGIfWBbVXiuS
28LqzUB+YlOE+D3VQbUA6IQ1C907RFHsnBAsB5bMRBtTWdbIKBwGjia6uHvW31sFUda8AlPfyDLE
8Z0T/vlcb9p1y6s0SwUuZ3rqZdk+7FYp4+PF8Mcn3AiSLiZZb7dnrh+gh5k7f1pmgKCjmQ/vAwSZ
UCxEtxal8vwgnUEaRniH2UC5H0fYGO9WX8vA6C70b6o/dVD7YJVdpIZJgh8qdaig6j1rYXu4PoEE
KqJgKMQG0dbhnpcRIXtrnBJhnLOm5VCSa2qGkYFaJbHLTcvBp6GKnyznxqGtiZ10AFLEZR1r2o6t
i4z2p0UUf6FeEFjPauPQxjP4mrr9dSxoTHsQXj4mvs3nU6uFesDjF+tmDzwDma0wO1K3+W3n1Zwi
RmD0N+ybsjciL0fWNXzu+dw4SvpU6pxq7wT1O9UsTH3TxutCtGnobK8rJ6c43WQb7yD3fHf51woF
7ZVK1ht2ztg2jloNDp1IAQOiV4NRXT1TW6JBWuxl+B4bgzQhnkQik5YuS4F1XlN2igu6Tz3OS1dF
5BwPXaaQoxZRSQXrC0wrp5MCDTO8LsKyqIMBgbMHpQ06QJqBXn8j0YODc9WKxLSmUs9oAP2ov57Z
Ysh7YtUwkraL1+YnSwr7I46wCRHWT12yOuJ5iDbueBwhe0Lak85TP4TxUQZLdBRZe/Y7ki+jhfWt
TvEpV5lG/Nqfk8ux4O8wGMDtIvBXv/reJWmDe6W00FdlIYD/qJwjpxxeU/UyGPHtMT84M4WsEv2F
iSOdhkmo/41U5U67erE5vcrgyTnN7xRxm2ThgIG6dxXExNurR0CIqAyi5IW+BCWFH6B4PB7Ii+EV
MS+9jZKGlMHYN2Mxua/Bw7paUqw98fcAEJ9aEdC17m9DkBVo2qbZAjKqvH4Y5fqiiFH2Tousm794
yJdv1fOny4lZz0XE6zx6ZEt7VpmpNG1VM6J1ClCHfvnIHuUMPs8itfFnAxqvexwd5aMHQT7bG6oB
+dABMN36uHfLUraSLjTuHvJECE3HU4r1gOKgQbqDaYFyAxKgCfJAGvLc4L06XLCH9uQ7WupIXVZn
Yc098/PsHQXvAUZqqXNfK7jO9BJAxmXXyv4aKBXD2VQGMVLnQahB5qQi/LaBxrDhe1BLuMPrmi9C
5/U7SUFrdsEBjfrt4/7emplOBR+DKbjycJFIHh2RKu4v85gEgbMaNTZnRYWlbOTYmat36uWwqkAF
ArAO+xuq/1CIdj4rXwLYgZYc5JUIdHUN7qsGzotVq62ZH+7RF54aVPxMzogB8lgRJbU8uYcfOQQd
Y2ztKE9RsBWEKN1HMuMZ82JGogcEANjFrPeSFz2jSSlKeRji85y/BUGiZUlzIRSgcIGhOcQsKFHp
qrkdng02hcABaI9ccGFRW7IysG6kouAo3eo6UnP2lc5os/Our4J1qtISJUk4yqNZI12JPEAcZvVr
dhwUSBROR+wCs1ewsubpmjmntH3Q4reJCojs6DhnbtaOrtPQOFO4RgxXK3cCLRFHpiueYROmap2D
yLdEEO9ysQSOHUCKmK+pxaY9rU6l/iKdeFn2oJe98ctmdO98hSOsUH7EtCZSMQLSYvQXAOejMnSD
PjYqdjkkp1WsYvzHqtzyDj3B0q7Cwf5+jLJRfJ5fOyKrYbcDh2b/SidqoQqM7l0R+pZM7srkzhYC
9lGlb5GVL3YL/9J+FxmUV476q711AKOngELGD7ZrVJVaD/yj+2RuJm2nzEeiDG1gPSPqYRUFmA4Y
o3fAW4jqsJ9ljS/m5GCyXf5QIF/7DM+/omkUYQbmaPAKvay2+Yxr7zZF9Dt1S1o2suKHKqGk3YSy
7WotcfoirQikPwZTyQmd/d1pUaGSgQxgS16CIKdseXLIT/cEdVhgrgyfThkeUFiXlN3A11nT+u57
o1o8yuEKPNOCzGzwomG+drYqF1+Udyknnclrd88i6flz9x4hUBcDJtAQ0O4CloNH/ibgbSDFJXDf
Y2MVv6lGPW7COLWiaQn86/uTVfUyu4o0b1IzA02RlIaaew7uw/dMsVTIcJd6VhoFyUnheB8MeKxV
O4729/9PC1tfwOU3C4JCYKlyWsza24za2q6UeqSVI/4I1+N5tJlqOrqCK/IY2MWoyYBkNyRSAjgs
TAo6XQ84yrYq+9MyugHxwByk+WgFCodVtaIa8gzRFg4Opdbgb5hGIPRpYbPzhb3oajd6iR0IlqX0
qpH1jDNGgXlAzS2dE2C8diG+0qk44eaj87p92vQNz68dMn4h9SF4+iOfuHP+Mf7EbqGEX8L4zLhs
a6EOud6yiLadUinNkVSVFNWw1k/wpzg2kCYLk3tkTos/A/SnpuFVYrYMcL+YjzD3qayDnwPd15+c
PizcKm5uBR9jrQDnERX24SQcnWaq0N0dxmtI6n0u5LyTGqbFo0wY93BSJLjmayRYSGNHIUkkVowj
dyIP6MnhjTiKZdM3OEeba0z/l99aJeAzHbfLh2DmxcNuri9UQc0ZNgYIHqqZ8s83cTxqnEUm2oYY
vdH495yl6y2PKEtJ4MRTCBdGXPa7kyPWV1jq/YSoHpA1q71ZvQfDwL0g+05AZdz2eyAU/n3eQKJ8
rIrKLj9Nh86+v6YjMjQtZhUo/OosTLsiraLM9rWQSYWbJf54c0xzc5WqDngmyctHC4h+SrB9lvdi
X8poh6mELrBrznzYMY9QewXRidgvMf/mIRVX9nV18wa9rz25DwVkOu2n5NhpmmVxYhpEj4ZveJfD
OnJ+aEMf2zvnDTvDHHYY0ww1VT9/fXq1j/VAD04Ndu7rK0tYntkCdq3D/pQN65Nl3EuqSFgU2PLu
xrtwUAszcpXgTgZmjxjI4QOPvSFLroUl6BpvSfoGbmZVKD1t/SJ2T8fIHn0ZHRbcPVpAcQrN1/J9
xvsK8vkNH6SnX1muf0CGbJV8RlrZS0DHYwD4j93+eDcNeLLQr7VLqWmE2g9elhKCgMspon9zlqHQ
kGaQUuF3bq1hu/NNRATCC02TdEJhds/DWmjjCsw2oihhbVlL/EYHnsrgMW1jXPEn4gn3Hwx/SckI
u/lwm/j0jUstURT5QjBJhCgmaxV4nmxG2Nb6u4aPBmepaM1rcuFEagte/DuBNC3sV2KChNi843ET
nxeqUVeGVBNksEpuo1RaKxEYrrRKRGK6ersmOlkUAB/KZJV2zkK0TZqYPUpt9Li+dwxUGcZyUXnc
O+/36j/OM2pjYqopi/2Mv9zUw6hV9koBOrH8EtpEJblx5Y7KMS8A8sXnbD40jrk4sJJ+mIGC690G
wZixpACVtz5ITKtKSRAE3xxwVt61+6P9N0ajiJMsa7pdW3M/UW9CkaDiHOp2U5t8o8xtIfxrWEbp
0wAIt+UnJMSoZsa5kL3l8ZVYjnb7Jw71EdowIx5vfIQR2uX8tSd6ICbO3PXHLCboyrZ24yaAgm2o
piDx5pO1olVOe8LVPBMPAhWC2n2NifNTPAtYBZv/pwq7IjdtE3T8rBJEuPd9mR8IR/RwUHGduOIH
e7TY+FX36v81iTKvYn6sDh6qZO7o6WiQdm7gRD/pkLGPjUoPSbX8gzhvSrp+fgLYWggmzE2gHx2m
za811/X2sTtvmPEQhiSqArBeBu43LWRLkD7kk5O9yTaLe5dfI7W/lNEjjPwF+F7c/Vz+lzzTlogR
z+lqm9LmJmiGstzMwLdrh0Si1WVSc4GZMH7x/fiyEvHC72POTKpx8Pn0TFAPrZTjLfCwZHILWwq6
oiwiVAMTqRuzzhTjPzCGpQBToNS0PFev03Ozc09VZp3mywbOMGrPQ2CainRQB5TvQRuURgpLRDpq
my4xwc9CsX6DoNnbAbfKjafjKXfSTwqs2eaBiT+Wj0M5L8SgBLEbq7V6+3q+6JJ0oJtW/OxD6tcB
p8Zz/ZrU46Ki8on5bdWaA6SgpnR6LYfeqa4f0uFmSREd25GnalV9kWMju8jjxjctaomb/aKSH8H/
lsLpaMQbZzm96dVKyxzFlQfBYO0haj4t/f9aGx7LaCHE84YPuMuSPzqpHYA2oqsR8bHllpREXdAq
GAXqqiDI+8UPGz4iWdH74N5FBDbaPSgZCtZC6WCMmAdyorI51+wjvrm7HZM35MsfuYC1U9g+ncr2
EvPs3gJRUn93TJqjlTBi2hKqDvwKZX4kh4830ToMzwJTOpyWkB54ZV38uvvymUGXqKGGNBfnqsby
7wBOXWtNsSsuJlMLb2DFA9s2d6uK9vHdsGFCzSNKuGBH+u4DGa3svycjosu1RIS55qmctAT9MU9B
2H9vfdvtIpGKeGhdve3y1VLeK0dbxX2Du0vBu3gDlBqYmqKry0r7DvyBafqHWiTljEsf/Zh2Uw5j
GH/pQkhZaT6LXz7bNWK89x9Hikf3tJTLI7c+VaL2WnD+dOrY88TKrCFl5Iw2thtVjNbYkihcmVAw
39pkIU95f/hpXf0EWCB6aAo6xw/6d4id/a470LcIjlPy0ns7zv0sdL2E9eksSREHy5DqBAIAXQl6
F25RsQ5hjTPBcOVyv6+DsETEIoTqvLvR7DJbqFPgh4AG7uXH5nclSf1dm7egiG1eCp/lIhdEqUVG
v9Gym5xIwRlhk3li+jcXp5+Sy+isKs17NudwjxrWRzbD6xc6WYRvZLbFxxdTcgAKmLh2yZt4VLVJ
/OVmw88k3imtsEmmO1e35UmHF20yFvDGyVzncT1xzNL/HhisqQznfY6twuizosjNqgcVWLBoK9YP
+VBKw2+LwJvEnMS96CVAYujBmfOx7LZAh4XQ6ZI9VPqhl6hJ0XkY1tlY+YHf9rbPRKEHnkwnSr6R
xssgEI2QzUbxFBUciD3vBJW5S3cquQw0Zwz/exLBfWF5RMULAAs7Q2fLc/pUMMBVwLZ7CJYQRu6p
tkqMq8A/0KYuSytECfO0EZvuctZmMn7AXxl0ZEAt2OiEMCEfGwUdQX8mLvsm4ueMpocIsxM2OeoP
1J0asotyCMXQF0q8bGocpuXdGq7hDzMqFZFcPjDvMjOFpq2a4HJdyZCVCknq4p4EJgKCRpG8av7u
eE9Gl/sOk0kQbfBfzmZrUJPcCJIsaao4F4qawtK7RaGRTBsgm5MKU8Xg9tTc9PnjOEwLaHQzxibe
qKtiBPnjRFTiyCM8uIb7EgJKFbgWq6NvYANcluWJiErXxWuuupf5wX/hrYMYtF7+bDSz2FAgrFBQ
zlcVjhp+ntRXp3RXVdVM9QuWIsqmGPRJzC6dZEvKlDPPLwmauYATNBF9rOE5EEU+NzJMwpJ5wGZz
uK9DeJ5BT6Dy76LgJR/igp6HfeSbSNCjJsHgCcQ0kT+22hxkHPtNm+tRTh5+iYGfdGnPYKYW+MCl
lmL+Pm7KYc96RG/Tl6b+TPBOqpLLLt0ojBq2nsveggnbHLjUw4B68ttqTXoom38WQY2+O40KD4U0
l/B4NZ44AnEqK0RKDD0/Yn4WPWYSDatme2UNV3BbNHWsZWDL5/OV415JHfpsMJ5fauubZsSXw6OV
gdyI8OenLaJjMiFfObET4ATGVpzTJy0jYSJnEbyKY+UKcDOfIxml30bsIo3/XEefO5+gjHep7Mev
UxrFRe76xfjOXmGsxnk8Q7w8evpNFM+aSR7AZPKq4oCJy3UtJhATpPyndZ88ujBxocjJ1qvu5J2D
OUfxK0MMWsqd/zjhbH9uUl4jDcHVSlkrKYitJLhdfWvFbh3atpetSd4XV6Ui2skqFqj9gAMSLOmg
vpJGV6FtJt7q6tATFUpdwdxJ08toJ+pHLIoqHlf+JuFt9F0rdECIQEmE1g6lMBiCfag3w9GTwitl
0Iw+shLWFztmzTjvaNxyhVpFUBDOlWIGRMnbQIbjNCQS/Dj0Z+dYaLya9tSzwNfxxdHT94f4dB7M
xllm1ROiaHw1fS3GCHrVeABJhr4Am1j42nDnZXBSrgrCAD0AX4iXNynSQja+ot90hJwcXtf3Jxd4
Io/R2dK7iIR2Dc3u0ptdhkwggqr+YjAl6Uf8g68NCMcqT++cGjIBFzMKsZNHMuWTceZ/v7aaZsW/
oLlq+QSA827WIxbi88zW7fEgr+Or5GZezxSRgeJh4wfKDKG0VLyEtkYVMRjbmK3nV7i098hwexw7
260mdmX01kD6CwM/dKeda6W5l0kMUozyL8sHMZhvNThVJDBVYXTacfa1MsvEIQPBShijT+Crax2Q
dy0z/lF0jCCYEEEY7NJlGbSdjkA5WuerwcFl7DIKjAQJlbFfXrY+HvMIHTSXDXF21H+C//ZsZq01
++DOB1kdIFx6tPp0jDMaeoaQa9KaNvB1A0VBL/nNJ1Bs5gys1ME4u+AgQ1dtY6RK3sMpapWbt3ce
NzQSGCea17GcUgmnbqhMA3jBH1Sf1zJrWWHPEDEKiNrgys6D9lF22QhpaMeD6fk3KwJXQ4Fk95WG
89LB4JSkCcxtFtKKmWSSdef9SwywDArGGiDHJjFt9VXMy7h/HNwCMJvdKRyX51UfWvp2fK171i56
yBX7UTtZRRqNkAXiMohsLN2ci/5IMzmPRtRXGM4SYa5xRDf0IXUKkUE2zGMY/1AI4zE4XTiE82EA
lruu6O/amIE/skAjXeBp+f01Z6tcciscl/ugd+SWCZbvL9j9g1XknEkUval+2KKnP5oA3JvzWmTr
uj6OFWNtwd6p4aFgf4RqFF17aScKw1DXgVVoABBzsBWMyKUQ8VERGQSan8JVDf1FSXkNfWjmE0eD
n+vx3PGYG8LkIjIt1Tlfjs+135De/KC9IB0c+9OkgPcNatcwoKiVfsPS4rETmRDPWgriGN9f8A5D
0g32YRsF2zE1EKltm4FR/OG2+j+NlpLPgUA0qH82YIrtoaGn//PrxNIdgA69o0s3nKOX595fuoFo
xJ7tL/D3cHwKZIaYXdVxrklZOFwcPmApzOr+L6Mu/KHeTDJDwYeT39rAqlCDXf2OgNy+QYC2fBQk
uXaZW22uSE09HDJmf4hOHgPWoWmb8yrv3ps4Bz0IlSlVzbFr3vsuoMNOiPbhnVDhZC1Fv0zENI2U
3qRyQ++8o5w8kZ5x5RNCdLHplnx8d9ThJBiCCxLwHvFV7lhB3DZzT2i1HOQeJfSK7cE1qUcoAE+L
NVJV4S0K1KwJc7RfsJnSwx/0o7OfMDJZDiKE2pEOWUQDf5xaGCQDl9NUoinDJy13DbRuoh2QwaFA
Ykul2iwPDs6QevFa5QyC9vQjBQbh7SSwEbDrKozN14/1e+paz3ImgqmD6IeYCotD98aqIm5jfyBF
5P/ESjinZ2gPpUOhsgq4QyTJgZLJ6sbkefWL13YKXQt3zVH60nq6u55oq2Nh3zQvi/UgzFO0pvf0
qG1CR2HbzU3eyqWExBTbhswSD19E3YCkaCkTl70QdOx2QyFDBBspHaWeoGbGH2oO5GwJlLMzugfk
dUCAbo1FF8LfL6JZ9VSrrIbA90lP3cz+jgvDePEIp19SWBc02shRFRVxJ8dvTeUMixtW01fpAN8v
N38iywPP+fjhESUq1lU43ta/kCuC2VuXhhsA+s5kuyaW8xLdm+EG+HPQcaaH01vIRt3wdx3NRqH6
UbQZKFqjKM78m+USxcrANL+tXu7mrW6Ocqo8Ikmn4O4Hz8mtir/Qk+DDwclvpOSd31zxCvFbDjdj
Gv2SSHDW3IJnAWJnW5y7zwROItK5cGTiTP+eiVPzjJhr6+ZA1Eviv0VAtqiylTNsJ+kKS+aYuPfa
KytvOTCoIKu4X/M63kJ54bCTSGexMMbyOA2MdxffkBrHiCVQxvvwyaDbJUmx3ZZA8r+eLRndsv1C
2JjZjuRNl4xEFyISTwyKZBi/qPTzoWajiknQ6sP5eueObjZ0V4tnpEXTJ1Gtpur0VkQgI8/Da/fZ
xzxu07ttSWJssYwBKGqG79ojPcT9bbeZBokMpAa/pfYYv83YIuMzE+moyjCwFbRJdOsPavashyCT
o3rU+f8ZvO08k/7AcNRBoQd967unmSavGPj9pCcTiSmJbmNbAxesk6eFZ+OUn1eSi8E1jtAoUAPT
QWFU+ZH4knaoU1+SYrg7DWuQaVPPJa1QFwvBnCbqk14jR+SSpg4ZWW03BEdmvNmk1hRsFQdyDc7f
UcdGDe2hABW0Obkm5R9KSd1l5ZwtMaiv1lL41z3DygJWY81mwMUzOufaQ7v4gA0I3i5Za/z5xdrm
iCLLYdOCsVFKWTvqu95Vsq0B84RmC66WeiuNqqGlchzjyIV31C+bw5GWy0z/w1rpO3LQ8n7AkOcz
ictTC12b7vK1RtbcJ2crXfvTgMEJKy7O4z72Fp2vefd7zoZIFkdkDPSLmwCmFyBhPPESmBZXC0e5
rdvq+ezF8soMKzvLHMEojjQJDivGz5nJJ1f/rn5iSLPgmce1zFF2gkxrZDH7UeiI1X+Tg/9rcMgn
l6IWyQvvPUhnHfHh+iHg7PVFASyK7qlAUWhb1/IN09SKzjwh/oTlITVvRA/hi33Tgy4yvsg1akdo
K7dE79GYo/y8MN+bvFKp5cfdIgdu8Mp+5IzF5TEF1S3Z/2QSv0QYDgAh5XxGyIa8qK1kTR/RDlTf
L4mjYLRj+YD2Q0S5A6Bmvy4PFOYy9/LVqQDYBpBYbk4xv9i4a+O1fCT5CMukiL8RmhglbxiPpl/U
2vfWM4OtIxRooZM+EDHkxfEGexr/pg6BMqkAPpwyJufFALNfA12Wq9kZDINuVgF68MusmnDnehil
H5AhtLkPihgjCViTJtHiQ7Cf4w0dGUQ9SIqxEvjrpy4J9R7tfk2AeGLryEdYL9otX60dMaDS/TpM
n39zXw0zzErrHxXGRlA00aXweGrGjUXGGCAb42ZHZf1o2r5dLAiGdpcerNXjEDCcPCqUVL6sYUBy
Om3060VcsbKv5Tc0MLMtHzlRpjQBz4nx4JJ9ldoMMam1S0Um1E+eygC1xlfH1k39Kxlc/6Udq/1d
HYqEem4Sjod86LZgCFyfL4jOj7VOBEtVzkcsqydtp7hHQ5oz0XmH54LrrkMnlp+IDZwBmCpmc3UM
S/7IgzKWPQNLGjiAlzVJ7nyC7k/P4GH+5tmm07RUhKO+vT/4HTckRqkL7wqKXWsusI9e5l6KTx2E
eDx7AFRqsQfvvYZa1/AhWepfbPz3yHHViRwhvPNx6GfoZux+jBGLmf7lubGRgGI5OdUSMuhxg7dE
MUcETmHSyoZjYZiphgkUk1Sa9X6JDoabCGfVRnJuTB+RnDDdEzskLJfuoxpJjPbVH9QexLwRAZo0
RgzeEBE27+txm8ryAhjxyq+Z8T62/uZqSkMUgQd1rf/wpYtFwubw1pjl5fEVYEUcU53rZifKibjt
p2iIdQeqX5bABJ7sfZv6K+Gh4H5CskI8tHhdgdrN4pzDMd8cMWLV82RSWh0804xwnzByljBXSDXL
39ng1+BaJgmX4bXJdspEQqLOstAnZh2lPJEaxDHc2etUk2kCJU7hMkgY/QVlhGGQtfq1spJdD8z8
9vW+9OL6oCxFyOlyVQtqj1hSc0eCL6fSQCyFsg27o66XLawD2XND9dX/RcxCRvLeX1u0l4tZ8Tw6
KBuaLK9zq2CR8ynU4avgrWfNv5ZwGpyNHifJYW0waO7T3axUX+YrEGYKhpL19W/bShowbqQ1B1qI
3EzOTIMTpf3zqL0zYdNhusnPiEyVotSNLiGv/yB49A7bx8WTsEJHUShCKi6zLSCf+8WBXpZVD1JK
3ti2NngcpPnpfevZhXFPRwckmzBeIYboJDfk93eaiuMzVriHcZHz187WWKFTdeOTgDOoK/jrwHKE
Vv2R37+F6FUZg41N32mptguMfbPCLYKrqDHxVa/Q479M641uxTrSJmP1ZUC2X/Q3sYCAP9IZ84rF
ja74eFMa7Lyg8pUmDtwi6KXe2g+uFDyDYlZ1AN1jDo9kTm7FgmP+Voc5hJOrZYT4v40B/IEtizdE
IAciJR07qjzW8fsoWASMbIlCG2LlBpn+nQAF7BFGOC0bSj4RZlSkgxluY0GQp6TVKEc5luM8cqie
Is7yYN6WbA8OSegwAZHppDzvuBppy3oV1/XBgjeSKGpl5hOfwQ8tC6otFh9VGSlnoBozCUVtjFbo
uqaqH+2KasVTm8TKVUeWktn1ShYmLxQZHv7r52dbiqOo4sSB4/CqdMUpYDUQ70TVqoM170RaOuSF
oIwmj3MoJbfheaN5Xf5C0roS+4Bqm2cEKU2apsWvSju/t95dlLj5kstOCWM/8wrtEvPGpofqSxke
xKI+4swIIfniJC+B/0kV1UEaVj5O7C8huPNGhjG3VpkK/bwz9GTTVTkLI30Ymzq6x8BY1PygXQ43
dVzx0kHM4UVM+4g8O081f1Jkt3e1E5/79bMpneRF4iObpBLf/o9DDmSwiJgobw3jz7jkaigTt6nb
142UkekKP8koxixzBQsKlWBTM8j3axIBWcz7l19bbx5Dp0QYaVTNd09KSI2Ri4Co4Y0147iKBHoz
w9XUzddZXRBju0IFz39W7vJ3pq7ICqjEdFiSbsouCNYFni62BlLLKXsIUIJv4BAgCTa2bbwYU0El
kvU3bkLe5mjZJWoVXx2nz0BhQYdeLyAWBk3EiW3p9utOOu19fx0n54CBtjMRXE3pTBYooRgbyvAY
54TGp9GszKDkHhZLB33l3Lj+KrCy5xhZk70zYupmw01OVYOgSX4ZJylY/5X5iYIq6vuAEY6VmvgM
deV2WG95/bA+tSdPcUKjIQVkr4jXNKZ8S1qAABbndiK5f0f94S/UsRMtf55lLjywYeCF9wPQxzNS
Zjo3IDSN9DMj8evYKULYvdSlno+FK1kz0iteYKeMCG0h4tP4ogXPXjGvlo0H7MAaB5fy8xoXzeJE
alck/J6fNxnrVhS681g5oj4L5JctE4+/tBtIGK4tz5NZEHd1Um92IKRzDVp1MxlsmlV8fOK3wKmm
/8TUsCZFaHjmv5Ku6CNYyRCR/FrK3p+4Y8mic/JgyJNZ8CVeanBGsO4qJ0T/TG/kg9Ihntq1ncuI
DsRPBFnsrH851BvI7+cNKR7I0aM5WIOnqeWfdDq+k3OHOfYBY2TUr0HfxIW0bhJirnm0MGZn9mqO
Shph7SP+/OIuVq6Whbk6xSIPANNmuT4fcBek0kShJi3X1b5+leKlVOvtAGAq1T2DxpZqn4GfyAeV
GJQbIZ6us06L3XZ5NgcC6NEe5/TvayvZVo/4vKaQbhLciOWGaouBK0mNyFX7W437wWS9U0mmfT0m
gUbXjX0xgV9f7hBoJh95/hhAVsAtHOkYINGfekDWmjsjO+MUFG/JdwKz44S8OXTezA+LJcACqdBj
rK+pGCy3PxPMQ62ZrEiupBSZ0zGF6wS3fqXP42xORBzLjoYS3WovHQ4fNF2jZBe5bMYCW08lNSaX
cWaAy5B8jE4Tcy9vMmWnPQhm+G95sS0oTMZHsX6Nnh2EcQ19KFFhd5jeioFx5KWXOGcZF86UMw1g
ScehPqyVB1inhnfplnqz3I4uWKEopMisgsLWDaByykXk5dtv7kPRFlF+s+14hIJ/34fMREqFC7Jp
aoF7ysgBl2Yu9dQgBhVQYbK6PkDzuIiYiJdA+0lqMN6IL1ZRK/A7MuxfldBJHcFzvVTbnsV199hq
OAlD1fjm531lLRlL4cWY24+AIKfZe96zA0O8H+6nx854SysHV8M6dfFolMIJItqXFJdKsJrs1XDj
G1hhMP0P5PJqVU4kn1d2jTN8JkfwKUg7yq73Bruvda7kdgQoNRnJ2MXAbqlhB21BtD6c4t6Q2by0
+U3Yy3zgeeqgxfXJXdWRi7aWOiYkRL9gcJtFeAFGRzc/jXDkPG9jSd64yxbRuAwAvLaDyjITUQE2
t6aNGZKnjMBQk2r20wCwBbNKa6GUpNUfJrmpBCP8QXyoC1K3eNr/Qmn66aiqWTkjAjG9YNfxZS8V
RwQ3GEA1HExYLHAdrSxCqzZw11Hha5jotPT3pAUI0zqXDBWIkjFoL+xlB8cH7fLYYv5J+H7LXLMa
NQaCuEHlh610GMDZ9I+2ZUV0XFcsyXl0L4qomLL/ST+yE5WrBVETON17Dd9ekcTx6fKqkZXQC8VM
3clihfVd+64UenHyI/qwkUAenLLquyVoBIDYu1uv1Nvx3wWj1Mi+kNsER103/p+r1G6J0cp6HUOV
WLGI+T40kzsKnaVWy0qOO8dlmTZ7uoI9BCB3mtEd1tCFYAy3MT9t+sU1ebp2vlbs85SDc/opDNDp
6b87uF8txHaA/Fzszthn/O26QG8mSaHrP8Fu5oVKdGzjCwOU4Xt3VvyARHgVVV7CE7Pj9O5742qN
9rRI9ctIybGc6EOI9xKARN+3zYGQfzpGQSyvBb7OEPbRLrgeYlwzpTE3VnWCT3AUpB/GbzHRtnnk
muhW21zIKJOv3ztfdRXIlaHfnjdzscbAReeB1KLt/a70fFwC7jf2iV+m3Gx8Pj8jHgg5MoWkgdpG
vsX9VyZC4+6DaQd3uj3JqXZblZTCVLcjUGE5Vx/0cKj4fg7hFJJupSXrOrbWfSghMUvCwkttZrs7
wLBG0kQThEci3XH+3zO3qj37bIN3OjHTRHjH1U4c32Z5E93R3HXN1ds540WDoppk6vPfq72fR509
jC8Zoru4ywq9zIMYt2JCo3E0Ve2B5taTzy9lIwvwg6bH91MXQ7PRQ5XXNMsRBwlNeyV51ZtQ1S22
miXzju1xf8E6MedIP7dqXCLsK1gipYkZGBT1877vMbKRn4zGto1bDifQTndKPDGz7j4KDDtd9853
nnO+i4TBnHRLN2qKMrfmqTrAKffXwXUwp9yw7PKvg7OuHtePJuDnBvkmScwsnZ2RFpq4Z+syWC2W
Kg08MGL2s61mQTdi9xSH60MpKcmPBuptj+dq78rgwpRmZsW9rMJisJGun07e0NRy54m9ehmSh7tt
h0k4i+SsUf/08x25sbyeEhtUHvZuysiDjYGPPWMzfPBsglYGVLx4LoLpO9H+MrLjOl+X5SCugB6h
yVEZKKw8lW5xJOO61U7IkOKOUMYysGGhVVrudInvRCKmJY+DkV8SL1iI/j9OKQZJ+CMrL7etWNWF
1JyvDNcGGsf66x0d7ENRw4SsxDpvmOsn0atDLCpXz9SA62avhp2z6n6DHRtGAg69OSwSNh75SMis
Sb8QQRtYNNqH3JhHu9bEZBuCAON6xgjoiu0Z4gouHKv0mZCkiRCLHK5KQPz5PME9ZBi6RFF2BZlk
ywjBJx7/3qYYy6y8LW7DqdGyO4VVX3fk8/Y+sPtnVeQyUsMBaZLkPDJM3F3WFqRt7I0fX8GQc/UA
3gHeSnTAaDIjRiEHBtdeE9VDSlgMd7n6upabxnfNlkvou8fgJLp60uTE23zjCtOiE+OyFsmcnMg4
JPQrRty8yRKHEPsCilcrysNuzjEBmJNrcst4KM4w8sxUjJBxCLGzTWBhF2Bv2pFN2REV4kjOUt5k
JkPYImFdxfPpZuv92Oz3a7baRel+lHb4uNFwsyrX8L0RoQAy6qgmBRM7A6JWrycubivMF98+rcK8
DyPhiuoZNOaMs5G7zCbXstDzDOWs1zHkq0O0RyITvGsXy4Ihy017DG+57wEZS3HbatHW9J5FIMPA
SbA95vq7klIBtrrOcPr/YxWIpkBxObwd5puuPYtyCGhVI9tO3zNn0+J2KZ2DxmlpoGndK2imA0q3
qALKM9IOGImfsBI9d+jt31i/D6sn9zf51IZu15L+CI5XfdGunPThkiVcXKlFGaxz62L/Uiy3G1du
dEjd1y0cDuGvk2K1YkgeKvC/K7Mkq1wNlOAEb/1+vsoLpqDz+U3QFYaV6QIr0F0WIoYrrGq0YNnB
uG0r5fkQsIxTWREMSnqQFu1hdNjNRJfQ9oiX2qJxUaTmB+q9FqOOpMowZNaA3+fvifEVoQWhzbQ6
0F7o47vq6Lj4UQ2mXs06CrURMumrlYThbpSgqm4Q9PIA2Eji9hK9IrlUA6O10quc5/W6fKwYPsF/
v27X4S6jqsRlFuv3PGAJyP95oMZa2nD9QRSsrM8Z3AXpb0iVznNjnNWBDcxIujH4y/LJvyjDmRcW
ZluYT6GthjAuHMCiNfsW4/u7cx9yvJCm36ej/9egS+q2J+S6TzqELDJRFJgjuWCPOqY0kTNDZ8uI
b3cKsCHT0lzofHuCiR/fCn4W6OgVpCs85V2653b20FWKyN+Y5COOj1nJZuC3BAlKdhc7Uru35+sP
wDKgv9iGWio8cSmfW0sHw9bz8JnYSZ0/+HJRgrK/IBwbettQonme1SmA5cuHPQydmCfXJa+LmAwW
uLtfP3UhKVuPKkGDyqi62PHR1MiB3FwpIVHhBZVOdpjxmReQsHC6Az0nKq9MqCz6FDh19XbYfp6q
4b1yTCmAAyZkym2sdK9o2Qa7c9Tf7Kh2af0054j+LLItCIaYkzYIfFEi4vwXCbZLbU6W+MsYAKzz
LTF1BwUciBJex7MbO3Vr8RdeEoQJGahNKuhOxMC1gEFaH9YDYuafkhHHK+f2WZBW6P5pQoedacjO
CPiW6xVdhcQTfJipt0J6QXRkwe2hJaNaOmRs9AGueU+OF9Sc1P5eT+q7rJr3rzsRTfacNlwM9Tcd
trZzwxHgTA/bypvwmCiBHMS0yAgmqQ9iqk8tsdh+jrgWLuTehWEhUJba4Itm4fJlNNlSJX9Dnx+5
n6Kv/cvLUPXSmhPn1mPTHcrx8P7bYnnsP6/HfDpUe8vAZ8GAEZQq//2AaH7vPDis8x46t4FwLmvq
kbk7332l+XyMA6FHie0e2tXjXfikNLLGEgoX2KEpGo0lqtfore8WcJ8a+JsbzzU5HU6Hof8V6B6h
3KEqOxwjnX8B4ceqkGxLBE0bVKgFAwKvVYQ7/CIqFBQqbcfRTkP+y3iVrJfl0QOQWsymkhxgenCG
Ljam4j3F6ZGi54UHo3ph8vCqk+yUQtohVkl5RhPf4+kqHE1ZlVqrpS0e/TeHB09Jn31B9ZDbn6Iw
tBz5LxM20OVUMo7+/F7pcEwdwWUaP577CYgVu6zamwYXD32SRfpTNEX/lDeVSHWXrs6cyqnX0KnO
9zpPtHHByZFSRKHZ7EPS2u1iVroxc2IQbm6syH4j4+j15TC1m6qRnfwGA4qi28jX6EwhMhCNWuBG
F7ZkUHtk/f/lJHu99d3+Trcqxs6DKLQsXKEBxkNXEr8nEXfYTwoP3qreuP69xoi2aZF0VZGhHhSr
pttuNuSBj5sLiIe461qhXmsmApwxXKaLVpTp56sy5OwY81MmzgHUsb35iTJ3IznsJJqlRzjYePon
dpTBME1eLHaFSFbUPyKj3ApiIU2Loi1XrIHOHuswnYUs7O9VtArHHpvRIBnalfHdkzxJaRYmRGG8
aWEWdsxqbGb7G0Yb5/7KdtZJ91fVuTBeN38RKnFm3b6yFiT/eIbLy5nA0SgpOtcOEayXcbqn5H7a
VhDOnHtoKfvjj9prokkpJbjkKD+PoypeOpt8dPEU7BFEe0AsD64F4JWXhH+y7sgg284RHFmMc/Zb
ww91dG693cffMCcxJ/af6Odw1yWSwmgm6WPu5irMcCIX3W2qyUzsKy+PyR4VLTH7Bfo+nytSsLZg
UlTDyZNJSt92sZGjR/IMjpSIGPmYF/246nWo29RRNTeYB1v+KLXwoGG3RhDHlyKMNPg8PRgWsnfq
tjSjWJ5qGZSQgwKVgT9XczhyL5RA6Yvmkp/ZfYX7fnKrTFTomB57Hd4TXFgLS5/jM5E6Oa7ipRwn
dSXyL10jJwWnf5vfhlrkfOIRp2MBJZBse8PMTeiJ/aip4y2HSaH+8MjRJxrtd0BHx/eKW3LhJJBK
mahB8bncZJwfiw6FjMd671jVOJPAYnMW+NRvKlQdCD7vHhVAYEeP50GXY/EkWL74M7TO95DP25GB
MCUJtRXUjjqvqEJoE8AJ5p2GJLL+L6qWAZnLghMfeppjW32oTA6kiTvAm3qlYIka7xvPW6DrhCpv
MI29e2S4UNyJCw0toLc77/8fGde3Ywjg6FC4HsfiLefr5FXmQG77F4mbYDHslH8MyjrVHcjoy6Fb
mtr9Iqjmp9nLcHgDz9snfU0ASJ0sZzNWrFvn2K2EF81uB6OWlAa7kIKTxzRbPLcxNb7KRxmJv3lI
CykHdp+cENQKbqxLGfVVlnyplR25T44zXF4FEdDY2AUN4tEKlUT/zmJC5uJcRrHgtM7o+/V5GYUE
MAUq4oVUwwbLnwZohU/NvECiO/vvlrMrl1GWf2ecVy2UMaXV5zn1Qog0yq+092pILMLg2IE5lYTy
iaAqtfpfiO9GcsB0TIXejv+03lyRstZiz5rYAY9CsQQCFvWFMbQQ/NZ/05OhGMgl4hkiFPgcKR16
ZcRJlcRf9CsZJaIr2fd6SapFFkRuXDiPjjqptMxIE9y5GAiJY5+xgyt6o78f1Z6s3l7SA0gNGy+5
Zjj6smJAj8f54Hg0emc9MkbSN0kPl5jaBLq0lfaJLgveSAocTXru5tE5nuKAJOlvsDeeydvGAreH
7UoO//N9A3XL2qwyG61+th+8ZQOY7elgNgzZdnZBXW+n9GFFCrDRPTlbGJfG1cKW6j5HubZcBBAF
SfDuDj82hnLiO0LnAlbUoQEKHJd3q5YvbwG6VH6Xe/Eq5RrjdKIGliVLOYnbMt93/TuCXOXpWzc8
8BObHTQrIua3IodnNd4Zsoa16e2IEeJEXccCDzRjlZzXsPR2SzKx7d+rjzFvpW4nPRNNYidw8sXT
ZCPkHg8QF+L67XfVgypLKsz+3NJLnSmf3HEWFKXYdv0IBJaVKqz0IMtjfMYcPq/fo5E2YVYTqBig
6eAZMhvIbhEhFwqXKXc2qwOzMHEHZd6U7iaFxr4AiKIzChscOLmDG3wZs61BHPScffH3ZXHcz0sv
JMV+rQTz7i0V7S/7rfpPIX69iPnhlz1uuoP1dgMlZwv20xTuKmOMoZvLiNlM6pn8FJvXlw5KA/FL
X+vVBsNXJeOAaZcgRDtqg1IiWZSAxGC9LhPl8lIcdl2ujOv1+G6fXC6b2qM5yZ+VsjTbY5ihHtz8
Jd9ADC55UrZG0T/qrVQsc1rEysJctWdcdKJPqpU3ZeJddk2s6AQYorDfjiSXkjWuOVpnWA+b1UaN
Epfm9R6P9T2xl+wZIzmndgzOq9IhPaWVNgATFlopQPcqngN3wgBXrujqYOEvps/mzg0bnFQcopKL
N7xSzdzZ8/fYjzkf/8u4fqegXEwXDTjWcMrQTSgaqkx0UnqjFBDvDaSlYifhNo5ALC4uaieWwHR0
vHeV2gK7+Jq0SvoV3ZbBq7mmHqMLnK6gFA1zSUdnsPRbzU0E7l9dSrAom+aoOXxh19DL5bnAgpTa
F7Kxw7sdEjijV+tyF69r8J1xavUciDIRh5xc+R4ysvDZKQkgILIiCt7ggBBUJHIc1jrEugGcVfSb
9Nr8tDYYbtFbpB+f4Toi+ceFPBHzj9Ot/DhOSMhA08LE7jZtosDcZO/nevlBHIYxTaLmpeKGC5CC
3h1A83qEY62ZBXIPrjjF1+7vVki2HN//urJpJFy3zriBXu2t+2D1Y/b3E0SbiEGKchYCzfbd5hUE
iG/1xEhuJ3Afr0h2NmaCZp8QQLwI4g1fR2VnKoEMEm9fzyy+pkpZP0ds1eXzG1BqAWqp0q01f4aH
aKitvSJJtV0C4wrIheSPR2se5mi9OuQQTgjEhSvFzOC0UgvH6WPcGRzcMP1KSp3z8fz/XN6pt4vH
ZZxE9Yp9IuGewJI8sCXSKjCLR52+5cmEpGkU6Aulo12+hlnCu38KUt3UTMU5bK9IYEFLZ7zOH0BE
pACF6KhG5J/nJKe87rwMwaeLu+3wEuhbJY6DtQ4FhzL/am4iGovCtyZR355nizuhMtkRCsIbiGic
BfVtZaTQuJNvQ3ajbZxlA3t2RfRveHIJQpVFrWEmhcHivq55JAUTTxTgqUsLXWDe+ZYT9xqWUJ3W
/dOqhKKRMcju6qnCK35WytJuAtS+PzWmwueMVgvJdYP1Fpi3DM8tWPVx+RM2teItef4yKhx7GJ55
2zp2tUZoPWV1E0C4lSSmcy2ChukUJDV3Wgh9AAoKpv/0iPGhLFtuob6LI71UW6XlAuueXJ04Hn6v
pOG0Cn/3PZI8J8D2j+WeXcf8VCVKuIR0nE8F8//Pw1mpFxjzJk/rT9IL3vzqeA4RhT+VGrntSO8m
kl/jKF3lamMH12vwHVwMl9gk3OOWt62qEi0eLK7VHkOIXVBadvLmRTDrZyUmNWqZZ0X3xHSY5Tb0
u0iU6uy1B8CxyDC+uSA3A9Btl2erteJfvPhoDl8Go4CFmUIkJAPnFc1cfQv5uyi4czzw5l7iDKah
Oj0jCYIHQ57U+hfGsjkGDW4DETwj2wki1FqzznrizMdxMba04NzvrouJKj+70NH2KwvC/UzjoM4O
toYBWqLDWGdh5GylR7QgXN/CDiHfqKLYTrYSpqM7++Jmu9VL0yBukTmKQq6n8ytX/+oZDx9iDBRe
sNpc983WkQ8S/4Cb86iboThzMmhsM205KQvqVGlK9gI1yoxEPzxZQIgS3eKSAGCZx8lHj6dq9sZB
WVMeon9RRcw7mja6th/nJMdn8lZ3gzdl+3BFTYvDkg6ONQUE0glBtG1dMyDRDLLbUOn2vJop8APo
IqJ9Y5u2/lVl1blw80+5S57psFeT8CDOcMEKBLzXc4VbON6Feto7iJpX+JoDWG53zr0gJ8QpHHe4
+3bGZ/Y62TvdgQlU8NHFVeZniQy42ovgoAJzTNj2UcQjiyBOrATVFM/RaZLKPf92DnjMwPReaT3L
LGnnIr3Pc4MM35qx4OPtB/5GpGh99WZG5Wy3SzhJUTq1YGWV11Be1XvwgJaKhm3I2aXP2YatS7fz
hTgOj4IKPltR16VOyFHtxp+l1vFL2GQ8BE/H+tA3gfDnhQ7Q0JgUYjsZOA1TmHhcbqDBKl/uJ6pE
94Q3nR+KaxG/a9PR5bkOJ6lazCMRc4JICvch7bUl+MiBUGHKP+xQ1Oao5U4HHUNMSWekOfz3JKzj
IQStlGNU5nV0rQNW0lh8KGtn/sZLyx8hxRTnonzikqS6GKAbeSN2hnSJojB4mDo15JIsW3Xks1+O
XIB9hf68/mCdpe4nFtS5QQC4nkvb0ztrjXSSldm8TMGTeVgxcU1n0afRj+sIUkIxABDsZxXpqI/E
gcvLlO+dl59gVe+RLB3cYzIjn6yoTEwU0R9QGux6eWIVzSJLvIi0vTG8DTZBIEEpNUoHJBKq3lWM
tuw1FC34pz0DuedNBQyUMBG7B1YINSxHfi8RsJ3XaBgQFboTb7nk9GAkfuoXvtblJz9+RICDN2PQ
1ZSVtETbgZRcZLI0ZOy093/55q/Y/60j+SvirB6NCWQgoSAW7nL71dMA9fHKP1p5xrb1sQyOvLUO
hqBVhzFsEoXMtUaClJ90db5Zi6pM0/KGcL27dqKpXgcZ0Y4uLOdIGtk5BYXOu9lGm+76d/y2Yebf
NG3bh+2AzenPATlJ7exx3UYBRdV+ocZHjk3AomSeGgtvUZOlM+o+xJ4U09bxIieOvy9cWocl/S+h
3i8cNk05CQrR14XgEYtH5CXXBqrbghPLqjPjw5Rrvh9CvtJZug2Dwsmp/r1dk8FR1I+9yRw0diQy
BcosjkW0gI0QDGkncJk4PMULRYKY2b6Otg6ENZCvybe2Ty25JAlAJNcCHFhIwfLPtOP+121AN5QQ
Dbcx150iR2nO4KLPACSW1XnzW7FOLp8n5lkZbnKWM1TTJOVf/bjOkZla3E6D6KTjmkssuQyJNx07
+Z2pKjUKjKH1eI53BUAvUe4l/WZKiVMKflmTW/kFGMeUGNzyAmJoE7VF2mbQHiT7e0fBbA7BdII3
7b/jKDpN9DhXI13NGruEXQFyzKoi56p29jNtpISKGxsYQ/NMIHRyB36a38I/REX0ZvQXfAbCcGqp
9mMz6EgCuZ315B4eE9VQJ8mGtIG11OeGgZqsfUk4ZpLx8iVqG6TQnwbh+vsqmsNS2fPo75QmOB7f
vpY9ASTDscmbNTfZSSM56GJ5Nfs7anclhRLyNmJIV8/U5pSu2FFxFJ8/BlxRapg6rytNXVPloDO6
CfVENR78XkB59n/q6Sr1xky8VFgdpjYnBve0yYnDSX0cLuZDYxJF+bprtt1OKBTCjSlvx7NjxbNd
YMdJx62QfNdAF0BVkRR4QT99EkFa2fyL6yqFK62afdcOt5sBlB8cNmgxGZ9jjLlBqyngxcjIoJBu
jxSsI9PrzNR+fJtiz8bh435qCKqlHGUEZ2MufN3XRttq7nXEyUo95v3d66vUar/6VSOkjnb0HcbS
+tLyAsEPOYmp0hDk0C6JfeZdar/0TIuAbi/3CI2BLjy9rlRwdbrAXE1pUn85K9iSWOazZPELOAOn
uNAidMud8U6ecOPpOBHoDEMz1OZkUva0LRtAtzqogCzlUiR9KlFeEvnSh4C2PAUJ3Juz0KnzTkqc
f0sq5nKWFgnDZiKwGgn9DJ317waFgtdehzw4byU4MVBrMr7JtHIiw+hp5tdhlhyex4ia4/NKsC5A
8KxxslgBFZQcsGgTQ3ZKabYicsfEqFYF+YYM7cxeVpuAUoZrPZy2H+j1ahfrrSUtiGsb31KEyXak
ebNwSyRimVvzcsBYwLqOqXlbFEOaPKvQOn7CRFCkxJHUqoxVAdDc6rFT2A3vh1oaVqIGQj6Hibxo
Ijs+UbFUInseTFflKfM4Bv7k+drB4bshqjpF4YOM77qoGsNQcyg/EujSnbaGVN5+zlmZz2ksJBoY
2cY2UYqMoqp5YvlJK8NVfydCX3+QoSaMKnTSmtMqVXUr0RqToD7/V1VZNCm1GuWboDh11TSQm/ne
tbEVYUZIRg35VYiOmogUMff7sZWAtCt/iK6iyQExe6icJAoNoAVivvmHGIxoliq4BDLqY0ddvcIO
jNmX/Em12zizbn951RwXZ3lOgL0tVMoNEGOIPoI29OjWGJJOUJeTJJ1LH4eiFUugFoZN43Es6WGx
uA+zNFXzZ3hDYIM4cwYCptKHlZp1EM4nsN2nXOgNpA0wwqS3Z3x3ciiPqE9ObKFBXjT0tSXp1wlY
oX13CFgKNVyyaj34dKuKu36m1UsJMvS0AL1JkWemCdAnWd+GhQua48BJH5/rT89CVe8t+9KXnTqA
sh9GPag/4erT1evJvWP3CF6Wb4Lz2B3v9K83i4QqL+wvskDcxh9vYELKDSkq1fEYI+3gkiivdEI4
xaWi4L/EYb/Q2JIPEGBtQV1m+WRjoSXwR6cD+5RgWXHmkGHNYXvO7N717BPJesKnvEU9H/a7L9kN
VU9OgYvIoxiIvfz/vcDBEVqIAMhcUBoMaQQvmWYlWAiMVBlwdBW4KBGVH59XEc/RdKBruPTHSGkx
rdfACte1LV8R3LvOlXdFSWzPyIHSkpsRx/HsVhl7mjcXJyJbYtL7/fBJPNxVjzQ6n8aNAmGhb3p1
KCyiJe/ZaXv8R3K1yh47KJLOZWis0zXd0Si/M6XrmWUQ89+EABwSCKVNSCBETmiYA3oXhCSQDwcj
1UII1Th4Wag4sibF2ingOqPgY0UQ/ZUu1kqKOB5Zy+OQhtJWlLRZteNFYyOHR0Sg5vcf9FvzPiwH
6qNLanBiic35L3R1ewMyTrTvgKwLx9p7Nwh67UCIWqJCR7XeGgm1ARVamwpCTCKT+hO4A8nyV69v
3Txhet4GTFK/Qev3bF2EDS/BkxBnO7+T5KCcSMEZLIrbdLECIXEmOUEnNEGo9UCdDHhYGI2tYl4L
g6sJJlHr5RBznjZJ5v5xTjlsc/3IVAhpyaNIFFb4YdSgNXE0ZlgVpcOG31tRBXowE8ORF+AYzioT
q1N1HxEuYwO2kJfdlcrU6Q5Bw4IEKASbfqz8mlsP9UNB06Lcy3m9bWof9QClNzXgBKdi7Ff/e8CC
Es7MtDwOoHlCbjpZJGusnJ5pMnsaFC1FZ2qv4FQP6mAVyN8yAB5TC9E86cEHhd0nELEmuvDs6GiT
MSGc3WfsjMbHnvk9V7XnJtZa6LVVw8uHhAVbj9o+ineN6bMF6i7XJLd9PIkIqXSxgi0TJ77RdBpA
vhcbcJpIvv0e3TjSKvKzYTD/6ebv0v3v7/Jaj7sTTEEFFRSPrbstVQY7GTgbsE5x71Go/3F36Fr0
fGpknTulCMfNn2T5xIPJWamdeNP+0O6mXNYPy29R7Wz+GIYFexkxf1GpsPKM9FzLE7ys84GA/Kc0
cfzUaN1k6GwdTUQ76sh7AE/6aZIByOilx7LBLkiJpQHpDfHWCcg3HN8pUMUjYr0Wn7fYmuJnkhp9
0Yub/kX5BrdnCJoUzu4X3ib6YkJTZB4pXwWIR86wTguH0RnTqyR4Yv2oNADo758PVHHZGEGwRV25
Xxp8kaBpCIspdYhuyXc/51WEIuroSCCFm3IN0PYvOeM29xOuZ0xkCzNaOL59teSIEIynaxS8whxA
oKKwnzWzQq6C6hC4o6z3LqXzhVimBaDS0FWMFBBXKemn9UH41aW+EKNQcgyoruscxwaYa9AP7Muc
8OPtBoYdiqHgc2EKUfCyXAPs1yh9fxuehaIWgrF1oXB6qsJNZ6CovjZnHkwiwDFFRLspG2tkqHc2
a1VBxOyU0jBz6oEb0CujdYrf2/AY6CIVtJwC0ZNgxHjkJb9kQbahwZzwhfUljyZVp+rP6IZho4Kz
dsO0z+6sbA5eLCE4Kvrz/gBh+T6+iyGEN72YKEIPqV8jz0JQUID8XTN1yj6ok6GfDOCXGFb7ABYL
t+onQ/T3bEHxRPoKJEsi81QlWTKkNLYhRrvfX+RhFDJSIpKYkhCyzyfG+wCvMnxcZqslALzLD/ZC
rfBK5JI4iDPgbdMKw62zNvBhqL/HDzXGyQpJWBQB46O6bREMolfcoLhVW9rMFw/3Zffogzs01xIg
u/YAnA5BzrSmf+AeEdrVv78/a6xw8zopNCne/4pJ/TjAuQoJAsIgklpIgqhryD5azD2XdJxjAyOh
4Zi3Lkod4aIR/cIEcY8ffhYJiyqW3Ii7tw4GSqOPVBlec30fDwFQvpH9rW+kuScjsOyJGSqRlDx5
3/vPHqDpi5WcFKyZZmYek3d/6ae4bFBp1eH6m1dox/UmLAxMSvvJv4SM8e6ro0WfQVgsUSCUKyqR
FbFYbuGfly7zsgDIDCOj+GBZs1R1TrIgnXMhqynD6hN24+9mtvg8e2TY6g8yyhHqfa7iDyPA2PRV
Cv1xIMYG2oG+n/v5KrUBgtglgacpKT+oH0OiRAoDX3hkrdS+korURDLXVkBF/630qivAzNBdv+V8
K+66qXPyzaalzmrrmmXbp6tvJKP4s943L8Dujb5nKwkYgX9iPXjSJUdn9aSxxjUItKLLOsvFLN5U
KxiuAGf5edB3p/apZyvKg3t8t1jxIX1x5eAHoH7WzOBxBp/H9H7zzbA1/6yWxDKduKPLvS0F3ux7
ZQxvB2NXBShZtzty1pnri64VnKLvIMqXgHGukEXyOS+8FqsVtPrb8O66E+B2vr9kxevnV3DrHnV8
OFPeWWulrpomT0HekWHi1OJDxTJ7Cmb/N26bArDuTYGC/ljmbswL8Qi8UGVfA6N+Pt4J2zDk1z+z
bEqoEFk7fix4FOb6SFPTs0Aoy309XrT2jZXeUT9HcL7bJH3bIvNgGfi/aYxUfMqtzrKJV/Et7kQG
aLAxcuMImnU7xja2WrH2NcuTecgGFYldpt2SUBpxj0sv5zMqIgDRc9hENK+wvtBz7ppdrRzohXiQ
RLZgY1li4RMLZ9Zuii31vhF8emvwOB20BAk1dQnX+38e4Cpl4Bd0l/NR2cvH6n7sOnrJa3pk7jrb
E5It6GL9FR1RRmq8QVOAmN4qSfBEljsNyvyonjHpArj1Tht8V/81iFAEB5vFFPFzOSsNt1YOJ/5W
nBtF9QRPQOS+Fn7BLEeiq7Qkrj4GBi9RyGpx/xw4p5httu4BhqCsS2cGU2ENwJFL5SKSKckqRceV
SY7kUNf4vYErmXFsHtd7m3SHzEOjoW6cGsjdiWNI2o8YPgMKNsRcybfwXX/3jbOXGI9pQhzSO0v7
q5UusflymMaYX/iWewijsG2eyzohdBkEvABk7wYBoVgsKwU26dpJi+I5chRQKyH1IWn6KTpUXsit
dMev4k3zhCYPrpb4Mje/e4kCY6UvUCIcxY6md5VSLOl3qdNbxk0n2Q7TGhwlksbdtGiFLurJQlKO
Yg/NTL8tFsSgmmezNmsGA+efWNMg3F0ZMpI4Xzfd2emtLvVin9unoctpSsiKw6Q9pqvA86kqmxZc
gHaAKZpF9qxUHoWSP4eNkcdvl9j9qnqlhiQ5UjBZ3qbwS0ooE2K2Y+LflBaAZgGETVoJZLqcGwrc
6j/t/96aqVMHA/ZTGKBjpt6nUndRZxs1LfMPgW2sWCPmgxTwyUVxSM9zhEfs6OPcHex5uOCIA4W4
Y8g0vU7Ce5b3aSIQeNd61LF1M87F+CjH1t0P9O9QEZNso4r3sql2CWBWIsRh2lzPzQGzK7ZSPm31
tn6X549QE6y13rntQ4OpDzE4uWtke2QKaadSjbABqk7nnjCw0gn7dIK1CvKN4iDZH1Rc1qPaE0yN
PB4aIoS54kYaA1cO1C8QZ9FytXFW5LTjpqZt2Hv9R5GtWur4W6vDVT2vKqaQE8bOceWeMYqspuMD
p8Sh4nrJbcTUZetO2Fw9XzZDbe1EyN2LpjAcPaiCOeIVYTlgs97kL0arEQhrHWP4IVmJFFnEkGoP
f7NXrIldjNlBC14eVspHLZQikhtwAf9Z3QjP0dIj7WkHFuq1T/X/z90N327Ff+SMYwF6AyxrZXep
xZdVdwUlzSmVlJPg7M3kpJRrL+0Ap5J5erHrHSCFR/IirDoZHTq5fm6I9fbh9j9FmBctt48q3FNS
YDbir3XTWYPDymrKlVXxyrbQXIPvv64Cw3Z8iKH7Q0Y8sjdSlSw58NcxAKS3sTCedWV0UP/gLaRe
/0fYFNUVuDGlvW25k3X+F+SZzYivG4F0PJkOrzdHZuyGdS8PjI1F2wTOFGU4csf3R8SYEQJj3PPA
U/CApm0VoyRJ9974jo1MNdd2a2OG0oltRfoEaCQxfJwaMYjcRceb2Q98Kod6sGeUHLwrMbwrtfMY
Fk8j9kodc21K5OE4zgksCLMcsPV4M0Kudhhgk68TWNZoMZUorXBDlswDkvjglIBlhgICsG0cshmk
rnNPvNrTxYs962YoxyRBWxDj54HLjNXrpb34ACKzfWd+QL1UKsUJLKWVrJfitHWLrb53jaePRZ75
wAaHIRL8OyBKJ+mObJ8qzA9ADPaJyHF27PIhGAz4FPx+6vK7H6E/wHzG0RvieBCuY7D+fEcrVFAr
STmT576faJF2uu2BIF6v3tHQFm2dFc2LzRtXcCjBwi2CaQq4VpkAePyil2x/EOYbzrWK9KDB0EUL
OjCEb1nuvqV+R8HmVFbby4muvB24+kuOwo+IrQkX767cvSsJMbJju5MV7OTlKxwdE6k1RHKhFN7f
3JKX0l68SsiRe7BJhpAyj6tdL3txKtyY8Fut0XINsiOtggPRcbCUAP19W4HviVRXEZ18b7sPN24t
5LFeOcDj924ttvrm+vTVkcPQbLSUEtFGuZNkC5MhBeaYoNfqQ/S7FMsYZtteI889ppPJz+nttGPe
HAWWt/71UTczoHJvtEatvaGmTF7hJJDEBP8nEvy7Q2GcZrzCCKGT/MO9rNWa1l8YgtAejlqaosSo
+4EfconSLvGZcQK9dbgngWFecPr/lvmQmQpz3VyFfzV5Et5gRccL1tMGqUw3OMrOXwqcNKGjbaYJ
1yFt7IfYZ6p/6EqgtPPma+mnu7wQF2TPRcU9oQd+iDzpQdA0SNnJUoStRwlrIq+QL4PTEL5dwvUu
ymDwBOUoJLQbbN3rlDaTuBh0jaEC8heCA2nesi21bp7V7KIfipyP+DzAdRc2Lk1Bcsc53Ne6HBwV
fOBwzV8qz4zb1HM618wuBiwzYZWkVbemBWW1muNhLAk+hq+JUia9VKrv6AT4oqI9/mhNw1hAUxbP
CvpHHTqrwWGTpz6LNw8aS8zrHU7avKJ53jBLvWonn7BJPX1AkL/XgyY3fLCGPLROSODNH9npSdrQ
eTTYnZdppwytRUAVRxlyVVe724oaWyI+Ib6ROOcdl0aROWkHjxeXQOasXW0amjAOKps/wAx/6jv0
ElxOxWPA4n5ahldeYMge376ykaqBLZ8tYeYYHYxnzntdLbs145wCHREvr/v6yBMWlZ/BRX/25LxW
SSgamISXhpnvw3tS10Hou9h2WYKwsyidG5MLQB6rby+iEhB2arBdAzwqb6+xwjyJL1s3Ct99Ymw9
FA8GzKSYIYPa3ESZ5xEvjUrbTXhrNPD2REpNhzjxrooLw9KAaavXp3riAaIlKCsreI04J7dHdBwb
KVRMjEwEHjVbJUgVoiStpADMs52y6I1Ihlcm2oxfH1sVsfcTBxgSiz3tWbbvyNWUWI9+7HzMzGNc
JdSAJdXyhL5IcmMui07wJxdwX3D4d9YrrQs+JrExgvp/3T01BCAbqIBpm7kI8bbEPO1GWXjMCf1b
CyeYMvpbVlYwGxa4cGlYQ5fZu36vJKxtFzyB31j/2OB8QZMkEKa0deUE7Rsp1S6COVsXyiBb7i8z
10y0LOC5x1AMHxyQN1fkep/f2p/nBgfklmNXNPFleB/hxSVwFUUdSvfuSTxpiwhyk2L35PZoXQ1C
U/BZEC3Bzmu/e/bgHF7gbXvUzaIRGkyko3SlfNtPlQHX7qLzAPDCixQKrcgFieDE1xpyO3K+KtkN
w7jqoOobvtc4BRyhMzhJ7ycC3HQYVJWvV96JvgbZJjdmcRru/Vn1VksHfoEoFGHPQumDRZebXwJt
uzW2K4l/s8MartZD/khpG8UrTPo0I0cxuDqHfGq4ZTc7Ni90huZ/FYt+zp4AAUih1t1eW2map9gw
amVFmnRqzxg3gsWvJljTG7Rwgha7KbdqVsqSeDMAbqIHWtKnqTQ9lLsPIb++S+oxZe/aRM3iGLoP
Hlkk7bUI0dnI9vvQ0UrvtHTCA9ez87ZokyfuMcOehZrBe6hJ0KhkHo8DXj91DIOAzK3SKZKLgquT
ib0kiJ31hf0DP2uoIaPdoRgm3aWDwJiO1nMh57Cb9nCiQQKsGeIz6TLYYSBBzTMxxKvlnkzutfqi
4Ps5SQCRCoJPr8Er7lMUlf7SC4Csj2WGXHL3OMjsdkwNG/J/LbQMA1e39gTOJRN9gCnwbtdCrt3V
/gu+ui1YpWM7Bf/32h3RbGS7d8Plp+S2FX8756ZCOAyrGoF2hoe/d8f//rkMaWrChcY91GWneSwu
DnWt9mrvMBPcNsTbAWO0n2n8t6a5vWHsVd3hmNpfgvLfeYe9iB5PjT5sijcOcLyjI1y1bmwTZLOZ
aRuKpfWjuC2ELYDtj5240IPcg0MU5hvi4RB5T0QDQjharcxtpgHCA+2LfZzGQS+8qokXmFlYPD1E
kKgyg8OCCrCNf3Q6j+RuBqmCvbsQlOj3mzQf6cjtMtyOX1EpgSXVQIe6j1uCeXQ4hzJqGfFlnshA
qj1KnezrtXCEvyg2vIZCeMpA0CT07FOb0HEHU/mF6u/QeaiG/Vop/xrogrfzMfSI/Dyjpy2FU7nu
2u3jJWMz2cefOT0wd5RsBsZbJ6EDPjd9sYOz3Yj5MRqi0CHZAV88quvIYk4umc3fdHUxkc9GhWgx
8fV+YTT8cKkUz6hHQTJkAG7R7OfQtC0vV4NAvfqnBSKcji90ALcTEvq6BlgeO3a507qrqheCKTtW
XmFl+OU7bBdI9fWkxSYDaASfXeXofSR6jO2cxXiIBKYLU1ByvxjfXCCu0B1SZGfS57aF6Uqbmi87
Jhs/4Y9gdeuV7dVIgPl52gXvDWa6PHXE/QKlYBRO8gKsBkC08k6VH0VrXqLKKzyN97YEctQpydVd
e8g2P+wrwFNNKDS2gzDcoNyfuq9hsimgQQ9Vxz4ch514cnMmuv/V623e8bkIm+SQHbPKx7L43a4Q
muHLnhvFhFyHwcr3HL/qbgli2dvOloe4as5itU5wzqjWYYssnvHKth7atH6dchYVZo02K4jt7aTT
FoJ3Nz6hkQYDAbXVRbmHUUcdUY8xAuZ01vNBG54Bajb/gsoOb8ftUCPq6J2U4nJLQFesy0WbPMSB
0I/UZtFRQJCYyaCeDXaXssm1rw70YTfef1uA9MAIP91+xTh9/+mLatDb7pJQFb70ECkA0vHNSnUH
69S/WMT/y1jWZGqRXJhoO8j6U4AQEqs96lb0EPU2/byNfRJHr3yC1Ui+pDxx1pPS64sb/isnjpDR
5cFSABVFETy8Jccr9M35LYsXYGv6tGpsTFXjjux1N8jIfSffbQibxypBYNetadyYxvLaVT+3xwR0
XciXsyTf+cadcuF9qd1VIntnFnVtVH9Q6rK33ZpEI1OMLj+9yG/jnc9nRONdX9AUpXdReHKBFh5l
n0fbsi0E161r3sa27f8ag6vpAFQbMY3r7rQOl8CG+5euprrUXV26PZuEndk+df2xPyij49hK9rHs
1pwblX+8xtEFKflqnll8tTScVApC7qPdNJZCjP75nhPntoMIhJKRN2yIlGbKvVa2YsJPNaLbwa2T
bZa8dXMeQubLkDPu9OIYcqrLfaw4funuFMnV0UWX2PNKqPbE7BMPHOT/Ii70EwPJMeFoHGGtK2eF
+aGHSKjOO74JKWTiyfX3iKUfcqQ7uQrv3Jf8Baa1CVNf5tUGBk99K2Yi5O/IbGW3blHZDqCH3KKA
VV4oNr0RymJf+g972L9CrsqZlsDUU3cE6t9KyL8LFn1gOpxSAtA7g0reC15UEydbmsHXs7cJ7ZQf
Or8ZbfpJemxrd+xgImvdWG5arXC9MMThvb7ePMaNB1+PZ0myOMknZmIwLVx1Q23EqNLEzOnZWff9
wGXZLNTImCqzvjIzIkrjn/XhfG/G0kLFBCxc3j6EkxPXiQD9rT7xfI3OuyH788UqwaQKuQjKg68B
5HOEZ/3dmBA4nCmBgtPFdVhmM9ICrBGFAEJqAxuzoTamXDUupXKP5XvBX4ZU+ljvKu0VnYdepX+c
3RJupCVRWKBYi6vsxPQ8GRd/YY87MCVhGaus+KbvgCOlNHCw+7KLS5wggP/a1Sxc8D3tfF16Rpl9
JMGGog9Pb8sqdBrvcAfg+vaq28Kr65Vce7Bnkdti+6a0hPbK2KSST+o/xh51NxBKrLZOLJCfaO5o
3DRY7elG1m08+0F4HgRqmMpBahA5YrjvM2pJ93rrTQkwpAeEn9OzKydnM2JrZVvgkLYvv3JeQCs4
KvvNZhtQeA1UqT7PW+gLi3dHNJFLY/svk0jU1kkfM+NLvRyQF2x1RcuLA/GPrtyoamNbruO5IhHX
IKAQzjaK3VggfboMmh42KC5S9Gc+0kYG+Et+LJEMX0NffWmVlU9iLhsOz2IsgGnDE8c8hug+BmeV
YE2iQv3rhatX6aYOhQWd1Id2Iz6WOs39ubxChJGJTqXy2XmavmXYg7iWkcWXQwMGq9jpOsJ1uTnM
95nis4WEHtz+XEyF3oc4AOeWByG8Codmtb+sIgMjuXIArRyDCzehP4f0dQOTfd27YrqPmHj0NS5/
mIKcjTuJFzoiyYMdLkHtRMIT54HdxWoofmsxKY6axeTqZooXuBu2GPvyMZ37OXiPgBme0tNtlYfr
2JyaPwo0r5MFAljpA3zm/1ohTVALo0Be2fcTXeuHbnojDBEBH53kuG3dY70QPA6GMqGIGdfMeyyZ
ElLuca0p/IXml6j/VKtEiy4Jnq0eyb5KNTblDg7twMswCdaP/da9pXR10hnHlUK11vq9mTGnKFAP
QWOUrGJonFK0O+yVb9kyXoKLJ1U33EssMjMJtZ29SHBbpXGOvb6fw6NSBl32f8hRqgxDNNhoQBNl
qEZN9+TtO7LVoDcuM+uQNTXad6iSEzbgQViR7YZzDSYO9hV3c7la+UIFKR1AdawWiJxANhw3hYQD
2usIb0UogTw6AOeKxvcokwJns8by8CRdEYGFC7o0ZFTOj4eCoVpSspAdHaOYq2IZzhADXGnr/oJ+
SLlEG1PsTvC63CLsy0mIfbGW6WbY03ObY9dcl7v5BydBIeKbtHH3FUp5rZOsTjDRkClcaKPRidnQ
sHYNqXEGVy3PUHnJGRLnBIsRjX0p64hMJQ/VQMMtRAJT1cKfS+c7NWQzNWRZg4YKq8wVBRmiUHf8
VDLLFpTYM31gxTpEmQ36mITQlKG0i7VBG7GOpfTCJoOTVSL+8E9k/tzeRZQpWvH0cYIOG5mEXySL
s8vF4jVBHjO54N5SMiQvwVtsPA3KKEqjVUYDSPPq3wXotI8neDRFLvCspk0/HGCY39sb5G/eLdhE
ZVCGJJHmo0nY/U9DrMItCjynjOR8+n3j3IYa0QOv8A4CGBWV/8UuPCXFjrr241O2+3wCwq8yCrsB
KnqZcyw4Z9Jx0JdYIlEyhe/PuRzv+HmPFY9pD9ifWyj1DeV84zKitPd0R9Sp56h64+R8fLcETnp+
c9+KK3+wWbYXpxlH2+I27yT5y/DYtC1YmCKr587HHGPEOc2y3Vd1sabX+rRj94HI2NAMfElGrNnV
ut1APbxsWhd74ZT+BJG7lSY2qET/mEyTKihPCBknh6S/Ja/MC18x9o4OMmyRk7/5ION2IZB2H06/
y/94ElDglAU1wAiQZztOecOA0q3fWjseru73M6TacsHcg3xTlXSrnSc9rih7Lwi12oaHFQPkHUhY
7zf1Bb9YfNqO6PGCgOAn6VSWNHl7Sd0Wm2q/i63PUd91W8+6LnRE5ee38AYlgUaws2uyITkNtisn
cRbV34DGqmZPuix1zXcElqh3qZJ/VFnuWgP0OZRS84cAioA+/Pi7RNU/PaV/MZSH1wTUHDvRn8bp
YeeVoE2AIvdEpoOcqSzxBIDCUol91UrOjvM+8+RIkJRhc+YGI0fuIRZMCfiFK+To/1J/U3V9cca5
yxNxrkLR130xYkmb81YbXdDxLUapdWNUL4uMZepMA8/IBquZUvcVQyvsaMmLyt2fN4t3VOPkHN9J
5HbxazT2K3PUMn2/lsR1fre4fDg2CVV6pSgpEfrLeIPwONufuK/Z4S5Nr0WlPmMmH0+0StchcAMS
z2LYhAwsAxsWa5NFhNfKYJOJ5F8dC9USz/uDMz1W7F6iDvQETQdoJLtsK23a7fynhKYdn4g+jv+Z
RBawBoPcRPS1UiK7bsxwgBYnzRl8e3X0YI9jbkb2YqyyARJ1WLmxB3HvmM5t+Xvg5ZxPz/v7Bi0m
4r03W9e26hiDM52pL3II4GvuQrUJg0341t9vnwuolhKRKl/gphrG9nlHoHp0GXI+ivBTxeWvWWYQ
zMwEPAgohRk9TwML+hAZO1MLxd8Z5wMt3RDuu+9bI626HMccp3KG4L25+Yndy0ODSjl+f4JFsdAZ
+Z0x5ZAR6BgP0F/5ioE/1Y0xwKZCkq0HdDEeQnCvaPer594t6BqV4ePI2AABbfbgtLY47REMkl0Z
BwUAJt8M6vQgXKkE6Z17YgIoayExau03teABk3+Zqdxa1HFuoqasx2n+ptDRbVwVPqiwPYP+PKSB
1xeWnORLJlzQ/6jTnmZ7DgepstYSakBwOPjByPXKhWK0h8saimbMPjSbiq+/Q7GXv1hdcVS5CAFK
4UI0WNOvy7l2pU97UQ68fB2qJMHlYlPxtiUAJ2tJVB7t3W7nMSWyMuWI3GKf4l+h4kj1SAe1TRQa
DO7AXOLI3xEb3pyiJ3BtuZgd96LWdDVlWctvyGWwdP1N0xfm46hvMO5646qQWyjb2SlqwRj8U7ll
6nnttDA7AD56labBopqW+paKDg7OumC9zo5CqyMugY+GdeciyQERHl3Io+ijygY38zL9NmNxRt1M
3/VtEC8+Qls/3TxeP5iLpsgT+XuftcYHKrvUM2QyNmRvgiLPWvB/oajiZ4bhlLsA2fEBclzf3iN8
AcAbVOg/y3XtW/gN/0B+LZG3Jda8X69YcWVlkCYbKm2Oj4ETMIvIXgd4tHkkGjNonLo1smTLNCdN
DdgEYdljST22EyvDnMdyFQIGLbxQ/oaTG5mbqhv0Vu8/hPhGND8AR1s/3dcZB40emwLNVYO66vL6
3vwIXYImllacV9XFRSVl9IpEmTZwXAs7c2U9tsKnnwOtO2qoOecfuKhoz76/9oKcdyrjFPfPXPVy
fF7wINHH1FqaJJAEuTxZZq77jR3WifNkExc8LMyFSDsrRQqEmanMLfxKQ8Xi+QzaBTPHknRcU8aA
XAVtskbTjC4+O2fT6rUxTHvWgvS9gYkKqQX3w6tpu8agtEQ7Z+hki3Gh9cYJGwm+MXTvalN6JUI/
K6pMgT/0FGSNzHSiIEOWir5o2xQ7cxVboGPhA1SgtNjdVnGr11WQuJ+/jZ/XlhsN80PUhWu+64u/
SNAzh7ELYdZdfynl2oid2SoqVBNysCbq5XdP631QZBER3F22NEyyC8nW1dAgai6QmcHhKxEGdjV3
bFI17zHV1KkABxqInungcascMH2lNyg2NtSNVgP8jubMNVdmDPVbt3o6o0dsiLpcsTtX8vOqnlRx
+Rkg2C2PY0g/qWXP4O8ghINu7fANlb9RmCSy+YO87ZvuxQkQG6NJ1UwPyFzCOQV4u3686amECCjO
bwuckgnmMt+pg4jBPLtPTqwy3cq7QnoDSfrhuxTtcAN7xDYoRqqw0uaMZsybAMo6CnLlqpsFFL8s
01s6vhjm7ncgTQVm7aCscx+kSa990Fqx7piBGMI90Rw9c1QF7JxG2lJWlH+w7CeXJdrD762S5mVJ
E3xAnCQpBll9UQYEaShXBROhWYooVzT3TcJbmmafPg694VUna2/ScDCjaMlXADZCbvcMUTNe3oX9
M/U/B8XEXemAdfCKwCKbBcqia90V97RRvMdAx+o69YW1TWFdWxPHQs5aAAWcn1nuzvrGLwRNqmjQ
bkE+7FEm82EFPhWaFhSKWtBqS9JIhF5eplOccFt7RgWjv+JzrEAnoGEOPzBzEMUA8eStx+rA6eCK
2eAHeBi3GtchdTIYC51O4cT5oQO1LUXi0RoVUivV2OnQupQy2OafGhqJjWMbeLgjZdtbEnREQwNi
NDQaRfXy4pGZEeGdtH+4uVx9PVtUhSD++ZOVDsx4WWZbuzN7mJzOZKQUsWWOc87SmMCw6hRJnGu3
2w59sJX7MvvQPrUG5YlShxXwUzeAB5QlBpjG7s9APkGyrl88eU7hAkxGQkM+Jux278higGCG2/Vf
mdkbRannptpjN9IJLdYLekUd9xPTpUjJEALXA2Uvy99gSys/kE5OeJUveZWiealDGEwdanldZxnR
NEDIB1KL28sPKyGhSNXlRT0sAAzUdlAOpCn4VPE9ZctUhOUMSjfiS5s6pkwLPga/19uMumYn7x03
7gNZ8kOeccffkduOLVi1mLVczxeb4V6eyeUYB9Pzv9sVbRa42j0+klZRMjd6FZm9YkvnBqAmp0IT
5S3JAzBNW+dv4CPYc1HYBaUGDZWSq2w5crHkLpB6fnXtqu4JpYPol+Utg8C6hbtar3oFWtG3Z3We
2UCAF+cqU4x51lP4s1aDXxzwsWnIj53RkBgh1+GiME0QSQxKRfu9mhNLvxwz2MdzTCtohslunsRR
Xmw2eFYYho0VXs1BTHgKSJ+NgpIoncltDQx0qDg/crhWGbqg0DTp0eq+0cgFBLPZe82NfK0deGD6
oHvxPNRDIi8WabibO/A2t5a8G8Ot/db3IkKXKzuFNyumDmQ91SEohX7P/ZhdM28DX/JIeQNK3roa
vO+Mm2bxdOgf5/bLmeNW5d84gXkDilsxvIPSSeGCyJkKevZM11/+Nd0pOT6BziW0Bjw6d1wzqweo
DVLOEn+BuL/u1r4GMPKcqEjpMV4N8pd3tXJrPi+4Hj6yFvPpXq/imuz251p0u0d+KyQQmja4FBDe
nLrvtmYY2X+GfOUQPcie/7c0ckXOAWXkCVl+5N959lttRcKanWRclv3uPF6umAKKciBxlEr0Kg+9
maJSTNOLsYcg1FAS/DFaL261C/n71D/zeVU2fEn9wEUEIIoNzxfiYA8n9GQet2znRMOYw6LEiIuJ
nmMJnmovhdtBy/qYO6QjcFD7JnVm+QmxQLc+057dpdmnjVIg21yJvas8PfQDYK1nleWldH2Ew2UI
wa9Xu0+iEKa+1rSj63uDPFRZGD8pXYved5cvPG9g074+rDducf0MJvSq0qJDs80cE7pVgnmFHiwl
t96ATkRmtF1Odl5gwkM390NupWSbHPfkcBoh9Vz2vJIP7ZArTlQhFRE17nwdFdYzWshbUODTzMvS
CXfGrvy9LTzCkhYA7sfbIZSBI16g5I+5Se4C3DkNOiG4Y6Qc2bdPPnTEqCGGcnzrN3B2lD2kMEpq
VG4LqsDyKX1beySZwx8sXp5WZOoQ2X04q0QboAa6l0QinDzzq0uM9hVVZkYtGFENcnjDhyTPnB2r
B94C4FraHRccVQDSCMJB8ABXbnVjNKTsI/Y3tnvvlcE6+pC4zyo92TaOGws0+uNwm4t7QCdumFle
PBPSX87ieEn35tjpFJoQuYIQIS3iYqWXzAPA6iCK/q2OZ8EBZim5v/PQFKEFdXmvia6S3r8HEWU+
aiLhWoN2lrNVxLnNkDKS0dTrlwEBamQ/lxlemal1iHoMiI9saIYlofqdJ7MZmIdeC48gdbaoBDmJ
lYHHI5/Pk1VmgMKXbmgXu4GIGKkbKlAaNprBiypQzC0xyRnk8PXgmhOHIGSxgwBEjG8JrxsARMLj
o3xsGFdHfHrwhBbDVZAH8a1mKxiwOftYFNsAYsaGR6WUS7YwUvQX9EMmkDtDatwu6mP1Ik22QVXf
+UuvwPGWkNoKYRcpU1DRnPJRXzOjSdCsiIjbeB6oFmnCL2xZUsfO5AqmuT4lGqEey91B7MoN8knV
eyrQuCrQHnHnK2zo9rr5xqn944LyO8vuj8rrdLnf7UF55nvPl6q7kQWrQDnmEq9lNT+KHsn4moZx
OACjv+cZV8ClPSML01RbFOqnD0vnLzncHYR3ahBkUoGlR+Wsh0Ps5sJ7uL4EYjFKuURo6+sNF8Lh
fYxMIrrj7/WX7qXwOpLRTHccDDmPOYPyJcQleINSyz2r3TX5A8KCtlfqVFrVh0y7xbmckVQcmt0v
RFr4oSW/X0+wD0CLQZxLMRcXzRPtFdwluKf14dUDL1oE/GOuQlRE9/rYPtIavm+/oHw9Lvm/h33X
aQoE+CjToXPyYLZrt5QZjpTypMuv5+2Tx+WP8gFiNicZTHjRUN60HklLwQZeR0v3fLsfxkkvSbsU
/nyYIFQGza8mnAmmHBqYmVUuqZTYXHBObidaO57zoAIPrFGgBE7Ju45PuLn6wT5YPDbZQdD+nAqq
NOpDb8UJHl+d+hhX2mFY/PPG02FrkUP12QlH3SymcGEYVoKgWE1SR1p3SEFaOCjF17pCopKaHBvl
TXwyShnEOAvf+dVUR+jbDucwhRMlaIBPnZwXZxH+mAsq8fjBglzmYcGgMOellAGadZMEcrHIEEFH
B3HPSPZ/SFcMU9gLJ3ekyV8MqiG8KcDe8l7b04OwcD6v8kS+/sXXFzIjRCPaXosfv2uBbGrB0xz9
Zz1XQuTmSnuQFNodZ51yKGFYSeAs0hqxhtcWC0kC3QnRQX2Enbc3/ORM8/r3mpysp1bwyDqZjhFB
kxjyiHj0YOAdqGFqlDDiSWHQgI1jp50yDSH60HvctmgqPx094wzVQf+do2fMx5YO2Dc1x9yT92dh
tkFARcPBspNSF/ejHThJt+INXaiXudWb8iXlEFsyFGmu129YX2QY/gjxeY4CglopJBbMqpyMPir3
bhP7C2gBIcfvyKJpz6rj5pT4BSFSvP3J4ZWg+JFQTALZlbYKN+YlRoQSByKE7J6JkV2Ms7CzDrRd
ffW0mla2iPRgiW0GcGEdIhAKxCkK6pI+IifbG+MqxPCI98lPBthHCu220OPHwgs6GG3lo8cseRi+
kjJBk3X7wIbmz3zLgfxTyz+QMlyXAF9vG6FnWFQP7Ad93+D1ZikWU1vxxQrNzuMHe3Haf1pbp9/9
n5MLNRLvC7OanEebC0Y+NiAYr4qRfYAYD+fVglIWuZtJEAVHa66GWxkyIjOSPUnoxHmTFAV2bSUU
3JZXvHU5FaGaTXt9Qj90+Q1PRkTfXKx5TcuoTSI3g3d0fF/G3FhGuVOTZuOP2mU3kZ6SLEdxA11a
p3UYfwo+ec/XmwdcIU/Wx0HZ9ccAcbfajFy2RS7qukDqsdL2pgmc1cxvdX4ZuzE6SyLu2q5gaJka
eneHFhIsLkx/2RgfHzLZMx970K/puUbtI5WQoc78vi9eIxALf0nvUoHTjiFQnBvnq0qQlOFksRvV
ALgmiFDwCug2TdJojTsX643pvg/icjEhQ2QVU+1O9xyQpOJpg8bcqZHJdIgPWC/gEYZfaoHnNl3i
poh/Cu8F6na0GyLUgjnMaCMJaLQZ/ZmY8fwYProRP9I8xNU3XZUjHDiw4nAfipiX1MGpU80YALh0
8diuhNTWusrv5SxMZTqoMI/g5SETLeWtO9kXdlGuZdI2f4gOaCNlWFBNtRXRTDxWfLh1PqKgzacS
7ZukR6s0v6UsWzADqJhMX4ytxmcnFst+VCKVeRHaaH2+odvrxBsSOLEXQ3ni6Bv+bf05C2QUkQvw
yX0lTpUx7D2ytK2cSlIMzvAX4p1fTQfr32X0ebbNF98pORBWjfTVZNgzwPhVNDvwNzUqVvmGL15/
rrIRo65EdBSsWSTfisJcLazKlLYah9hRSOKUitNFEP38zAmMdpLFCDsMNKEiLR+T3txZRVOOXlsb
vefbhzfwacEqdD1SqswPUfsmYOsG/3K3WRjxMRZ3j/mV045UvQdSgiKKRhMyuzC+0tJoTD578X5b
D0dvB0DTShhW4IRW8yo9lN+fm/jejtPxfU1UA/2PWM8Zh2CV9QdtHK5R8LyeJQv7elFDXrYkMUXe
gLaqSki9TgfmzdI5/BBSwFwYSyRUKVIgsAISIvEXB4uoSzdlB6Icu9MPOEDaMjBoxX5BlfimNg8x
oqz4hY+W3PIW74wI2wIH5Xq4Y3+z/d+NLz2AhIvcrnz5zNNBvOoW8BzzABi6c0fNcK800rSQRutt
F9piqDaePXyZTNan+Dqqtu+v3K71URw0Y4ya9fjDNv1wILKLmg+a0MzliLgjZwFbWZFDLGX1n/AN
aSsK4sKB2/YQlKABVLdzfMfIDxZ9L05B3G7w9XG4Y76lAVk8bF9iWkEFNFZGQWme4FKEvhrAYXH0
O9ke+/tLWlztg6Nmcszh37rq+67/rkZt4IsnmzmKhdnKz/hGlxSn5w1G8S0WHsOOaOV+ntrRXxrO
4qoMq6+AGoYS9+z24V2YPPwYRXEBqDJkRmE4/Besm9GHd/MqNIMATcO8+hfgXWSbFnWzb49N8nXh
E99M1Eu9x8BR7doYFQxA8nxnE2EaIQnh5WYp5V9G0oa+Om3UeszoK7m64RvCLKTCrkC1id00wbCl
tpoBBRb0sSuXoQzIY4ztI7Bu5mWoUwrXvF61nHOX2GupzutOIoJKlgmUTPFAi8cJxmllvZl0zzm6
x0zdtzYDAdO/n/WA87VobKZuySUYmLHUUC1fj0OcllcYVFl5GWBI9HzLa5RTJ1BHSBMDZz2zmmPS
okxIwtXPwMJ9L+0FRA1Vu/noeL0UNH+6JAStRCmaBMQDrNhrbUqUDTMv2ahYsLarqWwB+J0Jxxpi
tlgeumFh1hgIGlW8FYUaSXv8LfcU3YpJJdmOqs9DiJvNxo02NbVSnsbNmwbkwqM47CrR4ZgRzFC0
QaX0a5rF2lA/4h8/eWvfIYNqhD7n+Bket7jy/DVS3OcSk+AhLr5P5YGmJ+DpE6KySt2CdvITWmhP
tsus5l0Bwd6gZQGPQpw7ba0gF0+cagRV9oAdjbE48V87SX1FNt1TukD1Nvi9zaKoLYqLSJ7urImX
tJbtF1B1rBhlMIIdmz2XUQm4F7gIwxJJM/dkZ4S/2KfJ4afyEpeyjmbA4dd4GmCUHstKo1oEEtHr
ql0kHKPSlg38+4XfYGI6UY+W+p4Qvwz7y0WEYZ8MbyAOskuHLUk5NH8AoggjCoVyDHeHJKgRVCOZ
AU72rENpNKIt3rQZkKVX2dx4OnALr1J4Qe1w2jxfDMjhq4A/1uzwZX3YFMlNmZyaZjYyLmsGnMwd
fhLS8pI2hXnx6LLebRdpvXJxKNYX6kU4ttAHnbpQBQBcz4wtHq6mYbyIXlzA0cy9NvP03P3ao60F
wbhI1kzVp8TLTPF0InLDZktp3IM91zXlJ1KPzRh1LpSlprfC/xKEoDLLresjVPn66+GuqyrgLdJJ
b5nCRGDNfd1JDmGHaZSVhcqHjoxJXJNHmUHUGyE7o9dAlbEfLNbbc5eAiCpTNpRa/yGHn/h0Ba0p
L6phg0PdGLxSxp8y4UVWvCE6a8zEIC1VI9fhX7QWX1BjGl4y509XIH6WhhnAcDhvUbvJvEC9lvKZ
IZjzJMGzp1N1O1DZ/65jjFpNIsT1lX8B7kr8xez9bb9BBZFIhVSlx19b0UIKThEPym9Cqw42ZBKC
61ZfpBsKOzKWMItmA5pbS4L3+xt3B4bMPGW0i/8CejsnIQnv/P2A5HVRG8ny9oDYqXtVZgCU+3mx
oat+l8OWTloAgnyiggU6V6reoY1mmduX+d5jUPw5m1vlTFbHIOBJ1gCC3Ce6/V6uM5r1TBqn43xx
F8/yZ9N2T5u5luRJYaxLQW66Vf4VLEWQAK+loKiXf32V7nppG9Vqd0MTZoMnQP/z5gB4ggyjJwHK
B7TfX6DSu3g6wujzRV6iW3DUGpCiDTrk46PBmxVJL0XM5E7PAzM8wNxGvbqmlrz1m4kuY8L9q9Wo
+PfPuK4kK0dY3weA6X73tYLhK0y/DIjesj7o9dNd3zvv8Fn+Pl7XyX2Do5DFcC+PrCNzOsbf3PLp
hq6Q/YmdCiHnTh06WQLh6aOLZJeQfB+CHazcxASfRMWFrYolCYU9mxd2qZWAoOB6yK1gU9zkUR8z
e46QTtVEPl/jbHPSPuAL+msEbiZ0yXuppsRrRxqRBq3jn0cs/1lI6iX+xQ4mVLdz2SLi73jfIx+2
D0tA0U2MBaFCwGaJ8B/+ywaE7ycwYkkRc6ZteOi8FeANEkSvXikip8zkhnJn7LXV5X/2gukEUab1
FN43TNLBML8g/aWyq9BnKxR9xZWGy8HqESWS+yJ4/5r61mv288ea/0jtWfL1px/K02jD1sAzT4br
cOrtXPB/YpigIBR2VnBPXBbF7Z8yzy2RTT3kTBBj6HfZWcdBbudQDf/F8/D7C1ldq1RQk6CiVL+T
HAeROOSj1N0fDMAWO6mDd6YLVhHVANiAm+yrY7muIkg9N32Iv3j5Xit2OP6iwLXWXG4QjoOTvDhR
GixTU+QT6hkdfBd5yDxZchTiJwk4Yrw29Vt3YoO/O22dMYQYvpg8WxD/qSHhHW+GP5wLsqbmn6gN
gXJKUDu2YyEhdjWtX769+iOLPGZ8fpr/lzdebn/m+G/3KHrC/J52/wGWjOpg0WTFLyFY7A0MDvkn
giEwvL0JL1rmrM1++zmKPg22tRNT8IvyDJurcaz7sFYGc4JMY4EpTJh6LDKW+YA/pqnBAmCUoqQ4
bRIjy3Ma3HJ8DuGTMhl6cB6qLKxAAfq0HHdB1RcsNdF/16p2epuqdtk+b2R2nb+1qE+EzR/qGY+y
jH4FFEYp2vBNOjsARB5jBrnG+SJK5fOq6HvoyzElaJR+aFXhnY2D/QMh+te/6+DD6GFbIdHlsQIF
iFKlknS6XrfQsU4q8qEMwh9kZQNY8wIbghVDB8Dd+0VADw3+K08F6SKCIbazX7tHzvA1gDPjn0V4
VNoxULcxeozu4EZq8KR9GF8CZDYAeqom/1228QVvAHMe7hJXuoG9RFFLpxtDEUi+WBZxCHBx8tFi
A0v4m2W27MhxyUXAr+qAz0HMO9Xgm7AQ1yPFeKdvY5vNHZoFNxXDff3ebv39W2vXd/7v8LiCnedn
z1HuEOkqIxAspVmZfxhbHQMpS10t7WSdFKk/+U2fPgRlL0V8Bgl7lC46aF2D6TFWFVAmu2c+0cMG
3jVbwu5LVAsNEizB1F/furT/NdIWFokev6awaLdKT314WuGP1B2iouxe8Yhyz9XBvyTsU928yflj
GaIOUz3atbStNTWhNqHuIbQn3KTjAMIFFe7Z8SZAheuV4RwM9nbYKdhbEdFvvV9A8LujRqVZwMpR
6PLz2EV1hNy1UvOW0ZK0/7ciJacQWZVsXG/iuFadCpvUdoj8fh/feBlBtTkk+TyXJ0VvD/KYGeM3
o14e/v83rWCisItJlcv0LVKUhHBLs9fgeRz+L4pxbeqU9aSqTNQRLS+c5SUqyMMMsewpjXCDxbtc
Mn2THX0wYbJjdtg4QhKy5AtVrhXMvW59zdH3A4YYpm68UO9UYe9V4mQKbG6Qk2tiizcV41rPCyb/
80fWai0YTrq3C5F5m6G0S4So5UQ5EyLLUzcQv3pknF6uiUCUeSjzfl5iiEOG9oWQ9E3vAAnxj/+q
tCCMxIgR3OOOsPMaPsAKPQuzJ2jsjOxYfsh0Uhw7HQaz/bb4y4Y25W11sEt6Cv5Rh6Sp3MqSP2vI
wk8huO9/0MgkeW6CnUsQjYWnL17K+XZ8op9t1248gDRNw4dch6ZFrVm9tw66SqOHfdNjzSRdCf8r
WB1TRfOh+VFjS5TwhIBRbnUXWxvhwZ3nV5pckwbzLwe8OioKluAnOtuc2wEOB2s10NYrAKOfpCQq
xgq6mO5DG9k+fhvCSUewFfBT94H4dyQEf2TxfD9tVOk4tcv2/aEf+/1SbqX8LtbDG5CGRMlR7YvR
ZiHAIeFqUHE1R+BIpMuPTeLjyOGHLGkhRlSVT4OKPiolEtijyboHEiBDuA3XLQqbV/BeTxQKLiHM
8S512ijR4SsZVqfi+k2L1wxYtVKxv9SctL5SBeOtfV4hX5hlSDoUI/ksT3CXxERc20Ni/wRGro9L
wnUe5R4sSfNQAqqpxGEi8TbtjdOzTy5ztt207DZ5senZBk3vYDoFmegpOaoprIdnmaNsDbyuikmq
6pCJOcfiYr3IeQ01yYhVVV8/nd34l2njUAzj3y6KnBAxTLTdDR6j5OrxO0xoxnCltyyjlctvjqOU
sYO9aTWlXIeX14MmpMKJwiJHJ78+NUsOxc+vW0u9kKH1ScMG55N5bjzxVRw32ikZ93umAJ4D+1yU
QugZqvF3uh6FWKYh+De0LdBOubuymPcrvC28OACTzyUr4eXY78KN33L5PqaLNUPMGfnE+uIYPyPb
YTnYgs0WTE8TT3ghoAkaGzGcFchQV1ALY2H8PEN9scEhyuCR3s88g2ysnsKyKsaeJwCgtzu5nthC
8MRT45gin85EX6G7wnnMUXVzRnlR7t3To1ys1nSgQdMPZxQchaetFxrh6kwKMvoN7/VyCnOID2II
sS6CvWz+6hMloR4fiE22gNqL+6lrw4ElW7+AAvhmhS7h+1XUTG4zHjb5aY820p6q9EK6JUThu2hJ
8NsqPYrRXhxenJ2T6T8ybv+odqEgdcwbvrz/xxO1Z+HVONpi/2qwY8BFGVLfeNiQ3xkPc0lqcUYH
FCSZKg6MG6xPrC9Lg3UXQ/xPFVZsLINariMRFaZvo0N7jUnNEiRu4yeWyW8mbcibBsIzK69INI5W
JxDLygiWTvJSw4muqgRlsBPhO/39vRpInBHA+AanUH6G7iiq6bGSqH+hsaPhqYc4f2t8lj6JDHry
XyDo4NjnR2z4+IE45EGtCPKpw476LUv/LD2nxSOjUySIWwF/Y/0PLLYNFRWfhtZP/98qY4BweKAQ
45F4UOtykz4CNX9BrO+gta1TwLnV0HhtVvz6fzkJ5PP487bgnDxeiMSEyCdDl/XU7nF/YO/ACS2t
/xc8MVfbWJctJQVtKG3Bzq3NVcRf1GTtIMSa6OjxLOCKvwCcxJyC0XwVnRzdrJtyauUo8k6L7xjj
NrwrT2w4tVID5FggcqscTsXQWr6e4AHNMwgt136ZonC5ypJ2BNPKHEKjse75BOioQMqFkjqEdqKA
hgrSXkwDrb/upP0QDVuDKCCV0QeUuAscXL2VsTM+pUD0LCmwcauK6EqsVC2tAdysF6/q7uwMcE2u
xif/gHIe+2S4GmnTV0DX5Z01zSKXmotsJvaDfTQUGKB0LF3GpvBSyFtQN9OXGVGVkYzgtKtH+yEE
bqdYD0jr9jsBcT2HxUZWJ+kjNHJgDiweqR4bqIZj4o9JO4+TcL+G2l2QN5xpW8vAfnHuTRUUB3lx
UY3pKiYINpo1FXG1D2aPpwMbSrQFZZIvG/u49iBLAPDc34BaBk0BZbV25f3Pnpk/lQ2PSx/ccGqJ
R0RtaQc8y0WyeWwfYdnAtUJs5fDy7ml1dGICT0YcJevG4d1DxP2Fu5BGI6G0Sfo+8P493YFZATtJ
FGFhxsQH/18gLoKvTpg1XYsxcVAlwajY5OBqAs6ZoYltq6ekZGo9HOaTdag2JfjgRw2nY6OieYVs
Jbr98Qi2Ef7jKN8Te4jlsH9pLaQPetu9kbkhY7IuV/Nr3U6gu7JN4k9Ylc3/5Mfo0cheopI3xmb2
sn9E0Oi/ktZO3pMF7YaC1xXotnvsWbg/ghsJjGB/LWwsrsBX/U6kAt5x3s+B4IdKIziC4Gq1b/30
KiE4A6oQkHOgQGmDXr5sYOp3hHYoWKE/Kd0abJZ2jWSNLs5dIbqLI0fkmC9TF0JMa+TlylmpE9Wu
xDRllV/KtYiY9oQs90oPQdDMgAi9NpmcCyLpJHO73KqJyLZOIfjVMJmq6izcr/AdbZ7ShrZp+6Hu
3PWbpGLKq5Nu3cKWY8g9zOqGkAyOFG1nWI0vc6k44HzS68t1cPrJsM1LkX39nZk/cSlLGUP7FQGt
X8XJeiZJEaAtw7vdhv9efqGWTxBrDJUJ19vCtConSxaMRjRuxDW0Y8L/NXsBP/XbqZNufyJKbZQN
pIKNB672BWOMP0h/gJ1jXnaXxDMkSjAUU7YiV+HDOPt3eCgj5F7i3YNlymXZXQZHzCsza16vuGqz
3FhH0F+UpsX9MKu/90mdtKsU8ubION4nak3/ibcV2aoJo1rMc44sGLjZVhNFrBZcZzFO4hHIb8Fh
nrgR/N7c5RZQ0/CI09WB4HWXtkQ5iuTQ+dBtMhmcCtqOKRFtkbLD5JA8weg++80MBn3KynliNlVI
rMFQ8OnAZQuQDB1Nn1yeiz+nXb5yaR+JcHrhiTXEeQpIrgMJNHbZaiO2oqq8rG5hRM5QrLyigYWe
tv0irGWWwLVoxB6xHXDng0cPd13/y74rRuSzRkXHjSyYoI9LcBq/86yEsyfIVm6XBgo9otDTWyxf
n8IWv4m38TuITnP/EcphH90IeMXHlm3ErUKKfazwF6+W+pAJXtCIxtLoRs4ErFtR/BENNBavUTLP
xX+Y/9Oq1gzXrvQcOLhJPYgUF/x+cICbMKyMKouuN/gY50QwjkuolV4T9/nmNCjmbsUbsIjZcoCh
T1kgonw0sAM2hlr1//VmRda1jBMtHBPEqteOME9Uu0NbJh2afpaFHLKRfyhim8u/mT7wnj1oBsp8
THIPSNzyntHREf5QJgZ4vtwPksXmIdI4OEZR7275E8ws0Vy6qUtv+rsit2p7/nBQ1Izc7WHwgZtF
wtirP8p5XQR8V1J35w1GlxRz8zlY6YQbwNbaEeEHGTOcwzmyll3qhFXrgG0pj1DW5puWyzxB1x6N
P0GvPmXQRw4XMwkM879YV4uKeTpVTJzV7q97KGTrkOAc+1HWDt47H39z59PdrbdohVSkeowRX3hR
dbwdgGxcYB4enSSc5f3oeNGkMjcqO+ZiAww9m5ZC/DifRXRvxEVp7jzZwu2walUAL9qioTwO6kJh
XUuufPJpK7d/vFcv9ZnSjMzuHfVCkLJ30ZVhDkKjVXH2G64faB5lLK4gxkvxJZ2ecPyN8g1kmptj
+C0GfWaEgMwoPhx/RV0Ui1zL4bHmQ5JfQRnhv0F+8IYRQO0fMtOmyZVQne7vCQTeRm5IPmvEGCZV
R0yfc8WeRk4oUXb9Oo9BSTOpjpEYL9wF1iLg9PawY02mns2aWo3UnAYV6uExqkC1CT40PMj1mAq5
tMKFXUlYNxoTibd+/pj9PW5ck5Kg44WF94CgIwXQzNT7Ontqg4gz2qiSs+LZzyuMt/iTu7xY9g+u
A521YLnqOYAtAUwzVGPmJT5eLzz4Qmc7e3lzxS6u7oL1klVsUOe1lnkV20F/0yLFB2H2g2CymKX6
LeYH71QEIuc0596XAg76I7HRP/6eQRbNHj8TzGNo+TQjnPCVQ/PXl1ZJuXV8+2QhVyGnyLciZjjT
kCnGEHwnCUzIt/mGWLOBSR2xm9LMfB7uZfqeUp1++b0L3OERsHjpWQjM5rm1IvtEJBJvgEyizON7
hDQpHMqyRQJOcbExONAqqGtdaU/ijlf4+FZr60EA1ZWG6Ji92lLN+Y+bbRx4FkAkZr4SuD8/lWkV
7WbH+SB3mvqyRWvScGg55m2coyUx1/rZIbvKVMQXWkJj9Dd8bnLiNVe6kdWQ5p0TdXTcr4mC2srI
VO4fAI0Hy3jnsNHVhJ6H1ZFC33TPJ2MtOVhsIa3TYyEpxqnYcfDbjZVSZafsrCWnaZ3KEZH8FUoR
mE+IcDb9lr53EG91hy9XnJnGcp8ZzSxfhPu45RPDP1CWUcPTYww0v+KP2kCW256sIkwqnZuoBacf
s1wfT56PqYtP8BZ6V/ezspGtUXouj6PEa2LiFEugUJ4HTIZzvMlsid4rqyET5QfExAHutLSDa448
izcSypGrZIebipCO6eUDb8acKEjPg21x5YEBAHmp095QITzRC6KCRClt8k2U7p1OmABAVCqwmexl
rpyRm3HsanSL1nHV6VAtTi3tQagUqv3b4d8FI1KHuJlyhJEPr0IQTBIosfNIMWi/2nd85cXS/zip
q6hkmNFnkvBMPYR70T+oF5A6pWoBFvdqiWDgrIabDqSC6RK7dCeBgzjWPZfC/QS8yj1ttgwXOCVw
OxXEEWihi0KheMDDoKDpcRcupTruaRXiKCPY9g13q9lxcUlhDca36ZlbZjh6slkJ+3AvJD9stlzv
OBhD7DcrVxyEBVfbik9ERSapxzy0x33N7PJ0RiWHylLAktpd+C/mpQcs5VAH+++bFnqZpUlVIw/G
9Cz0Irzx19WfqWLNSpLYVQP4RnhjNwVGvscFtCB2VKRQyeR4xyBz84fJej/pjdnupA9eOVqX2CfP
hm5HpImVKopygvKtAFGqy/E0nTK0YA6LDufCvOhbc2A7iCNDzJ+uznGMQNoqIFAfxCl+64sK4Rjk
ytG8hMEIeymN9EhtUqt0I78XHJjxbMI2M7p2OzmwylCYkIvVgraqmGW3gYC5g8TFDegkiodHfWdb
T1/HBGXUyhowYt6P8K2Mdp1eDPN8B4tJ0KqLeOFZOMOBanHVbjRiV32ytjwBJuoo6Rv0LMb1n8Ys
YJ3kYn2QQbKbvO2iB1saSrRcAAKx3y9JhFVZ7LYTl7BkkZbZfDxQBIZ6sEOn1V4Bl+2h0eyirsLe
yveIdZdgg1dnQp5E+Abo6DzXAHZHu05CgpGeatLEf1Zyd7IpeRfkT8esKmkkmTDLJU5kB3iuLlmZ
kP+fTlQzGyRT65JkWVb2hZX00ct7t9TtRjVY34zmsfxg41OsjRU4mGC5gwpE/VY/Q1rrg5G19/zx
CDRHQtO3hVhp3H2z+zF7XiXLX7AUvvsy1ut95QlZtvvOhpc5Gk7Ots9byDCc6GUqU+/JJUpheAMk
fO6Dcl7FTtdTJkFLCNGdSAkINEw+T+4J3ku0jV0wL9x7hhjDgQgzdXv4u0Xx/C/og8GxohIMSteQ
wT6nYzY38CP4HbkkU3SoPWmpeg+YyKRsKVRueJu/n3HA6JKgz++AKmO06ZEl+G97Ciyx6Txn2z3m
YG6joUP1+9tvNDJDAIZCKfoZPH85IqjFQX5u3lsZKFcspFGk6i8LLh96l26AU2n1ncHfdAk5z5tB
3TviB9EXD6XT/efnA5LqRVZDUqX8D8RxDW7g12D8cG+8nB6aFzlFCJ87JZVKIf27DlBEeR4UJff6
XEE2JA9omKUCfIsENCB2Aiz7iOzlLJo56Sfl6/L80mFoH7V8CsCvtZL31DFTsVN9snwj+96h//Vq
x/8AjNBvdRRSIDHS5QgGQzDkH2vVjerb/DztmcEo8mE49lpjJv58tzn1Wh5nDot5WUE5ZAUS1uC3
nuysvrpTKVPUaOvfa3FgAcSxIaXACDw3fji/BJGHjV75OGK5mkviLPDC7vCKEGCEBx5WgQKxV1Kp
xDgP5YHBTXo0rX96Pug7dJNSxheZLwADhEISEg4T2nm0wVHncikUkLgokuZ5SpMi/CadqsDUvpiU
DeJv/npfnpY7EocC7ZexQ4ab+VbFG07XJ/AeCGbYzaAnxaiZPHqB/xohEBeXUmbPoraPPaXzSFDO
NYWgZ5o6NfngVR6EC+6MgbMfPpbvA0kwSFswB2LVLnR4h5IHR9evtXnezGyAOKhRcfUrodrkEOej
hvPBtOLz9Q76cGQTtxwslHe7sNHDZJlDgbezCIR89MD5cVy/kb5A5cJJi7F7QlPfJ8I9YR/08Vk7
LWhxkZo0+K5HfGMqSHgzDnxETjUHQ/ee7Rqna8FQsNn3TM2l+kv/8wzSFIPSsGYcEUIXvnHi4ovI
N++jSJtJPZ3mRF8m7o5xEm3Zxi5psj7GCLpYOHHcW4b6lxdVdNdQQ8x/P78yITOVRyzbZ/ghTrDG
4ey38IksNd2b6eIi6zkm8M7vfmvet3Uq5Pr8XOstG92z6cbe9nBuGbMLfSX120wshwUv2u84fdy7
fg2PCPii6RwQpc7H89uiL9ZtVVNt9XsK3vFa8v6fe6fKzJTfZqyxBNY40kVZjTi6cC6NlGxdYHqV
S69SkMaayTlybKQIMsY0DPFCPqAYFFeTzFKJJqcaBoHXD+RWcmUQtmkRZnQLhmKpcEVMhMRixIxY
8SiXPFQGJUGKqrj1xXnH55AlvnYxtBjCw0D9R99ZvqgDXrQXLqj2jebXKkqyNy5MAwKOyFAn9X9k
cUQ6/0cVtsW7wJMPPe7iYW/GXbsVZYke76M116BrP77Kyq39cegZRlSeZTi2dDZjMwuPkWgw+JDZ
LnYLmxoU7eL8b6vUMgpo9UJtI9df2gd17gEtqVQ/9W2C+we073XcRALYtMlZHeozljVLrR5xzHpc
JnFckRFuxxLWPTVmwJtMpZj/ydhEzSqfDOUU/wD5AD/MsFFm8lR8I+e1AI+5Inpb4tUTLzFyr3kH
JLNBR3NKlzDRSJvx/9rp+eBzWNaKkkPFMaIQgRmsQr1jUAZ3ZIWVhA9eNpSSNYSTWGoM+oVoev5N
wNnWmt4PxkQB91ofRrbcyq4g//aJLZaje0hZ9zo8/zLFJGMhWEQ+O5gZB+wGvoEkileFL7iwdMam
xq6YS0hbCg9w2qI7Tjjane844Z3K+LQAbCooVyNR0gMnb3bTubVWW6UhB6TnxjcWndaR9D+7V41l
AjgG+CQ3UThfYj+uDtuhtLCR6A9ipPqw4ayOi0EqPNvYs9QT89x7VBMYSgbclPbNENHwpDicMgoL
Sh4YLRGViP5hBKUnxz5ga17zWuFtRRSep0TeRW0zZaX/ThjQ3vnWvBptvTVrPuuAIP7YWZk6uoch
D7mT1QRUQpLEMySCqIdouFUicUaCVeDDG7L09ulpafaRNQGhvhEQPdT1q3qOzWWuYFDL95QXVZyy
Ns39cqS751EzlOwy140ddMLTHirBUbL9+NlLLcy9c+W7Cd+deEOHMQkgevliN4l4Yjj4a3M3i6u/
QLHQauVfsd48/zHBIbm0DK5gwc608HHYErM6NleeRBBZ8Y5BWkZ3CL83HRMYxLXlI5u3ZU4djASg
ZujR6FDIToJmjROL6ggUvPM/ZnqmhPk5WZiko6Vh19cx2IGPMGAvVzhkyYVqZE6ukkZkXzAxx3ps
y9zDbw0TEgDWg6QRp5ydk0VkHYYuoM4THu5LpOgT4IyIRBn/KyWTQ5Wpu9Y9S+2wqOVgw6iGNPKj
+c1Yz7H38JqpeBEDM3T85iZGz7YPrDwfl3p5N4F3nBXawhDjNP0wesEDJ2wELNuUGhHARytS1AnO
aryyLTW+yDUZAJE2ge09D/BMYFu09KYj0GECv++Ysx/9+B5ARC8BYJyNaVJv/qKQohkuioMyfW9I
svtGU1FQ8CtnPRzXeSgd+DU08844q2fVhr2LHud0QcRlCevz6c3qnNYTItecIiZY1kT5FeNQYfhL
TJ7Xw7X+xnY/n7CIBK2xSE2cPXEWUjFTaztA8gPsiNu/cYRtvIMHpnXCLX+VjZB4mS6ujmM0nm5u
G9SuvOqhW1NlRUXCVppOdLYPBZCY85nCqHet2XENQfGY6BA4VbFyHaIWhix8kZTtyYhPceh6umgW
3ZumouNMaF4BCy2/fKpOvUubMDJH0sjbYOgJXG5Bcrcd/2kzgi3aVVfNkH7DcSqgO06D6Aozl+98
3OFfJXR8iAjcaVrLtwmqrdOZqokjObHcXxFsVKYxDOE5mS50zznT9KTdJe/g2anrahqnnuUx3nHx
tbdLAD2EibbSCR2kJuYSaDCXjfpIxZf4LN7NCWD6GeDHaIE+Aht3SRgg3T36lZo6ouetjD2PL8k/
65B3ed4M/MULSeGHGmTu0+lhKaPMFTUh9nMpv15Q9bwv/EnS5hl74BvuI/+x5ABYIU2NFkjS9n3A
JPO6+iCXJ0tufAoDjIPT9iSzoghXdWhXNxSqYLEpx+xkCMyXa784CZJ03reZnhjo7gtAXX27FS3c
JbPsBSXsLkMIc4Bj2TTZjfmlBvMsf8nnqpfqRDnPE/yf9MbUQrgnLSrggL38cQPMViHgL5HqoXon
AHVMEtwroZNFxJ7UamDflSbV3FGVLUqkurfTkdwJOf55XAXkgDNX//O0/G78b0Tg5RjWyW10Kx4Z
XXqf9vS9UJeCCdfsICPgCv+bkACWTW0s7bpnfZk2xTSgBWKISw92+Ml1MMPNNIEfyR9l5tIhPLzo
z9OMp+qnt8xXDfF/uMHSlphbl11ikPDKQEI6kAPm27EaI9AUGDbIaBBmmG47jt+EbqWWQRcG2QNZ
lj9qPQuz4n9wWx1FEFnggHPYCs6muqKfFPtAyWSGa+bA1fSyW0Iph0XZtzyz8mBjx7/5rm6DPmPT
c2GLFpoNiLxY8R9p81z9jRLXcUXbRb/RNcsQUmXSklALq4szWacOqqF9L11nk56uTAHgMfeI+5CH
DFsCwYf4obwpcB/r4A+KZgFYgRoLKFT+zvG2x+rTJFh1HiZkeJdoJvhy0RES09CSrrAw4GDJmXi3
g/Ylqp+BavrAFZdOTwZgVuNHKHOXeGbiWWxF3tSza/KuXSHlJrUdUnSgJE19FIwHeIZKpGyC2FIG
3XMv6KlQDca1kmf3Zz7E7aqs6geaH1bZxXdEbs17C+7tHb6uIG+6UA0kNW2R9U1Daeq0fHDBLpZc
eSYOavU+TAHDbtVW+qtd3jxaMVz2yvU3QrpPVrGmkXWCGRPOXyudJP2UFISctCxvt4Ek7uQK8BMQ
cJbOQmEq4PJhx6Uc4IRrdiEw4Mw91b9U4pL/1isxMkA9viXosxBUWGpethglnPnfBNTv0qIy0L8Q
SJdQvGI2HgqpnYZqBnzE3kqbQMinj6NF6eodgBB69WK+yJ9lsmtsyxwQernUmXIaZM5OYkoRFReY
zfS6qyc6k7PaT+EW68/cvKj3t96Pz8KvtCE5JzjlNnOtwCZxofBC/0OvgbAvMR2S7/kAETRFRpU7
9I9LVsQFQGYEa16GIJW5vcxBD272Gxr6YRlsW338u80V/BQotmggZUvMBU34FwifEEn9iQvZQ9s+
fFKpbgWH0n71b7HgF+zO4AECgRzF7QVCpz7UPPss0LoaSqhirfMRIiUZPO+T4ofifiVO8ndhbcsq
+1kcQjtzQfovMaIvvybTQJ9YPkLbuS+rcWFkIOa1xzCq8Sx+SKiUf/1jjoVhxPPT4zsrRl8dWy5U
xyWFIqrtAgeaxBW8fHZuWXxbyKzmPUk+6tEZeMsjcY+vkDvhJTiqQf44ZuuLrGAQyxh90RpaiaSi
yGWWqDgksPim5AsZicx+ojC8ByY+lThRNeB0ohFpGj+GWj+yi5UbCwDwvOBB5O3VSOVX4PDoiV5n
v+xPnvzg5YoX/t5vUqll7DK4f6f1g7Lh7vELbyr0qm4sZGo5QYbe48QrrH6BDSWNUJ30Ov7fyvtc
dMCKePvv2K8l74O3M4klJVDeaSGRnqwAn+bOZQjdBVSW8HViOdedZVeX06lde6sTZwGCt0a3Si+c
/+Lo4XxUs+by192JXd8Trt6x50YF89MM5ziuGjsidc4T8f/d0O7JU2kg+ey05kAuc1X/uME/Up8d
sZLki/Zkyu9qHg89iu3YJelnUgDiYIwe5E6gS9XDuQ1t/2WOn3YeQHCEbYxWhR4qAhz/RB6oDQ5k
YEi89ebfPUVfORQYesMeleUM15jJObjs3Df4TU4vHb+6bertTcwvgwgu2gGFO0i3aXDqd8hqCyWO
nDWcFeJA2yGn/gHdRSj791yz3Z2tEsv/g+QFrQ5wJ2r2OSkQrtkH6E6NdGe/7aStSy7N80VBQUxY
AS8zbZSq3/T/VHcrOQDO2GVNPbOTnebzduyY8LvrgM+v0UbNMO6YzEanKDcHv3v0utvaW88+B5jr
yy73uFethJe3WZ0WaJFQtzH1/5GShe+SgoNIsgdqf7acopxkwQNZEiGKh+R33tfq2fEcHZu5HV8Y
w0+z93CIcSJYzDOtSjfslVY1ijwOxnlp/KLWJppLYnXwNG0nrg33LzvJI7KHfqtrn3BkPBNoqZ7D
hZQd+pRunIWcZFXFx686YQkcwaXEWQaKpSVnjzs94a7O/Tir7+A71u/+LZqADP74ClrfiZlyiIOs
pcOdZlA2wtswmhgTtDcsEegyomm9f/v2py9GTc1pOc0Kq/0kPSyatJ5t+2zeJBMga4rNj7WXYeAS
rrmLIsE1CaoDCHcr3ZYzGFbhf6KRbUHTPA6GojLxEssqssxU9LoVZA/sPVsqvZQ1Xmxlx3UsH1Do
3mNgA37noM8oZLZ6hrsC7SALtD1Et59AGoIL5kfj+c1Eb9ngLrRidClPQt6FIL7d2Z/1QdZQGKgz
m5XXWTtSFT1o5bmiUvH+NJq67WBGezYB6vgmEHGkvcs1hbIAEk/noSvmn6C56LGHXDaZf0nWSr6Y
00ytgYX8tT4kS9VntxsMZ/Vxso3sMwd3oDKhxJExWQCc6fbYiPPxqt64MPOvQYrBQvHJc6/mFB1H
Tt6+duFQLebnpAnPEI8pRiaLbRLNAWTssmaqCBA4bEEHwkbZQL90+swBs5oAb5utIJQjSO9g22Nc
cJZzSkeiEJBaFbbYdqzU72g2+PUBuD7mDdXvKIjzrarRmDWf7S/dC7DUynrYMJtxuUkzXBHxRlCw
D4C8wVh4knuBPYFkkJ6+LEeOMLnyysjeJx2QWdSVxzJBYzrol2Xs4Cy7P2DV0FZ5jF5kAN/DHcRz
sl646Q+nCT/+ranR4NLjp0YTsz2uZj/iw6T+TZV+EuuyYhgqxtQy49RmpUzgnFy1caesWH0xoA8M
7cD6beCqEQ8aIKzPb/mN4qjPORiuu0k3C0h94C3DjeDdoz1+7qhGMyZpkLtTHeUe9KDw6nUvpwC2
CghXH9zebkR8HuNzkpZWFP1Xbv/lWEdGRFbjr7/RiztXhVREg87o/6tSILHmXoHJejqVkKexYi64
hIGTKO0R8WywedchcAF4fieFMLxQoO4KkuoX9A6qaXhbvJg4J3/jv/ko8c0XN7HkZmSX1UM9LPTY
EXpOIx+fAVCuC5H5qmCospzhcC2j27iWf7AbexNDWs/sz/+1ppPHseJyO+bm9awVBz4xVmB5OLCl
uCuyb7a4hRNlL7Gy0QL/9XreMzsdUcJ8TTd+e2LcV6g3qqmCKWDWxPsVDtoIx9nMBtjzAGRC1DHy
xZqX9/39F10A2qL3jp7YUe0xMLpQTivx86itxoZhbWD6A52VhxTq2WzagsOvGC/3w+kmZredXHoH
iBcW/gdu7bWwugNqzvCy6ro5eWbJkL5uJ9N5H+PX0XGCtgb/fhnIk8UuR68n3sRt1LqaJT2E0o0C
3Cst2JXy+wd8wxp3suyLkgXLMncqvwLv3wY1NcLvSDhxY1Os/un/GA6BSEWNV2ExqJy1xAC7JZha
lMvWUJ+/MbS1YFMYrJKX+2SkwFRUuJV5yH0L5QZYzFzzoNfyr10DO9uKTUAOFJgfnhXofYr66i88
u8wo/yGqii/UZ6+q+imAcW7uNSm4ddAm8tzvdnFRQeMnT8O9+DGrMGvyx+pz40rrKiTU33qvupXZ
c468rADrid6oeGkEbEtVPqN+UJS76fN1LMuWxBXkxLmjqDy9sOwTz4ktuwOdByvlVV6HQbeTXxxK
N94pXI/D8ypn9GRZLdK1fh0dkrOkgfPhrOvCRCKkfmjkHdsGNTc9Ax5BmdHyupDDKceHeiNZggSO
cFp18ELOAzjAdH3u1AM3JkiLCNce7LxEbnE4mq0940yyyrX1+/5E+jhThtNOQ/j3G4Kf3QD0fL42
i7JOcSDSjprAr1l2eEkmCebftLPNMjOCMHpfTmZVtZsF32UoYxcB+Ya4Hv2PVVeHFG6jcLiKsj4E
Y2nJ0+rdpeBJq2fNPE/YtSWv8zd2cpTEypko+dy72Zj3DbR/b/1Z+UIwYe1zPLZ3LW50xgSxGm35
8Hdu4QS5voenLPH4dKhl9ioCaOOsVYtzAl6VdAnItoaOcuTOfHSiZPbUu20EOLVWHVd9LES4Jl7b
fJsQWDeKM+UjZUa3H31WshBCdJQFZSVrIWwP/AaxKbzkD3nAKcJvcVY+RQcD5nLT7j/nBtWPyDxP
a8+2Qe1QyQuVvBZiuIyJdCc8eu5YpUwi8WpsEy2f//CmtAPsZjGP9nVQUa0JeZfpuMmVrktUaRUa
jLkg/C3/o0OwW1TqEQQNJAp8jCfFfN5zy7siZH60BTR5NewNeAZ8lDTc/Y5kfJyBgSn9o03gkmZV
EFRSwDdE3bekBYrcOR6GQQBZybey6gSw7YkzcHzcE9r0rT6zgSOxA12ymOYLE+hfSoBCQwU0AxwH
8EcT7cfyaZQbR5S7RiyMA/0xO/Aic26OCCgomMa5n+7U3CBrSlUZ8R1z20BNtXE7NwWlgv/842Yo
6LqkBN/4ViHAjVBBWLj37naz6mIFeL8K9kbS4QP6AmFxvTKo8P1i7eUPvC8VIFzKVUISdMOloxMe
i2wx/aQbszbk9JdN18V4tFNGTwbL95uQgF3kzbZI/6tLWHXXm8LoMIUQIMZtCkROhWKNmmV4ueLA
6i/G47uEQEdkjB/e6HOq0U2awrvqPhqRMY3OZuY8B4Mcpvw5a8ZdOoNPR+79FFsbs2rIf6z4at1p
jRIsjnh4Ub/ZW9pyFcHfC44MdCuX/UD8+v7YDjRDKIk2MJyMWjpeHItzITSXrq8aRqiolCMmbAFO
DeQYInfAIBcdhh+j0ZFdG0a1jDeYiM5LtJ/PH/TGfBNTCWp48b66gpDQjBiXx0PfLqcAyrDG0nWg
vrdIFXFCyUxvoPefce4yDhU4wAP6YQwIPG9WPMv9ok8pUcyYRL5c4gO9Pc3Im3K2kr5nUkQNoJCp
/S2UIuiLrnYiURkKiEL9wvJK7nvfRIp6m4cKTu3NNyBb4YFB9Vng0c0WTE0snEbfAsKycYlYfLKN
YgICc0vZtblWxmPHiui2tbqzeUGF74KljKLVHxB4FCVmdQJsw9eQBJXckzwdWeNebVOLuuS+Brgt
SwuewfSxaYCAo3H1ThXnwBVVVKtLgOgMbTNH6I2HFufmDxx41mE0PnJH037oYdBDIt2HCQkYoGt4
itIh9luaQTAJUTao7yO3xYpMS/KbzrzbG72VFiyOJe3yfzKITa9vIA4c/7tyy96DDUMcvVrJf0T7
XdcS+mKMTzY2LaRAG7LUs8um3phq6IqdJKh5J6B5KpgVbYtG7WpKik3M9omTBXzuCZ9PWBnLL2Ng
p2X2n3NBEw28xKabKAE9s42wypBTwzSijH8zd+01QOXr+l0jDAAcFtQb/KUXa1JU54yTx10fNGDB
+6hz9fSbOZ3uVePjm2dJ5MVOYLA7kJYVqqkB2WlaNkN7DGsNCuWc76e1i43cRA1xVrJt+5NXN7C/
DetxZztAI4BCehKZAWjNMJR8Y43UGGgx8UI2h53o9B4oyWN0GGCQ62Wf+rsMT4ia/bFFJRYEmzmT
8t6A5ikUjN+61dcHnKnuuiwf0nKPvYgrZfxMNFhatjRSpdprTYs9SH8MUltmnUAhKdKLKxNkHSK2
tGpTxLz8jOVUktcC2IaAyprhtlFRrhGRssVFdjBHPP6jxObJMcBCJ8Ir8aL6pX6Ilawez2N60r5k
QUVkXi0m0VbjTBFjwlqHWVxukTi6xVjTMqivLp3XNbGiwwg0CSLxpNL/9aGvxOLetpOEDPIRRg5d
ljneT+FSxKbUF0g1BQcp4icTbST2UkL+GpOo4E2bBMm32Pbn8q8RsGApZEGDA3a5XHbAYRtXEc+V
YKrfL5pDapuaLk52+fA0o7PqNmD64GnMI0QeMRg+8fTa60OaQ292abdvKJBDHXbQf862Mu40bxwq
WTDLVxqKqhOuwMJv7YTimuz7cSsqXcwUbujtsypXbQfQ5V9tG5GTzbngHDcjppowMgbIa13M4f0c
HBqm9Qd9ObT48OJAc6T+N7K0iWkP732FSyS7HTVmQsVG9f3T0O+9Djs/UMvKD8RqeHsrtvGFsEao
BmCXnFNrU5bCl9+7aaUeMlaX287WLjhQ6jt3FkgUMn0s9gzEd4D5xinWs93YExcxfmFJN7268wRW
SOVGuyqHeKkjE6UcUY+tideEBW6foM6mOcpOrZDkcPlwj/EqaH+jSKzRXAjcpy5Gft9goWCtHOsW
YMxUt5eo8bFX7/mtUeN6JmrAQp6dU0JVWQwKJfEcJR+BZ2/3BfcFkmmPahgd/YwmugPfe+G+yLnv
XDjkMiuDzBs84iQiX9ChHd5tydSzOalBmqScesX7adrj7ESPACFn/FBiYlepwKV1PMP7+qthyJI8
JZVSUg8W+7jAU0xpWsTGST81NvDyGjLo2YFZgySg/+jmGB9fbxrZsjeWJmWjJ11YVaLjBMLNSdij
RcP+ab865r7ylbVwIeJ3iVsdy513elUFmkr1tUOQFODx0e4/3Ety5k+5IsZlKqFPPCri5Kt/5J/x
VtVw7YtAtrFI+JZXTi43MeiK8GcRsKlUPfJ1mpEK5iYL8950Q0PsCb4vbWUBgsp+m1VKPNjbg83y
/GoyZx57qd6xl6/vAb5HC3ssI5WT98QvDqQb/+PjZLLFGIj+r2TfnTxwJa3KFe4BdEY5u7MOXnhl
K+A93knx7BXPcowHCVeqEHK159URbm08l/3pedPTqxthA2awN0jyTimt1OBLhgB/zNlDeXzxbqxV
ILyl4RebrbUOGoIYFi21njm3qmTYhovVy34J5LMekYE4llTHMa1L7G1jOGGjs/0YVyuj8ms4mFk9
oNxCz5Q6ktMMnwQcjKCcFVYRYo6Mj95hxK98//XJlHzZy82UjT5TTmH1K2aWYJdVWwjjdl25NOXY
YfjK6+P+nd/LmhdffKirEmaosm3h+WlZ5g1dQOljYbmaXWp/XbvrY6UAg2IM5Ku6GdSVejfb0EYk
ZSS2tq++PsM/wiCb9pC1mKiUV0BmaywDkn8+is9yQylQRA0tJjJAmjjSR/GLrjSJlzy0dU1r3L0a
GABnuOsp1EU6x4GrvAa7Hx7BMBISqDZ1R0dXLMHYTJwaeWz4Gzn2DUaIs6LoCqZadsOARZghxAas
TNirQyqsFh1rYZ5kWeI6giHIODPwqgTX/4XkyFIGGeTCoT7gFQhLzNGsqkMWBwL9STfw5AZH+mXR
oHskICuHrgQ05Z+Kp69LvC4jWfake3P3enIGzXMdM+iwLwggDaRyVlC+ODeXT9awFpJkki1UWpam
KAjlztzpMZfStbgZgKYOYyeWwjkGEu87KlqdY5vQtt/0LpsI9s39Z1ZpzdG4rox1+dc3+fVQAhqi
r+T4C3WHuPgxrPPHWvo4jtSzHi+XuqeotbKaXVa/LuL6mn9T/qLX9mveRkxbD2jvVzjVNFAAj9Ga
v5WMYditDakpKGGDBW2SL5grqJuYLxkU2DHYr/ka0ka42uJas564Spfpftjl5Z2a6XpfIcnu3K7E
i9/r1/ly4VS3bkkF6oHuF6YtuThTZ8pk4qSln5PgPrUYSTX+qRZJUAg1z0KLCbETVQATx/DToShF
n9M0BjzQp6W+av0sXIGIxPooSAELfkD5X8ig/sU4FBboBaJ9loA4sdaPEr3cDzugSd7fiDzLMgyW
f5wfGdTM1BXO+KJVspiRgHNU/RU1ef3N3tAq0EDe1op1hF4FBShmYWeHOQa0p5HYMXkpXR+USen5
++GvrvK9PV8ZoEccgQHyu1k0pUXJVedYUlI2CkV1011xA0UEfXaBHM0NaU0Vi5ddbrZ3e+ivb45o
oMgZx418XO8sr/cj50oWVKR2wfdiAuxA63AVa25jCDwStnHOQuCMzbnV2EZI6sZkgZwyRqcdZ5R6
/zYln8L63KAc1ny6LToru3QXDU3WbrYTIfMSj0E8UCH+Me715ObQr2CggRMLAWREgVvx8PUATRIg
t7WI+DUpbDgr2XlgGLHE6HImRPU22FeKGTHDCkiAzIky3nmSZMCng8VVwtz91gwy0mUqlYOU6jho
GuSpGgEjg68OWqnOG+UwAC9fdesJCyZizjY5rboYngHilHjwj9QwsIdoYhFPD4smjIUmss/rONAR
lKUSLSIBCByp+ZP1akHiO5JgxkM3SoT83YgOo3FiA4upYKzON09J8QdgjVPPgT6ynh3wWgKZK0tg
vxGs9kzFF7wiBfkFj/Qx0N97hytQ7e1yVPbs4mXS6M13cYCHDsEiNJU32iWcWorHmKI9kh0scvs6
2k3Q8iH2WEzDPQtJ2zWNFu2FlEGT+IoXq5Hixi3ATVE+YPpYQLYbbWHrCkke3OliOxlJGsuZVKoK
9Y5FBwkO3D7qsn3Q9Ubx1k+W4q+q4Ug0Eepo2X+m76KQRcIv48qDpx205mrBi6Nhcg+U8x8n44r0
OGdmmNPuzh9R0yPVQnZeX6GJB6AEhM7LDvlDq6Mtlp4/ATqO+y6LnZGlwZaiu1WU4BaI3J5yIZdK
+wXtICIIv+yuF7kACd+8yjQJ3JVs2gDqv7tImjSYEYMElqm7lY/c8yIdQyDYjaDRQB5wHQBZ4L9j
diV9jxVMqRgdXR4ZaxxwFEmzF+Ax2F2l/L59QCHZgla6/tEkdIX0FcH+gmN9WTEsybvGNCVF/zT0
9dPHGVUvYD0XwaB83qYIdx+1n51GKaIqe8VqldWWdpMZDRCGt5CgwzdVe9jQZITCx0Y5FbG2+u2M
vSsiYAs2M8N0u5X9UTtKV4J5B1Kze4mDOVfe+ov2zlGbrOd98z0QZuNkW+573AH7tjx7N2mF9i4H
toZKuEpA/pBxaZc8d3vhYUot+lhsh0JdPcCq8Tf5DtnmrdvyHuY9yQirFUBDOjoC1TsJZjs2oUph
RxhtVtqR5XuIAoTnYyXNtyEKOZiXAG1x6aRq2xP4vzjvd6pjxPP62xSr2f80cLcM+xpTlY/cY0xA
EZTjXO30C4CA4X0s31fKfeS0eCRgi2Q8ByvHTyIi6pchT0e0nwQCMp+C/ckCBrdl4LiDhO8tjx7+
hY5wXyYk+anVeyocz8Ei0kM1g+QphlExUbr0qP1DJ5IXGQZExk6tx/yq4mJGQVmZgIOV4hAlGGzF
+VAbBca8QZV41f3/Zp/Vyhh2ydAlSOON/0+MsxRs8VFP0bukZpllvEKogneCwdR96wjX77qlYMCM
iFk+0dX3GBFLSiZccB7kAdzdabjy7xEvEqPWO5+QShAioolJhZ/RyCTKeh+zi8NEtN0tA0DsQgKP
LoD20VJpVsZJSYx8tlhz7RMjs0Fp+QFdYYP0GqmfX1uAoGNmN1zdWvsMc0OlSaDdCebQ7+ROdqF9
BQuz+Bhn9ryE01i0jvVq3L6V/+LoerM8nnkbw6nBckJwinDqDpX4BcQWTYhEozP//ycuhS9MyHDg
Lo+MIQgp5x9jCw8TYxtnmmEMec3teczLL67pVxRHamsR4cOXoHylXLsYtwVwJC2HizgF7dYETUR7
8QOI2FcsUG16V3fO1nRLPN6YOyOm600OAtXhemzfEthBYnAJt3xpDyXwrpO5SPRlFoznUeA+piye
0uA4dtFfvIiI6cQ+wp81y9/HY0zvsOjcgHTmPy3RNP7/zTVClNbw4Okr3XR2fVqsOmu4J7dD7+il
yY4x7g4UwdMFYJO+JDPXIq3cEddoeZQdhIS27pLCruix49c8wJoeAd6BlRRdmLQNgskxp/7VAWmy
bjWfFtUeZCOL9YCWJN1W5YRQaccrXbUzW/bsxK9NmCNqPhYxgxAC3qXzTystxqTrt11aeqHffMGy
XyIXQvVo/9LJVELr6b0lq14Twhz2x64TN0TVwx/5O7v/nENEcpedHwVtIqRurl6kyjqMumFplNnU
UtuufEJBdWWjwioCYYsDmXzbhPV2fMH58kWTKkPLXgHETrt9wBmBOp+DMIT8Er5kZjFZ4vR7lJIE
uKHUP4c7Yu/TkDO0orHoHCcSFAp2aAWC0uIQatjV2y5tB9SmU3QooNTuEwR2eA5AvNKFvIvUbVGY
EMu9hKIWvKXpSLeKi/hoe4E8TG2jQW2WzvQHLlkaIKj/Ki3LXZ89ujgZWOAQKdsEto7K4fq57e36
d6GZfN3nBFbye0MKWVYdvyHN/VfvSHb0+fI1G221mDwGMEO/Z10D9t4uiEES7DYSxokuWgjzRz2e
dhDXX7BZhm5aKGiSGDKFSVs1n0SXlHhBbg/6q1tAc25Qy4ybjsFVVnDD3T3J2SlJnfF+balC+bMc
T8WOl1puuClcCwWLKwM3auT5cixN75Wu/NBXi1JdqSq7P0dO1ni6P7/BIKNAk9Biojd3iPVAUb29
tpAHWG80U7+J8eI+7J3idBXym3fA9imFs4nFIhGljRkEUZXSwlaOCfDjkRQ1lRli3NFpsLVlIoDP
s5M/EYD4R6GFxY+OnModjXzEWPWL6LIXCaQB397qE0pZGb7WIVSjjQOdcFRtlm//PHSD8IKn1i9f
OScIkticoEPj4V+foQB1SvLnLTb5i8Di9eVqNWF5TzLdjpPxctrtu7aMXdd3K20mnGDR8mn7X6Xw
pEnd0jwKMt7ikFKCItKO7TA4TCSfayhlHeYVs5VUAgg90U6fjRSgUZohEt39fuBWAV8aqFpr3BCY
JloBbSg986s7KEqdpRC9h1QvlOA2Hgs9LFbi4vsct9o1TneiUTuT/E5VTS2wwYfkJWxVC4p69k6M
Up0GYdEHh4VZ9EtNvdd4X3x7/vxUZgDtLWtMnSS0Lw5J1ujRmEgXsUhswTU0MHtE6bnhkHeO8az/
sAEal47VUUEMCIUwB6RTZQ0UQ6CztQOHx8PSipGrxJzYp4k7mLbfhjJYp6Eu4HAEmbJPEcDwqyvs
8Mby4KTevtaftVN/F1TfQq24Yn8wEOoxyilvTPNAOWUa2FbH3TqH6a//wxOu1gOU71SO6XZseHIW
WWmIJiKEk0OXPGVR8GYeov3GLJoAGYchGhgae74YsY1UOT9ZWBQXWbXgi6Yizj07W9DYsyjdN9GG
hQasaKXgEHgby6CP4ciJe80NASxC9EQkQ0U7ijdX3kF7shbB+vHXRCjuJOnkVkEjDikr6NvvStSG
VmerEVUNYUKqQyZqwddXxNOyWhBsPSqrN+aGEnwfZOTys8MzrGEyNdyj5qkCnQU47TNJ7mOq+Vd2
6SPmI57bpRjNJEYcdkATjQxwrSPryONwwGI87vlcI0hkVOT6OJaMqW97lZZ+nn0SgSkfMnDKsu8M
lG4NLJPQwdK1qumzmZ2FtoG7OmSIJ40geJ66ZZEHDvN7snpy3InSTe7frsjvGsF+orFvus8VZ+uz
RtOoB8YZw9IPpqTyZ3PewVgxzLXUOELS98OdQJMm20j246+etxdzaLFplrxb7S+8Aa9CP+npBORl
rgP2eZCD+BJlNwZP4x0ZWLWt5KBmlIEcg+3jh8eLLz3rns23Ieun42SKg2EQr1T5txXZ3txDSJ7f
q/WgkrCoBr9BL74YuBE3PI8wOhgRBJ3jw6laM5PNmdgU20nOAoeESJXesBrYUOVpdTay4aFV1gyI
4Re93O0GX5WQAipNDpPfls1kOQDjpl6VCjQZObZ8+k6Q580rWBc+QATlKNub0WsIrMCkKKbk2BB4
hTi5Y0J/MEwBUTnllZ6NkFiKcn6HRp6qNj+0l1Z4sWBkVUyCiROqD6uO1wgGl+meRZMsBVn0je9X
+xf3z8x41cklLjLR3tRC8wIumRNQRQLPZa86nvqUOEnCqAaDRergxjd2rhVWPSeHNxSrQO47eKz/
tCU7xLNQoMcSuO0PjIr7s0bkA4I8f2s2RSJoH+ddQphIPc2krMK6ooOpcAsF4/Lyd/3KIOSPiCJG
5bUudBS5Ksp9TtG12+QePD98kPkx7YbbpLo6eeqsSIfHGSXF8Tg2IkQPwwdTWvW84sjuoGdw9N9t
ArR6JbSoLjSHYVV5hBW1lMPk4ZUwuRZmtSqMXhVlITSv97YtuAYJupySjK6PsN73MuQ5l+GKt5B2
5d4C3/xUy5eICiYbRU0AxrbEQMoyX3rJKO0uCwY0dUTrJg4vca22zBIudez1CB2kpEEms9iduCx4
MBbdCsQHQ34EsToC7FoyeoaZNdpuremEEYswd5jC/UKz1ce31woLLgQNjpokWH9Q+hu8RuZlRuJS
mAmXGuciwiSk+bjMs3pK9NH5qDehMjq9nNAHgKW13TvV25MuKda6GuMyPUfblN2O3wYce8OelKKg
it5GQVIZbV8Z+BipVo7H1xkaOkp9F83Ya38VWe5FaOZli68FewE46qjSKLZczOpN0IWzKMfsJYX1
/vdcXVWPkEdzLuanKs7v5DDMV1BeQRFvsn2OMhyD/4Tteq7ESCrEg0462K9dW1VemeQCkmiUgvyM
296xce/Sw8x6bAZvQR3GvKFjGw92giNFdERWf0P1nmXapth+QmGCpF+KdDgc68pCcGwXduiYZAg2
r/Ak3xZGm7n9OeI6lX7SwxAk6i9K7wcOg/P2EsVDXcN0Ri5cJxHd8sjiSsCSJHQrQTJnzhoijYVy
3RjefoMWPE/zGp3TWFXreIq2EGw5sR9XhV3m61qfLAbtu4PMzSdM1Jq8KNHkUYWHvEkIu/BaZo9m
eOi1VVq1SoGmahYGaFZTNWq1qQNP0nZNiuVe77D0Kdyorm79dzklhqxJ6kuP4whL2br3Lx7A6YkR
q9cG9ER8zet/clftgyt9kkkapL9gIZ+5Pat3B1tEkQcKws1aA6HJXAL3REyhdGXK1/PWRirUeOfz
t9LxzMrGL/dWniOpUTOUraw+97XSl6+ob2ILTFajG+zwSf4mktH91ONfMDlaBH8GgZAyyimnWLfo
wS89ul4eo1FkWST+2DKby31CSLrbO2nx+d+9hqwxfkyrcidJ8RuvH1GuCyYmHMBWuUo9uGNw5V3Q
Vtsb3TvlnfGZltlJirT//X7DocPP6dc+3m7vlpZPpid/0mAvTdZ6ZkMbvb/+fC2hdAsNscPdHcml
qFs6dh8Sc4Y/HfTuMcOav+560Nqa4cHNzwVZwvJufMz79D67p/4HaPTviHRKM81FPJhU8/EfYMG0
hdKHOBLwCG+TMOCfxnfIBZxtiGD+47p7zumJtopU1CEGFgsrbew7+11Ji/rv3vv4qObRW4HOnWMh
jK+9cHuneSNPZQxHt3rxTuU5F5sX+mvBY10mC1RHf3wwrNKz68POwvS+Lw7lBqT0n7We6JTMPa89
8jfTjjqwdUgfvWbuX/C/Zdi77SX4FJd3Fhr9INuRTiuBCrv257WVeHBCOYlq6ad2YUdruYKLbhf7
iaJonjU+6ahu/w6sUmgwf5uqvKQs+jrF/YsRCs0ACv12pNrSINU1thEDF1IuEE22Vb60+mIJe7Np
ZDTYf5PvRvTwZvbuNsNoe/PpV7patlzY2alBa2fAE1A9Ru0rizPtArDmkctJuJsbStxPjlr6nMzA
2c9Xql/W3IEiP623ai5i5oalOICjgzTN/5jiqzbKBTc9OdkZwTnCcQvr7qEEpp4GZU9ReH6JXZ7Z
3CaqnJGpN8FtlLxKBDWDh1/ZSD5R7v5X2GEVCF9+RMfpqDDS+RPesmxgcp3nreQ6I4ojL/bX64IZ
e79iGddOeSY7e5tiSQu3CqXV625jwUSWgjpqw4lvdsBu74VKFvqSekW03TM7XyXu3j46XT/XLs9T
QHRZJ9myc5I/G+xkeaguFVfKaIRblHw8gVYkBQrl1DEYWP3MSM3TnwCicJo9BUsI8QStKCBKAl4T
4FNbQek9BVP1y1ZI4QREV2Kj8/Abs7nR+csYOXCEGHHU67Wbx31FIy34D9q3yQG6HxN3VklwnQPT
DomOIEXctjgQVlkvCOlH1JGkhnom44w7WXRoMFb3jDV2U2mIgKeIYH6fkcZ/6hqrAIItPDGlYrzP
BBSZFPjnwil7XCE8U+l9PEX1jYNNnMeU83Ml6LqUG04qOQCzcT3Vxs5O/fxPSSXjhfkfJKZCA9B+
pq9b7baSZN1fUWqsRGLGblwdv1XqJOTDMB991iXwca2ePsr5BIRNi69wZh39YVP051BJjfdsZJtz
pzfITJXA64IbSyk+lE/r6g6TZmGsDbJ6SGLdg28FItGfwUjE5exTNSn8UhlPhC63R1r+R1cK2U2j
UWlKu7ftHvXa296LkGnJHrBicKQQcRRkIdTAxya8xvvx+FNylj+VPd7sRm+qVWmTHM7g1B22BkNP
C1GxwFId2bYylfmZN0evNdisht92nOsmIjO5bF530GuO1qN08k/hzNJkfaE0Zt+CVbjB0wDE6Nem
1lkcMUOdtIUYuTXHTASfHvAVVMcmWNK9/Ir/xy+tjCSVUJwUtkZj4DiNONIX3e82fESc+nPhg9t4
t5Al/jIHTDQ6QSwj23dnUE4Kh0DWxMzbKO7isthBwCDmOaDKEP70SoMWaX1s7vVVBgX4/VvruJKv
cV8OTBYqqRIxGECD4oWzOGYjUJI6O7A9WAWsgtNgG0pqtulnjC6sS4YE0NtJxBu4gD34J9UqOTjf
z6HKf6G8kFxTr4O1MZy7277EF838qJDMwY74UMrWYS2HJ0Tn4jhlEvw9Ms5oPJnkzkSU/acNx1Ls
CKwv8nc1bBdYk00zDQZC7/Rktwax/qfuezp8caQccTBSdRI+DjfZaMyGHfj7ERruqy+n84LPJ0AF
Mzl4B7Oim1S8VT8NBkJYUJNgBNEgU5wV1HdfNZUjAZkNHcPtjM+bE/nRDo8Ed2Dy7uIObOyT0Mks
57rXwJHyaoFpa58xMrot6K2vAxPqW9/jCg9pSlUKxl6RDL9JN37rkaiCim21xy6EnLsvX7SZOC0C
3IhNq0oKJ/PdrAYNu7JVEsxIXqXm/k6AQ6IsCW7Cf/Dm4GUmGbreDLZErDF+6k+3Gc67u3Oz1zv+
8vq9oOsuxAJNVx/qY7PKtdcmWpWtfskxDBYuLUDaHxEkZzogGIvUstBbmo+QoQ+/aPg2q1TXVvfG
TTSFXwwT8OQN4YI8vot12CkDi8x765GpKRpiO1OnIHsTUxlNo8OVaj421I85j8GnNetUr1vXDKux
9wxG7CVxWzm4gUkFqH3RWZg5njxhSZfgpddBTm2Bq4q3m/3/O2GIFY32KQZYtWY5e2zvS7ikBQH3
aQo7PxmsAsyC2ojGarPmA18X2oeKskAVWV77qrTh9yA5h9OzlREFFkVE/rr3T68ic3ki5CDVgglG
nZ9k+laoD7MjAWXD/v5Tj6NQ4e65UE2lbWvrp0gu/8yTZ6IwA1HtWlcszSUEkYkAfCDqoAyoeCJ0
ZzLu4vFe+D2AIGiTPgfBsAGKGJY5IYGliUS93x6vkngyI4VpDlngShzF7NKZG3LwgFYPKHKP8VlP
Vh/huAVwMpVj3STOktvqk3N5H2YsWgJUyc3f+s2sA/eWHxW1xnzgCQmlQEi0D1EAbDx7Sow89wGb
teXfboMwhsIbjHBTSs3v9B8mc+ud0jUPJqA3jJ7Iki0046Ec7RPplnfUV/x7xHgUtRdFgbgNTeL/
zBg+PGZvYBiNPSGtbkX+1uUJGeC9yal9EfxaIhFKOXz7zt5CbKppJ1/OiISJRs0+J0n5C1uIotDh
PTQdFIwVcZ3Mbq8zhoZ2zlgAHdKBtm6SG0F8T63UAatnteimhFlbgUbbRXnENCWZJ3ghMie3S6oZ
HYMPBcRc2f0JYdnxDuaJiP57OG6het8NRcFty2GLYzNNp6gDXIK322KjFuN3JwsEKRi8EaXiIEZ3
GpNTsSov2YdqWWl7stS7ITFimNKjrQdUTiHdM9OZY+jNLO33Mm0POTpQ2V2DJ8FevfKnSvF150nt
5G1CFEsscexU4Ufbm44oAHSprnLY2Isp1NXtI5LBWH26mslHkCsC/8wfShSVLFSggrPLCupXU/GM
3cngBBkJIhVatEXM7AM5lDEsVNEr9Lh406j2KORXpjsBRzcX/9YdJfW4q1F6pBr6Aj/MGS0kkgYt
nL1eUTwRvjFKEQxJQlDVjgW01KYArwvAgPZskpE26+uyaYSJIBJNzAqwwKUCwTcq2rjje8ZKgg/N
M09fhV/ZAdcqRufz4AiXcO/ppibfAIxqwRaZiM4xXmsVMJXJ2N27ZbbZy50JVM/rDZLcrLFb1+m3
VUNCuApPqXYwJQoxAKhlTHH3YSZ+8GXbeyVH27esQKpS7P/n/igcuzqshHniyEJMefExxJGEmESv
LWsDcNbNnYaf4PwF/sFhu+kPMLLxuANfi9neQXyjfsX4Vpxo2SbjQT4xbyaROeLTG7r07u7gzoI0
1qhaGxqQCW5/1ESEJksxGxc9LNNugyQG4elw1bjf6fhpezbH+GRuxOv7egYbTe4t7ANZvd51dd/U
wLeqBj/ond49EEgr/L/ENnNhYlOO77V1tr8MTeh/8+eVpp1hvtGFAP5EiAdvYj+45CQYEGgL5E7p
mELS/sMzghbvDjIDyXqulg84ATH7vzLQBiCVcO+TMXhlTrl+oRMUe6IlPFNJbvvjtStQX3/lD9Qr
uf+Zcdl3vlPBFnERtCsfP0xpvckW7hPuYFKutanwEIkUYQIu6laUe1b17QxlBNNDGRUG9ulpSsFA
50GqLnuxb5OuEJoA7969J4hBdVNR48chyE/1DCDSTRrHgnEQ8d+4rzqbkzVVB+RhfQ5dmkLxBqOI
iP/nOi+6kxlIMtZIBZnfpSNgVeGS+uFKcZL5L6xsLgjBIQKfOtLxRCpcWorN4BYA84aNryc2avtc
YQygWm+3XHLCFaEbEBurwvrw4kSNxVE4vlQb7Spwv9SDdaIGIHYRKlR4lIy/Xu9PsHbyhUU39243
Zp+ZOyhkjAs1la8QMn56DwYbSJf2vJ0lN5g3ZxAhgG5Pg1b2M0zzgyod3A/TkQH0CnSYCnSm178D
z+rZNmJN8hBnvNVPX3MfCMuAovn6Ijl5BN4h/YCPTloCmW1oStQ9UdEHCpmzjwDoHO4M8ZdOHMKB
fCUTLLTM/5w/lvhXS7ob09TLSZCFZPZxytAbMosxyDCY1wLjbOVqP9IkPPEYcEG0FVTCcqnIKjNb
wigdSsLG9CSfwFN/XiMZ2UehWH8nQZOesHKNJxc0AfXVnKoRk+d9IGuXbkT0HHfJEZl5wVt9ewga
TxFfg6Y9o1GE59tvG9eNbypeBat5jE/ALGRZIz7ghYAHSkDClao+LZQJ4vzoNz8285kZmwYuw3J1
F+FMLllQ5yt6Al8b487KdXKI/nvhkLPuF5vFKEfvDKWkokh/aVd0JSuLgwu8OW19ZwCUZaPFcUbJ
fqPtbM7e1QNnWQk0KcBDXe+Vpig+pcHjc0KnydjUZWMTcYJHfBUEQUbFugDUukD9bhcPAPfvK9uJ
MzSyO6VGQStXwfUn6unay/XAZyz8wi9ewMuD8uel3a/G/dKyKb8CzhFp5sSNMG2eXUYtTSjzV5ab
Wtb4I7B/Qb7bm1NmLROdX5KdON5HrkFJP8LnGU1hZuA00EyCCC/37D3N15PHqz06OKRHCEKslPX/
rX/iGJ5X1XknGOBv2RzhI1lZYO9mfcSnOggzMhccS0gFalq+F1HYtq1PrGruY0tC/9Mr6HDrhMkv
ioy3MyiA1MBA2ZovgcHo0y3dnD0WVFYUAlF8z3iNKQrcXmAn4BBZLo8LdQ4H8i9VfyoJsIh867c2
VtuqKxQe23pznHg6R2C4OSzCSDhIBac37MdGY04TIA+t3K1iAGyBKIsCqM4I6UaZnCaYcdAkmkCG
fxRgNATQvWXbYJJ26v88Zt/DtS35x8gMVbIOfhbHtZSW33ZyaIL7SbIPXWTC9XWsY1X9GdZXHxNs
ZaHHcgBPS7SQHl7nVvn6MXdGRHNPQflkxN1UDKIyceV01IlbIYgHHWyVGGlVJXagx3KSCYgIXg9H
Q0QpDBF56khzGmfl0sAHDGDpcKWQHgj/r5oxC9VdGQdkQnRuHxHwVLyvzfJLuosZ/cIo7jaCZlwm
O/JEKeXqB8Z0ESW9ddv1qxP48H72TSyT949DAVP3B7asfMKosB/guceky3sIGsoxamQa+ZAHNwLf
u0tVMRtCuG3ndNKNSTE7xTM7foHBXy0utXY8Jg/dVa1PsnIUrc2erYT1bgeWE490ylHClscgL5Yb
vE4Y85mipyxSh1KT4xgAGToF9urmGQwSlQ7vaJ1ONl5esPoia4gM5IWr3O3UBBoU1HBnJEOuxE4q
MLT3zCHkuDVQE6holhGilvFHxHYuvmFFixjyx4y0sY4FKg/O9Atku8cnyldE3ibmD1ua6z9wtxLy
cOcr4r6VSuSCTJh1vhCW0Z9I3M8vwwV2Zk7m7bZSCHI9Wtw3ijQZdFv2tQuSQIQFIJcGQSLfcyTs
DvqiceLIRFjCOXnrkxqhIUp8gkVZhfB5gW+GdYEI/+9hAh//9yuSRtEqRCfCF/91ewxQtWa9D7oB
kr4LGOevAlQpVHhYXQUnPEnlVYkTmvw+gt4iqwqTZl2XewvtNMJ0BQ7jZzmfBXWp6eyWdYKuC0vn
F8AZ08uZM8XM26N/SmHYuneS9vyfinhzPWk0Fv6xft1HCJOkAKBlmFYF/fnUrywVvuMnhnNafaEA
l64KiD5fQcKSXnObx5PY/hLpBtty/6FxJoJsTaZ6mdnAiWqP+Q2oBlAojwkhhBj0mdhwstbu2pwp
N8Qtp1JkocsLR4rEebSjqUe2qkcbzwe9CGgmCjN13miIfckNtUn1r3HTZ4qFDgK7qziuEmyP1+ZK
J6fqfJVfclKzbngBpJ3bDA1RXfytzxrGmbVOL5wn4I7RgHtdsI5MyKVOq3Ztd9zAQdR/fZe/KHiO
TLEMcyTDkQ+wMqk6P7Zqj3+0V9CwBCBIYee0fOBaQfQ1yRnPouM+OgoeWOsQvS3AX86RkEwcbOYp
8rtLuk14C/GaMRRAtygvBkU7UviXFt8h10wANNMirwku/NpwiyowJgA8E0WVUuSD9gwhOY7tMsIe
BfxDmaiZr8OQ5ygv4/llH8p4jZGTUNBqIlnTO33VQ0B8BF7Iemu3XdaewSaeOU6UktzwLD+Mzx/J
ULUOxw1adj8VC8+Lh7UHOVtilPhAajCPmGxhX4/QFNIMa6Qs7Gy1BZtkv23/67pDxop1KD67nv99
7Q4KOMivR2/EZMlzGe6siPv3FfwShPE04cUmbZhg8LyIE8fNd1AtOoo8hgZ/0NXze3o9HgU/OgeV
dY683uej3Bg1FymE6PXO+YkMjaaZvwURp5n4BSATk8M6I94kq2qyENNfwL5JM4SVDyzwu2pfRD/Z
1jn6jy/r3rc8Ep8IY5tQJwXlk4XVaU3inuL/hob6GWR+dAjNR590z5ZkjcYALEdsPEK/Fm83xAlV
j3tcz+UEysfnffSL2ipiseYDuYjusdJVy7kPZTUhrbikOany0ZSyiMNI+RMDcAGJlLZHWxJ3kyrb
afGYuLWdQtipLDnu5rh0vzUEch57CJHFWqMkVgnqc472w0W4MSKrxa+6ps6dqjiRFqFDZ4c44SQ0
kI+Jj4C5KH4xH8cgsmuUYuhVD+nH3vLaBa09u3GnJBZAHoqso5uwJzGry80WIIDmrJvtXT6YRKUS
U6lhF5GQiqXDaiNs+2NyV1v1lHpeAf1/169B7UHishtrOZrdoUMcFdN4ZJvdepTvA4O5/gQxXyYR
EqkxSIiTSM8D8vPhmPjWWThIPv0qaRPx3o2boks+WkxWwN4Ra5M3VuMk9MEGE+wV/NtrhPrUXEJn
yR0GLnUFBDkT+uwXD8RvWjYNFcn0X0Zhftkl4YPM9ZeojpFxR9hm97XpsmP4Gq2gPWoH93HwbWOQ
6jDUiKOrWGgqQ611ZBEM06+jUvK7uNfmcN9Oc1figlA1mB5q/70zL7+aibyHPtdB9A8I3yae9S5y
ad4KmElo+xkFMPRMYspaV2xbGJZWFhb4ir9bSa2dCrkUDQF0adFMvJtxDPLYK3dFGCGluuCwCLu2
Dr8znWb11c7yIUeN4ALT/gNpXBThITPkhMv0+qWs9g+F8pBqX2RjeDNoRJws0mToGqGdmZmKR+7b
eBHHYHTZzwug9gBhx2aZQHw/Y1FXaeHiVw5qNZ0KLPIettSoK4oMLGJThkaZYKSKyqxvzdXZdwZr
txucEcKpEmv1xiNCmksEMTgy7C9BylXleQsUtF4H9ZhcoyN0Ezp/mDhJ7axLXwFncsLzpeLq2gdZ
NIVeq71Rfz4JS5gbOt2d3EUHeky87eEkfIuSExjHUIqrPxKaGMFnKpE2eyyPc4XCzaNvCE86i/VO
EnvAz0b3CQF9YAyJFotbOZL/UAgb+t0y+qomsnG0W/t5DWYm/4gmn20OV2veBYpndy3fPILs8e6x
M6ODq6GKAH/QLslf2ByzAA3tOPxgWGqVe9ukkp9GMzrziO/hCa+SyE3O09KiDTtB4Q0iH+ULIlmh
KNIooQC5rOlmZG2WGvltxqo65t+EDwfEdKTNojE+XHLBuiFXtiTOiHKnxG4WHXfXvjt/Tb+jdCYY
C03DiWuzhWnj0viYQDQgfixLw/9wTaPZyOwQa/HObe7we5sh+ISbiBfBVustpSyYqwmZ7+QmRmse
5VjBucgyTZfPbXKFWMW9zz1FVzVuv4rfBVs/ZOvH95aKmbY2JiIh2UU0ypHOl2XTEzP1RR9duz4y
KlVsdFWU0OBDby107jLUFT1gWTTf4HzHNBVsprLgYFsdOxjI0iCgy99JLRf14lAF34ClvtL/OiFG
Z1jLDjpJnkkvWO9F6Kc4YfI7xVeVYz1EM9p9exZwIyG5VxmXQ53G/EW/B1pBSq7roJHHlWtrL+PV
xSz52SIVfBgDzkc7rFC/Nq2N8PJWIYKLAzNotXvw23r9bAZhlLUi0V4SAWJvEAT8ZtYtOwz+yCli
zJN4WriRGiClnmVyJbpU5EfyWYejjncUCrnwNpGkQWyObN6SJYVDwVmJZ7WSIAg2dZ+T6D4DbGNe
21t0foT5dbCYIRl1a7A31REIh1CIz0mT6+nt60BitkVIIgu82KJUWa8xPk2gX1EhWEW6MQLwxgfi
k22qf0zBZnI5IPy2e2ixWMK29AyOybCrFT31qXxFKiR7zkWI32WuHrmFkCc3H7InWcx5sQULEq9s
BQIEtzKBjJHU+JBh84J1fE+PdyEBQAESGmRnIKKIwGf5pHlYryPxemnkKhdV+yPmjnRcjn2+g36e
VKP8ON5esGRr4jmHFDP784Pn1z7xKQ99xFnRs3iWn8IboXw/Zuiwp5Ha2bIt2DsCPX5RCrRsguZx
arjhK4nJjnmijmdQYbkGFkvjfa0+Ew1rsU4dSfxgwKt0btK4BN+uCxpLvweuSLHlYg4A+9BbEQMl
I41F3oVMbqitWs6keDNAIA8tT8xcFXDbjhaF1k8d/EbSXwC/WOj+KiMSQUtUZvK9108Yk1NToFGq
nZRNPEOwiwV5DzRRk6KexbM3hRt9SHJWinBfJ0EOXDCCWU3SGukQTx3+ipW66O4TTnOY+rU+oVWp
dJNsj4z9QXQbix4/wGSrcp9YbRdUusM9p7YklRzS6y4J86lmSVcqyaXao2hm/TtJpWILLvY94AhA
+e+klQdAW5H+ozRp/3QXQAS35oJ2yq1Yn5g2eGuhXxZB9l7YW5PLkJi2P4o+X3vYzWeJJjXaRdeg
spSRowwlZywTm6NJIULceaQd/aePmIMtxWx2/2Y6AovmWPATj0FzKNQYtNF/i8Ro23NIYypBWbA/
Le8CVvc88SceCXQbrkzIeFtBYYb3nsKuhhDR3EjIfxC8W9Dz0Z1HYIOAariVYLeuy70jDjz0T55J
LJ4Lsx244Ujs8R9BCo/wgXwzcDfXIVwxFxazXUpnAsMFUWRttOHo0zASMR+ndJKDlJfpDxmKJFDa
8WLAH3OU6nlm/KSFG7pchFgXYdhSDj5dBrsfonvZOzwIY3PGI/YWPNDriQ9oAkJn89V5U/JzNxPF
b5hUuuWImCNQtHzkWNhQyboLBZo4v84Gm48wV6ri52MouIaUci054CXpGIO/ZdJ9z76EdPd1o2r2
Np0ZObWf7j28QylviNf4Bxt+jdlMieMxsu6U+248wjxuckwotHv42ufr1A/xwUN/x5MNfF1bBE2Q
NhcnGPyIR0YBwWA5r9QyUROvF/a9riEvx57Cq/9UX8xnxTfNxxHJMwUdHOInNd10FjttuJ9pMrWQ
hbTyOZjsl52VR3lHTW4rE7cffrgPORmKrbYlLdOHeSbcuPyy07tRqG6UCV8bpuq28Bf7g5KypEoj
uD7yKZzod+ghrwCIC2FN95VRrEkc0ErFXQZGgm7csTkI2F30zv9KXOaIzEdXjHqhbdYd4+E6F0ot
ypBxKkVo8iNpmV/e/jG29Ff4byXi2g+r962Gx6EaoHl1/sVbOKV+Rc4Bi3nW4oQ0R6lGFOiHYRH2
0/Xd4K6XuhWY+tq7JTSovHDcr5XNcB8uW74WLM8yLIcGcjSY0MpZR5X3MHD3hWZHf4SnxY/7VyPj
9Z/8sPZHwByFa9ZcedL8Nfn4A+ANhXFZsyc47odaNpFUBLGdaCeNLKDeh7wt8sfMkzPsgFfMoxBk
/TrqFbXHb4FYQarPLIrJfn/YpQae0XgJwXBfDk1qyIm2uhvZy/HCF9KfT16GfvFShWAb8MiGBAIm
JsicmkJenOh1UAhEFUcLrfHM5l4cWinAf3uaDBQqp5tJ7DaGuSVRt2fjTsPTELGdsKhE5ZVk3bSq
Uri89U2JmElA7akfN6URTshvT1D99vgwVV68/Sz4zScTlY91TWZ3271PFf//V5p1cXhVKWiUfGu8
DaQi0zHDnEejEpg4N09F2lma0Gm44VaMKdfLCpc3acpqj87SG/U2BI4bfpszhSLeNZVwpWi+3wBG
AFo5hrlv/CO8U8123Gva9kGpbi2S/Hx3IpESTDInQp1jatc7gcxIexWJQ9LV4gZt15iOJCyfhEfp
1FaOTLU2sUlTU11LQ0V5sXn/XmYkajPlTu+vr+NkTatyQL5GS6tfzhhlkhjq8PBEXf2VjQjei5j7
hQ90ef7H2OAt3+nLu5g3uEaEMEehYZstU3F9ebHnGS09OfxwB5ehySy+T4CKkQaYU0q1Q4nRjITA
vQ7QfqKK6nS5kruyTH7ZltaxdmMGJpBIl35GnfVBFR0qhrsX4ll1WVYAw0Z6Flp8a+Si2MhW5ziA
K2eWIWXm9A8gBeSgjYsdEVr6pAPK1caUFs3NdbC9tj2Wmc7g7PVn37jPCc/MCOqv5d5+xo16LQzJ
Ili8AwuuxLM5IbHQR8kv8YstiR1EtxL5Hm7zxSlcizf6TAoHyERo2lReeHkrBAOI44kHf5WDsppV
pVK7DDKXxeY1CxCdIJrpekenIn4HEEQzt1NDXVj+Kk2wkU3+vF/IKQ3uNDXVBbf1iC/8NeLxVCw8
09CpOvFimYXYfQcbbKsf9lOPNBa394DTfMZHUZcqGeqpsZboHsxEXCs/E8abYeukGhNcxc/BNk7h
YvzY6De9Oj+HxLwnOCZV1dudTKjG/XcUX0NrDxTV6so/diLkzDmTwlF3PDqswoOjcO8Kp00nxGcC
HUGjI+x0/mfcusi8OihStxmNCPTh35gawqoVh2/EGE7q7QqEZa5F7iikFPaatJ1kHDbOxjGfwxoZ
o40L6dz8QDSt8kO10x5V3pcNYMZ6gFJaqM3BYB2dXLdQmQgHeSE2ASwZKYxwtgSS764Ak9vwARXX
78hY4YMBo0hilU59DYlzl+CbxmbaiZ0wJWmRcE2UmJsRAwpALNIfEG1dSzjeRMXB48k7eyqYPGNj
qvYUMDiS6p0xVD1NDrteLsTmMQaYhFVrJ+zk7yihf6vx76Qy1vFc5CZBlwJJc+49ULWwOFCuJZvp
NTtBhVMyJ3BvbAO8tPB0XH+/9PtTSl23tEhF4oDbiniDLzy9K+PdxTVABJKreQKmIRiL/lkqGSqn
85bcgn9rt4m2m20VWh8uE9xuBnt1PKfbqjfjZ6OLBCz9DZmBJapTV2ZmJYOdHtTBY9ss3M+1rWah
tNf0da2pd9nIzD3gFjygQnlvaZzDXUZ7IBDrrRcRcarESXwHmcgWqOAjTDbizTZLAI0lknOiQlZf
lhp9CoKpAIFiFZetVv9qqduZZjrMtfFSW82XWAlF82JBZiAdRg6/nk0R8Xdt1THG+FY8ntIQlQIl
AeeZDPKrTq98HeeGfnhvPl0uEDlM2/VIUBwa8LXE2jZYImQcp0POcdhr77ajmIJ/bZ+ygFjTt6U5
iqyM5nOZ0I8CBPWzOBEIWOnidDSMeyYD1UMN2EpxvJoGL2CfpV4GtEmuc4j9e76zk3dzd7EriYCH
d1Gd6NdCLc5s7vEty3rnEA9w4yWtr05a/+WWjxlnKcj6n1e3j00es7hZ6VCxIDijRt/cdn54f1b4
Mb7yxdm4D8XT6mQ78Au+u3hkuNruOfHdOP+/gZw9jCf3f2CiBSVk35wSnPSJXtOk+LWWttzC5Wv4
9fejyo2KJWwchYTgNh2SVoD63bB9DVJ8XhYaGACCC6jp7WEWKjlhT66IeIeIcCU/41PEBwciK2Xz
QAOeYY/HLmTC5CLhRE9isk44dULNMbd+v0DlniySxo9Z2uf9MWr0zrHG+QS+DbU9AtDVA8SbSHd0
OkAErI2w3hcH2dgPEqHc9YnO+RiYVNQkN8FMFgNvPi1tSDj5aez6u8x4G/7mDgEH++gULo9GvRhs
G2dVJqGxkiyOjz3R3YyfONVZ2XbT8zk+MJW72r1bQ9+K9/Ao4b0KDkhJuoWh4c4qJmYveBAUFgto
yeiciAsO+Y38d0GhMcrK8dhEeS2AGsa5nvEleQu0Ruhj3Qsqn1+Ijtc5IyJuB25S7tE+pEiih4yu
RWZUYKJqJSVAaDLhBVpk2LTgjgkRfgfaZAUOcyyC0DTG/rux5ZYblCmDVBuuhFxnfafPSHDsjLiJ
r84Ac+iNwC2hHpOsdb+9I55iYHW+ZBEsTVGRXAtIei3xuCAslugIDNW1kWlZB0cM2Tb3QzMRn0ec
Z0VrGNc1EHZwduU3I7ErjqNaM6bKGZjb3UdtBlxgSpyJyC0YHiZIngM5T/zcFbbEzRWj8RHBtbG+
C+f3bhmCbRnBFiTaOaJOBGgloAoFZ11upkddvpQAIgaN7k1sgyuLVpvz4fFB2UkPwTPap64nQYz5
hv2rm5PbAWK6dXaQ9hMKyg3f8gl3rGT4un3beLDL9uV3irQgRYuZUEXT7bZwTYZBQsV8C/vz3wQC
GGqZQ+ePLTRkN89Ww9EF3f6w5t4mRqbwkuRZzs6cAMqQS34Jm5Om4dvBOVpUzh7MwC6l65xYSH/q
crszyQeYu+DO+8jQzkrqiCqGvkmEgz35Msk9c9Q+6n9Bqz6+V2KCZqiyxwkBI93u0QMFICpcqHJ8
mNiHG2VyV+U2A+w/0XnEwvNov4u/cPiuIAIq+QOt5g0D/w3vNV5yN1nPLt1FFb9YInESg2W36FrQ
lL8D+kjG4TZiw7+sj/0huT8zZ29SKYKhSGR3N9WzZyAx2FU1TfCm6GvYLtdaqMAngEK+LAXoNUOB
M3sMFXhG8S6KRn9yVBeR8/YOAw1mthm/2PCGPS9OZnMHjazsxFp3F64JtUG24ryBvt4rShnNpBQ7
03BRs28ockzuhSfKdxOuraqdhy5BME4uh0ZWmHKYtX9/Ao29vh5PjvlMeuHcSLVPqqo/4ymBSIZe
G9sn7TbB7xqkSEPtc+RyQC3Nz0WoElQ1nO9L+PLXDs/+RcgG9kexwC7SwekiRQihjMuXe3SIwRlH
Bh9nVKa7kza+9rN2vTXRGlZaX03DJkL//lzWTvIZak9YJg5DIcVAREO4ZeSXuNRKYkjSkge0A0iH
RdhyuK6BIDZ0Rk4msXJBDwD5+kg4/o8ehgA+n7OxZYgoU2rZH92JrgxDvO2EfNk6I/J7wMJHGwFd
YN+kxT0xEpKoObFl2pEKqvKPEROwOxqwxfZpLrSQ/Phlh36ysGT9yRn8p9CwhqAvAfN03/PDlJhc
tlK68omnz+qbv3d64F+8ivX2MlUvMJYiJVvEvKEtc0T/1A8+jeQdxY+wfeTChGBlHqyrOWxF3f0T
w8wOQdwlojAPUdWWQ4BcSS8q1Xk/U9DNPyK1yFtCmoIMJiuhrYmEPWYZuuxlVfR0DZ3aIpQP8LZC
NNabjsCh/wJhdLz+vDpAxyaqfREJ53q7zfz5t33YdBlNVb8c0Lkqn+cbtI8wX+ST2iDmv7boMz9+
n14JYQxPwzbcB2dRuZXiXCTa/QG8iOscqudFgyENnAnKKY+DrfyOawpnKfUOLWbgL1II/ccM8AB8
u5BXrsSUm/15G8S5uhOWhhRaODgXzf7DhnOEK314ksAKsooSkxwNBMAtI8Xjk1kTwZ6XDlkFtZmd
PK1Wx5ctPp4F3e2EybFvsIz2uYD9sWHTVWsv7fglBkHSKGq1YK6PQvnn5KL14R7br8PKrxTNMR+R
5lRMksj8R0/kki16oqeRhB25OiZoH06vHM+MuUIQuMsiF9sXKO66fYTUHqkBuwAx5p8VI8hN5mBF
u0V131YFECukMpSkR4KGpVrvPUxhBr9VpqoYFpFeanzYNqWjng+4B2BCbAykGplxxEs0zouzLV/3
td55JpEOyJsymimx3ihMC5SaBUOWOGC9cPmudGvlu6Oy8trXydWEKXrY94JwIzVG+3PMfAqV3tAD
yt0qmoRLPcdque4F8Vv2kPaTPBwhKgLOnxcy+O/hX2VV08j+crtcVuP/CepUJYL4/QHj2xIWxR7R
TfjQPfkrp03yllG3mB+BvCBidSu2z9BYd6wC3Ay7X3n15nMWLM5ItKVVudHmhW2u61tJGQbiU4GU
59CP0JKsiuDeO55N+Ii4WjDGILnVr+SYz1+gS53J3E8IOk0O7JsAFOICQ3a2XgLgB7/nVIiBRoug
iITUQ73GD+QwtYm3GafhZvTB7AI7ga1VrIbBQGMkH/BCi9XD9NV6LgUDeEX5M8eNv5J75xTl0UsY
UZp6nIEz7CJ5LWqtS6AK1Qb3nfxhSEL728GyWYRYghV7znvc0AbPEUXmxoOsySp2+6SMa4c4+9gG
4ZapqTW/BjSPUVoCIL1ohy5c4AcxItd/50io6sEDxmqKP597y3kLjbaxl3VmiUyZ/pMdvYeEigUL
HOllEKwXqdc30CeD8PudF0b5iko93XPoATLWgp6so1A2TqQCsKSX6kM1kfDiSpikUiKt/JrzsHvO
B2Z64jdI+IXXAn0iAOARe3j2iGVWRb1HT+hKjbI5QyKOWnk2Luv+T0GeX/NDpG+AFwCnxbqmcdKT
F67SmSR93XlQYduBbsZaGyE3zB4w9s98gmtr/dz8dJGgHtM9Ie3slJjhwpHtT3iE1tR2d82VYXeU
N2HsM1Hziw8VQZ268xT6nNZ4U6hRdKT++sJZd1it8N6AvvPvKm+W7VD/82Y99p/H9filQ4NsUutw
tDWVkv9+y4nRwmT9+jmOp0LKiL+rMSyz6t0UJ8WfkRI9kjS3kB6OmdkQMc9EPGkIsvi3alb4PDbU
5hojdTpaYOMm3pP3fruA8/haxxXK5s6XYSLDU7kOuwCxCXDqnljTHv0F43tnXvMMj4zCdTWVxEUw
cCWTwqwItGKX1JtDLY8mb75vKqY2S6mCuCKJ97tj4URFEdmkbfM6aN27eqD1QyR2DOhe66Ewm0Z9
iRsXWg+zSIxnZ4bxHdpUaA9TVBzf2INHUTFtq/gtAOaKOrkWg4g09Qb9ONj7gfP6YImPMzdrsldx
yQpHowV0CUrxh6cgs0KmAdf7xR09k/nu3EwCvFTVfk5C+T9IbmalM4918818PxHk1kQ3oBA3EI9X
SeiqI9gh+/nfuJ0q1IsLyJjROdZKPkb1TGVHUhz4zKcHp1KsFQcSB4W7hiG8BVBpVgZnBu46tgeQ
ZZnHmSk7OHjPAy7M4NyWWjYq8q2oykCtiqWMOoxKBJiLLAFYS1CZbjud+qWmmd69HdeKZuwJZRHE
oDFhtDQZYvWaCyV+F8XE7nwMJmL+RknuMUgitUMqDfDTd8Dl/fLs6TABdkI2haKZa6RC8NWYPANI
AQ0pvGLoxrd9iG9C1X0qTL/fGNZatDydAxM8gX+jvjy1IR8jLtZ4uS/NXFEed0Qvj8Ow8vX0FR6E
JYNuqrGMecbI7DfUb3aTjiBb7WG8GdU4Dy8Mm8ZqhbUlKJQDPd3GLq4gjlzJHKTDZjGI4UhjGxkd
gE/DY63Ba0HqUp/npO5mRm4niu171SH5koimvqjbIY4+ngd+IPEAGp/FP/diSzygHL4VfGpS0jcM
Ut+Te6JLdFYaR2Q47w09yJlutoy59nPkW2TBvR0sfJ1rKU+JD0pdrOpyqfgg3iGyf3C8ob8TTgBz
ISHYoV6vEHc6+8jqH6Q8VdpuPdwoG9WUdb/kKYuqPTylRGaD5xfj7mAvkmfxOdWQJ35uipdQtnXr
3OKmS9zp8nKzZ8R2ac9rL0B9gvfNeEIIJUwHZqQL+3R9I4UAivXRMKa8GgHKBiRqfLw1w7qqXj/Y
6XrVF5izQx1aHPa3O9nxWtLE/49BQluD54MuVSY99OhVPwyGxd2Lsx44uHypkXH6q3SFUbH1iQQg
XSE1J4Epn6t2urqh0M/b7nmwTpuSzOMcNRlHLu2H9wyvf8UOoUxwhCxD2+mABtkv3cflVhw/ATkD
zzT+nW1Nmq0BiyT26Ivuzn1xjTJToASDVfE3HRfMwfD0RG8k3v79Dt7uICgwvYRTh2YVqpNgOS/t
/OEIvwvWy3/FIVGikUjx0RQWseMsdK3ZSSGCiofwY45uLnR0TdV75+sg0wYGJP1RY5OtfIg+rXvs
V2AZbkaV9WZCdQlazWpknrQpF+1AcuaEb/cibW3AhQYQ+rStD5zCXVbpp2fjEqP3wM9ccwiJOGBZ
MFHh50WiMmZN7fWIQ7gRDZDzFRMBJNKYc+EM3SYKLplpZcX0DYDAAR8m4XgnKiZgeuq7ojqSKhf7
LxmPmhh9clAX3HbraNStbKt+yOaPGgTd11kGBjSQYYFOK+KJEP+cD4IqxYcbl0R82ucUobcNW5LX
idq7YL+XUZf1+FOYuSlsojAtqmKOrzCpeNZg/IWLw314fd1SsC44tEXKdPyQzWxPhYPlGJ6VNyok
ED4lfZLDLMouHT9tWoX9MouQpoa9QPHz69JhiI/DIA+pjytJBWUIgGfW+BoS9auaiZK5Nwd6DeY5
VHW1njvcjLjr1T9qySKgsNix/rmBGaJkAW5P3HPc1o+ueJRiIUPHMy0OHneTJSYN0ye4h+HZ/bFS
wt16wrkZViWuPrfAFY5l41gYRJ5gGLFuOl1mfGalpRjcpl/y7uZaF2NkXWEVvTZXFTwXcqZAXB5D
T2ZcX/Ln15k27TSDlcNJhDwylrue/x9c976X6zLDLvNoLOrLUbUSVoPzbVgtA8IQ24+hWuuqu1dt
8YF149E3hdZDrkiJZSHAqmkKMJZhMuG98ERFPnLaRIb8JbD39tZQ4Z24OnJc0FWib/se+1jKnhQe
w4L7N9mr/YFf/LTfnfAvK4n79iDlFRWw8s/0ZH82ywNkhxfwGpI+6pXM+sFzRBpwkr8L+jd5uqU2
aW3VAQ3aKifOzQxAaM8RSBdOyvluvlwrmYvSOuQnpbeYPJpg0vbDNTdYtkkMYQrQomBGbaja7762
D3knn2Se1Egb2AGlsLvth0LKmGYH68VwSkYlscwRVv7R/aNO6dbzCPynIT9m0Xfreko/p0/3U1Gd
Y1whtvAkGwYh6trfOuRYsdQ7aNCIvjN813IZb0JlAra1mHHougxLH+XbaLrvAcR5QtS/iwsYtbMF
cFIFuK0L2hr323Qync3nZuagPg2wz2Iyt/C71TDt8ukyGq/dhlogxHrYN+MkTJu7JX+891zvUmZT
RBMUtuIkL9F8uIsTFC9QLCIcPHP8nAld0WJXmynch29oAjsT45Gy2IKpfRh+cIqw1XTKpVyLXnEn
6unLPb0IdPNLp9VBdbdeBaBbP6WKLdFxQ59OOIAHYbu7iSgsM3cZEC6mpiJ62/LuoJ0ZeiANRqbH
dWhLGovbnKXQlzJK/eLFmFmHKYBFTqOmS1VrepO8zAgqLJAo1QBp6v+FC7/RjVnt/atFEFblOgHp
8Y15FexV1pUy+Xv8b2KdSVtn9nXA9UWUcXkjNiX/eod3jGvIMcaM35ZXA0/VnC/jM208HT8jtYis
nwO3PlDJPjx2gAoQm4JhPhXTQhKKmUH7iO8riwh8yMcL10dU03pI6eVEl7fF00di2jlKCIsFpB6J
YQCGbMnpnPs/hSxYWe0SIzk4DKHursGw9hR+PQQfU+jrO8AIrnDvFrPHLDFmZjaDm2ocfgCz+GL7
nRIKS4gESZN1BUCnRwHPyOFnAQBhFaBwHDno6sJ7oFHl1T00NkxN2KZU+y+EmKfKsICbD0a1hb1o
r1ND7BT90FkD9prm9Cotje+BJ4I1RLUJpPk/zhIyBpB/wZg99VHsX2C1x5kfsZdfKCpOVLTDkwIT
zszQX93HfgVEIVQGPTtRqHlnf+DUn+nZd41YETMFm9iwf6NaBj/sivHUDUNJUzAeZUgK0oprwpk+
RAv8parwFrUzSG+K2zd9iLq1TyTzpySPV1ze8YLHwrHrq4hMNXHDqFmb/6cmunIjpsn2ay2sUgIj
nBroinh/8hVw+4rBUPDmEdIG2CE40qX9awNtE1hSTR0qgPQMXTbGzMgR0XI8v+yCtERldWiuR7qc
dE65j2zfEFktIrUBl/GdG62049qciKrOXKjby1wFpZB0z2coQal/FLNGnnHIEfkwTO3CqQWNaDrm
fRLdksHk3oDwa/Y9cAIU4CXonPLCjlw7+35yDDBojX2HF4FvB8qwetP0fGJVEDhilF/QTKimlzom
cX2BcsNtpwzM/IeOLaLyp9PIPmDcZJg6p+CmuAm6uR2/w3VBOz/enYBWqZF/960Qbc3A3gnpQkQL
ioIEqbfDYvnYmXk7KihlD3kLfa6s6qRRaOwv28P5uXIh1a5Ej94xlaGf09aSWY/jLEXi3WbYnNK0
3pAEX9GSAWbglLhh2viJRRH8n6/zptY3nuhLjyaPJGKhU7f9/9O0PoPHeDmMWCo2K+CdUG/wfqox
xgFA/GdTXBvi8qOmVMdTkXZt1+GzYZepILBe50bHbRFt99csqglCnf1sR+iY1ohJMnPQK0Yb/wae
sqW05Gv+75/xCE03caGlNh3EFCzZ0cOzru+XpsTZlOLiKxvvl0MRdM1RJ+uuouF/qxvAl/VAaBC2
yQP70yqTqHq5sDXsSi7Y1vLM11zT/0t4Wr1giUZgETehrImg0tx+sEI3q945mwruFbpB+3ms/PtG
4MzPFmZh9BUft/R9O9rFK4kVT+4uFAMw+HCaOFH8MpmBaNMS37FgGr5unffHLhhhf8YNNte4lH89
hNUFmmYEn1ATifE4n/VE0DYthlreoS2WLhSlPKBChP6IZnxNqR3ctsZm0g1VjqdwNluGP//n+rux
GXVwGPnDG96vRvVn5NzCMyMa72quFxcrBSj5/AQAfOa22JU5f3Av9QfMqG9jkIJ+wSdYmoBirG+S
Gxo+Udl7+TmJ9WsQEk0rvSBwAiEShdHiKX7925bkMXyAN6LQZju+r9bSuaBWrKV4yylIfjYjcS1y
3f8BGTXB28GcB7sxkXP57/qe5KlT3OmhIqnvp3OSevPynJq2ddCQRhz2ik3yzI1rG/15RQgjHzXw
l7llLk0tj0HTBfdzWscIvw33rczEEQTSlnjEAlBZzPq9cZ3qxrtNPuMgrmbMjy5SFJGJ6Ac/NKgY
Adyrfz6iAz/Q49mBV6IP76Gw626/rC4pbx+BBFuwzCiWlUduICXj2rBwB171RMqeECeO8ojolPQM
AmqSsEzGWA24nzEFwk6G+yBaX50N2E2XvIlz3Qe2+4ZiqzITquJaF/t+PeQVcCSsMvKFm0SWJ/HG
3+gSf84jaRnZCvusQHZEtQKfv6YkzTcG/msud2CFQCtYXTeF+p+a+uznG2aOszY9l/v8PvXasn1h
q7WnT+N1+xO2ObJK7RVoxC6Ol2A4VxO0EgOGCuFnM1vLqI2LsJOIu1zrttCmvPZAhxFt3cCFDxtd
6J7Vj/rC/Sq4QjsTMFYweN0C1+nqcci6VBx2VWg19fNRaHzXCjEMgavZ6xfNNzcgYYR3axmU+2eW
/ncbMJ1bXdRTg6eOcZN7G3BH+bNKEotPN9az8pDPgK+45JmE7AEITSwfRXmL8JlOHn1QcfEXYMQi
TaraCq2BDLpTHVbkuwXrs3kDuImVKkfz5TWw6yAiIUFqIYxrsl6j8i6Yy4ltWx8vbJoz2pzBBIbk
3dvDfFW7VyL7wTWlPjkBtYh55xBHt40tc2/sBuA94mCczaVb50FtzovkBliVvpfB7kMrJkd+JoHm
65bHpkpTrUuEhh+CqHPtGNrQe8MjzAZZATEdNzQA42oohP9UtiuuEoK01zr02CL7jaiszuIcrgzc
eKVxsAZT/yOSqhRgK9dSXCydxRpHJLkWW/ls1A2F1bcuvnvAQfzeYOp8iQIfyupHIouvpehdBVeE
U4JCl04w39BYB8UIb7L9PabryeilxvliLLstlA6QsOgQH6Ufh8KeS/pSlsJKmQXrXlvJeVgkCew/
aYNH2bC2+KcVzQMvX3FLTXSEUDiH+J0K36JJtirO1gCo598WiLsOQBTV3mr5tn2L6RgsUgCVPEaP
r6Xze8y8QlwOYIUfKPr0LjbbTWd6RzsoGabgQgjcxGGdq0BAi4ghtdg3+5VmEP4eHVs3/smwo7fD
VWoSemMYRNlhj/rk1a/HPLBG4UR6IVVnk3p3wvw0hBHpQdtVJnuUKij4shnWP9i4nyWMjveXN1jo
v/eB3AZ5HP6WyKYm+SbRNqu4tMcdsWGYV093kvzZGZcvrSln0S+dnXr2z+hW4vlJxrpyzGWDLHs2
cLuNZ0JA9SiOZzhCpxmp81UZ5fHpri1N9zu77X3NjdppA8wcB35wpKp/tJQQ4ViIo4U7yhQNThaY
Fw2XlZCr8+RKU6NlqfuCnd37Nrl9wkbqh4sYB45lnJwo1UQDMZ5AxvIjf02PN7dlOu1F9PtxRmDz
ZimwBpRFV0FujX+1G9MGP9OG1BaCis6gjEHbQzXAshK73GEhLDC8Ht1MxcoipjcSjFssQPUBdGYo
xETao82PzXMzQbKhITAW+2ubYaofufe6nwYZME04yYKvSDLR7Jzkz+VNo/D/D4jK/xkwOSobEK/m
j+S2IjxUMfTInNNRb1V3oDZJ8VClGul4kvHq4r68aJefCgxessYCNNUsJ5tJdsCpYvFAi0YF7Eb6
SKtReSx3Ak3FvI1GHVRt9tOM/8kqedOzh3E7THbXPn/yEPtgNKPf384bK6N6YQ9xjI61+dlQHaJg
ZNLX1QajoeSafypeXIT+iw26EP4gMbnfPL8gVMQJTvPola7A+graAoUq9oDNaBFq0JkawGpd035O
2PJRrrp1eQvcNTNhFT990t65ZD0KtKvESThnfkUNy7jbWMI30DJwkMomROI3ADKCu202CSZkfsRj
660mZtqFK42vpltHFBSALDqSimC/mSt5CUSSHGal89AIS7wmH7l62QXWTeXd90ikc5bxQ9ZmgpJk
T3++MEoxAx1yki/jsvDX7yHVDVxEUTWpsItSVprydQfxB6fcrZGebw97wksVkP9G75nMBqniox7n
2YYNuNKJrobY6TvX+zEapPKXF6/+TWqImx8eRbXjtTee/EVPrByLCEikcbwocQ27urwNnfeVvXSW
iv5k8ubl30XCCOkl0HGW8QZ6SHJyoOZ7LVbwVtW2WWrB9jVS7QbCWH2elg+QZqHcaS3gllfd8cNX
To/a7pkI5W/f7WyUCr8PC+vXeQXlGjZ+BrwfaJp0ZxGW1YrwnFLYhtAHiavdml0DYlGDYj87wW5I
gTUraMVfOGrU79PmJeiXzO9fElOh/y+VOI8Romc2ETyB03wkyYDtMtvFZ3KtE7o+KmbY69Tqg2lB
l3xfLdwSv0rGxCEKaj5H7ixQdYn5XAwiO9P8z0yz92ayoLjsOlkxrAS8w3X/ZCavYzkxxld8rScR
pKlzMIONWydzsJQcqj+ziqZ8g/f+feUP/AVLvPxCsoqFulLv7QPgalB6tucpz4Llh2AjGyQCTig1
Wg/xVHYbemsYYjNwkPRm01HrknaRIJ81CCMFbRYlTkkIpHe65x1zbf9q3N+AIs1Tj0w0WhAaEvEq
XvpMYDruE6o30kjiGBGMrzMS7ztAxGE0bI69G3cQxaYTXi6ohlosMhz2SSxuxPILIHs5WsdJ3F3r
AcKxGfUl6ArNxe77j1HfUNglhNBXqzsxxgIwLdTMmbYDk+iIYS/uOBHSvl/0mmZopoB2C7B30i93
gUXvBd7hFUFZI43AclEncJ8A+H5IFaV3IEGAP5/RP8PxBHamY3Bl/sIT2j0PPKQ9owe7X19dLYUh
yQ193l9gogxhuu9yP4XhR8RMIrpwMF+9OqUe9nAtTJzHX9YaZBV/a7lMhkrB5Pos+01cE8purq/Y
LuxxUzWiXjAl2GYG3F8v6492bOVsWSfZm+T7UpUZPTttILLmp4XU/ME5a1SWyWNipYK49nosgBL5
oIyJYlfPTe4coAmMtwfFk8J4dY6uI5nv3ivvx0CwWqrI3RXtYl3E9eIYB3LtpCVCNS/22Nt9nqai
p+tprScLXR5GIqXv1nnu95FdWLFnIs2Rq1efBfaIrY2b7kXvkVN/fJ6UqP96iie4Eg/b9c3kunxa
yT0+LNQvw+Bf/Swis8ghdjOp//rfpVGTSui/wcaxYaOSiLGdpNJ+AuMBFa+Slo0jvMHtnFD73kZ+
5g0DeENes3LAwOHVLIPX8ozzx7OclazWMqG2xUezaqcd8A8KlsWUtgTrPsmCoW8m0aZ5Q6TXacUv
cagN8xH2uozAQUebSmzADXhC0TqoPlbz/jFC2HkXy9BBGl2D+kK/tacvLshisHe1TwYBuodiupmh
FK7ufginZ8p6yQksspZquNdeawnU0oKnEFXMbQQAlB/+E9YwT+uTrIU42fgKSkR++BSKmfL8hBLw
w3fVOMn5O0DkmbBWg06M8J3YNJMjl0ZQgSoU1yrG0UKFkcmZF48nFgI/9l5qY4FZeOlzbIsllYAs
lNp7NaEUJeWdGvOdOfPWeVdmbWaXXusnCnhqP+efyrxhq5MHosRUiVg+l65B+JNOzzNYoxHkIdUu
Ji+sAGbazbpp8LmQ+pnkdC79T4Wm2VjYDXuZlDp2KuX4PFtI2DAUA9JmtDZERH3Z4E7GX54ASbRR
VpG44VWGC5nYMSSg0P0ScpCcCFX4aGfXZpZVeH7kk09HYinxT4bks0SEBxgEMxn14sQnSnkC6Uy1
IABn7VeHyf7MFGAVgmO7AfwmzO/wToOb1aY/65slyNDJl8K5cQpswu9/yMolJazm0zDyCop346Eu
C9U1FxOXhINYUbQjLyPIF8BXdC1vstThEzocwb4FnRBGkpuazkbw0KNoZlgBNuO5Eznjpc3ME0Ls
KzC0g7PTY0j3HLsPMjyI/2KebYtBFE38lcPsPiocrp+f2AyTyClSmBEA8nbed9uKQsvXW+cNCBQD
Tt6Vs/rBsu2TEuhjLBIdCgrkFOqcHXW6RCFo2cuFXkKwmt5OQ/BIDHdAb50MdBzMAaMzFCR+rtPA
CskA12OpOjDIYb1wMmhpdaKqmM70jlyfdXKYfeF7OMxuKD37bkEiIH93Wva/WHvYRqmzyOFA5DBa
sbTVp74zi8blld4T+9XyMhQeFcJzqMIZ6OPzryy5QF25ylsoNsTA2dwbV3AOhjQunYAukpNOx0Q6
65R996CgM12kfAc6DVuUUCyWoiCdfbAzjzMHJVbf+oW5MrxVlVeJwQst63xSWA/jHr1k4fCqW2oD
U44c0DFsSDdT8nQh6lf+zaatNMYlANCeus6RGqVtLudgNH8WtvGUIBx/BufWiVW6cfu7sQq6YD8f
E0eplwZaZ7mttITHGB6F7go037pfBXDTHsxmzgBIuO9vOWBq2mImvFx+X0dbwqYYkGEqCpN5r7pb
eFVX6g4HBkrlT7n5o4qLMnDvtJkj3fHjVljaZ6yuZMoBk7b2lM2pZlh76+dN2Qr3VWHrp2AjipPX
ZHObySSwr27oFnI/3cs+oRztYM3qkCAK4jl6DBGfc81+6rVskyrJbnW0hV5qVni5fOPD0OM/h9+J
RigrcdpXXk0HLvxKWE7yohneaHabHwEmTP72h7qhlhiDCvyv4wfslz9dOaDX7FFZJZ1K2d8FbnNo
BZZcLRfa5D7FrKABhwGjAELS8z2HOGlbZwVARchUT0HjYyUlPIXNYuOKdMfZ8dyjTItItImtmW6h
9uL1X3Vng6qjDAEQcd4PLjqdXr7MBJ14mzLw2Wh8ynQCvYdtRv77rl8JOp03t2IrSASJCKQJ69lL
Cx5FyQ7pox7aY1w6HdNpAHZyNOlm8+EtB3TuiyPhErBPBZm/LcNwRV0EpcPCB8i74gzInQRvJTwU
4KSv9YpEPfbbgU26gd5ugFdGkqwJVAsusQVX0d2Ho9xue290rNDoESBuoICNO+NYP8IsNZGwSo69
5Ukx0V+Z7lUTv9UA0WTONyzBYmmquGN7iZIFeD3AZCxmTu/4zEjEc/og/xbhOXowRQVpuDNfBo6+
5XfwOq4QjgE/K/zR/a5JG61q5Cz0S8euhICmcUpn48qpIvjyWGZhUjlSmf3TyKd/k6EjK+HPbAF/
u/w8OsjNAC3OmsmHhkE0sqEiDjNq+j8oVxW7MEp1TrbhT8LP1ipwA9isHG2ez38W/mX4wFoTf+nR
AG6n6pIL1LlS7xAubtr9svtIdp9TYayPHV/G37yJzr3eV5Cy9DhmfiLhaUid/s6ldfhSTjiunz7i
gg2TZtz+wFtM3qnAYBRKYzv9NYUKODke8FyPJAS1lEbk1tpS3bYP/FZfRlqITcyGRXVHt+zNT8+T
hL8AZqk+yiAW+oWTs69xTIfHQCZzm+G13E52+5HU0hhAPOP2URCfQ7WGMS7XWHFSUx8eRbZKtbC2
KP9Qqts0nI7wkxFs/kMyyUarp+YyntI/WnfvnigE0tevRhHhGLVLmr3yjRZ+jmSttHjauaDhnTCi
mbkrNnEwy3f8Len7ItisL7ETxk+DMPvPPE6bLvOJnQIsIKlAUu0jwDKzVy9ACDRYP+Wb/Rq3yOZF
Kn+Ihj/G+gElLQOCymjSTsri16CBvQLykL0y7Bab/q1pwpu8KZWpsKr20lwF68M8s/ekHdWKHnId
LFB3xeIz1T4Lq5ulYds1Fod9a3GmCn/bMpFfO56UuzMEBVsTEbQuW69kETiaOajvjQ3flTNQv581
vPIcf94UNVF9iuOHsUbXz+C0mIcqFQJrFTmDXtpUNi2vIeSfOoqAmMX+ud6zFN+iUM3FrrKDf3Gu
VOCF3JZ+tzxDEcpfP2/iE51rhHiHMXNDm6w4xE5TaoLdpzXn4ks4eGK6OCmBsqATNDLvIFLLXoUZ
0GOdP9Vong675BIE/eQFO0NV8bjNM5HX+X6XGElI6wZVzYjTWuoUpESDOVnjTGrmlUYFzUBhgDYT
Zrs0wuLAvEIWImUWd7olEPlNUyjJqq/x+2NKjROOI6g6NAtBeq6jIoKi1TaSixt/7/3c3gv1Psr7
4KN8Nw2XNVhPNFgHTDc/b157IbMXrWaIWJ/mbpA4YkfPBjQKXd8uA5MTIOwuYjxgWwgVRVb5K8d3
1BTccHuGcfAKQcdTwrFA0YDNbSQ5Y6YJudCGevFj9/JMswKsaIUb5LU4rc7cjuAZMV3Tv/NtA0Jy
6sGvchwj8Ryb9sBhxV1ihpwn6HAhHytk+X7O78rFqRif58bcogMMznCVW+Yo5kKxWM5/gVInJ6nP
2G05fWeELh9rCaQCD51mNCGhkmOEj5MC2c6iTg5wK4+JPtsW1WGR+xuHVJmfko7oGrbQkjx0Wq4N
2FsZugHG6GeL+eAlK8Bg1L/zQApGssx28hwQYaxmg3E3VvXO0nwCTRJ52m1b7EQKgtV04/KMeL1b
8YSXA2r9/RmQoowYo5NcyPxfHCBJeN9AlJTBEe0axro4lX2bhpXZ8YLLUgB9nR6hjjUMCO0oPUO6
DX6bkJpMqjYV8OGtC4AoeurS1ft1icVp+hAjC3bLt3xA4pLJf+YDlBdSXmng9nYAwfka5osV0HU2
JTbxGur7gBPmPpvUwP6njDwkqxfV2jlmir4XJe0PKQRr92b4C5SejDCGsstqPTMFpX8K04eDWfAv
NNpJb5wVM/GR5a6iv2AcaldKGp769/qfXa13wq2HIScSR2UU9gviBlRLxt4fU7kiX82Y2fUpy/3D
TI08NXfEfPg+fMpn/y6Pjax3qyTfxWV+tFxday9BCrf7+HG+YDmz9lu0xqxbvYX68hTfLVIiEaUk
OnK9OgtojkH+/gvmN4qgPVkdTalHQUByCbFCWO6kgHNAPl/vUJ+8FUPc0zKZ5CducvEqPdNJR5fP
+cb9CaoRBAYVbWrGNdMhUjIVZPZNaKDFDd3hDMlgxiSciMjeQQBiE5ihtdLAhxVrjUphlaMh0SdC
JxL09E74hpGOtJ3PUDMTopKukueNPrRAT0oHdR/hi4LwJp8bd5zcozaMeaiuSkcBfRxFzH/6K5Ph
QcIHxJIFj8mSGtzHVIl4VOhVB/GVXkoJi7O+ci1CYH5Mj2R2gGgKNNUZ68/U8Pf2jYSyk0rLKXB8
+egbcGSF4Uhj0bmeC3E621aI+IzQHYstu3zpklP84/4q/We2oYbKD/brp+qNIWUG8yL1p04nPb3D
6BtxnWfkOUyCjppO/F9+5YV+8IIKRpxrzCL8YtO9Ri4lTmxENI3zocKlcM6Rw6PbRAPHNWCevRPu
dQC25duEtrW3fnKbcaEODn1QDvCuuiJvWV7l9IaDo3LMcXzQUuixB8z+lpmsi+dkPIjaG3pFWSvd
OkerrLEB6eW5UaZdrxh+NESkNrX3qxfSvLA9KQevBvUfDxe1i1xWL5S3FfJg9QRGKek86Xo5XWpV
Yz72k5dgyofeQUWXx5h0HrNeWBO2ZR4PL9RkLOcNirR2G4dMTsVTxc+brDp2+P53/ZS6XpUth3t/
yzIH3IfzSb/cZIbBYz5yjtjNFdWkA6z8VYz7UMYIprO83/wAeEQKESNQAvMwNoHCRIvb25WYL80C
I3O2IyJhITPTikHtNNqwEVBNpKI+KsEXnnAT7hb0Zg1LHe2wjqn+irUYPyeoQVpPWK2Qg12+10ha
9n5l/az2yWEv6SbJXL+7c9r267W0+LpsX1lTxRZ5Ifzo4YgZfSvIkAkrx7Jv3tfTSZZgQNl0pDeP
uwl+ylLZfFbeV6urb/Jv7r6Q7Ichf33bNX3a0YuRSgtkcy/yrD9GeAKELTKDP2DmypMsSLp731Ng
zHyUEEYfRdr0dDdSIUA02grdSL1NEY4JdNyVqwq+KzTzGAp0HSdg5mR6XitFl7nbvoBku2rrjS4x
lDiROpVxHAyVIhjYinVz+5UCh5zy+rxxMfgk/9up4KhjG720oi8JBYS5JpBH2yUckiAYWE/fiplB
h3MbEXNQ+O+cfvQOJ4YGLy6iucMjAcyGqTjPtcAwNbphPu9snjsrIHN6RE4ziaPzaz0h3jZifRF/
lnTH1xBO1hkTw7VcIXouSf8CBjBbxbHmXLCBcD0EF7pIdFn9trNQqyQXXEvOWwGWuBmRZfznlxk4
q7lfu0WG3kOkDmpgPJuXbQVMHqXpsenHoVBuFwqe+XqkMYz/+IGN6prGn/ewxXTVa2wQBkrOrCZX
axzNoCHJhva1hUphz2qPuE4HHXkYvUl+z5X1n7fnXgg0HuFIPpp9Pitc22OrFafC+NS/Ssg8cR8u
UzGb/tDLPbJktqwvTQgoxm/etFqj53hwac3A7sqfAgPvyNVcnEGtET+oDInEDhI4V+5wb+QkIzMs
OP5YPL5lwt27yL95ERXd04w1FrQk57LNGBwXD3gezXk4edG+SBWv9j59JxhE5PqwGlnrr5Sp20G4
Fn38NWcb63E1/QJnZXgCChIaiR3v5sqCoAaZA33fRzQFlS1819Tz/4enSJiKxosfsN/ZGQgymPu8
QTJbAFtxm8eiE85+EYndKDu8SDp6pEU2ItvuyezgkrY/barCcJ+uC9rXBQ6KTAX+YpnFeF/F1Rux
gE4SiqCd8PYi9MliPsOtn6lVOMWEzI/9lZVJViefDFITmW3hzPwjLxQPal5q6Cw44CaqVuZT4QeX
8uKBtu+twC0p43Rx1Nkm2896voJ0rVfM1fDQwK6K5sQUNK7nuz7Ow+FrulAbkNrIS25fxFHz5o4L
5atOfzQUlDK1pMLs7j20r49YZ+rdQWcJwpBz+CVOv4lE279e2Hiq1qA2xzh7eIUyXsihs0GrmN+D
5W8mMzNvyuieXOBO5DIBDhJUhYT12gig+d1aXGG7JEVBXWAVwT1yrR9fFJDdy7cno31ZhVIgNXLO
36gUCbLs1EGbxUO4luAuO5OMEQ1mdSUMxzf2WPLJAWMi0iKgDeCDkTXbXSKREIHurLX7brktw5nf
Qxi4V3KkLM1sSbaVh9hiJ1RzNtKnU7JwSVtKObiPgok8tleoGCeBOQ+22khHSSiuy1jLdgtSS2qB
WFE79CoaL2XVrjKFMCQ/LbbtwabdJoucBGwyyQ5y5N/yZbmRfZlM8xYJBb33SSVMjakJZ5chrSsi
cRTe0zJFzObG3yS0TRylqHMvR/qbaq6v7VnqdBIo6AMPx2ybemNK6WcwNpf69OIefDUwdofjLFo4
Uj7x/GDREfW14C5VER2ITtfHqceboIVRS/arWcKh0em1VIY6w65okU/nSMAiaqr4MDV7Uy58REF/
lb3X421+0A12ejEh5JPvC7RN7z2Nrt1lR8EoyXMflL9+/nj1feO6JmsVIWlFhssH0ahyx7+m2l/g
agwwRaPQGfHOVLwaoR7PXF0UlsYayEuiLJp3dyF71xyEVuU+PpQZE3H4PbfPRlMhncfKbCSa9SnP
iTAXAOgtC7nZIR9bNcv51yNzXHhaoR8PuhiXzFYt9kmZJKHpTDV1rXwj8XT1SwvfH0LFh3TBQzWh
8T5309VcibpPl+h6nhTyQ/rJGnV5a14/BJqhMem2wsSdq25mddRHm+GpcXH0Az7P+LH4GJ6N+zhc
EqQQhd68o3V5DrvjnPEXscEnajBet/9rbx3+SrIU/7xO7KBsjLr3IcFsrEfDGNu5JwJC6T8WsPrm
lWwCG3DPJd0/xbJZ9eWUciEuHM84X8sP7Dtsvx/S448zs+UmWMeRarYaVyJeVISNS3H3RqPR+a/T
INDjYB/Rcg5OgU8xrDcWlV2m2xRnWrHfks/48ENPfhmU2PD2M/4GBJ6c87Gqqqt0H3Wu4mHtQS4v
oVRXPIRamIDBCBa9940QhnXJ3ZCXUZqYiFZkb05Kc+wcs2d2EiRRBqNCtqCtaXk394N5x4SH/4DD
Z6a2it3ek/nSQ+ES7uu96N6J+VFA98F2P8Bht1dNZVn+/993LKGl2fG9MqQxF3nLIZk1VYq+RZ+x
HJrEQeM+Lk8Q4jY7yWos+6M5X6kwNLTnCLmUA16hOAbs71c6vwzP2GBXUmZ9lbiFKCHyaOoYJCw5
omzTxX4Tbr6Qgb6jo97Ce1glTSCbkh4wOwFDSuEmmxGD9+C/+t8DC+E9GEE7oueL2/ZSpdF/C5Lb
OM9mFhqJtA85IQI1DT90oWPRI6/HY0rbzL/bgYJ9CyLM7zgxlGHE7SlDUhCEjfRC5wgC7G+7OS2q
LVoI+NjrKfjFYGHXiZ+8ogIooDV3C/uQwqCYJWY8a1apDD4MDwBuG6JWjpDkiGHMTBxTepJLR9rI
PqFRy4g4rlUQoeuhiSatkbhANMiGpKpxArb8OZ/EB756elv9/Nffgzi7VIAIYvxoN6E8IkZ2V6Ws
BtSP1ABIoRDYLkKwj6964+DFRmACyMBRliNZD5oUtNrrjSJZdcI3OXR/yCbM112s4k6PFCdKPJTk
NNPqoW9c9nR/qpH2veDTx99fwnmizXNdRPoufKs7/NhQSwQEM4RtRenBAlcazAf+8Jw6mEo3QOjI
mmGHQfE5N6KIaw5p8/62U7cV/89JpOOSq6qXgxRVMISsGRLgIhrIWSQ0bKledUepwLm18H6POaT4
IIsdL5WxBCqQENvS+lVObWqH4yeBj6GqDJCGRaCEt7JzsDizbXO50narxQwGmRb7hNN+OMzrjr9A
+oze8OCOnudFXMpDnF6uOA8eW3XhivzC2iKueahKXpRM2QGX72LVape1aXJ6mqbbOxaVapN6Uo/T
NOeLGdsSMDjydGgfdvC6VI5+dUngJM2dUxtrMgbK1/VzcDbscuIhv4kTiqppEQPeQIIIrXKc7nrh
0aReU9MhEPLO84LBW2oHMTXYnZDtv9KT9Mybz10gZldvPYTMX6pNM2J8kPXKCIAV+YJrkpPT5/2B
bSVQsqBv+4fcPzcDDFBCK86xvaXSoZZ+qYXsKBDnwlwhKSN7tSFcHc+p0ey5M619mbUu2pp6D4Zu
3FnAH/UvqaIhe0dRiprKnohAOUE/WRScOWHlui0XDT9QZhw5dVBfm1fqVCK8m2oq6CdLNCd8td8D
J1aYL204pw24FN277F0E8lomEnttkP3YAgv7NbdlpiWEiGiLooDli7XqquuNHgzD35Ovq6SaQWDU
t268Dw6Imx3ucEaL4D1SwHObCWY+qRbjzqBDlRPEuXJUB4chJKcroyNLJ29yO1ShXkjsSTXvIpaG
BfSggYQXb7pI5vtK/8goAVCyou3+OMsGM3aqoxnz+F1tON3LNTtl0XGUZWdd+SEphXdLrZIc65T9
8AYDZlxPcLFaVU3Ie9f+jLQUZ+OlrkVUgpSqNo6VynIXmJlaFUwE/Egvj2IaJiaJau38Ll6OLpq3
yJ5OCDOXxNfShJmyeFk3k4ums5CT4ZRTCtr/lOHERq+CoCh1cB4yc4VlOysk43KGkCdsS8Z9KRqC
To6m31iAeI7mrWzX5Orm6Pq0DsTrNbI8u6b8zMaieEQXVvDCN49gnKahKe15NVHKXDlJGKnr+RGc
2iqn4hiqZ3NFb29oGdXiqHFBPbcQWT+feHw5WonW+1DzGxOmCCHObZTyCKI5+NiDBMms1AOMwJHO
QJ89YzYrobXIQr3T9ycsjwQqCOnU70HPUGJnKXD1e42MV50kkH25taQny89VyPnAVBe+vWJJYZ6x
ac1l5PHVIHe0gUXizWlyZwiavnEVr2sCZ4en92ev/n3mPP9cxc6agRdUZuK+deDAvZB2YuC7HGjC
/HB0/XUIm0Uj8jpmi62RrUnZ3p4RdjOfpp8eTitNw9o6N+Au4dRBicF7Yz5opEe9Y2XzzjVWwYi3
crr+xPA/tvVtwsSnPjf4ek4TecM/2EtFwHqAQisMyMWWgs34F3Tk1XaHwBMQWX71phCvNFrepbTW
OjpaLUMxeJBVmV+uMhCAtmg10gGHzGuWoXnSAdMIBmtit9mq52OsP7Qq9ldl7BQ+HAwQrTEncYe3
VqbmCTeVqkOYYx+NksUUT2m6nOrQmgLZDqhceaYMbyxPep6sOLC445j76FpBm0Mug91ojoDfW2SZ
sFZAjhdoyrT6ZePDwQ25y2/ULheYv8FesY7U7jJZG/6sChQ9YbOOFEt7LWj6gCXefXrPtt4LPu6M
J56QasD5s3gjUuNu2A+mcBndmm0L/IFkNeXNcaKX8YLWft446JwVRohhyrCkeYZzPvcvWxeZFA81
rM2iSi+vaJ48HZsArmYsfIWLj+jNhVc4kCEqAt8cr9+N/VSAbvx3BTChatLrkmUDE7gw2ovb7n3F
16O0D0Ujo1ugfQOm3gFxTwJoFpxZDihBRFUhEdIIPOy6q2KGM3pLs9PIDuMu8p73kO2paklQIvF4
bhWXAZBhBKIeObqYAbQty1HWzwG4lC0qeRS56PqJSuEJ3GwUYXhK8xdjII/zBssAZmQqwp7qNyz7
ki62wsjKuKblB+kyd/sWXVxm9vUxf1WjUCURvU7DHjsvr4JAgQzAHg2LMiIQZDCH7alEzgGOCDYa
mkkBH1PidF6vj5Lv1XbJEboEanE1QJs5425pKqO1QdAz91XHd2eOe9OQ6QqgV95Cc9oGv0r+Jf3R
gKFCyBBKjtbUo5zwGnt1r3TGw3AjmVAU3SBcGppGT5veKtPPjcwXWN3KIBuKU57GLSK56NFDafBR
gvDXKHXs1gnziiRtc91BV/rahIA9bVYE1n/R7h6t5WPh+8jlOsSBuV30vniTEWjSepjjelYwfwMb
7PKRSLTPwL5khDgppSWWfK2qn+4v9XgdNif4Gf1B0WOAyWdtM1eUqyK5GM+HEyfdtHTheUyCQb7b
Qac5i333OpyLOAssKGkdgzfLe/rtoSHysv3QiSRstfdDNQiA+tFuIH46NNmyzQfz9sIFbF0/wIK+
HAlpxA8aj4boAruywWOuriMkHzAfB0AJg/x3gSw4248gvTwDGfi9XbcbRpJBiw+V/Nv/+XOkqVHx
dnXp5IOdzsG+v6FN1GJdv2YHjZJLyF5JBzGugc3oN5bQyW11GUBSrfoLZs70LOpdPWVLZ01zIcR3
TBRtV6gkosPEDnTtVb/PbDpvfZDhO3h6FxCCRs5QGByyqKRBL0W2/icJAD/CFEMDcY8OUH1MbyX9
swcJTIQYN+crcieIbrgQIim/H4FOCQxsLvMrqq1qRXt53Q34zjDWxClQSteJ+JDLU4DAVaCyoxRJ
26RPzDdY4+o6pbq3pOzlYEjEmMgVdJKJztcIl6jTJjAxjbExe51D1YWExaIEEGf2GUJ74UUUNbez
vSlO147ZEoKTXNh3OB5Ro66U7xjKCmmBwdhIZwen/0XEfbbsXAcWQT3xhWbMgpjzYuF7w0Sk4zNv
wcfENf2gElFpKcF8KBrEGUz4fu7uMGAN/dptajCZyZ2JVQKeAxBQHSv28DCI8dBeBMdyuRVWgVPB
2mLJKb21S1e/9Rq27fTY8/Ka4JgtlGG2/wOrlulV6T/8waqFikA8pxptsDVPx7uE9870Xq1ki6qF
XMT6JsHWix+L09RP/FYPMOGixLX33DfYREifqyfYjAdpqovEAVIqZBHcRFtfd0ZKLGycpRngwCO9
GoGymIo/2VOp/HxosuKGLx4eANsv8j+WiRSmZV7n2gqwyqWwKHrDRdcIpvfCTa5ZuBdndHEbOJ4+
Bi9O5c5CWJXCvNe9jJVtFJcmTDstDsWuOmFGGfEKa5lFQidqp3k9t3y9lteIo8Y1oeCVVVFog/H0
rn5+T9vr8wfCoUjXNrVpN0jtka3HYqrYv2CsIDH+6darVqxjl8maiz3ljhXCbxwB5egBTL66y0xp
UlmeZYgd0LSujBAOCZu9Gz/ak4cN+WUA8JWZKA2arBf6fPgZfd0mLJ8yKcX++BKnn4yGes5e+maa
wM/OMcmtl3JyzMzaIY0DN/Ml9xgOUa1GCexULtQ4jUIPpytMLJBOji5gNlyOqq6oCedCJjkL5NRN
C+bNOoesk0UIFEUzLy6gCuFErSxOH+5Aj1h8GBdXozXs/2R72bJbvOCevIBj7RNiMg8Nq29EHJ94
FIt0M6XeGBOJIa4hmUjz4uSwBpUiVbYd/KEjYv8TcGYqfxWEQOtl85DA8AiWf+tHf62wvxnpvh+K
wwXNQS0UMK1XhMoe1K/QWlrU73iinGsKz7OAQExXnNC56CUXDsCgzWrAu4OhLLH2ztE921DIJEOU
GHvEbmLSVfA/EwQq5vj/RsvvF3/B73NFHl2jGNXTlgOyhFdNoAJ16eXtUCTgBh3l6GMcdKdoojE0
me/Noxr2J8g/H3GnYYTL6p9Y2qKZ3onGNgeqa857Qm7PJzelFW/dCLxH0ETMaRhyQeGLVvJ48mgT
/Wkaclx3Sn0YLXieKkBcGlGg41uhesLkfO5j0uI79n0Fp4UcOaMXE9Do0vZZ7Xburc94MRMNTCpF
BMVetY9KbDIk4xdVX1KgiHstNawE3TWGm3RRIQUq/QK41zn53W41Eb8HvSsL8M9XVRbjHjIkzs/+
g6nKPmDhljxh+nFR9paj6b7425cZway+S9g78NAa2plN3LpziAaE4O4PMGPYvEdRug6P+NtY9NJk
J72bzirXKTsDaufHpGa+Dq4uEhpuaxmXHijKJslR0PpI4SiObYMfbBmGJicHPbLLbXh1IfjJ/iDO
GMXtPDh4fxv6dNMSXOgkpsfKBGhLvJvi2YrQMHQpRbR6n9hi82qzyl7Z/xTUSD5DmBcNMilWrve1
84fCpzFt4p9odeQQMeRPGmVy7vEl7teMajpIPhlBoIXmQ8bwH36a5DVCBJw9Es44ZjgNsd7c07n5
OPEVXR2RqzPIrMrWOEtnw75uVq+RKv6UPePtDMLWL8F0xG6ZS+Jlm0ftCxtahxOrrkDUalPr3Asd
4MxsdXkxJ/Pk68BnVkbNgKVvb0GDcbN5VXSNsVqn3w9OQlYvqH2fpwNxlAuqihdzsJzZMaeQg8Ti
Q39jXPJitjHmUHsJMYDOWDo3b7/9PUgzmZKkgLaMi3GZ2tyKPlIveG9JsXt5cMn3CVqylRAaA6p3
YgA7YMQoAYM9PbuDBBmQS7Pf7nAXpMVs+S5IgWVaRSP8cDZUT4UvYnK9bFz19b5Adu9iih/2rR1N
7YNggYYydNTT7gTCNGqkXrAVDHP/sR1x5CDlPjBFZ3elLopJ0jzsQTX0BOA3WkcCUr/3Yys3UeK+
PR5iT94iTnCdIgCARomhlwKN4+rTa4V+CK7fOY4H/NyzhKvVbAJUUK5rXujSgzdJDgX7U3YynvyW
4+jZqX4436lQ4gnDwHQvgDgAl84n5oAfSUrj1b2J0QB/XvuVvEfqtEAvFdcAhWG6pyhqI0ZRwPJ2
2pHg66lv3Y8hDpJh7kxH5zT0r0zgVyHVokYnoxHd5MrwdA0jxXadysLde8Pjv1R1huAcJ9K+Rpjy
yeoeUlxUFbNDPouAMA4XoSAin//v8rqU1ysx37CLuKdHrYwc0E7SgnIQiWB1053vkWNBcIPXXkYO
klaOWQ3z/1nrogwbr89P7V50VUzTYMOb1Cq80OrUFgtUrTkMx6g/9prBsabZ4CoZwrakWDpqd+/8
N+22+/W2jhC/hlNXMew56AbkTVxeZcjrQaId4z0JnMH10R+KWk1lVnbnCOC0Dm5kNykJK2CFUglP
ORhU9g2qeNGpRkSRT9F86pD/3uok/82TeGkxy+llf2bnaGyjqXWW1AHw301wgODsdCoaN82NczeU
r3obxtnDDR8zWwkdVGHIM579rO4V0FKu+7aWLAmy3/fUjD9eKCfeYjG+fh26UfHxGnBMbEIU5eFR
1LTF0rRIMup11h95D5E0qHUlK/zC/Ua4RiB3CS1BF2dGcUh6eHg6fmZ66bzAukhPFWzc6ItCuOAK
HuLWwLPrFDKgi27TTDOevxfRRIB22tIlCAX1qTEFRvIk9BI61Q2WFg8KZeSy68bmlm6F8DK1ieVI
vdIDpUiD9CARJVGIj+ZmpOQD8eTg8PavEMj7Gyx93KTZeyVxZx7JPlv0Sc2JksA0dtLCrE/QK2Lk
+4XWrMExC5Use1hV8BX2G9wzS8CEF53aTCorY8yC4vCqmwOYhuR61wDv1PhJZbnqwHKF4yFZTvcI
tf74sJTFF5rPUEAd3an4Mt6WpYCx5mLrLCoHtXzHmUnt57Ub6AzQknlGAzBVjDOza9vGBSG6Y1Hc
BzYU0iavxb0qrYyPEbE026YLsStmQ4zo0Hh87KoB/wwnVUuyiWYCRGwJc2NbMGHGeO20vBBkPHQw
iT86gf+uPIsmHMLcyB9kdEP7yWlmTw5mPFENREjcY9VSNAl2hm6YwXmFbo3rt644Z+fQLipWbALB
DfRnwqTX9yE4NCingChLxFTURWC+CCmtk+qx1hBUl3ywzVf5dI0rLsi7TXcFLXazgj+/Hi38wZr5
J7OaY4jH7y1K8Y1eO+GK0Ru3EMuLSxMVtopSG/CGWFNCCh4z/BBkOn227/uMZQd8iZB4wuhc2GxO
JKcY5xs3w9onwpucpXVGK8+jpgIFGdjC2HCCEUtPF3238fiezTUOTkdhfrRdBnv9rvshGtvyRLrl
DW2qWRlkIS/uNJA7yJ6d+IyrzMETS1RqzPBt5OWroMsblSWFXAAhSO0CGmBjEEgVSI4NDlY5Tk2W
vcXlecY6SZ+2B2UFG+cRkqHG9W7WKJnRg5rYEF3CMZMIWSAl6Js3B5wM9tqKztmZgfZ3ISVBYIL3
w8xDnD6ZO/mG4qmAlbVCDgiTw3pHMciqU7rLsttMdOE1l/eMLmEmi7Q4wLzHscVCOoG6VdvAAxdO
mOQFXvhvk5GmkUH42lVR/y0bHJcpHK0pWZ83vptG8V8RKkOh3fK3IiEKgneJT/kPPsJWNAh8RQVz
GrE3rJ1lRG+m2b7DNmjcUVvtIgD/p7A5PlC3BlSkFYaTXQNB01LeYZ71CWFvooMRgAyLRbv1KFxY
yRCQpUuerp7+pqMflUWm9dxeSFwur/NBT9NUprtqzWoizpC+RTbu25+05n+ZmiLmTnXgWPRaE3hU
4A7vpVllx16pX0n03uUD94/hsI9H+pRqypnzJDhqL42ebJzNKq+W3BXdnKWlefJPA1gjOe+ubOlD
0JfWQrsHSd2Hsr25HvaL9yjszQccOdz6R9YBziPEYVIt7nUwNsJm/0QkutqOpS5xbx0OTdnwBNuG
03lsZpGGWceEzAKogS1sWZa2VKfwXa7Z/mNMSMzDiJuujLQZWMIvsC87QutB66AawD0sXQqJ8hLr
945WFcGzk3E9Q5vhWCmiHWrWSuOBCs/iDcwY+PH9z5VKg+2WEISN5f+SGjlTr36lhyE8lPC5l0ly
+ghEocoz9NI8EbQZ8Q2PAjYxhmWWRVPUWUGOpLs176rV9bn8ffP3EMwPvhy46mww/3g/AIcqo7Z6
cAbInIk6QzATw0jS0e0ER8s0sTgI/8WHPfgOjtXxiibO2fRvfW3FEREi7M1d1TAYKnZThmAXNgGr
gKiQs8Nz5mZVZFVHDLH46f5xYzVfiPRfRqLU7aGvdsa8HQXA5O/eu76IhIe6XtkRrpbFHyROn5qi
foiuJrcTHaUuA81YwDBkJNuzel7LCIExIS8Hkd46/7f5cmx1zn7GLQpP6ElQLQZicyQRGRiucfPP
hoOsFUB4RFLKJ7TX+SeaGJiqj8aFurtoly/+pwFEIJsT5LCZebq6rlP19RVSITNNPjN+IXF+GaUg
SGLDMo03g/c6YaMil+m/4Gp47JHKfGyzEcHHvBIz5V79Kemly7mG2XO+bdDqTytt1vpdpI2OaMHr
PnBwSvF9A8sldQyBbSCJpPjrXXWE/EQaEycGQ+X1HLuyn+NEFtQWVbTgveARzekZhYaytvi1AI1A
OmSDOGlnh5FMZqldzwL264ekQCzCKWByQR3QTL/6UgkdRHiTYDlf25EazEvLXTPHKnUknfll0iZ5
hDUNpuAxmPWog4hf2HzjUcLhqJke9KHmNmmEUyIXHfzFNEInpQ+3+WeuL6HYaGHGP5Ym9yWO/Di+
GHT1sVddU53dM1wZYSfOshT6gbSqT+aHKRlZ/3XkyboaLPjWPJcH2rs1PDQXIljAfrVDQLwYG/TZ
dVQ9KvmEqtLPENKG9HkuLFijOw45PD7hr8ueRyt6I6+gZ0/EFx2w4SmUlpheKloMvrerLY6uVTDY
GMm2fHRhqnXKqlXErHhfcEneDcTWeckT8NIz8DpvebRTZ4ELza8rI7VHixfk1wK3aKdOU5o46V3A
fAGHMPe1inaK5VMcpKopEHjx4/JRMXDYpRdi3xC7Wkr99c7fqnd5Prko9T1VOjmUV2qMfpvkVMlp
jSk6dPLuKdEIxFjD6fjKfeeXMlEosZIb+6WPNxXn3p9MLAUezvs7/50EXW/sEvHWYtnbCp4xIKgK
EqKhNFekNGgCyOZP0zPAzWnZbXVT/oPaYfn6F9ekLYg94/EVIlNSi5ZFTpvx4Q7fbzeiA7URZXMt
Ku1gxepvf9SkGzh+HeBpCJHIRpeEWc2c5yAFi/MrAGGlsiY6hVmlfGC58ZgvSPZdjk8VdLlBWIwG
2opAIkkyRsIat2dwVbWunFEIc9LWaShAjJzOUeBLdk47NToRUG+3CXf8w3Yzm7j5NRW0P0kEl/S2
/lM6zUTVMDguDE64b7Uju2bE4tO+WjDIBWT0wBb9FpFy7kZ3y0IL69XDefOzuTaFnE7O/MLAR8g5
673SNKqpH/bDJ9Rla7zzPxY5r7X6cMds7TPFM8GuypMP7BpJj5ri5R0vhVArBFMmeCZmOF4xk4Td
aPQf/clvcfQ79vIdZ+e0QYhcc65535T7lr08ZORa08R+ncNeF3PvzvAlvrhIhf6zPI8Jiu27s6f8
pYwNArUSt+4cLhPIJfYorpQuO5j8WcJGNBlr4VLkmERXW20ZtzaMt519VjR4EATp+QVbWSnloahG
M7f6AxBVeYPMGm3jMQsyGg9dSEQnR1WQquxa9TKwmJTW0leEnE1nc1E0VrXWJzrWtbK5IyQvJPLP
6Bn+nQ29baX0sxUt8+CEW2Y2voQe5S5JByc6elx2LtbErN0DXHHNvZrTwunBD1/V15DyEp/8uL+9
2D1ji1Q3htQ/3XRLHGsJ0YWx5cCJPgFDXdNxhYDfYwgT1nxT5l4+bAZkAzkjAZYx82a2glvepRvp
40JRxV0lxXFxBPfK8MmKqxpohbd5fvIG436w0wm55T+X1vvJA5qJw8kV2wTLr1tA0ogdARQicNpA
R+SeW8Vs+nR/spHMDi7fIdqqACDyx5V4VzWTWFm8PgGbvMixMAp2RgTBOJiqeYHUAjCPQY3JE+Tk
uz39q5Aw11agzk6l8DUcQWhgXcSEOsGw1AW+ncbeydarXQs5JUQg0WUS+O1G7571QTUfGADVBcNR
UR2uyUF1RPm6YrbiyKUBM0+zERg/9nTIkGaPIxSDq9EdpwZihET/qIpZ7z6i5FueLNXKwNzFAm9i
96sTazPWajN5HDheUOYYM7koxxqJ3Uiecf5kEdFhDW1XzIW4MVuf40jXLoJDgLoqd/7sJKJK8jmH
rQm/oZXrXnc/knYlAUdnDNSp5Vcsr9YJQJRjWQ6mgWFwP6sBj07VRILR5VADkBywSQT3+z5u1uXV
yK9W09wIewTljFYhQ4lrQDOk9e4rs1ZV1NjL0w8W7SfpB4LOdD2yQ6NMXsQCwjcoA82mxlnWZfmx
j3F0jyVUHRfy6eMXMcs1ZHNFt1jvxpqcKUC6/EDFSB07RTU0fhbrrfQx3e10M/iWUNPFSvjOKoMg
9lvg1Jx/iP9D9MbkQWag+9zjVyXbhvDZULqFB6zvXSw9UW31MM/bcJHQWRoB1UK4lNZeFyJ2tps1
NzPCeGkB6uBdDpR9vyese+yHUvImEOCSoCDdv46vaLo6JHWTZlDtSG2x+w6oOtLKIyLqTXaIpbm4
t9+/oS6QtwvQnG8sRCReemImfqAlKivKdZXh9YoinUcIsteXtQ1VdB27tarwLPv7j6X3If4nrmQ6
o5BjG4ItMOxntdZwRIRtLb6P3w5P7SM0g0gKW//PmZIbdv4UFinEYOr+JKCHSN+8afK4p+b8MzoK
JY4wL8InHwoosSYQ3uC3v7WL8X/UKpRJ63jIMp4IgVw7xSpUBOlfQuff8AixCxp08YdzcB3TpPU6
KoZEFT9I5YFBg18TQGzhVmjou4w4iKyMvJsqV74di3Rpfnf0652ydvPuCh/4mkSlyG+T0nqxhwIb
c9YNtp5nlsfz8q53cIiDzgEpVUB50ncVf3VsJC03OHcUxYvKluT0io7mU0tveb50kMBowzqgpFNN
6WYvx5KLeTkesp4ctmW2kF+68A8gL6kyB2MAgxup2Oik6M3y89yKsfP5t0ySYkzDK63ftb4AxKE3
cM+2erbPdsITf69fyiHueV3DDdMK7JeF/d1iDyieH24DvKJrk7c6j01gOK0c6NO7ptjZNjRp62g9
xkxQjKjRbTfGwsBOv0kUUcr52o3L1AQC3nIN790FRzdwtNeeOx97ia9gzkp5RBtZHF96gGKQIJk7
7SuFBEw1ivzdnjedhD/eOKEYmdxDyQzeaJwUGsEHAADsSs7Bf2GVIhOjHlE0ZpnJSwUhnevXAvFf
okhmpaX+ChMKidrevhpabm40qd74e8D9Dtv8LXab42OGvL35a9i2MRxUg6ESHqdzZkc7/aOpgJDq
m//ZbyZEmuygFXhYanLJaHpOnxKmAJ7M75gfCvjz4kPMakGOx6bjAJ+U93qz8yweBazb7OyMdTRI
UyZ30zo3JzLsk1tElUF/c3q/pHSYJh+S1+lXkJTUa7/Qk+OlLwzfY8nkbMh2W5eKqXaSD+P+zHLZ
FOj/+ueXIfSxfsMelVbDk0QpYlErhV/puIdL1cEGfe48wlRstKdaCUL5yMC/Sbo0Lt2LvgijiY2l
Fe4BmVRV9nKnkHl40J3NIgVh2JmbXmzevkxRLhJX4m4rlzc0mavSMiH3RGnlRqMJOz5md4lGx7cg
qaRrCQ2hg4Abga2gl/21enoga8rZE3dqoAhAUzoTB5dXifa0z4QwsnD4ZF0FECobZQHSWhQ09ov8
C2RgsS+JBh9Y5pmlaNco25PkWQvx7nQ4b1IidGgRsxs4SyXWt+UZiWyJQNBKYHcGNEuuLyzKArdb
e95Yw8nEqmRBCcRLcIGK47HqlcxlZ/JTlqu/H3G7bOqwcexkC/pTbT5rVtAkjcMZaavpfJC1rBd6
arPrnbE2GAIrGaIjYYnGDUP/rJIoBL2ob4FtjvDxWb9qXHwpVi0NI3Lk3+8Q+T5cX3zi+N1mK7aA
KJ5+kg1863pj8Fl/mBKjBPa70eTBkXtrteqUh0t2sjHNeaN9cbnT9SInmICCi412AshzL3gKgRUz
cF+8IIfSTOhg1Yz1OVtrSKL7Zfw0IaUd86iKxd/QfA1JAxzAXaOh4SbUxxQksoQzovMcKR31EKhX
SQuPPFOznAGmjNwvwBZ119nJxJqDe1GoE7UmpVNkYp3u+IUAJ8f4QmTi8x3d4ZWhlzdkCHL3I/Ig
T3wZLl10t7YqM04NujKRwqLz7zzpQ3R4Cphgo5DeAYAIGAQ8muywkCp8bI5lAZA2pNjgFbvC1f80
sLSXJyyRi5qEOJczE7gea4Yw+c+l2akx6TqW1NBUw6ddkgQddutO2oAcKdoxQTcGSQKBegco7vpD
2IaQMQ8RxGxcMjXpYkfgq6ZG5VlP7r0A7P88Qhx25sylnIfuY+k/9WaYqjqMX53VJRojUV1SpoPb
JyHdS4Sc7bW6o6rst4h3rg/AamQ7TrHhRF9nWYJ8hJ+lloNzluiYSq0aWI2fuHy0sl93zHvEPz/8
/4SpbknLJOcXQfX16YJQF8aVGrQem2rcAoywe131Y1whKaoTxJoNVCQvbVX4oE4SZpAu7prz1pXU
WJqAVMKmj7pH9iEUU/MEbbhdbhmjnoIyYlbu9mdMoj3WpMxg4nHJ0hNpJICJVS8ZSBoBR1/E9XSt
GRes2mixyyaZC+jU+ukulLwwxOV+YpM7oHUn7p0ZaAARwFJAIGoKkvKGlID8WompTWWYPDvhO96p
Hd/amK5mEqQWs8oM1spW2/DggcaivkSOZD1yC1JHy6ZxOBhqtFfO8UKrbI3KxAoJJy4Qsdo9uCTR
38iwuTDgGCKPifjPSxrQWewrYpqVgKueJUptSSmfOYIcjPK5dK3o9OtEMWSGUCLDxRsAalnpiBkp
AHDENFKZSaumkR4EKnj2wa2CEVX4DvhaCVCb2WfqVmf3WWxjS7CnEmAxygke8Tl012WSCFYOGqw3
/kZQGM6eXwpY2Q8duzPEitu82MtZGbjjuI2YMVXjv6URhlkeK8Y4d80lT4XF+6RRZsyU+ev7Z5Zs
x0ykofu5QsRoE4Y5n5QTTbVXUAhi6mFWWie7U1esn3tHjAYhz26pM+PjyniL7Ey9OGilF0btvXGL
VHlp4uXjPUoetl/HsumiBltXJQsMPALnVrRiN+EFWJs7k6/kuGOFpIrEp8Y2cospMuS5lt2PLQuR
JCgKLnev4MZ5C03+82+vw1A9F4xXvyym0eHdZsWnO//m5gAur16yUjGUL2qSwjuoGWd3UlmHD/2L
06prDhpqqUIsZPjmB1Ajhtb7qNLxasfsOK7xUBEc3LmcaSFS1P8UiNLYQsdMxESpYFsioEiB2UOd
RaVuz27pMGBQ4sOJk8Sd9Xn1PbUeLDl+KQ4JB6Xfnhiz6qwb2TA4oOV5iuoCOXPjbSCt2it6DhHu
8r/t3hhtI8NJk72oE/ITAwkY4xi7310GPg5ag/Vkyr/dPk66S97e2UTnY/IGU0cD+Cek8bur0A9W
p5UQZmS4U206YPlxiTgZbz/XSWXN32Yxg5ZFo2YK3JA5UBm8QYSkuHas03g1rv9CJOEcyhVmcGL/
YRtMhNI+8JBttOko88ncCh2UTVZCQpa6socd9r90AEBF+nhKxNvS4x+ocVvIDQWUl3x0Tjchy3nd
QlwuiO/vroTTdp/NedgYFd9FTBSD3n5yjYZQCCfvIdyhBvuQibd/7GOihbU90pGuLP9lO1c0tBjx
PRIMmPfXkQfYabA7AuDjbOS7M+eEZeMJFwHMdL6GzExUO86Mk7Vk4hCQDyH8ZcwGZipobHgATAit
9G6E0zmMM//CZ6wVugdabL3qpVtTUMJiyetL6cB2/NmcUc39S5F2bTmggbQIhUW5N5jMHctP5maT
9H88YwV8S8KWaekd+B2w9GYKnXwuubNwgas3DVv6mbfGdZG9U9Y7fBsTW9SGIcDkHsp1jsZFHEzj
T7/oDF/BnG4dC+EWL1qeiIbinjCTnnb5dpnRgjR9GFm3XptV3fpJBiYM1y+wE1awuc5yz/fnIzsl
qjMJkXIM+4WZpzjXYicTNJEkcYYg5OBrwRsnR/povsl1svUZORRKhWSDjTdXborNKq0blzI47J+x
TC2Hx21hN5/qEJaZlICYtWuWgbLIRhxW9PR1IYj24i7U5r8TnbxtlJCfkrUtcnsBN3ilbAMQc7mS
jJF3dbsjhKdo2FX26b0wSgy8vASdXHUd2BJxK28ExWNYsuCgJVf+EmnIhbut3f5jkp/5V+/GI+bx
pJ8Tv+nwCfoiDw6lr66WpIvbf0J+MoyGt+C/gnsFqIs74/GzyOZK/ae80uBJumQ0kHHNSzsWjy14
b/8H7ci4wMC+7nDiUDMGB3CTerk+ikeMW3fbfN+jTkIfZRRrL4h+OqIWN7hCTic105Hlx6JAyHXK
5JxroJiValD7vzVJ/bOoJbORJvZf6aK0htvlG7vkK4ScqeyzavbaKFnaqPagNnPSIHk9nMlAva0S
aXgkbi5mPptx4Pi0pS1TuRZdC9ksZU8WWPRdvB1dy3jg4g5cT6fjEUDj9sVQldopsiWiTI9dcECN
VKr6SiSCilHJ0HRhXFr9gjCYGfmPp927SEvAlWfNGsXbcNACAMXIKCXnWBLXJq+gABWC5Q27n7ZL
zKC1tMRLXMKwBalu9sotz2O3IQyxwZ9qCm1VfLrPixIpJUrWfM4/RV2peg3EmcBN5y81MKuKvROc
4I5MOKFTYO6l2xlIMg+unp2dPoLjLVYIpCJK7uYEXosVf0kXiDQG71ofSMxLnNa7pkcjE9cFLI2B
q750LGRKpWgSk+4pQY/R/jUTVVodub2rqqnFt5kCvUkYuQPdHeP6EHmx+s5OOHNsFG98sNCCx1DL
1cyYv1KAz3tlMfwXQpZxNUIcPaVnib9bJMdm9w53Neh3/GCxQFt4M8tahnRa+HdJMPJiog3GAvOQ
UJIPVjSxrsV3eUs+8p5LuKgx7R6guzl5VmJTuYqPJuVqCLaaGV28qxj4Zf7UwfTaj5wXicuuh7SW
b87AxHghGwgO40Y2cS9LM1R3bB1bdqyKBywlejrIJZW0Z4i3AdNMwneYqly5qhVSM3sav3hRFPmm
kReZYcStZ8DeAJoKDM3luUuAxFjLtNwmk5zRLrPFK3ENM7MmvbDSRYbqFykNBIPj+D8BmvhTJ4sX
Sd3xLdDcXgZXC3JRWPslFefgUXyL+ImoLKbuzobOydQf00a+FT/4GfJDFqxzEw+TvEAJecV5uvAT
zaUxHWErlVCSi6zFHDJvkvSoZ/3SQLuSxZewUWBol8aw95+IwlqbHDFNkBMYrI4XZNGSEimbtlcB
V8vqldYV3YP9S3FLsCXl5j30rom8DgU62Fn7teNwdG0avgZ9TKpd1Q9xqDnMlCGLiQ5ztlCT3iEY
JTJQhWJUhjA4hjWfW3ckjWn7YbFYQdam6W1osyblHlAHCApi3SoxjU6VWCOKj7F+vEnkKbMdhkba
UZ6ZNsO/pLaBHJDqyjGSIcP/jNrV+Yf6v3Nwo5OYfnWsej6zxlhGfQnACzljQ10yDJ3bbsqWCrSp
WVVxJaaJ3/91FqUJs3IA/0PQ21PGo3f3z0zjYm9x3R67Eh7ZFEQT/W+gMvQhQ1Xo11zNCTiekL1e
1qNJwBkFe/jUtJr0vraozGFGmCcyrOfSi0Q/IuDFQQpUr7tznq1ozk8AsAOJRoSkiYWr4vocv1Ug
yn3SxRSxajagDXXQJAUJNt1/vqy+Q36VzDwTFghp/XyED2izTsn4XR+GsejwtNtzvY3lBAmy0xEl
tZI+gBdBYmAS+vPSA7u3JUjR0myH8tvFuUZx2d4PeuKrCFHgO2jveazsQV7Sv5fiallmQmPFAmmT
b5LE/QdE29IUeExBncjfAIQrN2pThmkn109AlNmov2nRRi0I8+oHN2uJf+Wcxmpvhuw1wfa/V3up
YFYe4fbR22ZJ0weMTJHFV7JUGA23XFpZizOqdN44SK9Ha1QN3LhwOK2ifugrIowBgCh5p2+mtUL9
rHP/r7Nz7IyUqGktwTp3ZLpvEkYXj9Oe4LwpkKkYRjYBoRxKd9IXZmQ6S6gEp0fB3kiVP1MCC2za
WWh5OYhksVWsQx/INGYUX022aW6e/v5Gbu9AMcwq66LyvOrXETs/rGiyQX/UJr6FcYAeAjxyQ1do
MMZbhvfWJ3/9D6jwLVbYdKwGWD+hYiURAUm1sKHy6iAsHH/GKGLyg4NG78mK05H/TrNMnCvp+yPn
868+ITJPA5qxGaPixkeJ35qmqua6CDO56EHL//U1vphLmM69GsKWnBc4c+LnOH0iehfVloN09WZR
mTvhrMLkqX4jZpG1umrnhGI+v4Dk2K3k09k1JwnnCxHtxD7nP/x9L2Xlr3rcnSDjinfqnessZAgK
GhBIa8T3b/kOaJncHdvu3h8hWf7ZSz5eXiC9y3dbyCV/qclIclCcywGJHZFZL9flA03jqWJnbnEB
g/bldXbwmA+K9AjKopjNaTJiq4Gqo5Xu2HWafx1Z9LLauOHMlOGY//Mt9rs40VkGSlwJPR87pbEL
gmv4QoL4PA7QpAcxkBPJW7j1UrIS7lQDoMbux8kY9EoP4qSSmBjny9sqzJEnFMEwDkaVT141mSKb
PuhC5mUHpqOtxmCWwVIZJPg+9NWdCjSkYBzpRJmWCnBjIDWMnFX5jrCq9reAK+Sfu/spA7UMvh2u
eES9pDhdgY5pyvuIRZwgarPG8ewRCjPIWbn2y8nrmtnmrgMlc5Gf/c9iMZ0vsyPnksAEGNEPi7B3
jlejjo6h7n9h1wqHaILMJj2VqwLH0SJXnefocktP2xghbRAIgF2OwIqHaTlOoJYtqG813cNfgxh5
0I21fhbW+qjjUI7F9ufvAIVoYi8afB7/IhmN1g24myCfIMZFYlgB8vujnTVSGrkdeVw7suv8rBWn
ndcf1jFDsenuTPmkuFR9eOC1OcDVs9YMnkn6PMuGfsLsnL378Yc5RxnX8eFSUyz2Vd7N/CQBN0xT
RnS9Z/3kv0Dy8cF2e4/xBBgDbs1WsDn0tbchV0+jBIaDxLaWYE4D7sk4eUAvO+64L3iQnakChCzb
gqsJDMXEAE/nC5ep9nlhN9t7o4ef0nbtw6W7pK5L2ab8jU53oMqegDwRFZHEiGJU8vYG2JWjZqXl
E96NFpZnngQjdkqF25GqEiI/86E2HxaiH55pIePuKi97KgovBMQaIUCkCXIzOW9h4GDfK/j+bs3O
DTborm7q+ZPxw48oIOiDZPwAylHP0oYuswKLY2bpJnZRyTpUwL27/C2GCBungfw1Cy7AW7iQFPDf
JogGuEQfhaaVyI9WlMSZkzYsm1dk8cZ09Oln1IE3iC+1ssfS5EejsMF8v/iJzYge3ZoX8j2r7Xas
FgtiOX5sJcEQd00+DemegJc2JEcM5IsSf6HHN5g5qJexNPDxC/lQatFdw+ZgH+adZhAyDOmN1Jw5
Xs5lXypXzdqJROCY6F/9gLP6f2j1NQ3r288cXBE9nCdgpbL+/4WNT8kMDtQOafPmktBkOtD1A06b
Og8rOF9Sf2ElzcaUPuKC58I+aVfLs8OR62cCF7pUmwatukswHlSY4C///ADmpUjvf5GAvow81dLj
5BVlsndFvgM8m3Cq9/6gevrdzdjsg8AI+YPdvU7pf6dXJL1mQPrQMWrC0CKB26IkPKPPp4IS8f2Y
6jhsAxw2M79OYJP3sIywB8lbZ23566dcn+j2/AFjYxs+HAKoTnS7jjmGaw/+OF6rv5OuDNZA+nAT
N68CC0VZCED0GtqeCyHe2NmALzje12Yhd6LnU7AkcQRw3ue8WrOcvJh1db0urpQXzPuZCD/LxC18
TQ1K/rfDTb+3oA99kjWQc8Xh1jX4Z9klrwhPINZpAdf49YxwOGyaGSZPAz/M+Ms/o/EjMiN/TacO
YiLZcP7ft7p5FGhY+e/zUSYTOsUkewZM9x0f1zp31rpBJ0JSLGbbHcRSYy/x4q5gPFmztfR0Sygo
Ps5vERxCxgrdM55n3X7uPUhzs2OOebNYVRr5TgQqjLMeggl5GZencVYN7X8OUdFvX9bwJBHTQtf9
kdklYF4p6ejcBds5oUWm/oKCEkIsq1E0xw71LR89gIo6enbyG6Vl+LTEoDykDyOh6VWmWvy9O/u6
bVi7teRSWGsvoXHt6yly8hbGsamhp/AXY1o78BTyRMGjo5BAZumdlRwYYzcj6Pemq75giCJ5yE2x
sm3gKRMk7bIkeOY+WgMMPG315plV0gNTUF4OamoZntjH3FhZ1+7YeiACyODgvtPoBQGBtlnFsOjD
vo3U4WfDt57XsPQZa3bQtmNlhY+zmaSH5L+25MjnHKFE8JlQvWAGdHIzEbqyo8IV0OKjYghRN5JV
wx5lrJjLGdqGtz/4cl1MfkjoxBmZdFCKE2/zGaYke5A7g0qHs4q9RG64841UBUmq+ODhtp2FpSuY
XVWXXZTvNmkYJwy1uVassaGtQUblnJOuDxDLUbDMgsNXNEs5MgR89e37jjamMPMwhOcXTI4GNmZc
qdVCXwGmdK+3Q8LJQ+eESpaxXpqlm8jYRS+aoWWU6AK6F+4Oui8lzaT9bk4Bk21VkXMIMSN5760z
KeA6tYGUve7M889KPNl4TdrH99eqFOVsLItfuqmLzDwvNqsBnVMpH57dbKkehKbSZJRhc9lbdp8l
djZ3RUUbIvCVrQQkvn8iYAx8w65QErg9xN9n6JcjiBQvV/1/TjZwEXkK2Dq5RCzGMNoz53eKZTGG
41nPTUIDsaGAMio/blHGaSc14ZpmE5BMByjl0GPjNYsIT35BE7bRQ40y2Iz1ing3923OzizkVPiX
OoP5ZmWnZJkSynYDxTiNwkjrEJIEI8aLsLL0ejKSXVENrdyereRcPDsNl+BsiA5KM6sKN8PkfZN8
EopVa8CNi6sFj6Gtg8yAKwnC6LAYutOTBB6LSMOMqNxQjO6hnpCXsA2gx5vBSIGeoXdYzhNmQfPK
SgayU7wwJ0O6NA7xAAdWzdgk1KZIVw0Vn+QddyzJKOAJOq+LiGmodQDoHdX9yIzE6LP4kRi4LUdS
l1JbcsK2eMbrc33hkQ3nbNx+npMDM/gPjTLkiBOmvTPqjqyf3LKm74kbqlb0953p/V3xamPHwAg1
b+8xZH7xPW6dmPe709Z7FOP+XA/qjUxxRCl4AfH2z2I/C1fmB14y3EcbrcMh3Ak6/m9Ql2D11Q7C
lqLZsbVai6FG5TDquvblO4LOuuvF/KalsUgsLDRMcCmxh3/i1+JbprSV+3UPCFJhVnmQ3jah0k4C
dCus4r95pZ2zSkb9pG4fNeQwyD7TG6+2X3gcS4JAV4ddWJFzEXMv0sK2L8F2wR4/1gmJDNT3Paq/
iuoDkSf8k2SecppRcNo4dO5tKRy9BuyNH4kyF3KGWqqT+1mzJeTsKvqOm5bKCLj5KEoSJc184pPf
GGPlxeQ7BKhQXuizfd6AAd01vwX0uq2pWPNaNDEX3GNr++BjUeds+yMwpBsygUNCNgfDt61V1hay
kySIj9zT6diBfF6SYSkDrIEPhFt6RHZukVUQTqfi3UbHuKkqSPUqG9ZZps4n/4NKDCLzpnfj7sKB
Ks66kuG4Lqzx4kngXQF7KuZ9cb1CtPqjW4WgPn6jKwdhme7PxDP1jajnxQQK42ghb/H7DVdbYMNu
+vGQRLPvEdxwrFsjla5LCwxgW16724EGxCScq5iGQ60e4tpLC4vhffsCsuNnrHfUAY0htrUTC+KL
xyJ0w1+VliADxv58rDfGGKEhdDObrB3LczL3wPHtYdp73fVqbr15EyLJOCkZFtZ7vLdARA3qR/Pz
bDcKculm482ntItpQN7Kh4GjRLzYtN4nqERIGjtPwm6nb6/6ndYzP2sKH5l6bHn6qysaQhL92JLE
A0KDMK4w+PB49OYsJR3irZKvJ0npV7422SI1vCmVHKW4YDz+r/2zl/NQnZ5tFqSnJTjwoddSNYEr
qcwqTpcgHnRPuNzgSGEfl3o+yUwDh6kDXSsongO/lg2xRXROpVctTFccQ3/VD+1PSho8gdQYRl96
IEmCfMWLHpQVVkeHbXUxRbraLf1Dcbpjk86QM1w/pvv8Q4T4KJkC07/enUW65vHn4tiFNuxCN4gf
GmczcKCLcz/8qu+5j/s/BGaZjiuXZCwjihc5HVmROcgFySoAc/LJQhD+mjADjIk+hK8YJSg+JrEk
lIMy24DJ2dEggZRJIe1UaZmQ71BWkuADoCXYL2bUoGLjx8wLQpEi4ebPO5gxveqf4mYIuw9xWVTF
z15OPbOSDF0jmtES5iadafw7tdnzMRGi1W6YMLnyNL3ZhtQVJtcLYM6XBRVmCB8tqfsaY5IiJvv/
JnlEtHXPVzqIEfkfGtBPgHMN33xEizxBRkjNoDIVQgxcPuGQzFCVE5ckXMRq7q7GSBqKr8eUbuQy
Oc8DN02TSv0WqjJI/OXf/z+osJAJDFx/ssZbvFpPFbs6mVXY7Tee/4xbKrXByrdaiywVDy3Z6Vnz
SLeoJlfJX64o3oNZKLxK7VIq4W644fj16jLs66FQjCGRsZpQMhsipkNcO5aElAKNIweGObU9Ma/l
uwHcchIhm925LKZKOvkbTYSgAdatyCxmaWY6yHPb/FygMPg/uWVVP5xj2RUpx8NEcL+3CutrDd7u
6hOF0Zwex6IujfeyElxiXfsZZEi9biPMQyGVLQwCI+c/bPUyKQyAd6gWp2vo1EFQFt4QMEYBGNHR
93dQMgQim20wg+nRUcpK7/hYXf9TekcH8hsRkQvzpl3QVpIMf1Y3ejDqNDrUwbZ5GQU5rcBvrAm3
mZZlWW9eEdtwsGWOZBOunAdW2Wk4u5jxTOFCX4Vhd7TPCGtvjAkY9owrGlBpMPpQmYlY0iJ3i1WF
Rq+noyvMAN9bRF/TmgpzBzDe3sH5bZaxHksSxWSbzVCFjo+ZJvmL9mYi9A6oOw37pJc/nu9Wa+Vk
IdyPyLPtvtfZl6gT6MVl+4A2GbggNnfmce+ihDjC3duSyjUYI9e62n/mqz/wXyFkSVTecAuJMa2M
iv06s8foqtibHUDmm8WR2HhwfArKUKVg6kMIJgo3sHM1eDJfffq3Vj5ou4g3/+bLfBasaJXsrQhj
tSjAvSlT+7gm+liXhf+EKKaWvjOE0IlbZ/7swAULw7Zu3c2qRsgvihO0gELxj63RtmgI16g0h2iX
qguBJaCUUz4jc66GhDQilN8sVI8MQx6FjDHuUU/9GWCoG/Ur+X9yl40jUYzv6Du36Qr6uNJACcst
D6AJro5u1aIYnbPl3b+ulYCawoxItBfOy3hhvgh0QKDlp1EpOFmdRLx/wIhcs6XAFzQBL7DWJ6SD
+F3J4QnrtKjxjeDgsZflDhsVQp8KWfPomzCvVQccNCnivHy5S87tG/eFMM6yGTsi8e+GWEaXgWX4
rZKONaOej8Va7MCMgj7gJVFAkP2xkjHnX7/EFjm4PisLcMSEFUf5v0u7Cn0eExsmrYvpHvW0iOaq
ZDT8zG3VH3+iYxr2a0Jo+4hs3iCYn/k8LWGJqaWMgHjZ8Y7aPP8BxJRSdh9avi8OlWbAWHyT8lwK
Rq+STMvFcIP/8c1Km6k/g9rmtNvFnvXo/Yr7hWyiegfNZcm/pQZiQ1nu4fNq9nddMwLrL0HN56n2
Mcn2uK3P9o0fbVZkpMOG97BO5TSuPiN1ktSuqS4pBg1pgAvqHM07TduIoS77R/TWuGNf7pEEkKuW
vZ0pHo4dXXT2IdDUqZXH6/aJCDY/G6ccWBmGPDgBPDPuFju4rulNPU4HDIldFt/t06reujMOA7ia
K3+Is8sfBBhkIAEXktHOySakFks4gJaM2mMImi2CRl2Qd/jExTW6XB25AdLqT/DdohdSDb7XPFWF
Qr4kAV7tmh/jBy/NLoEoBHp7GGFAVA/+5IrgcqIGXog0FleA2UbC5q6lC8lQbEqCc1LZ0qW4hoiR
KnGQZqw/+oqUAU6xD1YSoUvC8Vz1gIwsgZOtCeaBmxEJ+2byPEyxQfqP63Rcs+l2wMaiAabNZsGC
pxXr8tmhp8pRsFEZzEA6VQ/eyNSIIPyhOyuN/NgomzAdAylr3w0+PBFbzOr2heZhQ6w02Kn8yfMx
zK/IOjMVwQLz1eDz2sTVSncX9384VJ7PmTetJJLjpzCIYT7SUTOGHraYXPtgpEz9gFc9LA/dBsen
ZYfORhUh6f8FSMgoVQbOY1+/z2Y55yBsKKWM92SMoQ0qY+wpuMH1bo4pYjs5jhcyCelpVYzW38ky
aQaApZzRdncG4xL/tyCe20UhlgFY57KVPt9NY3j84A2r/T+gcfHZd/GKbAEiGm+F9xWytt7ZQykO
6JdxHo15iYRIMFg1ZIhAboLnIays6mp6fmfKlGk73zGCFMgizzBrqHukelMou3hDt4cWRNfeo4B+
JC5WwtU1qQKRVYdk7Fu8Oz24BJpo7+GOGjv5UK4CZQNODhXKXZ+giorYxomRDmPG6Hyy1X5uvnCa
HwpIV+iNN9fTYh12KsZ6NE7AzyOg7BfgeCyk4mVAw2/6vjD3Z6coHRZ34JqONgLE8udd4NFBNxTA
fbX3xgL0jP6/TGnexNaMFUI8GtWCDYltYS2vUeiHUob2HbAb+VUA2DNSeu/OgMvshZNShMapDi3F
pGjkVGmFrI5N69tAJdr0LEUtro401/iChHoartNk3vguq31zEdurGnjJcGyIr5dtuqWHpVwfLHIT
4VFmmqBp+mEHx2fWmp4+UlXQ+fydtbbQ/Hy1TXJtNwz25CssrKgm6EGyEAAruTfR4PM1JCJHGrQs
gQPbeQC4L6R6A7Fjz/dVVBmEDEjVkwHbRg+6gELL5RsdmiZ1fYcCkY+WmIJl8UI60OWxM2CNIPk5
1wFPa7wHg8Z3XaXHFAYR5vLD7MKFaEIy2XIUI6ZtXQ9qA6xSJIv0rmDFShnJRX3ttKcg4y0bnB6W
IMndzD5xShiiTTOwXlmFpORKflaDBeTk2I5UHyUtW2AJNnFZQQYtZ0Q6xUbI4ew0t4qgG3alFP3q
PMhLXS834uaOrk4rBz0w6qmeWnN7rvsqrGZtXbAdcHRKL3dV59sNhQo7iwc0Wu6uhSaCq6VDsUuf
zwd3S/b0xf7GwPP+gGsR0riQFmPVAe4FRhpkFIwqZuUnBTTdTwjZlQiI5gpezVsnYXxA5Zkd7Rzg
r52xFah6/tdQKmnvgmU0yE7TEA6Enul4fhkH/w47VLWFL4lZOnuHfGREAh8+XUxXdlspVJRYhZLj
VANzT1Qg1I/YK2piVXGUyYqsMN0o2dGFofwtmw+NmCbJQcfGbRad06vsyPQgazaIMkryMa+IvQ6G
boW7mjhkrMW9hJRZEZwnvsNbKuHm3XDEW6NSxnuAUWolq0ZJtNiwWysE0szuWiEoEYELJfn7si4Y
M+RjGcNNtYISGx1FcGi6u/e8r1dssXcZzB+piZuM5CmA08TCvhTLgekE+i8bFWpBgBT2KuOyNRnd
LziEGxnW57x6NQbkNuJOqrcgZA7UtyFrU0AQSjXxyVP/hNTThm69wVfjMkKwXuydxmX/10aSLTOa
ZhINrAutDaaFAvoWGUldtRl7iFBmhG6FPCR6l1vRlC0uZxHWALgRF7y7LnkwQtU1f9l89ygGsNsd
jhqwQlwidJto/9osInPo4mVGXxSYwbm+XqykS4OU1HJGkk/t7zv5geqd/1j4uUkRhEeEQo8nWfub
SNorKbJIOv5QFnAAZ8RVjzAArv88/FGBnax1MjJFURkWxH13PG2kDX073oON5BGVQJR8lMsP3EVC
G9SIPJdm8EgKsCrG4oOTAyqKzl2G/3eBrz8EbjI4goowNkV73tZhU3RYg23812XRaP9lHXSvBjFA
jppsnc5jytSbOWnnzhwNhmbEOFsZzllqoShaRwHIWckFQ+r54ZeoVAzIK2vDYanFbio9sib7G0Eg
N1DmCScWzrF4JJRISDkqgTzh8VvRnFw6RXuZPNcVIqkTYTIxSYQSq9BJpyx14mci3jnb8YwXB8zr
pbGlRq5OcvZzEAUeuzydCl4wiZzt+5F4XT6hJFHluPHZRHPV9kKjT+/5uxIClr3ngT71AKxvq9wH
N1vyIyReAlivoLMl9OvMDMtJj6nooWThjlrg5kwPCJF+Ig6ox9xMSGScmGgGkVAKPdVB2LXKEB4j
hdkMZp8wftP8YeG1u76pnRra5IWUGtlLainFVf1ts9+ztCwrFPQkymB1wWW9EQJcLTmZOUlNx7yE
JDXFnxlaKyHcJwfHWoN6fz/aVCRjpt7isHdxOs9UA0rR8BtvY1CVScTvECbXGU+En1fiG4AwvEbq
Yxiypz5iGdhCfdlnJ4J1zBv4A6dQ7EfHAx2dC0G7dSJN36uWOaLkA46xkoXuzFBV4u16fIwYc/KO
gIqChwC2mtCs/f40/qO5eTUH0VRc4SYeGixljDY12mowT6lvhBY7k2fVrSheW/rN0d3ZxEtK8vK1
YkWgEu+tMMDzji8X4adk6HVjdkWDsc9eof3bkbyERq1RmluT0AxI+9P5OdGQ5GPtdxZ6glx95o9n
L3I3oxfd/bZTwIFdDAphRECmR7sqCy+sEInCT+YvWmwJL+sBgL+mHdnaFuDfZ/oR05FieRmj3669
iPGgmDYjxGzLy7gJB18rMPy8bDizwKUj/ZaIOFrpDHEiQp9w3h9jVtzj2u1shLLdGyGZYlWcBDYR
s8JZ29GjyIfqXlia6Rth5nGGGqtUc75YL3kaJTnq0W2BU+bsh4YrNyIgKBpcpaBZHLFKvyW536Pv
VRFvUZOJOOtgbjhy4ohzxc2ZLTwfJj/wKWxN+tivvNzG+XInSlNhctew79zKM3F0BYBWoss+UMWa
+wbxy+EplJnqqEpHy0WgNtdw4FrsetSJMifU5VqpwFYihntnJaA58v5IpylxJY4nVVvQfuMRYQJz
29uT2NteQpukbNZLPHbLa9ErPzzO9kbO0BeUyPNJSEIKBN+zr593w8YJxn4zHMaV5aT9ogCqlbGn
4AGkhjkCDZDDtDlr4LXnnXvM0u2I6vFltm1fb/2+bIEz/WwPDgK1DXRcIqIdz2wg9UORtbsOfqvw
cPVAODaveeEDSeEzKJrNjbpZtM6VdHEeOUey9+RurWBYwT9RobTTMSvkQqo9HSe6Mxf5hTT+JtlS
VVXj2xw0Xaoi4Z8kuJAxzx5PWpHgHyG7bTBvkVlE4+mocmn8SdPjWNpg1xtzM3RrJMUDSftbWlDm
eMcBcEDVqsE7jp39gSt7B3C6OA2des4CS6rgWz9rdW/EsdMkYlyz6824Eaa6WlcTu1MlJKrj2zq4
WVZ6auTpJv4xCVM2xLmxHrlQkElm1u8k+bVfVdIcLRp7w7nyO4g4l5707WMUbUn/gpfvZY/bx6f/
w6XWD7tG7Opy2qyU7aIMOp/3zcHqiYTDSTG9cP44k9VVPBZ+QTypa7/IMlW9KoQsBf2mSFMK3wbo
c++GYB2iZgDNB2e/lumbG9AZZFh+s+9FzMTRybGl52fTQ8CTGubM/OhGhLyrjdv1SxbH4N0UW/Is
b0fuPAWL/naPShegG4qQKtQFd0FnsOvlM2yuYXiTAmJep2l0pZupuZLldObZH1lr33PozFMEDpt+
/bdhLS8lPb5DfX40fYjMePdfk0eG5enPM81/uiDlSBV+yTcJogciVKMutC/unjy8+lc2yCwos9E3
bsnjB/ViOVrC0LnJUcO2UqqcaM3NawfjO4HgHPuIBkMYRHcVhPZUEmA7Y5DBoZ0H32892RPBPXgE
cHmc91/lXeBi9QZB2EkjMJTlws7HE7111PGDt0Z1u/tr3bqDEJWNus6HyW4Zu/3dROqal58r9Q0S
SkbLRGXI1YKY9BdHN0j86YjU5hRxK4pBnbWUcFMksi03v+oxx5jCX46qVM0zQIzz/mjFa1NnisPJ
uqz5mBv07Mf+EelxgoyywvE3SeayF2R/Aoo6sKu47TNrM9JgYn9Xj2EBP1LNTFKrOiOfRYrVktI5
B6iMTSzAJmSPwIO5H0W53h+1U77bH8pBnbPe8bzCwoj+fdLs8pOYDJprjnTFsfxr2SBJmO++EBss
U6lc7uxqFfuCWmmDa9VxAa3S+e246YWwOA9J5DWGck5a9ARpW2b69BXcEknaiL6lw0SbkCScL4Ze
bVCZAh+5c10vO/wVIniIQeOHEMatoP6WVOJ5QWkzh+msvsT1pAWDnHutayz27xT2UcgJAlN7LVZs
s8KXz9U5FXoKWyKWAkiIpcXqueyBhs++1dDrQO9t+EpHfgZuSt0W8U5t4CDeGfKUp7nXfregZ7y/
JUkZ6ZMfiQDpoTuhqBkidoVXUvzovM0bBBySbjXzZVHElsNOpYz321DR1+mR29cT6A5XEeNa1V8v
ZowE3Mzh/up5a6XKyohabIaukPExhotBlnZ4e28LZhlWgUQJxdiKDcj2Gmsxke5/rmn/wN/fzS6Z
Jz1ZgVPhFjTc9CcPa0FNlDd1qyqHHPuj0Dc324JfpmUSWwYIJO+T3okXsvVX+Fc/vvITE/4ILhpU
QQS1ST8NrtPru92Bm90R+yFM/5ajP+Ry+WMpXNA1QzX6sqkjrgJFmmU3MpMkG2TPQcVrRZMqc4cL
WDlyvXrG/ygujn6aS33h0M2Kt518A5uqePDsHn7vn/0p9leKAXxfhJLWbUX/y4zeRtKRkibhpiyn
j/ip3DnFpzOCHe5FE9sm3od9LTO7qSJV6dH/Fr0isDCl64b0Ttctd6P6n/aqXs1oHOYgGwZJmNEp
Nzm+5XtB+HS87PAQ6REl7gWK+JQFpmlhJXXDb2cIJe48IPMW/KqE5Ud2mQw6ESmkQsqPQ0GX9R4D
p5YquTD7YEgLBf3zjDNF1dR99Di0zOfISmNN0MWKHrhgrEoUHo6ED7/DGLnC3wEUDn1yvLm5uPYs
gkiHCFoqRsSFixUA78dsyqc37z7Tlpq8fQ0MWYgHmLTq9aB7knin0NdXA/JrOlzH1NMQmes70m3e
vEplIfw4yB8DFdJXpbzU8pLZG2RVnD8pfiGPbjlGE2BED6DKihq+adJ3Yx5ZIpEEDRnqR/BrXtiQ
bTaufhbv5tXP0cWuKI0rlXhs6WnD3yZl6QpGJhZImANTsmdvmHkGKe3ei7muJosMbbUsfSWTdLDu
QhzOdFMVaQsvTBao8dFa2GLH4dIlcJqHu0NwRhFmYj4XIUz4mmW4XS6ZIv+akfKU65rhL7bICCQn
8n0FCH6ggPiZ2JlS1HVp3VGmZwOvzI+43uwGno+xV+x0xRuoTN4QXzZa+tXGO3ssGtg/a6JLQ7NB
/Giq72PV6SZuBvJhkTIaOtRn0X0nIOwHCOwXkrVdeB8PKz3fFbmsluPk4AFzault/PlVQCPTEaG/
9D5QPR/hWAVk7+aaUXkRQcTeNusNNBtonsYDYZnOxO873qS3XlsU0dLi54KtDWzDPr05tkHKHrWC
wSz6AGB+6gSWfySUxJa9ETXcK7bwsNk4fdSeCAPQqlb54PtNsMfK6+0tGOWqEw27q5tWE4JB0HiV
0odVo4fxX8r0Z/TLAnFHPRuBCp1P3iyZaB78lsMXYSk8liKjYvL6z3BmANxYu62aUU1QpaVg1ALu
BI0RX74AoBBBWHq0nGcc1nxwU+LMbI9H8bw07qy/QrND4kESKEUPxHn7hziYkUMYJzad5KUrd6Rl
FYbZoFLP+S9J/bDrM3EWMT3xmzQZ/dt4d/EzL+V/6/EodsZti5w46f3hEageuFeiaElvRKoaQMpB
WKZFGsysy7QIM34Jv2hjFXqta8SFrXR/02uJ2Xdz2o7piyRqorHUDTcK7mjiaSxwA0Ne/dPsfV9u
p/HIi8rOCcQO1eAndX6/ulZ7Q1JfTyNczv0QfNjfEGPafnIRYhGWC9LbAOr84SXGvgUT7D34c+N/
uSwvrZi7gzfazB7h8OaNtFcAHuayeEhkiCYi3azd33tgv+NSwSi5m0vKZEK8+0Tlnp5x7Om8NL44
3p7WYmTXeRxv0N/c+ALLHEHRd+/nJxIydz6eZQKKnvJa6+XoZd2sTJ2WCrMbFqaF/D6GGwdu4Ict
f7MTSJBd19iws6gryvwlAj12+sHGk6EtIE6EXPSCgo3lOpcxdyhpMXgyTdPqSnUnPTCnSaqO+LRV
Sbth/8hxWOhnv8GtYCWvY64y6IWVxwkWv7wZUYdPyRzN9o6tmG0loSTg74+OcXnXGMKWsx3DOl/g
pWqYjBRb/c13/hIIpSBg7WVeQCXWQCDJbYuirrxXpjKIHGqC5X+X+arymI/SYNRohegNpEhRInP3
oXm4IAdFAERHXEt6R3NlD0COpKFQMWL+R9kuK5TllQ/Q3C0Zt4na8FCCWmCNzj7ww6R8rHEPzJqV
Z/qBV/FsTLjldWEVyrTk3UMiepdPd5YpcnDz2SnbOsVp19uY6eh0gn8xr71MzRdO1dtXO1iWP2VP
uWulRG0XSRqgoHW4T9zb5pkhpNIYustAC/G7lh+UwdLWDYP+8ffjclb0MGh/Htz8f+hBmdrIzK5J
S1MMyErngBIIoMWMkBHJgigcVMbA7R/tM6I+Fvl923lRc9H+8ZKi+TttLxbOs/pxXGTqdEqxN24R
qQfnrWb4R/Nu29GqX5ca4yzeEzKLb07dA+SJWKjNDcD55vGTKzF/5zIrgAtDyZ8xWv/yRWLUgAHV
6x/vWs6PX5rpgOPao3h4UlLNcJnSztglu4ucp02aWwBkeW4siwBXBZYF+u62e3s28uZffJW0QVv7
vlj35ky/kyKgzIrT5kSFr1r51aaOFg1ryTGDlYLjiLuoEXYstVS+nA7VKIumd/ShG2cBNLmQMvjA
Lpnes8rsOv8JpoCYqycfohrCNXz1SYRD5ar5cqvkETzBlouw+2iSnCPvJdx+fbjuJgRWx2w1BPPr
XijvIMJNw8y+dUg5UkgvRc+tgow5rTBZJ5Pl3M13qcB+z78PtMCJCL+OZLTLBOGwoE/d88OnOOcn
IqN7s8UnvEuPE1Y+CSpdi+iSEBmAQrfAQF0MJTQmXNVBPDk9l+nSJNheMvIOq/uSXq9zffZtTLPs
nwhdQgqVBlKf1Q5unMasVyx6J36A+pXMiwYSfWmhPD/WryThpEAb8bxd0CSfDKLrocRv8irxIiXW
yUyy1ttawrnrjiYlvZV6QUUwovUcBIwSLi9Qni7rLDGfCiqI0jMOnXsc7+IkXVgndpsuzu5qG2nu
tX/CheYghlFnwbDSjb7vBgK9eTST/p/5oh7rdqVsXRecio7WZ3mYhStxj+R/MRV8uuPTOUNY1Axx
aPDRkHJ9+KHrOpeqYd/F3UwycPJKs/cGAjp8RHJvm8Tq2upme2XMcSCIUCx8SE5L+Fsdsxa0+ZCX
CNMbOg2tsHAY/tHGqQ/r9Wiby4KYOLGgqaoSDAuEokUhvlxL42oj8zK5XzXjvpGOx8Jf68g2yjjU
D/gnKO+MqdzZtoFW0d+PePmhBDgTIlHGBamEO/IxssmWa+D2TxKwCNn51qg2fUmUnfL7X31O2j2e
uXdQmB4ZmB7sNupzjrqNICkm6jF1dozg85yGfV1xVcg9m/5oI/KiZo9wEbIniIk7cv+QOPieknBZ
Nc5yPGJ6i/8QEmtXLdktFBYlFStkUcxgdmQp4lcvjxV/JQSjdo1FzTcKZ7G43sNOlaXZ0LqQqrdB
ojnL6mPTZcMHEosdVG8u01TiqS6ycjEVTXkEC3qO8gHnR6Zimb5p/Nf0OTphPj3Xsksj4YuZZlZO
XceclGkdFr2JiXU0UO7lZD/x+rLz8Pms/JfEy6ULRpmkOTnK3CvoFdHxSXA269Spd8MA/4vFni43
eMwD0VDLtxX2fA5zWiAqNmuyXizyXtMgHbwdUFzX9rmZH/eJwENFwMKDcwUsU1WTl5huCk3K859z
bERcr4U/K6d/XbwHWMBgP9K5dqOAMH5YIJlHb9VHL1h911CuKUdk2OMlKU+TVPl0pZrKZ2aIxu/c
yb7k6bxtq0xxX3IvH2t5yk03pj6iK5l/ICTNA71BVc2skk6bXgBy6vZ8OrVzr7oWpcrg8JoSSzd0
6RTkEnhIvSrknBYXkaudEXYcP57ctxBdnP2UnlBSYICZRKSSEOrErgAFYCYJJPHDCIsqX2ti8Pxm
z+vsiWqg/iHTfEcWobDpOvSkYCcN2KoqvOkQ/nFh2JLXq6fidmo6Ckr00lZdFuwh/zy1vEmN1cKW
tDuGeGnZ92kNg8yNeH3T8lweX5hq4750ut0abL+C6X2ePA+KUaWj4Rv6FlmjmlnIDd9EbEpw9mde
4mYe/R9Z9j9humdO+AiGqvC2E1ZKzPe9ENhs/0QUh6tFCgiOxP0XE25LQ2BpC8NPgPxqGOk6ZG6L
3yVn3WF+DToc6CdqgvbcDcmwFpL7dzS7p7Nms+eitxGoWPbn9fJwGH5n2Besmls+yvAHN9QxiJhB
JLEAKRjGUB20F4HATO5U+7Y5H1BdbhQheQ7rUrBwZ1/rHS69S9sarIQbK/bvaiqrUj9yx0hdt1JK
gJp3x8Dp4uRWLHq5G/mc4NXJsRHpKK0o55xSSxnKyYG6so/brZI+zEYaj1bgKUxsbw+zr5FabnlM
Sp4aO1MgrhgKjUCH4EgKYYImSEQH6s2iQ7B5mizS2tzxN6Le7mMaOwf8CH2IzSql3R1NA+LCpSdO
d27hiUf5fp33nX3ymBnyPrKyDO8k68YUV9dLTw7wZ0me0KSKdKvDii2R6OVWQSzLcFhkhtVEVIjo
9lDWXuqYzpa6pOWSfgbnz4K2qvohavVfwCQzIDpPJNQdBCsTzafXPQ/xC5+GLBOPBvS0qZiCS2pW
+cQ9z9yDH0inUu1+DucMya1px7zeWNja2PL7qB040l8QBSpPzQe34vp+ZulscvNMPT9sHVGM9d7G
ran+LQvrNXuHylejvtQiv4Qgi2bz9/v8JcPiO35CGWb+sB8hyMSnGwZfynmZ9aINq1MdXNR2Nccp
6nNZSNYqgqe51RbxgPQVWucTfoU4jh6Nx7ogJ1NSto8ED8kfmZmQ77TNB58XLvJbIDB0OSHW6Rhj
wkM/xzErDvLE+x/iYE7aJGEjpUfA9xQWvK2EMkN3hIeEOnLuSOtNUrnb5/AKa/MV+TCUKpa7pibK
XKQWqxF1aNI3BH5Bfx5GI6UOXzkF6eitDkOxg3leE8oFi2F9s6MqEMe/0PwLpPYRKAtK3Gy/9eI2
1YAh4csAiaKgvk0h9XmPvc/VayUgDQXalyUnLEWtX07h5M8MTvnO0FkKXvHFrxU0m4BcDE4MAc65
Lv0ctO+gCK5N37eu8IHNzj9MJx3YnQ2MK3YsJz3Pmv3HLegklPE4Pg50ynrIA2oUtz16vUHSKAdW
Mz46Z2j0h1KxqKcQbmccGfa+8LDoBFjD6hYJKv86aqO3IAGyY4CmrBg22IMQBhW3u3Hi2vfcGb3m
JYEiJggYC5OO2t6DNeJkH3jk9sP59qvkEVc2L+iiFcdpIn1v2p/eCcPJHzFMGYtQ0l5mXh+uVQVo
XfhsiYmPUxBTf3T1iPxyAPItjrSVBt1g9SaiV7i8fLaYLhlZeMppGSrpijGDPUOGiJPdqWDWmiEf
yyMLw8aA6gtMKg6FsEmsVgaFU0hCHOVtw4T6P0H6FXAUaU/DGV5eYIB88ZwqpX3oc/fTRf2v0LUY
l52e01K5nlsCeKJHUc4Zsqf8vELyE4QJA5Wj9nzL4CRClep+/pKXRBr/HWBXgLr7F0aQNTN2PDGo
JcSvMzNpW9PAl5zKHWXpKjAwAl8CySVOfs2Ef1aGeLPzrytYiuzOW89N6XVKZrkgOt2+wqs0AVn1
jbSznICJAJL5YQrvQavSECiWsKJktdCRYzp9edUAckDuHq9lz+cOjMCLR469htYpFiAzLpXORNhD
soA2POV/JI8y6n3CoxBmTlnkaAVxVHRywRx9lg9scLRBfmWXYvQ+14Rf86hqWH1nXt2P3/6IV/8R
vOpXChFxqMa8x45z4FcU5gPytbjQBuaw+Rf3w4BVyk7w1DaIYSGVZxRrJeNI8W+jgsdpsUKrGWQA
vnze7y5xFG9Omxz5jjunI0ltlmN6jkleIFa1vTPCJsQ4IzF0xG37Nc6q2JBv2Za+OdwWDqSaeBdI
Tsut26GYQVehRh1wGkFaGZZDAVxZ0JNmRTTNz+OkV70SF/U5f24orhxglnLB52ns91m/zBMc8Ym+
pn9WVVdoyactIj8VSZTcBDUZkGRY6i/0WFjxNiIacGNmlq3kYWLV/i4XBzkcB204E5Z2VBIFWivr
rpYSiV1m0yiO+bfR0cQvUBx+xVSjI1fgs0+zAx7V1XimpRcOtaQZ16L5t9raruL4+7TGPtxhZgAj
1ITc+ojBiKJb7OBd4KTo31Yc3+qYryvAJFg3X2bgL5dYyirZCJbVzDhypqnRPvavsyF737vDJyk0
tra1+Bk9d1jclW5nZFXZ1kH+eaS4z0xLh4WR+6Rv9X4kigYX95+23uaOErax6rVdaTWteIXeGRvH
EEUmiJfHYsACH3DGal8g8d6a7Cf00yyVqi0zvhY9awD2QwxU8oxqt+ykMy5IUwKZwK6/11w339D0
Pw/817eTmkGIioc6TswZu0iPT2egAPa2W8YJxQAuwfP+E8TxFzYuk7Z8Ye779FxocpvkcndLfPhx
OlBUzINbxwS+uEaBXu5JonZ6nPheQzjv7mevCK0pgpJIJFUWE+eSKY/712NEY6cmw5JhZaE7+vK1
4RwQxtb/NeqXCBDtmbp0f7FNYB9P5MpNdPKG1kIWTCSbKA8wsJnlj2VRmGEORTaLY5Xrx+r8UAYw
aMnl9IKXg1Q1LbCnkgChnP7ycXnpc7dDFaUwxABZ6WxTYd6oWr3BjVqgAZMYP4eeCKhaE/0wIKzJ
CLRYOZxB6vP+626avqJfFORs8O7mqfYkvhTucXaCP6OTVg1J9SNVN7A4xIf25XPd+MwXn1o9ebqr
6j1YbvWtHaB0JmlfaT2fLqfBI+HCgHujWNFjWsh0j7igkgIz/76hESPtqAd5tb8d6o1mWdB8jOgs
1YDtzBDj1xmGJ+Juqrmt2NeRfalgNVWSKXtOVyQcz/u8LjQkLZoGUNSX3N/Gdo6VzFb2ME76n2Lu
qFpeccOwcl3jYjktvlZ1s4xv/hv/y5au/qEFBBxYaeWv7o4Tb+rtPslh27EN0lcv/029NORn+Cm0
oHVSzj9MbxCV2mRIx33ChXxv9Jw0I07AVd7aMdRbos9rmQVO0oDPdsthIfZI6UI4GzCx/JoujAGa
1bIcb0T9ZLr6K0oHe4NuV15I0W7dh3pEk0Sah38uvIiI6q3mcHyiQOT0Ln6ydltEHxqxfimOqPgH
KCWSZCubNKxx0T4IaWcOFg6e4ePSsXnmHvUx9qnJM3E8aah0bxnnlm/OrTZdluXze/MjMB0PfLa7
kvcq+bJcR0VHloWO0sqLSaSDPqcR4t9J+ZlckI2sQ7iv7qB5kAIwr0Rh3RuNO+LsgEwSqhQY7Mmk
b/QNjet7QJ4Elm3Vmzlr/Jw/nntZkGZGNNZ/a6lzFVQsDpmqvCTcfu7v0wG5tLsxVGADaum8aHg/
b+Ok37H5/0NggS7DihPTd0QkSNjD1TDF8/CAAZftLiiENbbWeHdrLWwonGsPk1gsSf/4PEK1psg8
d6fB4XbhAVr+R1ncgYn9DpPbpogRf9XSx7Lp0XQH2StYAzMqdXf6i0yxe7kAksYBtYAB1ArGJ9I2
vrXYymprjHIE7roms1SQLA99AXgSj5VATi2eizaVQYWKWdzRhuAXirGrrQdQ+ATvMH6QzXQ2ubu3
RT1LWafJP2Qd3NLGuqc21jL/60PQzOVhn/PjCq3wlRcIlhvHyv2xLcfiUFOewcyp7kI2tIryJb0G
epjB61jgjSVsGNi1clXiiV1XYnZU1s0A/TMAzlhI0UTOWWNx2yavY8qX2R8r89278WHe4yhwsmxE
gdp51Rs+MH0AWb04TIBnMOUVQqyRXUYKVNmVofW+SgESK2u6v5OkNmxTOaFosubx+AfUy8/9Y14+
vD3PH9MZNRUGVW/4tZvekTtFknLrCsZoudQBDy6pyvaApPNfQ5+4fBnqT2sRc4zbLf+7e0KR6UlO
dX8QEejIEBPDGCFvZwkXhsbMYO22vOGqEOIRidII8hvli06tNAFak25jLNZ+dpfobHsxDiMD3o2C
Rd7Rykr3+cwf+00Z+b5BJIBZIcsFqWsYKoPChTrfhiQWAdoJyKU1EbOsEm4wJxstcWFAz2PBCP/J
j5PcUU927grZhTJ9iRroywWisrIpk4Z7FetDlkN6KsKdVXCB+uVZBpxbRzMMCYuAQ0dSgos+pi1/
OavTStYOY61HXvtjlfMb2fv3HfP+w4PkJeDcuuVX7ec0oJzo5y0+JxXcBRCetfOT2Lo9yIyaZmM3
A5XLptYtz3C5Olr7U/0pu8J8Sv+1ailQPrvxLtDLZoU+Hj4iVXpm411X8Hhg3r0+hRVEye8o12Bk
llMNokEaBVM5tpznHkvd6n8nWFVzzVCckfoODUutOAyMUn0d/R6Wz3hqxFZOeiX24N/gEdP7GZDk
VQllaPE/Nb+8JYEF+sPkEmeInsGAri7lNmaxgl/sUXSQC1NUGWnGXjHQSwQBzyBfQL1u0N4yh0oM
5tTt1tWsVkdKjom4As0G3qfwFZSgv+ySuVhJdzQ38CXym5wJz60VTz4ophOw4Ivq4qyRwhs6r0tX
peCLS0G23NmJScznhl6DUCjnufhTM3waVHTZQTtw0txBj4KOIuDAp46ZZi5NtmJLBP01yTV9HTwe
ifPOSKDfvaGIzJQ1RW3ilsadQu+39dvEknVx2ZvpIyBGR2cUdJc7UDjnm5UU+wR6iWRonaXYFhwk
uiQu16GIz266OBsAzIDlqfruFHHZnfk8OBOB0KgmgqCnyTeGH6qeXD45wv5srigdPsY5UlOsnlXp
hBMSZx8wZq1jhyfRm1ZJKvt/UKrzg5uXIK5I5XoEUGrIgVxiOlVzeVYnSBJAXz6D372+7oQY8en0
T+SNRuD+d6RAWIP1dj2OgsGWNsrHOcrAqDXXKee80mC4hLVucYNUh2Pg3GGkxUurHoxMYACH3ysd
D6yn05PnrYYK2/d6UNjCX26JvCeQsRiL0qHcjnIoJ//FUhCoVIWFx2Et7RIi0cmSroA6xh21WOpN
7+0Zrm4OX1lKoTxBjhr81ajuSwqClbKT8wyHl/QhpzV+3bVLEfq0tcF4xVWr9xkGS/j0fCs7PwS7
IpU0P5SyHc2JkhwmWbQxrCBgK7vZYBK90JNeb0fn6pZVbWaz6lc5213MZgb1AJQWS3xzSWt1vXOb
33jcZ+sL+9SX52YBOPr7zje3lbUdkBwSfovcLRZq56r7JY5tYiv+y9AGXHV4rX6gjD31maVLYQCK
Wl/bAwugYMSwhhEhhe/6v3VMX6fJ2KwveDjNSWh3QUwAPXpAK6ouUYJDsBbTslPWhgWF60z8VsPC
Q1ULtPSYyZDyyKw3pYSGOmWnMYgOaCAqY1Wovw+ssV+eNdQ9OILuL+BiSUidCrijkf6LdXiDLur4
8/8HP/RTUNwsq1S+Q7cdhWHcIXOFNYzOw/W3yz2WL5BsyQgG/UW8BVBSdsto4GhszzaT3LHOcENf
umyB577OnTIEWnAxvlDebrY3hQ3tl0K2koh8OOc+SKjBfB8P0hze+d5y2Isfs2CVL1GeHlI7bWzD
q+pGi8D9EKZNN6+iCjfWc+C497xUXwzmzqAZbUSXf4FMkBrLx6xkxbcSK8NHVlqUzbrs6JPIRcu/
KpbE58GnX+JptoEoQ4v4UdBr7D6cuIDGgVP7uYc8i1UM7oZLFpFaILUbHZo4WTqxBVTTXSqdiepm
2W5uN8A3QkVMf6GBNPb2kwUuY6S+bVJwNoxLgcSaimkggqeoKjrqFhv66sEFTY0HgyE4VXZ4UAJn
qmAaSx4Bzitv/RezGqRUl21Ih+5iI4jfu4+nXPbmRBiWhD6ZAC8Vll0szMHw4a8CAE+91u9ftqyn
4pFVR+KZILyaH2hTDm00FKe1+hCW5sstWjazIb7p3NtIHw/Z/vRYuHa9nb8PBQO2Ikg9i7zGBsVw
SVGYwNJRapE80qhH/FfWnlvFWwK7hisCy33+/d/7MGuBPpsDC0PlsmkzBxI0Fbr8Y/FriH1dC4pg
Yg5hBCZJsxTeujXLXqv5kElIuwoY+K3JHtCkEFp5vvUGY2cPKVOaGzJfl1wQAr6/q/epSs+XZV7l
HjLuEi4d244UeUuXpEZvEsHS42yMBKnFzVTNL2Op4pK6sDDKn3RIwJTWF/JErlJ9/9XNbTLlpC+u
B6cdH2jaH++BadUjjCLrNFSZ3rpnAyU7E/rjqr2eoTNimKr2hxJSpD5i4f2cjuVH5R3tn+YcflPH
z88Q22rPz6DsjpaQNz9PkSNLHhp0MMWsWqQA/7YGFd/N3JratHfapAE2AVb9eZfwtEt1gbsMFZaG
F6GMs6y+fG9p9efq3HfTH19VWtudkvvoME7/0mTD71ZgE2VSgW3OuEs2GmNwSd7m60hLj7f4CcAp
x/YC+WWYjBAMilrDs8tcf+NiXPGiZB344shuVzbOoBcLiAFCqbLOljOTMMr0/v/wF+iiTQhyMi75
HAHdrLVlEjc4+cTp2P4QaZz0bymSas5Jl+glBGDV6Y65N+jf1LL/IWStyKto09GuRNV/ogVpsyty
EfxcY/tjuaihPbWzGnU9Nu26WNOd4X+ECXLxBps2HVft/HdKBDGEx/tVHqFIkb6yseuaRaXKWfgK
ntLHvTqog2sSGgPk3sPl90kLu9t8PNzLKwQrTEjFxVTN//Lufbj9kc+mNGBGYGtEjxBpkR0vNFQE
F45qGf3Whox9EmRxUZsjy7FEw+E6tv7X/k0jBp0DsJM5pk7JP01ZUlt7muTG95xzEH1BcZ4Nyycl
Nqg94o5KyKwa5+Esndt8hEeCoBDHNNno9iBqbnYfWk1KVXdfr3I9jgk0AD4tEv01xFMPQrix6MyX
9g8OMBJB6sw1LdTDYdkZ0+ZMnQOagn7eeogCEox0VsaE+8nbylepwPOT+okCkpoSA9ZlMBonKOFn
qrWAvBIZc3KjZJLTD7S+ZHcleotJ+YXYhG2xzQ7OQMAiDLFU6R0z7GVMEO3zEf4+VcZkywQQRdqU
VKyovwwXynh/qYwGgcjp1cqkO+IiR1mCm1nokMdE0YKxXroFsC+KFH3r5ABtqvvBBZEiVyiyTNyT
lNqYhRTkUvNUQikcVwZ4xGi4AlmthedSeVp07Ss+/wTtNvGP/SFrRGl0ETqV3kJLvDLl3s6+9PQH
pEvFE5z7fu74pXxkfKtVeobi11A/lPYRgETfXUxoPhBMiLzhOwPYbEEXQSCrN3Cmff3oXN+57+aV
kq2AmZuJevxjRxSeIshaOGNCZDHAWWr1sZoubQBk5stCmBM7T6MMozT9RT4l0D6B4vwFRfpuvcD9
2erNQTnSdFgRIhz6MPyTraRNuWNbsAmdI3Zor+9lkdOvbGTzrXxPtRzAmsjzCZ2Pz1qf/rIRnyhV
2YQ4KpwcWTNSozo9SyK7Fs1EFUBwAqDoXG5xHNKWCMRrnGR+sWz5hXvkidnRhT30FiNk8uN8ZzVR
dDuC3F0FQNVWiAFpY9vVzMtCullQ2o71jNPx7lWBUBwT6bI0ydniRxiny9Sp3j6Wu8wJZKWVzOSa
VAXD/1krBA1BXTDrihskgH2+oYe6Cxn3G+dtBcF5wNMFgN8lh4avf6C1jWLHfjGOgUXv4qiMtJTH
tNR4V9NTHMSZS7v10HUhVsYThT0BbMHLJ2ntCoq++2TbKOxSdRQbUZUfET4bNeYqOAHS5dSKTKG5
SFDNczJafz64S3aF/t4CZh6oFp6HisvKDi2qNhxs8sM9vKJJYICayyrDzZEL+7/2aj6G43od05wM
2Bru+5FoOqkxdPJm8zh7Asy5InlJ0d5VqglBrJNppGbg/jmkXiHeXgfOEalr8AuRqXriW8jNfbq6
QQUILlaS7SXLnGth305oHtI2v4LxeYFMClK8w5U8ZDaCuaX57juJw0SJdTrs1mpUffl2dwFNpMdq
kQPlaQFmnf9D0JLlqHiDriQKpHHJeIcDrBEuZ7qYBYT7LqUgPnyn1OvSgmeTuUwXj/qc1oWG0Ys4
w6/gGImC3isuUl7qIEoLLLAlvjee+Qif7ZkR5iQexzEVlt4ABccJltOvrto//LkHZ7U+2LuO5ECI
PcY9YF62VFYu2AGbpll2toxXLoH0DmjWJAB7Imd0jqbFx+iAOTs1S/IjcFyU8X2NunSbPAJatoct
gY30gJMKfByMwaEiXq4RZwe7ZGCwq4R8m9/g/ImUZ31CqeAq1qI3Eb7Xm39a0VKTWvVmvVmBz+Qw
gdiUqeBhf6/AbkPvp2w56Rv2PpWCfFzHO34yhPRTlGKEe/dejqump4jzYHOS9BCTlG6tPTFN/O7+
1Rlbyh9C5+RkR5eTUgIJXoevZCe9bU4USQpZ1zSa+SyScUqEFZ0SbKdX0Tu3s5QRlRZgQw2Jnvyo
ffhcXId+kyodeWo3ztR9OGvtzyljQ/6ZT0JMqQAgb1UQ8zAx7CkbbMNk13/1zT+hS8+1pJYmEUL8
1ZY7TuQqWrfpY0uf20xnNTmSr4TbGUQmuE2X6CXINTE6lwwcLKlfwtL/euPuP5rv6hNUIoemo6/o
wtYFH6itHTUDBVvE8FqCWFn+jmjFj6GgfOZoE2HtQIe8DV+ndiWR1FwOygJCKLYvAw3xvOP7nFgf
f1pyE8Sy8eVg+zYo9/HaGEpDdb1PW3oDol1fTMWAFUNW74RhBupto7vPtlFp/Yv6k719ev7ldL8F
n/jokftGmslNr7HHgScrk4jHY8hjg35v7jTNsZGYoG8/FCWFYLRilIFqQ6Fo0EmeEzk3VV+SoG7r
V7N3k+SveArr/RHOhV2P/xjpy/AVgbInPRkJ2YJgvQ/kvnumXwLkA0Sh5KpuHReB9Q6Sm7WHFQQ0
33QLFmEo1LzMa/hwnLyGpqA8eovSPZf+ZbFMk47qhDhz4viNBxRn9plIkcOlVRRqGG5Yad8qpRvc
OgUPXC9xrS8P28YeloaSh49slCL5TgnzP16wsCn1odTmwQfS3x4YPJUQ4EUrkjCBw0g3oqRTU/R8
2oJlcfeZQrG9HtWNZCsJBhwX26RWcmbM+ZHIx5ID8qoMNf9z6KpYNmO7k26G9LZBeVW1/fZgdhza
TgkaEGYFs1rHlTD6tIIp8ebf1VaewjuV0Sy05gawT1cm8u5hjDkMfhpH7bSOwNd+MXJxIH9ekWpS
bLdig1sAIbnImrFylq498sbFbQmb/0UFuWcYDVL24viRNtIPi98vjqZNeg4z7IcRqEq5rjgCyUM0
/on6tx7h7s48m0Cgu9pprXU1YfSl+9cEciicDpkszzxz26VSXWwLr3KWESd8kr9j6zhkc1/BRQ/a
ITqCVc7kg0SRfN9laQ4rPtAoGQLXsazdVNkExtQVuCYjKP7MIVbF0ZRb8cQbAP9yr29dpDAPAmbL
/tILonfD9jYtKdz0YNV8RFgIwumLNmrMxtG0IlHquTO6+UY8RIab0VGpmLIfWruGxqawRjiAM+tk
C2ZBxF4qxfvaW3Xh5y2wuDoFQGr9DjsbAfHs3BX1TE/MUE2Q0vGVLAjlYZzG1YV/gCVspq8+3S4m
c4I+RqmEYIQQmauTxwGLbDaOwQ7/W+NYXmsLgtVEuaEjt460otjWIOwaFfqlJNgWUGQma8f60/LS
xlDdNlX6vyVyVpJgpu9eftmw8GlVWyHs7XY9kSi75KYWzpsXzDRYbxHyvPKMLAA9Lc7P8ejQQAK1
tErfteuKWt6fW4Yy/VLer+QqIIRUjwB3Tzj2bBldkY2ZD4VEi14NchUhOQzqWxFzMvZXJKAfNZDC
qIcYxeWolBfbwIBX9clHlbGKNPBbBkEZ+gsGwnMvXJPOsXHQPrkDuyAy2JnFaj5lYT22Fdql8wub
+PngH19bUvicsmG+h79/bf3i5qIkUneVm8wSaUAh27an7PnpIP5yg2Ii1GgaB4efY+ijU+HpCVnn
MhO3R2NlqH4sUtVwccfmFG78tz07HUOKTPgcIfbUOrvWA5UcrHZsiiD+UXoTMMQ1NBsxVd6331n2
gwoxcfqT6gnHhbS61+le86d6Kn6AkY3O64IQDJA6g6PeIAmcjL9i8FlLgY9v3eAJ0QFS2hS6B7yx
aYpF88z/TZe4tT4eLZmtfdedYS/+24xvrmJ5PjaMCE8QgwEvLv06ygYmS8cQM9l7LFba9VoZtcF3
80GrZRTPqFYKxUlLkGnMpB2HEe7hXn5aObvzVOb4GLYsHuFzuow5HLeuu4g69i7GvdN2Ztlg8ZvY
w4kx6lvZDexc41DKBFM9AGursoxAMGaWCsIBlxTZSBGDeD6dLX/mjJbs1Wv2RMMgF66t7/W2pJPu
ENwdJeAkTeHneIcOGBDG5TA/Sv4LAIqF7IPha5ZY77X5IcWj9XPsyfPhuSMgphr17ufQc45reeOs
WyFuKs38gPaZMp/f2jd2+0yyF3KVGsmV9+wazrf7p6DWMU8Qjw4MV2xP+OIlXl5vC39kn8wGnBoK
8If2MOAqGeLaV4KRy+VowfWkmUCXcGC4IlxUBxSJnZQtAmMivrufCJLS4ujbKeROWrgHvfS3gNWC
00hSlIDIltv/MD/I9X+hi8BjRAFQ6mgy2OLlHTA45E8sIiGhEm3k9l7EmS492HAkeU6717BU1YAC
7XnH2Yay0zKDZ7Igw7vBxw2CoedOGTYbRllPGZt/4FoJmzalR8ze1yasrBYvfDPrUnfWIssOWhxp
PQ/tzlXfqPGuFJ652kpqB9tBhbAzxEXx1hAP01tqBDdvo02aakzOF0UmAHEQ37hhy/ROvSqAOcCM
5b5Iru4sKxN6Vk55pqm2d87Qhm3lZC7RXvma0TBf4xJiqf7eP2ogDSxHv+KKb+qMfkAcX7xKyCwK
kPxUgvvbmrtOSXOXEsQVbrGnwm0kt/mydiqBZ7KUwYncdwjQGU2WGcQvQ6s+KbfSbXUjuxspOLZI
UKcXfRAwnkJtzsNoNT6cjb9abQD9daZcAXuXLfv1cgkycGNPgUJYEDQhwEdEDKWLI13GAcEMK2D1
eOxgw7NmDgFujyp2NObpaK2GS6RaDakdVmvOo97Y8uQzItxd3W2zipvukULFBlwvhrNVpjIbOCwF
CuXeTVSo4W9HHMJya28ecJnPaWRcggZo86WBhYGzmWHy8IuaGHFare3/ejsikBf3XQnCSloMhlg4
8iHlJgWOtAvZm+qFpMhQAcGBMFJSPBM3vGc6WHcbHgTmaheVOuWfzMWxmnLJfmHi6z3IPVK0Qz6g
ljBkuC6pkMFksUz29tipqeySFwK7GA3s82qts2z1JsP4OIrPCPbNJR3JFUYRCg1Y7WZS34EZRPos
eD5eNeqeEQlqIZVambQeb47Qf1NyLNPEOB6f3hMWE5OagImKxM/xCYfzJfSC/buj9Rgb03Li/6KW
pAd4ICDG5hdYGXsmmCE+NZWr2JC4WFI2GPgUlmGuGRanSp6Z5lo3If12Jnii8cth0brnMYiMpReh
14kZF7UXKBcjC0KjsR8cP6DUmoBKWh5DLI1anyZVDcCln/jgFPT3zWFigqrdKiHPqY+1CWEC9Pki
/UwZPaddXEYsev2M1xEMSTpwjnkrL/1Tvsgd7kb39aCWK12sR4V+GN/cZz35CZ5Mijem9VmGcZTB
wjk8FbI6ntNe+zeAEELRh9ldIKgzOGo3m2LEg1wFBTaBCkaNGT85Vfx9wdm6BwAbKLg7bPV1ntbb
TooYicUfpnfME9x5EQ38SYKvg4gd1JlJqh8iQm6OieFINOiRPgQlM24/u5ygj5z7znOXLfNLbAe8
eCBE47e5VHSqwOpSQKfAAUsjxJqhBW7BmN1S1SuH4zlB8lKvLrCrBCI9u9aZmLjMyfC1/tR72jDR
K6SDVO4AZwJy9xoADkubXxog6bI+hKqiVbJu/7Alff1oxMc/Mzlfr1Vaqse+SK6PLAqTdtjmuUu1
w/yLUCG+lkBj2Fvqw8+00iFcaGO5nN3da5vO25ep+X2DEQAm9EHbi40ukZI7y0NdjPBgoYwvq9Fd
7FSu7EIw8hBrEImQBkXJR3X65Jc0FgVmmaNnhl9ofR9wKFm6+7TSSxj8/H6xodao1HT5ui0+taJl
ozWcLiFJQ3L+UgQxgcMhJ5kazXuxWgSF1czgdLWiceshMajuz3mauApcWEM6CVyLHhOlZhZP6nNN
RcBNDgdxhA/kJ9n17yIB/RfaAL89a3GfKtJ3jjbdqgdIYAmW/pfD+pKlQIZih0B4A+6c1y38TW52
Smrip25UpAfBn+4qnMZ0+t8CFQp8vCP8O/fpD7ZO7rS9LdfpDY7E2LZlHVyggBL6AaCb4c7wLZBd
+on8H7eF0URHrPLwvrw3PBMhY7qUAhx97DntAYNVSNYoQE4PFQKCri8HzhWXtwmYxFaai8Ncww14
riTBMgQTk5/RXcBOKKZ5l/aNhBgRzM+T/U9ratQKr5MaJ6JV4BuzsQtj9PzMADdRNuFEDSxyW02c
UahHELX4KCYIW+JoCFKq7hYlV7m9aBI9NDwu85hzaiYjJcw1eApTj6NusKCZlUDEAT1Mz+71STv2
XQqRTc9QgD0Ai6uC9nyf0rgTAoFL9TuDDT7F2ERtkTIOFacyhdRyljKCgmVQmYcHKqLx2XHnBS9A
S65Bpo2aqECBd1RDUmHlDX7Xb0uWXZcIxem0hGDstOw4WWTgYYl/dYrESkL+cNmQhCx3OM3eYbnc
ElqkXXIDrVm8uF2WlHP/xa6rfCdWSGEyz5oZCT2Qb6psB1BpATel493LidQ3ifSgHbl260CTKbQA
WixPWnXSlZDzTcyJoKrKgg4cf36dBlonX98Zl26DUCHFGPxdopzWgdlz9YQlpzus6apvIOWIdpHF
pgboA/zR3q49ma1dukmtAGTFXnrNdSREHoxqwagyWQHdYV+m7lTLqlQbGyrRnUQ7JhJz+LR5+eWi
JEH844/V9e+HC7MDdDptJqpn/eAMVY2G3mmchsBdiCyuWxrOcfFzjeuThgk8onza1qLp5Y2x4Xwk
TOATdnrcz6C8nmcBp8SAuy2M/ut9iFGhYN7ovIVfAmTq8zHvJOwVJY7OUeUaMCqAWMYbid+f4jgz
1I9gk4ZVzTNoZBncLo+d0j35lFChF8mSRf2wT6fqjLpRmvFHagVoo7kbsODFUnwnFTVei1DNHSES
o0Fush14BzjEOuxAxZr9I8Axo2sm+hSGO12CkLWikft4ImZdo90SaXMA2CWj6Ep9JVLSzZeJpOQD
BpEQjP6mPmNuMpMeFfXM9zaQwi6tJAOzttH9qQKpEBuo4XDvRoddfmqp280C6Y/X6tPOklxK9ubr
cI/wCOvkeNDiKlfwhxZiuIiSY6t6rwxDCMoAPScYR3+ZGZutF3mgkL/lGKAdjiomX+COni6ssgOR
vc3JLpJHt+eWkyUGN9Oq3HpVgpqCtYeSDxwwBUECivn7okN47ij5GgFdYptq32EKVtOKeJVCUFqv
DwGG1bbMFBsoc3x+YiwT+BH6tLYv8rW1efQ3SrgIoqWx/zAWVv/MH9HSeo1ol2tery3PT/LVllgy
RSfRVWSS4mz6nwzMV/E22j4ZEhnEgrPwb/La3EFNaR5VEG51jVJ+lFZVUfdUaUC5lDzoBWLNz+Qk
ocIyewS+pWABkr5lGCtK6HtQ8Jxg85ooAKB1lihlJJ3JvGi7rocb5AiNvRHlIGj+m9/PXqn3PC+f
dyX9kdAFhMlgO50OZqWyRJrdyYrtF2LbY0ZlP6MBjapEvmGHr14FlJFb5US8G/LBADPAkGfyr0fg
p0K0iKnfc/67yMMV9/xsEQFZ5w11cNK0h5fXERPk16mulJBj4Iz2BQL1sFcsBXa2ZuOaVIreVA6T
dmT8jtaN7VJN5uaVKyg5CDnNZz2pV1oPf1ep3mzwLjslHWEdZ4BaaXmhT0sSbe9YyIxcZA3Tqb5x
4zR0ym5OS6RSZNys3ISALVqJAunQ7kaIwCZTybLKwZNQUcU0w1KNP52PIyyuYW7TSZimnaEa14/S
l3/wOK+u206HrohbjRUC5D5Ce3ACccS9JCd3tdimOBCKxiAOaqKby1aQt36i8iF8QXnp5Otx6x4l
rIoo8k2HnQDZxlUEma3nmhS7CNnkN4YIPF/TdwkMzU6BYopJAzcpV52PNULmaq4Kj0r4tzrB00yq
eBejVQPDn1KpKLCIyYK+jADMK4CdJBZWTifO7isbCpucAB5HuPKGrbJy01Puu5IAQpQYra82ix0F
r5r92KdMI9q9R5+PofAScLPYN4lALN4nCTy7RHlfqytnvDTFsrOGyvluUq9Ssr6CRnqpklVuDul1
vcntevDuA3ytH9i91qGedzscHURMbdSsY9KO4EvW+NL6iTNk+Mt16bFxb9kto4qFtFrcjO3gJYLk
qebi2ICh0j/Qiz9YvtWea7KZqY/Njg2vwVp6hfJJUrq5kS0BxL4Bld8Azb/7PZDkjgogIs+Ic9z+
auZ6rim7nF1DbLLRrJeFcIV9B/5X7igpbX5URHhRwBBYrzPJIkHe8tuQ/Fj3Vwd7Lv7aUS9sscnH
ApLuf8zolKoMS/cCJEYtWHBI9jueV8zgEiYH8ezw5v1JYSJhfxIYzpAJ06eMBDoMbND/qSiBS6Yk
u50A+SbHNGql+sEiVY3oZj9LtacDNvPhY9wjKkWUsFT4eCds93MHq9CXaD0bduyKOOc70sDoHcDQ
Ywj/E80ze2+bdMpD+x7+R6zY/swb0O8RIRDm551l8h9il7jknXaHporlKlHe7sRrp5OtAnayQscT
Dl+Qam/sMF8g11Vgpaj/clbFJhLQzieXBz9Ty5V/JKwwhCyMP4KsNx8V5EaaQdgnI5ZAIrCqxhhi
oUaBFPvlrjGD91A75gcWyUGRctnbhxkGKuZkdJPAyeSh20KMX1Hr2NtTlwA8QvLPVyARdtFMtmSo
bh4oM2OQnMW2oZgQzt6Hg0TUGS9K23DwkzfAp0/iJxvHQbbFNn3Xd2QQ8bzyDz5NY1Ye+xjwTDYX
Q1Gb2bzHrgEYGEHFFBtdCkBUCX0H3R6iAhk+Jag378GEertk9mYlGk28dT8cA0wPaecNfbNI+jWM
+Z5ZxtO8ldAN9KgKhoReYmugo9IR++muwp3mGuxvWG3Z4pI6zE5KLYL34OBQVRpCzPrq8ObK695s
MN9ecTrO83VjMtGyC1J293zzyTxQvB3CKB7l/kIZqi/DfVZbSbxe1ULoPVB0CokD8DbFlH/OBVi4
W/FX7eX3M2uDnZdgQ4RzWtpXHnF1TnypmceW8gwk0rewkjIveAusi44PQzE9wrz6Xq2EBYQFyvDm
Nob44NO2bmIO5fejZxzAEV+gdnCC0yOvXOy/qxeEdnbPQ8gDyj4+LAWaXeNRsbokAvCNCmXQ8IYn
kopmO9iVCmq2CnZj6G6V0qCeypx8psFYlOG+B68J1y9COjmJMvFes2NyR13JTw5Tc+vqj6baMB4F
AOpYPij0Yk2LqFcPGRGhFNDhCzU0PSk4nMpzA7fONtiLAFtjPySEMJiSEIJqBBMkUG59Pzj1wEcH
ru0Gwah9HPjoQhxp6b/2elZi22G4wfW1xM49vFk1SCYwG4+E9etSb6438EQ7iOAHGMCZx+mYhqyj
GJp7Cn2h7c4O87KkkbFQsn1Y3FU1yic3NOyQVuC6O18Hfng1qV26dJy4+UXWYzVHCefE1Ngf43lk
woMSrA0sO6Lx0hqtbWIcTDHTkeHoybCu9KlONAhe46Pqr+K3VnIGxZnnfVoTEq5g7RStPWlY9r8z
w1xIRu4Xz86ulAL7kVQNbva41NAmw7SGXU1mw51mk66S+QJTxvztdvFpiuAZBX0lEgHQY+fXbW9F
n0zltBof42oCXyVMhumNx/FkXcKw3TmvZ1sJJgv+ggC4ZrPDDr+LEprv+6DjoBfAYnKWBFcWk2zG
mNQZZD9iAtsE6vnNLIInlcYFVuVPFHvxQMq7Z1laZdnVHd87Z0YesOtgI0kDq22DUV2VHXT8V2sG
c1f1ErIvoOI5RaQTpdvsWr9EeuOW4i86pi++ROM60X8GNogViEf9iIH0cLEW4KpH86DcCWZod2Mg
culLtYrdKsmTUqLmmyXsOSXGrWQqi2IZh0dZ7uS2m+jWTlV4LoKnTgitj1QqHlaiG8D+BetVidT5
LbCJL1Ool3ADxdjnOkg9135UVnH2Nab8eYF4J46+fFEK6uejAGO/b8S7iZ+Ee4wh1HglTzU5EsxU
IRp3bsgL+OgmzzohRstjF2BOFD5/8g87/jRKbX/j57iDbCRvAnPRmjaawSkdExhJ5Gk7e3/yuf+L
5Hr8FL5WiLlaICZMxnVNt9abjpkZU5UmAXXCN74UkxsnH29Ed3bPqF4x59YgG4RGUCQNJi9Ckeq1
l8IjeTakGUBSc/iTSSmoUQpyFgpNzW/tWObBmQTwlIxYJUgiWdjH4ztb/vBB9X/z8A6ZRkJHlvBu
5YFX9ZGH7cOcV+l/Ipb/3EA6wAgJuuJS7RaUPaPxSMzAAiFcR8PkRdaBVEa/0Te2DCLj08qBNqEt
HkLP8NMqNsQJMgoFr3MTRQOvYQiIPlDFktsTqgT2hfSC+rnerCCRMHSAfw+bKJVtNPohW4sChLKQ
iEPE/wgopcfJ/dEz7PzNlJDjTU91lF24QNy2zzr4UNQaSs28Sih4OlcmJD+t83S4jaqI45jfKvM+
ell8A6V1eiluHJNVpIczrhs5OMhzgkHR6/+DeNW5TNukd67xeFO4tXjx4HTZieZuJz4w+y03bgvI
WwtpsG6/iZoG9hrqtto8roiHlpldVi53yPOgNzP0gEqgIKyFjS+e/AqQIwunzbVC/nlt21PzwcxX
ocxdjcmhtH7fnZYZHch63v5l2xS/rt5KWz6uJcLR+MdCpxKOhRLvTnFIpNwny/boiucdJ+lvr69M
YpaOk4cHToqDn7f27kQP9up3YPQRKD8wYLdGZ4XUdpd2lEcwA8gpjT/ClJgdF20nHl5c5b0GF4HY
EbbWQ3ys5x/r1JKUy563uBW+rXLhZT3YoJcboLQJKmxm4uO0/CS147Q+GGgG0Y9dvjouplEnZKdu
Ptcc38MIZzfzUu/s0YaIVpJnyqXxAWWRhO6100hV0xnRJ0kTYVB3d4mNbU7t9PIwq4SvL7UAmlQv
7063lsrVswQ7mpNQAn8VjIc+ACDijY/uvBMBzAPI4b5D0N9XTXXZEue+omfDvvoDmpHh1JYdtf7/
8V/unzRh8sDfG3rIAh5OCa2h0LU1KOeQwI1TR6lKGKtX4hh8EfgTpb1SKpufCrRCvdXf0xOgJSa3
N0pOw7S86QoyAMBQ/kp4Qu5YuQ+ylgllXKXtLGTMxsqtMT6aJqubdvn3BiD72nC+TlA/8jgHgjFC
cZiEfT6ZC7OlP47DGxIUres0iNR/JIcgGzGDKn3srsXO9T0EKJePL5yyfr1SllPqStI3Sep8uEvN
U4A+mruAE7/xE4sUsUN9HeXPuNfJZgLdSC9QMx0IzbU+EgmVijKsLWnZac8SVrj6Tgv7tZialZDv
tRBVwDDIVV5WG/rle4DLEgCzS1/EeQWrxhKEfVegDX6QUlvzm3ylIX/Kla+haoP3TEOlVQuB+iN0
GJD/WAWi5+8eBu5TOcuJ2sgRl/F5bDCmHiLvw16hVoW4pXSCAraqZ3uOU5GThpR/8/3CXdWEB291
H5irNzFNv4mT1cYmpDFr1d5dqNMW096DDurPcXRlCIuJk1uj6rMVmG2xX4BuWaZF01GXPbhpwGgK
7lpm56NqqMqFg+wPAFjTOUAiUpoH5E0iRLy2mpOmm9ZZEmwsnDMt5Ktc5LpFsO1XAjyZClfwkxGx
eGBbdWQfMIJbFwc3Gh9WLGnPBViU8Z9+gpllq407gzgC8G5fH7ODPWN0Wby8t8pvkSdzGVvpOdQo
S8OmcEV6kMR8YIn5r6MgidEVKbvEGoSb+8LwxpItsZ4Y1YD6QYpj5O8DbkmvULCndv45wegU+epj
qUCmyC/du6fMQVPFbNEfoDLNpNNwazbKipwFqJPXVkikArVq2HKzj0LhqQ/u+c7+3L1dKUXdnXXc
7ujvUarQHfoqN3bwJIyTm2J+CV94v82f2tNeoggp5uQvPIYQJBlZMhRxwGk7sfbNc1qrlp+FXf/j
HbCsA9/GsvU0GfeVCaKiiKjw9WyoWzhIMPO/6eMNscd1Ym7mkohe5C6Y/B6XBfTIjsLyzKGvqUCl
K481oYzuLYPV4Krq6v7g+DUT9j0fa0Dvsf8CiXeurGgh7kWOr/4u02bKm0cuu9SqScy699wrrizP
befs3dCAc6nKHJqUYCFve9/6bJNbew8kiJFpHhjXykH71MWecdUuo3mULeiEfOEAXDQWqE15JcsQ
fsfNwYrYEALZR0H4jokFFHXsfJxwE9kk1uz3yzeDz1pcJYiYv5+JFEYNOhP/+oMHoDR7Q6eBXLCD
Zs3rc+OQiteEB3MOa4wTOZVseXLTMRuqRgdZUo5uqH1HHmfgqNBnJIwaZ3wNv0n1kp12qTOFKlfB
2yUVkmuIu3fW2f6pkSGEXrprwoJ0kR8+juKmryV5qv5VJKeHc9SC02zNA5ULwUnSdWSjvW93sEAL
V3JAId7RHYojqcACmX9uekp32aPEXcceicBCtaWIYeK/gAosW1gfYmllyz6zUx8yxYYW8+BZht85
ROe5pBGo5zG6pV51c9Uh2ykgGIatZaYgxpu9dUhB06xqBYUyxnVYFKZX0zTe9ERCpsoxyIDBpd/c
0KjwOb0PnR8uf/nd/QkfJUJPZgF2TCWDtn9Bu1+NZp1X2eIQ9DBNDCxbqOIEFpEvhs+2x9ylNukv
IVw3fExYx2PeYR6UDdSMkHlkQnb6of59jKB8+RoULeMtz9qIryGy/0gFfSzwVCh4sRn01SUKX3w+
XgDI1x+hRTAc13D9HDLByxX5OC11ekiEkBIJ1EkFt9M5XngWh5FkTqc3/hDqG9kslYsLO9cmNUuu
dMxzDPoKaHbDvKXzG+z62hZZP9Lnw7jnVP1Y7OfNEp6hKAShF6movE5WyMkQySTTKly5zhyc21yN
Bmqu0woIk0Y0l4cgl+rVYEkSL+n75j8AqyTbm5DaskuKHMgx+S1H+zpGGewGqf3U7b5lMxMeHnNI
Nx4dikp0QDBqXb5ol1Zu+OEz91KElNjY5UQZ4QpjlYSUfx3UHNQmWIQfz+KhZyuX+eXwhJcNUBAf
kb99EgzvEhn9N6u7JueY+QwDG16/WZV8wYXIY72+Zo1KS6T9GDQ4JXUik61ichB6RBFbWKivETfQ
N4iTf4pQHicyfrQy+iXyC6eyo/nfKdYTvAzPfhnCXpsnqEK1Kq5+OlboIkv3FkgLuT+MCN3dIqSL
ow2A6alHD+GK4DcdTRKnCCDrDA7QkzqgKV3J+Il+KJdeF2LccjCwoI0sdpNvE6F9AwpHT1QlR8bu
Ksy3GT1+AFcw/az6VOqxs4hkJKcZjw+8BB6wvNVEfqgGmlj8v9lqiGRq0Iz7sXkl76pT8yVkCLQf
xIg6tLDoGKL8eTvtV5TEe7t6wyxTuV1Mp6O+RWqXydLzSPwdxl2lZJi5/7hpwIEIUl7rprbFODHL
v9Nt376knbVVLFon5pJt8t7okGVypvSk+Ulvk189mkHVe4vOS2qnaIstCbJhn3umzPLTJc9c7TYQ
4S4ZOuqBI/VlVaOWEdk92BFwh2bqK2SwA7isaqoNmZ9OsH2lyGCIavwRedqfO/dVsiRA0Y3qh5BU
Dis53zxUMjq7n0pJ78AM8tke9pi23UT/lgRYic108CEUBOpy8/r8gYosbHS2CpQodIMVj1AGZgzj
H7xI3kxznTetcaL3pZcR7hxXihX8JdUJ6eSkY43Y7r0uNwU4Xdefg4y7UyAhA44IHlZmnyvovfyk
xti9f0nxdP86ED50JwK/JJfCivwwH7b6UB0KDWojQdIEMmGVQwVySn0lgnGttWcFi45T78dfBT9J
ZBX2Ss55bJYl2lS7zyIlV45rCsyK/oYJKwRerfAedgTezbT4EDj/y6EcMb8bYXz5hyn0c+dvhxK1
pHshxOi4h7hUJ7ENprWWA+BsbdxMDxsEMgpxdbb0Jz99NNg2Nca66Hnx4fK2KJKSFkdV7bEEJ+fW
y3yBj2d9bCtP58OT2HObNbpgKtL/eFZhiNnDR1U7TcbfHF0PNbVvloYgYwXPi0Hqzc+idW8JQnpK
HyZr7zIynNjhVB2yuatkKsS5f5DaV09AfJZPE+ORKAB7wmVjUbRZP7tY+Ho5lVWuFH5xH3a6mtsd
19UnaXkdc70nyO79ojOSDPkc6R2VtiIslmNtpGGI21qedq73nLOixnh1BggFg4SbrupD5iBHYWhK
HFdcDqg8mo7pKsHkIGelnW8LJxwuiQAhdjk55qI8pz++8dar9FigVjo7nmdFBa3NYvQQriBrhIaz
FMDlLJ1JcJq8FrzsaCnlTgk2OYi9vIyw0o31nrxAOTJj9RzMsLf3VOb0iOtCtytndF6AYfNduxSk
VbR3GvKjnT6P9/fmjtbB+3cNeDDW6LOVdsmXE4YF6Kl1eSbLmL8zzWDeqAjr9QUC34RCOYkSSpNG
R5d7hrLkvbwckc0mhl5JeDSKLbjLcUYzDjkoetn1air3+glYy2Vlkc35WT2eZF4AXFZMcmPrZC29
E1UyD0Kn1jISPoxqabZc20x78JYUUuTxBdi42yXvSgqicYuLxA/8Io7OBY8FKG04Y9PBYFi/59/t
DgED2VJR5FACl43a4k3QXHdbToxAvfHpa8kKX36C6oRK0Vd8hianPqQncnks6Sw/hiXrAuY7wqAc
Qj6uq/YVzNtTy/9FBzPUtn5g1CXoBTdYXTBx+517YkIyJYO+1JnAjoU6kolfVLPksBeIIQrD34Q1
RiWkfHsl92F6G95SDhNcFl1bDLlKioczuVuBzjVmwdQeE3jiBNJdUMJnK3K1PSP+wdc+QtqJaXq3
QxwMcY8htsIqsG8RfLxkcwkWQJw9HlEjMcGi2k3XnNfFKHCQhGPy9eo4JyYe1eApYD7RWkxSmWHg
SEnw+zzoLmglkwcF7QBgPePAh7043QkuADtWMgEAIMUbgEgAOI7B8GdwsajXzzCk1bZdcLoE3c4b
g8AYgnbgbHMQ17DVTwGn2OBkf/RROZGOL0lYs8Jg58ltzjyYR0IjyT2YN2spO2Dr6dzd7SK4g0+J
wwv4UxP1UfamRor29ntsejvswx1VbluAIl+kTdyWWL43uwkFCPJV9bVBLmfpkUSm7Mbu1fQ94S6N
areJylBS2PziPBWzTkT6vogKAo5VZtzeQ/KAcPR5Ed1KPCzQqELLB1auv4KZHdlnshAw3HfRYB6Z
y5EfLEpXOoOZybbQLSHu8TKQtdHhH0EjJ3LMcVlunB6aWGAzLeO8tHOIG/0bKZ3Yd/aKebwoXQu/
zGwYTPOUoRSdQNNYFX/XezrR36ohso7M8F1cj81dF9MfTcKZ6UU4jhW8WuOe+rOYYgrxnomb0FHG
GiVYSImP30gHboQAsF6XgSgi2mtVdXD3uFsnb/lpJgGVnVSiUOwJ4OegmCuqC5Y+Yy4M5yC/X6pV
ON7E6NGyXJSLqNHa3zdygKKWj7I06r1iRH0BFAZFzh/8YpI+xsBk79yk0EiqQdyO1cn2w3pPlk4q
UMFdlKDbWTSM5mu0HKnzR7po8SPe3rXZV/3hOui/RaEEUj+KLZiZWDgblb7A3MpjBdsM/OFdf+jv
Egrxdrh0wiTk7SO6U0e2LoGqc1qcmTGR2sU6QoPg38aUJQa3evNwSulki0CGWv+pOBKCyu1WCw27
0BFlacGCf45MFGohofPJnlx7FxLjnTUHSfHZgrxfUXMafVCek73m4UKQoJ28iXkZkCcqlmzM3GM8
gzf774DAgYcnClei2sD504FcrGqlppBF3pp4GSeYnjE3eupZwHaUvaHvspLhMNIDbXHlQpP2tbkN
mvxNVuf31cKbz3z94ES2uZXbgefa9hQuDG4OeoP8yJCO0A+fRK8vYCkg6a+DjAOBWHyHRSTBtODl
QVRPvJqqPj2Ruy6sWp+7roPgraER44tS8epdL7HeyN4Ls52jX/uBRwmh561w0QP4oauA5LB0W3bS
j+qUfnd/CKkEsYZ1oCiSUsggvPhPrmFCbHfsUUg4ugIa+Po0pvNEuO4NoR+bWS2ZmW7MOi+KFsl8
2cOnAUfadkTs4pF2v4sICBuWU+vLwc8opr7z/2kYMvBKK1KpeW+TQzmSunnbyx+8NA/MePyx80mF
WbGhC9PLjFrGLkTjpc5q1UVCocmO2rHi6rytT5ENqPoQoXYE54uhN8PuGwFoaMO/oIkrj0jjJyah
pu3pPT39S0rhJNhVXsft/aw7A6Ih/5XDC5CzOG85zzP54vq0j6NJ3Le9d73BKaA5y8UDAVMm8opk
bs7oWxLMubkWJZadwIe58caLUYaoNegHrx/jUNvKisdeuL11I1jP7Atf0i6xPKphpMpI/Q9HRWRq
o8fdQoHbI0WVFxXAiDfNlXQEquqG1MMevqDCLlOZ7BotipErr6mG+cnJ/DRs+qus9IwjhtUwduOk
rWxVzpRh4xNh9iEDmp4pCQGPWmzC6yPBBYb/GM5gv0FH0H2Q15vrRfbOf3iTt17TmLS9jyUM1zhC
b/Y3hKfs+W/YwxOq6snk6VbEK3eRRjMgKBkPAAe4x9KedwpXCjkdXOLNnfAABqF8DkfCVs+1sm01
QnGNGp2UZ5i8SQZeo1xLW0IF2PpqLQ/+cfci6QF+XUzXn+ANofZ5z+MjuRU8hz5q7IsoydB+zMEa
8fA+Sv5E3Kg+Am6JcpIaqb8R1IwTk9PIrBJkMqIxAaffOs/o6xBStIZPDO5tBGp9Z3WhYXp37uj1
s34OCZjaARXFoCI9QEg4lKsMeDwpyQP9oh9Wxn22+ooSpLoOeZLRRjz/Rlo/Q4PiV2pl558bWESH
Sr0MZS1JjD6+to0R8eizs7tsk09kPtRfM5BgiIQN/iG9RRWsAVYOcb7e0aqsPP1Ma9TIoDIgh2tu
pYvf4LvgiQ12P3HDVj2RhHnubaXNF+2eSCUFmn5NnoIhvZ2soAGKAeEGxm6WLbhl0Ag1oNiJ2OjR
o8DzTmCoARSgOxpUHvB33zSeCUnJyQpg/UYVAVsMpATj+z3//Gis897lU37swtMjgEoJmeVWw0LF
Y9GRV+eEJtVB/rrPQH5ffDve4/A8nJDwTdbO9EQXYQx6S6KExzhSthpEILqkES6nVi8v5jh5l3kj
EVKxiqDx9yStp6YANOFshL6yYfI5atYXbp5ZUMPW+atm5cEDgLY2aT82Vn+GGJJ+u+ZiKWHXmIbb
sKAQtZFp0VkPymKwtxKKL7sEws6OJt3Q27wmfgL+AzMNfzO0iQAD8QRY4y7BNjRBnLXiFKf6xlfT
zXFt5j7RjkHw8OOGzD6UZmxNnAgrdBRqwjWr3al1jk1aD8LT3WQuFxnwnVRQyVrHHl2Y5OhjYPT6
F0SpAfy5inmKcQHJQtJPBLGfo0fQ/cd4f1fwnFtGW/U0F64pM6aD6QfzIbDRPeUkTdXQ3sFAih0Y
DlNXfRh5PH2L8d8Oj+TPQxDeVfPuHlgWfvKIvqL11mWqBJKG78Ue5g5ddxtGgsAC46JceqpN9diT
YT1IMwRFWSVCXVl67LDODoir6gjfF444OVwh/eLpCnuv2KZUo4dNFuiut61EHM6iqd0aH81Xp8Rm
Srj3Og66SkvbDSCFxYcP0YDwfaiK1FWK4DdzTqD8wmYBKYnD46vR9p1l+wVcyHVQydtOyNr3AuWU
d1mbka+JP2mINfRs4LMnms7CfKSQylrbw2ok1heXS1j+fi081DVdJTmW7N6+ahOY7DbVCKbUfrbN
u2opabQfJtbgJHOY1rwSnKcJri15Ikz9OKPLgc3e169luKPjiKcnHAqSgEVAvIBUEiJxUVmE5lgt
yhRvnP2mCGFC+ULOadwheT+IS65awd7FOl19jP0ozPFmJyJW/jHKxnpfEcuMAJ8JIDl21eHkPl9I
Nq7E3U6bgStIAxPDT86urfUAceyTzuQQXREPPD/RsfmNPbgu3QdQvugm5KDC1RXOc4mf1vAMNEN7
B0lV/HVwadTstroQBj0PfaPZlMTH2yffq1fnYYozHdUvR4liSLXUnvTy7Rz4V31kmUzQY6XDylwq
H+7SqSEY6IgdFMy2pr61dC/J95TbxvI46QAD97eusJiurqFtYOs5lkegC5vUxVzfvUK1tRS8vmb4
Ocx2sLKimxDdiBw1dKC9VrqsQ1W6t9L7ROUEuc72kLXoATkE23gGI0JLgGt2NTsyeDbU1E3jObkl
M0kJoQxg4tIe7u5Uf5oC+HuZ7DqhhHSGxLUnAcjmPCcUzsZdCIaYc4iNhK9ZN4Boat+WoV/nFHM1
kXzjZLrqqNvdXkKiWppn0K0rhr662SNH7RwK0oRhGj+Aa3qXJdb2JEvkBhExFZZt4VBIPbC1GYqy
wE49oouaJRlkZin2vv6ZszPx7wgunEaM3qo19u0BGjzeMrWhGNsVaa6qrtLvpNG8Ew5UoiC+aUOc
krc4fvg9K+KAefDu9WskCGcwMj3B92i72Kg5ueFHlFVKwkxaO1vu3sQ9ZOytNaSpgSjsubYk1KEH
jTkizA91Zzq9fI+NeNx+0JNehafh1MAzlsjbAqPA/9FkWebt7auZ2TrZJqFXuau9KIuT4IX2qLRM
hdsGu+44Hr3phncYUIhRSX88wIKW35CBp0/zRTjqWTydaFAjnhq1iMLazFUnv259Ztj40ese9zzK
bypiAQAboy2L2W0aQteuDI7Xlxr3ErmvmIAKMSx15E5ngnSZp6iXY1SUjMZ03BIFqZmhg1ZYcAht
MIp2NUFpeLBGht5oQGZfWlghHcLm1vcANvBGr2Y8dqDHirFA7tg8foXcxGLmtyJRoEXrfmiEV6JM
AviRlD2ZVTqI49WXHSy1XZDGkCJdkXTDoWythj7VIYlSzrWNPOnB2Lv0x2QxnEbphDIhZfbfyEoG
kBmI81Dsdm4IHf5R+SRqeHLRW08tJKMWDI/baGSZqR+tk3F/91dOKkiLGdGflnhuU35qYrmhLlxz
c76ygFJ44Xvm54+hRLAEpd2l8xMdivHuK9GpW9GyNn04lJqczQ39Eyhry0hGCyS1dF8OAGcK8s4G
Jt6D7wvEa0Zm3orXj4pdvpQEhqDfhdcQ/BpARuTDbxmukvNqmhPg6IRcuYAxE79ebp/KhyaI0d6o
kXQepCs3jeeaCiBj5t6yQxoPzANwo9yJB5VPQwTTbkd8eYkXdsMsUZRomLfYXmhYTFXsCIlZZe56
jBCOw8Eat/Ysp/oIk+tk1jN6oifnEszITKNpVfxatf6nJG00uJaOtWRvKTII7QPjrY/u/DRkona7
xeml5gIoe7XieQoZakyB4hKsqDXCts1usxMGhf3igHuw4nPxYGyZtckqVgL3A4Bb/89ZS/j/ilqI
XgXkpSOgOhgOEArAgAvCYlCx5HHETAS+NLW+WgaUJeaZZUaPXRAypgWVl/d1rmoXwN3IaNb0+4Ya
HqJ4NHOfNcNgIAAxS1SKu9TpRGWcLf0CBQ1eXi3A7neyXo+quTvpMTpdgACPTl+9hglC7AZbhiJb
bwB+P9meKBu2921cDW1Bv5ub2HxkShPE3VYUzq7C3yCuKLA5spfezyQ3thesNu1ejDFL1uoxE6iv
HrUimemH4O04epMu7iVQNpXReZ7mWsiy4tX26MI8ebJQ+UtprVNMTcUPFSO3rbSygYCMi2iKSXav
HXRLlR7IIu+kVf9EDaK1fjQtOlpFo/YmWL8HGys5wqGnQqEctlohRPZ9Luk0T6NQDpEXZJyay+Sy
JJeDPaWgBIkZmMIiLwCsg0/xrx19fQlS98WFQcbllzGXxqRfKem/7889YVRD52qrSYrvWDmKypMt
/Q4khaXSWVs2/weP9sfOAJ8zi2wNhVpUT4FZF5jzhHmsG/A+5I+bit8KzDnX6UpjK0iX0rSVvhDR
fVf6n7SB154ocb+MmDc0XFqxSmtRb/zM99F/VJqrdXn+Bip62SrUX5tC3d3u5uIxbNHFr+tvjQOW
U+cFX5emWlSjX+cDCeOWMyarOod2z9sPE+gQj1h7ZB/i3F/3Bhk92Qg7HJkXKKEHKQuuHXgTP6v/
98XbFO5K2YmLVLUtWnoqDeeG1DpqfzmXVG2MWze6kLbnruXxGW1kczoaKyGb1FyNljijG9CcE/q+
DNyDEtG5abOGB6wwg2oISI46sQubKPB56pA6/+zKIs92+kUnRa6jWqES6LBvQaUe1Kwxkzn+LHNY
VrPnvhyiPRQxWz2mGwN9aV2DIlEsdcXT5+NhCUceJaNcfkfQEMyNUKClaHMM5sWoN8IvMhRFWk8C
3F77g2Q3tCQFZeYVoNAgEUH3AblLwiSK70QT6e4dpOwemMufntg3N9jgcrXvIzWIeBA69QHwcCVU
mRkeJ7yn8yoCwWWIISMFf8RNXb5mo/bokU1Zqdjst2twjUX2mmQN+BBTh3Yeol+kVkM/7MUd0Y4Q
/t7ya+2pJXS7An9tWfO4ztyvcVL7GA65hW57FRkyBjy33EDwrqacBGmz6VaZpBqMLpCkxw2ALG3O
Bb4uKg0wWp1iA+DetTRlRlCVzOgGgPQJrgCQ3uYd8w9gKoPMNQnSC88G8/DMkzkX0MufB7Pa0ma1
nD0MLf4rdXZt7Kkag2tf4YdK5teDUz+Obf0fd8T724n7WYlNMfF0gmuLy1pv8Z9i5nrEQzGBfsot
rZlsFQnX4ZlNiou3nK5QVLOQrKs+rB+eyiSiwvYhfztAPCFZsXGOrNcZ9i+C7q1TiW4s8Anp3sGJ
jOrZrazf80VAkmk1fpeCfPZM8GDEUN7L96T+BU98VYfpOPHRo39xEw1Sv93MTsbQdGEQ9QiYMZt6
9iIkMHsmmWOnhqrXcWWResmYAG+EHI71kU8gScBo3QaT7NTHH8KV+wpDUifyET78TusimEWDv8Sa
RXx3mY10/CGaMiifmd5BOeAQLQGSRh+J0tJAmqYjlvHobyFKP5w78JesLC3P1OmlL9wz91H9u7+d
OQ7qWma7JqDO1esn2nNwN6kgnCf/RVM6kgB6sPDnhDPAQPQxSZI8SLBeiOtJN7P3gISvaKDYqFaq
3Wen3+5GiBz5kT53CYV66f0bGNpbk5USobM+jI2jQ11vCWXBtwix3Yby1juPQwkndockr0p8kzN6
iYuA8yEgYazd5Rp7PXjgTjSiNPqsUuz+cww9bEXhGrhyas9U/p/auNAnZho4OKTp0U5Z8HAZC9Wm
7Utxg6addSpgSZZ2g5mcrvBCdmLQPkqzNqjnhWSiZI+WTL896LJHPKmrz3+EE0fUE3RQuzGnuCf5
Uq0MPzgDEAJ1j6zM4HQSJKCDXPQaCYH061sDF8u4IxqprlInJrFm9YV5Cq9s1ORKxcQ0lR9NYccm
jj8fxri9aPXC8upY3ow3mDDTV2o0NYlLvgFzCnluuxHEEsttb+WqLgxQxlVcelvb/B5GUAlIXg/h
ZvSJ3DE39FZat3CkQL/kt3MSD0xFLoVPvGNJl5GIUgTuzqUWDtiQoZJTIUdRFs0v1EmwfTn89dAp
2CwGUX5oiz4SmeOB0AqlC6sd1/RR7EVMVkGGT8Cy4eywSuGhKs6F9ZqS8WPxddrfpi1lVRgAxr64
1uPs5VLT6nMhyq72mo+/LXhZdtBJ86eh5s/y4IBRulCNVGTCLEcooBFlERWSzoYwysDcEEbiF4oz
MPY//T7kESNSIoBXqe8MQooui9Q79urNwcsJwA6bSFoWeSXdUZc8RKFxaiFw8BkTGGRvTNoCXQ3P
0EMVBKZlVdjASiNTtQeN4q3TbOJj8LVvSY8cMTFAtRkvNAox+AMvf/fEAuIgmD62F3b8S4AiCsQl
mCkzNWMClU1Spfd/jLGSKF8fux3NKL0479KpDtRDSkvyMD+84vaQqZWkB36zczL3/v4954G3l5im
eWiIQETdLOTHdNO7SYMP07du/EMO2louJW0zO8Zp343IEnWBiS+v35ou0Quj0lkG00R9dEsd3BQG
HZ3XYIBCP65E3HxkjIjrjo/n/wFxkdUEOwwgCCJ8Xv7LSiJK4EbAV/V3aGlBnPnmrPnEErZ9iB9u
KUB9QHpEq30SPbKhAmC175mfPJHns/m3PAzpQiD0I6xyYH6uyJ8OgL4bpargBDSyQAYC9nv33MlN
wfuqO45yxdpEE1GgxIfYDUTvivR/N2LD22kPZGLTxyEzOQx7Bb1ws8FVa61Hs2K2UGCCwGKbnR0q
8QT7WpOG6PdkffcTR32gLfvewkr1FmPTAzU9a9cWFKINwG+1PwvXAahNz6LJK+fmAWh7RlHACWEB
0oMPKGav4iygKK+zbmGse6n9usa+ZGOCaru5+91ex1QZTsMny9I6fiMQr3bL8Uknx3hIXCGYwpZD
yLOL2AsDSXvri9LzhiYU4rlV7k9qCTsIRIslW/NRzynDs7jsI3PcLf5ytZkBS4VQ2vWMIUUrCDuS
8Cz/0nUosYQHewwDdFPByD2XCHtVaomvBaumrMicfQE2zFXO7BD/wRm73G1JnLE5V72FVkFZRG3U
zH3XRmRSMidLRi885aUIJCavJXgHw6hKlgWwuzIBC9QzeN2PX17HB1/dTPJ70bF4FFluh41m1xul
ogsab4bFiAt2UKMDJnY4gMwbzaPsWnaBlhxLRQDYRjMIgNxql0jm6T/UgiITIeXruw/VDTMykVkW
pO9am26MFKlOqU+m6Pw9jnz2E+gXrQ0IQ3a4Eoqru1r4ALAQNMzpvPeieDIPteFBzSMXye1RyRFr
DueExB40o/1f6cq+ZMmZCul5WDYkKTZ7hjWNykLWdusvJjGboCy1eMJYQL8lqIitkRqJDDiGO7Ub
FdEviE+w41aO6HB/cocG2XSUh9D1YoJH3OCrxFjDRsMuxEtFj/2Ct7wgVk/Bwdi1gVWzPrbaJ6Er
CsjK+/utoDYh8qC8HH2EaSQLHkbcEAOMFlYZMlQiqCSh+2GvqiLxoNuPeJf0adU+lSSSdWdiOSdS
fimj7owzghYUDE48r7POsIcDPX4z50jrbA74BabrSj5VrrDNJEM6TjWsaP5dZAykcFvrLyMMwlhT
/o2q53I+cmg456ufiAIZ1BUYpz4bT9tnVTUP6B81sjA6nnlCyoaCa5zFOZBEHMw8NzZ5GUXRBo6U
DnROdQ1IgYXWMPO7sHIORQKxDP2nOgUdR1uAdRPBTuukvGIItEAGO/W8cfUKVJM3QG3YwW62BEmG
nbT1QIfdZlhPIL5c92HF74PFqOPU8r2jDy1zzPr+me26cZGD5jy62vyrrmQ1GMgN8vFlk8EnuODM
ytkWPWQKktPubhakRVSNhyG35kPPGyJdebsyW+sL8oH6axe0gp9V5w7IuYiIwC9L3OKYzaueu15/
WnvXx2N4n8vR/NKLAdu0fZb1kS6EVwwScj+3+KycGhudFroxap5ZZ8UweSPm7SQD/oLhrxLOk6fM
ZHDRVaQFFS1cNKTE1zvQnxN5AAliapApbocXpxiVw/6dld8xWu6MrMgO4tlSgNkBotZof6WPi2uk
arS7PZvOKvE9DsUGmDqAc15Q17SIHCoIzm9iCL4eh/Bsr01vax6O40M/NabqHBbAspq80TADDUFN
qp/IMAHDjzzGA3rdIkRAqR6390/5vqdYftVlRRzZ8oxREieHjIag7qRiJL8i7Kjuicrx8mglVQr6
sUT4AKXV6cxtmQyN9ZaqgXBXCXZEIHtZ4yPOxBaFuPGwAMpjyqAeWyE/KneAl1EsAEzoUa6z232W
Srt0ZM4JvkzF1AX16utRsqLrJTMd7qz+yh3BxU+aIuKmhNEc39wGIIQSPV8iqYYYn7bG/P9btclt
SlVqgMopU4JYyJqQuzm+PsaKAy2aWph7DMEl7/WtyuhWTXLaF8uf94zYNlHYVwt7hpGflm1LXCIi
RM2ph3terNyipTdW/UuxGUhIpOPqurdJaljUb0g9k+UPS4bKJJz3M/vFHVkd2trxUnp+iTk8+HWH
1f60PMyYYxjDf4ezCoaylp0QglF1/XDiM7XBlWSLNug39BTyDrTi6WJGyx3CIxh9vLCt2r8ubeKO
S9tY/lPgAf+EfRSSNhvzctw1fY24IpRsNb3PI1vtiP7kpkLFf49wYwr0rhj2V2V+UJyf0PS56FQY
bdcJbi6g//uZLLPvvctwAeHJYd//twXCQmdVWfXFGpND/smwvAMLpExfggvPfafUgkNtiPYgRXpz
TbW5HZmnusF668i9b5DNHzlwXGd/HM5SxPXE/PHg9b4/CBd/qjXvcnhBksrh6No/N9QyW6ysGEGV
3uQFsfeErEzJfXwLd1rt5EtaudzBsCvLmB/X8bswAnjrh+3mUq+YN59JNYNtm5lNoN+70kDL/qN4
p1/lM4fLXNRfSU4CpJIKsBRdnlT97ZPrf8l2KzyAmg17PdjoASmvUcvgFDtcQduAzGmiZ/L6xfZO
lOx1egir4lUZ4RlNuLmXC4hRAye9//WRzoryXs9Lh26zgn8hUWQJrwgAUb7Du2RcNflro9ZDJyzU
vRgZOS8CKtSjO3BcujPDksXWSObqxHL2o8zadJLtV1kYITJnUvnQ0tkR8XydXUlIWcTgpkyvUv36
ugjMQXMcDOmUEQgJQ3x5FrgiAC2jORnZlXtQaS2ZNanL2UWfosQN+es4u6S8TdT5za7os1Zj1Yup
cdRW+nGGyrmZtJQjBkOBl+nCOJxlmoVYkoBGzmvMy24l+rsHbTW9tq5q1AgU58a69HHBiNhyWgN7
ANXqko10DG/4KUXc3TNM8Nn5aq6RtNutIzynPNDqbHJPVopdUXWKQAZA3TzVFAaEME7XoOy7Lr4X
oE6MVNY2v4NF6QdFpEKCO0Iiz1mddQvXsszU9D7hAcnxGZz0/8uOlgzyaFb4e0cnjpH46TvnSM9G
7oj3aR4ZeBHu5Gd/BEed/XIhGwb77oY/WI0M6/DtxGVYG/O38z3bldkXFEYPr02s5CXkO6Uq/Oum
9k0kfO+soc88YeedVU1r84xECZIE+lfboVFfIhH72Fk9J+vbVinEiqylVhjoufKxwyRkCKAk9A85
0kpxenpNZIAYYtpjdgevzbxBf1Jvp9PCHdQ7L3PFqHydRHuh0s+DH/GTGbKWYxUXMUMbHOtQCZdn
04ATyFGD9e/FQoW7PJAdr9oPdmcb/mK0HQgK8dcWwRSWh2/+0qSLw4GIpUc9K+0obfNQ1AjF+tMb
iiGCMiDhEIXYwMUSZIL1lXehOvbPwyV/9fdt43qjvYi7R5+FPT2WId7JCLFRrOQ2SgzDz9ZHEyXz
AiHPltOTVd/zjF3upRRWIs5ZQFG0HOi4ttlDEH4YshUAvXZcnU5GA3q9WmzI8h98XKvJWH5n5q7I
tX9a5axl1+rOcX+V+DQKjQzzxIDhZjFxVcCczH5KMkf048ntDjFQjHCtMiJl1nc8rS6KGRFf2Fuy
RWsGTsB15G98hWmlWARPPUHr0u3V2necyHlMBTvdNT/7F3p+OtXJNt06jrJyC4CK5d9MSsJSGHm2
eaR3AyTYl66NGXJosAlNwMxTbTR+okTrsJSBrVRgx/5rlAmfQ0L1AIRsvhq62s8rIDB+HyCtXicL
8BSb5zCIPSh5p4ADnIR7ucF1PdgfJRpj6hMNRdTXlq1TWIiiaMgu/pu3WzWtDcPrfDRW9pl5FxgW
Lw2HxH9r5LyNUXqM3Pimo7fYZdvcQSTr+UE6RaY78+h14QKQF8oDL1Ay+CY0LsWiHtVF7gJ3IuLh
kuIkUjJRIhk7YpmLLLoCIHFvX/5smI/9INZ/eBl7+9HcPVS3hfAiwLRNgOQgZBjzad0IK0zKcteV
m1GlMA5pGFq8mdebnaQX7y20TgDMdTEs4zEiasmUMfzYTi4rEkff61fBi+HCO6cBL8L9rdX+r+ji
5CfFbq+/wIUm2GmqFIlRbtgrBSks1NIJHZ7GMC4Vi4zvJOEe+T3hR1+4SCVYiAw0Hhlmt28q7+va
BPO+G0lgJJmCEd5O/bbDA3qKy/W0YvhGZ7PtgKSB0Ud7amfMOXkOQfv3ZTFTUNh2iM+0xFbkz8n7
3aqm4li4jeGKGCDBfTgXing1sYLJ5x5fKFG6itmEaOxjX4CCY+oc000xxYEWT0MC8B9ikvwvqDQ5
PiR1pjHz1uSJkK7l8z21ckBbeBefVvfG5Vc2jm2DoVRdVorLKENtZT2dJC0AcXCuVLOtGECOfIJJ
EgKjGg6wkRj/Pa9GQtNGR8VhXKiAUE+9WEBbj79s73/4lfGlTrEWKMZVuIy2dkZE/qXMKvSttpbE
3R33B80osRnAdhqyttPYAqYuzeaHABiI/nzm0ZNFU7JgGxDRgHg6ijSXTYyOZGrcrEI4+H9Igu9f
uPobXk/5UbCnOOICWT/s8JYGtuNikCAxVtOFHWNwZTGlLAc0nCO1EVPYWWUt1OFE8TumrW4Ib/ha
Uk9Sec+HlLPVppY72Nc2dEWz5yqo31kz5PJZzfttoNGVX9kFyaLBoX+B3IHAHjDQYy79Epmdsztq
ehfUj2ctp9HTUjbHgz52iKVSXMP7jV0jiutZP/f92cYkrH3UOCnG3Tr7uwOTIvP3rIxe5af4BXBx
MYA3gGaHoaY0OFhCw/U2u/WhjC1gyoKmpx2JfPXSmb/xh3xzEtQaYOkxQD3Jz5Sk83Iy5dtEZ13T
2+95jw4ifkrPB0KhqXJlNbIBw1i+slpinT1xkYMjk46/3PIfeQ75lg/uhbUgpenxBBoqbZ6fWnJo
syZr9W14oCpQXsSUGWLKTC0FgrEtisEmyBfCpLbgKDW2CIGyzQHUv5O2YdBHqG9tfnKKa0pjRe3X
5j9uRnO5hhm0IW2tWp/NIsGbfQb2DciWcTR852dPkNDZIpOrtH11IjfqhXLDWACqLpKycYfVcP3C
Mpg++AWG6/cyCP/v4HbMSu9IIo3iYEuWjeYfIX3aIPRW2TpCRK11OmS9+xNuk0WSs+zVCwNRrLro
hjVpFFDURU1YoC8XyK51SPkYZMMZDQjKbvF6xns+DZgfUPv2Mon0ygh3dUuN6lupSLIaVy1n3Ak8
5SyXhvY9oi3/vgiZdkdSiK8b4b5p3rfjCKgPJOSY5I+TVfWY/yztwqEumEvtENXpAbB/hqvLcqqK
dMXwrHDIklfa8lsF/e872NnRy+FOBHq4BUKPCyHNqaURNBlm7sg38Y68ANwkt2CwkJs5C2djKA22
13c0+jreU5XZYY99XCyPeY48yAT/K/WtBnlKkhTHa7ouLbZbot82ZbDoe97Rw2evPGtRhaEzlp16
BQqBtmt6GZQ4YGX6uphIgpsBc2s+wp4EpKYzoCupCPiyL0uUzkDTjnSrh9nYfKL2Ke3Y8TEt9KJT
c0ljy3WiMfgTksIQ1F8t3g/4eC1CC/lhmOyYNuFXX+C/H4LoQN9by8OAjO9JiWdT2GdsfloJ2Cpx
Jvtq6SCPMYOM4LPZWrHc/vh/jvG7malm24wrYhFcHoXgGlkvrC7sd5hsYjmjUFBtrL3aBWQ/ZQ+V
DcR7Kyb+U92/yFFWm7qGVoRrL3KKgi1t32kzrtE7CbA8iPqIkwhNdeJuod5d3emFEoEjOZmnvRk4
eYq0USum+B4w93iGG2Jfa9F29SSAhLJZLzdYpR7hF1S2awOqzqXl8tU3bW8f7jAi1913E+Rec5QT
O/RZvg/q/0p+V/Tf3YFHedwzPJ8ubpFDDAA5+nIlodYA3BDp+icGNA3TCSmLz4dubPBj1gInSfJY
VNu0n4vKh+UjEKzv0jf45rof8XhcEKcopIPSrt1qzEDhpNbof05Qoh64pjm8UdKj0JrFNPDhQsqc
J9xISSIPkPK1r2XOVr69tY+wR9R8o4KmroW/GRJ5mu1+SyIxg7CDaa0L7vXbBx0DZ8lPRz0qF0Tf
tgPnGUdvYlxuxVI7kkcSFbPySVDP+kKpD0604IxE8cvyoGZstEFxgLOvHsY/s0e5K3xYhYjhrci5
t3pKHIyrT3ObNZDtd8Y5DisOxLGZf6P6C8EAjb0FRHwDhjscea0kqle7KEc+CN2b089pVvsMC3es
tjiWmO6YYZdF+mS7+c7S/r5fHJijqE8CJ9aDiv7EbXdMh+AMvNXOJj9loW6GMEtP1b3knwZlvi2u
NTeTFyOegrFjen1od+kdl4MpiXo/3GnTFTwDJVIeutWZ3jCqAKzfyRtUdbk8DPqlvfAu2vTQ2bWA
KxHCzdES3Qh/qCQrIw0UkyhMD9blr+b3jnPWuWkrcE/aeRHNSa6J1AuM29NYgrYsMmtlqDXsAgVm
VWehfpcTmlWmUJ/2BeKOfpjFJ3soqXtblZglZOS1yT/xYkIWkRkwOhKy8ZOVbxRdzd0o2sPK2E9t
O6aNmM7O5wb4Y+fpnp2ubQ4eTIOm+L1jAHM2Xb1hAGzI8fmITinC6M4qM+UR7AWnCiunwYNO0ZYf
QX4SA4bvOl6Z1LMwvwZ0dqoPR9Kte9kXlylqRvYYB87vaJRUIBpyrK5LU8Jm/+Oq9nLU5LYCwFpI
bn6m9EOI8BPAatIYSh08i4SiRuc/2uG7P8jmCnXKcXsv9hQ8txboLKwvMntgCmH2CKwHDp2GTiJ6
4CgYSPfl5vkI1kX2vBhkIIhvmk6wrPSlYrHlJ4HNHWOXNsMqB+8Gf6ayx3PmaE/GG+S06D7KV/AQ
gOxjr4H6tjK7iiYQxbrI9gO+Z5n/b3JaBXfFhTWPdgi/Xb6SmVlkp4/IAZlOiYnzU7+kGgyMB6Kn
5ZLXzIkMbt2MUvvATZ4pfiSNOGRIuMcJzdX8iUlWuPIQdcRs7e2nhW2TY2s3EM0J9nxTevIFq5y2
yhMrf+8fHdYMoulMpse8a7IVc6//oU64eAfiKgZUx3LubwegIEy+yD68oxKE5MaTElF7LhWBjXo9
NFF+25zHflzh6xP+kVEx37nIXg6SQ6iouhKO5QlR7KIm24Zl4BCxxh/qr8rLP71KWx5BOGvOPEEf
6TvW+fHTiKAc1tLcrY32No7GpJOOsupyXvlhO17RBen9P+otvwhjDXZDujVErtNIBnGBVSbvhY8B
oOOL42RZpW0mlMq4oMVmU7x2R3WHqnviNRqduGTBOKG+rjIoIhnMN5Zc6iA4oOKQM/VwxT1NnPzq
YTD83oyaRvDhaaH8b6Q0w7P6mPyDKs0emf85aY2rIkFmaTFd2RvuYoIMdo0hUvTlR3zSClgSq3yI
sNdrd/eDvBWVpC4fQiaUSjX6fSDAMkm7FgVxpbKMbPadwFD339XdRWzYpxu7H69stOsM47UefY/5
/7cNKoBPyWInWu+brUvTNmwANAllTG7ekCatA15g4GJFzJ0KsL0Iz7UIZk/P7JFLvmJSSB6X9f7T
EKqqV8XersSN0A5Zu1RyZQ83uNbzqYB9eFh2XdeTVW9fjOLvvDvqbHewq/AwjgWuVhtonTwuRDOc
aXM2RmJFzRP/eAw4uTOqAx/seHmF8tnkJhUTb/yMlW2VamJln4eBAPXIzTjPMPCboRvXvaslwWAf
QT2Ip1cEcbNKSzBIqmnoC/dhuP3PHAASVetyUQcos8xUyEHXTaXR+LQJ44QYhsLwQjlAWo10hVgs
fWCgFr70091h/Jk1vKaQlLDtRR1LatA0Rz0s5XE8Try8FydMsTVoC20yYCszbN0CLMcdEPgueiQ3
2coB57EsTL0FAAleLiwGP++ryNmavwOkysJ93makh6BIfc7+xmFf1oKrChqSFn+rDZq4fWfmrUPa
SDMpSA31W9NO/h4s0Mf0e2itnhkTaSgpBYd9v2z6RMYQXeqECzPc1HQgS8GBBAAbLuEh9J4BfK9Y
h4E+d8bvAx/irRHuxQenI3zkbx5l8wCUjo05SH1wM8gsy9WcE8cJG/LKL4RRasB72uCDi1rklraS
n/4pspM3VnwVSuuITq7dK0SF0az02jvEdIWZm/2j1l5dMsmCkzJQG3vBIgCRchUx4o9nAb7YlQdl
W44v/EM2o5sERgvRNDCtg7GAWT1HZwYH2ENCz513mquoWVYlpRDy2Ds4I8zdD78vcvqumqkTVLKx
G05sx2Yv0wbocb+a6Uv5j/0T968jxba+CVR0ZpZXJT7umksijO+PJDatGBj6K54cNxsT1gTK3DqM
+iEw5GMzAaQ9wRXn5G/1SQxwpcp+OIU1nNqipdT1Ke5FDBFBg3XPa8UDxrXBgoX+yflQ2yBV4J8O
VsisaYNZNgb7HPKVEaCdQVWEjXMqno2MV1bY493xW9J75WCz5drGzmhilcdTMOoJdN3+EKr0YvO2
FuCwPpFyxi2KGGLWpED8WvPmsA577Dj0nxaGP5UhRdY5PnL0PrEvdWemDpflImHdPoWts2weIPQO
Cisr+JNYJoW8BYBAdhyCuOkWMZ5t6hmWQk3XDnBNhWJ5gz/GzzwnDr0hI+ChV2OnpKUQ5P+ry3vV
Hko5hug/cbkxzh6+xmxASgaaP6ZWL3QR1YXoPkgRvf0EShL2bYLKTmrNh+ip00TgkYhe1JWEMOHc
989e/+8OaBnm4O6q8Ll9UjfK8gnzc/o4XVyffLair2zzBX1uChOmtKkcZlp3edIicPAoyEKmKq8J
89XPVONTcVloUlBQsDVkmIMcmEoPPFoQeaBm0F/otW+0MRFSQqRge6Jq8TSpppUQe8ALWNcnccX0
4Na2ibaG13Ote/4rCtMsn4BZqY6tU75MxyWFI7pwjphFQ9Eh7e0NRkHqaWV5uw9UWnU9DTYmowSv
YnJsfiUOL8cFwgcUVhrSEYIVjlnlDF3cVeuHW4qOOAsHATWyVFpeVH+USiHdlGjYJetDX/G7bF1M
jyx7JP4QPf/WyVygDBZh0vOVU7ZnB+8CQz4sPb/ylXjWfsykN/yTTRkPb2hQbqmy26/JOC5a24yi
Y3yYKOe0Kn3q95r4ZJJNJfXM0rj9U707+wVk6IwDZhdNkFbYI+8eU8WBwIDJkYRViAl1E/j/bTnl
FV3ft+W9o78jGEq1D2D+SD+Tgnwl8DmaCmZoBCsKLQgifyCjkC8ZZl+0ZPuSAlylK7rG03vNg/sb
p8DSKyy769t38f8eML+ESHi13Sjn32DF40NfnkI5KdpxFaDtbV2I+tMIXjANPv0EStA+Ca3k3TOL
BUhX9FvC1QG3+3OWULCmX0pvSpFDfg5iU4O5jdKFyl3vW8XcuH+0p8nWHbHnkpLbUmLyWNU1PE83
rPFRPPuQesjasPIBtguOLhez+1s6GKuEd8VSpE6RxLpIEX/M+Z0IM/0aYI3kfMAiibuglrnOHh6N
6qgJTX/0ZmaN9eH9KXVbOWN2aROJ6/cm4rmOHyUYndXTJ/rVU1n493IE8VMQHbZq8hcLlo7NQc9a
HYMPJtHWKP2dM1VZGQobMPAeoInM1XpftjqO5vfrzH8taBirXGyh6XGHTIuRzZIIpMBmbRNOT5/R
R4ihkpzD21Uv0Rylttx6NPWXRtYObLQe/+k8CkWJnpBqsI5C9RbL4LBs0An+XpeLxzYuzgTnNWon
QzGaPRG/LsFVx2Ykm2N8TLj/I3kIopdJrCTLHkEV0bXEbJbI8dg8jjPmANJmKeezSah1KL1Mix7l
PdLfU+gGumUQy3EyHCJgW06PYwUcqhoDWC2wOkkiw8pKzYkjmTPJuWfVvrX61Zl6xy2u+ONhZQuJ
DprYFaNHKZil+Xbw4hIF1iCnvjpeixLO6Lhat8dqVHvJJ+MnZE84vHDLOajoAD1PbtTKB+r2Yaat
uqeJnKw7VaGnDLUDpkotHo5mrzCgXcRTLmMnseJ7vD7ukBvxhQjnJ81VAkL8aRlgZ+hur8hHA3bW
K9GfSOmHRsLAstcap6JpYR+v9cHoFTLd+Y3bDyDt8EJMiqG/IsRYaQfbvrLRo69dV4vjTmxuPbVs
k1M+vSBTtngqLQkKfmu/JHto6spgTjOIJW5M/q15X/Dp1CBe9rKisTNjUBQmTZZeT5lbl0+9k0mM
jeZtHD/VaF/ZUYW7c2nN1+x42v817eNpdRlUauPEOOrWEGEemdK/01WTIctbvJZ3PqoQ42r4BfD7
uSkjL+JIgIEenhIGwfuDTNhX5p2biB36jJVjllS7zusgPXcIheweZfR2F2fKL4pWPutKAqpQKFYr
nYSJcTCUeXjswJAzGZzyNgZjPOMx8Qnl4T8nDdjpTHF5r+l1/c7Yf7L8/WZIxBDwE4DlhqZ4t8GC
x60QHymr2ucucbvQhiGa9iTFUJ1mXMoAMxVwqAZ6a+2bcprYcz4bYtiC29zvsNX7vgRJvBsznALT
/R45SqeBWkLPn2gJV3+PNmn06uQIZeKtxZHqX/bA1UvGpMQ6F9lHLR6f4+4qKqtyH3zLdmQ1gnHc
nLDMKqEXRDUIz1DQC0YXtCPh4AlAK8q/E16fR62U1R+jYrqvSRsbfks5J2R8ddTpmYOacJ14KZ/R
IXmQ0J1r9ilrQZcVEFMqUO5GlWW43bX1eVsxV+pL6wSHKYM9DMEdonjgpBleZhAn9sq46sMsWIvY
pc67ekjspOxCkE8i++8UPs4gVy6SeFDFaN1SgZlukeF4CaXRps1jzRQwjN8pyEGj9w9fEzMSwHXj
cOO53IQ5q/ONyZa84tUEWmGt7J6zgbDeFGYyplAt9VuKcOa4XCw/EUlIkxJmzMVBU71LWgHUiach
n0OSPiexf2SU4DwHAbQklNdjLTR6sH/kYdnqXi0Xiu40qyRQ2JZFxWQTKqJ+mpb9zzYM4ZniY8nE
g5G30qbN0vDmOhUf9BN0oK5aEkNDu0KT4lab2DJb9XTwx6rcmUiu99W/RCJgrcR0fVSCaBIK0v5z
K0ZS6eqXLrZl2qaDU7cHSXsSlW1I1TJuLna9nUN2INQfW3+3troLNx7DXVX1KnYpH6jWvEETKYVb
mobV32T2OuQiYNpd5buSVCKneNvgU4uc9QiV+DaWTF1kc/tFPGZ/mQYanVOnS3LsI5F71rxUJxqm
B+3n20/hctenLVSUQeQ4wXwU5M/MtpXFOfz5ShlsOIm3hrfoyhPZXxXhTh89uwYtou2hHcph/5xa
H+Bne3KQR9h8Hqtfb9cOytLD21oT0dopfjSrcnnaFfp83BpGe1YlfEU9ivA+WUjjUITC5gooIRDn
RKFOviGina/osvk3V9eJczSXmW9EYQwfF5BVp3g34jmjAF14nS1w+ZrPLTMA+4jXvM0U5LIgr8rx
jjjCLGqRQt/49k/+qG0pvbeRHxuCJz6wyHIsN1NLGgjhgB2B2eMti29SEU7AKOVixDKP62PzwjBW
+vD6nVFA1hue1TAR1XkT5xsL8Q7bx10evVV4ktT6KitCAkhA9j1xxV4HCfyWDRGPBlRI38sCfVNH
L1v+6zbAyX3WK2gXgocIC22jiDdE8nY+9tuAsYIa/RZ+8jUMEhEHs9uuji/8KkH8PI7TarL3ygrr
snSv5++TEkaJxXWlP1Fuq7yDcRxeRTzFCKf3IkFcOQoR0wWk0EeXG27RrbncpmfcR0TTHGB+cFgY
vAFcTOOYug0q4kWRoppcV4B6YnO4dLzFpB7MBh5bax13FT0dDFXfrqelaBZSYjROtTFe1PggBlbJ
2f/ZG7QOTInhFNKAnqGQ+nSFboeIxUKUAl6kHXvG4HBgu5sojOeHgzjKyQJJrGeeRj0Fg1ekjdWw
IemrU7+uxza/Uiwvb+k4PjPZxvTbe5zBfvDaX2tyG9cxXm4zcPfT3uoyeal6PjPqKf2398uf98ha
JBLvJOFNKmJ5ppwG5lIWPMMgOE2W/fFkd6tD7ELiEm1+fQhPmZsmYatYy2UFp+UOas2PD1WR/na4
AMCow7Iy1V7+Xjg+kVDrJpWRw9tGTqCNrtrclmuPVUtbLS+iI/A+EtF6X2wI1pjg4zn82qZLs+zl
bEVXUkDEaDez35djAHDzhhMM+2lgtEKURVs5nYm6UsdCOc/FyDeqgVwr0nfVz1mhreWVcFYi8lfJ
+gr/41PHFd/aXRzsBsIOXMUvoSOCw92XgxJXXsOJBbMvR3C/V52Lb+rUbP4UezDsKEmTOWZ+tluk
QimY/tPQrb2NAE3zlBmv7QFF8BM3d2XSqsXysDgAHZVhUZ0ZExlB5586f+46u6KETCTGXsN7Cpdv
ZS3zRpcwcHz7bt8rrsfRaW1Ug2BNXhWVmE2aTnN4r4Yqr9+W6kaihGxGsJJxiJu+Oxl+Hw2EjCrZ
Yqo2X/JNjVKIhwfLjDXARXoLquVdwmfLRJBR91cEMCMqfrHnnHK0vIa530eE4v9hYY+2awgQRNu6
VyupDHlZPHxGNSjN12BH5MEa4E+70k8pa/9K4+2Q9JvVFdmxf1nUr4oOmRPbO0na+7hOaqszuSdL
nUq6aC2Q3tWLlrmGZA4+aylOQoGlMF5T1SP38Lynn0B6tNVIdwpnn8NWPdN5UlOXIm70yJ2VjIbv
tK7eCqSXdHciMm3sUqOEYLW/SasUXY9JFU2hpADP220CZTtoDTBnrn/nLTq3drESVzxXpSIl/W1e
PiOwUwUpXmpeKFxi5bvfLR2J2hts4epCWcypA6C0AwyJlfz4DM57DnRExrE5ER5b01IHJ5Uo75d+
3AtJtK/VRNplCHQ6Eun7sNgVcRiWmPIaFzHOXKeoi1prRRdYrH9dZeXno0Khk4Davnl3T/OhbXe6
X8pr1WgBkb3JLuSzByS6MKSc1pH36zAfkh2FljUdXxfhgOfjG09jOVdUqOLE9ZKq6F1LKt8GoUVQ
p9DqZW4gS4ns4rYS8VEpq8STttzxsnbfv5xZVfQ7S6Ul3RuvUzxNzSSpkQ8YqboDt8PiUZSHxlF2
yLqRr5FaVBsT7Zx7jq6ih1hYc1rh2ur0yb0bJlQS8zuEfqdO1TCUjeUUsDr7oQQc28Fb+5j3JPx/
mNUtlxltJcMmge9AbPbevzVnzwq1GSgkMJmuiCW6zAaFoV0/bnElkhsXUEGi/fqNx6AWxkl7Pc6o
ZueLluyo/4g8hniScADniKgjgkGD2Gvfol3u25EeY3UlG2VwnDEFlF/HR7bQkpDN1xXprwV+WGsB
vkf7P3ExjSjfUakBZV56YCZ0Jlw+dWR6+RcKQDKOQ8hs0QH8+EPGbgDp9p8u93A7PNbdugUrjA4z
lhJOgQPQPpglsiAkVLkIwcflpxQly/O1029Zr7m+vL+wdVw9awdzAUEYnM19T+5ik+zJlO4KrvkS
3eIO+HO2koC/M10DibqGbkGWY8tNo3RwmmD767maE5ldZOzFAic4mGWUtCyPpVS+d82wHSuxGkBn
esmTWVgiSGe4kbvJf0B6Hh1Ei8PPYYNXEdCxNRYJ94x9BWm0ni/BRbZJciHeqHCixRur4d9gMJSr
Jr0QqV4WTgG0dWYxQGACBGw8WZ5mooB5oGcOLyhVthkq5OxWGgT2jkyEiBZmjKc28PN93BToBmEY
W2mrFNPS88IXf8+GCLfmXSNArxenQn0MvlfLOjlE0eyjjqNaBtDUGG0ydfWNscnH7F+NIUXo/z9x
fToncdKv9Qjx82WTIuquQP9tMqZfbjDSFrySuUn4kYT5uXPxzCnXQs32aP8yMRNZUe5lbRIVYm4Q
eJaoYeK5ZzIOI4L+l4hMyPL1NytYPaD9QJkj+2o3xgFW/fNXobhCiQg7xlpolz+/OuRIi27+HJZH
glKa4Vf4Ek0ZzicH5Rzzd7fo0XcYi7cInNx0ZYzz7VZTCxHTA9xLUYMr/qLkhaLYbSck6rnLTdVa
Fp3PT++xUkYRPOtWb70qLglnrTzie+7foP7E2UT7GF/cxlaLZ7rSGuXgXmKfImmquZSO3fBmwErb
FepaSknGVrXQig5izY63zfER3QUnTxSS1gcTDiuwcYKgg3C5NXHUTUX+uMIo/c0eU1bmAeuQqIh9
6wcmyqC+GI09f9R0NjqB0izkIxii3az231up4SEwbWLj2QrQ5Z3408GvotVTB4TziXLnjUpwWDan
RXu1g2yRFJ0ffxZHssodNr2x3SXMyhqsacmABJKojzeXzIctdsddDMrjC+aHoDz6sbMie8g6xxPW
ggSHioheBhm1FCdtr1ZiSl6Y13RMUDL0tf4xeCwakE2FjPjeRd6jcPMXU4qA3VnLfbNf5LrOfQvl
t0zTdoBR8wTpN2R87QEvaV7v7LdD+lo6bmaj6tEuimlUYIGj85bnEDUuFhacm2HD4COT9dVAe+ot
6QbmtdUHWfuOaGGER7i4DWKUuYvz4mHIIZ2JfwtV071JpLxkA0o9dBhblMR5h4SIjtGpPULV2tjx
Pnuw5oaDWE4rj8XV8Loz2dFduNrgKw9rblED0jCYKAgifzwx1nRDO3Gbcun220nBHt2sl27wjGW9
globeVp9b5S3tJJspBbblv/cfG4OcB9qGTEM1lUp0aN1zNhlb4D1G2OazbociejZvrol3mkBoxGJ
Iukbb7hI7U8pWFD9RdhOb2cZkrtc3WKBC+7Xl4NpiAaurKwR9ojV+c47vq29y8F999/P4Ffahkbu
rqRj8GoULRI2uvLU7J7e07okfHx3vuJnksAHkgESyK0HcRUN9QSAM/9pIC6SEmJPSsl8oz4yXAgi
jjegWyHk0cqvOAC5b3XkcRh7398qpWVXXwpzDJ8keZGFg5bC94fhxdLzp9mKme60V4jggW+Qs/9g
mhY+IDVHF/XHfP7qjj966ebHJLR+FLChfYR+1FPzBaCd2xvvHA7GkLu9tqFK6w8rBmWbIpLsunRC
+ZPEodOSAVEeMDtWq+1M84hK2i5sv/jGWdaM+PDQS8MqWRK5mWq3thSr/qoI12tjH96Wp4taoT9p
1MH80eMR8a711TziwZkbGvKw9kgEfuBAL5rTObNzNMdWeqNJq5Nj5DdnuUkkS4CNXo1QvbO2ma4W
IjmFglX/NY/pxPu8gjFZ9SFNl24k8N/Ova0CONdVHdYHMQkQjafDmKDEYKp/s9uaWB8eRP+bOiLL
uyoNn6dTTN/Roj8yYLBuI/BqOQJgtcDIRPjzAlSzLXW9TojMdleJMOcoqpbjaFJaF8Z7lliB0pyp
7qaAgLggY19DwrLl3c+GK1Rv7F0usZd4g2Pug7vCSBQEtD+RB5KiRwEUvBWYGGWD4q697evfPe6k
wNs5jUZDq8IIsTsO0/fKv6NlYU8txvPfJX1YTfuv9Nzu1zEZy40ZrCKc075A5xvkf2yOJQ0m3L69
IlzhFXvZeyH3puC02QfgOF+xsRtKyE66+lJyouiiYU7NZ+GIiRVxqiyL2c2vhEJ5IyKLaJFrcls2
v2Vu6L+uduPOYTNtJNsXEFOitMsNYxHRrKGk/VgrsLzPc/dMqU7IJ0axmsXXdJDO/GdgMuuH85bz
5ApS2uCOclRdMOeRFmELH1VxonxTbbICPg0kZO1T8/rpIkPPE9mUmUzFNA8Q8ZRxYW6NeUSPv7Ap
UYd4Bid9hvMK+qwOUG9s8JpTOK4movOOyBP/ReNVjQ+cQv2pLHimJNJ1v4rgZrr2tXpd4YLj3JmT
Fudyz8m4uES8vDBOX3kLQQZHm6/hA5hLKfiVhHqL1tK/+uw4Ds6mhufwtpvoytVUPr6VWA8L8M6L
V9Nc7k0ni0qad2qWQ5XLLzS7yIeP71cYB3AOyHOQ6XlV9OhJ39K2FMZKCes2mtc+rsj6saFZ7cVC
oTUTml8Jd3nyG8wQ9gc8ueHm2PIcvse7a9oXALTU/ZTHty01yuZ3nmZ2bKyJ6cx6YqraPTYqrcQh
G0LOdoLgWTrUJJVszAnLH4pZDOUKRFG6HcltmzOHpTkS+r3L+KQzA4JXJlr6cle272gTR4HRdY6/
FO5hYh/5Yyap2G1HraCH9Zh6/cmn35fAbry1MfbIQlQv5oRDtos9ffWb2lIJkzQaG4FNXhuielem
6aR3I+BR3qslQZBVhmDi4/zcfRtKoB/KFMBQQDHALdHbTeyDY2lYtr8rNPf0bMEvzABhORlyMm54
X9MsdkAmxd1z35PdCUOhvRji28Gg2ZsXssPzsyHCbPzYXVufiwN8Hz64LiHC6Lm05/Bbm/b9XPCN
va5YWUj9VvXG8rPObvk3Ae/6vbs2xDmQhXBmeff5Tb93ThKBL15zgK2yB3uutRqYDcx1bYVnANlO
3RZQchV8glbV22mcWwYKIvMwC8OXXcEQx7SyL0JAMVgh08Ts8OoF2Lb39n4Bo2M4cgr5gCs/iWYe
XcaBesA7WRddpK62YXjPyDn7tkETuzUxJBsOFZyk89QDw32OxDBT84ZPTYCnRva0zH4zWhJyQAbC
X0nCTgkl+H0Or3dIJqXyd4QoVDUsbl5R0ICttHEnGatgNvm8lwln/Dv97UXOoIAsK+zyWASOBtaa
DHKBJktqILLyQh+xOKHwPcy1zVDAMPcrDrmjeZynClyYd5ISzMgK5R2eb1TY9tH/cmpGZb0AhguO
Qx/uFgbcsGGZvxqiV1140YVLHBV9uUBuftBI8ex1El8jZSH+ubIzwsQu9PSgr5fOP+AcyvikX0nw
Ty9oZRsNZtykyLelS5kcQ8gznL/BZjRsr7zGlI317IF9meUG1/bEFFQp5VR2NTmmbsmrQYOzoxH/
DsXDjZr2gSObdNB9vPoeZ8YiJm91+rcP7V71WCAi/jNhOsRuHsvhvtnuuw1Mn3+upV4Hl6Qmc71M
sn8k6nNRBcOYXzBsC1eZdTkZAmSZbEs0E5x/eCk88P+/+WUx4g+aQWN48HEYpoFThVA0lY3W1I/A
/abYtLwYmBl7d8ECwXK/LLfSd/vTgtjHtiq0d+7cvJQXj4iqjY0AhDdXvg0fP1ogDVGSu9xE59ea
azs4fM33RZr5NY9uEXUdLK5L/TOD2vi79W9gJu6sYB+x0+IGp3qqPZdNQMXs+DZM8p0XpyexxaGe
DCuS55wCcUeaOlsDsq7waEEL4q2FGKU66Jv5e8nPAiWjZqJ+NpF5HttFpZQADMDUeg1sNuEbDWBe
RNclXal0WO12ixWG4FsdI6qUQSjB/bOyRKM5Blz3SsAKWEmL18eBEi7Nxl/u/ROn7MhTcYG5uolD
tyAJOSfQR0PzXB/ht588e7KJsE6pRbqPOywqGu1MeYwaG/eHkrq/JiEiBi5O1pcCyNVCbw9bJFbL
BYSsQUPvI5L7V7EJ6mJUGI5yuf+oYnryr7JT6Kgfm81fHvGHQsjOVI+VenkHwCqqS/ZToA2t9Nhr
PFMRVyhig4TqDaL8/BYiKlqCj27f+MUQZ2H30EHN5R12e8EqVw33K10r103RspFbB1ADspprC78S
1piXIfTss7hQdn7LQ1ashIXIGJKy/f9PLqKaTraNX92Ojh2w47A2wSKkpxv166lgeDmkAUTuCtBD
ofBCYMQK61FAC6M+IcyPCNBztT1AUCCxtyxZduTlvHv/4X+fK83Z35faPNPflNKFwM93WBmoHL3J
GcC677sDZCLsCqLCHr1P3/xahi8NMibKKceMoPuP1eJ9tVgcCragDDl4ifgnSnw6AAnfBZlujrJG
b66yFimz9t0PS4HCnPoMMBSKnWirel9AD4DC+fkUis8sEcldLM6sivRbatYpZk4+L5OwZdzFjuXx
3ED8uz/WlhOefwRRfsIwitwMbLVVt16T6HBLp4ZhAPtkK+ghYewrD+XwEvYk902cAUx6TthtYNpu
U6W+7QhAILQiAc1AGklK1kAK43dP2LZiPkorRm0yhO2jLStUiVY4LMi403VdDFmsbkFgbj4CnKxI
uJvZYxTjlez80Ga/xWCLCzDcR+XrUzREQRB5wUqZ5S/sJ1zgMc1TvIulDyal+A5xCrAkEGJ/DXvq
u6q0eAqG54eZBYMLoZvaXoseUmlRjIrEG2m7AVrGWgJl0wYte2zcwelnLkTNNKW3Aq0EHF2j1wEQ
5SrrV/jSUrEU3VU73OX65MXxEE901nvaKSmHTp2Mo2ccurHhP+56EyL5CL5KEXb45YegIkMXtqHu
tNs1JqNl1pZM0O9170CErC8LsOJrEEaMJzSL1onpplREKAmuKp4WCsfmNmv6SQ6d/srqDVtDqXkP
J6DCYllt7OSEKnr8xmmp2pODqUge6TNiSCZnbhfav+t7zv41QO8jXd3gScRAUz8U85yho8UY0Mdq
5U+K0diyB8SvgwwfA3BLx6Pi49LzJfO0kn9s9Io/MR5Ew4YmbZLuJZbKV3/dfavQEErt92CS+/3F
/SLyHUDInEgHu7hALaxHh0lohDKA/5Dr2YRHokAkZFvd7gWEDGf4Va4AJuR14fS3p9YydkHvlOpC
CTOuFwcx4gbJrC7UR/hlXEZrf1zkNkg/z5A9kX331sgo8F3dylwVklUZ3eHPz0r01XMr9s+SDmke
G8k+p+5IV48/Z0In6GHOKHNwF4Lq9arqjgBT7gNrFrBglZ6XNICOL4ZeN3kehNtFkht/5RxvVxMK
QBrTlevHEH2ScPi/dt7WzT9yspJXjJOIkzCvAY0t/lgx08xFHskWh/e36e4pQMHCcbS2Oz6Cmyvf
THMVX7yfvjimv3xQ1+YUzrubLJNcnSnKZ2tdSoBjwZIo+GjwDxw4A0Kl+cIBCbPcENW2KTa9TLOu
zkvs48ca84HlxVvVQ1vPGKuqg/c57ePrhgcDu7uOQJe6mMCzBoQHH+zVpwZOztuh2QrYdLaxOF6Q
O9YKcd7lZJGLIXW04DFW5xU9y3OREWmxwdkKpeQbioEUV201/7AJv7hDNvTRxcXIZG+l/8QgtoiB
hfxusGJB8Dm4FmuARj+ADM1IlC2d/k5HFVmW5w4YZ1B5WcMRmP2cVnBVq5bZ++F8AsUT0uDVAgxr
gu0lII0dlTkzO3KB6wBXNdF+Iy1qJIEquXomNEvsn7nmDx++CGXfwofmuh5chmxmI9U3qL6kNcV4
FmouQrKYfGHgzPAWe5F9U73L/uIuz0gVKH/A2RIOo2nIgSA1/vA0/lF/M2jTnI9A5enXKDEfKNpx
r6yZBnkxQy7qodlTc8CCY9RNZvmOTP+lKgBIDQOAFULvb9+fuzQx5n8UdaBdUSomIMjt1vj4XabD
kWvDMlezJraCdNppG41NfpaDU1T8lNqH31nWwDVsD7kPe8e6brv1S4DZWLgadC6AnDfrXdRczFGT
6TAPCNY4L/wq6GceHVu/CcAGhNWQHE5qUF8RdJjs0OL1HLKc7UZzxp1H+CqA32lN12UyveAkoo1s
EPiMDemmfInSc8NTe7lDIbeI4AvCfXy6HtvLORyaE8LpoGwoNKSz8ZMUv6eSCPcV/dMHPkGTQopu
dBs5Si29Xv1a66tdME2tKqh9uLyW6wIk3/ZEQLPJgdzJyXvf16zc6R078A7Wp/AkF9fAeEadPMl4
xR5Mg94dySJjfNCoHnZYjCfHHKskPwN3wDqZB4gA10zdwCoxCanSOmZAFucGMVuBvZymPC34T0Pd
VSGlkwJDOoLm3r1vehrzDuSQfE8pNo5wx/5CKBNbkhny3psUhfbxP6QRGSvhtOILakFMiUmSy97Y
gRf2TvZbVFJAR9SwlImn8evdxEyfrXjonJ5PiAjA56MBe4W9YsIMd1xXB6dfM5Z4k5gl+Gsqxqhf
cO24ss2Q4SBj+9DiiUPzpfwb/2tDZ4nvYEDGtFkZZ5L2aFHKOu/2uEr6y6Q49D7IfHvmF54J99Yq
Vhthu51+oWUYbxTHZxHycejCwfqMPPJ9ptsGyQO9/JcjxaGG9CNHKqcbStaDoo1yz5ndNyw02WTg
huyobhde4AysMEicwhYPed8rbYKZXqfUZhhRA0wvufFCOaCtFK8MI+wrnsFtdWDDybFO5g8uDbv6
dlIXcBD7ZT6lw95d+ENW3nedA0VhTN0x4Q+VrVg15tGWKirsGwTla1JtS4PDG/dEhuTtAvnuD/da
vsYhMq4alCY5jmt3hRYucPeSqj6yT4RSMYmRoaWMyeQVRzAUY52kY5TJ6ZkJCzOc8w0kTCq30wbA
FIob8aQWBZri+u69+UxjRpDVT4Z6XdUK2ZXm3mInozDvBbmEmntpb5XbAM0BLjsInWR5fMPBRCY1
It4Xk2pS07VvYdOWpl7vCB4x1YynwjCWUCMN2m8dqGGjF84OAgInNfyp/hIkHISehXh6ltsEia0r
7FdrlBa9Dpcj5u2A12N9kKY260S1FXJJeQIX5eJZ6dK3BQCfvzgT0yGi5sQtKNOx4x6Hd4ypYejl
kX774Qs6D7Ja3iLpt+A6N27yEHZEp+YWmHbJSow+NVsRRmTvrbdhldxoF3poR/bbD5JsJPNdkm/R
fvt42ESXzmnhdftPY98lzs9H4t6Ge/04aOXI25B7hwvMlqy64FBthlguD9oWYiXOa6ejBXNO7/iC
9xAbrRYt9DFlEsSaXpRxuzmxLXsJfkfqTKOi1m76+Bi55lvDAjD1ScbBWHu9vB4W9vPWd9IuoC8I
K6zJjqXNXA93YgLhtkJ/NRiiYdosA/bF75fGJygQoVB7g29nRWwz3p+pV0VxosN8TIf2bC+azaNa
kQcK1KUY38EPG9kpdtMPqxaPkjA96qgAd8bGxboSyhptBSr9lfAmmwWw4dEunk23QU0SoAt375kv
F8najdvrDrWXNH+tBakD9HeQwja1E7RVa27tqQDOKwTIActVahikp4CtXYbDXLiy0jHh/rIDpSlb
unaSOFczCKuCVrm9ln0QuE78RI5i+onZjN68bQaceQTztKoqGcxBJ9M8xK70QiUzavcMKzsAbxsJ
MPwDP4+4xhIGObaE1Uwy5g37VArruQkTNdf+Vo5u0zDmtQ+q/zlcjsjIqz+G04ra4t7XiROAcuj+
ZsWzcqGyUGcnU2dAYiSQ4EfuA0l3q2efzLSfedg8AAq1JuAuyYYDbpWgDzxBLzsVxOkclz0AJfe+
O5T8taOlUk49eMPIpJPr1NZuMqckc50ourB75BCMBgAZY77Es6stFG6QksWCaO6Dyo6yIo+JR2Ti
5zgm3KK76parRubtVucbLC5IX725JApJFw8n9c5H9aowSuywvRrwf4258nhdwXPpPBQtP9NuvAlJ
/ZL7h7EMXy19gWjGxG68imAyyLb/54/6OSLe+YWG+QvXxhuaIT3cLON5aXO56G14vkNb7UkOpp+y
IoCk2vAOkvhkuy4zIEL715KzH+MqSkdJ5HMkZVLjDh0rLKOqwEFTpKfOjUouJ9olYvElsHBCQMZ0
Ydulf29Kx2lck5a21FACMygzQR4BNBpiPU+22OtmiBqfKXBGYTKM8+8SA3YSESfeRl+tjx4Ff7EO
L6Q2mCbfByensrlEG0N6TCK11qf4TUvQAMlaSSnRVT6aCT13ZE+xOq/ha6UKWAGdxgER3j0y0Dir
7b/6Aw99VOjGwl6NzQ+t+SKIvCZPXSVg52deEdCtehKxmZNmLd+0x3hYjyyUR80/s7FZSs6Xh8C1
jnMMvuICT0IAt486pbOEan9EoZ3L0V4pxpujor3fawnewqNu03oyg9CMADhg6SXpRiczmzocB4jT
8V8ZbyrHE8POED64oiWOKI6d44wto8426TsHrFRMYTs4fP2LR1/NYBhSybb4P4h2z4lpwPl9+OWb
8FuGHPH0dVKZ9OKH98lnL1E/S28afEwFA5iIK4pP7QNxkoBr51cyNiIxMzkodPYfICm106B77S8E
chyfKboJOmgkY0JdrLHy/n3VNwgiCWXJjh/wzj4VpsP6tzzyXmR7Cb4A3WZGY1oaR6FOFOxmPQ1k
FwF5iLPdTaf7WHu9gHGN9p5HE8CCJHEu1NfLJlSYW5py+Vr0V0AdVKQwVKwqaXm7tAxaq8fVnur9
M0doEUEoBp0PsMneT4l32aJ2hKzmCa6RNspv2OkhhDcX65u2wUWeGPmm98CEgp3uNHiCBctTgvPc
UbTXq3VuEqrHCtu6VCmC202SmwAXxGbmSgVgRcAG5FGxk06ZI4KXMjaVPo2fkrUFUZzXL39tW9sV
h2hI2IJsO2QYOkaIk8aFRryrEGblBSBn9Oyx+HHC1rjSX+SQrxVhLVy+i4YP3nbL9rCPle29UE8G
RqxUdb2aHp2P3V1pRmLH/akkeF5OYzqUVFl7dUe49GYLBzdJwzKFgnMhtgA1uBjSurzTvQguAXYP
kIs8XUKpkliTlvv9wBsZ6KIOCeUZTUwDHaF309SIXyqUqTOGqKRYzs0RFyhh4TTL6HdWUEavR0xC
Dvgz0sOLAD5BsFPxSfRnoiBoY/nuU3tdDuvANLn5PlWY4YfCWLdy0DYL0TYLaVsVGq5OKC+tg4V4
XITQE8UcqIFnFdt/NGmWL/Uxy/8rMFCQdb5shbIu2Wyw7NFsxtBlX9i0sKRE3AGJwaR3NCyAo26d
QArvqt7fE6Z+o+tLbMBJdmmJT669tA+KFhhYDtzndGla3E3udoQeiFunOrvFCVoyN3uZtvXcbphM
IOnpUv3hCxFlG1tHzNsnyTnM3Mnp2uH4aLe06mhD4wNyg2ZEjRVCTJ7/Orz9JgCp7/ed0U3Yd6Tz
0EA4TrlAsHhhFoilOwrj4+1je26bR73iqRh4D/QcfaVn6oiXn8rBnIAk+rQC5y4B200J0cPRtEkN
aFzQZRkg4H8qBldYjotvjn0Ya6h53zG52+qfaEMXigvH90aOkA7041G8ZBmkPsTgyn8qRySQek/n
kWsjsB9Lrsb7HGZV09OTKXbieHtYmPcTPa5hLwM2Qow2743dlWSdopjxyKJ9m/66zCDQYUM5qz/4
++Z1FLOH8QEoC5M0UKZI65KGK1M89c6q5gzU45oCfC/z8e3s6aPjLzDemTaxe4I4QAGudw9WKBuJ
GGk4MrLAFABs5XbqRieHk8AnTJlFmUqvVKg4sTzcukopVS3ss4zJCULKucJfvi4rAmBjWbybq8Df
UZAivOSxLExTp5H7S7XAyXoTiykL48vRH7oSn/Ohoi5qp+hHTW5P3tUTQlZvIs8EhNVv2rm5bd5C
cVivoFT927pHDRa3FJUgn1UcKajqGxSUUzZxQDgoaeEM53YcCYw9r3ivpUozSZy08MfiK5oWMy9q
xQvqEQd4aq1p+wxx9i0Non5x4LaDRNqIscSZXTuhNRKwUjfQMT95gUp8jHXGmoWMRC53cRan3WNP
gNGtbIz340CPbN/fkGgH7R+81gqvbdF866EQCgW/aX5rHYiY2KzekODrqiyjhj2jBkRIKE6oGTKQ
q+501/xZf0abl74/9M/YdAh+YcqY5ezzZTJT6iYxi3DlOsS0IHMENJXRmB7hiyjfVv24oww2414f
7r9euz9VygkBcMvTXXEwlYvQFZfEX7iHZc3FE5LHiUEt/UluIj0q2cV5GI0MSCTQVxrd9pfbm1Lb
1ZfAlFWZk4dCLTssRipDtCjebVy/hEaNYZ0/RVSh+j2iZDHfDTmPUbg9V+Y17IFLhTqdMySf6pgK
hCJ8kWjuyi0GD34IMhKvnQkPb3MSmHkQHGrPjmlAcMOAPykMQsG2JWH/cG7MgVHOl/NhQ3D9/juC
jE6kGYQHYAkDokKUsZ/4TPWqVu6zO+pG6c/8AVOf7hev/X7CyRipYH4K4XnT5XY4SLTBehn/glzZ
V6uSAVFcTwomrkbbZIeeOk7lCbqUgaqj5t7cN1j5f8tSsRBLbYWiQ4v/SnbjH5PxMwML3RBeRRfq
jJ3QtDefdJMaCppnLLjTK9x3re/2lA3Gq2x7lgii++n642Zw+vbGY+/B3i/SVVvSp4ORkEv5PPiz
uNmasDAsSiUHExwS09nzBU961u5LZNtUXyj7dayqsLmVrznGWwghFYwvCgNrxtOfoGqdphbE+07Z
i2POr5gf1fLJEtdnBSiUTwiTcpiVzCmx5HtEMRzW7Dkqa6Ag7NsfbgHw7VWzggtK5J08PyFZI7kb
Hovw6TsAkC5/NdALJmGycV0IM7uHKFMONAfAmZ/zxQ4/n27rMEH3r0OdtFpbOAJyeQ39zkyQ9upF
VjpF9vNImoMjTLTRERUjVFlhGA5GSiXaoT/LH6xaeQjF8VWDZJpa9PqMgurM48AlPMaTcN686F9i
riOkfd0yQA712TLxS/jDpHwLnVA6dbX5xTjhvKk3o5cOL5oVDaKc/lknSBTQVQB5lyO7C17biJLQ
u1A7RJ7t70n5FUSwHRvCM8Q5aMWAYab/q64SHtSn99Erk3QQTNgm5xuMsWPV/TSMbEG4TiIQ0QF/
oYp0mUhFFmN54BSOuWcjC73zdcj/p95GSITZYvOQy+GwavdOLyCJA8dh0QYY4iuS+cBRZA1DWhNh
sSw84/DD8GV+aSfJyoUy/5UinNCOfiRa8h4xFTPVRAH8LgqTdfBgAbDIu3reyhGyty9I8SLpeMTu
PTUwmcf+Ojfjtv7qIT6GERpWGv96Ek4M8mZehi/9AFY9APtNXx9Nz7YiuEMSJ5nDpfDkJ3BLZI0Q
ohPQWwW7He4W3SsZaGqhGq5h7BsiF7aAR9xC5/PZaKGPmxBn4B5pjPTsbfvT787oSMUtNsBn7Opw
yDvvxm6R06kQwuyzNCMX9vvOupeA7OdMfSZl+f1oHyoPg9s1A19PMiu9plODiBVM+bAj5UC13tje
3ZP6XQOwCzzKCf0F+Wp4jIy2WquScbLfSkhjW2MrVMeohuZ9ZRN/q3Y7paL66KifJw0j5Owy+A/B
eshYqOwIl7/6H5ZoWNEk7kyj/rgkotD6fJwiBfetGRk3WiXMyjOBiMIGRzA2w3ZsoJuVe7NDWwAK
mod6UxXIVNxGxN19nzJCGEBljQJ4bwYlkEBqMEKSjE9Om4II/vQXy268JqHyBPBfHvZBAVvtvARL
8xGLlnVTrqLBmn9XLI1qkQDLe/fzQGQRBXVRd22VyeO6Jxu1WT7spUY4D+uYaZR3zx6FTz0dBEMt
gr86sLMORoWEboPC0nSR6U6zlVzy56+CsfAWdlexnKW+o/Po46HNWb694p6EDeWaIJbLVMaPS1E8
V4lUXdyZ9PUuhHry7/vhtUXZrqWo9tFwnl1vC3gFcMnOmf4bhACv7HcvUmxIjvggurZThTtvxX7n
XI6he8iqidisp1pDPswYz/mQgC+lgnZANUdO2MY1iK8sNPSCZucDLOYOSXk3Y+zKcyTwSPdiuNKP
VFaO3ZUBniEYLT47Mdb+OZBUgA3pwqukFyKP/wQb2KXFrPI40xT9clmuZfkAlPOUocjVMXbLt5Ri
BRW2YebhP5kJa8J8qonrDVDMmONzE6l6ezAR0RXcpV4JBDtZnPVLofkrXQkJ+xVNxSy5GdjB82Cr
LRGdHJ9dLLKLNcKZSwZ3PDlNhPgdsTmyB+Rq3j5WMtCUusjICf1vZx4TFWpQq5dFTcs6PbZd/2BR
0QgKYJpNofJOEzQlazwLL4YINtTm41K4v8t0bwm6WfoHWJsgqVbYAmlV5x9BT2XXxl282H7NJ86S
KXlYK6X2eNZLhw9fXplqSc2lJnDz5K++t/kR/nU7U3w2DJkKIyWNrYAaw4MtYytvgJVIXZCARMbR
SPsk+bXFYAo6wUj3KvEuebrmVldhSh6dfYz7gCVVp/JUewmG0LftGtXyYaIiQl9RoUXNn4/pB5k4
9OlVr0dXDxr+czgc/9PV36vnrU/3Z6Wq+eYcEN6iLwZM1RTLqNFC/4GAwTBWkNTdIma7umvgW+Ng
7rWjCkhpxgBkChvyQ9aJDel/2yZAi1ME7hKbbyjQTpJKQRepFOysY36y7d82zEL/u5uqYHeKDW9L
svvXZmUKvxl499pdG0Qp4qQqdJBDWlemAIeU5og+xvPySarnfbcAn4VfSVrdBXRBOW7ySnQyAT+M
0ONB8HY1HwiAGrYExh13NbruyivZ5aMA1+PgWYcHulKdHqkjE7DmhgZHrgxr6B+45JqWfF+60Ijf
mrXW2aMMAMOjmP/lxbL8k4i1/DERBzkXTW1gipavB1XG/dNjqb5a4pg2pKXJuTO/T4oYD6cunAmt
CW9E4q6Z98oBvq4/WXzvjzaaIII7w0zGukHbrhSKxbYn3UukuHERBTcokRVKHJ36+FocDfoJZB6Q
YeEEY8qmEXzDPq+T+HlN24xmTFJeKtqZexkI2RgQPCtWuRWgBjcuo52SQS07PY2hBJTCYsr7iwJ8
q5kj4DoFPeRTe2Fm35RXHdCj084OZ5dRf1Fyp8luI+XStD0e7yvunN6l3ExmxjGwyoU9Sr4OE2MA
xprmN51nbqFbR/wHzZ5uk2xM0E7YpH/mLw3zzVzW23WyHoaWQgvzDa9uVAZazN4mO3xvUcwM8+aq
FDSBvTJ9b14gzDxz79DyOWfonEDDGSDGVcVeCSLPCqNN+nq3OpENvOf4xo8Y/IsxZqQWPRIc1+b0
Fygo/zHf8hV54h+3NwjsgMuUaUFCSdCS0U9i34H5ln6ft+C0aYUdWFyp0daBSN7eqxGLdvLvxo8k
DKiwfrhshuWL7x4eKuHIa5H1Ckgy26Iw3YV67/2TP0q84R8/TFHR1pM7aoogE1ndWuyNGwpngXxv
+q9r74qo3vytU5kpiMzOiFm9EWW7QzB82batpnl1NtEFNScMC8RBcuaKbXidbBbpXdodQpiTl7tZ
YoIsfge1w8bSK7e35bjEbp6GuhTO4Zn+jflBVFx9tzrCnQ2Si9wD82DvjGGQTSFRT5HDuZJbpz+v
4avl43/9E3QsSsxMcoinnFLR/WYP4qjz5V25D8rQMJ3foRyXD45lhZYaAy792ZBLbsorK+bye8lu
ltRRhyCCmQJ3TPdmuVicxtYavhy+yq7t954Q4JGy/rEDoyE/5k82hLGWHrwnBtoYGAwB22RnxVIP
LlPqr8tAlauhsWfMwneHHmq7+m5lRNXFQKuAgQqaAEN+I7pNDQzI1mRKO0GISKdcJP9NVrs/spwP
H+YPnSqjMoMwV9wlTkFFRW+QKMyIFbPnALkcU2QxjrtCiqpPyp4pux1EYIdKTqjihDQFIFOAEqYa
WnJcsZs/VpTL+hOj78gqhNFswnPtZouZMnl4vIIi/pH/SuBlmWPOv4Hl1O0VyKlbDwurpLViA3V5
zggcCMuW5V3pBIjYSTO++lboh3eXxr0LRBGJQbQooF4cSqoNjC/pHpM/c1GyyGotdoCiL0au/1nA
85VJY4r/n/8YFPFgMJhIJw9KbmRIWRiD02wfw+eW8G4+b6bMjU8SbgvJMAs0iUwFz4FsTs6LTcQt
gyWdPDyAYfBCcHnQYmln//wo3umjwlhM9nB+uyMmUkIn9/DyWn26TDp3ZZS1y3zdfsj2Z2d/qbKk
nKxb9CKphf1Iar+4gd09se6NTRBP8C+ybvA41JyyqDdlv58cBQdY3P7TFm1T15dA9b3XPBs/n0dZ
o0zJyjrwvN2nHsnBJrl+XNKGTTNBDs56Sa3fwtpkzx3Bgx0BZ7kysr1CtSc8NTcQFPY2RRP504Zn
N5sz43GCXk1rK7xg6TLCfP0o3ykHtXnhvhZJyd+UP1FtSbq0NWL1y8NFnB/H+d06RArcolgV/zO9
DAkPTKZm/prz2QWYl72Q/06NWHZ3Hn2qEGrIbL3gvO7IU8Mc3D6vWpyisnwRHPewGq9gjdlrIn3k
ySlBubvj2ao4bbci2dneT/BqrvynvOGlfBS+zMb9j+LmhHEvOIeMc+eegSWIbA5s8QwODpNv9/e/
f2FrAjZEjN1tT53tZcMqV4887KUV2+BWlnlwjpm2EbPd6mZfU/G0OWDzja94leoO4LiGd7ODQrR+
TOfIPZgX9S8V/8w3HRjUIZwUBaLTUvCiDDH0VAflvBr5BPJK874XWZ3UwuBr4vvZdqidtbFE5Dct
5SSmOfNYJ8WFM7YnZve9JifDWyUB8h5xilU/6YE/7Qac8P25BXz/hU1WUzM6X4nFnS915x0E8C/V
YLnqjhD7ara5jpEIqe9sDwxlAURlALmlUT6EM03nWpGofWuO/x2i2R6hNUzD3MBfDHr4EE3t0lY4
ssVRvUdXyYIILt5mBw9f5xnoJXojCRX4JlSnmZIQ06TX29RUKRz2GbmqK3BdEzOde2uzMYZwbuCN
42zhlLVZ1TCwuHfCIUz4WwgB9E1MGx2hdeZirszEH6PhAZk0D7RlwLGtRu4NCeIbfBDsPJdVBEx3
weNjEvaMqqCJ0p1EeurOPLmxnpgE0+CvWfsXgD8GQC/hCTfeWZ+Ap59KlNZZlLQlQCZZt5sjcepi
tMM/Vq9NiVv5q65VssrvoFSrMxgTlP3j1KuLVCJcBbaCrFuYCRDUuuHOmbKJfCglijysGKI/O+qn
Ap+ysuqSyzE998wNo9WKXFikuTRexiI3gTp3GWV/rWuD+BMmAOGteCTsz3lxMF5GNgl3hTodgWky
zwCrjJA4tqrD3+jBE9xCe55nS7/ClyH52kuyPmpcrU8LHHkTlV9kI0+5fL2g7qnrqrAn5SZ6vDcv
w6GHu35Db7KG0cnyKdh4l+oJPbw+BenW1ZiCQFY7ZmQPXIGKvyrl0sV5lmTavmrZqJMknG0tIKwv
9C8kz8A6yPUhO05LGkBE0/YXv/0M7s4ornHBpalj7mrCunxkUQ9DAl4TILbUGUSuY/qwxUoqOo0I
TULyhlZdmvUv/yRiBnVT0Yl9XasWmfwWxGIUoqP6/Kg4ApUCrzkuRwzHpuGY10zBSAdmLZOzVT8D
UHuKycvVI5FxkzzlISl43nY67FKzCfLnPk/q6cXilq/rXJPwo6u7iouPvVLb6z24aPWpkuzJp+wk
9pPpv+HFNZxbWcNjQ/DFmmrOtO1KCsucfORDXB+3WIJC9iGtoMmtkChBI2ypIZx5GuZMwm9PeeA2
IA6mKLOoipXhXAOGNquAO5aR6K94txfaOkSoor4c56b97i8rlkia9WHPG9nYLdC2KQa/yU8XqpqS
1IHs/hF6ffS6lv0/VLgGyVNoqA/4JJTTHJgHEpcou1de5JWujUjOMS9gNFXuhglzuPHPqL1KiDnw
IWmiL5W+prhx9wAvI6rCA/6qTHwbU0zCgyiSOyQNaGDMolFadWM0tARPRmkirqwWkQO521jR2Zsz
hTohOnclGSDyqGgVm/Aorl0J8bkfgDcyLtY4ggawgGXvdkvX2/hmuDBMF2qRKSluDh7KtQd3X0Wo
yeQTiXyZW/tW4y/QAeb3icXH/CLIvTtRa5E4QyamwCU3I4vV2Gx7ieMNBR4Ywha7ce1lG1SXcnCC
+l1LcvWX+W50R3cGuAuIOLYPQQ1/hnuuAQCXBzrZDhmOTfrXPbNc/fEFWiVINSdKE6TGDKglGShk
pVyzuBnuARUiz+xF59zlrrmHPVsXz4Tt/2byLHjR/PxrculIyr794YAQQfQhhcymVP8Y6jT+PaFb
6gbABzAlSjncGSnclsgKdB2bAAofeyoQB2gpS4vqF4sQbfrL3OioJvd0Fl8LOFnD7Ck3aMk1WFGD
PdGN59aNXR7g+LrzjRNMEvLOof3i1Q+pSubycgL74t9e9f/n/WOxj9VEQs7KXNGAsl+bqHXy9NlZ
i1QovsaDpCZAw2RHh6FaOn7tljkSngfUuwMtWzEVdiVxTgimS2jsDxR8k3HtdvPvUzsXfxeVREQD
2KvLIedWXvvtVW/BtQBerJY5Vg+7iF8jv/TxbivSMbWDv74fSjNQ628walFEOyPw94HT1tb8Eo8N
V/IXbrcANisQSvQBdtZu5zUwOmapiVVyh8iEcgIEGVQurV+ldEvWoholmyWOT0jZNdxmExBn0mz8
4VAbWvT6VDKgLqfAAcREpfQsCPLKmRshdcZD8RULtgydN59uDteYTu8v1uJnvA1Lhx5/Sl3j/BLz
U79K89peqGQw+xZWBGZyMMyr9KHBTivwLCvvGMyWoyMIf6AbiEtKbv/1QMu6iGD4jka5yyL7DViq
9XnIwKnGJA4M9kJERRH03Y1vAJDwVDe3tl7sNtJyfhTCPDUXLBZJusFq88kWVY9yXSgHbssvlfg0
HhGrDxFkuH9tcJru1ot+Cc/MykAaUOiudWaF5b2w4x6cAGNuKfHUkHjteD90gTAuAK5GgIe2JZ0T
AKb8CmjLS3DqX3fB9nORa6guBM/Uxgx8/RmS7D3mR/UrsgNAJQz03cZA4mczkgUEYSvtCJbgKHnv
s31/rax+Z8lCFXMoQC2onyyqFW8peSasUa/ze1Ftug6qB2/edhxn1aodLYJAvckoF/GhWZv5TrfF
C4W2H86SeIgm9vwzfwEeDXLdGPa5pfJXSmJ4KK/4fSFAJe/v8sXwNmiBmZZJvj0QQ8OQVNBU1Ump
BgMYs/In2kueAKF2uJhucA7DB33IzRftPZC0JWWC68w3jtAtgwn0u64gdVQTBx/ZcJ6xqcj/I1t5
LEEq9D8rBwJzvVFk0471+xlttnXmXHhXDwzKkWeStEQjWXXz/uzt3jeBPZd5K5afJvuoV/YMXozv
9L+Yz5843rBwGIEFxZi4kCca9faDqgErP9JJd8jlDVpcIJ9GJvpA2zn8Fjx9cr7EyQ1sK3H7WZOF
4rLF5Aky6pnqmFr0rfnI2O1FD2TPCwWDXI0hOEOaVdQBKGPHdPHlZ+blNlC+DcrYTfQjg6LALGzi
qnPMxDyLa2RDk7f7W2M14LAGkMNIGHyhP7Lq1rR0G3Hndyyl8EP1C8OzvWaEG2c8eLnRQLxoN+kP
Gp4w7wjCxaGEhhiOner8CH5ZCMqlqn2GIpXgd55xtfBG3rujYNxOBIxT3gMWC1zvI02kKvI8MP05
wrZlvKVnPWRBsKjilo2/vw1MkQnvS056EHbjG3ykxVXjlz4FtxXdziOAZWGmkcWL1SPlHboiIqi9
YZ0gVPrW3tjGK3hTm+a4Adzpo9M1R42yCen8AUcr1ETRFqBXOHQRHUUTuMEWY0EXqSyb5jRKEvt3
y9s5PL6fCmsA7D49uNJqOR5COnFnBUiknrHwrk1NIEQa65GBngIqsUTsm9osoxJa+SSHptHG1rdd
YVL24ouPjOk4fjZHdb8xqizfBY9ToKyc/PTfBs97zhBPnWkwY7ZdgtIk38XQBPgEi6umpRY3wijg
yQSjSKeHBVWCyRQt50BMBsXbh/GUxQGanF0EgrF7sma0G+6k9VJGPQ9LX+RhS4zecb6jMwKXlwU+
UG4NcOHFmuenhizKvJhVp+ALcY4Dt7LbCynABfG6jUXIJZjspk2mrt2PSApBVn5d00OGITrf+yjs
92/L/X/PtFpZ2nX06z0ddq669uTuJ041x41zmKr/C33wxPqhZZ0/cSAHvBWa0+ITbMrRrPG4lAbB
luLQtuRXtU2D0ZUiGFILkVTaFxdddVTr6taaM5ckwliFUvm7SsqIXpZg2AN/lg0ISRSz4oe1m0fG
AXWkuCE1dwcjhnIcxjFHUGa+IvLCnFSLk3Ud84eVJy2T2etl4z6qLVro2Nw9YZzWn67j4IxH4whn
gEpGgYDL/5Ftg/NjkpnJxGsPhpQ1lf1tKNF37r4r/O5RiCOGkl/9TEHNi2jFpP3ajnj9oqy/ZZ6o
vTWaAQFJkMAabKv8w+vXsSBY/9bRJQGlhDOosyYgr82T27v1NxNop2pfK/tYP1pZ1zO5zU/I7fyA
r6yzsJB29wPYMI+WL8NUoAWE6CooTai74Gz5umDJJUXLjFUUWyurp0kMc2WtCTmu/7IYYfdI1a1j
kOIX+EtnPWiZm8usIcP0Tv8V8Bf5gSnflcTY11JVJ8CbJg6rGR6bbCn471WD+4sqQvTPZnwsvzMf
cBvHxKHmcuEXxojSQ/r243G6LtbnPAk24uMhAzzySomlJ1d4wQCwoS/YdO4LGm37T/72K1hbvD8P
ne+ITU4IjSYTUAGFkvr0crWjsq/Kal2sGcylq8Kx/XGMc5lNXuTztvJdlgcoUZryIoJSG7v9OzeS
83YxlDqxq1AaxTo4E9XFTNM4VvOIHV84P5ZqPQx2uUhycUa15+uZxQkms8kMqA2xYwOPUH5LS+9X
fGLFyMg7Xyj83Adi9apKpqL5+UjOrNluYFak5u9oVMzI9DHOYXMQ6SfsUjTpszxKz/pxRMys+mJj
G61lo9Vc5TMn/2bgJ+IWRpCdvuhLMxOLly9vtgqfg+rOoqqHH2SiFP5axJSqcMHqemOORMgGDv4l
k5LAnI8FSuCKO0XJy1AWoHynvrOerMCa98bdswFXskoEZqOC6ZOpDkTSt74PY5IdGsHCggyXNRiD
5VsMibrTkODiLABvAd9qEXQ70oBbBcs+Bj5ZMGT40HZrOVxer0D7Uo8Adt/FwqfYt0bortuPkZjX
ur3CgJb4TwD/razRJSHmgTav5maTP0mWha8fXCyEuRkWjW1vjimDvIlqiwdTS0HRurzAqHYcq9lu
2SOImTCFImsrLyA0DGx+jpevPzoOiRNoA+DCWMYBahEXUvC8xbaFGtqoKgNIPXp1no/gJ+nzVLWu
I9bF2GxSklRfG7vusYB2k106WH73YVIbAOwEGl+ypBxK+8WVtt5sruVY3eUhoF1GNmtbZQQDm47t
eQCwv0Bssa9xfKLHdr5/qrveKGTaLiD/S7it24gTEoj54r73tmlk+hGV3eJ4+R7KeFEmI2UEsxnl
KH8O4T+3IEId3jypPigAGS+BUJOO+ktGOFANZmYXXntyCYnesBnZvh1A/olvVT1p7NvjlT+JtFrP
N/IPY39pZJIy349/LEUnNhIvitoI3FD/AlKvM+o3Y3vrppWy7ak8Zaas0MAqNg/qqiarCsItUFP0
4z6duMlroI6MRrb86wJX3VqHt2oebvtDDPeCVBfW+o6dK0RX+2BJJN0X78cte2DYoRzcC4DGNvIr
rC8o+u7mvQR25p1XwCnPRYsYFfXMWEkhhdYkmW8XHaA4xY1GIb0VhJn4Nwt36Puq73lIhkksRZts
6eEo1kQEm88yaGUSE5nVNQG2gHCnKyeGpmvsh4K8EQbY90SqJrxpyxXzBEWxtSuj7Z/MIUtp2s8M
BlQhDe4YHagZup/z+ccKSfAPOy8uPg7JGBjntnps+8pHM8oawxG/tI8x13mVjQ5aigIfVNrTTUdm
//6RuKR2QlHZigp9YbW5ufajcUoiDocQ81gopoHPtfgp0QocLSu75Obv5yrBd4nb0rqyhS3SwHhs
16tEJuMC8DE42NPIKs0k1/eYBwFbpCkylIQZDPuwBSnJaJiqi9PFD/ba+3Na0N/Rrh21/P99NhFf
oZRjVS8Ynuw/oTGNLhmQUXKNg+H59aY+Hf5eZA9jmzqlh0bRnuhdWgdZq9/qE3yfPffvRWkckz7I
jfyPmUeVU3YkG+G9YIxVkYfvzOaSUSQzDYs8Bgt0J+rwtgyrc1kmHPTgKCDHGW29PSSR1eZzJV1T
UB+BHlSgK2wgG+Pe0ulfPFb+Tk1ktAfH88K8Yk5p5Y/JGtcbNvWbHkA5bxWIemsjrF/mgzk0v+jj
Nt2lVCbI3yQggkHzOScIvGLLbbBmsIz6BzLcvtrcCdTuUbx2QVa86h89aSqjpWNaaMRsC4+v/K1D
YJWh1e8zpH/8uyuZA9BPaoW9oppYu1Ofz4LFFwequGumQnYN6vLyg54qgJ56FAiKXr01RjeewHnn
l7BVRZ2j48o/MJCi8AlCRMPuTc0sC42VnvXWQ4cWMiNCZ4ZQ+dOukREc7toTl97JrZ4s+2joaXhz
F5fpYFjafB+ZMZSC36L/62+/MCSQR8iQqKz/V2ITIofKrP1HB/lhDLVOG3oI5Y/z+Sf6oWwbjG0+
s3EYjo34DXLBCNTS42v6j7vmZ8hy8vrzm4hHcdnXTUb0kz6uIYgTD3E6hxBMxtDNh36yM9jEewCH
6rkHy/q4Kv07Jp9/kz7UlcTvPivm5teBTYQWVT7+/YZUWqQ6CSaLI73Vb9hqJFHDTw0FG+D+pbth
tq00Ze054qeZ0Q+e1e5H997lHAkYnPoU/QSZIFBZtSiV/2nmGYbk5UUAVa6JRVYPc1kp4Y7udRPM
FUFlh6K2SqVoR3S0YZlXECStUA1AAQ7+5vAJ6MCDag4VCdiYxhUQspKUO4Qfd7iHGq0Vyg38wK1d
/3+aZ7NhFdgwSVG71fAsyH/qPUNc2XJIokc08fUwugteGHNHrV5KPULnCMJ6Z1HhFjTfwtI+cqw9
IxNpUS/MW0BiEPOsZiN6MEHtLiN2RdjXcitGcRpGNthwLtHAEVISvPXzXEgOHqkkDXsBAyvec4kj
3YD27XnykMx4I87IA4oA+HQN4Bfcgidy5XygSWneMsBNxc9xwEsMELIQnukCIJTxGdjQgKJdCXYc
d1IvShgUBfQM9OL6obvqnFNXIU8aX6q3ZuSpvbZDzdXUoaAJuMLsQ2O8sXaNmoulX8TUvlM3dVPw
oJwTZwYgOske7mwmX5rTGsGPyZVeimGitzuqBkwPXVboXgxu1NHAxiWdxNkwLKh4oI/cZEIAt2C1
qccL8RCDmN4yjdyrujgqZZwnlDGPVzyHp/TGkckF0SNhwtX+Ofmg8cyYyx0yldsNaEYcWrJ7Fhpm
DYGRgLat4h0biybroKRXe/r/9TQAF0Bock5AlsGBH81Tfxd9URNnEZTHdnOZCF6pr2/l9nezXCkU
ez8rmgJZ5Q7IJD7W/HPTIfPyPKuKrFYLbmE+cRU6kki3O3pRVq3pgEDwBVAjVJH5kyhv0OBVGLnX
jVDnmUs9WiMD6yw5JAJxiPSlbfCEbO0uzRSJUDp53koFKU5Zaq5U4sYkZ2ir9zTujBTiv9pNm3MW
RacnjcIADwvt0c9VK1Yj/ThQdNj68f2/V7PdaQw3VH/trNSSBY9ApYN3TzK+i7HTpKSpCoyNtnSQ
OSXnTwD3OXviQ9HIQXmTZDcqXBoEi4Stsh9IMDJ3FQS1SwzOfR9lCMSR5plV3gRrs+V7Swi8gfG4
f6guJXhrclUq1CGhkJzBHRg4rH+4vWVirQlLnq2LNi//85MC1+pe08TtRvHrRGUmB5UDmYJBnQDF
pdsRz/Rbhdrhj1Fp6OSsyp9PE+lYRoe63Msvt9Wpd56K9YN4Hlvk629vuq9Oal6SaUvhFrs8kfpP
jqAsqUuOW2bpLhLiU6ntEUG8A87I5vAtBg7lUWJpaFRN6foODV14IjLX96+NQ55nleuTQq0GIKam
9Y2CVoxjwkC7mnHbgF8/ymsecD9dp038wZqkMDJXbAKTALTXsa3LjryOxHU/NHHOK2FaKAy81yNJ
+dpXPa7Fm3PuyDwoUtG0H1V1iDgD2/PttcyvtQ4I6qbsEpu2K09A0NNxIlg/HB4ATO+6jGen4Gdg
+qWCfmg21yKtI7DfwLw+14mx4Sf62xXX1EvCs7pEMU7lWfSLzXBnhG1TwQGWLhIhUclsCN8PACcM
6WJ8ePiLpHi3ikU2XhEjroc8GN6dM1+3ptudGCYy7Fxw8f9YFYDkfrz/ns+BDBFHK9LYvbyeaMo2
46R6/m3v1nPsVOCGdD9UlF1b1XaKe1ouPdIb3X5PuZAL69FxQry9lRjS6/31Mh2dQ8dhoppFDd9G
p3M9gsXu1cLpj/g7ZQanKyKIcKue3K0Xn3JncBPJ/o1bbLj7yvx6JtAfvzlA4HVp9BUZ9GYDbH2z
mdXKHb7LRC080YOqZCuD3AMHbWSoMI5E05rTCLFXr5m3dMUD+GZBfWJt+6YKt78EKU7xRkzrUHfB
4r/JeKROmD/RZgPCYMPxBL7ax1zFpmsYE8zkYbrX72kRDneI2cEiDsCz7joD0ce2FZb0ik2KFOJ9
py9L1eB4nGbl4QlsfpHzbSInLfaX+CN1Cat14Efqymu67PDoOdghSTvdBXghBE8uVD9RijjFDBkp
C2YW4Elf0ZxB3RRyfUzKgxaOfmZBuuv56sun2FMP8Y2rXIBiIpIPMr6/q+oNgtyBoBkKwHzdh2nN
JSiyCjz7LQFAX5M7M0NHBBlUuvYtSC/fhWMW/+aCoopBal3Vu2GffdxvZW4nvGLdqBlJlvV0Nasw
UX4JLW8x2vf/fwwfRmZFE/I79Y9G8ldA3QOTFQO727kKl1e2F2SJOf4yZDCi97+vElVfWHjFoXLI
kFen/51Qsv77vltBkbvphZmMsTH76qwXU8TN1A8BUn+aGD+LDjgUkIYXNf5tPZuPIKGfdsiwoEsN
IHUy9dZdW4RUYNkA12T15LazdSUottc+MygIHVGdFfSj61F0ERVgKTxhdy5E8EhFweqY3ymhXo+4
vxyFwRbP9gNGqF42/YyyV4J7oo5e162wTrVuu33YzuG0wtklukyUC/QQlVse+O7/opxCCw9k1EQM
7czXvUZZznYw6ht42U0qY43BMngp6OhGZvUONiWLWJBrWJXf7GL5orgqer3KZF5S2B936EfylWs2
cm6ENBc0xkD8SFHZWCKuhdptQeu2RsShC+YlEHbBU8QA51N2WkgEFYURe2Qw7Hy4HY3Pk72BH3fE
8R+CAUpenNtyuZHr8LjVZYV+ulEzCS/HZuBI7zzf903Km/NFLFclFBfV0QjaNdypREMj3JwN675j
Dsh+TgbmA2dM+Z5v0hign0hbQZ3jV70DUZS04QbXG4AYyBFrSN/29cIVSp9t7IgWc6GIkkdDj4jP
t5Z6wNithOEjEu7e/TVvn7CMzdntQz2KT8GH5bR5u/6V1KrOaK1PlUs4Y4bA0MUsoIi6pq5jlPC6
u9OwEv4jZ8VcRvtAA3mhDbSu6PXi6Te9jlBM48ZnEPAgpOeM2KIsdJvSY/PbqnlyB/D17ccNM9YJ
QZfwzPL/kagSDVrlk9CbVNrDkVgwr5/+PNejDOvcWYDc+3rjljxiShUW+QVzoy1JAPxaxKyfZ5uM
l6IoA94XlnUUV7Hsg/yof3MmB15Qo6o88IUz0mfM3qg8yZTbccS9e/ogOLvQ3N9L6Lpp4/5Xr2Vy
IVY/mFRr/wsNADdyz71NGpGdFuA2mMGdjQjnHnMfPYIz68t75XdXNQsuNpI9Y+j5Q6JkCL60ayP4
OlEzSKOlPVvaAohUJ3xqdpPNeNFpVKd1Ej1sBoVDXSNihP7AHxxYzWBHFttucOoue+b0qJbo0gjU
yN4ykKoc01tmN7KD5x3QTFUiXf3qvh6bjVjodDK+8FzRN0GTK88kd+7cXF7zIKL+jFBmXsZ7WuBW
YnWZRX3rMPJaXQY5D8i+m/5Zlx3mZY0ALioK+XucMutsEV10I/kFFGCYsIQdvIHWfQFNMKBLigcX
mMsfBfxbKmmI2QsuwuHKHI1S1DybjZzNIJZn8rN/CeP/uCEN+PDZy9nRYcb8eUyuwW92sLxuIwkj
R8UX5YCmiaDT8Lots0SICMVysbdsq7qJENyRpZjNglUFi4F0zOpLYKYk4Fu83A3K1N5n6go1JgXN
/Z2rxpQoAnwdMSLPchGKRGnscSC5o/VkLCRajmyjbVHLdKCWlsvnYfnAZdKu8LZtvdoOwFBrg/on
hk2DhlK2QLdNSjXP1w72FG2XSkBFhIKAJHneUH39HBbR1NKRCzwQBSQ743tcwrSHnHz53uR2YvDj
a7uUzhZvEh4DGS45qVeuj6nPwRJfkf3qUEN805W86saWjui1xCs13n/6TMqZE4Ra1Yv0Dq+Jmc84
X7uQC9pmqqhg/F3AkWbRTMOuMqMzywO40+pFVWAZ+NIYNgW1yGA4dfpN33WXYeQbD4jGjnbXhkBU
EWuz0OOE1c04ZnUjZ5gBGxPkomFhsZhPCRJE2WBc3i4x/Rd2vnskq9CJh1Ui1OKbnfqGXpCP+b7e
m58gRaDJPk/y6ABR1mkQ+rbW6k1LtgZDtz53y9JzwTZbbogAzlEWO8IhD+5t42noViOCljabHXeM
P18CxfCQAg49YwWW+O5Bzj7tccD2d56mhE9LlyXal2ZiKJXMviycuLgqtdmnOJAqyabuSDR4kpqZ
mHPhXkfbAHVMaUyEJupZquvlEwEKSOPP9Kej6sITwtRQ1to4EQ7Gg9RnBTccv0MWs+PdMj95kgyw
kM2rfa8ZJ5XpFUnbP4hg4+LEYrAwx/C4IvhNYYw1p/n66Z1sBlxZY1DabczQyWnKOjHwNFV/3Go6
Aw/Oh+hqQZzQT2Ybbc7XoI9VFtpwQueLHgkl0n+SD287dkXcC0EmiJVUv4QILtRni5vtfafFURxR
FxrduYY8nHx9/kAiwaqh6+jm2X5kbHcTgADAKurcgiPSEgM65mQIOE0Z+wjE2ILmcfGymj3QX5/B
3UJUz8IT1dfjPiHJE5BoCJEFzqQADQEsIZ5tk6S4nnuvn7UlQ+B6oIko/m2NUwXuJfeTT/AkF5is
DUoaEEdw8oIx+d5nXjadjOrPd2OeNyYSujMrlw0qJyuDHzYLLQy1CQkmSu/KQdwUcQ7NLTYmkmU+
amDBFwvSfW3W2dfAH4MdUsXYG4ZrQHel5KGoAcl2L3FHbJZ8YQNPfjEJVXpFALNWFkioVwCfCteQ
K5LAHkevRFsebuDNjCm4vShn7R9iSFXvrxOeG6PhKoZJoVPJhKIcmpA2cANRvgfbIy6cWLwhvoFa
qwBvNNU1S2p//VgP7TQARomHzeEu/zkkhro6Yt72tHw/YmtwfcT29oIyED05UXMshur2zb/DDL65
IZegQ+O2zSnqFlx4VS6t5KP88aZZT819Xj4CllBtlmDxSAUqa5cLAe3xDM+fhbl1CeqiNRRqImk4
Ilhptc6RcEju3kFyZsGy7YvNP8wTL59/aMMhRXHWqjz0TYiYlxN3B4w66H2OXwr/KtkYd4+ASU4u
bY0SkFNi6qpPN3S92h7c/fXbaEkBL1BRgRZbM1xlSquVsymPhQAbsDxjco7rdpeY3ukxuF+iv+Lb
rc/SqYAfsFE+JEJ+puX29WSMAlv65OLSohG/qC/pzfXFcMjj8DPcpvtr5sr2n8i+RnxyyD6J0wQ/
QYCE9n61octkVd+kjNGOS7XZjKN93A4AQCzxXCV9qQjMFaDQsQnK7TSQ53lXIjphLlkHjhXBhP7e
z/4qSFAsX7cemzMk2yS7g8ZZZHHb657kt7BuNEdL2J/QCi8//lwGrVPnoKr0YNjmvQmbSUhqn8AJ
wL4hpcIZCQADm7seZr135qc8zGyYkIHC8+UD+Ni8mTLhNCyNgtowh0uKefLPNMVlz8wzFk7q9x7V
9D+jYRE6TpE64vTqTdNJZ2n2uh9BdNlBW1aNnH9ZM+pAbYMj7X6QQcuVOh8jKBH/82NnTFMRo2mC
OAbF/V0qH/YIrLNloOyH1b53fpvufciyoP8w01AGpJHU4bQka3WMo3cdS/jH9PJ9czUIJfxXTO05
npHTGK6zjYTIrzP2KXOInnN8P7cEtUVMJok1rXLtObZK1wtm6Y7Z9+5/V3s0qnc6+Tb+hy18h5mp
OHq45z06TSG+Xy79N+RlkAo1imBL71yYspq5SwNrQL7n27zvbrM6HIIUgsKeqrUOJBl8xGQU61RL
53aJ6WmygyyK0aS3zIURs2K7VoEpvooG+0B6SjBO4PZe6MMHyCF40687f9Ojk2wcn+uR+f3CYyU3
I3RTRpP+DIRlA7fw+M9qUQOi/+jbH3jZwWmQBMcH0eLljll4Q93nyDtVrqrFdn3+JqusFwWI46+V
BgATnkI2Fz9amEBQTjvwqQdVdP2VYGFRi7HI07LP4B6SB92y9CPm3vmR2ndzu/F4TmaqCioBtxZk
mm96ZFSlOIKlqEN+alVX9clMoLJAC8WoJcbLV49ZnR2uPZpJ8jedXCI4pL9z6KVt+DsIfpE0ZHkp
2s2Ro14dHRIa8z5WAMO/V88El2yH333UbXnGBCy696ngksTqm6lf04s1QvMx+0/dwLY/6L9s+kqh
/Bzer8b9rTjwOpWqvjWBrKv6aIj7iYy2dEyFsPa4cMw0jqegGRF0zaew0fRD93sIJkZpgjWWKA6I
BZ1oOYaK84+LY01w5D6iRTaVD0lUzMYJkwWBIRewqRj7UyQNmhkq11ZQrRgKKDoaDGT8zghtZEhr
ZMFngoSCYJUF/RpAcdwj3cgRDe7ffoEkfHWrhoHe6xj5pKZTWr9VKr4MoQF1fTOwd221tY4JBk02
evBnBmZf414bMtpMawaJJFF/hN6HouNoCnx+7mkta5asQHIYJsK9fJztkokf+4W2JKPZDBvDP6vv
7wyIWe2heH85cfGRdTUja4OfcZweGEpZwN4jQLo2rIN6ujetVzbJTx8iVpUen2BSMCgkd1MLFYic
VHoG6eLUFGLTyYfwd8cIctdkeqb8kFwg6a5sMjcEyuuaRXMDXf2aF32+xB6XItvmj/u00Nq2wxj3
vhB2YP4z3clAtCxdL2uWRzC1u0RR3GscWkznH+LfbuicFEISGos8VAapUfWvLjFm36KJbzXWaav6
8E+9cS5I0rwhiwVofchnXVCYRaF4+VOVZVmTbKuSy6phVlw6GGPM4W1iHSXdEFtP0CEknat8Yvfl
/WT+GHJ7LyEvFNeF4YxS50M+6PterwWEndF2UHWuzWLszJr3JsJkFSyCYu41orS2tA77miFdI9Z8
+8pnICX0Iyc9oVBdpYg8i2kR8O5i34VSk68YSZY7QAn/kww5++mUwMh0ITch1uev2TTtYgSFdbpk
GUmlok2wdTHC3ouRaPAV9v9yaIiV3GXsn6DOvIxQpeMKrBBhZQrY3uJ3RS6+PfB74E6j/FyhWUfR
FRCPUXkCH/JLH6LppTVppnueHH4XIiOLYjxZrA9O84nZi1/oQlZb1NaUHsJJgn5nxMow/+6p11bH
L43ZpuQXtdrciQsXiFTmiusH4pvzh6k5EMRJrBpkjKyLvNiiItIs4G7sH6W3CBEPvOmpIVu8flHu
1zv5E9IBz0CwjZfoC48GeGhb7mj9rHR3Z6m4rKtmfJp/ZbMVZ5w851BTUVj6yRRDOWZVnLNkAfwI
2cUuLUMsbggT/KA1raLqXBirud5dRok6Gecmfys7kM1DRSc/0QrUPP3Qiyh3VIwhwsGBQXWZV105
dkDYZdpjieQ62yrCDYGJqdZkNAGChJuIxudw/eHr5ZWCTBxHJlag9t83RppjO6gRpQJ5A+R77wMD
ENgoN1Nysdgm29JEC7WzBICrpRxkpQKTrcJLAgBZUoMwcAFQE9qiI7nu9fEwenqQ6U/7EoMiFm1o
GDvE3CNsMTFQIeA8L0iMYsSm8rf+a7FjBIraAFb6XHo+w1pCH7Vxeumr04mS3Hk2DEoT3QgLDluN
/0w2F6pRYIwaUPeAWPfkl+bqq+czDizaIVztQz8NrxdKmOLm3+xaT6CC/MCkeAOAZGEpPtjFDDah
huc6Ybobt5fJCgPQMTaHjVDB5U6SdJZqnRpuWrhnbCBuvViUtnSdZE+zDxSyKEqFKYrJYdu488mU
fdqDO75hwAqosJYlqHfP8tGE6kWFi2/LNUASH/gsOtfyF49ZbL+jP/SlRkh79d3hb0Zx3RHFAVgy
yxoIXU0XtGR9YsheGWUIc6nwSqHiAailDGjgACjNje5pyXFMYISgqhOGsxScY9JCBiK8Uo1QHaBt
K4Y3sCd6rJKM0WQ/W5Z+k/f6iVG06oELrILz/S642d8ChQocMYdAgSznisLXbNcxcZL4+dJK8WIm
TGZEmhH7CJU/1UZNn0/9QjG6lI8r2g4ISu4I4/fENYVdoF+LISSUtEoTSx5DfKEPCTroUVc6gMrh
qHRjEcbXQ8ccPfG65iTSYv1NpqzQYdn6hFRn5Mrcet3f6ReG6oHpLokBoyie5immtsfKqqvIAP+w
ufO4qFXeF5NLMv218H2EiHOlKQOWMM7V3VKsGYO6hOrplrCzKEnvBrtdANy709NR1TZwkZapVcyP
IrOwQs1QvhUpapvAPt8x7cl0LmIr84ASt/j1ysUoByIMORW+AV/gUtoCcRrJTlpjxLQ0n9ouEQIK
T5HOcorhoC+hWD7se55Jcscn1Cz9xwikp3x+LwslojB2tmeOjCytXOAZbl9pbeh9E+C5ENTHGG4k
br/142eCLiEo17j/GJw3sRf/piAl/ZLf/alyS7tkU4+lzaRGOJbrNuDMF0PRBxWVP7YjV5J0SMEI
Y2OhIJYRlvMHTGHrcbZm6zUiHzgkgY0s9lVyDyn4UC7YRSON+Bky8FAs38HPA8u1xS8M3O0C+DOf
+1z6SNFDC03/F3rhV+tms/mLYBq5YMlBQTG+z9Qq4WpSnYSX6hTaV9IX9c0Jpy76YZBTai9PcNV7
jKA17zPRffyQjgVDMwkH76B82wheKvNm7xqGQtlEd9YQRUzJIVujk5nPMChU2Tx84U2TPN4ZxyBa
I6taiOQs1ty6qy+WpaUeZxktsOg1fG74PG/w5DCD44Ic5kuG1sjkIA26srE0PFpF+9MotR4tJ2N9
amHHf67gMfSyr9VZVugWPgU8kcQUfSw+UUYUUn6SrDucj4mUYbwUiXKzhokDzvhxr492HMlEg7AP
61cKB5YzfJlDQnLqsqNOtuCpMdAcbIDFp2JN9PfWBi0sICYVAbKcTsr0HOTrSrH7S91kZZuw18yp
eP2hSQQWR6Q2clCqf9qS0IJ6/OxNzhO48OMF8bbcP1Zf+4FiRxRdfniylJU5aIJen4zY61R2Ei0e
IduF581s2PrnyNOaQ5t4AfxLEUfTAadunS5KDw92qVVU0po9h4AK2tIajmgUBtgWDV6RjldDhWAl
xC++NHtpphUnx3k2hrJEvgqgFraAJKG/WKCI3lgjoIhJB+C6EiU3HUviTu6BsVqlIRtMa7eP4BMZ
6kxMTZOOshaMNii1m5LfWod3hYLOyxjI3M/QNjqbCgRuldSvXsVPtEZnLUyasqfliFCMCNAL7mkB
+DFNYFUVnDTvZfuX613Xn/LY/bmHSy4okjCpRd5lTztxLRkzhEAXemciz7w51dA8m723iOlQsBau
zyCcX2KM9tiTQwBozzw2VuSEceXkqoR2ZUFPYeYl+7KhurShicss+R0B+U1VSytjPUQWxYPeSoof
vw/QISHakPZ5c3I4Hh0yADCh16RJF1Zbn9hAaLhJ750vOIAxGmwKehAe9wgwezuzSM+aVObWUHFi
t/qpQucz9qSMcIP+DI/eI70Tm6GUGUS3plG4URr/6bhJRPL+mCG182yK/qDOLt+cs9jwvwOyGDZC
Cu4Edq7yOXYi+Tq0VJoAIIgwT723ALIHDSsGoAwQmBiVhLdqris6SsM61fRNuemFZJZXOtnVQQc/
ai3drXlFu+rRsxpKT46Bu2fZ1nnE4bVFI11qhdb8XKa7u1ikmFFA2gYodCzakYHBMK5fXTzrT/cp
UiycvnTdf7haK8hyrOY7BeiYL1ihJPmk7lawL6g3k7uWpj0ECCWOn9YYNzZBSfiljHGVIr4F00Qz
ifwkmAWTKtZDd8+rVfJATmgJWo05m5i1UQgK2F++ndMUDcy8gaW6QP73Rrf8XRUddRruzrwJglOM
LXjZrQ2uhLrre2zg6FPr1SmhDSvNbCnJQR3sZroYpCz1FnKHb9AUcVo+RZwwXRjaJ+1ZNOhoUNkZ
ktyQC28sOlgadQL5FTViOiFsc93fm9qT9FeIrO2LnzaEVcy/M13QKD3ny/npRf/h6kDL2QkpnC9G
cx+NjP2JVnDL1zPwFrQ6u9dSDI0LV+Ji9Q5+bEBOTkPib1H7kZGqZpfMFaaoFZE3ZtGgZJJYP3Bz
+ZKQ5MAELl46hxxrQiDXmTXgzo5rIjVhUtRs2lKfUCY4oHTdiOLAdcro2qC7Uy4i8I1QMp4c9bCC
0wFsSjqX6hDvJ4gf0+NwPIYzZzvPq/qvxGo5oinvKUVJCb0BLZuNKg6LXOmcNj2Xzcw40p//Cc9j
cHIcPDy4wSsRRCD2T3ao2pXVTw0T4pr6tpwpzREKmnmfCbsd87zfq9G/pT7q45BDnzDiWAIdIXi0
fsJTsKyDuHMSDPewjedvxydgIlUlFRzZk7/J6Ll8SpwDS9X6MeECu+cX9ThQhHtiBwF0o/G1QLqw
xIyGvEK0sdoDxxHuiXBM3ZRCaXuvKN1vqJ7f8vMdgDqzzNKaYTDvBEM7iUfSplmAQwMP1JbKrx5M
TE0Vqm4+S4y7kmEkTOmaORAnsst7hy7Vv3gcdOJFCILwiuaxVr0/X+KO9nC6Sk9+TG5F2689ehd2
rrb9lOdzoz4Et2caWEikrNr7du99eQw8DnZ1bPjULRZqUKoukjjDvFEZGSYwPNDblqKxKBZalSBs
Y/zl/1A7cCbaxGEzz+gpprksuvPd0Zbnnl21Z3/a9d3hZ/oEzr/9kQUoG9003utU5bHkIrnjYp8G
VYSMfEJ0oLmMED9EsHFTqqsOoqzKbOOw2SZuGz7/lzavdIua3i6WQxjLaKrFtP4T2pOMtk/1pj9V
+A/g9Pwq5hNOCb7jt5kTg5WJ7dBig548rBtWgtcPob7/+cMny38vHYw0p65UfEK/EyTqenu8OmH+
Ty7aVP3Pq2ssTWp4tFi2MoOPs2GiPriu9n4Md0SyEDqsWq6f9IXnjnqLvACIAZGMZdZLA1QKmNou
Koy4wofJuOCX5v8jiQQU4Lzm6TDNhGbIai9FdR/TDljylntod4F7x5d0LnUrpxiSEJ5PslDCrRR9
1PCGD+qwyneFTJJfvpNR1mOgIH7SmNXOuBpv/hHNBdXy7/4b3UJ4CC4SG+2R7dnu5zobeWQ+lv2M
ljC/UgFRIlVCtlKPMH0SpR1ClRkxZEKeNvG2kRYnTPKdNIbZepYJTYPv3bi8gM3tEpye6i2RfOpD
IPk5G3WgxqfN0Y4TKx2T2iRP+Luw2+IN5rDo8Ck39RLUvjJxqNglesDPpR49drtbx6g5zgaW4x+c
/bCXfXaEKXlrU0cqfiChKHD33onIZyXidw7y/ga0j72+PAApPh2FcBSfrQmOVqmRQrCpEF25qQAv
PaU1OsXIz1SAp5AI4fmizH0DDLYn1FzKt3xBTdQsP9KS9tVw3FFxhu3EmI9XqJRM8nC4tJo3V1QD
9TeLHp6pQ0gUJ/ZiO1Xz9yh121eck/Gvgdn+8aFh2YKVROKr/LisdNt0Aa3aaI+o3UXMBweWu5/Z
BtuDeudrMlEiLqsaUsg/xjmA/mopyT5hT7iFE7rUU5Xxf+EfLp+G2U0/xvXVTWb92N+hP+I4vNz1
P0QTMnNDm/vmaq2dcQ6eRdPshCcSXC1ZVzB0DfB10oV8+B9j8ZPUMXJyzo0dhN+2IITgiPmi8lQt
DojvXmRWX0htNDBuyCO5gxq3VA82+9rlkm9FJxMS9/alndJw+pGQXfvRiJmQrkX1bKcI3KWd00Ve
duJKhZqg/qDiWpsXXp3P8iTlZwq6N9VlUBh2yF29IRIPymB7h+FWGVXKmjgRkdR0jckERdzJPbFS
kxSmG1RLNLFZFXg+wAt2xALE/VVuqWpHqP7jofZvOZaDRS/uXeUoUYqVGgnY8Kc9Nt6lYbAeARKM
bvJFjszr/gFgwyCHHrLVOUaMy7Gc5vffhuGdzrbmOumN/2kVWZptU/Xseq05oEDDiI6cbOOngUMV
UDERm98WO8/d/PfscsIurNFF6s5GchWPJCpQx9Loc5yMZmz+19xzwP/mK1V4z+eR9Iv9JCpRTgb3
AEdpG2T17vcxKE+HgMY+eI12H0awLclaM964Jlp7Or0Cadq3CVDC9OpVgaCOhBWO51DJo5dtVf58
lCLlL6FbRjhB+yXf50JZf2vDGRb5YAhaVu0B7tNNeGqKzvZrE97jRVbs6zv03dOW8ZfRqQWQ7jdA
6JhH0QVe/Q/C8owCCAQ5ITWRqbQZmOaFQmgUofbOn2CFJ4JM4NznRMN4xbxju4C0Vn4elTLgY75d
gwPaXavLmkO/LiKDoFy6Md5Ksx6ZCX9lnXbgDEtEBZU8p2s8EzfoOQ0ZtC1kjJrCMelVIfRcNL1m
4uQe0Sl40Pe9AvVFAUpPiDCxUfTbU0diLgMTPjBtPvE3d1oLKGLa5KariB9UJcx25Nj45kAfsdpR
DM/jjRydZrbT7Wzwqt2TlcCnQVnQbnRi9fPV3TyFpTRV6kYyGXMkR6XySG5pQsZDLohNvkGeXFJb
CxASrSoDQKOJ3oaacGcWKueuJhjlvtsj0ZCtiLwdiExokxbty6ptyxD2YDhDB1omKotwBVFxvGkI
1eh21BAErHzaaSfqnrZ+I5VacTE/5wwyK0oQNj69GGY0M6f+qTQUCIC0cAvrm+wl12qPE5eY8o3X
84EJ4weHe0lmaoWxkHYPa3JnFSkCgyXUgYVwD6M7g2qkr+m1/cQpiDt76tVy5WMNJwN+7K9MUhaE
JZSMyMTgiWGUesz1bFaXvhRQihOl4IDyMblf5fCWh5uanK3I74dbjE04/IMu7TFRGHB5QcYe+9jP
j1qg8QkfOAs3z7pz1R1NY5S/o7NG45dZi1Gnjc54wYqoa6gKafkfU3e09Md7o9L07t7qlXRy4VZX
I9B7qrsBpPG4yKziGOS/CmMAopkDQmu6jnioESKjeSmNTGQRgXSPybQL6VFyZqEg74FpLlusZCOU
6iiw/922Is2Yy6+gdInZm4/Z1T8ndKdBpfiatJtFAno/cdulIljmf2peeKmgkAfLVuvODck3G0Yh
cdbLMVa6ShnxCGcxuSGdinimBNAmgk11pfepTnor4t88lR0FEdQROewOxRuHUklBaP6kvopRt3EY
Umx4opTwDP3Z+VrEcNZ6l0pESw4SVt3yGiLodE4h2J/oZaUW4OCeoD8ZsvIZeOxDEvBdYjgSU2zd
U3AEW+Ies1EuBtiOR8HLWZ2hzrujHLORxm7NoxqxdF0eUQ+JnE7OrNiyirknnzIZhoWSjKCRKBo1
8L0AS2AUU6Ry3uHO5xjUUcGstunykpPZYz/irG9xxKynMiW3AONgkypzU3FvI4raO8mFPbVGoFPd
+H9r/o4iyD4HE69b8ICeXOMDt/gWM6cev4FLmpp0bkbyeOP7VhTmmTY1WA30lM8C5bqxad9eS3do
2VmQ9C3dPdsDVVXOyTHDNRl8GvRM0GatJVgOWPO/AmadvCBixv5N2cROYDZ46jWfoJkgSDz3Y6M+
Bsdkplf9ceIukPffkk4GEtfgyZbpWoRwNf/gmlI93v1NIrpDzxyQUyf4iPyi4uzILO/CiBQGkHQ/
6Mo0XBekBCSer3gWzRkeeeqjXABepgrNWBmdR69ib5g4Ar3v2+tfhsGh2l2dxbcopRzeNQtwgncs
ILAjEChs0SXjJuBc9KkYF8iMYFLxpaiylF+uoReG8Oio19AibyjJuWArZPEDrpoCJ7bY7fucaR2E
esShvf1+mzwTGPFXulOH3KmkoJyNecfTIT/j4R7IuWDhqrbMYn/5pAMDeJ5vs5cIkFbYt1FfPtfx
l9XBu+z01sGZCyuXMUjJm7fYzmt9HJ5t9zGIGwkAYyK5ZsBxLADzKqt/JWAYF193+5U2qArK905e
oOfSnlfArvSemv+o2RcbbOlyyFt4qWpdDSsR74ClzNtuQYLpdDnJ1RJ7IhefXtlduKA/a/i4i7e8
TrHpsOmhpFOwu/40GZQvxd3dVxNm7JixMbjX4BBvkQaWEmiDZYhbB7VWOVO3Xt+hucxkQIfJ8deJ
0FZ7oO5P0c4Fgqy5zhbl3VVnf5HI3BTeboijYWNHPj91h7bN/8Q15vU1V2qqC+UAD7Bw3q11SaYI
VDYRePomKSH6/Law3q9SRbTTcT69a0KfvANqGCFk4F7DZ1qo91Qv7L2vPPHdKUKR7x6qsV81uK46
k3dl4zytgm/GFW9mgbBdQEskq/Bzvd0ApmxHVOoLXZt/xIWN3KFo5juuVTB/8nqV+z4Z8hfJtYzP
Sc9o/Fg4UgBUlcBBBQ6y2vRw8Avveck6I4k6lvADvJaObZm3JvOAYIJaWsaimee1POsl+Rhltvah
yRpM2gBlg3yPUIc18aki1QItD+PsIpR9qsLqUExsTwvBiJUstPD2ToBGwvKUhvOufdSjO0YNzuh6
+7yQDllv1JRlm1Nl6KmKl36xJ1AiHLMlZz5QvrQEGZT9xS1Uwz6GPzGmZSE6yUPPLB7SyVsNdVSa
fTR1N3u71nY/53T20kBGLoQXwsybV/oy4VI+dap36w1zeSl21FvPRsMayPgy+cRLSrLmkF/7Wr6g
wC9cbLUBqGkPBm6sQKYAsUfAhJRZxTRapvgSj2UpAVKR4v66hlYPKto4cjsMdLeC6VHkY4JDqNax
r10wCWT9FMQu8ES0byfTI/x2mGHzoJ3M2pDfBw6K43R8kYjxB/Y9oII8PWiezxqBhAOG/e9la6tN
BerFXpuvJQaIKP8KaRNJe2Un9mfY6A4JyoR9Jwpq8F2vI9ty0ErAiTTBOzYiCqk/i45xNK6WMjRf
m8JaTjEiswRgYGl/0b8u1WBl7nuwW5gpmLSSJWlkIPd1NtNGOezBAcZM32P7Hz//Sy6QPii+XpVV
D3FGhfAKd6eArgKerYuvGcxdwCXNPld5Jc3423uACyGi5TtbMRKFxKRya2w84fLLMCnQOZDzpUUQ
2CwyVC+0QUGl9xomNRJq7fHOXvlovOYEqSzlFv4loMmkHDLyqGtnZ+e02chAs9sysHLWbX4U6IhM
aW9pzdxgkzb5FR1mWMYa9kYOCXPQtGLrCZobTpOk1+U9qlVdVX1yoCgKmDz3MQjUAoLV2bwR7eog
7RiMOY5QqQLRirxaxtz4InWihWjEPLyezEIB0SPMOmEIySNrRRJlt4ed26CY3MIxko5azg+D3fEP
bLcrF2vCjoC5QbBYF+vtRC484O10KIGlPKam9sL3su6uAxgcgPJTBP0CcEhw8o767+gd3MhAqFnF
LNv8jDazJMARoEoXKMqwt+rWxWXPl3aDDEPkFA/EDn7ZH2wdIJpwRUQ9GEATB8U0qvajGoKNbei9
G9OJ3e3ExFRdjEkrTN3Iwi+NezmyBqgebIL4Z27ch/IKWnH8stEuz7GYi97Hxf/+RO57IpaqlXdu
Y5mhhga4xc5sbKAaZ/hrcOGXmTW6K5R3pm2hjzlNeDymeHIg4NSDz537wVWP5qE20telBTPN7bJ8
wa4qOJ4eToe98gvK0hyMpl3XwJAZrT/BF9cKQnjMZqVEjFFf/G/fmnAXa0LdsvoMdWH1DOhKSPDs
89qGAGiahYVboxvfztq0T4hFT+21gfNzXUq/EPH1CJqsCULjFCose+koPBINBz3RjinSJ7S2knsP
6m3RqvM54huYyHigl0r4ua5vA8iLGP+Tvsl645+D/NlyU/jv/lO4wON7GOb+a+T13RfxvSsGf2X9
eBvvs9RwDz/JyfwUHjeuqDEY/5U5WAR/nrqUVxQr7CHrhzak0XH8IHUPoE1Go91bMPWnqR6r8HYj
qDkHeBdEsvUf2kl/5JMxCw8FEzrqHY0G28LcChvMCQGeAwsWF/ikcaNaT4KHrwVE83UQuRzeEK4Q
/D6a1+eQajYbJCNAtslfxVjC83ddsMCvJuecCFkmlDZefe+LQpi4674F188FmmkxfQngV81H1aoZ
fn1llqlGkVkpFlW/wl8fkoAoeoVsgB11bvqF2v9oregMM5UrWVB35KBZEkgmn3T63OzS8ZPC+QSX
hV02/4ClRA9ENWpmEF0pYEYM3qIoXnzACYGrhvHIK9Drebeb/rnLkI4PEZtCaeHORrvdBjWBwvXZ
fw//an3T3nWhsjaroEbWcAJwWMWaWr3KCem7IWpjQ/I2Qgm6fi8PrHN5KvTFZ1ZEkhidY+KsQT1+
B9JYh4r9iyclnA3TUu8hhJuJASpoH7GxbtqUn+qOQRJa1ZKc/FgH9QLXmVK0hybvKp7a1Jbu2g5e
6s9hpLh+zAikBExkR/JeqobAlZfxwL1oYtvvjPN0/YhzBK5lz87AB/+7Rl1GKnhRLcKer7apbGZo
THxZbBW8Y1uc4C+9JQ7JyPRxZq3VUejXXNLCEdJA3Xx6VSlAEAS/ikv9jFW5pOLmzhQ59YUa5S0q
uubJduRs5dMxFUpHm3yJZgf11gAnlhKaLgpGTFXuNxKvtKA7T7S1B/dGS3a9AOuV1rWYut+18mc+
wq9jDYdH8AUb4wRLo9QmAoBnZ1kNjJqhSQrcRrjPHFNolEp5x1Ks61/VCkfzx6xZ0DS13J5JWK7Z
//xrQ70AP8Vo4WxJFF+5lrXOu0mXRrHyfqZKOsV5/4H+OcMXgzp1zD8kJ1NmxEW+TxbacV1nmQjg
c5Qf4UgaTEqY9Ntg8Pi/DEBDthD9TRxINpGvORw/oFxlUw3TVrqI41hUFCqBDL0NxhBxM4LPpWjT
nnbn5UR9fvpdteE8e0vAVaMYxltlulaMWcSr88ZwA4K6BsJ0F/gon0FAY7jWDQGnajc4tCEz4evf
RKkJGho/nnAfbCHAP8hPrwU4qqg6PBOHlZQ5rqetJxu1LzHO13OoR/vhmcBALSQ4sxdpDjEOUF0W
Rv8kqv460NtZJV0yyDyWmAZf3rlB86xHlDsaNTd7Fp3Idb8aBvo+gJQQa8fcopC1MMGs4I81laa3
ue7HBnGARjGzhW8UGKKYcah2glC8ugCrZ8tnPxpZgb0ug+DfDw9lmyIEmSgfyJ4Xp+aNJFa+ZqLo
K6ffYJKGSJM5We61YZK0ObHVdXNKYaxPnY3zNyr/ZpAswm/k6XkQT+Yy2SGaCS+AlF1KpLRjpqwR
qhlyfNjt5cK9laYGiqwGwLSL5R4KMvSpXtsezhDhSC97GJmEDuKayxTSkc0l+Y0q4yGSRO4ICzv2
LJtzytLEUbIdcW8zSKGBA4ukB2FJyec5qnc16qH7NoqTG5HhsGk4qB+jlCd9mG6j7cTO/uLurgC+
fOllHkjSjRZI/S0sfM+ykQqCw8/vCui1ABdPAXURab2YWIrYlDHWFKnTpbNE1SZfGfqKkZywC8To
7Cnrhkl5V1jqKglegXCkMDIGAjQDUrS0TV4d6l8/D4F0dzWxSxaXuJFGd8pcFb1aHtoBc0EBKemo
rz9vZCqPZY1QV5Ur+l3R2Gr4dfcIv5gT06Npy2D6/WQMGVpeH3KqQrzj8BEKaARpU6LP2t/VsDql
ncnp/sHNwRRRM5U5Vt8fwLoO/6tjgdSkbPZ/BnH7/8qTXCknHZjFPW9FSA3/rCHcZQRN0ypkXw6Z
46JCMC6hT2nFHPEMl4vImLpbpL7YKbSVdYGmRGWDnXM2PAMwI8BKAwTNHIHXSY2jxrzS4UoeCWeK
aWG2cTRHMWQGyU8dweu2AVXBKizCvXZtfVSIvjlUVUFULeJEN6LrusOt66efxWAhCQFoSzj/N+GW
EaaygqJ3GyFms1GDDlyJFQZyoUmC+Cbvqc+zg/JHPTYTBo2PNwtGk0YA7wBW5K10xTR25w/oNoOJ
8cUV9pwPw/Ip7cVcH1204lBISLfU4xq2TqkNdeDCAhPtgikqgtMvjzIgbj0G8qdycpYWgr/BdGDP
mFiEYh3eRAE1jI+DxyK9ASsGREtFX7rq2yWw5EmWnjTl9PI9aIwS9Ok6PLJrpsPf9WI7imwYYLxb
TXloDKk0h/hoxwgc/C2d2vz7ITARrM3Iy3PbiHWqL5L9+cXKgNMauQDExaBNy8RmcBndBT+0hGwF
62hBoXp44WhxYTGESCX0UNcDoGvgnXl9GuejozNx/FPDmvJNxlZGOB5YjNlCzUm4t7kG7nvY3bLA
6Csj9jR8YU6FXPLWGPL9QB8VpFXCDr+Xqor0zzqaHmRsSPtEZc2Z0Qfb/rO/JCT+4UNwSRKvgaoL
XU9N2NyEjD2JgivzbMoHxuvEGTNgIdeW0SIjHhnLeEsEmT9yOVBO+moO+3+XPQeZGjYJwSA3NVnZ
kX9i729lfD+ruiLTw4aFE9LwD5Yt9iP3Czf/yJAweQH7CVCeFRnIUTp0FlwnxaFHX7GCxnCDnewz
XZAkXXU1Gb9FytEsRH6hrzgnan2iEEhFb5D+Fk8VawOMFeyzRqkhtQNb/CYWUX9LzyllJGDbiwuO
mg9hBc15XOyt/Ow2dIDxXwqW7pFIwuKF/B87eb/S0ySSmBgpaT80iXhHnrrNmbsWU2Sdd3HQD4AO
xzowP6r/NYxsRdHQzC7XYxL6dM4HMv4C4f3plFSl1n2HZWeJ9OkNuhzhjdMB4mGdZFCARPv6GjJQ
gQuoqwpnQCw+Zn2R0624U1GCkA4HnIIbteXqc8MvnMga9XuissIOpiDlZAnvl3A6Y2UowTe+WPVg
u1YIcqSk77MXeOIgyxojgKDd7JPlFF7Owg2MfJQXfo4/c39uodh6pQ8R4LyD+lFQO7h8cPzCfwZr
6+OFNcqWMRaDi47E/9BCSJbrNgoTnsSRkzeP7ymiBgXAu1J45ry2VkRl0sfNBfs7TkBn23omMpn3
1UGqigLFedvh+ww1dYwOYmeyT5IvDrFdvlPH2SUaY1lFs5dz5Ivm5n1jzwScqFEb6KQYNnoXvWOD
GuoADO9FiK9BuUoXjXULuzi80LVC0ccngmOG+16NB6SQcWFaAKkk9uDhxSyrmuxgYNneV+b+YR+2
w53Jr9cMBekWcXnm0hbzQINjPYZDbjfZ8MkHMvO0hGwA+it7iUU6jxoVwTPLuYH0GuFhgstoIulg
n24I9Gg6UymY1HcZzoODXi4wzGhYIN3j56gKEY/agV5zVRFnIVdE7hSRrAcmkykQJQeSlk+Gkecv
ckNSvkz8U9npt8gP8pG0xwwMl9fELjZSBDzDLN8O355qP18U9dSr0PMiytqGrob7p/3WfH/0qg+w
rAgHD6bh9dyr933Es1nCSNbbDEI2gmYA51rP/eMGQWeD03sAS+zTplRaZ9uxQOQGcVmHH6eERk1p
mZhU9O+joTNQas8DGjyTGUaunFeAbQpABsYJV1PHroSQiM1/YtRgXIFTTJWloHHlJ7WnTIeddxsg
sOMKiqhrA14eiQew3s9FIVBZ9gxW9uqeg05t04uffi5os/6tNFLpY8A2Nh+RhgXj/st7MXluohIa
SUmG1ITkpuOMgB3nboS88duigb9lDVQy0iwwtBHxyrqLZwbwMDvNs+2upbA6Lt457e3lf4y2IOjh
xFkOStJWBT1HN7+TE1QysJZrR58qYda0L8nH9+VPsdg+MXUK6iXp+ByTTRv70fcMIjpnx8dbodkE
TvgorqhBWP2eHrS51VHrCgXjyl9XDmBLMpM1go2YlFDydB6DBpZeW73pgjGTAPkrt+vH5f5xamdc
8C+pDJbEGoXZT1xwnW4hH/HCOZN/4iivIPfpDzYM4bHcveY+/XNT8XVZ2ZiwcZzGx+rwo/7gI7Yv
GtGffzy29fbjaI7xM0doXQyiI+KOkjjaVmpBGwm8cLV+xI+pVqiv4tRCiFgr+MfGYZBlqL0Zellk
hyiayDPRcam8dkaIBQ1j+7TiTEe9JMUjprZIceksu4Mn44QyKBHP8k5x9XJ/ht3hUglYWmMdaiVj
mUyC7Jm2yafINBJ/vK2AruuZFBzeSxRAAnJfPM5t15WKNJXjWdvCGr9JzmB93Ow14DgCaN1jCtGx
lShr9Ju1z5x8Ll7F+gid12MxdzFP4maDkgXydaE1kvB6RODrTj4766jJRyWMfUXvpIykmucWTIuG
XVq0uKUAsEHhl88S9WLNqHLRz0qatdjZ7h4dxPp6SjITHDWeOmnjlnARo7AvRdCtSu/Y5mC3vRlg
t/aABNWn8I7QSirbfXbZWLjWJCqJEiP1uaE2tPKMvB1j44ulA9j9Dwf4A+CCQ10Nm1cZnuMFv7We
wTqqfrTeoC2hZUrkLkzR3dVuaxwIfNsn5pePXnODKpk6uXJSNIHfLqaW4RtZBhDUVDCyJ4/PqjNV
4mwFs3AtYHTr43OL4wpJv7EQ7HZrNcL8ZAFYKB9Triz6GzgcLU/PGaeJxRXo5zarSQOzeRUjqxyg
9A8bP7vCXZCy9UKg9vWYPCSvb5gTp16yy+HRAyZnTThupq3jpgP2tEck8Samrk1EU78GgmseFaU7
DgqLOptahP3aCG4YAh9QNXYZuTm+7jeaOZYn6vG2a3UrqcpP+gZpKP1mHBbYQmwcm9I1Qv8S6pt+
7JSwbs4fC1vGGKVnYLTniBV8iQuzMfdYqg3AQb1syC0xSOVrGICUqMN3/QgIU3Dv7vXoJBn9T2Zz
VyVWxOkWOsadLOIBKfYyw2fXftq3rwmurE53BImaGjJv5gNZahixnM4Pwz0sm2DOV9M+Ud+od7KR
KD7YPFC4juT90E777eZocUlEkoSXLSgAG7YfUguDNLuw7O8Qrn7TDG05X8DWHP4oRdi/FlCZh275
uuq999VQsGDqY/W5nJckGy2LwP7b8DV58RqsoWQVCZ+3JoLzW0CZ7jJsJmwe7XWtbUtrme+Elh5N
bBfr9BkvGpdcLuOoAfvuWvUQRgmgyHKsDAB3bIBACZJk17rVh5ChC+DSnmnG66zrWp5KIlpRi4UK
NS2+ObuGh7QMFaIrLnwtlenGjYP2m09ETsSfLNz7bSCIye6qoDM/MYaC7UYypT28Z6CZnddRve9N
x8Q+cLMPZ1s/j3Na9ytmLoGOBUBsxJ2SPCMiG8VTBVzsMkxJA07YspuYu6W6OIPOtnM2BjYO7WYZ
A1zFrlR7yrHM5u++0cBB+DxM8sZ2LxPgO0tfkC/96/zC68/ifDsK5twa8hUd4S4PDjuNuyKEdjNF
VqdU/boTwrxZxLEsq1koLvu4l8Pyk5euaf9BkxZUd2qhLltKH3DCi22XmkD8xzgmN7NksmXhGeBK
pphtdquyl7LrKtZIA7g2kF1MZ/TnuXbJ/GeIyd5dV2zWDCxacKamctTuQxQDKQ/vwAVnWC2dGO0b
SR/QH5Do5GkapaNUtjZb53vm5yxFKZXeDPmJJRY2D/TCdWo8EmCtXPz1eBlmKrFanWvnzdDvvUSN
nPcLSlWKkDVxpJ3NHLoyRjT5iH7K+oqkHD2tgysZ/iB6FsYP/Epsjfx+j9c4KOB7PW+40HmwdJQ0
0+lr4+uovn8D8cYzx3qqE/AsVPLf2yZvmWpBL8FrtwMMV+MHKYmeMmDMDehBGlM1o3zErK2KwvG5
YZQVUWTLi+8J7lj75PSQz2csvYs9gHP+uDFtPexWr0uU5gzXUc28Rfd/lkkdHD/daP5bl3v793W4
QATsABZpDE7QdtuRtciJMtgulb2D9m2zI4GPYTHS0ukFRpY2TGokddYB5YuNrUT3TUh5892cI/nV
byxwJoUIYApp2rsT7QNwWAIsTtGM0mn7Au/OZbBBUX2CiDsbqCgKbo8MRFQYyAb4IpqUr/aJf5aN
AFiKya9oC49PLZ9dIqAQ69sAmx6fYghcgehykAEvZNkrCgGN974XPQ5XuHDqK/KiDvA2kDMl1lw+
LjwKK/PMJy24uURXuNlNz7KftNLdutTbwTLfswfC4+v+D+8HcnxwRTtLK9/Nesw6zEuipeV9P0NI
1hzhyNFroVEBvv8/IOX7lnZYy4qN+iK4ArENh8nzG4pYZh5HUZ5GRylUvPiUeEt01u9R2wAE1vdt
lkhB7YqtOAgt6oXl7RKpz99qCjbhksu9scrHQ+lruOXLI2Qtsn5Vk8eWQvEXdibox6BqlbIF5yGy
lEyNpNssL9Dc93n60VVCrmPZGSUBDq245IM2+jOFYWJjqOiLY4S6QjQYzlPDPzDpEt8UraD4vNeX
JywBOLs338C3six2qNXi0FnHsO3Zw4vk4bOv+ljXshNObv3zmBsLSkr2GJ0tWsc9+SiWb046/Qm0
OWLZk+xp1nL+AA58iJWEhmtMNNBZG+NwfoKdqZ7XE9yN1lwDIf4JQLaiUHMFnMi+D6QVgWqg3j7U
jsGUo9RfnvzejWQHfrENsn1qXbYQ1uf9SMMGCmdaEIu8GWjzN2lpLkAWOkK0Vex3H3qLEO3I+scV
wA8tSTIsKDD4obgbooefQMI1ro9LRZZl5z71yoowQeFyEwTMjOWlKWUCYBpuD5AFd+HBJttrcwDB
8ME/SDZuwmvkvToQfmo92unnOkcsdxU8Cl3uhe0fY68lxoUlW4zxEKdyA/gXGbubuNM4Dm3R68U8
adWsPoBMKDeYTzo0gXEqXOwkn+BGRsa8HjxVuvfJjhZg9BMQ3Br1xiOTy8Z3iUmtjgOCaff5Cm94
aVmCpHCFXvgZ5VN1bWs+5LYa8R9OI9UStLAPYe5VGhUy3xafky1kVpuFKGC70Z3zRskiHhLiKnam
FQiWvWbZ++L1moNs5RILL/KSfXco/v3c9C5qcIEJq2fDfeJPBKxAyyoLbn8U+tbD+qOMcAJ6Wo++
xE/+eNbSEvfMiOYE9WQbIqOC9saYY+fnc8ZjEtbGMCF+WCa5kQafCrh6uUTT26MFm3wS6GlmfXjX
Jui4THyhImBCb1tyiK/KIW2vNtD5Vs7eFPr7ZwxgLPYuREj7kF5dOrL+ZXP91v328EKcTw8vpbV+
zP6pcw+U8VmQ79rqnubYjHmg8BRa1ef36TrCD4ayPNryr93uOLrVObbkVSkAcSn74y4fCAHe1rnf
aJGbeH0h+xwKqcPIlExLGHt0szrCRGGpIZ0mqiu10rOGuwA1KbKnyFA71Bvtr3yVrHTcXdEY6lRj
pQcMvOQZWZ4+C04P1YZuyBXxQ6VFzjZFr3T3c8S6H13HO8L9BNZbsQlsHxo93wVQ5H0ETS6uDOwz
tnYYbFxB1jiz7M2zSR/CjpCuS6QdhZ4QwuP9ddsCajH96jAA+LDgzkvIbnEfUACP0TbP+HOTSlK5
sNJIWCezYahVlqafBAanO4xAGW2+NfsTxj9+w6spCXVX0K6g2VezyfXy3v/1MoNePPPXPy0lfhak
lOiGzPwX8d2wUWUiAAxLv4Ps0VgA4R0/kNRXw/DEe5b7esWD2Bna9OymEyZe+BKrFiQx/jt9OZTv
+wZZgG/lVQr8/d8P+4G9ROjGxbaHlayknnKfQBwfHgze9s4K8hotEePF44vr7P5IjCOddSd0D47J
aTDFS8D/OahGra6vSrCY1yWdfPnbOBVczv2P00tRmD4ZvRx4GE81lXdv0emQZ/tSIzomhR6Taexg
FshDlF5Xx4fXGpCrgAmr1iCgfY5hcTY9nIgt53fecuRtmAFyj9MM8Hmqg8y/hf26/LzQmtrn/9fb
5w1X+9u9+2rxvE3wfxP3kAHdByC7MIoo72d/kJ/ODt3U/bagm3T9dViAwzVvKQFd4818sgLtl5R2
zPHg6xYC90juPTzFubST8D2m1TQ28Fb2Rt6+N1Kfoe3Hr2V/oj60ABWz5Aon5mxJuNqh4EfZy+pi
kqHaO9C3WKzGPp94q2IJZeBIOLL1mxSE3CcsUqH7U87gmmQ2IFHKqp3rMHyo9/HWKrEclGrS0BVV
/TOYKznsBP5lDfjY0aQmTiP/6LU61jncoHsG3++pO9140kovaPmugx3HHFuj6rvLS31kacm8+pyv
Y4plhhQ17aMXewXMnv/6uI4enRjw9Ne/X/cB+1H1ERQPqOcFdaa3oU8BeIaPTID0TVxLUc+wM/GD
LOn8sNsnnyUOWxGp0wH9pt8MMg5Nnsb5vJ+oWvtbL3hr742XMdhNl6EbMY6pD6UBqsxNKD9ypOVy
/yGoqHhh6DQVP3DY6UJLYqQ3DwYRq3OHDGRIGkqZ17ZgeOoV0S55c0Bk5z08JoSxPe/wRYTCDYA7
Da8rvBYEZ1DSgzlHfu19eGbPPLIUJauWs6oWKLs6plEjHBuEviLMWP62rHAHXo8OKqNqGi3AbA6y
nVOJvw8q3oRZlAcXURL5SrPe79nbdctM/DQVySSRObE/OLt5qwB34eu7ieBYZT4Q/rZ1nPYH/zNH
g5nW9Jf4mPXkTUKmixbXq0W2y/0QgW/4X7OL7OVFg1IgwQFCCDD06kVhEsaCMLIS2Mt9U8cjv3ZA
VBV9pLuso8b8S2fIIIzjpgQzqJ0Sv5mb/oScTfds9dnjpCVyVxF3I4YFmHAxBvP8NSu6ElU6yEAN
WIbVtK4FqKvelLkNDSmTF2z1E8snrBHe/2L5uVF4LsplFPIzKjbPhfEFrwFkoyM562aZVcCTSGFm
3W8RFx+moNcLHKXgDzc1E30AU2LRHrGvj55ki8AY4JmWYJBQDJJn0Jr6ngLJ8f2SMq6lIGIjkAeR
el2oGEO508l4zV2fAsaNMkjbvQoTzXq8vvXbD008bjsg3c3MEsfrFpBUVtpPyBoCWTP1bXuJp0/m
LRbwcUtDb27lNo249sF4aCxFmhNbZpmJn+gYAffFn5+qe1UktFvCaWpJ1p4E8TyDuj9B+B7eWTfk
CJNuhmR5jXFYuJdc1OAXDh2//WFmm54j8kbba6b4IDnPrRh0XRL7KCo98KpARkszIeSY5WANN4UU
C9x2xVe6wqG0S7+EjCFrMlZu812Nt+2vkGPR56QZlVXYHo9vlXbSa6Z9s/Q0O5H/LdFO8hd7EbBe
JvvLMtlS8vYAH49t/d4KrKkXP7YPAXCdvZJTAo7LP2+X93UhMTtz3zMwrNWxT/pQ2rwvM/E+uv5+
TQ5nyoXnF/M2/US0zToVpyCLB/OthMr4N3UC/fR6N8O9QOkbE67y+Ld/gy7xzlUFwNhInS09UWkT
GjNjTsfJcZw44VrIfwE2LXYHoBYmh/PImoulxY4c+sgKHEduZSR+j9eLLGIQY9y7BKe4/1XLKmwl
RPn3metSsG1gn0StQCIbu/JTOPfqjEjO4ABLWj41xEkstdgYsBdGUUOV7yi5ZXOS9rHhhPCqf8C5
FjnMTIsYZevSQN1VZg8D5BdzsSAMOWgyMNMS9cRRdYZmGsZ5x027SM86OjUftkI1gPkRW8dTUOe7
6rBkgKxWNSziWgMiophwqux5DSwA1e8+7KE1NXvI+UCQwZsj6is4HGg+pGAfCewDy744dUTH8vGq
xNpYh/dZE+ljthcNyC/rHdEo4TuL6sljNp+YaUFGHmXRaPB/0mIVC6dI+QIvYDZSKyVv7SP+r3hc
rwbD6KjPJvMeadXwNytlfg1tl44QkcSfbJsJ++tHnRLGn0w7V9vd2q16yNkQ42S/e31nutbpEVOF
2USnXAjuSn9LPWv9LOWP6diOT0cHDFGTqkysMZjeAUGjyxLKpHl29Sa2utzlj40we5z1CtArWfYE
TUodBkCQiqK9RR/StKCk7JiEacCBmTFd//Z96iqZ/1tjkRo9A2ZXnp5bz9JmI6bBKWj/QotYhOy+
8GKrlC6E5Ug8YgqEUqVG79XWeGs2v8iddfQvaqwljN9WdlV9ofv1nMH3eQObO+/aJgE4Hc4IOgBK
PZywimNgoKZlTfqZGW8SlUPuKGqpVmx2VV9k0T5hTtqOsUDuhtXTDvVPdEhrkqOrZRi5AzGDa4It
SxMF7f+x3qBepomXh8nIv90EGFBOgMmT5UFhO5ej9ya/jQuvLTXhUmb0U3iPqLxLMbs88xuGgNZ7
+wn/1Kq6PhgtB7nJMAHdiupE0JK8Lo9sezLuCRtYYTTCVfApJA0OmyuPtHdBLXH9nhvNlD5vrepH
nYmYiJgvMNZGRXByAuaa9JVPrSCNpQY0lo6c2Eb5RwI2pOq4siQAQtEKgG7/YnUSlt0MiTBHu61q
Wz0BtzDpz7ra/OcazKtsuLXjKg8zQPERP2O1jwKAhq+wYls7efJsocVEehX5cCU3mBsUrInnqwum
l6a6eOO9DD+cdeh4bJApErdzY+ktol2cmORzCpacrOZs+JwV/OW5cYdWfCif+hRVK9OdQFnZwCGg
bnkjtA71n8MpGB308TXkoNSiHbWHr3qxLTS6H1BUAK2F/9hFEuJUiNm+dpYfVoY9p6D8tjvJSllv
lTdkFdrDzwF5Ss7eW98GdjRX65qtra+m7xhOx7fL/1k08502j82nI2pUARcRq5TSDaW43ERzFU5x
6zgQ4hirvH66EbZcvXaFQ5CbhgueA8D4Gc7OFsENqhmJUwr5F1NYXV6GGTwTahjZMPO0upRbNXvB
I5Pd1zNNIkHbL2wCMI9jtAsmb9k5tbvYGYD2JJnbh5o+j95rYWipVl52waEXynE91bHMr2gthcxR
1BhOtE8sRrJKIXe+P+M6Mk3BmsDMkkHxnUVf9SwlwlndIk+HaJ5+IesZBm7uIsR4Z5Lwssjpyv2r
o82qIh5UyyGpr200gN51UfbFdaWuYeDDS/o+buUjZt3XXy+FscLlmkVbhcA38F57yrs0TvfKGNWh
96h6+lMK1AosDt2kmGEP4tPzqq7/3JZ4qwFOQTCt1D0lA4lb4vNyR8YHac4BlTHaDzAvVKwKA27y
TuO5S/IKis3x0OExHg3Xgw8OBJN9BJWK0R1dDJobO4X9qthB7xcZlRRXHTLCNSjBCVfmOJEVbEJM
8jrHqcpWhXzDKW7Giy10phXckWsbDLegxKRcksAPZfv9IL/UDJpYxDuBjNKBHwdxGPcJIefcU2LI
1jb8qMQONy6jaPP9BaE/+9wKeKrcu9kaS/DnfwDh6QTF1y7a3w8NV9uZSLVofqszu5buTOUqARkm
VRnaPszWfn05Y90NUBXNnYkTxSF39gu5BwvfS/51duU2FtWOXpE8dDMYQAlLMbBP7kTMjmLtrUDw
/9D9hpgK6EvmGIY5tXxFKqRVrh9kbMP2cwzQbxNnD7IhAO0uJtkL5+H0sXAQu6/p+YTnpNzGyPT5
YnR0bwasAKwxovcAGL07Oq3sTnMtBf0YE4MXVDtZ7G37AA5YPzNRBLVdi9g3PRs8ue7oPsLhBvZN
npaLrL2PtAP1iN6SJJ4/YZLriQzTvRg+fAcaY2saC07C9n1QiKXGJtCUW393T1NUYg13cajTOq3l
Pjl+O9s9PErgUZyzKv8u45/eEmLEd7SLJnqtQY/9lrxw//4hMl4U/DxXQGa1kP0KqCoTqDLQqna6
HNkKIf3JWALqKsF3ZElI6y48DaXUs9Mjhz4sUgvejxG6DLXNRjGVBGCWItZ94LZcShgXqqbxs6j3
mjbkj7COQyx8EV2GVajDcBm0aPiimm2fFaI5c69N5PTI4z9bdFWH9D2q4lJD5JK50k+hUC3KtZ+q
uV/Wn1p5ndOE5DuVBL3Ue2lJvsF+Mjwpoccl4oXs1B4Dn4u3D8siOEfTFuoJ/REyrdKos9uQRsCu
0c38/0ubTYZ5p3rx9AfE7vlcQZyz37tZsjN9Em0R6xhoGQukJjDifxyD9jcK7Rv/t/penCe9lZCM
UV4TSZ9QLpDA0aBrdBYgI31Kqtc/pi7gHEbPC0T9sKR6WFEje1Vt8gXOB+2cgAitWplUUG6ymRbb
7h8+EwJtr3WjMPOsZ4uUGA+bJUrq01BQ7fWWpFMA41sD8khLTgJIyNUSFfnoQs8x4TTf0x5JfCPx
hhnM2Chy1IV0t9VEM6FdX/WFjEGfzrCk5fABVW0Jr9YRX/ohRPeT/xlulaqBXV3202Qxx7qvJFr/
Vj2CFejJpTm5uC8D60g61e6/eb35W4ieOq1kIg0KIX88NyaCs8N50Zk88lEaooX31jZxiy99RiIS
5NaTWKPbhZ1hXnvMqORRkc7sbsOA5xKpNV34AHMt9mCOCoDDZk0kxtYC2xHVTn4A1x1ImvFAG1Wo
7h6aaWbAzZR2m8vQrvVLlfnxnSnyvK9QKQBYKf/EtLPtRqQuXTspyq73aoKqTsw03XO4rBCrqNDd
7PtmvcpSNlnmJL3t80ZyTzSXnOayFt6rb1b/meNrkqpy1CTmvRdxwNfSSReBMCEG+NU/bkTa4/jJ
r95z8ZeSOKPznfnONvkPTGg8pTWN8rNrOnkF1K43rrW8w3ymOsNiSwONEwHUDzwIXVqbXw93or/b
5QlrEVYr1CShMs9IU4e+oFkaeQFnfQqQ7X5eC0+92i5C0Z8vhncOWS88o4y8IqRZftAemvJ7SRhT
lC2erL9Hpec3ht9DDsWD3F6vqPN+1JDeXz6rPz98CPSJWLvKxmQXlJkvFzJv7NWlM5VJ3RyoLsgp
9P6uzXIHri27/Ke0aJxfJaIgUjFUHHG2dijh2Y9KHBl2xjdD44DRe1s7tnGVavYoImG1N8JJdoGH
R4L80M381y7SPTHrIwHdgNigED5OV6DGhWDVXQuWxgVXpXiwehNor9SlhH4b6KzntyPEbhp0PAXZ
U4Il2Nz167c90qFAHilXnckEQfQhTmRYozrXhcQPk18S+AROMpvNgrS3QjOdr1GNNmcJVPDpmsJN
12VUvqyomiOO+dA7ao0Hc3UpbNaEJJS7ADG7oc+A48NnI6hLQilUaDgIz2imsRQjdjykOstOStkS
Jmb0mxaPWSJ5W3hxK6PyF0Lc/g5I0UlPmBXrMQQ6eGelBFwCYPbZF8o2JD5YPuA/YlKymNXihuYE
fz/vDNtWx9/j4sqwF7N7FPd1eBQsnlp19PkcGZE2qCAHlueQYAy8hofqhTbVp1Sct6qCEAs6ioL8
qJEtogURZycAQBmQcNqMN41I1Ck4GS1PhWu6VM4lCHayxWspQd77qKJeSNA/SAVLnifuyZXo2HOn
CcrRy05tg8vBLz1NYxCMccac4HbeGoXG+wK3TWBJvZiIgjPmfLMXdlTw/QHKJZ2g15R8TAUq+4to
1scFpL9vmzVVPy8P2GmIoOAt5h/0pZ8vSIimqMIN4/d5QrCIhQNuzOYr7OVTbvw31IZ4CwJe+wAd
MihPmU4hDrR4hmyRV9V78IMwU0kaspG2VBXtQqBNfN3ZYt9H+lv/wAf2mTbQJ9iW9LZ1gSeTbUeW
U4lnsrYLn0f1kd7nPAPJBafZoA3mH/fS38/psebT8/tpxOree1ntuMJOdDkI6PVQi9e0E1+dVLxR
SARX567yKlrohNJ9X6CXsdLCo4/9fZhr8O6eccoBF5FR5pevGMumnTl0ucR0X9VQRY8OrBLR0TII
yaTn2d+/wRpkN3qBuVliCLU8a4pj7iCwlEG9nbjzaPtnIrmD5Gy3pT6ki5z4ip7NnZJ72qqKpeG8
TGCNKQdjsQ0j4JUZg0oyPABKhYtgjDqcf+ytrhCs/ORtLnHY48wy1sToDoBWLNCuBp3vz0ZBONOh
0CvqfHKoE0krkFFHJb6FK9VCfk2yb7nd6reoaQ+VmYp8Y+AQutKy14VGyhLwf/YolGXxvn7IcU6Y
bsmTRnr3bpwyDwTF1XZHqa46HSRV9xzHej9sstguhRM1FE62eAWN94+3lp6GA53pSuXeHq51GOG2
tOrd1uzWMUZUzINfnKuqkXXClkPYippXN2ncbbSWBeQAPTSknF+XP9ytKiO8e6GfgjEunWsbPtu4
NMe4eEfxqszinPsMhj8qbwG0scdt5FNBae7kYmfaHXKWuMxkMQ9MzFlX4gLvnpG+ugCQHqDdlBXu
9WrOxDLrLaiuU2ZczCCsidzSPzLJMXrd4XJfmcMaaPDAD5jVWyIw6nJ2Qogtrbk1za1Sy5w85kcz
E4nDb8M2pQ0O8mDz2BOfdtWOGXr1oQ/p2l+OzxrQAyfRtwWIzSqo5eJTUnKneXsvcNeuchwA8wB1
Lh3OvGUyiMVfr046OcQ3Q58zgM0mwIc92aMU040By71wPey+nGC9TNzBwE1y2S80tp5+Q3pKtgVT
kIp1WgQ6Iv8EwcrM25eWqK/fhqiiLrOJMPpFGRHViveBM+A65Bm8/w46eDVcWNzNeQYhmsJOKXVi
KUWwDisI++mIdVXCj+iDkMvwm7cz0IW3EkPbUu9HBYwOzTCtY7AanLcTmvk4Yr5E3IaIiYjl8oS1
8aLt2u3QhV9vxt6cBXpVf+H1bcS76WGjHuSvcn61oOquZgX4YX3776xYB7tJPLc7BRgHqUKBhVgu
CpJVrB5kWn6XNLTj2hJ5BRGlGxuzZDkBlh7as4LswnYrwbJwvrLVqefGoOhkaHP2w/dOQ4/ywf2W
qPRMXBlvB4T2wz76W7Jw2jORsJphjl3nAlxRd5sqo1jjXMtzrG6dFQp6SqkNumQR7Mfh/bjXcVJ4
9xiZm5oekKGIoQnIfBSxi2snUhKyodMjtqiSoMUfRxrqaFDjlZckStPlD5ksUa3f70FnnoCxuXCh
U0NzWqTrhH6DMltm5ZWfHPvKGgpuPrbmWXOisWwOFVHwQfSqp7AVKCazWjF1SZXu0/YI26HSO0z0
+aCsKh34fyRStlb8I7GN/+HjpKBKkN43ebjCEscFMl7pbYz0DHFAm8i6YGJJ19eRxxLsh9Sb3tN9
z0wchVsOTfb7kimAUh/Ldqn/n63mNc3y4sBS5HbbxI0dw3hcQV9B55iyzJFzw103Jj0Ao+JbDlaO
gXwOCeBzlFiNpSteGae3WxiUJpr+VP+w3WoyhUfzM78WDPUhrBI4chg6knaCFwulsLYb82P05VS6
GLW/v7WKkzkXHqTB3cYbFYUVk7iBP92MEnHe8eNJGCk50JLmRYffDsbtDZplHfLuceibxcC5Nsva
ujEPwc2pb3uENMcdiqiMWPRiblHTFj6n5GETPgSTR4HrZXuoMvfOSSThmWnpkJ0i+sga6CkNM7h+
lJkI1s0Wd3FtqLTjm+W6R6mVJ7wFcY6X+oWL9DMhHP4E/i74d1zCLHGC/CXwvxMCCtzKNg5aRBOK
nTwfAmkclSSzoa/7Mnel55wzvI+Evm/plzxsqn9fTGulAPvNiWblx6QDpIf9OqPEOdNqTo4bPZyB
6Vl0G2ZTzIv/lNdgVxPH9z+M27KWCO242XWTcy6yMczNdDVadIvJFXsV/ZBc2KlC1+njQKpNjDuv
V72wteP933XDWmOnFUhx6nLVdE1cNz175wb3qdZt1sft8cMYObyOvt7DdXcMOVW/TQMVQWB16osG
byhLrJr4JajZ+kPFZwzyhWYElFW2gQhmB6eFK9d2MeXh7XdR0cbGHu/t2QZlI+ntGLohw2rFHM+K
45hLPtl0FNEzEZQtQqZ2IGB0yKxI3i2K1bjSigL1r/PgbbbTGErqoVR9tqKwy3dP8A2omfemmadX
yAjwQYUuroc6KemWvbzzVcuzCikauprlZbUw8lfWiS5wBkqR5pOmV4UaWK+pYSi+CV0aQ4sjpNFe
rM6L0IGNzXRRXnPQNZLjpBR2r03RoxpQwe/nZZR9a5i/PN/aJ2ZcOs+mFSBo0iyrbXQ2PHf2QfrS
Gu3nnPlLBvZRJ43YfA9/Cg6HX+cm06OePXz3bnAPKY4+BQdOIV7i8Mx+EqWwIFpXZ7/VKJlkPuND
hKx39VLVStnvdjKjmeFrF8xx7alq76lFRBk1uyOUBYZCML/ooCz2PKizXyuhy1jFznYI2VBUhmFB
dPk1VKY7ypX5gUPePI7Ni/9oJgMMSiEj6oYiRCnNeADy9d+qnVfPhQb03Zz8OFVdR8M1m2m9GAIy
Xhfwgg9M3cyyMz4AhxyGZHSX3zvtVcve9x6nNJMMQEzvsCs0srClLTbM0Gf0f6Sf+PSodeE3+eLj
zAS/5Bl8B63AA+o659MsFYQckYVbBXrgNJDcSCXPkwjrcZRjqUqkQakpmIFKKiMLYBarLGjq6RTg
1vN64JHg54T8z47BNHHgwISKizGyDWFPKtSgHomfIKE7sjaXBZADOZEVDNPmg6vZ5c2TzuKt/v+S
bpkYeuzFLtyTpOoSoVf7Jf4q6TkcSyWoG2hKkrvX0KsPA+jJlirF/liO3KelD4sKobq9iZP+TIrL
3gSsHgNwbQT+zBBroGpvOcdBv1278SaVncqX3Y0TF3VLb5h0JgJwlrpBIP3bR6QxGl3K/zu1sGuT
IUY1fx62gfxRMb2T5v2HQfG5trDHYGv9KTF6G+GFEwN/sb7Q8yXlCuBLeFcAUwQzcCAJudWZqXFT
0FPRZmB8KMrfQ/MHHbCaPAyW6CdhwlxtQbOWSbyfV5tg0z3AnBAkLLt/GuGJz+GydFGJyYzzF3UA
e2V07XofkjtCYeKprGEkAsz4T8PJuK93b6ekM6XllSbi8d3BnHZJPc40KE0GzJpHDIe+bs500lEL
OqpwbG4auk0JXOT5e2AuCkfiKCauY7CgSGXfjlHdRAm+LNNxNFuCrHg3oq9w9xu8hroaMAx6SU3i
hAcitk0NnVAvhSBGtISKbsDwEcdl+Ww+kLqZ65u0X8fUxJsaEcecVl462Igu73md+by1IATrUnY5
tdLdelkfPDolaB1LSYZ/531MnG7MXQGNOjTUAu/FFKujhCjMdVWAAGl2LQr0COtfg7srjIVExeA7
LRs1wYFfiRf6vh5Njag9ENr8bfn34x33R4vErhY78Dx0MpmybdiUNouZUOL0Sw9YEBkRh24o/i38
43pP0H4qyd574Cdwsss8JkJw4eym9fJ7HN1BHkMVAPf+SO8LXhFFruiqC1iDqfhrerksTCmnhFVx
h+jui2Iw4LU3s0teSjLuPOdWvHi4LF5q9FHIOVrVGZw6wvHsL2aD4pg1lqG5fNPuBy6CVIhZvvw7
gjTMxUtZQBp6k1N8P6DtSbEsaikFUEL4RRNaNpwYt8UQfH3DxQthBVb8rMsHiq2jWR2BDJxI56Ch
R6NYEqgtf70GlJuuGYnLgGPzp9pbWb3x9tPEbEgrBvhYywVE+/1p5oVi8Jl8pHmi2gaWvbATee/w
O9gY1Gq/08G7qTbGz5yQbVpiyfzwAS1SF/S9bv1JI02htYU5FtJsSV/cDghTcMGI4/6wkbviXA6Y
tsgL/r45mCX+vHgHoFdPPuKz6THip71iL35c6H/ywL/zmN6fo2IAGc/U3/NyRyFHNttJUAaTSYMq
bXTmR/1uEmpQqyNPGeokwNUlxdH17LFBRt5FqFucG2G7El0JIUQFBQC74e8x9UnJGYnRRW9eg8AX
Wudi1WdaPiiGgT2Dz0PvX8cfqtPsRHtiLV/qcCMaRiovwpBZjKr9HvqvRebcK1dxt066isx0dKqE
XvgTkndZL7rjk6UScCzf0VPzouvUJcGTu+A1/j2J5Iow9eos6INgFeMeJyQX4Ts5uuzEkinHXp0d
Rr7RKiKJoe/AQSo9OfwA4n4rVSAAQMJwm3gIiN++nEUaTS2k81/n1FUx7dqKKkHGypX5zu4ruime
JxnlXvSY+x8mb2L1MDns7MXsobQDjxWn/ZhKFSrrtWk8dgCqHr/3OlMFm5zD7JTdD5V/paGVaLrh
TeWsKHGl1fSmvqKX5YkLs7YOCU48VMMq+0D7BofJ6ezwXDfYISjQzm4WF7ACLZIcILAc+u/wSh3v
EvNl8QuuH8RKOSjfYcCNM8rEm1rQv+WFecp/JZWvtXjcGok9cgWz2V8pwOBqZ2T2eQXASG3TUGhS
Wk0TZfnxzNnV7p5J2yq2xEzze8OEuWVtffJWUquASIkxvTXMa1Wul7etZ19hz36/mYJXQ5WvLp4k
n2eNzArIIWTT2MyHbSS2h9KtBpeWIQSTfAYGV+BU2XkZvhcK81V7QP0C4lQQ+M/YcsxfLCQ4xhbK
9rbjU4tBZUe8W/SPghckcXIi+wSIFWxmDPhmx4A+TuzNOXlNwOjGJuhmR+9bM87kpoJBjWFl73TK
h5D19r3IqtRSKMJU0BnWs1SoZEIQPIvgrCP5AVhEJKU7fqUJ1sa97J4mLHp++repDSmxqggpVi45
JR24E2kka5i9ztLC28CTjFfkMvov904A4cGBllTW77EV1lpaZBPD+X6D1h1tWPJDK+VCVaAvHc/D
KIquWiHI5tHy8SPKO/aj11bfHug3jMdO77hLXXGeh/AeSqUGUkAY925LYlsEtbNDFOeMaWU9UrAV
/CW2abvmfCj7BrAIXz/xh/EsttJJbXw153k8y8/GFjknsITzLm471v1J+gHqELgvcnn28YCSGVO1
mwnxmEtsEjLq9tCYRr1LJXPBwxJoclBiFBzI5p32ALppR8SiLsJXi5KAUVkOdKuMbK3xSAlZdpay
3XMfAVlV6IVdCmPXQotN+yVVjdq4lLJnXX9lQypZ/0KUxaYGKroXe65GKYL4xLzgDObS1J8/GfY7
Kcv2i/qngE+F4ALyEm2ZhHaUDjFSUsunxHey1jtare0Cm7cZw1bukc4YO1Pd0zQZ2G7WjPWHQ868
yTjP1oL5vNCvVtrc9IC08gvNNCV9vDMtQS1LWZPozk3vXFDg3iXs2tw1bdmVg0fEusAkEymehbuw
TRqadDTQPn/jbevsnUcxenh8L20fcpIMOgb1I8Fd5yH2puR5UCYPQRS8IMhk1a9GYbZfWnAa1cjK
Z/q2WokN+cW49iJ3kA/gjbf3thFR5pFLIsgiABTWFmFFsFhRV2n5zhr+1KDpg+4fSQXiOFd53bQo
FAqullVRUxzi2ra8HJCOGlaTF+UcPIi1hVA2FpwdLlmjKoxPFAB+oeI4RNn2/ji+H7uzV2QjKVoL
AEQ4XOrmIQE0yv3N3F7A3swDZqeYEZoUg0DOeq1PjXyoEFel6bYO6ZkNpQDmC43Xv1ivb5joTvEi
oNISamv5TcznVeLnI+luBSH41933+8gLk0MNnPsZL1k1/cdKpxBjANxo/hZo6opb2q3OjfFzuOGS
xGmn5j1M4JXp8NriwBRTmQcZklJMxSupfm3NkrXDam2fvaooDoIFOtaIJJPSgxV0IOvExEaBLKGc
WrnIMjbpQ9kunSg4/n7YS8s0lHWSu6stQ708dXK91bMBORfZgq8yR7lE0gVKL8iI3Fx1/u4gDArm
b9OuHfaUwzyAbWwrrEvLJR7Y/V0aLaEQzAf+0xkLLXQs+v+L/TOKdBnS2T+dOJvkIjyE47kxQS4u
gxnen/HwtmTOUsLrNfWWmQ4dIk+t7ynEkLScKT37CAYYO24JhPc/QbZlZwYxdaOozVlK4dkO9n3h
12XxcIadG9khuVOVO0DEnuJs/RTfnpKa+3ZU7vZKYgiKmtyu3Gt/oE+NcVBNBwqBAetZuqeIdEBa
KHOciF+TO42KcjUVTBGHUwse3p6z++DUcDtJCQ9yzpnsWvoemLZVJ1JNi6tSEQANn1kVYf0W80lJ
yl3cCOrhpuceP1Bz62i30vY4kzGTXbWzdptE6q8w7b0MQbCtDH5MSpyrgroJBWhYostNSxbrgJsM
Qc0s4sLgKJoCkJIVgEDYxjozPQaKhDqd9fdxTBOaAhZK0uXo2hx/OYUiUkyiOT826bMbHHczycj3
7DUcnXkvL+QduGuHBq9mR+9oNS1wcZCZBvX9/tWB3l4pbq5XrgUL1pIx0xBxTUzrajxvV5hXoBmC
NqFXYKYXVe0yg/UY6GgLrCEzyyhUdpOFFDySexNgvzOKTaJPkZ7uAhs5TZqQMYagvvk3GDJd4QHE
8cNWgAyN100/cNaB+DuS0TQU1yC/kawg31D0PymjQAzYeMQVZy6Q1l0vlvbu983/CkEINz0jT3sr
hOvsKSS1RSahcBRiR+qdG6TXTh0BjIrqKl/GA992c3TKFbNBhE6adCBsEtaDfOIIjl/3cG7HVGyF
WrGa0XbHtb2ywZaas1Nsjzm72lXDZVOWdv/lel6EEEytYzkSMno5p2QVmNbBXiel8pNoOjHohZxK
Xcaq56pyHVD8fQ3nY+KjY5ENRuYwgn8U57m4n24R1Xs3RxS7Fp3koQR4U9oyWF/GZPM2BFO7jh+5
YTbVgvmkazlLw/GMfCBIec65Od1Ec8wg9vjvuFhO7U4HI/cpA/iKXL9u8aM3CJ3G5nS/p12COV/D
oVftQ9VJV+pYGl5iu5dFkxMLDrPxKcCttVRxs8f71OgoQxr0D3KNh8ED4/b/+ipqE0IuzqDY65AU
Gbxn3EVc9Zolf+ISQMuDEA3jYePPKAMaD8nb2JYNbqcX6oHkwc2or1UtVPhzq/Y28mqyHG0cP5vK
DJ65iZFc6gN9uXkVGG4P8gl7xu3WakC6DSVoUApbQzQYVELe0WY0hDvS4Y3PX01LP024BiypELjr
GUcxxuo5iGkaZ00xgYbgtTs5pZyknvDgav3oLlcLcAkeCkWShdKLxIGXNMR1+ktgPIViFCeBb9HV
Gik2uQw2kG6iiAgOBuvBhmVMiqACV+1ncycEeesTGJyF6fVsjtQjjoH3bJd6sgbLIFjwmhWJNy5U
mMsGnrVe+fo8WJacZnkeWIXSRBC018022vPLjPo3AAW8h2ZboqFz5b/gI1xVTPr+59d7hWYAdanM
SfRhd1Cc1cJLeNgwdSzU2geYAzrVER60ZHc43fOGaU7FiqlWlln2d+bRj88xT6a4WIdR2NBColeV
QwjUfLaQ4N7J3vsVzOiBJBAUPaspE0r+jBCF0RiBwVOorMiqWBk1Bk9j/cZ2vGeeBel6sDqe+7lL
VXFdPBZuCCESDKN+W1A1cAiAnVNtWiAHYLMjsF65MUFR6HvZc6x40mjmcgEQoFLTIfD1f0OldYvX
gq9uLB/+TlsEUKbgTpJlKds7mV6ZNV0TBv+PMczbC+ttFBkLlVoZGV4i6l67A+jdE+wTKd9Prm8G
HKIyzF54u3BAi6c3KHCSXCvlS+rkArznchBXgplE+5wwn02ujmXdnERkni1muPlPRVfv320KXum2
Sp1lN+pYdL6H7WJzeJwf7/rx4N1qExk+uUu4/J/YtCutrYockITYxL5H/nINDd31LEl3ZLN66vGg
5bgxTi9njVnRlsan6fVQWTJRg/+sR/WyNfvxsCyNd2mCWA83lnjcy1e2qvrL7hGaqrKpWoadB7re
E1bQyHGE7GSYLSA5IsuLm7YMVdP2Ekj6POBC5eUoF3mn810jYBH1YrskZtW8I3nIaOP66qjWYTKq
lk/6OqoIoBVVSrA3OkIO1KRBHLTZQBaklsY9rR+VOAxG86Xeg+GCFMxYWsSz/8d6OfyaQNwMuhEM
APLDeFyTydD8slfm7TnKJCN2PVt2IsIo15vIebcGnotZsH0sulcbOm19CUjohsP9gvNtsLfvo06s
YLtjv3Y6r5VgUvwhzFwolxmRF5PXc7O2KTOOCRTVUqpAhxIj3BdBl602MFR/Kg3DdyMZQR2fXgOQ
8A9vR9RTpe8t7gB+hZEZMqaSequlMldyPwUJsPCVbs/K3sZNhQDDTQ/+jQfXAZP1KCtJjMuozN0/
7k+YnxV+62dRspGqs/e3TE+89B8BC9hCH8D5rPgsDXniQNFaysTfcqcFKgHpD+IP42yeXDvHs+Xr
CSfRF3VaiiJE65RUmpA6t+nKY5T9WdzB+DEiMH+lcVjN71wKJYJyeas8xR3Tgiyu1C0Vn45RDHca
kyeKzM8F1X2PSvQMlb8TNX1YB7wgKKuqEH/iGN3bLUg527V8IKeJvYQ8eSzvqpPxEIH9Eg7ch9jR
6g1V1tx0N0EVRncW2FoyJhegqyh5feywvv/IyI//0YGOged2XtsEqEbJa5JvtU1Zr/7XfdPyylOb
YBWiaJ059OtJVH26Ddi0k0h4EZNHdIXlUHKzIUnS/FKX6IVgKsLVRvm/KAjpMiqvJXzxkbQB0Udb
kVE339EP18LHnHiSKdNRG+Aws3QOF1aqurdk0msl+rOesEP5eO45eAxVxCbKnQMlq3iwWcac5jfA
3Nh/t78XZwzlBBdqvZFWVMzEcBvPTpGT5ZXMeBFcBjKU14WUaI4GCG8iApDGniLYCnij/K4KUIx6
oQ7Mnoml8MhDpk5GbpgOFRTsP1xkOtWpGuFEVLgrtL08DC38xd1kanGwsXtSg8fWRavTzmcI/j5W
1aGSeVMyA7BrgTsqdPdctVOTcYTaRdVougR+byJhk4cGjNyoBTD+rghKaIFbBLUXXRwGxIUZ7Dzg
zmsyQShOhavH0XcygcuJhgF0sDMWOW+4E79yGAegMpEXwIPpPNVFSToDtRC4PdERX/mNeqkvNCqb
/LlfN26EOgfWkMfRkJEOYXA32Q/2nbwAQkT8LY83AvnVByopWBAGhiivoccO9UAOIgzTEegNLyAB
+Gd5KKntTrDvYTvXiBgBDKB5bLiMz5lOaiIyqnJ8heRqRghmd1EYkeMy8UZYSsmy5+ukcucbDRRa
4IXKHmI4/0w6XWybiPwlMhsVyfBx8/4aMHverHgIbXHFhK/ubIxR9J33+yiDM+G+S2lkoKSi46yd
0ABJbaguArf71ow47dDJofbJOejb+/LUwiH7IfnsiegAtqwlQgDiVLHy+iW6Kfe3idnrI/ILgTgz
vaiCzuH5AyyxhBeTvgDe1JPwoPGjmbiWiRswOKPKqhn/ZuhU0TXyAy5zNVgqIxRjGi/KMZFrYOwP
bOwMj99zE+smfDOlk22kvjuQAQuTUhZESiIQpizlIs/exgh6sW6cQbSXUxnHCffUSqoZTOQpNYAc
XKAOM4onjBMIPIabvxCFwzUxMYFZCoYMLOufPVZMcIs6NciKV4l32c207v+HeuC5JNJZ2SBhF5KI
yj+fqKRX479F40GWxgPZdUmiZmiOdIUxmyUOKaznDCwKuaZN0d5Zg67QTCqpwQiRvBMmTdgi6VNS
O7ZuGRrxfdblpIsoshrX15i807UJ1z2TI9Nxf8yM8GG+QrQ4cNvzL0J6BOwgXnbokPBnxCFx/AJ2
LQKH+lr5gscuXE62lGxKkBU8o9i7v3QpoKg119ENLmdHCnd726QCFFEdZU1etJgcwS8JOUOWHmMs
HKnxq5SwsW/n7xwfl/CJGMabJk66LgKpWtatRgFxHbnvJE3eREikHJ5BYcfrpe4w3uqX5keehktr
6qXXixrDF2+ofDdl5/s5LhMZUEGt4FY+WJ+9FF0Z+xaAuC/kAuI5l82fYA2sLIrPbRoJd1jUJE8F
JolsLIQNyoqfIIyVEPOaHQHEd77/lyTUx460rF6vKfP+9jy+0t92joqDIcJNm5IPfGqYKZQLF4A2
D0VmRLXW38qgvJAIqRh6YURMZd/fJYnlghhmB4FDczhKnCKZeOO+oqHZeHdjmiIIxO8JKks1hKxC
A4tPF1EgNzCCsuxuUdBGJoclLQhDd/wTgenB6UCGngpkX5WcF9J1DiMSwFpD8gIXGXlhXfIT3go2
WinX6oq+NGThWy9m/wjJgkFDXtE2bI0AyfQlF/Y4i4+s8f7fbtfPbKQSFJHwRtzotjlmUNOqBb2J
yIejCtgCcfxd5CjN0eHF1GEI0gtcIqcpO4nK0iOMRc5oc4damVp0mEDmN98hCU/Q/x4lmN7DkyUQ
4sKKsaCCmc50YjbGSPRsHxRff6fMQ3uCXHtYexpMJ3FDJ3r48I/o9Rtws5u3xoFLinnyHRPjXzAe
Sq5PRWkLBlNWeoP71OIQb8P5HEEeI9beXtFdx+kZ4OnaWXAyR/3qHaYy4XkS05J4o3+TSWmgqYbl
XcFRHJ4ZocbnbXc3roc5VO1BHaqVJdKpFiJL2VOg042XvvNcvYgaEneVho3s0X870LHKq2R3CfGY
bgRN5jW9E5Yc29SvauBIlyepU3B3sSeSM+1EKlyrj4l1wHT9UVPYQ9oRk98eFQlqoVa3AQdMGGRV
RSPIUuZ8TqgOALz2Wy174TmbKX5KnNRDdEdqc24YVpDrdMpnH2dF6hikLbt6oszOnuOlwl09Ys2V
isK5IDMdATSJ9TjPt93K0R2mqBPz+lYKQNEYwki4+7IVIyiUbp+mAGA8dPpsuPqfKJBM9m9JOVgf
en1ec30vEF8rV/n6/K6NsG3e1o1rvJce9emZ+oDouxDkAE7b2CaTUFSc0Tq2mBCD+3fhvAVyiquq
j/7s1RYABGkzMEHmK6AHVXwcjY1jepmV1cpFvb2mbnbxEU8wCIkclApQt37hhXkknHy6luO+U3Np
9DcQhj+N/cHWu2nuYqCxIFNaTwqHFIIOHk+/DfYRfSn/KuL16Y3Vm1IYSAPksPt78uF9aGfwPZIS
cL26T8wYRf3feXqrRPpBHnwfhDRbgb3zBrkwnJ0qXUXl7NbvyZRi6ddShn0hf+X9Qhe7Z6xsId3n
Oxj3meJgly8ip2jXr5M7EPjxj6MGpp/oKfpXp6aM8KB09zheKYJN+ZvV/E+xW/ASiI60e72H6sH5
wwCALHfliyAEmjiTd2iSW8sKLtYYWX+oGUEqM0UnUclyxF6bDZsZwbEZmfkd7qWXUuKLLEAFN1aC
d4LaQP3iMlkR+jX5RtTy2hPHHMTGGwOOYW5TsCHNgarT7bJOfRWGBXmB0uDuUTw7u1g5d0vUECuP
qFDMQAz06/EGxiYOukyDM80ul8+zxz03JNuTOYFrRl7i1aDloPUTuBoRzcyZUDKqfAtQLLEM1/Lq
LFL6bO9w8lJzGkiglOpTRZy+n0vEzd8WADtK1e996qdwPLDFUiFZK9ritLuXmh2JxpJDhxzkdzv0
5S7lUS85gy8Kc/BQ1wPwB5VdtZSxcidpsM6TZ1srGFgKUMlWAzpAIYRkTIGVCviejjaHapRqkMwq
ded2bh16Y2VYbUoNK8Ir924QNNDjlQlTwWMRc2QDQvEXaMk+62CvOCT3ow5tfwu+rRklYOG5Z25d
qAJd/S4DKLmaXkV5fCLFB+NQgpRbEWyFKJfvxHtyH+6INDV1fj+p/nVzrjIez3ROrhLsb+h1PNlX
0V62tJMuN/Bm2EY9uocF9PAz/WZra05A12qwYR2oB+sYJAuvf22V12ev1OjUWDFVrErSZ1B1Qd5D
IzvzjFdOcDuOomRE+JHPh5TtpHnn9Sf0V1JdB8GUkz0aGQCkyMMuXSVSZW/DBnrl0NJ5+6MmQ7D1
RyJ4a40PvTPIfTIjzxPuXgOMFA44u3zhN7NOpK0QFhnjQfB9rUlCqdPShGwU48PXVNYOZBPCYEPh
6OX24VsoL82OqXIwZXTzy8o40KbBMincdbOXDFkJz7CpZXUanFf9uGx8lYrrELzUaG3iSucEQ6Mu
UlXEbxrXsfp80SmK32t7KCQ362D+ZoImfRuLwdtZC/gsfPm3r4QdHObjmCKtbW3WCa476RqmOwov
Aom/Vfy8ka0z0qovBYLQBJrIvQ2SkClgKrjSK87nj3IP+Sq8fDv6kmI0iao7L5YHZ12tPIR6D/SZ
zqilvPJ+qsQ1HWczkD69mtq+N4NB/62rncd0K0mRGGGnVAme2BBBzsUZJi39UFH8Y4Hun8R9kcD/
gfM4i6FIeG53LpQlpwU6FJT4DTsUmahCM0qeF12QksT7G+JiAQt8pOgdAuIw2a7n9cXKMh7NKGEc
+JhVq1x5pBpPRoQfZLZPly/0sEI+eFinL3abYgfmoObXdr3xha69ddwRFJYzORMbzzuN6xC95LTu
hQISSKSo6S9SQZaT6dQLDWvj9QvP8v71eJB6ktcrkAaZ9iqqS4nkJm3jYsov6OGiVQjRxUKnJKv3
pO+2K8DU+ncL5m3GHsv9sKvho9wJBYhDDSVhP9iix7HD6EHhCkrSmqgnz8SsZRo6b6S4svm4yrld
OENNVxe9IxsN0mDutgGZThIBNAA/UA/iIc1+3PUsn9wZJ/WV/e1xqE0GjUrgM7QtXSsywwzuc3j4
UU27080v9Ho1j06rbdH8PCsSNbelDm+fyx4rqHPWGkVFhs3o/HFFYsGnNbD1UYEQmh8GyiZIO7yC
TGILvq2GnfP3M2KFSSxUfmO9V6Wp31oGAELmpqXKjXYvUzyheBEwetbeHa3K1/pG8utguPG5GAPU
sz2p/O8SLTl0HsjJbTmRvb7pnMipz3ZhJK2wqkFRfPHN9ngL44SgSdLAhK14fAnFWDxk0YIeMySz
gasZs3L7ly6r+bY6z+f0t0lx7puBUJT5So0dcvsbdXtCiwHrNwJNbXNZSjNGOo07msi+D5BKwGJU
h45GGodzSv1BvJwL8hBnTkVCFH8vsKQyeQzpDhVun0tFslmXoPyVOeu2fkBrSDobT2K1TXjsp4t7
uFcRa79LmZdNWdilFuhfRO72QLIFetinE0xuifyvYPiAo0b0eFcPL7qMXoteDwdoMhdtWMkF3gLz
ocwp7a+qOW1uBCVWr+ic4ljVs88DdMSdlu/Yl1ZHHndbo5yAs4evVswDB56Hq7OqXgAN9H+FRh+m
fPN7kTiZG3PYiYP1IsotxHbqfXcL5EuvEuwxH2LWkIpQ6Htxtpnt3xCN9fQxb8GF36VhVdiH6Ubk
UdbUn5l5WBfbjErD3Om+dfsHIgPINgcpQ7oaXTYcPVg1IEkRW5EER498sWYfn2zwXrOilxkLPc+6
kmjD3zpY4RkjvVoD7h0ZkprLEYZWHdDt61oKfkFoETAeXx4UrNxiajReUmO2iqv44pRBjuO2g8lr
RJwRzpdcP+YhQiNBgRQOS9zTa/8N2jcgbCGUIlJdJa8BdBipQmLQCp4nQ8VHJyCv6XjcptlowXth
FAiQWM1yPLpQfNB2/YHy3rOsNTbSjxmnBo2nYkokJ2S0x0nm7hr0ftP3+FhJS+aLNdpVYDJKhwuc
bo3Hr70VUvgaRPJQ7wdXxpeYDcF2x+LvUWHwFHqL5wcxYhjzrM9oPAYK2C8u/ViLanczY8VNn1t7
Y5X/9+ZRQIKLZXiZcf8rl8iYHMt0qForXzMAF5MDXTWBXkEl8QthQdCdpZY7nVcwjn44MmYzn+Mm
6qjNF2Dm7nslCCxXqpoCIR8AYncHCHnsh6RwvAnXWv0f2oqkrAJSg8sjppEsWSylDnfpQYAx9l8E
WLHyyTLHzZJxGZH+TZbnGbCO/A+22excT9iHKIl3Yr4fXy0hDh8/CQ3fH3oEtPI2YKLBmLze6i4w
nWF6p/tJaLS3G5XiJfz7dHuoL29CjNhSUOVP4J/qerUGj2qX/YrEgni5MKvkR86c8NI4OVZ3Sqap
0dDM9I71SJA16kN1TqJ53y5MSs2PWb5N4sJHGy9V3hZKenOObBCVtfZr0MPRatCFASax48viMrX/
/uP++mEtY9XnqyVSJDITft7PwuqtzE4Gj+PEyFyyHjI1OhIlO7Ii3j6qSJ+Fs59CIHVoioNMv4jx
lrW8iL6Ch4+elqwxhTOjQ+pvFuZPic1qxVDrq3dmdzH0R9EXi/BL0wZY8q+Nz5337E50vHcV7RyK
SvHm3Yqw0MxhqIyJpKsQ5yFfSjrMAGQVgKzhgijilQtvWDfTXzUJnGpbzfrv0jYqHrYSWIZsCUXL
kxrBXu0i+ZhuOmgY5SqExZdZWi4fr2a2TA35QC0OCyJQKD77giXiLvOKnGrF/dNnxD6wuJuk9nRw
N9mdD6uS6eRVXppTuDT5byzy1nyj7KCpq7MFOz/k/aENL4sRMrIv4y6thWUSX1hmnWkhvD62Xt+i
uJW70khsv/fO+xhBt2uTtOeEQ5aWB4PXK3372Ybq8VzozIT2qQT7XclyHQH7jtoII/bnZQAL3pES
RzPS1c1/xS0HuKsy2TByn6N/P2CY+6yO1kNiKoMqYgvTh61abOL2N9YOuJrdJl/qg5PljbTsI6IF
q1A5zK8BXoZ9QjWkgOjblEs7bVtxApElW9CFx/Ki1ESWEovWOHysYTXxUAHhJCqsS4UVPbSR4CVX
1ObimCozBcf5moHNoN1C1VrQFsUO/VQuKYS/YDfbwttyaJXjVFgBTDn5Au6Z1M7WcKCLoH8nak86
oeIzxNiDcQQO7jcfFFiPrNSjIvtS1DIMI7NfzzpLeOaj/O/wRlQscEGsmjM52xstN0iBIbmeQBlr
khIajynmWnZdm1TYSC4D7vkqsEp4HRpaPVPH9lOe4yblYJKC2pA18B6tfzzDHFl1jbX2noF+A28x
wx7LZgmymL52ueecc3iLlTL0S/wgKhNCWqUBjU7ZDqh8nDJ5KXqM3tjRhBfz0LEDgDkebcbXgs7x
HWC22rF+24iiMLXf7wMBZx/3I3bYyNp1cAi/737ecNV1wmJg9zy5bU1rW9wo4W5qhYY0NGBt7Ii6
ZvogI1VT0fhx5Ef0PkApMNXFy+oBaUaLDRcMSxEaMs47NrPvO73jcFI13SkDTEZwGUaWYh8OY0CO
02utc/yQDr5QskvStHYRy8RaVW9ggSojkC0bLNKd5vf3vwVPk8HrN4v3temlIbutg0BvhcYZUe9z
wUDPgFCsJZEp0+ol3mp2avEnL6zrW3k37rTS/B+MFaTeGrueH+HEHLO9ysfMafsxXNYwbu5OBqsz
aA8i5w03P0U1GM5NTMumVsdBw5w0uSn3Z9fvmxkV9hih2Cshdbc+/tp08YMjKMnXPWtAX7PFma3e
Hz74dWLX7+mpXAk3mzR++c5R5YIqPSa1Wueh1KHCEjC2e5jIAUFbcQJixwzq7FvBig5LfV7AsN+5
aRMN4ELgnIA0VvqXNRYk3ueDe7BNj4ZdR5YusQm8EaWRwYRMyw40g9Jx2xY9XJNsky5YUTspDOre
lHNoHBdxmKJf8s0E1J9sfPGkD4OolcsF3BhwrMZ7ijrDlXpqP8k/EUK2UfsWV8H9qXMZAi5Ituyd
dXJA4RiHXpLH/A4JfsTC6g/Aml0Lokc1KsEYpf+yc+isq12lI8Um26DKzRSp4M+jaIUVs7iAQWtM
MKGxRjObGVnCUZIiYIDV8Tv2sqvivunOzUjKVVIKCyp8LyXZIVRZXHY6kxSS8Kok2Kfpe6ECO+jq
65eIeeNMR+5/86FM22dIQr6jHU/NyIJscXqM3mie0CqWhpmOlGUN/BY4klWFaJ1c69cRIs8/c041
FcPB3qw3El34GppK8bRNqFROLkly6OomJ0gHLyf74abQva/EK1xQMdxBPUuPFaICRqfXuUzmCkhK
jxjaOxkS7FhYyC/n3UseRcKuz37FzgFPZuCKm/6DrKErJ0XGeQje982ugNGtuDWgUyWtpTy+VcMS
2fjXROVjNd7xVh+7gWdpueln2s0hs6wgMR9ub63gL/6h+8LLKODVbJwPmurTmDoeAVkCL/z3erAV
U9RomV4eTLVgRvlAQ1HgvLfgnjyshkqqP7oxToxQ4weYhD6WZ/HF0c3RSKPN6Qk4/ah690hKe1Ji
vTWZ9yG50NDHGn3SZTWFI3M8Os7aZvUiYZ3DZJI39F+Gn55Ugr2JH+tzQ0Ppu1YNRko1NFTe9xa2
3C0dsayxxBTX32lDRdZPYylyvIxTw40YzB1n4RaZY+af6fdHOHsXeY2pCHG/rec/HekM0g16MpMA
SJ0F+91vBo5bTucL2xLhzDUcEvidm4I8D0SsgsutBxdAEI3cRCSpZkO6xeHgaHdHtreCnlhFeZtJ
GWXOkCdhdUmgJF13MWiWmEP7G5/4L6Z65tdHopLI3bfFQeZvn2nCPrMewPe0+MgsgahsuS7Ys6gM
3G3i3KTAeoy6LPtYXEXObdf37xXBi1RwKEdC/25r+HFKi4h5PdkHk1U47Xll90WvxiLHWWIYFH4K
GA204LFZj/CNdw1EWzJ8Tv37yhYbK60u/RFKyv0EMF/O4AwLZYzBa05jI1lVAl04E0zImNzt7SUd
OClK6wuGvIO6YRrcWssLWZCj01iVppyGR5ppc2HJojxG/W44WbNNmVs4NZ2yQl0/MKdVOyf33ii3
oEYGU1Lyh9sbJnk9DYSfOiQtfnzwfublv2Bn5Qu6Bbx2gRUDAaidJBw37Sd5IM4DosgCcMW6wCmG
TYmDaZ39Ebc01l9Q1WwSZDCkf1TJu80rjhdFa+dsNniKfKHn1CPPYggFZJQL89OjfUUWoMEHkI5C
g2Sop5RD2VBfvQoAwJg9YGZxJhOTEWEpFstDrkQwTXpTiYtlWdGiqOWoxRWlZv51kLUD8iBWyPLf
MHRWyRK/HCFlOcuHcpFX5E7WtPCbQIcZbhAU4QQhlLVjbKMPCpuwusGkeWzXpJEye1z8VAF4LNpu
97hepMbGnInyd+KEalc6zujADnmlnl7uHF+1I8vmtroAH/zGVEwmxJxNPHj5cfApQIoOR32vqscn
MGhNVk7I/cOng5RCyEGqHUOlCYZ77An79eq/LKv2tcR8J3Oywk8+mv1zeKV9+QC7XsY3iSpuZ/WA
W3/HZm2d48xAALl3UAzrAgc6tKLG792LjmwuwIGm/2yarplKgISF9FEZHfkHD4aktAhHGy79PvSQ
8C++UWXvBJUuebXuoQbUYpYwwJfKL2vBBZc75RFBIgdH5GoVknstmlVkmNhgqH6CIKmt/hlsLzyA
Xb5OLPN3kHq7/j449IIMW36QWtdqiMTtsK1aTgx0s1Wy3+cfVPmUly0xvw4q6s1XNKuxUPzFAkSq
vLwZD5faDRAo7kUf7tYBxUkiJIV24dKcOBN5HsWodsntki1Fyssfl6UH/udHFcWzukDXPKikK3kz
LRcr/gTLoesFutxv+cnqrEUccpK8XF5xCXmPsWT2skRT2W+QUlXab17y/nc0daNGHYOkiUr6m9mj
HFyKIbrCdSFn8YO++Z9KhsmMmFTDQwS8TKzEPY7X7fLFZJM0FRCcHgrc8Rn5wYndXm/Was75i1SS
85GZw9Dw9C2XgmZpFCXAAFZmayAO5kqFcJs/rFTXYXjvVsK2kgDsBZncYcgGk51QXdbOCpiGS2OQ
D7sW2pQXYV4kN2rjHAyQWTRIGe1UjDkvo66ik58de+H+zhOcztVt0kQLzQWYfka1T10rFadyNl96
tdY8Cznw1wpELqlcieveEAu7Vt1QZD7MovtAAKwljg8SB8dZZ6Rva9aPi3o7NrF5xg0yJx2+jipL
kxShXDsGQcvpY8qfrCxmS/9CAsBOK8S85o08Vdo1l94dIu/q/Q4YfAXXATRQV1OGTngYb2MDR1SA
e4cFyy1LfSM7XxZtKY4RytdPTYj88Sy7Mc4287nScseg66H2nJbGhmcPjCEUK0sGg51X27HWQA4i
h88tkhaecU5dfI+JPt+LseUs0E/VAlo+dGsJCGHrAINhqvbvC4nySpDEFEKI55FEbbNmGgUe0L7B
+29Kn/Qv9ivwU/NvNq7ChihAvuy/YzDaIwJlK7ppDKGFHzpwA3B2z2EeMSoPb8WZQGqYj2Dmx2Y1
koySLVvXkaw6Vlvgia2FH30v7j0aUnai/2485UrF9f3R6XLYeZUWRmzPELnsSxuu+8sylPyVzYLb
q8u5sgvW014LWXJD78s6Kn5OA+W0NGAPRGkCyVyunu2xIw6oHUrxbxFpNe+TCRGWl2YUrUTLLcpU
bw/j0ln5ceiim4ZhNg+skk0+B1EC3xnyRErEsBbWTYeVOXAPDvAw4Bhs7KdIgw5TIs0iSvASSFTy
oXdes/lHHPwlZ9gTsKlnsGwithIkzTSADI0p7mrjigmbc5ksAq9bTqoY7B3nzujpJrKiKxr8Q4a5
itpEVR3ES51/Y1KFq7Afu2O19LsvUS31oXhcs0lpVkkVUpU8RjjaT7nvx67Ksh+Ka+25tc3ly7WW
Sc5qlwXVgEQJek0DV3SAdygADS+J4+Pv4PRy89irXCV0yxogpFTZrLVonvtosJ7caDe2KD0/600L
1U0MTnEoaM1CEAWD/UltntRpiX9pR/uXl7MtoyfYEe0+z6umpWMFVIzkvnbo5R5j6IPWytVyRgUk
2Bono1BcVacA31r9pMv7hHBZETBXmjjgaGe9cGwC+sc28y48hotcgXymxupw9A077EVU6NfXCmbd
KYOIxe5cUClvduJa5Ba0OeSqcGVl4yQ3G83EZRjoBe64YKWfzFonDIAwPDe/wbRgBnwvfgupcbxc
IrrBoFV1QIqITCeJ0bhy/GWsFITz4nkW09U2+9OvSMjidcCBumuELtBLM73Z89bLIJH5SO6dZ2y8
ZgrH8paJm5dTY+/+hLIv2mjnVIQ3qU8BCV87NykYO4OcdKZujoxurAup4EXO3XytXdyM6Z0IFAec
iAj2+PTU6kUbQ1kQFNvVeoxZKQ1GnAoXTD+iLate8p3S+kvxDhC0Hu0h87vvWwNLIx8K+389+hyi
J1uJ9Xyif5Fp4W6vDun6h11q5BjWoI1Hvp721xtEyfNaSJ5tFutBR7bjhJO4mbZmgVdKMC8Qag/W
HMBXrf30DdKNb2/rUV5c7HTyXmAhtqely+TV+F7K8VcWzYLHbU+TKVQ1p5Ou2xsFpM9MF6aj7d9q
7A0Z0NJVJd/kIqkrPkSkHf6F2ZRij/ZIE2j1PDlUfebOF2kDvmH5YG22N2qrbFfbvkL/ZwOEeGtV
NehhrWj4wkeunYsnqzLrhgK4RptLSudKPWPHmxbHJGyXqn7zlwi3nlqbtskehVvHxPeT3zgL9dp0
ewbftkbxcud511qt++qYMWDL9WcGSIJ4E9ukjZF+WxeGDnZzkvYyyp70byXw9MDsc91WpCteHJhZ
60jd2j120wFpCo6H+w8rlhq96vGZhemA0lKVWlPZc5RgTyrO6UAYWVtX2Z8hjK62kodWmYBMeOIM
MzWcXf9AhinV0tggLtOjZNlA/ow5FPqcwnovXRceL8sVkFlfIUq641B1sr6zXP/OHNZSGdfsaWPP
BvwqraDMXXM/O6ndlF9t+0mLjXarQ97SuUyZzz8nWTqYHrkkLzzGB0pGc6246KBAoKEeoRWabT/m
qicqJDZoheT7v6QUA46gilldVRnkMgslVmdBhlQW1woHkyZGgSWC3/4YTV06N1t0E/ve9TxFvaIq
mBM7rLGITjZWImZzG+TaHk5ECzK4QXjm2oZeiKMinPGTsWni8bSooi1OnJBWzLgXOF2PSPikwX7x
/ebpzP/ZDjNXFuQwbH1itZYZ3G8WzU3DJH1TtFf16q9UL5SS+dZhV9E78erXowRlQHQyHgxYwSxD
UEeljJx2TmPDdgGCYmKvAHz3oAewyFJrTXMF4SKj2Qge/a+8uIGjWjXuGW8UFUSHZRDJ7q+v0f+h
ENiJIp5Ini43a3MTe5o+NOTO0EDKyI8/Oq1klDjZwcuathaPv4TnXyf3fysv1FNhXkKP1Wxs1xsv
+cGqiZGisMIgf0IDqWP8N6ELjuEHm6zl4+6YLx8YwtcfHUK8pcg4Y3SlDcFKfeAYBySmkn94YGgC
2y/p1OHyIOuYUudaQ8VmWfbqgVMguxb2+MK2/1ra+X+T1u8Z5ITZ5lpa/6aFpyLjc0Q1XDBQF6e4
7rd9Tmk4yF7SSQfyQKPtVtBJ9pXhRJ3Gmv7dVY5xW/appsauJqdbLs4TtvR9ubFK6vN73At+Q1Gk
9yCoG79QA/XiOVCbsb4b4rJkCAi6xLNnBWZrxWHp4hEM1bBK6HbUP9ho5aac6muHEEP6JflMWgOp
vC3uRfO3hBx7WmJFP+VWm4trL6jMd5wMX5ZJzgA7CBbajaDnaRYZoLeH95vkUOAU2xncLmsmAD/G
UuwAKttCiJ/htpxihWscikNsisU2lB85YJHg3nDrI0ES41gk9YWWdLHh6WO6TXb7QDIyrR0wBuJQ
5iZHYg+jwq59nksyDJ1bwEbGTVBMqRSYiIQClB7EpwWt9GBUOZZD9KXe/rM6qXX0lArpwCzjMJf5
1fppNy6ov8tolNZ7THmD2k1qcvFBgLGzisJZRDj+vP/3JEQ/t0/eb7a5xJmCP2yYyUAhJlRlBW9C
G+clpcz0DWtKkhSz2lD3EBOjp4W2V/i6TWmCQtSMMWDu5q0FgIe4IxbOWd5/+ZJFYzfo029hsQAX
hvwg7pLc4+Rcw3ox/fYCzFAA0ZyrmtcEPGi5MGjc8zG9txnoJuqDpe+K9mZsVQlZCSqIgbAFNZii
zbe8qBpl9pTqdimvo3TYneDwk3ZP3+LfVRINOYCZXlAx/irIpo95oUd15KroEPeDrzKKmJ+hsE1I
cWOkPQCmr/k7jDiWcbDjLzP2BM7VpsbOQUFO/s0UTllX/T2N8/D7Z0Jp460xNGQrZAD483zeDwyO
dwzg1Q9Y6Q5jo4gZFGHk7lyIG5iaRujblS1rG5U3v2zSz/u1cjSswrfLGwFpUSRyO31qnTRSG071
86sWYcFTOv0R9sOTXEszzaLJDL5tfn1qdRXGsrzFOardKOJAMryp3GFoB56l5HTls8jhZBaLgrA8
4yLAJWFt9UAJnyC30WghmQOi2z9K8CVe8k5gx6PJ9zt9NztgoUKfgGog2tRy8+IKREu3lzxSSZpF
QXaKvKwT184SO85Vjf5JqIvy3w2qhPUabqWLvauJPy5JHRFXWLLJo7fJ50xHmEj+2ZsjABpV2BjG
W6yyrrLFufF0gKh4N8j24RysOOvvHe1GJcqFM9vYf2llYGbto3RoJbzKvR9obtIsw6JzHY410TFN
yo1Q03SdUDWV+00S+1s7xWf8xJ8Nl3X5LwNPaE8VXXsTytPt4ur/iCjs3xxPaf72iChr8OWpYuCJ
iWZBAxiX1mIp+yVvX2ftpuzHKMyY2Otj2vfok9+0S0VWSBVq1Zqxz2QFODB56ahlv3KeiwKHOA3C
IklOhlmtZPxQIA1jlUvT4beHobi7Z5xMMUh+BuyeCFr9N6X9RGEE/deJ9ZVZah2hOu8gd4WKyFiR
UFbN0O3I+Vt0CjcirfYNzu9Pw0RhOMRKgyiO19OQk7YJ8kOUzayRsy3ZwZ2Yi8W1P+s1TdTrTEBh
UNh/UHZr6nVf8ViMt+S+jwsyQPBV0+YTSVivWiy3H9c0zaNyRt8p4yls0yMKkbH4iHJClvlYMHSn
7WAvzfnmuPv93+vOSAga5aVwULGrfxLiNk9wRQZbBjLjhqD9R76KhmFuhm/iYgQ0WXaeEX0YRU6N
Jla42BbNNbaIVSWZNOiED4TzN1s5i4JeVFHVWcEtBFKZLXv3JSztt0eRKh28S8SH5tS1mXT/bWCP
/7InHgMEccA2PM6QIZ+LOrsmgh5AnUvkK9FuvgMxrxLmfp2Euarkis39QJsQpLGV3X6k3fMsBJl0
wg8AYt0/MTA3DJw6v4COeDUYFfW2xoQ0ISeeJrzYFVHc/YKhQcziR15XAg8BhELRF0JzXyWZXMsA
QJTOquvWVe1Jz2qWMw9HqbJSNehzBhKEdzw7gPCsaxfHKoOF/1u8qFqyyki/1KGD6fJ1iUY6gWcV
1qz/E62tnUgbuyy201npO3Cee/ka2bOUvvr5IHN86cBkN4hcG6AemPKRBIGN868SvrrgO0BZobCQ
9IXwgi/Vd8j58ji2ejZTl+pDak1GhVS1PC50JosddyG19gqPS4wVds5ETdRugIYHrQFGjgBO963g
Ls/wZSjD1v0vM0k8PJ26bm7A8C3VcmG6mn2+GiYF5e2K4GFsbt3wd6OT68POAMwEd8UkeaJRjSnL
9YXEC2xSm/MUXPPXcl5TGSM5G/8hFprra37X9tzmmpilHfvoehN77xk68EzlFNF6+dNv4G+Wno+5
YoC1rmOxauvAwRL9znfqnt1j6N4rGXni+LhCepnZVTAtb/K3FAv5bui6FCe97Ku8cB3yAS6RWais
WNp8clR2/G2e9xqDCr+DD6HGbQ+XX6Tk+eM6CA09zTOZJNigMBytPzs8VjsDjWfEw6H2XagB+jl8
UwBAC5Z9+/giVWRLhkC982kqEibLv2KfaAgKu1hilnAxlt2mVdGt6gAPFYfD++zI8mnMApXVrsHq
4v2C/rbQjiNYjFMC6c/DwTFtcuN6PGpQpXxM1vUultok8WXYnGQiRANWGrY+SX8M+Uv4OrARDlE9
mc/rfW+5yX5plk313qbyTbLEeNgQaXWcVn3U5eZDp0RwPd0zgpB+xmGeDSTYOad3AgaGPjBg9Hrs
kvP8FTZ1reoy6DRfKycZJiHOdwTUoP/JAZMNAM/HWe6yfS0TmMj6Xx4mUIjVhfcVsyWi8FkCWqQr
+wiGNrtVJgw6fzB8dWCI+ZP6lH26/U50Sr7IevXrYs37g7FT4mWiu14pfaBXkNtgNVwe6+37aAyk
ADhcW/3ycVUEKqa5Hx4KZul14uQCZKKwT0Fj5HoXp8qbMW8vOmrZszHjYZ/k8mLCP6/jDZcbRsn8
gWGrfFzemdE+rzmkbEIzpofNYYXOtbiDyx+oqJ50Yy7k9gnsgc6eaBzPdb+Y14Nnznw30m/YSuRA
AMZgr3HCCCBj9LK1NhZtbvhxZQm2Hc8cPEH/8coBr226RQFSkZJqdRp+AY7C/Xi8hutVOxquqACt
Dg3J2n9dkog5ecuYNDn61psex6xrJdf/DI0EE+CYxKMjc/xw9Vk2wFq1mROnOHlh3n+z4A6+cmEp
92314nERy85QeCcdV9KiqN80LRk7IbdANV0ATNl81gxg61dNyIj9iArsnKBFvA7PFihj96sKoI20
pQj5dn12JtsfXEBzL+7SpcEdffM954Ao0YLDDUieUQo1173Vt/7l+6EGMfWyIlcNymH+ZqUMThb0
E1fRCWxCWyB0sMrJkVCXEAZ283t5e0KFaZReILX8Nl1eeWsEefTvGHfkV9FaxCm+MGOhXifznCws
/9WOurJRXpp1LWS6ajVoTSCBBmzcKCIqJmBEGuL99+rSaxezWhMYIY5c88JNjnhtI61kRDckEk4R
jRfML0qUDWSGQJaN+QbuupOxRSmSV1pyZs+xcThbzcwHsJ/4Tnm0+4T4c2S22NQTo8tqwCAjMjZb
NsHZn1R1i1/WGxWhwCo3goRB7EowuJ0aQZoT1mjk76woG3GiuAZUbAvdh4gnUtnpvXLToy3coCKk
HmysU/ouoBtQqkL7ykrQ9LqkC3hWV3EjyThRH625EfKm6XoRM0H/O+e2AT7+QmiONnvOwOSspK23
fgRV72AAZIqD2bXcyePZKnpyrtWwAr9CzO3jmJUJL0gEtimULW9sFxurIdzeQuPKEFARXX7G+s+d
NRGDJTFcR3v6tWpYdT2GTnm59tBZ7u9KwUuD+LSKPrNbuS0Ftyos/fuQAPBvE7aNOTbU9DnTo2/I
4X6zwomhC2+16rVeP+pb9LgDgYHzdixAsiJf7BBkHmlyG1elJiFhixCekY618mE4uyYlKfGl/OD3
dbWLqA0ikj2gIcoa9vE9yc8HJX9/He6Q3OFzY6ATYTFNkxS2TLl7ani978C9MjInzkTWdWcLKUzp
UugRBbZOkdnz/EEJUnf/sjpXYL1K4tJhpS26zqnUjZEP7JoQYL9nF1JdDFthGdkfCMywunNUYR2I
rCSa6qfxpRO5pKVjnAxuT5+FVSvxuKxBHyWJO16HTt+vg3trD3Al1OlzyLO0s5I6x6xOzSwc8wp9
JwfZFz2vmw5cPNsZDVrLCeiBer1TpcRFUh9MWrWa840poKszKkAfdapcuW8ZCl8AiYbYgIL+gAmS
Fsr+Yh7bq54OnmrgBfQr6Hk7C1Cn32IzjzuqR8CoT9qi9Gh/69Zk18oVLHtGg8iWVaUbXyGaea5+
OIbjBDmlVB+BWWQKASZcM5SCWRKdi1CIcpyO6V/PrWS5Z74mC+w3zz+0+mEqCh6R8K0ZVLmVoQxh
agIwFV1xW0wUT+1gU2jcnCHBzsY7vyA0cXBVdm6Wfv08vmgkcWh0qoEvgc6qHtBG5Eg+f/bDl9Mj
+I7yAkXB2I4lj7ytTyfgWtSj2kPkGpIMJi0Dl3nrs1FajF2ZOfpD1PpYQCCRYNEDJmwOOaHUv2UO
13UV9fy7mf/dAv0CUefCn7JP8I0n6Xb4gu4CdFtsq4Nkpw7jcq2qBkk/j40qEgZid6u6BTd37RdU
rDRD2roLRgsZpHxhXyXGGjo7OEBRgLkEjCjq8tWZ5iB9hLE4ickLIYG1769CDN7n73Saw9lKmOIf
v9Paqaf0cwQTzXDjxROoJL5xXyzLCaeuisu0d08EUQnNrGU/tIIUngenG5lpGPUxhuQ5L2nXWMqB
jWDdy47BqC/JDKvStzwY3DXZclfPP5pWhO3zrc0J6Ort3rEBUaqQ0frLkIebYcaWO8PAGxYJ9Dph
x/8pBDMyOiFlHNJTVeef5MhZIHukFOEt8gm/aykqajaafT+hXoiILi8vu/kNn7zDj40YPIgb36i4
RUJsWb6yBkD04jAF9QSL2Gn7qVcN+mpgt0dZ4IQXP3ctyaeMyv+hbZc6haxZLvinKQncb0ANRqRl
K4kNDVsgHmV3HMIlJTLOxyO2ZytDwk/QCS/JjQFNjf3tP/Q8jiGotK7LY7usW7aYaDxXi9sb1SAZ
YN4MyFz+yMws1CxF0dRc25cAHZ8RHP5uydhMzYRNNwT/0cIFvHU129IUo5Q15/A3IAZes50P/PFB
srATPatm+W/Mx+APdZlWtoR1hNCU481XjfJ34M0wE4IyCfNel4wnBVifyyEOpT8Qq1RU6n7Z3VBD
lCUWSWK4Vha6xas7nvYkGtmELxJ1lkk5g0VrvopVjK64l/ao8BVr8uI9osD2Ba0TUKRI6bUAc31o
Fo5SjBzWU+iIFBQp8FoJEWoa+ZUQZlhDQrVBluc0dNTyXtEOH8mrtF/Ffd5HNigBhIH4mMC94EDl
e1EkvpGTEgXQKoVlzLS2m0yWlQ8OW2ZJE9g/OnhPON84BL5Mt1EFWzh4pf8wx0bYP2UYjC0Ou3RG
Ax5H9atBVGbyyeQB21hnHiog/29ZZb633YKq/NquiQbHFcivBszHppA2p32RgLp9WwA/02rSQ3yi
Cck81GK5DhCityiC4J8EtkOjNE1pBA7X1X1oMc/MmXqjlFwsxphnn9mvmL4ljLOePKlI8yD8g66l
rlzmfEjnBLvS1gEeL0uxmPa+Wi0Kjc8IMnpaTtfqceOJz/5+tzgdypYCnb1Jc8xHRWaJzH3RQ5SL
Zp7oZ+PmIiI2SSOnOluHnNjpjWb65A6pVMRvRsLDo3chY6uSfZj79YeZDyBhfwDkGQh9Hup53+yP
a1ulMgSeaaK+D5rD4wMK7tqxV3wEPOd3m87uzz6tHX3Yx4I4GB3Twurs/mcYsuXoSN9dh2iW8iD8
UTZXUt+nrDPGubRaamClqihFku3DA2MtEhtmyuzK1tEEa0x4S8A1Gf/HuiUlXGPBy88YefRYGd3/
0PwYq+5uBjTlYl8AIrourB22K3kekXZT8WTzsdCzevhTyiBps9QRbCh5wwb/fg8/O0fJaz3iLYpo
Z+7Qk7JBpwj6yvfF3YmZLnno3h8QK9Lx4D9b8VQ/g8PiZKEMDC9/h+tBSV4RGNYAqOwowBOigNA5
FMiF2NINntcJ1ET+YvJMz6obvr1mvBsmJ1AXFLZ18wfJVtjLHGh5Hy9CrlfDKxvpE0l7X5z1kvNN
Wzb+6F/CpKkTtAxHMd9jjbr+PArodAvcADDvbWPIO2BUcIEAgfleb/GMp/uZEZIH3oRVvs8mvjyx
IKEHBFw5iWQy2ni4JDgnWxLqc4FyQP3MekCU/R7u46/IQPxE6T+BV2x5coEj/Uf+AWSGJL9agEjm
NJLObh4NE0e8eS1F826E+zJD1vhtkdjCboSI8W7RwfLhHrZYTmF9bILPGyt0Q/JYHzYteuE1VjO8
P9njOIsVNErXx7zy14nIhVgMqxgvpnRo1MLC3eODMkHqMSBOtC5fi+vyFLdXjFHJmYVLYHFN/RAu
677+b4/hDnUUIgYnlTCzxsy3cot37ye9z3WD7EL4nb1qVZsOz/Q7sEQIzROUc45f5E80VJfJpUSo
5pm+pHS2x8BIuuqo1dDIXjHNHOLsaKpzLOU3jv8thFAkCe02aSDxX8Ok6EyQ8bT1gJPY0cOtshet
pCKDrNBzEm6iv1m4XOcVFMRcgM71GTS/+w+yVRRsBcIxgXPJeFFkFisItUvSDpbtcswedJ2kvndo
9yP4AjMauawefxo5nXnv8DUJ8hq3GoTp/ZnpwUyahohTU6tXl9WQ+CXagTyqMUGcI2Qush23TLfk
OE7uYuaaGXlEYCRS17YXrDksMWplsXti7SAGmdrdqne5C9OyayWozsac5OduMVy7Zj/ovT5kymzQ
c9octt6ix/9k3qHgCMmcxRgulmOnS/ORqC68PhLlEmt0/unt8UfywtVPBaKJUDGj3i1ghWxI6yOs
kZtNQ2UJF2cDNHM6GtUNEGmr+0eX4YuuldwuBiQX29v1swDkav2oP7NWCZZklv9zIGYp49GGP3LP
RdHk8tKoaCK8JCxYhPRUkzrOK8uAghpsPKhNxBNwYIWSaZDvDK6jiMFp+qbtTtiVaoQI3YZjaToB
PViaOjq8vk41S9qtGntoA/3Dn5qJxw+4u7zFBq6r9jfncMFNEBtYiOjqlYL10PRjnUZ3rjXamWGX
7ewsGmTrsVBOlvZaHNzO5Swop0VaRO8ayfqTgbT1MNOJ4WqfWz6bYs5NqKfkDQBAQiB2RlRxDTFA
qJFNJNQOIfNfyso9DwtcZ6Gbt/iGTAKkRYWdWEZyfpObQorPmRwvfJRa9J4RhAZbxTO5/MXtDv1k
G3F+30OFPu8QTJzXi+e3dab4DDgr+PVcuG4wPv8d3bk/Yw5x++K3yThhfng/xALYc01xU3hvXq7q
qAMtVyMl9wJWfCbyZnCVgFL76YLkXYkjglo0nZo/ML4QzUWQEml2iXEdDbQQcs8FZkfMD8bVWcPL
pMdb+qbB5/fMiKpYVT+PFQ+MaqtgW6Zq5gwLkrt7irIQqeEQDmmd8/SBC3impZvEOvUWJ8YPQaP2
Yp779mOEdny6Cbcw0xWBK65BJWr76nqVMods6/4CQO+/iwSNUSCEgoJpp9ra7RPw0bwdoY8neODY
totIwRPBequau2n4/rnKJMXo5nOFnX6iA6qLtdxpH2OAggvuUqMDWZO6RP8MSbRqXhDDC1pDy2jT
KpvSqJv6wrUEXzZIe9Bu76j4AQBlsvepiRyxY7pmkFAOc7YEbkJ9ZR6dt+9YQupuOp6UrSV4Dbbh
bWyXDGSwuDSlYWZTa8iLWvBGgu83yGdbGUYGXRskxR6bvtYzo+PDaHReWw1AizlqwRADtBhAReod
p+9Ii1hC10gxZMoWbXD46ZykbysSAQRziKuhkgYpkTyIHDfT6sNwVfyEvCKDcZFaA8g3VKL6469y
BxevQkmUk+SFA8jT+kvSVzZCkDzIih3kLgMJ14unzHmhIOOjUOxNXqsKX52vPEd2oKd79h/sMYpc
8E1F/y4CFu+4v7DJ8HR2ZBA5/lj395yOXE1KzQoiJaBX+bPU5qMIwy8V7yuxuRw6SMNgQPQ8UD0J
M7xK7drgvoP0MtqFrVc05LCo8LMsK2oHNX/203pIpcLvxYMVc3GgWlA/F7SHXPwIH8Xt7NOWZKTZ
0jQSSdMzSadwdCe5lZgKAEHb/IEMU6w0tuhgkUSM+sWP3bzM98M2inqA845ZsjWsD6q8g3ckDBv1
n6oGYdYrLtyvNGZ1tczWVyrPZYvEciop3EUuiuSe1no1kTsm7b13w5l0x4bxiOqrNxoE8ftVhC06
GKWRufUC7Jflbyuye03GteLn9gms23VxpC4dSwF8ZPxVHgtcHVTndD3l7wcn/oW9S5iItCbmhc+I
BbaLM5JWiDQwK4UUBG9rwZWEP80Oeay8d0XpN/4Q/MBvSNRV5le++32IVo9Wdh4h4GymcmC3yEKH
gDfCbo1kIfk+u45Zq5Q1dtDLJeHJajcTHPpVOygySyVpgT9MbrTEVsmQfcbm615xSCsVglDOtjAp
UJ1Vs51BhN9cjtZJiQ3hQV1EYjPy9u+SSqQpoM7H0RwLFJpvaMqNVliARG9g2KqJsZBkXZ2i6hPa
xtOtHN4yIvs8dE7bwNUQHG3RPkvFL1yskvtFkqzXAA2snYKZvIrh40CfVF4mcflwl5I2i+22bcco
RVlyaYHmQtEO5Odb5smDivqxBwwPXSFklrt6dfAbZNdXTn98O0pCYL/XME5/+CItmdoWyQF2JgkY
h6AdY0VfTs7q5In5ujoGAVIYOOnjcyFBJsqFnGoNpHSysuBKQ/wHRY2Vf8UxsmRIpDJmJP4iI0vb
fbe8mqLf6RPmhzcj01ZIxlKYv3M+E0IS7HELTn8uQC9y43z2wr7Fsu6xc0ZOioS7sgmzublx6Jxh
hyaomXjlIe6WHPzHTa79ba88xJHkJeu1sVuRjGZ9xfFe7pk2JUBeOuRfNYmCoLstXqG8I/q0S44c
/FIMRsDcyEc07WrU4TeQGhQLIpkuPKUUb67XO6OsNVoNTBOkBaTxbWn6JDjnJXglThw6IZPAb2ju
KQv8ZPg8RfPPoUEPR//tVoSvht4+9s6oQtXUi5YQ+TmEsjFENWvM9hDavVJxU7lMm7ZhwMAtxSfB
OQX/PW5KAPkn5Eht4y1HsF3Wkcwdmdy/usfUpRQbIClz77MamblvhV6VhUQvVhlTrUrfizXJuPtU
YSzEFG8PgEMU0azjJiDGZTsMlCCFXivwIQmm/pIThStE4pV3XWGf3VRfjbubJru6TzEk2el/ZMbk
pqaUD4FoqxgZnyS0WbncLtkmXEUQLJphKqF/cuKh1ST3IVdsNpS6TZW4QHxzwrHteSmWVZWriGyW
K3LDSj1h/qNl4xKRXnZBJhV1dDHdeJHPilhpSesP2SC4HTCJe3ixVYuNoNco2V0UAGrAOqMaQaRQ
tTMIP5h5dqVEHmsuvMcrOCaMpHwh/7VEyv4EsCJKKRe5np17ISJ/LbDgsYXrmfWXu1zwNIfsDSBJ
ZOjdNPsuMyGklATXkZonBF5HVHcMPVvhkg5a3EPJkTXAsDPjeESmedaKwRKRBCogLAoBC+XsNFBu
xq8r1p/zV3+r/BRLL+D8hPbBJsN9XbmTpBQQd6Xo4h7QmfSiBqHglEzLkMVt524UlCJV4EB/XjAV
/KW9A62DBDJ1TYNY5wQvpft/YZt+a21F/AE7WXucnEESZqmFbZclXapwQKASUP/OHGIOmN9hhEvA
iVCrFX5xCKCJRFCLQCPGnAP6DlBOuzMqZ7/Xs+SWsNEhndZ65NTw1kdcyodZYwazqvSrQt0bsbzC
OlTHHuDdY89nTRsLEk0IVU14kEAKmEfijGmPcMCtAgtll68ViBaW/YyV7fJGNo0I8DVnD7ToOlE+
2Cmitnd0tR4AAP1moEoSezjiJHH0z2XLcBmB1EDUpNhlVCd1jYsQ8wbtiMo0me+m0Od6vk9cYOxn
u05OQWMjKnSyTXwQsC/CEtgJl6lbr++bMs9U9ScIGHRBv9v/9xStno34ErSk23ZSHTQsw94Fdm2e
EoXKRBMrNXs/56+IIYYrOYDOVOtKerAYzymmsQO+53ltVJd61AbsLhfqdhGQYOJNpB7jTGH9F3Cc
TettAllYiAG6bkdVOP+jbAv+M+1/KAvPYdpBinyrGgxB7iWd6qll/V4aasts7FWgU63bWAdVz1vU
PvtMDMyD6jG+clQVQveAyKPNxtrXlRMwsHSJgU6xsGtEp2gZmyvN6n+lQFLBsKCLCbksV7k1265m
gsAqDSzs2+SzmFV9jUeiUmU2rf9oZYoxBaBpiTrtg9nfThmE64vt/4lL0VAwNTNW6vCLzLKhHNBE
9G2zODukQAhhWWqtLTpx/d3RuqBGrFRxX/AN88/7VUbNmkqHMfObq5wcXee5bW9lPPWttHCrTAxh
9VlU9OXDwg+BiTSTeUVpKDSwPbBxFT5VOc39dszmnwBUbTCXZalmbgFWcGcdzLL51fgnrmrhQ8Bt
S9n6Qp+Rg1vk0x4Z6g6DL4HXiQXmdXJbZ5JsovoafkONFK9bVKc+80hPxKhOVoFxp1e1/158HJsu
8mYO8bMwrLnBc4k0Aadt94GZWICv8b7g6s3+LMt+WkfV4H+0rznIIw6h8y1G93SS6FLdwaAfnDrr
uhue7krkZjU9fAL0yd4Y82A2bVBtoyK1M5jAbxpzPErffX9y8lKTyZjNV8UXpiVaEzdUAhLeO65n
9PHewxPitL6Zz4dhVGgl1QYXGL8Y6xkdM7PFlJWhbKFMhNVdYzHV15jcQLRcPZyrCAwJSsd14NUm
5x/eRQzEWRDga+jM9x+5ShvMURs+jASntQxc4HqZwxSnGIz76l1NJNJMhQcUokPWn9LigvQx+Itp
rvv8LGeHTkEzlmRYAXSREKve4FBpiaF7TPUTJet/Jl03YAsutmJhQaQJms1+gHSyBuk3Bbtp4PyC
kAiU0ktYhvoDL83kU2yjC+h98ZIBqYn/pqBRcQ/ce1S1MX5JyokXT2k0zxF6OR8iIYyXGQ1ai/Dk
FEdjg9w276a2BXPU0dNTo45OuCThZSqktiw/QuIMIs/whzHDXPtRxMTkeed9R+iN2yqW8Y0mDcZL
n5paYALcjoFLaKTqqdC1SkPLlRa8+kKPX9yl+XTiHKQrFSNb8ydXGxt9ZNMM4bssYl/kklsh597y
yDbBCMZFJgXyiKPcS3AWoygemEhmkObWbwHQ5B9N2nCvY5L9To/ILGU+MfwhgEVdsFqLy7r3TxpU
MFRJ+A8bgcWaMJyc6WUnDlLJdENA9W/pSI/2x3yM6WMmDVmy3NUwnxY6IxHD2P5tk9T7Kp2R3xTT
KYhSN7IPcJwruXbhzBPCfqufBDDWO3ZDHnx6oa8jml9zgiFXV+/YjviBMzslxNv3ARNKvVYgcz8r
yTKzjhlQRz9c6FfA/vZTyejwZ8Qh5LCUQc1VEGGp2hFdxF288O7KLfXx5x0XJM+gdEQswiBto5xu
BNR+iC25HSZIZ6lpyTanyH/spGlcLBDH5fiAc4KRYvRdj3gPfR7fj+pQQOWviiauEccwM0nKlGCL
T1VlCB46S1Em86znhfnZnAKVg3N2DNfvDubP390+s3dqxdjn3OnExlHW35CmTrf909T0QVmQOJ8h
mjYB77xIpx3lZsaXNS28J8WPF10fshjCmNbueVIh5s6e6oN28LoucTP/FIH/op+a4CxTPROe10dB
G/HE11AlZVjX9DCwUucv8T33E20M3kdpO970U1C7XZtP/doU76evdFATJBMFtuebWlhi1syV2+Z/
8J3s35VMDEklzdG2bGacnkcic17kR7VHNDq/YQ4iQMK1op37PBkqKBxXQAbVGllg99H7IkSuiLL/
gaRGnsBSFbO/cACNNSornXfooXHcmrh4tCJ6xEPyGviIF99E6hmiENxbY1fs+Nq9+oW0o+R3P0tk
ePsLyHNp5aJT4oXdIimttpU/688UsJyUra2VqwSMcTFK80bBpRPZNI63dP3KkcdZmySIWx4tPktE
kHCRDNdB7AeGB37396a/8oPGSjg9Ooq6JwMx+ZelRH7vlauaMs4L4BssEUthSlHrVw09wkm6wXbA
hyql0Mrb2pkmh0Bp5oJopBV93YbdhaF4AInuvW5u/2TPFJTZ1g5nEwaSmJUhkumoyYPa7SGSI1NR
nJD7/nd6n2pkgHfVwXcgSK+bwFRn+yIZqR5ZlAEHQLOsNfiLSn0iyMIDxpe5dmVrUq/MG+VCzTFi
36DdLHZ38KppfAdK0+kPNjSRGnDGVHJ4tULeFPstPjO22PueQDwe5hr8wh9eXFsnmRZRKUFKCe7V
p71n8zssYd8CglPYZgeK9lUR9wCPXGrs6tPWwS895elJkS61RAD3xJKrf6L59jt6ebLroiCYCgPs
JlJz0kEF0M+XCaXitG8QMw5IJ7aqjuVmjOEt/E7I+vmcbiVN2t3Yb+VzHJysrCoHfX1Rx7funkCO
kx3NeRpl/O4qBl2JrreEZi3cFvMrxp9nCzDa0S1+f7Zcdiu5sGivecGNufh4Q0q1BXYdBkeEJOlx
IZD/hnFepQE+lcrz0g++5/5q7YB5NCIgVxlh0l/yRyIVA0PgFg6zTsQroGBs/04B9d3BKDTI52Oq
hYWUyAO3p/GlIwIX/7hSuN4I1nQ3ZPjaaW/1ZXiVIe7FCFhfY2TSLYmW0ju+2c4AEIw8f9HSwqPo
e7OuvtCA9I1s9V98crf6trRTQWcLztzVK8YR2hui6LdDU0r88KgAZjaa6zosCX1mdWM+HhVk56y/
KmZktynTo7fc83m1XK4VOsRhKsjYNnJ3yQEXBrHzoCxp8vJaJwcwbFdm93w3next57vLqysX5YxZ
dtnREBSxrKa6YGZK6wWImWPi4pk7XMeGl5FxPLqcI6evOHa2HEibNPrN4zkOsYBq+BLO9iaYKU1r
3xx8F13YzE11bJzTq/DgTsd7rMd0YRb3wDoTkXcQcB+t1IiVW3ybhXCfAcRfOxTziRLY1CNtoh1a
A7LWBL/OEG3AV6F1tg+NOaf79WtzvMR4AwJLcW46ZaoWwjgVOEtWzqs5yx8DHdPKoQZ4VlPLqplp
qSuNHDygSD/BQmmH0UQU75Hi6fEwMSYOcr31CEdkYK1K38MuyWNMvJQfpJe00MpN1Iyrs3wm6WHm
VeBAhZpWbiS8uUTQBCEMu7izkXr1GNnWv3EdqkAq5w7KCtSauvSt5A1PmoloZrRFI2CjVJV9i2fy
MXkERhWM8ap/Sx6ERQXHsVM9ylBTpd2wl+AdrxEIspTgT1HncH7W7++ML9FPsdbL8x2KnrgiAEe7
QI8+Ox98db0UAncRI6BtVRLTnwe9Ouv5vgmbOcGp30xf8bVVDxzk9ZiOkHc0GnfKqk7LS4uIo7/r
2UpZz4lZp7G9rhuPXoSAHd5msvPJ+n4Qd43I+2ka103RgEpwsMrbuzdGeGWJNg2lIZME03Q8BOx5
U0LF5m0ROU7JuPO2Z/nUfvMGFYIbPmkGAZy2HqZ5yf1cXpCN71konuPTakXKtQEDOim4YLMm3Zhh
/2YvNigvNWkdXS1Pyx56DJ+K+B2Rsd/iHrikt26iuZhGWTsggRREXjen/5qbpEj1UqDu4B5R9TV1
QpEjIZNbklxyts5yj8OqYEeQV+ojI8JnTk9RbFEcKHF0tXEd8KenWM7TyEJinfEzbg0PF+iX6RTg
+V938f1B85DJ069yVs3lxOdTKxrXHtdKkPZnTlC7eAByPC1zZN2E2lUkprQBlcyTt2f7rmpY8jHw
ppY5iUnofjGVsJ/s/i/IkOckP3qr8nGwY7nLLTl4y5bYC3mVGtl22Dl/g23f2kTUfIzhoUDA93Qw
zYmTwcMoMVghtbuzU9pMb/2euYpcwcPXo9mzcKfpxB/4CLuXnW5Rwmy1Fb0t+JwmxFZGC4Iz2p/A
y8MSqN3E2cvcTsNIbLkY8cxHYF8WNDHIDC2e4620a0dU33S4Vk+REGrRNnX/ZxJpBCscn2yMcl0V
eI3No33leijTPL3V1s/qV/asfr2RueBm692mV+/uMYwVvxTbEIPUB3JIUcdpO8fkm1Aa++Xbr9FE
HWvoG95GSydZ3VeX7+BMFJljs+AHV+jS+YZU8atCntRsY+pIHRmh27gGMZIAnY8/0Uda1FljqsLS
EksNrgvsz2GEuCKVOOntfr4+Hm9NmcZVWJu9uO/oKxh+T5oiE7v3wbqrpeFWh7lQ8gthWFHmCQTk
TPgqOzTBkoT+N+KECAE3ec8AkttlIaG/GddLTDL1+ZmhZOPwN0nJl+yelcZHSwnYTmv9f5+4g0+f
5qgcrC5GQpatStcacdwRLdeVDsmlk8dAurlD+0XpGNvm7by4qx5Sdk4JzEdEeGAfJwtArHl4fP+z
kOBYpMXNO2QgT8MEgRhvtDk00g2G6agV6ZkJTuL1pa8kaY+4bppU6BgRucVp/lVluo88sM7VSpKH
F9cBW/AAXaYoykzkU9ItczIOVEAEF+Mj1j5Llo3lS3WWT3BtIelxga4EkJTUX4LI2JMv6UGXR8DX
qVgYcfSkOJxvbx4vuRWihHxA0aoHCzvi2qufSV09MFEn3T/J1L7oC4cHtOwIU0z67pEZ+uB232nJ
eNbnQ/8rzWiREuGP+RiAPs+rHNIIo6uF5s7tXbDNIijcpxh71ztf762xg9tUrVqm7ISIf4x+nqtq
B5S+XKBKn1a6du5eKPSSekf6FizKXVj0LvCSZdp4274c9LohM/UTvwOzgQNF3Its0V+qjfzI+M5h
BKJZb59WF0PE6DB2FRalX9Fs2X25tnsL65Jk5E/pVtj3V9NEw00UpZpLrufzgZltIUz1BiHEA8kn
oRlVJ+nbXQRsXqwbWIRJz+HF+EpCHx16PSHGeTYYaVsMzmFtSe/LDnUf+gxQt66caum71inMrn0Y
Hb5NWm//1cWZQDtNuL+ejIP9vNcJs5pHb2ruEdyQJrZ9Zq4dndWbxyRL7125ohNXO8kiTIxhWsDS
FeqvCG0xqaXgCcjkLFp4vh8D7gtNarOvgBmMPIDeE3Scii4nYxNt+ivIzqEXfE36xpmA2JcGb5k/
VwRQgmshzHQUVA2CqZ+ET3zMMq8cm8dDUTSGmlMhActcsr+cM45ymzy/9I1amf4NHhgXPktrGy09
RtdpePATVQvuMeHAJ6EgtQfhguZ2sFA0ZaCx1FUFSXo6jaPqm6/hjtx+FZhM75+sUQFDlxfSqRXD
QFuU+k4uQsaiwrASIMmuBGzogWOirUmgqH3Ctpc7MT16jJhqpQeEmtGAVfv+0kP06O/lhaZ/gmQ/
Ib5n5OS9Yjhyq8zEE5Ke/5z5Y3qJtVWmPdmrsIBV7vj3N8+IFBqjX4LeHe6lckMGVW2ta2qH5Qhz
xwKCsGl5XjTPZu7vggwgxTxc8uqoiGYJaShCPGWrYtYlzl6BvsNaiNyKLidw/BnfosbOPPw5uFQu
S5rkPSgS9S1p+tTEKe4gePBDwLPX60ah3BMkRNM0CXCJQX/vUXGWOdIl9a3U+R17Fh/O8vhv0d0w
WdJou6lDqIc4kQ4RFS2Enq6SAzlWlJ05tOEHGYZn4m2boGqhD/lo7TcHp/KXLIrhlzU+2MiIRv/8
OhbF0uF/So3U0mFYdCsfwMfb4SGQASevKDTQH2HoEyWxOX0x3CTyeMnlNNW6UxfUqPmWX8BxzOt2
dNyVFSkISjppDYokSH6y6SGIbjOHnzBfqKcsMYjAVtqB6pRikUfBTHOCSJSohsXpXONaB56llXUd
RnI7npOL2mmDiZy+nOUNa7Sr7O4pr3OpHBzjxeFfAB79KyrXec7bqzSElvqWjOsd6AW7n6HJjHjJ
vdySYJ7X1H3F6Vhk/xSn0bkadii8rMO8yuq2g3MlYU2ftyCLtQCysS+4IQIno2H4RozBB5VbLr/5
EV6UCJfAskFvhozbnF8qiAV5sPK1mkW5iHmRqXAdiy7ri1/smKbxwu+0Od3xhbytgE0N/qhH4R5A
jg4kjBrnLJGiGkqy008toSIRrv3O/oKP96aktxA5w+lY6Ing2ZBxVusn7ebiJSLheHhAWVDqqBDB
ntOI0cvi9uHkIn6zPhg9rhsqwVfNge0rp6cxed5TJd//jtERfHoJ/mteRYB4bMCY7EeamOK9vXRl
oKXMxnYqNV5H1VV10GRAIic3SQawezV9BGQJjAyoYiXloEg2NhLqoJS3cyv/ivnwMmM3RqugbJPr
ES1jbFQqquUiaeqEe7uvCOgHExG57smfVkH1LQULg9692F0J0vhtwX6RAFPZwPBnLmKVoysuCsKJ
G6i/VuAmf13Z11M4kHfN4kyAP8OmuK6cuYItyBpS8s0Q2dlPYSXWi+/dEz5HwZ+dT8NSjUnUHyNI
q5m30mzCYP4nrskRbd1Zc39I5cauGYDz/wCYewcQXEsO8BYyIT+ik3z3oYahsf5ljkKd1sdMsVvQ
x1SlqGAg6P4bfurFc3vrlcTUiQAzRQKWsHdKMcr0UCCsmn9F5X7Hi21Tojm0XIcZ391YRAo4iYnF
f1/e3pIVmENuf4PCx7Pgm6/gzhYQhes4a1VzEu2kqiVVrBVxzfkH4lsN/X9gBtn7L9tXWcuQ6ZOn
qj+1HbVieJ6biEN1HK7QnMhCMZe/+HkheR7wBQ9LcF/Mz23ayzy5Ql7PKuccVFcE5xS+57zwFl47
Ku0+4MKhdWmT7GTZaqaV8Jh1mZzG5bF30kLk4uNQl+WUB+8n/4Yh5rAO0saPvHRfXZiMFfIsPQ7V
2hJE3RqBgjjEEcWex20fmE29Qa2DWF5mApSFcj+L21TiFKW8gKr7w79mDYIfc6G0dPv8TP+L/sQU
iYFhsiGmmYRaEwXdnC+7tPI9t1p+fCC6oymmOBAFheKHE0RFRzHvtDtQTKpqQlWNT+z2WiAvh/Ae
ArMkPDos1z/n1722pzNRLV3S7QEQBSAOHLBf1RoXbT9+F8VAP1GtVJNtTyq/UVZ+Noa1SWYVR4Xo
rFJT17TmPqdpNZ6e2Xz2HjnMAcqfgPBcwYhyyFdfvhhPhHSShv6Qjdt39ViDJ7Sfomvmj2+71XcY
t+YXi0rYTtMtHurDlql5mmEzUUpKWqwi3/mIwWtwGugU9gkjVV0AqvNM3U0iFbtmy+MYi707NoF9
5cbXDjXm1HedfsOYdLiNGzeZjVwcMu3JifQbrfQRKYHd6E3bSA4fZdsyov3UgiZkvHS6kErwuCe0
3SRBjaRmffEDKmDUB3yA6lut326L7zaGZ89mw7J11101W1Ork2fcfVxig0tfthHRv6l/gtG1tagA
BGYAh9V3cLFVhe/LvQYhNYGUTt/RpQli7kTKEjoWU5dP59hh4D6UWy67zQyRnXH/MJf/L/uCb1fO
FC8jTAH8nhLzbt9i8nDk3ahNFgHkugrqOExMSGOYJDTRvRqee6whyyg8gtnhV2h9OUHCi5+jyJGS
3I5L+4ky43uPKPdAated+zU7WKH+tx04fQdE+R2kdA6QLN5L42bvqRut+teeSFU+CZ1DBtiQrcgO
eWFCw4B2BlOuJb07DnvTUNXUuyRdPQbUSsaMznp6LNh2suzNbEOek4oP2cOGGoC94OJHVab3hUVw
Wk8tAWA70xQfnYznMP9eIZvLxd5gfgfG/lZwJX/gKgy7OpkAqmFdYVP2SQdb4rU8I00FS1IWSItD
bFlEEEYV6TF+iTNpQrTzoQZvm+pCE49eJN1tJyvQPj797ors7xjEw1+sF9A8Q6lLMlocfegFFHeM
aYdrMv0s9ai8cVC495EVRzD1545A1l50cDb7FDJ/vZ0rC/J6L1NSK720hSc3DDKfwvKwIDgGgGwv
dzoPqRCesNlYwGqR2p0saffJMI7qTrv7u8y+XSIs6kfGCNbLLKyJkrQcCQfWVXrZvVp7ZzFY6C6n
jIMsLUlC1PfIcilmzY6HPc8zAT6jRfR/Zd2xL8lviJJ66eG0tCFg3dvVkwHOa4SKJDBZBBXW6XEE
vaoPExVYAfgsq1CilnZ/vGxgNBZn/DYFU7Hnq1e3D+bnxTE9uUfx/yn+s6PgBjgZtxwFN+i/y88s
eL6TMvugDJUXHa/AZDKnYK0+9IMxlIgl50eUFTHCJeWlNOyU0cYd3pIlQ2N4C1VPoP1rBfCaSr/3
3B+qNIZNd3vRoPA7f8Jt4+vB+0nIkaHMRZmI/g94wwh/GWjNTXCpBPQIfmNncsOEcGBMeLF+6CZv
1uqSZsGdnfRBmCs29gLALRxxtYH1I8xTSJt+FI1jJ6RlPk5IOcPGVH9yGwpI4avF21zJ/1yT1Uh9
aRb5HM7ypKi5sLCChAZ0eXwH+0+jQPsYNVOINzeAPc1i/VrqIGWX8nzCu8TCLcirdbPhzc78E99O
/lwv803///uMAv1FCsHK9EqEkVjwD64YNQFIUzJ1D7ACBERJhp0LIVoc8BB0YN+4zViSOmYAkoxW
/k+8lbj7rrp6O4jnpKfWlMGWdHpyTvXQrqXqgbd0gaQvXGq7iOb/QMw/Fq/lHIVvvT0XAhKXdrEr
z9Inr7ozdQfZ2zt6HSv9kY7JMyb2PUAzFvkjAy8UM5GmiHGdhLHXA0igypWZIxOKLSNcVZvEjcQs
zZDrRODWGlmWwJsUYXvxIEFxDWDd6dGDSXrtAcK3TUddjzaVByJzKRFsgCn2wMzL4VuT0p7x49Rj
G3G7Rp6UkdnQuvVNWr1UG5nAuySPw7KOgF3pTmW10ts0BPDYTYpiO9DMCeiyAMUQ8aHiUih07X6q
CxFdnCrelhJK6l99EpktKKkzKv8eQzhJToEXtiaj2dr4ydPa3C0aGeTTLwrHco/reOzUXqnzd9dW
Joww4jY2tDdjgVizuWlm+JKsndrC0teUzWLpdkdrUS3rhzjl+vMvj1inB5JbLCjWG2QNlCg/U61F
opTzlmQ2EfyOS23c7f4ULg7rvPR+Iw68nbftMZ2t6JjE3Cd9G9Y8vJmqYTBhpTDI/Bu6zpBbe+1d
zYz0zOQcNL8DsOXjswx6dmcewFVHm2CuWAx7Nr+4FoH5aHpXBy94HsdiHaUW6VbnLo5Nz74Gm1Ku
mXwwSCMkedSuqd1zRcdZhSgtCMzT/wY76nC9QDVUXo1HVzhWqSZcMSzfX/y3Efa55B1DwBV8JLay
F04SA5+J40btEjyk226AHmhxjV5swAqtZkVrPLHfRTITt50CFBkJ0kEsCAqYh8J0Gm6lxZl+hFEB
a7bOWqZBN8W7CKh917zjPO1WMAZBx1MACFixMerqAlzQGpKvFlJKCUA30aAlT55dpJXEyfohHHxt
acJ8DBiL3lhiV+tXWE7VtCGXt+u6ICks2OMBvnYUbI6DUP8aQj+t/HhX8dA6wQaaplANjJCeslHV
IBzr7HIPE2E5mmKboh2PDM81GqoxQ6dFEsxx4t24jDEys39mV4fbW8sJaZu/SulN/N7pB7zUwdwQ
pMUwI+CnM9RSjjf2hL+cvmk4fM0IID6RttiEXg2KeRDHWD8KsJWaoIQPq20uSqbMpP8rBNnJ3cZ8
tUr37FitmdRnpHKnErGNyP8gwh21X4KxjKwPx6B2roSvQGl/FLwUtCG7fc41uQ1Sbz5BIs47RRhh
VliQKeqVlCFpalS/S0A/2C0vzpr22Dm7yX2ivRnS4DP3LXSRXdl4VqusgXRrYOI4a4EW/bQM/VGx
WtiJT1QmxsDkQlt1qSvLgmHx/RVeKc/AJR7EaEHutZDdanVN3TapBoFaKPQjOuUXDh+206DZdt7g
Mt21qbgdfo1oGmdH4NcT8She4DiNW49PScXtQq/zr4xOlEdGDvNUAtz6Oww4EtjJKbU0MU695zoF
4lFXn3HiwmuxWl5Mk7JPBX4cd0XpAoyfdT1b47CQ5ZIm/QSKSdJaBvLaqzjJx2lf4ZQoMB9UUUW0
kztHjvs9m5fBOlA5CLoiWmkJjO7Rak2V1DxPOlM5yJW3LMqhPBH6wHHOE/YRovY/5Fup1hhwlVIU
ShemzLP6n34NyNw8e1KU+XpKLVBOT6xHQyx7FU7IG6ssIZ4nspP2v2R35yuvPUdoub3r/3AynDS9
m+/Kv3MrN4yC8So6W5lRNYuc+EJGzksDp8Y/gwDiHVUgWz8nBzx32csAtlsC9Ov+FCdx0E18076H
/g9XfOp0TrZx2vYFmg3EG7xytV1MP7xYzq0nOVQBn71gokttLF0pQIkfd1jL1wDvmdYglpHPZcx7
eVOBUvU44XPphcD6/rt65it1mPfxexwhWmdSc2CK0VK3nci80hAXMYrG3Z+g0IPLyBFloBY+i3gj
rBzZBsZEUAsxFKcEd6vN/p1iXa1pYA/BO/C0La+D5cSqIXH4in6cg+8Pg1Y9r+iPG8rDmWQYAB9k
PQ8fyCtklNSy4JI5bJBJ1iiyO6GUSV+sjDrzDI7zPiT+vs6TPPokZt1esOczo5xddaSoQn18P48P
tKpHV2BEFlqF0v2XQ5eVXC1teEIeTho7YkgrmE+CJ8XBDAvdmEj3wNA+4XqhMH6Y/M4NZOTsJ7cM
jlfuRvir+HvZiWpYhwoFZxT1gQualxHZs9h96iUkGuzhQB8zsUIdbyjtmvbla9uSDvk9EJzs8Y1k
PKhye42bbgSprXlWrN/+Drj8HyNMC+qdGAWaOFqvefwRYiaI7v7I0FONAwbU1CK+JpdvWz36mSTV
SIqrkVD87ggh3tCW3oFYoU61Gv0T73MxGz2DTVTTburT1ucRy1vqJnLXJTJpq5s4LZoOj4OnNbgi
NMwftl+BQTUE7fGeDllSkwXuB19quH8zT2c0mYxnxE+cRfKOuklS5r6W2LkKgngqi4mMUVoZtCN5
easa4ETNYYCCaL7agF6oe8AhNn5n495QzMeTPy8XeOiBjOS2vBt+rA0W5shyceJaWDEOIuClNWW/
QSEA5k1jbGaPA2RBAsbLuTPECE3pzdaXeSRW7hPlyy3qHrwhCHfPvmA2CO8fh12p9JROA8zfYfbU
ZLBcugIkf6Sk6/svKcftEyabq7pJaFopHvkRrwfCch1vdSvEf0utXsocYj7YnWVfQaFD+ff7ww66
oEHYuIx6b1be+j4aSFabBsFP/oG8zQD5+XQONEWpBJvONchNzb+6VyrCA4L4BlPdYLjQWLMw/7TO
P+T3dC55qFFKR3KiCg+noGpCC0Qqm/LUY/sU6BEZkNb0kQlcBazlTCBn1Am8zknSggh8pYmbi80h
rOjK4LrZps/ycne+jzrATQxqol090DHPOOwg7ZkcsqFMusd1L2/nIUf0yQlSyhQNX293b1qWtJoL
c92/sBed2aDrGFqhpiOj8vjERSWxMGuMYpi2Tut8OKm2Vd8VFxaKXnasevrjJxRCDNKq1/dx69lx
wUEPQyGNKtAcVlYEhVoClujqw4foT019e5CVw+5pD0zFV2GypISxQh1mhLa2cE5f+Ej7zCsxS88U
RKZfZ5s53cfndGzFye9cWni/z9hSvV59/uUv5veL4CwCHVDHWJrusJjA7d9r84OI4XvBKwEBt6OR
g5xrLPKVMcyM49ncO/LJKUlPw4xuu8beM2IliXAAAmkL6tgT8ca+K8CHY0U7pZoKq7IAZFychELE
vp+xjZmBVqN6eB1/umEk5kssLRxpTnxF6zxX46v6+nVgsc51eho/wo0g0zZ5SfhoBPg+bZdRndtd
5Bx6ETFJdcWS81PaYZQk1MkTL4c9D8+nA8goSK7jJx3guqepGnucvy7MS8cX4VyDMlzUIoj5U036
D9Y5r9VRPboocbRXDt9JyfDeJYJvZisjZvaomUq08y36eAx1xXa1tI4QRjGvekyE3FBnrQ09M6rU
/FvuqFH5BV4M8KhxWuNab3fORUotvsY6jcixnCg77QxlSbtzXl3/VaS02kneDyLm79YgKw2tOQC4
rc5mb6KXAoEMs0KdZ2tMXhdyD39LpA6OLYP2Ff///Du7GL3pN22TGOAkz7YVxXls8gLCEBx25jby
JJT5c9Zve4sZlevZfpCpvLOlJv22UyefeFsOpVMyNEnV4MquiAcutFCujo34LuNdK7qex11xw1+h
qyktYGxhi5k00LFckHmSjXD/XCzpiI6br1QOBzEviqlPLfhuSmhefYFW2B5CNVZn1Z+5eALCBZ4J
CPa4tJDXNNOU9KZhTptjanGTY3Afd4nJotI2Kk5PqaOYQZxSNgfJHXjIsHjxbDNMCHm44KtG55Bn
DLtTJD/AFqj4LeH2SuwsN1DkNLD+o0cpgetI1sJzcRstKuCT6gs6LXpv2o8lhwJk42AdPfKkeOJ5
83B52P1t/EHDS/o24YgrA4e1bcVCLhrVb/D2qRHc5P25J12Scwdwv1UmlkbXqpMl4ubVVwOsX4A9
72rtFrZMXe1ti3Fj1se5jpiLyrFEdzqAwd0N3xBxJFzTOPTl7tsDf/IzJ9yszRsPKXEwWawc8n1W
qVDZJwJiIMRBA+TTzUGDjzfVXs89+vIX51FPNj5lHi7P8hufDU1MJmeBnGkpOJ9dVuBUrRBBXb1O
y9ttzXtYWhzxTKIDagNqu89k8kUEPuQmZb5M3p10pvLeoutO7Zj7l6N8KKY4NQXSYnVVbhDB23lZ
1cxPVCIiicRNSuNw1wXxepv+8DfjS17SW+7A8txhbyKnIwB4KE5b3S35JPnudyc6YuBUNtsnySUv
Cx2TA8dj7qjbhfnWi93v7nulFIVogDJPmRWcRRSDlYvAPBTxb7lPDwbYkrzK7JhrbjvFliw7TKvu
1+NEJAcQvPbRNwsTN/bK0H1MoGXZu7CbuNk21c7Vn59D7SGQ2k9WrupFYX7c7fsvoCl1Q/6fTkwo
DRMoVahNacVUEO7C0IwX8f18hiBbqLIHXQeBnyjJcs09B6xt/mTP1tG1UGi6c4n15LuT2p2xPDLp
wbtaCnFehbahkiz8ekh59vfmG2kl6jZEWyPf+0Nw9LgbXKYFGviQhN3XoD0lNAP1Uy2lulLjZShh
5urwfqvFi2K+OA6eC7NdWNT4tY7aMEUJLiMdMGKLDnkX2GrsmPZaVFW2P3X6g0hHAJgYBVH1ojGP
zwb5YPbGzaT0AH0ROjb3T/avf7q0LgDvQGUlGfzZQgi/8yy4qMQGPothYWi89g6x4yQA/wC7R5FC
p6pqIrCRQXHdvTBqXeBV5KfsvCorvnz3lZ+nUKA0w41H1os4W/N1C/eaDXkoXDEV3+eKS76vRe19
hWOCUG6+U9TFsKh5pq+inXcf9VqVbtTPcwTUY/sNUka13Z0flEyooe2lZ/GneC/+a5LkkwdaAJQc
JkjXz116AhvLVCjwVogFMDkdVMo6rmaOBTVotdcO3YM+JlJLL7byNOcdaxQXqNZnESMxNgSRJiwq
8SWH4ZXaf6kHHezd0szEU66gD2IHHJQWEXJzpy7cluXGrrOzCMQqZ0PitAzrI+08W9+V8jfYdLRh
szF3fpHyrfC8mRFL1rTwZC4W/XmGv8jGjvNQJK0vm9I8BiZQaW9mzBE4OnH8S5qEaHDCKBfSyr2w
CFb8fGopSAZWx/PfS8feslJcFn8xqYxFImPseiiivwBt7DnyYi7v/sbsNZ7myzVkUuVO0THb2EW8
/8IDcOFc5h3Y3RpOkAxk0bNpVZ9/nuZ1lUhI6hhRHrpwOrTifZWVCYtoJamg7tsO1R8ybIk6lb7q
tLfaE8aCTdO6RKp8uTkfWKBV2buY41EsO4LQg6SZeEfrpCyzMY+VbnIXnET4/RrGFJpgzpQmFm3+
hOS2O/pwit6rBoiJNvExI73a0lpG3QanMaDSzwG6Y/SOkdV2lkWviURDeYWu4w+I3QK8JsgNfW4K
tOfvzC7xVufPdGUEjMasK+UrxrKNNqaMel2uAbrnyVflDL+MitrWnYdjWU6+LVURvHs+9hBBmsHA
qQxcwx7yyndL50CMi96ApkkJicyHty0dO+MCFueNDzJiN6dl3yaosYqihy/Lj7uZD9UHwpjD5Izu
y3rX4cgLCM6nikW0TAYnBk2FtgjQhNCc8BePfViEDkT+qZ/4DEkqihKr9+XTazgGQYCw3ZWYBhbu
gzZeJFfBntHJI+N4Ym7pEdi7v1MyefCMkndepnllSIELWiRs1Y74+b9RHNOSDC6URTpjzWtoKdHX
u5ayZiQ8qa2xN4sf/OIyOwkpXl45nzG1NAZTymvFgtjwNjzPpB2aUIeoLLEMwuk2BNQa0/wvxjda
WVi4HgIO/UwWUesyG8/OVo5HZvs7tECfzpwMWmi/JaNcC3uR2x7+Y5MYZiMe+oO4ZJ487a9s6NMB
+W5q4TH8nMnKZP3lFjVK3gGpGjJl32jFL9dI+4PRNKFyrewHb24LKKy+7CHTgHxXzORptcMgcao9
kebIsqGJi+zJxrxvuRls+CcgSZVtN0paAyiiM7ia7Y1qXENv6bKAgL+psKnlHsfgtoXNimvOfs/1
EwKc+SANFOrLBKrAu95o2kb9y1hwPFYhnJT7E3OyWDyfcJAvkC1q2T6fW2Ep7xXuYkQDt6YNMhzc
n+apQ16nPoRa7RO18o3Dx1ph99Y+xVrdiwtPKgxib51zMrFD/XQ3o4TFypU+SajBNb7/24WYgPrV
el4kT1iCatadyxhynmw/j1ISFGJILxpyUlspXOqUvhuO/dAKJ11NTbF/3W08SqxQn/Uw+xMyTLgc
RGkBw5ex4Xg2+zz+kQB+L192GnvAKRXZtZhXXb8SHODONQF6Bo4GQE35iXD8EOlYzV0vy707gdL0
3xQqTfgkkrX1BSeGlUW/FVz7KS4U9l7iBJoRKhDQ8NQFenK42driAUwn3gqvMle9VeCtdGfjvZ/Y
PyCebdEH7u5XjS1xg6pL1QosCU0FjgfIBqI+XbIbwWUoWhg9EH+sPjT1mP40/CPkqzdoioJ4LLkp
otecy6UuEQTWfG8+A60ZiaUbpNquL+OpHwejUJbjzPS4qImhMEyKHZmQITqGPdO/vRiF5RoAsaCm
QJ6nzx9ewEAdk7mwVTdG77RhUv9gU3yTJuqLW38g1hGMGKj6vkNgNAxGpS+iDZ0Mrxy8GQ0l+Zjf
MYUvhpyum0vhkA+oW1FN8MxI4RjG0VM5kuTxCVNPeO4i80rcX+J6JBZPBYnsdhyLGfS21aEREA4D
Q4xuHGwwfihhiUq5XxgPd8C02mW5MSF3I4+8jAZWQSSg36o+TYk+epEEBRFmvyTtsGk563ahgI17
DIUcv25CjJTJkkcqSqWePHn0FEcpD126F/rICvNfdpUC6K+RtNnLWy6JF/0gme7nFmQ5FIaKKlRt
aCy7/RcfZTSHZr/3ho+G1zPrtnPB8Wv6u0Y3Aw/4GBSF4dRPvYgWx5Oc1fg7vH4o+l7qaoidBTuN
Cu/cs1uCQqp72ZFst1GY18rpL1rZt7kfpSqpovivB5pXl8wJJ2TtbHWDdO6/hTemCdDKtr/zjiwv
W+CDfCgbs58jsRLE+eWo4BtrzJl8e4kGFlHAA+YzdGX3rTL+6aLxtJhSg6FxMT7r+gKX1bj+55S5
3A2oiL03/LQGac+796lhioEjTORVB346n9tBMX16BXp9Iq7Ia0GRni/cRjcJu2Nk7qeQA7cs1g6h
2qU/4CrpWT8IbmU3x/Rx8rrtuU4T9OFekhtTm+ykKTjYCmtv7kOexWx77mA/2qQlOcf+VApS5M/G
Qd66FMmsmb2ZEPDHGmkoi+MLOTNdKRHGo0bhLgUc6LDd12F0cKNU2gxX7ey/wE4cOxizlaNRuDWp
BskoNsd/g0BP8nUnShnwcUjpNfeeEy68hDSOGDPazRKSu7PZpQkHwnwk0XIRrNdzIX4erqPsq9Ly
tqc8+8Keft8BwHzpPKi5ZpJcfiVsyFHrcgKyBcg6S29BuO7MfcVqpruBdR2tfE2dgU/dcJAlQ1BT
f+i20mTSr7Bbz0m7D6OZTYAHsN46kXtcqlf3slYfKH9PYCWLbO1b2hYX7ORemaERd2yN0ROehuo0
T48Ks19mblLpJOwWu2+yLIuMOX68T131ErQTY6qiHQqt+nAO+vz+w8su6E7UJCv9+NhjURzMecan
73hq5QFjVCLHHN+mGw52EzaGYbVBLHG4zC13rJPx5ynd4jQ+rRkgY4tF0pML0OmwFU9dAN7K/o5h
SJ2cSJ7EPy8EDE3CSJ5zmiWFZZyuYRYrtSIPwrpu/d3IJr10GEfMkpRJeyAJ84xkz9PpazIsSpHZ
dSOoQIxS2Aow5z75qfK+IOHy0xHBkEt5wRZki3dGL3G7WZ0lxuQ6EGKirVLqZSqDoYTc4eTf+RJ3
tR/HFuHVpO+s9UpiRkuQP5BWBWoNFx1DrOUGP4CaH2RBT4N7IKRg8nwHy3RqCLxoyXozeIxsIej+
2CoyOQXzbREVESztN6EinK2mh2DoEbzu10ccTKW5Btbnhqj5/1Q0JFWD8E3SM3i0jUwg6HMvT2ep
MlEskGUePty2qcg0j7QRFJMCP2BLhO1tEogEp6pw044GMRUYu+8L/vNAcFHyZ7gBSVNDo166LKZY
3OkkfP4LuV22fn34BTyHUQfNhez8LPMP9d0HqgwFZ8jetgBAEYKp8fLt7GVwa9ZuPdxNeZDFOWai
pW+3KbrumACMVMEsTkvJk5TtRvNZFPqGZI2cVcq9aKcHbSJOVlRYzu18aijA6FoMhaASlOXa4AcX
7h+5xTuf4uUTwqvyypPsOhgWIDU0EShQ9YePkEyCF6XwQ+KKWYwP8cKumCnmkruGUiZm1ELrpWW/
bIr4grLBajt/f16E/Vcnrvca9Mbsb/PrEkAQMi1cyUngHRSW1UcIt4uQX4vhx330NksLSLuHPryG
TQ2sqjd8vzA/Fh+Xs+I/0jmSgZ+Pcwz1y68E9jm5VaZVoqShVku/Wxp0/pbs7qGfNseokpP5hvh6
f1mmQ/WFJM850MZClZTjIz1fc+HqV9UkL6d9qR0CW9LYrfHtd2LGoWc94HZA6NY6qbB1UiwEjkNF
uPcQF1R50nMwCtMCqcNX8Gk5VYjEKYArxMwSUcom8VxFPjPY+P66vMO8HDX3xJ0KrpIHPg6Uub7m
aiHo4ATHxhdaBaExCl9CPlmYh8elf8uwcbxUYdvqFljU9xzsx6dVix3bc+Uwse+zxzgMCS9yYicG
nUsVMpqeRSV7pOeUTqBvD0FsCtAndvNXzG6ftvpTw7VuUiTuIWr61SK6ty/FebINHoOGpZPtKIq6
q6DFRbL8IPjYZG82rF5xsSAwYu8m2DJrkapWQsZmAoyQSLBGpq5+1HCOqJiIZzNr/7fCXREtg/iM
lxHQBbQ9TtNa7v9h/98e0t0pyc5sFo98nTA4PZZQvPyByVHyHa6EFv5f0SgKVzrnRdmN3TDcoZ8Y
n1QsC8lMsuHMjgXbkOEmYfMyvVyq3/ytLgLmuFO7ZciF3/dSa3+1CQMz/nEAxRBE3sWSEQ3EtyQP
n1qzeCEkldOd3r3cc+AQAPAHR6/q/TJm5fFhhRdDzPvyuZRjMxfT+PTIjIjz5wCPWrZIsM5lk5R8
GuC7hW90LZYPhadSrHLGdPNkXQQ/vLTtrR2F7IbKutzmfHBlpLcfY3aGsHEwwWSlTMcFkbnH9Pcr
qx0FJK0TG5I7Pg4QmLw+z4voTv7HXigeqCE65rsW6qy6RVZmzR1IOVHS52NwDBWgzF59j8BPBI7f
t16TPrBlwejVkUs8QdpUJhlxUzc82Q+KAPGE1RP8FvxKcWI5N/S0goS46djVRYHo9oPNzq7aKEKl
/KT8wTcwTS7ToyINRsSDsSQmDFnHPfZewUCVK1Hio7ajOCd6WQr6Dd5RPMuZcFirRcqotIp+tnl6
4UPC0rvAr2g2fvLwKGs3wrRLXqvUNHLXK4BqPpqHKglFZTxsvMvhfjQjDJrCAlFpnKe0/vo2WcVn
4M0v2gr9ueYs9u/s9fJoAaFnm5mbqBc3O9Djth+FEiDWgitsomx2gwEa/SZQ/RZfJc/b6vLND6nb
3okyTMRu+ppFE+ThCfXP4eNxqhMzl6bP2XmBg04WVKbIxziJw03qhZnO3rpv0pfWu2UHUCjwPDY2
nD31gUQP9T9H4mCiYlpbbUAzGoJmlRB44bEsO4KUILw5SpVUlFu1HHAYaOEqa3Yh5Fby5Dt87F6w
iGVGrrAk9Ux43fxMrZUqCzOdA7vO0HmBMut/DXS28GNwD5qYdCZz9x+4jSA6jU4q2PDDLfg8gzdf
824Z3l5G/E7Dbl9MnmWCi/KuFtFZ+BKlUdcNU1eKn137QKxsYdNPY+y5HhituZ/yMNzvF6sDn8t6
cjVLIV1oFMSK0RGOaEnckV6fwTEXR1RtDqXrjeJcKNTQ4oEJzFReb+tAoG5pcL3r0p1ttjQTgVkU
J9toLnRwvvnJhO8JBwA+LVfKHSER/jC4zL1mbEfBEtgIvghthdI2pVUWJk3FEYgtQQiH6jr+sbEg
rxZOoEsQqrtS/7abXDs56UQ2DgQ9fY8cV6n7w6FMgjfXpKp6q5hhTD5nrfTE/hMQxyLl0pO4yBrq
BqWA8jOob90uvhPyf8ri8ESA0yLul5n9bhZsfw/3zA2tIDnkdLiU3DrQ9QFXtIV6BKJW2fi0YBul
a8/aDliiusLE5l9H7nixkamxwElygRZme7ZpkkPsArmow8b2FMr09o4QRukTKwy2Ue241fhi5qig
zdYMnk7uEbhDeqK7tyeKjXemiyWMuQM9tkADg+pf6PfxlZZHiOkEx+8t69UID5QYfGl969KTRE5p
DxoHWKOyXIWw94TpK5S8b3GegAPr2Dfcrhebsbny/u/dth5uT36m1Yk1/SUL2RhCG5PcLA87eQZ+
F6Vni70Gc+7x+tED0B/rd5DMA07mv4wKlQMCtKBaV2NqYgCUZcJ0PTllF7/7lUhr69EbHOYYBz0c
OFCtFBpK/6/tPaps0WMw8kpuM0F6pL/ASkRVr6xZ2UrPUXpPsYB0XdVlSzCVC7X6ngC7vkKd3gdi
V0L1EgN5hr8GvgYhsQiuQ6oCGwRJvRC8GnrtzVGUbX2UzfTgnKkJAg5cQm6SVYVur7751dc9ga+I
O+ei+/BlgSJFeTcECCoDZjGq4fGh9ck9mR29ubE8qPJrhGQoNH3CKfs0J/qxg8Em8SRFUMg9b2x2
2vfcGLnKdDd4ky8Dd4nba2JsBuOdqjhiMHetZ/k/znOh4Hd/qoga46SqoIn9ErAXJ53q8kC2bQYz
4V7BFgxnXFbn9PbyaH/INZNJWdIDGWPrteVytg3bZzs7CFsSJD02qTOtHi+chd7mC3mDyX1LEjmP
UyJde+XgUl7PLdYo2yBM1gyzelqtHJCr/dHm0PJQjQcOgo7SmKn6PhzNaRZepWY6+dp0XKEYzWcT
gAUTarkb4jgHBHGLCDy6uOSOW/JIEj1JpJj7Y/FVxmZCOs5UyTDeRBtvbFtDIV+oQIhyppDrm3OM
yhIbEeVgq0wt54zpLimyvhykFjYjuoBDi56yJkj4zs9bZWXC/W9Am9W4c9sdZWlHcjpoyCyKkRTg
28QuxmFVW4Mb4RIHeiYSmlTW3gFl7syE8XBL/8zTZu2lxmKETyk9X1FpdGVUjGDm1a5Aovnm+aMd
OHn2cPUhtj0ngBfPOHrD7z53lTEo2Pi+QHZ7c2EYSLqrhUbqenBr4BnAqmyhc3UgapSVe8f+rAvT
2Bb/UrDB+2ArLdHPn84wjt3q0JadHS08/t8yxZ+6KZKxSbfWj8QT8C24bqLlNh8beq+XouSfFe6O
IdXFvFHQ53Oh3vxBPqog6fd5kWVr48dAQ+1qHLFAwknVnvF4cQbN2OgNadG1ArIzeULiwFMeCHJr
Dl6LQ4OXe9A8QWZjutMgIPfFw97JJRoF5oM5kJ4xdAzWdR0xiVN7EIpAhmn/KSRBa0VjGGF4kEiR
+AGdvNirygK43viXzQ5vQLEWvs23WzJBOlTE9SBYpDQIZ7uTca0NAMEYAQJtO0HZGBevh/mXZwUQ
L6iEB0WuY4yh/TbMMjODXmSvwGAzmAN3tIqo+ZpyF/6LTxjT7lBdPUpuReb2WlC1gtp93OqH+HG9
GWY6f7R+9CT3mczBdLOPmSRfmwRNrl9sq8GrEwWOPfAr3ZeyynqCsDO3PvU2oFypJxB29AgOXcUG
aTBcFQp3DCOWYkoSM9K28FSTCKLI/tjznQSXgPMgMNj6U4w87THGMjKsYR7shJsYrlghUpgsphF5
ZloL4Ar2iD79+eCn8O8cBSIXE5Tuc1/LE+9MqedCE/6/HaTRiZPLkTmNZAsNu65+FrSfV5r3xFhq
YONoaQ5xFAvseSyY/xOVePHV/6ydJSkjVOif9d5561WYEEOlDi4GKIYXO3CZFYMO0e+gsCJzHSaW
baofCL3Ia/+54D6sKt+bJ6Q12xp174QdsXd+uPdnE2UWbccskW4I+/1tUxnjKWRn8TT3DYP87g2F
Jyqdhm2pVaWxvXiZZzLctuRgXNC1lHJ8FgHDWXTnkBpPAYBAabpN6HxUv1JlW68KZC+LQsze4+xc
aaexQ4dz03r7EuSxQyedOpT6vAdKBEwviedkGxsG/u7evi9vPLiRN1kOclTuXaC1KwUJvNHX2Tyj
mGZ8BKosltJ/ZTUiL9dGDjBnDglGrakSugjD98Q8/VlXqdHiUqg2NqdDupF6zAonhFs3En18Dokp
cPoZJXQk+qMmT4YQawre+ZX59tiOD6bAHhHElYDI0OeIZb8cIE1ZfQJNPjI+cGtIYrWRzr+KdOB8
mWJRr4qAWqhe9LXM2G0P9kvbVVVAfALL2Tif0f3sETx8HuzANovkKuU1YWox3mWwF3AWFoFEk10C
jXGFTu90Iae5L4kpDXr30hWlKDR/slojg5PLT6+EUishV44t9k612QVaZCkfFDkrA2+UEdc3Y3S9
VqaTYNXX6ORWGVaoGYE6ciGwhErCgZ//yn+zsvs0FUgNv6Ife0EehS5Rf2VvQl3NQ7kV4tStY1E0
eysuy24/ay3juOQPkTCx2kTRRIoMbov9X69ONOtd4R0CwPbseU2UuFYW9v7IA4Bixxv0AEjg+KDm
kVV4/472WdgZKOL+jsvPuqaY/VEDEnBTC1Yq4xAwyJIPiGHG2vrRNMmSY3ir+cXsD+UCA2b8YO/Y
YQAhaERcuHJ9vz5G7hj3AV1cu/qMJFYz261khWp2gs5Jdffxgn2ZwoRF0OPcaE7dsNGrrj3X4Bya
wi7zp7Y08OWd+1/bgfixO2KKO/mmygbagZiljVagEoD4QiqiCQSrDdvwI86cNkCVGzz6tG5cIhWb
iUdbCAORz/ZUh6EtqALc6IZuqzyGRnjjwFUmVn6/d+Ws315ZOZkwBlxFjIjgIPiqpWjBx2X8qYYc
lqkJ5QYqwo2VwQzmHAf4RMMgR1XPeQWVM/16wyslDjJITYet9NDz3oeOREwhG4n49kcsH7JKo7St
jb8uqTwVfM45Y3xVQdkkFV/J/P/3+FkBUrnMVJlDH+ONbzKwzX0vIt/bDxPOf0eBT6FCME5h3jsU
qLr5OlWS06AouboduYKh71D77ktPkFCUJJ7xrebp37sqW9+3XaYVizmfV0IlzluW4w6tdBW9TLkW
+u7AXGl/vB4NJqgn0CMiaKpAvcVkb2QMv1mQA3AQfMmkoBUcJRbfY/f8sMXpwGJzegYQ9R2+lqsx
kmj8TkC9J8ZA+BgLg+NvCo7oi+VtocQlgXCG+BZgQDIoj0JidgG/gK7xOFVgIsLkuhOtLsgRbGO5
eCNVgDZLJ/QX1jILD52ICQ2obZICNG6xARdF30oc7JKxxjSAMoDuMGK1AL5F9PnehkJl/kiNVdAI
GNMHoWy8qOq29reVfOsmhUykpAZl8CCWoB45QVkSZH0TLU1ALXO6YMk4O32xHab4h+wUdtRlWnGg
wDF253ISBqHiVjMphJwGv6JtV8WXRvf/UDm1kRkASCCor+CCtmobxUsoXRxQ5YKsU107OWJ4/O/f
F5WW/GlAkZwGRqYjtmZV8P3VEcUtWFaVDuaskaTGY4bsxIQr14ZSuiUztzBaL2aMhL5OkVluKrGF
iynPFNqOv4vRv2XMK8FM6XtLv3F46GWPly0B/KA8Oj4xMNp+Em7ywy+l9t3rGOVxd8lwHtGsZo34
O3e+q9iaSOv82L59UmhL+JzOJ44OjtXl3EFUXRtreuAWNOc8KsvB7Oucw6CF8u3Iwn+IKDZzrLpV
CIaw/TK8hGCKCgoCw3miioi0CNVsavbSVZL4cWK+hXfeXOJmTTVAv6kIpvZ8f+U/pHZ3EvUOe/FT
ELLO5wlovvkMeE/Lq0Od3RiEWDQgfB7TbuXHfd2JFysSRLVzQTaxb9HLumaPRlkzS+n2+aR2u00M
0Rjr/or47CXg75RF4OP3q9bt8o4e7sm0mW0VHNcff5QKCzmD2TOOmEzMlgaG6bvUw1UBzZTIO0di
f3p88i+T1IV7C4irCPZQzyJkTcPDnUN/zBOnT9fDxHHNoGKZC7quS6MkKSrTpo9G+ui1uV18e+WZ
NhJ9TtaeHDtYQazx6brvKVDj1grzoS2i/eNCL8G29G456/MucNcK5cC6FepOA/wn5TjqWz87f23l
xEcc+DnR/HmiPIRoCRXLWm7S6MeaUVsWRSEPN8VToxWHcd3DWnMyM0+22KAy3GPLzBgCWWUz8xX5
KpxVamnzztTm6N6pDXh+avFNTamGtTreSVDNGLYryLgrLsxcU+SwSm1M6wHla7PwUN2DM4fhSR5j
Ba1sj3Emaw2lOSLX/kvJD1d6iqc701LsOV0jvvpPXlBalS+mjV7xvnfHBz5YGFbHWl69grBpneif
9DNgVXrRXbG63UrWS7lYESeO0UzKczofWgdYWv4+3kZvKHu16+3rQ9Wsk1rma32/T3VnTFaFedTw
oxhUygxP17ScQi55TnOrOfSNnRN4mQRPOE7LdmDnVtsQt89/ctXlzk2XmhjVnc1H7eANTkPMrc1B
908jYZK93m4y7AUHNE1DPCQjlqNT1oBRbJ+hT+IE/IUZe47sd5a1RhkQC46M18pWIj4/1EwQo0ag
YkqEb+jh/GXh0o1KXmmCUJGaXBHBhOmj/H75/RfTGe+cR+9vS7Tzca5fmzWaLodNJG4acQM/fXVV
VMHhaGb+mEnGRLSw/xVwabfWvu8p2OjPzVq/CxEN8480RrJKiFc+sBubKLbfPozcUKY1hckTWj/h
mT7tPvsuZQkdh3IRrWM+T8eYHqfSyJ0tkr7XzfYRyVgyAZj5Offmq+t7V46Wi/YlzM6tTHkzb34z
VJF3y/5nhOLfm+WLdUb9630k/QzmwwdH6Vn9iWUo7sRseWsgZCE2FTruQ1wWUqx4/rNq2YPS/ydt
qDe0MgmMV1QMV7xwQs4Ai7ICS+9EosS5yvM8v2m+ehJeBPdZvS+JGd3Xyd9UuN5rBaAdRs147xxX
F795T9ufnTS667Q8S/ZO3cPoVPuxynAHu+kO7I+UQRfMsdcmD45cLYswnkn8n3xO/R1v/nZa6y68
+28v+GscexHxy2NZRxmsPXaCL7NzplJxF/Itih2TJLDxSMBUFOEbvUsbp5r7tdlxhK2VAPinAZFp
C+MYI8NqBIzCL0X0QwFKODR/2JTu0Z+Fg6P6pwlP/FfjFkByvM+FWTL3sOSMHG4YJMG4ONnC+hBo
bfz3maI9QniCIcFKYwphJ5o9Z6k/WhJ4G0iyy5Kc7bhvjfLr1A/zJks27seJrtegUKe8EAocouhb
pBUxrp3l9FI9iVlIrGk9pfme7LwG2qTN42zZMiiP9hDJeNCeEpxBJAsJonU12DMsIgCj2c9odxyx
3IY4iQA2ywxtlhH7Tx7+Ux8c6o3HxouOYaXLe06zd8kh88ulQBi7gr72ohMG+74WSJA9ACaA8M6Y
qAipES0bj6pyMc+gCVrSUgSyVBkvMKfuJjH5qeYfhNv1wwoaz4PSAKwsgFsp3GTmRE6ZRLRAt//x
v2/nbsPCZ00LsYclD78LCMT8w2NltGEJwk3IMRDzblaIHyOaYyvrjf4HOusDbQ7r2VaI2gjkE8ha
pmSjWW8ADgEDRnb8wwyp+SLb4zGGmhjCfoiELJgf6uvG1tcpag/0WRF5bvpGn5RCTjZkQ9NznU7b
lCuhXa5Xp6RivTAuo3hszK0FeFo1UmxlvSADU1La89/UI0f8yMb/FWhUnZ9Ux59PhWqIF1jSYByJ
2MgeaUII73OPQs3vPZdAK+IAAmmpTXGGpIu6F4Kt2jN+xmvZudErzuu4Eet5ni23FVUhwr1qZBi6
MK6uy/3q19E5fcAzvSCj2xkU2jBymwTJ6kixdNdhekT7xFERNYsQSel51QKwsNNqWLOKwInLn5lD
58vrwBoYkvco6oJ8tYY1Of2nMTVD/Nl6nWg54gIlwyCy3hYU3eJJVlFiKxzUa3hrWJ0LjZZKHDMO
bEpbxqqoXEKAioeTI0cFK/I6VEL3fTsxI2wk/kVXxHDlcv5aRgx1zam21lZ8HfT7SGsNdOiBkoC+
UiJNqW0KAEcUzZOZKnMkKionxpQmZThNLXQq7M3sBQcAgQUtRZFgSNQ9/X22+m4vtWbpkla9GjLJ
ub0wuOs2xt9zSdR/9G231ASufxevGNKfSfXB75kdpeReWvTI2iw9hGZvWWBMjOBw9TOUwJF8Wd3a
S7GJt4KwktvcFfRJ3ozOR0yc9yCMkYSXqdLsoJ0Dm4SyHRrc0aurpL6U8GFB174cyrzF20VNWZFF
v/CNdq76e+Ujtv+uSVIdALkqeH8i+drhfabocOXefXcIYJ1ph1R8w99Ow/4gfIz0F1iqo+bGIOIH
DBpDKzqXKHuP4UUHEf4qO+ZiMdGu9ISeDdAp7jOktYD1/FmOVMfeu6WbfZeN75M42342GbmjkPHh
fyF6IirBn8qhnYRNe7QrfCdGws8mEUvjeWV2y+5ds2Fofa6s4ljaF/W3hCaBJx4bTW+cDPS/JX6u
dZKMCSPa0i3G9EGE962grPQJ7InPl+XMM+Ctqb8yD3IzaeLzyknT+D3mdeVzSGduYQGRJnmFzBEu
4SfhlHjjDuOb+KGgIPcYDvVLK572XoFQXzLmFmKJV+ARwVRN0jlDSlsTgQawDMpJEPrHDiJh4SxS
ThvqQBb/EHwR5ahnhDQfzSM7nBMr+zVXIS3tXQs6iu04jYV7qy6mKHSJV7rcxPl8P3Lb+H4lvpmn
I+s3CRpiPuoob9PGWN8tmUFxeAqJxvJcRTdVM1XOkJjW+V0cFIRSKKlXyok/xtjpgJwQ5L0Qm7A4
Az1k28djxvHZhvcBPVkq4YvaTgJlT0VPMmLFjNI3o7k6Gk7O4k7x1qHN/cCdkE5PZKF/Il+G+RzF
XBDufQuNgI3XPHqJFmkPvt/yfmQQ5yRDeLMNdCr70TJ0bCjdhHGVyNsrjiwuDZOhVS3jciyqXcTQ
DrbLMcjAiOVeJcLCaUf2n6IuwPCG+nY5KNBgvNCE4OR0xyLDDFPkvHNqjPKsE/uN1X7glJ3CMtBg
k1SGiuijHTJGEB9ZGHbQqgart1snsKe+1/QzJPFq0aESipo0IVSr2OTMg+81C07sjpar6xBjs+YM
vS7Wy4KdPw1EWZdrRz8Af+hmrEr0oNz6C0dD9TsZQtOVoO6Xuvct9lovJZX6zQiQWXbrClLaUuUt
7A//nqQKEy8lVau8pEA647TnMtqldtmdZ5ryuCLtDiH3tgR4vul5AWGiQQ3jqLQk0f94knULoCG0
Bq0nENB3rGr8EgDQBT/pWUnBuHRGwkUvfrSwFXH4eP8Xdghly0kvi/bUtN2V75f1XxSCw2DLxT7r
sO68iJb2nvnjf5sJi2+CYyqv9lpOEpIntmOoP4VSgN45gWn03+1yXj17o9qyM1IIg+X9KGFhWXPB
w32U1qOwl3Cl8cf82ZAzKZq4hrtO39zghtclPgUweHKS/S9qMUDOLNCcCMaYrfaAsxROQrPt9ev0
QLurtB/7Bvi5yYzcsU/kI78rXQmIiRtknSKYczYChBpdeqZE4TQeNf1LgN5o4RbHZlkiPWFSSPum
JkMRQ6TOKYBmtvoq+upTPBgxXqpT7DHeeM3/9mClECD0qtxGT93Xc7UprJa46snPGaEpOsu4rMvz
jryRCZ/6wtYM4nEU+WfP6rTZHqEyqPlIXDuIBlhbe/kop0t95veSuIkPBf/qMJr78PntP3GXQRNF
IWKBRFZrawZZhBF4yXOH8UNbAts9S+udr4vDBk6z4hkcnbuKvMMPz+M018+qo3/2rzbtnYdVSAzQ
SMRgZIShge9dShUSrXGPL7+V92qbctH7lIJ1dqzDsIDZMOTrzSOAVu6VW7qk9H7wxdHXZkIN2jLx
kDQKC6uznKIM7uG+HlgzQQDbch1N05iqA4+TrE7nIRF1JGn+wnwA7aqFnrNBkmKY0s4vy6v9Ct8V
fjSvF9aFn+NpRWL6UmuGRWr2aWC+DK/ebrpq/zqA0KXzKCFwr2PaBnfp0rycbOz8hqeK6ZSkwsxZ
e68aVv2KVwnwrtM1yDg3lxfDyeCMFSE441jiVcEhj7c1Cf9QJecjOIV6fp0cB2Yg5oFelD30KpUy
2JdYcvu1B4NDeWpVyWHk3e4plAI8u7Eh2LD8aB2IwKLyHqsjCfMES/EzphJ3xN3dH7vJKW45EwwM
6cbb9ml7CgPBUWSumL818HZwEiKexziNAahuzgTl1I6LXWb75MTo/GrHSyQybmuINEE9ptcwgnn+
dqfNnXRXN6wwQX6KgM+U9IBzjdWo7nyvpjSx1AYX/bqNv3qrqrDlcLmTy25kBVNAoVEYZEGek17N
kWaURcAuiuDG27f8l8tBxV/b6v2WGf6kWNc/vmGD85zQ4U1D8LHqs3DroFVtVUo20/TkVJ/LlIMp
6vsgeQX6nRyCnjt0anmlFZIMicmBfwAaP2CZDlI879Ur9lTaQ5/d2Vrj9a2KgbJrMgF08nuKs2WU
JEPlESxm0HzHGlHVRd+pJoYqZFj2zaRfnCzNGjc5VY7N54xcHqKcCinXDv6JND42quinSQHP7JpD
wocHHHntX74auidWNVr5VgGZNMc2zdrEl8rnbF37qtaq2ksbRS3z7atz+LOKwmKdj0E+p5teeu3h
DOisLCCvANLWPrY2+edEa3TJIQEs6nNKmdKQngdumYX8Yd4mzs2ZX74RAqt4cb2dneyQ0A0fjqo2
3OBwg/yAMy9cd1OByY32W3oyKbCOD06LFc+DCmJN/HDiAXzSpQ/xuOE8NczxRe9HpfvBCrNuQxNz
eWoTc6ToL2JNQcnn405ejiKTGEtlnCEWHvlgCLWcXRYAC+KSskPTzLtTzEJczbDdkEyxFZP2Wfkw
qnBmMooNSzVPp+4J1g9RjtGmWgVM1Vpk9KmYRbtEklRQttg6+jz9dFJ57uVAsRWmTvGbTNlH/RRb
QOa9QHvg0Sh8bkqlIzwrIL53bSIIP8AUwrNZeBUe3/EPTN50xxrjf0F3K/vQkPbk5I2O5VymyFRS
hsJIv+WuteHz5QEOwGkvG5AbakRws8etc+jKqk3ZMqTlH+CiPlzzuNXb1nuSmlAS1rHTzy6Lpilx
xe2pfOZmc6zUoAkR9NrfmvVhopt5xrRLZyVka5zvlrJ0zp/r5hWLI/yMoKoel20Bu0coMTy5vt3d
yPIksqDu+wLvclhpZrIaG7v1L8ptu4Y2yJCub2Q/5pOX5aq9TFE7yhd60eQ48NuXA2aJWwCgo6Nw
eYhcLdAfJyjVSJ9e4u/bLSTJLJf7TDCgIabeUaTcNGi+DrFkiIfTnFTJo3Z5J+Gag5W5vD94jRAN
2pE0myJN1YqMFYu+s5V+hJT0x7qqFrMyoBUbcSTAjUYPNOcY+AaVu4GFWok1l4P8RrimivIYYF9F
Ycwih5qv7dJbzGV05lPF4DGX/8Pw1EOCjNC7rQC6fPYek+fS/+Im5kFBKFPUiGUqKBd+aO9+48J1
YNCJZqToOzCKc5QpKtnpeEwXtTs+n+ibqAnRSOyxT4cCHehdQ4kH8QwM1CBTnbSlJHsotdW1XBP9
RIl3MWJdj466v9CR3T5f+mqI/eBxVuAI1OMnE5SRIOLS1bK9TBd5Nog9tYB2qu+v30JYcsTpGPlC
1FkpYTtqWdKLcl2EuQ7lyXaKs2CdVQ+1gp4jprECHFqkNpJajy7hGnPNR5RwuUuOUYy4n5aZ1PtL
6Rdo7SRe6zR8qRZNJOMCjSxU09Ar/QxBERstZaYy0gSeBlaKXgpuvxc6ofUsok9QhzHKbLbhwe34
oCJFmEQPG6ZzH/a2yNo1+0t4SKJhBkvlAqjY0MfNvDpDx2zcU7BXYSB4mvjNzjZCCYd4m16Blp/J
EBMMBu/TkN33ChB0bYGUZUVBMLQfof2GEnKQengvZkry9fKA6VlSUurT8TiY39z9GzYWRLYOyHIU
ZfAjJ37yPG5+v24SYD+vFSFY5p9eJbKswnuKc+Ffj/GhjUP1fdVt/YO0xamura1T84fBux81UhJG
ZQFKO9X4gKWhJCzH3uvMSRVgezV/6oeNDEkeFF15nqdZsSmk1GztVxKXvOPv1s/vH6XbrDY/Ctgq
PxdDIqUpber1poa6xKlwyDs5bYEaZW5J+8ruUZGInb9x6QqrPrX/3QRzBrWUup/u9jBEs310B2MV
T/+LmyzN0bgvbGHH53u+Ogj1tZK7nzMo/rC7Iegst35CGXI50o8asbuz0Tp5M0Nl9l127AcAwka7
hI/TUfMRNn4liRsaMoLfgsjUT9GNnE6qUGZQ6/YhBkbX6Bb+6CZndg7Gs4tl+OLdejp2sIRaJvFr
MwK3y/IDnHujVDq/pMQBc9S+Jxhf2xfTg0qcDClpi8h/ZzJXEuxS0zwTbwME0aKozZhBS5ZhSV95
zst6nBwuGtVRr61uYjnzjhJ2IKU5W1z3fyo8RsFbHWQc+EdW9P2YjDNeM0QsY+/t9DUj4N/KKINU
EZp4iKAGKgOUduFpC7kMIqv/nqzwAH9/cV7HFNHkd/9hRMFP1tuwCXwScUviVXvBvMmHmVAXe4uU
tzg1n7kYrbsVTdmExQ1TtCZFxcJoSXyPiEhPI4PBc4MUm4/ySLxkNSUas6uSpO3Ms9AOOFCiKa89
TEH1L6APnR2c2Std9sOHr8spPuoMLHfYypmbbpLdY9EqpmYc/j+X/d+eAy225EhFIIwIiN0OaqKt
k83ezKASYWADQ6u6Rd67Xk4q0YPxD1Fkd8T6D2WUgbONR7SLFbsvft/bNJTNJ09qFjnCsL3KrR3r
6cyH/M8hToaun4sBRMd9NQZAX344UN5z7cE8NfYwws5G+lCNDNLxw0BlUvKKX57ig1NZ/mI3qHd0
piiNWZ1jeI6l2HRgAyyN0DVagTFXYqr7fSYe8r6jqgfG80U35FsVkUD0zwDY5DYGpZEnnEZtVRAw
nERu+J4WbaKebc9FjE/5kXZeQvJpcsoSadJ6eEDu7yO7MEnolTpyoZ5ooVjtoKLTzADEs5pd2p0J
Gg4eDAFg2gfnbe0Hxfaok7o58Rkwxz2cbFOjLdnAAX09uYuiI7UsFIvYd/umVbjBflZlXmeaMa8N
4na1hdom1lPim7yN4Yx/EbKCGP9HOAn3vwZy7uNSpVtniQa0SSWvVd+84ClN3Hl2EHvNes0ENs5t
nPtzCx3p5ZwTL8OnYL5QCa9U3oWZXEh7L1YTRLiLeui3bdd235Ix3xYtxb1xd16jpgYoRqSsgrM+
1f5lCx7TkperQ8ut2NPhLAD0bZuvr3lsWNF7LfdaTF4xDZl/685JAcbfliPRmcaYxpGjj3okFbEx
lFVqlZ6XWvLn0yaifUtah1AGGRViSwMpEjQVQ2j02CA82C65yuMePazs0XhRMBrGLDhJA2n3dS2w
0aMeNhxvroM/ud+oYJQbSpE+ps1xO+GswchpY8M4euoLWpkoLT3Xms2y7wzsvqpZL7JiCWfCpoJe
6LP9yQjK5HMXJcBMzGe3S8DGqmmTIcDkDodmx121RwvQNHyKpD2HVDWl9gsyI0vUaqony70JtTjw
EuLF8qMG1ma250KIZ6th0KvhlbafuTSXWKwRrAZVol/bk0e+6IRNGiD3XENyvRvkDoiN2KD1RD+2
/qageVzVqZ75tTpLidV3mxIaDKASZttnPyZ/KEB4gKD9qaj6Q9LVusp5+5VgVDkWI0giMkO9gW3U
F/wXyayXz9YYS+KbJ8rR9wKNOv3Qu8WZdjT3+uxZnI2r/pYZYzhzODPgX0sGS2yXH+E+t9+7DLWn
Udp+VwRsI7G9+5lRVBJ9FHzfT+3P1HtCTmZt5hPyeVB3CxL6MlRmH3lv5Ez50rRC9u4ytmMSZCo3
QbkDcOqdeHgQFkIh+op2aEey1CL4H/vRfKbly1Zjw0HPlrOwD6HGsAYuVlFrEx5tmspazxMwfyaH
8H2IFg1E3FqwrDeL54SRTOTCT75MRA1VTsq0xcyy3O17cfsoL/5F2xTxi1u0J0ZzsGyVSTHb3tjT
c+LklnqlbP5c3IYVmnYrxbtQlicrhu6LFYv9U4Fa7dlDDz0Q6P4tAeLzOP3MpBd8mMPEt1iqskK2
CB6nCxVXrol8Fx50tQ86ywkaSgXxk1N7swjiILfPhvrdVsbyljRftBM1EfmxyfKbQYkPvkAyH6nW
rjFon7rre5JI1xOTsRkVzamJnODv5TaHgB2scuf6tYl2KvIF6amrj31FFGuDpaisrsX8uoeJ7/1B
Tl29RBS+bcdFvkyN1QmCyJZe6G7DyLlq5291wnPzRGOcHVrAAtTeJ8mVbZ9hTZLiWhbloatCwuyl
MqP6N27dTNwX0a9TP0jLZTE+OiD1Q32iIDn/oOPfN+i2OhZzMm/lPE/ht3S6CLkeSGILTk1trIz0
KSkFJKObPrjbforvR/HxUDEq3dBQvsEhw1kK003H+HH4AUW+Acf+CBqIf/yZjaUzKsx6fiNG5o4k
rh66vHTWrMYfGQigT4qea7rT+A8bzmWiqSFH8ASMSAT1IyANgPcbzRMvg1mAG3jidI+o2MwSyTRi
IBD+P6n7WslvXBhuve1d8Wv5zRch1FMMDw5ERtyP6axLvE9/onLD5IfJCoYvHPB39ZQyE6qf4NO9
MDa96hslacHEKxw5Wl9j4QhXTUYXk09qwDl1fEWv8bnyrq7KAHe5PhXSa8Uz+dGHY7xcJlNiMRBa
oL8wzaSO/8M7KGzIoek798gHOgysaDaIAymM/XLQIE0sN9abMgIeg7HO4TJlHV/Lvrs4mr7deCt1
JXH6TdcTJXpsS2jgs18WsaMU9Jk3hVdmQRQVyyCif8+A3ARlkka/Gydbi5XatgQYz/6qgeyTxpmL
KIQlCOVzllZTTE9lCxzXECfPihy2n6WoD6i9DybipNMeMm6ulIBJ34ElhnDk3fDPJwJnvaJwR+RI
3quKqTFS16nNCbh0AGIqqUbiOQQPtDWVucaUVQAvHYZaSjNdJR6wcLsKp/yfHpC1gW4FjmghwzXG
oyQltn5eoEO+ZxHYPXTIfgsXnmMhVUM6X/8msTS/pXJsW6W5fHTZN4C6a4py7sPgLFyKNTw8Bjas
0jt+pw+ATFvtIngURm1AjDCpyaE8FamkcrTdi/tKCAt35VSlV4LI959tBhfDUtgvCG4lNPamWcjk
KMY+fkQGKXCZC91O/+8gFwAZTwIjK33gqQ7BCQJZxVeF8DiYQI3E79QogNGzgll9yy6xO1JpF+gt
M6MFYUSeE7+iYWkVPHdedQTnxKVnwis6zRNnPOFH5R8NWElNVMSNKO9t9F+/zsz2bL9KufTrLkN4
PmRrxSZzKEsQNy8WZzk3Ide5BHp8C7yFD7ANLOBXszElU9rjdtuST3fIz7GzHOUzHjpVp3zG948Z
jiakNvgPr3bni4kpBU5aEsYt0RG/gxqb+fsws//eXMtNlYyYjTVAKUmyEkXTGLjXCygcmlymvqFK
Q8I7/wZmxoGP5+ENCPc3eV+4iG9aSHT1Fsv4GLH8MhdXrM01mkGZpUwe5ISFybVY5K+uINFBwjQ8
f9xIbo9+aqDaBTvYIVKLcpqMdWhoSpZQdANiF5oY4HZ3WBLLpJ0x3HLRX/P5DYWKQdpk/ODNfyIt
TN4kTk8xkqKpyMwokHmRoZbPROtfte1vm/pQ5WqufO3Zp+oUnjL+P/XAAnrgtp7u+glBIunjJONv
lU3iqsVT7mFDQ4smlniaU7H8+m3Ep9R2/RmPHZY+9ZeCIF/oPdmIPvmakT1un8wqKD0AVqxLcGJb
VJxxSnU/1Kw7hkm3tiYeAXpncFJJ3NpWUrZQJgdR5WkdKcPtfgy5ZGh6HT5XQ/jaN/ltXqZfx7LA
NWSwcWA6VfMtHjzYvHFxs29ISJblqN7X1e4DSTzAmAWO+dT853GijY4IQkkUpIxvF5xZG4NxsNrg
dF7GyrxfxmX7idg2zFm/smiVuXHkYJe4SVvZaCY0pQ5fpLn0m8s/eT0kdH8TXQBbdpgfqTaYXO6x
Hz1ZlKbFs5bKZBMYqcAil7RVjQhoqqKwQWPrCYbzPguZLW9bxOlOBd6hIwp7/qizsf+LMz56qmqD
E8qQECg7xYQqWPNGo22ays9IETFzi1EA8cqb6Km22nyus01SPE2SgXJvFv4AphE/hObInmCaeUsF
2exJR8RJo0l0PdBJ8FQJm2Kza1NtTaAU1VB9JcDt8MQj2Ewp6oaJpWZ/38N7HJeY8PpW642ZuKfn
1HHy5FaJRcex+KJ2Pidv+0FTBepWqFSE8w1d11t3JcIYZwU7OiSp+dhCjO3ncCZ4YI20j2J02+gG
gkx2cqiwcg21n4N83Kj67PlIr7wnyftT42mcZJ+J7NvN415OYk0wrkDB3V4OWPs2SNpoC79wRMyA
tqFfT3udTIGUENtEuGSTURI7V12DRiRZVTTBHbbzdAkPsIwuxxqCK726ppWpqU5bESRLHjlgcucM
CTUPjBetntH9GkRbKq3KOAIU8DtDXAQoM0nYFWvDLa2memMBgpQdh6zaeglNf4GA/I+gM5BUp3Fs
eQaG2SqWf3pOyOVWjWBgpGMKobOlNJzct8NZ8DVDutW9dxLkBFG+Quo0TNiwTmJLKREU8oYMqMt1
7QSRXR85IhhuZRTvQagksQcF43aCtoCyRWqu+aX0Ktio951KBkiUU29+UI8iriXeu1XzjYB2zQHi
0PgotLGCLs8Wa0eq7YyuYKpHw9wCLZiDy2AFuOcY22Nvby+BeoCkyAsjOi6JdQhXL/1lZb2NPyHx
3itWX7CrdZFM7QwxCa599Kbzl6lzkgF8mAY6Um1HqCMbmjHalUiWHXf+DN6zZ8eilNTJZJPWnGuU
wdsi5KCNs2AiferYsYPWY1zlgkZczZNktw/skyWp4UTrIEVMyE8hY69WLnvKYAmbrfnvY9HdzMSm
tMjOj1r+hHv0305FcuZNtlWehzgYOrDeusissbtfTL8HngqzaaDuj5eaiYskHUi+o8TEWfXzNbRu
DU00JIey0Gb95RzPSrA7cD64+13h06RcJZLlVG+RH8JOtM6Q6LpMyd+I/JFOw0RLy9Oh5vWP3W3F
kMIyuQ4bht5PKzgRQa3kRKfK8ZLZdPP6goW7oSzDzBCNt3hkDbiMZlrr02xbyc4mka2zOO+HDKd7
+wne7Hx/ky/X2Ij4wZkzi6WAAPiuH6x63XiiBkA/1jfR9QF2k1v+zS7oVm3TfUnET3TuakFVgA2Q
1fig1TpbJ0Wi0Ig3+BE36iL3jt3gG+dgebNL/HiHqW5zxfsBhJUnRLJ+ps+kme8o7r38KyN9rlSs
XAwauKJM6cmAXya1k6qHM4FBKAWpe+jumywIyODM4rHe5uJAZX2Cn6c8c5cCFqiC/vmF5CilgHpG
CuJgKbD9K6An5KgjJe27EZX0Ov0LPMDvDMlyjCSKLPMTPRn4BLzMtlmdKfLsMN13zsq2Aeep/lOS
d9IPUOzQXtXLXi+hrio3Y7PpY8z3tlYouAkA89fbZ6oTN+VF807FgVN2ZEAu7JN1k+HLWjFHdb2L
zLXbjxeFEtmw/tIXFunMUlx/uyJDMQ6LC1OOBa3avek7aEbt6YcWeaV8tAvrCunxRLZX4zy8U5SJ
6/Nulhn6WDWB4NPen2dyUmfI8abF5i0j1b/F1E32aUcP/Dhm8rKsw+Pc+zXIJo+XAav2WXACkUjo
8n5nrOEEVfMgDHSXmJCj7LA9OXfnEfv/aGI/aPy2YMM5+xbZSQmxmrFCzfzZjwk70xN/F7WNv2Fs
kXdWJOYvJPtPVzYfTZQ9WAEGE64xUeA8Ffht+YnuWs6rytYlKX9EJy+r7aPkyqb/acTc9NAMWgVd
GONHK0XMttHX5ORvhNWuEIr8rtHT/BfBK1J8sbtl4Y0050JLd4JobibfCf9OO2vVd27jQTMNt9oa
6RtKlmTmCZM6t8toT/ZBjJpf03Qfww2tGGbkM+Xu+91NswfWQQF83C1KFj8NEl2F8z6HIcq1Oojf
zZbo9VnPGspE4Ob14op/4nk93xW2r6PZK0g2ZDdVzReEUQ03k/DOIl7tKBii3H4v2MYgVnOh+1JD
Px3pgsDy2uOdGq3bUxSY+VS1RmGyERRSPNF46Jgxgv2opEwBkQPhWchDdkXxieGLxVzVw66Ee7Gt
X/nSZT0keLtQNaYpM6Cr9Aqz5LoyDhuyfxPSmP3hz+JjCu3unP9+/PX2BL2mZ3+gaY/t6Tb74yLl
5gj1w5rKJOx4TlaE/MM9O7sidEtSFi3mEbwmSFPxTiHlCveA6ktkIrul55e50I/5JJhh+ii5V6SZ
hLHA65yLANYz+JtRH9k6pm7JwhtNaEaNK6fMOVq8xiKluqlrJJ68mXTPhwemdFQMKVWfmf0Su3lx
eQihPGXvtmVq+W+lb5x+OUrVfeQGKDYSLLAR95Fve72ar3GiaY0Pb6uTcGKSVT3M3XQ8tCVIcout
Cc91UlmhXg1e3lQ738uPFEYGf+tucBd48ddAQOazn7bPcisvhFT/fC0R2IVrQp0r2083wfo+58K1
EdSkpEhG7gPb1GFtSlwQbr8JIMHpKE53C7VAe+oQCl5f8UqPg1Z21fSkUP1zubqIs2nPDznFE+CY
VaS75AQ5KVWiSM4Cz+BQFtOuzalEh2XqUDnGqGCVt85IEmckaK3YJ2QMUTgiaDRHyRfeaRMEdE4w
UPF5LjMvkBrIzjq7XtCy0n4HaHv/FgKMovF3MkLnxQyU00cmrHr2qeibsdW3BLytOfuR6tORLIRw
qqxeBSOoUQYddg2n6zL6gL7w4G66PCz5LIl2YTRY5PKvqmwueHfP7FjXBIx5lGeL9fMgxaCNkSeM
qSB9REK/7xGgkgQ5v4DCc2V+QEIkPOs4517KJBm3XM9JRC8eWuN7CbV1GnX3EzLCLcpje7wDalnU
WNnsyYWIW4FCfQp7G9Zemn1v3M0ZzE2geW0KRLhewxQ43eMlRWVcBRKk10pRb+kQX1UGKEeZdH18
dIzIhMBPvREafX0c8My6kDAR6nuonQN4TihgqkzJNU0tEIfgM6cGp4NDPEUsqkNzOf/ST3nJKRBx
9fLDBEkaCx6V1K1CDJvN07cxruQSVye/r1EvPPtVilJSJ+AAlwD0SO87JTZN5H7uiJz/Z6rqrr8U
5Zw7CzJZ9DVzHTSO08nc1ONjEdYdI15ScY73R1iD/FNk5i7tHpmeL8tcNgOcUwNwCAGEQuSMszPO
kcHJkL+J+GfFKeGMfgw1O6hVX49qjpkvQje/ieBofPugT4V1rOPvVjIh3jxDwUsWxQiYI2gurUwV
x+Rr/TXSs9FxwwFDTMKvG09GZhEm1GHAzZsdTz20Jrk/Q7fyviqQlbwLPEgKY/C0yhWuSAov6B21
WjS+wK0B+k9yQhJdh2K5E4Y/+0jcbKE5PxqPReufqa+fD0400SbomTCwa+qHNrHFan7yuRDR3Lz5
2JELSrSz0eXHUJmStEHWr4er1chBeWoZnGJ42nlvGZKST0MAr2GBoImGopDGcKa8kwi5DbOfLhzH
ZoXR/Gv6It03RXEOAj2KbNceGan+CcCkEJO+Q8JyBjkIunbxlrJNlFEwPIZ77xgAR2fpVSnl42ip
ZkZ8gWaF9C8OGs4N2zeQ7sgy06UrTrkURmBAjq4Jx/Hk4zbtclr+sHV9GRSl9mcCBC+JIcx/qDgD
qNBzgdVis9bzA5sbgJXRVOH0pFJgkHOArdY9o8NJ6bXTlBSRP+aNRWuNzECb9mMN0lBoZU30nuGS
7aR3p4Nsp4cUg8pa+PqPn4dNhEe8fcPQEEjwRd4kBJhR1pwAt9x0t1FjFooUJSKo9UNot2pDLzqH
Ju5GKFYh05WGptIJDrygo/vULbyBGiJFt6qAJr9fLdRj9TuIwtjl03nptSt2mRjCnAuhurOFAb0s
43TcrQ6c5kqLvcxHZ3c85o+ev1rcdeZSqF11Xr6d1vH0k8MbGELm8wnlq7lI6Dj3czNYAwlglxt0
HlGZ5JNt1VBpy+vtYs0qEBgkpB19joY7h28z3unX6ZVHiPql6Sb2zBnV+mHl+7SN/JJj3szjhOo2
G1QZPnOKwjx0VOsP8Hkz43aUAyMGyh+D1i+RQOvfaTK83rcZQBEBfBYKOuiWFlEWKG/sdU+ipOuy
P/o1T//9xcNGmJMcbJF20hpUTog2O702qv31ajMFC+4deXTo4J8xSN4F4apdOKmim6XPUZREuuEG
utipMW89dQeE1L8sp232qlRfVBsVB/Mp6KmeMGLHYTtvwnNkURwPr7V9fdVxk48L0Oq4e5w+gAV1
EUGm0s+aV1UwtPWBpzDZPONOXJMhRfhaz/yzlnzDBvq+/yh7IJ11tdzH9nAdgSgf7OfjsyN5s2Wy
2aJwvg6ktF3HWjIJHA+yw4ngm8JaE5lFIxRx+piHvbZJ+BkMrcCq0l5xSQe2Gi2cSFRfCU3TRrIq
cQsmnXp2s8vbLjFVPN48MqjD12pmA77NHqxJ324OsSE4JHBMPnKekr/neeYB2xlysDuXD6B2Bqm1
MTvI1n2igZYrtNkYdnaVXDT21DVXOK2chRS5kfF3sJhzcqJ7nhNvnnb7E89zgSgMzZq3NX5w36B7
55n8hxEAUunRWUI1Z+UrnSRDHKTkW5PVIwA0QZ0DBx+/u77qKOGWzbR4qDh39AQXZWTJvHyrEjBA
is1gntoDQYKNbfTHkcJrhMezfKQGQdDaHVE5n9WPm6OCFZwLFtnwDb/8Cvxwk/vo769+yGhxT1q0
yfZBv5NPzCUZqWzpl9j8I+UYCEk2iBB2PpUrEAbLGSmtcmkEiypnOcxpggSPN3EpVoKHI7r8O/xT
CGQ/CfV/K1kFKeVEoEEhzmixxVt1TYxQFz4CiVS8iiYwG8GGyd49gG30Z99VcYIKEpVjBlR0wJu1
Btp29m5wZHNcllXf1kDB+mzCLDbvCNklXFSza3YpERvIAt/NgA1YEfwCeIuf++3+Wj5r05/oruyT
SCVuoVqIj6WgxWY8CMGXeOuFAuE3N7b2Ywit2Ob1GgEa/eSUPe5Jdj/bfIqahTwVIpkbyxsKBwD+
+t25EPtZ9vpX1ZaXfgPC2Ta00MPLR/n0XjPtxFWCTZk+u+9DuB2kGJCcXuk0Wkxbt2dyD0C02y9w
eDOmq5OU126LzFNUTgP6L1UW5HuaHqqHJUTtz9XJS9ptx6AIm9qc0mnGgoD91eWIC9+eIWKx8gHH
i8nFPMEBLW/IDJz0Tvz4ZgwjBWqvGBrDxk+fVDw2CBhH79pb+3CtycVAQIR1IiJXYXklWtZDs/sz
XqGgDQzqIVUrZur4kN/XmaHXm61cCMsKQjQewUuHj5TI0+bD1TmgThW7JvwD8wtq38WyYyiJ9kRP
VzQk9Y4ih97CFQSb43FxeTZkn6RdVr5bc4gvgYft3GWOQ3uZH2EnncAG27JDgrMA+olqHcdNPzBh
PWBGmYwOgk+Pdi96w4D7YJrvH+dMnktKnChCoGVu/1vuSsBtCmJXkto0rAhBZalenhKvNvk/+jEP
DQYSDo3GjHeO2R+BLV4B2KjvIniIaKgnvDIYjJermcb+/pWD2dsmPjpNvHQlBiVdcMLZXWd5Z6dV
OrYBhapFH35KuF27hvoP8YEOJ8+KQhlTAjST/b7tS4k/OT6FBgBQAGei69FeeqKM9uqmj54VEp2m
s3W29n9rMsXaVjY2tzzxmC0ogiQEta/DNBk3Q7H+y3wY/AGIc7WT5Mo0JA2fRiV+ahhy9LbLr3e1
Rj4i8UFlRwQmH/uYMiOVFtsaZ7NzLtLL2QleIH4ICMtK+vyGR9XXSxQMXAz7zNrsoYJEKsbQTjoJ
jc/iNV8n4s6HwacbMocmvNLtu3mAYGBpSPh+ijrj+QUjvSgpfLUeMJSmeMEoqpYbSY5hv/2u1Srt
Hgc65szuWwHCa8YAx94/B/Spzg7tRYoe8KX77cSDOmU1Ploy1nDWGAhwmdA226A5hbOpoG5iEALl
B1jLiZL2x2+jPdHjFxs+dnpLi92O+C62XtjARx9XvxK61STeTclwUUcRd1NbX5f9RwRO4HQDXShm
TPSnrikD7MUVNkbBHEZxtvgVGIuVR3j+ah/0NLLh7crP5OuUzb34UWcsfBVMaq9PTB1BZcAELxA5
2P8nM72+6RroD8vKp6hUYZbQxpIASQm6yAyEEFRS478xLD3ID4gXCPvx204Eo0HSpSKIvAZR6v9i
zGAoGx4Jjsui4PvsWMqm1Ui5YggqsloT/5UN3UFeSygWZfkoInL86I4TQ0NSwqi9WKKzqftCeofn
timqr8C8kV8MUR8dcrwlCv5zTS+pgqTYEQhjChoQdGYVWstYdW4r5AfAQ/WNVxQj/PUM2w5oDeMZ
+70l+Lo9TNw1ajCY+EMQu40LM0in1qp4x7wdutTBpsEsLg2OOefEmCu3P5391+Zk6xJ/rHP6zY3x
9ONWT46XQowlT5rQc3VtH5CL+PTWfS56yoMtr48JY9SvmPnTg4HP2cgor6EXQ3wfONItglNPQeX7
Uu5bZBEK+yw+X3gK/VXGAWpFc7WpQqS/M0sQNA2W7NiOkuygH7H5dT7wryzQPhf6nrvJVfDpco1Q
mWhmFELFHWDVFEGeaFFceC2kzgUFE4hu0rE2hIOMT2WOu0fKfiNo/m2KiiO+hhIhNeJCAwUp+Puq
sXY04+Q48Ed7Aw105GcEtafJ86UuORn5NYyPsWyqUPTsrbz44qeh/4hpauRbs4v7uPcRC/DCpblw
FNpDC+cuDvN7rgzT7XtlMpO609KuYVTkNiG4qa4220NoI28X5183xexFR398bOmZQzrZ0SNBv0+4
g0+ZApQHAXTDLwy+F5wbh5tt1pDvmaPG279r2SHvHLzQ8Tif9vkddCN7aUvq+Alb+gVIxtqdSUFG
ZWuDf5oVG67wG1H6xGnejGiE7/HSCPkuSumcfbpPyiht2NUqFQxyWB/QiVT3ATldNg1RaJSClHNd
hh2QUttm2/eNLfmgnXkNQRH6aQA3YrcTgcHSPWekXLGpoOAVtkCFdIFZlvSECyG8eP3Ph8lt91Bv
Ks14mV9Tx8vdncDQRVeyrKZ+tfL0Ng1glUcFjS8LuoqPdMU8GA7xwaDJpDwk8mrzOqb39C4DxJ7a
vLV/YnOSWwrYA2q8s3MiMWJaeVabYaMlNqpv/H5e1iWfc+cSfTaW7j7JOLOGWyip6PmT/h8ywcU3
wJLIzqcB5iGkJZyoWU+3UyMTOraKadTtiWtkb4Jgy45AoaNjxMEB1k8/1OHNliOHaAKVojMgk+YS
balOe0MimjCgUBn1Ku1MPLgzOvrwMG4H9HbeMjgXfkMBJlITrieyW+WtvEyXF2LHwH899DeTaUmE
LPUoyVy+UJt7vYT4kc5pW5DIgb/xDyxuUbJUgLxFJ3aP0OAKslquoJyDYUCt8QNQJe3REn465xsd
DhYG48noFDpiis66ayqrO53f/0FAYFX2QHI+JfBj/wyUWDyuQrXvkUf4n0XxGfJZfmgjT9v5+eXg
76YJyzaNX5ZcsoFesgY64JURJRo0HsaLB6ARPv6w3YEt5M/DH0KhaKNKofQJ7yxmT+z3M95NZkeV
/WdFQlUxBjNEqEIPELArbPmFCN0CwknlE3cDfIdwDvcH7F4SzZ+0CTJyck+oL7u8AiYuN023nW8N
jfJ6xjIKicneLFTjWbKGv4fWTCPjPhJPdAzUw4FzDZXhnjjIVf67f0A3p4xJbcGEqR1MaNT16Sew
key5QajHJ8KcfXuidtSRhjQkdOvtjIiVc4mrZKW3aHD8MKvSA7wTYU92NzAHw8ZV7rRZrIQWWg9A
3a4QzcAmIiRLKp/evpD2d/T0OGO2uwq3Z5K+pgQ5+iJ4T/wz5NHTAMP8SghrA/i3OLw6EVs4Bq6k
4we4F7BiL1VKIsCN2ALC2ohcBQpTLRQ/61scdcQgkatsLoAN4M6qdbzew9PoC6I0UiNJ9h3RIXqA
2yUg8pBab+h96Odx7AFjXH7oXqd6NAt84EQEdkan/nLzoGNl3OufC/SPmysQYgYvkZ96RSmiJgK7
ZG5ixUoFtTJpQjgQK0ULxZQV/N4pHHGdVdeyxXVnQSSv35YikjWZlbj+li7MC1pbPICJZ00QzeKb
8aVm3sXDTVWcRYh3MjpEam4cJgWcFZXdU8+KymVs3OK2HPvDKUHIncyQuyWt3S3G037vBlR4oWzK
fGpSDJdZzhIj1VcXcKcdXQgwSMUxjuS39WodJqSv3qFU+VATiRoPKnLVk5gFbqPlV/EnuN0m/mI9
EA8Evxykh7k9p+ylBqVITCWUagG/2NQU5E6ilwGMIs4V97eFs5ZpMA1GAFGK+99MX1Tr9q9RdjSc
dZFZHZLitkr8gOjbUiskuBgtkrfS1vW0ZuUJ48y/xONsnDm3UvnRkuA7cVRS5mRfL2jmaYF01m+Y
3nH5puFil/kdH10a5Ivd7yuiOTU5U/jdpF0VPzsCJjy1qEPaFtK6S0QZw1k5RhKXFLFbCnJDtu6W
G5Pzxmvu8QsjIS1uexraGH4ZgTa33SksEPIlFspz7R8DvQqiaY5lBA7ImDlEbp2n0G1ANymJbzi+
NErlsmgnBasz332+JLkQSBRdxwBLEFzrlXAzeWhi6fRHZ/5oC/dJOzNonLRFlQqjcYEEKdO54yCu
oLB8oYO0Axalw6N5iB8z8ilfVkT+pf6TMo35iPannOgpVolVrevo6jEkFQALPEu3UBHKJSzbdZRB
oojzG8gMXvI2H/WTj9P7D0R5GOLUdCbRF6alRTonNMcigPHTAoOXzlIBtqWgWAn+zmZje0zq+POr
2TClZa9jDMC9AzrsTR4jX7yhFBGi0cKE34Yalsyjc1vY2Wf1GG/4M9CXN/PMQBGLdnlYf6QKwtk9
vFdzQzALRxRFWmgqJhcVzF3ldxhb4ZeWJpp/6dDGk0DGmLZaWTfwWp9Vux1heeSlf3BwtNe76Cfg
RICSIsiSr9U59kEOWBy53LBFeqqc+wOcxICNGOCUA3WstHs8ll3m3AZvlCDT2oc4rBi6y5s3mdwF
gERMcdH7bX7FQSx5xu5g+JTlv4+1U+ONlGQH4Mx4BPIVWMXa+MXHpOgUtBJ/38b+znB5+2JzyZSS
MEyMdLh3+U3G4WU+BSeYiSj9kcWYQPNDlF+vx8Lz+/InT5AFjlRelnsNPdywxOKkSn1fufN5wCFY
JwfVy3qBoDWNhhf6RuPg20+D5RUEsg75lx4LYki3dZXte3S1lj1RN4hmZPiklxoUblNrcIS8bvC3
5wbfuGkIj6Cn1qXrk09OhOVPMMnw+EnD8vIMAxe2W2/1tQa4X31x35qeYStNXVQLlMxNxaij0atj
fvg0KkW9xBfybrsBNkaaoBvXkyrkNOWv1o0YzMR26HsCMwdXP0PaMhI25jKDf5jyj3pvdVmYj7Rn
cY8bj1dEEk9X1PDcP3omL3H7Hc5b2zV99g76K6safEprlGpAuA/Lf/TLiuicXkHyRzPHW2Rpu6sl
TvNQJ0PahIXhQrwGtBhE6JEAJ0tlbkDe9aQBq+J7vz/8PZYL7Cl7QvvipcgbgE69/Kje959CfXgU
Iz64bzZpnpEkOdTiI4jWfa/OruTAeEaCdpXb+xth+PR/OlGDwyKAsuA4fThsb0B4beRV+G6ckI93
xATiXzcwy/5Viz2dNrZUMk/62uOKYAQJzMnfmJgAhV+2fG1msD+VaQ8Qo6KLXK1L8qDH8hPeZ8/u
HAvfikHloSNS6RaqAyXdZKI9ZygUIhbRvaRw/VhoPyEsvf3YA577cq26nW8herLTwALLGrnEx5t4
kMR748wOW41fG5wU+Nd5YO2//oPANjrldAjXCKmQ5XurFDea424wsEkZBiW8zAXdhGuYsSVd75AA
llEH2dW/jZ5vNOhZI5bgPh/qQnIk7VLrKB7MxMlHvd9Xv/xc1ncH1ElMeZTy09VwJugtvitnmuQk
k/wiC6J5a+OEHezqjZIhTM0V3eGmIlTL/A77Wph9OUEISj1cOEpJzoSuPvM/BoUu2MN+bmGeBc2/
raL0CXSyiGge+ujX8l4xsuId3Bj0/cTgPxBFkMaArecb7rLQKlIz7AjV40KvM/cluLm1zA3H3kfQ
tduXyvWG8oP5gY1h4DEDLWKoYLmUeQyX6v9MI77t9cXSOgVf2IPAYrqkmxX9R/L1C56vbNmLlvQQ
r0z5jK8EHwcHoaAkRLAZoRX54bFMP0bxvkvVBwOzb20GCxbfeEsBfOZAArBk8c5UKAETi0JfhnEg
F4SNn07mgmbPRpYdwzX6OIUi6NKuYYYJmCZAKTW2MUdkuDUp1pmdnAio6p+gGeUO6VWiC/14u4os
Vgz2VdVqh5k/lruro92DnhVaYpuduCWEW5hg0E70mUTn/NJsf/cBp1Sz/sfsLIQf4RoXObtCPGnN
6F4MGNLQ5jHII4FnCp+P+v3ByTQDJYL8gtmkeJE+9ayyHOljITS1kp2WGeXHx63433/mtbIf/5St
9QmZ7651wihpKhAmG0rCTGSuq8nbiwrXp4E3/kF/ai+y42fEpARfYmGn9KAyZReA3bY3z2wiIOMC
vyMmTdoAYejMzRg+xAUhqL3fiDXc6wJJcO5FG3YfHx/SH4OyD4m9LFg1xnchGc1oceHm6rY9fhTc
uh5Op3d7xPERXr1wWN6XeUUe1fr1MweEkvlwTME/nFimP2ND/YnUg1DrLfVRX9Jl5OzPpJHRjDlp
EhnTv0Mp8RsLbd+jQ8yRTKHXMqgC+fO0TTkH30B4YballWF+Jmr5Yr1aUtzlBEEsYalkBe7BSbL0
H6ACyUQCnNBiMBIt0K4VmO1VXiqwVCeeDz2Vu/M8l70+cE6V9ygnoUZS7rBD8BHAp+0o1aDWM1It
fvuun30azinGkg7+UDq9OZdXHFbl3uMW/OeRocbANtn6bDQ1D96w04HdhUJO4zQ2ujvSpoAJV2v7
2evHYM/tcstq3MttNyVzoiE96ZXKqfJStRm/9VWiLeeQLkH/j+2gLJ04/8rzojWgywBHCk812pr0
A6mSv4ULYsAmkNjfRdhl3ai/dJWlB1EKGqro3NTxzWEv9d2VamW1AaS+6NxSjjM5zvJwCcpnL5jU
5ELcWlhTtmjf23roQAHZ2yrPr768M+NNQWaP/Pd55n28N0/3y+E+qfFjVSw8j6KCaUnSLTLyPPGB
Nx5zCru/6rz4mcij0YP0EVE7G8s9PA5axDWoJFphZL56ikCib/x3w+DHWpW0iFPxohJa7xpy1VO8
crqgFw4NwfS40c/NuqMn5nwRDTI5uhSGYyLRLYpkU7Ge2UycQ8fVGRCwXgaJb109Sg0pURUZU2mo
6rDCQZ4bmQl7CHzff2X1/RO1pFtcqSd9BjmY4U4qvPXirjQueIfxHhUJ0wyZa8/ytfwy91xfCBDL
YRhw8f7BVQX1+RO1AOAhWtEbojanPenWpuLzo6MVIOFtDB7SE54/YlfQ+nAd0wn4a6Yc03ZNyq5A
gZ1fnTyS00ZDstKNUpzKi6Rm2LoYTDUgcafDi+jXKz+vCCnMchVQDYyGHtBr8xz3sbweYkAJPZPW
3i3eOgP4RkBCrLWARiEHqPaGz6UNnYGC1UG0ibzmhx+eUKZ+/RZr5kHcHlblPub4/x0ITD/lvrc3
7LLjDqf/OiEJM28fXR0j8102nAod+8CPh5BZZ+OVeYPp7m8RtXjZaAvXbCN8jSFbHekuYqfJss3b
yBUVgIeB3uSMKx+jJvHRfA/yqWmsYPyAowhrcy05Te2+TBWYQD5FHlbYQpatejZyxkBYVCMhZ2tR
Ggij00Kr1leaU1Zz25jKuMAz2IeCaCYnqN15AiTWUEj0VNhcthmr5gHkiNciop8L6+RGGB3F2m+D
/42XH4pUMGutBgk1rVCybGa5fJXyMaMK7wIph3mrjDSqroRmGJyCQZxXpwptdQKD/iD8Bh0bOnTA
V75+gK75zGcAEAdLnMw+D0MFsC1Yy52RAmN/FkWagx/OgNfQcLZbRfWnoRX2Obt5t7WWZ5Es+OH6
xkh7gdCu9vTYRk8earl6dIAQvjL2T7318ojVI6sqaztL59HtlU0kV1sSRdoFJ/9yUBdC4mRmX853
iIoup8GWOz2um2kVClY5GNUTluysUcq9etDtax8sI5YfRcqBQ6FbeqqpPAXv8L/KGI2gfzP5lqL1
wT4/+2Cz65nhHZ11fMcssk7KDVpcoCy3LQ+QRXNldFzxu8aiYK6ZimPFSnurcBGZkaOkI8RiSm7I
RijDoh1U4pJ9UF044oav8AIKLgFrltT4QUAYoY0naJagmJLdbmq1vGi3nb34NlV74aHk/aIvwFZk
DF6GEiStT+dTPzaepr0EUkRWEo7+BxyLWIl1r4fsivCC/fCe2mueBu8r4Wx8tLIDAkLeG1Re5wbg
AiFI8TnNO7Ym7rKZ6T22VLTx3SBqapXcqk4cmN2aOZlWsptoiu6ZNxavcew16PuMlLVenb1w3/qH
xQy7GNp2VI1x6VF5zpLpnKtJt+8LZ7fCv8EFXPBM8qzrpYXs4F3UkjeZb2tYAnIIyOqLkOAw5PbU
sirYpXx1Kix0cCFytmWLkUOw2GrR5LP1tlomHw8wgdyXCelJxp1VKyHfGUGTxZDKE9Xa4UAqxJT4
dmV4bGmQ+S4XWVvrchCavF7gXXPsA3mjG8f2XCKe9xJv4a+Drgdilfwh3IvyTZeLk+O1LUbg12fj
S4+hqMTyjaiywmZOwo8KH4R2ULLcq0VoVgync1nppmgxLfW0wnuCqwSu/nO1nGplmcdyV19jz3Ml
aKCM11wyjcI3B0rh3cL3m04HK1np0iDaEBtVD5ys9Scz4TwH4F3vdjZAx6q5BfRvXxlneAgs4nL1
nOFTJsmLVzrjlCFKJ7/0zA9ub4Z0izm9wPdJJFwOMCCNOpU/UoTEtaHoAOiMZUUVLG6iizd6bapj
wuzR4MH51dL74RlPXhtXbXrcibVYQFMVpFd+UEoIEgs7UVc/kAmvNuxNp6PFoquXOkKGfI70HvzI
eX4e3pfZlh29sxQgoZEi0I4fJvpoWP1y2L2eO0EtPLkjJTNUU7ixlw7X7Yi8pZG69+jFqRe+EiOO
CDOScCDecQnPuxCeGFpWJzvVPr4SEi+BTsLFq4UzlN78X6gl6ITZHLUrOq40kKm1awpOfgSr4inn
XjiloehLrXpwy6lCF3m7kgcPY7VWLotPAZ8Clk3457jqxx0fGQSSL5h/YFtaHdkQAxpxUBop2FOd
4mu7ugRkVx9yexxfJI4h4LPvNAuYCytUeLVG9K/P0BCDOXJm1k5WsjU1WC8zbQhZD8UR7mnKbJuo
2g/M4RSa32fFZHcXjNNDQbwpySRQTHa3lXgfiBpb/bF1ZBNtDe0lgC5S3UhysUbOZQCkx9WF9h9K
vpSbVc3UV4sr/Uo22uMQNH3ElvPrq/pxypli6ogmYzhiXpNcbzC6h4kZKsCcUyBn3kGSooRiAmQP
ZIUhFpXWZmka0KcirpaJKhq5Da9fiPWo5JkixfmJKYtSmJajsIUB9ziXRZZdA9dG2SCBoXMe40iJ
Gv/plXOjAeZ92pWmizclH3WpJPgOSQ2x+EQufNGvITkxX9IJ8YgVRub74D/bB3ZvZTnyN8J0gMXz
JNz1Iww+mRQNr/9WEwel7ao+QYR3lRqQOY5t1/GRPXtsu86mequGsPQWPfqWZldOJau3/8kWMXqC
MzNTGFC6Qeti0Q6MmXzNSV48o2DNQEoSLXQgeeUSzKgk/dr0xZ/AePQm9MZFCV0jZKQ2kwvWCJe1
LOiWTVFxzPz7W9sYiUyjAVIKFca+yAX0DWjRyiLwTF2MLvk6DHYQgRs+iTyzWgz5+/R2fjyW74tL
Jzmln09dFC0BdIQxexa+kXyYhWtVuo5pE/84rZsAJxxUSJHOY0e5TOpS8/InJUP0ndlFXfJu3D5k
A3r/BQa+xo4F4d4fcVVWvEsDoOza68bPdSC/b1nPa8hBiIlBZ6DC5pSnp+14/9fqEiyCY/ybvZd7
vol3ZKaDIXvNflRXiSiY+K1fUBMwpM+ulIOA21WW7ZUbaOp7zgqAzuk01b8+mJfmFppA0SxLfEr3
4HDF8/T4G009zjXAblT2Hdd3SnB9l6FSJzOtEWT+izpi62s4LqILZZb76T1Js+E1Wo/NDNEBQYxT
BtvtQDbQ+q0ioe2dys7zz97YSWd76KOUaqcMffJCdnkg/aek1U34Vwp+EBvGpMyGjUo49A8ewAdu
nhVC1qtS3KMvYCvluaC2RcLgRnAsezpIGvL6XP59RbVw/SEJw9Tgwlwe/Kx/+MakILCZZiw6qH/W
QinLKPaIyjuIizV7p2NzC1cEIpDXTxqOiXekbFdf0/FFpNw/kiKFygjZHW2KMKFzlgC+kEBOUT+Y
i8y2SOfXlHYmcrBQJqwlE2HXHK5zGXKmLtMR/vTsgFS2bEyofCG7X/Xyd5F4M/7/2pH6KMe1WCSs
aRT7A1KPUrSUs5VQ4AjtJ9+wbZC+EJXI4ItfI9J8cmrvA7nTYO4HvWuhm5+fTm+jLP91gSvmzJrK
ba6BviGhTin/0giCDvU6mMzs51RZ6UPo7+F023WjNmiSfGZdHVDSlugU+nLklj7c2Jd8mVj2XeqM
gRoB0H2XHoxOBtahh6y2/jYwARS+9CPqM0iLcY+uh1Tb2MZxC0jxZXph7Xl6fMKufnkhHdqIGqOO
z8mfkWtdGWDQFtZdxLVJTDnZkgq1dQmC2o4r7iL0UMgCB06/gQ5LBqWmny0u2nx+aJwByxZUIUs5
aINcjnjlnSKxULujJusxa6esS8yYHOpozCk75e1BYnmW4pF0k2hmfkEoa2VEI+7VqKiPTigRaNoZ
ytZ0RSLXxOWl4BAGOUapDixoeJDHCWnIuy1j2hzoxZNeZrPYwCCKoO+/Sw3Mv3ZCrhl8ysHvLp4N
sZAxWRDIaNvNbqkhCRbKsjmfdZLITHOjWYUnUBHYxL8+dOx2NfpTuNVGxOR+Km0A8deihkxVc48E
70uuQ+hSC/Sum+p/MwcmiZE45Iqh5U0qhlCH+/L4xlZbABMgqcRk2BvMJFeil5p/eJeKfozBdQdZ
ycAdZWvFdPOiBn917bOQTwwMHtKS6DgJDjITwnM2hkmc1qncLGUAuD6JlzJBKv+/PHyiph0P1fPK
MgQYxbSiSGsv0KpMFMruILaDlPGQJaT3xFZk7PsJz/X/hV72ePU2ge6JUtC2aXlgWkeCRzMjonxf
fqNJGWBYHh/WUWHbGi9Ie8qZVxloPrjBFfhbtCNfZOWLu1pBXdQWuszl0R7N2gl9cPUPPc1UK4xO
1orXGxJeTRqJKjZMWUw02WlNMLTMTnirTw6D1YQzGiSaQny4CzSaAkA4ITA02AjULFfXQwPQnUx0
SyF3wqdlfvglCF759l4ahwZ7DV0vdDWp/WltJfrEA4aJhS1LDeNVKdjhtRm+DXkrqnY+vE0SGuGs
w+z2ut4KY6Gq+DmJrwUkXVgslK+n8/4IRuoCtp3xlG88ony3mLoSqEl/0jcy/J7pAH2bClGpWUFE
DJTfN6o+RZK+Tu8RRRqa2/l2Zb67FctEGY+sdRED4g7FkbibpLBe6szC0ADqCfRd49uDhkZdDd91
1teDetd9FvGsj7du21bSEGEleaSiSMDZlMpRgz9snuAzQq/LEuv5uN4/XhdQQKAzNuod9Kg3wD7S
I/ORsdNmw92ELZLGBRJcFF4PIQ/MR1sgMbnCMJE12ejw9EDZYYKuUgqMrLbJOg2JvIvdoFmXn5WK
qlHwbKjaOqOoBmI3nKNVzp78nLNIyApwv59YZz7gzvcwYlVTNx2ZzXViyRaBvySLOldFg4NOCZEt
z+pD457Yamaij/3WIIKa4GxkjRx5pR+yG19YlyPMxNQhLlnQ6hnvmIt+E9J2bGy2Rq7ZR7uFeX97
5pk9fPT8RBUWofKwNpgYqW6RGWXn6N/OIBwAgMHRBhZxppj1k7GeBKfbMBmncaiDZrH9iwDW+v3V
fOMuNHYxAXE2M6P7UDpjG2xjgs3waD3Q+rSpQTjawOK8MAKc80RyWE0F6xjfbrtsBE+dqsylyfgO
wJ5AFKdphE8nHxCyh3ge14rXPVUC4VuFqj1H/C4SU1/qhBUCiRnaNL/wBCXxBcbI5XLfhBMrckWw
WCjPoPCvj3t8wsBwpCD6G3kro2pBCl8QchtzyB+4KC1j3nCBVSuVrxjsI5Xks8fYmcLJzcC1+Lv9
+aLTk9zIOCq7mLYndRazzq4gtCU8vpDzu+guUQ2Vtr3yEANiUTBG1rpoIbUqyMuhM3BYNBfJWk0+
N+sPCiNPZnLzPPpCGpmaHZ+hB8WH2hRt8c4/f7N8jvfWgC4+cu5V4TPxQpx6WuY2kVImFOVXMuUb
69tx4NXdTyHavXaAGSVB8QCoaIAJSaaCaTUiojoFWRSWLvtO2jMbIZuzoboP56rSAqP0lXh80h66
InCuYX4EkFyllN85fkQgb1VT+GqKgdbjgBZQnM+hrmrjNV1Hqp7YlpksEgHnUNL3/QZTIRW99SlG
xNLvs4VoUyrYzS5z6nMiAUYsehPkh3E4ty28pZ4rhVT+vnt3wkSBk4itFfNGyFy2qp9G/T34r+/h
7QV3NAAoVaEIwJWesWt6hzt/GuMOnXaJ1nlnHKvLpzKthGOd1u+g+r589t+dh+7jypUv85O2o2G4
nF2aCdjPyQBWHf1oV2FHUccIEh5QNTrzHTrZIWBqIPn5GMY2frSQa0fOxcRJvjD73rOriNB955nw
jfpfAz9lIAWECD7aytsAaO16u+GIwhffU4FRwjn7yoN7bZuXl2vj+S1ghWNdTpuT2WfnaeVqlEqz
8WjNVmchOmNXt/Tg3hXbVJ1YtcX8CM8JeNx7bpp1pZ9QqvoETIYPd2JJHnRdvuhkD1/xk+LSqCnc
mtFFDtONkGF8ybOVlxftoA+NK4OhUfHFbHnnYZVgIKuOVkTCPc49/7hKrRCDQYW6keCCd7GqyoTs
a1IMw6GBm8xiuerBPWfa6FdwRAUhFucaZfF+UUq1c9CkdgKTHRUr1iylenRp7TN0F/fJqDLU/fjE
Z9wOuD3oXTOXywvfMhs7kyeNH0/sdwPpwtGNVJtJ0ftYUuqdC2yUQnNUAyyybdspvhHDGvBkt1Ud
Cd8qltT4stCvomYlr3bqTLdLsdgqmh78pSzpqua5Vk5CW4OHbS795RkCdffSQWf8h6A02VgWpYhu
OJvtGlb10Rd3wttbDQNJKufHNOYxy+8f3fyWkdhjh2tqatSHmIpLiqb0GFxDmdBY+RURJDxGTT+e
C//DeVQA7qJSBzTxh9CcdvWmAMGG332CAiX9O2X9WaaBBJaFiQEHeWNyLzKvzn5smz7fNCe1jZug
F+RPnpu9bWz+0WLUYpT892+WPLo++UiC4+OcuQYfZaacvOGO/4gfC84OTfejnBlYk/NjeFVuVLvL
XnFAYuP7As4QjcT0KkBwB9P+Msc4DfxG7SLt2fXPbvcHFho+scFPMW4nph1WorZqn7A5mzLg678n
ASVshLcVExhh7gKszn59YEbkNne4AZdf3xzsFayhveWNikukfB/ghErQwfJCGzHv8hKoeeA9Sb2+
/fXngCUAZwWkT0W6lw6Z8XXgGLct+xQulzjmhYr9VhyIv6DTEuYCCIxhnVnXMDBjGJioyI3FNVdd
q8C1LKLhhFALL+G/LlE2aEs7JOVYVCppsAIoZ1V8RWl21wf7dFK+di+JvZ8mxnV1AePLs6aB6FOy
XxufMbUgaK8Tlr6mlP8DHoVF2baGGuR3Z87USbzng7WmgFOvzhwmhiNKuiupo9VsCMYaJ5WoOY7a
LFc3zgMlcIbR4T4oFxe6jf5NtORlgjW6p87rxLQ6yGz3J1Qe7HGQqatjklDv4lrpkcTQ2dENzaqy
1SsVcOqw3VAuTXXhf/J+2L75rf9YwBH1x1Oehp4Qm9eovhXGyLqgYDcJ6FcW5EruFAaHBb6kiuWc
hTscOPLupryR2NIfk1fliywOL4XWz4lWrln6GxE7Cqopmpgb6gXVAp29WuO4/0Fq6GC4XWYtzDT3
F14cJW3TkmWQv8OCI6qIWgZujWH97fRUV69L7YI1k6D85WYkmwljQYLH8bdPR8uGEAsImea5Ezzh
z2LtTLVBFD+/XueBhk9ispOmzFSqFBWUHdzVALA626sFthY6I1+IaaNuhSEdqRKdjLu5J6ibmuWr
5rBcA0mmlKJ+2DPY/BEUzgDwF0MCgbJ2uLGDn10R8uvghAr4+7hpWmGKpWrXcTloboiap7++HPaj
iy18jfDIlXL/XQKJaEkp10r4qLzX5TTDoe3rp07dIQ8VHUPPzoDPpSuykdPfZsBxkZUyIAWdpXHx
i6W2wGsVUQwW5xdJO+EvVkf1b/lLLETij0jbsVH9EZb5l6Wn1LsvTHpnYIc/oyxH74M2X3DPV/XT
c03cfTmaOKWx8gJUQx5r63jR7GpjpVlrU9NeeePz+Q+ppI0O+rDTyKnxv07V9RrqZyHhAdcFKuZI
A2bbW5y71TepKx1ayI6grg+gfn5WDuzS6InfZAKwRNbTg/i4B4DaBZgja3Kyvt3ClLTkMbrY810/
Zol7v4peuYJzOyRCs0iUhd0E7PhS3btGfC1+VVY6BBwOX4S2VBKhEuRuIgPJLYSRB0n8wiDTvrNX
nFnJzk2riH2hBxCYkTdCUOxDr61DTYRAIypB4gGgT4f0i6PtJbqJAEyhlSFBrGZKYOlNgWJLARyW
cLyTOpEl+HD2f75oLA52ivBo41IMQhViNKhBJiSATapVpy/+T9tkWJ5sCGr4OA6urQXnO4XX39Xo
xEaSPR/FVIy9VIqKZkWhLSLdYt6ng/f5PWjDiJQvaP4BE6rD1joW/SJqlu/DjLsOmgfeg5v9j9Md
X2qJFebqt4h5TAd43aBj50V8zQ0hjVfO0tArVVVyKrPj6VQH0EgAxBYi5C/9t3PTrIaRnB6oxPUr
QOrTVog6QdoX7qrmwpczrF60ksnjOOWfFTTjURi94uz+ixlXDPFqr70T8humOjsJsT0uXFbbX8sF
vPyYyjH8qb5Gf999+362Bmmqeb1YSOrUefk3sL8hzWflQ1VyjbYM3z7VZMlK7b/qBN4pUa60JEVu
o6TnoXzFhYmnMSR2OKipg67MvI/Mww/MRf3JnEPN4dXyjDwp0FkmyXDZtL7dDaIeV5fzGPsD5feX
SfA/56MK31LML4Z6XvUMg4Aqt+siVUkSFsGo/TmqKV9TaWRGdu+Dx35NwvVkT7YZ6KiO8gMhfyZv
A2ydY+IMGpN5/ZCH89VeUSm35sLrJRNLlzOXPXs2+iqc0TBMtsN6iTMUbnqBEFG9d/AkelMwzSMR
dQwV0VuiaFnBbvdO+Xmy1I+ahDlQpJ3J/HukWFMH0zgWVvHr3G3kiQRIpvB9A4AQ/mGY/sxE8IKa
tZQqbmCx4Hg26Khj6e8JCOsAjT9Cok+RvGIixX9lDWBzPf2MsXzyoBls2JLv5CtGl/DcSVBHw4Gk
bA/jTzn5bJUw7xgTR0MIXnThRe6QnGA9Kj5dl0OqzO/Z+ZgW/H4yPAbbxSOXtg/XjhQ9HhLYUEpf
3sTmwcQrPVBFXja11WfJcaVNKG62qjqiSCQhPDLV2xQA2AwV2hYmh+sR74pn0KSKRuWCw1J9Me11
AfyEsr8j1YWQwb4rnUZafzI39zJ9G9j+nefro2yMbEZAKv0c8sXZULh+72xb5KPoBFR0Jfw/lIUD
t66CvXcD02B7NmglBdmF9SSKkKEkbmxzOqemmslq7ACKJYYoGmb1P/YLLNN8Ur/ex0ODatRYwVDW
gjC9h+vHmk824rvRpJz+bUsK5CpbtiI0vPjDeieJnwe2IEagCe3ZQhDFNj17XHkSaEXy9YbHEtPt
BJpfvLyUaAWFdhBK73/S8Go1O9EOUbVgmCMW3vVbkzW8eWsHs0l3Y4DvF4QlKfU1+pEmEG7sXyDd
2TOZLUs5HQSDJVkuipXRtry582+cT5HVmVLEv+KDAX2cNjH0axuGG/tJbuO2gY7b2afBcPzZEOpi
3YfQpPPjenDWp0Gcax01AV1OS0N9Rfk1Jiq5QeM7utdGUjjOcWgPSbv6Cn+oUbXPUIRsEUj6Jf+a
ctuAMXRSXU2hvpgMuD/EE0OMF0swRGthJFeYp5uJPnLJZukhwhGRpvgk7cQA2pX7+15BfB6wpwUH
H7ZOmhYcgRgX+YrN2SjOMaRMDdPZO0M4LTg3ecW9tTY0iIIpasL1IlOPdunsMNzjA3MJxm846fVW
eBQXASGQX7JbWKfrilATDp0mguMSSWuzOLEGX4JVmq3vxTqmmwOwuoFpwGkBkT+xPBICtruy87p1
HB9zKN/CWLELm+jYSTTwDFejjhPLjeMr17lI2V/fCXBJwItdI6BxFr2YVu9XUJlgqBDosek92SJu
ckS3fwHwMQk1DQVC1r7kI+Uv0CrjrDs2OCi/tJaU+7ZseaUZuEuacIyIivfrkbPEzd4HIAUjzEB/
q9V/X/KlAaTb716XiPMW+owmrPxkRk9h3w1zfjJtDW4SJq2/THiDkp6K0fHePxqIrBHTnsz9yVr8
7bs+ycteLA4IGrhq+BNZ8wXCP/orEnjpf8Vf3QDhNoLaNgfjfUtW1FVI8hJrz22h71faqylfLkhl
S4M8aV/ynx5ExBBwrEtmn5GkaVRViRsdefPFSDXfNVOY4PyascbJLuT2DqcVFbSYzWh6kgf6PqXf
nNvFtQAy49v8GwvnwQNdTUIXhHL35DFb5Bb4U3ccMOyDQGpgrYzfceQwunig57Hvl5f9yp2ee0SA
BhEwqWf9gDHCHn8X7kWMpg/laCmG0sdh7gAk5KtD4Ok+phflLqixe5EUgY5aH0dBqCB7hS6sv1DV
aLU5iRaeeFOg8wgQYNVmnOCjyMkoOgDQeGZ40lRyFIvySLURW1WSfQ3z5HkGNx1AItcoC0FRAIgi
X7IFgWeJ4JdB8YvpePYJdi9J7uLlbO2ZCHQVgF/KoZ0182TgdxECBQjnDa5M7bNhKVPr3e7Zw5U5
YWSJAKuAyRa/P2eSmX0U7rsXqyS5YqRXIl6dtbJyGm5SvNRovPyJbMTPxcEtyx7O6AoHQVxnsC02
H31Pr2zSW1IWMQKW/WzPhW1/g1T3yw1IRnCjpIJK4n5vprviFLRo1aBqhJzRrGSb+4ywR5DBD4Ga
iRlzx9r9631RGEhqS+lWaH6QN0ARpt6qha94H2nyqqfvrCr0lJoICplhSZprvAED7ILlFk8bvcgB
hJcw0y6NHoqJtpO3IWYGWJvZkZN10L9oLci7FNaA7YZCqL9wcdF18DVvp+D0jbz8I1lpO4uAhMOx
iN9LlrjAM6Sy/M+cKG2QctIZ389MNAWLpAqOVHXSLBtJc0wAtydh/apnZ59UD8sxlxc5VvD08uE6
EfWyEwbTPWMrydd4jM1VocQiTNqoKRnB6NIaN3FeVkW9rTqhcOv8YTYKIDuX203uTbHR+0E3+a7u
SG2O26AlKjfHPA3mCXIOcvnJ3AymTyY4uK07OMrKxFQJmyvIEuNfxTlfFRmiyY3acfmHpWnh/0Nb
EA0/sUKzaElvKgteO2hMxTuNnCqPS1wNQI3zXoGShhAYgzIyjlxy1qw+pJto9cIyYffoJoYg9E7L
j7NbksFYHckg9pBDGzDW3OjTA5rMwvEfQEpMqe8bNnOLuaTyOagdwF8S2+u0wnTgGGfvrf5p8owD
fcYcXuRzkhdKI1i8Ohos3fakYwbwdca8vthoiNO9t3FoVCHNlS3KGNaVingO2MaEJ2z4gJCH6MzM
6sV0bx88quqCPopyrwbhgj0qNnGnBDq2iZnDLZYhCncWu3qQVmjUwBOzEMYC8CsW+jcl8zZrs7du
M/cqw34zmQFRsPEqnTO3uT7/axDrpQnNpVbuV/NbxQuypPnIQbr7BvsBDBj5xFrC2LecpxQ/a9ka
zeLITgWgrmlrvFb77qI87l/77MhbAl4G2wbng98K+IWB2cK7mzBrR9QNM7pMNlUCjIZ1sysWq7GY
QlqdAO/ju6BdvoreqraTsksAPgkwsy+ilnuN7K4QxCy+l2Q5FOKZbCVVxNXO91BcJecb1I/dwQBb
xKzMHa4O+m+gRTxTXUX74AMyfUbVd/qyrHyFRKvvNNwfJosIP36up3nKwaKmp7xG1S8K6CdZlvG2
1sdgitvQZhWKyDmdV7x90PXUq3k1ReuCECs5vOuO0ytQDS7SVir53ydxf3N5aFI9KlVraJZ0WYEr
S5O0x8aPfRimzgFWKEZPjsI4ytZdq3ruVJ8FWstOkz/WBQ7ov1tizUAxXQ/gU7kJ6l+ODmbnasNc
r+W9Nk4QaRXR0uTvJ7PQSTiyZVILT8ZW/v8oB0yDDBUGXJ6y2HA6FQ8+q9lWzghLACcA0R59/bkm
Ksbqunn+uvU9p5o7C6iNOM0q8+M/MB5UXwyn+B7H3g85H38VX4OCsOGAP3nDoR3A1gNvDeWQqU4D
gTj5idHkYWM/C/XVFDh2UfKCwQE/EYbjkgt8q3TEKsvUUJeZPax/OtEGa24Jex4kZLcOvU3na0gF
NdUXCht34tMoJSrEtDhLmE/XhKc93vWmBXlep17pnFQjZX/zRPDumWGyuQ2g1+ksn935nKV1q9Yo
6FTZWUtBaOniQI6MxL7GLN/kz6rN/pWhuH/jq3cJDmPPuxeNI4dXIgtsXd67mbhqT4IEEkJ5ip0l
0zIQ0JXeGTjTUfjPI2ZxpMm5vFDI7oFLeE2vcCkmL0Oe7YBl2B1B1xyxZcUvwASXr9CtG1RcutkR
zf8d5nNJkKh+FDCnAKcZ7Kh+btzdPjosvD27v5q1U5a1E9P9S8qc8B+Y/qo7Akw2qS9Zn2XFiOxv
DjUjMPA66c+zZmjeQVCvUuqQSpHXdI3oq2HXlSYtDHcLi4/oy2846MlR+aEqAlKbhRMZw4SFwquh
k3OFnovT7VyS1Yoj2rZ3JkQmwrdMjDPWtEpLdl2g/kKAb0eDz0Z0iYgn4YMy3Va42b6a53e7BCVJ
ntQ5ilSSPlxBYBYWY9E0PmknUAemoiMyvBo3t9V4mMTOLUf60XSkg5vScqGT4je3toeCgKqTDzt7
O78xnp8vdpwUzdBzX3IUGItLVxlt13r5D//X05v6A1wd7aiDXgbG1z7qge62/aHS4/PPhd/C6tEA
co7XIURfl86+KhJI2jTx457TxiRMItspJmppXQXHZvs3WWlkZywP4h/3IQRuA9ybv+WZIZr8NBDk
GpacDLVAQCv1a2gGpZ95OQrmXu02SfSrjxZ4f4SE6Jgn2xuG9nY+sgvGDpdpCrG3Zb+xTmnO1S24
aAwaTFXXDZ7Po3GwU9gVUjU0gw7CtZvDRV2afphpRsYWKz2YiBCw41h8oJ9SY2bIoKqDDEWqLEtM
+T8SXEgDcoTXZx8HrNhqchntPRMQryLwRAWyTDCTVS+Y1PZcU6DyZs0SghH6jQoMxZQaxzEoqR81
DAqIG4oNPDVB/1LN6HeopV2PN0JmqwBSfIOU7ZLs1rGVM5sY5RBm96CYQEnRuMWC0KNfLMFaS7gW
C8DKudmmjo7PX4r4kmdqrdYOgyXbG0JzkLHJfOFbEKwjucNefd5fG7ebwTwRCVt1UN6YuOnsEa3y
S03+qa/3ID3aX5c+8aVIaB+xtQqvsanXwvvyt8Yron7ySB9kgCwKfVX2Z107otbTFQmUFMT8J0Dg
CLyJCgyHZWxUPd0aXqdDgFoJSGruSnSgVV9BasiVsR6DQ6fqHKvNtWmOirHbQn6DlGqjeXbH/pOF
YlEg8ooLgiKcJ+Q9zNnRpuBitUAWnp4JkTxO/AJU5vpbMGnxFMcdz16toU0vf0kx9BEro7273mtA
4E8GKeKk+zmsUjHpLQLH1woNDEi2JOp4ZwFsPT79V9O5oGh36CpnAwzxvheOxzqw0tptk0ZWyruI
S27vWIg75xkn9uJvlxGw9dwhcz5NWPoC6oTt8B0E6qXZU999OyIxgGiRmMfK6vOFeIZ8IKpZwHeZ
iBS8VQb0bgHcIlo2FyxOdv5l2icEIKYzdateU5w0pv/z1SfQgjH9e2Q1eyi8+7E6joO4NQhxGHb9
4fayhdZ5PDjMkYriQAXQ47RYoVjEZFxlTkhlAIRqVXmILWPIZEvlu3mp4bEPWBOoghXseVWiZk86
ZdaMyk8vX5sPc1G1Bz8J0k6kbaFgiaU3jluInoofsQULmWbG5NlN2WawJq0EP/Fmczt1+3u9AY6V
Nn6LMundKhOSxx5XFDwskv8CEog2am+Iyd+SiBQxprNBgjXgtQR36HKuFgryCTKrWS/gUAAXaJac
8InAdHEbXl8vWzluRf0wPbhbmtfbOV7sT+WMAig+F6QHtP71hMX6pYz4bEvHuD8BxcoddYj1OBzl
kC8AuZarfnBXbTxdF0w6cPwzRM792UfrtBDqmdDv9aHIfcKMoKf/AfOgMwqgix/D/TKHJ9CNk8gC
unnEJ4enX6hT0x39uT3wWf422y7ZMrWIR9EUvwIjV5py+aBU4iD6VIhb/6Ax+QFFWWqhspXdcjeS
t3w62f1+34O6ktiNGZKcvsith//Y7tKM/tA0dfPuqDcsw26DteG0mLmIQeh4bm+kbtKDD5AtgmaL
Ps75GU14hedXtZ/C2hPgMrSEfM/ao0+ovPGPHjCY7eY4pr8K4URb6CAn1uAqSVs1No4IMu8HX1Lu
1opEHN7QgP+eOW6vIEQJMp9p+yEo3O0Lw+6cOQBv6TLoBJ7dvVftb/RrmGdN/+oRIkhfjCiImoJM
c22JxlpxCahFF9HPRRfCXckCJHmx1/FqRSH9mtio1zZUWXC5qi6KVaJs633rJPyHzGcwffaCzsSx
K05hobOoRJiEqrVivZfu47Aj5B7/RrjECXRPPcjpD2ntWz7Y32eYlJQf9ufZx3YGs2LF7d6XuIrm
Qg+VCFG/FFlk/2QOOrB9u8dbyZ5KbcsvUHEQzCYIC0srxcZVA4ZVMn5Tyf09eTn0MAS9h5hP0hFX
X90wd9lzaTNFrdg3qc7hjv1o3YvfRhbXI+dyU1C+1qfb+0t172dvZpQUjgh8DjitCG9JrdY0d/zw
Pk+r36tTdOrCmZEzQ/h+3/eUDUSQ3UcnrVSVjy+ikZs07aHXWOWYXTfGAG/H5bYLZuNPrqw7xTkj
01GpaB2RZ12M1D+r9h1l00nWafRJxP0ek/7caYFHOtsFH7TRqiyJBkmJYjw7sL2lFCdYU9ARiIZS
EFg6G1LV0HAb1pTG5yTpv21H6MZzFhFPdfAZoN6lOsA+9CgLTka3gN77WbYy324+A16BzmtezI3k
1MnulEr/91Kw3Ab8rsm2Dh3a4BkWA8aCyRVX9IN9q/2hS/Hw1A7VGuzPtvEuzSzrB7PQiOfh84Y+
fEUaY0l4YJLbHP4vkaQN+TQPPbS7xesTsUxPo3OiDIydg/2UbpGopmp46HF1141bDGp0VmxOcKsc
P0g9ELTK7EcjUphPsPzGAAKm2b+k3ARyXKGg/di63TRT9IuOaHp0S+chtI2tLUVaNBqUA9dDcesC
Hx4jv05yBox4xm9av+83hrbmD70woVoVJP0dfnk6kGpGctM34PaeM4j9FsOsI3QMBi7mzZLpo0Ud
c/cRJOjHCNQspJzU4KpKpx61RDVmeHDe5z/OHonEtP5EQXpg3wQN5pPqQ/rxm/df7sH3a+Hx3Sx6
IrWwXcB7kFseiVDk443oCwFuZf/dRKIGqcO2EkIsH3EGjpb+Q/f7HH7/WFyU63nISws0J+eNJPJV
pgNWe5tIISpoI+b0P2SakAU7aqJPCIzmnG02oR60wbyDeyeOVQkZLCn5sKWt/kAMVLso8C/iISFR
TrmCQv2nl2MJeDf4FUT/LYZFFWJ0aN4Z9zqsgRwNM8ugqMDIR06kQ3H1GOMitPQ1kXFLXNbwkhfS
VPJH5nxougjienSgel1akgusEPeuX7IGbXcBnx2M6Vjqb3O04urfRHjNWOqnK/ZF84dCOlsBiMkG
R/8zMvb/C/UlNgu7Y7FqXeOO+WqkngiXb0lmImq8gF0NnqtbthYFcMUwNFe6qxD1O0xWZjiW/VZJ
uh8PWfDhn8Lq4tVZBLNssGtDJXV7pC/JCmhIKKC7NkBpTC29JPz6bEN9u3TQ/xOGYU6lYo3TVx1u
dTZTNBGxftmn1v17R9H1IdfQR9Tc1AM/PfEmR7rHyHebo30GFleGN2ce9RKpqWbrdRloO0pVIWLF
UiAydQvDbd/8m+EfAEqYDIinLTyuaFHVuvKn9np/yoefN3jcft0RXKOdj0SCIfWmg35mp/cA5K+e
U7Hg4SVhj9jNi6FxqdB0WGSSsaWJr9NmS3+c0GnGsJ57CsGqQ3NSWiAHKPt314d4761ufq3m3Xd7
y+upVUQdFlThDnB3tOv1Tr8JR9+fWpqoK2Cr0Y+fSPMCYUIVq79ZDdTZS4046PvJKWOlqMHwon0N
TGBiAqs6SbA9nHAfVCtHsI3E/tD/YvAWukaNBZ/HAneKHkGKVfqEDfndn6Z1pOlehsxPlXilNLZ3
NZ7G9j4b3gDyvqHv5HS9L7T1JSylkjalNNbzrSF//BFYbGaLtuhP3h3AvpPHkq5/oyPduRa/9gX8
th00iJjDB1s+KIU2loM79VfHJQYWBXAz9Ry1kNQZ0kkdCazXeDPkGRVWcy+MAwd/IokESbFW3ijn
5tGm/rDJQvPJeXEZJ1ggc3ixsf9aXPgXb4KCAyhbAWGJ8UY6G5tG2+MlUlcoz2YKcqkqK4QmHQkQ
p+jNKasaPoz0lslUWsf5YqDVA+dXu8KG4WB4PzUX20RWyUmrnJrCXhUgvWHhq9ncY4/8cy2l2sb6
Z50jpK7EzGD5eZnNsaOiXEEIQoWnsALW/q8TE1jKKGH/Erq7t9Nfajyccn1nlnEp/ET2zE/DkxMc
bGxZqp5ZrEKyg37/E6XW8kk3yTK8lZTX+Va1+wkuGoCZYWx6b2H2YGS+zwhZu4iRyUKG8cqWVNJB
ZPJFqMaPLyxUJm48HKT76uV0dqOJYP9UX0plUFDdo590mP3TvpFvhKUppgr9H4nfkPbMAXZCdE0R
gZMSaJsFFEpsUunls5y8tXbeyDLmWuXVj8xr5mukNwtzJhi3e/5tU2McynPzdC0td0Mfb3UVqTHa
hLJlXY+23NAfH63YYSx3MYQj/HEraq2VyQyRhz3AmfNpsn1KIeULp0oRQpCd2wwOMd52KOnEarqR
H7jFhI1vUdg1kTPD84Y2rIm2aG99RHKzsAPsOpTvexqtFQ1f1aLuD7ZR6NHY39BKna40HPnSH9H+
z5jn7boXajeYxPrxoxCH2oVL4gIphyONq4NmnXTnZlfWikFhTcEvDKi/G65xFXou3kPQvjxMxz3/
lVpyF9MLmV0scD0CVDXVMkfgQ9EVpwG8PJkJYTPpboyA/RWGbQ8mjulXMxdAn5bdAvGFndbGaZMR
bhgnUR5SVbISeOIupdDwCGBQcUgN+Y+S1H8l4+vv+UVqEXbFtHuX3uZlT4qiXh+9c7uX83LUnPTo
GR6hxjbEaFXaHwV8pxvnO5nr1GFtvyLcWNQ4m/LpCO5Mv/LSi1EKvcjqaSl97a7wPYjE0k6y7LL/
Jmq3otHjq1FlbsQ/9GivrtHrbLr47ZDqEG+772uptK1eT8mHhDOofth/itPomHI03mkUxgXG66Fj
BaMXCuKncldt6wF2/YFw9wu7Y9yNEIqAIu2kRgqmI56yfex6NMl58a9Ef+8k/kFGYBZbyULKel8P
usQqQpqi0DUdEGm9VrRPUiRXGG8xMqdXaOrHyh8pFh7CQ89kTDRHL3v3riwHpVMxXcWx54i6FytQ
XCC2P/vt/WxxTXlCMTyjzmkyvJJpUK54/KunsQzTSp8fAMngjwUATUlax/9ae7477lkgRgx9BdDJ
UQ1CH913+XDDYlvZlQYnKXJWwGm0gBYTc5Y03zlMcxKZTxWb68ZEEucWvjXuEVQrekrh6+Al9j58
Ohuk3MKIizhlmvW2tZrMZdRQrtI/sKFGigM/Tr3Cb5NVvqfKGyBmulxYV8VQOMq7BFv5t86XAgvl
zwx3fOwqBy3XtiC+iVONlkc52ID8Z4BBHA2vhSjjlu/BAp9wfAjQ5XWmsArc5JBH4NuDCVtJf2KW
oaX6Fgprvu7Ubyyo8GuwmeUQ8jImQzJVnqtQ5BB4/DoOR0WxQTPp2D6/7QxP0dCf+72Aes9adZ4Q
34Rlfq6IJLsWuWyRBsGtW0uXL/du0xxxkcKqlQX+ppi4u+3Zz24VsXh2QiRDdQjLOKz4SYyJcDvC
5N7PpaVs6yMqwWsn6vgmix+2p8M6jpndX5yGM5VMgkjI8q3AyscnmB0+6DA6b6PWF1zW2N9fS74f
0eNrPBnRZjT/Y/K5ohd/rUS3whV0BTT4uzBBwF2QKep8SS91QNrumuvEPn3T8BwY36Cta6qLqsak
f30b1tzxV5B0eyUp3gkNKsLDOc4vn0uY0Iid4Hq4Ovwi7l94eeKYfFcXW6WRxit1DV71I2LtS9PO
xf+bwVItjz5vmXeE0+hYNJA8CR6CykK69vIic7q7e82FScfmWY2hhliLMUzkFrsnXn9JXdXDLJAf
DmXOVWqLV3jmcXg7b9YzMhtY6utBkvecvmWgOgG+OHVpF5upfYlRnnomxkaKDErNWqbodHZcAFtC
bbqsZb3OorZHqGh7tPeuJqEG09vCSobatlQbplTBq2jiCFA9bSXXSsDs5diYcFHlFAUAte/IQCQg
hkuICmHm0o2QMKpcLGMMYE3/Eme3AZMMTmmF0sfvOkD6+forJVSKp42sv1ZUx39pt7i/qda6iCF0
NZO+UHlw0zlpZuHkQ1XeZPEUCPcod+l31XfgBs1PIpo031JQqovyPQlPCZGKBAc/bBsUbZQImBYx
D9O8R7IGjcE5Fsk9pQpuaqqRcodpLgbQpsxZK936/hrOn3O3iMLtEhSXsq5BSnw9VK9vfEdgrCB1
2JIkKwjCzWYgtOTzMOhACNQmNqhGSq28TnB9uIt/z8WVRys3dGujFHCM/G2ertvucheohg3eGP4K
93G9m7VMa/UrHzhuG+RGLM6/RnMfXl5vbU3HvK6YJggbPu9YU55l9R6BjYBz8lQCY4MOBw9rLs3b
8L8Uf8A8tLD25M0/OakM/MMf7tk0wXqcFvmj+NfK1Pfym8puJBVlYdH1vGyxo/9hw6VNCe5Rtyjj
azpiNE+FI0QMeaPPneB4O7EzKIJ5NVT9WwdeVSM/i8WzoH+orhtc6OOHYa+hAl0FBZeAKbCzcfgh
gGwxEDTTd1LM1CEWrz4/BLOd5wq6sFyK/fUYWWP/2+kvtHRocvUmC52T/gvNptsbxBJBZ4l9npYU
EE5HR1IolZ6ltF6sSCu1OFBt65yeyxQ+pRw1zRCpKBDoNSRifDUr3r22hJs2ai9uyEdltOymXPO2
j78znIvLF27OEXqdkv1jGwVDF4Y4GqqfTmiBXrE9OE9a5zfWQhulxUidtnb7vHh1dWFtpk92/hZX
f+YsP/cK9rbzn6hgeOzQZZrBbthV7oysH5/oeF19mEz62zRGM3weHvDDKw1AcQ/y3g6EeDtbeSJv
S0XAec9fXn88kVJmEn6Jmfg8XXK6UEJr49NMDuOXRXHM/ut5rn5812pB9M1bJFIM462WKb1WYyg9
Vzisj8G5LlKy0AUJIDUC+kD9FpZyc09m+BdMLBX+Nltuhuc+/b1SmJj7v4eyf/uetVrN8aRlBmkh
AxrMooZ0mOHDfTvRZZG7ObqZrxFZWsByks1Ws2zkUvsBspMNmvDtafNigH92xejSnjVcU91Pe6F+
mge44qT5IddNi4gV/B1T1wze1yNV6N4N7k7Xm01MTEZhfPjm0lRh9+LG0S3swrXrSks0S/2hf5/E
UaZZ3cjuB0k1SRdkb9Ti2g2Ks3T0hVDyWp0R4IW/0ZMzwr5gFI5+v6GbgmVEPxRKicIy6I7wx+bQ
rO6h5hDrChOedTtZCS4egSY/4KBfFWK/QotDB0A16/Mo3pjmcz7AYEZm1/mIBCJhgZJFvzGTqZ72
eBq3oOt4zARnuB+2ybUl1Xa2Eq4LoW93hGJdnh/pWV0mpK4XeRG0CUmN/6Qq5vbn1FH8eMps7X2l
/V6eQEo2932tGCENI/vOQiEvpzTHKbhCcFgou0MiTC8jEtk7s6xmLnIiOrM6gH/tVubB+/OuQXyB
4QYnuCz9jqyjb/W2AWloP4/W3ZUn/VKJG5MBrVPX5ek1iRHCwbkeRVYKsbECIFkdQYT0O2yDpZ4K
rWJ+oyEXX9mxoiY5RfVesyDPLdVnfEtbetX4bUONkHwOR5q6ggTLLoTEY+KfrTCOSnsEP+U3uBy3
9jrfGK61F64GBH2NbpHUyzgjGG2TkDLUorcYmiyK85TbeEA4YExDlxAOtwzPNM82k27v/y+UNRki
218lbz4G34Ek+pC+3B3RieO32lGj9TH8/pfP/qxxDv2nCimh/esuVYBmQHpUpdC2JYizZqXKeSAT
ybZb41NG7YDEJXOkpfpZeMKQKSnY1ZW7lEBb7B3nyEo3C+lKyUr5Zr6JTivgkfes7LTL1ac+bjeg
sKBzWR2D7MmnpfQO/WpvRHkk1cqRTH7UKOONg8r001kVU+wxKaCXV4eeTRRYBkyaPDtbtk2L9kp6
O3UyhJCVqvD8rurK9RAYtlTFB3Jqq22z2a3etE6MWzL9i1wBDIJrYRazzIbPUDTqzdDX+BXCgjUy
7OHhrzSvACkEJiTdx3AVh2kBlxjGxPpVuusQxu0JkBdsDegVYjMJdvyW6eloNiWeAFsvpkuOp7xX
S+QEt3eRsXUZBXlIbmgU4k89jPhejB35A2VKoW/5ynQ9nolYAkaae2HF/x0WuwKFmZN6rEmrd/Ov
hZEpwpID8qrrG+yibYish72VQHpwHpHW1Y+l6QHu1CmHWutmChCJz89T9cTPW4e6gLO8gVpPq6JR
HhCoEMNqlCgh7sAgiTy4lCHON9Q9nE9Vq6wEnRbwhJZrCz44z2mlGfxuxzipV6oQK4yMFInRFPg/
vGSBsFaym/vk6/d7P09NS38zT48m/qUgBLTbp8WKGSUBm8JEfVGU2EMRiRIYrM5XKtErBS7zqH9m
+MChhjYadGhVjIbUVv/F17t04SHD9EzuiQHmIemoe2IegzlVJ8QpSVzwJXtFbH8dZClja6E9J0Al
Topil/4Qxyw6tC4D4P43tmTFHxRLhbj1RDOW1f1BSIPidNBDINec49vf7FLh7aJ4/7pjY55ZDTvi
9fv1Bhi27ogKCtsvI8I9bjWzLNukEhfj9Wabcrq4GuSv/3Fw2nU9sguc1SAaifC09VU6tHpLW9Nd
1P72VylTNvi/pgSVfESnUrsZFBPKqc5ADganujxKLdL3ZEa/unJm0dtdT9RTMOVqQAP59DERMiUZ
d7roC4II/doyaDILivgITH6od8QQY0cm9JKh+TIqObX/vL11ZFvWVj8iZnnJqxcpt1TxudDNlqCt
GLTd2l19kG2Z/hqvMyM9kVFKHTJcSkv+Zs8nHphNZMlmzBgm06PGTp5gX1uLadkc/W0LVO8QBWvE
7DIcTpFwa8BFgzRMRqw5tHIApgNHgr6b7DWkT5fwcGz3Elj3tjy1m480Sax1XDrAUV7d6GRXNH7F
VpCVv1MFh/kg08iQnujLBTZa8FiJU3Tlm5wi5pupCi1Nh6MsicD1l+Lp8pjzJKzP6OnjlgruN8QB
k4MfIhPsK4GqUsqvGXEbaEc8AABttOcXESr9WcEKwHrtM9A6H/MznaGrgjB5tTZfij+d/6RK6KEC
0KWXslm+fhn4KzFcUGFQkuDES6lyjlbXFR2+e4jWg5THrRss9qVJzx7BStwBNKPiMCKTSegRuZ73
r4z3myPaAgPQ9vkVGoI19qw0Zn8KGbiYJJA4eOvXit77owcS2zuFgOTduVJ3DwUrF4NnO6BgGo5h
WEAPyIGyesQXX910fpC4LsTOvMLXL0sphF/pzOOTxwpLeKS8Evd2k9ZrAtp3opna/k18UNDE3qah
NVxZE3/ywdJOSV9Ct3dPwnG9zMZYLwldmJfl37OR5UVZqGK0dslBj138jXGLeQwO9QtIAXIF7Xjn
8LC0HXEiuIg9Rf3OJgXCskxl4TNbf6Y62iUJbCVyzsj8wQdn02s0hpvGbRrXkWzOJEXwMTk42NSa
JaXI8nuLLPFt72NAKhiXSHyvYtl0d1HTVbDDHaY7MSpJnfzF51vJ48Y66G+fdw6OSGOBMNCXXAzz
ToDMuVRSTZQ9t721cxllAghH3ulmj5PBW3My2NnJiGqSAtZ/HnJp+qDgXGklJQy1GCs+/P8SFKLH
iLQoNBe/nIRzRXsvsNopir9OQ4HiXP/WaY5tNCcsUc7rssvw0Gr71jte2cqHgFJFz7PvMGfW50+M
WeeOHhZbCSy73l/FjvpsUenOHyDUfbsxAk8YNsN2cKqUX0dpfX5e2f0+hYgLoBD4zej8XXhIfhr5
o8eI9Qr/wPAiftrZl/oqBjWdsfkqJr1FiH3ni5wtv5ft3KvLnVecTVxLoFjQ2s405/6GUGgo2XXm
25nOpDnxftP/OeXR22LtK3V045kofTwziadpvBXhS/G5ms7UySMhGouIKb4t1k1QAao0fvhi8XA4
0yrmXoaAqkbZHXOE+DEoyxhVRP4QybR5Q8IVNPT2C14YhTIrj+yfRZYLZoYZ+ODpwnfC+xCbJbBo
7L/KrskfWenX1/+0+TZUHeXkdBRGxR8vfhE+l58dRgfMgRo+gr0wnOkqeCjO7gjyjoehiBnhsgZu
uTSn/vcqGft1AHzOaZkdGfoA7RyXrv/HppltTODsoiAQUOQSOBSAQ5E/zdiVPJJhltPgdfk7BxDn
MOlUtqUrrn56yyDNQwpmQ/Rx0Drt+d8zpuxo6gfNLBPu1fKg9Lah7lQUkLRjwU7OHHhgpNZS3fyS
DrfgNadoeKnwQXiwL2CBPkpigFsyWEp4kjiUUrDaqj+EmJsYvFXjLH+7W6aTWvptyEJJFHLx5hGd
1/FzOQ9MrfK2alCvPO76oQXwyofs0Lxcqe/ipUd1yVtoVYEkLeppbLIpUxmSViuzYI3IzKO0+S6H
YwH1tMPvi9Z3ZofFK1RT1/exBzvCkBl8n01vBJudrJYrhuPPgvDbjFTW1eA7nj4BwJHochqiIlN0
Q9nEIN+uF2IH2B4c45V7Lqw47vummu5PFgebNIHezZ4iNQ1qkblJJHcNH4/4nOiEk2LpBi6r/Enq
eNfg8FoaaVflfqA9pbDE59emz6txS71P3kFCAuoDCsSAHtWGrDMk6aXZ2dd0dHrznOLPYjSxKUPP
3/Cj2RkPdFrHZdKbf224PpnW2oVfXnU7cp3egH2ye93H6mIMZH5e7+Mi7rDoX7TP42iv6dDEyGgZ
en1hZ4niuoY+Fo+LyxCerlfitB9wLUw8opDZwUOCvU/CgEjril+nD4+iE6VEz0zQedCs4Hz9NpT/
t3VJFUGtkiuk5mFK/rSzZCgzNB35ZJ5/nI2GZlaHzW42LkLyvjcb/fYTfNK0TrFQF/Sx0D1Ed/Xa
NxinTDVGPgMNMGYXs9EUpp5xsSzhnc3cVBBIdGR6HSoxbWMtxgHBmn9GCnhqBi3y+8SchyBTkXGx
wMmLhO4yQkxJg4ct/NK9vHVuUfEFJVrrOdsP9Qwe9eK0wvxFXWWCHmroJ/lBWezFA5cs6gor4l5I
gONw7coMNRlsZE0Uc4TxJ7mGkL6byQbajhz9jz9c/v0i7BngpE/kNp7Hz/VxL3lm1nqBMpFUI2+W
NgeVLBtB9VB8edJHdMKBPrZrdX4mFZmNdEzyqTMlNCOLzIYHXDGR0V2JXn+vfrjdwHV7i+51VQWD
BCHqQ8ysyYWNXNScg8cdKqLcSfGk0AcmPfKSAyd5fgve+KtV4wHPVlcKNaQJ95pqXL/gxmmnPUbp
fKtbKM341en1rXAp0SZqWTIoJkXFfA6rh46DSC9LXvjx33r6Pb7buRK3tXowHBbBPvuk15lEOows
lDK9PsGf8vBgRpmv8wHj+hFM1bXD5Zp7lT03Ax5cXY9yXHhwDU6EddYi8jMH4EiJzXaZLPyCaKa+
k80hqH/eoTzC3R7DDd1SeqgNrltNxJUSyHc7H1k9tfItzrgWNsPsAghOBnVRMXhK7SXGEEnhAUj+
lyKEoQRklm/jBcIr1eZdy7adclTCQiQ5LJ0dPBEb0kiWARPxvT+JgFDNYxJ1nCSl5xXLD+MvpcPj
r656L0ndWqAaIA5TEfReWAxS0LTxHoUxD/bIQNiqLMY4pRwX1y2Ur+e7Eo4pMmnylv/ztq5Curui
K68u3QwNsRgzWkAZrahdsaK7isrbwl6zkSavt3fg8QcLTiWop21tFsmTD22jOs5qpWk4x3aNPeOR
zFbpaVcnBqezUn8DAKUMmtTjaL8M1jHrAeFCa0He0MmsHoavglGd1Guriw3iLjgCF2K0nOt+qOFQ
2ZHIYyNd+Pv1EpNT9ZpCXSrQVsVEPVCmwM/wq/p9Wet2cpHm+o/UjuEczmdodASnUya6AY6f8Vk1
vlyJ2ivm+iyQ6PyRerVrAPuFVBTJ1vh8d8n8Iispa5QBP30ZNOcRNvpF7RYt3tNbV/QhTPBw9+4h
xumRO9LleYs5ZKrqY4lFeIuTcIolT+z0ghEGed9z5cuNImlV54f3gOtti2k3oNWYt265QEprzaOE
ra2weqEMPjHJ8+kf0QMlmbn3jTKVtg+wLEadvoANAEl1fSyeVF8EoOijT4kbjWZn2JOddrSwzoN/
rDPPQQe9nuW47HCZ3kduqEO//AyFrzU6ySEC3Lwb4P6O+7MEKHGxHPz135rMHUlp8+/HWwqc6f89
3rdLRL+5ubUA6DznQES3p7JMnp1VjIy6HKjZuqvr1zITlTHG62ziAsX+vVD/PdY5+LG+XYgP9/Q4
/Y0Hb9i/Q2GGNtL5WFCK756Rzb7a6q9Ui8PqXmHoKLSBnTtg3tAxCZHobya97UsXHdH9H8mrKEik
lkAbYKGxPkLL4x5uuL5Zh3Jzet59blTUZoqZj4cFoxYVoWRjy2dmvUtODF95EBPEn/vFGECEvqUv
aBqstKFC4cS3z6v0xwjuwyioQWJdEfzeIYCXY4XqsozFbah7n+VDDPn2qsiEtLlDtLHYWPcXYX6g
m4Tfb/nt/NrGJLpPB2Sj9oXCC0VGwoBaA8JVRHkk9ZMZ4EHP1S153eol9SNa71ElpPVg7HmK5/87
bHYjPLLair8PUkKTQFNYZEdiE3r2G8kDOQPF6m0gpxpjOdfnEQ7xokdByrvXpszMn4yY8iMdhh4u
gIjn5j1wdRB1mrHJVDunSvYdsxMau4NSE9VlgA6DGK0MguVk7aNE8g19qj8VnPzH7ShrEfAif6G/
jLsS9WP8oRB8pX/Mn3G1U4hVY7JQPlQ5u6tbRxpk2tpw9VqF/tmZIsE5ZkcwUkt4/a1aqy31RXao
4R5CwHJ8VPCRs5pTsrOENVurQ73uz/z9PBqcVWVv4tF8KDQ8eApCZ1vHPMqpl1JQa7vcUI+rp4ze
ii3AEBuN6PKAQTAasY+DkXIEyb3CXVUTQhpRUehsNQHHsZhemSwd1ITveJPlAqcyMo0zhRxqHir5
Y54t5kgYuxD4sXCGVFWOGI8xvcc+DTqc+drLzXr1rpAtGd2abTt/qe8vHfow8Dj6wGIDadAX8wy7
Jhr8V7pWQv8ld/KZIAC/uh/OFCfVQacLRh+lhq8vZmmu5AFILmJxEtqUYCrH+az6srzEpsrcUn4x
rjBdp1AhGVxCQIbZKxmrUtvy43vxoOcW00XJsveJyL/BsmIfB72tWMtlkz3dAYKkEkHUFB0H7sbJ
bf9fmmihN+JQ6mTLTv3wOIfojMTOuIkPu5dUS/4DA7pqL8Bgyi72Iw1NybZFP0/MHx9+H9H4fGc/
ynCjabw7LkPTlNYe2PN0ZIRXFHT4iVs3VgZAe11pXDX+1Ikb1PZ9IjMmcM1cmgXlu2PC9ajO7Ap2
CVSLcYLtJ76DB3yH6wWLSZChX+zUrM4pX+fExJvkXqoj5yXSmteff/rTALauDR9X5jAyW/8d976D
YXFn2gngYvQOU9bzD3JdOwFSpklnREQUEOKc/Zo9k/lj3ke41HJkycyupvd3QMigOKFWF/rCEPyO
/z4adr2JmXTgVhgjNop/SAELfCHlst9+D4mQH0p8su8UNRFZu2HRXpXu1Gmen3de7jAbfYXSiD4k
cbtINjcsuq2QiLPRRFEwfeWyHbp6BbvJ7+UCt1pRrDXO95vpzwoBJ9C5RXfhgjRh3rbetKyWfStn
NLcuuYMKtQxbkUskHACJnpyTX24UgXqCqRyytRJMs03UMzqavuksywVKwQdWa6q0Y4qa8WIRW1L7
aDXwCBW8z07bEJEJNhZ8XxWrdF1pchW0VSuuxHEaHSXKTJ5DTRM+ku0/IoHth8PnR+kD8woeZjl9
RNlbhEWgqeC73p+kwGzD6Ind75w3Y2Ha64Rwhn/GltT6/kObmyr4tV44ghFyNDV342wHFxAXYbnz
7+ejl0PqF8obqM1ly4G7gd8iiFKd7syG6Unhf82UQhztQnGkm8nSPJYYxdbXfIK5wTX1v7s46VUy
RL7zD4HLkBsFlhbkUFKGb/Aus85uht5nA4n79xIYF6TyLbBm4Hq0Ez5DyRaktCHLlsmc1AernMsz
mEqz84VGkxzi3kE7dNxhnnkLbVgc5N0wS1oxiS+8kNSf2ozl25r1ShQieo8h+hqFzF06YPx+w+SB
2U8xbMy3vZMgKDelA3d1i9tZoS70QXFEsQbji0J9/snwpcLrd9JG4uwEoBk6ngrY4wp7kNrKxguf
WbFrK9OyBfnxh87EQOl80mZRpGKgaxo6HzhA401pcVrTQZ5IltpLr18eHcstevCk0cBOEakWzHvY
VrOtHrupC4l7qJNZLes/5ImIU9ZoBpTODOfaV0lUsS65UfIPIxKoBuhVC5fh/hrRTyFlBjLZeZO6
b3ULB6o5FgNjf6rxt48Lu9+Sc6unez2H9XM6RZhiMV0zSifJ5F1jUFFUH5spxJ6yhAkNedwZwU+w
9c2TiV+EeRtDDKUebm+h4Cu9cOynQTQm5JLhIvbF6ObdvEfWZ2lobzfETT+7F7CvlCMF+RHJqEKl
ZXJO7O/Wrn8iQIvNBrf1epUGSmrhg3lJzy+FcPaOH73NIDu5TkEyXmJ+6euCEHV/9ypcF9dK/YbY
96bDPldzi3FWrpKc85/8Lt3yKgS5rgYgslVX0nreGNF0vy+z3TaZGf4cmn//F1m9bay8mIpLWHCq
+pK26LzU7RWzNRmY5UWL3LtInToAztefzGwM+S8u8ABnIQi8iLoGZwQ6bfce7A5Kn4oaCUwbqOOP
FLXFDl94Gx/W86jcstz9QsneVaeGTHWLcqMGcnVXoJuxlk+E+vcJab+oN/cdTVqjZHEz/LaKrFk6
Hmc/yq/tKBnrgRp68vJZ80Z5E3ABtze4nelWadQgEiuUsjc1cXkxypq0v+yPa0CDyZW+FNbroOvz
Gfik2GU7ZDOYTbXp1OlScloZYu+fj+rsvdWTReGfN8UCkXJBqeatKVTuL+eVXidijDPME9P5cfZk
wffKn7A9si1CnfwdzUJVc4Wp3ygvqqvKsaQV9CVARyV+LmorgrhwLMvStmTAvDC0qojff+bxxNq/
ycEVwUSRi5x+vp/eMt2lvb9ZbBxw44RJ8SuIdhJocX40mNmOe33tkF6qD3pAcNy1N+9K1EU33riK
x2Q1nqAlpopPT5v9Znsuw9hKgRvO2SEBbjuOWUebmEtQb/wx8bvrjDAl/ONplNZ9bKu4iN+WlyrH
7ZRxgnHCgu2CQBAO02yIFSPYpXE2QOvQ5ck/6EDBO9zlQq/Q0EgxejFcexDRHAk3ND43S33hionD
kHQKZf74UjmDVrhmYgWLjbW08SjC1gTJbkMJz202ye0iZQkCNL+wdWsO1g2uZ93MruBgWTFG6En0
MuUd5ERJk9YDLqVcYOYQSE4+PwMs3SF3ropHuW8lfNvrxBKM46CcD88WeI2pEFC2drNjbKb/qgi4
B0S03YRx1EWsazWpxTs9uYNPAFZcfd/QFlxuHysJPwxA4nyJ1r4WlMc10QIUspSZqkzkVOTiSWok
jHYIXel/M3DG+twA0zoLxvTiM192nXKT8Av3OSTnpoQbFz5J6n0sKVdcCBz4WjvzQN51wc8vJBRA
OkJcldpVY0ooQkL+AV3rBFNVAqDngCIpE6Wss/o5fPyU3prMnwNegwQnVoNZ2pEd1bgY7wMCHhNr
rScFDIeECKm71UFr+FpW/LVWVYp2PjKb88gAS5m/UPp69VjA1yjYjNeouM3iYGfdSGTY8wR3hLE3
JgNAu6YxxzO8SetvH3iXvkqY/XCOPk36GdaAXMS8dYPlzXk0GSVHcbuW+wg+06vMy/7gqAmby2Y8
R6rKaapAbIEOg9obczPEe8vo6AAuRFA44/i5Db7EGnC3J4XWlP90tOSVVfUzeohtnbM9UTJwz+Qi
o/wJRP9xG4rRpzb1oSWFoL8hAgNevwXMP2GGHk+hY4/bGeYSRoBZ984wyQf/r407XU/dVmF6CitN
uTwQLz0XAoRyOCBDNwngjVceOjslVbXaRJEMRWpP2TarMvbHn+rUPDG59/ZUNBsDcOisgDQUwI8U
JhxRVi02qqgN1Dsg6nkGTwWN/WVb0234VtNbKGVRZt6kEmDIpfODAzUleMF9d7ZuqFy9h5Qtt995
Oe8wKJOSoN23yvO/2N79uIDrV8BUZpC5swohtI2KnaWkmP/sD4LjC2GgCwv0eiypRKczg2fnMMQ/
0tZEa7l2uw4+5Fluj5npwbSOOZIS7aYXZgt4s+GabIfO3QRZD97EyQa9t/VCp5Uh6ZxFocNJ9l8L
06mwlkBj7Sm+YmNEGr1exjIV3tAxfrZld1DWgAlt6ghDt7NDR7cfvd1Df2Dy+XM4fsdBbrjiPY1d
QNQ6yKyFolKlCp7BCxcw+EHNTap3wohE1gBaZAF+biD4K3ChpQ27n2lFmqm2axc89YuhBicURDNZ
6iFGyJ2+Ep6HZnOR/UI2PGjxkqDxz/Ol8uVgEnLk+y+qY6zhUhEnHRaNtCfc697AZQnC98pvmTNZ
mTI65l4Bh4rpYT+2i/Zkx1MpLQ/h+SXkUWPUvVg1FKFZZt0GTQ7bQS0laWxG/8HFiSI5YM5kJMEX
uXzLgUe6q6mGChnFsEC6tM7IYMCIfZOakI9D/BifNxXRl74fcCDVUMYMSNpDfleJ4P9XJ9oL7jYL
K/lT0oU2OvDqFXlF+u8GCfpMHGjOoMurR0XEpmgIej8I5h7tt4g4a4iKfcj6cMXg1b/S3xthPv00
r4ETyFsgs3eEj3oZDtdM/OfeNZ1xpdU0v2D5aa1v3RIyeM/TjiW+uMdpcmh8QE/CmLdYzEjqgFpO
axPVzqPZTu75xG2RuulmcnyhGrIeEOjn+b5mNdN9yKlq7Jci7v178jZhWoO2A1cMg6zWY5z0RaU2
r6jfT+yHLM5gKc17k2aF0OJ01/lXyg2v9k/s0XqC/S1pAYl0+9pnL4H5fWy0astTVq13E4Yopx+1
tMoTRkD1OY9kFS14u06o1uL7Yub4DEver+mRmi6GviFCB25xc2ytI8EuU+qZABRD5JgP0phl3pb1
YyOhWff22gzH/67owoibsv2D7v3kjDg3wcU2/J1u/nGxzjfcuOyjvmcDADdscGcs5jW8jD7A4+LA
I9tr0ob5sP80SXPEPDpG9HkKhz16iQEH0agIIvh1MXk6kxlSiN6HHip6xyDC16XBWcQH679EZYhm
5QZdbcXW+6leQeOA+aw2XvaK3dGyEVob9z/4xdhuhUpd0aNJiXp2n7W3c8FetuJv32Vjvj+P7MOt
0trZ6MLjThaZCpw+SrpVTJhi7CQf84Rs3mO62L5BMyAP0UTLQ3cRtaMHBgtri5SgXN5w6n7NNn8x
UP2YPwkSxE4JBVV6VXoXp9ZJ1FzwBowY5rN1dbUZsqh+5TDfWdAfy48I7AquvH5xLpx5AY1SE6Va
BZdYWrThJYXmXTgaJqAdNSfROgc0OFGqS5DqlyqggTCSY+gbVMLhGeUgJrKLCE2XewaFZIh1E2GP
FsWIsjcVL3W7B8okux/KPubyc2p8RsflfHbeqLMdVWVcNOCwlhBlS0KessttRzzyQZPjdjAPc6Ei
wElMzLYmLxFzuIICZ0GSNawDbKqv/61b9f7mUyx8R7eMzGP3XVaDFgecmz/rB6URaQ6gn0REGewE
xX5jfm4d3yCQTWR6cd+OKrA9Ja6I6npNHEyi0/d0DQZ2qAFQNO/amLH7O7j6+FaAocY7Eh12ZcJo
dPBUE5l6uBTgbt0Ig5zTZFEHfiSD8Y8+k084FGDlcSvChde3paBYPJm+S2w5pTsup6oq2N6CgeXR
7ceoY3iHHPuyRSlnDedfoANOFAa/O7jZ4HkT8AQQw4/1zIHFfuPAK05KEpEzRe3JY/9lf4+OB6Zq
8PB4iH6YrUWrTdsF8FTIZYA9NAPRVd+cs2clEznfjvnTnyKl5h3H6FmB8XwPIc3ahV3LaUqBqImK
sbjcAmRCuQP/DByIS9NjOg5D7dr5x47adYw9A+yARHZ7uvEqVzlUy6XWfCuoP90SPXgNcjejlS+Y
pLwX9S8RMZZL+6Ua/EVMgbn/JijsPZzB40lRT7DViAZ6SD0mI3rWJKi+LcwZVdIlRD61Hq0aOzGb
A7j1zb21ROzI4pFbe2WVdEsVEl9uX7j2HTOxiYgk2jC99tTjfWNX/ri9CGF57w0yHle5jTjREq/I
3dLsEkIZ4O8ay1FIgSp6Ygewn/z645dgmaqFLE4kwI7sbwxKAYRp+RiKVx5G1H83x3aBaeBnIN6Q
G3O5LRhbzjJgmilIpWSU3fKZ8+HDpYXjvs6tbRj7foJAG5MJtouPLAPcmjTp87RfcGP1jBY4FtxH
xUUy9ZmLvdC75xfNkGx3z8fgj546HXTxY4pyasxjbNGbbS1VFJk0CJHc8/hEXMZiFv5Z+cMznmgh
i3zpXbPVoOJ1YVRByVLnGaHFDAx8v8szYyeiccxkEiDC6xmZ6YIm/VWkBb2UaOyJ0uF6b8jeA22u
m/pFbtvawclcQ3CskBDwxhQkImvJNcDLfqTYXayG9X68Saqrud5LClilWVmyQDHhc38Q1Q453t9f
ktXAt4TewX67PzBwrQAx7s8wcwRxhu/BaLNbRN66CO/UN+3o4U/QC3IQg9g4gd9Bnfo6tWJ6YykB
GIu4TB/3Yi2nbCfrupLPz6ukwFTZkZ8uetFjXlkZ+M2qTXON8LQ+oT3NM6gzoyv0p4LzdMO1/qXn
3XoChsUqxWfqmUKsyd7skFdE2B6TqKh8QtH2GDxvxVnt4zhjgg7vavJMAf5JqrwyqgshhySpWcDO
zBlmUsR+q7MkCHRKGSzztG2ly9a+oF1WE1TD7Nsnp0p4Jz1FWrA6B4a+IpF6CvBk7FeObLsSxGv2
912QFbPlufaytwTiq9TBo8q3consB41eAvGKBeOh8u5a71amp5FkJjxpapYnaFpLN0UJaqr9HF4w
x4t6XkY4Eu+JASTwVrBZmfxIYyEHGn6ece9up2nwTv5xOvaEDiLSBvmVG9EKXnB4UdMjEeLsestn
gBQqqPhThLw03edPHUb1aWvNDFTu7YMrLsbCfKr4bkGVbkAPFarypYB5omaDb5gVBo4MARBR9/Ek
+MqivRS7ZOE07Cp+IkZs2yxsMbsiOMZAvr91uQPh4094UJaXghZyFTwLIHSh1tHirZ4ZEC902LW/
AkFsXasAKWXfiRcSk0Duso3GvM6S9Cmw+0Ph353pSCyXrOPckF/Ph30E89fbJ2XnayPXZh0fcKe1
Gdxa3cWITXQjrhFaLJrqbm9rywbsNaPxcaNo3NW5QAXz4E9T45/pZ5qT/OTya2OpZQ/+Bk/JG87v
O5DYZYlBl1rt8/CUwwG29hZ4EsvZmaOlZSBB/jYvJd+REzO7kcgwAu0fBWoB6F9FjIXuz7a10tdl
YOXdM+kdO/aGWgOr8zGieNWVowhzpZzw0ZlLH7698YfHU3c4tjlYqME4yAsTVn/vdUppgnE4rLtL
gBvJ9+ys5IMmMQ/JXgnA9CMCM35+XtvFCCv+BEeYCO9VImtqo8uuhDv9XzXPLZV5VzIHVBW980TG
oVaI6fOz1ncU1MGAYXKTXMobaL09/cdK7dZtb1+yo3+gqPJCZirucDpStP6riv891JBSNpdW8eIh
nUvN866ZZXpfPxb1eccDhHUT7lS0PCTqLTSLqngUMLxGt3fvGOfl6JkKiaj2T2vQyKE1CvgMNdXC
L2ygjAlQ3BvMyBd4pnPIQJrglmdfLJ3Eeck+OTWh0w5VGyWjRgrOfI0gIu2dB+KNJ5Pgd1J9P0/z
/z/wDkSdgiKsJVDIgRXeASAvIPENZJkbhRS5HoOGCCvuyCf/psiFJEg/047p/4O5Ed1/8ai/rPkV
gfFMtQR/SbtnfxsQrkMYNMQP4HdAgBhW4PcHhJoDKhm9tg9EcPjM300DPFvrQdhEJ98Ov4dr1MYJ
5QkSXPmIXERtkjTDxsNGX+0Fei3or01RhcJ+rIkeOJf0liMNgCBIGD8cYNHBmXjYh8p3HbmNTHbJ
1rvRBPm/n6Zb33VifVUJzHyN7zT9zliWhIDva6rVaAI0Xx/w2xWthCa7UGX9Fo/kRYlmwTFxeqqk
8eqgzoEiv9XERWJhrTLTcKj8wzUqp4z3x7zJfGfbe7QJC4TIu4BS8kEa/CgZkTrE+YKmcPHXmP8Q
0AnTMI2CMQcfjfMJ08JSd+FFvS6Fbt6PAjPoqrh1HD3rMq4AJzu90sInBe3i4vRDGLTN1qLhvTS7
M3KMbLdwFrF6HHOYU45DXMqFdYsAcMAkfeZkL4/aYBvJ2GrcBmXbdcw6IrlOwyFP8ItZR8OexYr0
waTj6e+uSJMYNqgBFFtXlNnDfjlmsrNcgChqaxHSvMUpTUclHYbHwa60Z9ktAv621+xo00Y/1of1
vb5LoGbpAVJjLu1laxu1sZCPR3SUUmLZyJnUHroX2y/BCFW33eqzKM1ujcMh3kdakARZmEuuDGXD
Uq2zpCQ1hJFxFIRZhj8Cxyi8pjjDAD46+CEkXcQfUqSRPSfEQK1viLWL/2i00jQUhqO+cne4g6bj
mIfOTsKcYTEN5/cUxRwjKSpbFT2gbHGHo/sFEV6aqCEKc/KJXl2uOtz9aAxtbEitZftfHIdHucAq
6TWfbnEk6+r+nyFRIYMhpqtEGRQifA9+E/ftT/1/8sBuV0Ye8yMUVgEff2Sj822vMU+2BgsB4glo
3BftL0+ldwp4iMs0FRA594RvIdA4P7PsH4zeNyHHrX4tSqhjIOj0oNz6PzmHP7ue2YGbByh923LS
s3koDJnom6Xv+SF67E/S7sQ5/7sS6ezmQUcbMB4BpzLG5lCofUxz9dCI7EA1u0wm7SNKaaVFnQ5p
BdsT8QkXHXErnIkkJ+9ZDTMQKZZCvb9YbpY4djjg3AKvYamU8/b7Zy1c5CDif8yfShPUL2qOXrno
dMs+SyBwHFQF5T9SwLl8+H3QZbqAFYDaSFnBxwO4YXpdG1zm0YURwNQbSqEEipdPUaNA/JTdJdNa
l0jRw7t9LUbLJHGPw/xixqYpEd3NYHyedCkkCphzX2GWb3gO3E0v1meU3c7B4ORQlSZBS+IC5klO
6i2Ybv97CmKJuUjJTLURkU53cxO1AkSlsvJ5JIbYQoyyf6u+WY1PtDUDD7cWiT8NWebk6Pkeas0e
PPeKVtlTVxOUy9GhPjYmr+S/sc+7aS+0CgqQqJFI+B/aExKnQ+lGI67HMZVhtq3mfvfMW+OpSSjD
j0OAKt1tbhpx4RKzGXAW6mWrqXy4o1sXNU6xVbTq2XpUWPCGUOVAcr6Yw+PraU1cVN2Yvu2g+9on
4P7JL0plM/prNps/Og9hyaxWyl2BRlKCJ6TM2DXeqHT4blOtqeb4yj3SWAlPUkHakXtCDqB4yn0c
lQR0GQIDQDKGLxPCloWV1GIVwQ9jzlGFTUByltJF8nE7h7tGCxCIqNV66knEgJvnyIu6MHdHiZNs
O5ht7Iizq9KBCDarx6GtMVG8XHVClth/VwsAbzSqmm104DRJKPPOw547+qhzOp4J23CQJJp+UzU/
rDnhdTba8xXxtlZdXnq+Y/ukX2Cnn0+Ncws94CSZSWrqKfitsrCiSrIvZ47Ks720FCYaJpjF4km+
olt9rVZ3W8ZDHYRT9NNrsAj4ZADn00nYJ9kSoGsp3zKlQu6/vUmGqGHh0XIVmEPXc3T793V19qU4
oSNhoagRCkZ519jHBh2ylVZx00LIhVBC8v6BX+dmV5R8MEPkigxWWbim+d7Du/a+f7Oo4j0qaLuu
q1Jx4fwF3L8EMQMzVMhxWrgA/N7CPuXVcg+176ncCGDhIZljlqxVZ4tSdkozzOpUPdtyp7hF2gaG
Q/xbue0AnkikUci/Hrnhvv4fPtctbNIYj0LAMvWwwxa4hAIwAsDOAV5R9G3lZvdiVrLaG3ahdXXq
cDdPghU2OzQpE7zhE6x8gePPwabCmZSGGY2MaDmCfL/e6SDmPVx9cwhVGu2gd58GOK1gBtS4125m
Z4fgCsYOAwBBCXyQBFFxw7ZXEzzVb5J/43FdAXr9Xi6/kwu6LS5JOHXGrBIWgWWkP9EtKsTBt16h
ukCvX+fFv4TXGe3JSf1VDdsoyLuspQdUmImqK0thoDBoUEzK1ZPzgEM60bCCf5eEPzL+ugj9+JH1
4GBSZdK0uxejvsj/5R0p0dFfwlcxWN7NOpU4jVxIVr28Mgl0iGXlPkvc8FbdyysOwUnDWs95MX00
YGPGqiN0bLkawz9c3PxYigdagn96amJs8plkb4yrvLBzKf19x0KYBZ/2EAcTYzk036hJ+5d4s/qT
//FU74HuePmEKKIzJFXoDgRXCk0+OSjlBJeZxPxDolwC32bVhWJRa1X2HhUl0JIH0EmfL2LdrdWO
+12XKy6KTijO8ocR6jhvvQo2rlKFFl48VGxHzhlsuGK3wNsIvqffyceUGoW4VXfyjaqYrMtAmeI4
roOAyhQJF3AqeGkKwBiOwf58FGC7Ew4nIHjZbFLfQ8dfeaOpI3EKMVO36M8GCkmQCqBj6dy7ulN1
Q/5O36Xa/mFoBuEfxVg78fiaRq6xJBwJn7iC/syONyAOHqsIBh0rOErFl1kUgzTRD12s/xEvW47C
vVMXX3R/5qWDoNGV6m/ZIGLDq2fob7SKNI48qkDPBd1DFQTIxJHqzrdgHZJo6ey2p+qNyZ1/wPH2
PfHRvXiBYR2bNJSvq4dIW3ELFacm8Zhq38BZd4U/jhwvzDBQcVE1dEYFVgxo06XC8By0agDd937l
4lQQriRBNnQrKQ2jPmeNqQoe3yNPzeY7J3CWwtOfK32kvduHnmafjFdrUlsQWtSdwdplh0xikwVw
B15w7mh1cjd2o8lYVnTD2qJQPQQxzhcfJsaKBlSFAz5EMsWv2mwKi5DezKLjNTj9F/bGBY6yT6ao
5P8pMptSL7IMWCf8ULqSRj+hOBd1oMzwE+SZmeVTEY30YRAbqHakq947XXhArQ2tT6LklUXIckU+
Sj4WSOTjLAgSO9JUJYmHN1HP6LE2qOXUj6ARjISCkOYVvRDY3ZkhxnueT9s8R3wsUoHN+IOvZFYZ
44IZUMatbqmgfNbNm3ABgNV5vAWBrknSoMvnq1qF9DnNybWCZKTh3Ta0QlbRYXCNuEfhU83qgWvb
Sbm3lCsMBdcuf/3iRzWcOVvSisW6RTq02fAaZrCJy6dYGGFdIR/N7u8TxoiUR6BoQ49q/B6m6F3t
wCYXj9n14q2S/5C54sKNJ0Fm1EUwvG9aLd6/8eeR6ZkfrNmmU1lCTP7KnXWaZxhdwUMMzct1jEgW
7zMemAKi4zujmxvzjq9hWlHO9eE43Y79tAngwTu5u++ebF884qki7Yk2re+dZ7KBWixGHuaj7/Ud
hgo1LyOi9YOKT3cqgEal/qUBjpyzaG773k29kPuiO5tomFhL8YapGhW84DivjwjkTiLLWQAZpnts
J+H09m5w81wrFldWBjPCliPfhufmU3WBMtizWK4YfgII2yidpfej0iF1J6907zqCb9c5vFTco6sT
lEsaKxDiaGD5ZPvN/f1Viyy1EA8/N7LOGkWDABKTqxQAVCEQ++HwT5CiGP2yeBzLQ52fpftJBwBk
4eE+MPuP8hVWarYYx6kaDB8ZcDqS6E/+AivA9UDhdRiejiUTZqCdMjER8WdYjTMcmvCiUFcgWDnn
/pdRzILKLN57FTtcORlKRnYTWICk98cINyh2OxZGOSaq2wvyLBUAJ7q0OvK4aZ5zWLaziXAk4Q5I
kqyKayG+Jg0jebBI/97tfIlTU4Ct5wYlX89jTLlIe+HZtdWfxMoPfJungE/IyoYcWUnhL+3fOr9V
6MnFJOlp6z5Lpa9THKw23udDSbMmuc9El352BSiCOQkjLzQFWnok1tea2YcHVIdtlpzlFrSwO+fy
ph77ql1JIuKL63ombVTzoHZ18c6wsivB6b2TbGaYvCcTVXsn24lNgQ7QCY7Ma+UkyxHHoOAZOMoV
PYAYCbo6JdIDwADyD3RnIdBBwJyQwAyZ8KWkvzk3MXHrxkL3VeA1gEo4RI6XPn6BHHHyu2nyrGq/
0pb1+D/O2rylBQ5GVPAQ5E8as0jQaX/GE88wFEgRijl4BbZco9mfAbPYmV4Uh8hh/PzM23sI4KSi
ZJJSTJHLMGsuuY+BOl4909OZgSlQUuK8tc0/pQ0ItmwvLS92oAzgpkTGs21117iF3Haqh+OqPoE5
xXhNJhj0sn1bnESXrmK2Ox1HX9lI0vWOmRQkQRwTmU39SKmQ+TvD2CNnpx5Waforc6Y+y3t/VL9M
cNDHbt303D9fEvpXbojJOspO3D6N3g1ljttBHeA3SJ3XSt+2LLpnTkq3kUzAzdIjeDs1zRo1bR7u
HDpsqP6qTNMXzKOfmjxdTuu5IwOYYem7ehw4JOvmdjW2eUQpSpcqnxhyW1rl0pIOQZngXzluThxW
0K7OeGgcAxeZ2ACEFzuvjhIvWeVHxzdtBTuk6AqNg26LwGAY8lVgIRuStUl9innM/DQtQ+gh9h0G
Bd+ux43vFKNv9dhibXaOiwVVKcYQIo4Iph9gMEY/gYyAaceLY9N8PYjG31VLL3V+5yfzMABjhkRt
faPX4U0D63jPMMUyQRB85eX7CQrIQFps8qHXciacW4g7BsH+VNspmpzU4J3VYsrWbJAMLvDgHz2F
PML4NwjuK0Qi91sxh++Dy2m/5qKoGTsaA1580WH08bUiGmzeUu8Xl+Z1IsyJm7S+FKM03K/89iN5
/13aZRYiFMVSwhCdR19gi9Jxj10yxU2DBCdFixvhcZ0kJCHMMe8IRPFO/RUjc165HiLxLQKwx5WE
v1bfziK+k2v5wxUhUJ7UMaVp5rZ6zRxBmguFqiLGCKeWmrDc8Fxo92bTRKVVdlAZNKVgQjrHf8Ru
4I0+qK2EhcLcRMTyc6NLc+2DoNo2euE2dIOVauCl9gudWbEDvQKRp2g59OnGCsQVhDvRArLWgsEc
xMMtSWKmctbJXOfovA1mKhJ9qOfZWG2/8kbGt8DgeWFYSRDykmfahp6HEnpjcExnSsJMfq9fhb/J
z+C/kqCKzA5iahVqmCpuh5gOb4Q0b3lr+m3xCGDeTKmz2DbxboBrxylaUw0s9ii+4vJSnKuDUq4z
gK5VY87I+uUj/o2FnEiNrHOSHiDzkPgJsWgTQMEdJgiCysrCpMC6WifMAXcltarV4DVkD9lmNLri
c7ujw/M7x1vXOOsD46CkJdug/46aTHtFtE71WZI2NXgFZ4w8iUm0M4nUuSBfljW16FGhkrF5vqu3
ZEVUsjZvj26KV6f/sbJMoKUERJLRBUCNyLrLZIUoKahgJxfmlN9bGExuhgNHytifg3IsnjM+Z2mF
rGJcBiNeVPesFdzmldyKwsFDZNvAgSQ4U7C+GMIjLWdchYDHtrJGRwSTaXI1wTzAPJt5xwUuCPfm
k9jSXDDPGKCR1d4b2R7VZw9KjtOgjioBI06a9yZ+7idpNVLryPHQVg/zN8EIPnKl3eALS2i60eeT
gr1brCoF4uKTSzy7n76dRBEMYDWMhmd3d8ANdh0XzQadKNpzVViN5Nl0kaZW4JTGnlAqa4fRkkgN
Ph6OG8L9YFjRtcwoWIpyr27qQoRDRE1JU93svJV8OKPs6SbAP7HTJFhILbAhrhjPuSR7yGlpr29G
5p8up7ILVONqyEYqi4JOc1eM4AmPBwgjPhQjvFGu/sYMTO4S7Piv0DOohCubuw2pAxn5sN1f1+fZ
p8Oj4q4jjcsw5o3ZrfXJ1CityRgfix2+xquyQyQ6J0eUkkV31FkM/NZj78s5BMm8eoLS8ddrX/if
OMo0HQAEcV8S6tGGn0zSmUsnKYltvwJ2nRMUAkjIPNT3fHQc/DLfBuRQM4GYrd3j8fU6UDrMy2Ee
VlhYi8GpKps835a+aVm0x3nNLsbVeQArMX6eUbHm7TgRCnhfLEEMmTTGoydRgv7NlSrB2ornAYL3
+e0yE39j05y/k9sAKU5Cyb5aID8JqqUmKDITBnAlur3QdTA1cB/wynrlZpqdOkqxNf4ChwwBDJT0
h72o5WibQJmEdYxnZEo7enxfUBV3dV2jMendB3B18KJiNFRfDnCiyOWNDZUFVGI2KVpdqw3QR2F2
M13yhvX3yC3X3/CWep5SGMhdAdFkXznGWW5LFDZsAUtKaGy8kuhVgJilzIv7DrNpwuzAu6XvLFgI
NN7lhEyA0KGgAGNciTPRJBwDFdQTdZvAvxviFtj/O+sXQkWLv84SpjOGTKbd/iE7UdqNXEnj4cLL
BHKEuo1M5e9LIAWhJpbUYh2KYXn/i4/LAnPf01b+1SnRg3+BwYDxkPToZkvhgORbSop8Co5Lpid/
tAzewk+ie9+ObDFuMcqeim92OVG9GmGGYOa/Pbf8agBRLei9yhBXYFOUCrb1ULKF6sgjbVE3Fl2v
Psfilsb197JgGUZRn/hRRYR6pMGKMF83oAkNmF3D+NGQ2ebG8IiMGMgEf/PKqauKnCLbtxBXfSrE
E8NvGriEGIn/sfnCnlBoJToj9jcy+yP0gg1mBKyu2Sbo8pz/BRt2GfhBHxk1QSUlQhdpugDDTWcd
ku52fcUV/t1XruMRdThZZ6GBQdVUipLC3z1OWINaylboZxSdJP2RF6oE+jp+GVAvrwJ32E5Fs7nW
MsqLnveoe1Nmt3/K8Hu50MG8GFCPmx2WaGYSXsb1R/XEuilY7Is9S9wrs6NQq+z7H/zVuTh11Nhg
mOcdF6sjVAoqSMdsHWv0y5sM1rYvqUHVZ8KzYEmTZGPRe13hrQT63i5+dNkljafFNmUOKxrAgCwJ
2MQLb4mITdMnolb8zzF2AfCutNClpDHFWb4WNmebq8y/qLJ0GJHuPKzoD05gWp7KpsrwZQnFoq8X
kKrObE/q6MGen1HssUNsFtZyY1hToXIKYhAlIBFPg9ynzvZCsf1ivF6kYnJGBIDUdLm3tcFnDSN0
djxED56Wy+vCvoCH8bc3dOy/qGzhJC9Ka8iAJAIGrTUKPBYq7MF8lPkxn3+PsROpCRqkexQrgASM
N+vwj8F3rwi9ippvL2GNixhuNvwv4HUoys/EhJighhyOKPADsAHdMdJUwGt2gjeo6U+tG5IDXUz6
fMyWsW01mEH5cVZXrs37x13MQoZrfIyCPl1qyNaLuadac4r4x7S84mNuWvXzp/0vnK/gcW7/ynTo
ViXbhPh5OiTu34UhiEI+2rPo6h4AfS6KFvn+hdC6z6vx8g5Ah6yJGRI3oQGEx27vcjjF0LafAutv
oAOrAkq88D0+nyFdhrOfZuuO4XGC1vV86+YEhuVahm79gubCEnc7J1QEA3UmYHoI0eddDNelVsNk
+VpUNVxVIqdFHv62VdZekpGkR7XxE/twBMwR9iv5rX+wPaQyKxUMJ+XD2PNUmnJMf0IJsh/sAOgI
Bghf+TjjjKJI2y8epyNCkNXkuZhzqfOMU/DW1Y/kpcSxMwbPoanUVYNRlAG/Ln6R82cqMclQnHpj
MtvDuJMjN9C4Xyacb92Cy2LzMayQJq9Mus4rgGkQ9Vhc/smQmh3dz43+70Gtr4piYZV3nVD7b3ZM
FRmiAVZrHMnIOZWTiL7sQ5f1JB4sgpBIhBP4PUWrc3b6xfuZW24S9Botlw4QZkGo4YJvm8cHV4to
Q2FIjJ9bVd6KJN4sz1yIIaY9qImLsw3omrAzveV4rdoKP9Oej0ctYNWEGlV5dAhQUT5vUs8pI0Bq
G5vogYvI6jua/3AyU6H+4kjOepXXSAatmEECJev8ecYisl5T+tAiGUp7SGJly2AN3QGAOQmh/Wwq
rFVMIPqKzC+XtL77qZC8xRbK1cddbNxQEsZ/+Fycatjho99+wF6kquXG14K5zbHkTULV5BFsXDfV
k7I3KDjPzMYRC5SqH85Jl3UriTd9NPz7+pFYIHCnlYrqxt23iHP9sI8XPyZNoqd4qlaFu6aTTSRc
V0n4s1GfDU6Sl/sdAEaPOROUCz75n8kzrFTysw2/VaZP7uhXqJRLLaLfryNEDNQr8ps8QPxQInVr
tOhy7ZeQpXCKyWixTLGfiNfZ+ud1qhjFaDjrmgM3RqiSGDTV1gffaey6ufKJHtYP9C/CsYH/I6Gd
Hm+gLRnGlJ6co2jhm+5jnNM06/jgmKzYj3IGi+oDUz5HQj7O6zcqwq3byEE+GjqcMpxvOWa7VDIw
C/Ub3VYWKhbYNYVqJTjfO/viymKZGH5l/x2ecrQGwLz97VGDw1sJK71Em57mbfLdKv4sdG8H08sv
ehvuK65KqAVTQtIVPAECxF0xvMsF0NVC984JLErXsGTTYdmYWARBXtb/cDuKZ5NFSsJiCVR/UC3H
eaiZ2TSllV+CWV6TblTvYMZi7vs2SFhtftvlR3NGHNmEE4oaN5ucQtnb2K7D9NRyGm4hXpQuRekZ
few9vV0ghCDCTRZzh+lErQ2JSUnalim54UN38DWMo5CM5Hz/WM+FKuEHY+OAuGPRWB/MD7paGyK2
lBKZgx2A8+c719NhUqaSZb5dKYyiFQDfgQN+ZrKMpYpWyMrphHC5AtvMSEi7CTjVtOSvpy/qKVy2
oZsjsx6qOyJXpMqpFt4FiWBHV8VDmxuVjFrvK+4svJ5JgNVRBYS+qhrLVJOu0cFl0Oy9mitlY6EZ
RMRQEsj9y+J6bsoezQ1AXxTIjcbFQHvFgNft6OwFCQ/mE3ksP2JGRW6wl26gRl7Rx9rIBaibEb43
drK/FhzuArb61h+lXQpbV7bcdlpJ9M6O3M6LSvZ0eJ2bhbOlVoce+Qt8HZ0FQ90ASa9NaAI/9N4V
ivnCgc7HKBKQinEs6PzpFTtZc4NJPSbA+TKtla8bE25i1ENcQBQa8raWfJG/hV7DKDuXU3kRgHQa
CD9onXzDW2TUwxoe41ijQlKpg0hywgEayMJKB51LT2jynObR+vQWmPqsQSg4AVVWGDX04Nt/0RbM
XMV70N+sx7OrqtpleKGl29C4wvo0S6DyFPi7cKx107/dQAFOGwV9hDn1Nk4GPbmV5c6AdAJ8P3iw
W06uUCVUVo7nT5bGrNdVErw/ry0ySfAz8GcqQlIR7s++kqXASvwOsUHVSdVnU41TjiX/767Hy+O+
zz5w34/Uu1URGvX9tBT4Azh7SNkF0bqxMnQlFGzyzQev2Uo2y3VjHxmTH7fSbOV/Dzd05uJT2qx6
1ASaSb+kYDU/pYJF+nKcUoJdtaUCzB3UD0u1tVAXn4Xzoj4Tip8ZcCGlPN/XQeMFCY6ry0NGYqjM
khtFtdhiI4nRXlsxqUhiov383p+crKKLhb7uHxKrOTDRV4pp5BY3DptKHWk02LcohU8YiHgOx0xo
I//LIl9rvsghU331Cll3WR95+Km9vCMxUpo/rM5DpBGpLrut+mcLonBi51Hig+D44uf12HuYf4iX
y0fWb/tNHoSnxEE55Bco26bu2pG0GKFUM+LEBMIwaLOOwKq5YA/iSlnCOg9BpVyv3E+dKXu5DrYq
4ig0b43//SKGDry/KyQMzGi49vDsi1fHDiiHTSvfk7xcbFNxltGb2Kp18mBi2C0UjQmvnq+py3Qf
z3qIpVxjq1e7ZAZ0C4wgYjyQ6JRdXJBIuET/enfUAvhiefn8Z6td2YPI/h1TEj/7QR5aA6nj78Wz
BoNpTcwhtfjpUH3mt0zaUF5L45jr6p8qhujBJVVtGgRyN+wvxqDdDahxKTrR09E+ixHnvYztizHm
1rz5R509ig0uyvEksaF8SR+GISsxCG4pksQocAZIA7jyd4Z0jlLIcA+/GNDpIdsL/lnSL2lLyBTQ
7A9wOLTzpAitzySxCiT1/zkPKRVt/d64/2a9voCv6AWEM8z4lDiXaOtOCj+0M8O5n7BI16XpoRv/
aiafcdyYXTnJX854mK6NqYJpi7/Wc9LXYqMFR5wdJzJYEyUCfJKG3QtMlxvQDP02SRAxd/vf6mv9
U1uQso01Ntm6g0GwqPxNHwnckU79Ok+tpooKhwGVTbw5Jme4xGd+50/4eCaIp9Yy08aQcxATR+gh
W+lvn3C8Y3Rs9uAMHVmu48FrkOlF7lhYN6gg4yqVzgBs59OVkzZCpD8TaFNejHFzTR6e95Km7BDz
9OXA0fb8usHmbjEKtfob/AsNLKIKjiIZsLYDRjVDTtXJ4aW2KfwbrepMuO02pdl5kxhoqlBXpstO
jvCKkubtstL8yJgAyEGf1ctcbBPQcTTHJWDoBm/M6GoMDPe3jF0duVlY4LGegoV5wIb/CeM4+Fs6
PecXwqVWFxZyYBtBrsxYlR8sB5KkUOBaAc91A5opM4cKT1A4VPrLsHD9K8mXlkg3F4kGO3nMaD1Z
UIi9IH91J0St/YbZtzPn3NWqH2cXIy8VDoh5Vf5ulVLiud/2IYcdP1Ux9RcNtHBaxtmwnCMTVEnJ
GP9dtQoKGoWysm/egcTGplwDA6cS7KC+RuOrFAk2Re09lsKHJOeAm/y7Quir7JEKSmfwUQjOkZgL
QiqVoMR4tB/RILZ0kcLELeNm5fiHWotLv039US7xydqk03eN9D1p8x4bbcq6tIpDaZLv6SmNNQ11
Ezu4S5bvrUL9yF9rLUWqdAp3eOJQ1pjVdFIXsh3rUfej8Hwulb3BkCrixZCSdu1xerH0kOcH3IBc
NApBYHCJqK8quqC5jSe7oxo6zXt9W3Vs/BtufsMX5249m5O91Tnv0bPB3ZkjodRAYP1gTw4Z8aCn
BKKmz46KqFUJaSAw3BuQvQfeSnS1eFVRxnq4JlhRgGIzg9TvRYAH46tmWU53nlT+X4dqeWka1YQW
/+yFMsHEboya9Ytdp2SrzUzXNtn5m/jzpaE9HQ5vIYoLz3xkEKM1nCxoOVyqOfuxqQ/6XisHYZMw
IXkSWQ7ArmNRhrQE9GXFwRuB39GQfAg+WAn+Vk+DBC5gCHGltqQSI1+yo6li6gFRfeADz5LCtRej
Rig5a3F9mtQcxnf6MD0c5hhhD0JEW9iLRcx8PI+/VVxEzOz0YhDxMtLKx3iTfQBXZuFJek64W5S5
V2ZGw/rD5hqRnKoQVRPbiPamHHxyhsnzxoKjDivk5PplSlGD31G2Wl3WwojSn2idZkvvPv77Negs
gnU/4yICwY1WDwvXmUAP/sy6uUJ5/VQ766MrUlowocQ0qrabyehIMHK3FkmbNY/S5ZVhnPAMZ0RU
Z6p+tLevDT/A+H/F0WYWpZPexjrU9xMeHekJKwkT+MPqxmkbqZ+WZCT6W/1YOxHxyYrkxawGQVSW
mJUr4rGD+gDGrF9moxH2i5BpbCLOgnAP9+T1Y8DSL3fiNCKx+YCdapcKDAMnH1C1eqC+NH/MRxJv
uitqTDxJXq8un/hm9nWS1/JOnKnFmVJC3Y0Waw4kM0RH8sVj9HC0SMttWo28nICuAHTCDh8ROzLu
FVQ1B6fvrl/aa73IeW70MK8bPXsIOHn51W5UYZJc2Yt5K6OcMKWnJTleTfYBYzH86H91Xq5fGh+b
coF6CTNL4XcthwvNSyFafQNzrc2WbHsNEy3n94iKzkG6d+9rE27jI00NHJjCncHeiGDk3DV8g/Av
+wS8FGoq29EQos64LEWuaDx2QM6Gf3LUyk91mMlCcudoKFhun6a2pvkykBNhK2RFl0NYfgCQBJF0
owttOkQfISetr6IP0U5c1fFSx5p3ghNTa8gRvEPSA0+UL4rt1wI4kJqqOUrtX0ozvzrQWCjO4vVi
vu65WQ+Du1rbU3q85Z0P9Ha0tRhFUBqGlOJ1+9XXJk8leb0KT+uWg6CfSw4hJk1ohal96D6QY+Nu
EetLMDam5iIAktMezlez++qe1w0XQQSygvFaf1PaHR4d0q7IkhASI6+EnU61U4FXQT2rRr3ZtQfo
UgFmLmQadcUp5twxd6LlQwhQ9tl7s/iXJIBUjWhkQakmA6/ohD7o9JftI28/Wj0fhCKENfVut0nL
yo4cgH76ye99kbINRswRQKanPppkmrlzP3zHMix2/TNDyfi7JHqY+IPHuPzBtbtnrfLRFlu/iJwN
yuvI+3dGVbdXa03Rz1KO4yHdRMGX5eOgnJ/3+rYYYnpqQQg4yq2nBweTovi0RYo0XDy7QySg+xPq
aZoQUvxfH5drB+uoIx2aywohclUhGU3xE9y+09r/MNeGtCVvS8B+eQ7D5JpaLwRnXsCq49cWaec7
Dj4EANKh6MNgLb4TxX/C935oq8FwRWJGXDsyw07ZJ+M1VNXi7SrYAWg0yTi+oEZKg7Al/fqfMnlG
zUfJvmdj5KbPakjTy5Rywp1FjrumaxCUgKsMvRnAKfUdxXceThMTfTl6yMJsSfIl/FNWuc4Ky6Ns
oYNfYALciYG/1vIfcTcvtLUgGbeq47aJK6j0VeWrbr7drStGlyF0RFDUwBkGF1nzzxqLFrwt6pbE
R3Pi+GgYGbDvpFsn60b0fXWPpEYwdGHS7VsvgBJUijq80NvgLbFxlWO0KRjY7TNBPF2aenlRtjyw
kGsP5rcOpGtCPWYM9ssxpKRzrCETKCbOjE5jbO/WRCiIEC88b4jRkuZiUIgRNsHxS/Jha3Kq4mjx
Zw6VVSeWKjPyRAxnsf6ZxNYqfxanCqNuT8M6NjASZOxax0tKz4NIYegkXvFohE+u4Zdo4oXrtnNc
ytABv9dMsdS8yNSOFu55C9UvLN20iGhMegqd2lDuDuXgKS0qvEngahAg7iI+EESlPW9f3xG6CuyK
fqXdggHmV/5jhx70r9rQVW3KXwxsfqfMo+dX7JSPw81rB5S9fKO/rcwPPu4Q15GeIUneZ6auQyUZ
CXmAAOwCGAJ4SkpygDL2Bkf4eOTEX+nBTDTc3vvVLAsV+kzgPewm7IoS5rBvEFB+xRG+IRp5CoIP
Gb1/kbEjXwwIdc41hY8yXtn0Fg2/+iQsFPQLodXIMJWO2Z1TiXe6v3I8Q+roYrjlIwSPI/+8bx0n
2vgUGR36wSj6Vv4DDdZNLa6SV1BR2fNHfm4+SwM/AZHNifIby93GsxtmM2BQ4mi+f1+o0xiV6CHR
DWVOBxMN5dfKskOXpeQVA/xHU4FuwiWkQV1UJL14cRVQgpmrxc6FMBmiyy+g/uougCVigS43pYEr
f6HruzYUnELjXjSYECWNpid4q90GhGdFS707ypSEs2iDLaA7r0SAv6xtDDGh6+M6bcxei3rS84zk
LoemYgwQC/4Yugqtx5Z3+oBKuN0fAORRGz2tpjN6P1hzxVF+UETEW/kIoDbpLBt5Xgl4eHE9Czs+
LKXjXWkbEpn29GxzaC4uNMQcZavucTAk8ex5QPvJBT0NVo575kmAJycdHLADS1Y20wiEECSKM1mU
4GFHDsLsXwiWazpLiBXQPuNZ6b2ZBbAbHBCat6QfbcEWY8orzV2SbUaC3qzJmrGP5fhZLpE34Aul
e8VItrCxeOd+i5SuqXStxyYTHVPyi4D5Vk1LtHDSI3QzPqSa1F2gNiYahaFYhd3BAMOZiL4YFDxb
09mY32SbG0tOLfHfuiauRvTsrVtH4KMtYB+4CH0mmoduEO+BiKZZNTqqelkyv33goyi2P1VNMSa/
h8YVcADrLYrnDLE2iAhNqJXnAPkJ/Q9x3tXmHiyvSGpNzgdt7DrXato9qKgdu1N91ePoPC/CnOxw
DzpKnsB9USekcQXAtuESjn1bwcBGT9AU7B8rwWFiwb7ZTZ71/HlKshKooAFy+Lx8iJqk2phQzYJi
FO6+Vtw9kWmFH18T4rp+plg4EKqSrw8gnIRw884LZ364RWeMvbnx/V7mIMrPvPluwQOxgAr4c6/r
s0V9rEgtffTSdZgNfK6VW2m6u/dDpWRlMcf/WVw/L+LXBoOVBG2uxxiFBnOzmYDBUkKVsHsFO2X4
baP4bllqTU0E8mqpc8HLsKykdREI4Wai3QWJHyiGWVn56Gmckzfliz/4qPBe3U/EySqMvSDiBjBD
9DAeqnZ1/ZaZlGS0LUe8fwhddvxTT+wQcEJdoEcCzjZjlaVmMI7wzUZXqDfReBjOgGNbgRl29CvE
SerlSKjOq/vvlLBaX+Mmhu57LBKiaqr6/5723SNPOjCgwV62Ftxqjpaaj1KVPWhWUzzrDQbV2Y7S
EScQIrRWOlb2ofja9mxz6otUrqrCaHKxKJV9ROeM//y1yXxHqC1DG327jHVzncZDt4Bcdh/+S6ph
wueltiEsy15dpg/Y+SmeA3z31+aF7UC/XcJ4MhXi5frY5hNujnAtpn/bNSHwtkPIrgACvpoZ3OCm
XmoV7RE26wM2WxrmbsZrLy+6FUVF2XeFnid2PYZeddIx9NBAwt5Bl3oy+dP74OTkOopkHpggLvLi
yWk+NteE+KmwbbXrygB+P8OsD6lqKFiZK8N70J1dpI1MXJCD504cs5R4EWm9TZr+EOBaBXbpYz21
uZQscBGyXV4nBDZiV/csZocnxHywtSXRGZBEDcMrCCN2OJbTIW7VrRHxGeqczOlDtxe0D/vwCxkz
Ais5IbNS/qs1p7L5Cqrp2bwiLjDOY3owWQUVvjOj4es5OOtMlNF9JItAgqJjSEbElnDPXQVoMzD5
juNQysl3DQ8s+rMOJtX2x7Q3iBJqJ/2M2HmjawO4y1+MtK4CDhdYplP+Xl2X6ZuWqOvNyNRXORmX
++99ZqVXLY8xS1Adwh8kuEavEQ3T4Y1zMXLqB9UbytrKiwusqPh/FbRuiB9xQnR3V/i0i2yV1ewx
MkTQnOZ7l/vyszH7c1omNOjmNXCqhPxn6J9GTRZMb0mMJa8wvYyWR+LREx3+aei85OIF78bqfNql
a6leGMxB+QjEl4HDBw4UA6+lfb0I35yhh/UtxftYq7GSFt0dRpaLLW3XmlzmCDprh3Jd76vmg93t
KCdmdQnjOC/K8Bv1p7ji/bHwhn80AukwghCTZj+ws6he5t4T2R/5260OT+GdLq4m1kMD6gl6xedj
mtBvCkzfL/eK10fq36fds+rX3BIWOeA1dzf83B4teAYq6mOqA4mcgMH9iOmLaoRBpuOO0cwDFbxF
gNwFM56fl54WY12JMcBEw+JReWLQJGTqu5z1+q9MFE1iCY70+M8arAOTZTmegy+5lJUEWc0tzoRU
fF6PJQLC8Mz9Gp/f7+sbiC4podUH/8ZenZOchHa51GOyP1uQjA7K1O6kpdg4u3nebvKqDC2lnwio
19YkmYNL6d9dSp0lJqXtwPkGLjPaNJTNo1YRnb3aLAIka20plqgvGbAHschLiqrK3jwrJEIhtacr
snDzRQ0J9p1kLvmo3d+Tk4hkT8fVjAnXnWwh4PDWwSEUFzSJSngGlB6ffq1DlWKeQW2FAy/FenXY
QSOqVkzy6ksQ/kQM/HBz41W413iWYd+NYUqfXkhs5B+FORJZAyQgzep2300CHNBWYPK8DdJQVoVM
Rs+QpNjwP9YBcP9n8ANdQDSf489WfC9r2JZQaZjQO6xlilGUEL/kZiIw6bb9tn24rPUrguG3Xa/Y
EMc3+gv/NhThz3FpJKr3hgNuifeVZbbocV4cskygQGAB6EeVmRJPjhRy+IMNbLK1mumSucZ4HIcX
YRznfUZOjntiikUMFk0biYqIA+P/CLS9XE/W0V2XClzVJd+yNCPIXE9UCGnoiii2/mtKE6R8BqDH
pn1IPGUKOmrAhNPdrU6Pb3SC1DP02MsbOKW/DRxyiCmoKENsT2dkLGkAOtIwnEPKvQwDOjS17Gy8
Houb2h5pXdISiR5iTtn6/JgKni/F2b3a9u3oDKEYBQTqixyZ3Sbcu7FwcaAhxIVuBgCcfzLX3aR6
x9y23jJEu3In7Uc/ogJBAZUkHCGFyG4c++h0tmw0Y2K3h96tqUJfELKjdJeNq9Qkro3i0mw14Kju
6jYBcgjr0ov2df0dTOheIcKRnTXqy29ZJ6eLT6AJzAguBZcuvxdPC5r9xW4D6vwyMJXxk7akIhL8
Hv9kX0LPRIGJvRAKckD6L47jhq3Aov/FChMeLY0BQ8oL9rQ+bZh3ncRSsjIZdmGfZuX0R+fC/60Z
tl3N/OlEDr7xwYrI9SyEN3pnQ6GByYUNLtGjrXnUKIQ3LxtmLEKPII7v4rp9g64K/VejM5wLMO7A
4sLbva8uOEKA4jUnKFy7VUSbCTlxqK3B/BTGNnRNQFHrEflrZtMfJjf99dCGuw77XjWUM+/LM1tR
svVGYv4mpvfB+6RN71rmI5sPR9x4CLuSTUwdjhF6GdZ5rKGE+his4/Aup/7Nr7FI230J772SyZVs
vmwJFjPnl61JXMBdw7o3Nanal5BrNbxlxhjDrsaCLWeP8BH1VOLjtURib8T7At+qVr8t5Fxs6OzN
rGhkgxnrIpiyiqBxenA7Agd5JgnAH3Obo1aIZwNSwah9qcksesRYyTpUAszvGVXAsaNSltqxd9s7
CUQWJYI4ElIz55/azRMmgWYMSNLBitiVRKmv+9+sewuAsr8Oh7gzct48Vn5WaZ8FabvaDcDTRigV
Cc33rMo0WghvpxWEcY8NRU0WnXY4YBwLR2uvZ64eSRyesJXFFxO17lGl8qs/KlRGIVYUQQPY25tT
MU3O8/T+1IONsZbW8TuPmqbIal/r+Y8zpwsh+UXqS+6lhcowLg+AjWuupyt5hG4BimKPgOZPg6gl
apbSh15BAoLkjGNWRfzy2SBGOdESwfxySBC3LSntmOOWZsJ+BEpLgtFe772MBDhSVJGeOzzJaJ58
8oWVVHJisZYY0MpptFZRVlueGKxjCiue8VDbsRJFb03rg+UVL3Jre0BKEbkT3+xa/aa9uBoWQ5hD
R5TM4XzYA0PynkjYPm1BuLCB8t9s9HSclFmjvZ8BMMTRlB/sTaQHGk89oqSeXVZjBGA1Rfmb2gCu
+BfQQvFHj1ott0Wqz25b00R/Z0wKxZM7t8PiPs7gvmItWFKO7iWsVzQ//RSGarvIuqH/M/u5Mp4u
PUxOlPTzJs0ZEFucDlZ8LFyyo+tg8SkolENvE9quANMfBCaJqXtY6DcwshDSKmnavGmO+Pq/Ya4t
9dAYTG6gE9EC3D7XOlrJNTbtud8ekfSH18X4uRhE0Xq3Lr3mLqx7u9ig/IZMObMkBAG0/HV9m46c
pHQoQRjtlNuAxm69uBEPXr1spFiVculEU/QsRbOpc2gnH5oNd/zvOiaTSKwhOgzyMDCk/PBrEJk8
b1+WpOFOC/I6eL5/CT+VXYa/S6nKydKkb+beWdxE1wHVXEzTlHLVmAzFI0wMtUio6lIRAmA2XYIS
vnioA4rImj1+YdIEnhvL75/4852WqwAK7R4o9MqbzRmaB/iISp68Z/lRYdXm7IkNtuly1+UJXyjS
K62J/wnD+CHKWAvOfToUlE/YbndFEEqAVfaNtR6unOYMHCp/QU/1dbHlYh+YqiJLyFtPHh9MoZPN
qAD5ZJYdhzB3hLipwNSzp28M+wnJy+4sn9tBLQGJTsVOxtiXL9eyzNqdXECnL7hInfIIfI8UAR/q
aQwfT7nPqD/0BbdCMa3UJKRiFAOsv30vbyR5MptRoVSmUaZMSd1fPKAhuYkJrFIdqV+1FALZwyF8
x4SkfCcnlnj/Mqyo+ZmXNBqN1T18qZaHmjifRs6FWh+qnCrtymmZro8rtJBPTr90gEIn7BGv9djr
07G4ZWFSaam6E16wn7KUv1Jh0H7wXxrhKRGUv3ilQvdiU5OcOxozA07vNbdaczYm0tOUAiA9BZu/
WhxTJ8yz6ZYi6Bigjrdixa3u1/dGlh3i4QH8cRBcDX2yPKVUUv+v08fCXdzGaja2eo+6D1RTkeWs
kOtApMeWqOirU7wWwnSXr9zdWOcr+3JZT44hsruCuE3swV/JECmfrV99W/Qmme9OXveCl9B7ABWa
aMeWKXGNqNHBNAKtYTWLUVWU34ThrcAZKr4OrWwkjeFPgqvJdu+HRYKhsk6q2G2Og7I49rh797o3
dNsmE6A0hMX30P5ZM5K81w1t0YeAyCm6xtBZuj6H1U+hKlHZfPWxYY0ZlcZEbjqBnIrxpwR9Nj4V
wWjk/Rqm2etaZWdYl/yJDQ1awrgym+7fEK23gi9UIY+vvepUy1bTYX2qC27PD7k75KLt5w3XCFQ1
6H4upERcXKrQTkQRiTo/13eDqkyoY7HWsXNywIDijfKz4nUjrdreT4yyesJTamRAQ4w2cUpiPvXK
mOBIDR/C1c6zWNrIgYUO97zWPXb+exTMJkA5lHj7VDh6N3FyekemR095CyvC9XhpL6QBIuLM2k9u
Z6RkyySWtRaI3fwtfiQUjc8ICPPIeJsGT4b1clXBiV3Zn4axU+LmBQkzTm0Et0VP3WG85uGTXAwJ
4sKwYwSSiz5wU+pw15oeIrgqKs3IxQkHloGWCSXh12CwyWF1w27/SkT3Af4/c2bA9e4r0QGH/nwc
zckW4nMWrx+jNhJqFn3ElRAgCgv0VGrN9wWPFz39+GdhukUifySx18mhpEZYipes06keAbmU/icK
xNN1jBAc82z4Xiw6SYD2XVK8p1MB8KNnt5OWXD3jUMeDV51YrD5UvhdxIchKSC2GuXfJ0kqXDw0E
RRArmWtn/zdBG+qPdYzv8Nfm3ZwPvAW0L8gCv4mXszysASWkO1ek18na04CCOBrMORp9H0Z9khZt
9AUeeNjcOQ0R42UGqm/jzVJy4f59pw6jzi41Hvj8YemaR1SPeqC5Tq+wRC2kNrY9l/j4bvTmuicO
lJ6HJcW60WM3k0m3sMLGqCP0h1QFY5+o9MLHr/JbXJzBtnVJNZWVf4xyE9yg1qUbbGnxFPds0jqT
6UBiiqdDTkFB56P17S/NJydOoMW1skgtDa1pdTjeTOBrevaWYI8bMd2C2jEJOJA6GZBAC38Mscyh
MyK1pNcqYZsrVb6cZvy9R5nhwkL7PM1ES1TczJBTd6MIl5fLiEoo5jg8llY2vrmZO5RZPjryFn+X
qYFrAJmOrzBHnPIY0tN6ja1MAff2xd7er8R50N+YNbG7WroHqq5Mq1Q8X3gFpuiHGRFpWtzBR9JR
nMsFi+m2RT213HsW0383zsQMZDDCldKhHnT3pAn6TpJFmOF8DUXOb8ZWWbOg3KLPVDUfP9gRzmH1
WNTBOye5um83u2Cve8TuYLXpCYgQ4phyuaNo29oxNEendg0khWXdYaCr2xC0Perx6TrIMBBQ0jeN
niCtLH0O5veeWi7gvi7zcQJrDHbxFPuPSshh8gbQ0wJ+Dvj40dyy638ZmRqRgLOrAXSue6TZWk36
vFkVHZKRsskkunEC0pzU6o8s2E+hE8dE+B2e1CUKW0jz1njtaJZXlybjS2okxsryVW9EPWPjWrWs
BP37CP806v5eSBkAEWeHofV+Hv10d6ry+rk4WEiI9tL9fVvKQnjOWSNi1FXuQSRA/8rXUTZsYKFR
bQ2OFN1UvVAp1KdD4pGEseDw90/rty4Bj3ywzST5fZDzy0LugqkPG8fv0gDFozBf1+pOUpJvRg9u
UONiXxeThzZBLE6jF/qxUyPx7cJ7M1jiRLnASxpo1P3dskbVhtz6vI99lJKoQ3c7VxKceq1CTRKs
Zojy43LPehgbEVn/5+SYvs0bmdcP484QSZoy5NoOho2g12E7aMIIRdt4YMYQYUAcvCial3psKbwC
nNYe77q+afvIjbMn7IoAvKvqusU989fZR5NaOt2QUlPdtQtsVFkHvJgKZGxsG8H1WSyt1I72JcWc
F8mvI9hSKNcQ83JZC5GiRL1WAVKd5IV9UecTy2UM9HYXGVxFrWc0h/0wLfWocOpX5v/87FPjgLkr
KTv0rAmOyviVZN+Qw1iH4zTnPCakzdSHxyE3s+LRliHgsbrr6FkRq9mAyv4SGb3ri2SUh4fhtW6l
R7lRSA9+q9Yw1/uKwIokZedaNLTdfP97SNu5NWNzVuZgjEkErQaMChimLrWDkem6lJ+0QSblmvgP
ERtYndjBURsZKFnecR+z+dxF4esqeG3T2dyXujjAaurMTulOlLyUdB6nlRr2Xw9F+0w4a9IdbK/Z
G3BCCjMe2g8sZhaXVGqCFec+H+DFsdbvuuWmz5oFU+5wt6kYEtHGgxF4r7his/i/5jdmEWLkLxyd
O4WlP28NDhXWa8+5H9qay/nhdQbXY+FjupH3YiEvBttsIFzbLbs2RWn76NJ25pkhrqAf85C/Jvlw
nodKsY4zz9woK7MOJZG9EU0kuqDJq4Ojbgv7XUyhpBm9/P6ItqTUEolYIiazcGvxvlIupLZnEcnQ
uNCKwMCs4stErfFoEdf8SxY4RQBI6RksROdoxH4MJAJ2bekVASGHrmu2wTsSEQaJkNSEBVfP6tBg
w7sFXnyITRigp2FOvLoMyQ5C9RN61oXeGe8DTI5jhiUoKGoPuOaPb0UOclEQK0c/MbpJODYg+aMD
eDWN4nueLcdK2btvkdBYh+A6g8giulLFmHm0A7W/fYaSIgC7w6fY++zZrStmxyREcuiIM0kFT/NB
cQjQV1HUBbIHzZKsZkMG2UNYYoaJxHulm+EmyTFNY70iiwOSd1aOEEl8SfeysY6fM1iP/uWxX0jR
6cCK7TtWt1dJ1X8+a/H2mXYNdpVkGxPpOL8dqhnFEKTEGGc5cSIP0UWhvr+TrvRJ1pbtul2O4qur
cEZXADkjqoj/Q6+ZsHYKJxi3BQi4YTjA2BQDo+zQOkgpQBNtnk6Aq8+86VPU6Lvlys2FIeuedfjt
w8CB4rbgGqY1mA9fVb4YXIzMPnA7y3KyXFfBmRpm6isSx8wKsStCGkeOZqDGC0dWPcqrlheaKdv/
r6gvbuDEPpjQPciborZMWqSTs/tmq6Leg+HjgGEFXgYW/PXxw+NAFPhS22L8L0p3H2oJkTIoGeaJ
0eszfBPt3SZesBrHluTnnHjDvHY2XmGICqP+A5RyCRULs9MZoU6BztvTEn5b+ejBldUBO4DA3DYK
XQ9us9GM0x/L3dAeUbQaF8l9iTbH27lVkTZBz/twkFQrhqMOYvdWKO2IwhL8rCFk68W9Zsj0br7M
XVl4PJ4FGlxJ5AM8mBjfSvqFIQ98947rrW6PPCNY7+hy2PDry4EuLE3n5s9R9p1lLahzVloHLS70
2ebhSlskEOuB99pk2FvnBhlzHt3fl7V0cDZl0EqOoAtlE6Vg8I4RbY1bl9v9h76CKdlt8oooCXxv
vHLbko7iiAYlwKs+XEMdMLEqZqVfI6sNvx4vnZogqsPBsNCFHtuv7FqEkKxwwKjWqV0f7yr0hDNS
rP6IG0y/Ca+arQ14TYmRWKWXQuhVrcoHVc9ih8fksDhb9xF1LGPO2M5QcPoWctsXqiyCsosC7EDp
PW7IHPAEV9a0w5c12bGEom6d6c8WynGvwdU1CM/Q7wzGuT3zgTva3ezO57qDlLGxmwXnUgMdgvua
oqyVVOPUboJDoIgmoqv2ckKNhROKD2/5pZf0USO671TNvmNDI6t/DjlzwRyFu8Tf7PKNO2FEBzCF
8jj3VqmIeNbPoKwB+9sD02y9O21s/9sMhzUYNGWouxnXOv7gZxfC15oq//fUbo9UAZFghxjiG/4i
sEU/nVeG2yH8mCK43uMhaKgzYqbWQbMTrr9QIm/M9bN7OSOzIJRQZ+fo1Lwpjic9/YM7zHKfTfVN
JkTH3KMfMK1xAjVC7FAQoP0ab1ltuXfJ76rzxJ6jfA98/Hzl9PDJtSmmeXeJ4JXgJwE5j7xoNdb8
iLjELZr73VRpC7NiUQ1sTK1asTzOKHCfRooAUIM7Bq4OBWlsJwU1OX7X/ZOoFCND5QLMY9mBZK0i
xFy17uCOE3zFtOB5KfW+De19OuiActNUK9Ngjjj8PO44xpfaxuEAJ/fTjpL2Q3I336E/aXIzYWss
Wt8cdQbp1pmpXe/JTVrPLB2ZrxXLAtF5lS+QDtI2SJQHckhdNDdzPExICg36KXtch8wfmh7h6b8w
g3LtNmCRwjWBdifl7tR8W4nRkppXojc5DxZkiBgSGuh9CxyAuj1C7luf0Q3jixLvxei2JfhrC0+1
HCLe+YDS4jovCuGRRA0yapoqdibjtW1+0qf876vM5Agfivc+SPauQEI5IQgR19DQqBz54cau1e19
TnUhY0FJjqK0zDlTRDxLR1Jqkh4UMemzYIKieopS864YbpsGOtXzjy1gODpG5088XNO9uBzJA5B7
lEYxy6LEWm5QQTuzQrzxIlZe8WXwL928BL7J3eS7mx3uODtIqD/7udrMgT9G8HQhIN+V8itAVE/9
CKYhNYPVx/lP45kCenAP1HgHg5EBNTlBcigXzDonC1Imx11/QfwxD2jTbRzV7CudXoJehOlp46w8
YVWsEHMmRmU2jcA7SsKC+WpbOoUUwj58D2cSrr0xfJE4LmYk3Hs6Or/mcKqlV9/IVRYuDHrVauXX
1KmYi5TUmzVBgvgBPkee7vR0wTjbeCzU769MDFBObYsyuCTNCFsVtwcJlS7OT1ff1/foRWKDxD9f
DKHtNdFxai01fEVYhRrSM7VicbTiukFzVad4iga+9D6M/09MOlrpGMWvTI2eEJNhTgruPpmRGqkp
3oe0Dy0gVQGRI9pKbdeRwoedzwX+UVVKF4fR85IynPiPI7K3ircvobCPQ6q9qSlkQt/cjxLzPdOK
vTbevByjVvg4zwfapvmRg4CepHYFT5LLztC70s3zkmm8iWpjo/777RkMyDRnBKZG+cgLGzzLsK2j
zrZJh3yvDtJACnYkIpwjyHdN7Y+Cp6srjIjIcOuz3HNFbkDqTAO6v9S2eyTh7QUleSrgsf9Z/yy4
Jzab20+Wg+Lev0FnWZDE/x+hCzvrFveD5OfwR1tW+O5/lZ0nKN8s1wnlR4M3aNNoen9jhsphEpvI
5VHBg78168C2HuMcqd5re8dQUsOoO8SnFNXONYv+NtBAVGIfJRIFgqxnq0l9kgiSm1X8ggCC4GsE
7pMKMg+J2nLvbXVSzcsJUCpQPAtYsrrD1YEV9cb3topbTPT+B28Qv/NysvGn+YYYIPJXLfm9Hi92
23e+1x8Kaxe8IK85ndXOLhn4nmZL+ath4xsvl/SOECwODIAC/Vbgl/e5rlvpK+7b3qwyp7kPBN6G
A1h5/CJ3E1A+GmjTs97CC/AhRVUdFffUF0CrQ4tmIIipnb+VYFVEx4GLnHuxXkgSkg1xMQoLdeJc
pVBWukN67nbZ/43n9+Cxutai4uy17cMYMswGgYw8++lhvSVh0b9or5N3bKe17N4VY6eCdt55Lx2a
V0T2Y0mDyfn7C4WiqqnGuU6JJpNXfgTlsiNCUp9NVg3RhySeP4c3fFdHcMAYqJ6MZcNEceVwL8aZ
kKY836Zx6lhOzTtCOboY9jZVh7LAbmiKJ2xT8RjPf3+M6GFmR5pbLFgY4csQi0j05Rw7WzNa1hYT
0htdsqT0ExZCxZbeD+wkljkefYBAHTkquFQjwbLW/MQ+K4VB7SlKmr4pT/oThqSr16WnOVS0Qywe
+f92BeS/1mO/PKdRTnEWFi6MxryFyin8MuMKPONRzViQvzwKpBL2Ur62CZO5I3JCM4LJv71Two8n
qwTR2sjiwbbuHslLTD6qyyLQythEJ+ve8cJnEBUbCDo979NuoFAEW3jAaPlKwtVtQlP2vTYDQ6no
KoRDk/e08ctqTLSlMOxnJdhnZklvO+m33ZuBRhHZ/IWxjlezEvewyvNW/jef1G0oQJRiq0OthruO
Md86U0A8BSOpkxN1UL+L87+GBlWhZ7YQhp3hyof14ovQS1tQO3uDRh3kwOP8aVwtlQ06R3L43DGI
TV9lzJmzlggXlr9PvPzI2bNeugW9OSMNZPgCXQgFuicvJ1CuBd6U9OF9J09jSieNzg6Mx6BAnhlI
GoYK5Gbj32oNYTVk6zkUeb6LWnFtEpWD6SQQdSDQK3P9khH97p8amb2Hy4T3uel3kduHTTYa4qlh
P3J9rBfAE4MNeAFOnPpxh5evuXS0VuX/NqZFaV9Vj3uBIqnmr1mgte4PI14vLNMdDK4MBfLqNDtp
MW7Ll/lQqC6Dml0r/VKGhD0nP9uoYD6qGOMypzMTV2mxl44lq6K3Mt/OLAwWRldvrgm0IKKDF8sM
HHVv03/txbSrhes3apC4q3YLoaiU/e444Ez5RX2ufQKJDMsPEo+JrN91oDiACCYXzyDIkTYdtrXi
fYUTUrXDGlYAqx22O0uVYKIOlCXDh++ffva3/YdEEKF4WL3gqr6FhlStBIFaaAVq/r1YFixxqPYs
hcfYbWvzMkd9RBokMekjLUbaJAeIpgSlHuXMfUesNW7/vadQDxQLnYRQHldEGBIbRX3T4cd8h3C/
uSqSj01NJzRHhDui5+kCDuakc5ZKtJH2ECN8zhZ8JyBYDDSrKlz+diorcvPhz1Ux46E3htfqsXqL
m3sABgUKG3H4Zkr5FB/UgsXsO0UP8qe3SbgMGjGNhCuBONvt+TR5iENNSv/LZLnl4sn5a3cWibXy
nK710SSyeWmbMp96KAhOmboqdcH8xAzya2ikCzmp24dna9eWM2p62jPDBOCrlN7GsODo3yL2Dr5/
jCCloB+FoAuwoy8Q4J7u4oGOW+8URX5DVyie7cliDjZvPz396XTQYiokP+3Cx0buwY7U42T/VGjU
vRqyis/RIgG8QBGy4eKo4j4ujMgjx42r3/IRptv7ddI9nvIfvTvC4RGYTtDMudCkY9gjpGDfF1js
N2RL+h2ogDoxb/FNc2PVsmvnW/K3o82wsEIY0VbFuh5zrgEkJ5i6vZasarTAzcQf1wRjC0xs/nZs
DcI9cFXmE5J/wiAlPbwneMWGrUncdWYQlRJZ2+/pnRKC22y+ysOfMVTQjVRizn/mnNCJBn7/ANQE
fVUjhm0KQQ0+UN5MsIEoItLoL9ZQY0WvJU34uo3OnoArZC5G4rI2eA/GrrissiLRBUdpjIl581e/
PPrBjWvAA3FFjPkA/wYos7cSGoiCbFC/doxgzuNvQufjv6rKsHoukmoSOjcKwYQbCrUw7Fx6gKTg
DEbHZT4knjZuURgDtYb72KhwWWGhGq7UjfhCF1No8OvRX848DwUEUFK2QN6A78HMHQ1WO5ImqkG3
s0+8bxTgS907V/27Qg1iNa19RQtfLUWy7VSKyX000cGngt3+Kb+xlnI1OpDhzhioTxtJqtVfc+Hj
sngGza7MDaDWB+7JB5lCiyJs9aPUdtLsXO4xTGX6xZAEyIxNwCGWrMoxfkG3j9gtAXScXjBF+qgf
kZA8UhkpfRjzamUAodUV+ZTqJTB630myHxTOmIepB0cJnkca6EBsBi7vkStuWRAzRSCQ348A0D5J
3HXrrinNkPsESd3bQHe4IWDlaBLMk6zCeLRPqO4nKdTDJcF6DzFgRenaXmx94Ga4pH5x5z+2WfbS
s9WE1m+xorc+N48+GaHcCEkKp1B3o8tjc/o2xrRDMfWJb+n7YcXEkT/jbn1WrezX1HWpvNqckirN
wtK0EnHFHo18VNdP+YwGF77cCtu6hfPMyy9bAW8CVrUSSGfmXlONYVGXdps9zGhwqR3FLHet53Gs
NiRjqBJrWnOlYJRKRwf7qll7GS4BuZGe8LODe2MFV4ro/sLLrvwRRHkwC0nVAAyPA1bVojHRUPzH
X2Z7hMmHmrt3zbQObPnYWKMlb5ia3hsmD6UiERaf0FFEzih30w6pOq3jIlbeL3217DSpqda/Bmzv
0T8kU6iW1gk0aOtRKPyjDerfD/biUV5W9HUGEFJDUq9q3XUc84gDr6ve75WqyEPgRANA7wJrS40R
H07x+n69rNcWo4ipSu932xOv+Ghm/Q+eqqyU8su+3tIuh8SIkvRg65Eo9o0XT71K5oeS6dtPUAyM
0RoUVftViG1QRz6I/l5JjlY4dLPLbRCt+0lVdcuTa4OaDKzIz0YcmrA2ynVbP6c2JyAaiLL6R5M3
C/lTwbxlD6tb/n6tBXtkJrfCQ8LrHvx/Sgq7lX4Y+ap9MaGsl6F+WOXMVQv1jlPSSiJrhQk4DD88
2kXMvro3xgZabi9iNAhvOjOZxq8UY2IQ3jVrR+/RRzv6rHoKHanmHKZtj7MXVPx+YVizEg8K3IoM
jCkUgpul/3Lqz4YZQjJbRMp6V5zXV1oIy1tFl9k0JNe9uiLU3dHcOoCLHEQbTIkGPm5x1774mm8C
9TUhQQOqCGrEwCoQlCFqwQVXTOpUIeikS0VK2pSZMhwrjbxC9X/jxlbBgE2hBLhPg8MNeakh2eX3
91XZmFwYC0hP84NsaZIPDFvaLBUiaWcJfT2NclTKcuGlEGVt1PzNVRnux1wiodnyPDPSgGIgRQuY
WPUsa6kOWVH+BxAqcqalcDP2o5dBdWpeDAaDZ1U9ifH7IzjcuLUy3fiAYZ+RhMrq7AekdqQhdSkM
a++6BKah7jqdH+Yr/rt525idVPl8ZhwrVL8U7hhXWUODljqQ0SBfy8RExw4CudKID2iS5hn8lcmN
V9pKu5K8npoklAhUimYx3/AHU1GsndDs4GqeKTQOxL6SMVifYRXkGdm/EG8qmzl9Bw2KDB3fwqHQ
YfrDaFRwN3CaF6KHd/47HefuDbjCi/Hng5V4HC+4tGf808QgQCPkT55zM0aFQYDMKqdWGTxah18U
MdleK86+bupk4kkmo9tKDH5V9BjawdREuzILif6kZ0+4q5yRwg1IbDO9rDqcRIqTsf2CBFpohjb1
qikBvJggLHAc3QTcQAPs5QnZDBlzpFDvLlkQx+j9tO+4aqsPT3LGPet9+nG1EiGqQ9MPsyXdwvEY
5wUL6eXKXuDJ3hy7jtjPmasAXHymFqWAdwimLlYODJFHjp+ZCoaD078VEtiCnjuHGmAuwFoQERoA
7mDG2osbzyFPjPutgTW8vJIGrtfOOkopTnhX2jd+ahk71NR/x0dSZZHnjwZ3VZ2dHcFN1b0nei1+
fga+qEq0P+hdZ2yU5vpyz9SQ6k28SirU8n2/gat1WlnTu2PL+yWgAVufEFmXQh5AI084GAFji/8G
dxf0fkWnluZoLFLWqNChxcDgXTYNjsfFDAglrWfP3gEEwa6DTYZ134N18Y1M3RVtM9Sf54svbn0n
WU0BOcBv2dSprJBjBIQDM+b+/6y7SpicuvxMpHhFggN7voi5AAN+B3tpaArL3N2Y9sQEBJMdf1mU
uPTw8MLu4TWkpqHMRBHlV1LjFgHAC0gZsoQHXFuJSmbrP9lMuHk6QZqTowv4Hcr/26WOd5sP5qcZ
mtO3jAlHe5lFAclNf2ZrIRezwp1ltI5kkXydbPIhbwaVN4uTgOspkBUa//dVR9D/4HEvOb5x5drL
lGcfQndhbHgIFjaDv0ra/rdsbQ6yfo4Nqpt7eDEAS5RUW8xeWxmQ7nR/DopDRs4Xem7pEnW9TOxK
P9fsFLS7fvUpIvW8fYQTLtNKQSR2MQHdRQjBs4lgFAWjo03aYVChQqKgwuLMzFJTDfIHMq7G6sL9
P63uddNjxsCnL4j17FQI66WbnMINxl4hc9RVEaD5DyV+/jkERz4i5TULwANsZZTq8IBZ2Mq6VNFB
f27pQ0/AZX/peLkEANG2YycwmBuvR9dCzGO1pJkxAdt+VkT8oDsLZTftff40kQ4dpxXSG6tbM0oY
7e1l8W78AwSmuuFkASmyvyG4s3TpdKX51GlCTidGnn12lyqRGyddngW0a4HeqX1DYq5bS0ynmGY/
KPcj9M42mzXAdulPIf7DfAz5Jt/0q8XASjUvHmmZISSsLLw6HzYUlDNk7sNqUX1Fsne/2cmfEdG5
QumAgc9GuGDF+X2CfV6toCLljSGiHenAFU9cn4jiGMRw0N7uATRFrBCYymh3CDKQAQ+PTtRTha5m
t9hjfFWzVj/fqmYEV32suGW5MVsD63iDit93g0qTZD5N/718cwxPGrhvMdXumS+G3psmlF4zuaeK
jpN+i3hhOsmHplLywph/bDqG5IpQpCpM4JbwC27dPH5T8lKBOnFW3tnODMCpxHL3UcIEYOSz7U8K
jPohD9Iv+el8nVRg4nG2EDskZr5rFa2HE25cJ8SBHyiYu8NkVk4LTzi9U8ph8SpMFYocOeGrA7K6
pWMcXfpLJPOwAGKKgPILxy+O/qtbRaGNIcvEqbo/OLWF3/PYidnaktkmLHYh674PAyYtK3C1e7pB
NAt/yhe6rdt5MBIsJYNanr0LwPudsHijwMEIqzj6i8407mElb97AruOdBHcdSC9Z/hLGvnTW4/86
7uZWHHk84G8Qakyf3E9WaYvSr0/+MewWQnsDzbZTO2a5wuwhtIg9u6Zgj9qHmwo5L0yZnLPGkWOY
3nXHIJk4Rq2uGOXhu8IAKJwrec0PZfYFg3ZQfrMfvsz/albJD9OJSEZoCjYS/eRqwe2SWZOwus76
rge4DwYLr5dolRiaEGfxw5R8xPlcu86biRC59KAxIP2Yf2WYJ8xYyyJVFulg5a9zvU32q0tQodyu
x1agIs4BQak72beAD82+cKix+qZ6x5zknH/a2xW4fGJxgxrRSV6kKHwykvbgsf9/h36hp0tmW5lL
vX2UhO1DuLa+wjB7QYmhk9gEyjsTuNkoj5Y6HI3OY8ZKswQSEt6pEZNFQQYLw5rRJ9UqqEAuun62
2q8iOeBnFVhTc2T2BQuPh6GWMEnW4M1yJTWCJolidaSxCgc+7hhVKD6ZdHhojppPTzI7TzVYz3H2
7d9aSbTVVQKJ1Q2A94/VSTtbFHgw+hLE5tCTis5oqcnr0Ql+7TECTZ2mDhT2a3Qmm+3mTwctXJPR
wZLVkybJtR5yYyxjRvaMXiP+hxo3ktJAnd3C6RgoiE8M6ybTz4E/ZhZJidROp6DKUz8q4rhNkXJr
QfFwDVD5sh500jpkO/3FkSjS0Qtekp04ZedoyLDrBIHWLtU0K/AVxCSoWmqS/coUek4DE8UizVMc
/xWJrTOfftJpbKXMIiZUwJfegrd0uus1R6PIws0rLMhQo7ao1v4T8onQt26E3vSKCOG6YkKpQLjD
DbEJ8OY9A3Pu7cK57oJnKWd5I513M2DpTpSvgfBDhY+sukUVlpC11MSpFeSSgdbU5qgYnfYbChIj
o1a/4wMDjmuruccpjRvyBFJ5h38249gBgFbEi5QBHZd5KqwBHdOq/gYQ/v1G61bzSD0kOUG33bFu
6AxtV6ezV8ZSDeUEhYdDDhyvxl/vO91nrUDpSRWUq717xsYcDimefmU+Mzledhm2uLQzd3MaV7/a
aqnlhrFiTNOFUnmJMsts+KswzM+68DoiF0UfEfIieAwEdjFpFgPSJURk2x/+ZvdpuwXEs2up2a9C
eo4WHI7LDYBPnZ5rGdcKAGwSJmcj2cYfJeqQUNfWtrcRpGuBAp+swPlabsJd3xy/P3vjsgjrHEMM
F7CjEvDzpfd52pSMSE8m1znmpY69zsk/YBUSyrwXZ44Eh+5ukP7HYSsE//8l2fmYSfgX0p+NDfxd
NGhKfoIJVOIiawQuXI/wK/cfWzq6186iW5bCW8ElGDlsvWyocUv+VsAWD8EWsz27rQGSJIVMTc4X
hqGKPrmwwK1bmv9SGZCB7LxIZAruVu8GKWhWfOewlDQuJVlh4plsyf3krBDPTJLTz0fhuFAxdap0
YUZ/PLeQQyIvaRsO5+2H/9FdCtwdtN3zt8CCHAAom4SKwZrkIocgV4k0zNL+8VZDxc99HuxRsf+f
IJrOw3glRNR9RIJR0ztCBbaUggqPyWzm5UlMH0tuWcaBlaai4vTWcP03NK5/FvJ7WqMnesUFY+WN
tfaVqtL+SgvtL+47l0M8yg/D09aFQooOPJkLCPyzZc8zyt89TZID+ejQrhLho1w2OMqc9cZDDXuc
Uz/KlpQKCa3dxlsNEDrITRU3FgNvzUqZc9L5bEMpfnUvtnhZ5uj1huAo27AYoTpeTXPkjV+k994Z
0hqR7JhVUEbkzW52Sa+xjCTgK2mkQ2QB72F4s+TaEwqlCI5A/y19xsDNW8OzxM1N1LFJdQAgIZhN
tJm/VX5d8Hx2bsG7ph4ujGZscZmb49P20AqRouKNqhxnJWqE/K5Jtf09xax1HU/zb7jKGpwRMtyY
6yAbNkI6ZE7jPcWxvlHSzrYmnKdH+W75fZOe8MD6pwGQztQymOK9dLyV/MDfMsB7vBAffBUKiRb3
PQ9dU8HKtLGkbqkgO0n08A/n9YJmyREx3V8HZkT5VJlkXyOSRDnyS7PdyI9l9yT60Yzx0R11n6MD
L5tVmKOlQ2t2KVn3W4vde0cE423D02TcevGqZ/Xh6hYWfKhkLnWa6Frcn9Gw2582HXoO58bcKrEq
QQLDm71Qb3nLfmxyWnBR4aBeSf+G1Q2PcFpyjsolhfXoCfc7MU+bX9ZWvxqYQGAyRLqanZGhCs2s
GLZ0hoxNmRIHoqMMnJnAm32MJx9rFTfYKBVlaBR43C4DTFlqoe+WqL03Mut1AF1bn7Clt0PhwLtU
NokZqJwO3MrSHGh7/lHlrHnafKgrVBp/XlIYp2ow+cJBUOcjZ1hKnp5bWajZd43k+YHIboMQpgYg
7ZSRYLMgjffm8nu5Rt9+kfMBQUqrBew2GuezK1g+Hc9Nst2R1OxfOF8OsZ/1hvo+Yf8QI4zwOOMP
w8AzqjkMcnmxHTYHuOtVoC0cgrQI/CsQ7HSJb6xoHqONVg3n7MZ+LHcqLX2z3NV/GQ2GQ9Kfz4r2
QPAk3atP0RmkSGZKV+KElMEejrZBPttsl8oj+OVy7bPi+RfIl3l8KCc+Y3y1b/tCNE/EC/ayiccq
7Ziy7x9w1bhCeK1XNjxGq36ejxmB8H0xXyf6rYviztj93W4bMwJClNnYEnWS/gzA6sGyeUKXvasU
H4TA0zp4RGrjExCccmIxOkKtqoACVIAxFmAjDPpmXeckDh4VlqkZLWKV0BMN6ddGTwLDG6eZvXpy
yK8Or9sJlzR8X06X2RIC17F/InrzU/WNp7aPjxDpsZlZIZhPrk6lN5OfkitKBRd5a1PUBuHvO0Jz
ZOC7tBUpHabchSfkn97xtnDkna8TE91A0LyRaO0SKAdQAgCM+Xj5a3lBUVyQr9ojZ+LSDhLctCo/
zQXR+VZU0bIYh+7q4J/MsJQXooZ1/glQltoojTFUIFWS+al+HARbkNl2/DUEsrbvleOXIdWH3TRp
P1HLv21fX/liSKQQokGLr0/siNMmSt7eWj8j9vIojVl1dUBlghg2bisEw7iKXeTBGY+I2F2+a3hV
rQ4/guYPhROdlVPAwCauuZv5xhpXWg51U2dZ0NWCRvZPSDV9RAY4cVNr0kITdFbLZoRAf3dXmERm
A6/Yj47E7tcaarlC5pokEsYnTLN0bky49ulA73tcJGxT+9BNqyV7Xa2iXLCc6cqT3SYwAQpiA+5O
kTxoa5q+jEnxi9x70uZ2gPrWpxh3BlBZauVtiwtnJ5FdTrgzbZj3dflmhHC1pByrEPp71P2z2/tq
x8DmEXPl4u031/QYYmdpZzLTCrQhAYLaApXkENaXObzgyrcw/DUAeaK/WNQCk+XxUK/1d0eY5Vpc
PMpHU6QhV9qhgWlHUbYoIZQCBiJrallMdu2OoQylfNbBglWYUJiLrgGryCfPKPPgEnVEUHcZHiPp
fYm/d3mfa63KfTeGjDsz3ArB4B0M8WQ2IlR3kY3NTNfqeA9zORc2pOdSx7vbvyRjwWm9cZoDSwTb
sDSzKwuTIr7mMpQYDhJItkwsaLFAu442mEfGpAskZXbWTR+/ZrS7137kqM6DTvGDfgHSC4RleNAE
xm7lqVcOSEw9Gekkuweg+XKpMFIGyVhRq5t1oIa2J6JuQEGgvSIwcfC7Zn+7Q2O3uLRxJRpEge3w
x3l6rCX4BqXvPO5Jr9a2O323P3e+z+AB1zskfoYv5DtHlFmeguIUsv8GVUra/caeyFei+F0No+YH
4vVdankO1aE/LvG/SnnxmBt22T6cAKBEsJp1yiMCTI6b2XKFfSxSzeHGEQ00rqKkte6+TvV3AQ7p
LRsgncAls5+8iZuJ5/oBwOcY77AtOLn5EvqjKhWT3B+NI8kfGtRZfOz2875VSaCq4dRihXxrVHgJ
anPydz8VfJbToYwF8VByORau1zgpKjlMVvpXJYy7g/7r97taK0634+QyK7/D7XfLstPMbIZHDZTt
JL5eOABxkfciiuDSPO+Yqrpco067ns6f/F+qxfGf3MCU1IYy1gu0UHp4Ozj6UMBbhBpRnnTZ/tgM
m0SZUHKivggFdP4AmhsYEqArvSOjQMRhcf7+opZGP47dSVbyARLgP6b36klSMs9MHiYQWf/7qIc4
9SNA5oCVY8CGgqRAsKUM9hHIwSKiVTHQhZk166qT2nsXjobZAIRMT9ftgUE4M62owZgQfIM6AHxs
hunYdzSwtl9gEo3XWPZOkSwubC3BYuhNKQJFb4wB1XzrIYiy8C/YT4u1azG0xM/p1K0KEizHO3jm
d6TqcL7tUrszzjJ1fqsaAQZaZVZqea7L+JQWQ/Rmqm83S/si6SsE0O2lI7er6AfTZInFb0QUpden
6bWzqiivpRrPt0NCJw6dHllI0B5GCDhpHGRJalQGKl11Uv40Ji+br501k8Szg1np75WC5S9Q7+e0
ivfh
`pragma protect end_protected

// 
