/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Fgcvq9yodAEyu7zsWWZ7LwHLqer2uRdIROgj+b6me/wmyj6mu+r4+a1EPBMoGlf2Rxb0wqrGm/yl
7FT0a+0gf6RIUa901Ug60cEq5l3MsNjnNX0EuQ9QHnbWnPHO5sk3W38XYr3s1DoIymcMyzWSb3j7
DAgt+R0iGXGbLJHe2UuAgwrybNhjpWacbybFOYZoLu5Z50wmOHt3p6J+gVbTwfuHK/f+KnS4VtSD
EJxx9+hQNEvkukNe5IcvkATvsJ495o97/SdF6+o/UvTHUZ0m3la3MPtrbbqjxbRc5d/SBaUYwJ/0
DSKgI3IBXs0nO4MGwCQX4Cy0xa1KtNy17Uqy4A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="YyF30NSJW4xBU1bz6CmJ7uDDg1utz4oEiyNQAWYk7H4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1568)
`pragma protect data_block
3JkMrY1IEAXvStruy6C+3vLUqgRo5Z7trVAgEQIgtyjcmm+S4KTCQH9RJZpn8RnZZTW8Hh5Jx4NF
O+P5uEGGmEuw+kJa6VSA+hYK8cc+x6Ojf5lARRK7buCwqaffR5Yjhk+ZRRknNhQZZb2QmG6FX5Em
rBCUgPnRiNsFECrnHMl0njdtrPd+ZfEinxVv6BbO/phr6W8w4C/6hPYCZMn8iZWh0XolimDxELdR
itucT4Mmw8XsRO0SoJnlLFzWYTZ10PRBWUTjVl+4KqcLJV3EWvvHuINpAsKS+HwUpnDbGHPOMmTs
hnCjEjjYzBZvu0I9VOmpZmSyt1SqBQOFpUfyoOxXetZucMwyAw8hhpVOUrB06CbrLn3ajetfcWNf
kupbMOnPLXcimTzyaSBoCf6IxAywFmxtrn6iGMbDVo6xcAdW9DxX9YVykLNzGbxm56DNNsxTLchu
vmoMTbExPXL9yVtxH8V2DOTLtAVbFQwmMJcOyGQc0xOVz1Q32tYk/OKtRnE7T9KHNa1LT40qLiPo
Te2lfbyNR+DfeftQl4pNLAKgpAdoHlWf65337fZzVAYY+EzhT7Ce7tgc5rthdmR85QAQRhZR+Hnz
5vH30kZwQ0yynWLEBgYLP4J0M/Ayu/ZLBy9p1G5is+V1tRc6zYXC9DVvv69lK2PVH09tGrIkhVSi
yBzCgJEdcRmZSxXh0seqJ+4EVGn4cF5Y0HZVqbbIx6NccddzwnBDJIwbOGVtxjh6CIDcMYQSVWhY
g+cEMEL82Ezdw0PRzwUbqUJCJXAjTEwdXIH6cvkwyu2Jt3vvaRRlhW+9Mnkv3+d7ACDRsceOeGGh
v+KvE2LZ/TjZ3MB2CNvr5eHy+h/J5BHXqR6qccs3m61B3BkDERNob77/U1ojk436UVAB5zq8lCZ6
UUh64l6dGIQJqoCHPLnI9CpC2uqMlwG1lV9IJLxgzKdWlYjhTj0jfm2DnZ3JCZ4LcX9ZTnfNXKMS
QHNzYJDKQHiaGSXJhtKqCq14HN1oyea+b08pBB0amvfPGWD10HrldNAblgSWH7sqcESF20tE7cp7
k36fH+Am+uAxnMYbhZty9DLaNKviHtgZRELz9Mj8AK9ZC2MRI70ffwNTU2BvtScoElqh7AU5XVz3
P8EoWO+Xac/5NoOcbnVn8QFYKUK0ndOnpvIN2go6a5HAnc6+MIw53F5sv9OPOaBbvn3VvfGGVwh+
YM/5PKErKQAUzC6E9b6/oJ5LfwHUL/dTza7ZZz9DZllKM317w95NCtFzVJTB09SGWIklC9OTBQF6
WsT3ey3M1gmee5cyntxeQCj9QtpvjFuoV1Ti8yS8TzA2n2ur74TmvYWbJv5QKM5qdh+l34CBCxCX
NEpWN4KRmDjQ1naUx0rDZp2lPhYToINRYBYbXqYlncSJyTcdproz5k1B68r7CTfjNpb62/3g1jGv
QIhRFF/35HLl2ii5/CvXYu8vdjl+/5zuahk6M7/l5TsFJjLoJq3j61ZBZkZWJssBJaaD8sY9EOeu
eT7YmrRPHtmBO/UcDsyIa3dr72OwXkjWHWxkp79QSH8ECRic2vks7oDepvsrGUJKj0hIn1BImgDn
Ybyr+5syTIE6g9qeBzc3mwlJ//VsC7TwYRHj4KRcUz4KybvpKclPpmrDAiTk7+8u+rodKdoqgDRd
toa+O4V9hIhYy5jjHz60tt3pxdMxlHLFl7E6pAJeq/fguByNOzdfb5W0vWC2vYBxM5ia4V2/LOtd
41aQyv80DDzwvwm3Rk12JFafcsOYFhfDNniov+thzu058t/XbYQTljtDcF058O/EEZpaZ333HLif
5dNNvSidJ4ERJ6DrIGEe79injgMCI0elH33/NeWBdvrEibao1AiSzZDlkvnKyYq73Ma4F9gOoJx4
7ob5cEgr6atgHrApzCvWtsAYw//MypudHd9GJsIV/Wzdbxe8cqp0VDTQZJ1qVMOpBn9vGjjSpe6G
72EowUYaXc5aq0qOR0ficwiLEAVdL0TnX4Xck1lelt84WiMycz0lzN8Tr6GmTyjRhlxDc8ec2l3M
+33MoRrFtIpEqH8o0TbXTMbfUKGDiuVViI3OQiY=
`pragma protect end_protected

// 
