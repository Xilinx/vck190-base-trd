/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
l4gSYexUXlM7ifAaBP6t2MLRFhQaRe7Sma+zo2L28DiA8DDFN158h0/DaBr1OsRaQKqTpiBWurc1
Kc+8TD5uaOBbdGAOqQnBtAA+GhRIwIir9IbLuxBMnT/JmOaK4MUYPqvoRzrgYyXFE5yrJmMkU220
b8Arh6+dyt3Bh0bC5r9kA89v3D+ja9uQnY/8oodAq0Q20j5GmOBNL7A1mEvLof/A0UYhDRCv3pRO
FKF8KrYOR3RN8PBeGCM1EFnr+wW3J99nOfKe+v5+if1arByO/0BxWK1JYTBdcxntFYOrk/8juzWe
cyuQA25yLLNZSsEfw7pTdA4YqggvIwnYX+4CfA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="nooMg7GjkDsMTPG3DLODBuXednbZgjpzUjgowzton6E="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1264)
`pragma protect data_block
OIw4y6hn7TeoR9JbrM9EZKKXH6OR/cL0wYqU9/+OzZSas+M1P9s0Vwo1ZdaoVsZuUBR6fAl6u5CV
PYDcwZJlyZen5Zan9VWIsoY4oZsb4p2DekJskLPKZaJ7I5ep9Xwj8J+nXRKG7PIiYFBhLbbAEqjq
J692CXdn53/agB5BYYk8n8705EPEdsj5u12MLKWZhwnFByMu+asRVwaPdXW8hIRAVJpO+HPRuFkL
Wyj3Ur8k0RmG3vl3I8b9+aeaFDrMqLCu8lU7BKuW0IZ2NEuufGfSTDvQ9XsMMB7/aIdIfJYiXxSD
FwrTutKL4GJYI30u8Y8XI1JrpK45JfExStyODGpKg/32DeKtSy3J/0vOTEh/n2Emn2fxLqqDBzyk
hsPjPLAskXcCy2jt5Gzmsm0+KvsALYb0GCd/ByziEamxgvj2Jy1fo2dx7dTBgsDrd4QTE6MdVH0z
TXUvtRwgm8KOMxUsxG2wYAfSWNBu36LUPIUWbDCG743TvcBHLjG0S9OTF6/k/Xo0lac3H2V4Q6Ud
OtJmEXWdwhHCDzZJkROoQkWYjCQ6Tuist4LZEeGEPonDtif9WvpeGAIUeoGhS3UNi/5kbTOCp2YH
ZfejTzxGbelzhU7T81mpi3lX3pSul6dggq1/J9wPi03wQMHYvzjjzXppDxJ5pOvhBsYBJQVRUA3y
r7W07Pw3ISZuLIEQ3OlbNJrFYQrd+KQEJjXvRa5L9wZ3+IRjlZqgjYEyw5KOYU1Mm+ry9oA/R+SE
VNBmcItJqdjbDevLmM0nq8fMYv+aiGvMWW12INSnkQV+NuTyKe1KCAFsyMr2PF2GgYsva7iBvmpF
Q7Q/0RHeGpN0Kqf7kBGBpV/QkQjYyHlSdPZbe5AZUSwiOHx07HoHTAAnf0JtWGR5Ew0zds/2iloU
wjOojpJsPN7F+ANchCCkS41660vHg/08yCQmNmGS2IPjGwZP6YQtw7W0il4VB8tDinDCYQgKhIzF
ep5CAtu4puJZ88Gq5x16+UBamCtWSFAhUGXLbp8HbhpTF4xX0VZNZFB8KJfYIBdQnyzTcK2mqwIh
cd/u0NOVsdcmVDkyZbV8LRraUqat+20pyRCqM7+XrR7pE3eV7an8K307r6B8Ss1exDsD0PneoMm7
7QvL9mvNOQXKFPPrjYxWHrXH4957WQwYsenLLbJncpn/HbQb/jPyLIyO4nPgn1wdr4WQBpr9O0fe
SLkace3h1+GPHp6XworI2xeZy1dbiVaCVS0lUK31vjVpY+dQ1bsfkWCV5rw5t1saBfNIKoesZm0l
EnKhMTxAQQMGCj9WpSXFzxszGCaen/doCVY39LjFOezSTfHJAkCRTxB07qMQvCXFdInmDPm1czQq
mbI30QSltlUPqzd7Yav5CvHt4F0cPe9olJhuKSEmeRPctjOiqHXCqMdd0QXxdfkU0uLPKagx66ll
qs/GzWADRcVnGf8N4GefW2P5FMvlr2RoCsDnqEbmG2nQgziL93g2qQuspAzsHzzPwt7lvi2Sb5sm
g6f+cM4EnIjbWbh8kbCNSf28rO51mGhSbiq0EANiJlq1iS3tdTwEZVgT/hkxAxak6GjPiTg/z/6k
aOIHLlW92WnF/nsWTFF2XiylFYcVdgvpICuJWknFZRUAs0HZxRTOOhVCbBwAkMySzSZW3L81v5ei
Fe1PVMa/UjpC/Q==
`pragma protect end_protected

// 
