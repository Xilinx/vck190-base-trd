/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
l4gSYexUXlM7ifAaBP6t2MLRFhQaRe7Sma+zo2L28DiA8DDFN158h0/DaBr1OsRaQKqTpiBWurc1
Kc+8TD5uaOBbdGAOqQnBtAA+GhRIwIir9IbLuxBMnT/JmOaK4MUYPqvoRzrgYyXFE5yrJmMkU220
b8Arh6+dyt3Bh0bC5r9kA89v3D+ja9uQnY/8oodAq0Q20j5GmOBNL7A1mEvLof/A0UYhDRCv3pRO
FKF8KrYOR3RN8PBeGCM1EFnr+wW3J99nOfKe+v5+if1arByO/0BxWK1JYTBdcxntFYOrk/8juzWe
cyuQA25yLLNZSsEfw7pTdA4YqggvIwnYX+4CfA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="nooMg7GjkDsMTPG3DLODBuXednbZgjpzUjgowzton6E="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1397920)
`pragma protect data_block
OIw4y6hn7TeoR9JbrM9EZAyDfRG/MgbqzhzcuW1rKRzPThlodgOXOzhDXur2X/XwTxNdoEuZdURD
c0Ps5XpOrjc5OloZY5oICOQb+6poURIA4nYZ20aq9GSo+1Ywm/ZQuvkAhcnJFWXbbZFUf7Cg1dGQ
+98H6k99F/OoLOOyJBUEMvxe+5X4+aqjqQP0ZJZ31UnY7s8gEzDgKOFGrLTJpVI/j+FefoGV6W0b
3eFQCMRPUpE+e5DUmh6GsoRA5sWO8sDNNeJBwnYR0X/JNCFEhV6iNTw6/93pCj12lykTGfvsbGcv
XiNt8xDaZ/qmXWscCENhsigrVA5foDCEiR2v7b6tXpelHX4KnibOS6eeL5AVcoRrQyiULlu8lw/q
zTME1iUyRu6A6MMx3DR7pnCww7kF1FgepUNnxFiqMZYiWXQrEn5fwUYltIH2xywJMVGSFU2uCfRj
SB+z/T0onnj8RYeBoKI6j/asfdbLtmQ1BcOWtoaqw9IoC0pnjmJlNX/nHPaJnwyvqx/Unr35nDFD
PXsHoCbm4oN95nqS5jg2Q0S7Tcf9jSIaSirWqBceFEOPOzksLJ53mTT5xZuOaWEELj2DhUpA7zkh
RCY8KUJznw4GBVihzJa9dF0XgVPw5vx2K4Ldrcx5G1NNGMj2a0XSnW/4//pt09hNliO3YH5biSzr
MGkKYvQiQujESaaFS4t45ZyLlNfUoI5EKbyaEyEDRWypcZGhBdmL1SDagiZm1CiSO4tIWNSgzGOe
ysQvXb7AaKE+6PwdPfLCNTx6bMDGxKVpm76ULa3ZRt5EgMCsRP3DJEDh7qt1ZV7a1n54HmdBdJP4
Xbm249TYCxWp56URt+jQ3K/nnmK2NaNMCrAwMmM4FR48mVi8lhfBJVEhvk1etAtAKXx7GvKkDTy4
ejrAXhWU92Fk1J9817UUnnXp8osvshMxm1qWYXqS+9+ArZeaY5ug9Kcrz8JF/ypjopRHzw69BQFj
COn3b2KZE1VKNfhiLHx5LpDgIkA+Ole/ZmNJR9pePIqzBvqns1lBWCc0wR2i8ZL41tiJc3CAvllK
neNautpEsTCLji+bsN5LovyUTuOpsaYsq9yZMcmd9UkuSR3B50I40DQcJt7nLL1+fxuUDFTPPueC
5WzXJ8ZCq7nQirAVEcLmzSFARd/fcupwF9P7N6UncdJodsxWnhsw6qKxtG0Wj0VXw3Kbaqv9kYlH
yg2+sPo+Ck3BIaLCgAuWmPvUzWlDIvmR/k5SB95DfCl7RmBTIWHx+LPYwZ+40ucIEDkp36bHNyRw
ZAVWZlVBtrEdNSWeo8jQhVCaE5J/pH3HR1hqA3ZdKtXIXilZpK/Yy6AD1f//nIy/JxjJBAHQn2aw
WSKOUysU9vYGJ7rSo2cxayBkA1pdlEE05IseU81XmEzS/kq772ovJMggVxd419dLfykWzk0D6A58
ZM5F8tCsWBXg8echR7ohjTaZpV94Sh/vVp0pIg43yaUXFElgx4DAMMBTLPfMmexnW5OhWXkioT2n
iqJkYBUCStSc5fv8qnXhrzJz2NJL5m43WWxLv4NmdrfLg7fatASDvczssfNmuEnaIhbMpKszzkRi
d0tXkuKbmwg2HlNDf10Y+pOGODFvJr+c+5JCMfMB1OI02O3PDMz2TIuG/Gp2lkILtUyO/txAyii9
nIgw5EGdbUHSe7+525B5LSQYYQE8Wfn+zkJQgopUuNueppy0zAXHe4/XbYjpHEJGkGww2EWufr4M
GBChWjfXoUUpCRsRar0U+SQ9V1vhXEdKsC4/7tCBi9LKSlA0bl9C62fcpbyq+u6acJb5UarCc1XP
xl2+acYs+kQUhqyyBCt/hGaQedziit+wTboUmLcCs6j2Nrf2oh+fuCoFJtu285Us7kgjZCVsqzPj
BpZhum//aQChwKK1EHrLbD5a13VY4Gy/d5uL/GVbVJDP6iDclA/Coa4o7PISYp6kEZvDrd/3+z+s
/FxceDPRfeB2sGKFxON8lPT01niQvRnvfk+Ve+MbnRxn0dYweA+aLcux83DN1De1xr212WOuwvhk
vZx4RUsQROSIuFfFrCev0gNUoPYDiBjJTErHTBajjTHsJnsficaoTWqeKZk/NTFMkyMxiuOrdIe2
66/coiCIG+xlIBLbgD/VZLe3CW6LIKGYbThA94+5LNDoXkRZVg/+avWqJuPM4UbqtpCaHGoDJ+3R
sFOLQz+CizrfqVlZ+fk2NiG2rlJ9ZrM353+RC8Gb8hKbnt5xOqDrwt36TAyClz2tqSTK3nZPb/9n
0xyCCvtGiFyu7v9DkdIPelXQ+V3Q/J7ZWdEeDrGgl4f93M1TBaKlwwMLYx3wx6Dy5hzlGzpSBqTK
biO1v11VH7UcmaW2dm30kmPXZi9fQA2/AOor7vNPAva+bdsHOP1vW9iuutavE26PZP57lk1M2ghU
Xw2/AAjCIegBl/NR6eWhD6XITTyLSIBs+f80KrLEMXd0w7hqf6SYhXZUQc4vfdZn7zpCjDK95MsJ
VM4Eq0dq06auOiPcj9vPeCL0hJJCFIfV6shAUJNWPFWg+dCkUpCQ04Y643obn10WP6kNAMkfSqYe
RCqO8/u3JOIBLT2/fV8+oyTcIZK+Od/RXh5abbDXIJx7f2B5+gssvdA23hROYpxoZ1Lta/KukuyE
wk9qvhrvmEWWDJ2HRSa1ChQEJoCJTlAPkXTlkXEwMTCC3nnJMHKkBx96iU+0ie38Ucyw7+emvcC/
HEnyUy135NN0JbjzDpIyh1Ia+S5ohxQm4jDptA4U/0JAdxO1bh8SOCRdfFXini0SYhVHnMUDubbd
DvYrp0ENx6xCq7svdK29tCM5LdMwZXZRhk/wSLydlBwzRwzRXKz6d6/2Atmh48oD1FJ2xgAdk0Fk
C2na4CPTcfRZQh7YcGx5Oeyb+jIy+WTkxvQAjVkjoPeLaIoPyVGRl3GvS69q63ckZiPngUycE+FV
VRAlwrYjEpckzFFr3Wdsza5ZluyUOcQHCOuMCjYrBLU1MxmIwq3TLYnK52S8qdHtfvNgLWO4LuDE
GnYCBFo9LoOvzRmIKeow4JVbswPRPkEU6665Be062sjJnaQCub9zM69ygVSU6XmQZtyC4XgWqeAF
9a1fPYCsJjAx8Xd/wCtHmW+p5FNCIOk/TqfW++2oydI6688A3SY0j7SAgKUdiBITHrN3nUmD3efC
5htCTS5anI1pn3rK8ftSaTZnxCun/zFQMLSvv//hVlYrjuAtbFmGz8OtoGEs5CoaifG0e5yX/JZR
IJefOyC+WtC1y1Ec82lDaVtfi9IIViQisRtSBtamHSL9efsA+PDSbQS5Y3SS0RqAeYuDuRLa7iF6
lqgfQRnR7xA2E+yEsqe2ixDDnlxm7qMJdoDzYaIy6Gdq3yx5CXan8zT3vEzN8xHk3ZQBJLVANMRF
Te3B7pXjVc/OFIeGzEKEzZvc9ik/RoD8WuwsWDg3vXxcb3/KgZGfbNFCQBGu2Sr5R1bm5tOrsuiD
jv/ucjbjSjxzKZyJkHDwPESE3+8o/rU4+zugmx4aZt9Llp4t9dc4FTID9h4qsHMVskT3uz0lFi5u
JL16MLUrNtAxcwjaYE993IMFNLanQFOlIqbiWgmrzn5VpNEIPHfiVc/th54tmT+QrmT+4BDmIamr
aCtXr2A4w6H/hA4o87pJizmFkYE+IKjabwdRkvnKcR5ayX3lNKc6ORHzmI/z4bwpm8y35ppsmTQd
pKAjlHoda1IzqVRdd8Dem09hbHXN9xozbfWJ8DA8efd7FWVvYriPutaDK3yFrY7gDilkV2UBzAP0
yTXFPT3X6okk3wgneiVv3SoG3QCcZiSqj2jY48ja4xkJaTmzGGKhslzd/ycgr0bU8FyTkyp8uu2T
VEzRlIzPWH6cm/UPwDILPhGQ89E/eIjMHLmZoPjFjHSS21w4uvl4fJzimcXpP2U/UheSxjptGFVa
/feZ7wihAPGwh6rNBjhB3xtCQX2Nx3yciu3cmGrTErS9uUtialad8r4YPbY9FiqicGH5IVi8kcLj
AVX19mOK6Gpuaob+1uWtKOjlcBCZoYgjGmrbgDq8mxayYZts9/Tn0vsbs021aC4f65CGRdl7Q0m+
rnzEAZLITtTbkYUxvUTr2MrHe7FKn2h0WE2CUZBDA7dbCBbJGQdNgYE8LIsYYZWga5+cotFdRqDN
HrmZHYh9I4v4qdsXiLzLJ3PDBdC+ftp0IQL28rGoJUgyQLdEr5tAMTNUdPcx8PbBP1FVadFqAdvl
8IeRtWT/uK3Anhx2WOSbRoHKPe15fRdKTyFf3gOVh53ufWcQQqSfhhWmwWoE4n9RBWHM4P2KzoOe
LCpHM7nQAxS8c+SefkbqzTeG5Qsc+wdSrtt493ZivAX2gU6Pje/draNxvXctmHGJTlsx+hczrp0Q
AfGxMzYUiY/NRB20tImAGzoovUITZUnxiiFt3UK5o0hdKVcjd9PwQtBkPeydtEfm7wI0gbGiSyX7
gLksXa6Qu74W63CpSx0sKxbmu/nQJUEskqaxV7lZJsdDnJCSJKGhcgkAj2x2SmEyeH11R5O+y+vy
HCeeWXJCgOYEQpQAiNLFdUgzF7EZJc/ACxJlI9hSu+T7JT4aWG/jSCfYhLbLXT5M7khLhcvGHWfc
dNFKXQlg+ZNERIzggkVXWviZ12XxG3kwBhFxBT9OVxAmItMMIq80FNo1t3a5fO+88NOzAmC2rLYE
BGPPMqmhrp1Ni/DyQW0Fui72rTy6auMTK1/nOty8jiyiMwNihNLqeqCUYcR2cOgS3RXER2krOj8x
BXE1eeSZOYBGO0ZX3Vpj5yK8G4t0kc8YAWgC9pFNaymgPTqmVROrbq7AlzFDEq/RhdtWaRE0ksPh
DSYn7IY5KTPm1s+Dj9yXzMYpi4apADZPQExYbGDQtXiNy9XEKpCLc2xa/FV+KsmvgI8W6Wlhhyy1
bbfyCH0aQwX1d1pb8qdC8jYeeWcoPmgD/FynsfX3PRpqD1zA27lh1kCrDGCnBlNjrLBIOXe5ZsH1
F89I1fvPMASwd/MEBvoysK389cb0zMIguMDx1Vt/VxNEF2+mGV9Pb/JTRSIdZnG0ScJVsP31AdTz
qAL8juF7BCtsZhnR0OuqsBTEkmYllB6UH7rSJetgmr7sqPNqpwNNVzfuTDuOOUuHKT8EXZqzzGDP
7E1B/4kXqbjtQxPJACWjIg2I9/sg9bhuqXZiwDnINe8QarYwmmLS63kSCcS6ciGW5+auXNbTpVdD
LcvdPe3SYRiJFvVCEfrCQ3b5coReJEOLoqL7Dt7vHfjBfZBSdxPHr1zjhY996kTF5XxOIXPALy7S
JKwbLggvhmg0QvbzzBdeFnAFwynwm393K9hk2W/Yr1rwqVqmSecnte3FfShG7j3uwOitWIy/K7Gs
AMOrFbtc18MNXzMDdrnRSa3PbCByfOPZ+LIMywZiJl41Cdb78mZ8t41g3cKmyHclEmMdmNxsCQSM
5z8xqf9cU0Tkge617zUf3gr5fX3lN6apZnPBea/YjFBjFDXPc+0eRWZ3gsMmId66NFTKGA90iECx
XNi+xOQWceMdG+Ppautha+5/+7B5riYt7VFOC9xMTxn7tlMY1Ns25ENcJqRRBLD/nTlXCZhcYi+T
lf2zDwDLSW2SN6f+u8p8Wf7a8vwCr+jJwV+ojvZJBq60y/XcZkuB7/b0FtKasyvMHhaFFGD3+ea5
p4NFgqQh0Xi1XYI/KXGDqP55z5BQVM9cpX9sdFfs3c6X14gOeEwMhhhVJC3c04c1LPzmwa05LbHB
SmV788t66Dnljw0/E5UsxIO45D7zHGm6mCQUKMpZ2PHH0Fif/gTYaLYnsTYbBWx3hSrF4Ebk7kXm
sTa6DkJZzJrgEdmYC8wQZlLuLDWjY0Oq+l+qScFWkkdVWzFbYovBv5wxqRW6P/2RNoxuuLCHG401
wy7V9MAw/0strGFENuB/n2GuglFrehYnPb1iv2Utk1VKj2szTjo1l4Oeho35uASz27JfO8mpvcLb
jstqvd53T5duobmmXyZz0BwaRUDniIbCYs5BPtHaibCM5LWUhzUdoeitv4NnzN4C2DPfoS4Ww0Zz
i0ed0yejE28YRR75iBz0zZi4t4PaeZdqw4x21RYgm4uNm+JzKEeKy5FY9/qiOsRztYhNZ6qO6wUb
e5vT5BfzQxi9SV5kJgy3w8n6UtKjc3TCswtOYYE10nCuAG7jkCXSUhY4lEI33EIiAGS9T092s3Gq
CGkyLfllSnDw9ovvzQmh+cebavftHINWCaelSjuUj/XFeW2ePWKG+TByDwPpB0MO1qWN6WAHKmG4
ikMIM1cqY7d8zKMNOlzYirFFkoExCPUzD/+wKD5j0dMunSPOrW6hrpTROntK0MISYWDXWkeyn72P
R8fA5Sjs4WD3Luv+jaug/mhbtPPjid/A8UywpurQu0/RmECnYyyS7q8V4NdeoNFr+A+CrNCFszKb
+aLRv21xh1HGatH38/s0wFuZrJXLH6wJKbLZ0wVoRxmORXyogVzv2Cj0pmIQgyxrzXNX+BRQVdy7
qOPWxPqzuIOwdS2apd/xsu2sP7/StRpbuUmedz8wrwYrxnpO0M0nsfs/ptDr/aUeesXNrQjc8ESG
kp/xRrbaFyyJfI2eESbvqqbPkhJGrzgkmAD4MdwQhlxdqf6fWbefjoyk/F2Y17v3+UOXuW7keZiC
8OKNsLtD0j7lH3qp4I6Dl9a27z6Ph0idPY8mwmjGriUdrZEfmoC7ZshEa9iA2fVcz/Zr4bJNaD2V
kdyBzKbREGSfMYPzX73Td4hhNwuaf2Lf+1PiCCwUP1h3IIlvV18CjFJ431rAV17GSoqzk3pcGgsz
gMWf9GfLJByUXoAy+wo+gBFYP5k3flrLqI6Z4FYUWu0e+1GajyEo6WCb+73FF/24/DjZDORNJc1J
oGVRXvLlreoNxsxoGF5ecxx2V/XhIiwjYYMMLiqv1o8nYVH+2WloB+x8m0/vs89bhY5yk9WJdYGf
r/sSRpTQhsfC4I2qHxddSgaLIc+egjgymTkPhSk4HuSdptVslJoJkQCHkiW8UDg9M32BcTMf890U
Ff2LUlHAqeBF/9PAZPYve2WIpt/yW3mBGE6guVwHhjnDA3G+5cGhcGnB71//w25BPS/wXiRH9hsC
YWpGJqUk+TpsFZrDCpn56JIDm2wijaIp2/X6ao9P6VKf1oQVEXfHg8Adt8aV8K90+fISp11G17GP
bgWitIPfsHTH63h63ilJpDaZs6+N1ecaQBxBjWqG2K96AemtNh3mtD0YMyYr4cZ/UXWkrvYw9beh
z/ODX7KR0QIE+dPscRWFQfsZ1sD/+kvGWLqZf9DLo+67TIiL0IF812q9ygvydBTyWK8dBXf4hJ7I
EYQOw5Wic7UgDwAMu7vaOUNAVwnaB6lOVyrUk322o/8or8Z3c3y/FJ+ckahXSKXfBnTKABh9Bwgd
BtcxrKjKK2f37KQO4NSCzUIRLYsKqgqmGQsqNd1wnaMMdsIa2ADVeIrUbRdd0muBeqkNFQ8CgnNO
Nyspt63mJ2TSIolJl9D9O7qFfrQNJikWy6fG9kUqhK2QczFT1Ls2nxPho/GC47ngpgOcZRKl+L8P
oPNgMaKoxfQNonYWVYbV56onVYWOrAJmB4Z9b1OelzmrMw/xmarZEYOzYxO1F8I4aLbILn6j/tR9
lvXxpeGKiGWyTT6BU/kMDcLP0MpqiIWFoxvN0fQ7+/zeiL05g93XeuU9ayotcm7FD+ZA+eSswkaV
DgHQWWpwLhMb7/SfxumN1f6uvM8ZWIT/dVE9EmDrvwQbf0C3mfMec0o8fGRVo1p+fCFBDgQjQBB0
TaUVawl9HCziVep+wf09pQeZL1YnX8i/y3cjEgsct+ha2bD6+lFOh3ml3J5ML88nR6gYB0+TYybN
M7odvNYFGMetylXPGPriUZt34+kJYeAoxh62hDBQXk7k+PtwaRi2c+/C2l6nljR7tK6M5oejXR1K
0e6Fmg8SnFZf4oARUQyRw58BUm2VrrfJrMIUoQJ20iPTXAjEpKBI5gC+lTHcf9egFU3J3GJv51DD
D3sLozJpqV4zSk4RzPktLiDM44soxyFKY6+hUNFsKGSk3qfhqfZkwGrFDfVoAl2eKEEMP4NPuQ6w
VgONQdwW61ovQS2b1/Z1IOfeoTP0/Xgj4enC+0zrU8a3zmSL14Fvda4qAUV2IscnSgGN4ExDpFmu
iBMu3i1JuNKwfH4fg9XiwjG0H2b9FMAqOBQ3RCfSPxOeSF1kqOEmTnJt2e0m73BzLsgilQN8RLFJ
QaAgJp4e+zgriuU+FUJdtNBHapX428CmqqSwXyI6xESxqZfY4+vobvoXuFPRuLEd52fpH7wUGi9m
LxWFszDW9Z3hshhKSvun0VI2UKioj/Y25Q4yVSTQFhw6YUzGdTbbZ34s9htpkkh66NKgkSrmkzra
NMb3NZ//ais3M81KWv3Ef68B6pxTmzE5vPlyLiWffKyWlyyK82FkfzwFfwQTqnswljQQM+Zdc7kb
iActWVRMjlBQ4CesVx/UYQE+LsKP7FMtDjK/d3ah0jxBhJsAZPPsd4s/k2OdS0gD0itDN5En2v6a
eCaKbOQzE9zt07rG4ULJooQh/xxDiQ8ctGF10zmz3aHo72oxLbP2eHVgOMvXqKsMk+k9eICwSMdK
yU4F7hHaBBeQS9BOBWcbj7eMOoxya3KGAXga+3XlbVECAiKrupdlSE5bTkMCp08PCYInPMFVsJZD
51WC5l4LMs4diG3RCHe4IMQH53W8Sf76YfdiERFmO97N8rkYivXbQNzTDzK3PC2VxOIPRvPymt16
4SbQ8j6NTZV9oT4iw9jkX0rReJnrToqeUPE+A50CuwGO+lfr/34ul19f7NfypnOW2XdxenGbypXX
obGEiDcNlRFtKzldOFGP9LB1KZCzJudb6B/Lpopgml6VbFMli3UN5IXYwCam4IJKbDlZlCfi4gav
IgP64vZ1B2maCaqoCIkxfzy9vv2KCNKraGr5uvnIsIlaeYkjDYf0ak71OYxiBXCCooWb1dmh7VYC
NXguR0gSsMGe3CwQ85hZxMrT+CCuSTz/ve1lkeCwJbaGaxnsMYCKAioMif8ZBs6V4wyYVSaMzHS1
PPGvGom/ZCYGv0AJiZwT5DC7AOKYQbDLl3s4IOfzbyAZ45Q2CC5ML/is7zWd/l5LjLn0N9aeKgLq
Z+o9TkQL8BfPxY9mOjPOCEJ1/6jouuP6MlpcHA5HaBa4nedpKkRuw5+CNnb6pvU1U2LsMQ4QMKmq
gPSreSUpz31CI1twyITIIfFrWCdj22tz+Buk3ggIzItr37/udg7asBvt+e674ooNpJH7rI9JmOBH
acsAQxaZW+r/gG0rC7g8+GEQj7yL2ZlY/Be8YTWT6hev8irgQ/opi5pg8XhajCqwzH9qc77fUBzl
3G4cxv2CBwGlLgjMtakDEbtUGeco69G2JmEbr6+pK+iglqYZNhrw3zWcqFN54BRahfaQ+mzIwG7Y
sUph/v0+M5pqH63I8LgJQyfEceC8MkTzlxibsv/5w2PkctO0K1netQqi4WB4Uhi6PlIUFjSSCDOR
zqJFfUaoblyKxzQG3c6iUJJ8LzG/QJhdptzZbaZPZ6h1QnHY7m121MxNuj9aheAkfMW5qZCfVo/7
yPi/BD1icdYGXx6dR6udl221x9G8pNhkhjys1YiZroSY6Df85nqKYT2pGqWTxLyff5zgfd1CQAWW
Rt6bJdQAOFzn1MeSOULrxFNe4ucD/h0MnghytRJW/8hY7cXM3nI9OR15ssmX8BHFmjnaTp33It3U
sfA7g8JRmeWGW6TltF9Ud+GiY7e9qu55NB9IxvKNhllPyMvEQvJmtRSyNPvGUJLt8mYoNiE2axDy
S2E2nyUgLNTVB662zMc3hkRVqaGP3NUV6mLkqW2s566YhO6E44soOJXc5mhzBrMuvRLk0NCor+a9
7t+VIqAFUdqspXdOyTW7F34TpkLPpAOez/YTUWRg4Fo0x5Z/hSCYlxzVFC8tLY8Ww2j90Z2Yz6CO
S/lgtI+9XfmuqhoeHASAIJdXI5L/Vfk4eA7l/k/Kt8GcQL0y9+bGIbNAbj6oLio8Bh/VpEX5PpK8
RQACv1g6Zzxr6X96bnDvYHyaqUxT+t/JNeUBDStp96rmv1cTEctce37Ksf7jMRMpjG1anLLDlVsx
tYouKTrHiojTmgL1FQsykxVZT8NPa6u3n4hf2fVQq2fRYq8zvL/U8munvhq+PBcigoButykLL8xy
QrJYZrn+5lX8irD5Hv27MOjOvtzdCcjDiMy7YCNi89xim3Roq7NW1vfr7Emd4CGKKiyROpkWe2Y1
OS99sfBjDlexmp3CojhnW/F7weo4YaZOB3VG8x0D7JNb9mhZXr3qS7IMkxi9kYp2YyHHNnaeyXaM
X+TTIR6WktkQ/JTAAht6mhA5mVqf9ur6g5cQvIGJg+VU7aHGXOTuRQOQgs44jnpzJYwOHogO0mfI
VsebNZcCvRRUR02Dbi538rdCEssu6+Hgu+ySDcZY+KPKBNi59DUVONZduU/1bOVWui9FAg+X+j5s
QoKP/bzZ6H9OuJxKuak4rhi9ztSdZ76fezqRUFmg9Xzm3sw9kISfGpEFidwjns+WRX0HT1Uu30Jv
k1BDFwRYJfrBC4kaT4GS7JF8tXRN3WroSvpXyU1wFBy5j8OtmE2vGZSB1V770PLHinedUXLo8qdi
AuMiDRPnnVynmqFtP5y+j354UJA9tLOPjRSBW/OtdfjWMD81rJ8Jl4jA8yqI7mkXJPmjL+xJgpPB
6Fxcd5mKP2/SeJW3ur8zOkcXbSgPm+aIBVgl8ZcIa8Nub+eLJH/rGX+/9TwZTYntTskKlzQ1w7pa
X2nDXB0VGjCUWpHDN/ughLWBj+2rpdykOyx60ZBNhurvwa009n5J2tYrMIL54clXEJdORw/MSHIX
cn8+vm6A9p9UFBw5/2FDCmXvvPXlTYB48OCCYQe1+Q8WW/GoNYYfR0bteEaAHwRQGlh0EGv/rBom
bOMEyZwT9Q+U8knkg3UTxw0MJkmPSrmlMToipXPrsT9bwx6H4Prs52DFWceR6VjM//OXCqz00bqD
QP6/wNIS8kPW6zSYCcCa54SY1ZOFKF/VU+FPltpq9q4C9WNoc7SdxCkBWuy2FAxt2qgp1wVIFYJA
j6Bx6+9v2q14rNmyQS1F6iC59FUxHfbHjP439yIcHFXNnTSzSm43kNwLK0XaEQbj9iuIrPIsXIRx
WB14qx21nJL3eruTNGXmVXdt15CxfPbJvcARGwDvrsb7SEeSca0BOfNAI2Y7QRtZe7Zc8ZfXW//s
LIg8IH/cQUIKxOo9rOwNwfKbWIBwQjI844F24PlW4GvGEoL3iYoq40RL0LMstOEc4qYLuWQZLRl7
Uwb8dTIUKHf7ZyHRFMh5uEV5o84GbKc3D9k3O2l/j4+JmcldGezPC94Nn6wuxSQESZXqvLalmSsL
olQXWM8Iwp8gygE5VueOUoow3kte437O1IpO/aCR3iiMjOkSvbyoOhDXLEhV0CO60VrJ8OxWNAcP
CZRk8qS3xH5igE00/1ara9xIYusSnh8mX5NLrtE6R8fTotr7lZF6rObiQH0Yf7IsZuLzcPcM/avV
bmk0yQed9+3OkfsMAn/ltg9xyXD9BkJ5zgEtnJyOrP645n4EmyeHGLm2tnn8eKL1IsulygRsTJ1F
4uS0YjUNy2y4IrjeTs+S4MtjX0oQI11n/L+Sat2JXO8+GfiqAjjCYSn3z+Nex5z7LlvGTGkvz5b6
XtAffrAoBCvBE9NRWtaGwj2G88VP3Xs6kr0Cc13NTPM93SI1uKOa3T0N/IkCLDdzP09c0s9LlHn4
tggrNnsCG2wiYwxly40SRfGFzzbKqABBRVEJrf//y4r9T+WSE20pNPIcO6KfR+e69TzM11NAThOM
WqlEcZ7cIqNviHFyB8ucY4zN1tzuv9DDI6DRB+via/9Nv8lpST6+ksEUCc0NpODA6Puk9EtE7l2O
1Mrzk5bkR5a2Y0QwPh2ewHHN5i411/WvNv/XwiMumbXjXILv+zIk1Y7PYfZcRPPT4/eAwrzLYZCG
luZXsapJRLFp+7NBIcsEJF2NJeoXiNmrikiwwXqKNgmaLx7XX1C2AbiFbbiyhUUmeNVcC+uS1CXO
V+NbGnHsBrkE+oWuDvA8MUxo+Z8BQDyTVSZF2fEoMzp7u3aYYmov6OtlvORcpPgO4dUcKGtTdXBI
eJDwJTl9tgrshNGfD3OJGosT83wLztczKZQDMV9oPWD3jolCfItY5OJeoZVSGSjucLswTCG2nF0q
KjExxQDMGZZa4w46gF11oaAJWa6Uy8kJaj7GvOn+hLGEorCBc9nyupGLJnLToHxi7MV1n4Qal25s
cq9/+x2ZEZbznwWdnXQ/5U/bI/uv/E0+w1SDBIjeyRy2SGLVHBiYKIGH8qVavkC9xBL/cdfVNv8/
8ljKidQHcHxTK+IVehAnCKZN0SwLY0ltcgFhu4G2qpf5zgaCOUHZgd4zmNnxPejJEmjrUQnLtXov
G+Wy2NgCTBxXyljHPPgw2zY1aqvXPTrghqukOi+k4YdWtZeCQ2lqF0ob1eVmYU6OlEDUmwIUlsso
W+5nJPj/5l0D4lZh+auJHoQtz4JYooajaMCSG4VS1brxgEQMSAg1xvZ97oSqVGyBjQtOnjYmL0Jb
Z8Py9wXBVDqdVIZcqCalvNOI8FI/ojzoRWPqI7rOCLtYJAHNBagEwU6N+5SNaXxm71UchPELDRO/
1XuKBqCI0JxStrjbMxwCPgOLyKQQ5VuNGUh9+GxFnuB7nekcVCNUQXW5G9eDESga7QCiqTnhHwWA
LdVvxw6KPKPOXyuGVkKwq0WIYFWTuK83pyb6ZfBoSeJNwXt0sRYRLB0AklUfjs5uzfaQ/GlY6Tvd
OvIxH+QrCNtFdom/rzsKxFeN4qrpOiP2mut62vJUgL42d//xSn1vTtuceIdrNDtpfwxM3Hp/yWH4
Sod3LELHyqg1HvYnqhW7X8xsWfIzNEWcFQh/TXn8x+ZkZ3IlKziDCjR0z2ipl0phZi46a49iUvM2
jpvvCJ54s7GASiuPxY3kGkoKOw28Kbbxb7TRRxEYXdpGfns4iuM2jNi+QuFSkKH5JdTTRBeYyLYh
YUYD7c70WMEOC4GGcInxtCkX9OdnOojyI/f08E88gknlDGaZXPCVf0YrNhWwukH8AB/tt1Z3N2Uq
L+2XXT/ABRrCNo1zbMYCZX9eRaXRwpwiMf8YXD1no1/IyLUy/S0K0jy0xn9ev6RcLWBWvpWRL6L6
waCGM3f4XONj8nMbrC0UWjjpQ7BMkwnxDpZ2r/Yikxg059GuqgcnPkQ9Q5I4L5pDJ/GM6v/cYz/F
sWKoHy9SiSsFy0zsbHlC6Hx+c0UhNkj6oh2sqxQoT2dLytYNrH1BBI4g57K9g0Gh6TR8TllBkcJM
sTtpyXeoaSOgMtuQUYGfYXOgpF2vMiSUWR3FPd91Pn0QSec1wVBpIMkHnRyFiLtu+YiDIbH4RyV9
O7gegR8s4XaeuaKmPWEhqkoC+diKzew1Ik9kYqydyALxZbUlnFpsNS3sqMnyYhLNpkBijQXDCpU1
iNAtURRWyn7qmxPndfa889VtxXibcuLOSujBwbrigaMUYq8Jf/P5AWiU4II3YYMh3Zqn7IB2lqRO
42+mSi0RHH+9QHb1WGRT9Izh76niXS/NkQR233mBeL1S5YmyvHmacv+RBsmLn85bVVZtBULSE2LX
CUnovdBhbw4vH0dAi1KMWv7mDdzmsr5/BUAHQG21kP+o+M0opEsMiy5g6ku2NJGMdgh20UHiwEex
dk9aMth6mEdY6Kdd6+nYitDcQrt/6uKX74aALKOMEKSfhrYhI2RYsx+3/hGWuMDDnQazKtyDrjCr
pFTE9UIwbMpkcQVassmMWMnuwU4jASZDJ8bKvM1tfJv+omtsghUAyPSbgn+vGQ4bDkOcGcX+L//O
dQGRBM2N9Pxwo79T/3XE+6VJvDYtX93uMpVD3J10puPHda23uI3udLfbirbH7HzQUk++mqa3ns8g
yFrMZ1w+x3w/8lNrAyAY5cJo09EdYY0JiVryxgu0A5hB3766wVmMCi3gOyLFSHiDB72yxnmdagDw
rWReAaMnWYpfzD2sJOv5PrOa2Na54rX+IcioOBcy/koKhvsW9Yh4fqABBt0io2V7e9Yr/Ya938NW
6TJ8QkqzfiqFuqi7sy9/QWNToQ2+X7FDKzoIj9Uz/i6D2XnpKIGIkjiC4ks9nhsKhHCxW4NjC7Lc
yGj/QinnJ4IgDvoeWtPE3Occ6WFttYClRvUovw0lrbPY16M78nbEIFBr6nMxpXBDU+XsdJEwOBgI
ED6zcdt07x29a/GwEehumo6IQnBrRSg9LjXZ0aHUq6xjCmbiQhwUZ3ZYOYfDROi6FmwrGcTZjrB3
OztTC375ttzqR2wLMSr8oyrajMiS40KJF6QhwuYYmIsxGFRkJjpn5qRqbT6T+13MgfOo2VKxsXm7
/CQbIzIG4aaKKPm/RqgSZAgwf/gb6qmAy2f+g4GHxQB0dRMUsvq8IvhQmS6apbrSxOtPjI1hMsIa
968QT5PoqDjHRGGh2WaRIE3e/iDCYm0LGRHzkgwjkDFP6O8L7pHlxtVIHq3r+LIzDd0Zpmlqs/bS
ujUQ8YxHZpGjPakA3lzfv+YBFBlt9NPFUaZxtTQOIBFFGljilEi3eA8pfS6nOTRr2vaF6dOosvKm
Tv893FtG/36434lC8pfwIInwpBYJb9j5z6qcOsvrYfUohZnKMDeY+to0xSIcNuapGFYDMBEXDuQv
1fuWSsSsToUXewFUAmqHV5/+Mjh/VqmGbFmZxUs7Ilb+zvlLhxWsEcCe4beZOMRMnuFuYwCCrV0f
j9PfDT/J59FCUtm/Y6qiwrsqrK8zLolrI7y+rbl+2OFP0ZYpZQKO4k1SeckHZ4fIX1p9YpE9zVXF
WOLhfoRb8j/s8bcY7c54IaFtdgC8iStIyBRuLgPHn7YII8WoxZkAhSwVaqhmzpwFn6F6HRmGl8q/
NgAedLinZcI16yqDhkfM9HIRuLux9dHq+EJnYHj8sIv5I0Tn9J76yCGpf3elR7k4nSDJt4XiDG1P
khUaRSS+ZBpcFNx1FQGgPO+UqJGvmRyp1jrQ62c0q67mf/1yEBJEhXfzrXLZDv8t1FlGx7vdTDfe
1Z5kFpN090fDQyNBcu2VKATeZxZrRMNFpDv3htqPt/5GyGuulgelB8PQBz3XYYlfBOhe7d18jEb8
l+yuI1Qb29clSE7kUJJ+rZ5aGZCp/Tup1+9h/FrJEYCThdyPW53pu7P1gPPJaBQNCVokhW5Txyv2
BvtViHtHpRcW9TqoFtJ6qb26keYtQawS4RfF7UvC+4jEfdJAGlJEv9eXuCKIMY4wzCDBFr4Q6BFI
5yJOd1dK1LRKMa0/dtrGSdxb10s3c/f2smeFqxd+EUZpVxralpKSm7HVaSZrzjq/yzlXBeXtfEPE
L9dAaLL/yqLjsFzpJDL3Ry7saeja18MT5y37HjYyHxt5VLR9uA9Q7zM1qMJA/ioxjKFyHBSOPrz4
tng5e/W19iMJSNfh/XCO5wjiFI4duzSKItI5CP+fh64YsO2aV+sOZVrxqEIlTAejZT7MfMwDtxcU
sn9viqH3JMm29LkY2xqEtQ9fAjy4MnOtuqehUxMnWvoPVT5MIrCrkULCqFTrgICSrCPmQRq6GJ6C
wGksoiO3Lh1TId+eFOYmcuFqy/feX3d9XfYe/5PJH3Z4hkrqIHCGGZlzFwutINqDpoQE5/VLKdUv
Y42eRbc7w+RNOnaK6ZyoIQLqSdTQVWMxhlWIDAtpEm23eG9bfOCo+jXdX1PMJpHojffd4ADQ9pXM
aZJp2HiEyJeE6SuInnpB0nzoP3/VK9WmPpvowC9gpXZIgtASLPh7HNOOuEQ7aaBSo3OLsoSmR057
0QFjpyMSUGuXHPKRHIzls3pdRpYA4gEi9FPEcWvD+6OxrQPX6t0D6Pz8abn2IcggQUwTsIOkGofI
TVcdxO8Ta36BFdin3Wck+uY6rb1ULVcxHejROcRcPpozegwygyd+c1sH2cUb4bpTXhKZiysKGWXF
7itLq4KvpJPRkS+LbHa20TD889KedyAQxZmtrS2p9pBKYhayisz36VXr/ccfLj8t96st+G1pSvIM
R90SAhJHwiuw72ytXdrKTZUC5qLOEXPftNyiOKKqE29uY7yDXTcvJc9fquCSrRVVNt/RZVqBr2hC
KhEBRCbATqsD0uIafBpNrcA7jKZ3hR3+HneJI9/fdMTbnTa80Q63YcBI/9xSfkGjfKcW2CUDSP8f
FYefKFNzdqWkNTLg/fYbcXiMZK2DbybeArdqMmunRjDOXit+R4BXCQlX6Y1GmOIVVRYN9y8wkmyT
0HqAyzD2Mt59nnhiowWGmvQmmByCJZ6m+jgDWXWtMPO/wPH+i54EGiLKK39PQqX7qJlRbOTe8O3H
ngODu7N78Nc8WKlu0q6Vj4AnS7NpJY0JUKVvGl81Gx9lFtkWHPDLquzikX8V0qqJBzvog12LqN8h
csPCOfTaaFydyA8VEizR9mMjxLYeIgUmG6vU0hSmvMoZvVfFlfuiP2G85tc2V6RaP1uueKj4HiK5
Q62+NLVFMEHbPzJ0yO53NCEjIiYmpgq7yzMW56C6H3UtHBsojDTVjbhYNmnYy3ZOHGHOCwiuGIIJ
PnPLEUiu2wAtEnKTbb3tx1hfy379g/Y8mBzYAqAgAe1q/Kf8VFlY4SYp/rzL5RVdEXGYfTnSwRut
bJteky6q/OkbgGA+Y4HKdi3TpqcxA0C6+ERolZSJ+T6sjDZ/W9YeQgydYR+j7jiZkFRk/hRLmK+v
aBbtFBuQUsQoBv2XG88RS/Axqolsd60SYmsKrvwQvvEXnLlLDPNbfSRpfUI1/giWTxdJDCl54fG9
ZwSzZGpbjJcFXEnHn/JgMkx6BxT5MedCQP+yBm4e6MPsTsFElbaBHosD4LU4shMxNmdCQMOEE8eo
QeuNTZ8JAWMkp6kY/G9B4mjhFrs3/+Pkzg6Elms2e6QV8EjGm2oy5BW5mJfTsF1uVhq2u9bi4ydf
zL4LLdX1OE3iX7vctQFVH9SQKe5aoQhwuqQE4X6lGDKB0ta61D6MyV4oNK7N/KuJ5pqo3q2shmV5
UwG+WpoS9xnhJbIdhpUBukCgGmZ/x/aE/kkdZAhbsQVvimRl38dzalz6kvkP78lIENxvwcQeNU8x
4tUfzL0Ge9QIKovZbj/PcJQNLOQakoRpKpTiNsaaQZF1EKk9NNuQl6r9eqsyUF3v/WiQC7EJs6HP
jAyzoOe5WR7fdZ+Ep9GX7gBi0rsNteR0mid627gGLTu2UrHi2WjT/iTA93DS09sX5femFOi8ncdo
q60EwmYn/tnA26nwdSSPfM2vd8geeCDD70je4e5FBax/WMG1AKSuDnoq3MegrrVBgThoit8Omq7D
8Uy5TUGydEGpRNuWAiRhi68EHceeqjl2rdu+96ac9V9gF8BtI04tCIv/JOHlwjHFSgkSjh2Z3H/U
mdlzxukP9OwbJzz/ZutaN9FJRklYlqOmcUrFZ4zCM8VWS+OTKBXXavt2eIpF2imQsPw6vjvP1s8f
ofeTX9hGb2YAqSao+Rr6WRl0EZnBDI7n9RVVgjQH8/muLDytf16LWkCsHIrFPwk5iTQu7PvxCJgM
jxcWpXFhQAvQ5cF8nOvbyi0TE62fB2P+dnmTfnoAgtO7GJdCW5C3L75+A1yi8Vmv3SoOZ6ZIZh+Q
i3qrS60ADOnggsg9l2wstbNAShtLdm8np6P8oIjwXyvvv99G7Tz1u/Q4CDSjqt+HfMDAJcGYU2bw
5AMg54AsdXkETMPIcyPBWwhv6FyYoI9x+HaDC4SevAA68lom0S70GLahpAiB6TWtt7rlQHBm32wA
tEynet/qYfwpoNOe//J0Sgzl9lg8SEpvbv+bwMdUtWFQrzKco7zHFwo3cjs/sngADJXvKGxcF78j
vasXsDTqwibZrk+QqYRgDpadlTUObvxMFhlnHvK1VS+ETPld08lEXNBiOm2s0jw40cvfEwcOJaqj
H97pr6rD9D1XaW61jUQFkZznYCmYgnMmKPk1pyH3TnNfhn5nAUFebwbz9Bj6kpDwlvkjPenFa35O
zwEkTWUN8YnAdJI8gCTZ5CrPwaHMeONcxto8CbyMu43UigBWYKfHPO6h7KS3PD3vvAuVd3tQ2eq3
0I7yI701HcQRT0ydkxson7hWUzmor/z415zdes7AmbvrNU7DXW+cunkNcJWv9REy3wMlfE6OVWD8
kaJRg3NTDTJ5YnvUijGICbaCRLm5A2yMqfdD2OS4qF7G51dGeKwuZHg1oz/wXbFEMkiaUeBAE9N/
5SRx+g3ga9iwcjmRRzsC7Cs/y6BYaWkwVmVB0ltGgacTAt3SS6J30xGDGT0nFx6fqmA6g27AQJqJ
31Wkdsh5j03VvcoXl7BXa5uLdytY27xiSQ6vLMEKO3R7czruZeUh96194yPUMPi5yu7b2Su3ZYgp
hNzY9oGuGdU0GL8E0SyDvdSsHu2F3boTPIMVeBXeMk6mm1n78cPwWlSuX/GiRbebSCPgQWwQjxK0
ozg2sghqySINqJZ1sBPGCtkdB30yXZUFNvtvAfoLiaOEjL7jZVhvB/04OL+y/Sj6ZZUPRMqvcBT/
JAp6RMt4heBfVAlz5W/4fMZ7GNJWczs178VE9znCZHluqUpPoPzw9yAIOlKrjpj8tptNJokNf/g3
/Hnhapo89oayc8Xy5VVZL231Y+ikQ1Pxsvg951VUy9VSSj4e0dP6ZEnbn/aVCR92Zds09UMciX77
fFLVkFHpU1/2w++vfz3CZ4w0hiDON5H2Gm8TSgAGHfJpkTJ7ngvF0Wb048uBzqxhKqjVnsbdFUhT
SvaMhikET/XSqIDIK2yj+CvQhoOzbD/v/J9MUaM49vXEsOzzncb7WdyDF4VL6PRFNMKskkbKUE1s
HWL1q449XK7H2jSV8ta28UnNXkngqtETyZaEFY8TkAeq1QNzOlxZlrrihaU4UhQxPfJM/WLnh03l
p4rmNpLqCU/U1/0xF16q/qcqaQWlDBKHIaYVTrR47cLDr2umSI8fpDYxkbbnzkxiif2sDxPAuOi6
5bBxH07tWOa37RIQOJWhG0EjIfQMCAKGfyFbhS/NJv+/qFw35smtjRwdE7QGfavONFZJuQHS/9M7
bVl3TAVZxvELcs9H0BOpF23TkBQxSkwZlkirZ/O+D0BwydJWHSaLjBY3hWQgcuXng/RIU91aERVi
2Ta9fb+LHILpNDthFC97mlOBHgb7ig65DVza8sc6an3Vz9BqsuqDI/oYDuSqiNsqwFrKGk3V3jyH
3QeVWm4lwpgJqceFxFgPVtKAsz2uJ9KbyMgz+tIPwm80ekUxvEJKsZV40gfHgFWfirJasYHOThZv
iNOEO46fUxLMwjR3Rn+JhALtTVB1EBWLC0NEiuPpe2XB5NANNbSNtg/BbNX5sfzY4aFvv/6w/RDW
XCwwvsgPCEi2Jy6JEMpJGFANfOw+7lD7rF63AihWDBAujfPSH8dTq263AObzzSDM+21ykYsbnZW1
cDyry2Y85WiFtr+X18VOTGgwOU6imWJjyeRnn/HgzHJcP5mcsb5q5iDw408FhIsHDDXDIxacp2Gk
W/yVjBHnRaLpG9NPtlFQAeDYmmxSEVlbKEVZ2g7R8NT8wohbW6DiMhyVWI8IipCAs+o8FocszYBr
QGARfFz/ESdx30HjEpH/9pbGMHxJ7gSIT7pXgt457EbMeLx2MRCnCgQDx70IVDOu1alVVWoO/KqL
DH4Z5UXzulYyaQXWKrgiaqkflHv3fh8LECxjKIDdvBCusuLMLE8W3ckQ2i19h2hBE3Y29jl1K3jb
hNF0V5ocP4PEQnlNNCVwxB7oQDqk+O1YU496hMSaQXXq5g5WZAjmoxO9iR4Lp0CpmJL+wEIwE+C4
T7gqUdw2XCc96o/ZMuQx2GW3RqA4uJrXVaAYzGkF4jnjoSWd+tWDGAEJciSukIHo9TiSwG1T56g6
j2zOzyPGtK2ZPv3wbkuvn9CblwRrccHG8Q7RkRbkBoKAmat3DK1WYK3/Q6klaK8tynMyMvGMYimM
/LJL1VGNDEzYO2hbY5ndWd4ztTOQVzPmyO/2oPGQBhWUomm9REhqUWQFDQjb0znJqkaFgvstFzAa
BVDQ8GuEBY7KQs4Ch2vnAhrt3ihFi8lCOZy653lJRRMM1uy2IFHuL2tDsZCLg2KpIFJq0EIzfLY5
fcMtKIJXnPEO/hiL80CTJLtDfOBfAxLsRy8jwyEOCYAYjjrtsM5j5oDb8i5z2q8FWsIDMvgt4oE0
zD8hLpp4xbISHuBHutYLHGPjo8HeBhlCfdDUXV4FPVW/D16lEQa1Pat23Zfue3FCcNn5v/MXDwlB
5YeqFO/810gUh7Aj/OsqBPijN4fPtwkRkyXKqusasJbDnseWsH/I27p+F56NEeu8uDlEOWNWWscp
cjG4EWqLCOjxW5PismODc9GMWJhq/Ay1Ei+BKuijehqMO1kwVTBBeuecD44Z3peIO+1pEooZg+1O
lWXV+fT6vXh4tak3k3jx6pcAB1CjgUJtxwF0lR2wEJzEcGa9zB79LINiSwcRYuI5RQVkwJntRVoL
6emsF/fy/XZsPERih5Vd4jTh9fM4cnE4ceb78+bdakpuvMIv9byKz6HuEpEmbfQLPlZqnSVQPdM6
1iP03Zkpk5i/7mZ2t7KPwH7KgATc6KeBCkxtOgiKD0f17KSokSS83AV5j98wvF0Q4/SF6xNZT2a3
GaPdfFvZjriL7ZBO6DVCZnpLnrqGcl8zrwuHmSpUeAtoXWXYudvMPXZDuLW+gLoCZVzAWL3HbEh0
u0eWzZS741f5moKabriBi6qN42jXV9Cyc5OVHPTR5uPd5iIH1/ix5cOHalEl+gYFEMzK8ZsXZTyv
dXz3RM5dwauME3Ir/CaSXkYxwUeZ6e2a2DBum3NFzoWqkys9p0duJI+iSKd9KPqCFGx1XKwtuvg7
jA+OA+fF2mKSNH42/SMfT2LIxVsMblgBME7nmfVf+WfekEvQ487azfZO4VKz5EA15kVNVm5yi1EQ
V0Ef3SNXMHpOnVUFeP8bGnpBM7lAW2+Tt67MhRApVqL7F66lTvE8bewBnqXmDeDCUA9EN2Iu3Sb3
c4UjU97VUzc8glw93v+E6dySkeyV5cBsD+4yLPQkqI+ufxGWwbH5GLs24WklXPU/DJzrsrueUzsZ
z+iArIZ+nJJhqWr9ANza7buIVfr4F/YAltuMhSOfagbvVu5sTCwLETL+tLWMHcN9Cx3lpT+u900o
xeCwTnKde3pcffsg9GupEhI7pkelX4lB4x2YfUP/qZ65rwZK/s7MIvrstt9QYgmP698WpJSfargG
11oRMOW+i0xAfVVLQZoXmtwCKsVpcEezqFLHX5r/AuvBXmLwk4CDaXXw+Zd74ijlIo98wv/h0CW7
NXWVz/DPuq9LxFrb6cqfMkpucgrPaMhcfAD1l+R4aIbCN5uQry6WsqtCKJA/s3MpSXWw4gJgUyha
Gt+nzwJJvjIjMkkL9QCWH6y7CrXGyJ+pSsb1E4rRmYaiB+k/NwuGJhDmWgSBnOQMxgvNKHLl1cqs
7IH7yMJDC5cJLunIeal9OVm9simZH1EdgFfzbjONyubH+VPZ7At5Yeqt7UHsJ/6OsXqeF7506VuW
U194kO3JOibjl1k1WgHVLali9W7Ql0GAtqCtnshngK8KafjOvar9fcQvN9LzHWTERwYZsb3lE4o/
UiKETzeuT9iuirGiukTbbqZN2vllHorEtBGe32a/i+IgzVhrnXbzgv/VmJbphS+GmIxnQPzRZsQv
MKtJ1rx/ZgN8J6ebuGkDBidjRd4NDSTRMjtgbLk/iASxP1vpXrNKY7s+Yj7YG0rZ7hiWtgM6DZTG
WjP7vMVS4TRjF4/XMoVTAWwk7qFSHGD+LQsvGGNtpEI3EI2kSpRsCgJY5mqaChx/9zCtgSNsrrPS
A/CW8x6TrYWHr2oem5c6acFHiRKcF02PrNRfHX4bvhCCQptx38umxDMYcTxaZzcMhHLQkjYuls38
V0mB441/9MQy4vw9gj+Y3f5/QEJZy+6XXQvnmXzxGFuYwqVNtG3KKn5fWt6KbBVX3yFPtLvuIWx7
LWPWrwwkpBZ3sgXbxXq2zTjqlMn0A9339b/nP1EMQbHHc2uVv+b//9tVtnvyP56nkA3LlnLe+9js
ZuP9+AA5MAppYFbYgO0+9eyB87sCcgMFthFOtfcTSY6rg0xKtg0ISkmc6goSIzsxqehqSZFD3JLc
R1u5Kt69JKiAtKA0IIrKNxh2BSU0Qyg7Nl2eS5wAeyavUKfu2DG3RoVhUxgtlS26S9dM591O/gsL
eb9en8RPtZjtDnTLznFIk7bHbVGBlFzSXYUZiVyMWVAtR+cu9hFnmj7ekkztzeGtZgri+9QJJJlB
RlnEKUbDfInmzOZI0eyWBycFsx3hF7b7w3sRDPTrtfnsN1OYZh8eOXrcuB1FtrM44Iv/3P0+iqty
kPMe8nXg34UJcnKIbHUqmr+wH0YFL1No1kdqnjl5+gtVoQ/N7N6ttSGKgw2qLn/JmcoYHyL1mQ70
LfJ8N47xZAoQfF2/P2n1iqkXlekGJa5ILk9iX2FihW9f4/+88fgmh6kBxle6DHyLZ2V0x/+nEf8x
NmTHzviAwXWjAR/doGVqavu0GosMUCv8Vmyb+fohQEmI4CaquTAjYvwYOXSz8goS7NtGlL6d5eOC
wn03t3h2uoplsr/PkDIptVG50ywGKKYzfNa7AmBv+4XiWYtcEwr0mjL90NZ/K8cagQQl14ESiLFA
5IRP4KxrlNeSAz6II/ByGRIr7O5UIZWwkV6US7JRmjwUXcNPf906btJS7izNhaxqf1IYUwd83xU/
GlvilfWvXeNXM5mjbQ195PumoE0FULfP2FQXiyJW0JULUUDbY8TQlNKKM2n/h8uHl9khHiTlZcb+
FlmrW9ZPL6fAHg9ZoflqX+F34cDAflS1UiFlq+oW+ZGKD5sg1/4yIXpbIF41F0gJ0GoxAJt8HKn8
CA2Tx2rztJkEU3FJGWTSOmXEXtPp5FNQ0pmuopwcPhsEsuMoZuhlx9FF1x6wVZvxZVSEkbswRcrv
2/Eb7tjA7CyMBfs78HAPTpF7+9LZmuD4QY5BHmvvZr86saTqRugr8G09Qs9ippvKJ7kptbaEkea+
tSN0J5QCQWwdxDGI8qbcvTWfOjTvEa2CBnV0bikIWjo6TxnyAsUXYXm1yAKaGKRQjKML2WXFndMI
NF6kbm8cL7Tkhhq1lEL4kgJZqlimr9Zb2xgmCAKABvVnBgEWUe8G5bO8lwXOkWjESLHMJeFs45GZ
NbknIqOZqbTBsCYMGutit5ASsT3vRMKSzq2L0GGuRLdjRi4KApK+16y6OR6il7A/dt927XFRaXKo
3IvVPOWcaE0V+I8GBwv1DHm01kOhHpZdOqUTcqlAPy5dHHlE/917EYnICL7f3+fG4TSMyoCoDWjS
dsrMZr7D2yHTbUQzvAP8qqBsO9cQ0ArtBNabJmDn4KT1ZenDSH3j4qBSW978CPXumwZKs4Uj7MhP
h1W+edtHQU3M5fWGntB+Nbew9+nSBU786F/jGNaAvsbiI6pxYcUoAiYW1gjCyY7QxRcyrsX2JLAj
2+O3DxWOvnAE5T9Gx4SQmEFo7J6bx4ZoJYJAnMbIFqASuPXfh71nQeRBHn+4u7W2pZzXj46OuFkw
q6mbngAHeG/SMd0H3yQMIUj/Yi+VLyAMqseTAI0nczQNmL+lcoieWbYpYMOrabiL9HFGpOmgL5nR
bMO1lbbo9u0gs9mGs0STbqsCu+47BiVWOwj/1b6w71ar5v5aTaiVHPjHNaA30gTCfYUYeKvQwZh7
aNQH6MwWgU7Ff8WH0zbJuSNi7SOFEC3W5incQw2mNXBtEMuN0aRV31G0TLdt+rbLhBDojVPjoLPB
c6fKSlch8z/uNHwy1SeUfhAHcJVEbEgFVEuf+PswgOAp2BP3NndVw2OkXMk89KCTEXU/GdsLwZN0
9rkSsyBM6rGlfVYJ/V6IaDzkB5EBj4yNBTIF39KaIH6eZj8ZbMuAqRx+k9o8KVjr0IfoCOJ+fBt/
7FWKBy7QmER+Sde32nza04SpHSE3/PU2QNDhHeRgaEfLu4qin4YRFDav8fzW+yuxNNeL9Hs5jzOH
f+vZLBqdymyMcbooDuiEsmaZnD6W1RUV83jaCcp7XRznh0/Q577LABciiZNdNybFPENXnvdTIHdc
6G2NiaUc5+O+52azVFfrx83YPJ8ZcBRzAeiphAoX0nBiFFh2zPJ+SL37KFReGVZHGD5866iyOBzh
3yamN46ShZo0S+PXROtlYhv7fx0sTA/GTvSjs5g8R7DCc/LNydrzC+jyuJV0Ipmkw6HHmXRUOSbV
OQR1aLU6I5aAnVAalpnks2MZlwHi247veSS5ahSblMtVUJ8GxN6QYOD9tkA/IglQFbZllN2kblXh
UXJ6FdC9qI/1B+qgUitOxEEaQVVF2eU9tpTWP3vKcMNc8cg4Zc0RrmF88bCOtOuD0toDZlCf/YWs
M3KOt6rOasDE+evT8qQ84afqxiAe8pROYi+Axh+qKEpU2aRjjXYR9z3yJS2mLvOk28UXiwcPX9Ca
Nmc0WYbMxVRGuMIwGs03Zq6CeTQyF1pHpmUzncEf5SyOPsqIxmFzTuJhC9481Uw5TdCjYLm8mcB4
wkrbuF3aF3utH6Yk/FGdVOJPDRx0quXJJm7t/b3azrdZRfwRteWFsVtmbaypEALn0mrro4/gCR9P
+wWd75vUxhtJDBBub9HRjNASADR3GKVlXByc2CkIcgA+TYSSgMV/VzO0Ecr/aFrOp1sCRY0UXOVD
SIt8vXm61g0/bcu62KMd8tJtlScS7QiXX05FgNPSUMO0TXAESEu/j+i+2RP1n/RCmCO2FzKCJeut
aaLO6pKEk19mIEViK9Ttwi6+q4YeWuO6R0ylMho4DwZ8AurRtSqm7GUPYKU64T+rVkizk1GRlI3S
4PtaMdJeLn0v7ZLoxLGwrpjjEPaClX7ytCojougI45bg4/WtJeIh61kCDrgeWw3Tnc6ZQHIkW8b2
Mc2IW1nGH6wzAhrw3crnEWOE7BhmYZsyIPUA8M2ia4jcr0Z63O09CFAeHxqBIJusT1N6sF28ZOqR
hqzfnowj6VnvlY0C/dIrhj1ccwOZbleSt9VxpfiDQYY0KWwUAuEwq695vEssHf9ldeN/ReDhv7cN
LNKBM+7KuM1cvWY5zNCxlhYaEJne6dj6GCOvCi5OJrAxV4yXRhvhiJyXz+fJ/0pBIIz0NdXLmsXl
PmH16QK7NVwqVKQo513eXxq+10jJJs+SUEDeXienFrbS6jldRKeTN+6BZzExsTipU9MvwTkyekJk
YmPYz6nV5HtMpH4PDwcr+8cdDt6JGoPiMMwarQxI4XQlFOK2JtxvLoOaFaHzmADzNcdLgdAefy6P
G1OelNWonai61Q5aNtEzcXi6C2xEHjroQgFSoFPQbka2oMuFRp5Xfzb8RJ7ZfOb3uih3Xd8QMi5d
QYkLYyK6vteSv5VilCiDb+XWyE74l17HolU81i3mk2wCKD8guLVG3DU3Wsu53Z2xoPxV61D0OENm
xuuxxuSUbvyUYbFr/dVJuJEvGT/JvI63DS1rxVg2XLQwD4J6FF/EgARUqfjuWco0JnCEbpXydaGm
VQgx1x5RzYJc4rOSMmC8y/ymDOop7Iz9Vsm0Sf+JSdjCzlLMC6f2Bq1wX6o3AA6x4O/WGPDImSRU
1PwNROakZkK+yg3KXK3haLUOnNN2GLmutuFyrQk50L4BJxrWSxJw2hN4bBfg+4JYWbSPYOABIhoS
atFKb5QC+JbOmAweJs1z8YGJJke3J93cw/FLxP/r9RTb5kV6EsNUWzdN+bFoZH6KvULPfTPou+6w
cVNRHNGQcyYShxTbmw3KGOJrQRR3vAdff1L0keT14CZI8o9WOYTA6FWIqIBd0ugVM21lU8m6hJim
XSegRwXl2gZ4c+mvokeA1otc1t03+588J8f7bGHbWzLQYmU+7P73cmqVWGqMY5NxO3qlYsO+LOqn
WhzYV4uDJSK0mdB97ozNneYezX+Hh+SsJR4hFDCEg/2qRFKd7Zl9nsWW9yxZaYt6/7XMIAC8Wmv/
2gyfS6FvMc/kRn/zkEpDnoaTPsXzyPMEtISF33yl9UA1xceQuutc4GFV3TiFgJ82CkQKlVDdLuwd
F4RpLN7zyXYf6aOA7kEGm0G5w+o/ZKFA3UmX28a3AeYJ6eneS2WVUpsnAiWNUvPjzMv3NA5saQPG
sD4xSywGLK/v7dpb00ucz1LL7zU6tBYN5lm88cu+ieidUCR0MmZNCvTztm8jwwAvYgYwoJDgCBrn
pn2TTwAFYf1v3DW7lj1l8a0PeaaABqoqjqXJN7eIkynYn12stUk1DGIK2xFLTCNFQY8FivghV8jE
GhGqxJhKGxIJhNOHF6ZiBDp7vre4x83ft4mM8gqiyu8IDaX6sQB/TgqqUxgUbkM2cmqivhYhlKXZ
323aC2mHAodPfsH+HALsBknZyHeJvlsyGucZvEKJksNIRB4dERE3wrrN4zXMZwYrUs5/7dmHN1TC
fom44nNIZpjpS4Vna+4lf/d8/IQKxp1uEHT9W2NBLoHhpNkT26leFv4KmGsaBaLp3Md8BBIhE4K0
R+T8SFtJYANCtTu+LmO0yRlpeV8eCmq+oBEZsIVj4zNtb40eaic0LS84hBxxDUonWwlnvBbqOS1e
Tcs1XKjFiFGaxlm9rDrygR+D1N5xDYZom+v2S4Sf7tRPvjmcL+HoLKwvJnJ1WF3vO8D4RnVh7PDU
ZXe3bstJ9+qAoWfns+Cf94nQ+OsE+7L2aeSdB17f+SYNYnQSwJ8lLjtLxA1ugXxFF40vAZwWABRh
y5vR6DMrnowUSMPaCvCAUpu8bEZ8AxCdhwpWLN2qzRR82c39SAbcxdR7izfP8u2ZjwrmehnqFWTZ
tFpwlHgpTNxUobrDM5kOQ9kVG+XZPui1FnWEJ1rWHUhf0Bhn+h5be8BjBkDPSRs3omOUj1YrrmF0
aKkdHDq0hoxGuhc/X97uXaxGy7gF0WUMWJ2c9gsuffV2fnPcTpaL96uESnEHnG2qKF63FQ5F68H+
cg2XfQ1+DcEPxmw5HEQmn1i8OgS7NYbzisQAs5Y1C7/0zW7WVANpcmHEcJ9NQbFfsoU0ap4sa66y
pdPhAoxNJGFwm0FELNJA9oxoqpB4md5fsDVnTV13mf2Vtj0U60sYWEG+BPWv+UFMm4/u/VAWtoun
ahY/ZyskElRNUDTWbZgSx8aoa/DpfRXLdFDG4QO9TqWzUtLN8RX8yUTiZfc9g6XtH+LT53lpttcJ
eg4KT72A7pKFxtxMyM6H9MpIDUhvBOFZLIzLKIG943M54MdyB6yXmy0Y1MMZLQABvE4e4f1goTKF
rxzO/lJrqgy0iHqwBAqg1LlnUWpwX4qqXrnG79KC5LracFUXVRVkYoUW55bzPB3ozgH2QwONc+7x
now2FWpt2fM1qoE4FlHaYPEFOufdCpHWd4O674CYaCWUYFe9pqBeoJAIjsWyGP96yMHUOOKoa0J8
2ztiCLhLBuSj+nerjf3efuI+OZT5h+67KD9kgeHdi6SOF5qQv0ERDnVwSC8nF0AmMFcUaGbSaRDV
PYWnEo2JFPDk8NplPi9R7d2g5t6fd4Zdtqx0wucwV/URnQWQev9IzW8EkQ3m7DZmgtXeqnTCfl0/
ZAw94FzXaEgD1Mt7Up28T/r19Uz1zA8SToFOQmq9EHOzMYiXGvpntICuYzQ913eeKzLtQPuC7Pe6
dE8Seb3rMPT8xjjgNe1zCX8+ukbmVfGElsZAuy6GrYwBVggHFkMvUjn3vKQY6eFpWRJELbTGJym9
pkMmQndLTPG2kggPWV0AKyhDlkpnp+dSm8WHt2fcNF3HCM84pQHz8svfVztEdYBG6nZKxTcKRes3
ma7LiV1GQnvuKpWFxIfQeJVdu+IqU1XWJIfPqIW8SGmDituyugSSVysHLgowfEWLSgSsYtP0L8PI
2vAe/Y+eYZfWE5cL2qLgHVIy0lDpQb8V44+70hNXD8iRpXHqOxsQLIEvIKniOnUzZIEYMgzTdgnk
BmdfE9gUE2gnp2NYXGWSGMg9dV+ywADIhgT83H/fEhNTtlwHZzD8rRxRvWO9lNOuMnPJrhb87IIt
9E91FhUeBbHAPeOtNXy4Wy+IXzBMF3/XisRq0PQ6FrNXXiUSYhG30tBZGerP2ptQP5t4cKQ+BdSX
RUCu1MfZp8gT4KaJE5+HtzYIsD2VOWOaaz0FBcVRA13+QpaX9ECGGqC9PBaoJPoT9bR//fsRdGxg
wUosrbcmHEWggE3eXb3Q1NC7WUfS+ULZohKUHgQP8wQLD2T5g2HjXsv0JwIUZXRN2N099vsAbpGL
d7QOx+te8XPEn6bxxpk7BJR6rqNzIxwZVG8oXfOhVBFF2kJnM+W/ukvc+DoLS8QJAtaOb7mcC8r0
QSR7fukRcEUBCwtEoBZeIb+DeIYHJNK2nhbCt2egCKQn84cwt1lacXnPH7A/RuH8CFEgvI6mmUbc
H38dTPc9oJVManKFyq9zJgkjucX+XkbGm2P7sYeANdHLHgpK7dJ3n6Utz0A58VLejAtvbo7e4H4Q
LyJvtGGYRFileYT9/70r7lgXhwC/2t/AA58KRNfVE+lBMpH/tuKf/05nVVirh//OSjtdlpuHEMOE
c+EX0h0D8X5qa68ExtVq34BDgSOLpKTnjFH4lr4m/qxQfRQoXlkyW30L+Um/4bxixaUkH2zcxXPl
RSPEWtBteNj3XJngf/nmdSeuLv5Xi6/vfv/9YW+fhfBCFsRKFZcz1lGRjzTXuzOpyvxfdTQ/c6nw
iZPu0Gs3Gf1Q6d+IdfDMhfKwCOYVd4rl9A8RxfDdd8uTn82QAYSr976yxD5Z1Da7MjmgZvsP6nwd
Pfg6iUEC9s4O663+unAFtdiP0uKTUfpodqbUOGgOxMdpZIhE+n1C3w0123KzBfd89r3FRV+dwIAL
5NY7xOX8G0VS3Pc4dtLRw3wsb1Zv4ie0HMlGFdIT/zqVvxHM9HGgnBnmcjaqs7HpK1extaGGdZBh
u4+faAN2m4+lPr6L90vxSvgx5e27e8kuMTdlr6hY+CozANM8eQMd8U6IvxnF4isTcSFW9Cx9DQPO
oJRpjNH6V682DhzLzN2kUYGeS/YP5vYhhFuS64oPlqRAJ1gCuZhmaIbqUdsN2Fj/cLmCMMYbulcJ
CzjSfH26NDw1SgKvfC9FXWxr4c19AZcl28oGIXrYoE/hnV0FeakGfscmEw8Uj01quTzAIRy1A3W9
fIhzq/hYhzHrHd2q2uNVZjHj3AGD8V0e0rqBOQOoFx8R12Fyv2opSGfMFEQ2/Az6+ihzweWa3/uc
UBb9KlTZwh+0bNmIzaPYDjh3gaFGrMFwur7ZHSyTQQeSW71bwHLTVvhpKTMen3tbtiF3qRa3GqQF
+Pvstap2TJXkKr/4MIiaKeBLYDv7kGntJisa+g8v9DVXjbXws1FhpfOxREBGc8tJZb2dZ/vn/MIn
8ioWR8Gv1X6GyMFf6XxBfALsSXsxCFtbCTOSvXaNwLrfx/u33BTU+/3qGu6QBbsGHembOWe0Ealf
jJs6rFpBEatywXqlrVLRWm76WWIWvWXZNKo+3U6V56mXNjPA60sx7WXeMqyPydMxaWka5nkTxc5e
UukS4/PuKFOSZohFSUtdXD4RutNnBeUqTVreBHwNODeKxOuB/bgTFfKTLUqp4uvEYZlemf2fJ9aV
S/Gyjl8waCPIKQRlDcWhMy1uRFKwaBzz+SxujUPYPxy3RJuDCagT9pw0ybp9AOKN0/5SPJMC5qaX
fDWIT1G7uAXrs8vU48WJ5HZPWpa/fALoyALMRw0Eszxjsi7H2f01Z95OBamc3nwHhWkVFuvLv9Eb
oYFf+YRy7i+MfIpYJhPsXIKyipgNGAH62lIwkRd/EQ6XgQqQp9AZhnWk4nWp/GezJjo2vup8tVZu
bYpBi+2FMVA2dmzujUD/WSQaQq4zChpmS+iqA9rVAhELncrPkAaF/hYFSCMkPZD8Z4PoAI7VEkXl
fyx+27Jjf4XOXJXPY5AuXEDzi9tp+CZLUSEX/Vwa//WN9mEZXRwb262rP5YJVcJqu848ufMa2tcq
uFJz1Hmqe4XelfPSNcs96UT/qjkjNvOL+kzEKpySMAdOAD8QINcvY+EU0z7bJjQFuutQnVzW6eSV
Ze+m0YPHa7xfeR20rxgJrsjhpeziXY7S5GTQ2fuWOBCFAwidS2Rqrm9bilhPGf22hLfBepPxrqSL
2H159TBNVUC96XoIzxztfdoqeY/UH9fqxk/+I2R/E4XNIUdSPSSQahQIvJRfc9iRnJqXUc+bfhpo
zyDyyd/YPFPTp8T5jvUoSMTcFf11MNdEMm2sZ9yp+pxxuGdLXHA/lTDM9PIFMU3hGBnHtsKoJsVv
/qRehuGqXz6HAtIOIccpXmL7cQPrNc5n5ZkUbPAkWleQ7AJ7hWvzArzWhqFw7nH4T+MIKXnI5I3Y
9M+qBKwWi/OJZyo7ILnIcM5ePGEGkJEbyA68EoRj9Bk7oCOAUGZrAEAhLFWsC8MHJvnEMGE1kkez
sk8nn7ZfzNiYDv/ZuyhvYxldI3DtuJz/dIpExcFTlnK4XK7IIhdKh762IAt7VH0SJev7pxGJnn7T
ZlYPOSvqvY2whfzaKLSd09+QOuTeWf1fIBJ8UDan0yjH6RvKH+RT8DHmub48FHcTgyi8VPWB08jU
Tsiy6W3WldZvYwI4sbQiy3XhJWCG8yu9rKEhby9NeCGGyxghzOr1eSr+UywpYs/wgWRMCIKAl755
z/5GLECzDyKC/tk10jZDPvCbGoLofLtz7dEGIxHfVE9RK0P90xXxjQS3jDTieEkA69Yznkv/froF
FsB015kvaU0CjkkgLJN2qT1b2i2R+9ZsuDCFdaR3L6NcOQIdAaHD/l1ZwrNU5P0eOsOjcmrT1fSJ
66ZO0fganteuLRKjvo8HfHGgWuMxwN2fppfdPqB5ik61QeFUnL2SBFu4mJjMSMLNQpK6b09j9eL+
XWOuxAMWdBKyJnTsrG01+ucbfe6SXZXM2b24tlUgWnrMC9ItgYjGYgdIzmuX8jDlC1U0gsbCwqPD
mnxD6aY4fN3fNCAtOouStgYGeOz7e20CFaQlkkMEj7AFy7CnK4bYxQVXrWqUU+z3wDLtSTBxjtCh
9ZLNv/GjiYQuMnLPLdyQSCEmwIjZzzohL+8SmNYK9Hjl6h0t6iJi8wEC6vJTBI8yIJjiSDUEx5tY
RB3EkxqnIMCl2ixdLukrvS7AstUs9Pn7vlLAv6pMni1UCa59KWfdYVDxrW6s3ZdCgPgPDlLsLUyD
SdSVpGpCAhVlkHQ22b19CD+Q+8z9BSX5QMIeZ4z33+Eyh5ImkEt81vCsV9bXzQ9xWmvbB9mkCZtm
LGUhoPMOcUihgrUSeuAxv5I7DeArKZh8MgGsC4wAaQ+cwE3Ajeob38MYqoEX1t833i0sEqLavCeA
xRpwdDV2R4Wlvxm12PvzdpUvCI7gyXuI3MdN0RAzt/f77c45uiFACmqxjuLQ8r7L022AUbb+teXA
PK1xJFrLn/Vz5oNuXnr7SLhm9xKJ2phTgS8bZ0eSILwRH3j7l696MrXb6tmDKcApRBY8hWmhx3NX
wpSB7tFk9fPZpylSb/Ky+NaQsTQv/Fb1F8xKTXWEFIqbldH/4r684WDwUeKNKIYxlhTE2crdpQ9n
MKjHnnnXG0UA9LUy9R7pHFnq4jbwpRJIDAXnhv5B/JKJVZis2yvv78H+nPyIXk7Jb5LswLY99uQg
VVcpiG8gpSI3Yj2MwbwQq5bb5i+tj36trh6rIXfngbvZwgr7u48s+e8tHJCcRyCJttF3p39rYrx+
Xqj0ijiWtvSodERRgLnw5APHMpa7f6c+AolZLhgacvBHkp8dE/+oUsjdKeF2nhSF677lkxQRatVL
VKVOA+9OB0dEEPU3KcWJzcvCDxWBK9DNDQKU6+keZmW2v3/mTFsQUbv4xMYS8Xly/yjOO8lUxcbh
GLJhB0kGl4j+thiIQTReINRqliVJCSQyHvfD84aQXOxnkMlskc+B4HT55BsveBnAunQwU5RD7b5g
WbAuTzC6ZBIxDwf1SEtAq6+BM59OE0Qjmd1qPaWawppnMaWIj44kYATIFEbqxgsGKEeqxf5oRkBz
AjDw7uOlsokMTJORftrtojyw07EOJpNjv9eXoQkes0TTiE0ZjVCD52dgWqnm1pvCpv8JQ/hGRGmQ
+KYmjpBwZ+bStDrKs4PkNaSLs2K3m/3AbFJVshozo6HK2iuK6WXE/7KJHq4c6Cti1kqkv1UmAOe/
7vKNfIaLHS9rkBmKXjIE/uM9l7Kt6k1aVQLxQdED8LKzvcH90bWk8qHfWSekPozhDMSwnzeT9lKB
atKQDxzWvo+GaGxkl7J4ZkEjsAqxdCwEVobAqTVaoTAEru28ll4w+WItvFjRP1WgDjJpfGWEkg3t
Zhko+arc9NaqoSeiRtoH+vuQRBl+VoIhfYL4cgIRHuorCrOWWKezBjNLQkZ7hI4oPhpsQIlqCM9i
wg1Jysqgph5XmZdRiK5v5R9FCObiQ52nbzVUwIWaqcb5o/q+V32miYXg5F8WJf0Q0lNHwmRbAGbD
K6B3wo4XVMZfzRhnK8lBe004XY/0bXYAzAgcVQ8ukiTd4ih25IN4xQNKIlyJsQvZKVRvhKeNq/ju
RWayICRBhxcmwuAp81iB15E/6uNmyUYN0Rxiv0U+7F3dmDW3XeJSZZmsst7xLE/uoVhZjnh1oz0u
t/LKqsKAn7FBs/9smKW1xcPJfEI/oeot2/35A5YEbrIP/XjnZ0GxkQjTaD0u7GW0SEpCpbrCEnaO
sy1UqFXe/LgjM45vg2uLxaKl5UiqT71JIu4rR3TO60gzL+xGGherxBRz7eVJfpXhjRT8jojhme2X
E/TtoslEMP5l4DUO+EwhEewl7D5oFGiLuXVchwS7S3t6I3ogUPeSWdZt+51HFP/7lgYElDbZiw1s
S+H4FKRR6/QnGfwg/h1pPlUwbEhw5r+mBIAGB+4Wzq715nkscqhzhULmNw8tJpTkf+oQugAlQJqk
xhDuXx62qKrRUGmA41BAAf02vn4eUvB2+sioBXuXFIPX/TF9OHBy5ZlpXAiOQtMFDC6YDtssF4Jo
Yifiq9jfUe8WNZ6/VPOIsLOTInCWzzjHt6JFP8Wi+3KWMRHgRGYPXjJuMXR9FewcIJJPYgPQmHKK
HE+7/qwZ4NUZts5SyIgYPYVBENRgCJ08sI3ce6uid+/kFg4vpNDCrCevSLIWX39EKmZci4bQddS8
IdUArs4YPJTonQnYeC7GynVUHRFJqNu+Fs5/q/9Pq08+cNVa9rHslokUzlIWEo5D/8UoSMqtDtMD
wWl0buAXXpxQ3f+PKfN3ajx+hzoSyzQuBJyPlMzbzCbTamh6poM/RUhpMEcjpFovaHiyV1klfARw
HhzzUYgwJ+XrN8xjm0ZJpEh7+gMbRe9eG4pYa6H1Z/21u0JjFquhgWYWoep0TqdSaTV+Qd6pJcHG
mIa2dzG2Uw3GIJ0FxAW0+sOZkmI9zNwC0gAPza/AQtqtl2c84cwQgJN1FhMQH7HKNixL5keTXSfb
3pr/zjmon7x7z5X0mmuFNPocAKJWBt97TIokjXtjHsvpRG/1/+qLuJgEnnDFkw5FZRvcbcfrV9rO
StqMj6bZTbrXbYyMjKw8xxIICBQGL0gjZTX5UrBekhTPLSlSDRmNMdVB51frc0NvPHLTODW2eXIy
hHkUti0ZsM9id2FAjerIIgliQHxcMMd6GunWrdSfMcU4r/k67weH7RfwR+f5WxqDA74eOKX0ETOY
BRK9lWT3slkvxQq/1BMM+XFFJg7TVYo7Ic0kMqAU0yBuRhPUth7jnQ6IaWuM5IgKvcf3b3U01beh
fWFfb3pY6I00U0o4GjYcA3L7q1FtQmLd6cHqZvbvmQHy1E9646ytRYMPNAbReJH0OdCBkIMpMDEU
kxE/kEYBb2hUMsgR+cRIoK+5F9K2ftIvNXvPee+IQTG+P/51hvzQC2FjavIcD6JM0TdlRuo8n+1M
lf67NhGnhLPECTlsThHF2Pxa9ndHhTjK7D1TWukauYqfrQeyuRGLLZ1m8LxEQCc90BlBWH4UZHYB
TdihQEiRw06ksTlWZ6x1pRTfSFBWi/gJLYpUvl5FEY6DaBGaFASjGnOI2GZ5MbXPfeXbnBOteMYx
OiMXsp+8t42TVR+X47rBEIO0w6jr8XDIhQOSm2HmD9WQ7LAhkHgEFE3XJG8FgN2LYAzXfRzDhU+r
HcIh0fM55gU7t0BN0EiRpgE4hAww+NWSE0OrhC8IqmRi51wwHdjvdiA2jKwvqTt9xzvYQqp1DSCW
CF3xyxholWpdi7ugxm+Zt8oWClSDfeXBsglbxkkxmfuBijjgtAIE1rGDydUlpwyzI3aR16mhWdbF
REHujGsJwO9UQBYAS80zjNFcXrIShQMupsfdCAjQYlGBCFoyg4jBINC2jiTNMFSNWGARP4QAkb3W
DFA3c3vkebl6ACaCA5wE5U1/Tpqo9akgv4SFFRF6e482dXOnSA57VbpQhckL8L44kQVWPweJyUcG
NJiTQR25HDr9DV+BPuGm054XJmnd3/bYGJeyAnmPXTN+6XRcqDvhK9owi01S+3LGPHUVoQjsEUtV
ZeswX0HJkoeGyWhBhdtRefWlkSpwUi1T+P4u2rayDwvjCl9rdJRpvGZTpnJccldGYHFKZNc7vuWE
plrPKIUXzFqDnXMmLg7UVJhQtawm1kkv/EXCHgJqs8n13Q9HKpVQneeZPgbxMuzNIQEeiSiS5cGd
9ghvNZB1E7zalwiU3apsZb9hg09jvWfU4tt9A564pX9TXKcgvVnfF9dKgtpsQuf+J41F67QKmXb3
qGd4U29cIwkPPdZnPBVJQ6yS9188C30GeeI00Z5JAyk5ZBBetmfS/p6GbdlpCJlWTvvwnX+tVKvD
DJqd+8qgHNrARbmCjiyncDwh7JlHThlOtvlErvSCVFB2rVuizg2fFr8RVAp3iYWOEMqAjH7Wu74q
XstWv7OCp50dv+6oJQp3kveraXtra1r8TnSbR/AFBw3q2vkkSJD9U8KRObxhEHrxxKGJmB/gBiOa
iZdkKRBrZpAN7GLh4iJHVYiRV9wVVqoV0w7NSFBfBkFQ+sgVBWo3IgKQJpUwlFKC//F7AYeGPNuo
WKcHZAC1GMupYscU5r9v20AfRQShjLxPjagRbj6zZq49PmsmFdwmcph+lD6xwojX2U+CHKcAcVSU
DXpBKLUldZhgHDUEgWR/7bKu/t0MZf/vildNDHSuiehaoKEqn5ri8SLCiJiyopmS/PqZnkgU+O4j
eZFU+GnDxKBuxyvHv3qCPTSGEs8IhNVP+3otDLtiTT2H+J5w7YGODzx3u3UmFxtPSgZmOvLf7w21
1JiwRznUiYJN64zDJlqu3mEe0tTuEfxJFleqUVscP+hBy3JmQWHW4FKyjO5SAkWmUFzsNGp+dJl+
7VL5OK5U5iJ0SHkJg72TYWImZ+BRi7RkqQYrhnBwI0m6FHsfhXpgu90VEroMS7aWIM+Z0ioRYcV5
v86hUM7TfaLQ0xvbaV6WIbD0gzspgRm8uZdBphb+dbA+vQ16eVeo0ito6oMqFknOiEyhdddHV06p
Doss5bhyd2teeWaev42Tc+e+WTuFpAa1ZWDYDGbtrePMgbm99vFPTq/CwwTOo5T5/U2TR57o+Bjx
2mnILf8T7mPmjgjfeZ8Ci06MVY0I+e4KXTLC6S74kO7092OPGDP0eubuc2+wgLItO0SuHUkekJyX
Tk0FljUsZ1qhFNBGwgQT55lPKogFwW5x/QssQthpCdHovSHgotcdcSY6OzkXP96l3zsPLf4pcPzh
+4ylm1GzuWqU7g1UhQ8SdUgRJn869QOuh4DDuywd9LMkoHrE0eJarNhFbCugPTCGoFBkU3dyVAhw
gdO5RodrUvJbR+LDwB2QlJ+ycMZfy33+Fm17VMDvF202m6QyBpRtbIccXwXEhmJ0UZgtHVtvUPX8
ajSbWhnORf85zY0d3Dg4Qu4kpPMfZ3dpnVAtEydfVit3xquhxrLF1zHep6vkuqS14/nKS0qxdPg0
Pww8DfknHV9hVF7Uku8cnDVY+NZShoqEnHXHWWmPgco6sdXTJJR7oLAw4qv4bRIvYa9d+561ciTO
u7p27gFWHLawEdYW3NkCvzqwI27L5hspLoY7N89o6FJXPk9YADii4wQzbGaOIaQMV7/2oxmmjQWU
EYmGY1S0VH7E3ZHUtSloXNBXudK7w8jno9I90/igtIULqeDvNkJx/u023JU2+Q4mePyrZ371MNCJ
CVRP1qUTmCh0VUwPxk0raDXjnfr5d+Tck/QvCT5/SylFxfRmyBOPeOeZwVISUbG+244yKEioZUK3
pEkKZ8rOe1viS4y7V5W7f+VwQv6fO7iLdZm3OzlZeWO8x+baR4QlB+x+bfigvpaCffCPueOrhNKh
uZbY/MqL0YiPYJhVaIa8dM7etdNWwBCKqAXaWnA6WcHNeCKojYXnVbUKywFiXMuB7hynFYtD1wYz
ncikvfXF2/v4gB+jYzFm0vC3vBHhP27vABioUnYRZJHwl83pg2OvDAeWUl2VfeGjz9mrMKJaW6n2
6rZgEi7gu+1PR76pjs6dw56rB7qccFyZFPZVIFOY+OYHPO4jhot9NOy3qeMCI6XyT9SnjnJlg06K
XxN4ZjxO7goyEq5d3RKsCq+S3KgTTUwthWrdFD2Cc42R+K2xmN/zl28fnc2Bt8s9iZ5Mya7jmaBR
L6rpd5s2h1cH0YmUljaW1bb3AIPtWzTdbEEdM4yKraNGuD7zFff7AB/x9mB+jYOByM6E/BQmEJuV
WJAYef3yN9/eEGkwEK8zblymMxKtHOXYgAAQjrUdXNJJR80zorG3NWR3yXNem86/PDx4g6mgZGyr
CVoPhUdFQN21iMn0HQx7S5OI9VqG+/M//eNG+3P+Sr9jTxg99QhYWrJNtrriHT4EbjL6QX4CPW04
dKAjOl9devUHu4lZo3qjmIreID8ZPGp9gGCQEF8N5ptiGwUtIhgD3O/ihfnxYu88SOz0BIPANUyL
qzKBX2vrbqRT+uv01jgqeGUKPOMeM5xqpCXTMkLFcl2QQP9bR+ai/UzDMX5rLFCzIyVIzMPAaNfN
+sExe/vBnISbSjGTiz4sv6T8/CHyKwXl6x/tr3amUDsstpvACRzzD2laveGOdvIC4R2JyCdUeoIb
NGjepI3hxyI+I7Ajreh26Tl8jyJWTIRYWwSt5jKJBjAmCNNDdY4pVG5Dtwk+MkHm+Dxel8ywXhpz
ByizcwOb1xggaHa10D1JBvxmD9ZCksVUSKvHXxjroU/Xij5YA+Zep+4ZjslbfQO8TSTGY28rsb78
Yg8WBCkL2UXmHEjpgAqkoh6j7IXhT/gjO1Ems21sl3NPXi0z4BvHVKCMNSnlVNFIK35imgc0m95/
HCFMjewd2CzXiO3IkUQ6Wh4h4G1Hr+qdfsdCa7G0PJeRGvK+RKUQ04Lh78cqXD/JSVsnxWTjuBay
Zels43sMfV3Qns1EfdhIqdfbRwonCou8CLUD2JT80kQbCJ2gCMAFnbxASSc5GEYOBHoERQPHDPgd
TVnbDuNc9CBlt2c8N8R6MNRFuIsdArpfkuNyg008cx18faFGr2xpt9cGRE/puiBo79IVscCoImbv
TIysXpLs5QZxUzYSDdXeI9TbBCARzN09IK9pyJ1yle9gVqXvwScSQuFCmB/5dgvLPxDXb+3AFav/
fxxhgPAFQWO3VKuswxd41wML8CSu1vICAkgihzgJ8WQqk9MRGyOvvlJnalM0AbZ/kIyu/CFHPtKs
eXbHkB71YZO2fZZ1Odgbmxu9xhx0DzgTrq71ZkPruwWzq2feQBcIl7DgSLL+hOCIeFeAAHQbKT5s
hJhMstmoiP4szfoql+B3Y7wxp9jeWRvrN333gllfEiJ53A6pUFgq5EiKjIp1GaAU6NfnVcopo5ph
redPWXEz0jP3D3jgDd0uItrkZTeO5cztzFY/gb8usSab8Ubs32hhK7C1prGOXFoDQC1yChJ5fwLL
nZmii0NsVg4msGzhhcYTuor1q4DKqax6eUXulSLMxPi/EeQPBr065BeXEUrBxAAnNlZj4ChK2BF3
AlgaMQ76EIvxVpKPhDkbPHXQp245pybDRJ564nuC7l4ONsXgkgF6tz0Ly2lI5XZQCa+E/hTQz1sF
q/wowi0MtH12rT96tX2y14WnsfGjiuhCzSpkKvDegvfE1BurXpK3hebRHCWXCvs3e8M10HVkCNUv
x68hlwvl89EHkIZUDwVwJJIN/Yd6gzW7sGnkyYY+gp4ANvJtbYirPrB5h42ZeivqMn1NyGH5Qfxr
DzTQhA2IsdluenSA91QC/HWHWIOB1TQmze7LzZPuXTZRuqBI1ZmGU1DPehMUuBBi17UnYGZKvmdG
y6FUwMVIIXF07X0cjI9AMPQWcdo4wng0JMQYNbct3fVwWJvUGt3rm19Ehl1ySh6zmf+JEhSbTcfd
6/YKadSPwcebWkgjsV/XnQHNgztxk0FMNVyxu1jJA2tU1FKSsuq6UrP/xCy5wR0mZ/ccRlEYpl4x
Hz/CURrjKw9x+pn5urdXONl2PEIXTgSvnndejKBRl553g9qLDovEUP55k1v70yOZ1kLMhFJ4Cqtl
yWkDlGPQWXwmH4oHiZzEplfyIs3qapofAq6mntrNtLg2TFY7mZi7bdzG5HznkbvGc2jScqon7qV9
XwqEdImDCvcQp4LiZwQOwGSTBldxp9/NJnXTVK+vUDGWh89Uye9jLUb9B4yuDhIKwuqIyVwhSh/e
BNt654A2vKt17pI5KWbo/Jgf6ODuk9oO4ZTVutkSy54PgrMYZ5kJQ4JPrIQ2wdpAs+bvVdyKyait
e9Po62L5JyljifOusjlRN5/Nk2W0mwyj2LqfXzJHlwri7reqzpxE6TKuURT397secjoyNdYehYAI
WzikmeHrMKeYZKg7/hE2HaiwaGLMQXAKllof/ukmmug3RfKasIv6oE0gyD4DCggU7QELlM+oPrGm
j4rilOTVUR/LLba+J+pQfSqITbBvghkSPH2Zir8gJr2Ley6Yvn2V/8GwkcKcs2BLYw9zgKR1bgck
5x1Y3v7deLNSges6Uk9A19mOacBNMHFYNJDQPAc2JYA0fStBk60E+YL3STiNZKhPlRz3CL9AsTbv
Ry+yQlJWheUTF400abM+CB89APIubgFOPJQLU4oIG42T3DEMLL/C/1FaaRWl1YJ3nxWPoIFLWr6P
qeP8HAzOol47+XmwGMQozoQtz2m9PbpTxtom1m6gqehobBvq87kcYpaBnprufQaxK/X9OMPsH1/Z
dsIIDuV1zwjLg969XMODePRdc7VEb118QGMIzIY4OjhFt6agucLCaEcTPfkgc4eUa6mIK7gaY7eI
JYXe/YvGoep1aKcVfJi7KtpmSNIFTSvVKdIjix2aYTgaDlhPNNN0OAWYZN+QeixXgC2u4dxNgJrq
l2Hw4yanyjaMycPN3q+TbrM80/gPrOpBNZrTLe/cnWOszQYVoK4H2eCE7DBSQG7jaTCamG2m9rAh
ysuAzae2u0XaCAlEi3uTkDM++T9VcMRkKwQt+4QMPSLzoisix8bDSh7goZaLnKUuDOsgds9TetKu
r0Fk/5jvtisyeW3FNEK2E+qk1WxIXRDE7XwNinlavHUZW83RAAP9+GjlTGb8VNv+kawkDEwm3vE/
WGy/EJjV4J+FWdpcZLqN4vskb4x/sH9EVXGLN6rDOVmr6ZzBpbFjNdQm6XqeP0JRukGN3+2MPjdh
OkFtlKSzZnHVMJssZJ0BVVZDmSPCxYZ/d2lUiQRq+Fm7dAoG0Uz+1qCGrqnIOX322n5s6q7uZqbo
K9AXLuPfLqE8MbMx949Zg+KkVK83vaY+NYkjm1Brga3dMnGL71mRTVZKv3/DMZ7+oloudGh7wJmn
u+dXLf+u+5HRoYhBJ4irnZ3C+qxtJmzdDRe+AzisxtUGsbTtVGCfr53UItWVnIDW9pvT1gayedr+
fYKhT2fk7vgTd1yIGhnMyeordhpFdr5WqROAPMlHf7yaXu8mMq2ZoJRHtzw++0SVNqRnyLhEOriN
sYWPrs0e3PYXi8nbMcgmIcCxhaVtcEdxXLllqlDrFwamVIdDvyns8/OKdFBWIGns89yTkopJRAGs
bZx7bi65YWfYUGmKmBGGCweD1YqTb3KYzvSM1ixHtZ1YxaWhqg5OjCuOz92xs54gB/dCIJsPp5YX
V1b+BaKMN3M6YwL2eRypoLGRdb4psmgXYtwAHbbXQJoCl1NRPA03F3AL+JHicA8PILrITFMiQgsW
fTpV/DB3ltEgUW5s58VTL3d8gITKdpve5ERq23BZCxAfcyvglSYNlbgwmKeLXjpWVABOQR92DBqU
gj9FZpum3q/Ts9ur1qa/3aGfsD/iIxv0UxALDUrhZBWMTohAn1M92JlXZJz5rYDyN8hLEbmLIZOP
1C2qov4Ph6zDRZbrZTYAnopE65CoANk+5YjdjT6204nByVQyNDJvVJWFuK9rIOGTrCIVlezD8UWG
5E+5IpyId9WBzCiesA9nUA40Q7TpDzgC7+1FmWx15Pl+HO94FnmJLDgww8vVVXacr/0Fp1gsOMe0
gcIP55GNYBxHCOzirvJfunHzV8KEip7GCYi67IywpadcpbUWv20kvta/QJVYF8R68vAAriQvGgfX
TLLhR9bOwlZMT574/+XS3ccHVoTMSRgXuX7Hvi8om1HGt0hVOWGChTcthTIr9psyexbh05ZZdCSI
9AKm516qZuFfPZwV4zMDPAKMZ+Fu1sjoMcEqKW15zKBP1f4s6VErX0O4teJgcmB1Rpf276o4Mf02
IoOLt2MgvHeUsz7nRB+WB3nw/+H9+5AhW268zoldHvqOacAzQlHkms895Cnow/Nunb20U84gamcx
81op+rRfo9FZZZe/fMzI9AnNIg86D1h8+7tMHhQxKiwbEZf1AdTLZENX3J9lydjnSQ+si4FCOkDC
ST9jgGF6ym2ndmWqEJ/dKdSWVPMSAfTDkGrraE4TePJqvychKtGMGK2TL25/U9uJQ1h2A06VfKZ9
fEgeezrQX9OKKcBuobtjttVCdS/JYxdPwGq5+S/x897yu5ZGnXAk+MJufD4m2ez2vZm+fHxeuWgC
SRyv5NtC3Vcn1CVs8CcI+ov3Aom2c7F0nlsSGDPcKPkBax/7qDLvSqTiAcbRlOTAKpqPU/W2nOuW
ZxAtl9yGMLGxpJ2xXME5MvO2dqioit0Wsaj8jH4Un/1laXJiK1drfuiVYHeh61cxVF4rz6wtLE7U
6EQGPoQDhKsi3OWj0XJLtbp8E7jmCVO8U3rtZlavYRs/SC9t/SltQFvaBZDB424tagC2jW9rxQ5L
d8schLy38OHUKZwo2O9MkTaldeZxbloHwX/AuXuYkHlydSsn95QbGvQEKDvu25cIBvqR6BCNQggR
zlNaVI5InSD8JGJnn6QSnX/QiLMuqyCQ7/LN24YXVb6DquHA2pOiOsJwh5uqK1KHRekYiZcdjO0A
kJN02QomXXriF4RR52vRtNay1jeeGN6fJH6PljZSiarV79zYwpIhrTMgSyUJcFx7V03szgrhz8eu
6EOWYxrleW2vfVJ+Ns0qHs0W2OE0jFNemXp+Cp2TQPk4zDvC2S0CAIEzwDYnqMgBjVHBZ1nCr71I
rhIiSsKB6I3UghDk0HtyX3f1zyxwyDHxqQ6RMmHinFR/YWBYSeaSn8JlXtBOowqgGUI4F39gT8bw
lZrzwor7tGL76I2N2amr4wt3ByCMFZ2OkuR/duCb60GagKGxBpava1MkZMgL5PajsliOe4g/a7uX
xQlDTqb1/QwbakrICYJ91/TAwxxul1puoFrj6tNTLDRahWwy5spCHZboy++kc3B5L96mHK/GkZd2
LcIzapXgUQ++/M1ZmSjV51ACouwtBpU8+7BCMxaMS63b2Zb92uBax8uMHUc0m+nND8PKWG3ku5lK
dhUYPX8EwKDuZcOnFzRytXbamJ+d+8iYY66+p8/S86NoCo7aB95vvkVTIFFSwY1bBwo1WUen86YF
sdPZMWpBucJ5nFCnxle7R97SODYfneooUGox+mlbIpRtktHVbn66d7U3G8FPt2XOvpCYHOy1WBxi
Nzhw/BHFpntJ9nQb3GRXNXM+eh17siTy/88KWh5ZHeI85M4SlSVgHBGDL6UvMgxksTa0t41CL5+W
jQMxxBst9rHCs8AcbGdFArHHs9FCwCZOIVrsquDtzGQTynvRkpfNt5mpNTLmcNBgDjRX3A44m/P9
kiYnRd+eWIkazN+6ZEeCxCNw5x7D3sQ+DaVFXF2oLCFamtvtkSqcfVTpVXRlsiux4w6u8RJjY4v1
6f3FBnJlMq20PIJ3QLcTYWkBO3NlpXbndH3ER5iMf8ds+RzEbc/rODY5gI+TfEQi8ziaXfQiviJq
qXkHwyabf9c2BLDhwDBo6QRhhiD9Rfl50s1S8+eSc0UuYobjbw1sb4ogftLGTNmeBf5iOl93aCh2
mC553QNvMnWeGBQUItjnzaqrd9uNnFTmyg1qp/tmzyjCOclcondm62vNrqcJxRfXZjH6uyCT0M0A
vSbWapiG3i6mVRp12qRITiwXrMqffa4a1AH4eIt34IUVZnnrhyvDvh9DyaaVpx+JNIw3qoynr4ob
pGItZ0VpuxiP3i4M+Vcn+WiVV7Qub5yBrErPchpQQdkfoRDLHRhpP4A31OPq0LzCHMhH1mlBPdqZ
BaAzDGOZnf02ud+Zidvw/h3qiJ8gqb6rapbX+E56LkAps4RrSqPuAiC3SwFgoSNVzxJSoGdo+ZQ9
AvmkmDYbKWgJICVcKdWTJx2BEgupIFmo7zOh6vyCTkMnjgp9SgjaEOABoaSm7Nj8YEldUkEoUG+g
EeUXnW5X0YTR0RiWlmCTuYO0pQdnUTsGs6tgKgtie3R9/0cZjIlnD57mpQFCNrI2ec0jPlRbIj92
YoU5j2LzltjxZa6jlA+PoT5APu9LMDSY1yl8oor25zl8vry+e1aJMw9wBh8BoF/lMGDK2EifBcd+
nY0GYAG3bG/+GHccr3OKkfwPFByow3IbKRTJxXHYttDxWDMCb3BKNkd5BicyZJgcb5ThOkQsU2pU
YdnOxJddgrAg8vqvngodVG6BqDr1gvf067P9mgFI47UNLzTfSW9o7EeuR34vWaMPElPfjTs+VLpp
SH52sFLoW60Tx5psml0Xnpc3zdMVUk1v5kSaaTlic6IxBBqrWA6QG6zVpuJhy4a4fWnUg2w/lZ3a
h4//Uh2lXcwf4OadVwgAcJn9LmsoqG0Gq7W71Nhn8GxG+RcrW4jOD8xB/sxWQv7ETl7e4rjCN1Zm
QuZKgZncg0r/1r/P1Iy3OtxWOiIk1TfMU0XHlPauaSq81yeEQw/1/rWfatwbPKDRftQmyhv06wkx
wwgJnzcQL4wiSV3b4IrXZh9a7P1RBCi1KJU9QGTWjdZiYWIWzep/OpIzJmdDocS1Kr41nUFun7oh
L9aV02BMagU1bxSu+pkhO8SqPNzEe1s5XYNMwr/uuT/kohvnCpyIKAbQodw0llE/uo3JD5CJyWvl
dyEepO3qWnJdJL+uC4VouOmDC+frU1Al4pnQpnyfcXWrERd3hSo6OE/7MGHbZl/BwEGtZOxx8cX0
pndg1US6Gkgl8saHPaVwVGHwL9QhY9gPZ3MXJ0dzqwxu3TGk2C5ID0e99rWoB291zRyZgqVLbL3n
3x5kmZUXTSynlQPsaIvjA3j7FKRVfpPqSZpbVs5UEF4uEYvYXHu6x6bn/Ag3Ym8R4+uLLTz+bueo
TyNeR3w9PI545InWfzgFf6OeCmDlnp4nQv4WPJ8DNXiDnKu+dX2czjG8tQ8+LMVwd8lwQRqpAM3e
42/sMAJIVUd4TV5SlgpA+gDzhH+mQ/nPAFDuyZwAFv5syFRi0qsBKdjy8v9N1Pl4FOZ6iKlaEeE1
iaoEXn0AZy18uPBoaubKWEC3zH6bLNsVm8GEqE52VC3XdTOUTpJ9j/k9Bndc0GYuq3xChrXtjK80
dy4+ClW2jeDll0I0FvV+zfT1eoL+yDYD8XTRqkhaFXQTQkd/s/84ojA+anc5CK0ENHl54RtZj2Sr
m1YIkm9RHLfhcCdbXBD38Qb+I5Pygk4Pz4oJ6nbVykqSroB678tI2hTJnLKx+1Nv/9g3kl3C8TBq
OoCTjhy+6FYz5YZdMAzDU1Kuseu848u9tWozHJVeaDOZspqHWHOujmDOznYE4pBFHvnV8AZZ0CY2
OhGbunxA9YEX3cpUgPZjbCGrvwvNJnsCX+MGIcinZIb5eDZc9zaQV5ZPhAPq5hRs4TOlZ8MvefQe
SiKGSmbwN9ybp+mo+cQgFG4PCdePZ/HVl4T6n3dItN55NN/ywfKnh/aGoLnxMyp1un6WFGiNsCKF
8f7OQPT8HRq4W0UUxPRcgaGcvd6YPUeSZx0YHbGtaLgWHOwe/JcBje3WyvOzgGApY2PW3F85E8cK
zN31N+JOA+AMuZgn3C4PruDQWYAhG91TDNDSm4Qr7UgSHONht4VU0y+Atp5j88UDl+lhhJ4IsVMf
lhi2oN3BKrwLwwKEXr/f2aw/ECJWVwkpUDlCO2cb9yGbD6G4729cXNLhzYeq8EXpI4zTs9RRVQ/S
nWu0B7IXLkfhDY+aND1Tusd52yeZhGiEut1ROBf/xTbUVtbOnbGNczu9yUecFHeyB4Do29+reLFQ
z6qX+bNJAV0I8y61kledsYYOeG0alBUWdYM4ZKYVLT2UQzum1AyO9tH2Jhpbg4Cz7/iZAJ3lPQBo
vxtSiIA+oHAiz36uFLcTZ+1T5ybut0UKV+SX1ZaZ6Qec+Oe0az2iIzVaE18eNgOQJ66Ez+DV2lP/
eUXsxzLS1D0nQUEjtKEFMJQegox2Rq2NJXyiZLBxGikj9GRiYWKTJwS2I2a2NfDSOTvpdOqg2q1F
GSJ+p9FWh/ruyi6VICWXgT4beFD9p3CaCxgtwdX8MyXguRKwXu5P9JIhkslnXLF+CSVoQBpzIR2l
iLktxX/8qN80AoHnhj4GInD6zBBaIxxq37E9FSHvBEbqIS8rTGM6CCvNCslDvSuWn4dUU4Jx06aT
8hYfvA7/Sv6t2zutXd2E7nazDBC+OrDs1ZqqXZ2abXqNytvyo+qR0bwR1nArzcJ40MT5Hfz5I1NY
HVz25XDHoNpjpSRcma4avJBt5XFg9P5grxZiZt0yR/Jm1l6OBq33ikOTcShvjk+RpD4ssEqaYZSG
WEVRn8TDDWn+zmhjUpkV4G06bzpZFztql83B+zbSs0FcJbkfOskCKIry+F8r+bps2cjOLrVLOYvO
pdr7pCLyJONfkaronxLjVEtpPQ/A8CfUsF02084yuZdRZpzLhDNPvaegtES39o91nKcbZCpNt2Ku
Ileit1fDSWgJHUdkHM8MUMXMNineXNz98Iz36DjYamIZFepClrU4Xhhu2wtZaysTjyegY/9NRmqt
4cLpc6NVEcDAYMHOiiJRRC8jMudAsSWNo2gSrREj/sygrC+erWgDVGTpUuYBajl3sx01w8BZPekI
4xB2SQNekYrObplttKJ3Lgw7ZzJIsQeAS5KPSK4vhQvZ5LWaLwBCLDd01BU5cgprWBLbAvMQfLvv
isPgcY36uiAOEmO7JOelwIJd2I2a6PgVaXHextM39nnBQmpjRkWc2Njxh4spmMvDoQVGK6BwME93
Hs1ZyuggCg2tLJqayKZDRjV7PB8OQ9ak2OV9W9E0K+bgYgRCEaRusOBPYmI6gZJaGvMJwt+3G6x4
AyAQjSx8uFyG5VhoUT1wKCmy8II0OL+QoZtSV65zoV+rziaqSQdWUYmKNyPuuPlNQWCQWySZs532
OZSu53vPs/Bj3ANqDjLcg3GOO4X3hwOiN7ivFy8Q4t/yBHZVmIrol4H02z9PUXvU+TYYeFxWULmI
9m4RwVReN+2W9bi4+nsVixQi6hgeqvxfpbtV9eDYkhmKCRKeg/gJ9O0bUp5671MX/YQUG6KBxIxe
NzeYgCUIUE2ZRSmQ776gKEHDac9Dctvc75rTi5DzoqDllcAwHSMx2Z64yUR5SghZ0VSw8V/F9xN2
v8rjIxA0af1ZsPItBHHqnpMuErOH1AH8u2VfFh+KThEWdRYXC+BhvoEWz1KLb9wRu7o3eX4/3fm0
3y4Rb4pwZwGz1RuyZldtX/Cu2bpPPkiAmumWxifaMQATqreAdO3xQy3bAT47EAu6JeS9n6IJsTPx
PhVNF5sojK5zoxgnRTlzvsVejxpMtynUkC7kv9+78sx28V8+5RaOvUWBn160X1YBvInTPYVaAd3u
XiL0h/jJKN0DobA+Tu9gUUOsJ7AfVHuF9Oj+ka+4k33KZt0nGHgeChe5IMZQR0hzenLsdkqHWQ+5
mqF8O7pfaJVNK0+rSjULLQGdhNEnbpdBVINC/XFUVf4RSAWmkTI+LSORYv4FXMrrzFn1GPHqlI00
7iSM651Bl0AjTFwlE/mUF2cSRcxRGAov8FD9nLBfHw4KOYNYBuK0IjDSPT57AR0bX85CSFlpVE/i
AK5RqY5ZfzIXqfxzOvWCfiiGwXJp53FnRCrlatkD5A/p3yhpjQ/ofFT8t8JqXStg/bLCx41LIOAC
YPvUOpohsa8YTGTVc3kQRJWZXFSC7zSgNQn2ue4cPY3oUMM2IFhmhsREqZOdssFFG0smJ2XTIUtN
+BbBL73qgGdZUGa+Oi0jZGij3QoZi54G5syj0GV7Z65gAxL9z61QDaVAFTKsfWTiapLc9JC9J7ow
np+kY6nLUyhBRnJmidf+s6+HPZENUMw//g/97wL2Lj8gu0xcPlYh1ZxnfuL5k2Jc/BC7RQjdG0oR
/GaZZ3rwLXDC/MyGc+82g+1BqVJQiIkVW8pgJzuovIrZJB0WLHB93jDgCWE9ynRaEvOFTUXS2fGR
HENi+LIJOHWKxHBimkgrk7RmqlkKfkckhxIK8YfUNqoO+Imo/Ym164mKtcE0FafNBl1zZKclZTOm
WZdWUiP202EJ3mJqYL/CUHGr17eyLZhHz4RmsSHokVjE7vfRpcM3V1KDmmhr7Cu4YicoN57QMRch
CErexKBHQRqHCjYPytwf3FYGyoRxouNlaauSZnLFLh4LKIE7h5w1OF7LAXzG3e7gElTrCpjSdWM7
cColefzTNzCW1Cxzt0aFc2a9m1WQvD+XwBi7Oj8HvzqEFUaRG5/DiOiqcDhaNDBW8NW9OfkwW+4f
7LZX/JTkHufCQwALZ0KS2pWMkFFd+2rlZbe/Cj5Udhxkc6FibP19C6nwfx9UdS0wZDxDtTzStr21
y7nXh2CYF0V+j+NVGsdvstx6i6+l2XJHXSv/mB4xRqTsC3M6Fpm54fwKatSXZ3Royn7PQqzEO8UD
NdnkvtYO/kiICzm1JvnSmT1ERz2ZBBlc9shW94H8CdC+YDPAh1RDqafgWvjgMmQet0A1yGS5p9iA
8AHLJ2g97l8kOI+2q/xl7TDeyFJuOjIThMW+GQslBgD/238b1/sXpVhqdXbznvT7SSw67KrdqRzT
weBJiPbaso4Fw+NjPV2sb4LRPKi2Y1WVE8Dza0kl2W6E2VKVtbUMtg81/w+hW1IqudgV7kez1A5l
07qUaFDPZLlvVjJhPPSvgbykbwCT9AHo5NAgnOnyMuGc3nJcaEiiiTkPtAcBbcO93N+Jfjc7mXcF
8B9fI5pnAg3g3AMz3KYrA/YTxPYBwEbhcdiL0uq7heI8wAh36sq7ZfQtvc3zh0JCQyfWlYnzSyfo
1NHOewrMkVsHMD0AiQ7anO/DrKWLJ+uAQSRPggKZqawRtXCcXUd/ABhpSQz7yw1INe0iAuyE3pzE
b1qK0iWxFAf4exc8IKZvZRUYgIwrRG2jqvnqqzfEY33h42cpJI0GIldD7wm45RZQDhtXZ7OzL1EC
OcffyPVO38DjuBqqBzGrktOJAs3TcNPamFlGMAGpix2Q9QDw7yXTEGkvr3fbktCqA8hXD2Zl/gvy
cfRWjmyitJPRXTDI6CG7m6xDmdt+FSOxwDsuLPTCs8AJIt/1egyGBVFaWNtj7ahUXSZyd8cP3NIV
SLmg4/VVR3iMZ9+wzYNmF3GrHtC722uWHohM6jotuMSdjaaCpD21hYHjN9lx/bh05NRivHPksYJe
DPLcL6FLkmN2idDNKMVnOjY2T9C3jwVdOmg20RACC2fbh1lxPNDBJ6sgwVXviCMPZ6WPTJidnvNV
M6Ute/au7/Gdn5Atv8W4d+zVRvjLyi3EH2kN+FhOO92yR+9gLIPGsyQdmGEaFhdGgTSdT+bLrda9
NGteGa7NsJ0IEdziVxauSTLpC8lDdTu8fx+IOP5bUqN0qT6BGoqsZWfID06Spatss7mMio8kqTBG
WUlUAedSwPgZdvUPtfBLdnrOWOpt3PKklxTrq5yuybIqKWI2l3oNCWAkw+7JGMx5rC6Zw+8zCq5x
rQ9KP3wumP/CBmApS+wv4a0IhsyUuMYym7KiqboDSh0dIvShBQiRHjVYQ2FAA5zunJ62iz5mbeXe
gZa6kPVZ2GZd6v4wICSJAwQjZv8WovJHBsIubDWzZkzFOi++yLZ87en74LrlN1lXb6t1PijquMN7
boKI1nXh8ExfcyV2KYbi7Hvw4zecLmH8Yu1U89DbexiBNTbndkLE7g/2+v0+4vbl1ALvs2N1nkbq
F1dN2/lFOskiVBQw1ZEwj8m65TOA6MlVYwmvyXwodAo4dPbkxqJuHFJGTQjWrIxRDLP9MdzhcmOV
thoDBWdbd6N0lufxc+fspKhS2Rnp8KsbK9pI/dQI0uU9x/uKqpbL8sou3lQWtSv14AwkwBFNBTpu
mQMFgx/pG4bKjX4YmHu1PxQHQSL0ZNzaNeT2p23LAUw49UcDCBUSSZTQrupzQ6Goc1GTESCSMZkc
zkDvusdjn6QCNsP6ap9Cd1M4lFYh+gQCsc7MXp89Lj/M3hX8w7Qx6sUjFh2CBhILFTT2oaxNcwK+
94jt270vuNj3J+ST3ACkMKI8pxAofW7N9lYeGOfmGaUHzFck3c5KB+Lzizpa6kuhXx0VPoY3Gfl/
9K8PuHu6pGdNTM/P+fqx7NlIrFiszFdGb2AsEXfWnrBefHXIRecyAc8TS1ADxKcAeEDDRHGAHO6d
O/fLh1MT+5nbg/QssDmILqDvrzL8SsWRszwawqHDWNCGVHB2xp73aXZO3M1C+o5v011GESp2AnjX
54J5ZP5S8kpGSuSEcoJu8O+XE+Pqn9yurezLWKpo60Mqd4kDn+cQeZd8/k3yr97jIzs8oigb1nvE
pREzsU+SXn5txgIPtJHlwq6XO2jpYTWCuO9D9WYR5Hp1EeA7uiIoOIiooMY0mGmfoFqnl5jLvkAl
58lkET39SSAAdpEogynQXHDMTwzgIt6wDqmsDGDrQyCRKxgYZPdDb3iVqqUy2PIUzO/LXguoISSx
Vox0BAqyBH15BPGZjhfbiOjNQpbf7VEhxq+7uLo8/QRAs8eSsIFqNxRyxM4Dyu0BM9R/ImMamlza
ATSoXK3IQmmLWNaNz9Hsox3Fn0DtAYp0NM5u/8gmZlsDC/VSwL16HChzWq0gqk/Ty5okBVBQZUGK
olfAMrx5HOpPPCf0P+h7ZB+/oq2zp0c0fIuIwU161cl6JHVuXp93r0bB2M9jyFWGLo6RDtaM+XjF
nrq7twY2rNbkZmiMWbwnJvrCuvV+JrDMkZFJFyjfkpgvGKurDGBSrO3p8NSTZS3kyfSHKPf+v1j0
9sZbWqqOMDUojprAbYQsnLj6v64dkIlzUKzsgKagGS2BGnthgEmypXo5tcHQe0wpaMk+NhLVSHmt
BGxz+QHj/DGbW4P2WMIWZpZcnSgq1JhcxnGm+FUX5f2PlzJVCTwYivLv3mhm2BGt7hCyI82cmrLw
fZZPkhX1y8ZbwB6D87s0JeftMN3NFK7D8yVLFWU2qNV4fJMjEqfe+rZxsOW0gBhTSozrFAQsQzK+
U+ZUODyDIgmg0vj0gOfvFS+nKwgShvHYUJCEn/dfHnhRHel9q+7QxQKnGyJRYsNZxEwPhiXsS7nc
XZ7lxOyPLCwRXaIPJIC+CJzSen2tIzHBh7hV/NLvhqDMYw8mX0YSGWrTCZL9XguuJtuglnApycKl
yUt6M6SV6M+DVuKrkNfl8gII2VPsw3405R+ZrIcVxccC0MEDNjdixy2pABZqQXC1RyAPuomwZZ+t
2Mh9FbNwuwzLAg4I58TOfKrC6y9FNkj28Et4XBok9VCJjcEntmI04oRITmsrd/8JTOWICAtNOH14
BpWNq9fD4dB1aooW6+lzfeR+1PKof/32jblQAFzCbc+pyVRlBl8Q8hprL29Zee/0Htw/SrrYSiKJ
LzTIYf8zF9TlBu7mIDEl9EfwsntAGxxmUcW8qEu+fdWzXe30/G3m19/ShBf+LOdbTHYq8/jYCpfu
48balhSoT0gnsAhJKttbIl+VTOvNSj8dbMvreiMemYS9Oe8kSa0nkZLBlyPgE9gpie1wHIkziTXo
+1KKBUdlgv+S0FDEeonmdXzZE6nNK0YAtawo1vErLYwIMuAgp/M/aEka/jbuBE/dEpdwQ44QZvql
bpQQy0U1I7nOV18eD2l50oOI8S5VMwEb0SY5JcH57OCp3vPGhuEn5a/F3Z2Go+I9Hdc1CB/cd21n
+EWE1tg6LtmQ8zBMSO9YQUa9Xk2/15UL+dYWmq1TzTlkeYhyc7M84UhaUCiSFOlBSkz99ATVyUQz
xvUcKHK2iGX/PrY9elvPQt5vgYyJVb1wom3Vb51bH4tv2laZ4n24bSQ4SvBVcjWzd/4tDjEbHBM5
UGmxjoy7Zvm3mE92i4CgECB85bVCU9Do3+lyXZ1ejJhj9/ai1AfxYXCJsOfywvgy4Er3axfAm47x
5ji7I7Ej6ssp/cXLsWxRZ8ATyIpAqHYNnmo/Bvj6xJ0JBiSZB5eqDQTdMU36aVdbuy9F5QxScKQh
zJRnpVo8uJ15clJvMHzrTfFBEPEd8uXc2Pefk2Man3d6P492gHR3igqQoyYOCfVbd2p1o5di8Bcf
dVYVXpQ0Gr7vyOaUQFV6veKkzANpjS0ixXVYk4KGBoLT1lCi3fa/KSe7kvA70vmyErVA5bd8Za0I
S/k1MnyRW4/0FtjPFjipFlVFS5ykV/Wsd8nn4cSJEpLSQwshi4DSAxXveRv4pK7Tl30XxuIfi6LE
cgIAcrT6ga0oFKOGa6UnKPvAOcKyl2LZpHF4xncWhGfdJrxwqygFLr3bj74H+wPBRPahisZsI1Vr
jGkx7BbsLLOYkT0huYZw2GoykODGMTaY2pPg+dRLXAeEpdWSaa/VNY9xHE9R/LVU/lsQjcowjt5S
A+njEByxcA1AsYA6nY4meHub9FQuKkVDv+k/MwiqhYj9njqMQ+rdy5LIdKT4SI1NnGQEhja2lh1z
uvkJ4ACz6tGgFNgvuNblpUxpENefRaNIMjGoXqKviPN8HK7iH5FyJ0LdAynGcWLbF/70UedClMGz
LjkhCPC7UyZV//Dc9uRxyeWNL0W0uA+uuDdVkcbtszMEd0IVaeATRunQEtnX1vCX64esjQjIa6BT
hxv1ag3s6P1nQvu+ZnyCd6/okP+JWDw1SdRXZ3ktSjzlkHqAs61GfMAeCb8JJuEO6Z9Av+2A0k/K
dLPgv+jqMUlQNlyRVhRgQi3edBpaNUkipRSqMSRo9AO1DLm/fZdJcxwC0zsOvavntDhIKLLkiX8T
dCLY8oDsHws4ESctaaAMbri1bpAXZsebTDQC02IDhE+n1m1FPhMJjSNYpsL2O8u9gjA28tVv2B9a
dHLcB1PmXLOyt/2X0fvoTjzEEjOqxLi1hihCr3PJo6OgY3NcdQvS1VszSQiWEwq+EuE8X/rLj3qk
gOA/MBzSuQo8KwLx5MfgIX8/8p7xBXyrWHfHW6FEice7x9Qh8qjKJuhx9PN3bImJ5Jk/NHmDopXn
oDEiguytF8KouvJiBpBLAuPWTTrq0KsrDLkX5Jqbrc7ZYYaBPC4T3yLj2Pc/N51At1ulYo0qo4ak
4DNwlPDGbhoBA6ip7mk20K6omAL27qINE92/jCSm5PV8an6CuvY/9j6qxyG8kfjYBZ7tp63+2Lhe
cwYLM+IR3nGiqp0zfjBJD5sIg2wuu2CDWfD5wWkxz25szhwEKwm7Tr4hyTA35TsukoBkHixr6Q0X
DwsaCm9n+KXNmJfVgnoXJo2kQjJVBxv3MJ2vg6WFYmE9GAHyzCmtSzKxOS966CExPpjhso8wQE/8
6IluOBVum32mvYeLO0Ppqc7ad0tGH7UFnmDmvWKD5vlYUgWKervDGcgG4PfuYGrorlIAxlNl85BT
m1eFoKK33BbWdD2b1qEEVBZMq/yEvv6oqu2NxLextkYml52Sxpp/SlwghRt5gPaDnchcRbU5e3rd
2TosagSKxex0Lu4DJs+sKQ8ftiun0ypkRUDdnbGkyEG62L0PR5GL4XCtKVb0syrhbsNg8hy8Fhd2
ZZ2Dps0wE1ADcdHYDmXwi5MUiRE9oZThss5g5Yyb18dj4A4hXXhSOEE/M7R9+2L1UAIo7cLc67rl
cZ+GuTeh9e66hNAePLluLHW3hTVpnfPas07MlLFenvSZjOx5y1K0VAFryxVH4FX1PAVcI96zFsJV
so7HC3yefq2gdvyv1HA/1tjsHQ6uT7vW5i12EdZbRpjSWJZ2Xid94Nm6SBs00lt3FDX9yKEYtcpw
y1HJuyFU6gdsGT1TQH2OCiXk0zImpALnbobpWom/DsaYXeK5+/wMeqjYoJqcaH8tChqXR6Lp4KDZ
gL4Ei5tfG+v9dAL+EzoT3hW5jbj4BBDpRxvQnUtaFeghy+qogoT0kpII6HPH5SOtbNxN2mMw4LaE
0UmIP3lXhBGlYzB09DN//YpMMalRhKF/OU7HHrOe0ZaHM9ywGBTK4f9XQmhBbIV50pRHxv0CY3kQ
MsKfk+PtXYkkJfYOvIK1RRgi0pXPuWZ+4hmrXKMNhfNT7KvPz3liJPupg7HHAlewYBbr++uRqRLf
/uQrKiT6vtflN4/y2TxFP76yGG+1Nex2qrNGoo1XfxPmy+qHruhLtEoFGeN426mbUsFnhQC1ZcdP
BiMF/RuHT0PaUEblM/zO76xRAZ4ovsaWbLMZ7+D00ujngHQ2hCU99SjgmwFmuoKA8SdtEWTwQNTc
rEBGd4IwH5BnvKuOSAFLAOkFw88gI9XsRzCF8n40WaHNuuuDOukDq8efyFNYMEvaye+29n673M+M
VLwd0NcrBIF2smCc84sMrHaxjXzdbl/xqR+a1ptthbFe2MLXf1ddHranUGqpYlBnFKlrSh0fo575
LUQihTzvcEIJtBB2WGKSY8FyUbmwM6qZWOR7uD4i77Cb/k6wfY9BWx54nWUcMxg5Idk5MgKiuqfX
rFXBc6aVjHRUxHanNRKn7jvTo0Np6bRanQC7kDZ/FwbemL4jh0DDVunCLHeHuzfIickM7VTYWScj
hfab0Hub8hwDNNQgDaDO0ClLKfBdjR9psFtFaX50k9BsTZ+4Z3sCEj1SkcU37CE6FkvxqEySGjvK
P1fQ3YwBFNtK/z2K1P9TNYr9xD+2s4oFWpNWdtmcyC5LNsmOyvRvRmdZAjearEkhj0tlYCd9GIjM
nXhrP1DaoUaiX26+rhpvbcwhCh1BopldnnDtxUU+eGn8MM3B1IRrrD663Vm+Ll7ve/dOw8s/RKeH
vIhhJbksKw1xElXpwJiGN07NtLKld/xjrEZ6s9d5mJMrVqvIVQ85undElVXN/THhrJtumAy+DG9q
qByskESq7hLUTmRMdCSkBb1WKbK8eQ9xKRL/o7Iq2leqUOCvx9E03SQ4oJKcLsFVqpw0A8XHhRrD
GpRd8rGvkB7n9PIxYPbWqbdJ1SRX9uQjAepB1P1uvNfVJheoO3uKv3I+GA6tENNfX0dsbbKjcqO2
uQVEMoiinR6WJIEz9alRKFaP1klUYVxLJ32Z1xyFY0J8sm0oOBhlTUoOCBqUCYQIVCCcf+pdnS1V
gTfVH/S52kUGOhTITdnKTttEh+9fBLqAW5do9QPGFswp12obrKc7IbWW8ilUnzklA68wzdddcjC/
BEPxeV0GA4xvXiISCuiQDnjqqs7hg5gAUQ2fO2Jud7L2R7TCfYeT/t/arkIQuRK0z9z/JjmbIpye
0UAhkzSIFO0NkTS8fO0h87cbRpf14U37uFDVkeXWTla6iBBy1G91Lws3BZnXLNlrKF7YvbnZaeOE
V8/XUADeUoqzVGoPBoQoVdSzArmqVNWPfy7cE+OI18kOt7kS/UugTiKxZ8ow89DQERK95qz9aQV3
/ln1huQkVGcrHUBpeh/Y3w6Is9Oi2hXNe1MH7+5A/Blz24jVxRxEkueyu/2+r7EQHS39y3W/lKjm
COHAnarOVu8NtNj1h8gk7AObWcOTTAE43HDGezwMOWwg2xYwdpig65KRNe8xyXywV59gETfkGQQ2
pMxIDDWtRbGOQ9CtSBjZsgHEN6ddNy/rFMVQGEVjgWFpRNOkXoYWpIkqZNzcclEh+h8bJhrdIyfR
xGiivvs+67DchVIWjhiuQusXRycw8MloXKh7Zlge/73CZXvNlCNXx7NoB6zCoduCbMdzW3cYFz9i
2jZEQ23g7HgWaqaTIdBhU/VXfReonVVUKZ5AhELfhyDrYKOcc6n+UJ5ebjpo2DOzYcFUXeotYgi9
BSPlyNQuRZr1juvdI4eYob3/0ew5WNmT9ZCP3/vAsQZzCQdoC3s5vyErHOrQMxT9VEItTMVAjbai
C1wjDdX8ViAHUt4ru4Qfg4YDvFZ9JZxtu/4/HulvAPy0WR704Tt6TymQ0I+SkWj9Idz971PpB4c+
QJpWcpnGrR0ZxqLCAtQ1DURxWVXOtJbSICBlgA+nx7O12rzLHvuQs35Re9ea0BmUCA9qInHgu/8b
LNyCUZ85OUpAzfb7cFixciVaK7icaoUwPYRVCY3ZM24wq72FnVdhDndUlT8zkcDj6XWk+AlQbWus
R6OSPWbBQ3+Bz/wWrTwyf2C8Y3WBY99gWMTmxRAkcO/0OvrKeFGUZpXJK4q4TXf+Le+PGGVYyoD1
UbiQFn+kLCxG4K4PBS9f88GGFhSPeVIHZvn0Q9st0I7npPSKSiuRhcnX48acKbAcGA0/4y74KPvu
je1NhaRn6aV1ZZVBLaMcVtI1Kl26cK6YBBlOVyyyoe9aOEdnMDxNpYacqXCfrtkagdkiZ+G9L5Pi
hciNRd4xZZWHUCYn948w4Ji+npvBO7VF132ekx9uZWfNLBJ3S37u2uRf1T4ob0GaYWzZvotHDu3X
dpbt6lA3lFmU61yAZLaiI4ym7CsrRp4T6HF0suHvmK/N6p7JfgKldNogFN2LNbgCTndprv7Gf7fY
jJR47Jubp7A0DHdjvbIYwLcDZW2UghfvXYLAupateL2mSYNC5ZeTvIm/yqQkBYNQBwC5TP3vjbUF
QdBB9b4s4OMMmLR2HYVQXdhM5iNgY/xCSMcPn45Nn+y2lr13W2IN+Ap4FLBcRlkgOSVSi4GIOqcX
ARNGsKXabz9MQ4r/3chxJosMlFkzqfKStyAbRfIprl72Ch4rW+Utd3iVLVSdEBqf/6f0Cmz187WJ
3FuH66dV9TJEU9PM2kHcbT6a0YIjViRgmV9abRX+mn6jKhAATaW5h/5zE1goegeEJbwVzkNs9QIn
BlaMIQbjJAKG3v28eyNiKoLwvVFXNntuw9mheUkaWZ6RqcUikWzdMEtF3VEyiAwt06T/b0zdUgUv
wP1M5itU/KNg2ZDTSf4DX8pYmMsb8q/Q4AIITO4mHK0yTQYKMM4W19OPabIqeNeqDlU/YecC/Nbl
bL7S6VXWGQP9Vihd/K66W5mh9vXAMc/3PQylkzgqCVhm7lQDUIVshUS49AoTSbnHdUFezZokrQcv
mOr/pu5fBly0CyKn3sdsofFK6/IULCDchxMh3pAJLC4X4CBkrcje1NnbttIDF5IZEEhdLYNzbu7N
MtSk/mYOpauIUyprpDxbdYH4xRWmVv86x4Lsd6reCPqwWfaZ2d/pP6pCaTOiesr47xyu5wD8qtmX
aepg9w/Aulpvjd6slWDQOlOHARwbl+26eQQVFldYw5Y3ldme/yx9y2dNn3BSprd3gr1uubTttwhr
tPQpQIYLUt//I+Gw3HE8p4rO+AqifG5KRhISPTOJ9SW4fsXwLprt0a2WbZqmWaCAQtpP7XHW/wvp
FkU5M58s2UGa01cflpu0VZj9zsWVOkhY5Gkbbj5RBq/BgY5MKjX9r5Kss3uI9hSuoeqHkkqMY7xY
huEIwNwjFvih/qnT5kQ5x+sqG6g883RFiOtmdrEvSWjjkrxvZDv3d1qhnv1BOexj+SZ5JQwOnYwc
YHE6K2pSxVcbPuRRX4+72RdYZ6QGq2w+BA25N7nUUbg8eJr1dPLAJA7LhZg5PZFCwpzXpiI9XJGe
ZKy+2Luy/kQJk8FC/d7wa51QkTw/pqmOIE0mN9VuTJawhxh/2KZ854ZCK6eTp/Ad28JU5ZLWKCQm
OhdC6aXSiAEG1NE9djWhZlhpSTkWbO+rmtR0kLUvHw7pS84jU86QptQG2IcCxsLBTfoJk3trEdT0
FwUSZa8c++FuxPsDuh9hu2FgZmDqP4VEFT7faLHJER5m+wM+p9Uvt4XbwoS7bqzoppqWU61ZKA5I
4YEswPQurqU3W0ZTlUczctQ9gHykhwEyXDkL4ZaVHOx0Gq0kk6VRpIwQP+cs//KLSzD8NI3Gkpsm
X4lGMIlV/mdv5/FusLSt3mzuxEKitbDidxnoC1Qv3KxT7quLIxr9U8++c0R7zWtzRpmo+mPForVB
S1O7IR0DCmucm1VsUTuS5Iljwln8cT+5CbrsNnNcffmmmJTcN2o2kdGaCzMoyzLdVnwB++ZFsghB
ZFIRrf01AaFyh45TTemXTHcdAyTYQ+1qL+ppU0xCYiRTxI4ORV1UBDSQ0oXdQOudCemqIN30ztOc
OAYfF0Rmqsu3Zjh5P60r6PkH/yydKCm8SScgBJvtrx9rFdE1YLWC1agwYjNfpHNJsxjueknivxhy
sPxSMp9gmNtt7BGOfGjyigz97PWImfYkMpBKiFyUAbYjep1y9lVpQPO6/meoBRl6DkHkKDWm7gZZ
CAJLi1Po2jeUKclHwgT/wg5/hAQ00fFV4QsYII/WxguZt0oKkeHQp1iegeXedXMcgUVpL+RDnbsS
c3fsGwQbRRbTrdW/ajVMP3ymD6gaX0+45ZCxpRU6+jHnSMsBRel5NEferSU0bmmMw7+YkvnyjHZd
u9f03A7FpgmFrxQHeeV7znvkFwc4EcCy1QMN1GfzkUu9RL+pK8Yrhw+hL0XxxcSvUHfm32TEQUAV
K8CPMCznmHmQh5aervskd5YAXW60HU8vd0CABsbnXuFhV9jkDHwlHvhZhW4K3zPUpotWqSgaARr9
DdbMWgl0zyAGk096FMd04SJThdgTgpaYBsa804lnW6uaxR9VIuc94Y5rFaFXEVgdDMu3byCprLXj
5+z7F2yrfgW/Mg8LcWHZLeiyvG1RkFLxc6tlx3wNEpH45OK/Bp1uW/X9FvrjkOFjS+wlMhsWNKz0
+6iwVlGjrezZXgHDuk4Mde0OCKG0xFtN5dYmlsTBH9GuF/ZMGEhmP6A0SgCHXRgwuCmdL8VnPKDF
PH+r+W7mHMrftEIaY28l74eN7vx9BZNeM/rkAtpZsES9TJjowIjZysByby4l20+7iyDGzfodDfEn
Kv6ttWciq1yJhef9H7FiH3+ABzzqy0LABoqZnl36mBqXVm4Z66LvQv/h2rllAf0bqD1q++VuTTGZ
spSCfmeCOhvFmVqz080/WlgGKFNqEH73oxM+26gPvnmad0vOgoFs/C7xCIVcwUOTC5xWErn6hJvL
0pGSLNBBnabmYLTgDTTKI1T8Cl7HGkSsgUJWngcBUgt777q6AC+9Lrlj03pwuZDs6C7dWTeVP3NJ
arNsCRwy4NvwmH5Reigl2H1LbaSBOwlxTQh51klZ51doRtUDH1Nl9xWB37DdmY7w/eEJnhHnfkwh
rNmgdaXsg/fJ0tI7zq0sDM5z/F7Iy5UtpwmXxjSZdurNHjYlIYqsX4z3JmD3XHZpPzFgH6i863NB
O7hLyyPe/n2bvPEXsELCZqxXdpi3+H3f/L1Zkh8+U1EP+xuPTQoLtzDbgYY6g62bPzQXPcYjI3fd
M8qWHc5OmZrHYqw7kKm/MrQhb6T3NpOglWbfMiNs3dgRguhi3re1WpnIe7U4osSIrbHcqixSmzax
W+5R8F6SUN7c926G/fD/Ky2t1P/BBN/zd0BbWGv4vBf9cRs59ynzIvuCGMarxGW5DctZKtfiO2sT
vH2WOklnflKyRlx3Vizj+v0JQbTp9OYnFHO8rKTmFQgwQZWsu+Qw+k9xzGaZbFVYD/utUw1Q+NOg
sXhharw4rY0hCZM8U9Gg5/U36Qp0b6eD32uLSaCAgY7vY4i5E3cDBS6xIO/I+b3Rjm4ow68sQySl
ze6Br9qcMTxmPpCY+uggVmvS0bVHoNwkUP357QPVcTGaoRAit0vfQjiLSfJ1YVueUZYoimLTLQPA
fNyxETzOmE9ybBf1F6chf2Y/FQPwPDdpFALhzxPzMfRZpGAKLK1PSyo9DeLnUd2KpzKyzRrM5DXc
tzHv4s5eCE1Qk4XMntUiuUKv0OrD0BDtH3AgBcyUW57dh8Bt1lun5AmC4kQMRH2a5m+eRTcZl/rG
R8oITbI2OBXin930AnSH8N8lHjbiC+QpbCrMUpdH2WmVAzwgv4SapJEbZ5mymIAVhdiUeA5bYiqs
BreQp25n0bb78ezRPCue83N4XN80eoPeFXnw2xL+wj9GeV/5MOLF47RHAar82ccx4Jg46JdeoE3P
Fyv1z0UPLUlyb/gEisFvP/VuQbJ0JZZaEcj4dzA4cAQJksIku11EJVIAGKeBIm/BJY84QP4reyiB
5eClj4pUNDMvo8estalgv5/aJY7sg2BOivCcRShSgbS+LRzVSJpvqMnlwNg2OoCSBhDSmPwCiqeO
ObRV1mwQw6DMA5SgiXqkdEay4T4QJtTrEv5602/zgZPhPdH7gOf4Pm6kx3mF/0AtzWR/p8XjCjNS
lrwcbg0dVXkzF4I3UpKOCef6xXttDK6z3r5O8csFOvE0NMzMMrAe/XNdUd9hsRbxrgeyulwdBvN6
9YfwXHHU+l/ugNFBOJe/wkrrw6S/VRLbR5obdWZRaBITE8g2LIFiGOzBqOq6Nnu5lcPVfKx2zKNP
4cxsR+thHPEHxtO6l7H0gXnWbWQGzxM2JmpdBXvzGJxkil3O/pN/Ih5fSdnoBd4foYktg3xuS21x
8tTcXqs3IooOS4798+vdwbQh9AtjxgzsSxh0u4LD0O4EvcP/mc8Z9H+TSV0cuvxlPdynzMS1j3ov
oqS6TzxVK5ORd8eOol8eoQTIWZ3HUXfVjMoAe1kvO+NN7Xa1fsoPsNOdnPcjZ/SF0kEb0W4vHorM
PULlSPffkr+vNL7+3JkUauo9mRLwGmgKiFihG3Ca/euPhR8Og2A3pQK+rlBSfNzeWoRIPGttg7fL
JNgXu5A0jlSgLAyHTC5p43OoCSVgXzWDzzhKqaEa8oDRwlFo2Eo6nPGKOsyCm6rAjVRE1ylSQPcI
rBnKs8xLh7KYfeYOvBKc1ZUYAZ6gdeOdqpNGadNgUjTvvEXeDdwS0X3IUmWxBSxvVBOsdk6D6sNi
A/roWag6GrdecA4Zt9jtzzcIpVlXu42iIro+7CrwO6fwKLiwcWGTt3lvY6udup8tXjLMm6UEImXW
uPEirEIqtqHRPTeI8KwUfodUMaWotGWi3jvu4BwLl7ShMqBb2xnG0AWr6c4M21+xEzlwmGJNHjFT
PRU/n626lpnLwLc5mMbfcpIV4M1fgTFmCPZEkrFEkCDI9GqF6pvbdFeBlVRYc4QKq2fTiUsyS7H3
cDDYVzWQTrDh88DdsnrKTL1g+43v0TESQj3MIBl0wQFib3WCAPQikl2tTSkpB0c6/EKfhnOG9exB
/1qiiqD/670xnWwIUvXfTV+Jmo7Db1IHt53eWUUXIuG2zw8fm6XK7qbQjZSLov0hTHB7E7urJm/U
GeCEozGUElyTqMgobhZpt7d/c52zeWQ1MFgBfeobt0nKPRJX7/lscLfYxS6QZNJXH2TOOqCFPnrV
JKSvuphFxa25yq0EerNZ54vWYX9Ezywf8QTJNH568mXA4SYZ+bMue6pjT2ayXItwwO/wg+FCtf/8
untdfyyBcaKsEZmewz52de4gECcwakoO7Ci9pj1WHo0Gr+v9DWcJsAh/pRzh1xIQNSm7ibN/l94j
vwIWYydDFTJMUYkotAnK45SsIBbzov/eGYYXfzVgUszRus2HGMQBiVWh6ToS6/A66meV6h7vahWR
Cw2eEq5+PNLsbtO1VsEYfFguajd8k/B6n74MxbQrX1K82e77Cip8L6ReJ7YcYaEOJvhReHFWIeQh
0aGAnnsNGImc5It4vnHP/ClX+XddPTHYBusb+CT2uA+jTUDx91IGg0qdnPfazNi9v60+gbw+Gt9m
7UJwoSfvwvlB7PG4Bfafoh/bx8L5sJUp6VWtW2TgJMOiSEsaI7luEQrLa5mmIgp0CnXThuVTde3f
A4gKD6A5CnNcrNTMcYjafZpMrzc9L66Q0BCxAr4Drhbm10dml4nF5ODtz04KIXibpU9lzQai6Kfq
keSi3RvwiudhFaA1ngipLk3rKOWPzDN2iX2t2zR6xHV/Cioyd36l9HfjTUyass8e1j0Pe7458khB
kV91PLdURuPdsWUPDOYeGtPEhnFzApSxWnNJeytJqBACzW6gd13ZvUbkDQZJ9abL6nnlhxgqNlKB
oMweWEMU3MQim0BNJRvULvBsX10YsOdV+BUfqoErWkes+43vCYdq/mnNndt9tDZvUQ01tpmBrFje
O4Dw343XqyXqPEHd6fgplflHo2FWcreJP65t1ky1AIljV7VLSOnVipyRSFU1QeS1GBpCuktnzSqz
7FGOC5u7Af9VLcLKY29NXXzmxHwiBrimycKLKJCx3+9bq8pXP60raAdHPYRtIHXt2eRgPsUojT7w
jdq8PXENP8p+g/UooZQRljAmz3R/iukWETvrYq/2qsaoAEfos5DnS3YNL7ebMOr8afwWnwUJ9ADX
mxVprygaZMCYRIpDbq6r0WlIbloN/OsYdxE7x7RyKe1t2p+V4B/CVZW+odmBRCo0qzw+/NovkzHN
X6xxXA/k9cbot4zyl1gYTdnowHl1aKrFGCL76tHytXjuxSAcOx3sHf8NgDEhaKvQ9TxTpI+E8isQ
VoYRSiJk4QdH4Xa7Vus5oNekh2i5FLH/EbHcNbxRO8IT2XVUBwuJ6/aYv2D6677FpkWWNUh5iPQZ
oata/yfSXPR8P1/rEhIx2aM80U3Kor8NiyDWcGhP/G+mNCgcvcOL/KfEEk8bw63UzApVZLvPJleI
5JnG5NXmmNrTSHQ4DIndeYLtDmAVy7pfC1gemc1iU5zUCYgC+wFwAqK2jXEL3IEvMp0OvsVutmOi
USYaB0XD6rRmEpzxdCtNEkTzMqWVKzxTNPXJnyXJQgggfq+rtmEg+sFRzzUeQMcZhM0PaLSwQo0/
Yzw01tTxbCK1RzxJVmUAvdWiqmt1Nq26OceAKkiK8pvw0s4h0pqYPh0ZTk0EUt5IIinRsFAfbt3P
8DVWrDjFfxSV7b11rlJ7PIccvFeanilf8kMAHbdQyo0mhag5bAvRbrJ+U8I3EUkgn6B9LnBzlpop
o941D918u6yxsL5aaR4O4SVRen4n9+3ErwvPzcKnOZr0zNkEvnKhvVcEz0wn4EeHUqxWb98AXhkP
frae4e3Vi1TaYFkx3fOkDKcTWKX6HfT7MFa6X15eYlVNnLfMpK86E9/K66rqQUcx8Q1PvqdPcWJd
Iy1PmyyD59WBaWgW2i3+8aZCfN1B7bab3FNUteR2FUNqZKSvDQGq5lljf5NMP4v3Z39ZyNP6+OPv
n+2e2z6u5OcwzV440/HiU3SBCRSrt9lAkZnfZBXvlgAE+jtfrXmt/sXh0r9x4FlkWAvreo1mbFBE
vgrj1MbjpspMGbw2TXKQf+DjRAU+Z7uGTY2hFU/GF0aey/eAB4G4VUHcnq23wzf9rEvccmi0qqwn
Lu8s8LOmJLnKWNIpQvjgjaXQ9PyMCsh2GNA9kj7C/t0hTXDSvmf9VIcnoHJBSqGQvyD7uXXTH//P
on6Uv/jIcH3WL0PXa1ETjqVmFL4EcTESka10WSwR3x0rx2vvnwUbEDwP6aH91q6y4Th/4bPA9inn
Zvu1Pvfi1bhcHqf326qFIugcEGlJMQaUQ2GtetF3wpzORWMXP7rbTHp+QQf/EihLv7eiPfytUHq8
CHqk2zyh69EGq+Wi7RVci8WRF0ECFjFf5j4kw8QyRVKnym0Z5cNU/pA999d7i5WYR2Xoctmgqmy1
lwChfeP6BmGKXYUkRbI0uwu2Kart8MesrQdAsup3rA5zmx6IAQnkJEQBb3LQQcaF4597QyJjQ5R0
c//z5BvLgOn5gBlkE+Inquzft/NhKAc3VX/SEZ2yfA5cw/ZyAWQ2H9LxqO8TV5M1jr5J2hHs9e/f
1hRp9+MWDIBDRWxrTLCJjnmiRNRYtN8/ti5YCR7D+Mkx2EAlYZ/vZBPbqwZNgwh+i9CyuyiIHfvF
sY6SHY8UPuVYX2c1OnCKBbmVjday4XSeepAN8z7ANiMQFDgzFsqIiXci3c2irWM25ReWQvQj/X7Z
JWEx8JhQcHEmu0juFx1BNrU+XqRPMNGHsluM4APhoCCBIQ55NahqDmftAUFO73LXi8ipa59NJ/VC
oXkKvY1msUHvC41VV2BHjKrZg9CS20ktc/2UEPnq56xkJBHRnsLzBMZPl+lXWNRbipHKy15xgcQi
Lpw/CCK9OPDfsT3p+TH4/RbTvhcbNrxZnMJ4bM/+xB1jrLHT9I2I74KHD81A02jjeaega364aonJ
BJiVBCqHx0d4D2dXvoPP2z9iexDJxaac9ApIsh0/4des4L7ZY6IIoAEx4bcQkTrSRlA5IsJA4saI
HtImGDoyiRJmZyWec4nF7JkFxKVp/7nGyJl7LMN8iFEYkjm/4mpJy006/J18JmkwKIb10Uld1D9V
95XMnzMGWPEj8pJRsoOeoee+MAsp6z/axZPRkEiT7h+COihpYJfP2wcUb32IndGApKQw4Vb3vl7e
fOuY5zNfpQ8weSU67FG3FIONOTSpDjJq6eQ6siZ/Ri8R2TBQdxw8FRjb94F2Ik4oxBCnlI5k3pg/
eUNPskD9ckKE6Y5PP9mrZZ6US0fDsedidrpz6g1QW9/5uWdT8HZykzP5DBoTkSP2qo9r0imivwZX
ZkrA/y7LQA3EnOD3J52h399yCldNDwSHIKGjSE+XbYjnIaundjq+pkYh64zJ5oW9vNzI+LpifjLn
jNGNcI/Mebw7dXbNwgogy1HDAJ11eitBgCo7WC3PNN96Xo67buHrXuBs3xu2q6bB7/+hM5ZxisMm
iZDPQerN7e4Y4EeMCPX7vc8e/tKU77k0bqSBpTuCh0jd1rcyaUE7qtv2+HXSxA9JXca5goOLNApc
n1jskmM5k+ovUMTs8mgC+U6QaJfqEVioindF/JT9RAr2xuyHuK6Ied26U9ep3tJJH3Hi13D2lww5
VoJimN81rYWsSIC/7o4cEXNNsz34cbg3bCLB2qgXRv5H9m9p4+XH9ZuackUAA8JMySh78kUI80Km
5QJPPkiq5IMde9V1DVwS/Lp7aee0R39gan5T56cBJK/UEkx4df8kpu+dDKsjSSRwiG4L/KGShkmm
8Ur/2v0fkLZ4tCpuysw0uBVpcI5RuEqTrFAnUbi7ZELnM0U2bz9t7n1VhEDcTylLHIcfcSKAlzUs
zBrx3lXh+sdjijjLN1i/BK9zLmxJMdwxMutYB9X+tp9YyMJjbKBAj5v5FC8TetLZQ1n/4DHwGcw/
WWa1aC7L4sscI2ucWQmANxJBA7BnDSh8quvP/HSE6pcUYzKmwme9lQscfKIoQDb9Fc1FnwHpgUnp
byiJdRg4By1KIMnw3/MFY6KoYLRc02bCg7w6Q7ld2d3l0gxZ0N82NgcT1Xzz2vvTjXjOtc9JU90K
WiBRVIR/KiLuTPpi0bRpMYae2ibXguhEJwlH+I7WHHNspF8Kydl8UKqIpS3m9xMk7xECVEjivC++
LUSj5Ba3S8z8UsYAF18lswQMf7HwnjfPvg1CDjmF1ETfqXaYaX8WHSKBUY1/+XN5KXB97y/iQsyO
wtjfRSt5QZaKfR4ljIdQ037nfjdbKrSuT+ba3kaLOGAuSJD8w6HSPuzoo6bzPat4ZiM+RDcQ5lAB
SuNa/PZqnQrItYQLt6HHO7io5jtllUywHj5qUXdB5YrJp4prRIR33lW1C6CbuZ6o7NySJ6P17JUB
fNTyAHn6mq4Kd0W51B+2mm2gzZrlrLO7A3+a/0Yh2DvPWfGBAtEfttA1UjVv1jsDGhTtrYrCcSE1
iH2gbjT6eUm3CweXhlr9wORt3OIToHE1MBGaj1ISC54OcQY5/NX0yr/xYsm8m595ATg2lbLRCRbu
4An+a9TayRSPSICbJZElca6L4J0P2zbpeesk9kSR329rkVfGdau4bQC6SlujPoDv/0mp/Ifr+qg6
o5EkF7Xn1pBSn4fCZgzgQqomUaTgi5Kbj+VVFMfOR8GkH4zA06hr1YeiP11JYeFwhVVP+J9p7Z5x
oTZfSvuwxlG+i48qm4e1E/FCNBQUSLDg5oNO0qrRHRRbFO44yf+rojCx7bBP0+Y1+X1Rd1P+5FzP
EPgjqlnj44yiksvyv+jIVa0KD8H3I5U8yDecfOG1Dyy+hzq/z2/6WzaOYwwj2Ezsa/w+WQ1A66JM
fr15fIpmlN2r6HrEkeNNNOExT00lDjbuy0QECONhLK9R198tEA5Lh2h8Sn1m//vV9vSXdFOPE/3G
gwEv4RQ5sVpdoN6/x5Cn6FtcUn7dI/QFBXwrw8DL/4P8j1YUq8U8wUDY0M4Tm3w6M6WT4Y9CJCTv
QiFgQrJGJeXjHBzHyZxo37iKhZuz+kRfASld7yP2hEGl+/f+LRUm3h+uGT8DGBp0i337yqT3Vuv4
QsdyV42GiILj1zLbKSpgC6mjmqAoXolL4lNz5Yti4xGTIbhJ/PfpGYmibe3WkJDEaryvpOv3VX96
NValRXBu0NMBZRUf6OIZ2IdDfn92LJKDcKcJVp8snWvsVUOcpKhlVscVvS237rdjNg5oNm97EBYo
MmQQmphiKvasJgB6kSaIebPMXE69q0rphYuo8TFzp0NXWtsQZAfEikzPLD0AMBzg1KC3hoRQtKXA
KxvGG5TimKVz39PI3C300dYfq7AwePrrvE/bdTXmpP/QF0rDssNxJYOvkp9pZ+1s1ts97Et5yUT8
BSjcxAA/t7BkDlfN46Iii7fThrpMAFOMsfoU8u4Nu1E72qBTVf63Ee3IK/pnn5JOjNb9hJH5viHf
E2kM2UW9D1/eMlOBYWnMxHPhhOceKdv5ldyPs6Kblb81DTkHrBEfTIAKScJK9xYKMYxTD9Rm8zcW
peAXYaD8iw6LE0LSj5Weq624bCJxtas9BikbKty6I+AubKffui7Oe9QlDxqbVGIEjC7LrEVacr+2
HLVfL/n0O9rGhvxplPXODfXHjXKJgxYaFBrJs+80vbUnvNW63lWIj5fCvYm9bUx9c5KFb56V/QG9
arLEya4vw2zcEWCqPXdc+kiZZAIWH9xCiAIWaPaU13tABDobI55XYN59X/RXCdBhzeNHRbhLDjyo
q03/Af0C9pF2SbPsdxNwSx46M0eB/qx/yqD3UP2xvm+3Z8cONzbGqb135G1TWWgkJDL0Ui8+5Hnc
lV9/Bj/ajoXpejhP2aceFP6s3BGZdRWzV/piS3trxCo/riVR4UuxFiHgeaNAVSl7rRJ/K5dRcbTA
tuhbepuNa6DclAjBw0UiB1Rn4bw+lJmJA974O/y54/V8CQsXA5PBxxFvHUG0HgB2Y6bnO8XIBSuN
xQOs81N6NbqQlBHE6ualODJbLtFlFVFXGrfiIYwbQVuVYJrbh+VdlKPgwbjbPVUYgGTI9wa2CvOO
0UuGauDKHp6dDYV31j8AH3N+RguIlR6b09Inqp39eyJ5GFkMuu5XosvWsEbIfao9MdPa8SumgV9e
ncOnjlYnzw8i4oiV4R8W8W9JFsC1FBhCG6gRJfaVy8ZkZ+H5LxW0uO8OnzoMQJ+qsTJ65CHzs7ig
jKYnPZKBrJTxrUCZTM45hidmoABwJzkxqvgbuK5cp3NAts9Yv41ONjc310U+MFkyzirx9d2vqr3f
e4jhxZ4iQhCTKo+jNR5gSaeRH/cBrrDPZ2h9bE2nB3eG4MNCkEHJxFCJzrh5RCTYE6ZtN8gibg5v
ew4PGCGansntYHAuEFo6Ckl8QtNHNG+/YKYhp4dnm7nx3pTQ0tbo0Tk2va2lj8KHzqX//qixKDHZ
HTr/jxwYnLzjTsseDrtkw/LbnzqpTl9TYVguSp5LNpoj1Qn65xDk2mVtG3i5hc9gni3EUWsXlP1X
OnTj6zhBXbrzUBEvr17NTp930xMC+iB3UABHnDp9LC4XF1HZJg1B9K4nuCtuaS6E6I7emV5CEHM6
cEzeonUWy8KqcGbA0YFdsZqnWrfWWBIGddudIEheor9PPQWsyUTo5M+xhsFPlAolWX8KRiirJ/XZ
gSey4S5IbLGedNz43WAQOX5XWgn3sQ5wkiOVHC3U6e6hQzRiJo6bQfBdXrDEzUxXZDzFSnhwGSNd
6U7cYa5b3REnOPFJ81m1JsuVIVrrcnzyFwE5xGMdAe2kSWyFNnAL6ZMAE0A1v1xubbj9v7yHMP4E
5pgDSUs3MjUHdC7aWdJN8g1yfghZfN5mbYQvW8fRNEh6w+4vIQRUE9M9+8wz2tg8ltyMGLWapjds
rkec9ChSj67Q7FBb9nGetOsCYbwmrV3oqm9dHHVJJSRMzKW5034dKdEkh4Mp7ovLUpl3SUl+KMa1
BDl4j0u1A0+Dp93alyQCyl6n5hJ0UpxHpbl8VtC1D2z0CtzTDtI1I6xWS+DDIOwonr9P1x7UXksc
AUxMDMQSxeuO0/cUl4FDW+dyxF/SVQGg9mEZNFqOtuEO3a1npoteV+Mt3jzokv6NDvXS+2SfG65x
2S8sJZmT4+4YpfOsKecBty7W8l+u4boQ/UnjNV6XcVyc6YQ6+TLm/8/1wcuzugBt6x1EzvuPb44w
LGRBV9Vwyk/Qjv4oTmHpCQCUQ3JTngmHkC2WBPO7NZRMmY6gcGX+3lKSvjbAOtxOLYPlkk/KQfwk
l3rbzyUAK5yfWir5HmOQIDtcWp5wHDGt0Qx3k064D7PBF8wDiDxRGb0zPsYOct2pzqqRxPF5fJp8
eYR/aaGAGZv39NgCOb89CUE7Oja5ncIQK28cI0C3gINhsv4+C4Qd+/3s15WdKmSSrdXk9ffHzeOI
rCzB11o5CV7dp41fr8LsXjlW1/elZ49X6HCsU2aJrq7XdM99z46yl87A9S+WssOUJof8qFAweDKv
7G+aS0LsTdM/2yk4J1fBC6SWtniosZz1+5vmCJuEcb5aHAhXtE084W6ZytDPMfqUDKZQ5vIDEGPp
tZwsAIHbnn0dA4bfehPa8ZQjAKTL98ls4eTb+/7QjkI4HO47agf7w4q+94cJtPlMX2dFAnwJIkcJ
vjvUXxSY7awork76ftZS1Q/oDqZ48DxuDr48y173yMFhpkJ99tr1AsgI7lFz3HurXDW7R3FCAGQ5
2oRkTR3xLI92aTahuiitrEW4D21jG1QNtZfUm7dEeX2jKz7S7Kkt/ckYyaLRXEmmCfik/8hOpBmS
B3ieAM6MqQfBFA8+49bzmaxq1Y6JrSEZY9qDCKY9OE+iO7/Hi6ov1xOqcXVFH8AbPJ+UFogLeP+C
PLhNu4mNE22CvbGIVxv9MPuGPfKiI43UzFmm7wE5noxFMhMpMDAMpl7UbCBuw2+znGucruyn3SeC
X+5yKp7j3GKSIkPxZJWNdKCF85rCnki2Xxt6OZUBt5PskCTumniaTFYVPT9J/8jaFQJ8/BTt5W6a
etc8tLMJQ2pAcnyy8L4GXxY4SwsgM5Zl4uXk3bOiED4RKbMxOn8rRTWXb5phdAE6aZiZmAfRQal+
s6uz8Wo+Z4Rwe07J377HY1ut8GFma7GtEFtkxmqD+K0mPk8gmNdVfNL/X8WqynoqkCN++QqC/Tds
ijb4EJTbUALcjvATk/LFjCSJGHn5fxE/wDcgWMCT/JqEhZU1vjuFUkPEZcPr01OeZZ7oZaByTXma
S/YzCwEtHCw9BtSJk6j9IYJV4VYieKxO4G46ugNmIg28ymmWHxV1U+UG1ADoyd5cGm99eiRkzwEe
cHohgN6YXzI20Jquit42FPQDaJZ/PFBCsdHeJTyCS9JRM8aABaw97C0rRaeBZWclZv4vqI0VJEfL
G84uMq5jGGZpD/GBu/SxMbcM50NRcL3lViI9u/U8Ju4Ku7/gvw8sdpzS1o6unVchNz8TeljDRBvH
F89ny5S0uQd/x0KfUK0cWhWCY/2sx78qVKvA9qJDicoS01MyZ08P6CXpSHaF/M9Y0DFPvd2ERRZF
amjzfvTIt2NwmjqK7+81w0ZUjJApIVxWs0RP5l84sUO+lc49UNIhDGaCR6dlOOEgxloDnKx3P4iX
aiEBH57DIvQKd2OXpPTpfLf9nmdpIm8HrevJX3xrxqIiaLxI7eER1sQTUzgwZgjuN5V7hScu2KxP
NsS3UvJoLz3/FoyWpc36sfx8ixK1s+ArnnH5BtYr4WhSB6RHXNWkmNhBfgQ2WjVqWm2VqPOyPdyB
/img9OZ8yE8686xBNnrpeNoaVvOnmAaLfQOTy9URqYSYqOjTt4DH4fnAFbVjloeogJm91Oe9T44S
icYvu0yHBjeuwnuwK++lt6URuc6A4KpcCijS9PqSBSzleO37g6evzO8tvmheGcu6G3y+3RjVgWMu
Co+1MVbT9+Hhty/CK95E3zFurB5Eg4rMRE5gqdKJpZ44wHu3IfTJKHB3+UUnNgAitB9AIpyLLhSM
zrdG/808o3xnNmEgc+vbe7EdYwKYZmr3rSubReuDAbm+xSlW5ZoQ+imUnfaxs+NcuiOqYPDA/HYi
3RgIs/8N9wBTk4D1UC05mq+C6jbBazxVq8JJivV5AJa3USudhMbU+e4fSo0dsjjRglxepi/02XoS
Nd8H5rGtipRh2T565plfIs2HHanj/CnUC5GEe/mk4oeCOLw4/qN3n0WoEZoeFJX+moH7LCfQY3Ja
eUO7k13HlAzhxg/vG3DPiScZ0NYX86lZls9gY9/NaSoQVD4q4JvO37rB8RArs4A8hXwabPOAC5p2
JOuGhJGVbwe3MLofyULZzE6UsUlH66roVJcORgsVs8sZBpMLRsnVm5v8d52SpLld+MRhsFuUwvcP
Sw7xMMOHtBTBEOHfagq8qogweo1XFrAzzogaw/iMTX0lic75lPKSWWGX7Lz02oTYqknk/huws/Is
32AvdVC8bgxm/bVruhEokxZnPGEvP7YBYIrap7XldLOCt/HYQm39sVj5gs7MlXz+AxvAScTTyp9M
oB/Q9Xb+Tvrmt1Qpgqf3+g48zSArO4Dol4PnewI5eclVQLM3PWgjum+tJPZD+EhFUyM/CxLcmfTb
0Ou/k/nIjerrhBJQFCHcX7RioKZkoPSxvYEg6ELpHKU1J1cU5mvR4CRTxa1cYqA37jqV6IkyWzPm
JC5UmOUcLXaTnvs2MKaSqvexVZQINn0rzy8GyValXFXWkYNG82oW5GxXzDkxROsYPHlO/xSsu+Tg
Th4V2O84OMVe+vig1zXe+lz7L/fG2uKvRUFZIfENfnGR9svFNOB9G2O5tBozysJhmOA4Ns1S6kIW
u0+XhEd8XhooItVZ5VhliJW3JYUm0/qbrDYI7HV3nzdspbXOaw2az4tc7zkPkeT9RNo/8GkMOobE
d7TloCILUMqtQLLhGbOvso2JqbY/Tc+R5guBv67ehTSONJMQNYLNmxmhmW8UXufILMwdd6h6y9oV
gEyRl4YkqZcZHNAXJ1PkKZ+FMKpeBcVxWQwHZtdCydBix+u42xKiTtXasTDaS5y1gqshghxUQGC/
P3h6cbuNAlYuoXKNHJWsRInQnyn4A4QYKKPSFXsymdmF/wO7W1BrA8ZMX2XgDmvGPzoQ7Vm4sEz4
O9vUXN53pNniqd/MM/+gZiTXMQkgzh+Ngf57TIvZuSdALMUoY+j10rIXTLeJO7z5oWzeGEZgk513
JW/YG4jk/X7bY89It7M9yfg9yMAPQ9Loh8oL+i4zQjFHeT+o+FnPZ2fLrjC+bW9Guc7a7e8+4/xz
PzTL9zGmy0vfzJAx1VwnCEm8jTIbJyv0EUzEzAaOggwQk9+eO3g6LRoaiKt6WLLORINftafS2KXA
EmFK6d1BhOIaPmlkF2qfuJJwfqzoU+Y42zA4JCuUpJbt3qhCFYFhh/Gvs85Dhy7qg7JiWO6OIM/l
ZuUHvdBbSAPOnDx/I0zs9ag3s7QgmqQELNYHjLynC7YLLCVfmCuYM9FbJD2pq/qt1FyZd4THoZQE
QjsxzcbkREZEbVx7+7RB8XIQdfrRZMEj46MvH/MdvVQddAXUURGC/0Obuus0FckD+2GZB6uTKPU0
yoUZWO1YFwaU3FGTS+bj+NEQNyL0JfpOwGN2wQA38owyehbqVpCowj+QCOlKLur1YgBPkDL76cWp
L/0QgHZcFK8OufnvU7FZUVO4qiHuV+FhmAySPdvqwl4hM6Icb6XZU931lWgjzhm1qzLEUJtIW87y
+EtsBhsAIO0iYzIIwPKvDq/C9UL/rvtO5uCLCY+NqSxCjaZItZFu8xrZO17zHy/u1ayUmvJmCeWR
TievVhmWTXs3/6ujNAiCHevhpBneN1hs0qSlS6LzS/QxmGm33IYtljs/oQuTgIdGpv/j2FJ4MxMz
BvyrdI8NSzrfkDU53RRxljY11NWaz5nrwe2M4FfhZAXl3QkaTlPB5YUVPHDQ4tgV5j6Zhs8ehVr6
ppmNiqo2D9xQ3U/Z8q8gJ1qKPTWfa2XIZP5PTei5iXb6pS5cJkWWMOioXaOmmyQz8ef3WYm/vNxm
f12wcpItJ7T0lqDRbrZLlW2jk5rKuPIjilLfBSAPS7KeivdZOgab5w1U8PT+67yjDNstI1ZEmVvZ
dOnLalD/9spMJKXSDusWiM35stTAQCjyGYNK3f8cUV1NPJdoDi0dEvtth2y0E9I3iIQfMdRcR4G6
ByEsINon0scnnh1ChhVxptwHr4ztI/6law55+zUquAiKRsDDJ9UYrPmobmEEOJY3NQTRPLZrcOVq
7UtU42iCO4huQzjBAV95uPdGUyF0G9KgE2MDxRj+RXoIIj53Fw+bybr4ANeHewV2pLdUQMhfgM6T
zTJuVfuEEUmXW32HS/MgSgGWTAsQvhMOlT7zbysdXePDRVUZqq4auHHEs61cz7lW7MlvwfhpdL5G
fli/F29xH3BPUJxwhSEoEeOvkSBHoA/e5AsVOqNBJG5MF1Rto5R7oylMSNs2Wq+PlXGo3hnwE9TV
dmLhO/pkt2hWXBQugF0VpuZkH0u2Mfa3qKd8WtRKTE9qAIXNrO9X7U5C/HqePvMsdXy4MsfbXbf7
HifvB7ixaRZNKEJ7PNwVn75KEYhykseBrShhUr4MbgNwC/Yr7eQoBrYDG82n3I+B/cvTrTRrS8oV
2rXpbq8gGfIEwcYp/zxTS43KcWH3ZKFjduxk3uJSBsOjHxLWvKKtZUSU3FPVCw/buUAq3cxod8zD
Yj2XJZUUIohewCtHHB5fja7Yx7uqU4A8AJX+LBowoQ9YbM3uoc2BLRmD4UQOOhZfwEmkBsT/TBYd
ZSDMREHO1jhqv7wlzzfe+1mrpelNPO5sgw6HMgXAkX6v+x/DF+Epn0Ryu3+YYMWKH0pWUD8JBT80
fyqcdy9MI2yIHkhU/3pR045txxPMnVyED7q8BdWtrzc9tcgQetlSkvdaHu7f2h8ILh8JQ9ZksF0d
c5AoRc8l5tOMaOWqkWPHkBtqi+fGaWClsj23uxDzDvPQTFgSZEL8jY8uGW/O1UGT3hbBeCoVaV62
RHYGNdyYe2BxcL979nU5q71EurHgpsqX3pFX/x+CxEmP4ckpPftbgCg3WWEyKaMA2XObps/O1FNi
VX/CgivVfFpvqRYfMsg5n+UlTgE3Y5XPNz6k1FTdnVe9HXzQM8Tg/tK28buy94pGsJCaEtii3WCa
A+ys4d7mIRkrGmhXNAOvXV/iwrLkzpBc11med74j+Mlsc5pJYoa3aH4pIvCCL9CzxwK32+rQa6F9
sx7GNT0qXu3PqUZ3zMBhjMk+0vSiskBCq2vl3DOwQJYsmc868V20L2Rh1+IrmWp9Zm9+bwElLp9F
CgEv+sMewfP0Fykne9185hKAQVTNtLjJS4S1kfM3zullsd9Sl2nVAmlATAtPy8CvxFGjQTO8dBQm
02Fjr5eEq9CfdWzc0u7TsjEvJr+2nDKo/7r97/NSvbcgENIYrATlshcikwiv2orO3Ah7SJ96Vz8I
3QjGwriPrKKbNwJtZZifvdKeSwmYf9uphBXTz7eSUeV3ULkUlIxWhW7cd0BqjZDqVMkcSuhac5lk
L+l9X8yLoLclknDHlGASGqqn3I1ULCwvFRi+fH0JsgwXwifFuaDAsZL1sPmpTYiIKSZ6zKWaNKNh
dwwORRSo7PW55k4ECp+B/07mS7pCCX1DWP+ywDF+JXxuFYdOG+z7TOziA2zbo+va8oKhdPbn5++K
mZweDkRGkfiQ54fsC81+FVbu2xTPInhq3O6/BgqZ/0NXdmNThZrwUcBFIExrvo1M7il501iUhn1s
bV2jIcPgJLJzB7/J+VJGD4dKkFsRigCzGnYF8yCSiilN5b2dOja26JK3pIVUJcmRcvi9rGQqnGlZ
KpBqSR2YiXJ63ijtfzxeuYbnCNKxMc2PcfSH88QgNaPLwDpdifW5NFHAG/f6QIH+lZgKilPlJb6a
zV89kqHGa7vrFhUVShb8zXLdaXSrIwzEIdjYy6Qqe+/tkxKd3kco+l3CU5s3eg7YHLvgeo89pa4p
xoXF5FUpNcw3dzhTn8V8bAiZH7XejLuz/u7LJftcUugdnBDE3YdVTd/qfid4SKjxGUddU4nbKtGG
wYKWUkD1YBUWwf9bAWuKRDBnTq8XCDfmXxNWmnhwDqmKD8rZw8bsz/9nVpmu7cPYvWkuGzPt/+pG
Q+/ZFnIhzr8642qAnD4pHdiYw042zDZpE6nsQCZSL4JGlbcTmepF1bs/1d6zogYiN/SoA97BoLiX
S1WolvRUSPLoTy+mrOlcp+mbt7iRtSPCcobMWAYnFCJFu+DofBetDkqC4qgtMaEjfw4k7AZoaMtW
FgYL5sN85vAQ9ZlwKHcJ5J8O7CRPFCvbIs4naR/ADjBt/y3tclhESd6JjXsXDZTeeF4K+8XFODjk
5zIe5ygTCKyxMPOV6ssssRBSwxgkMobeC4KDshu9RJGUIAdniK5xYXK5SyqDA5s0eZ0TH0W0Oi1k
sYXDqpLeMBe8x/9ROohwm4Fg0qra2J6iDPkzJn4tXigUlnJVHlw/jhNESi2egW5koQIg1Hfsp4/f
zFKPGUBOFn5nFgaOKyEp+KgkyVjiCFKUce53Xkv3x5kt6g1DgVMBCquoEqL8FtC+r3kdv5aggDPd
5clGi6mIHoc9kHmi56eMCguwUi8uZN1VJSImaF0RgO8Ben/RVUVugaF00uKPypZo+SUBlVOTuhog
Oaf742zs0b6+ygXoewQsY9gWmuy3LMQoiFxL8A+sXDP/On5o9IKpALNaXG53/tPOW/Z5Ya72hug5
JAyvjrGCm5lBJi9oId2cV3EK+4d4TbCzbP8013epmRMIZqCblza8ckuT4sHy5HrDGzpH4PxRpNax
0wMXAa0HUBaB9VdUtP9MrjmPX60Ov7yX8pE2e4Rza3EntijwDZ7z0T47du89q2B9mi2QXEArKy/p
4GkRTFgYiCEDySIYUmxTQ3Rsxo1BO4ahxRXdvhMq9N1EgZdVVmuXRRT9sPqHcLpSphcVFoqTvclj
YKA9Emh4fnF+mDfNPg3U1/qL6MIRSEYN238OrS3mR+iAJgxeTuyHdBQl/99M0MGNzIXCgHVDDWc4
ScqHDuw2PIsBLUn/wCEwVZ3EJy8rTOi6W8IYE06WdYmTMj7ePHCzL1gvRslnXdlilq5OM2TsmqXs
hqYwqMKkbsisz+7Yp+akcpBl0GhTecw7Zkji2TNdLo8lbS82UOI5rZD4TkIEtFzCiL1mjzYGk+p6
Uaf3P9A6oTCO0EGf8oCaQbVtuiVEohm8u+apV3n1nhXUKmvO11ygE2aw4xMiF/yEb+Fr1emt5MED
uwRO9c2JQA4TYYE6I4nGKxWTk39L7WWA0G8n+H7uwQs8BtoNAidOdTqyGhQ3oRK8NHL6DWB+C11r
6+r02zZeJjkTRZR2MF83XHoegtJHNZ9Du8J2wSsTl6OLYXk3tH4snAMn/nAvzRRhCZH64JclBXij
K4Kxp4JUd/dEqioDKTuW8+8LUUCrgec153IvwqNPl7OUYyG6iooR/b9HPpUrWa6x5o7DSE8y3CAT
ebt+Is/ryaXurQjYfANnbRjkaSbSAcVFd1h8OX7WVUPuOUI0qk+OqN+j225Uuzw+6pgY9mHNqSA5
ZClb7kV1UifpIumRGUO903la7Hq1R0A69BZIULfr/S1kcW9hIq5xCVbfxs+MWP6rc3ErxqmwmUbr
PRpBh/VgCagZc4UxJCE/yNrr8qb8znIJTOWeuFotm0cCERzTQGYwb7/PMt8xipEwt7G3UMhwmmVH
6IdSXVAXXR/EPs+bRX6U571u5dAQHg1QDYqybUmtofFWrnLBYX2OEAQOEthS20V5d0B+y0TTHPj4
ATa0md0px5BKZajLnZ/ULRbfl/EBnQtwWJhN3RlkXe2O0/vlPVgcHvEAWGgCTAXNhXEKYJ2YISSa
yXYNfi35ax46ERT1nWeRQ+hzwJpSJASOPXruLi2sgMdRF6UGhskWgyhhRtS2Lgo26Y9JxrenEaEp
pibFuYVJ3vFCxfrZEirhXSbAcSryTxJ5vIlIpOC97Z4OICim9qRqSZVnJU6adwrR3AqCAuMDwG6x
IQs83bferWiILc2cqHQYPrC0YChe2emGc7HIOgt/N/8jgUEJN9fnXjKeSJFUTQSmqh3pDZTPaCQq
6jwR4rb2E0zMC9G3Ns9MS02nxxQwOO3gc4XbbV8gYnxcio8UHRt1SEg2TxZTD3VR2DI2fguJENv0
umewyX+BNWcxuDD1pnLI3ri9zNTtrwJcxH5xjjgYGBHdBgyMZnMRERByEbtC1hQNlkFBxGZxCsdd
L3TCZVqhlgLAeugL7nkLQ6IYsRcM9RGtFBKj9cRKaZsHdGzYKY7GqUA2CS+v7QpOFqxN4itBaQ6d
svUM3ysJtrYTUO0QyvRsgBvEIk+KOo4gvyREjZzhsC0SrMV6ZBwfyfn5WgeuVc2DauTe+GQthAuC
YGn/ALd6XdByhV2vqm2dweze5/8EpG2mibWwakHeyBfEFKa/32ML/m1lqq+y72BqgwRUjoGPqlRB
2qNKM8Pl/0a7vfTcecTdOhKTxdt0gA5EWJMihK2ljg7XPv4kyeSzLgxgwOlM6UDrAwQMCkqcCS5V
nTEQONwfqHXej2FyEZiXjwPZYghCt3XRy5gWLNt82VdOj7WSXNfMDYPOoozvCLx9HuzIuS1osFeZ
e/egmwj5uIodxedbqn10Sj11pqcdBntlxNJ5B9MxcI+9yt0BOGy+cmsY0SacGg7slQFW7Uqipg2/
WRO8ri0FXZDAd79UOjY3g5HGlL1K2ly/2/RGtqMetz1CgpzeKPPNKMzRtWze0GwuhBuYgQrWWWD4
LLNtQqZskp0Wp3qXcLhNKPt6Q1XE8D/eeS2QjTiTkRvNUb09W6zMQWByYKlDeLi7VumtJNr7Nfa0
g5f4CcaYdh/W7oXFLOwQ/UHgIpxpBwKM+UMRv4o30RbgGTkACy//a94q6G9Bo1RNuwQj6V3kz+C5
lStBe9803r6kkccB15EJeKJ3aeYSOHyx/CBW04aT/4GJb+ZcKfY+2Zx0khycLffg7T+DYRvWID/f
qioNhGGIOsXwv1LhFnEXOHyuV7VRKvOOFTOifWqycVudGtq7qABWSV0lKw2JKpJtw1k5LzLZRF7u
NmdYNVg9twEGq0SCjYi2gEX7Pp1RhL2aNUT6sLMbH1vrly+b2H36UbIZQOQy4cdGRNHa9iZ4TV36
aaz2Z+mNOSciUGTLVol3VYLHL+0SmUejeMb4T7TXwq4K7OdtJOzfoCDUtBhgZCcjKIDbg9Ynkqsx
/jah5fi+1LfS/iyxNdlpmd4RMz+e/czy9Syl5q9O5S4h5B2k92CTOJCaecT/pS3XxtYB90iYE1qr
Elpr92nhMI6ttl/domUFADMJLJUFr1L33NhnY7ds1lwhB1atlktH0MiZAa2X6X8Km+M9dSD9wJpQ
R1dm4WEK8PF1Gpjkg/tCy3cCmn8HdLGe6Lu0JyZQHF7lnpD68dTWVPGfeazzGbyaM1TA7PSrr7Hp
quw+aIrY/5DnyK4+v5zQ8S8DaSU1UM1jLHwfico/wirZYuICigJEyqEympIHQgeQbbHRnoiaqkMt
QfX8jXzonyhVeFRvFoZkbeZAe61jQch4V8XjpOkbAckfpkIhzxBXbd1E28v6NX0v3siM35HhHUpp
AfEFS26VHRCsWdl6sX8H5vL8edP49NuAhoWfOjRbFxdFM70AEn1TtlSynNsQKZIlQ6o1o4xuIrFZ
jLuS6xo/hG4U3ShEf1ckHJS+va/QQBcLE2ZQpaURmfihZTjV2P30oODqBBvOJxPAHUY/04FKerq9
eR7gwGDgpMyOg2KZh3xi/lTmTK9ePJhAas1P7cdbRx6eE7azftfblGanzmrGjINYIvO2y4bDiL1T
xrvfvJP3wrQ5cmlMRR/fZsjKxSIHZ/yBa/ZbKYy9LqN1Mon8WR9K/ChhQc2eiAeiGs570qkdkQZS
M3pOZWaQX1H6UNBBHsiUWRK8p6iTNHlUvhuHCJS4blY8k+hkurUMBvE17DVlaPzuTeHT8FHeQvmz
ut3CyRsYWbiRStzopafEsKkpSpIo1RkRCwlQC4JrI7QoGDPWBxEtx7UXd9hYuQ2WQGiHBFXU01+4
0cG9v/SqcISfaNYBN7CIvCH412oIW5dwNxooAqQsFLcqo21XA0I48sC905yCV0uNk727C8vBMDS1
JqSC/RAnISu3IPdw55hWjpcw0CgcQkKnJ4s3q6XWDeRDGmUZzTwVxKOmzDml9JE7p1DGZJi4gn0y
WmkQfAPse4Gk7yCaeRNQGmmW8o+ZqkZRZME9Uao05rE+UJ+WqoIh29EYdTLj/Pb6h58QEP3Fbp5+
FeJjGnRt3d5dWUjqlDY23ttubwPe5vG2kgjkxWN/f6sz+uhtEy/+kejccW89nka1CufQCZpxGZq5
qb2eomolgzyHeFNmLe0s44jfSaA8taKcpoFXDrrqHqDThNQqMNDWrjH7/mSdHp9axoCnAbASXiyi
C/VL0BtOn75lgt6VRhHCWNPSI1KIruIV6kb/pnn8CFn8zHUmviPKK9GJce0W+Fo/qvvJheLICQAM
X5WlRUhy9sAh9MgTM9Q1xNqaNulTpQNj4FJnXvpkog+4zwzj3RrEg+ffoj1WYB9STW3cg7vn0TO8
5BQe42JGq43M4YRJcl1zp2E7UpOCNg7kF4DXYJEbze5405FG0xU3ezpp94arLdUfSLtWEEDOTLmj
n+Ak95JEbHwiX3woz+53wy+00ss3deI9BeydYAfrqRyZ77+2Wqw82ep2k4qPa7w2SDNgVOa5KQK7
R5MBk663y86BcMQ2OQNCj0Pca+mqrr11JYJZKDEsl/Xdd6EraHwzgAVzHvxf9ZBx43bw4NniAit5
B6rqtSb7SCoDZN7OZhniXM6CmWjRSSWeWHpcfUysrzZfujtIw7SbZBoOMoYp3jcgdG32ajUdUCb1
E7GKJYnGXo7kTUVBqVYJljycnMp1L30HX1Jc7grYLJE+pkLPwNdAaCa3TyYRmPNvaSqMnB7vwO5F
X5fhqYe8xAH8aazqo7jnSBLCSAQIZ1A4omtNTXpl/xRxe1K+AoCYPO1IlkUOHuJvC8aTfnpcxcWb
9OlyrEPwsw0kYz2t00xWVApxzzKIYco9Bw7PS2d4VRwS0+1lhvuavU/srweSOZ7BJlHJykPV8Xx5
xMfTWKMKxMULSP19qWsb+ADjhVMJGlN21oulJfTDbh/1iWk0PGM5N9/H/PEnrc2o/yr/cHfs78Xg
L44CXimKfGlGMTzYAgaCFNYLM6phnEsmf7U4MWc11Sge9pgzurw5eqWe/3mteVh6k2jdEGf2hMOk
YO8GZF/w62QOqQI2fHoZeEG8IoXBMdpnZO+xpau25dLnRphUg4y5joyHO0qe2uoo6XfmbbfMRRil
+iafv7pHduro+dXL8n6u8DJcJEbx6djm3QaE9oT2MRFjuCQibUaPdip8d48J4R7JB37D2Cj4heOx
b4a6R345mF+eAXKxhR1jVTmQBxbUITb71pBL/THZ2xmLDR9DqCDoFykmx/jBcN/sZXfzCXJk3T9E
oRG6PBnKUNTP02N+HyBHhdm8KGNo9MxJq3kK1mMB+GJqelTTvx7dd98SYSTOswS9DHQ1Gc924oAY
je51n/eEGsa45xP/7L57cGxNvUpql8HEqfv3CBdTv1TerjWyhhXPARVHmFVVrOj17+1AQk30HZi5
j2KFF9JhLqncYktwneLVob7mW4EXQDG+b0WR16pakW1D6soBh9y0DBVJPfuomx0+kdx7+mm8AgyT
QWw4Rywk12qKOeVHG6J53cyw19h1+Bs2UNCs3SaVIV9mJ7JNouI3mDasl9aby2Jxn4dVeIyloYjy
Bbt2XOcqlxC/hCYu/OxddOGXz7HZ9giOW22rTglCSzYD4BIFrBxvpd6m//7r88Do4Dxk1WmjTB17
1dmR5lLN88xLWH7W3q960jvL4DXFCKl+uesI3a+472DlhRD7JinaAoF2OvZgtecHNtXXLvAepdXA
Wc7vUnLI1p/qfH8aJ2lIhLffGzPP4NPciKHm01XtpKigcdjrFHrVfqLs18/B85zfsY70gZMbnecl
OOFDZgedP6hhEcmRIle56StXeczlDJK9QWPE45Z8601fIRLH2MmwRAvrr+QmzZ+zaErNTyqp6uDG
Ivqdc0NIDCs2nbviPGnFz10u4zoaV10+mlQIf6nIBZH1KIh71vpffLa49H8slFT7eIDJl4OfCCDr
4wiQES1hT/tWJf+yr8buTHVPzi6841DQNcxmGAltROjqnYg9xhpGG/gBoaLK0L3dRbVVTeNa/2hY
Y5mn9UppR211ikg8YCYXqH52bQwYifmRMRfEww5FKIZTv7hPWF/ull0CU1YRKr6k0lFIgYqZKOFk
wHlb87BlyWmPWU4Q2WnSSb2XZHQ0ovM8QVHg2Mdf4RcOaMWGFwaooUwyheY878VXX9QvutZFZV/P
Zip+gyIiqdlqmrP63ay85S8iTgNY7//XewHW+qBEn+aVxMRNOTcVqA2Rq95Wbt8rDvzqQWq1tVgZ
SrTlvTRUuMwaX0KTVDWVZ15JFPYSIzc5cATYKP3K1g84XsVc3BdBLcq9vBkp+L3LT+YpKeuOZigz
5wNYmOSZVKP7OUHhXWTDVqD9ACD+QJF4g1txH4PoR4L/9qJkvC+Ko9vSy/uT6bO6QARSSM68GWXb
Er2oUGOH5EmPkQG6MN1KMHXZ+uED9H2jxGQLI8EAn3v857TQFliLroUuWdELQ3ULbgo+LmmoT+LA
i01nhX4ucfm0qXXuw4padBBpzmySzff/900BZXfxwxInc2totx1NhiI9sI57kSXoNG+WhgqlWMmG
Y/tZNHBwxCL6lbP5a2C55aLnWXQOziLtAGAAdnFl0w/g1TJ7LY/c82N6JPOSBVG4PGcDKuhRPagS
gQ8sKG5QhvflRPkcPYIVc+4TNk4LrLFHFnxcXKtDIQu5lhjS+MDKLq1eNds32mjbO1SBz/3SlEmV
oCSwOc/arkCgbFpYaiC3XDk7krZODqdp7MGQP7vTSHYtXtBANpsQnw49yXKU8cseZgQtXz90TwPc
FOFp1s3UCd6a6t4mcCwpa8p0oIzQCqrp0TrZKJpOCiO6nZfPGIx4Y9O05RV2PunL+3RgRdz5W8NI
8Xv28yMg1/8tcLFan13EehpKN+BaBZXUHc3jKiXkI+vjx1V4o9nTBfbsoqkPAxQPQDxks1qdXTSg
JbpJ17PA4k0qozXeq2SUZhNSOnpUZAvP5K9VGk7a7eKn5hUOWzUMUgMjdBmcOUtKr4qjm2K9JinP
bTY58aDzoB7K1tpw7C5CidFb9JaX3by7OHHhm7eU1s/mBRpDcDTxuCvBc7Apz2YXXcYBjYnk2G6q
SyZNVGfOj+qpy1lSV9dTpASUuHW4XOROjkyWA8thr7bBhUfAi1V4+b+Qp6fL7vZKdJRp4B1L7WCO
M0vNCOhWmLFboZncR0D4VVyf2OoNWEISdia+SfBTIvE6bxTDnLdRLiDbW/YM6zqqiKoeZAO7qLvR
BjuBWr9oAnr2XlI+NvsL9bN1rOcx1rpsL6EW2FRdT+5d/57+Xmu12Mud2APQfH0Cy4GNo90pM2ff
JUJNCZ//k7K2sE5DwGMviu/xpQowZ623WvTvkI2WExQvBnvw2WvE+hvGEMYNdLWQf+tBHejCSnfq
CVf8AaOM91TK+7ikgH/QL7lJnKzKa9fHPTLlvQijJPGH309vFkzVXeejbDtaf3R9LD8mrIB+ZUqO
q/Hu64p4qbNKAuoU0gIjwqLMNJ15t5SQLPdrLsGtlGGPHxEjMW7Dx3UAVDtLDVxNqPA0A6LrADye
l2xtk261JLftOTvEBjVnL8Avzib5uV+aFG7TfK8hK/26NfYr/kazYW2XjZd6FZg6R1Tt4j0ImwHF
D3AGFgoUsZ1iUGLGHvskRF8duEpGn/P1MlQ55JofoiXfup422kxy3tA6lQwCHwvwiz/lc08deqBu
kRd0zwyYwxtZoDH+lw5AkDTHoCCDvmwazowh9Vc+Xidx3/1soHOmrOdLXsHo7If4Aa4hvhr/wCRK
TRsGvaOnB7ypVPJn09fZSrR8k1rRyZtc/fm8o46S22IOTvUSnN1H5plqGVtTgchdse/7S3OhiAPz
f4BeaOAf+oGMMdQeFQtkHU21krXuX/HOffgxk01Xn3zLlweLh2yOUX1svq1ZL4THagMtYUBnZJw6
8PRVgE6bdZyQdZAOvrtiqzj+uxZUU0sZ/aooE+qxEWGm9/LPehcNOWhr0sKSKHwQGXslI81TSH9f
mkhm7qj66CJVS3RwOzHbpmzi4XmD14fiw1ZbXm96j2eG2akuH4U6UWvS2eiVA5e4mmjrXNB1iY+N
9DKLq9/ueMzZDdBPE82cN7PugO61PcbhDTPmlS2LDHU8PahgKlt5nFepdAeL6uTC4VoePCV4Hfq8
5uSiDM/y/zQjejK/ikVIQ0RV+zO9hVGdhpC7HJgaobTZZSU8F1ale4h40yK1bfg+ajlZ90G63xYA
rgVdPrIayeC58HlW+uoB2KlRMMusjViJ57JezOfSrPGNJdY79HoZMxVjBY9eDaahoWUdFfmMtuLV
smoFByNo2hViJI5aHACggVtNojAkyGwAbfTG3hGauYEW0dyYq9SyjoIItLbx4ii2y2SWfz0Cu4Tl
EEENQZWVD7MROBhH868zhPOVIivvyrHkpSB+xHpsonwI8M3wHQFg/9O4Jrzt5dGb98EXgQBev+vE
kKlq7ToQ5kbgHFaHqrvjkhQtMw50KJdiNE+RYqE4SdTlHyS/XrLRrhhJI22KUSj34O7wo5fpbj2i
j5aEIkuuf24tlkVy9dpDuK2IOJrtHvU9O2Gw2Gh63iZ6/NYt+40KHc0mfX2VEv33kX42QY2x2UF9
e3O5S2LbLSpE0MCpFcNKV2PahhHaNinm0Dp1BQ5uw8s7e922+QW4UBSYPQggG9osMd6eEfQmp6gJ
hcC34kUlmWZQN5Dy95xZU53iH2ixGbkFIQea/ULYvsbp10zQWcc5aLemLFm4VOxm4cWmzj/3Dq5r
mB5xKbVWJbPJvGb0qJNyY/1cM41fTsvW6czIDMhfF2/27mhA30AhnU/IiiB5RhmR79y1kWe9Uf68
mRpMIHxf2ziXek2On8ij3L+grqtT8SjCzrBuOA3EKxQiabhUKVLg6+034JLvFaUf1C7ErVpzxFVI
XX7PgXY7xbMLSIkPtSgyR89MbMuKMo92y5PNiwEjaQ2ENfY0QP8QX5j1eRYioyjzslOqCE9KtZNQ
CfsqWw5N6GuiqatKCEREtZZgOsNXkgMeYsE0XMqwUtoff1kPjKeMQImOqtDZJNIiaqvTIgfMtQtQ
IlKGJsR1nUi7q1Tuxrjlc4Sghuz4vMxT9/tc8Qg+kHIwvITAjNbat47P+AKPiMccYEVuZQ8aOYI6
QaQzBWXwsbUPSSNUudyiuHO+mRzTgLjyT3sjGxFeMkzq/t+s3pxQ5/K5ESCwl3an6nKmAz8RVbvn
L0bPZ5XuC8z2Ecm2b6U/HvZRmgpPmcyOCCEYmAfyF1xUvYKR010fVZNz/v5JwvjuLa4kx9bKs8aP
lv3qEXeFw+uoKp4qiPuERRdlLtX1QH0cohmhNClr5tIEKs5U1moTQfZ+U/fGc7xumylxmPq3j/NI
64aFFL6pirJbXePNz6p83cVKDgJfyeywiNE/PmdIW1CbV/GhfKWFGxD5ohBqVNjDnUV+Jb/D0WsJ
rnzo210e7wsTmCzLf7rCxdlzWzweHSj4ifQmScgEpcQ8kcQGQ6QyVuFYDBbFg4AMy+JyDcELGwsD
ppOi9yAza8oBhoxngKclEAsuEeddL6GECVdkmItZBcv6MNFUBPZSbGJAbi0FselKWGl3PtXrVklw
uD9nTd9Ru/TLys0NgDB6ebkoaKiJ/SMSlva7+Sps5hRiVcPCQTV84nrNQy5LpRGWEdFGCdNVW9CG
RYwosz4LCP9gbY43ajNiELKpQWegOb12Ti9ZsmMOa/fCMy38uuwiwivs6afp63vGw9ZKVAmFPFYY
Wf63shpl6RMltBJGHxUkPL/rhwvkuu+zYgMBNvSaGQ/d3U19FduHIXbPe36ARqk0SjcNa86CbH6b
esRkE+8fg1011r5XJrNcuwKE0hen8RSs+qGbIDzIU8eMsATZxEekxHXmevDtjZRFrIp15y5xP3At
K6ez8xBf/OVmj7+LTSQilUN3MZIHdynjY1RCNgIX02JuPNP3ieMXOPuMNHk6XoPlF9QSuk0A8VY4
TMELZ1btTyaFyZ5KLPApXldqWUcQz5/CjuPzSMuF8XS40AmCEa6e7d1uhbbjFm797sJdqKfuvEZt
3uZgn2kVn8XrcntKbk05BFpXxu1ZXXRdDPtQ7X0UXaxDEtGmNehGkWIhJhDCYkdPKWf23VKRcMvI
v2Ycwiyub6TtHuJGRRjzRFevRudUf8g3+YtxB7/rjn8wqNgRDXFCug5cYLDsfs4MjIfAN0rL9XFd
UegOrD740TkS/oxPWH0Nx+I4IY6/AnT9kIQMiz3MERFZY0HHBWCGdK/VZ2gzCdZ3VUVduE9Qo9kQ
bVhhleZiz1xoQNajQlBUnEt+jZ1jhE1YE+ju3K4nYfhXy1Wv/7CzOdJ2nS9/AHLggXXFLQo1Eslo
7ig8K9nkoLMqf8zXpBYlCu8+PNW/57Mias/mDx04VtzsJX5s3+Lh8o2fI95/nipwrE3sVFhoKT4E
0qybxpLzmoRJ9xjjnud5TeEe6KOJ/K6ZN9JjZX+a9yGTHUGkaXoW/RqwfOgWYSzRYu92bawW75Vh
NTN+Zy2BJNe08ViH4um3z0yt32N4W+j4FzdItHU6KwxH7jgvM4AH2/qa68757I1nEAPnMwOSF3B0
uVlY1WIQEtVvmMjahxy4healBl0irMinN1cuN96u7VgWEjfYkySJ9f2SPaxE4N1z1spQMu8Nzw/p
EhGjaIDg8AM/wNFlHZjJkPfx3pbycp+Aideids3A6e9qMmbeQC9+/L0d3RQ3KJMXLdP22nRLnANN
Rd7sGNk3ljBsV7dERAuCbW9b9XZ+mmnGoPxpM+zKMzjn2Z4HM4zdsgrqvqB2H075WqnCfDZf9IVW
Y2VOrFHf2QXYPxHXoKo20yO39k9G0UTpUstz0XpSXvOw9sRdT0uW/IG58/iMIeF+iupO89FrbJLU
iKRalbnYcg+naGAOSEbrNthq5N1Smsv0LQ4QhubSwA9lTrR4Or+anFqqIz2MFo+wBcjiXn6BHYPd
O2KUXVHyWa6VmozO6ZZaORUrxd/mw/QP+40vLaLMA33RI8xL+kaxHBZlUTwEaFFrS/q2gY/IBheb
lOVgEHOyWmWJ3H8D5GypP9yrcR06W2Cm7i3LWJ+HXUSOL4mY5eG1hLPqHBIJBVv/fDFcPt2d6xFP
dmyfhEnzHAfK5JWyFCRhy/JpjvLQHi0z92t1au9jO6h0T1eRDogIv8g9dLrZADLTTHdmj6Sljf6L
XjnAPPug31V1/BvOE4inn6asGIbHlmoFM/45awOOGa5IzL4nXtn4G4YjCgBiexu+PuOFaCEsjnL8
MwTWuh06Tq+Bd+gEJQcd9oKKGs046yB8X5x1X7WKr/1bDL7fD7R/lWKte3/ikSu9t2E3MaItLP9Y
0mPdJQMfS4Njkp9sw5Vx7iO6I0MkUbeRzE3n10BJ0CWztsG7nzNovLb+0WFkGSlFsUzZG7HgKyzy
ZHLfL7l7wYnNm++lPphkrcC+zgxbu4asUIG1sjLGI21ctehahrruBKyB2YQfhTlCc+UXyOWWKIV/
Xp66dCjO04mb7xu/Gu63gSNETP4iVbYHWKn7JxMExsyoPzlsbHf23aGYaDJ+x64qL/Q7XrZWjVqk
81xVc2XkVuYKwm1G0TDJ6JKphl0MGNMa2tdylkW6R9b2t2gSeLXuyOqvGUibEZ8d0Ck8F8kDfYMO
3taizE6fW03Y3O//juHm5dAJxvP/CfDdJrk9Y5hu+qre2vuGlPFRpwvvHWdEHbZhtqU9X3pqLKmz
QTpDyI8/uELoZKSsoktuW/Qx+8G9rEM6hhUANue/fEdpxDVVQ6LjiecviG+9A53DI4m9FTy6M3My
EiLRrsEK4sAT98dV3eDLBu063cMf833/8MsIneUYjOHDBC1UHJUHVg0kVkHh5K6s9tvnSoHZ1BxN
Wf2xfZdkOC6PNpBqeBF6TaadggaBW86VPIfufNr4o2ZbdyjnQfCOSuxIpwc4aRLgKiZmWYxvsQDL
oZYRhZ7om8MSYzzFHCuewTYoCI171WFqTIdhQ0psppYM4Cs3cywPcd5fK4KlrMm5Og9d8lawMt1Y
qMgSThViny6GdRyWpOS9QhF6KDUayIuy9Otc7CIhsUILgKQfgJSh+81OyLZuiHi8Uqgo3uTnnvqF
MD0PEeTA4+k4qecddkdXl13CqxG1duIF7b21gHWhumgVEm4bQmOykoYWE9lKVUVyiZU995oH3jkp
XquZBx/hUil+4MY3cSFvXbdYqOtu7xWsEHhwb8aYeeYbm9j9WNTfCpAI6fIq2HBI6RoUmEwdlplS
AfCbyPwNkX6+EsQOhShgx8rFQfT66EdFMHT/0LkjCFCN6YTJmnbb573nxo45KfVTbzkAFj8fItZM
koJEDurwrFcua4vmk3fB4csE0NR4QEYagS9RZ3x6hrI7w+SlnSviMxClT1oXXr6Ovs2KUiChlWS0
YosPiqJEy3EIO7u/4/L8CK5fae/m8JH4FwrYp6oineAZ9Pks8wSbzJJMsNpW3jTeJ8nRdFp9qXEP
oCttXrZ5ruVMXzC2mu+uS6GNa9SPfhPECCkSNhrtFjq7daxBv4Z11ON8g5Plxp/jSupw8GqACvOc
nYIaN1GGH82AOZ333X9bx1egDIfVN52T1McTcproqSCs/2amOAuBOWW5f0OfpXLvs+Gzq2km1AVk
lH75qn9Szm3Gr9M5pKk9h4lc/TkpUsoNI5BIQ0pPhLsCeCEoanBPuOMmL5tuVYcEXog3ensQ5Vez
+Hbz7FryOSQQLyGs1xztcsaCxYi5U2Joj8L8xhE0gx+eEo4W4yEZXA3zvmkDFkGRnQrsr9WA2z1a
yNiCJEWsiTdPRSskbD7OpUA9FLJpLgzMi/VNL41S3I3jKUMvsaww6ZdMUgEXAz1I+2VLX/8qVJ7+
FtTd+2HheB1XWwPDU4NbXvmQIi+W+rI0bmVQhHYe9AdgpROcVLlUwTH8Rx7crzyX4zSMO+4YJ2Ak
GYUvzBlyDjPTkNEibRTtpY3UB+t5gDg3XiJNC9Gy9Yheg7A5oybkJQY/QwYs9ZJzpRX1zmaTxGxE
kFMKFQQvWJ9qkRW2IO5uVH1N8VKvNZyean7KSvFysqBWwEXTrbNtvbW/ksX1dmCNhTFsHRxalpM+
kH9KB7kEafTOBHa8I2MMW8tDMkwSl1+hWTjyxrTBtdEUTrTvSa428pbWj+DpBDenL4nOsTtH9vvh
Ev1kYvAYq5RPFXtfxfa8B2oIlD9odgGo/2Bl6aPdq7LKu8DuefoK2dKHU1RV/LTqlhiSotOYJeff
NqoFNT7oHHZEhZXVPtcE9/bN/mKchB76KFGbO0kIiOZ+kJD4X05/t6SfmOx5ey9BkwhgymWWAeYQ
MV0xHq+xlTPJkkfO0rvuF2o/0g9NPCk1OswdVxJaEWYS30hotk3mWck2XK/SowHC+yucyuuw8ADV
V5np+jQQUm6jPppZbvunfnKZmfgAzUCuhu9AfLy6hM4vrVZEtQKMbIoOpEQzir4j1iDZU2dCDhtB
Dj2OH6ghGHAES592fDhGV3wL57aRZ3EWXdVzgquP4aIDU05aNp/ID02CGM7kc7FpFSIrgjE8LPuR
UefJ4Eaoj5yCWj8X7ElLEXwpUjuosVIH/gTUT16pwNqVSthgYvZUYspaCjBWraFdrs982uz7kiga
XhCFPLVrTv3sgLIP9MJXCk+YljftL0FCnSl4PzBkyxwM7WYzo68g4QLlNqeLLGpDmapHWzM52Jc9
oHGYzv9MA0byHnxZ9O4ZJONlGqLKM1JzZJ1LQma7plnjbewUaHueQ4A6GdkGAmoT+1A41+0jfN9m
urlyee+rKroj6XxouXqrHW4x+9SrWLioWsAl6AF0PUiPf2RhapBK+S0bQdtjD+gjSF4eLC/k0MzJ
kLWzkbskKynStFcw+qNjswi1ORRW+PZaiGwbn1EpcePm8Ewei9TUn/OrhTRt8PENzx+J22G0WNS4
FCtCUbXzdecH5ui4rMaGlE3D64bnbnqgYfu839oEy2bOZrPvN8EOAKyjJOHBu0C44bf4XqyWqXAE
BD3c2NjXNScIzWNxaZtfuzHsI4EOfY8BXVm+EJ0EYzk4OtJaNYmviPt+OZY0FD8t23DSooXrhvKK
+7hvQRINWBlugF2cyWAcGWh3USMqFtPdn3FHCRq6cztWeakPm7QSCL7ESk7NeYyshUAzHmJefsRH
ka77TMqXyoIxqmBaKvRVlrKRTuhG1nrR+w2WtTd7VLBlHhCW+gpglxwHCLJUerjQFcNIDvqTX23n
NuSCZcoNhjg7p0MVhPFWChFZq1jDO2dXDs7N/Okt4UAJFa9QRQcDBOhOn8+cpKH0xsSEt+yfPqK0
B8G/VOMq9aqCGVeZG6IYIh2dRR+MrHM3twyU1nzbqE4FqtB5bxlKWz/qcj4rl1B2+fUixLateHio
FU+G6Q4rSGDdmgO5akjVD4ZnCtAirj9eQKHtpRXjxkGlN/HgQr994aDOfgJNg0JTP2fCFNspkDA9
KujmUQIydjR1gS525iu1OdJISdGE1oS9VCFlyAy5tNJkUOPDY3ov1veMXEk7euW/Bp8e1N68s3vQ
pc864feQhJW5pOPxKVvushTeSnxNzpRyyV3CoXehC3LNrWRwsk8KSnkXRRihvSNQgw5OTbnXAm5q
90rnRbL4roRIigycSbnJXmpazcXjJPaHzs8BVy7rfSY4gTA2UTi40fWCuyBuLuxfI9ab40mKlhdy
gdF1C3/6N6m3z6hgYES2fBJc856Zx6tmg56SpAF0jn4T9YZiqXl4Y3WYcA1nPDKbLXsxmGtwA1Zi
Gnnvyo5MT2vKEgOglmM7QtuE1uoVemQChJpOVVIQiS6D9vPEh3ifjElU4/8TGczbAnQJxVKxAGqP
Bk0Sfp/yTvx1Aa0+CCkz0Bj8URs61XlNyWxcR+yVUIq03lOPhatjjeEqJeDW3/EEJiqBiJpqetkx
Ma/ollHxJ5L36qQDdLZm1aU2CJGqZNQ1akGQ94487CF5ItNi2k40zpX4KQi8YXxehO5uGyWuHyP5
aIoDo8aVthg87UpPn8bsZvw414+lkojFiWxSR3M60EMMsx+ob08yiB9N0/1ZXJbEL+YxjnB3ATFd
kmYg1LUOSUtCfmVPD/3D4UcQqWLn1OWX0zbDQ+Qk5gnrXVRBeVJYHxPJuRfbH4CvwhBCLU5/Rj5R
TVZUrsgafrjgABINxtRTFtnSurhUQtKxw/g6fn0eTli7oAVqOeuzT5SoWsPf7XZ/OiTgf6Rzu4nk
R4kIhaPl8QkCp/gvZug5drwkXWYcaUbczYEy2pl+4MrtF0SE8TrjeqlksQL9IpEeLPWGqreg15bI
6MCRuZuzCy+kVVtG2I3hQt1UFTTtoEHueiInT2ZgUnBySi/rR41Psav6Gt6KsQPvw0McAca8SsXe
+TQ5LItrQDYgnm6vQrb8A/UObo2Ve1EBNZ7zFwRyntHcSd3R+C6lYRum3FywFsjFkUKwtm3sk3MQ
bHLC6TEY7/RYJeyNov9FMDD3lI2UIhXHSM/g+TB1WIMw3MixWfJdDaKSNxZ2cZtfeD+0rz+3KDY5
dpFw651CsgZtCGzXLmO5qo/Xj45AAvXPLwj2MCYbfwUgqKJBM3aCkkhdi1V/gyo+8LzSYoSa6Sg7
ZtC1QdH/p9MzsNLLMaYRKpKFXGJvb09aaS+extW1nNu3+Cd+ZSljvRAzxnWNh+Qel2AGwLyZObYP
rVA1AbzG80K7kdaCx86y7H4vGCLytKVLuKCS7TJvMlWxUaACPpx2QDkBaYRFTERlKybC0X8EJH3e
WqQ0YXZdC09FjP3mt5imuOyJ7Ss7RZ4d1gqsO70HBWDPDNlkC5FLPgWudTMq24UBONigz4FQA4Av
Nz4k+MqewRWma28y/iuGQ0B2y0dMatNW5/SKAacXI2CoeAD833lfgoJyHVD0wg3nqYmj1ewBJyDw
R3X7vD2xBBlKWrGFEIFmy7m2dcPpMUUMfJbY7CO0HDV6jZqXjeWxy865irgj5AZWO/N4A/KZ7ZFu
qOW7MQrgymEsPq1wRhOxMWote/Rc5vSTb4kafYcUSHpo2aLttHUEW11CjOVclB1bQaj7aguAhZK/
ItBbV1ZqAABuqYI1HpiLS4R28SmOFT0FwLCqixGNEp1rOSV9K0fmMuTi7HxlZq7zrY0MP4x4DqOs
OKen9qGuRjtS8zrz/Me45vu9Z5Gn1P6rtjpbc6+JkXPdcKq8Bzcd8sNqXobMurQ8MSDq+3Gq5r3y
daBi68BLLKD7qcc4FhHoP69l41bVFL39R0hdHl/z06CINED5HycS5Eg3fo5YuK2xyo2nFhdrLp85
4T/sWwNzCnL+DEsrDzoOLFvqzcj69W1ClHB9Z1bBDOIH07zA2scRk0cmcyWPxueg6V3s6NDYQM/B
ff6C6nTnHmcyCBC/7mJovN2iVx/LhtIffm3XWNdVcSEGIcnUe9ZbJPl+3EekT05xW3uGwXgUdnRb
v943KCeS+GA0UQGI0eTjw/jSmm5XrOY3EshNLqfb3tPpm1d50ATO9i2PPCVSNhpeH9RIk3DEhinO
1MDKJyduFk03/ReacxfjRvE/TblpJkV5h3j3s0gvlC/SjbgJpGLTkPWtuZkbexR2lbZDKDJzVpfY
Li/YCo19ce32Jq88q/GZt5lV1vGupKDAET/4OSpwXmYeYsFTIw71eLOIrIa3PrzwYazfhNHhgpbk
PP8UANfDzqB6ZqyFLV2mDCCOSkQk4F6b71o9MmDFPauacGKMGyNWnQSad7GeevHPBZXVQfK0l5KT
rH+IkHnsQXvCuLJGY1VdPm4/kKFJwBz0Z1oURWmr5laKXuiEj4LlSVjyYSncPQkuBSUzGsk1L7nY
kePo70Xh2sv5JfzkbTYuGsSt1hJrkD/3gKZZgAaVndxB7AKITZYfFZOGzHPDjwXTJO+C+2WXzGYg
/eVXNQ6Q6dlfT7d871jKsRaOc9iq+bZdjiSJ62gauTWEW41nQpFE+7nGaQHjBlb41RNAQG4TJT0a
IZkWAxUNTcaiw255rED3F3UoOJ3SWWKktxuOlMbraSpsgM9UoMCV27F1mCFEzeHRVRTGEmUMMPsj
oW5AICPVmxZnNWP3Ue365abr1I7kEaeou1UeAD1M9W4BngwlNohe0vdbd5bFIzU3EKV6usbJFIsZ
uugMkOpBPa+x9615fKl92cRE9UDvryrGzFv6gT6TIdHJp74CBsFUDKWp+9CHaXD3Qj32epLShhrh
4HGZWR8qcUTI/+uNrmWf8Lbj33qvEr9oubCnrJvTUXIWUXJyVnpdVVU0NLLz/7rBwuQXiP3wijGF
tMHHKTzqRnJw1Ej7s4pw+/tewqWtJ6OTlv/Dflf4FXHb04QC0X7rbthGUOMn7rTzr/XMAqbVTv7H
cEuNubJu1OBR8jUeLiV71SlSFsp42VRmV1hJHkWQU7rKmEykizKJ8YvYQx7An2L6d6Q3xwOnfJ/1
FNDeWbikNeqe18+6hC539O3wxxv3X5dcqdTfzqnJ3iiQmQHR9896oMKutxwRoFVZr0v2/UBw61vt
cEofUGG4tXx5JvZUSHt70FFSblHYYbsHF9a9M+QgpofrhTb2X/E+vwpVA1+6ytxfBx77d2mLdinM
xMOQsnik3adqB2ZwnT95QZFUsSPRvyFgNLYakHhMCI3JIvtu3f39ZQV/iIPnHDDQyKlANZNqtkw9
YoblkOTvEaCu2HGfIsRvdj7g+X263aGQz0TAP1lgpBXRcFRQH4zxTQE0rkge9nrQqfygoRFJuH66
j5uS6EzsDm0i7QRAfnuxVyiq2E8R+8e2Fab3NyQp2Aj+u0/AvH0zxeUDovQlNWQB7s5XF0bHB+0r
NwzwAUwIUFZxMiB7V1xXKMdk5v8EevqrFF1wMAY6J0bf4V4nh3oLy7KGzHpiUe59MyTvGrt86d4f
V+heLQNNrNOXa8lKvK4cpQztlBT0sSxmKUtjd5z59X/nIrFW/HeoFoiv2iAUJvbzld8sWKytdMld
g9ABiRvzAatpugmtULdD501s+c5puE+KnzNO/3JlrX+vkelqN5CDIlXZZ1y2YL4x5H1te9ANkYbi
YSfP3E/DJLArA6hsfoZTjeepPgZneAIv08DCgEu2aTBGBfaUO27G0Fsq+Cze6wd14KvrxwaZmUkS
LrJ/3izD4zAT4nHMTO33Y2eOUitGtsnjfgmD3te/53ZB8Hqx2FEsgIo+F76GtfLkWUEHc2bKOBM9
0c2vz/f+rmHd5LbRF2M5WmIbQhqBeCzzsDBzLmcEJFtK4RR6xQNBoq3qz9jB9rKtARkkJV0z5Avc
lgPB0f3cdf8DUMmWSSgFgqaKaEyRpMwOPUgDZzq8V39d71kOU1bYVrVM6WtNpK42UgrI9LvPIDuG
1K6NV+zCXeh7qKzCteHNWk1/wv9ktN+ygqcgeE7OfWem5v0Z4938RjvZMqu+/WzDNsbv8uV4uzTE
FlMKIvm+LrhglRHNLjnUS1CKU9/SVoMlsoLXeB/Cfrx2nWkPmCssZqLV6MnGM7AZiYSjGRXvli4l
lENgmsymwCGbiPoKZv0YSSzhXoa4ZpJTz8vj0M2Nt6U1v9+vDoNYRPuIdvXhSQCk3Ra0n4pFjKDY
uYFEw9gayJD+Ri55sDDZ/w0/motyWsfUMSE9/NXRJ7kKLQ9ujhXDqCf9ExH/jv4AdLQ+pNyk1yO8
6OvnDOzPRVY7gLN0PQYP0hDflVlh6lNx0fdUCfp5PBgOE8Cnmqy8XfQa9mM0kW/R5LYs7URT1d+3
IuLZNlMzwrdqvZdLDb9/SdovJHENqJPdZUksBr4B8ou1GHRIAMXhWvkhdfUrnHLDs70ppaDOQFv/
vgcH3Go8QRcRaC8Y4F88QviarXP01RTfyyPrQuJDpwgTpkd8Mqp0prpjjw4TYmKYVHKqMC2cnwvq
ttC+sdCofMNty5zsvzbGNTpWhUJUHTYQDKUWYYgU6V5DaPYSv8Nn1zMy4ZctTEInAaSx4KVU+rN1
bp/xXpkCAk+tMAIByQpwMj0EAiEpcYGaH7u6/o156V9+SySvrmVsWRiEpO2ol9I02r8h7zvvSyGp
HTdlef85RkTMEsXT9fK1OIw7ivAsvI2ObFXAfzfSmgtHTC/IcWlK9tYTr5eybjNz4iqujTMY10Q0
154HI20TirmVBxkRggcpS4pmXbwqll9jAduQKkrgyF8rANaEN8kQ+TiWKnb85txkCFH9O+mjGyp6
TJGBwLAzrj/jkgxCFA3AzOsp4DHs8ukCo4rR8qh8a84yrKCqpiUUAqwKUcrXMzlXiQxjCqWCsvTw
iQ9yoqjcI2huXS+Ybzajgj2XYY7B6LiyWuHFO3DV157iGbz11+AhyHqICORTB3CBtqxWGE9u48nP
EzgxxbVxmxCYpRBuMs7pgHABkM49nne9R51ZUv/wTW2Gae/O2fmOGhrH7AZ9Sb3KLKDUIGkyISRa
GGTBkGKzAh/q/BjpdrUJsg3OwCy7rlvuFyGp3HwLosEPtMXXyhLLK36T5jJxpdGO586weMK1sBWd
ZCgynulsvcHy9PmnCGQOOBRp/7njhOPTtMe+9AOKaN/GdpakS84MbFX8SAzz9ijrZv5EqMmFPJZ7
lwIsjs2i98Fi5cjs8v1sgtWGTeG+yeVCAbt5vmK9qgJTM3ql80cYz4PHhLdCbW4SSbrqNO4c9Qpt
bAfjvWQPgelp3LjAZ5yBuiuIII9eyURhYYURvo6aMTJDhfH5Ab1cQVTlu4/+7xy21NCTd0pOjrLG
EjMx8Ui8CjWscDM/FHSsSQ6dXvHGDg02dgXb4rE3fWe6LBz5sGdMxL450nShJglpAZKCf9VyRar9
LM3javMGvosme9peMAG6roEBgG17GTZq4RjRLbR/cgSr6I4KUj2oANbVnK48flMS5szq+xhtoLsm
sYjc6cuqrw3D/jNhRM/Od0//YlczvSwY/8foiy2uu7mCtLqhgwI8Pci7A3mBaVPNa1bPo0BQt7Wr
h/lgD+P85Z6LHRRWzulhhS37RwtwZ1xhsjSSAuwXKcksUtr9ncXgzls3BkBioMiR1aE4fH6O53ch
SpF+xyLltShLtABqEZiihul22TkOmx6+GlJPFZlqQacrRjjEJFWbyUMfDtiJfNFk4VnJahVDVYvW
p1k08Jgm4VtO4BOk1nNbKa9BhMo44qxR0zTNAsSpymWNosu6xj1kHwFhbmjI69F2DNBD7PSghYny
vUHO/iQOWCJaQ0B0vaahqFsPGLPH9lH3HQXD+eUH9kd7fermqLCSJmk1JkV8XFQk5NIIXWwVcdMV
LHTbQfVGwdlQ+cwcn8HEKwVBDS0dH96EG3+LyOm1XhF+3oWkZEQC/dM6aenG9xjRwPm4nPrGsYuN
stxK+pD18TmVaPDOfxzKr+t/7w1wBRHSuLMLpPYflwQbYcCqWOJzj2uN07Hta5L40c8mcLj0p6ae
vC/7YIjundJORagM5m/tH0rLHrTegBoYqDdsQSFH5cQcKRbXvKNI3VBy8eq8d3xVPxZsyQT6Mi5Q
oaly/TDnV0Vykw2ALJkhNR0xWw7zyvlxh5Cv8P/q10D8kUvuE80E0dNJeGrFPsnrBxiOpdv6wQrv
G8bafiVmsnLbxATF1LaAVCIMfV5r9qoPTCu/oxRdjqmek52zsXRA6V0d/2gTMN6eJL6HxJhdZziB
/BXXX3Ez05TzGRZPQZXFwZwFrkWtG+Ljho1Cov5BIQW/R7fF8qHLxWIIGPEbJNHyo0DyGGD1zfUL
ykj2fYJWrcNb4Fn4LONJgqZzz95eduzTSRkuhwpuLpq1stmVYMSD3KnyL/jvihbJqnhIlFxno9Zn
M8C9du7n2HtOeWqJMjbsq6kRnPVdJq1YeGcx4dygZFM/dftAoQpoTHZsyHGV3LuotnBIjPvY988K
5a1NvZ8503XGh+xa4mNbnrfRgKS21jGMcdXvPrwz8Y9rYU6vbDmqrnsEuI8fGj7vjlE4JFdskuNu
w5MX/Wsy/nlhpvNd2vQtcko+t10iwXFUz26NTHusFq80Kj9ijbjHezAAR5ghvmgmx6N9NwFmMAuX
6UTKYJcihtMoHejoa9wgEXo1NZA/i26a5O95oHv9Wzzjny5QxMORu31Ns9WJZFNmvazfnxNvPKmr
BmOBZH3PjbAm2l/FIIHozbAiL2Piex8tgya7h6oSdZ9dVvrgZC1EjG/X+xzyFhn0vIVWlAVeddbV
W5s/ogWRMYNN81ibfL5s0APbmt6sO7TcKZS+km3wdym52sPKbK+JCE5y/aesFvzmk4PV+dXGGmqA
by5exy9eACEPmK2ryjwDGw2OoQ5vP2NMZQimamkYGHybOPSuKle9AXquNUQjLLwns9XMT/QQLRBZ
hcsDvfFgfTdYk/SUSWCbKZrbvmRKxPaK5rZVi9Pbg+T8+az9Bfb3RYMu0O6OHwEE8QjFGSrRJtvC
W5iO6p72ul/FPOqm4aA4Ao/ERs+krybWv1kbtVMFCWt/1D8O+kOx61n86xcuc/M5baqLzo2qA2H7
0oYVrSX8nKwKEvcw2wtcjyRhM9frxM7dM8OdjPynf9bHcgfcT9rBdnNbjhoiv90BCh7uq20oD/4w
HtU+KLTmiB9Yvojzs29DSRpocAbyKpHIq1mcgMzQEATw3OiHQMa2Sq8gZ/5y1/kSFjBDOH7n3DlZ
ehon7f8fPpiHCE8s43q+YLuklOPL3FfDDI4jekhnnAW42GyNJsyHutvFeFbeaoSJJl/IMhQ+U7Me
OuFKQPszcnj8qAYNVs0J6wju7QOxphE7bAksxPSJnp7cDhMD4DGFcL0t1wKEJ3pVMD8MSFXEghkK
lH3tjq6D6zU6DHZ/WpiGYkH5HNQPqj1csYtdwtdc3T8Knkubf8QR8vVdoKi+fwqkm5Br+N96IHCs
odzi1zzpTjjnL/9gWQ9+s+WcBpIWMqfBaqjwEEXlU7nVG5zbP0/+uIOFUiTdLidFFOv/gvZC7MXb
kWSK8NoBVhzLBDXNxwtYhZoCejT7UNWq9CDNs2Ox2NulXtkLxdOMmTSfAiEiHjpItVKo5D7obKtg
J4rB2DIb7P9AWGC38EniToAQRURqp+XGrSw2GMeLZPH5qHYv+Mci0OZFlNVxEw2SKHjE8g+30eut
e/lZFCwUMlS+awPDhSRpNreDXYDbuge6Sa//LOo/Xr1dW6OY4uBldgb/KE2DGsxILeZqC2SlSy0Y
qKSBSA76XHY7GmDTGHWo/VPGRnUbc6/zKyz7m+fSPmfeS7Z6h0NIBodz2XFRhtmtVDNPiinP9Pom
lI9G3Q4aXP3d9Xk/PZfQ297ubH8ZhgZhOx6FuL5MOMwtz8/TbFm2rsWtCrNPV9wCdEs62aT4+DKp
397cwuM0LHLaaC+eR4lyInFYlTYOpEE0LIa2vHPi9RjsoEBgayn3HFhBGyW5lxsp6DwsMe43TLnW
oXRGv6F80xgBeGjsTMYMUzZ3KJ1FO1a5KsQjdeSCqZUt/kjpS1yIcopgNQA7iivMVQMWl+8PIPiW
VR936G+3i3Bxv7BZKw/In54uF0Zls4coUL+CeH7uYocygSORALfYrk61WSFoM9mVm99Mijot49Df
XOi8eTQ+yjF+kQAyL/BQO6pAHD/90+3pA4/zZFQijg7m5M2fOehjEbgHFdOJn6c0vG9KfXCzpuam
TTk4oZQBQ3ta0CTvVTz38DCfNq6Z1q3omne29JCz6S7TGmQTB/YEkhw0x/kIgy/TL01uhEbiRV6K
1mIeq4eYMaHCgQwAl2jau+qhBUCuZl1J6F/WTm8CPHjTsB8Gu7WPTU64I/e/QynGGqEOowlrJdEy
4fSNVT/bKi6IeRGybcb0UPTJ2r49gHoKyhVWp7vLhw7Z3nn4Md9u38YmPhmNB3I0Y61UWM4ma4J4
kOaiNOYAMP0raHD0AQ2RK0I8ZvqMWD257UQ9Z5cGhdr5DntClNv5wMyCs49jAbhVYTZAu/YRCNIl
tGd6UI5JLXBlXQ/Twq8rFXomTrdTZNivxahtoQ4V9ZiH3HOFL4CNGJShw7o9d3cRGlYgXqmQ4T0+
Ae/Q7092qzOulK1a3FBmFqLW+q5ooJxCuOHEHMj95MtorrToK+xOVNkqYeNtyl7fS+wGRj7aHvP/
RKD4RCJP3AqpSPuktlloCeIp6HflSbqYCvDodbqm/3xvKiZaULtT+/C9sXbDNn8QBSLQDtNNW8bA
59FNUmWvXcNws4K4RHxcvPyUaAb2IXEo1bhbEpJkpu1rdPsmeCFtTRFQUDuXpxOMvDQaxy//BNOO
nltowBS83wNI/NDD/aZC9G09B1lgJLZhf+SuAs346PLPv50vSMf3jwOIILYjItDRT4SvaZ9tnDqM
Sjzy33rhnz/TIyxFgyzd1Z55sziS+GxiQ9kvE0bnEvmy6Eq6d1zza3VOqoZmuP4I5M4vY/TNJuE5
ZJmrhY4sHGIMD5TzsKijt5pG5Ixa3B6mlOVCJeh9TuLZQtPyCfcGSgVuTVWq/KSaaKT3gOUu/GTj
ilVbfafm97fjrQ9V/dO7ywkbejwrKzo1bTTMVtN/CCOw+VXahJZumNTwg1VHLNgf9HgHhsngtuvc
wXgjoR7YpZkVayqpbFm91vYYedL3ESH954yKL64earvy54Bk8gOI8mCh0M+A2Qev3FOORKCX6uzp
7uTmEHntMgsBlgSixAdxRFlQldZ3cMno1SPo7H2lb20lgx1hrkP2IAQpQLFoea+quXObPXlszvG4
ZQ83ZuMFXxqtDJ3pbVaRBhQaBxQEBo3Y9zEgf3xGjuERbdNAA2ebPqGgf5htHPp3E4V9v8BmopO/
VJeDT1zHN8FWQp1+NruyIEuzj9R6XcakvHxk1tqwZUH3xl5dyUku15G1mdVosE2mxvVt7K/1G7Md
hZE+DlWhd00aFgYLa9v7vE/+TuOxemzfzzPlc/uQ5v9hD1nuInJHRaQDRQ1r5pHj5Tx0s+eJROEi
3IgfCT3umkJduncBE0eLh9tx5IlFAQ5bOGTZtTi55EZt3D7mB37t20AC2fW5rMOMzThjS/pv/x89
QbgvaUGh9+0NBlTnAxW7tboJQX/dgHxuaQBOx6qzcJTN1IVIeFke9weq9bDQXWl9G1h0OPZqpxsF
2toMX/lLaL77YteLWWlsENbupehN8QEE9GdbgAbmXeB5YEcVVQY9zvDgBtbgm3wy6Szz01eL6/GL
eWmbxYI/2r3DxjkQj5e/fDz8mGNC49rRNum9MWvcHlP0hY2TJK3s5cwMU3tIM5P2nmEaHdCDD1sL
ebRTHekSmnwgxQFSb4ow4EqRq1LmNZ55W/jgObpAenZT/sGCqQI/TLJu5rnv1H7U5rEFLxS6RzMT
ChkGOsgYKguvU31+dWeSE42cgwNny7LvESsHNQvg1PYgWh67kVYDzL1Mn0MJucmX/XIpCP8OZ6HY
HAX8GCU/ghLhqtmUCM0QdzNwsJUOT+20/tOLtdS6+6U11wFIStJGxlMZ7kygknJdSOb3cie7mNbu
gayxNJad9jQwarbVqN9m6O3pXwrdgxrtt6rTe73Aiho55Iv/9aZYVeC/6rUh4wsPTL0R6t8FeoC2
PgIVXiGJLBWysZVDB6aSNLbc6H97/Qpj0qMHh0GUuhQRAySFtMEwk7QfQ/8GpgMcQXxV77SKRtPs
ydewPor+R0ZxWNTJhPUb+m6MkzLr0cjuxanMRX7CSLvnsh5vrMBAPBeazUWZv6pgiccGk7tn+k00
Ln/8IwQRYBWWbhEkBznyjOF2clUvGDTrTOdl5pFr4ocfjTDSFhjt9scx0BtbZAjhzO1cEnS4j0cx
bLKz4OKYdZ+iqlOJ63pJ7bU8kw08/6DErn/Q4F3g/rSdU1vzzcclxnm25ErCbINKcCJ0ZQ1/0ziQ
PU8ZrefwZvcklQlZpS1jTxlil5/e95QLoEPXMO46Vo9n8WyHTT7hKPyu9gUXNeBA75HpcgpwsD6Q
zzp7ktwzUNMLFAR//n0w5w/KLby52yf45i15VV5g31rNCqW43zIqBddRXsjXCbtAwgoOCtP6Ts0a
vZ+C2NeA4FAEhLFkDVxC4hilCqbq3WShuYQHb+kfCcgKrKaA3/bGATIGcFyJykm+dy+LuDkygys0
sdbeuP1FIlM3dD+bPdYqyR7JYskBIJhBAtjQuUrdC3QLbOu1ns7rOKL3DaBeeLZ5y1kkGudae9c7
yBM0mat6raRhV8M6QQV67FzXokyF80v/LE0h6lChaqvgIBlzCzB92j+/kNunTsSs9TxlTpbH0Jbn
Fm35Gcl7AxwrxXRszvaerdXW2SeildUv6q0nW0Gbjcj/ZUimIDeQzGL4uo26l/QUd/L5X7G/xy8z
2LTI/tvtUgwtl7AlR4TnoxybQWpFJ5QRAG2AIRkOygpN8571vTNA6akL3lwXxKkzaUEjRx3dDWeu
s6+ldsaYz/4qFcsbCBEHx1UwHSyF4aiqA5RS48WSx854WLFz75IIy3Il6Vvm+SJVEZDAKFYjJTL2
+jL7DZA3hhSqKO1FdLXobstkIg1Z1/H4LGdVLhDAT3mzZ4+U6+KV6jPrnFXGLEk8Vj6rnmn9YQgg
dAirFwC2n81UD0jRPf3oUofmmEQgpYtDQyykI+gPK4S3Skd/mluyhRrFvPn32lEBoiQzfIajfRE+
Dt/P0SDQ+6kU6PVhlhx8QcMz0Olg2nwOYUkoobQkcbL7qRhRCId24mUBYixGSpdiLVi7cWYKLb3W
Bff2qsAP8eeeKWMWDw+4WOYTqSl5mXPC0aZb7hcjBD9744lIvjsfuYyW5w5bnNPt4fAr+nN2WUT5
usgoxDTGQTl9QRY1ST1SXYJ7SZSiT5aHpSsS9LFw4iGALEFIJarE228SCS6q209FVqH+Oc2HvDxE
1MpWxznOXfKFoYZNYEStrfYFsMWsF4fdsXbly6awxTB5L9Ar88O31Qxbsxi9hhAtjs0qd2h7YrzO
VgVB5nfMwO77XtzXhL1YhARV/FrLkkP6nK4rhHL63RPaDNYLgjHejmSGazIDfOIMeSOO16kK4QZU
m+DbXWKNLwhJvSqBT5t3klQ4axcu72Cd4CXD4PNjn5eLX/LsJ8fqsJEe3cOJToajLgEWqMHi0pbl
HOCz3rRo0BfDKJZBMnPJrpna3xOoated2Hiiv+9CExH7fMfcenW3uc3M+zGjB9rqByZPhkS4Aofx
5v1lYf7O4MOubjYLJTfNoSP448Gm+iy8hnAtCTq87rss7YEvzyweDl1OK7LOPCY+ghE0CDUR6yS5
KTvxKM0+vheeTB55DOY0phDap+WyWYkGMknXjuWNVVOTXjKalvKue1VCQ9hEF0A88eFlJu8xunQi
biUJG0GQGeVQXY862yy8vNDPmJh6lTVvOyTiNlQVS7ONrl5qZAY1JQ4RSgGqCZvDjJ5PyuyNm70a
/BgWXUs+xavHnkBZYioz92vZ/mpemldNFtDDZjMhaXCtFImX4BEdpr+hekINYKZsy/EOhoiPcy5d
4rWxyTd3BF9jILzS177rjlrP9M32JTT13crFzWdAj7WP3SnFiu9l80Ku9jzBabIi/tWB0TUAOVFy
x/3Dgp0hZUQ/njgptaxAxpWWKzXPmo+H82reI3Ksz4WviXvHK9gC5lUG7HvXlpSn+hGH9HQzB1Ir
IhekUVkID4zoC1gR2bB6yaAqlALaY+nzW6x/T5hH/5wtsMlU5krasLgfIOb2jjk+pHhqgKy2mVoA
rHQlSGVcBN/OnOiC5sQYwy8yCP7/3QDSMvXtpDkdRkKzHnSEoQFjdDB4QpdvH41uuAUvFWYLWOo5
EnjgMDAXfa/yIM/YFwzwOyrgdNGCii+BlgCga1SGlAR3dtE1ZOgVM7F3NGgpVBBqRGCWEejyvPae
JYsYvA7t9mnIUZaM7Ub8GastKvztmrE30HJ+5DHyrBIwiODy9j997VOboT4OVJ+A4VthcG/q6nrW
JiznIbLvPqdEN1W63QgKmyIJwnKUTR7/bchJ4C0ef2v3/BfVAhi+CLVf8uS4wqlXXUeYNG5552Ee
XkFSjf5fgOe550MD1ekDPbgAnGCr+4c0+f7puTIkmr5t+5+16mI8clCwZIeydtlbKY99Xuk16kK5
rh/f+A92oY6UqAUCcIm6DkB2VZ+y3aL0wY7oWULVulHvj+9geKNVkZyZIl7IzbPuErgKfOILjK1F
ZBf8MrtjLMpBURZjTycENXAs9n/Au7BGy8Y7T77RrfcyHem1I5B+5NUkBZ7jjQLNW+dIuztMJBTi
noDjFx5qiOl3obslVznVJ62roWMBBWxXaoQQOL6rQbxs/yQ/FSWegrPHAbIWXg0ZEaHgecZJFYkI
WxdydsZ9QXz6XfVFt033575xB9Nr2Gw2qbGGLZJKUjeb8gaSuEelQW2nGKnHgscb47o7yIEFvrsL
iJMmte5bbHb6pgPnz+Tn/fpNoHR7noaBMR4fdtTVwjgIMjreT3umkcAxerzKjEfPVLyaZAVeiPGB
RLTHfDdU0z/mw67FVgSwwFs9g0ohPDTwFONtXaFMzhMogNQdgcrlmGpKkYnHTOJdXiDRzBQwgi1B
2ZUzTN0DWHn40xhOT8ZH15/LqYBe0/s/4dBWKrG52vaDr0bGJCnWUKeZaXFe18LLR6QmyYGaoKkg
GqN071jMba3oYEnS2NSdrenEFmBqHWQqN0r/WsR+0S1ViUoY0dA70C61OVR+dogLUMql9hmfhke1
SUy+fLwmvgeAeLOZvqS1e2IE9/Qz0YoE8pXBoROlpTQTz7xONxCBQtxTtsyX+3Dc18aT0JhVKKxe
oTQRv06q41LP1koDodxFZbkq81CEvLy1BTLs0hDs8JFQSt7GnDfHZCB98H2Y7TSu5VZJS6lBFGUu
rItxx4M4sYtAgE3LqxcNQvB1M1j9tiMczeVPBPI/pV6x4e8Wy2kMZXzommGy4Z36fr2Bf9M9X9cr
qZRVPihE/jl3++svuU2aQyFpIpD65sJbaGELNt1BeWt23kVRkxGlXmCEZt0eQntXaPxbCYxzpYlP
0StfjQG4MuvGfSBnp+ydaJP7Uh23uf5DaCd7GKaRDaDHRVhrsoUfjhhL/vpSwjuK6DsASXmLx9UL
BEPfO7iFGq8T/fylsvSwSF3aKi8KUQtHZJBHeNEOMOGuJn3Mx1zIB3lN9m+IC+FJYe9bHe7f9CyD
/k/2fMsU6K1JuqZ72MChl3qPx64vyNlabyYeIeRNIlug2V6K0bjWVg/kR5hAzQOimxZG2I/HafHR
6stGxHvhXxFaU8KYlhFOCVnnn4mY7kxtlvgnmHyLozTQI3zDGwfmRfbvZSU9IkCg7doQshmOULk4
dBaC8etcQZsNm9nAB69GtVgPMDvQvoEMeq6PqCqQIObI04ZoI/Q1Zz9mqtgTp6cs5NPxqr625Xq5
Uo2H6Z/wRSez5KMjFrQLtP9qWdM4f8D8zrpWDhMvaXb/rLsSktz1wTeaEZFpYiMZ5PML/IUgLgQ7
OqLmjps+hV2p3BmCUOr7gzG2gnFa33kIuqErMJz7GStGU8zqxLIlyEiyUw3P2YLWMKVst50i2KUN
MhW/x+m+XK8TazJmwUf+4X2i007kVZ+40yN7wrVOrK54jx9utOFumRmaBLui7HrQlcFlCmLpsW35
Su7E0rvWsGJMsD3I/vehi2Gz+jMmXGPD+rNnvezRq5rKQdgVSNilkgXAlgAwuBJtN73tBbxIXWAS
nlCq8On+99+rqWNCZV6VbhSNN7CGu5jTU2o/3wkROg4xAO49jg2Tb38Cshq9pFH5y+shbi5ELSW8
AlhwowMRxevZTiuVWq2RNovobPjmQ9/D4IcmQLINQ/2t/3yXXYoh2vroCpikxL+Nz0YHINvoR1ym
ukl+f6cNvAkm/jZUyVk7B/HCxQ2jmLK0CgwqE7DOeOVRasVik+T00H4iW4TjdYkFxVp3/4/bTyJE
9B0P9d3P1pWr32y1RlEZW8+2sL+qhHFQGD3z3W3PXplYlFlQprI/8pkS4O04nk41/dLdbhBTvgGG
gBZtI7LLZGr9yuod62T+KyoT/maAQTGol5D8OEaIS8MmLHo89D/DBoT14HP5jHiRiywoHrM5VCxq
T1YtopjKqCi7XVUQV+XJiVb4+ncqYr7CyO3rtwBlTpXMW8xbeCQx2PhP9tM8C6Z/sygZxsiGJi5K
9ktWMdKQAeiLgxqmoLBIme3pc8V4okJEN2v2BByfCnSBNAvk8wurXaXrSfGOrbqWrBYIDxufxcFc
PoPbE6LvM+62DWEKiIvqCHZen0kGJzO6pfAh5li1U7F0fV01Yfa3ZSwwchBo0BtFTSMZj7CS+xmS
wY0EnYq8q86eQvntyLJv9RaAJQjgxoZpA5Jpr7tGs3XRadovTge/6RuvuxmAVC00TheLzuNBHSJN
bGhP2PsZ/zFxisUdDQJdQbHBgDb/HkS1YDTEn11uQ55Avet3L/B31epZXUJiaixAA/zvyJbt9EQ+
roqtu68IMuF2o9f0XzIjnHGKOfYvvBAyFmrqsJzMUKQi0YYxsKXYIv47bohTv7j1t9GHFAff7Mkl
Cap4QBlbCtHpkF8SglT50Lg+f/SFqn1mdVcqJ0y8fe7GGZZz7mhHmB2i9civRAy1yW3lExDICcVv
Whw+NjvCqP2uGw4222e3e2W08e2plYYSogz11kGDn51jJ9vDQWzM1/LRbCn3egCvrFGIeJUddhvp
sDV6qAzwFo+dUbHioIfddqvdsvlFOpiOsDOpHgTvjTHZlp/jISe2w2ml/ClPJqQ5MYRaJqtLvq5C
ULwiHGGigvP1e0pd4jFtlHPsIG7GKPPzmSM6Kb+aBK9IdIr15MkiLy4OfS1uAJ708k9Ed5Eyc0r0
7MN3QH7Q2PpeWUs/LjatWSns+mAp8SvLXGPTVo2nHjYi9I5ZrL5HSrTwX7/pUSAdgbbpuLr4l2ST
CVQlvl4W6cNeiI6xEqs+sXPbVZMq55TYpZJOyZnoZEnhyY0xAq66oGJauzMFMMLlgOy3XTiGgY5m
erS6tkg3PRghd1M3zvJSjbXgj/DOw0/PcletcGEvObpY+ojl5BnDVVYkGdu+oNPhvfxWdjCtPANq
siKEWczjVIlS05DqB6gqDXL8G6G3m7y8/In5krd5g5y8dekHwZglrWfMimhLp+7VWBfBMXdF4H/5
036UCfExJagQG3OcOcEA6uUiSlrxauzj5172QYwRT5qBUJBXxTOMe8ir8ZCHuZdmLAAGUlucMDdc
C4RZA4U021S1LQgIG9jLt40kXab4qCpC7IUeUHXvPbvHOf0xcEud9xPECHniK2SywQ1qkqZhzYnn
tshbQU0aksipn1MjkWvQAzWq86dv8KE6fbzrclj01VWRE/g1YayC/Zl6lqEDKOo45JJBuas9YJFQ
PGW7xcQ6BaM9lRUB0d2LE7ntyxrPgtIAj07rJok8WAO7pQl8CFRLys2iwm9x9ovhc1CXgc8MIwzw
9d9swub2+AtabKZFiIXGhcUQRFkL7o4nuWbJ/mTjb7XdJ5ddWCpx/g/FfLFNncGZff6UCHW2wB7f
apJ41f7K1eihk1gI5MGg47v6gu254sDGZcAkKUy4A1Iqydv9ksIeh8PmzWO3mbLBsCpiQvJEOSva
xr+vbHG6L7KUL+5R4B94Krub9cF7J5e4sBgMYCuaeYuBL91GmmMDOB1e1YcqC8+WjxdSiMxR+f92
L4ZWSFTjFj+uCCSIWphocE0pNvXd7tV5Dyl94ChaPRfa/QcDPizLBfIr8cltDWNiJFVj2Vx4C6U5
eBAPsJc5ZmNe8cywZlfFSQXzgijn1ViswHTnMUUP10wiM9Qhn4WZwdOyhXDxn2jCTepjlRv+s9Tm
mkMlX1Wd964YM/1a5DmEnVMkkTMh9YHfs4I30oiRtKTZA3C4DTEgtEZdbqXXmRZNDLp3ZoJtBvsQ
4WmermFclwbCInuo0LaQAEfQAVEXoUcqDsFJyolsQvQ1O9c5rFi97zfZxSo1G6U+kENNUy15Yt5C
UX8ctdQ7fW83718xqbKSQ1eZLB7efxLElylcRJlnX30UdsZ3j2XtaJjCwohIYDlRPBDeFmkSwvug
67VU1oe7gVSRWJb8idvB+UT0WYv5QOH5znJnJwlJuF0tj+mVWpOWDaaSjgXwDFmUf8bZnAcBhjx6
OuapsqhMBQbl0rund2OXRc//D0WU6E7lGpONGydFWRwbCLfNGJM1yZHw7gYWGYk7T7gEfZJ3Sill
NiL8319/TrhyQ8Y2ft+dT1wZQDs9GyKDNe9bcnh7hoZBZukSE2TFk49kiJ9BLu9/fKHHGhWMulij
ENgG+clhsLXQQhEE9YHuQ10op1KX/2Tgl6yHqI2ZddhWzb5otWy1MOz4zjodTNzFjSnrqEokCTqY
V+uT+wNW0BmpktKb2auS6lTA9jKnAFZniIKm7PSDkiVKto32RGC2Aq8z6XzS3ZG5tgzP5LJrOcjW
d2HaaQ4EhMD8Bx9KQplmKch5k2YqagzPnez+rfX8N0oBWcJbfFFKQPH53iZKI/VRo8Izwpixbm92
m9mPO8mM7cyrpKJEvLucnZxFbRUPlZMLfGVRmh2J8E2T9Ox3uXNqziw1ChVLECg7Swqd7n9xVr4b
kvaC1cWgpbObige8uvnjMe9mIYhL92i+iBUE37CihSsXt8pmT/TDSTY1N9KTP99uPZ/gFy0QOuEf
maq7iJTbhAXc0I+InvgkCPp++onP0kymwlfv0bInzxYYfd8H1KAK49gHQBjTQVy6jV1KK6qKFmE9
hGK0vZejuc1l0GmqF7Et8++tTCXAJOMveokfZ1CPlYTt3ywWYll8640IEZGB3q1BOw4hkxHs20I5
SXAmJ5F9QN6I14zsBp5uACpiDxRlCj3CmwrEo5wwlkLehZvGwpJBFsCQsLU1l0OQvZCyWHcF8QW1
HotR2qCdI2N60c2Otn9HI7sw2BkqLeD7yaJLMg1dxmr6kMsCaYtVninhO7yyLj3XW77nmN6jszbu
hjdgTtHIsWUA8+Sqgii3jfWpFIQC0V1vc5QkVntOyT8V6igvwFTC94lGhcyp+UJwBR1uZhgrH+2C
cGXk0kyEV7bJ1TZkSaiTXujHcn63sThWmqZDuVSW2ylj1IRy5NFrsi+Bq+w3mz5f9tcb76ba5Jza
VqpKwLDpEZTf4PhxN2vG3/Eu08TQrsuWcKOrHnUFbObbZe0Oj6O6mtPmVQQGIfMzacKbOJ0RPQ++
T6NgQlzS0MJ3lglRhVYw1gqkCL851NWqJgSagIcbn+eBo9WJmyyJJrSRGKtGN3fZUE6SEJFwmUDh
KeO1cP2YIh92oLACiWZcNOww0f+EEQ8Yex4zb+XnkvZGBgQ4ol0FcpdKllUkDOTSNmG6OMXOveMw
v47O8ZJamSsd+rddcAY+U7KJu15s6h8rciN18W0qF1ZfDwLI/ZGNmlP1iJcf4XK2Pdi90TJxs5V+
Z469vOI/ouGYtcoFJ5uI0zR72WAvooGhP3bKNb02gT8FRMqT4FVDEzpDy1Eu1NrxD5nogr/lPH3P
fR3vZLKbHmQZlkjtiH1HZzz5pEuBMuCzaMxo2UrI4M4zLqlaVBAlLmNbcKSDIfV1uKuFvWGwZ16e
7uXM9G3dz68Xpel+gNbcF/Vw+5+paOi/LZpY4ehjr3JpO84SUB/OS3kl3RUjK9ARUyU+4BfNxqTj
NnMgPoddCdaIDUpGCwtcRcpDwh+k52lgtzjddunzvBuawY0A/ElzRU1/t4lqLqEH5t7WHLbd6SBh
VUg0PWCOYTKV3sQ105/JOtYPcvW3UW3VdVCzJhUnRuZRzlTYc6kTRQ2sM2V7oulDN9n2KAFjO+WK
QUE/onc8IZllNsc3YCQT7+X4pOOB5zNbtaORBE5e7TrhMKEzncnBPbg9OYLKo3j5nJ2cjL3Qd+uf
++L1pGzH1feOnvoQK4ojW9wVUuhWrEmnUdxaqZd5grOdWhBKwfLeOMVoiP2W4koS+zrIr0UdGKax
ZFoqxzI2sDlZQXsH8ckmQ9inxDlZdLzcpdN9ANds9oneLV/3pTKufMMB/voAW6gJeCUgrdz3aLc0
Xua1iDtPIjk3uPlNlXk1Sjflf/S2rjMb8wKFuONmZUiB3/z60+qpNehg2G16d4recy9pKJEINxml
M2LoWh7xbGmbftqPT/QXNhKZ+6OidenF7+7NVjabufPWfQPkrK7UEL4T7ZXPxWAAFwG1/0WoUDox
2JLxBd4b59u3nRU6Xinuip3War5+zVYL9jkvMrIJf6QaXm8D5mWLbmSAGrprMyHNQ7dRo7JIUnuz
SGutibSf5lqrNlbz61lJdfQq6ZLxX6gFBu7CpOp9IdN46mcYDH3OxmDTY4WqRtrzGp483LvTDZiq
SsVcar6ORe5MYrjkTRYlS7VNTagI+svvkOGPAIu1Ukou8VxZFcNWsSbt3bALLk/fLG5WZ0IUlWq3
pVwSuve4kbjJwB0jfDnyYVuRwlqDRYe6Q9163iHEEBJOK5aLut4eeQ2TSEYFQl6P7DM5p1wh36n6
MG2ye8WKn76VCq+7Ze2Fsg1MMOjd2wtPTOKWqB6baO+OnBNRYi/rYLLz3o3OZJ6w4y7FO9VeNnCV
/BgbiSppskUhILczKwMrWOMA6dBjqeD4V622o7t41EUsqo+yy+v4WftjanvMe0/u8+w7qCSduGyX
M+wt7zlP4PmX1sKYsqnkgo3WVouxYQEZwxWPvEEIVCGhw23s/kf+XoXuEKhCmjnLIwO/Th0dm8gK
2UnuKHeZVEpUJsoJOrzw/eCXPnSE+liAMwu92gDo1LY9t1GqhRl4rn3W1ZODZOxyo+uFD368X5qU
RSNET/wZuhpQKwlH91f88y/LGanrEToQRBc6yLU4yf0uE8xyO8bZCTD3cScvOcdds47Jys5Vq+OE
n8rt0cyzfvnuCNV2cg2nUXQ77PhDj+9hoBoqvqx3TMkxqId1Y3IGyq3uMa4kvLbg/dJ9oOf1qLv9
z4MV4+8RjVO6tScrOp5lxeUA3Euzcpn7+JpbI23I3rbjrjBBpYwhMl9/Xw0VaynMTeQN1HJrvIm4
OVeFrKBjlgIcOhXZ2/a+dkeNC3bKBsaffMzUtWrUb8ifNPwLGnzxU9CiV0P5FH1kR65v8yxyCYcu
zjRtE4/KWcUF/eyOdtbaNK1z47XzjZfAcRGN0xGaQ8sxqXYnB6a2c87n7YLt4+V9Na6Opoi+v0bw
dfPtIqQouBJXeJyFJkaFnFT9Vy7k+Tz9oSzCxzRPLVPqlLi1dzyz0a5Gh3liXZlKKqICZspfLTgx
7o8KafQFH8kJR84d3zwJqtwHGS26u3fteok3esBDDkfiJDgBxcPiWfQYbLPcyKgitaD4XnX0Gr8u
tB86oGTW6R/BgqoRejVSIATe7jpLq1/RTQ+8QEINBHZyxXYCm3lA/0JC/LfXiF6H0PytNLOPCvBJ
9ShWQiwEhXeocvmpOTEPoB4eL+9Qx1WX8Oso0/4nsESlWilTt23rG41ZJrnqRYTpdSljsAzlFxF5
K4vw/ZNgwLW2zgf8A5lPn2CFRRaz0fkYYzhR0XkEUWIcl5mLe2IqkBjLxrvn0JzxFMd7J5UgrZb4
uwOBOqB3XnzuwNbJCd9YQOqC+MmYaImCzuBEpncpFb1Bs1P+vhhg4RwNf728HJfoRAoyzI3IPaqw
ZcUrZmACsUXTwI0O21aCDfbehfOGhG4+/9sVFvWoLsJArQ4AMrxhPMmK+vXtxC1P6n/SsZ2euryD
zhL68tFz+Sk1l43v8JTAydV/aDv33EPR8JjPirui3m2LQbZvQ93topPZEoI0542FE1TxL/bPXdsD
gu9aSPNyBmm270oszp0ROZ5RB4rMKLTAz4AuQ6bKWcTRU2GTyhzBncOuglsOc84JlFGTRTNi5eK5
SBYgw1agfFh5+ZVMw1nt7KrBrWADTkhB0k1IFUH8oDCCTz6LpBoSljYZPugwKHxSctmFoUC1cyUA
Mq7f9kLNiQT6tNmguPu4JEYC0w3cWiIE+jsQvTTdGvuZgJvgGZniiM+t+K56KRiYisE+5j/Za9Xv
5OGgKW7hX+N1SyGzbhwaw9twsh0mZqXtqW2DLrsVlW3ibcgiB5YWJsTFcZPv8GfQYmsLb3enP5jA
BUhu1fp8xEaWRtD/+9dDEmBcBS1xW9NKHj4Iwxo3Mn/RlQAzK5ZlmNfccgAqZ4dfSTLU/cqmcEi2
x0DBHTuOAvnNycwbHJBSG40v1+KioniTocvgQjO+n/gKWLLqZlSds9qMcbnD7zfLKsRl0KC+JCSo
kMXJZmfh1gPcDSvzDn8JZjKFcOnaWDMEDGsFd11BbdmM2fTRpepYnmhP/Dx/PmGqPegvtjm2gp/U
I6R3sEAv36neZRJknOC+X05SIQJ2xXOzirzTlREMvvIzr785ZfUrb7MwJ0ZdDB27RmS27rbhCQyg
C6C5koRptOoZgWATmhlc+5z2Qv0quOAW5teh5jWCYVvfWCUvDfjHWMqgtVns/hwPgYuXyjcmPDTE
TK6VHgPhOhjHNJieJ+5mgpaXd40nd41aJ6K+H4wFkCPXL4b/XUhL3gobw8DuQgQN+oX7SyfbVD4Q
Fr0c408l7t+Z13vNCWptXfAo85yZKda1Ilx32spsCoVO3ykgaCl/FvOfJsgH+KrNAT/jftHtqut2
mhVdQ/SI1ALP6gD43iNLL+VPONt/aOhTZ/bxc2lAz2lmGTceOf8TWrBDLansUiDIiNjJ+ckiHtT2
YfV/QTgd1o8uYZPYdjzrUNHh18S+BmBkX73v91by0JVnyFfeDW45yuP1RB3WAjjl4EHnh3ntFWTO
YGsIENfWZX5SIP3qazjU51nfnpoZao8PYNY8roQJwSYHCrRHgpm9cnOVaDPLORNN5qhxZ+LOZZum
QzPUAlRf3FSsP/+5bFiRZO/eMXNzWsJvJBxJIPspiGKtqXuz6YozMLPOM8dANaURfM1yd1kSIiUd
AZXdl0j96SmABjTAb3j6axA/xuFCGHtzn/7WZ8NI6GKYM43sPAubwdccslEaJdbviJ6pnanMof7j
9WqT+zv0OKSAN2D40F5J1/KNHPBKNddTaosho7NKmFJ2t+OVgH8lVeCJbwi8hF76J3t09h20zXnD
QrjN6uFZ5iKfjlDeT2NQbyrigLh0iEn5QR175M2mwTDrncvx+tufutJF5cdWoe0tUGLUQJnxJIgY
Y9mskqrpc/fYasUaox+mhmgLjosrwo0goUdQX8EGxpelRul8JNwRELW64Ls+o9m9wL5mA05qVfYr
rRdVTVjJh8o8DPWCbVQwekBoDfKAjjZGbFvsOEHWfG9oxm+b6svXbKSV/7IIImcu1DZGQfUfNEDf
xTYe53gl8OOOHa582jQchDqHYnbLhy7rOvKt2OqiH5ldVFtzkzTGrmhtXbWZ+ZQre7DbbPijwYKN
Nv+2O6YuXnNyU9as/UB0EUtVMTov+34T5z+lo4VXHjVOLw8sYC0S+HG5vyQsQfhYlD2J2S4dRQJS
Mw8DYFfrZu0w4ZF7qEmq4WKtDOU45kRXFMmxgd5x2ywqPiwWfG3Aqq1RP6Ry3Zu6cEdrRFlp5L4C
VoEj7LewqqzGMvP5+9POR4aLw++53AAUOVzDnsAnhULSKz4KiXi1/x0DlFn3m0zEEh99TLytpdeF
wJElxAcaJLCABBAtUsoE6FCa3P2TFfHBcAhnYxHsD5E5GQazP4ksJvslbnalutMBEE0GE8m4PQnz
GskJqMdtio2YVn17tVtzbTaCgoRou+/xrKb48ixTaKBZiASTv4Z+uvwp5cBLzp9SDy9aOBJ369pe
fjBVAXS15OJ340jncmRp50L9hq0FULv4OavGZ4E/03/Dl7SFh0xwe3Xp3um1aLAaaDqDA4sYzm3D
3Rjksd5cccWa+Pxk+eKhebj4Et2loIsBnsE8Jx1r3WDdIQNjy74g9acW9p5gf83YGSYHMlPqSwHr
/LDuG1LRrihyHInaX3tat7oAUJx5NmUcO07hQ/GrkhfvR2VQko8fIoaBq7J2o1iNg7R6/jvXdm3x
jtxK61T8x6oYJTqts3Lsg7dhpNqYSHTjgmV3vsc4GXBqwSE1C2IacEdGeUzeymJbddVCeUyBF5i4
SsG2VzzblWxwoPCO5cvYPtgspjIRMrJmBqZdHXRfQcbCqaTkNC/NEpMKUOIcVnn4TSU4Cnxka1kD
ZwieT3TdCtuSatdUu9b/ImT8+kIsh2j3h+p/rmLLrqmivNOIlpNO9HQc5VdllbnM94oRtFcyer2e
r8zK3RQIeuS9Y5rhQXeWWKN8hQPb7mdjylo3+HYonh/NbyMk28FGPs/ddXcLC15gv95eEw8FCt+z
HfZW8BmIGQB9mgjHxt1WaXiehFEKfZYOhdn4+jVoi2nMtZ7JubTQq15w/S5TdamXDYGCSimPFF5H
nktlPqsySXzhEA9bqfFme2+ZhCtkHz3EOtK7piHWqoEWgK2rj78IZtY2xuuV6kKPZikhhV3Dj6oA
Ll7RIxwmrXvDQYBGIXhumDVAaU6vp7zuUznbEgakorFsZpmXfHjh5zvmBm/3qIUEAqphgIJuYC7M
YBl4iHHIJy3OzUTsEmYcIc1674tmNLBR+WFl5YPigc0vOTPjcEovTJwrJ7trPd5gFZsYBkJ/0a4V
/WXYyH3IMA23SRVi5J7WZkd32mJNxhbvgxN4tZdMTl7/xO53bMexnAW3715uACVU+zGmfnrzh53A
sCRmBIYlwGVnKGRj5FEm2KRcOU1oZQRVsnKBIVdaXvXTs7z43Vy6b8sIOtm9HwHMaGP1UZwZIg3s
KiOr0C5NWHI8igzfrGTnun6UjRpv58cJs/e8CwL+yRV3NEV9cmf4qGZPIHbJewRGhaNXnj617KA0
BNE1TlN2yWK5uzL+6D5viaCbLbSdu8qY+0rEhhKZFO2BVzLyphtacNj7ja3honvgfiArk0WQbgit
I7L801RhG+p3JCadX6q0A2KE0c1fSyqnXNHPgeSQtC98SalqpHkHVMWYymAM7fnFXj49OamoEQy3
gC+JuN3Ldvo1HKV2tzwcJJ56f/W1SgX1TlsJQSLt6FPdVtbiyEE/y8oKzRVhkvcOxrNCsgY2PRJt
0YMvMEowrTkOgeX1/iXsy7n3Z2DnuKH0jyOuuoZZ2CggnM3/NbbmV5z2BtENR7WXatRbQ67Me9aL
JWRVNCfqHkbCydobQ2fd3zPtacIX65yDptQOZLzDjbocTvXdn0WLeT7JIW8Qzp+R6Ia08jttDiWM
XWtlOll6iuxDwGQEufnmT7iImo16tG8YnW8FxKIFbmE7m805jFlG61uyU8wG7Mpwj5agE45QTSef
KJ676Q7xchYsl08Ci2P1OONzBIFMpwpaIan2lvf/Go+X8/33vRY3D01Y8A+tiBRJxra6w09BtEjj
/38QoiEfQsAWcDDHoYE20wfiio9XtiHE0iOfJRv4cFFgt3ZvGfjak2E4qNPEmxMBJo9wQx1mCkOQ
l6gKJcaaTTG6vM2u2OfrdwyCd5pJesEnywN8J9CZXFYqJiqKdna3VSGgKFs6+s512Ca+J+/MLMC0
8QOZeDjvK4oMI6eZq8JxoZLXlJ2rD6F96zxncUrHlBMmZdb0eoA917n4wg3i2iyfxZe1IV5SGwU/
f1OJdoK1GcxkPnC+PXO6uTOZ6IG+Oh47l4giWnDJbZGOD1ULjSrS8oFEkgq1d33dDGtU6pHKonyh
DlsdnAMOowQiMjKTN+LFAmaW2LkJcKKvJ34rdhP9Z8kueiSaW29ge1+JT137LgaxlcqtYQuOQcDA
yKyVJuq3PNguMEO7tsZqO/zatj5GhVcnWhdDadxQ3xA+xhJQsTSrUE4oy0rvvj+/JtkumL19DYTo
NfR1aORO0CHL3l58AQBqyM2f+EhVTxxkkuuMDoCZ9D7gds8bKEV37B69xBdTNX9zkBtwwd5/YEgi
8/YZdNZqUTDLAh3OXwPMyk4BxDrjZzD5dzhiba76VqkuOMplSS0VJ3TeMZNuiV1Z2T1RYaL6wLOg
QQLJlWtIsV4muOOnjRVEE/X5IFRlWg+zFpc6/ql75HrBizA34uJ5bXm3F0XW+lD33veuhZcvK3Nb
Mw1EgR1eHC2d8GomFdliJz9+olcaGvK3uSn96N2fGHJy1jURP7tdkJsxGR1w5BVTJkvXvz+bN4G3
FvJycdj+tUx/d5B4ZHNVdyoPOd73L+oBGbagahwL4QHocEmJcJcY0wB/rgvzxcQ9ANUSoSYogMNH
vv7M7fLFqkonR2AyMj4YZ6JBLfwwbnS3TdG4PQQZDgoSF2lEkIHJ1YRK6Bk7FKmJj5wfgzhOHy97
hisG0meRocQvg1ovGsQHpNWTJL4YpmdnIawRfk+khe0Ei09jAJSM0/l7IIWD59pz2IXP7Tn6oITV
zORZ2PZ4MZsOzmc5zwTJZdsWV5ykS14PDj7QvNK4eiv2xbXh8CwavscuYjwYvpUMlNBqlRRS/iVr
pchMFLLj/jdD3Y8zyaRoRe+TacRqDH08IPu+nMPdPGCxMyaDVcDYSAMoKwh7uTgC7oAooyDiHHgy
LaKLD/Y4nFKicUWvwBVd6OKzaiY/mBsgXaKIMtKv8n37Pu52v/HJHib6FbnrL8QkbTuBzoX6k4+Z
XQfJrYfRSDrlmFJoujzp/Zritegq7ZTqM15oU+iEiw1C/JILQF9vFcQC9xCdVAll64Or7ewItdJ9
nmovLkFGkt8/mHVvZGVRFl+r+3jJHT6H5j12xuN0yYz31Pfv9EM2TaGEgsPC6O4aAeF9DXsALakd
CZ7iCxPbGooXJd30S0WMJwAVqKnuqJLgZEzQX26RVTDOLTkv2OnSA8eLhL6ctKXeAR+0Gj6JRtBH
Y05KuZ+AQ64eXSYEBg2xMy+alLeKGEd+auRRivF4vT26UjMrLtrketUs9qstGkfPQmsGwxHVziKc
7c5tip8AVDIs6xE6sUjYm0L04KaRNRuDQ2NlkYiFp2lOSFR4tTXESNoLRH6dxzpRPMhfbs6k4nFg
FCqPjPt5dq3aliRPL0ACIo4GNDVmDWOkSLqGWn05oTUI0GIomGyaJ6nJbuhnltn4A1CUFai9ZK9K
1wH4gS5rg974+YRhJ7JhPN5BXlJXlvLJ6IORGP36E+v7wXX6t8JbqvgWGODkfrbE0Zi8U60iEfqt
BNbbf1HJ4iUZNcHeA5aP98dgFlXNJdtzdFyM/QXkOrryeDaAeBbLfDkoPeqGvCZZwLVe21P7vL5B
M34Yia/Qam1A62/dlre5Bw1LsQncLRihFpMLCX7Rqf65Ve2CngRtyJG4PkVAHjNqJYqpPtpiLufF
YIlx5t54SgB1iSQvUW3gjNfvz5bshn/aBfrWNzP4xlUilStyDuxpYSR6IxVtkAE2ZkF+8xooh4yk
LB8d76TjmQZXyMfzHX73Cfp89sXdIMkkMagXGxGZNVbNEZTRzsNrnZnxhnxP6UngBKpkvzvIspqP
tSJXWwgSSSUbeKPiKzocsvF6MmeTwN72bdwoe5NDxEmdnAzmoOwPdyz/WP5wXNGZSOsiX+LDFlRM
UMljPbPuAu3JllvOZpfqiAJWKIrJWyFrA11KnKab7IkPEuv+USDLISnzyCog6jlQ9XIIWYRPGZuP
SHHFaNjPg+pzd0ZsOUkNvoo8fWNoAOa4k+zGP1jhiY0gy06XcxfN78agDPYiqPyMOkAQudIdjKmg
1LX1lDOhoU51ecQ7Ywu+tviLdpY0LU9gDEd9xr1/ctcxTXq1SB4pMXQ5aZ/NRbJ7zDKCwMIJU6TD
NSlxzsuqlerEbBrxfXFuNPZV2bVIuQrjhkGOp2WfanPDGM6zMTvGn4EDnIEUPCk+eftQX1Ru4Mkl
t7iEvypGHQRavEpUJ0xKNaZn9s9lVBFFAWh7dmS0Fe3CLidU2eH3brkU4fOQtv3lwkpmzpPTJ3h3
kUaOh6khTo5ccU88DApxEcdTFti7r2Yg+Kp3yz3UWdHWQaNryCadF/H2fsUx0zNvBmHr/PcEst6w
LbIgLpszq74mpUrOZrqwvU0ARyNITnYTleIaZ6P/WCCUY5Wfor35h4NUGmtikfNrzBozJIXcJoW7
wGuY1irMFndfGWPr4hgn9Ugz3nax/BsurQNnUf0DGUvSEAXI+ReriKmAaq5aq+kVjhA8UXaumMeC
xr3Lf1uTmye3kBK3zoePfNCa93x2eBjyhJHHuKbWDG16YQnWWAQgZzkENbmMDeBjaOBwb4OhGvpW
O6u4xRaAAmoW0xEKy1CzgBbRbVoHgqG2wt6S6xHSZM6xmaYt8HBl5qwALFm5j8FYTnn9qBr/yaKu
euyb103D8tOlyHefd0pa8UcYqmc68s0e21yx5UUJyp/eCNPwIef6kKwjC0OVCwrLd+E4ILCTO/lK
Muq2QpBG/0IaMTOR5VpopaiLbnrlgFsQ8gbk+JsH/V7P0v0sWBWP5VijupnXNQTMyA4dUEHYEVAN
bcihxa3KuJfB/yjoGECnx8UyIsRmdEB4uqX8VBOtyjlDfdDV1eWItsuKzhWooF1bZi/OWoCbgFaU
khBIrqlYwgpezLslWsdEL4e/E5EftM2ZCKwWA6yyn/e8osw6iFAaXLv3Tg9arRXWDzKBcODo2YjK
W/BlLDzlcFYAYxOqFpIvt6XkMix252g42D4SIujbypKlDLVhTv2rAQRf/P0J0PEfcNbH3WGyFyhx
Ww3McuBXKIxhktJXMjw7mWeFw4aOLz+ydMOTpl3/RVfLBiMhO4JTMGiBgFHSjID3Clntv0BrjWn8
8C5nsZMk8Xef4o6/uUiPrxMBqQRyCftUXQpfMT15U0JghYo8pIcxQmT9Y74Ja9EpK59bVz4AeNES
ck/Lw72wOcXi0OBRaQkAN7bYFK7OH5jqLFMWvN59y2SPK6bi1FIo4S1H8ZY8EgGxxjlqcOuV+AwB
htNrygWW9fp9E4xpoLlLsq5Jd6kzsaZgdwuty6vQYkk5anSbGP46DtYBk7fZ07/wrgwKNbVZp6ik
hIasoUmH1QCx1mGe0YNdOcCHbNF0ScB3aXBxEJPmn6JTcBsK8lxcCzu38pk2w8ZrGUGDNQaFNeaq
A/H1oHTryZ9ptzDp0WHjavbjw+zRyo9XEXNqQomxhqLsOC0icdqlNg/IMaFmZqQjfBdq8T7tiMys
L9y27JjSQEXtmh01/nx+i71jc9smIPLcPbzw6AyfmtjcwSPmowcIrgnwRuQCMxLr3iLLuOEBi/oH
tX51dSZExMVhvgkDpujU7VKPTT52mnc6x0bKFBIg/IYCyrGl4pE/wflMgh5wWl/qkGLzQZXGyr7n
5Bymr7E7Kxmu8+5YBj22kP8+G1IPH/np/bAQp42J1zb7akZwURoD/gZy0EGlaDLAUjzuvNgk1BkZ
yol53qlC5C0g4UDGfgPpT6NDt83Ywc1IwdAoMBqPI/5fHqhpHHFjcwo81JxDNdbmLfzlQo70Zo7B
l8uuE7WtviRCS1ETUAsTLvojHBNfGwY2aheiuWnPVnYY1fOYO2b9uFw98nj9azyrbt/M0E73e6Gv
cH8rahd699qLodG8o2eeJ/4vsSpaC+56JFIkAtsUbezWnmZ721o7gXWHTqqKXscXNhBVTpJcD+hb
xR3FvdazYCAzXsm0P2L9mFp7FLuGb/my7Wu64d6eBohK6vf8HEywyIo+26uWkYx0+e4yvQntzUt4
GuKn2CnnuEINYH1j+qWAJPOgw6TDyyS7Iw5qxypEVIaoa/doLWbvVtqJUH7qp0JhA9iliqxt/KDj
TotOx5KI+sDV7mawIrNcQqaD1Lu5HdUvNaBZalEw5pSkI0CwwZu9pgrtvsRy7tI90np5DGIOFeUw
L/Vz8O9qMRMY3KzFh28kS9TGWPEeWz47hsryXibzSeIe20uvE73z054DHnRQRBAYwcnzmMC04mSX
4BwVcoXvCL2SnFOjl/+26gba5YJfI8F3gRzcUJAAzsHyNyDy+/LTEyTYYN8VKk74O1QaLOy7CRZW
3+u9+NkH1/lOIxNA+xUtS/hGOmCn9l9n9G2YFBqgC80PCFiIReuy0QZuBNek76ShOsutoJn0Wt7+
qm/Ox9X0YD5gUkXStXDj+3vqJSKr4d/M+Or1hPA58KaXabP/lttCaZi7mqsR7uY7gCQVi7+jQZNc
IUE5CHmzaWB2+Foh+viqk1upgqs9wINKU23tGrCXNugtOquUxFsfM+bVGRR6AAEVlIzXatauL0n6
ykA3XxaxJ8QgoZfRBz0q7ReO4DK7sQlkIC3nhcCbRCUYDNMpPFcwJZWIYAgwINum9ucU7EKY61Oy
rlqxZGtdFvoDUWJqgbD7Tv2qZIJ9435oOjY67mKa3J7UdyRogi99ymfHRVjl025XkWpQcnYC5ImN
Ppgn5BFe96e7zxV+tyomzFu+5eIhXg/ItMrDVcjejF3TSqc7EXA2vYLcVFZzmOtTFt3ivBMyE9R6
NCcq4DRfVDg9BWPa8jrtpO61iStaP8CFNFFyzF/TWGxKDpJj036VaCTh68peoFnS4e0f7K1NC9oi
SCogDbQ7BuHik6ZYCubpExM6+ydaGZMfM5eA6EpZef15DIDd8CI2+wffG4byxYucXkAtDtGukVNb
OEPa7OBSyRv9GD05Lh1ojwnBP5RIr8IOqNHvt0CC/tpTRg/MHkLLWWetzDplpqZQ+3THtnvr9vUD
51b5RgKR2zXmY7QiIQS4yBoQqAUlD2Chs1j0d05hF/3g+JBkBugTbyV46J0D1VF8FcxrIhstfAu0
6m23DMrV2Yxw7/HHXM211SPAl39exmYlzJOy9ltknTbw4KuSOGYfu1zO1p4w+m9RPelUMAyoUIZN
RL6qBJIK7BaA2IQtn0fRr3IBRTyXpiYBON9Mbn/onv4IE/MuuqvidU6A0Jhf3KGuHtTKin/vPAAh
pPeheNcNpDtsigtBTwcXAcc5QyMwDZyWKXG9qguXmCqBE3tln3iIs9nSF24wqfEVGO+NkflUYorD
A0JRE7dJOturuqvS9n7SUZZ2AEkA/uIx3O/hCFWqYffbsTUFdA/7uBLE8oPg4OooQwH6H8f3Qrvx
zKNRj8d/cMoJre4K79CwZSVk5wu4Crirn89Ihxf6/F1lasaEVVPUZyqRy/UXFXkYRh6M9CXxm74g
0I97ZH41V0RK2QDM8ZDoOC9yYGqfXyJ5uwjP30xs0QJMVbCRsRewuzG/m2jhTgB1nQR38rClyO1s
E3vu3mLrBybKm8LXEWqR7FVFyz6vZ+uL+J8WiwfPAxEoVmA+eUazdI71MrcsZAxOamhl4LF4Fxxd
6Ghm5E1E5iX1lPGziCNBHl7N5Jgefd7nY7tEd96msYK6jZKKeurdLleD6hpWnPj+lv5PBPiuVBMi
Fd58NhepmhEhE/dvMssCSQmxGhIeclUgv4Ou2D7Y8+KHqpRFvCVGMbKvVcjA7lxMqZmObYKxe6a8
kSD+3YrQw/JMCoqfZnSVWmaJ9Um59mqXPsXq5eBHOdX21cV7Exo99xxWxeKUu7XgSmixOfclfLXp
vtrO1VjmhANSu/TayFJVtmLqmXpvsRuIgQJN3BxIsGZXDAVox0ugivl3xxhJRSh1VkcbBdLvGNvo
cMdLmAqrDNCJK/mFj9rOLK9fqE+XvTkIy7Q9rlNrle4/2apkJzO3TDi8HIPqel/CjwA4I1IxumBX
BFzJvNcCnPmFiVtGg1NdOHsbtwZ44dZO03kcIUCpyZS717vB4CZTooRHsxrsKpsVnGI1jX0qG79o
LNolMqNqmnIspbnTY61+jP1W4W7kxpX2zTVykcSATXLafhP7Z5e6LM26XlRC0HLWLnzLz6v2DBsf
r7MQyo59Cgd+MOZ/IdSBaUqV++hutgO93CEjUUBTjX3JmzX9Itv2YC/0mKbNnddFnXEI8tR0tmz7
Wwj5Bo7OtyiMJLw2QY3dST1Sf6nWTuxo4Pv+nNZvXahDerWwQTwb+/+pCGBAin5ltn7p33HHpI9p
T3ix4QBs0yU0m/Cmsb9VpzaqET8hSGVcZITIbH/e3T56mksEdxp6JHjpeeEy0R0gJR7kOsVS0fU6
qPuRF8F56yLjTbReNKfyh6hjFoQCkfJ5mxiUCRrgmx6/P1HKD2usBDHvz3lDHSAd4BITCsyiwWsa
opJeO74AJZU1xT8wl38/mIcU+3NN+FSB+v7R5PifxHyZ9zyfmCbn1+xnfoXbP9PWrNzq8HspRenr
/HBSJeS2tdhV0GRflxxbmrcNbsGsbpqmG8ADw0byQYKXcZYuuWNwuMSycpc4inMBDlMXgwR3S3o7
rmzJCWvD1jt34D1X8WrjgN+eG2FvxEvqzW+kiDAp6BI2GqBIGHtXkiAYyr78r2giNyLJDI0K/TCG
yd537Ojy0wDwtgFpCpAByZj/KA2mslUDDrFBvZ3xFP1iVmai/JKom63rInvb4/p8zOwdOIYBvDGm
iUNgQUQv3YaMNFJ/SbiVXI1j75uni425t41P7tCklAp2RZSEnwyKFReRt2cp7LYZmhBI49ScUv5T
d2YR7M6++5wOM6xupwUSyBoHlZe6W9d2Y10mffDT8rvy8PXPfQD6ijQPoS9LMLxmczBOsWJj8o4X
FwbXHHvB2VgpR/GsswBuZzVeZPmNRmA7orhTyPQ7nDBGnH5I9FhZ+DtA4GnnH+btBKnF0zseKZfL
biEG8EAjYjFOwLmplnVbIEmj73Wt3iDXMR0t/StC1oT3067zFjIjSbWKPSO5yCSjBpTDYfGbBjxf
eJDKDZ1nVRsRLRKgsFgzaX/IPXjJWYtMuR+JN6Kp9GkPwkj209S1tCJCOdRKcjWUFTt8B9CfFPiI
uyIU84MUkCE9Nf6GMfgCKxzYaOxrVijavJmK1nEanhOSOYecj0K4y0BSVs+YjigqYp136ctlpd/d
Pp/ZoR0A+8iQ9+3YxiTt8Ux1RAEUJzJwLMcTRf3pF2TI3VNYFWGrLU7NnFdAmnY++xe4MbhxKp/H
MaTeS5iExuQBCmxRkCylA2IL60AG48ge+jLQwoFVPGk1bkdq+ZXxZX12unylcNYuLDnibeP9tt1F
WXNlBt8SKaUOOonBwITIgoZOeU6hfDmGHMxhy04tK0bfjCmbSVo3ix8AK3vPV0lECqepsfwdGT6l
FUcpKNozsLrSolWbU6YhhaMbyPxQTzF/1SDRY9O2dyPByhjKPKQ1h3gkklMZqwauUn22vQsefOd3
v+WtKHmGy4w6bYo+5kD8qAvlWeKmkqnAIcK3c/5s0hZcdGYn7E0BoV6j8bp2Kuqv7dwQC00wfyAg
j7GQI4Bq8cS9Kk42IKYQJ6pAMDplclA647vMq144CQ7psP9LWF7hldXznAS6Iz++HdqvF8Uy9ajQ
gK35r6pEyX4VeThFz9oezAgi/rc8AbPgE3/1RNqaG6b1ayr0aM3xQDI4tCh7HkFRV9qA1sX68MFT
QamZuKSXPzZM8wpqSaVCxUW2IHYoT/xQDkhr03tq47PRKj4yp/x4nQi1QImrJhypoY9pvu7iwD7x
AkdLweluJu3yU9WeD9VZDlDZ0r3oKec8YWzfa3Xr/4Dapeju+cvEOCIDRLVsDQ85L09aX3q1I7DC
PT7iOXKneWxfkasX09Red/7LmRR9VvAMxxiodVrnfwUee4SsSFtLRc4ZzXmSevff/vyGvj/xaUni
B2EEQMZOMkvCKmnOifzdgBqsbekvZ0ZT2GAPSz28KZr0QuKou2vnnFwbT9DiT6lHNgcS2fIEVTXd
le2PXU4hIrjY8/PzRRvqFuHpe8cIO8MlWCvgqmdX6V8b4LjKxCXaWKNxkDxxLkDe5xqB4UX4G6F3
N9bz71JiAc6HhFoaQ/ehrR34qC6nCN4mBdgDOkjOanUieYPefeJoa6lylRXTr/9tvYWVmG2H6KwT
8q4B2xM3dMZyDhdJBbzOcQ52LamNP8UfnFr+/YyggGcgQrleNK/K8Movua5o7m1EYSdXtR5qmW9t
2+Y63sqpEt2irWmmN6+waAUT92MDZZHvXk89s4wvRDXB8WSgvRLuAedWQ8IB8Y9ho+Wt6TVyzlBk
BYS4kHaCA8eC5DCLXoSo7m0Syw61aBmMq8esBx/ecdyVsbZRmkRIeY86jJG5PBJqJSowAamk7D/T
1OdKUxtVHUokFRhH4FTNpJfBkgVWRaf4c2ecDHTfwyHb/F88AlYElP08v5M5Ja46mHmOcBRXZ4FY
89Poz+NMGZNUB5mVTspPPNV8bVmeXE+9SMC3Ah8UuUkyXBVO+6cwMSPjurBvHjUevRFxBdWN/1l3
wsa2tZLKR0E8kmiInygjpitsbFpiglmAXa/Yv7Y+mazFRi2P00mDh0iVw8yeWfSdBekulB/jQP2x
1+62ZJFl03rvLqiguWMHQypi3v7cLJZeUXUvKf0eFn8Sz11Yk4P0CZTulNUG91unlPTcU1vqD3t6
aavTJnyZBP9kUIp9jdXXzH7T2yBuGwNg+D72ZslmpwiFofA3pZ+g1oOWTydYtwwSubTvMUNKl4N5
QNqCCtirmUFnyx7n745IJjz98c+AY1F2pAu3fP1m4yBx2RDevQEizzLsTr5BY6RakAfVSMQAzyEd
3aWmcbrGTzcX5CKGc9b6ZDYh9JTP0mKRxeW4xETc3K3YwZDj2iJljwwMmi0epcCXw1n1Oh3Z9MSS
aRU6WbyS9ZfiXtEUsYLl3Qd8LWLPAS05UP3pZfwviHH2xnWBKlw8FiWUj7kg+93I2eLsMI5jKJHx
UR1goGw3Sc+si18MK76XGxuo+jYQwcLRYhjQCZYQu4GEXqaNv4K21ZNMZNlYH1YgS/C+kQehfnVW
ngm8C0XwOP36lQQLhNR+jT3IIsySA9bLTwFqmM9OGXKYhgqGpfHcv2p1mx2g3+Qd/Fzpw6jPc85K
j9XDpheW8pkMCf3DKX18b16dVGbu6Tp0Y6zJTjRKJuaWBaOLGTvhSQaiFEBNmu1YzVKlnbrpsmZr
zp9RPVMYWp9WDHvaS2vJ1qjTZJFYnZGPzBQ6neMBuVirGSgK6aETUIIROyLnQbwjcwUVwvaQd6jg
vsqKcVfPI2fVOYcwqveWqzbtOwoN8ZTmJGJlaIZdCMMsSF4noSoIbHpve13Iq2153qM3JeeESQm1
FfW4IZgHatPPH5u/FNB16+epPy/aEpjUWCdDKnG7VzUT5DcwMt0ob5kjZvUexxOpaPXljY+xsn0i
dk3e10NLdd7OfqnYD0/Lj2mITY5bq7EOAqdl/r/Fo9n8guPQPDkmrObVg6h3VedfyfukEZjdqBlH
+dU90e49qkaDxeVeu8mTjo81FLKKdPikRy79DokaC/qSv6Ud556zAKwD5HR1prlpP7rgHD36epdX
WS0JONwI/GFbTZ1O80gbiYSQNiSwUwdwYyxwGP29/KNpQvQ7l7RCBYYReFlRowFdN9CCOjV8JX/x
0MtfiOvTRkXcG7s3pKC1GRnUCjUlAjbVuN+9yNbRpN43NWynwuTJmYd6XM9MHCRM6g4y5JR+5v1w
gbTr2nERi4CrQm+XVldlQpCmeGQBJkHWfyEXb5yHq/6EQEMXFmkzFeXX6POYRAdaA3C2wgrbPrmG
zRFGVFgmp1zsQIW6wN8QKdNCqDuH+kwMwfdC2dyaO+TPXjYK6N0GlX6ZO3MAFbL52qvmzilZxH/t
DcZLVscPhXLQDjOXpcodX3IDIi2Eo1iv3d/sdsVCHGJC09v7/+0R8oJA4XFbFgOi+pkMTk6Dkelk
x5gQTNplEBZid0vOtrjWbp4C9VUcY/0Rvu/bmF8O0dk1Y4fldNbl/pdgJSDIZ3MUT9lzdvQ4X6Ki
5SiEhuyCTZYLjoGLeNfYvVK3KfRObSOFoSLqI1/zNIzCNcXOhFKrca+cxfFnUk/47fE46LRvUO0B
booNhNkQAYScf2SRgIc9VZqweulez0zFV5ZaPxwQTd2Jh0mNPvrXqLhcYA5QxE5d2mEF9YB95pqs
G5FnVd/tgU7AQqWwJjmjOv3Uqzftz6amUqdHsEZELeK5mBk/e4ombVScgh5hYX+jvf8vfnkYtP38
0dEpfaFQJWSax0xcM6N4/I1K/L+dj2is6OLTi7Bxd7CCQrbMSdB8ZLXs891n+ekyhbD/JCBdbHVn
QoBufc+W30J5T0H91SUUmjGmWadcR67F83js7q/MtGeigAXPUr+C0NglFhFOSAY4wLv4nTbChAnx
GLlgPOH1DL/6sV5TLKlLKg5ioOUc9LF6H1/QZv8KK6JAQ78JeLsKpLZ7goMLE91TzqvaCKy+sviF
D5QD+DKG/BoQW8kQSTfK9kcALEnga485FS8zwZ6YzcoV3AU1WNwExsOrSDtXQAbp6/qHvjTvaGov
/V/tDgAjM9W/qxGuXJlELoqQ1ThcCN3dr/usQG4Evs5BavGRjbCo77sEeOIMTjPrNxPRn1mynA7Q
UBxhCXmcjE6ws5o8rmlPOOfuT+vRILmy045DmxVDd/ofZvBelu+TTV0VFDikefPv3bZ19345r4Ev
k5VW1iR2X2aIefyrziub6gb0Jqe4kqG89GkPwWYbFOxN/AFnuToFYbitmKEDYrsG8XTbOTuGX97n
GBc/2UskoYrpXn9wQ7buuLBhhLhym1kI4bry9b2b9B1b4ioFwAxxnAsEiFpuJz1oaVctGBpybn3U
nipzH0X3ViP6Xdi8WdV3G4H5waU+X41B3n4PFg7MgK04+1rHeFm5x/7ToWGbRyuKMzuNKWPjs9Aa
DoJFbCQZPWvm7F22bhNtnfjj/qA6weLViFx9d9x7ei542SOUPsFGGmWZ5J8WU5UGZ5Wwnq/hatwn
5TdGvLiTxDbbMwghQ9bhFPmHDP+g1U8TM9oZy/NMuE4hrvevwYFKWUlbLtPMsetbUexV4eo7D0bs
44q04awUVEmxZFShrHN1RIVvF0fjnSbWHoI+U8bgdawsKV/vQI4Tn1lT7ooXO22JZ6T/rMMZ5kfy
1JBAFCoDtjGAy9BykboZ2RGRAmmuD9ZQq3lAbgJ7itp+iM4GSXRfLeAIZ8urzM+IOEGbO0mN6FZQ
GOJdL2iBhXqqvJjjO2aAxTXSxJZdV3uTm6b0zDo4+25HQ8N0OlImBR/OylmnqxCXcFOk8sXVbnle
GMmKcxKAxRJ4lTu8ushNjC/uVYdwn1YBrgd9qoxhAaPPL4G0tYaN6X+8xH95Nngn2VSuWthONLT0
9zS/EO3LzY2HZ0X/tNZ5hiLWAF4hqnBXpacvX0gcxdDvna4zO47fnq5Z3Y87zq3Rk+ytd/aXgB/u
JJsNKLtwwQCmKSzUx8JslMu3oXwnA44AMdIDKMZF4onvpoe7ZW/HlVdv4gLyJy88ERZivvkdOfT+
HPSADz0LBcm56q7XmfiA33MUP5UvWWJZ5nLDuJIrX6cs2ZMiB7/B8EZJywjKgNO3lLhxuYhI+Ogy
E950QEOiJEAuLoU4rzTwNKdE4XHQKF5FNHOLcCXdBlZfLQvy76ecghgNGtJXJWyV+ATVvQKVS3lQ
ZeAoCuowT3K8Uve29D5kVCYnjfNCob/z3rLP8HUfKC8OxrtAs4mzkAEajDsz0vWirzSqG3zcQrHB
WL8qGvtAFRc9pJqvkQi4i8fsyY4/kgyln4WlSXLViqU/fgrb0Q1+KlSOEfuA9VJhDuOiac1EiEyn
gVOIgO9bRXTj/56peknz+gxI/IZbvEFU6BIQAI/ebbQ5ghyM4PIWvQgwNfvnXKOTOJ/mDxJRHJDy
eYwXflor7nlFoZm0UINQnvES7EkqoZo9ddX/pz0LZNULP92stwdFb0V9VzH5ps34QZ7qUuUL6Ov4
doLeLML9XyJOOj+aJStFl+e8ayXdODTNtl7+TLmyrcrtbdFptDG7WjolzOVIbq4FM3tOBvBGHtwG
FAKvfcwKNz7TJN7Wvqn1r8RC/eD2fknt5tB90pCxrxMIlNb+oakV7PI18bALhZxeqQ/Col/r3PuA
0w9fP8TEGMd8naBS+sWgorJRaqoULiCtxE2Snd4G8T4GlO/6uVjZle48n368z+md4UKm8DvKUk4b
R/qs/Lu//lf8AfEWUgxkjoRwF5lZyb0SaMLyrIVQJax0mMUyIiot/+Tm2GFHernzUBYZHo15Rq0/
+qXImhm9wbCRVhbZQx2dbYsTLMPxhVQOqZplqbrd9TvsODICIfccF38JmjKaDtCMnYM6L6HAkPaO
GMQjN4FL1dC8dYEET1dufb3ggeQ16tMGf+msSca1k3xKL/WNSpYfnDU88KYaM93Hem3ofN46DfOG
3gnxySP2zsPTLxcOWLBMM3rGrHIw0xyXNBVnPRrN1NGiFGMEQtaVQ7h9OGC4zJwlhV2hhYTJAYds
zmWMsrcEuoI8TD7UVqsd1WEoemJhSoBjWx0N4TiEh2Taa+2H/TawAw8cJK6D/my1TiO5fIpo4SP8
de0C9/2A3ReqSloRAg0DSaRGPJf9LWD4//xoFREBsw7sHl99i81Jqgruh4MzMVc+GjmnmTsFWJnD
J6KYvf1rIWK9ppmf7YXRhIfb4kFC/2unvTHSEaPYI7SSO+fMRrriD1XPx2dCdcvpSxg7Y5rsmCUp
7qGj0oNIWpydP/iib120uIXOr+xGPiUcTppFDD3W6qjp/XwxWx0+MoPMd3EL2iGmUQMLNSvLhiD0
Fe+N4SYT7fgdcOFOaE4A8uA4JGjDXPubXAGX1NjHVxrgUKrtTmbJ9Yqn5VdqHfwO84xlDVLY5u76
NRpx898BbhwH/mqsOh+Ysmnr9KOvrjzIvD6chseMikIceS/sgzbPI42kSqqB4n36Q+Pnin6NpuQe
S9wd3lu/2yU9EbAAacq7pcE7GisRjsdBMvpvw5RzaRE32Xji11rlBdlltk7hRBxy/p79p7nrfCGJ
AwBIB9CBEZ24VZG0MbZqgC5fEdb/CSsjnAXiB+lBHriV2+SkAACne3ELcVDTyoDtR7skbRLujMrp
BhjiAtaDIzabaScgzH3uYSiCDNeFf0xEn3nn2XvqQrDl57CqjInKCr7OgoG955wg2Po+n5YLwdxO
4aYiaixmDbXFMjnXN9LYsWPOTp06gjUnU9MqOAq5EejHZLblTyPg2i3Frz4bH3Qiuj+FopsgX9Vt
6fTLQUJNa8Q7dWiaN3cTOn9ltoeIw1iX4OBOkBp1KaLbPSjzha23PO4vV/TcaG6WB6wIirYKhX/t
ck6HV5zuc1BuYSZBNGDQLv/YHZ70tIK/zd+CvlAWx58pF2QIAidmIYJS5JHoSbf0LQCSApAa01OW
gCWL6S5QXHQ0LBtCjWT3jkf6Add3SlaxzsFi6E0N4A0eWFSupiybUHh/Z+P3Rx+zoK6F2FgsexK5
VJY9QDoeY5kS9Fs0METJMtU0JL7Kq1RLOb5pzmIHXz/2saIXNO0zbv/1vwiWEuVGzzyUyrR3KXvc
PiLHWegnmSF5oi07L0SEStkMtNsKzjWT6sRm2q11kNov06W2XZMNstiICa6407nPiSnLgNGBRER1
lPczFVjT+ZeR9kMHlq4gzH/T6BQvCwjKj1pu6JK5Vj3czQ3j59eHuZNtwAV5NrsSflQN9GCpIglh
VX3IDjrNJ9iTtCxa0zabIIg8lyQ72SMyXxM2GovPLK183ldiVhOzoVA+KkSan5b0j3Cjn4GS9fAZ
dJkFUbYf0YmN9cRQ8jwrpu0ehaN/wRZv1Yc2i3iKECfRYCKqgsYVUYgWhPpu9tg/Mx8qY/QNJEyn
9Ejfv+TgaG15mOYrM0oveXBkYGmBz9lAM6oQ3xc70RynUkOj0BZoIJoDtAKAo0gAbXr/4pv8k9XK
GVEt4ki6XkVanb2Rx+rMdKvAnOoW8a85iUEIco3m8J4gUlEtdF2wV6eTzyNuKWL5f5FaFZPgeWcj
2C8x54702oMqTdbJCw1oTApT7PJ8OAlO/BrQDleFwvWDQTJ3Mo/vXTXzLxZWLlHLHQZ/fVTxKtDm
GM2zVZIK0qvWO8tYVx4JfHR2N/cVfxAg9GJK75hYOdo8xRlDw+zoX2piOfkju0/zMTzp/gbWAi0X
mabe8brYNbEJCB6t5CEjodc/8UUYI8EOVsB+kPBs0BsetB5x6oWoCxJ6Z6JhGW/dLhrLehzVNJ59
G4u5zsrBShl7BInDO2pIzGmlrAuJa8+AV/nd/wVv1w8yEzFMhJBaGlFGLKKOeLp0lTGb+QI+VhLW
CVKWtsDW5yULXcXy0ys5nOs6twIpoj0AifPg6nYm9vG68T/jFRyEdqZWXgOXQzmHgAfx3jqHIUf6
MxsffqaLNrG9lWbCx9dpJgr/HWo5Un/a0LxflXXkQfpRXolU/rLy0qs+NCvk+vPGOpJw1GXh7+rb
X2bpMLIfaMizsnuD6p7TMIVDT1JF6P/RzXDg6Y+ggswFVRDY4gbLQNpDgpxx+RZJwyqX2SysEib1
zE2nlV0YqRmeDV5eNCu+U2DyQHDE0/9V4Fp52vxAbqD7e/8U15BNOIpO5oMDUY4QLvcRbRvdSTqi
orSmwvBgbvcdr4GkfOyc530eqPa2fUwW3vnQXzXl6vOXi7p6AP7j/DeyZdKUH6/mXFMkx8ntzp8C
9jzftGliSm0ZkR7pheAwK4Qvoj1b2/BSURoYP7nnRn0kOnO2pUHtXkSa/MP7ZWrymu9ah+cC7/3X
9LFs1J8/HctIw1f8epz/RTH4e466y53TvqPPt4I7M8ieoqe95UCzwsAc3J3KGCCVCLApJIgBnaUf
yBw8CPPCFFeSCpIkzvmIxpHBiF0X25HDbLDzrZ7U47vo9KonlCDXksyjRQ8jVZIRjpERvPzcIDV8
FmRSEGvs1Yn5cUyDEI6XUYPwUdMBJbxnmQTMi9M4ebbiSEmdSDg4++99JzbEbaHB4HDZ8KzHZbhc
g9Zsgd44KidaeTYMPWK0/U/rXKH61uAk0xFKB6yTShPqWXLH7ibyXOlyVh6lQDzvhv76TR/2p8Ze
GrQEHaqJWJAFGY52jrEsT3j6oaZyj6CSSCMS2yVkRP4lieMonm05YbAw/SB7hNwWlwrcFh3Pg8lN
xd+p72Q2X5wSoh//C20ps6sNpUw2vlq214kvgRoZOO7uTppJDZujjD+IpZ42fVkRCpu8PP6YBftF
M5wepzzCqX55R8tRWlWmJS9AKiWDWa+swSSdPEa3eWekkDioyv8gXOVGRc5Y498X4Hl9TQ+489Me
nwptr7LnoHQY8fcNnU5VGAyIk9neSC0l7usLNge7wA2BzvUXe8NGdwU2dgrb1cPqAuAN0QTDiIch
ZaZW/u6vdGyh2zybazZ17s98piGU1donAL0lRIogvSx7pHL55V7BzjIEZ1SzNWaeHl77teukTSNa
lXVUR/b2sRJCg8vpb998cNJKr2NttzEQqiXXCOM6EwUf8Ue0KzWu4d7TN82ma1O+DNe92mA41exo
G+FtXVtmFo7N1YWOnwMrGLINqKYADWsF/v3HaiUsPYX2u9RZMffu/gV1l0bG9VNgwCHnE1kRV9h3
8IhHIK3NDvGWu5CiYrlnZOPGd+VzBIG9IfeeJx7/73TnkFTVYG+DHsHNDC1sKnGWdAHQgJdYY9kD
VEN+BFqE8jJaIC+sGQqocdPdy43zuDizAPbhxeVqaLsNxS3Hic3P7sdZgW9AIQjtYUr/5cE1cM2z
n1ZpVWkrah1BFaMzNwscSYxHQt7hrGOGTSasXwiswr35fFDhQ9WSUG87XIoubqckcBD2ijJjPdxT
V6SKDvYpvf85voIdHrZ295IfNVe1+0y0Lz7MHP7Du2Cd4rT9ya3zKV1JsQedUOoWO2qXbrdlQ2Tt
GccJQCxM6hJbfQGqgv8r+IZ90yr0pqvCyKMT+cYBlzOQwLBDfMEgGni1mhmI0I1hxvSRFfpVK0F3
buyNjjm2drfkhy9xBpwpvC25TBGKeZ298m+N2rn363XYQ2uAOUaI1R4VY1PVccnqhZ56RzbPrrWB
o9aBxtN6vllMZyptIHbG22phuhie2Ku5jtR5kvBYig4nTEninj7s4ppJ9hwQ37d0oZ8sFKA9z7Ec
TFuSlBZ1pdMg4yhq/F+27Ll9ujJyhLaCaaiDzsE/8pO76N4PyLp640gxNSmcwiau3L5ZhiWNwt2z
CNnLw0XIHk7O7HFlhN1nQn9e6JbmEteipiWBtGQuOy1u9rw/ZXRE+RcojXYxbiYhzFYVzmjXsOdf
4ChL/OkrgdAoctwhDuI7Ow3rU/Eiy6fIlHNYxg0zPqHyL4nmmWAdJ6MBJfsy3792VGnNrBYfxGEz
Q/HfW3oFOzEOwZmPwoRKwE4k7T5X2GUhKnuS2gjNh0L4jtdY1ib9neBPqytjP8cHLIPHaRGQHDKr
55t29peQj3NZMqeESb9uiu0rfB5Doq9lp0i9n4a3DBYzyn8Zsve90ZrxLO0wivOPbQOFXig7Xs3V
0u8umeRgB9voh5GDq75WGuKm0C0p7N6aNmEM8o1FdaG3JIy/MMAz9Nzj95FDWDlKSYI3N/Xyz0bO
PpbgF/IL0HbEexekJ6bd5snjYJ3qqQ1TrpZxnnZ9hrP0B1XmMlIcNNqJFUoWCHSmr4raRWAS3d53
p8eHknZusx+ewGKPCHPas1ajx5OHKNzPzcFmgIkILAVhQiwilN2Au78Hy1sIxqQPhaXcpEkoJV8y
UVo8FvPjCU4OntsMML+2cJfNtbtNV+EM/6cHgix+jy+avM/8+u8Wl8QVAjmt6iCryJhbIFiu5tZM
hIywaS+XBhCt2vV/1hj2uAknvLRPRm4qmr3Yxi70t0dHolGtaclG60RcBan0bXj+GoMp7VJU41v4
2ZPrHAT9CCcVnmFQ0gxPsuE0SANkYfdCqESqLZO6zBTI4sZCTyyfxX7iNdYoIaILKEun5HiRtTKQ
mpINw0urR/lt9nM071qNuGhfpd19UNhvdLAvAgewKIQucTbuWGTUlkw8IaiGC6MtInLipdVpk47j
ByQxe29kGGXaLCkFNfBYp9U870W0kinPLJPd2rM1Ue1T8lr9BdkjvOo7LTVzFTGqXlM4Ag+lKyX7
9mTTh+ttGwJcPeLzMVFoiQnz3tq9p9S41iDvnr/FO6Mg2aKT67/60cR4tZXHDtdquZ2yn3UgmYe/
7rQlncQmEKTBBow2X+gsuAHDLsHcNDDxfwL6vbayf5dr9Fz0wZJZ11BMAs4hJC0+LWKQKBFUoR7i
NKd8gkwWv5PFeyT2pB5CSgm4XgU19Jnv5NgyAHs57EHy6OSb7+nCerMOEBpN+/QPP+RXBzntFPRN
g9n/K5k/O7Wj3USExvrL3kJ1GQwHmTQKZoXQmUHVyEY8ruFt5NVxEogUFe5+EFvMtbuz1HyhcfVk
vaUNbnBrxI3acODX3BZPL/NoK2cNfE3IYG6h8WvlwDEzym1DuDsj8xx3AlEXGs6vHk02Y5QEZveY
wH3zHwxYEG8To+VmHopwEN36f26mJFghekhPlCfYvFYjoYVz+cmaGRsItlwee4rBy326LdSgKI/M
OjT/Po/OlLVkTWWL9As8QBefM2zZighuXSole9JAWEl76QsKchq7ePhWN4bkhpDC0vxouqDm1zbh
CCLhtpieKdilBPP8w3PzGCdx7m2NF4PRKJHQnCqSIoO49TIgYliqSSMGxsljI7yGRHqWExUAS07h
iLGlAhMTjxHwLE/C49zNkcuHc+NmCiAYMteRHxLXGcIRIji4jzNIp7jr8bpZMn7Y7Pi71d2FC9lS
K22f5NoDjJUybJwvIN6k5hNrO2dClkytXwNLevnNFxbKDBYMyhp+w3j+I/gKNw7rvhqIwEvPzyWS
Rs97ptLyFHW83ZzkH9j4HH0yUuJ56cvzGuxddC5MOE+FBgE0ec+SgUSY3ux3FUGcTtlti5vGf+K/
DY6KGIBXpAO9ZK1aiZXJNszRhZQAN13a2IoDG8E5qNa5iFL4Tn5qZF3uTnUu3RjqDPqI2N2/Tq31
TXHe4LAB4KaQDD6MMwwocg58bEP/fhS6Vib7BbTyQLSjm7obBpJqYNIt/QUyVvALx+2aLZ67jft/
9SUoAscCk8cCRVNNY5Pue3OV9VsfVUl3hFNLwgioqanxd7BHnI09z+gG+wgquIs513pVdw3OdOBf
pBo4haNE+II9qqZewdmQ3UD1+tXU1lUpcB03/iG8szGxy+1Bec+RnZILJGfmTLT9ODsuegwfVfeg
LacHC4vzeX/yW6smYXIyMOKBEYiLpowwOBvENN4d2ni5oYB4i8lmRbtoZl9KdYbPPYG9tZQ3J2SR
UPorWALPTPLnkUD/0DCyiLof4qQ/QBUZEyHf4IW+L8xWZra+4AxNcVKzSJUCIZxuSWwy14FE5Gbq
bVgCHE8MR7yOtpkd8b9j6DeVDEp7jwQxQnTze4n81PVjlEPjXcZXOcWk7RDPE7HvKqrjLECwney0
ThYpvRiA7vlHHkM1SkjkTNvNfntEvwazg3OGqVAgJ+e37lMwFyLtHBdD+ibRIZzrYGgNnT6Zt6hM
rJnvTc8lV1mtR+XzzgnEm6dxQGr7nyYPLR5mCcqWLXXvXpF4EFHUZJ20fL17DaGY8FDAz0ptYVEC
AkylL4i72C3COYq5wtfHLPWsTYydw8vnt9iFkr7cAPaCSeNK4PjpVyE3pfGvMW8tQl4s/y//lwzP
frOEc6w2zUvIwUjeyELgOlpQINRjWZFFuKzY/QkGdODKvFJxROl9qUYYYB/9vXOKv+id56BffP6c
tCM35uWDVhYGcVJf+tI6m6dO4rMVNZrxNnBfs+Ri6+eCIO6/4oOtcXa+tkv5XIZxA3G1mqBKJOGj
kSdgMw1NfYe0hvbRLL17Y/3mEbB3PrtKbf90wB+2USnII5cpty+FHwaHDRyj0unuo70HgW8KT1qi
uDRPR7VwUIK6E9V6QnG5n6vKQSX+y/nQxZ2Y6jftBNfDkt+GNUVy1FnuqyyTyUxczJ9xzi9ft9rj
yUXlC7ZSEKTpIEwg5bjLnDNxTYwNut6KtJOlhQQsbn8VJQQTyFXKB3Xeh6HJNunSYbYcNUyupOoL
Cr7Hz7me4uqw4xSU5z/Zeq6Ac2G9BMggiQPpc6sYeOItD7jSaKaoxPDJqluPC04Wje5vyozDdaMU
uajfIdh+7AVrM9uy3A7WQjM5AXR70l9mtJDVfi56KCc2kvzdb1/JaSD7lwyjvyMp3kYvDJ5oRDoS
vMJoQYIbRQNpI4PCZ7MXzfu0FZWCgE2tBhzmDF2kCu9XoqRPb9aYTg4dcNVOKn7Gt5mFqw7PPLA1
fisPUrk9OFx/RPbBmeR3J0iOj/aFoIhHnLhMWpy+/7rdlb8Ty5ZmhocWTqD219BbFm7LVVIGwLOv
4FMCTviTOZ6Q93Wp/esqefsenEEEEdPkX3tD29XHZbn6Qk5Q9N2G8hJ+DMM1Rh2oya/bHNCx6utk
XwFF8nJnp7XotAOPa8vGO+QYjEJsJ1vnnk3dOHfrnO74Dg0NBKRa+4RNbcRN7wMJM+Wsd168JGMQ
O+Zz1+ZGvH0JlDC8wQek2ya0QdB6MhA3FY4/RtLYy5gBVxhMLoCgq0qIeLmbzLQ6xXI3K1wvSeAv
jE/Js2xVyfKMVGuG14QrVSoJfDhhaM73s4UAFu9v+vRYICxP6Yvry2Etv/8Di9dZSU0DWp5wdAst
q+e7nVuqMbclu+afy1tKzCUoU00GAOu8QAVvJE6tmc9Fw4c1rsxGq1QpTorHqgBQKoNWibGX1DLd
5bfVj6Zaa9DfuvEJReSgY/zqrelIBlcElv92jMIvbM/L4nUmsdYGqxv3/xmv3M8pP/vURnKmgLtn
pVutcKuCxXLpNl+y/hnZKLMeRLc2GLGX8UlhzlrXeT9ZsC+EZy7OXF3M4iDD8/k4/QMQYSETQWdu
UWcDBUTbPdiEBYWX2fYjr683MwHjkoLPBQEjFtczmQhMGQR2nxc07Vk5Xm3JG7nRAGlehgyYqvy5
+BcFUf/YpKEjbrRHvc9at1cLKvZSBPhkHsI1NrSvdwDYLL9k2dl0j5T6FoeX/vupaH+9mkZ8TjiW
dNa0L4n8mqsdr94/28h2RCXVpcSyz6OEiqhdUY/e5hn5Vv7eBt4dy738QMTpqW9WzZq3sfiICgzN
Vrk6koUlD2VgHdl8MCfDkIx64t+Dp/DCOLxAPA6QHZTDwhcgyUYIRxXbGTJ/I6J4oxn7C5T5b/QZ
xv9i84IcLBxJzBxHKz+FSVggNac5FdwxwQYONl7a/St/e2NNRVvr75NG4mhCUPpQo1RvVfrnfjsz
aAQO6Zqgnu+8gGssOFf0Wsyc6h8g0BelBdx+xHklSglJg1IKAj9Y8xnD4B0jaDQr9yDTt6e1awNv
USGKBMc5japlhSYNK7ZjtuOjhIK2U4R3GRgU/+LnU4UJcG8F9q7pzo8U77yxEfcKZviYO2Zq+3KA
xUQMRaJiur/IKhPx/NVO4vAc3i0Ppm9vQE3P8wT0nlS4xmuRmGOF1NKIar6yzmFA4wzyizqvnpfj
gepFtrvvYMEEwjErad5Fl3ksIHqNBN99I9RlcT9+8QkuYlThch1AQz+eSwH235u+na2NjF4PlUjX
qMH/wa/jfgQjb6gdV8gl/tEh8ULsj4vd85hQN6pljPyof1Rt/QjnMsJTeaFRDK0wqoxfrwbGG2uJ
Ld2iSw3sfqLjxXJs9aROAATssds1zsG6Ws9ggc8P6rHIQUAbrL1RbVJmZuINHGTlpo+xK2rlu88d
BoJ6ot2pI9SpTKlwHbeX83BQwl1J1ZDir1FpJHZZ7YDAUJMudlvopJ2QuP9sQNtu+WexOPZdPbKC
JnPfqsSfsnYfnH//nqkdcz/0+7B3b89E3QvnsSVxs6wEmgvJTj7padJDljmu1Ln5CuQNqrdKdic9
mWHNaJaYG7C/jOQVyfl0ZrpdTY1XAk5A59g8FAV5AcgOK65LSAhg3RitszUS9CyejSUxuNPIBzwR
t6v3mEWT4jlGT3UGjwuwMjO0kFls5vHLuK817Ywj4hdU2WN8LRg3+XcwwUVNxDgN4UFF5Qk7wdJu
FK4xdeQvIhWSs+4HuKeoj6+KwVU7p8+l2m7SuitDhnyHUcEbOgz7BcvkEncvh0bxIX4JdIQVJDM/
hA+I4AuE3kcPAednJvMFjCfkoKwuKh/+Y2nTw9k+fVTpbGG2bX3UToiANPxm/mzV4cACgYaGgEEZ
neIeJULs6KenLCEv3liaQFCWNwWnARRGIrojOmGl5I2QxPnqKV7qUFnPq79f1G7Ba6jkXQDESiU/
ZUaToQ5FKew97emFhRXaTHXCZm5L6U9MTkZ9GsE9yS9mBLbEI04rK1kB057c33RltUbdDXcWZUXo
5HlhNtGsRATlhyDZgG0yrfwI4oqa/oldYFGA30X4+ExbNFXCfsn3lXNgFWjE4aHrNa9x+9IqonWS
K+V1DY61bDVEzQ+T1FUXKcV90GVnIIqGyV6isTKNNrYX0rXNYC+mlNseNTHpdE0Wsvq7nB8zo9Fa
NkACizvAPNvxxXaE6ttkkhnGqBsceXpgv4gGRELs+0OenaGn8o9VH7/zBSQWgc31EDzSRajrjL10
cYSHXSR5u+hXtsiSNTZpf+yUnqGEV41SgpBGUv3HUHI0MSkQtbceQfx52qFjTObIM9VBfnfpFA4X
p0c3H0WKn2OFGioRnE2eDZAZGM0yiW7NlQ2RtWga3Lb0IekLIv/VJxGRn22Bx87GB28kkXQsdI9H
R1pVo8n12Uu87XkVmviBKVGgrDy5MlWvfNUTXWD+rVJ3DJYMvyoMSVGp0jzWGh3iiJN/3VX+YVwN
lHD98qs6kRgejyVAA0YY9mnbp04b+83duRjGaMiXTjBfe33LcnycC5QxGyUz6j9d47YKLwB3neGj
boZctulVuXq1pqy/ZcM9V3XEPn+qvhfWmkcZDKihN4LEUfUg8GowGuPkop+x50DhRWqIL7tDB7FZ
ATAibK+2M1XX2gTtXitILr2njY3ColmW0DSliWJAVtKjg36uhRqlbhfQ7u7X1N9duYl1959j7hUZ
2dAbhZvf780n11r6P8mwqTJW74CtAbjV8SqZ3z3unB1os0XqjIzQvneXu7ML5YWeciIRhnYhQf6Z
X0ncyBrtyOjjzwkuus0JA5ohufrx/sMcGCw8z1bhxpawmFeexUCg0N9Hdu3hilQtcQkC/kS5PKXj
LTXXNu5TCcqbzpVrkqqXicKfGPM3hUUI4ZSiDiDJmIy1kpb/2KQfm+K22CdjVQEyg5RRWL2M3LXH
mkWr7sElIwkHybaeOuwq9fE5Id8HeYxHMo6Px6fWIz/LJaMEm3aFfJZ62/3KKnIe/Z1XQBf2YZJ2
ARt7Zdy4lSB3mWO+8Tb+LQ5EfKB2BmdfLderPLYKuZ9bigpk96dwjgjQkmDV75gBWRg9m8vdnv7L
ggIin9ekkxb+4Ugi8Bl1B/+WwYJvdNW6YtAgYu2DdH6ZK58NNPpwrkkGM35No4ARAWj06L+gxktU
lzNo1QpltrSGWRfrpRUQIYRP3cUr9rrSLkIupH7eqrlXhsayzo07+877YDuhvBhPNqyCg5r55nMI
JspA9naUKNFXCj9uOxlR900UcRloXag0TjUB28z17tupl38xn+qUs7nSlepvI5ygVFTsx1TyjelZ
N9XBqZvfv65PE9oH4mUlA4Qx0qIbsLKCc7RjC01eA6tNtPlCcWkMW/DswisQBmi2ZzUw/LtWL+sV
rN9MG7gM30xjiTp7xyw6+PKhaLjSzy4d2IONTS/HywvF2WmXR6NDbcA/Cy4nR3Sqy3yw14KHfKvQ
eUlNwioudQ5rGkZHjSGWotHusFyqHGmls9u4fmDqBrJMAhKFuLZZwgugdPZi8nOFnQIrghjFZAd1
+2c8dVmO0rsRqD+GCWPe0Z9WPkZDc4w8QFMr2/kLTcJvZQJiQpLgCfOgU5SVY+jXNxtdfvZZDsdI
C7zutxowmzIAFdOJ3GvKrSLaemcx9YQPVoIjX6MUUgbOmS+2IR94FspAIsIYyG/XbMrrODhBAaNa
3Oj6lgeqphYcZlk/p7WQpSB8TjigbAL5eWlRixgSkWtEGPH5NVcuKrFCYkILrfFA1bjsbm6g0dvK
cWMqg0U7H3h0EJnMkvf5lDrrcxnk+t6jQD0trOIjLKppN2JNKSmWHXl9/x+6lXBUJcZW/Pce1wQJ
DjLn6HyoTmpPgud82Ku+7x6SlVKOhxBntFWVYWUd/GqGjU/GzREa66wHUETGLts0MnxswOL6qjEx
+E/a1wfzwM2EGAPb+WlFAK3yINvgaXQhMMCkMCeT5UBUrlaHLKI6GSksQQltkJmZLeK9rCaqHpTl
u9iWqtXQp1lmVs0EdfHoCg7DIG25wJMjbx7esqTTc1xOyxfXtKWHUJRiDmO39Wl9dk1u3cdrSXim
kluwW4GaGKtJzAuSTM+JmIHPYUSJRvNmRr9U6DQ7XUMublpgB21Sv/1pWHAwqe4eEuJ5s1C/DJ9K
+qHAxBuhbNJAX9jhtMC/RjFetjOlQX2D9QWcGZOVBeUHwLxvvOotM20q+lfAt8BQzaOxYyk1OOKL
a2NMzR/Ukvp+xQNDgY/bDFDATDrMiwpmiczUxqnFf6HNMQXxGaV8smpxOoYJBeJmeVRuIS0u3smK
h1i/ZYinls7vilD46ZrBXmi3mUdzO3ugZgbFLiYEWJSZLZ2YpuZOqY+EL11O7uYiA9yGIDEm8eEp
6MoX3M7U909KhluEbE54qUxJfiM8/2Mo4qJlBt4XxqoPp9bWUhHLe1DyG1Vy3kZ8d/mTCbq8uaQU
6O8U8AC0sHpD6tQZK+d1s006D2YoJR8GyWspBvTQH924Ei6n9islHHAbcwmf2S3pd+AHvCuz6iwb
XI83tfMzUoJYLep8b4uyjpnkE4rgA3r/1QzvRaLbr9D6iV7b4oJ7KpxO2AYw95mV2KIu415seGCQ
88gziNLwMGFG+9v8MnjRKrXyGOB3LarOElG5ueZhWks9lZ3mDbHBdbH3EqWDp+VQrAjkKrPrERNt
GYRI0k3hcgrDKfWYj4zcN/krZSfPv4jNhNrggbQuDqWRpuWiXu4xIjQ0CGjtjIjbcFG3OjBws603
MypGozVOvJtunmaMOgs0M7553rfnZr6hYD+EhcocTRE/GUOoOW9P5oC2MHqg71UF5+yK2R0Rnntb
W6/KlJzwsABSuMCkK/nph2gl0zZ5FNJEBpkxj8mNwdkA6/vbzJY2QleOlENc4ecyZDosrIGZZ0T4
kO8ADFvuTHjU7IDuSsn7RRhsSA6bxbZtSQ+5huSkssAYN6ceQ451MNAkjzkQ6qo4I6sf7cL1N1Ii
QwzsmidoiZp5uIA8wbFddDsOa0mP0KoYboaVCihMP+s01b/WWNlKHjqk5NU0z3UJtUEKo+tiF4Es
SG8cmLd8plsrp9z+Cla0X7UJ8qBCM8qswLw0PaPNrNGjN7U7L2xHDNbji//ulEy/f5NQ3xTe4KUK
0RCLMh03X1/2C2JQP9w0V3ix+CDKqGRNnTgdoeGqcXqqdL0ChLzLlP+f8L+Ok4iacGSr2KvqLjxU
eH+TK4foa0duTjdpeCUATFLEzYBZkWgtUu+lx6rVos9IB7oUTvwGgPcJrYZ2cUg8evxs89OE0DL/
BY6SNYcqL1k47d1Se4oh2nZFKjo1PfCZtibYh1PlaFqCngHhU9Wonxy1chnD+BrxgQH2+WjGH2aF
YoGeksUyjMgEQvyrenPeRH2nK7Y5yKNxvPpHP3SIGoyO+KE+WVUo9hACR/Hq29B61WbLfrBmgaIJ
WY8/4aPXlBpdNclQ2cjLEGuvCPIwfiXgg/5LdDDFZgzdio+9wY1UtV4lNCBwddqSxxZnYhGxxKGN
VRy8xxeoVz5KiTt3/J1CnMsGvgmmzTntbrtAxxdro1IZystJjXDdxLzWNwhH/dnUvIbB5FxKIasy
4pHDZsKxeO6bG2jdfB2Fc/uMWbuD3MKRyEGDXEbgOij0bOtOQTtXXcs7kVUG4fSpv3K6RKrN/Uyr
JnHuSA9gRn3ZRrI3aVt+iUAkaEaIQdVb48bcyvNGTHgDzk4jioil+Dhlt1KD8AZlBAUFWMk0XYmz
dO/TgXNr5lKai2NqUOnNhfzEpyAWU7JgzV9CDH3Pd8sKJIcUVKP7tl+eyE/drn4tg13KdSXgAvvd
W27rsUgLmBGS+mNxcSVpUwiw+HxDP9lxdp9N2ZnJujufiuww21xsvbGExHe6IuMUEu3xJcdyBzSD
G7CLfg6Re//oD71kvzqR4E8hA20ybfQNjbZfo693tLlqyrd8jORv1XIjp3cjJCFkuM84WoMb/T1L
KJCDoVOOXXmRYXpiuC7UI2du+AP8FC9mYFYFfNmhvY49OqCJ3LQZau5Qmt/TnwiqgiGPV1ibcxBv
a02FMsEOQQE9ifumXTFtSopclUvCUM6WbK96EiqPzte+w3Fhzv5AGo77KTsYcNLwNk2KN7SnxmMA
H+9PYu2Jpct0IN/IFHhLwfw5ylDv9Bv0xnFGrYiEGJeX/zdnaQF7pJetvItxThd6cnoG8ptpSoUc
x4CdYDbCq9/+qxtvqzOsqHOKNZTjKJc7K11v+jYHYv7gf+SI/qmXx4BJT8m8QwBxCKZSKxiBOB5H
Jdi9mU56xJDYDbzxg8f9BT9qB5Kxtuw1+W8eVKt7IBnOHMLlcrMOaJbPyxPI8QhEw0Segti0/nT/
4kfsTW/hE6+jSzT1Do3eN6RlmOFXuS1YOP9IBgEWNhm/B8mYaMHTPdEk9O9Mr1ArC4tuy1PMbRxR
Q9GBouqZcu4g3tNoWta+tw3p/zx8RvReHqBlQqwLQSH32A09QuwL7x2hD/Oa0RG5I7SnYasd38Rq
raYiXs1iQq72vlFaogXGCN7iNv/A5LCHHCtSVI7ox0V2RBJKpfXaHzsYITe7xYv5kuBVLW2BWEFg
v1S2bbBPoop/g1IRy6k+hozqRFyvHBt8nvmETpaYFbZ5Cx+XWpub+QXLcOFyDoibIFRN0CFcs4jZ
g/2NMGBDpkxfORTl7F4furdPpIhuE/75yC8MSQ8f0OIIP7X3WV3OzWXdZd+xYjQ1pwI0SusWhS2C
IDL6wvIJddrSNKs0lxMERwFo2KjrBobFr4MnAWOSJA0iShHOObQKWlGINHL/050d/33GEZSAX4y+
AUJDjNv6SPBJiSFfXBJDU7L4v998ZETv3ycFM3DDkR3Kns5ojvpBqApHnEV9KrPyQIYlnIcuSMsR
S2o4R76Wic7F2rA1Lfa2SR8dEILpdXrj+jXgU8pxtLbgv9VEfdgFJz7tvEGGXicvgD+gr5YlR3H5
RJIgbtWwqP7wwmQxCwf3NslgST/wIlfxN0siugWhGukAwOylTv0l+ZR27pTOmzTnmC3/FWiNKUN1
dqEQplIbRjtkHGgRw/DmUhoM7W4VFXSZ0EopWhndGiaCSd1d54Cix02cdWwxNhoLLp4ru3qkzYlL
hICrrEfWs02Oy/5uL6uKQIzWK9p+smV+UfMmozh1aGAq4zLJx5vKIq6twyNS9PyXp5VvrzwZ+Zpo
GVoha71SYwBJbSU77JZp9Ym+Wywy3zuBQyF7AP9fsiY54B8Y+SR45Xra3aIxJzUL0zCl1p+4PA2i
RDZM4/3fDePPegkW9ppGjCKgHdINYeSvbHqDKdda15y/UE+S8Kj87eT8PrxoqR5Vda4ZIrKQPekU
X8lKiMsn+dOc55TEzPgUFjfmEZMbS7pyIHDV/MKZFKsbPBU0+cbYUUYPW8tY5xRc6gD5PL+/I2z7
X19ESK/HLw30lpjY3u4AgxgnDfEc0napnnSyLXbAtcC39dQC5GKn30t1FmhyqwXKHAOO+pfMVNCC
Ple5lUHdGv767ryU0I17eKYG/111c0qUq86HnCPZK9hkMTn0F2NOjl3lWCK4UqknZnKj75U1RuFC
tvxwZzSI3/xZV0rTou3nb9ewkxDqGMEcJ7QlokxxYlwZKpS3kTKxfRo07sHXHWaWbifayqxk00/n
29DihKfekPYrUPY336A34Nn2bgNP4fIQyt3OIxkwyb6uA5nWViwS9xpcZZAnT4044Sj+UsnSgWzY
CRLRW4XJ6nkSONNDh479sd+fZ2wg5cwW/dXGg7sRO4z501rZJLrc5gg7pPslQyLMxcnnkz5LlTkT
xbedrDlP2ngiOWEwv8JiBBKW7DpKLRKmnU3Ubh0BGhGgv48K7PITT6cE20p8DL8JJGM4a/uM94Sj
+LeUhn04Gw15tENEMUOXTO3NrzTddioBoiYXuTxFqNcURierfLx0MC0bJf4/DIgHuyZGEAe24q6T
CuzT5ixXajnr5Axo7KxG9j7fGAqA2pKHZug7+zKAFEH4hThaLe2k62uj8lgo+Jjcae30Te1j8gzz
HIx9KSj2mK/JNQosrUoRqKtlR0Mbu15dGWVDcg08z74ZtvZze5rgG06IZB8qGbgy7+4ZPtbjMnCZ
Gawh6KRPVwu71UVhH753Icf6LJCsZFQz50EalSWC1cBr+XkbRItXNx9j59j2uovJs+aIYnlWDj9x
3nab9dg3NjVLogLVYmagt7IjXUWzV3IEZ5m92Ydb2XECxRlm4rf/Eb2aY2omHRn8B6w356TqBIBe
nUTAyNJGZ0p+oF5y4ju6CMxHip2Kwtl/a49caWZicsw330y0SN/WClbdlBd2+cCT8cNygS0e/Wqr
UwgF4zZW7GIbDtYrRIYaIbckHQOq6xr+KXix8Ct7OiscBMQAIneJNiF6ROb1j3UHfdK/3KbnCx2Y
2V/TR3NQBUiWT6Q3pPDCxN/shOuI2cRtpGaMhS33ms00X0Fstfd3RPbvVCxHCPwhzopovqEHNmRW
mbBhN0mlng+4SlFnr6nJxPFx9PU+UClokur9DzN1Yu5ULfyDbE0bQQRHEw2vebFKFOhvuTEVgKsq
KM/W840GnTfWuyDTv+mYtRgwxsDItem9A9ENdk3sHpom9nhsnMlVywQTIPWMjwfgTSWeKbA7JaRf
1vvgZXgb6D4ezeR+f1TsMX0/hi2k0dd/2QGjg56BWIGXZ9h2ERI2v1ceugC/KIJn3QfABjhw3wla
lzV9Yov79vGhGVlHviavfUYUwbKH32TnH7dvBa0GaNQxf4FbidG8LwR4MGq/XkV/yb2Qu7/Kbw70
AhFFCyuaFbdRpHAd1KumFeTl3UrZaQwtBKYsffzOMreQOGULEADDgu6MEVvZofLq2oCbY4slKwMl
4UlfpIzEmHjxOIY5nFweQmRTclV/dzST9yu/p/ZgeTQvPwi2lW8SDoXKlTIpsCtGixjQukoNvZdB
IgI8qyeKbUNw2B3OzExocBdCBnscHebUySZ7WmDqqqgqgHnLTn8fCSh/P3raih5Ix7bua+7/hZau
BtXsl1FNUTECK6sLN5wfuEFWI+jv47CwtVBqb50V6yrUKduxaxr79TTmIyofuG9Zhs2pZS7kYPfZ
tkisscZsdZJ2lDvY3ZNYioDngAecwM0Z8t7cWPnZaYISLLvvr670VIJlWlvBwMTro7s3SgYbxWcn
+8o4BUL+CnJcckXKB0Z+bR9Ha1S6cIApS04Tay5VosuKVouIh85GBcLbXO80/HfEzLPGghzkZGzD
v6+vLRdvimEwXnUzVO58Bz+DLZ8jXOb5FB2cvlQPsEjNgu6nUKfeL8nZfDp9SkXudM6cs01DfP2i
SJ2+3/GcnGVp54Z4C6ZgMVS33t9mxC7wEQPOjdFCardfAJQ1ZnApFgqPzX5v+yRNWEY+T2p3fAHV
TL28je0RWS243+k7jl5TdqbuUcOXxsaP0J/lfkoK/6M3tLRhNZ6E4VwrG4eNcPCEr1wIrJZ21SfI
qExKl3NQKHbrbG2FzbvK3Mq/kepgrDG3Kc/tTmPn7oToRDFtj5pwD3nC0MgatWDp8RRPqWygop7W
3FV218UTM5ftAEMUNtm/iH1704VwbRWkqmoe8Ukpj2AU7U4cd0gAuEf15OCYDArxYghx+IuF7E1f
Rmkos1xQPDQ9IyBRqGJrhQgZi7j5vwgAd/ESo9QTgmKrlOvu/YBsBzilt7DuSz2bBZ3ygIUB4nja
fTzIUsk3V8IzC7mwoB9h158dO/69VQ8TiAq6KclaPyUKvuZIJs5A6voXsY90u6r9CkBeJDDR5A7d
sbLeK1n5p3jrG+mCzDUS7LA+u7aoA96Xxki12Aqtf6DNgOstRbC6bmqxxhZ7xUlgmNQe9ghWpXIZ
FfSYpKzQlBFE9fMhINdmmlf+dwDSc8idolP0S08aYngJ5d1yYyfhfdiYCG2OXAvGnTApLKjOTphV
QGfgJDSJueqd6H0EbFfH8sRHKtgAo5vHlOs4VPHXfNPWe0aqR84fVF6y/4pp2Qru6dICABNCYTMp
D05jpuyRfqBB+WY3xosZDtLWRWauENhIGBqWJXEO4ZYZYkPhm9Lo2Fijl8Plr45RKOrz+cVKAZwo
voFtQBZNX/JGDoF/FAGN78OZshBVp/iECHNInHrUGMcVqjkfxsgXWQw3/+4fsbwEiE/pqKtkXpwt
i3nppePFOr1jgiWmEgwTvQuynZT1fDgZg6kjlevKL+VlVpR4mRqRlWB/BszwaMmQS8XB1o2kuPZx
C2BQOOPxsRAdmxX3eFJ4nfmcx9pxH9hiNRcIEv4YqTTi9ZMBnAvASWiNKKOnyUiOfK8lpByDlS0h
42y3eeQ6lJlb3QqEdv+lkTqkmgfZyQ9sgY/CHANel/S8CU0TaqRsyazRxWF0rpVvUcGCFq0H+Ssr
bNEbeEkGPT1tY/tHnsjWwebxWoeiGxm5XBhqNWJQ5N07FWViQIBOo6CGp9WEl4vukex/YU3yZXsw
5iqeI/CTsgFn4LAf+bi8GnTpr7m3HFpoSO3fTAnHw9i3aT/GllEI2JFjQkAOCqpBTmBVxKndS0Qw
gaEN45i6di8XSEzeHj1tW/4FeRdlmZZ4QpAoHh/9l/pVdFUlqe4knzUs7InzSG0792lz4CLj1/hP
oE348DMbjpgu1F5zZ/HIwW1NXP6OM7mpnyR8EBMscORw74GRxkjicrZ69tQGMfKy8N2MtkHihDb4
mB7czkKfD0lsvybA7IMjqo58oyZ7D66iuZ7xCDCbouIO0ukP2c5NVSMjciP4BteN6BsH8ZQO/zDY
OBKE0J5SchDDyM9mUZhsl7M1mdrN6F+6kH0mcDm6FOpo8AVSuh1/N61FuVCvO8vO3wcLqxejI+Y+
JBC9g+EjY4R3bZymv7v/VtR+pifwLXUTMGS5CP89jc0opjZ3KUVW4A2+hkCCtD4bJB0Ae1RgcoCe
CUOoTfi8G+F9l++q/9hJfak6hbC0Fe8d3h9t0GgPkE4yhAVWbs93E2yeb8q6JvnpYq3JTj20jRvN
HSODrus+V7llIZbIvqlP+0FhypZULdOxlfa/tqrXu56NntD6/r78d33vHFs1Sp4R8dayaGYkPEFT
IRKOm4oZHHEopCso5SevGqbPdF0wOyK+rLha/Zxdi/+gDzdU46yGelnuKrvPMz3Z6xJsdou6QfGg
dtwhpnzVWr5YJdW/2TPRkWCGcA+uDVOilxfNCzW1myePVbMivF7AnaMW1hv0Y+T3GHTCtl+fD5+o
8NCJ0o0xpUQjfUDeqnVDShLeCOFgBnjpCXbIr6obQ7d5f5TNgbKHJy7pPDDgQC74xE30lB3nxrq7
v3UygYI8LodSQ+UX7n00IEcCykNyDh4ufvNGUGbruuP4kNt+HDTNN/bmFi55iyExe1nLweSwV+/7
G63YIp+bdy0eSymxQRW3y3mfIuPApwB0ia+B/4Va9t6hAfANe0S8swU+ZBdHCwaApREvf5IYZr94
JwLrq1ZWxGrGwYAIJl1iBaVEo5dudHetauYCdhP3MQPU8wgDc/dqs2nud5x1BsbCBwXPZvdYOFHp
hZyBUBw2PdmizsL8v4lv/Mljx705i1j2fXwoVsyKka0TCTk1ln6LhKGS8rkfl3OzhOrJMX+O1lLu
Os5Kf9DAQRC9bYsolBsVFmv2HUYD6r13z2rBDHJa2JGU/kUFCEbvhjb1ooAhQRoyVnPEyIiqaniP
EAWH+2WXOJ6ISKHdwsQzVr+yuV0VTPPVNKh4DktH7HVwoGfBrsbVbqCtZanHER7Y2xxTR9wRkyG5
E6RugI1RiNwI1V9fhJT7RHT9IWqS9hYLIjzYNOe+Vt2lBIQ4r/xRkvzhnWoCDDpThk1EHgK7V608
fx5jhKpjzEEMEgEKJu3zwKbUfMeW9HP7muwJgQuDPpxonenQkFnNDruy8cubJwNCDA1Bg84lWRkp
61yRdUb2gb1AKSMGA/+eBLTm/aijTk4urZGeQ3s0VaRH0TyYfwB/uB+bHZG+nY/Hsal1trpC6O3p
qCbrdN5Aq46kGmswbVy0l2+CLd9Ws1BHX7KrQmJICDgQRBilnY+grEGdLqSnFRVn0aWKWK4H8Swg
oahUxkcQfFqOOOEZ5FB8OqE4Gv221Snl8hR0UiuIZ0BnXabKWm+t6KUf9cP2AzTsIYmEa65D2aTl
lVHBZUxWbW75RAhvCuIX5+WnOOi+eH5EAjaQm6oFUfuTTVR4bMt1XxQ7/+bqsO1GzN5mPvbTzCHv
fSVegN/+A4Xvb3RUmp8MF9KGDNmJEm5m5XkqdQ9TeXX+bRcnMtCx6zwIw5DRfpk7zSfDQ1KlIH2b
o/pG/jgROgGu1nXPF5y/HxxAQIONqCpWc5axmts9boJ08VX8tAQeNs1r6KvLqQZUxDbk6LjpZjqp
FIfD9hiWOpZH/TBARpeWzhGzBwLqYRnv1XmGIpQ7A1bvjz0wcl8WWInpX6BAgez/l+qNbKHjlPTG
lZYTFuBDb/DuCZg7mRijoTDxY6T1S7TZxZBJbyZMsSKoVlEy83v/hi3pZxhG+ljpa2jzdPf9Jf+Z
9KVuTwv6eBbFOfupqRYV3pIpWEYf/n4AboGEL8LpFgFrZCzoY4/LmgoUcQi9mEHVE7tXgskPKMv8
072OCGoaD/9LLDHincgbmfqvYDoyKnGMcsDQZd+Oe6jgblF6UQdPa/crTBuOV9dsBj7EhZH5nRs0
4BFl4YIk16zQGA/bevMCRV85PIoLDAhrRmzGWsd71JZPruSY9E5Y64LdJ829mp86XIdCM0kCUbIp
1zmt6WLZIyNLQQ1fOYWOltqZyt0CEFXq77blzFZr78FnAoFQWODCL1eSFQjxywx1zNed6luXiqhB
UymM0Smb15jIEJrC+wXycp8eksNVToGXS5ymoyL1ivtGNpJZ9vjQS7yJz1VDiI1jgOXSKCLLJlyI
RzEAOrWPX9wGIk8ODM7KpB8tfLhG8BX72/NmJLF1rKdnZgTWMTjXtX4HBSK/vMvD5kGXx3PM2WFu
C1dDqLy2xm6aQ5RXepGVXSUnjdOIho9zHsxH7lq/rpEAIAzaLYSK0XXUqbLT04+YPm8QrTsb0wv/
HulxM8lUZ758uBmpg6kJPe+StNoPOrcP3yxlMcAlHzFpAIJhV42CMongaXtj1wWtoSDyxHIWRyeX
6p5P5qxHIL43MGpOZWI5xdVKeRQftMdGoAl7fPfGDakkbMYbj8QktX9mRI5+/PPxKrYOcQViU6YJ
2gsDOtJZmFza44wvZSS6XFxLzJrAg7v/UrWHFVz7OOm3zJevHAmBIwfQeAX97YtlXl80MRni5Aci
O6NElFH5uLuD9V/tBe3cw/mdNDdqJrfqCUqbDFkKtwdn1w9kEd6scT4OM9NFzB2slMZdYuWkrxPT
nmM8M9Y5+ulzdnOp1JXIwAUuDGueGqNtH2n6QohYmJc1dr5S+MnDUtTr6vYgyrFJod1LwtsCyewl
u67sySB7GInFcNdl0PbGniMRKYRe9AA85bbX1KigrRxqPpor6kLwmDVkEaLBa9bczqjRgDl157Fb
OdS2C+XBC+VfgYgDXVpI5d+m31RgAf1NggiDmpyYxC/xRqvydtQXTVzw+J5WYAzBl65BTSuJ8Ocn
qTpkdXAP9QmEE6/1Wykc5Ccn4rkeVPp0xoKsNi9YFvB44gWYv7jY1QxAcM8r/6L+hNBZhz9T1U29
/wSL4XErQ+mDdOcKWcXV5t722omkEA62qURekd654Lu5q92Of0duxtPjQXq9FT3d5x0VX9se25Cz
LCb3m01TwRjJlhfuM6E+mhDgMubM5DD7+YMarW+AC11S1Yc6xjxIoMKDAO1CWi7YhPX+pL6lfFss
H6ktg62BgxYuS5A90yEYvKolSQWtwIGAYXeMB+MeMgP8Kf50oQJHLaOYULEWDttkDhSClpk3aIZv
s2q3bdhT/C6nAeeQttpN+13IWPBsQwC9ydY6WNxFKMomfH42hhOvS8zT49ElINJsyvk4Jl/FBF60
8wnokprWlLe/Ihi1V5VVZE4WAWFRf0JN6XYlASuKzG0toAbF9f4OEz6N4oHWqn/NxCdBwUJ7WpQN
lyLkxaew4QyIkBzilqlFBn7QZZPc4PJEmGb9lu+PeD8i+NV295iMLRj5nU+GtuWzK+2zqqLbM+Yi
6bk5YoPmz24ZWEj36eRja3UkJgXKJzWwLj0srZkEMEWy0K83QnBIf5xk+w4FaG131PJvwDNjHwDr
yldadN/zz7yiAdTjbKZS7haCZ3JsMiydge6UNlQhsZenKlzR+Co83qHWCJq9vo5bXgS9KM8SCRtW
NbGdhy+ovimL8SPKNOqjS62/VIGGQmfigV0m1IYYI1L+1k7IaP/ptgxlHwtdSSckKwOTXyQGHnD7
m4lkFVvkN623uQzZWGLtY1amwy0MNTLKS3tPLoMTWfwa4rbE0hZH1n4LaKo6FKHgzYkBv0ArZD6e
VyM6McVuJ5jopcsVamZ90gC8NOXywYX66+QqffpePMIHJrqPY+SBaxO3h2i52l6impviDcJe8kjF
kl/YfsYvI63O51mUjC4dgw5ARUJ7LtyBIezeaws52h9/Zww7cGXwtPKqVuR5u2xY2gLPta2KpLhd
fD5DmUsQdgHRCNd+jo0Kle4dw3I8ml8Ybz9yZM71jdRNFaYUoegNLMkj1gHjjiM79+sTN8OAg5LX
73M8oEJrLIu4UfyLgUMl2XfZUYHhcW7OL4WNp8f8KubWls4dlEX17f0Wx6+drz2xIDtSc6N0CVz5
alJnJmN7FREacWoe37CtsWEWiODehHZ060SMyjjv02Gf2CTah0E1Xj+1LlEyW4OmecbT6LtrBTza
+CCkEb5HVpZs1gj3A9a5J8pVPvZQmlYxSrrwG151iRQ/Srh9hCptPAxVIaUz8GAzXDZOGELz54UP
xt3uTksaD1aD3EJIh8lsEaS2CejuB7qOHfBnCr09ut5qbuQMJwv/zD63kr/ORQWcTm+lOFgWxjMG
672pcnFEgwTSDnqQXO6JX5vS1VWSMPAIYlZBPsi2N3Ayd6HmUXYGUHgri0b6ek4z9tgvEhwrIyJl
+HvYEFcvdal6N2/Ct4meBO6HnhkJ/sZp0VgQfEC0kljZc4J16o5wIRu5wZZv1JwYl34xBA/QBQQC
qpuG5CnAuFW+Jj+NjD+lNkwzg5+e/sOM/PMiWRopn9Kloxy8vCPDmwXeoEBxu6QrK+2ZnDcFKRgR
MzCLfd2nDr6KEmy+5TpnZXN4OKlX7vH5TFDdI7VtWd/GhaRlqZ5aTHD/tOy/l1LFTnMoPKFl+cup
Tds4wp7Ru9DwIuLCv+/LLlQVMWUUE4KfGBsTs+2jpFx4TaTOZXsfJJQspgat8SX2HCx28nxNkwMT
5wbWsGRFQoPw1Q69ZL5v9ChLob96CSSSpD6YnIe0tsWvzFxAb0B8gvuJ1/yq/Yoi4y9qDr58w/2n
BE2MgZWEPc6ps7qOo1yvYePALUqeEPfjrkekcqnZ7cdHMBtyORC4DZMJUvZ4tsBBJPXMF/IdHI4U
Z5xPUco1vsdAQEe1E0ngYwH37YSjyxAc8JYbBjU4wzUw06HHefwtv1dQyn56SOD0ne5U1WjUO4Kd
XWEycon9ogQMF90piKBg9Bn/icu/UBpVGOZ07CGz3sWiQhXI5RQtb3r2Cu0w4zPwuUdiISRQH8QZ
vzW5nwir0rxjYBfodWjgyR58m2AbKcU5tBOXP0SGivzNCbECGvj9mxuKXzso0c8liGgaetNq0oLr
9uQ9G61E7HByJqBpXOIwXidS6o2zupj8qkXQ9zyNQ0bVPT4i24asp7L07OF3WktjGSGqoAeJiqob
qrytFn9GT0Cf5ZEAVU4t1fE1LM6x0OPQJXB19z0A+wc0bKC0VI5ms6nbjsFXvxdAIgp3+Ih/U4cn
Ukanmo2SHBeyXm9q/EXSt7UaIQc6ri7Dd7nVwdCwC5TG3rR+yP5hJEhpsTE2vxkMbHEnsyZqwlq0
J9dNlLBo+kUX5oRB8jDgJS2SHYXTE7v1OLIA3ov+P5loS0ymdwegnBjhNfvKUPclO5G8GWxFoVc5
vF/CdaKFmIi2uleG8Urn3i+fesaO9M+hsdWS3qN45u2aeXsautYXifHYBVWJuOAj4hI8o1qqp7Xt
Wjbjz3DCl0zRj4g3sCZg/CbkW/S1o+ENV3wy2n7vezbRLAU4wCGu9uZLyzoIk6/bE2lLBhMm4TIL
pwTMzd4JWm8KKXeyLerW20jyCZPOCG4B/pbBuddRPT/gndymbHRMkYSfFLwMFkAEemKbpzjqiBm5
C6n9S+SeouF3EgA41PxmmGPgW4m6VGRVeygKVCuPnnfxmOQwxtpEfaf1NiGfsXYQwb6eI2sewKhv
g5meJ1hrLM9MvoNuizS2Nvi71LvS32LFt1+tgOrlk76xfrHvt/ulL8ro1rDeaZGQxevQYkencNWb
ZUgkdcAtZOh5lfYvC5fPC4hd0LHh7u1EPgJBe47DLwasWCFcI1QPQyUZZX/ArMAV7ln0cRyw0BBC
pnPWLhHlvE6eFsrqb2bQJF9VieYyluRUpsRzPzkp0e5eAC0kvcUA63dIQBBtN0irUWfZH+v2EpK3
Q2grILSsMPQJIqG6U5153cArioANHCrNoYQrPohja45kpE/hjgzgeQ0ZdozBgDtn5pMfcixTTioZ
n6mOvxkHRVV1ReNGCD0VUFQugcoBKSh9LLHVIludZ2cE/IO1Wn15iW3WWecVfaUOXrWjyTHwx0Rn
9NQu4mY2KRc+jAYi3Lm8iKSRyhwJZW/fd2YPphxI6VNxaWpgSTbIJBdyMpB5+Cg27TMOUrMBuaYx
iUns/4DBEilCDjQz6UbBSquvpES1D+TI+/wUPGwDAwkjbT2sJ+SzpTo5oKwbDw5pxPdMPdmiimMt
6bTHSwFSqPQf/WflorHivwJEXVupgY5amAF41XDrn7PwofC4rS4FMA7cYMrgZHvh3DGEWjkbQklh
6saNZlxUUFvbfXgopbkQNO1PniEVPlfpJvlgJiDXuxDvHKCXuDHVWw/s+uj13uoUnsIEmB+wUOo7
udTw0Cfegi5Ee19AYKuohfsZnKnXTgXTDXDLKn+imbH6AX0jVqI6cAae9KbnlWrx4qv6W3TeRSgH
QhO8vKfYCPaLjFRNoh+AXk/RIb9BPkun/+ltqry+9xtj81Dhii2r2NW4tAH1SUjfiWrjxjet5uYQ
lJXnSzYoErASxoFPrKccd5Fl2w2a3/hRm+Em7KWV52IHWrA8/RmmFZGFfvCY0j8r6yd8LVq8wqn3
Htf9uIagaDU8GIYVc/NNaAgWgtMLVF2G0neIh7L6y5AjzeWa+5ePiIdMs+YuLDZDJDd5arlYO045
W5hnrbcMIpXpHS9r0SDFSS/CJSMUH7azHKnPHdfdZa3HmU0ME2P2KS+8AoHbD8HuMWzC4nDn/ciM
6B5+dwYDQcPZAaKZKZWEZtcCi+g0FZzYknAN4DlnpnHVTVtIM6rE5gjrBfSY11rR6HT+vuLUhqcG
Mex8rueFNZuBVxBjY8afInwI9wnZMkhJCIfZ6v1olZpGZrDpR2VK/RcCmAjkRIvQxn1S9drqxZZI
S4JtiF3DDGOEtq/0nQ7m9WVWVR4A+ckTCBE3NcWDB/BKw2Ty5xdCegN1KPPDqhAehup4ccJbfnic
ouPUA1D/yABROm5JZEI8MIVbc7xtpWoF4TbkPCBE2BYgG5+1nkVyoKSmEi7tkNWBt1qq0egjIwQD
6qB6F142MJUaxdcJ+qQZuzMieooIQ52UeSxzFaSwzEnvxZOhu0dhHnpYWl2PnO0auIwErmAkzoL/
Nn8/iPuvBUDUncwxol2JICgvk7R5v6jETCP+5tLUZRIb68T9/ccAX0luVBfqeSWZQlY6SYOw5ny5
QbxVCZurPmWGgXApA6WJ4SshJsxLuwfuorAT+io4GvFm2b+NKw1BmCaMKnMnnMtJHrQgiJ5NuXie
DD78UmHDs92seL43UIEE97UigmtC4rxL44dctEWKIg61fsSgN/bhR2mDwk9BdJyqomSNcme4P/z3
SDUlPUDTVrIhKw4EI1WD0e1HnVz2q7hPivsBfZm6ElgqBdbzQuJGg1gYY+BbhuMVqU2q9QShgFa9
dlBB8+avqM/AuUitg/EEi+CObXNEZBPh3QZCMvhgQioiK/LUi2BNZdodGY4riPOA/Dc0K/tqx3G0
j6UcmWbgpCsaaPbYMI4cm+mG7i03rZrTY5jK5fbjEOYGrx/jCyq3RJOsDescZMVzClLdkiKR0+y4
Tg3YYTWgmkVmMlRKwzeSoI+on20QioTjBXigsR33A0XV/8Z42FjJOZJN3pWpRvZlQfQW0LkiBPQw
qOKZRTKI75AAnRCUQNKff3HypTnsJ1Z4KTpw5Td10cYdlKcSl/jSX/Jx7mvK+KfuGiEFS9r4ivs2
B5uNLCLmWWAWBuvB9u2FtgQjjoo62lkBsXUrP5b7oz1vo1chXs1fSKCw8MtuNQdsg+WUlCscsHAs
qBO9Tl4C4SkNHClaXi9Ab+N8BKvGuVBQbvdGrkWksiB5XwIT7QEWGLxZ4z8RJ6fw+hXvhj792rsO
Efzv2/dvrMkI7PfUc0EdmH3iN97zXyroRXhWyMoM4vtBDCD+6MF5i+5d3RmgiJo9aOckSqcJustX
J/kqG8xu6rqBpFe6p5KY7k8rzr0FyKBLkRB90jpCMD5Uf12uDehsNbjA8I1+TJF/gTy2Ku1K89Lq
ZBYLMyEpM9WjTPfQyHOgBQjZVq1WgvxPk8yy3R6p9oeEIhM1e97Q98sjf5GXS2abg2aZm6avGB5Q
fepVHdD/LK5TzQR4PnKNeSxa92DlNuAdwTiQVBSNhNGTQefruPYm+TJrT2cRY64JZOQI41uv18TP
o291uOyvmKoWiQqm548RqcaHfbEOwaoostm0tSEvXyrialczk7EyiXn81Mr2qZqC2vWj+OR/bhZi
NkCh/huyBUcuHyetFxfIeQqZO+5yrH3I8GQKLTWLT5rIrYZMXktMJrk54YXhx6pAD33libvQiEdn
cHgRWwZiR+0S7GtjwzU5ezsVBXKw1R2zUqo7BY0d8eaovDt3fJe4kXhDpYl7FNeg+asD8IYwVYo2
oIXJoBTyN6mxzIlL86CMQ54c0MFq9S+iNklqC/S6IM4rdy6+CFW2Sw2pgedkXZ4x18uGyXHrTQWu
noIEZrmFS7428MSR5+VXLJwMYpHITknQR44BUauTAlz7Iug72yRqWt0EqyUrUgmCpMmVb0pfwesN
Pl99gX17D+tHg/rDQPSSgX8WJkal7W9qw/YpMbpa578TRxNhXfJPJk9HisWCWSwF3SicyP6NCuDh
lKGf1BgNHRNbSdtYfgecWUyuvoG75bcqggtbbEsyVyXMnYDM7UVeSJCIO3K0Tz+xtHjkggNqZGL6
oVgtMKnmZrkjr5/gQZF8+TRlJiihsZyVsPa2hvPtMNFOeYWwFHH50KkPADln3gtHswZb5ZNw5wj0
fhk+BlJO2n0I54mo6Qy6YH710Mm1XHmDnsbuTy+Gnf5RYrHfjUeVNDU/dS94FP1ZiNHaHpbQj7o6
3VNG5lstWmXKNI1bwcaqMcUVAnGDHyCMwc0s2FqFpZRdj3yQ0PKHUJuv0DzgMrkxU++rHf/CxWbt
frxvCqC2Yoylxm9Mc8gNGhlpmWPwzni99PRWD2K7jzIFkchEGGyMuUgA5mpjXfBOWllnXadMZ1dZ
mMfCZA1RJ+/Qpjk9V7xcQHUSq8ZFaWDn7GgT8A0mm6iXi3gCZvnLinn/tf+qVkw0tcFlz1+G5+pQ
MHbmtaTfx78DCwmGgJDnnQOYJBlcMJWR9crH/hEb0uLjU793cvTfccxBqG9kSyivvrzf5qVsVfaO
zZZaGdk9XHUC3O/vZ7CWjtrchORoD4QPiIHpfym6Oz2VSWCj7cNsuR/m1oSuWydEu2F+/GyftbUD
1Lc3sbJp/eV/iDRpngQ97SeFSUWVOl5v8hjQOQL1a1Vt26sQInHU7fZ7nmq5vGT7nkKYkrWaCra/
OLw9Wh24lp6y3D/lA59GBfXE99mf7En0Ja+FQ08seet9yCnYoB7Cx+5ErNVUjfbzdWKG4L9GOr/r
tY9iy6vA1HH7Ci7FmoGlPRzeVdOFF/BeW0LA19o8h1+VWx6GAwy/avzSsgZsvBzrK/FVfwa/U6ek
P7K5vn4iTkpYHnrA36Bejdn5WrtbYKLOo2KTx1s/Uqn8LFXtK3V1IXpTDHjcMhcpPJtT1VYSXbkD
6lu8k4f/HyELNH5RKE5rV7pRLwxH2G36VipNH56d5Wk2SmvuTOjsGEEvWrVVtbxmNEMT21u8lkSM
ZcMfvaI3NayBTMPmxdxDxcsnmB2Te+mroldUJ2K50TsircFCN6iJitgaflB1XZnDFoEV3dTm1CSI
8GlEk2pdSaIk88LAviWN3nurc8z1TTM+m+2grjVsWTmOvJnSLon5vLyQKfq8fVOZQ39WOws69WMd
9WA4xF5r5pF+fASDP0ItixL20Ir0rgbX+IpatosHnpBiJCCPj+sSQinslfLW7rSCbw7FCdlOVctl
WflMovLLc86P96oBZ4z6PtLOp2GX+ONQEnycmvA9J6KMcFrAvF9TS7738AMEPt6KzfEHf1AFky+7
TAZYbYHiOnFDkiKb7vOqdqP7Yphfr3oPMzZ3lVtajlaF7k0pJF06tDDVP2/2tV8VhWlPGklpbKR6
JiBi2UZr4vGL01ludQJLLYUPxTSM4yjsUUm3EKHVDZz7JfqDHLeDDUG7gaWeIb7Hhw8klBkQ7t+6
v0qIZGWfaFT9Y9cWUMZIrKZP/9/1iIbRAs5xsFiaZlig5otHM8Ca/99Un3rQtY+3jMHFzT2GAMz8
g8jWXv2iVAzAXg17RPmLgvVw1A/zXHdNCIeC5lIhGuGppgyXqKXQp+XLhKBE8s4+66riAQxrjcDU
bRQttVVqG4WJwHluH008DTLgTHt5qw9/ZyzXoVUg2zgs1bv4dvgopomfZ0Lun9b/8YSHVigKPWJw
pdni5S/C5n9nJ/sN+ehExeyKqD2D2AXjgfnxl+ndaLC1TAeeaAabW2lZDdw0zcQJmwgEWV+lWBqR
MkmwqSyTcvL0tT4He9mlRRDfv4QQ0tXcXA0ekGElINy670Quy8q9fMfEqKlBqx/7js/oMznal4HY
Ll/DwqnAFwHt0RFmurUTLaZ6HVqwctzt9pncS25f+gPDnAjQPTTeve3dhmU1loeQzJfH77phadej
WQ7wDelAUjiBGpVu6Yp2dYfm1KupkCbeeD+z6Zk8iS0At8ljbg5qiqMbPZh+LZ3Rjpl/4On3dguM
PUyvTer2+X5rW+Ol5ye452Tbz68cVYpif75MkNL5WD9t0C28BZiNkVrI7igg3xTAt76jAC/mxy6t
dPjMcEoTezPbcKwzQtOm3WfkPJlZKtjoSYfw6tFpz2No8Hpkn4Hv9Ir2rHDwmPbCU89y4V8Q5amp
A/ebxIf2rwf2J9qEcYaEhpZKOrAheU9Eh55uiUOmlyIJgZNOxmLJXThYnhEuQLtgYE9Mr3WA8NBR
JIAJDizMiMJPDCcX3EfoFFEYydi77qslMmKlIVcaZ3YWNQIyT3XPpYDczMIF9fplFogcs6PuQKTV
Th2EryoepETk2SCidmPRskRQ8DueeC+13HvSBemrjqxiLScrHC2WqSLvE70I2ubO/SNvedcZ3vH7
Hsj5AmPU1HyRqrqx8mBlcRks4C7NEj8uxU7k96j/jdvYt3uOWVer8PFYYMSu5gaH89Ok90rydPlQ
rojmjwoFhe5mNVx1ou5j7enqoZm/8vWCI63Xk9hl4voNnFcN7RTMDuNRuhEYxd9NeNX+6ZYMwPB1
WmfSfEecmr+PSldh0USpqGrqmXS1skIGjEiyEV6i5j3XpKLkMOaVcwGliju2LisjrP0seT2+ArAK
taMVmW819w6T83e3+sH7kPfFnIHMJ4Yr5DgHMwPzoLQthVDTcKPHzf9jD3gRiMMtS24hyzEhaaCK
o6TEORoquRtgYmJlsAza5KwrKCi1ajcXP3r56CqHQQ0GaBM33Ustj0t19RGZDMcFGidoNsmLH56Z
e10C4rImitWzG4/3ffXGfOw1/sK8swZqyde6yTtVal6S6+ZppAYIXpLZISfi022SRXnxcNs98pP5
VKdlHbtWpY3/eouy8GzwPRS6yFyC1Vi4Pu+a7oNrgivcJWVxPGL58gYBWGQPKRYVxj7SlpPIM8hc
M/6tZOI1k5JIrb1n5GUM2Dssbw55bFofRt4Y3CGqQQ3rxp6gIWFPeMjSp6LD7RCBre0eHjXIkxZH
ygeDC0YRIe80u0Pv5azPbwqQ7jmrlUhqwHd11l4nuqFjITOzh5ER2TsXpLh7wYsYcVBJj3qfSGku
Zk3DR7oDSv6GtHSE4k4tcfoK36GU7vpfS6u8wcJk+KMwxcKmN5TZLCllpAmIoV5VKwSCEKMYzWl8
aSMTW0OvVPw6D9kf5IqOWxjRbawlVLPGmC01FAATJIQMXjmDBULKtpn2v2o+VoaexOb5S8nd1vuQ
1t2kgWJ5RLzWlLMHHHFYmlWkh7Twn6xasm1Uca5r0AhAIV31MoSUzazAqQk+XHMDaqrVT30SsKhy
OH+DTarYGxoLLYLKq209M6PKAt+6Y/iJiSPiYwKqiwYuWjRuTfbkKALYhfwZWpTpiVyZBfAjs5mS
JNSfSD2CZjy1nFxulSEzZNKLsJ4hq29ruuKZifqGO9HhXhmHtYMvrl1U0izj5aj9Iv8qYuf4ECfs
95u+x1Fu40eCQ1kilZlhgahoTD0fO9nXbmlhV/4YOoWUkUMDf22RDC9i8416iLvywvjgvANkb2ZB
XT/hm19s6+JNTxn6z52HH6KrD3gxinV1NKFSrBGL8qg0rv2NjYPidUe5A4RHM5t1K8Vmu5Dmli00
BBG+rux2trbljnGFKWOMy8nHrwdesgk7HnsgmTaWggyr66QSTdWP+8ZWCTPxv1AbS5n72V9uKDvO
kj7MV+o76gfPu1Zi6tQLdOpgGVzRiNfhOwZg2ekVO9NgYjfbMmo6nRVSlbaYoE93vCBO2DELQAw+
RK6GFK2Lw73qA2Ww+EX/7R9DEJ/UhTpuhvAubPFxCFka6aPo3ZhmAuKbfhRIWSnJKUpRAP5qsBtq
xsnBWMCtClDsRH9okWH+52Nn6ZAGg/CYJQh+oKB1ggnDAWxw3FJ60piyxkrRoZbuYdt4kDCOMTwp
new0yWRrnoa+3Z3RijUIlCYBOiw9kUfjCDoXYiBICMGDHAuiKT3rDcpWchZLogzrUQi7tDH5gq06
PCxo2QGp1eGXF0IRg1WCBcpGscSOti2h6X6g7Zxv8TzfUalzfkReu6DwfeF7hrco1pYlstuZPg8d
I5BxqGLXAFIGIkEU0KCML+SKzXyytuyqR5Us0sRH5jO0J6t7mOtfIAxTHQWVCcsrUj2g7PQjojz5
gH717HKgrBRTfa4ra87iz9Gl99cjev0kPkY1g8s+/PArrgts6NeyISIg5/g4byBTTyEjGS2YRmOI
cTwi4H9QaO1mvNv44PwLtnbo0/KhVA/CD8b5rdoa6FPW8H3zw+lhSuOnsdIg09+kcnudOmE7tjZP
CPsFpzswSa6p2stkYVdGvyutNx84BMGULzo1gNqOmYz+2WM9S2C+hqCF3CyFY9zhBgDsMntW6KeM
t6ySewnvhBv8KYQxd3nhwz9DnlNct9ycft3jEL5bGgy23MyE/rwOmA5S9m3CPiSGjfu5zF/zRh5K
rUv/hNqzfz3UASoCZpiEjXXc3eaTd7/h9M2BnZwOq2Fn43hS9g5Bs1bTcBVf+S61u0pwHMzICb8v
US3iYsCP8p4ZgmSGfu1Z7FTmvSyldIzvSVqcVuHIopsh+6KxOaR2UMHb7bsBGgC9L8Xjq6mbHK5Y
H+SUIMSiw1PSyn8jNtAOdJ0tYBuYQ0BTDMtchdLvIrCBJWuevFl8lHvjt3ewmYyAiqMbcHlWF1JN
J4hoM/mde9lly1CFIwYpkLnIhDPDBA3gju4vkWFx4SWPr7/MKTe5nlFgMfFwjIcPlMSj0NbwvibJ
CLD23K9sTSJqLf+qS6I76C41HXyYGWW+wTAJ5iSgVsFihAlAo4I6kCvvOsTtydg8/xmshvBDE3Z6
V95kJeeAQCjElHnDcr9Ox6SoRc8Dpk3e8hW7nHz/9kw8GOWYrbbgzzLzY762QtaLHCbrYKLmqJOT
vW9WmYHW83Fn0zeWs8Cjr+/fxuQlPjQOSmYehyMy8XxBik/XdV9ZE2HHyHZ82i54CHaqXQOTFS1D
cc5HgbrWVxCEPP3ujPROOWY9S0w2d/bSh+omzvqqSzNWNbErH+C+ruLg2/z8sQR5FBUZTibQj8MP
iLfhVA7anVVqy8QCxyKUStL/NAFaq5HQV8ZHJliGXPp5cH0ik1bRZcYc7zdJdxQgIWsKMmwzGzsj
5Uh6yPof+1jIN195GFP2yD7cQsaHFHHBHdF/pgyYa4oK5PbH0rKXJpWsu60iuLADJ/2D5U+boqcL
ABpblrPO45nfyp5MfYnYuDlrSnd0Qi5dT2MY3FQDU/lDX+NKugxT0ZVM6pR8+6RTOZ2UpJ7nGCIQ
VtvjWAi0Dm2H2Xz4Xcc1h402frU8lWONEOL627AaS2DjS+mZMMVRtUfUYcJJeLvzj2CrqbFaWn2R
1XLJpBbi6Yiwpv3IeE4Od/HILbAeefswQ4be+VvPjYF0IUxnz5wBumvJcGaHn+9xUGzIZ6pwvcqg
Ojx4OtokTwifhGk8ee7kMNArndHE/0Ta7bomIFQ02zrHDctquJ5i0w8d7r2ctWQ1s+CHbni/14RD
wd/ZX+9iwKU7pgixyjgTbN8BhrvNMoVIPR7TIlsXtzNlTCxXMRQCy0LDrjwh48eWYQ3d4EhsFgVh
tLYZ4mGRoMNrnaBhILOLdOqEKQ9+2TRLVnOUFmnzB9VssrFnmpxoS9HaVb4xq3EUo+Xa+91Voeaf
+/Z90n4CA4km5qV9JoiiPwquOKre/lXwMrHqkZv6RiWyWCXfBxwHdnJGFt3hQWTKS/02VfiFdHY7
YfgO80p+r6azOAFkc90ezd7ntzsyoHU9cdWiCaCTYVB6ApDZ+PyBiyFx7BpcqEKuqf4P1UiUrV7p
Easn8LOLjgr6vaGLX1iUs59OpxQCddJyXqGWLKZKE1oQk5QD0yoUyvhZk0N8m1qINLKJDQnqILm+
SSG6SWQbD1wbClJ3HvRfBB+WKgYRtWze3MRIwSoxj9sN2PU1QdEEbWa2pOQrQAUzgeRckZ5ow8Z6
EbwyO2+g3Nv35uhs2wB8k4pFWD4SHzac3rM2LBISG4Rj5kH//u6PMqj5p+T5YXQwZGHzErO5zbsH
17oCVzgZuHlvl+2JoEpPn/wKioyHA+nJ9QZEmRswPtQbt1bXT633IoEqxXpIiy7bHxxtC8Ew+TCa
Uggy3coxH/Q7RkyiITNY3OuNEKekKrFVhJhIqQEtYlWT/IKVr9hZJY0gMJmwaH946/Jle0eE6qPL
w5PQB0bgD+rGolBqlI5Jy7hxL5OxTkjYFGsEOU0tof/Qj0Lbo9xwvh8CSesVK4LgQPco5R62Bv1e
fz+ie7K0eJ9bHE0eM5vdaoacd+acTHo6sqmyIVmL9qS/mBDI0haMrSxq7nSJ+pThayGq0dSWE0qP
mt4psGabCreV2zOwkP7DdxYaJdZ7MUZ1Rj1fCANLYn9NlZJNIBO4HdoO0DwZvqBHF+36NDJeDaGY
zW6euJka94EWo7a2Jm3ZgeR/ZbYRAWm5omKT//UilL8aB9AJq6ysEcoPmcaZE0hliKtCBclm0H8B
ylxmU8l/QGt8tMuUPsBKLyweDsPWSzGc0YiSbj7xkhz6p1muhpUsUocrZzWhA00hoUaxzcVDkna0
Rb5meEiEBMjAp7ZEMiZKCm5Bnt1lanGwZ6pyiUyUFe/PXc7BqnSwV0Rgwlgs02MalhPpijIAXJHk
wnA3gMIz+ONwPsWrEYt+PbPSV+AWF7OSqDJBvyNdSk3rbhdMbBd5d80XlJzUvTJJiCKSqkoUXlw7
OTFcYcItYeHoPw8sh+/lAwmRrPynbIXJCCKwzcLkyoy9WcQZ8wI7mLgfYa8joMgKtH/3vgIVmtol
umtBMiitgNXz2rQTKMlbSe+RdM8joe5L2Er3nOWylPP7iIzUIfpde9BWofD1gg81jBLkkEH4Kgvw
a4cJjqGPNy1rR0+4sGgznHDUuHvCgT5wHflYWknDI83T8AlTynMpucsJEiSViS0UVqo3q+FsWT73
wdEcIuq0uTjegHqMo0CQ+TIxExknCqHvi5duRZh4ICQnQhpgEhEFv8jhecsjpvoDUvu4R22f5EJS
AYwk+MYHm5yENLOM4jwrHlrt3Hs+SCurN7+5Q6yC2hNYyKGYIbKUxScdTi058dWXBwyd3mAcDg1A
607iI6F8s/kQiMDNpvv93Rjgf0HI6t9uNwY31dNrkhuGoq+cXvfmw3YTnFGFt+JsqCJul7EFZa3G
DPM17L2/hUYzCC6ps72n3ZrHiVmL3Rc3ITzod0VCZnaZFd02dHk4Jyk7TMnl9MzyKv0kxLkxMHo0
1BY/eW/3Tp+s4jJD2zvU5DNWkbhn0SA/8AdnB8sV4I6Qio4p4XigY62u/hzDUFsyj/BiY9mUI21l
r+BKbOOkvcaM76K8M02S8LTNf+HkoqJg0aJsbh2oyT/EYw8qwN5SX+hNjk9tq9sBH5XYzHQPKU1N
keoAxXeQO8QF4LzW8yLrvxJ6EWDM6OZvvxMuTnixdY374csOaLQnogy2ecQ6PLYXJe42BRQQMMad
Lfr+jCmI/9BW/3WBw1euZC7WsHmp60ur+khJx+RMPffetcPZ+6XPm+j6yuTSZpw+ggo57x/AUax+
AGtVTEkhmuAo2XuJCiyP9uDhpwTJ6sHnAOKbugN6jeVtXNNjALxD0+ZvwM2NwuCXZ/LFOaOstHji
gbyRLm5oWWqp9vy7EcH6B70Wo/NAw+MTu80b3Tn+mB8njFOpGrlGSBiaEI/t0IrC9kDH5chLD2Sa
hdUs5v6Kyv+c2GiMirbBsAYH3Z9bv8SyibrODMUemUlY2AJPTkqSWeLeuEv5p5ZpqJPpnrV4K5zR
tI6bBf/wUQe8/YXPpYhfBZ8WWimA5d5nggfCE7HZP7svbLxELNs0HdcwobbNVbCtQqXWNVourNdL
/i/n5qNPBYAfviznoL2KMoFBlR5vnLBFkxSSnM2zpDxrliC19ss7cT3cw3x/9jb2svt+kaC0aiJ5
OZCSJR0jLy4eju6xgKq/KXi+NQhGxm69u6s1O69maqnun4fnLHb7QU3Cb5qEawWEUAdb7GEXVQoJ
opd0MjBkTkvsr7NNwzrPOG1y4Gks8MqAVlkcmzQVgo36yotHOeosS1fb7LmJahsjETKIpN0HZLbT
04tDolPd/oc2d4OzOtflJORVcDTohYqLP7WBlT2YrkqLCJYEDa1ISpGr2KxM1RTVOpyMY230NkDY
90FnM5J9annVOCZJVCuA0xF9Ub4nuoCc9bm84XFo2PmyF/IFXlLuCacZL2C3NLX+0ZUOP01j3iuO
jCn16xZ4T/VV2dJ2xXYoJ/jShSi6lrj6fBFJNlLjpRHbZqOYoP7KMj8qchddDqesMzxxzlGzPNTY
y8/94AJZICLcz1IixKQn8pDuuXY+Xs+45q4R7KS//xFGd1qpKcWfHVRRNiXRg/bbDdd7dD/24Vwv
T3uXcKLpbsjOAEwzXPSgxMziRzlje/o25dWhXkRmBgCAXIUU3PmPqxWq3kgMG5cYg6feo564gAS2
w/wVb9pXAKl7TR6LpGrdEvOvJFpaqYJ0ZBIFCscSdzEWLajMQurSZ6LBl8p3SVRY81HWHEr2upWm
8wxiZCemZKowyszqcUmb7tR6wigXUNr67Q9d/8GSwGdJkAO7T+COawAubufVXkL63WdDE6hVuqTq
yk3pNQcPDESxUgaG5rzJZMRPqIPOp2jT+oGT+0p+EA/SXlYfux+gewvwChVmsdJhdpxLg4iYMFh/
a9vUWXe/Et9FLgZJXiTbanjwdOUh0+gHuIte5GWEf4YgkvPflaCjSK0QVHNVZlwiKGg+DWDfX9rs
2aKYP23XsCxVHydHHEnyg97pUVsD5PT5ih8f4bjg6N429PJAL46XcaRfIoDQj9VNEjFk2RA1kurx
hR/7ProKwkd0r6P9XveF3YnLDO2Pgz5VMIptKo/QUukT8PLbVS+Q0Ykv56CvTGfSsYWq+rPVFR35
F/s+yRvBXx5Hk3JuqBZQqFrkcq0hecnMCOv88vUbG0UmwI9Ab2pGUGK7+pSxraoFNjHEV0Tni4o4
ESOafVvJcABIRrdazMmh2mU0fhk/AeDWpjPsJJJPq2htf099QhMgKvZNoo89TXH1cwxlGpM4kJKG
dHSXLeRI0evXD6BBN4a+kwROt3GTLb4KHgL9nFm8z11p4MDKbxx+TGi3DdWgae3uDEXdzFMJ9M7v
bnTjHGiJIHSef2PIEeo6tBehHO1WnSVh62kQqPHOIU8UyGXDfsOq9NZX/26j+Y1ciRN9bd6O1I6U
guMh8KfISzQtxpOKRGbqIUicEZeKmdUV/KoKP4Utp73MelI4QweswHt9qyZ5G19RJURYvbM1LfbV
ojz8CFF3eaBnNP6OM0VGpjfsL+eLKlDM7cDIIcF8z8ImEpKVJnq+LsyoPiFsGDq4hq1S8KFszEJP
kcVkZzJ9V+J5hq09OXVxpHJTZ74iELxQP7TRo5vnFJ+Bsbu47AO0nugbFSi4FpYnFG5/t66B5EvD
RKuHkQWi9kf4FTpd6b0kzQeKfXZZBx0U/x2Pv5l7AvkIbTxqqGvdLvp0iilQseSgT6GprYw08t5k
8Hj49EyKs7ww6IatQ1DLPCPgcLf4ppzsru0tyBwdRaA60RD8zrWanuyYyD5v2SMgglEY6K4BeH3g
wGMh4peo6Wzdj6eAUmNOY0U9Zd0VtQgy69fGJ1fWJtJ/wZq/wQseRHzkuQsYMN6ynKxtzR3ebwwl
S1gV46/qp3MdmPm+31YrzB1LGaroFyeVXXMT6UApscaTD2xk0TCGRLFLSKk9h3ZTgiU2VDB4PLTs
HioNlMcQ0O2qBqTI153LKR+pooauC7IFim5umCnODKok06nlmNYZOYMnxBBcb+rxAJWRPXUtKg6V
DKqooYfkq1RoBuJVnbFOjtq11Uf0VGvAObFkx6l+RcFx3orzk+OPi1SMA/Bd8JwascSwYtNu/KU1
aut+lrel9c/9dkR42abrb4yGBh+7Rzo1wsyTcaqOzbBOS3QKHkPL5udgMA8cK9/GLgqzzhDG4ire
+8phj7D/2DuHr+lxfKnEyhJHQtXOFoWtOAMt8OGzIXF0SVfuE9t2j373eDDghaw0SoJvwqyxvlpJ
mrp95TcD1nZHgMyDj4NqsAn/RxAzhvbywVEZsyUgtzOMStQViGxp4F3ZtB+r/67yfMFcQlAPfJ5D
hBK9qshiOQi6OWLvHzJbIs9cJ+6ZA5Nj75R/xWo46Da3FxZ6kS2WlFOJAr3XED483/X9bpqHPFhG
eoGS4ZFzJYF3Y3IeHD0GwkfFrnwzWD9c2GDED2C5pusMTk+pjx0mzneRe+8HSWdYklAdLgHkCnPG
ndfLMjgKXRUIlAITAn/hMpEjwqgpcvYsEANVvVsHBYP2qiMojSXu4kFXLnqExG78Rn3xUMeHnjU4
OG8dAcnQH3phO0aaSVlG4QI2byBjaC0vu4LQjP1/De8AEHvtEnzdy06/W/zrI+d465r89+I3Ym+3
JcjOCgM3o9bShwuonFtOozeAlt8725+rvZy7DmSefavgb1FxV9/nTjO5ehEmbe2uVnLcZAEMFwwy
bVB1JvWAt6qk4gecXAz4ByX+qU3bSP3wkFBXrFhgEfGc8yezXDsDv+ySdO1bLTxTyIK4Kylb6Pr1
FKvTFaL9PNx4Dg8mYmW8zKUdIY3dawnPQZEtyZ3uWgfSnm5R5vv4/h65rlw3C4nE0zhPjuzZJCxM
2J4EezO9vgF/oKFPriS6dJlKVsTy9MX64KqAewg9GJEj8Ly85ExCqXGVcGw0dznvUMU0zcIenCBn
vepFsyh18VtgImj7k7cXYRB1/JYocvEcRrcXMq89WvemS6FUYT2G38mh5mJKcKO4qmzGP6513k7J
3c6LRAvOjDS/X8BXdm66yqPVspqmsizxpItykBvKSrolLcIJuFWrgIDq4W4uBL1G/93RASsFg0QU
5t8dTniMpe149nnjmIDKMY2F8/CEuwuaO3E4zuxdyPOt+CSjB2bdZo1HMjwUpadwdwQi4rsDoFgl
U2oT4NuEkkSwmSjeGEhNTSmlvKaelKt4idQZnnl6UZxLJ1CWdgOc+mjxgvWYHxPIg1DhvhpJy3Pl
ew7PJYo3v34PgJbRzHyQsLI3eq0wqoBRifLZciVzNQ+ssJSiZgPIJ4/XL+5ux989QrVEscGRb3Vy
LzZgKKwf0GwiZ6vGUc1VmH4nrLqWGHddd0ygrTakghM/kI9lsXwf+sEUbGejPSnm10O8OHMWbGu6
6ELFWG5SMrK/b0WrQoL1IohN8fs95kJg24lNkVvOYRY7W6vEMLpRMCIaARER6cg8E7vHrfdqadKO
tPrukiZoSQzhkqBkn7gfA38WF7fW5s5mQ0mc7ei2sAxFN441WQ2ERIsuu8l8mAuGc/Nh6SQLA4OG
55s1MLcWXZIXgMkMhVwMOnZ//xA03eHSV0nhRCTYvVd9VfQWylLGSOqhyipx65TSdpVnM6ctTA8V
IXmJtDsOFWDOsdMciRvrzWL07MWMH7IjqC2WiZTH/iEqaqDPoXEtElfASgEKrpSWRQ4o13/+5vqe
jMumTl6M7WOJ20pMT0RXZ0tnPJC+LCEfD226PXyp3FufWvInl40NB/tzGcXsaQXI9+UGU4MMeW+O
M0KOp3CXNL/XDJk5Xo6tXRZbBIb8NePsDbIw5/Kt2nDDwShmFqKCXno99GZQ45sjNvh3enUjWAN5
gBaZOgTlGOMhQ7k9L+hluUdPsrrcnJMmh+tLV2uIuyMnmW7XmBFYIrjMJabZib8nJLr86JVRD9aP
N8SkX3QSMpVQPucHzVcuGHALNIAZ2v1HVy/SXuV6/GZjbwmJOa30aWYS7KIpEUdIrAtnVOUMLinj
8nYJbHKn2Ub7CiTWBGkt7tVUwLJ6VI39WXSYZkPZso+PrRSjs2XA6xGlugXdtGPIED5UWhRu6iwr
OdJVaDPcAZUIL1VOQ9Jmy1rxC1QYJwtdlSalVKY8RmCmnlpHHVh4sqJ6xXecxu+2py4JCs4zy6J3
R/DkpKhCmkbjqFCsR2NWavJKOF/kzEPVy+IwgXudXdiX3Q1DzDInY+VG3hccvM3G9AzSq1Zat4VV
LRUy4Q/4PqO02SYg0kTI7VNyOXzB4RcHbbOAqK5aoqiyoTACQI1z26egT77gt1GNMN5C5dxKJAGY
MNodYQ+7jigEQItuPcC38FiKbC7mLiMbX6vhSMHdCsHlysojTuOY2arGonY6KgniGViMRfdLpdys
9Kyls/pPpCdmNKJNffOJwsWRmilrMkXM1tanTC3LerQunYeMnkbyTjLUwK7dD6VTJO0iDLozmXLG
p/RZS5v8rI2aSvTvX9KsYoreQQp0bD/9jPuB4djgBSwX1Yt1IL+T+Nz4vNIz9moMHqe0Ot4oDnqI
ud5JihzEuFGDzdTrqmMWcXozzlkOTN+Bw3BOTFXFuyyEPAO0MQ7chZE0ubDCvY8bSvCmqDzMBCTI
o07JUIdzIFQo3OgqxQPGrabP5ql+5kUQom6tUmXBb9YmZXPyNg82gIo1vRUkPrVIpvB+4PflBQlP
jxpJV8YIFpLrIJztjaZuVBYIeJ+GFSzRF8CVkFWqFxQd0X+Ef6Q1R4d8cw/yW4UHpx/6xc4IlxZS
eXBIHnwUrg9S1oSqcveZ8Nt0DyMy3IRzz5nNYMMJhNg5zmcRG0zGR4V9pxVzFzbPAo43gTa8lB2K
C9MmC4BX+6s8VoyF7+1KBhR6Rqnh/ju3clfvod3hgPRuMfU/UwltEyraLSwM07Ys2rqFZjYxVryf
nABYR9//sfmSFx2uR2ZeczyHOTOcwDUJgC1OZ6ZSrzkEDDfMKnMZvjDzbSbWCdic9JO4kgUnKzba
HbDgnEYS28pAcnraDxUrq5e5zMtRvh4dq9yn05dknROv5Fi+v8x/Do/woEkLzF7vysPHamBEcY5O
0K2gCSyRk6bY3xnY1ENhdII2xdLUY7zO0iQzVTmQ7loGF1EZ3rk1ZGeXQXFVP+/YkPlp1DoPwyvs
JdVJTX0ScISBeiussgI7TyCxw9uxfEM86XzokOgkwEpGnd0y96ESzS2SgZDacblC2x5JYBb//R/P
Y/wj4AilwGRtODy1lVrnWgANKAk8DQ1KByptLOZ/hwlVcL0g69qe1Xxh9uK6LBV+SDJvylPXg8Lj
bvAUWQ1uxZbkBs5Gljy/eKXC3Hs5QOtB5pncFUVsu1WFSfnp3ml13lm1UaqbQVkhqazXP4xLrnEc
DOJyOyTXoBZNUJcyElnbP+LSpn1Yeslq4J4niFWPtrv1muEu7nUE3VyVivZ6ncpbwN2r/oJeFifY
vtYR52VffBjHmEN7qKgReclJALWZR0pP7MEQ/PnLP420MeNxOXbl78TaVRGsWtHZvkCBXJGi+F9L
YNx8rx/bumVlfb9tjaRWWHOKsSyL7EZmkKfpztfXx6VqyfmXDDwukAXq5Ayv8iPIvPsg46N3Gwx1
AQgcoEjR8O3ZTyqyTy3ddZYvBXIu4YjIsTcK2CQhfzA4FDaDn2ANOAqBC5N+BBfl5BdvkedW+sjS
mJXxqxNNiMkujqoDS8xjrUT6ub4o8vjLidfAIPUK35e3LRiDet9Vh+ZwALo6ZxLd2Jx/C7xLnQit
6SUuUFGdQrD+hZgu7fgKODxdP6J95uRjsTqoTtV069eXtpzmmntkhvofd722BRCoqw1jBcwkfMfL
xNW1IGKwetF4dGrjGA0DvcTFPWh4MMj6BMghxbhWax9QS+ruk55TWIzs0cMxcKaE98TcIZniYHNP
C/ECjlK6Y+Aezkse8Phge+ldkLFK3xKvOSLeXgt7frUnvfv27Z/JBXYv2nCN8+1GhoEebsxxSbtS
uf8d71WX7wispqdoMrQrEqJaKfVWljCH/oo0KtR1S++Wz+QFw/0FDPaQHD8KnoAvae37N2yniNxK
WJp0OzpQVzzkFWEY4+FrQ+sD9wZb13/EKF3XTwttDcsp4WPS8cZT63ub2vgbnzswmRA8Dtv9fvq9
EpXhJOD5IpdEVCvcsf5IE2cbuXceV+UfkH27fdYsVuWLu2Rffo2kdexPDZp0Erxpi8iOWI9+P7Le
NnPUC0PiWPrhCUXh6Td/sFRek0dn4GvJ8LvF3P35itnGUKnWwJ5q3W8ty/nHDQ6rZ2Aw7yPeOzIK
/dyRai5znppp8AwKkh0y1K7vYy7QPtsQgxGhbBhVCfFJFHZok4/8axio0H/cIMNrkZSFERQcSZOf
ZU5oiwg10YHi/0tAGVFk8vwFkOzijZ5RJmZnZaQM8mPr6sGVCwqojwCNf7yomiGKfBLpZbqkE+7U
DUv9GXfv7y3G4gtLNFU3lRDgMZHOdHfegJKYQLLnPfSJmoX9x6AuWwEGyTZy1Q2ZLG3WrsZx+KI6
XJtJABKHpXRTc/HCjfNf/ns0OP1rQ2OcjmqzGznjLH4ablAXMC22ExT89wOchzBSRlBovtSiJcYU
exmz2WuEux0L5ZguRwMdg7T7gMb8zbaJzoH+iyUQC9vGfq203khRXBzjCNgfmgIS28SZ8m7wX/kZ
v+iXqBMi/ayzIe7r6dgrI7jB6BiYKUZeU3hnSNaN4rcSnnS0DNLH+P7l9mkv/uEFRDZZuNO3eaPb
S7IdSzSavan9Zi+uQjg6q6W7fM1FEAkSulkzJsqjYTXnDY1KwygLKfYbJKEHfR7pB4id8qrDutyZ
F5xaUyp3EgG3tDuhwuDIhAC6sO4u/pHSDC7K5kBui4rA/CmvdzjKgOWevApTEdFChOL4/ZOcaQAM
GtvR7Omoy1DPOfLTA3kLWghvGlaAtn0kVNaFjfoLoH4sx4LPQS0K6wZl/aGCst1/15VWBV2WC19k
J3p7wRyTjmfMlDnMyB4eFcDH6oEzRnKGpUXPV94hgqCUX9zTyvvF6JvD0ivxeMerkYRsDiGCBYb0
snYwSrFZg6MemzzMTDcvfiZ9rKPN8SIZMle27Fp3sMqKZWz76sEEVvxyk20Z2e9VbVAj0f5McBwY
2w4Jut/y8hyrgrNvQ3di2R/qp7qhM8Le5t6DQZE+bKVVnsIEeZqvZBcE2dGKHDyYqHK+KJeQexsD
VC4az2RL9f6DthvrWUutlGV89v1oI4zey+8WVlPmRfgHG3otyFb5+t+6nKChclcmXNzTUoxtLTQh
d+P1aKZwfvvHjuo0z0GyFtvg5njqltDvMm0lyZuk0R/euiYgn7tzPb4gXpH0kOb5VLH+d4EJ094e
cQfPlcVp/wfngXJUm9K23iJMyhBT6acjZbPEHSQNmawoGr8yrZliD4YHMPkhRajUwu1+ljcOe5Ue
dR2RiIOAH/0/FrJFcJYahdP6HKsQg34JMaCbYJQnrCBkao1P9J9VV17G3nC/1mTu53x5bJO/aaH1
zk/Jl6ypu2ZEW+mJ7jtEatwU9WBhAOPazKm3GUa7G7W8KDrRarTV9OmGzME8tiXjkJnrgPW0aD8L
nuuUxd0swtT/EqSTCHrR/v+VQMvuaFhLNWJ3v5J4DZqRv1tei97ZINhZR88zz6zAaUgxKd/7l+8t
Zj1NFjQEF/tJyTu026Aae9LafTHzM4FIw4hoB0FluAv/kvO82TdZnAeRA/KT3lch1qAvW5YnXVAB
mhc69EGcPmLZSB+0ILVp85rQ1fSgrLMCXMpc0A6aRgnFohn3iJG2iBpBvQmYEuEKO/PVTbv8GZbS
k+5jjwWq4ncGk5Bhjcwb9KE0QVjMPZL41OVNKu7jLBq5m87Dl4sdZmuWflutPbK1sBUG2x9yd7PO
COVRJV9Ec0VddEGhosRTP727NwDBzRitLWWBgunGagwvnwo+hdKjIZRmfr7HkEEZ1GM2IRjI39pK
tXQiGjOssxSu2Lr59Cgk6PGyRzvlme/xhMWxcsWVKhCDDhtvEdEhkb3EMYkFLV+ua1DyEdKk7KL9
/dz+uK9QJf54LFwlgI8Az3GFr+lyDPYvmZlQuufnw74JzMykI35Dh2dhTUOXj1V7Wp15RxlPPdRO
v5X/Wto2tP9mWw1f4sNvViRleDs914yxrmCoRlt/p31DGlyQzOk0B0O95bzewqH8IOqciDEL+g1l
8HNgnpo1AawAIRKE5XjwYIGUfq6xlzTRY4/IrbT7TooMQv/8hKoxO2JE9zJe8a4ejL3BWeKXb9wi
8HkuAk6KNvkzYfOqqbc1agXmRUewWHGb+Yz0gkdcnOLhjrnJ791Qjx4nI/LdyvyQqgIyu4NfsFwr
XVB7TVCyCLNWioJoWbfOpcLL2xa0W5enSGPUfd2vrU8EoEoz3WuWHfjsCSqolT0BjnmeL7b4XSJo
bSnrJwdTK5qNqiyXbB1YnGTpbdCPdYWm5mbSlzWosdSJFkqctMaKe0yaG4TGDw7gfrx91tyvV76X
Sl1Qz7aEP0y/721JVa7E2/tbrCH0NKKfEhDgYCYnF91X8HVP7v7fAO4CUne5xvbbdZzC87/7Xu0R
JtqifPp3sQXwfI1wsFA+rEDOhCSfiLL/Jn3ci+4dXUXLCxl4gwM5wc4mbSq9E7iiZTrMFNLWLP/M
zx3A63UIIp6XYrRPzajCN2euNkbZOc7128WzgWceURbcteq4WWAlG4HL5jJ5RYWk0kK0ZtC8nNE2
7dABwgsKBzYB8XlZqqZWR0BJ+anyb7pB1gQL7VTJL4qIX8ccrUe/hMHVx1edkPed4KhHuvRoDOQD
14HzNSbZvljOXzI3YAfyJYbUSnAWCIrz8cC7bBRkiBlaW502Fw7wunwDhUtv8fuWo69DTG70vKEy
65QSnirzFSHKcrOGJd8qWz9LUWdA3W3oone3GYSrlBJAkqawK7mcjiaXhDJysDImuC8iO4XBdeW2
quZGB+wfvGolmCYGSapPf0MoAD7s1P6xEtPinHKVv8tsQgttZjWCmvNbn6ryGzkYsRb4KFIedDyN
Vg/sYtDta6yzFCmjHDse/nIQu96oSor23pSr+JkHEHN5Yk/sYAwh7r/ejlYDCcRt5FbAAfkHlsqi
kESmUorQPChVoiaogIOOOqFw5DmM/yYrdksWnLY2gwGPxZfDFq0yq1c6DB1JipcuTrzi2d6NmgYh
LxyAKecHoP9yUAu/9Ssif/5gXmhBxOEwo1CU3KSm37m3KCI4/4cS5V/FmtyORHfen1ITk6WrYQDg
QEnLWyl0SjUySZiIkryF47Ux+wcFqExdFkI06TUQykd9gnUZHLQOzGNwfDZje1Jf25H6Y0xi9o04
Z+cUe32aUYKZl5EXQkVnTkCjRLm+QeWiyL1wcHnSFGwgqHFTrBO3Wao/h997G7vazNvorCkAScxp
MdRy7FRBxkdl6a/LWT2u3F5X8ql3vF/HqaTzFQNY0skzRDyWbf2yu0YpflQAxXmhpewxy6x8KQwd
h4Ympz0ZP/Bt8FF96ekSTJamCmAu+HiAUtDHcUjKI+gpLq4vL3fJar5jHSTlRJitUiiUDkRxXaEX
loKuWAOniHkZmjW4a9iE6Qev+HCys2EkLs3vldf7+R41qpLjqw9aZgeN1fjtLkKtRNGu1fHTdBNJ
HVGjwopKIb3swiq5KJHm9keaOX2MFuBCGD6APcAMCSf9/RYyBWsN8RYs6SChyVkxxF6yNftWlFuG
bU8J/eN0Zi239wJL46yc9pjg2D7hnOITcIjG2tPHuVuDuFqcpU9Liw8Fd/xe+0Q37Zw2gJ5sgIFr
zKRT/fKmd/tk7uDo1Wuy9nwRGUsk0xZsLzsl46mUPcmA6MDOS1dqj2Woq1AvjMR0QYB124VTUz49
PIctyOn9IF5tEnAxHp8ASdddugR5gUkCoWyWr2w5zAVn7XE36FaDNfq77BPq64t6YKZRo4tGwumD
yDpiWAR19Jc5Sbuvg6N8LF92ZZO2DyJFlp5x0PiNaH4gQSYVA47MB5BEo693F0npZTWbTaN1qzq9
4Q3zC2tYZa9nqVckhmneKrjMB8ZSHL7RKya56tPEAbf+hqx+2TJbBaqPGZlEu5LTtmYufmSZiDq2
mnN9sokLA+iR5LQCnk9uGtWleTbh7YKZtP58E/u2u0x8cnk2h2TwQhmTPEEiQN6hbgZHzQOiBsSV
uBAuR2AqfyOFvNFSdyjAFKkJLlSXPr9PxpMJM9H6bAZ5xQhhAmkERQN9fGb7S6g69Jr2fQ9wVNh0
r9Ekj5LbiCMFknHDqxteo4pxrS9Ug0W3IOgjd+jneRrUz+YbBNzhQws2TSL62KtJdN3Y7QkN/pku
C3/L1hA6J7/ay28M0hXsf3WM7HKwekMOhAyJHWTzcayo3/fI/627/DyABq3bYChzDlQ8UkVlDNBr
1AMKLJvLHmj3asAhlKSAaULBYgp5AW0rzZf/2gdEL8kObOWH4wpi9YE/vk7J+M4gX1969/1I6i1u
nswZLuvLXWJROySIon6R5vhRCnL2TWrLJX2rCt+DaFLuy2iUzD6gv7HGmRqbxfcIJf+4rozfD0ch
MiqxpT1rtxmiP0sfQ11n0GCgVJ+J+QsKFItJsDQgTSyCDfG2ZrwLYhOPSL7i6mtkVEBWiWk6dCvI
2dwkWOge+ziRaWEJRIXPf7WVqM+Hec+TQ7ptzw49zrSF5d9PTS4IULP9OIjNP+T+FEfw4beD2Fxe
xw7srCYWvbNtPSag9FPYZZXY6uCxA96Ih6xO327EJgjLbekOl1pT5t6dBlU4i0Mvp0YuBQg5X3Rk
/NoqFlZhhjcQfx6r4DuqWhdA6q2q/yvJkHrRJ4QOIqeQDG+7fjuflyeUjsGhRQzqQxdapmPLOgwl
zYbOg73TTfxf5a9l9ancM5f+crtu6R8pWbDYTlBGWWd2R+maj1gdnPBy156rtkLI+49yTNOhKA/j
uxJWYwarrSEXr0+o1rH+wEpGVin3/qqWHky8xonsKjcFHx0N5IeZpSiFlYNh6LdP1DJ6MiBbSPMX
5p6LrjERmV+FeO0XnbAsVZQSjK9wyc/LYgCqR8nu831GXPx4iIpK2FuljtAxX9eFKQK2eXXGAtBR
frq+F6yZ7M5jdXKBDJeja03++6XAOP/oos7+PIcgpvxvKYiuqkfo+dKPYOrHsXzne1+j4EC451Gh
dhfqS6YW15h6iIiV+o3v5Ej+4ZcUO5HAF0NubfaORnFaZ/CIeIAcDmFHE45YA+fd+VhK5p7eMCsY
K5ZxqiF4gg1m1Ab7OMuQtnvlTHw2va4N7Lr5lWziFor0lRK5/N854jBLXZjZjgLwPM9L7TRNGCCw
8Jwr6n45i0qCa7VPXSavUsksZ7tyUEvT/tLOeKi+uXWFGOzvHzhPy6xWxzTZLqWh25xcRUWX/NNl
kcxNndSbSsLiNeMXyi5egoaGr7XGAIXeUy0d/e7XeiR6yLghO15L3A1+vH3MjPIwqvesMUjGBoca
z+pNHErP3/IV6JM2Kx0pV8OYrN6Cuuv/1hrp0HD4rnNODkLeK0YAOXMll/FCDlflPpdX3hYRPCWK
h7bhSZNrt7YW3oHJff6C9RI74OL/rwLKZt398pM0ngVKc1PuozAdDCDJB1veHHuZys+ge0UkBTsJ
iixJzkh9cLj3JPy5FJ29HCW87qrczAxSm+sjM7h/VTEqY7qf9xeHxcYrteT/C3SMT7WrGUYcHBcj
an2ogx9nz9hunyTLZo9ZdhCXjX9zmbAQpxwQ0ANALMuehlxlbSxWxE+P7S55lvLyBkowCd5wR1I0
xt3OTFAYUf+sjSDVk78MMVgrMycN0FmencY/CMPYEFSeqOloekB4OJpCmBvPdeC20U2Qrgqxj0X5
rXLsi6mZxnCmR8JHpimVbKAxkPDW3pAYkxsuDOCe1vSKl1tIqOLVcMN8OwQVBJUjap8R7pIF5gQ1
gpdIabBKjkw1Ki0GI3y+9NIQZivop9DBl8S1Nmkyk3M9ANh4sY+tDv4a4RDEhYl6iUK/LJHPKAg0
SWydlx8qLdiIYoISe9pUJq9OKf+0oArzwSPoDxfcKvL/qAfrDqQEUGBrKnfIvZvuKfb6Kj5d1zNR
OvyOwmqP9w+ISd++Rx486su7JV1C3StKaMCBEqCAu/V9WjG4aZuHjdHA2NHiAfoqODXGbUrOgsZy
m9ctca7UIOzQnKCN0j3xLMmbVJlcIJH531wUPvFODZqdAlngqPu2YNXxyxo3rC5y0yBAqt6HzkqE
aHI+6eKr3xIJJXCOQs7BGGn5PIPLkDpgZCc6SrFqqdf0TdOnVFqwjLxjVrBNsOBzwYqXu/G/XrIZ
Cj/r2hZleU8+zPRbsYX8c/8qDHZ3ZLgUDHlvvfi3n5FXLKjU+qUwe8LbevX4RfL67b6q+QosHrTy
sJHzjEstu3cOxttm0yUtWJJ6gubYGKIlf49QqBIAroeT9j7pUiwP1EdSM682iUQw9Ha2YPkpUbrn
XdxRy+9IQuFJFzZpD4fPnGiTNukXv0Gd5VF/o3I/TmxMcWozM+W3FPtGPlTU8J3W9VwNHWg1lOI6
mOZCCVC8d5R6hzlnMHzN9FW9DckaQSR2mqEiH0BEpfdpRNgljfhoA9G6edqEypt+EhqoiROFwYHm
FghRocIxkcr/jclhAN0AtegfwzXwpbud7N4mIMk7I50eUAE/WEkrpAuYXsM6BZ4PS5S9XrgEGQx1
GH0g7KeJgf31p9o4xr9T4a8oV8Qk6gmJ6zJ0BBy0JPJOUjSn5m5xjs5qLeWgT+EbOXOSA5/CVRk2
E2/99ZSNDCGNhdvTJcXTdg60q93bIwdsEXlueQLwKBtZ4yWXEwUc9YCJ3xkqm04Rqaha/EXRGbee
m3/o9PkgX1hv2lCs7H+DaxyQQ0W7it+CTRvH8OX9k23xnXocoSE3ie75Bk6wRLntx4vasbJbNWRe
DEWtA6KvY9LhNtZ2Kc265czi1dMoK/w5ASKQ4bvhJJDTyXMgo8FA+HTZc5UkEBJW1qpbM04S25ql
dJ0I5XEknNpRFiFvxPSr5f9DCglIcQN8y/wzT2I5XsLn6gkT4cTxLD1y8E7lkdvSNpdyVKkt+7NW
aJ50qf/iCn12ZNrNC5y0qtgXU744XdR4O9Nal/sAM6RUNNiwX5NIca2uT3agvQegDlQL5Ll9DWcy
ACXPC24EISjPjwBC4bQ9MeKrMCiRGGcEB9UtICEyjBt4WSpOWYS+L221xSyoP8tuXZ9wl3vq+6IY
jKCy5NsXEf8fB/4xcWEyXoTCBawS7W8E9/w+HzYdeXRVMejV05OGEwA0PAknaGtT1aifnF5axjUJ
yrW+RGPtq/JKwdmqbniwOlUOyrWlqpckizG5lZtXbtA+fEdV6t5i9zNsWm36bsL3NpNan4KbjaTB
K+u9rt5Nh2MWJ6vEg1isI3YHMusMj5e1EQy+LU/Am8LGdX/tZKfbKKN4a1elXJ4fglwq49f8GbrQ
SRMf8sMjCqSM8kB3ko6ccIjIjPbTy5J/5sFn1rFDLBu2Fp0TNq7Ceb4JUcKk1FesXPTaCgq9tCd+
1iJj85RL5romVZb/K39jKKFwdvThRo8Kgc23nEaM24AAvZZr5Zt0vNolQsopcFwasWlD55lZBMqN
NJnpGFAELciwzTU9wVQeYAe4XtdtkmtwhRs965rI67jZB6oH/Iy4fxHmmHjgsGQj/gcbxTHgouIZ
BT4vKdRAkyJa8U7o7EyYCuThulfbiFS5e4P/0V39+XFTlJEE5b25CcN3WPXLWzlLyvB8cE9lzau/
k8UcwMvCLbDHw2cgy0Dpr8Rh6wLxQGz8lxG2LaMes5FZ7o0DpsFktlCMya+8X94IUjWXYA4gVId1
xx52qeHUXCKcFWLpkBOb1ZRjomxtMuWZSwRgDQaDFAiqbqI8JRVEXJNPMCb2Mzyw+AfT0s4+y7D+
zs3gmjI/1UD43+VprZzSv93z3XVT7MTQQO1k7/fLZn7UR6eHCkzvCWEe8TQcx6AueUow2rzqXexN
jrpdVtWkezPOEyXYLEQZ9eWAkyDXUiiNWxLt7Fsl63yxjoGTTOi4ttUFK/5R11dTlgcqldPGPsL/
3Tt+dl7VztLJ4iAdvCx7asCoCYt7P/XV2kIdhr5HNhFn+JR877nmH1Zf2Chgpn6BhBZ01aGzKf7B
6e2gqZS22UZTSSNEyo3C+ajldYttdxojePp31tYp3pn0MbRFEIJKbFM6iJSQzT4ALltWkyJCYdWU
JFd7UuwWbNzvLXm2rIgABTDF/nbBJmVXa8rUA7l4apu+gLBqswGOp0tAgwmq8jCpIZBxDwLeyNXi
+sMHmWJzrYBxLh6VHgnJjk8RylVwwG3v2sK9T6/n/dNKi1DvAXoirIyQcHVEuhP2tnzbjvyFJOkG
ces6xF56E4qWTEsneVMEcKN8o41ChJC34OTUFpy6ZBq1zOkipCATpzDIuBbwBroxgXyb7aDKmDts
Kz14f2b+Yumxg/qzg1lG/HlbeDdlDpUCaBqKKY+Zlxry2fR6cwVxuOjAWfkgLtebs/X+5T1WBOlJ
sr9B5SKvO9eB4pdhAWGKh6FfZeiqUs15eNu7qXzy5cK9JLRox+N6jHjBdURFzEL4Pz9KeGsEvOVM
hmfKxXTRfYnEcQWbBKRgOwq9QLJ4nD80Z3ONCcUwL/Cev7wnc5RFS20oVaCAqDesnLCJQmEozdJ7
skRUlPQlnzcOWW3+8vbdwf0TGjlUeqcIjiI9IttlnA/Lv/eNjTZyLFLCUhou3qTtDp21SWlDcXZV
19rTPES+Aoe92VITbujlOc3k/EPX6LAAk0JDNYFvDz4gV6G0qE5Vdv1mIhxdKL0xkUKc9nUQjvai
4pM4/1eYhKmrT3xyKYtNHwzWD9L107+/nBfWYRgiwUfYO0MXUBQFppxm8PZ8I41sp2vYbW5RrfRG
D3E24H9FI+F9juQe1U5/396q4FC9fRtFDpvQk1JdpBHfLH3LOFOG/UozGrjBHa3jndK+RBS0lulh
cSw7eqbEtsx/wyBrPlwx3yxsoI5dDIhIAS8kHQUh4HXMHZxtZ0G6Hz/eKCMNBgp0rxPLwyJCuJi3
rVvb2+ZOGM5I8FcKfk2Es38wfOwObmHbKevayO15LflBTPjljafSyqE6hA95XLw2terESOvDMwLO
Pu7V8jEVdY5TVxTH0A+WFVi0Zh+FMdt6NeLH1k+Ujh39QYbrcsKiTA4p37y85lpZqRPM0XSN5nIE
MKiVkhVIbL5ohMZjJ/B04+at9vzAQi2QzwaaTOWNT53KD9dIwJSgPfxfQV4hMStGsSEXg8pfZoni
NJG6EDyOCFP37RZn08WzE9CJUL/HllUt+vo8YSBd5LeJnuNj0eQ2haldICzW2LeiIlCr85/jcByc
2Y9WdZQAXlpGpgwQ/S3DGHLFTWSK41BFL7LvkJ7A0Qxizeww+DXQPQDMJEvNKruCme9L1Pza1oWY
ouwWcw1SvzOeS+RI9EOk8Lchi1/Z9M8lbjfX5NAn8xuhmPQIuo3f/r/JsEnqPRDArvngwy+/mUEk
49l/9IVnHIYdThRD/4WbpHzPZod7ATK5OSrwEF1UPU/tFGKjKQoMi19PBlkSADgISqiRE0pS8TQ+
V7i1ViCI1cL6zkyWjetCO5VJNpWNF6LKNHqSpjKAAn4VW2Oa2pLR+EMv2dB/wcMCLSgs9cZgyVuN
B2hNju8vGlQL2LnMmEEmt6IDT1Js4HDo/JWhBCz6xTjzdZFktCljAOSmZkrX5YzFqVf/rk/fPAkK
s4cfil2OpB6rRKCUqbUjOLwkEnw2u+6bhcLJAayZkqiaTHsJq43UYTfBiH0CC4/4Ztl/hdc8iLyU
168Gxmc6I3AHlXWHtBhaJGNsPkmxm6Wrp16Vp8DQqVVImo7jrStOWu8jcdSE9Hih7B97Rz/1+o5G
xjsyLE+LU3P6DFtEuKN08K8EZlCGHrBYYzrzY0zBJFe1k2eKtoabdmQ/aZynuKqcZfjWNBwx27uY
rDVcTpB8misgTIxtVgXBbNqOnI1GVCdD3MDQ5frmt/H6MD/v/yn3753O47zwE4WralJTapDSlewL
eCWKutjNoj1tbs0eEc5AiaZSZA2/TFpG6D6OM3tOhoLHpHRUE886plmHIxgyrztGc3HivSE5974V
oo9y7HcI842K79RPwQdG+19s4gYmRXEWE/MO2YPYwqsvDAYHYVGK9Yv3NqXj3XBa5nC/RVOeG3zS
dA3t9dU/MvnyYoO6A5ko/VWGP75NPsaknuLqw+Gn+SV/aCSH8yFZWIPphQ5dTd8Fskw0Eo3cip2+
CUJMAnYo6FJHlaHnFGMcdN8sQYwNU1uonbjVha3CW8scL8OGgMH675CKKd3YzB8aqfVmwUsw8VQq
WDCPrwKCSeHlbAGKymyf8ln4+llckS2hSYUFMGSRdcdK6D+CvSTe30meLSK47Rv5U90p1y1T1Fyu
5YvecrHvtQqF4CCyo4n9cGeri2OZX69xQVEjOZ+c99PxZq+acHEnhlPbNbaqzXxrMY5mAcjPxurk
64Opmu/h14WUuAkj5Jk25LI2+H2IxUNJlPOy49WAYsBc4UpGSg7L0Q70Ho3XiqTBBEwl4/z/R+3y
7fdxumoCuvMfnLP/F4/sf9zkQqiWTbm24kDyV2t/u3Q2soBxAlSqzLngwVN6GSj8jmwQmDkOr+ue
0a7x3R1n6scfULocELNbu8ToQoUePvuu16+A7kXY5oaphc0/iBnLaJrgnHbQkvS+hOwVbVOI8iP1
mUQsHANppXZVWOvCoy/5ud+HQglF1+RYh7ZxR8IsmC4hJDTTnBZ/6ncYEff55WOyowWuXHDN/1fB
Ee8CDcfMHMHJ1Hl96BkzSpR7Ha/flC0IZLJe8mU565BJfzRAEN0dNbAfaU0eYL5kHFGmknaiWgrA
7L6XPtEBCWOR1tZ4gwFaEnpm9ngO7hVTlYLsGfD7nPsGyrC+N/N8I2V1tPCE0kL6YhRBg7HL2/45
ow5lH12y0XzAB2n1scFkJANLB/sObUqWsRmXJRuEW8ywHgWrWQSliYrSlNSa6vcJdWnGPQXxKdIf
liHnIhytlI9uNIJcZpjIKO/z/RmNsN7TfbQJk8kLnqLbAStjZDVLabREe1KQn9CBV6W8PtnyIlY8
2W/RRF2iqh072jBITvxce5gvhtC9393m3MNdfA1O3tAl3NKYUKaja0MO4jWKTYk8Wct4+u9s30o6
kECE+nu6Nk/j603p+RFAynm7jRdvCWRRgc5c75DjvYGGczJK+ZQD+F5OyxHxRInTvCAmZFYLIpwa
bskkbLsCbjAO3jfef5h3NsCzAFxhFRFyN3C3mmwuP6z95lxmfVHvDRO70/biTv96cY4h3YwCVJIk
qE5X8xGiYsmh9zMQy9pGwHRdqFaoYxQ7JQ2nIxhOn/sXBsZj+k0w/OdcfcfjDmwYfhAN7w04dYFn
j6b4OoFVsejqhHuw8C5p/9czj+dfEKCtekUm2mBLn4nb0J4ofxzbZrB6Arat+7HRzBDNJeTDlzhy
iAt7G7l5wGzy/GYcTsYdH10upq3F9tlUA337+WbtmYYVQuI4hm6CTDWVtPftb7QIo9vFlZYe7a1+
iHJAjjfPAtH6PdvtIDVWnPHPZhbX9wzJy0LREMRdm7aDO22wX5zzdoO+36b4KP7OELnFanzfYscs
dvvOvHrw+v5ebC7Y4+zXPxi/R/reyrYvbL7NTWxE06PDoybO7yVRhgqkG/UnUDwLgDdeWABLPuHb
Ngo93MkNgnK+vD5IZ+BOqGSnbg0YYaAYU8Ka4oGv3As58d3iPOYmNfA4K4HkrKvr+X4m/9FyVqhd
xndZajTSujUp+ay2KpsmNoPrsHaX8YQRDlunegbuqJij8buEIGqy/vYks1AFQyCQSJlAVgKYQgkz
phH56aNFE/KyUcG26ZCLYzKjCbxQ0R9XAqgRRNku1PbAkRwxt6JxIEUvSEI0hcXxeUQjgGISBDrT
E8jMYiVrPoQZjSDIqDISVktMX+I/jfm1aLKKFN5psi+vT9nusUr44dzh30ARiIR1CTsNeKdbwdKA
YipKFYVUDSDBGNogjTZORfMkDrZ2ACuW3oyOxURlbx0cBMl8UNOSy3X+L7X9N11AbifeQtJ6GMZp
iRpBk4inG4/dtuUWWWRdSKanU+A2/g26tckv+7OZ6ZygIcCDbREhSEa29MsTTmz51p25wLXwbBJ1
+uAvRzhawakg5UCn995rBX/QL67vqjFJ8mXhEUXNIblf+uGwtqYxzzoXYjnronekXX/NiUgG/Ajv
B4AnS4sL5XT37SsuxzGrtMFXahRVhuZrgKjdJHoumFpu48GgFaPM90TG7YOauz3ubRs69zF52EMO
dPR8keFet3lOFjZpBpPdUPIaAUeS9SDZETbsUnXOOlnLrmJ8L+DPoWwypGk17aocVChrcokU2MUP
kcaOJH/+kDn8xgdVKGXaMaLb7hKY0i/0BJHYR7A6QZW8qDmCyqUGj4prFTgPcCASKeN2eStGCGVg
kgxsJYHAtpzAzA5aolt6t8S1O5698ot8g6xmd5JNW+9A5YyJuYoYH6dfpaFZrACpyk4rEIT3ANrC
Uc0NtvS8J+YHxPVTraNeFAAuddguAmtdJpZzxZmOMObc8WoM5x5tqOGdM0q7mq9wjzsI15TJyNDG
oT9G+y8XdWfi62do/w3zv7tjV7AugzW6NUErsvID6y8hoAwl31sa1ppZ48YfxjAmcFy+JP2ElCgM
S0BWzAi9+6I9vvrbT9tKkYflJAEiWMCX7JLKfWeueJ90C0+nGfQcriGcFDNZcVSpvGkOix6BMfHG
mnW21/vG7e1r3RWnRgCmSybC91Lz5zjPe5Fn1dGroBSALC6OtVvLjpGSBVAVKeoPoommBHSpmSqd
pEcIefuE5vybJa8RR2VyzQAxANu4Ub9Tx+iL9aW33lxs9np2Qzc2joGezELdWZz3U5bNvfGMNg9z
4fC7Z+u7bY4SOQTb1cQMTRipk8OIzz5Wg5pZk1cTZycM1qrOHyyPsCtAVVC8UZPm8D0NEbRaLT45
/wWfCkeBOinfXxKO/Y70ve+JnJ8cYnaKzC7SR1mXK8SI1htopEw7nbxPBucrxx9D3H9TRTySD41j
j2yN+F6Ry9+mDAeuXB/NK+zo4f8lf0KAIknQ2QnnwanUsQKx7DILBoxkZZUaBSzOyA658hSAm4um
E24rB40ReFa6Gman2J1Usa4BhmCfR/kcRqRKGhL0l7TyEpPUkxMFp1bJ3QGNZXglvMq6aAUSa8EX
q21ht6168EjgI1z/479IiPfdAYeELfELNmrTqPRa5wXL4saKp1GVHCL3qZHqVUF2Vhoyw8tYyDbC
QCuNzFkx9qMn5/O5KGKz7nisdYEs5EmZDnuyNwyohNk0/ws0RZ7nUBlrkwbt6RgTjakGuXqX+dly
FnVp6VplYa3YR23+8f8Zqmsu8iR41ApyW4UJ/4EGlBgIokR0SpHumfy9UnrAG3vF2KeF1u00XVNt
Vnk80u1jeM8rFi4FS/OJNfgVonhWUKX7ZmMq6qZEl8+156MJVXHjJS4cfuxGRfili6TcVsqUB3qp
V0qUYTExKbPpBauvqSr8H2dYUcjMwSEWJHdZgU8oUuF68qhDxRxlFcPNXGOOi4ITGJPlZxNjadT5
aXAtqkATTPsGnmjSu2bAbvK+QmmaVTu3tb15ndWQUQvsHVcdH5LCerF6eboqX5/i2d0R9SlG7WYD
EkxxfijEOCNeZlvJPfFOh66BQkXuDYBg3FgRCh3+MvCzH2i0oFhf7o3EiGJNYRLmOT9Xt5pxD+/t
FzbkxWeyuUQXO4NMaDu5LqXu1r1oZCYnJ+g0pQh1vOFeOlFqvHiNY/hfSB7Qpxy55i0BcDK7Q4p7
loyn9SEHTuaTb6XXaJWfmrWT+57kEpwb5PzCtB1lB47fKd4xCLpwZrHP9HObFsad307b0IzZ+8zw
7qgEdnKiiH+zMkBVMUl4X/YOHOwmboOvZzty7H9ycwYz8jcYQr8bCPovm5G68g10tM598VuXFA9Y
Bj1OhcsE3WPAn1oBqThV+ibkrujdLnvH2IRaB/F4HR+Sln9+/2dosN/05kLttc3I1Sn1kRXfVKZu
LNA2VeuHuKg9hH8gI3eeN+RhoFstcQXyxBClNxmbVXk+Us2dckJQ7eH33UzaceFKOQZpLezmDoKd
5A7GyxUryp83WUo/m3c6lOBd3/pk/aWI+CVZQ4a5E+uA9iAlAbi24qzUfNgTnyfb6FTI7d5LxWxT
vnTy7zb0EM1+yjBjqGOIw4tj2f3nkX0RxnS0Lp3unNWQQyhtvr7qpNRyb/SCo04OdERApG0uHL8N
gLJecyYtxi7ic1CEhx4vHGSf4T1M59VeLSunrXPFzcVKVD7sUTiKAUBNQK1GodLChdFdmGlHdi4X
Qir88phediwNa8AKWXAhfQYlSai9Z/19f8pSiAKeJXXNcgsD413CP44pvhY0ulAn3pTuJQfoh5se
AUk2asYYFw7LtJzJJrt/ojtem9uMSTQG5KHscba6gcVlRZ34ORrLHpoIr7q+VpfRlQXMdCCQdPVB
S7q7kZgIX9RCOCkWFw7i822Uo/bSHV2aZp58gnbzgWIWc6xTfnApXuriSR5htxxINUbc+Yzj8Arx
0a7eDG6KwpzO0E3sxWNRoMTJd6QH5Hy1XvPccUshcZwc9MBZYLEm9EuLIbwdhb1Uxrukh4UF9lm7
3D5SG50p86ABz4y/mFLuxvs4oSEdTzLTtWLpGuuSIG6FaQTmdJIHXeCQ//L19YNRIqU7UVRBJPIB
5HDNFpdmPPQa1IUVqmkYPZPTjFNUKBOk6ekJbkHqEjUf3RKyH2mDkSZoBI7DTFGKzUWNo3/p4abe
zgHBsjguzodPdB9n4z3BjV8gY3b8RRYXpPHREYAo1cwpvwO29fonEoccyBsm9p4hsAnsqDNOLHdU
gZVT12ofaoXBAIVPlPBxENoOTTBTxHy21/t7bFQFXEvYFlnJiEMyGmmf5/PqosV/VCdB6BgWO+OB
S77N9ll4KWB6WvtvTd8PUxRZJ6wLM9qTVlxbvPAOkQssIzMhv0Hde87GQJPGtdng3L4QMKveMBv7
AOL8clAICNfPWrmWXp4WitkMQpI7ox9TfoURhFNrGItwrYY4LIgiMY+1JQ1Y9yo/CyWEn93EMrgt
tPPKUUd5NVa8hvPORkxjPNY1T6+wLKCk27o5xPseJbm1M0q3hQhHBSA558gdWIUzmNfp7opM3RW7
WbAsESSTS1a4aZxt3rPVLEaROLcIpvjl6oVOO2ZcZB9XsMvncRiwf9BGSuZ5H4qSVL24Pe5VLC7v
dlpnh+VZUa3vaJmRzxK8rIn9hc6DFKrpJcZTmpkHa6X3VUwEwmNen1R/xqWYYyV5UygYez8yzQ4I
qz7s97CwGO1xqXwHrVTuf5ZxV1sK3Bqgr0yxi5C6tbJh3ir2z0im+wxmAZbxNlU52S0qfP/uB9Nc
13TYW78VbzORFAgvUztU4oq0adUG3J/KPbeDKfix1mPgDnKShOZtoBofVq1ZqouzDp+8U0pj5sSV
FaqIRDNMOx/5HNQu8EiK3joQVC2J1qNv2KoBhBtOkNXWcHlFRDA7DM9CljjPg9xHCjWDgnFbhnGQ
wgI2Z+98SLIKaQcZ+rw8CK3I6+VsDaDyKC5nfbLRudOMMEP5/+CpR91K2TDui3InbH784CH7StBR
3pT5eFIp6fPmJZ/qBbJAPQ6xevjhe+swzIqtdX9f4U8FACtUBjyjIpzslgL+wl7KH0/ODccdTIPQ
JlT35seh4WxRmeA5OKtcXNiQOVJE6XxGIbNxiSa9lzMrCK6GNTeE6HfhZh5YuzpmxJd7kvTQVhd5
ND9+1q+0n+ID2p5JoY4Yg4fZdi2JBBoGMQw9zshQvFqmw1KTb216ga/p9TN4SOGv2iDBabkFpM1S
/C6Ci6yccncaTb/OvlRJcy7JBxeEF2kf7UemMKe0Ek/ZkfDKwsExOg8quEyTWwciiJAtIUpKR2xD
ktoN9pXCvTpeIiX4pJMXkDdaQiEiF5L/84uSRKwolyRQRAO/XePVq+eLR/RuRNOuKS/iRpIo90P9
9fo6jVd0d6A9igdfrbSYTKe7HEWcGfDm1wtxeyw1Q5NNZJxellSZM4bdW6iYu7aENnHcRxOPABpu
o8OqITSW0wKkCniXl5+nSRuzyLCGNGleh6u7ZoKMGneoDVgzKL2Quj2123tBwnAOjA8g+8vymxy8
JsbqMGp2pOn7Je5WN0juWyvkKNrEZRLOqOxhsvOAlJyYwSeEoVDtV68un4FTGfnLlamsKCP+QSKX
z2RXtayqWyFJk8YsgUZBpfuPEx4qV5/MaJLF+CxOPl3ShFA0sBALSNYSx6p3vHLdhfywZopolm6+
+wtno8YI+mhSJ1qDlgZtzSFDgluUQpp2qvTlgzHBA3g4mX66xwPEr60HVZqYukCl1IM8yxHTC1kw
h3CXQYp1A6tp0kOF2nguLBMAxKhjjfvQBUw42YpE+2HQ1kIllWlwQPeTIwA9U336xzv8ZFTMgFJS
Ob0OeD2qHWQa/wFzDAuGtfvv1Rex5Zn6KWULD0H5mkRVWXuo8dqtmdYIH0kEtuUVjQOpAtWVQL7X
3J1Gnq+S3xA1SD4EiWzy5OH2BnKXzubSMpMKY41kd1pG2cOMODFyJLm38ZIBV8ABzAfqQiac6ikj
V5fdS9nwL5a9S/SU+hmgNF4ARXTDHmrQ8/D4s0wHTD9DQYyWmi/A/84eZ7lwwqt4X9AnwRn2BDtH
B6nlRIHb6/+MSYwvkuMqcpysLeXQdotloztlDr2bbt+hEI9SRibXXg4NVnpPEPjNSQetwpghlU/3
wcJFharDNfBB6BaJHxBoyomXEOziKgtFyvCg+7z5Pum1+tBsqbhhBlXw0y19e5zsptrMzt8gsFx2
RjDDq4gtrpXB9bQO7yrX32ccIkAlCN+A6nQKGmNRjfhVqMHlsQ1e1TLr78rKWXdHPOioMSReb54W
QhRtGGfy+ikuargBlqtVF//4FU7hk3+/ktcF3FL9x/4/+lGkL/Ez++EwiAO6L3hEcWrtPgJgT3cb
TeTGj88vk1pqBFE2OHBYqERpzlnbFsF65RYF21Fg1TaUpEibAmp0eeFlIOnurTu8zpLnwoIMzanT
XqM49SPBlumlrkRMlVOL85lQsXO5JVnCxuVXcF63jADGQkiuB3vKHVqdAzbAINn0KCgrJboAoVJO
SVIwOViscJXwisICmLNHXC1tT7rbgnqh1KBk1yHkRccm6MccnOyNY8h1Rca1v2demDczHUcyRDt8
+/9sPumzK9vrq6LLaEdRocKDeT/QlVX5rTB4WCtXUkmrYIVMnRTXHGi58DipaPsGaMKIJZAnGVec
NKL2XkPDqeF00EZUqbrNdNJGzPCdltZcLQNsZdu6dtody/kQjkCKzyluk+cyjnVJzhXSUz0jIedb
Bdh8A4VweJUk6k6mh+sJzHbTWDY3AYghZdgSRaGESalXn+7hfVRboBZHktF/SD05f3u0gTK3Hni+
nYU8pFLWN1cWMQvLpHIaPgGM2zlBoS3S6bTjvmzny7kJZkZnbC14+OTthm+TTN1zgCauiz+Wn3o6
SfblXhcIOa5MGapoWaOC1PQ5MHKvE51ombaqay+2oHgBn+BPCAcvVfso+Qe/Dyaqls/VoGnWJ5MV
wqv2Jln3ftiBFWEMRP+YSZdyqWB+x4iLGiO2Hxr02ButROUxAHVDkV8g6TsYSXEzIhgjRJ1TW76Y
vwvYS7gUbBRlK8+HhWeFNM2xPTXMz9jChCo4wNpUlG6YUMrZXUZ1GgKQucDajvTBjluYK0O+Az/U
6AWzhF8ZLAf6T46Rui0tHOYR9axqlq04ncM42ptUMllQ4vzYQ7AVW9AA8W+J+e7TBO9AdVKiQ/IE
88tK8tan50z059CauV4qZVG8RdJ6+lQXe+6J5+3FioUOieBeUMFBmMfP5bF25BcU190l/QV6GVEz
9MuEQz+0Cccu5LkBPO4AbYr5K6QWe3jrvZ4geLJsi5icIDz6c8OBW0ubv2ebdUNwtOB5MOdMBwh2
uudt4pKG4Q42Jn8SLdG/QiY+DK/Cmlkyi1hjr3fV2CfXkKuT5VxTQ9wG/kFvN/5M4gF4nax1rVhI
3Vn79ZnPPb8sPyCcAgfzQEBrA/K2ayGIvR/cPFrjUF+JzRrqK/K9UtnmL/dmRKjVMo0EsoNxBmrF
4QgQl3prsra4dTCGnV9kbAwHsv4ZtHfwZSqOrUMJWfKo+sRbBjS5tsxWKuu8w4ASHifD2dVIGYh3
z4ip08ziiPZnVOA89HBBinoGIuIoluZBpv0+KAe8TOX/ft4ba3N4zKp4aTng767lQr5G3U7Rh1G4
Z3ww7XPrRICbk8EoeZHef0CO/jWJOF0n6uogWnrxLQYQu6/f1Z5ewA69wygv4A97XlVAfVtBn6DZ
9bWCXB9Whe6lOb3jfNHHsAN28HI26X1JMCQb3TqgS7S+ih3I86v703zmwF4H/R1NeQhVqt9wL5Mt
mchiA/FXgjxwgmiKpfApTEyMALER3L/6rEmBFwM40Rp6eI3/vk94wdYoC4ZEMwhkM3BRfR3imudf
ZJjGFvelGigEXj58DXLf3gVa46itEZ1SeK6zlX197CLxR3dbOnVL4HqxpdhomGbAfRq0d5bHQWUm
mZVBan5Vmo4md8t1R8zmAHR6DWeJanX0zbiLw13uMM3ViCkDSIYRQrp1h8un+WhiHCQoQY5kSHMt
3qbq5IP1bLZ3C3O/TASOteaT1u29uTvwP7YXZ/nqhVeekwwF4vatq7ynu4e24BuUfj05BNGVh9Ze
IGokVER7eQyfdw9gHQXcAQBYIB1ZLwWCehRHDU3xkM6j5bf1QUWF2JZ7X4sx5TK29g0LxiHHA11Q
SuTZm7e6MrPS9vZLBgrw8ETD8Ii+Mlttdhi1gfFiehrr1KAH5+1EGOyWn3CSo04I9vBcM88aYMBj
IKmlh6qHlpDyqsSQaDno2/vWbzZfGL3Iftdfhm0bJfYHK8jOvRDdd37wvkcGG7Cs9yqcZ5Kof02w
Af4XuiylSRy9DlAG5ZbHSjOqdXEqRnsYAoVBlczBQdyaGQpGqa6rkWb0QhlYhPzwv2fYeQlp2DaZ
sFjqk/XziNVu20TFh//FQRG6ugUYGtYNyqJmHc5pm4vdguzTqhortZan0DaMwNVZaPQp1NrM8r/w
eR41Mt7xtxWs6zKR4dpdT/NvLZwEedpzLTFTb3ZaHHo4GkQWQ4P+2Aqr/4kLQlv4s00gTLPf0Deu
s+TyNwnuqE16Mql/mhR1xJzgbgHD9FLpS+ss6mMa6u8EK0jmX5rJE3piFAoSglyjNb1ORvX1JjUi
6nAigoey89bLdVwTrtpK4FIHlYTNx7TulOj8P2zgO+q3cMAGRKNZvANouj7aWoAlB5f/hlQst81j
E3M4myPKYnSxMXImZtL6aMWYPtGUR5PNb9By2ky+F4Gsu/jN5ya0elPYotR2QZqP7iiMd1vaTuHo
7BsyKp6PZEi2tjadH/sfLHEykGlObjqtKCPCUQv5NmsP8Mppdu5zFXGHx77xYklxE2jXq6VxFICD
TlmD23EC6SZwFvKueXWnWTdXiSaHSOi9LVb3WTY1lCLQ2mKsu/jHaf5oFLK+JCaF/v5hBSWUVBJa
gtD7TFOgmXqhm0INklEYNVx6hvW9h2iTPqT6d4vAiY+a0DcKTuBUyFcLv58N7Z0Pdk5TaX+LUykS
t/HvdcKoAjAxpUkEJUeIX56ZyqU0juWzGgb+V1q1g7juJvhsWDBL71zroM9cLxufuarfQJbb/w3R
igFuQFRJPi2S8BKhmPc8z9ftYAejw7tz/YlGkXCUgOgIXPZMut7BZJVt3sH/XrA2cYJqoXxr37i7
efZ26iosxB4T7LrXkpb4yKDbixoGnZdz39N7hMeV/S2+sIEs/ITtTAV0Qyhf1Is6JxOBw/BOyeqD
/slx5p4jaidxCv70xkNKvwtf+lowquQawsB9/XlVUU+42m1UArRG2cUKdP/NuCZbSNY3O6panm1w
xVl6hl/tPd6PaScIbwYD+sRGTbuLhB/ToDpV2vEzJR+p899z4VGKfssZuqUba/dI3ztk0+otZNkt
2ONK9MnwBbTLvPHw2TtMpQnnO2QJNgPIJenSc8XcWePPHiS5UEpWN9jI4dn0OZg3JSfBOuvMpKEu
Odo9s8GseEgh3rolnkt/YgaVitlCiS4kPjAzjtbWU3/P+7NwjIbli3VOgpSdjwGZsEXE8taf51TB
/qcTvmGcDyQ348XbFR7ZVKrr4U5BvM1oiBtvEkCImEmrAKE6R/0JH0jngZzqIx7zW4KXIw3La8Ph
+NVLpp++IjjP7GfFFkiNlcgXjkveklv6k+pnpbQZfN6Dtv09PRaes/MprXKmLWww5PksD0FaXycV
wtc215rLCdncP/OajxFFrLMsKe1mPjwtEhoE4k6g9VhCPsH3kLVYWZzYkE9m4itv5Bt1PFU4LtMp
fTn5dXUBphdCHSPXlrENv2sXxgY3u3kDbJjqBCCOm/ThJnbyL8pn9UJK2LSNIizx0EhG+5VSVJQd
hUGs1ePFQ5fHLdB/TtLzqnQ9ZGoTI0yVQi3pFC3jZ5vKAiPp+v9YKj+sasaqUZMGJDBpwBL8O9Mu
uPKfeCJrhzhDi8fLqTrU6AsoV7sIcy5aEfk/cRpmOj+XJevM+OgnXfisIGZ0cXC674Mn9CnQY5yw
zL3+ZCbAjsBIojlIM5cTUI0JPYwVYxTOLTOnnqawV2ovxS1CktcNA2WmwhLk6xSfEmQWWx9E7UHb
Gzbll/WRYnETAkBVF6dr71Pg4YpRyG71OKEfd15jBtfhsTOLtiVuxNGER7TMQ3M7gAQevPnbkhlw
XChNTnNg3xU8jvTJXthUIWcHqDckQOszfDjK7/GBraGbjrmUmdff9d7ynbaAxQxXo2yPjOl8pXi1
NtRaoAiLt+s90uF3SOn1IbasXGNgFMZ67w1Do22iwvcnILD+c4Chf8IXB+Vwmva49Il1C4iqhI5k
zENEmv879Dxucm8hV+JxGnJIzZY1xXdugbZhiqQvpHn/hzI7yzN6suANSPdkU4tqyCd6YOxKw7Sj
rsjvhbFa1/dAcxtAQ7Oh2OO4DvLvzgFzffGFeJb6Wuoexz7Huey4ZPVp7221MFVwARW1OJ1BCrGP
jd51rIY7NgnVrf95lUyCqVnFEWhUL3UcZaDMQkgyO1toaubn/foE+xDwSamyfCALGOtF5xImseAd
h8fwmGpdgj1opXRPjnFsjvuiUgspjM+m/sngiKHpL5zLezxc9sDCrMZfdhq9x08IVcaIIyyN8xxh
cveaf7eZ91ma+CgwDodubziHECMyG3FM5+x/n0cKjKfCa198lEq+rUZlm/UYIJbmHHDzGfXSAcaj
yMTezKEDHrDvSwV/gXGm5ggIkXNFaFzejeoKwCuRH5PdqbvZkz+aduoh2TjtJIJy/m5NcFe3JBVe
L0brbSJGIEcAm0rCO2EWbDn3PyXfx5GReO8Puq183a3LOAzFHXW9z5zI2qhBd16/qe77MBIsAkhr
k25A7GxpAG2ccUjLHPVAGp1sxINyd5KEsxRD14SS7J8IkbNnh6MwLim69BmqiKCfqmyfPDRaghNH
A/ANwmhG/CheaM4Y6LiX+3W431U/6ZkbhYGtILcl1cqWxKQuYUvZDdS7boncjHARqMW7ylQesQbL
/xSMRXswlsl3w5Nug/Z2ItI/QcIlTacejNCAp8HAbx1gly/dm5qzdg+wSOhci8G/k2htxzG70bcP
BtLgHNW1CUeRzYMIxQJfWD6LkT8stwW/5stxgRnjnqqJTwM4HVLApQquOoZuCFnM+kI3s6CpE7pO
sngODwBoiW+DqKF49nfwHM+uL0JHczH7U+iv50cNPWpIHNBBs90LzTPfQGxFxlKc1cO7PEJ+MzwA
k5jmsb6u3V3OaOcPofLoKG8tp1KheTg84A34c+7B6iSTUgNgk4ZZaRcTZZAf2lLN0Iy4dFLTvpQ9
UYx7kwz49xdYQCmoUqjew7t77NhnUyy9QkRaR51iI2HNqJ7yPC7XEkUDKC3RI0VAIEwRbNZMFaaw
g1mXniGfEUMsJddKkhzPkGZPMTf+QJdw6/mgooP03uZCoc/cIQyuP2WWJV6uCG01wWbIVElJge3x
26A1li8rKinYHYoRxbEStEcJiMgmF2N9Dd/iPTqYDB/RCszgejArNnpjO1kIwA45qfW3teKyz0bB
tTfSsAD8PQFGNXeWnkwt1PbWikBEJtWBd0ZjJoVk9RHwRTrUH7XlFjEbatAjnDnAZsGlotiwnB8q
lVe555v4mOpXQmMZ+EsMvI2q34F7Kw3EM9wYRd0TDfdbFtwcMs6JK/pC22+cGEAxAArKA55+/HoO
RpNtepdhtWHZMOAGyPfQvURcJL0s4hHg3CplJ9tbCYbSgqDx5GoidymjKNjNtbncR529f3wX3Bkm
1ND645CimxtYA22tQwexmEvxOD0hwk/GMiK8lOzlnfIXM3f04gyO4yAvPFlOmx6DmfVbESW9MagR
do5qIyQP+9AuSUNIPVJVNjKptxFIyBvVW9El69Imu9JQgh5urQgJznWFfRDGC6FD8PpUftLEenPT
mwKBj1n0/ctST0kIuAlWZxBzd/5b++gFrpOzDVWRaFOxDNKIZzwbcE/tqKQ2QpiUxRWKZQCeOG8e
Hu1Mxo1G4eAeqChpdX50yTaKP2U7WB3x++RwBvn14bvRJRDOSNRn+SBavb648fIaqXVH9gmpo5Is
vRZTtdxH07LdLcE/0U2LHIes6DFyR52zM5iJn66HQ7Age0rwlbydrVs2+r5FpwV8zTbcsruuyIvJ
nbngPPFA/dPVk4gcUvNoVkL9Vv14QYwC95/NlQPjT5TBrRyXydfzkkA0L111Q00UsLRhbSdOGXEM
FqPwJBuI38D+lFaEGDcEF6w0RyHcP1nSikcWSe3seznujMtgYm/LTSlAmHErjMgIy9fpW2eOYeLq
v9VvdwU0fpUv6gx5jNQW11B/zauijXYr+b/KS/+X9auER2nwGvZYUFpNsJv8v8Xwu34xgJ7hG5zb
VCpy823sCcWc7tMOH/ffHimmrFpKT7YJTrjR3cyxRh6MQYI3Ev+N+VQylj7n+RgllCjFzgLFirkG
pyupULu1Wrw5PANA+wM4bIrnXrQx2I/beihgLdr+n7weumdidHJDr4qeC3scJoJt1YkbKzY9IF0S
vTBbvpXqfXAnyMeHgcASRIPymUeNDdy2IaIeMkfab+gZOH62OWaDm7RhnEGnQ8dnv8PPBJFLKgk4
dOCNCBAbBQUgUd5KY8rKJoApAzb5B+HvaarNhvTbBuXtogUWDPcOV4Fdz8DdSZ/+uXfu5rTWazZ4
wWji5C1BQmM/If+pmCHJTj2GLF8gwXPAVa4Qha2y3Vt01+d312LE1yhcAX0CbjskicLSkRKO7wWI
gy5cHHvCuTkQAcTeSbVvjhKmXC4gDNEmHqjckaqFeQdG9SNuqzvrt/kpH1W+gO9auMycZG2PlPWe
c9nY2kkUf19oEPdZIV8lyYHzyGDzhIHJ/n1QN83+LADfWIbN10oz9Ha9PjSdTXjQCic9wUoZBBVn
QDic5Fm2H7fqx4bgsnIPNF1t/tgmzhZ27NIBe9PMMXAE9I7jT46mSYSG3WnAAVMkV5ti9/3W7cNf
e34mc4/wUMUmBwVEsSSTWn7c27gSTU2ygEZ6oR1xReIC1vgZyoEWXsPqshlacEOTHGTqHOBOpq80
tdS6vbGJBMJZN4TRf8/mUO0VIuvirRfQbiz3himOOlpAHw2Mxkp8LKJT6dIUEkEK0X8CGSAqiSHg
XJMgNKnYhL/5FgtaHjGI++l1vB+bUBPZZt9VOeyeEA4XSWDzSp4VqHxLSOySxSIEglhAV+0LEWgk
MnOMXaobly1ynXnn7Wfp+3TTL0VFiBBubnMFoJmj6lJ9lX0YcqYBYCYru4vleBXsXz3lTkoUS40o
9AM1R1rQKG8r6PQUvly8+hc46XRuRxZXZG/LvoW958slVY1pMQUOHZm223iuZKmcQm0ksGKJH83G
DAWCrZ3W58RZ2Oat+obfaPZFHqoEbZEOgGRVsymTcjkluYddi74Pp9UfD6toXhKoAl4wQJUG8jPC
0+osVV+2lp3V7BwTfsD2VJ7ZOQ199xT1+g1PqsYC0c9pa7tdv5KVvUyr1xyE2bVAe3Ze2yz5tbZg
IuQEwkQejLyZcxZd6mo6ZhdQo40+iXy4hH9bpRZ5mdzIYXsQ0eKdvUdAnulcjlsk6YS19QYVDqWp
2nRbp6133QvpbnpBFxHqmM/rnce8vr6fOvQ1j4Q1+axw00lVr9k3vaN81917UD/T+5bzWxVvUf4O
+MVslLW9A4WJgefSxWS4m9/GD2lQHQ/iWwLNRNDnlcm/eHL5fQuRLoDEISAIA/gO4pyBSwD4i+43
uBWv8TKsdI7O+JIisma8cU60fxWnMQLJ7WvqxYq5t8lD9+r2Oyc9ro37PlF2DtMDnmw+KI8PXOzr
UwVUxRoHbI8+jIQR+8r5OT5rmrUVXFb1KH9BN3f94a3cyogWExjo64OqXzRExN4dqBYknvYrBYXu
5QPhr9/I0GUbn8qdXmJi0y5Ed0wnit2WM/KsEeJKdrt5ErPKXOKw25c6CYh3Qf/elAHuUmQqOKwA
koRioJa7YhFFOZtF7bwTsu0vwMzB/yqkm2NYQb6zbMBtmPactdk7BIUTRZqd6GPMTkF/xrn28pe2
Wr7H88DJwMWy+TaEdTH6671KJ+7Q43zRyWEqVlJ7TDmeP80KOzfhz2olmU8Yg5UKPvktL04Csvkd
p8mcg9m3FX+R61m5vJCCOmA19Kp0Z/ReCcR7bUmxi52zGO3hzYeuaF8A3icvXKy2bU5Rdpg7jboM
GRAOiGmvEU4xtHGsEq4iN80J+ROO3bQZs1hf/LGQ8qL9/gcnAB4u0EmXiDn+h/3WrU7hsfH/H5po
KiL7vNVijPyG6Hc6H9+IJYmErQqxZUrlTvcLQF7vbfh4of2PT8V+DycKyICWp5QvBm2nJCf8tnIz
lHU48G6ADsaGB7cDos6pSEtEiM9uVADY8wjWN8hylmmozK5JLlcPuS2UNmLHJJXQUQeWDscbzig8
ydmrx1TWi1cBqhGXoisG4La3GpGz7/AwhM0kSlZSl0wwIYz4us8EKvHLmzZFrSg4RwEeufJXrtJS
bbh/yHD7Ju2+t1gy67nDxyjqp9S/fzupa+5xcNfltQK+KhGqBKYUlYrxxaXPsmb2kY2S/qdw2VTJ
OnhOeDM+kVz88ynXZg880ijZmdkC4g6JRUELdSmmJN1PkKfq6iWmDlqohF4JTiBqyKLf/JKL6W0T
IRTFv4Kmd2+TsjTksreEwtbENDWhLiDS+l+3rzRhNvNMfMX1kJ6xXqPJJaOGH+I5sFQ1krWgxNT5
O+Yep+SJtDuqLovc7K1CqHJTWfdka/VuaVcFTPB4xi4smaPE2/O0ZD80VDahJIzBAB/Rh+XosRDT
m9niXs9qyvBUSRk9ruVyu3O9TgsgNIpgDfPm4f87JUAZPuGK8kFdkTwnnTJ7P+uIWC9XaDGiNKY4
DC2yrtNpyQPVp9gmav0+zvBBDjHOuO78212Q/qwrRqWbmNFj822Q3oyeWwbMWtWhvaWN7QBVyYox
K8Ys7645dnlz4kemLyrs8SE/ODY0rlGZfJFzAvHsdub9BGKvx50RIxljKfwSLnd7W66WY3TtaIuH
VT3Far8BC2oydIGpgkC3Ogx+rL+DO0wbgtrlyk50rkzaJVy2qHY1RbfiEUABEgtw66eY2KgbsG8q
tndGvy8UcWaYEBkCOqaYDPp1kyiUTUOxO8joN90I4aKA3YYbPRSqxvshO1hci8e/49wHGL7WbSnJ
tT6RyHRfSSClgy4D1fW8BoljiGaJcx6h9GxAe96XEWZIErB1TO8/mX0CsTh3C3t6PNz1ydSoOwRO
rYBd/C31wIPau5wn89ie2yXP95pjmzMFLthkJAtDn8AxbdLwZE9hqKi69vwLz/Lg8/w9SA5v69UL
vEWfy68gcPEQfnnC6zijXo7wpWZl4YqbuJC7PSKhNz36oC2NByNXagBmjBOodZJApUb/tlGvrF/8
TSa3UZL8E94PZq0GDjZzNkk4ZLM4mh0n8DPKJMLcIT9TlaskX+cdYNLuA7xcIAlmpOX+rzfMmj3+
3B8xzTz55AX7yVUb2uspNsaNSlGcaAFruD0djNjb1+81cwi3cz3lPl1RAIxV9FbHqg9kcsyiVsty
5yVKaDYfDfs1q1EUpznrSNshfiplsugCzctmCqgc3+OUN6sCqtg3Ys4fzqX03RWPb2WUXMgXeNVc
MSLCX9BuvZO4RBlUMp259UfT0NU3zAryF3dMh1OTvYBVlork34rRdUOrcFK19dcqAbRSpArfkzJQ
DxmIFmQqDPK6PNoar7xvbE5gap7Wzp1rfpoAp19cn3hqnI4k9fAPYjJqMKyHzLg510od4VdOvElH
tAOkRHsuGv5n5IVvYC2yPcd2rL9EgTJuNzSCjBMuavqN2zBTxAlJ36mrtnyk3XRw1AOq6UGNmXnL
ZZQrPzl6QBQNCpdCA3h53ERbmmJvjl/BzTklr5A2mkJ6lQGiELQmSNdKkDCRjTcqRSauK4RSAjKu
Opr7j+8vyE/Znjga3/R4d+anUjNnO4mzDhe3Daw4npxloypAIlqUbB4FCJvu4Mb171zph5ACzyTq
uBpj9NZ4ljSGzl/24SIvLHHceS8LljfIya7BORn6y8oBJ+a2Ztjp8gg4RKibaaCMPq1cjwdZNm4y
IH+tbjt0ufuV5kftI2nUSZJOgTWpNv2uIiJyp09Q91/gMmI1pzTw4sKH/8shiXdx48e4fxTdE0fp
Y4Ai44DlUl2OxsdacarKOUgBxZDHsLNnS9X31bCT830ZLL/yMcoswY1T/5KME9k7fMRRh2adMr9J
jgMhxqbNevclaKV2u0kctmqiSJRgUDzWBIKBvKidWjgnjZYd9riB1NWgy1b6d/y4NgRWXJh1z2+8
dZbzr3KIeq8OF3fMxwrxqBDOLNYM98/OBr6sI/lfkckYCpzy/Mug4sVil0WvTtUHzvMVeYGQZ7zo
G4UDHy73aPOtOirMXtWyZVa/NwW1Lo7r9BqgI+sfT5Fax5J0R/91P4VzNeLueIvTQ8zQU8BrXW4D
Gxz4ACMTfydNQcMGbNqRcqdcYq+f4W1PrEzgXse/Ov2zTKw1R/m8qf5nuS9B4DfvbkmyKX3X5Pam
IYJq4cbb/GXE5V0qcmq1FxCAKNfCEv6y1N2W5KTmyB67NhP015f64VATfUsOLwE0yAAFDTw6pm6u
vrtmlzLfTrvhLP3UOq1GEDfLe0WVNJXMB+ByecbMOuwY/3xVABkvjYgyO719DChK2S1AzUdgwcye
SESepKO5t2IIl6yZLGXDHeCrCcT2/3tnkHHKAr9E6v33NPOOxuxxFvtrMcxTttFaMPpKxqn70zmD
Z0qVCIG9GN75gNuS3p3j05ipZJwTty0pWa5x9T2aaPdpCEgC/C3k6yy7+cabFQqx0pbccABL6gfF
rGWiD93OzfoO3nUGDj2k7blmGVe+hqwRCcLKmqnXw2ekxpMsRDw9NASYcRo7QEQ30NkJM+MTj69Z
clOTJHRa1y4uEm826mjBy1ftjV7fqPc9LKP968/+9dq7rJiEYrTYtAmCJD3Qc+PcFevh6khNUf/2
AHP8GZUfrC1KlR1fe6d/CiQFZp0pg72mOzRww2kv/VSiezhcNYcBSQeKdyVgJulDIVImBtZWO+TR
b+Rwon+OLcXpaNkHsLLMepvg1RKzHr7Krw38RoI+2FkM7R29JLW1EAbxnz2uiOz/Ekq2jZJbD08o
uIBfeapQr5Pm5gMLamra+8th+dLe90ga2ostrXaTJr02Tcka37H71LMlJPoadaLTYn7bAEpMFkB3
I7Wj5JDazJb5QW6N8XFaNbvbO8xWGpQZRdO1bH+HSW8DeT05+nw1f2oe1RbcWPZHLEM+34c+xi1G
a/z4jGC9fKdsj1J90SVOtzenlcZSjAXWvJYC6GukpQZM3a9VUfwXURp/o64NKesGsgOnxcNQ85yx
1mhwZd/crYV7LogZyxwxafg3KkZTmmRg6Xh5Rd7u5STF1dFMIaGws8UNPo+dya2TfjBCeGD3ac4D
7UeYzjwkAuSaFpTDGCcLrn7f/HQaWplHy3Dx+oZvBsS4zaav37A5GvMMQX7HpQQrsITxIip7QDZc
WZE37+DDYoYmK/HRjACSiRXbov2zUVnn7Ohg6WGJ7PfUl3eWa7iayo9Qwy/XqxOvSWibU/qRd8uo
8l9H8K4h5Pwebs262jj6dJSWOTWgpJ1s+67BniGlFVW7ijnaQx44IZhXaaUDjeB9dfzo5s/3x29+
ASLj4o2VxLLK0u6Xa0xXBA+CkTiebAWRzPefO58s1u2Obc9wLFhpW5gsO5ZAEXdCOeL4CINLPAXZ
m79KkOkvX/Xc79eiUD5NWcDL045z4arqY2Q8mW8n9j82htv6UVjS9jHZog4licdNMZueEHzXax1X
dbDYMuNwpsujiwz+xR4V8FcvMwB4pKY6dcqP9gJwEQg9AwHzZ56dULnwpWUsDE4dtjwGFjhcMeQd
dnzpDwAEd6+VogSjEzgyF1q6G0sZdDGQ5r/z8ECexnS73FEfXyG7ex8YHIw7awDAAZq+RR3jiXA4
xLMuDVQ7qrO4PE29a9pooDx63dpEMN+4UY7l/tOfsckv7Uyorie0VoBSm5BaQLi8mgf5ZAAKNPVS
xVpEUrDMQPxf7i9oIlpR+aSjPLzOMsAA4Z4FfCxswqT5o9eENmHquXq6KQUreS5+N1gYkpn6+h3a
ARCvT9QsES4OqcoizqkZn5me2Svvkoc9ChcWd2nBo8FTPY+3+AsQ25LMh3MUNoYsibYnHDRZamm4
DVIisbJgP4ZmBbmGkwLmWxIvLVK2z3WHVr61d78EZWtT2j4Kb9eGq/e1haqNvuExwz8mjCK9NNWX
wyOt8Vu2q68zJms0P18J4RGRlzopi9QPXv2zNgAmgrH65i++vWcq277hoxDRTGn+KBNB4dvPSPTB
gO8ibSCHwJHAjOiZt4Ku7H5zadhtEFOMj7S5aQcoBAmCmdQrJUS6lhXehCpcAUdbMPsGTIu501RH
RRHX/vmzAgR1X4rrWblN4g4Gaw5az7KQdb6sgfxvwUSr6zeJf714dCEOYqEHtnhOAymXf7TPmmPN
9Cm60PtyijHK1LSzt8NG28B2UNe0bmaZuV8yKtitNiD9tm+ix1Iod+cWh4SrKwGmYIPZIADSt5l8
r6f/qZwVjiKgsVajM3+Nu8LwCZzlTDex1f3hvI9B0Ult3gBcaWETmMdwObVd8V3AY6P05YsIADcS
jg5irIExZBY/JusVEPhjl2sgUvvxTY4xBk/MGdajrg63Tiuyv54LyR1qmm1P3tmxSZ4bzgKJshmc
4qccfGX6gir+ht0AgDKVPk53AaKrGQaE8l48dDvDtUG9axNdSH6JqGuYmOXM+MAJBJdt5lTKCtIg
EG2vqFLqCnkqMumy0W7S5kvQXWvzw4YOJdDUhz2TGaRGywqHVcuPBKoe3xwoKVLaaqmOIenTasUz
+SU6tVLTXMN98o8i2pKCp8K1jIBFFPJ4FkrzL3zrkShr1Ua9dBEe/4njoZm6GH98pd+s7VqeR3u/
6dkQocTwd15L8eBUnFTYfPla1Jc1divVxCj06jhOD3tHN+ptACJ/HGOansGi9UwKP1zgNmqqksGj
GV9SwhH8H2KF55Rvpt8Yc1J4ZMHEW+Zng8ACe77+0kksiZ9PiHp/ZltBuzg6I3SegH/aTFpjvmM8
fX3wxqoncj3NVrQF/zapuwXYHLh3QvLK7vD5oBMGs5sGsfBNPnsLXCd3Z0imnNVH0iyPFkQgQms7
aVkdeOEQsWiLEhRYF7xCe1Jm4HfSz7L52BwFCXhaU6youvGzuP/UlqWyHcoMYvnUZ5BhxRkFV/hn
PukBRwPvUUk0hIyMiRZrDoXdenRkEb0iSF6u4/Ytal8egdKufBzV5FoiU7+QXFPL3kBNVFCXYIFP
H5XMKe/Y/PDMcnoZ2EnHQCIkrtglkKj9nhK1d/p61xNTgO6uyFDAO7ZsUPzeVmsbkqV0/DtseS/v
X6Fqtbp9soZYIfYx9wJBbYUFbyyNdF1qk5rclsUHGPFnIJRYMuryruIR8In1oye73ypoH54/IPMi
k8eqXbcPZRNckfC+Fh6WyUHObTV/usf2yuO7gIznEl7E/G37V93HfOviXw/6ywhJgOI6fLBQwTuj
e0vdqTbj7STcZgrTR+KCPnMSMf5LvVZ+qYACHfcXL+f0d+SX10VVLvPQFO/Bk6+nWGQDbV+lqsT1
FxPaMYZeVCv7enR5lcPxzz/03/iz2iwEG36iJ0M8gwWl/mLWaGS7dofUoQQguXl1I9esSeKhMaS2
e6U1Pd5HBdxA8BvrFowNDI4f75argTV4ffL+OedcsAFGHeDrd8GKfy3z12b4q9mdKK/LgWXotq1p
dGnHUNvdGvBVkRFvHD99pgKmqMd68b9dJNxQOkDvhogdGnRFSt/y/i+delSSs4DaNDnYo7a45lF9
2npl1jdKXMTs8FcHyLH/ThZMCYTqdY7Cx8EZl4r2gjayzpO42L2cuJ4CibJMChabcrH5+Q4jbEQB
GdzTQGLWs7wQZ0lm1HfuYS039C1AwwHgCWMN9kbMyx5SBb0DM4NO3GrU8+sSvaIu9+9aDHn1shkR
Fpcc56GPbZg0Vc6xzfTf/JBbRW7Fh9UPTJN0EN/MyfuH7pkhrW1cuIrib/yazXA86nXnP/xT0kX1
hRDvQ9BIb3sqEkfo/LNUYkyuoiuQLPLdQo63mavfZiH+i+MZzpWinK0P8CChn4L19VOo4TZYSib6
BJptDS/jLPWB67Y3K4nKbST0YBGdkaTh/UpF2UcU+DBsvrmRITsW7LpIWTtsEuVNJc5h5c7RyqYn
02AAO4oogXmiPD7N6DxLXLXnqkLqTzqwLvfzkWECOa1eTHRTaf6VJISchbJNBJ8amiUXENmyRPXh
wVHj6rOgYOKq6uU1bT8kAzmPpVQhuExL+kgd+KxVRXFTy+EmOHLsKZjcx+DstsqN637ZW4q7+2K/
UGVWz90rPqb18d4B5/AMkLDEpBZ3dXMHgrwQdretjGy6EFMGSWIDgPP8/sQ9X9Utnm/nYMO3K7RY
QioX0Ws18Mb7hdSpgs2RCbE6CHEG80LCqygfbryGytrh1UvKvH4yaVhd3PP8Ttn7dHjzJBozVl+9
Ibho1AQIrhzIQCzV+KEWxGp8ZZlZydw1VFGETILPuHHVXqEdbLkGVlPoV6wnYd8Kqi9hK8tSuDM6
jZXxmMDWQYNGt4Y3gsD9nVQtrih7LyYx+VnozPHGk9ptIu1pNDCjhtWkMCwpEMrLSCLmDrSVhvaE
FlCgiw0+XowiNoTpd+3k93DnrzVVnby5QlTcXvffWTL8kQRPYlS9/sPsG+dwcMxFfLIS5QUO6n+x
HpqHo8+4bJr9QpDUmsJSkDQJpF575DIihTvigNDah7NwRZwARFXBMKBzb7QXz3mvIC/fZey+AdVu
/YZEW8MWRz5t+eRRg+hJgeNLabC1VTIm/J8iKAuHmg0FaHl4x0JSSjcaXuGL4EC5aw+rgjpxMOge
05e8uMz9dxlRhDUa4OtofddUmvGfHQlGn9M/fam9y5gNC0q26m0zeD1KzLxSZW1pkmHHQQ2nrHMe
wXzcUeWnwp8gvVeidRQWjaX2dbGGg0keJ7oy5bvGD4OFr2az4ZP3ruAatn+1NqPinc8bC4n/HHmo
hPgUmC8N96ap21YnvhYxlwG0S6Sprnp33nw8lVOMikK1qh7xgmQ7RE1GgDa7M2qdX6D8EegAkQLN
yD+fDJ/bhgpyxiVTdOhtJODoz+quzBq6PeS7SdwA5fRtKI4qk/c2TSeOfXlRaxkL9pODbqhh+vLt
qTUKFbCWS4eYU3OcTDfTW/vuwowtu0u+YScodW+Fmv9yK30fY72OfJW2AZ2hpkUmw3R1GreToqd2
rYjjKeCyYscFdguqG0u6CmsnlHZfUIvngnMw4XhUghekkbsWdvW5TebI/yFezTICi2l1Dsnw08oJ
PAblZhVvY7d4pKaN4aTBuL0u1Vsk17bfjrNbJ//LpTr8q5Jgs0I5exnMj5MrTKVO7LO02axsNeIF
xxKByAxoYGgnGoyAM67ArO8Tv7K1QjsEiVTqoT8zVVo/VrU1wKE+79uycXMUnL0D9F3hBDvZMFpj
6GUEfcTGl3ih58PZoDNs7g2EleR7et1idZ+0CumbJdyCaegp9Xga5SscfPPLUmZbjyKujzDCnfmA
lWFdc204HUmKwd86Rev2t71MSbc+oVIT9pv5tnpUYsgm9smTtaMFmYnc9mFl31IFW/ipLrG2pGyJ
L8KeJ3fH/eIQsXmDKonsgE0O4rDIFfy9B7g1TNNRVEfsXA/j1tB6BJ/1th4UtGW9r1xDAaw6pWBt
Dqpr8T3pNRMBZ85DOXY/B16x1+NGxX5wov8gbzRP3aE3NJyxuq9iya8xzophOrGChZU+nohJFhlQ
cF7Xl4sp90nBv9MtOfT3jbIYqD2IdhNuxFFbluT2hLnWeaazXErohZbYX4arIXzsHSR3lFQ15/sz
rOYp1fdTcqF4xA+RuyvVGMTNzErsywYFnVmawEXEF+1G/4skaChGBd5g8Pbk9/CsI5R7q1MOq7zL
SF+aCM0p7wzRKgbrqr2oUirU5UJzZTV8Ul3xgHscytqj+JGs8rrOycGqzQxYbVNAh944k96lEFr1
Dr63YYXXFKXvNfYzdsFBNDohpPPYxrnxOgEtiwxM0VQwCVwS5y7oOsnDXVmtsbrkm/Bro/Hsx+b8
9mDVQ/UbDdPQAjmOXRXyDreji53ES8W1Ak2TV8nHXASpf0evBMAf+PrQEWHfVyhoxxkMuruKNEWs
UFq6orAna2ziExtaUYHhmMhV7C+JiyobNwkh+3GYnTkMLzWbAbiMo9pX9bNMD6YCi3t4ipNnCQH1
f0voi/AeYUQP1fcdKxH2Ehug42v1VtOpXjf+pOYP1XqNNupmZPRGjCtcMeq8SkhQbf6XIjP7wzqN
zuarsLmQb6gJvZ33JygpbixgYcu0Wgac1HnXvAK29EuYF0LaEuZ07X4OJsvuFceezdDjEzz+KXOM
oTow9vJP4UuwkR+ITnh8kQ2EsgtZXgNzur4XpmEUg5smru6b+G3Zmj9ZnA2jGdhAopMVPzM+zRce
pnB1n/zQKlUB18nzJMJm11qtJiMjVTHdnOUxoXKSb8HyIqpwqAxjVD3FXlMS26N7xOTTjdZ1t7HZ
oul5IRs8ox09w2a/HsF6Q9i2lmDzGVD2U7ZL79jfXq6ogPgWXMMeH1S/eGGBk62qH02i0jMKb3cK
L+3cP4MeQdyZZBeWszfV9yS++uEXKr5oklghEFuUsd2B5uwyFu4IBB+p6JpGsUjqEDlzZBVPuTFH
yMtErQDtoIxBpikJFGrY5XFIO2kkfgznWtZyXQZpB4t+e9XHgQLAzgMGLpEKM5dwgw8dpeKkTn6N
JP30oH0YbS/h+YOTGXLQ9f3MDXT+Z8lQqw40CTLN35zUP6xhlfIZ6NMpYQlqlokbOcMlzYOvWLgK
+K9InVbCuCIWIreRYRrol+tVMUs4V17EUcvpqAyJxtFNoZdluXsR+63C651jIXLGAv4OER2dLHE6
WT4PgCsuyK2+npSivDfFS50ZxDKInq61Iw3CqQjPu7tl/4CsqgX8fNONzzNhsqQWDPxd8dH4x8q0
2cgvesluhKseByjfmWoybK0an6fcJVXc0enljTMsyTGnufldEXNUPDas4qX73GRQOR6RlmglYwAs
23uF4wWBHGlno/BBtZ7h893EsV1LAcjt0g6LJMkgomdwn9+Suut2ygrPAlUUpsth5eQJBkoO7Qso
wiGDz4+DE7IGl6jWp6WfCqysftQ10Ykx3uQ/UaM5FC5y+JrHQGKVp2tQZpsX2W32EF6KMdpD/FqG
Psu/gKG6qCmv3Pi/31nR0xOvcL+8iUgJ0/mFXJuCA/q3yfHdEc7mjjtRBbjzrrHqHX8xRphcm39E
YH8dXkg59EeK1AaeUqtI46hq8yR4ZoD+7OT+WmMRHvOzLsENRE1fWrNqpyP6uFble9EU0Eaztdix
XruSXFpn1i9ZMcxXmvY/xQzjLI7sX49tz09kLcYSZclIiOR7HRZjRrW9OAvuxrExwxvJsYmgUY/Q
jLQV4u+/8iO1lWf5/nVX/4KMOECG14oikUvpZMXjlTbyIkj00xVU5iK+ISqT1pnIrB9ZEeuvaa22
yUJs2NYLeR/uiB6rCvIMmjTBQ3VK22GbMhcFc+vawFm/E2h4whMg5dBYwRXQK6VE+ADMu0LRGE8B
NEA47itO6zU6B/RYgFEKOylAOtXAr3hx/zfNLe6JglJQvjgUmYNVJhYhw3oTWU7qPXEc97ms5Igm
SdO53g4ya9qE9IBAsKJyvNk+FYtTa1aVglEKKE6VEv48ov/uFfZbzll6xaS1nM550BEf4jHXMTsm
lsf373lt8HY8/p3ZI9Vqn2F5/jBIiutmPf5igMhIChLM6D4lNGCjTtpKKOnx3GEVNfqqT/LxJV3A
UXusJVyTizDeezW88kdw7YnSaQk8WTBZU9EpSa3xLJR1Sjrbjl4qAiV3K8ffU9DZoHbVUvH6bJMv
NPSU3UZCZe+XycFCCUxsxuRn2BBQW5Oz5QlkbGhOIbnFf3CtspNbHtlRzOVNMfyO0yPJ02ENgOtq
G0hWKrqQtANImlPcq8XEqrjQaSH3bD/v+968fvAVGqijlTQu9IakNOWvTDVMmAloNWsIZGfJ7G1G
Ax2yfgLSP9IsDAPf+/fogyGaRsA1pxXzJBYBdzkNoOI9EH1qZZkLJnOQI6pZophLx14VNqaB7dRK
A65QIZzEmHA0nVM3XX33Y/yKUK1NzhNtMoxcaq/I3Y72z+/Htxjsf7oj9mlNrMQZVR7xw8xA7aGf
ugJROYsV6f07j9Ppn/iE0Vhc5aBkPoKw4SoCsyauh2dTbJBjfdazERMLrixSeAo/1v1a9mnG0kWa
JpAo75yuLVzE9+epP6n3no0bzmn3sCxGmKcWb7szcQ/S60dSHDj/KHkxqyt/R/HBhHSLHSNJcbbt
Kt6vmUpuN1tO21BlEBvPp/+4ZHHtgVJgJQa51a4vZ9PxxO/d7vFDkT7l+KwaFKb1m7rEs1Mhuz+N
lqKWH3cmHhGwlYY9rDhUkYur64gdalmMr3RTJ7VVyuo0OPQgRJCAuuTBGs3imwwYDYHIw/Bx6KiU
8Geo6oJGuHBKR+IDDgn2oGs3M4kVZORuOXVGNKOksAFeeajnk+OjHKzcTV7RSn+BlF8tHc9MuE54
/OI9xnWDRuuqW4ZKKBCFIkRY8vQj62JOj77M82Hc/nzwlJHk9LTcl8Ie29dB8YdGp+JsIzMoS1Sl
fRmJ4re0eg7vm6z35ABbaoqp5iefBrjcLwRPiFt+jBFul/TXOhv9tdVuAj86EO9ZODtnoBnRMQgh
ypTn1EE1qJsSRSPsrNK9FR6NzZ80NUWQVteYymDx7EeY9WOtlNI/JIvZJItu+5ypnx82KVPDHWd5
0qn15tQ2oRK+yqzNMG/R/UUiMqJuqHSyaBhhbzdCkcq3FoF3i1UvOchBYJdhKWkZv3y+jPkzeuii
PskAVhMII8aZC/NRcC9HhUqf/fk9y/wibZQcvgUCxiOfh0vWI010HwBZeg2JBCHof2qTcLecT7xH
wyP4yXAlva5vR8wlA+L6d++6hA4eXGh6fWNXV9BsekHnoNxzLhD2hlcjznIJKDIts/C3Dca6+NxM
tk1UKI+HiOwZ98dZztgSqj+KpIdgm3YpCfIsXOwN2UtuhQrfIte6KnneFCzwkyYcBfYXZVFbk5oE
dft4uI2uu6WdnXvYnsdneb0KYX3L7rz8kGB8i14kmtC1ThbrxShcigtmL6rWWxMSTHyj6LXO0FW0
vbQrS8FGmh/dCvZb4dPapqK3vE1dI+JuT8UiX2g/8usNr82Bh2/ecob9VT6y/CeBf2B0HOCnPa8H
abfC5EIsx3rQSE9YFB/5MZwcV38+DYYoA/jf5gjE5TMh/Su+3HcsHyvwkImzHMf2iLxmxfQK4dYO
90k3cjxW5R5/H6hvRPX0nW7e6+EDWvNZVyabmL3i2eqphk6hOeOKjIeCPWzN1QFZZJmhot9wMe3H
6yX0atTSbTlE1xnwli8eCGEG8Y9cHt2YfyefWxfaUyMsmTX+TXfH0w6F8hUgRjfwgbXk/NACFbFh
BbKt1R3JR04CPnCoOAvbsdWFfX7OBTq6XRrfVYKlty9+qwIApy5StkovLVjbcLQ3BR8OMXwfI7Q1
y+iZr175fa4IoWMZyyP68TJbDE7sr76xop+iRtjA0wY2wYVWqS70IcCbpSDfgY6saEdE25smN5HY
lOJoMS2KzdXbyUd+DJGB3TEsjRmZqfDKHPCKPS4PMyWMIF+BV8Pa/aX7mo3DBm5J1Lv0TdZSjJoF
behMRLdaXlCfvdMmkkaeLnbx6EBAMnIIjT6Fjor4mdzd+HqvaHmQ70y0QPFoF4l+ZEv2RVQ7e8zk
mEeW1Ec6qpvA4R1T3QQYk5SxTI20oX9jDdHKqZ2kKzd1MC4b4CTT/w3/jpwyDa+pYGPUm8UxX9Wc
tL+Zz8mnmOmi5LOykl/6A/EeTObJOOSBTVdz9XIPPo0g8U6u8dp447Ge9W8oexePSaOgyqqnoK/c
p++bGSUgpJvMiYSlfEhvEJfEYDD3D8zHay0xStQBfA/FmNGsntshdS+jyQsveBmzzUfkkkVpme3N
6Dv0fYvNBzDqVCNpw4oI9GWz+Z2hyXeWgVO7bClTljtcT/vnlnPTB3u3GscLBD4Uqj1wYSU8/f1+
E+FXLniYitzT7uQOY3yFIEwmkONdJIavX+E734OH25YdQDCnpXaZyxFxge49Be6EeYR2AhdP7BrZ
4f4Sw0E5SidOznXAU78sXgKBFZkJ2HQc9TeIwJSKJYh0EjOw+kMnRvvIfMPGz6l2zpguXvevDc88
KDe9GEw7kJHWqX7p//tC6kuoCSTLCtUHJkjst2QlpbM6pjNKO6qioJlBYhpZQcFrS0uT87q/J8x0
Ewsa6syhMW2MbaVqbb2ddcwHRT/y2o/tLkKyIAiPGfdmdiNP6Iv8zZmInzpPTqUhxReWrtT0IjER
cWwchbAXr/in6MihUYhPGn2TBgQMqG8bF0+0vBVBFyWt8R8HNifT6YlvjphcP4paSO9AA3Gqu7Nw
TwJvyPKPuWwnkcbCqwUpxDuOyLxTpPyNHCBfThhHpqB03ZaNEYQqqu/06/TOntXg/hvmO3lB983O
3srG7eTXSeQxjCHw012wM2sLoPZyC/kHrmBXyVk2R2YMnwRKq0Ji8rPoWYLBjKQEezze+HLTLazd
TinfOb6S5q8yV7FNooir7fP5yF4fWTL11+sGDuw+i8BAjHsd6bH9A6/Xzgvm04OW6yF82G+s4CbQ
bqhVUEHNdc3TJx7umoL2pzKIqZZYLv16eienTYQyajSbDrB/v9AGZxuivUGH2nDrWUlYcmnnbwY8
g28qbEqsJ000i6Par4H4rGmh4yN6/msyTM2ryX183tom/9sTsNMhCM1xdITtl4R3KTs0EmJevAXj
2yEMpamNxbuLzsirBOem73IUOUh9hmoKxGdNvUxdfVnQP7+de9EcG1NI9pauJFRTJDZZvMDl/5Ns
RhMEwyuXEo0SE+w99TaQIuHUbU+xUuinkcFN19TgBKSqazs/5EbbJMez+h3M+Di77jNGpB77BI14
v2vSVYHEOkY6gfUagPogvCmXYNJEW3E2SVLA0NyoCDyw9EjaOl4aFbJzDQ8g1FlktV/gDt4eOKdr
vWqrKC4KHlL2Ekuh/x7RszNvXgACfp+2PznfgWSIfrkCPkR/YQsFoxX8IL69JShVlguopT+/bf94
oz5C9l/tZdsw8OrGuTkU7yf/Bpr8W/3oAke71xs60oace5bOpQCeS7Nixfq3SI0ARCsrEPGDpfAM
7sjcBd6ZEm/bA6EQSvl1XTt+j0CVajVmLBGqm/Y0AB8kO45Q2KC3sTdBQ1TCIG6eI07wT3py2++v
gHzsgsOHT0haX0p8K2MY26z5pWswtBUTm34k2cku10AetML0bjEtFbHbssZYp/zJoQF81JSSfEYw
O8mWWkq9FX12UjP6c1zM+AwfhH5bar3n9VuIiWDwpCFt2eRzw6me+by32CPgHGitgfi/i0dBRinx
kAupIxEk+2y40TCqAK3dM4cufJX7DXPe8umeKwjO/i7AXa23yKHN0CuIRhj8iJANekULzugJcRyW
aFQtPF/RB/uknpq2MJhsSwaw2xmjgwwI/KIWcq9GReKyX/la5YuAC8aYo0Zeevgt3k6ilNn1A0Yh
sHbkEqtv1NBgSyQI0Qe7ZKJH/BFbdtPLVIWHhE5CUoHc1c5PWGDfDMAprW1NS6gO8LZWmBJnGC5o
MVrSkFmqrNIgZ7SL8/nFX7o/JjjVvT2qv8G31IYNwqIUIWKKOEvBMQvlxODN9RMqASa53A7Ze9eO
p/wlC5oGvZYCk2s/eZVygL+shzq3Mb/kwDh088LxuOuX4ZacDWx2qteqxjFJwLLel8/P/WNP0xCT
HvIJX6I3S5HzijRpC8aiizROmp4zW0ZfmI1YqhXJynzUtrjx2N5QnQ3X9Y+A3pveNMEzlFHfT1XZ
5eKHcrqNKL+NZCBcv54/VauW59otISKXIvUDNvy5vUz0ktllVfFQShgsWMF2JAWyJYhoASGkvE69
w1VmWUUqPmKd7HUj1TMo0c0YkRu2vIxFrTLnPreDPKL7tf7CKLj3Px8A8SDAeo4n/HhxbiHUqxZp
704Y26aRwSR6AbmJ1+q72CbIN2EZrO5tVKDGaxafp4KQ/7zvPrvdGjZNMTELDjHaq67RBLWV378l
8jVlHEUtOHX5qWUg8Q4NTkpxtyaOwYleHxRW71a2QklSFuog3AjYwUIYrGqEpI/PY0z4hi9bQUmZ
y9gImQTzls1ojGYqYYY9vUbmtE05kzJcN37QIhzpkEmBzglV6yJLH6gfhcgodWKQibOlegGai/JN
kL45ytMDF07bsyfQhaAGCnzlgcj9Xtjis/a2Sble8nJIFbZbPhupbpPVoyKdqblAEgF82dnEtN5/
8nk9Jx09zc1XmXyoyU0HEVYT+3ryXlKIZ5t5Do0vQgtXmi+Il1GOZJocr74M2lfOMvTEZwWqoKA+
+zARnUJ7JnRAjC1dISjms7pl6fMctBoVO9f+K195+d61C78HHRQPZqIAnK0VWzVjXTGWr+F8mBzx
VshgEUmxDlbPQO6kgNKl1G75aiV56lk6zB2aCz/YoCnnvz++8epM814/h/jzp7U86xGjZCiczec2
mGQzodH8RuzW9tUJBPcJb4NHMl+TmH2k2wmADyqONUO49Y1z5DWmEjwQPulc0nZIAPwrjvKK1sTx
AdnEH9OhEZDb5A18koapSrZkcCLM0xzZOhFc4Cz4r4vBuEND7j8VmqYfa/PgzRweuWhVgB+qPvah
vHVQ35rDHwcAwsVkkD+To+m0L1oD4VlLPO5Ii3Q6tmKh7kUoq1Mp+9l5s6NwKUeZjU30Mrc6ACxL
9ude7MCn7deTij9zd+COPp9snaf5oliwzBgjcArJpTR3puF9ed6EI7QX2elQaSaBNFTeM5gST9Ay
9EG3cZb+fUF1KPMY2f2jwUYlsmpG6j058YWMGMdtN+593S8XuqRA75oppCswle4RFZn+ksXZEjrR
UPj6HpR/u9GhYVVpA4ZCyqb1gmMrNh8P5IRjJOF482lxNgRr0i6Kc8NCvnjsS+QlT9wSB7no5ScC
l+wTyXdHptpWIwQHCMyIO4y0UbU+eR9vRjOtCU67QcdrmGZJLiNpkGFYI1rXYEtTO3I5HT0Qty5q
BznaOI4tWaqykD71NHAS6v5AY8RGo3Zxsv70Niee+qEn88n4dGGYiDd9bioxoIQaI8bKo+BQUk1l
si9zRKOIP+QI16hvJ7QsMFTbCwrjiOKwGyQvy0TmjJevefkSE6XlnFNI+8GPPidQNYVXOCdpSN2M
r8+DAKXIm7gSTw83w4E2UAkQY2u/0SDMq46R7ylZKxioykwx8GmJ6AxyclexCx+lltbnIilYLMqE
19gRGUUSXq3osAw2wlTWtEB+XyV2dPi15vbKiKGKtF5xP9itJviCrg+96qclEcCW9NvGWJen0d2q
WT46gwNzPrmOBZgx+vIEgq92DgQE0ISPSlW4xKy0DWRWMGOXOVWLqFrmcyOe/yyanA8pp1j5VEDU
dbXozSt+rw2uRVBvCDbOsMY+MrUx2HIIjP+ginSPUEmoTKYsgq5VYRk911YP9XPBhHkaWqQeGV+X
XFZpjuJGVvG/OzJ3PMjVzIddERC2t5d+gF9e4Br1+2dSNtLtaU12asojIoaDYffFBYJ6Jm0uCww+
kfeKx98PrMn4iVtDCbLVDmtszFc3/4n0I5s4g4FgeYBvY006yRFBGtEqwrEb+oUJbq+IvdRAitfy
r0ml2V82EmoZLh1hWds272fyFyMATJWVGb3nLo70E/ekTmL3GMiexKgIB97Sc4FL94YwPcLVLJdf
0wFx6jeDMlXjcEVbgJdRebGf1VHJtLNOsUMq+fXQaqRydw2EGLDSyTKi8TJd312HKqNxig16AiWr
qEmmqHAxVhb05tVfidvquCX+1OylRiF97p9jllZ9zBKHpDHcI/wPqN2sfOv8jLYFVehWXabAbmRj
7aiGiFk5Mb+UH7BMQpHCwV9SRJ+xLUE+wFsBiWdwXaPG0/YaMA5gyvsO8JWLN4L0uxZtWt5edxAz
3DXXyd8O09LGo1fEQAq0hRUFbG5/vtswYcAFxWbMHVz8wEJL+srGndhvpk0+yhWYURJ4wOOJgSCk
s3yA9Ye6N5HorzV9nOFRwxDanmBVRv3hnmGwFAPavOu33AsHbbDu7tU7jBnP5HqNyUW0EZ5XevEk
wC5qRtVjvZX057ibJ9RPc7JbfCD4JmydySeRNraDEwL7O7s5CKK7IF5E+wr1KfpzACxvDk1O5RZU
w1aQC2mZiR8WPz5B7t91nNpAHMG7K23mCLdHsJUcbGgzXuV6uRzIyhpQ1Cqe4icdULAxCkN90oBF
lruK+/Wd4FWwBMP4XgZSdBke0uW/3nL/oWg5t9bawrq2Knc6lbKlMRRjxhwoufF/R0/C7GzNRXIm
V8OdGHgI0QzArzKkal9xFCFnG2RKf9zTrHChHUVV2RthZkBVJC2TCKSI+M8GtKVXeyi4iQYb0OP6
7fCjaTBiQ23s5a8S3SYbjKTz7uL0h1XBPI8spJ1S3FBHww89Ivv04zRZVtVKyx/aI+IkYqThSZ4p
tswwhYUcri0yrMwvnijxJ/hXeARcd5aiH7wU/FrcrpZJdW95DCXd5W7nKxtJJGuf8xXENXGi0Az0
0J7GsOS2UN8bUIbs6pqO63/c16FcLObGL+W9F0oCnlWMUI18sNcZu6F+tahG7QzmwLD6gwSgkd1G
RUsz0DCZqyVo1dzBewh8iFtG0vTrRSiR5L1kpwiU17P4lZP7CCCpaK4u95b6YdhBu/l/trnWV309
LcQId6qDytpS2GPgl3X6w9a+UYY1yufqaIHcnkbeYvEIx9XHnVxzePz5c+d5Ixqx71iCeE3ZE7li
k6houRwzPvq+r6jmd1DFjDJWWQadxGh3PGH9kUVOCQcfe4UOY2nz2P7k2MmOJ43+1LzPhTGJ71f4
XOUMXGr4jlWkF82CSkChR1h+bRKHs/MfMH2xU/RSFSWvWUlBYoHyhWvKcgXq3VxVMn9D2iEGTU11
JnvX4KUIsg1hhpbCMYTdmJuChb1iwrMUf8KEhGxPHGM55m6laVugwpm74Mpt7aJ2JaMBQkWxWo5i
YTWL5meEJ6ojOGmo3W39Zv5EvOMHp/VMjHnp+tw3iUL7iZi2xvQWaHt/n1R8BYpog+pi7XQcyhhO
uRERmCfPASDfSgQmwB/woNoRA57UcoEKraBQMG8SnJSi8wDnAHvjnMANz1S7v4saVPJIe553PwBn
cgXyuIiM8zRvuTbiaxxxz5yjLdAE+mKhA7ESZKtebWVJA+qXrWkBzzvprpmWsk4olPNUvktiafpF
iHPSM2ErA2N9fZ/f2I1euTBwXEW2ETB1udhLx9dWDI6T9dP+3UCOUOxvn6wBPyYAysP7I4DDRARc
+PCHvXfivwHfVj5Bo8RKIt2dT/d6BLmIAV9GvwepdzBZhZ0JL70k8CU1ztIJ2QzxbJTqqIYT29Eg
bIbaN96x0S+rbiuCdU64DGg+mmM9VgC79mfTN2krayynZ6TrSXLlqv2oLkgyKLJmZrbHlTf99Ing
jbwMjcIfGTkmD+BP4l30Q9YjzCmOAHvweJCeVwvxl5f/cDyk8zo1v/ddOudebeP6OyPEJpfl2ESb
bNB4Wh7RqAVinGwij3+mg3es/mWiwty69J4RQ4NqtkEOfSbzga7lYM2LC4XQimmmqUkLgc3gOAvK
6dyh4CXuIfZUZJPZM7LnqTzqKLoOq6fECBeuRZFz/ORlsmYQm5EKybMLG8SQ8NQwSe1HHT5/qiTl
G75K7r0WmHtmitzr+I9Uf1/o2oi3y+g2n+U4SZgmtwCgDer+m70rtL45J08i+WHP0K/MOtgF1Gbz
JIcqg8RjQtYFQ/ahtnMBbK9eZFyiA8017tQUzMrwyeKAHkOCgkLypgrkDIkTUnYfBceytfSAFufe
EO7IwdLda30N/0L7gnDnf4GeI8K6j1G4i44BrsonjgEiz6rOaw3/rarNqM5PHj4AUsOjh7BVPEXz
63WvGyidkPoCkqVkDz2EzxrgsWmhWywEhCRfrmQgFcV5SWTQf1XtJP3MOAvsRhwqy6/uLI78zbmT
EGHn64Yi0Q6qMKqPbVpmyIAS41tiN5Wr4pmP2p2m+F9I+9Z2KeUhDRPMG0pX/cJlTR7AIJanYhap
LwpHOAgrV82IMK12VawLB3gms3TnUD2ZFeYhH/r0vk5sAmF9LrD1OUNMocrEaRHk3nDErrWd5o3e
58oG0uWYex1HMBtrdrsCx3YbDZ6CyppFQWStDf4TJJbcIZOz46Q6pEnO7yoDNMMGfmqeXHz84NBb
NWQvEgbA8A+RKvEHJxLd/NBGYUPfJUzMDsHVSIWlfP4h6beeqSV/KHBCG8PqTwS+Z1UoqxMc6fAv
yDDYmQzPn3A/5+N1Ir6z87uQocXBMat5vrnDbxxtpkMGQOVAoMFfrMGSMsvGYxNpTKvGIS85L1Vx
0uC145+vfsHu/uLfo86yIrSt8vyWyiJRFrVC12lKa6794xzkW1vgPD5UyxGRT45ie3kv1nBCncy6
256eejWBpS08hK/7p6pCKBskNpPS20h6wjKpOy8y35+9cgsKPn2hz/5iiM7aERGgCzAHoS/WXjtB
2dv+2/Q1Qs/GI4eMqNkTuNKlqVXYTU3RB7iops8XUTAg4zJk6nifkGI7sS5mCQ6CxfTlilUSj6pt
2To9pJQP/FCHeeGb7xMNqWf+WtDjpTuB3fqASflktyA1OYRz6Tli6/nx3p9N3Y6CzF87Ko9tAhtx
wqDBKu4Abwu1TIJ/tq52INAUlfDhievw8jmiD3w2SQbPU6fdLKfSR/ijTx09/m0tYTPwtMb+f47A
SGBRBheMZp1LcQlsfeV8uiFCxHNynjytI63e8Zj7hj8fh8RZewPILWQfrbGFWhxz1EZ5cCAXdJi+
pHuy8L9nRuMP6vSN/Q89QQWEwVfAjmM1aSbSprzZfckvxxfdC0Lh1S4oJrXazeFsWcke0NO41bWl
MgjRaXb76eMTKXvo9AlZMpOD7sq2ngreYhCXeewmjbxaxkpyInV7DAFh49pTrgx8VuoAoSDc8Ssw
fnGRQlf/R0SaonvA7W8t8b4skNsiOdOd5DZU7dFXpFb0Y2gPTwbiEqGluYvFyMqiLQvcaThqrkOp
OEc1prdh3s2zOnsgg0fbiHUzpQTuDkAQyRHR/apfLYem8pQtBZ2PRs1wKOwQcTxNUKtmdHwdC88B
EQSJpL6ktX0nTqflXNYijGNVUuvNhIheIEefWIBlYefD4fBboPzN4Mo7092RDbvvkMJO4bYJLwgv
P9PLWvqFin/Sf7wXAjKNZA/XXPLKNnNQ2fSoY/Xs3CcYqe7jYtPPLXvVirRXLyDokVAucK0y4PTH
soKieHS/bqp/L4kYXAELjDqrrEVGngVAyOyX2WRF1r6GJViF8eoFhZWdDuhqvBaLa+s4yeRi9HH7
5WVxZcSBSASjup41gZ4nGGeT0xzEPajQUcWrMaHljyf8oEUftmzopaAIU8rqX6J9Ts79zurq99CZ
Z9OrOha1hc7KJvCZr7QrmZAnFzR2LU6dFKXzHcP0iYqjZKCRcWcPre13c7IjKJ4/A4PawHW1CW83
iCqmJJN4Hf8POvR6NZKYtk8h66L4YZb4IPhLB8hZTCV7HGvXl4dpn78qIWxznKZ2S+9Vzn2AJXwJ
P6PTvTO3wRof9mtWfhfqYBQMrAlZ7jDDI4hqfzuUUAjwTx4xszgxH6in5opZUYT+ZhVGfec/RaMd
oZVjsyPOdqjT0eJh2GhzQWz0LoPok5OQSZ2finyWnSzE5gis/zi0lL/2pWzU7YLZZtsR8Jz7gx0b
Ghd7yfdbJdSnzc3/TTk9R+VJm79uPvhO1r8863KP5FnI8hJuO0cI3YBf2tyXMYH+NDikD+YfHzY8
zjPdACteIM4yT4ElFvA6EqSnuBDNFdGNEuYzfabLLKKCbPibWSR/LL7zj+UKa9DjAW+VBMjFjfIj
NMCyvqtb2fdMhGP5Vu/3+onieOPRAx1Nu3CZ6q32PVjVsyUCmPhvndBSdLhcy3e2AJDG+IKKLVoc
XdV10dXUz8l5H73UPqEcRIm+YYH/RI1qouYl+PNpN0IeYYxG2nvnqQXICJNRlBe5BtsaHodgFckA
yWUhnxRrgUVEx70vstKomQJ64s/R17f0zfvTQP5OSjfBWkMNl2s9PJxB6/i/praLWBMMVaoP+62N
Edn7mp1dlkvRnjSmQqWo1R8ukFLIEpnMP0gH/ISR1cyNndJ6pmS2VFgpvaxIYV+rF9iPVhgIwsxI
qihdqS0dnVivwGtMd2GsqJ9/ZcBUlJx8nKEj/a4AxdKjrArwHHbI2kqnLUtuqJz0nUPto3kMuKD0
UaluWOvFR7NXrxyMv0E1AaldUnYL2C6PajC5N1c+sTiKghesjdpwojOfCwAiwvH6807WTZjTQci/
YO+GZUCwduUp1hKwU0zEKi5ymRc3rpDCXTMssl7kZ21qHqA3jAUXgRtCaPQS+/tCzQq/NDzheJfa
oPV5CqzY/rkUEhOb+csQR+YgNytYjtNT3J0ChSDJtCywF6o+eashTtjg5klP/oQWGgRv8xpL/7yy
9ZKhF1x/ptP+9x4QDS7mxs3FQHM2uoD0bgNVcIFdR78imJhUD/Q3ODqi9rCcyvs2o5CBxRFGh1fG
hQHfEvyG8kEoEsYNESZFTtrZOBnK6sH9MWUq9hqnuWgpGSMb7+H+i5H20b8DvSso5MhFSXfqiK+s
fID0m2ET+Ujgo9EGkYOHIz415/VSyRy+v5eMYOjdYGNNFfmQcnvIiv85CSGn90n6AtN0XzA/yZR+
VNNCVeIBtlshy8/0mhvaZESrH74/mob/jfdzw/SCzDeaH0e5vSm9E39LxiaLbw0+M/K2cAsPaN+s
CsZ/geGk4/wTc3kAQDR8Qeqnm4owOllg+eiaNSCKDd/yOiTt6UXjF05owDPMswntP4abg8gE+F3Y
lOsh+LTKcr3R0gXN52mTjrnO+ILgkMFUfYkG2vrJWeD/cysyoOT/q0A0BrhuwTGa6fKvNk54rxs2
BUbKvQtTkDihshIZMpBQ/ZByuyLzEZU56KpxCULrL1CK1shf3ch72EXvS9F17tCOe9LleFX5nVlN
uSepmRO8pgdVwYiDJD9H99Xl3jVRSjAn3ZUsES6LAaKVh8jaMO6R2gnpDQ0u7fQEL2ZV07fqLxBk
QA3trFzfJsqYw2wSBAlyorxgGAule56447WxhK9AMPWwSCEQtuLSCuxv9GBBWEMdxiY4rTmoG2Ls
l+cTOzz4+kjATv/QIUUfMAte1tMscO+tmxSXbQkb5jF1XH6OQ9GZ2DLYRyLgxe4Dqh7fpBkCfAde
1pqL0Rt/HML2/vUrV3HYwLPkIbqmfCiQra9YgRkVAtVNz36ke0xpw+O7fWy9Qo2z+LGZMYH8e7R5
g8R+zA0/ZLeAiHX5hlKmT0RPXdvwUB7X/QjcOhEYHai55NK/urNjgPjsWgt9myFfiUu8ojE/QWW1
d3AqtyKoPjG1L3GL4UaNsD2nE/jpCrIrOGwBsZOUNINExwGBa6LfM4vsLGnDj9s6rpwki17hlNZz
ahEr3vvSj1SWe5iOdN6RV84+jUQJwl52bVfIrXajKrXVxRLpQVNAhn5kZwAOvJRuVb8vtjrOjiKM
3DLqZMcF7bzK19BwS91PK6zRm6sCKV8OUyGV+KnOzCFPUGDhxFks2mmRJRga00+P1IwPIlfh3j90
xg7OpNdCyi3XMdazucBzuKB1K3N5mzc2D5DXusj61sBW1iHLXV6osEiz00P3D9QdyHJhfejiP2hc
165olvWhUYaIs6sOGpeFPnXgWjMPf8of6K9sMm9KFmiCt4nGH+kGbM35uLchR271oaIjGdiGY301
rx+4L7x5qzXL7qHkajgoGM8rw9q6aK2lIYz2ObQdW6a9N32WO62Yv1QCQHVvXgGJJehSMyTZdB2g
cW1vpbQohEbRkIx5eHDD8YLmhGmSkV7k8FJLf0lI49rQaVnFoXKP6BMPvkGIarGDwRm+bLpJjYWK
xqpXUwt1sh2BTJM57kOYMOc9AJ2NmoZOMuzHSeWy3gp2cyHln2b0JjoT28bIcCjTtEDP7fpGpjzI
Mb6DL4G/G/FYqx7QTf2nzmceVCCY+MW21eXHoaa41DoouiePpcyPQqc7D2n2MEtieFFSy7CBZN0+
CubLFv/1c42ED5cZ+5wh833Xr/bj1OBiAEL9uKme4w5bwZQbeoFKBO/PQvwWdrVNIM3sCIHr+8iy
QRcPYdL69suh4CeAgiZt+fc80tSQ9xchxVTuWKVlnrA9RXc56b/DiHoY3KsbUOrPz+Pe5r7HtyeE
aChcvTVmFQKKn0V3Zh5kbfC/DxOp8AUci2dm+Au8WPOpF55a51AS9vqc7Yd/VviOcyE/fpVQa1bN
dj7Zryi5+hZzOtSuZNzdoGmVvG2Tze3GqqzJQwNuRlXRMtov+vSGw6zy+ZoDZjjFfozGmLPqzAyP
/c4fwB7yIYa79ITXVasdhaOdRexZW6HFpjM7xppWZWl4M6Ys7jtMYorMgcFTo/5Mk0+833C3hyn5
URfWNIw+9zM1btsImuvLw6TZqxkwIX32Cyji9mzZPkPdbgFJ8AG52+HJnJajTc0FptEUe/8FfvwU
r5TfyR0PIf08GOfSEeN92pe20J8tBO52exOfQwgpuBOkmWOM+0AhZyLNxcZDr3OrTC4R0bMR3rDW
ad0vsgxeCoRR+MeUx8JEvaavpD7y+sdREjCAcM9/M80VZPFDc+p9MmBFFp6fAX3aiVx97JgbfFua
2FiGmRiXpOtZZ/cOWf+8KAoJWZ7BRCI6sq9i0SSxuSV/5cqUA8En3UkPUaqevDv2+X+SRpGoGs77
YDjmWK3qcXRp7/RW8BKt/zxF726AtYHbEzj0r20Xc+me9j8eR1KdKncbfa0Rmpz4WCoTec6d0gG0
zaPxFcIFSeat8FuuloGrIV/A/a29is8aY2zIr0s/kf4SN4rorp+9HSc+17zKc95T+zzDotEoAgE/
BSSx6X95RVn5gz/IAFfhDyG+qtIzXBJgVx2nuQnTQPtuFmox5oIoTCKQchGgZDvv4GitiAy7cc0+
tzuVWLFR02bU+HX8c71BenDyaCz1q/8ThEnCBLJBc7A0aRNs8sddTRRStuRYtKTKl4IgeZKf4l5i
Fuc62DOX6oAb8BbxveGt2wgeyNSNm38s18eCT4+HMb0BCs92TLlKoPKgqD2S/3bEG4JDCJywdSpM
g6IMj1neaSIrqpAKp1FvbqRIH5Wml2rIrhDkTc1Aw8wGxiwifHBftjiqJraC1F/Nq/1/JaxOwI8o
lVK6XSvAqEsnobXiRT3b+gYO+sOcgZYYaj6+bqyfqnYvm+S9IJ6XesGn3t+brti1OwEABf/oI+id
byjEchJs783f5LGsl6noKEahgdvqX6M8ctiLfqIBrW7CrGk3ivxTFmROuHQYPBytgGmaXlnhj7Lz
Y0PzpgOGU7hteCmto2mePdjbN3mElBJDQUf9WaEHmM818DzhZGum1naXtlQO40ECS1Vf29PtlCx9
efv239legwYV0gxNFOCXKIxzjjE95ZhAuZwSvr0lQmkw98XP8gHV/6Al+XihSYnU7NqyAWjD69bV
DQd763lyLYUQ/C0gRfufHvf1p3m8MiGFp6vMBYJHeZ1FNfjXEXeDoQzlHoXSY0XDeGlONX1HNBb0
GsEgIYa58AlnlWrGTTdj3WTBtld2aqZBcZ8OWvpmRiI20Y7Ssh7oNv3+YD3ehesIU8flRvddxxUp
fk0OuCKr1nKYqyg1FdEZcIOxGgn/6mtSm0bmKBuomwIibzaXq8t9eh8qMLThEZSqotq2B4T6xDBM
KMuYQZRQKfm1l+/sYijc6AkWz/qDnECzeDHjIRkPhpRL6qmzaCX9buu/+dPLT5kaaPOzr/XVPRfn
f4ULb19Qug3DOvk15wh0C/pVT5FaPC7f3NvBPHK1qwns1apICjSwULQAJOMEFu184c0o+3mv3vHn
hYjQfxbzwl7JhvuLZ83ctUmIV+D3eI0mqjZYh/WxBYp4v6bS/zc88q57VtrQg/NSKDwIZi5ZS6mY
wOM34O7K5o5Be/D6alW5gVRANPdh7/XPq+F8lbw0mGDKhJ15Szc4tEzfNuez3zX0Mi0VEWLq7RGl
DvwmQ3RJLTvb/6i26qGfaOwxt+BJn658v4JzG0WnXy5qvDkC2l9gUPf8Kz+ZiUCMQkoUIgtzaEgB
Kc0rrm8SApdDouLf9FH+PSiRT8uBvdXNv4NmSu6ez/pTIPI6xfW0g4LbcKhF5NRZ+5ITqiA/652H
n2m3D/0MpxnjTVqGLz3HfSclUGXopYhdFEzBbq0hxpMUGS73v2xqRuLx99j/huE0tm7jBHQNapmL
QCOTLGJn3juZsDL7rU97fFAa4tk9FG03mpzQSWyg2h4RE2PU2ICaCCLq5FclNmS5eecl5nwA6EvW
oTsfrNgG2KwlgtRwZD6pZ3BaDSJs4SdoB7p7BXiarYwppKP1kyENKHuT9o1M4f5m7xWLTe9RRmUf
96wgLstZDto7+iZNlxip5cO35i/amXTV91GpFkXgoW8DdEbKiZWXKK95K3NnNra9miH7RnuNoK1H
8cfubB6XnwuVaw3D6PX7fPsYKVWgSEQpHFzEEVJmTWtaMx0bCnGaXhsk9Sm+pdBXmKJisRXlDwi/
V9GTPmrgzcuvtjUlW91Vse2pJse2aXlQ0C3UrtSFMd+J5RzT32l/YwhaWQEfVFNzted+o3HMXN+P
gn7PiF4F+RVQs8ZX1VbQP0Rcax22OUWbW4mjw17ys8vvKvElQbI1YbeqJmHkRDEw+5Zgvz7nELZD
U5awOdUTF1y9NVhUGVm+SdoWWxn2VxBcixaXqQzytl3r07b0V+3D16ImjkchEu+DVDkkVFbAsMkM
FHwrR56CcwDT9VtxVwpNXPNuYIIgd2dcITfH8usZoj3g3qOX7kFr/1Kh1iJ+gthtINqKjymZN5tm
3tgrbENm8YNxvPz8CeP9ZWUicsXjK1VhZlaGwE3whvDpId/5XjVDNvByhBfR+5ji0NSk9CxxmdUW
IqVBTlI2RCprGIvkd4vRdAcRT4Kx/l9HGAh4q8qQpNZzNBMKZmvyBGDhHuQc/ZIjVeBPGdz7IhJn
Sl5bseJ/rJVKPpbzKoxT9tyHbRDYhr0b4yKk+4rcrPDb2pEq/fGrNN8aUGXYdTgBlN+3lCMxSBuU
6WFFBmQGIws3mnBcs8nK33sbolMLRbAD0YRzaNWNSe7i6Y0NYPwPx7S3Cn68beOU0KPuU68s5la6
8VQwxPs9ZxKZKxWzLervc1GAGioInM3jEDePKnHDkwuLo1Y2wQ70O6LeEH7on8HfBVQrk6M2Ym+L
x2+nbHl82Gq7h2fT/JeCdidVMBy69OF8Vu6lfa2zHcUBuqc8RbGHdKKYLVRIl2W2YyOvYCZqm4DT
K2pauUT9fUeltjNLJvaLxNYkp7E8LF9l7Kv6u9IP1w3Z2SwIuz9iuCwxBtT+jsqsRbe5tikaWb6K
G/QJeYAVWb7vh+WN4l2XgpUPW3NT+DgAA0i/JmGy0rxmecW1sOJuSKnvyEAGwSo/V9j/jPCCLnC4
kDCTcB4IHI1DkbLOQEnr5fkHeANwjgWBehII3IQ33qTabN3XZIUyxuWpQGHnbgmY4gY+VTwo2QVw
kFiht/k9+9h7NYu9AvFAPhuHoAJtIP4bfYMYWCpkFJmmmnGqQji1aN1MtrJzbr2rAeRQFvBcwvpl
2kneNXFzZ05xwrrTHAuyRWWTYPAVZNuC5wwNGg6ZsCPAJek9+BuG2+Wgu9aUBHwrTmpor+GdWuuD
YWUKVDXOBKaum9516ea23SCCPCHnH6S1OAdxpYHz6/OAIuohf+rrb5VellzCian1U+Ndz579VStJ
avjQJKy68nPSvzz6TRDWs6PauC8vqJV0OZVulbMz1vKlqdBARE369ygy6z60rV7gOn2N2NEaXAaj
vs+QwvYpaQt0iMR4uy5+Ioc6X3ag0l/0MwIo6ulfoHp7jBMx4kcMDT045DxMPDYJWsWHKwk+dNkv
v8+hcEkChDZ9nqSbzby9PQCFKMZDmF30GcGxNQ2SI+jRuBiYIPl/KYmGoFPdPI/6TyjgsXEWKHoL
RIHV6vTdWUavXsobcDwfkR+yeFAKaRUKKKH/x9D8AABz1f52ddESeInkRZlmHc1BPNjH+xV+sAhb
OT4XfWXWZzM5dqLLmDDJG2nT6JIYKKGzMBAH4Vr9vOggwqCEGns5zCe24FF27Zm9fpvnFuOun4VE
J+kIq9f4e2kzkKH3Hsd83vrNH24/6ymbHCGGoJ3JC5mp5c/U/LeCzeS+euGzUqNt45UMDV7gsAfS
kGxrpt6KyrpfT300bzyb43btRfrNabCsAxA0Sj7rB+Qgc1LY3oq7r8pjJk6wz7pgp+jyEIl3YROo
6QrHjEl6YM4zE2bCKBrYnXaZguKTjp/QYvevn6ZUCrH26NHNHV0UC2vgAkRarCJ3xpWMZs7Ew40n
XJvTacOP1NW0skQA4CW+s9a8ThwPMlzrXaqPgjtPLyZW/P+jdQ43QhTOYz8nSGHGj4BjCS8E2Qqr
lZZ/PINNpuvwmOUAbc2XWsuynNlqnO8+LFw/JPF12nt85erliy19pTG6KB+1IjMj5n7OhTg9aA4e
78Bro+AQu1kHgbdX0gMGqLIOhKIEfCX+X5Ef/3WWI81GMtrIrflxpIsE/Ke227ebewTu0OEfHuqs
U+E5RQVYl6CYu0eRw/VfDBKZm2qyW/9YsTyTS/mS+vXyidQys4/jEkD+jZtrOm15CWER2HXn/cWp
+CdvGdWF2jd4m+2mWxmEClnzIx0c7jhza9JLoRWqt2Jv+zfCsXcvweeYN0lXhI0Jdza26v8jzykQ
AqHfpMaywSCenYld9JiM1m5yHbB2ckBzzA9Xhc2RS/PcOPWM0SJhj2MSKanUg2jYHPKLAQponQeJ
I09dmBx8PbEl1Y7ezWj3LL7FqQa6RnBuVIZhI3c1yABYCoUlaLOW9/nkAuEZpWvKop5EUCHy7LMm
qukY6Nh8+iRqQWqyea1gfdLE80cqSaaAv8Es0q1b7kJLMmdI6toR9nvPJmfPrSIVy31Qj2Z7uZKl
aEl+RmULpJTB8QrRyl5tqPv2iEQzJfaFBPeoXjCK1D+usCnPP1LYVlUXjXb9OKX0zeimw1dF4zuR
qmqlJfuX057NGeBX38eBJfO09XDK3aRgdIc8simsFUnpCcSpVXtsSxR7vqOpC1OPw/ZOPEWhpJis
s8r2OphkEW2CHKSr9JoJ3Czf/iTGgU3+Ck+SbhmTjAfTmSewhwdigUPOph8HIcx+9ck2esWVzZ36
3zeAIrBudJNGiD2CznSK6df+wikLxbzVLCR+WKzn2GxQPHgL5hSrV5UsXquajxNYl3cmXqBz2j8u
NmTASEsSsX0e89PyDULI39Rt5iqdsOHmF0lzfVlTW+qjgmJ9boRt1FeDCTsZmm5AmC8Snh8+5nzv
zG7XpCA+G+NCsfqXmXvjN2fibVKjKHNggAsvToq4TNbg2c0P3ZrC+Y3KFNp8i3YpImkqIwtil/ma
CLNC9Tu6rM2wBa9Bgo1ctQlaXFLpiuWDUkG2jSy75ctLCAHU3w5LPRp0u4mrFn8E5g3Gg/ZMs4gv
SLeFcn8b8JXEkQgNjBYqxT5xYxAjLAlk0wLEzlsLO4vzAO5VxZqVSt4uXYxO/oL86IqcyNljDZhZ
lzIx54r4JIZY/mb0IsUwPVpXC3TPjSCy6RWY0dnfuLC1Uiyd9D/44gEWUSE9oWfXcePJv7EibS+Q
Z3KBuCDPrSmidOGSQ4e0i6vywQ6q+37EaKdEKHSOJDaYr7l8MfZ85v1yVMPkZ4UNFiKB5B1u76pb
dWKa2hjhxg9UBX6jbTIIzsg4tV0nwQ7GZ0INl3IHify4gtmxr7XjphSOCqeJ1L/JJPuN0FUitE5k
LNtsPPMa+7PVaXfW3EwgeAgWQLgs/5Isb0r5I3oWC1/5t3tDR0jp7ngV9ANX245+Zkx2nNVS9Y2G
d4RMAvnONajhGZ4kDZ+5qxzM0NKxYmchTsCPR9c/jkKX1xQTeF6+28rU5nN8rGVWg9xRyfePk4+v
UDRUFSNkbeBRkwMb7VBHViFKvMYKVQBzLB9UbLrqNN3MuYiea6CrLi98UHGh2L9gdO8k8cCbaSyI
zfMsUjHZ3sULpiqow8o0brYO36EELVTcUty8958gJW7KTnX1kmykKIX8zsQMSi/81u/1MSZSt5Tj
U53aNeZMqKvD7QwDXeahQkxbltd2m4LblJQMuM8JmqO+FU0QTNY8mQD++qRcZbzmcUguR9UhQOPB
4TbpuiEj211RYgZBFY2L4WaDWfIrfumYKatiJpS0SIUJ4hx0MtpEdSxI/mE1YjXAdIptDtalqmBB
qMybPUkDyCnuIrNxU/jjnL9KBUTeHDLItyOLyCZwUDkBYACaEIufoX9ko/sU9SEnmZKvUh5PDatz
uUDF7DfckIujOxT2Sm6lPI3/6VaUaWZkUSJSuhzZY201/vJs5yzdsZM+AthAghJplGWmjNYcYglv
cQFQm08GeS+bQUhMF6Xt64LUOYpcQg1dKqvvN0AkT56vInxxyGwqqOhcn+lYen8CoctGbX/RLFOP
4KfKIm3+R2cOGra7XrSONDZMqgClhdL5kNv5/CShgOJU18myKkiIVIPFQ0Wc9sWlGqRkYhi05yTF
hncS6b6fJKezGG1B9cko2aM18jWs1M9tN7ciigzvLb6k8U18pbbZYm5uvyAxfHu8eZ9WaAoAgJ5l
sNXYX9vgHe+7LxXSVTWV9oruW+pN/4ZnJmyb0JLRoaw8d7psy81vDThNmfvzVpdwfrWVWeJK6nDv
hTHV0iuRDHoNahAyaRU+lYR4k/tTNXvQcTk+bpnv83EZ5AsoMf1CKPDOw5vqqKzMzIHoJ25LeHjq
4DfZ+1bfWyvpmqlKHaY9WZNoeo/dsFkvVN/ZZyC9kkRxYDH1aS5CbxsuTFsHDFh3uC596ISWJh85
5vMRPTcMeYqpLc7X1uReD8xb58cVlpN44xUvSt5TqSgN9OkFNEcE9cy9AN4rU0Egffh8r4FIsmPM
j6tNd1ZQPlj4lUXmyqbQ1h/5KyjOmtXqAEAlXEUHsC9aM6NdAsuWMAkU7VIC0uZ5nQrM4VkEPJbr
AXmsbZXM4O5pYobEFlP/ts4iMUM8RhZCX0jVralRxH7+AdO+IehuUqtoelQQCGpOHyUFgfYcPDbY
UqJf3nkvTt5MDIpLhCGKJmEIx5BRphfGpxQEOZtLZ7R5DLlND0AhhzW2LUooKxSgMADjyoBH74xB
3VOO9cpjTFugh38RuiQjsKZ9dsNzM3zkY5s/NM1WHceCj1rthXHKmdmBDe/1HQcDS+lPmWVbThnI
ziVpUlk/hOU8eXqHi1kDzDO6McqxrfNDMnDp8BLzoQkX2Sa1cflvNctVyGsCVYWXdJmgKU+tzupP
9bE08el7AjeTP5IZviHyDnsJt/ylKT2J4BP1MhWshtsA6zNrY0BhZtYVUCwzuHSWh/fkJMOt8Xju
v522JouU/ITmvrcvzCo3EFJ8IAzI7284oKbfeeq2gEpDkylMMdGmvf48e8ck+oDzM1cRgc1/mLKD
xC26kuskC7yJgIzIbOblDuf3qNuJt8zjyeyVD8S+FnzazedDsZFMVUjaazgHxMGii/JqIuCIMT2A
MKfy8jJJTmsIFJU2xFiO+gMBC++9np6FnSThhxzo18m+nbprmS8FHLUlScXm1YsKUWaWpy123EMF
xMBb265oDvo/xmH/5zgs7R0yxKkicc42e0KOTHdutlGXBfi1VWayNQHUqQYwBu8rHQqz7aV+pTlP
4rJbXNqyGd1OAHIQc66c/MMLMo3FU+BlU0oKQJ/2GzpOImlK+i8s5WLtyIR7cLdbz8dxqjm/8Fgn
7Qa+eS334qaT5HFNOH1qQultIIxLDTuSN6l+Ai9LSKgx4+KFFRwIkgM++1zlTC3ojNYToBxoasKm
XneZrh4Nx4rNFzqGg2ts7uTocpS9KtX8egrel5gFwxeKuSlvz/Mpi07zP0FkoouQbsiS2AqQDeiQ
gTOeDLIyKtU/tyxNysME9Oj5Qg3LsS0v9Y6VIAX4B8uHG6LtI1Q0lCcZX2p/MZKl0WmaaH8JeapQ
clRO7k8D7rGq3Sa+GNr7RldIGrqT4oB+UhcgOCNGoeGMbccv7UFzLNsFGMBBYCaStw8mL2CU3+kF
72vbdHYdSyyIc++KZYphS360v7bBnPbTb7CtvhqL+Qb4cVzYVDRU0UkbUZmy+dkblfUQ9ZLWmS3K
ySIdnSpad0ZlscuWKOhwx5QGa1LMrxknkAvbjzSL4AHwBqzUxAJ3MNWhU+WHnQMJDQo47V2sy91a
6vANEzS+7I1IVKuGHN8YGd541Sg6I0x/hlu8DFg15pFrI4lvZPHp/BRvsUJjWC/gT+yW3jeXgloD
v/bXV7K6u+nELOK6J/b1PqiFhZyX+j6sGshjb3B/mgzNxqqs7QxqfBZCcMg8358IsxYYtCeOwGDu
FEOGjuplOhEfTvVtw0Gh5AEVcFmK837PeGb/7cDdPY7+bpeKV93Ekv4KdrWfOUidP1Gb7UQtPX98
evcab9P2gir6Io3rqac9ngE/K3jTT/DxjcBFviMhksWMyy7WgKFff3hBPzb3BkJ8zhcg5hCEOSGI
r8olgmY7Uni9/uA1QtSLbPL8ufAIt9qhrAnmnIcsFrYkzGj7+so1gUaVIlclb553u6qMFrJ6I8Pv
SYMKCzcJGI27l40avAk843ufnyedLAQuye3O7jgUGwIpwxAUtphowoxZQQqyPiccoEEfXEJp39+6
RMUpGuGVafYNkyLUBFl51rHYa4fcjAvhX+hedd0qdCnx0yNK4tZ4DQnv5OJvFL/3/ePRYaGkqELE
/OUD/LzdoRl2PeXOXXsB0er0fLOIIsskggMFSIu1C9MnIg0D0YUSTFnGzzsCpSTYBIri7qF/O0OX
DKBIG8OxwQKjvisI8O0XcL+l0ocCp2SNT8L1dYOjzx130bfGAoTRJPxZNkParPGUCYJpixn2XQ/g
hvw8qxpdgNNbDu/Jj4nYPfVykJV/K++GR1sQIGB01HLXLm+8TbUFJX+j20VI1GYLjI3Ias4tXcHb
8+Ar1UhJJ2Z3uIx3JtISNM2RMA2oRiZuWTYl98xe26iVpvpO0O8ERBj2g7RjU0MFqdhU0Ozisp/e
+fV0WEgMoeS2aTvbQLrHJv0Ciw+pHpPLdbyKe46P4WyNNdmCEXXhmpGpbq2GiYRoiklwpWsI1S2L
Ta6YYCA8jLwT9ILzy/bJnoV5knoB/4bdI9U1DyBEMoS5nnON/hVTHKHgwQjuIyzrnKDtjcLsmIaD
CL7WIBNeTZCKqP2+kAY9I1d644muFGxlEpvtvKHnFhJjue5aBSuvv7vVZxUV2E5nqPVanDBlYFI3
it0TrJtVvx1F0dEb4E4rAxw1SeKhCmwbRGFWCK53QF/QUwDZoy+SEF6KqDA3f6zv0dvPhUtBK/gX
MjoV+7a4A50hnOyL6re2QmUm8PvP+Rjvs70oFC4ssBYqhszsR71LQAPgJ7dnL+p093tV76vX53B5
MbAa9k1VGRjxLDLLDGxKm7RWH08lXciUihKQRR/ZeNK2MFscFId1izhqZ92Efl4km2DR7vB5gnK9
nuJE5Nd+o+jJQ/nvGZkA1w+Iw/cjsj1tLK/nJIgOeQz7BLh+3FYHewrKIUe1m0I5t0S+Zoc04Zwb
fkWpeYXpVpLmzac2SM7LvRNgL+CnspMcK0tg+WadbjUtf6OTTdLVxwrdTTY+JcCesxLJ2V4XYDa+
Hm5VYvxIERlAdxHVtcVB8GcXxHf6mnb9aTbg2QAbHG9OwTkfbBRUJRtksdtk/SzSXm4vpuCIKVyu
MvwoGtTkczdvTL9TtRTpJXjgRa9HIrxwqclIm4aYZMZu/OtvrRQ4eeicYcyVpT7XQQD1Of4vDiXi
zZYBayc05nFQQaG5ekyS/cRKYAIoPcQnFPzOZRTbH7gjJjICUC2tud5LJwb3fyY+tOmIsuCKiJAG
i3cA+FJ/DlsJiQoew7QxQCP6Vf1/F3IH2tG4GrZi4ATOX1aXcunajgKRRilsCfxgy9QuDo81NNaj
qaT81hAPhuiiezWCK63fP/UoivWUh5JFf459O8X81Z0pwLzePdM1w4knVh9OaB+7H0/HST+klGM8
GGtEWW+argEW4L5CQIfvchIZKsrGVxDdvvRtZgFj8azSy6gpioJAw1knkn2TY9EPKiVp8boKCwdW
Qei3t/a/xbVZ/t9SNDWGmJJdCPTjQzIe58JeRR+IrgebzElFyKBDNTzIO5hERox4T9KNotjMXJXf
ohLp4ZTV16PWNntOCg7AkOa/xSCleM3CsQDDydERA3LnjWqmjnKRMgJprJP0ICS6r68IBReomhxA
vwlHWXz5jh7kAh9roNFU0J5EBFXtAhZ7H9hINW+WA93uxQICcGXL/U8OsOz2jgejbJePFOJ66BUF
07sDBKoTwFr8Y4IUdj2/t92Msd5SwJ9JPLUTiRTiMo0juH5758wjclRTMdVMFhfKnyytSQw3n/0y
eOWWW2ZajG7m5sS7gTyx4S1xPVuSLhAzr7uO0iJuVh7pYlHVCZePJ6nismDmJf+ivydhOLdETtgq
J0vRvI2AaKB0qyOEWJc7kT2kzIPI3vdRXMt5VBCqpAf8UEeq494Fkj7/UqJe6OsXAUd8M1FMDLfM
zOlreHVS+/IMgE+pxoJf1X8cDAiMFm+mKOyBK/W4X1x1/nXYF4i7S5e00cK7m208ZzDq7dQ37H2v
ThLE4Hr0hZi0bqr8lJCSnQI0RrfYn6lZTj2agVb9BvQ/kRnp4yhSnF48iEnkKJTqj9JIU/xiwRZs
l9H8n+xpQyKSLrHo8Htj9/y6pjQukUjuINLzp2/+myBOTJ+4b8rhu3vjQn8mJaKSpGKasWBMV03B
BAv3O5dRD/BS/La+O2AME1HmCWlvS+vavo90sZ3n/LGjzg2FhhOCOOodMnxarzHrG9TYBNH622QB
uWKJefzu739DYLJBiIyv5Eucbyh57q5HVM8MitupCidetfVHuntVT9xngnG+EO0OQHTc2laLAkQp
M90H47YG97STQTz3hTEd8Ukjht1AheV9b9uvK4n19G34g6snkwCTbRwubq1+dSPdmAqLVgZusXAL
Kq9HCadhk+u43J8ZM4+nv5QHIuUujaBxzfGcVG2mtYQqONUeQ+SGjqgPRe5P0jtDiWUSlSkf7odv
xNwYsHEaCzrjyMySdWW5qvgiiYCGV39N4hG9P04fpcQptCIpsW3hG/P97LykzWHEv/q95mkkDznS
li10MMg2d3XUOgqW7njQ4wguQ+xfvt9C6uVX9d6RdkoEo/Gjfuf3Z0ZmHQteWnC0carlOY2pJwtJ
hZ9YxPxODwvber40hbAq862HwOfx38zUhhKIQjiATNNfgoP5Oi1Ae5oPi6beDRzUbuSM17N4WhW5
jQ6iyIk850Ags4Xr9IYX6ZOaUDkUMqBoKhU7gps8lmXuZKfr1fL+NgoP8rtXsm3A8Tgl+kO1e0Rn
1JuKZmHOZGTqNJtxsJ9UmcyAEVuFCVRwQBomtRnJcN6/bgQe7CK+Zvw/IiCsQs3RxAAhfGUQzCyL
ykCWhSerc6QO8FPmF1HrbvGEOYAaapItTXEkVYiqDqVNAsIIpSK6XK5rsYFWeObCbVqreb9jEMr5
Tg5d0SmjtkB98+L0KdUXa6wb2eHoWyvwyUmYtNkV5XXdmTqjqnhCDfkYwq93cbHVcEKqmxv4uNTc
1TcqJdAXy2sbiXJ6H3cbRot/oLwsKGUDmVNE11ssW5ysH/zl7Axd79HQNmaUARkusrugEhZ8xWde
Esw3nX047qTk/EfZhIxombAO39TCGpvEZS+FNpzYNaPqPm+oA395rba9C52NbT6b65xs0SV7woHP
fGKBbUH2NWcLOaDKGaoyxmKNUyjI1R5tkeQd7yDTB0IHcYa4rFfi9qR0utk4yXvSEVBoglvqxl2j
Z+4ZVwu0QP+0/OsmMoVxbK2seil14nJ3QkCyauuuRERRQDhZznu8G/8oP3movbRXUB8xlkTRGMTq
MiyF5LqwXzotWtL9uQmALVGbbSXzfoZDKn8Y0cCovh2si5YYuS2zvJuHL7clqs77iDYpcfSnsyDz
6H4At3clSasz/snnaTfYtLHK5UVpR/8YmBmpoetzWEtMp9z8LmWS7ztj8s2PGepTAN8hg3sWrhm8
KE1MgH7Ym4tkmWMVoC/KAQd0ngMUnKpaq+aolKWSsloE1RouZn7gOv9iwRpdeW5Oxv+6w1fPJKLd
g1inZcUfQwbyLxhLRlDZizec8QjlJia9qn+tvWq76Szc1Zh1qpj6NW79I5+jQp4DIYWxKPjFpp3o
PVMX4Rnh8aWcmCPWebmHaSY2lU0tdpNeHAbqvJ4yvev1MNnGpIZ7Qcp6AvXpGJYNczhF8Oyx4Frf
Qrg1wKXvgvaHt107QGayBmC4KzebiRQGEzLq5UazsXw2PuayJlXL4l+pNjR0zNTGzwz13/e2+BeC
bMhhNvdBXAH/ufk2emJt1I9/RZLNELh7Mjt7DWxw7jeAOq/hMpPVwLPL9XB3yE3C7QLs39WhEwic
mmcG6KZdoqCONLF4+vmRSFTL0RMeGHetIwtaRuWoBLgQs5Crrmfog1Vv7hLZw062sHyljtaXxUcm
Nig73JOMM+F5ljxuv5XpAahnrEdrs62PnuxdfPya+jtrxfLwsN1pkxXjnU1J7xHV8rUwYnCV+use
Nlf4IQ3OpcXFBPD5BLzpOBUjc63QfrW4c+7FLf6PyS3kaq9uBvRtAIvJZxiyG0qe3sMPyP8oqa7H
8XJceibAC0ztunXke5LpxzGsKAERbEKfdqaj+hkVP/nXcg+Yar/G7u0R8+Hua3bUQKJa2DEU6SCt
8kZFwehr96yTiClnw7Bb8OrwnoIyv/32zxer0PRey47QYR6+DiHfDGOj7CL1MMizSbAWPo4boqeO
vAxDfqSoOy3FA0029abHz2tlUQ+PIlA9SCCGw7L8pM+WRL1jC6RlMrxzz2f93OTMMF6ccDWJCkmV
YUr8nLPYSCm27+dLUkZmzXArd4vvnU7ooktCb+Z1bOR2/22jbjvD38ZgvrSmVulfmQRBgab+ukP9
KI89WmA14wAGZbu/+NsRIK7oo3klZBX+nLF8XTXj4GWo5jpQ78qCb+/MUR/lrfZXs9EKeBmMH/to
O/4U7tGFTDOxBqmd+An+zHFQelNtVD+gOXa+oPlvGcpp6LsjXiR85hZojqcmUUJEHy/BLHng1K11
3nMT1aF12MWrV5nFhwOa1HMTFm1ga1vJ+PLnzRHjjNbxuR9MQtlpAsKKeiHEnnLDvbutNakc7xDd
q0z7OtR/dKEZi4oksFaO0MCSY6Mqv6MRkxlYvg4W0NVJaWwkD/sZzFXnwGaBdsHGkc6GzEVQbXdF
vvSeIeuMh9sDmDI76QuQPF5So9mJcDjEf1vO77bCGA838mgTeP/Z+PnagZJxuNG6g8uPb+S6aOri
rl17L42v2XUo2SU8OZE7wOGDsOTj6D/nX/5n1eR6T27uFInG7oEk2Tp3OMaOuc88z0BHBAXMA21v
gBfAFfwTprCSstARBZyGvm/jdE3/Ygbt5QgPJm1x7PyJu9tUdOmYyGc+dmhSriVeoMVxm1zwM89+
VLPRP53nJdyyXSgj+34bQQmPMCwBtRGNThuLBp9mKReRySPujSNjg1Yk9vLRiN9ypZgnKkmo89yn
Grh66M0QdrUqDUqJ7Pnhsv3NKwbhahiGqH95KvGPHnxiU1vYJGEGSvZWURnNr7uAozkQnBWN9gFC
zIJjhlETqRoiDqBT2OyrAsvLKNZMRHlQgERNWVTzptHoQSOlzGlwk8crcswQZqpof8Hm71K7gYJI
8cALx64gjbjj/D8SwDb5J2PJ4ekHrvZgNfJnvAYndBmKLaYDIpzG1IzHv58TzAObquEynQqq8/sR
8ns5TCLkZfjhwTBQaZzjmz5eU226KBCuwkGVPL/qBUTD+t4leu1nxlMJZX5rETuzjVoV7MB8MvNr
AjZvcGiFQ+QpmqoKoWJiHblhXJ/S8hNek6I1c/ES+2WlcKj5OrvIYJJzymtRQQGZcbBJ4rgLeur0
S2oNMB7G+G2gBcBZIGoTlHq9nJpcx4ykcJma4b+sejx5Jy7U+UQRAvLHmlFqD+oAksv2GC7pjXcO
xXEgVL0zWE0iAe/p14cohrt7Bnjt5UUuSfIvckOLh/rbGWFoP7soESzksfOhcYWAmYhz9AdrZBAS
ja4bUjL8Mm1wnnpxVwxCI1lRSjLJZ5chmd9tkzsZGo5kRgmVj4KIQTbtZSTWpmqIbcPBZcSRbSLk
5mRadrpF/C8W11lqaal7T0UGjQhhURRoMJRuUqc4rdfSA2LGDkLKK5I/a1rUnGfQDlgYb7Z8l2OM
jk5eaDs+5AMQIGaOWJ1uUHGwvBGwRZ23Cyyg7gmul/mS0NMzg+e/cSfuwE87iSg/uUHO0dbKuPYm
OQAfIQqQaRLHf3b9QB/hJLzz9H9joL9k839iVZspXlIakyclb8m0pLEkMNb347DEF+7QZlgeGBSE
7hZr2wG0MswoPSIz8yo2bvzwa9t8lwKhaJZx520OzZzLOa9pdxxrPGeRYkrHmQgd4HvaSawbdAmQ
X1KGXgm7+vhNw8NjxoMZ4ouOiQwz+rpn8fXvJzecmnb4p4ZxIdEOnG0aUAF6XBJs5RPqMxu02dG1
TY4iz5geR84LktkJeIxtCcQc30CeI4NEKPxCCfEwfw81AsgmjJ+zAehM/iOzHzffDvQpbwIRKNVw
K6X0UT8C+dR7h7G+LjAw8pIwwogKDAOwHvZtZGTus9u1UBxeEjG73lHvaTTTkH6awKquhToKMG1d
C2vbG657kKalnaw4Vu/gZ/bgv+jwmQEqXbAcoTR4Papt3XJGFjtk9qo+yVsTa0NZt+/aRtyrMkuV
tL8YGmqonmKYEf/2yoEE+fykF0vGwrG4M2eV06gDATwjMYkL46/kPChxdi149GpDwO3Yu5FKMROL
99pG8E35ndMda2bW9q5VgUkwwaUjhetXQTgwHIMNGHieQuFr7i8AXI0Wni3ikK0AY3AWk2tu2MTs
tkfaqQzHMMATb8KL7C6Z+iKCi8DprwwgwuKzW3JM47M4PUIKiEVTtZLZSGzgoK2g8K5daFG9yTJG
r3otRwa/lLbkdPYxQcjrV8QOtvv5cMetX0SjF6Hvn+/jFiBLi7YnVgROcbrIeYFy2gIQsiFuEaX+
xeVAyballifFnxg0Z+OqzH5GIv7ety2lbSp9hYfktKqpnEede+Jf0OInjK60DkSxTN0Yauvnh1Uk
nbLUHVB2iYDobCcofQ4NJe/EaOk0u8mKHvIoPrcI+uTaUmwdtD8ZX4NX65AF6yvc5pfGHkoBXlJq
2zrN7tXVh+VNBAi5BVcqwHrba12Hgv9NHJO8nzdq3lzAtPfZEzSDjEgfrbfZ4Tt9yjGVeFlMZoTt
qldHUL3HkzK7oPt4j+53Tj7rnHbuxCnbOZKkobsn+mWW8WaPY8RH04XsPUhI1FuqUOD5v42iLL0d
RM7eloit4LGEN9kiXVYYKRCOO6GrS3lOPd5Xz8N8a6pYivItinsQSvcvCs72Ye7DRt6L/EFrrdQB
SXmcFjsMfgV1Jpk+A3b6rWgVzX/jAVnXt/IexzULY4IjJrGk9XlHJ3Q1JKFqr8UZigtM8lH1RIFi
QEtkIOFK5btH9xO97GqzAL1ujTJgztK2KSUtIQg3wpuQJkAI38WzC4vvGQTfxU1UAMgEePBi2+87
aUXwE/dhubkIjBEaFA2lYslNhLZ3lT3fWZHuBJOOrDqX9XfsrGt9WRx69EzGQlWfqehdKuQNb4HU
0PIHWftHzpnQ1JBk+YwnVP6I7LSJ/B4U9ERDZIsU+k44KdCSws3SV30Bn7fpIplnI79Zih+xfdsN
RA+OEbrUWcWJNmftiOvwkvU9wqKO9cNSNKyiERlVsQE2PkUaZAogOtDzSLixjvjQbz9j81kshESd
jAhiCoOLX7IH7X8K/QRhzXdCGnY7Sv1QWD0FWjz8sNNR0y/Dj65BapavIENEH8Kk0TlSofECBO10
Kw5rFb8NeD4N9SKdaTXa9XEBGhS/+0YvLuwR3NBwrTxUNq0fwh4MqqSYXphvNfmgJswljF94lfYA
3HqW6uFfbBrbqTE8XgCVV96YUSJrTp/69qQHoZeoLEIOzCgj9NH9F1vaNe0VA0SV45ZXEFHC1CAJ
6W1pcCJi7OkZ8ya93/ADGH8tROSI8/Y1HzAw1jEkbfgs6cneLgVwp3RDPtbERwMr6ozPhSJ3ZW1X
RjUO+AnX5CwlFvdZcQx9uj6+uL+IIuOW4tZy48hcvYBls4mqvxFUdXRi6lJTIcUY/ZlAugcjYqiO
s2ctCq54EZNvlloBxQVU9Bh6On9XsWZ1vK6UaNGtMiRURrYbncdI/HE2VbOQA1Ey2voVevb3YEmo
l+aEm9G0vz5pPaqXRH9o1aP5U8A0OtxRckVFOnm/wSnjY1Qx+qYBeAri3Alw6TIql+4qOWGML21y
IniY2uLhw96cFZdoGZim4LW1D4ioG/GdbaXk2HkrDCMJTlPaRNOawFkrIPVsHqO7DNyIZZ2vKzT9
+/enfMXtxnuldmqAok8KAICR77nlTClD7SYxUi/KqvGgH3kG+eiK3qVHV/XERVdD6sYc0WGVidcf
HZ4Xbnb+DJvJ1gx47adrYX/ZnmaxG2au68LnT317QEmj/waj6yq51bNPe6VcnktdmU8JFkszHqzn
UBLxcqxo9jZMMZHQfIDproZG5Vw6JLndOPzzo5apmAOb/ZZ9fO4fD8LcLQw8rPSyvpcDQgi/yjnb
QPO8xTPA8qLoGgN3o5+KZl6+/5ysfgnzjx9Kv6pKtNCX4sd9bHM9h46Znr6yHobBW/pDaAAn8aiD
do6o9mM/GTrWNgyNxAV6CWE+tkBr+gFTf/Iu47m0x/ieQNTvy51yTa7MYAGWfSUEV01oAU415ROS
H/c3MjJzobPtl3mzQHhDjriMnNqJrUeVZeaQkB2rZRAP9bmhbOW8A4Vw7u0ytRYW6akszjyIjX2T
YT0UshL96zjKLw7i8llJXzjsgxxzYL2CtjtlhOH+8SvdpADxwSdaMOa2m0dW1nhWYGXhog9CrYip
AOnlnAZbY7vh1dzagjPSdVvZaa5w9ZmuKKikrU4M97W2gWpScWNiK092I5Gwz4MD2tCneL8EFeLo
+Yyjm5Ye3E5AjUOPUFdNMzS136P7/FUQxFO/ShoRlejcGKUVRfhNqnCYxCVL7uCYFQ0VgYTGlt4D
Xw3GG9y+QBISeHGNDP0i2ickn3vaHC6JGuOE0rfL8jSauS7FYAPCcFn4S73XVoYO4/XqrEPX6MbF
NmGw+1eiWDvBa5zJIwdvRXuHg1YAKw3OSJXw+O+429fQdU1uWwYfw/wVlY1OSiync9On2Z48y8Lv
H5CSbQ1SiL2mfpBTGgv3OVv6FaxrHK4VRRWSVoGIGLqJp+hFeb9f7LIDZ+WLaHivPu1GIA4ilnH9
prFK7u7piUVs03noXTWP5Dhj+q8YWuMU9hXuZ0MdF9AlRr8VfxnplwHVMaKdp7fn0ejby/K3xryF
9nue+iRfTStrFzP2Qdoui5KJp1pGF+4sTQX/R3vc8RVM4oIsAp/F4nycS7+dZOC80cB5rg1P8uW8
6Jdz47sT+Zb33lMTNyetd2z5t6Q6Wd/0agSmdqJG+hh3LhSIMElbypzohexrQy588egtiW+59alN
y5IIATYiet4/pD8j3Phfp0fgB/V3AKi3fBn+Trl3WOv3YAYziRHJ1F0dAndWdXlWZwGeGJwYXn6T
6EA8xVPWK/I+UAOC+FjgvjI1dTHjrD+FWFU+Z3uL/SXUD1PlN+HIfZgOP+vmZrP8ARP+bKeu9Y7m
u6Ix5gyrS4h4b5Cz03RuZoNS/pGd885YylDPPM9TypmPEELvhM9dP9Ki0EciPxf8o5dbDijD2kDy
84damtX1lnaK8PTLHxICzpuR1sb1PSnEGhBWt3TOpo+atXDI35H7+H4D1Qa66MWkHgHW9HUAtuB4
nDoHNLkmv+4XYOBy2WmE7o+0cEI6l4uWh/GUWYg9ZW+pnkW7LtpEnt1JacyeOrpixIoo8pSvzAN7
TI2X5L4GjDH6R8lxqyiV3lADVQZyKJtucI9VRZkaJ0THuBIk3t/uLsy0KTv/piAlf7O24x8O0Nh9
ySURSYyp4CsKLX2ZC/anPeOnKbFycQqE8OnAE9we1fKZAf5Gln5OnRO9L3Bvz/8mpLcK/UljBEyU
9t2j0mqnP3rK0U7RlzdF5PoPwF3u8guzn8BS/lAv2hp47w2a91fgsH5LmXbCM5EV1iJuH1l1iEw+
pQpysrA9Mqe0blnyLoOCkFgzhqg+ViVUIzF+frcsX7IxjxqDA3wPXxmKd0r/9F3fhV9nG5yqLiP2
iJ/mfPayTLn7e6nG8XE/mtYc0P84aoXKdAsYmANJ+XLu9NxX07N2IBTMiPFjld5NTfTHfGtNAgr+
jxXneMO8ftHPx6mv2Ft6+kr5WyVOcjQxrWUGeulgjmKI++2SpoRsCdrWsNUlIzth4ayqchMeX9SP
d4j2HzI/Sqv6CuhHJw8CGQ1QTjdLpxcZ20X4/h9oZicjQpO2hBuIlX0joN1itZSxvUH+QaGNXVr5
e5e8+JYcwTlmuVSgkb/kupoXVM4wxFlbh+W1ibSrDxV5TkeRG3gxFM2Vio8pu2G+vZ4jp0KZRfgl
aSoRdNVzriaf29kAunfswNUIAA2Etv06kMhY5wTeZnv6C7XzCYw+IZlDejWhJ68QAaTrRfVz1x11
gpHvRvv77Is0XMErQfE7UF2rC1mI6fh3+Gm2Amv5UZYrF6mduXjTi0eP/ZKhKyd+y7y2NOJ3pwJF
ms8Qan3Q73WdbGDP4S2W7w+OKkF8WkzR2a1LwBhlGCqoYm8/yHYKdNnmdgS18ybwW/IzOjV8wffa
7lj1Nw0sCcCrPS0ZqIKao1gNi+JBpPuVeQ/zc7RgibDJJCVhw/LnxwoVcF9Vex0/FhkNcyYENSIC
cpjMUILX13jU8XjXWWhpQA04L5YYnDOeHwGORNhLzLvIFT5pTuMCaEbYxzX9GOsJBW3+hNTKNKce
1FVH4iAZQfjHjNr0OWSjk2F2Awh1Ozlu89sOEicBun9QlnkezoszguKEtclUZscGeDMa7cfBFEr5
tct4m4f89Qy0jeBq9KCaeTiOJcvmjZJQKfzR4tMNzjr82Y3fKG9C7q2bW9EDbUitU1t4sF+CUuBj
JuAVNpJRtRJMDCzKbtuwqyukDH9I7I2s3TtSFFoMxud4lxVEJEDFPa6/i55kMNOaV7MqYM7pbvYb
RvpqiQ8a2VyAyoTECEymFz0OSkNiOOKME/611N+Q3FkWt8WsuzE0Y20P46S9dn5+Ia62rKKA34Ul
UmeAKUoetpmxyV0dAif9Jb+g8HNozz+O9qFcHLJ5+ACpEpIxPXyRN2n/7lAQNg79WfaL8+4k8nS/
4OFww+F4OKWuQQEMNwzUoaO9kMv9zISOs85ysUeWRKMkAim9i+RGZZzEZGGcafatu61SVIbti11i
QyiA6TTF4rq/xR8SFtF1D0s7g6fMn5mOpF3sUWBDp+eo7vybEzuoxq2P/wsWbpxDn4+DP6y6ks2L
Kn7kE7urrYzeFB3uxi4DgPO5DcotbgSnE0RY2jbalFsuejFfD1dAaSwKWkdP+lHHyeTYV1W28DoV
nXSoSMkbCcU6Xj0BGXmVzS+MwqS7qb33LswD6ZZ/V7HZXNt6mcGNaOfELcLS94lvQmf82/pq4w0g
KnmPbLykiN2uHD+mrgK0XRFsIQ1Qj2fLo5oCCi9VMFzI2MMPhQ9Ms3tvBlncCchwY5c65ip4CJkp
gkHZNOXYU4mr7hrXkpJmEBujgkUl8Qf/U1wdrwa02BNJmQp0ztvQA4GlHF6wlGIy3iqh2Zvq5cgy
nGFy34agjOLu31lfGelbpFYL5L8TZ4oszXcrAR9jrbmaJHr6ffsK2efmbz7DiGLH84NlysUbJxS5
pORThw6011KVyVaL9dRcUkZ72i1+B4SkJq1YNy37VUBtZOJzrXYet/kBrMOEs67N1J3Mgbqoy/Cf
4ERVUVh8g+tgiSIEoQOcp/D3JkqX0IptZqH6bACGarVovqIY9TQSQ0saDpnePcCVL8KL4JxUcC0N
4jHp2mjjP1FvY6PYrsRa8I9x0AMWU3jDCJtSaapKi96zNzEzPuxutv9NeWzKBf/dd2pZxl7JTmKV
x07X+YIFxFRg659Y4dvzeb8s/fhTpQjJ/uvyMRb87tb4Uc8g3dH2UYgaO32rp6qjK8zPccilE4Mh
7TcJigO59TOxTAMGwABkxv5pwAuuLf6KTERByjMPMHCVBHsqtidXcYdaEbWRw73/F680jhy8ssyU
n/+eYgOc25znflYys5s7mnhc8oLVsEtTq5LT1ABMuP9HOvixfEDfxkS1ks9iOywzI1p1ymeegxnE
PnCoiMGgHD9YBubjXnOg4T04xn1+yDbvivweGaQN5nh2/ChF9gDc1AuRqE8m7kh/6pibsXGfx+ki
i6PSrab/PXsvnwpBES5I2az8ua/2JsUD/mtXdw9nf0+o4dvSBYud8PZkOYAnDswFxsRwRG+8Z2bX
fD3tdwy0fsXE4FZjX8hKBlLF0ShRElyWhhl42boLFRgm0MPpbkYZskD19hdJqkurElsCA2g9LUxA
yHO/J3QP2vKUDd8qLtQkwqx3pgXq6FvJ/OPGgjvjHV5OwURToK2i7VJ3sM9KqifgA6ol4dCqozEX
XfwPUZpu03vX3UZ6Jm87GUr364Q23vwNShg/8GILuVrqsCbSRvUUyqGZHU/0JCOBkI/LhzmUvCkE
Y3LujaYKC4Kg9o2yYaGTBCPnSg/5DTn6reQ40/E5Q+nf4P1iejce3iK0QmQNRjX10gqSQuKa0dxG
9/MtgzjMsmptMZVOIbENeiEoAZ6Ol1k5l0LkVVyWO18XDyIDUxdRM2E5Ail66x1NIUSRb0y2ln5M
DY/lqjK9fnB5uE9xPTrOrFujwFPq4QM58LkJt3kG9zHlxXi3V3JKS5iiScR26m23CDUeWWIyAZJW
IggBKHxGHTm55CStLTrTinTL9e4QzjRgaY4zlIBezWyPR77qEs1wzlKLCAmJyPKgCETupaRHpAlq
53COUXDxLq6cVLuOwdEPgHvLaJ31LN0MmSo1xJUeHZh9kxgUTtx3PfszRFUDJjq5frkgeWZVB8WZ
MGZ5F4NlBX6MdZQH6annljfsCgzlQWcyvRBi2hxizoF813dExWhaBTZ/XRu255tua5av2Y7OynIY
saJ8mw1MuPelxhNVCgZRl9ZSPMRAnfkVNRQ9R8+RAPyoV6LIc2GF0aP91G+7aJeGzOu6xXbuKUbD
S/eHW0LEGAu6uM0zsjSiNW0ZmlGR/uQIsplD+u3YhSkPOr5EQwMSQnwpEq6isz6J9yro6DAugdMP
ri6jY0rrGqS8NtxGjOmzaKxSy3AfVW24IvCp/bxfb313Wr8key7HueIb4N3i+xYKIOLVQjcVIwlR
PTwnVtgCpy/BrrGqrY16jgrHC4iNOGWDvgI9ZJb3I+lPd3hnMEUoFVVQGwG7SW4oDtOMwV7HViui
nzud9qMrjQ1R0diBsPNao4kiWsYMUZ9k30dwRRCG7M1XD5kq0tKbBEgCVa36PhWuzgKg6mKOjGom
v2LKZKFPjwLVVADx2WKT7wj8Zg5sdsR34pkQhjVVOlTN+BOVSf8s+Rz360g6aVmIPrRF9Ic0VQYp
+KZD+qVy/UvfXx59yWLh96OE6zZch0di3raFIJYNRSVltfGb2HO3r7qSsobqzxWd70sWjvY0Sw6W
e82DutNubpWOxttCl/ow7PO+y29Tg1VBelTMEU3TeahPzeQcid+ZMGi90jcIHh1zdHzIpaIv7ZmM
MWZCf0/Qs7S1fzsUJe+UWnrXolNiGIx3rJBNcQJ4w4vUebZoulLuqrh2mVHHlliBZTY+fGh5VwXh
P4k9AzRXGsXQua8PZ252fI27tOyFYXnruXyrd9rgtTSnSWqRMnrATjqh3TkCRjTYPU0s9hb43SWk
54Yg0ICgyCNFI7WdTIiTTbHZTwbJhU1bEfCOHRfHX3aKkNZkasTADnHIqiTsiqbtSDksUaMQK75+
Zy2LvjJJDBkfljWszr/hmI3U/9a2YQI0TsmKENUub+FCh2AStDlFvwFbMYaILGmQuGTSdAIJXxvd
/OQVJzx4jnNXFS/xtynwfphUznCvJOLACibs6avVEA8bZrU5V8lOSADmFN2xNCxRb4mrK/QohAEV
lHySnBGENS3MzOg01dqB+7PTt3J6X+wKpFCuT10HMGI8W70N5uk6oBS25cpy+02j+/lj94tRHMJ3
D/8sbsO95UqDZRoMS3vaiKuZa5GzP6FprVlYmNMzvYVzxNLETnVc/cj4zG6Jkd/OZGbAesci1DPi
23GmCfGbiQX1kVKAIJbJjsFkyss8oGGP2jm86lR7eEV+rZ5/+qgxZZ+LWS4dWEBFpIQGIBgc8ab9
katYwx997AI4nMFSrfSCi2h/ygwhORzy/BOrDJzn1vv8MygG3DpbN46pmuZDXGad/0yN8XMGc81w
w6Uswlf3bf+usRMT6967IRFkn5oxrBnkS2elhIDlTvrBAPOkR5nW1LPllg2maxsKBeQ4o8FO/hRf
jAkLlB62y6cqcjgw0LS3fanYxVzquOiRNGXdECyZzY8/SzjGEswHb4RCreoilNQ3c/8/Pl15Oe1V
y6Tc8eQqz4MMt6iTi9FeAONRPfoSzRdsD5sxEAgOq0Hpx5NWHzwdKtYG+ZmBlE96yyT7kawBPC08
M5AIuHqQZFhorBOFazkoPRgzlHSF/GCH8+Qhvw/QpfIqonqYUfdukFV6ZtHZDdXvmStJcWUGg3WN
O+iIOb1vy7fh6vhM5i3+kDbpHOByhY/LGSaVGIlPQKC7ZRVrYYYbd14v6QpKzY9Mf8i0xRIyI75K
FNqU06dS+RLkYFc9vw6BerCeHQ95FiWKrW7iuw5Noo4LbLKTIT1FqnlC8rsLmRhejrpzfFixoxNy
D8typjDIWRcxaprlbhkJFYapFliOGWNtvl9wlSkQgsVGQji3zAEveNbBf1EwN3zE/YosgrBPOclU
mmHi0/zaH2JW010z8h/4n1upvkGHwHbD8OKEk/K0kgzgeX/RKtpT00VfzSkvRsgbAqGODu4EEc7P
JfzvDfQrzXYD0au5WZCx6nB89eCAc69HJNPYr+gvBeWN4MxVReIimfiVJ/eOGTwWsMOT5tACvDYk
+MvsUdGQ5+dbebngg3jiInpX1CvDt6acL6JX5dpah6RcrU213fHw374EpQFkByFV5vm48H3/+xpg
hEsqA/8RZIxR7TrwsIrj5FpG1/JM4ikkAb9sznsV0G8v6EDcSnUkjVSV6FP4J3Kq49an6Rxj+YkN
2O2B4sWzq7DfAieFeQJ8FmFn/54T9G1byPwN3b02vz0McuVste5JmyhBi5ycMpKQZNWw0CMvXDaq
34S6gMqYH9LR5uFvncu4nH4oWeOYhvZSF/qPM6QpdkcW5vm7fbudpB9M/2EkgWxDJSQ9VVUT3BSU
nTenyw3D6AhKgiDnfRtpQ4Cx0oAzXaP2Gx5WNMgc0O4i60kzGqW7wvoLDTUAGCdg+BAxrf0rQrYh
BYrO4PcDTwfrVMWEK3XjNONM0FmHKtk9z7baEEXF/wIgiYdCCayWNrNpPDLjMd+rtYGSiSFs22Pw
EH75NzqRfPIq4QNuDOEd3UebjjhdbbTYoLuF3prOzlaSoes3nlq/1a1zKcLef0Qa7xYDr2kUFg28
eQ4mFdzHNANTTF0bNP77x2x20Js49OHNznRGCFOHn5N3GKQm9SdpDCpeAVnxny27g1iBz8Dpmcta
Ws+6QjkQQgn+Qo/EFLuXJDs3Q8lUtajENWpOz2TnJzGRk+8oWQ/jSQdm5z+ef4E9a0ci9u78msJi
913/meuv9TMFRkCWFp70IzIU33B1+TFi/2ZX+WfI8AnK9TXaE6iuyPRPmlOe0w5NwR+ADtgJoIJv
Oe3Tm7+sjcG9M7L9raMdQ5V032AgX4WBM6GZLwhoigIATfW/pWAYaoHTnCmSVmKtLeHxIJD/Rh3Q
2JezJJIrpL0wNqE0v1ig0nVPf9cmSY7upSy4ZRkC1B2myTYkA14HmrxCYXSE/puZB3MavDQnaTZG
1NQ5WuBxqLrRK3YvgNvYTjAT7bqaR3bott9y28Pv4hZA7QMnqiqc51IyLAhbiugVp2OOOirGvTmI
4zlXPUA1kPdB9rja2DaT9wz8ARmD2yOfQXkiOVJ7L+TUC2GrW3KVM2CX+hZ7MqZILLe5jGoAYAEo
iI+whOfC+pArVpsjWaxrEdyExu3hhix9rtySVecxikAOohnn3NgEVJYjlhnPBiUBd8JCQKsDIpt7
ApGZhpQAoGRoUq2VwbKwb3i7vi/HJlLPgK/rLiJ1kw2VaYJbjhccqp8rsQOWelpn8i7yJE2fVKlp
EoOdw9hTRhmsO6bKop+DE9/XmpWb9LXlMAuwfEbix6b08qdjcIGklmE+hF30VZr4IKBPE210wp9z
xV2R9G6w5I2Z5Ysj8NuFRN+WNlQQeIS/E+nJ2FhWr0A43p/JbuA+gwaNYa4BsEZr9xpcK5RAyNhC
x0WFH1aGDS3Wn3arLnCT7KiEnT0zQte/BAVoeQ/+yAtuoq65pyj1lKZzglUJKhosvQUqwGlEYENo
lE0ORvcVWQnK33ZPc+sKoD4lyuMWN7vk0RYCBoA0P2Wj2fOh//3XrR2+A3uX3kJirprX9C+5kX1D
p7hV/bRyCCaWFtB2XP316Rm5OsDjODMsBYA97VkyNAUDe2gIl1jYeFNXZBblnq7DV6zx4parh4lu
uYjV2sjXw9oH4pfjqNVL1NdIZqGUl5xkPAnhKy06ku//HMiv7tqmt+K9d/ffB5Q+gSHH/H2Bp+rG
o+eP0+pAhxhvnLd51DLVGTQvjeC0OCKXrZ2mcuqoDe5kKfBnQqtWJ4rtlmis6oNW9m8YL90L4/3P
/cpZFhM2lXKRt8lgL605XBvUq0Fzv69JaBca4Ilaz8dfuRO8NjuyYStrQ/BQbKKNH6ZNt5uGJZJV
7h+YrnPjuHtVc1oL+a0Lm5uAGUvaPdmSEknva1gJ3KqOq3UmdIoOTrR+ckpAorxjzq/QXWzZops5
TFixchSXc6OhXvqhPHsYZtEn9vNU2jzxjoHeLKt4sQQ+zmdjLycNEiIBNbPtZYl1nRJpFFQpO0BW
bkGVz4UJUT4EvkpvtqFfTSvy5I7gXcpH4XJz8CcnzVsaGVdsq71TaFr5N0Rnl4ZcFGeSSXiImzV4
HGHXLBIAsgp8nNc6mnZyH6OKZAvfz/VClEAnXkZUTHrFrH9Z+UYW5FdHRRlScCKrIAJnvUPrn8DK
FhtrIIGAu136IlixJ5gDEAuX98b45gHejiXdd1v5uV/5Yu8SCBDxOJW4eBylNjB7IDGcFj7BYU3X
z3R8MSrzpxRy9a+QyMfOTTQsocbcTviCLh19Ug2kcM35cEwTiGLEewGWMi6P1yc1CfnnOG5yigIL
NQBn/zmhsFktrQvZf8aqVpVZJfmqAslGUYZ8BtMOuauFB4m8sOCwJLc60f2SYdHbkTHAjzHdKjqe
anESNVmryi/OZ572oBs3fiVxIqugbaMiaAznNO+XwgYMidbgO3alXfDty6TCUMnAE2eetV3/ct3d
ozISYh6fq33qmVRew2U9jS4zMZ7gXf9H/FxulJDWOk6sK/ZnkwCbAcRtxYz17aTzVz0JicrxDm8x
lWHUZpvqIZKaT7bDATwF9EAHhQrB/aYNT3+sshALBxruNDXcJiPndu54Uee9HQ4Stwo0ImKlwqk1
Rw8weda7Kmkd/hmUShnoYUwRHsNVv3+L67M7iDuBVy2ANaagbwJJOERngebjzxecanaieQqBFf3Y
fGOLakqdxWKgDMPgHa8Jix8C+TkMt1L434lYPn0pOB8ti59AkI54zhQOLtn0+dFpFrtEBjwy1Ni0
AEpFAxVDn+01IzmDCeCDNKcZykY2TpD+LIOWm02teXoxDyxayUP3YMSWY8y6z6vrnNpJZxiERd2I
qlXSREATIHzKLMikpPIMnj2koaUCbrX8bEyJWtdKFgjmZ3DNGq8WIz4WNPcurVYodTRZlgCPSS8g
JZ0kVmgtpQ4zg0NhQ/XiIZqYq53f3USIXbeu2JeC1Hq5Q+pnd53Pl6EoBTthcSP5a6YwxiyAF1nX
YAo8EuNxdC315PqraXvGfOC47daqKa356rZ+3+ndKbvsUV3PnbCPFNMPcKTNz+WZ8iYu0Ge2p9bU
6TcEZsAv/afkierVKD97kFUMU3q8ckY33e72+n9xkaDUPDMbY52HPK1o3DuPuXJekdSA4RT+KUF4
qFKKbE3XaJk2vUVfwW7eZuqmAKPrqJkgFMTsxAMTtqjViczp/70mcVXIWY2+XvhR810PWkXRSUdg
KyB8R/CCnwc8ojWnK+xCZLxUrjw0fIRsThYui/prUbZA3cDi5W49sFcBNawXLoOQgv3FNXvjasF4
dhzp2ZXTo+UV9Fhkl9i9OjJs3rWTadDi0QTVFloy8Kr3DYqtp48yHY/JGeOGaUBXC4shQTrhoBON
RbRdpWSt76dB95Qk1QHGDsnxg5hi7X+3EPOk04oqtaW7bDpSvXKx1xk/d51khtFWYzEMdzVC3rE5
7Apz3WhphJEnXUhwfUiUQTMzQbl1RrHZdGBTLOzvkKyvN/oSwiviVn5f/jNDmu2rpj/Q/0VcrCvP
4+BxTPVHmqYDgHI6WpAvzW+/kz0JlTDTQqgAkfLCsvD5nJZhP+H7qwjy0AVTXe+sfkH5ptT2OlFA
eixe0yG4ep/Dp2+c0wvKxja62gE0uUzsZRi/quRr15VvgRTg3u4UmISThx7ZGAkM7BJr2kKw6Srw
04UkowZIzLU0RUJtyLTk7+p56uIGyn8A4N5GWNRyK8+LS+R8wPJXmFNi+p9lcDs9NyDG/5CokgUC
hb4cTZttdMTroZn7R+a9HbvX556VaJtgtROg0W6tEon/9d+Kk2KCmfzLTc7rorpM0iyFLliDgPw9
vdKe8FBkTCxH3Vz6VWht+NDn4A2pl+pNDyg0ybJhe1wNAKdy4mzeaHqrg1wtVUUIWGTas2YLQ2+K
nY+ptD8Kgdui2TyBnIgMKyhTshLw5zi/Q8dfbojnOWVHb4m32FUbffm4Hg2kdZDEVQ2/OoqaGM2d
SRwBpBT1vwlQXAXSWBVkKubGTqujnG9ysNkUKpvbkqxoBBqfdcvGTAd6nZpy7JGatufNo5Fdhdiy
CbjpeXm/gPVyCwi7OeehzkZRGfGyR9ILu3q5tT3M8ObXNfyuKIxONwoKkBv+xB0gXgQyBb8VMcie
gsTZSd0kuA4ZFQlW1kUZA890jX1lO43k9tp7Ku7xGOyblxWuQ4Tj3i8dcyVfAs/1K7CcaTOKgWQi
q+rYwvNM51j+HVpZ6A+PS2qML9w5M9dDp6T3OKlLsV5QTUY6GOt6AuYFtlcL9ksXVPBLfccWKsgM
kPL5ntN+T7glvfX7Yl0fNIGCkDcPfRctYQJrtbbZo8AEOH//YGPbpnyK7Yny+4W/DHxizaUEnkf5
WO2Dc2rYzC8jvkhk6zth7fy7vZek96KPXspPrIGFcM89NaLBdzeK4E3yQjyZEO1JJld7t1iQq5A4
9SXpsp4+h8Xjbapqkm3dAUe0xxbFCUebwQyuh+BDjOKH3TLp+GfUDgNLiiSJP7GovZBbjyh/vFnE
b9Z14QcE/6OeKbOI4HsrXTYyDcT0yL3agam00bZOji42AwzgdaH99n+kE4uMFQDIpMkvI5V/4d7i
Gg0RbYZi/06yf2nkgNbEDdHK4+OZPWpXZUtAxsCWnAkQhBV4B1huBTnKeSIa9FGopXwjwiMjlZ/F
K5t9LMjoD0A0u2SmHzLW27wwExF8fpt62ntKeaElIRAvxnapNDPEl+5EiYhEj4N8DNc4uDloRG1W
VVCOOoszjy71GbkWiJe8KrHS2pp/woXtmO6YaeKhmUcaEgqDF3tr7+kWt6uih1/zwnKibsCq7uEx
Ai8OVQAz/FJRyMNpJQiS5565ToVOxdFtWPshjwiuz/5rGgaW3bV0W9tFyLKUlMFN8kof7jcUaEwr
ZCZqr7ow/9l3Lb3TTFEb/KkE8zC3wECaO/v8W7WNPd5hf1+L4zhMdCb9pAK3vzlunAeKyMUzup6a
8CHPVRdlt12oZ44eqZDw8vj6c6ynlJ+bUidCIWaOde9Uh1PyagqQJtcRn3AzQ5isUxyw2LyM2gDx
jWVdjZTU+XD/0dHIAn+FasuOIoZzp6GSxHre6dj82QACzYFSivDcEtXD+lO5d3zXpf53ud4SGSgP
XwW9Pmaz+1/ZeC7L5hkbsB6AtoswFbYtVVNjWFw7C83LdxOu3FJc9AKLTLFg/69JNbAeA/WQkpbS
0pTuEIln1RhpeMy1DTYzsss1HgAjyXlImVUVLeKfr2oP1UGKNl72xirdzUpU3ttm2rrqXW8qJPdf
4wxuRb/aH4UMCOL3gyWr115n5AEqSXA4lTTYzFMhB3d0RVIn7fHx8I1hP2l4X+xujlIX1+W369LM
ZqrkaKqss8HxTFvogfD+gd74B2Ofcin4QnBQu9ctvmn2JZLS6Xe4DArBzyBQlxqlXBkEJdadnUEJ
EZrG/VCBUQRNBybDEMtSkQA/syBhvTMftnBQ7z8VUy/LhDKWplqdLU+K758Yqo+8vcSXuIBikoHr
Y0bqVSN5GmGcVzqbqfBL+KSnWJVBQET2YjC/JlRxJIizh/shze0gotQGkaJJv1M3uJRGwniS0Eu6
/3hIE5j8mDHVi1y4P7H6IyvOPGFaEm6uX3Dcx9GGqYJgkBMB42azforlOFILJNXWyJaWsjYdp3uY
rX75K9oX+Gz0XofxRMHobQnt14gkjILRdaipxe/yBmlsfAwZm7udrUlCLm3A4cCHCoi8ePiN0GW6
EFJI1lqUty6kyJB5nytaA7vrjKGrf3ljmDBWVXyqkas2QdtMkew+Xe3+LDv5ds8fYC12BtUUA685
C9Up9+BE/x1LJyLk32uFAN1Z++4Wpil/4UZwih0OUGXkvAKAG3OXblMhuLDXLQ7gJSHG3YxUfK6W
aF06q83l0rRtVUR0axUhySDl8Sj0BZFaz4/VfdWeZc1dyadC5fq6/CD+Tm38BYgbLjbYcuavK00D
+UUGc0/f2WNA/9UQXFvhXU6e0oH0rIsfWICksVrUT4YHiBs7WO5LQ87LL9vPmgs+cu/Hld0LF5ai
BvJdaDxrW+z8NJ3WNRdpjOtYkLtIAsuYaKEQREcKdP2WkQCFse6MjjAYYq/UcBEwyZn1ytvornLa
A1CniHqH10Mny51MX623YVGh1fi7J7t6dgJJAGrmUi03RCTHZLx08mlIsLetXK3jqvyyNWoE8ngr
tk6lhGdie0Xha3BpFowteskF8JdqksyqVTuQ/vWZ92mmqv+Y67oPHLg4IW5Nymq/vHDmlwXe0xAP
m2ZsggrGF9ReKyKZhwRtYxdamxAb1qhRt8ZDd5ggTENXMG37FKbOLrXQy5jLp2tU9o1sDy3W9nR5
d/zx0doXpD84JntReMPDkqULKfBY4oy44pV89jmsfckvNFUdKm1Hp+27mSUix6aS45XZWpAW5tRO
3c64iPIpefiv2AgmAasVEidKB95c4rTQwSVxQVGbVSkDp/Mo6k8hsHV+iqeoGxBNMTTJCy96yGAb
UJlYXMFOYKvtNxTac7LJlkauqKJ3cHHCfYIERXFc6tajeDDyApVI/53uAplxRaVOs1gyfhI1gPnQ
0/nyJ+JQC3nEwoBDjnRvEeSYMseN3ebRY5YVnkUwIzF9Pn2DKSK3s6BGuY+PwulFSnwUAy2ngpA4
WIVi3CW2K6681XVjUdQqJH2SjiuLTxy+Yr9tp2Xlzr4onxWI0VDaRtGTknxz2zrp2OknRTwOkdFQ
bUWRZMiGIqIsR1vO8IZ3ia9Suf79OjI6Ey4ZLmgPT+b1aIGUtIYvYwhIBEnBdJzsjxcOji/H4RaI
UxaAIxCOEUfbTsvTABkGjJw25yJ+WkEPvUvnhZxaEQI29UY4JTFu3oqZY/3+ZMf2PI+cdA0pSAYO
13vZJlulNYiNWt1ZzUEGCBZ9hBqg3yHk/Biki8DgNu5hXLJSlaebeBQIxkgGAdteyplnHmJBB0vd
wqGXgf46eDNYXcJyF8jrfGWtEa8eerl5x4DteQUXBlb8RRPl+zk6/7VIMyYds5XYtW3AzNfF9DHF
Anmz7IAeX1smmFB9ZfIqcKr+ShTHEhu22tzq60zWKSk3iZUxsXMuunkzqf5/1bKsLnZOzeyv36b9
7vH++YJcuNwZ2ErX0i0L7xwBwljZpOaqQJ+K/VWsuYCMyVvMQK15KxiHSdb8e2SqbHxX8H2ZxU6Q
pYFf8OLwXkLcWe+D92aXxOVXi3QX0nrFnI71V23aCNJTlZD9CQUKfv+YcsDOJwxcuj5ZzvKAHaLI
nVN/9/Q6Asut6Mw+c74QJzdUSWMn5EyOjx5xxO2uxlgPcjAyMoMS2tRvXRPbQ7oso6kG6T2Sbu/8
d/J0zT+sY97lr2n9Nsi2WNs/VIGFCUW4SZOveIrrxrMORSGdFtVNQDVqt0GGNOOgZEMGh40h82DK
7vF2EX9g5bgLZsrH3+ApQniOHXq1LzGTpHkt7lkPAv7nTQr8ifZAcVlNTtMMViprsNADffFIBOQD
Hm584O5gNDDE88TCjJ80PiHsBLzMiNaQFc8OTb04y34BDRshzdIvIQwCRdU9dbVCTWfsY1JkPmdo
pSf+Dvf1DmlRvAv3bbfT+sQDW4sgtzz3eA3uc+T2rM5wM2bM+VXp9WldYMXPUb7uysf/ErYgpMpC
E2d2uduGRnrzGHbN7TSTCIWDRMzTY6Y2K1YIVhuvDX1iWGax389RsHP+AL2fFSNyHuqAlW4lMBQy
u63jdd4EVR1xr6VjduvGQMS1OQ7C0KnT8vZ+qdhrwc+D1Sm3CvIaoUe+bwdmTDp5FmCznt7Lz8xX
O8/IzaSRYyjvIBV+L28fV9W0o3dSs0xfvklTj3rEP6SKQ7dU9w6o3Q/OYfh2KwRLB4C/MeM5WWHo
hyzxFedUCDIGBKyTTUnuNHQiBB1s2iQwWf21IZ1PGKqcopmMoQfm4TSK2zaTatMvZ4ah/0mBP+Me
LGxjB23DkyYkhPa5Bpd6L9aiPaqiWwvnlKvFbwyhs8WpN2C2VlCMg6wnLT0JvIm2CBPRplPO9Zk1
dgFwrzi6/Jt4uFon4711xNT0a+k+jBoRoIK32ACV8D5aid4Kc3Vn6c9z9ED5pJh9+obIM3pQROM2
BuKwPm9CakrqxCrqtPh6/hcnDlBC4aoDtmMQmivImLz33MuOBMdq1QnYyLAy+iHKEK9RZeKIwA/L
5PhNsdk5ZYWFOeyQOe+4QoerzrsZDV6BV5iau7yKLaKX5RCopxIHO6Rh+2LM91vyopyf9e3hEGwJ
PJpDENLzC7HmauaeuO9XOx2cLiOfIrfW+SE7kN98pQdwZaQoT7mcflNXHxKnka5TzJoGFEiJ5loG
Bh/K3g2o039drOL7wbYRzn4Zq/Uma2SnxEll9sSH45+hyPBNxlXG/EFXyyjmj7K42t377gXxBVSv
lA2dWqc8f0/bP5sxs/B+Pn/VbV3SLYv8flYHHehtCyR058Wm8x9eBImigWdM7vWK/eGa9LpYzT+V
CYMt57RZlpE4uohVHY5hIg31NBvBtshr+kfDkjHvPPZctx1dp8dcb0kYDMZeeyekEzpMg3CwaKwj
g7EcOyNK1Ip+HA1NR0NH/f8qh33nHT+KlhazqmfDR4AoMBz8PhPy/p5fmgB5bDn1ePCZULRVPWSK
y8AoXZvUBxjBmW2wr4uKZcPQWADlOBn8ybPbf9aeBiy7I10Wh0rJOcrsnl7JOyuwBtyzmPLrffI+
8xabQ2AHM1EzLM1jRb2HmkTOgUgK2b7xRe0eJ5XyVsZdaZUxojzk8XJACf5BhPCMb7VjZ2tC9MCl
Cf0S87X5BbMqh3ChL0xbyKTq9QBh2B+GAj5icQSpiI1KJ7B+hLHXGe1HYHfP+ykKHbPb0clpcUEV
Q9FiphhfO1piovqfWxEfWdBqyfqYlg5f+zwibU/lT+Ei8lWkUPbDmqjMR6vObwHVyxX8jrwznua0
AdeCa6lXln4hJRVT1ZG5RJd90InbwfG/vD3vwEe+y3pzuMXO4Y4nc/Ar+HAB/BnZu8Od2XnY+n50
00jFryjY52NHgkdZwUQoLsJdCwxocojuZjOLLpc/eikDz6y6oIr6rKUZZ9JlCtFFKaYbO8U+A1Uh
GLkXXuF0HJW6nHi9xuQGeWWh/NZe0ewEL3Rn1RB6RCIh7WF2h13Yv9wHT0pKnuGfJ9Ilq9zd19XU
jfBwSTZbHOYoNxhTlyRBV8XfJ2fRoQtaY+6TKp+bu7y2IzMcN5peDJrp13C+BW8BdioObsUZVn7u
lVoHXnOdBKCOzHcYoYpONEN5G+Q7WJGJUPI0+0uknpN+QbCOZMqjd6wA04IEnxvd9IgwJuixN6FW
dolHGAvfPGe/soSIVyFbqyrVvTD1eOLltrjYFzxtF75PpG5J7BIsfx/+i9c20TMaprulG9db7KRM
L/+oGa95PJW9QAbD8eSQBjySFlgRazsTDJSf/eyLaH54AEOvTHeqvou1471QXpqk0q0h0GCCETQF
tLX/7hKfumKCULeVb+j0fbXapIQs0hTv4Z5UDcULdH9r4rsBI1nmhUiU26GIdoeLpF0BMfCXrVe8
OyZ972inVvNAW+Utci8i4LC4Sl6nPJazICJ6X3jN23Gf/Unt+GKxaRFDW5ILlWCuW8i82PoFkUBU
zIl8JOE9Stu4G4d3I/2DuhSqf3buQFIbHjoBhJeQaS5dftTOihSJiawnjH7ln3xpK+yBFnC6u/er
eVhZYolKF6uOkNBogpN7HLlR3LD/y2pEWNzRpkp4lum4iDAGOHyuhDGCqBZoStYxj/3lV/xPM/0G
aOgBTYcnnfv4iPGiVUMwyluzu7jvGMICD880nLT4Kh6LAmGyTQccTq+TVfljRQGPpOXiYOdhMOtO
f4MmC0Hy4kNDqYVJhO6C9s9jgyBpUevV2AuSbVXpmcpCs5ufN+PI4M0BTgpglfrsINhpC1WIeCnt
w/mql0eDeZ7ofXhDJrfL2r7Ujv+mH+TGfKU7cYFTXAKBFl9D4gnVJWbsmDOzQffKydYOivlu7jWo
jaJaXRrhWvHwSQimenZQANDaUIsyX9t2IekRA+tm/aMuX+JK47nA5f1tqgNUbX2ZpkM1w+XwIoug
7AdlDSRLkUc4jhsKixR3UgRRyMxD4VFHGwqhinxAE2FZgM1XNPBYbpqrJyE59WwksvYJ5b81D+wb
VIpV1g3KHRznBqgZMLm5/48Lb1oa8x0rn7JmEOh0t0m32DgnKy55yzj/mIwh4J6RrGG4Q14+UMK/
/yFFy8velKp7/0IbDxoqYn9DnVDZNVcsv80irzwrNi6h6N6mhYO5gvXbT3ekVE98HIBGURdVVW7f
Bg2aPupS/007CQP99lf/0hE8blVZTRByJEJEysG0feb8mHPNBaUGewvQ3GDiRCD0cTwYYix+sWgT
AiwORd8jORlrT2Hko5pj9Om9KkyM59DIY4TJomvtDfk1RqfIDCntn130MYSQiB/BIUsyroQN5yNq
mKHeykrV65TKRywzKQsA3U0g39pc6n6tKe15ssekREV6+6XsjZGs2UapxKmXFeAMTvBilbABmdXe
Mj/l1e0BmyoWldKBzr3jsX+/f0QNwJZqli+XE45WaxYclwiQsQtkSDUR03Hl4zXk48Y1Hnbj0F1p
lu2CUFE2IYgH7EIS/s6ya/K0D99xY+Eyci8p/DAvB0SuutUw4J+jBDY/V3pCpyIE1ez54t0dqFxj
5IKJpatS0xOdIRql7FYyGz5EwjmNe2/qTR3/RMG9Brm7DAyzKLwDxoJAHZHPWoacjnMyvpQsa7Xk
W2qpJCC3vY4XGUUXX91pyWQhLhKsHnYGxwjDBXtdKbJ4m3zlfRpyZJr9ZoTVvd82hhy1rJgKitLN
Vmy9grsKylkRAQ9ruWvkY2S208BKI0/qNZ+ZqyxcQrw6CC0Q8lBf5IC3QdhZxSaiqGTnHPUJldNZ
ll35Bs/P3tiFgQoVNbzImtyxDJI1rP0rBhu5yV1de0EsTyQygkWr3yZUyN0MVaEuuT+u7SpeT+oy
XFpfhMrsqOIsyCBJGKg6egqJX7LqecNP70H1JTrHkHTZ7B1mSFSM9IkEJ/MsnlV2nO10ZF1kT2nY
GvDywTpeeMJJhhv+77jnEuoHi5aH10H9KTunFGnT/XwITLQHA8G1toQoxYUo1lJpAWDHcIqbEyZU
J0YGfxJImEKBlDOROB2J2NdyvtQzZwO3dfrHsUKrIPTcA2GzyASTtrWtm2lnbgazli/ADwv1kQ6v
WtuosnBfmrt6wYtV5IckE36Y7s7xo7FNgrBsxs3A8z27+OtQxFqhdLhOQagmQOCo2ArURssCVza0
1hkCRNi37d+T/63yxJet1CRN4zeIVk0PI5K+9Q0j3C+EoOCOhoLKGwqtlhm/uSvqDXXJF8mGNLc3
22whoqkZvkghnlacu6OXOeU7CxdKlwLmxwwo1Cp1Rfnx6UiM6sFOd424D13+pty4qyMk2oiEdXoe
AIpFeKFtoi39SsTGE4x82niq3fJkUNvnUc6X0RgfEX2CnBuH+EDThlfwluC8QpDkp0v83GLyOSH3
hDiyHcuh6iL0+/e48SNyhkiOTLR5G9CBGKkvUT3AokKAAFQrTrjhIqrhCyqw/R2CL7MMqtc4CGPP
yxzZt9pEC4AiKrXayTAsaYeFRjE+swutrtJxyQPuPywvtDdvTzx0undommXSkUt0NQEdvmJeptjG
fQ5IrcVC+VDHKaoFl4yuLIdQJQg888AvC6nTee5ddSHUY24sJQMbbjswxaLwG7d690hfPqf+JzMJ
QmYRCY5L933Uq3NElVJo5cygmEnRjLTUsUyzf3x1T3cOIdWxfe6ebebtMR7hxkno2nINlO+wzzv8
IQbEg71dVvQpSbm/I3SIUeC0EeLpxobobyVaNH8Q9s6WZtZ2ouTUqm7pfzoKvJJmkBqffiBj/Z44
hCETsJD+MtEpOXrmz0bjmyrqcH7t0QLvdukp1S9WW0S6YHSKsGGD4tX+QtbVwIRpH1Q1D9czpXwf
sSFxk/X+rRBiKEKJWQov4cUWHOBnTiPo3AXTjEzlha7hA6/i/2/uNvmVuh88ZRpMoC/PZmqNvaqD
+43HELslbLdNzcCJb4Eug7uWUq9Fulrz/jPstuw+gKpXIlHfn3EAn29z1D0oXkXf2l18Jld4AQ8O
YH8K0HzfonM+spzEcivUuPVEgBL3OFJI1OH2xfkUivDKTUByRiaNcmTYFUbouMKIIojWqbPfYrDL
mU61bLsnus09cCpu8fXfhyCwaxrPfpWHhtJKSxzJE3yG3CpWeIofbIG6pocBIpEoNq5gm/pTstsx
Vi3DGTBfP1Yz7GVx8uSJ8xJeYuUvxpMYMGdtFmghV419Nj3zNhTCRJsPX7gV0qbVqDLmRgxSpHcY
cHLNb8C3L30mi0arjQDX14RSpzWDl1tSZBJWGvR0KBDxV2E1uo1RMRD9tyG/LXVGDe15kKc02Vpa
m5mC3yZOAgsu4ZfHw/kDnEOdI9WXvCfVmRXirmuZG7KyomJfEbezmBv5mzcZI/S9naiYTHxfzpXg
KeOH94f/qtauQ8nRkibhMx1E1jEgVUWk9bX6j4aaSxy55yNzyFGMOOZx3fxvpaElNRY8vGQDpmk8
51tIGA/Z8C/owM+5y8APsSfv1mR6TfgtHpTZtvEq2dr6urstUPPYgMn2NiAmFXLU9vaV7f8KhJN/
uHdozNtIonz+yWHAecj5WevQDhIkPBZG5oBlImAkJAaKUwkuwUnCu9ptSz2zDqOYJIsj9C1F2EfK
JdIgXyi/9vvOOdb2sz1Vvpar18h6OZVkc1GcMocFu72xnetLp3t9pgWougbNzHmXTyTlQfMVQ7TO
GzHO5EM6E2HgYXQUntPgA90IuybuvGw+Mm5ptduQ9uBqLi79wHMDF589wDJZVa9pEkzHDKd3jM0m
6N/LXnPQZbKo9CuXm4Bg2IiyQzhjy6fxBpTY4QXYymQwSAZqKf+vloefRXSXMXNxn0uOYWWmTIgq
MGGSLSSogIuJ5IK7/l6QwhI4Qzl9TfmWoLIam/WToNTVlqAjcWAvsEE9BBtppKuDyojuQexd7znK
r10NYKEEuXJwodv07Xq+aiMFMyj6LwZ5PXv6z2S6tfv8seSOHYa67V8d38no/eRoaH9zoekUyEBp
c0g3EvsSs+5u02r4vSbCG14tFY4D4CuFfzwTrPArY+w9mu3USGA3V+MFHooDZXW2wv8a+qqiSsWS
G1hLojBrtXKJWcqeBY0b4bO0n0UY+NwBSac2/t+kx50cTuuFV+bRwe5v4TWiWPD9A4pWkvazAsTn
kARZJgSWouHj57dJ3aC0vfQd0OfMyw7lGHfU16pS36x4YHDvDcD5RAEGPRJ1gvry3095yxiWXTbw
iJ4EYxZvOT9TH7Q4ZWRyHcXEqoaNWsdp1d7w99ckn0D7qJ4RxY+k7IrznKm3Vymqum+leevMdXtj
DLICvrZ7+YlzpVATemv2FpPKsw6P5O/yCO8yNoRIH6wzMV8CxLSvRtqPJ8SdVL/0sNsE8h9MNRCf
p4zR8qATGUyosHSqmHNvUD8jRawTY0B+EGMvKmpXwUNpOhgBY1LUHgK6D07YmtdhiDefKUUHpXsE
hmB/EpVbhxQRN2nAaEfWoay2m3WGKMPjfg5GUmcIiMzEltvr05khE+8y1MYMoHi5u9GOJdU9siQP
bV0XPmnAgMe6AutqRYOjCClwXJWJAFDKEhWQX7dE8gqxS13/7EcuYtXygzGRQROwzzEWTeOYulR3
1S1pvUsAKMPIIkOH3eCQxur/TGKQ5bWZ5Rf/CjLhDM2SWTnqoJ+iYFU+4txzKFl8zOSaPQi/YFVb
bTxO4tW014DTCVYFdId9avG+jSH3g6steU38vTc8huSsXMoH6n+jUuGhAOd5wH9DRGr8IENtvdEC
QqAohUvNWXHe0gD26EYzAHTpPJDukH0WVCvRWWAbwJhw0Y1yBgBwSfB477a3PLONRqhiKdFangmU
zt9pejXASHQxjZmFVUHT6HihCd7cuwesi+UKgp+DKyvovqdD3qjtR5veKMRwjKTD983Pk3V5cOxr
Mt+wF4SMN82um97v5QUPMch+KGCR533EHQufaptVbBIp9jQTBQp9zuXpK+B1CxWztEJ4zF68rNDJ
DvcMfiDH7cl21DQHfurxoA6KtQ1m8OJQe8jHlc796IGomVAcPVkLLpeuHrQlzlBNCNiyb8v4k0mJ
G0aNT0c62/ViqFsXgE0SgaIUop77RAIlnZDMCppaCDSeg1MROIZp3EwwpyXLedydg0yRje84i+xp
RwVwSGfUi7gGKLOKH2/YR1bIfuajfav2fcfWOMmlZ0zvspKO3Ci61NuAyT//9c2OroaBFEzBMpsb
OcMm/mfGj/NbcguqIB7nYWJHTYUK51u/mlTnRgi/WZVi2TwitpQqzZOkNZI1KhsMrfAxMNRKA92E
FZcKsfM9sbnxuip5qC7AdSCT6YO/AX/a9btX01onhlwxwuO2PmQwzoDpp4EPxOyAB29cCJUDK2d5
PmPQzA8wEmL1MKEQl5ytqiIHQghgH2k5MDCPpaz2SvpQAJegIGCrwUYc3wH6MBloVq1pEQsYC1PO
CuVtZHCUZdbcMQfexjqj4/ZRQmoGrKSdf2U2cZxeEKdlUvhnX0d7k4rsKq/cJHTqy3TPKme9XAXj
qfEWZWT/9c8bFzAe9zEiSaJ4Qo25OrIDIbOd4CwV5j97917qGAcRzKtIRH53hArRQmQSQ3XYsc/R
aBRgqFI0DJneXBQCZd9tFj/wowuwMa76uVQ+awoXctYnJNN3qv935jGqT6VThY2gSHFtpLSLL03g
5zn0/QRJM/5GnJrcqP+SPJBxul4DPh+RBvFkXoFQ3Vgw0IzJSTC3si6Qn+ltxgt9eqq0Pe1Okag3
szP5vPjAXwZ806OIsB/BVunCum1Wjl15AgPQv7KMjtZHQUZFk9VfGyEqaKG8vUItZQh8AgKTAQth
PusbyVO82DNmhMqJ0D+1jEDoz/SexP1AadeY1j0J6KEORPuWmiTy55m5mUBc0y3haB5fV9gx0Flz
QLlbxDCS1v1ewqYU8oiWvgYbe/qL5BhNuNP2+uA/wgTDwYBUk5oiHi6Y/npLLMx1577WbuGCPgVa
SWs2DLrwH5N79HMqpxSkUKQSlRBlul4oGiDt8cQLNGSTmIJiqhsWXzBuR1sttP2dCUkvP4fkwhol
Fp0KJYB7+/jvCG+bdyOFs0czmqqMXKSrM/faSExYbuqvEDS2FeBtJ9XKZ44yBRj11Uy9AfJNxEIj
4hulouiq4raY0GemsGMpLrwh8T2loAHw/BqgdT74HHcywnQVtWHt/DjK21ikNvx+Ith3Ei+Igc3m
K2zzqV6wgazJSP3BmRPnHeK7VmCMIjD2U61vE1jzK7wf+BoewI6eOoGABsIK0so/5VU7J4UZhelF
OBkFyWNJGdCbEYdLkZ0A4rMTUamgb6fxmd+pNszBmMVMRtpeukxKvS/6sKDjpdYo82L5a4nIJVHF
YxoX2P85c3arXHrh1xorz2Q/ygfGDhLwb5DfHjNgej86SLV/h9fgAeWUcXcQhLAcqS7axz56Xj75
+iU4GeUKc7Lw+MhL/lMpkOAh9Q9yVpaT9higiRpRBPR6y9fudOPscDlY09/Hdk1FOfFUGLH93lTU
Rm/N2OyZ/6SwsNxKw7e338FqPA9g5fAijO26H1iHjFxa9vIyTafQON9s0UoyYBY7+Wca0NAPlEzD
e+Z0k+gnBzm2yW1uTXNBi4pO604h7zYgcsaA6ODXxpycyLaf8UJw9PkvzsVTZm95RP5vft/VD7ql
PqhCP17BnrU5cX5FcFaWNRToz27Gu21/0J92MFuAu3VAmCIBaZKqUbjg1ATmwGfzjCkskgzn3+Y9
EFzBHR4DzwYGkjIBdptNjBoLeFolcuDTo1KMTurM/Vp0CIK1LwdSTmJPjdcaq6PElVcu7tXqSoEW
75tX4RX885oKtpeV/vm3SxuH/q9sLUFhBIWEcogX+Xv1dEo+TxTtMwH73ptLTojGKd9JtVPKDYNT
UdDidJ8xeqo/XvKmGU2nMpsK0kOo447XSoh90S7EEgXO22bR756F+2NmdKLm74uB6iCipd3zYIvW
Z4/0aXCdVkxIbb1XYe8+mHnwCLNomiw9cMP/HF1lWR5x1CGq8eERD2yM3mTCeHDejwVqNgXh8C99
VbZ/Ob7HXEqfEwrdqcrTVTbx2+s801sgXNuWHvsT+qbiSGFBhyAkMLCTlmSjjxH2F2n2qzEM18yt
mklUV68oAVCe+K117lm+zbrM3M+qV7Eapc+EuMIDy7KxHpIrrxRCFW5zJcyrQkdOILTNeqzKm22O
TnPenvvHw8lVFR1LwWD+AMU4RJMEkuu8ruU/+YzXpwtxOMgeMqscN31EzS8vKhS/L+uHa4oiEjW2
4GKVF+Ue0Bg5lWN79jQxxarcBJGX8C6m2MY7Hb/i2ds9mVrlSwBr429CfK4xhiAzBM8X2ElZ73u5
wiyoCHOeS9U5k/daeyQplTTKT/Ro8Swm3YFh+bnGynt10l3jt9VByM9oFOFmLs/eWDHjtWUnlIKR
6AMlnzBpEDNd7yuPM8Fr2k/B9WUOOO79WI/gNW7Vt9XVVYS8asYjzQX8al5UitNHwAoeMlKPjYra
krbuaF6R2lsDN3KZF7v9PRVF8lci75/i9aHxciFrRbUsmQldFSLf1V1wadQVl5ZlAFfDQ8WpnjTU
Iu+/Tzjvg26E65tQ7cnTdW1rQkKw8JBBNa5HTxWSrzvFdT2IYIj4oHYaVhTMiz3z69BWOQWDYT7l
+Fe1/piNWIckd1fDo3oJa4tuZKRTmIDuN33msHRDXxSlTMk9yWTtQfPwnDvP24uhqEU0pKD4ayWO
ET7xl8UxQY/D2uIp4JJv5i2YNyOMvnYcqudO2T/Uue8SHo96XHkvj6TwzZ/2OCW6YlfxBIfDnOVj
4gZ8Z+Knvvmhez+RbE41NegsuH03fYnTTXKBoPL4MtcwUVS5c/yupNbE8XVFveBKK6+EKPnHV7Bj
X3uDqK5l0q8MQVa5ETtqYxd580MV6mGfA05FRzR/1AhS8wx9iXZmqNKJA7YNyKvU9TUcEMgPYNRe
E1TKchvjCd/RcrwaBabnXuRF3hLiu/2Tk28kGC9QAjOT4XVA/MXZ6ptimLl6Npzpn+OAGQMNHAHY
N0ECR0hxFh8ODAY+nHVgbQ2+ECDEbTNhat7i6RqpjcqrlfoFwrHxj/eAT0L+wGA9urFhPbtV2wkc
764zMKVMY8N7EtHcT4fqtvjQnKGlOo2C4aNidXSM8A0VQTfjRdKjhtqow+17fkaeFXFq1Mrct+Qc
LqLHBNMa1dFX8LMxa6fSR80vcCUlj4Pzzr2SHJ2gCBoEAdKwUQR4su/AW4lZM+E4B5oLJQdeuNm/
3QwrW0ciDqM0W2yi1ovPdc/9tKJGIBBaCWcVTGx03N+3fvK0tKKVncixFkyTDw4KT1AsqC690Qdz
jSCwA+35+ZeGFAHTzy74GZTfb2o3gtJ3AXLSz5Gfr5UM9VYQyHDTdAJ3j+EHodi5gqZp0Vfe+YUr
vi2wxdJ/CxogeZxlluOwjnK07NvrLzVJUKXQfRUh4laVLBbm5d/1ASuW30Kn1m3wsVdgNFs4sdQS
mtUiGl1dqyKEkbuQHcMkX0l19ZQ+sGFkD2uERBF7P1Ssg0AGtlWAmm9n+MO+FK6RfeihBQN4Mm/r
IpL7n00r1RI2Be4IBGXrMkAe2dA3Egy5fmAbN/QqUiKk0/wWWxc4/aI/8WlEqo2IOBRd3TjRNx/Y
kOGzFCR8ylke3VTQdwJM7nJRDGN2lyHcTkq65O7dWvzrfJrdB4as7OLh1R2nw+TjclMQA2b2+zT3
JX7tWqsw5/ab7EBdkwsIG8ORVDvoXWbjQIoIlF9JDiddaJ/vlVbGsE/UA2r2BZL+EPjAdu65WOEl
4Ahzze4EeBTdngmIPuvsA6ucJq3ArY3Drr5LJPwihpZiA/aNPiDyeC//zmNgG+hkv70rC3OpArqo
pJAt8qpeoDPpmUpUhyALfEUCAWNOKn8MpKuVXaQ/MR0upUEc63SfVhBYffC9d2QxkAbSiWhuiOj3
6EZTtjYBgdX9F8ZtGDHUnag7Y/BAL2MwtncyEoPeAw7cDFtynTyC03VUBStAjsEZMEzAOnF22FRi
V2k3gQPrO3Sy1UakoByAWIoxq4QporqyXNUAIqUFPcORiXEqJSNv5EXDwOp+MO8PfOejpaD64vha
pyQAqNbHV5b5PsmnKDgWbcrwNsD+v60c5AcIhifQnhtuuAXkER2418lQOSW3+v9KsY4LwY6e5y73
wlGLb3ypTizWKBrN/FfoU1FF+kNeay2HxxWDp6VK3tjrW5zXyqr/2pIpFweddyV7HuZBAMiEsB76
DSR2wYw8bTXu2Po5AFiC05lleQ6GWiyjUjqMH12oBkxnMrb8sLN8tqTnQquDmF9tJGnLiv+fBoze
XqQlgHLM9iFj2udfOMWYX/UXilmFSnKAMoyv5ij72FWzMP24AfdImaRrAd7SbQ5RLw63ECORKxuy
WrNvBW7IyzXgTmY6mF92A8yqh2Swxo6lEVjaVjxgUdytUgvtXHz1Lu2+PSPvoeWEFWRP/VegypzF
mU2FQVe2xrW/oYI3q609p/MKBxJfiCxoITSOPlaKKMwWlfd7ir8NwN44C1GESZLoCJViNHSoSELo
0Np4GqnJOZP36Ih01KRVpGJapHityw33vE7nlFO31suWc+X60+H67hFynA+c7N0h3Ycf+9jXQPc7
fbE5B/Og6GSy+waMF7PLOJN5t/bIJEmWMX3cGsHelOCHGSFGdVD9xwqIcuqL9ccR/WpBEdgu/eaP
nymMqA+1wtBJySFWWxoKfYgMx7nExc3s6UKnFb4ZJ/3Woi9110PKVmJJgObisv+4Cmf7iZv/7ki7
Ag2+9s2VWJzzUkIE+qedAlbDEg7dgI81gqVphlizNLdHbU36T9vVR1l5bO8389yVBuJvhUd04es5
3rJsx3EZkKOLIJG21SQVNoro6SsfjEp+lwx7KhO4oW+dt9LcC0D2hVQXUTABkO6HP1g5etJSSdBN
nqBDqPfWp4OKEnGOpigIF/6lQ6dCJmyqy8FwPmUDgRsarEiqgc662fb7+F6VIa/Bg+WTynFzfgzy
9T49/OQn5iYo8vUw9bO7Ol1Ix1d6zLD3wGpCOnvg1oMDrkOlaO9oapoCJjpMKDDJq2zMQ9yuFs1W
ydsFwWagyIB9G3HwTTsOz7Fetz7z9jFwnEp/BRGePbYF7QsxIwW4pKAeg23WAxWKFWXRXElzZfWA
iyvcgmxB0QCZOWZQTH5N5EpjCVwPIZaJxKeMGg1rRRV8KYvZdHVKddRkMADUP2UdGj3+NA/tyWY6
6oOpb/emhgvKhfu8SrkfRIgpcmgHciEB0jPdRl12GfCcMhwUByzYqFqQahOkDZNlai9hGzTpvHzy
Zh/C5blo2RQWeU797s0kI5m1b1imj0G1ukqMG8zLnTat6GjPbReCmfeXndliP14VUBYJipJfszEt
nzpMPNiXCF5V05usN4FoUUTNobpKcN/PwkueOwZTa/ceokRe572aL9fUrNbXBtozLVhQp1PSnP4t
659mpZ2eZ75QLu6m3jRBG1SnDRohmKyymp78zl/rm1IXI+foPNYV7Z9SDb5IHZmEVou6wn/DgRi7
qVpNekC629nh8Yl6Jzq+a2Fi8nFiM+x9+8aFzfaMErmPicOyVRQNZUQVKxwS6X04zlcHqZCX8UEW
0mqwJIH9l4fklixZ2UqK6cXJT+wh7VcZcq6sq7UldKh+LyMuVDCtk1M05jbstrIaqyk1k/eXbVro
vYIaL57kMZiDSIueebkl3C0+2NrzeHr/9D1SegoBdoAy/Dwy8hk67Uckcj8NwAvvmUQSMhndsHa2
1fnrJpwYkX038y4wFKERPZNzjy5Q9utWUuMNY4vLkk4IuQ2wvMdYzZjq7rPd1MU78nNnZN0597vh
cBSSXNlY6unVQNF2ZDDFBwxq4LXqTOIMYprOE1uwkwkLfLfbFyImm6HtSNZKBuy2bKG8qnmc8zGw
SRmLBDrMuO9XDTh2tEMfqVpISOoCX++Hr2BHT9HkvipL+e16KvIzZ+FTamzMN7HkXqLTkiyTVuHe
aB7iffrhsrvY6lfEEe1qCagQo722+capb/KUFA/FAv8cRjrgQ9jfxAo1G5Gtx1A/I2IT8+t0kmoT
r+YvB+DsLKkJS6JDNU6ffKW5cAJcmca6IVB75+8ZnFHVdwGJKK6dE5eQOA4Tjbm8sTkqwm9sHTsm
+1JBqmfcNKkyM0cg8uNGRjdwxzKzOxCxC1Hr4Lpv0ZotWehEjJCKqfh0JOnDL/0AOXx7cJ9WdeSa
u+/bQyE/srKApMngessIVv1sFVDjRTMyX5WQAgBG4CE09xAdB79oRn0UuNTXx186ula4/YO/jiCr
j8Bps8CEUCRUHfqbZbq0dP4CqtZMllfK7WWyHlJRPScKUV1O5X7Tuffi77ZvYJAilmv3ZpTpP8Eg
z3wh40U3DeCrZkGbK8pMD84CBJSq2n2Xt4nIIbpRgSk3lrfsvZkS7FjjeqYUTmk8OYK1qHZyaMk1
BiDRX9H254KvZkkfmWdrJj6j9lvAVdsbpZUxTZeWr536jNTaZ3VxNm40ZnaL5UsEM8oIhsq0EgYG
B7GIIqtJf0oqSf1b3Y5xOIvM18xjyEQLJ5LelFQa1WisTakno0eGteKdKN7in7WUvRN1AHRiZX1x
NOFxQ0uzQg01c2aImUMdMFWRIz/U5z1JCXPIpUKY+hKnOmfLIwS38DdXh62JT+HpmLu4N5phlcK8
MLSqu/piQcW3+6aNkM2iXzBA/eYUsS7bw7LLV1nKFVxsFrm5ucgx2w0x8Q7hbPd1tZjjbikaomTi
BdL3/kcN/VfqKgN4RkGyjQ+sRURrD7RCoXrW2YQK3C/7v2YIO7DxyFxtrKAfZiEoiH126IijCUHZ
d6krB7TX3S2kk2GwEWfDVg2En9lgb6CX+3ToHJ8WIrh3HgdHzgr6Xsz/bxKHt3x/RSSV+2YkU7NA
YJbvZN5kCpJy8NiV7XMqRE0qxKv7vNuRcgz8jT+TL0TQivih+FQ0QqBr4/pTAHxTz14WHHCWEY21
MMlEZoarZM+JZD/TDqCKBvMl7R7xQ+5v1NVkIZUftD6qYtLFwKabdEcPj3YHz4x44wN03VaSS5pz
Xvoj5OG2VA6MupMtk/TrxmZ43iUsVsNS7ZYdAQHQSzisernSN3hOkoqpOefIcEv/HuLUxNRMxQ+p
tMKmjzoBJ3tdtzEveV9ZtZDEzBbvL3akGbYRa7k4yJW+w+9Rkr6TmffSUoaAftnNMPJBSrAq5ngA
17pVJuG8pP3YhSeXINDX5jvBOCdNoFWpX+EwRiwD5JKTL+NhxAVHLcdYoGLXjTFYtVEPqcPXMdbR
l/iYxsJfXIXJVH2/leP2njZWNQltWYSnwU3+QJXHAJAsvnuW5aAZncvtbI8iNEvi5Gc1QFyWl4w/
7Je/BaT4lyGrayRKl9I59oLjrU306rfoz0f02gc/an0qNmVikaO3qvpHjnzy6+knk/QZoOmVZqlO
zg3Eaq5YXNcM6I4gL2Nmle30V3pD+qN1ozMd/xmGCWnsuSxcbp2x0CiAPb8HZwuLj9ozr06yWiiU
C2RWrNvtzzTuryHyPcM8HQkOKjIZjJGo+4QXXtzTPYbYLc8cT4CCWecTD8q7y2EcDAB6YTlytxu4
JjWcC3QE06rqHwde3cSvwNtQ4WuUGoq5q6DEqqs0fuohL4gYSVOJWBOFiMYtem+VcBocXeKwkWPu
Sk8eQIV5tzyUhBhDj8DLdqcB1C1137WWZfmpyaGSuzPr1COq1mpXqxv5PohXIojvfv3NqYvP1+0Y
IiDILX7GYr4RTBTcPptHb7AzWD5CfA3tnAsBBrOEEoaSZMI25EWnMVQqwrAOWr8EpUIaYuj3GJBH
sL5+v5Y1G6+ZQVWPfSJkcJxQObOsrBXb6gU4lUXnf9O53jHNLo/5850mZv8AnTo/JXCVUpwJdA1a
pYLN+lqKG3uODpSn6tHN1ieFGSw304LwIzl9B4cCASMrC5TF/QB+7URrU2/o6gDJ/iu2ugViyWR+
J28qtvSNCg5qAPiE6SANN6uvCwfqg2NF/8F53CAQ0FgpjGygTCwkQ7ZAizV5B2fHI6CsUWJ8Ir/H
t2nyUPzOiIB3JYXHZBBoc1hx56+zAwK/dBhJLHOxRkLFRBU3Ua+ECzk7gejWf1baSkFE4zDbwdmm
NKvMVJ+lPvJcI6gH8LPoq6XReItLumMdNQf29ROlUQXGY/n/aHqoDYfpvI0xj9jWeB5dqt7tHLK6
8ualzv8O1L8unI2nQaAimVXUVI8tic+Dr/5y/e1sss+SeGoT0aV2t7twmiGgjVWeaBZtFZ5Kbj3+
1wcCNSr7ppbaI3ABg5YSEnle5DlCFNc4UGp/h3k4Dz6sgTwV0hyxqmC0wE7Bj01TTxXXfTh8in7u
tYT2IBrtVU//ut3q52llJ5co9KAu/8gub6W3+E/XqS+KPA2Dbn2ATyjiDPjsZ+FSZtXsULvO8PL7
NzLuSt41ye6DDqpalLd5GbFCa/X/uoeTPhJxEZu51PJSC0G9TeVlsZ4FI4SXoSuOSP8hj+DhV6k+
qUaEucUC6338w8AnggylgAhFJSJ35xj9nvMpw5q7+fuJtecDFLdEbSX1xOI7i0BiFMChJVvxPjvi
IPhCjqH02DVscIEqkuNtyuc1p/xmjsEpYXxZPKfcIar6S41rdwSGOOPZYHzSXYYhfrfraW7QWS09
Wlb8sRr3oZUffEoBqDME4uEDhSypeA7bw+hESFH6gNQWSHRcrSjbsEnC43d/o2WVGh49VlJQl5u0
Zfcu7uEpiyIqVNQi39RfRlHIa0JGnx0D4K4ObtlhuG2Cd57SD0gjgHt5kPNlPRa5HK+fvFfv2jbe
HrLfkJGQTVIV18Hljzzl6e7z/dpL2sFZzTtim/V2cfE53akNt3pqWcRpcLg3Lxyhx28qlvWc+6sZ
sT7wSYUZjCIiWpKDEMDMVvmgo8xaPxe9TgNLlKQCFKJcMD0hLaQfG4PY+gFDfxp59hcBqalQYBRz
w9tLAiR+EGcGOZNAtXhgh2kra+Hd3v2F/gLyBHAk4dxIqN+yxkujRGGnspa6mRPAas9ev/qy7TyU
wfGhLIhgVGCWCvRVgIu6DhkKL12pI8qrTRQ6TDmlcGTxdVTjnAFy/R9wg91mt1Q8S+lUWrRrC8zp
2JYX2CduVgK1N7N/STDkcA+5ueL7hX6+j+OB8BIHEngk39FzFa2ShQkd+0YTk12AmBidKSz/aUJk
kIiC/F9oYT4ZDXos7Y8bhF8usU76QthrZFN4Pol3b95MQTym+sNaTmK3UatCqcRk+TsPZc8sbMvW
ANe/MxvPMoXtrMTWv7TtzAPq8x8N4HfM1o4o5I6j+NguPYgFU19iSgjuh6L9MHN/7g83YtJQJ+qm
w2bO8Ry4mxef9kcE5Zoo7lepv0VezzHnehfgQA67upEn2szETExFp52O/J1gtpjZUBrZYvtPdsdk
/Oug8uOtC/7Qb9Iubi6PUtPZg5HA5sIgEgP9JPXNrt1ZdrrSpUXiXY+5qzozSnRAGvtRCY7q6e7N
zJXJ2o5j7ipEaWe28Kzi2cgGzfdhK9bhSvCOpw2HEbV0eUGzGkhpwsTFHUhHoOp71yz5/SOWfPFT
c0Cx0cEOKqDrwSxxKrqHNonL7rNc+Z+FI2gi04c/aiVhNNqwXNfmaYV5BUrrU717XLpve+lgEqlZ
X/Iu42mDLzwZ9VLhKqPmua1bU6r5UEoQ1e9CFYAn67IcK9nHB2irhQICIyIwl6bW5wbu9jIc+VOO
mRL3WjuyZLrRZ97C3V54iaLx9IhQel08fXrGtavXX0G4YdptcvPQSTv9OipvijvENx82tVTRDbh2
ABY6VcGxHTG+rRY6oyFBuYfWr5B3YXo6cYYaCI4cAyvkbEM0Ybq0KOm79Pbk7K9iNNFcezgrpc3J
V/RFyNs+5tJKJFTcSZKwTI5hjqIY8o6A5Cf4iUvOu43Qz8WAFNJ539sxyUjGNr0Xh/bc3swQ0P7V
LLlT233L/uyk7QBlCpXZUxe7DpCFPWj3MQvDXC3Ursx/9xqNF6wdOG9+twAqwWsXTUPK0Nfc8zCC
XmCN91NcNiGkaHvz0L+azHvy0cnpOCGIgQ3uBZXMvZ7hnDm1bVku10B+yBjaFvLLJftEsLbzrLsR
tpIeNUPUEKeJA9ums4fcMuBOLQupbnT4KDLzUNED5dDSx3BKjYaCMmZqMfYOGKCup8iSg24qdgXT
r4tR138eq9jgVr6kKegSJxsTjjsbfUZfrK0Y3ohsS6Q2YFlivHyQAvfe6hcz/UlXO2Rode7IS4v4
TEsbicx8DOoC8ICQXDP4A4u3jgs/roU1eMoSEWcCRWQsY7yMYcnU8+IafVXC6LeaszuB1i//XJwC
fQ8aNL1P3pxUVyMhAmMwFYXLLehUuOSm64U9hHfhR76jRe5B7uUX5Ao9mC5OGF4B0Q/JfqF3UwsY
7PXSACA2tddwf+6prD324G80hDjb9jzpNEzxwebgmDnBWAtTLzWimSv3R82ENCRvHhAcvVSPZa03
6E4lj2nO9YeUF2BEZrWtSUsYDEgmVs+Zc8xxs7cBTOCcl7kB/ybA0xzRMBZSvOV3RjVeYnZO4mhu
ORXCoaUrqp7N1LCC7Oav/cKgL4Cil9tGIcTqwI0b9md4To4n0BS2f8kCJ/x9lQOch0OC7/TYtMah
Yng1TYNXfbUXfcSyWEGXVIayCyiVpMSUk+eOh3DWgHnff2eZHwTHWqDy/j64T1FfIASNGn0rZr9g
eK5GqG5cUBW23ehfYJhZKR7FZAvml0GzY+F4loNYOu4oTNf5pAh6N7rYY17aVIheDeOWGszZoQNq
iVRilCIzF7Z8/6Pg8F3Ysnails9t79jrdoUf3NJW4kAPO/gAa6WI+oGJiqpbv7KQkvos5WsQ8BEF
zfvJemVxRUgJeO4ExXttY7UjH8jMYuKiKpExt8F2/3m/6uFqRbuprt8EO0lx6FzC44F8KlX0525x
pTK+jnsls7iB1CnqTCuHlMasRKAD4Xl3o/dSQ1ADKiTl0IRcm/b3swFAYtbUbvy/DytGR04ZmFnU
yMrodq+npVYpwMck7Y7vz1w9818UlAk8rdVmnZkZT7Nb44vTZAK2UIqqhK0dgfescaLnVHOk0DZl
k2yMtgL2zGd8W+2852tmZmYBDJ1H2GBZzCKsP0mSNnRnf2ZUvScSuIoMsD0SfAYqw94ZkIShiOGY
rXTEZpwewtQRkfnumlbh/EgkFix+bkYWSAbg01gdTLwFhQOOPEW3vGLJqTUCEJhXgoX2GEW8igR5
jWvcY/9b+WnrZExcWWy1h8J1ZeqqQLPHehBHaxfYtrC27E7RQ9k6KUGUVOIRwKnKz2fvAadXmw5P
mjrTItCrK9XxHhNN8ycjv1vLcYPOa4O3J923hvIfvuFQS9TLDgV5pNv2exjNTy+hF/WWlLW80MGY
nPriOd9q5g6X393HzxfljE+jrLfI6vQvxAEyXgCIJShWgsuvJiLoZ8PDx2vwRPQjVp8I0v9M9G0H
N+cBtkhZACONNHgyBlIkZ8K/6XpBleO6PwjVMkPsfF6vvRlR41IuMwjI2jr+7mNS8j010aYOEorl
/jZ9lp31pUW3WCfzgfNUUMWxDh4+Gg5pfiZjyLtkWghM/VbLmQqJcSFAKqzUaXNBwng2QVW6puLW
1HvOi9aFmSQFrVu1Kq+kvrxuev8T2OdsE7mDNktHyWoqiI424krvhZTqBaaLqmrWyChl2DhTp9WE
RnbKYbA8Bs5YfZKN1fYlBMtieje2mRx8HtNGy7MU1Eg0zWcg4GzzChLWcYna2ExO0VYDD8odo67/
FNmgos4w7YUFzaQu3mHMDL1IWMxfgsMlPu5Xojs1tin54HyarsWQTBOdj658fmqKzRw6PMUfYElT
3bBLmJ/UHXYuWpENxyqhfCnZOoJPZdCzqub4aowHmqamWEmIF+ROQqNjeUacJOcIeGBWzXUc3IrX
10TIOwzPgeCuwdGgntLMYFzAs48fsqDZXQjCmg5VLH7PSgAl4yCElfPkW5XTsERlgNuvgVqNo7+V
LQpMrVREFP73VEsucpC/vvPEFNgI05MO8dgENn+hA2ON+u/6H9TAiReeXJyFFvaVpFjn6plDS2dx
4CarN5M3OfvKt3BMVdgBGsZ/082X8wfCjMKrjIM+lZE+mN2SbS/wynurtH/tJLZsdxU8qK/q6F0h
ZDs3qzw1yZXs60XqlhhyZy9pZt2ZGu0VNTZMh+YQimJbb0+BNTj0qLyVaK87M7C1i+KoHWVZdZUs
CGQZRseiztpCX9Abbjyb0E9mq+o8OdQqnEDYWEcwYtn4qUoEoATI6C/iGDJf9XTSZn+xxYBjbB8D
y7nVRx05j7dnoUjAD3hAuXpgYx4v7tV2BGOfKBM7EjJlBbVRjCJDyUesK3vsawClyq/c7q7Hh0KF
kiG737ROQ6V/3pp5uPE+It3QE8O+oAJDj7eM+fIZUej8iNbdududbKs0JRLSbTVDZlpopwKf0s3t
9vtCDtZc3go8Ro04RxV4vDh374AD6xvPoNcBaQ6U3vlg/ZDGw6bliuSDph2T92bGXzCmHJ5S8jl7
4mNP0QR56xahftewI/Y7KvKR24xkAMvCmqPh4STKtcTYi2IAsMwPR2v8ndBqJ0fRopwevEmiOIV9
teyfDXS0/aGp/+ujod+m7wxl0Oz5JK9ATREa2+UD1mcx0QfGKlvrbZTs+LRuMplvxj0Si6PC48OA
wxJIoBWr6U/y2VxEbSYoUR/rRDYIhiNhyXi0xgadbwosdv0XC+QGVfD6WXIaOsTZ6O9VSN6By8YI
BJ0NtcUwdEnWTFkKxdsRGbxL75BjaCVeUGJbLx5ql2Z63Q5BDYKT4/TH32hEm+xRofs7OR3tnzi+
kBjUN7CMiJeb3v5tDuIvG2TkX1eZotMEe0iZK2idFansMcqwPhX27JZE2UTIO28HhuC3NYpCNIrk
QbWDT6S8IIz1G8EGHKKNfGpRgThiXYX0mM5Lc6kqy/L8hbMURw9zqgzaK4/1l5r5vbRa30hNItQI
wUaBn/rF4p+hyF8ruOkbjTJg738G4mRWdi53cOd+PAgMi2DZ6gYvbevYpyGXyIn38/7t2vASicnW
j3WOhmERjOLbV7Ee6xRdk49i2uEXTBwKLILnU4U9wPV1KzUg5HnH/LtUv3C/rcY6AkqP8NHKTfQE
kqhLcUgwxFhm8lQYImlFISBVvU+Wvu8YUnDt33ejO/XMPq2loQt1EtEcS31sXu9fZ4AZuuzKmCxf
jfec3Zes/kxhthrGGf8g2GdG6mytM9e9A9qHrkIyhfYKDVWk7uuSvhINkIOFZTQSXlcFm44LBJgw
mWunqXiNNPD2s/Tx/Kg6gn+JaVxPR3l3wbdfGoZHmZb29n9ygssvLb7rWGgjFe66LpUIXIF/YAT1
/LYkhRhMKa3W0dLCH1EWHh4gIfCmd+dK8U4HRv9ixSolVQKRj9ZCkpwoZ8VtCyIlwRZmHVOvt/ke
gAO+GF+Zee8YBOHmI78uzzd/PaRgs9S+KG/42408jFT0bHZ/mZOiDDRVNnB1GXX2tO5DoB7WZd71
IZHVrPbId2L6jYdz1exr+cl8LQp0HMm4t9+LDF8+7b4h9YS7hrh+jlFzKNceR7htr2CR67Zrptzf
zLSVqAm1S1RVBPlTII5O8jcCAYNQKHRtDQIKHVZ/XlzmLs9XSd2xUkAXldn9U/YKy4D3gqUOraKZ
hcV3w5NM4+kRhtzDbAJiwiyugSh96ZcFfeiDTiLYh1HjXshjMNlL5AOYoWKJnXBw4kb7jxkXV7yC
RoQhji8d3aYs7o7vGu5Bih4gqkcSRUyOZUhO/7SB86vsqzZxwQ6oNvPS6SgW8QnVMqbP0DsSxKXI
xn5Hyajr6aJACn3w2wBKaQM2DpiP91Yfms60/PPXbXk1b+OoaqbxszFj9pgCNjz7r38WKycLKoUF
CAqmU5DRmS+8UfhYmVvyDgF/+3EBLvxFau0arYlZ5ksfAIUte+FRTI9jXYyeTKqLXZpaiUztJop+
aNnu3d8scy8yMsXlpBgzpRplvArNTOtf7li1/UMz9BGdSAwR03TScpMPrx1aFg9dlvopi1yo/tg9
mUAavIdKMhTPrCC2UPEgj0KkqTDAaG0DkZWzDqr7GwzuKiAgljcGyhKzWaRLvdvojzTu+h83LACL
t0BLtezHPTPSfXnwqkoczbsfHdvM2rnCT7Se0qNY524ezdZPvLL/YduNUdA7dnTpdQQMX0BJXyFi
sDewaGnuztKmApq4P806bTvPjEbKdeBm1Qx1RYCD2LDgnj4XaZp0/6gCM6KHPN1RVWUzFtQYfu2h
mURkEFG0xyAQ3RYJwCD6q2w3e3S/QUuXEKf1DgxfN02edJQcTbN8w8JO3baKTY8UNaafxT3stnAp
Zb3LqhiB164UXtk4kLt3AHl9m+pQ1+ppxyKPBvrle9vhJ+H+Oa06TFNLl/J76FXLAbf9lS0EB9x7
LZKTKDIOnDzVt6abmdx0ENDYsOsyvX/K4lYx+ba9x0AQyLpuo44ZKuBUfefNMsfeltX0GKhpvJlX
KcXuRRK3kIIhfx3z1MpHqZbKYf4UtKy4II+sFUiMI4RCDy8rm7MnNGDW7ZVSbs5DYJqiWvQjmaNx
1r0HINbDZPGQNoheExhn2nVhcFwQw9tlYmLoyH88jA6NzsUKci6Gw0Y39R3HvocVdD6ppc09HUcD
p6lFxsLH7MpJI1d6DAo8zd/y9E569kyFOzF0tELi+z1g6FPYjJkWkUS4ZuSJHBkCJ0Jzd57Zh+L/
lfULqjZx96pMEA0Er0rmgcIS3e2xZsVIRpNJ4joIqcCxatEonPUNKulksasPXctViuwvCb0mmds4
bR28VVvYbQ8FYccBqYB2qjhvyiyNcYHTjrDMl+azC1xCYlgkL+Qkv8ZxUnj1T7uP31bmThBVCH86
IOcLzTLZiNDiEQgytaVmS4A15vcEJ2yNEwPTkUpFAoHterFNbaZR7mLey/qXqoOg1a7u7YZCUvfy
sqPONZcIpmy6xiyA4nSpL9y2DfEum371+61+mcVmBUC9VRk4L1fhPX8kJT9QOJ+pBY2joXRhh73G
YcVoQ4nVA9ws0Ck5UkvYiOzTMHUSr8p+I0/PBceeq9Spqhl3PgrwNSf1sCtbhyr0eZLZUpO7SdbX
9LWw5FwpNvowUnVobgwJykt/QS8/Rc2tQYkJ9FhbsSg4eE1n5OT9GXXZ5ZbxjLFo1JReOEKIGlSp
a1EvNe1RMVWKblvxb2V/Su/701WKC7U1afoUPFGjGpgBizj3JD8knesmCiJRwY/raokEM2zXIyFH
KPB3NyAMld2PqDenL2wSMDOnErXxltmTSkqd/N9FfnbC/H0Y2iVEus1L/EbaxgcGzcBX8HHxQxfS
LVDkIkBTezIPQx7tF21WkeUylFjfknB4YwfAOmZ3cmFEWiBdQVPkfZ4bzPKH7T5tsn+N1hKoyEGa
tCxLjBjLTyBlbPPO3Dv6dh9qPZIaNdzSYv8s7WF4gWiGBk0PPyUG1ip+BvXCNxmucctwMi2QYaPM
z98+dCdF63yCBokgtsy9wKccSOLUoboVqBuZyB38DtAzxQmMWUuPLQ4XxvQk8OhigD47Cwy0JX7d
PRfBVOy4zfOVL22MI7sXXgTAp6S4CI/1AJZQJPaI4fy0wi/2QHNO3mKZRXUtTrGo7JjcRMPyUOUA
ompbURNFx83RhSP6MHZQAvC+hZLPT+BNzEv+yDTAfms2yrREO7LYI9csrsgkgYGzjwuIVeZOkeRl
JqbAkdNoyfT/75gAx6slskTuBeGn+QGbQ16XTXN2HYxiE6+bc/5aBM1lVwF83gPyXKM4fgXL7SnP
m20FZ31DW5IA5w9xRAgZIYfLY1S9JmgvTOxrqjSAOlpnnEMx9aR0f6rweE29yAiAkrqeddGdFYMQ
rEpRbe2isiUF6+T1oTu0taAyxHWo3IUrFNHrkL0ZDYbRJv0vfbiHdteWrYwjjfqtn+tAxQS6HYQE
2CzhworUMnxjd3CP+RnrjaT2n7H9O3sd+WFQi/376zWAMjNwlqNPGkGWpPiDL0CX0jljBtad6Nl2
+kngwhl7W01Z9DdgqsJ5yRlKvLrCKXMWEu/nEc0so5Jna8rpj89605ToWCQGHi3tm5beCOA7qQdm
rkIVE1hychrJ05BAUBtCmwybL+x0loLABt0gRWw9IaENSw0tNbi+0WUxuQXcyt50VLbj/7/0UYHn
Ic/ccT9Z7AIWvE0f2hcByb392R9dYZnoF7rX/yh7IEOI5dJOTcBYSA2jvq1xx+6bbLBanhEJvViG
BWR38BBplxgINAf29v8g11OsV6+WmZOg71Qgs4ahiyYy2zCzS0+H/7Xt9SMv4q20HVU/i8Yr/nso
R8wJeU215De6H7x4MoNVDQGLMwvps5r9KqWGum6tn6FGsLRzynk7kzhCUa1DgKnWLvwx/dpGmsU3
G+bHnPeFkHyjpFR8ILvFKnEWKdaEAav6z3mANZ0o+PhsaBnthWOMWhC3mCnBFjrMiANRosgttJ8c
OGg1E9sMlNJvFfe1Ay5+UA5KHByOG0HZjsKdgKnTi7CPQxDEqIGtXv7Ik3rpVyqFiWw35x6u6OLL
h+xEDWAmMGyZCzUqiyp4GjqgNJlSXEpNx+PqBMfbZ1LjRNQmgs8/UrA/RCW/o8wIQSr44mVackxu
qcP/6etB5vzXD3Olv7F6AFCiRRGgm4HY/2q1WLO3VFQvUEX2H0SkLttRjiyOq5XGQ+UjToRaG1OK
VhY3qn/MDrCohZ39ONptXvVL/zrhUqGYdgApgx3Z+v9v/lOX7oDY9wmNK6AsAxKikk8WSWCCnABe
yu4bsMdjJlaVmMgFIiOOtxmVvbDZPUv5AFmuy78SOMzjQ86fPGMdYJx5YDM902MJYTnUpjDQyniF
KCrbnSk9kOiAFEd74MOfgv+qgdLjCT3aVnwzc3yWXfI6Bu5Aln8EhSeoS3ftXssxcEtEut/+P11Q
upGjx1gCvVFWMx+rhDOicNAKUZkNZqZgZ1RiCJqVkuJsJtLV69/lwgjH9ryZ7Zik6vxVq2gP4jhC
GiMrOMEJsFvfcX91W9GA4qDsJEw6PTH3BGM78qfmkZ6ANnI4rxbNViVTMR5aaYLWtmvBS7QIVyCI
CTH4B3kvSzKVNfA9nGz+Kztn80rtC4qfbWC2/ZQ1kyLv2189+yrjRrdC1N9DEaDcIGiA+FJOFJC1
I2zWEXJdRAiupT6RLzcYstNWRQBwX9F+GgmEbtJWOjKRPpYdMCfeaSpK7P0aBxHpPtubW9ktrOm5
lF7r7+OCUM3IUwf/suXpxg14+6BAKhkmzmhGLGTBcNopt/e9X+nW5eLDtkORAiloJ17WmeiENZ74
cVQeGsbQLet9HNsusXTMu4qByzS5TdGyITspaXy1esvxzjb31ShhF4rSYs65mmsv4lCashnMul3X
O6ua5lfld2AD/A65o62g+X56V2PsBGoKSITRwRroVU6dDNTIxKrz9qGgZHcEDnb1xyjmk5HJ2h7m
kMR3/asC4shHolnIuFX4InObVK0S7vA7sL0Prup/HpjXMhQQ4QQpUk4bOGP0/DQyF6JeuY3/qnOS
tpxYIWtsgC4DlGssi9GfqOYL49RxeHgXQWAc0D8eSU4b6ZXzo8tPbj2q3DF71rmGULLg3YK+GLgF
IlAPU4omICNtY1j2LXtEqNaoUCHu2P3if7q2Ia8/v5TryS8rLsQOcQxPbpD8op/ELqduSGL4enWS
bzfFHhBCCXDJBaHq5n0tsiWRVH/dKz+DgLFJcCzOVujUfqyYXJpYu9NHYz+PNEwHlsvssfLNj3G0
qXY53bU8dzsng67r9XElOnLkGg3Mr//KHcNVf/BrkqF8UDhGgDkYL7F6XB/rAq9J/Q3uQndD08a8
XNAfocY7TIDbSK1q7i8akn5ObOSfhWom3oPwFoCjsevjLpC0C5buP9NcFE3lXbnqWzvDgKs+EW19
fFEbbvrk429PoGCsCfhNl8az+inaRg16VWwXu5igG2nz+hKYx+oGetEV7cwDNPNSmWlFz+l9O4mZ
J2T5eIMH7i4cRYqVlS9z/iIwv7Oa2i69CyDstoYDVbSpOvCN2hj2JFJaF2Q24fhb3MHGXYb0kAeq
kYnPbjLx6HcFpogHab2UjpePSJjX58orgVMRPTaPQMKpveOmAwg0rZ488DtapO2DEX7liTcso97A
VTYmM2F86lVnk17sS6I5GHncCOJmrsVRhz0jsfrk6csYtEh+rRB5Rr31TFaDzywAColqYTWo8hNh
9/qBfkPrSVwZPwuTR0BtYCsVRiPXyk+JGN4F/EeYmy+Bor2oFKmS4P6O78REnQBy5CE05rFHcL7R
rmIcGmZyodAB6YG3LFuLPN25iDPv09fmiLYngzfP8Ed6Pz+3F2riWV91BNlx5C/0ajx8ZAqdzibM
n3a6alTO5pcZtpks7j7KECMko4Nf+ikv5tzE8TXCIgQ15RKzig01yomXQn9S5BjWYm6v852tKqd7
GKjW9OJx5ftTf6Qqu7zmBxOMjOHJTgl6ncuvtNJSkjuELfEb88S2H7Hgbw+vIgJ4H00HNYOKP75W
GhrqYSBobB9jqhuqZLBC+QOQ90NpwfpRxX4vqCyZ+7DH0d6w02gJE7Eol36VQ+tlX8NsYYB7wqZ+
pHtIaNghLWgPjcJ+n0f5JE4Wu/g5mEZeku9bcrQChRI8DgfJU7P8ubXW0kF7svTQkWJNk/xUxe3L
llrfD2phaEhXfTDaXc48TtclalwJeNjG1ycNDb0Etot0YKxNktHVjRn4AV2+UEhQLsVQDQA706tS
u9O7YR0lRIQ/29bK2BRVATeqYlsAlmk2o+0uLyeKbgxyzAJ8wwM6IM4a7ntIVGSx+vFGqUMzOJr2
Lm6G2ps6+p1XWZ4cBcnJuZWNKg87bWf18KA3zYRahVpfv19SbEYlXJJhdeUnRyuCx159ihumGR5o
+2bkZdzkdB8iJi3DkmoQ3+kyVr+LVCLWGn+njxzZoVaePtaNiiNUiJoG5F0PQ3mY2BYTBc/NboIf
7cytAP+kB6NHNYiwMASqwVorIBFMQ7yBLSeh4jZKTHBHXJnqrbftxQuI3RfZlcOUq0VtIAy5tUpv
9LpeHN07XDGqCxJKz9r3JaCWySS13R1dl4ano+awnsVsmAf8gJh5IGHZknzn82+Ey0TO7wyP4UPg
OHRVk5iUZ3HuGPGjpDneU9l1sBZCMqmzfVkqTNVfKHi7Je5biCSlcuBh4PaaaKWJOk7azzaPrmN1
YDhgF0p503DUL/9UkJmh5kXuqt0eqKY8BIrArsZKZzynSCoFV5nvS6YStF2ibLt3y8eNdBgPDs0x
pdTA93YOO/+oEgIQD180iBdmLVCZdkAyKaCbHoedySbHtvm0DfoT/ztRGSZ/JlFCAojhfcA5Z+od
/3XJxdPmx4F8SiSQFMBlh9NSpjeRzLLSSC0NMTWtuMzp6fp0Q6TD1PPxcmK/2WHdBE1Pn01ZogfU
Xb4Apu+itdBSpc+trsBnDLF6k/req38lwR5AaklKPCbQO6c5nWS5bY4YtpdVLKdbueDJq3P+P4Xq
gQz9IwCG1ygRh1jLi1XpguA1MLLeoCIZve6KPG+x5cqvBdh4vUIuVm0CpiRy9Dc7W7gEvR2OmHGr
0eQ3XQ7QZTNbQ7LmqJmeQPxpYUKlYecsTjYDXTZc6hwFlCEB4m2H/pn6pnsn9jezVv64kIwW6m/n
61YiqqatLxQwj7mpHh327P+KvpGrpc25FRDgw+PPA53NxeEFiq/xluAlWX688Jb8Z4P2GHB1J+C6
Q2pIDKl2J6MAPeEUeDqfVUEh59bWpjI3V9xBDQlcPP9aB9y6FY56G6nBSvlpY/0akLZQqcdJQnBh
nda/tR3u9m44Hmx9cLi4xvWogDJ6Qyp9Pu1YCqC/EsiXyMSuZQ4dmFVKXOkKic4Z4alQX0rgqY52
OdQaZ+guu7FKc44yfpauW+IGvoYsyhp37tuokA4nKlEMLEr3Ziji9JfbvdjzbDMy9mFasN2Qklwo
w0xXs3iAfbC5P28qjljl3hcJelL2Uw7N2Qh9SRNmwTkgUprGzBdwNyw7eYhm2V/MguD60i2H4jKx
wE4Yiaj0Aq+x5BP04rIQnUYbbiXCBH3UpzGg1cf4wnC9iIOrLNNSWtsqUk2BowkHlTNve+ocvfAn
wuc3S9unaq7uS+zMw52uxszy1CHdR+tY5xlmrZu/djK1s+4Unl13SMmBs8LGPXXSiIZ5SszIVuZ0
iYe4SGWIxM5g9AyUTZmvPSJpPbixfT7/OMYVWCNJw27PJhO8fENeD21uRiM6+kxXfe71T92hK3gD
IY7WggTeo3igoWLU0uc5cR0MQqYW98FeYvG3FNYqnIZj7Xfj969QDy/SdejJaY/2H5mzzDCgVbRZ
uCO2mXcFtmV/t/HGnnXpRgCbmNwXb3Agct9uYYl3/NbQPmBt6GHvu1/b9keGDwX6hgQRT4FhxLd6
KSu0tdVmlN3DdFxZ2rK2i3M9NagGlGM4dcNa1mvOEKx6zMC3d83K6clXvPcf/cDAkHG7Ci2iFqpB
xXkoWcunP2s7WZqbC6QkvNQfQBVshqQEQbLeiYdXo4Ys3M7kwuBoygArFZbTWxWr8+NMU004d/aW
RMqDTbSUN3zrryY9SHFKQKplMu3gJ6JHitabKZNRrKg9gpjC2GZvA4giz2mXY/V5x1hQi9SzfWwf
f5J5FaDcOGhie8Y0gSgVaOMRR69dBlbPHECYWxBADhCicrQlzrySp8savIntI7ZjDL9yt8YrV1s8
WpAmehm8fX7T1/TRvL6jVSwUhMJVlLxCj0mhloKABVgTogJfJ8d/LV2xDfJ2OFc+STM2VKZRY1d2
dr/x8zSFzrBSO2WsJGJ2Ssv5LX00f+B6P7tYun5vxpJuQ7eueONSRjJy/4x+Wkagb610sn0x/2ig
ppvjYRvEm4LLiA8jW4bbGfGrQU46fOjXD3ocg2QuyIdCu4FTt3pYW47oNw6IJO2H2TPvHMaQLZtl
8ca68u2CSTKFVE46tn/Hk7hb5acV5evdzcDUltlfNmerlKW8Z3OHlUwJ3GI9PvqvccSU+kxGU4rg
s3OORXp5Jtop9CNwqosGieCmSlP32jnPx8SJZBMnyw6oUYmbOf8TnPSRTgDiHWGctje8sPy0p4XW
H3dbRINWn9nzVG/ZUt4Cd5ZsPXkhrpcg5iiCEdmwnqm5UfuUHMxb9KmR2+pl+B620ysF34ndgBkS
nxr7hqTBrLpHgEcySI++KyALYNtsKxnIYfoVd90HpLYhkPn4VZwtqTcYVFwHZ8rn2fOQW8aEu+zG
f+q/AbYImMMv2a/OVeLWViyA3Pz3bxWBvqq01dZcsZ5gPI1Gc1QRF9tfw+AI02r0Gv2OSAOuJfy6
tjO0eTOvpbBEJZXBf7GHLODJ2jV/zDbEh+VqJo/wbG2qnPhLDidzJ8nmGuV4t7oI6c8U/BKBz5i4
nLm4SE7RBZOmxeGj6Ux1aW3CHdONLzakNfhq78XIllPV/UrfCf1AzdQ8aZHYZCXo8dbjXkhy9Ktn
j+w3Rv2KNiQ0GNTchwF6TONamNuah4fnNOo30Y6emGG9a+vCBOXrhMsSgMwOZPOOUcGPYuRkUl4P
9PsWVPd6x9girvMPO8HPCQMT9r5equ5vdLQEF7VTzLcaHHPYwyHDsVAod3iwlJNlUOBbK7NTwZdM
aeCYEtGtFLcZwer7RKSvq9dZcOWVXpmPs4Lono0E/AXdZByalNchbwg6C5g5j6DLd6YjKcQtZVj2
cdKdxCybRevBbW4f/U210N04NhYZBEbyg5A6FHHR0nN7LsRg5ALSTv2lY6ctaEpDLoRIg2rPqnCs
RhhDEzXdHhL8ifCiOYLXp6FTTeCM7KTr9N9spiq3GdBYe6V2Af3j7nIy5EiuDGSKbJLoiWUfmGWE
m+rNTnyQ4Lh4oasg1OsWO8pJflfPN1i1aUin1A0aZ3QPKUObZCQzkdgsuofjmP4kD2bI2O3riO8O
DACDJmncAs+VMGPQfg3K+oVyub1ovo5IvKFkvo2Pw7xdu8Vu705PXtHivoZWQVpc9l4icNLFo3Vn
y6RGdjyIuj3peqP4Q6+ifbRq9o0dmbmvyUTSHi7MYg/GiN3Vexg430bxp5hvuc0s/G09nGciXrTt
5tjfQBCTkZ5e4rQ2okZpPU8BKWAwUgjpL11PM+mqVSgPQpbtXgx6QQ+AHMcFNOGXXD8C+3aTeQJu
KWpPh62PaQfsOHucLgGjV9qGT5ZS960L6bx2VMULtzA5X/dNTnALG7BdQDoQC6c83X4hE37qPBSK
8nhQ23IdxMs6CEJootVfMFJnKMpDXK6tpSRJgDVf6AL3L8jPaATic7JOOWw6co2LN+VY9ExOcolg
N/SgcLOww/gVdE+a6wViNMLHrQBjBV92V/B5v1NXdfxZi09kdCmpNbmGb5H6MffNnYf89cfLTFTP
dvugTV8c5wYYCxnWg+ph+GJwnJzN2TnBEvc4sHMFWgN5ShgXJkhr9z2tMbQ6aUVo+LkJ8zrvsu3d
uAda4EaXNnqGa1R5wNdRB8GuAOEX7WFdXwZJpc1yxKUOnOnvN5yvUWwVS0vLG2aSQv/B46j/DMiT
77ZAfO1u4HXv977xj90OLK5mKVH3NO6sMesAC5fCg/IhcIQjBqA1nZahA48FTULEclXeJwS1QD3f
TALUveSjsgBcDiimbFwro5XHvDkojP9/mBCSBNxtzIDDkjZzwLkDBoA4zdrFrSd85iDVJan6I4jN
Ta2+T/ho09FE+0nglWEPw2MrYn3YIpQCOyk0ew4JJj1ClwR4iACnff5LlMgP97Ah2G4tNyd1vP+o
eEgYrig+8hdgfdpP7usNgoMcg9k2ohp65iKSWHtwFzDiZSoA8/myx/FmH5wVNs2b8bzRE/X/j653
UQgxGfr4NKIm4nM5xXhqnwPBGfNRdpGkX/baVQ98fQNViwagyWupoGrYFhxXptm1Ys5ca5UFYWPN
QxRjb3nHvC919USjAcDvr4jb+jjqfKxT/bliw0RZ82DuUzDymK0ZnS4HgVeBT+vpWYj+3J/yQIqi
7pv6bU/DlQ1lzVre8VOU22x9GeTyp/Pe31BrIOytX3ehj1L3NLyu/TIpl2g75bE3G/AUnUP35EQY
kO2yjCwc8CdanGhzeIj2lxflXlRGNgla6E6ieFH7vlgM3LbKZTO2PhFIjN2duGZEv7rjIG1WGdfm
eH3nH8XgE7nUxG4TNZXQO7R8eNPjndfxoamMM0A1KexsAgzo5AS99QpeOlPPZxXNFr+oQXvJV1Ew
/ZCw66BiwtLwJskgAl1Q9Ez6dl4G4NJBy5dwWd+F5aHaiWlvNhMomYLQO3lSDRYSpZBNKqyGh8ns
nspsY3wYHlkV/ibUbhV/Cb19orut0xecJVL3axcdyKvEZabKdoANsQmsI2zzBmb6Z19jj4AlbJZR
MDkyLxy3Ma96jLH0uoyxZxa0qneo1naC63paBgil9igmgcqjYtPaDwyndAowBpNsSru/Yfrx1Ofq
7ynxt5W2owJCFUCNQyh7hj90tYJOB7cPMi9Sm5zXkbmfX9LRg+DXxwuRhYB1QHqa0YfOhlSMPcBK
10pXNUTaUKqBoJWtnQ3eN1gnop+7EZp8DSkuG8kOZrRTTQieffAkwV7QoWvR3bjdKQmNy+wr2PdL
+wpc+kwqTwfnctMO03dSQmgLCV0o8FH1YyXbIgvAyWJCU3w4wIYgMll2n2eHi9Jfg2CeWu8SIJ6U
L9zopdBASH62j5UcZAQGmuBfn9xQYQppQ+X9nEobeZ/R4vRAw/6ZFUIQTZva/NKOVPrNcr9ZemgZ
ipQczyyIrnxR67dpi6GrN9cBl1Xz7ImUIR8EsmlEWUR09VLdcc6BNbRZTjmsc+rzsjs+/Kshy4M6
EoMOsRkNvZki2lwWWVJH2EGy60HkcFRW/fpAHv3XpIREOtNYnjriqzLa+jmbzWEJbFgPeWovUeUH
iSl10b0FdFhnMcOEPjBkQwakHjKfFmi1VruEy7CkU/pSTL5twDv0Bo1rA2Jy519znZB5YPTle3XF
UR1LV/rOgXOGVk1d0WpTa/ecbxdnI/blbFpPsp811nugeH0cNKWteqzQ6pPNhgH9+2qXRJFfvZxq
AiCx9yP4wAH09SCmMrdVvcmhlKgdPrntH8Pf1Z7cfZzV2ouajEiHNMsrzj4KkTt5b+p/ZdCgyncH
FN+18HMTyOZ5lnhR8EVERL68ivxlLxJloOm/7RXjoAEINeae1lBKU8pZ+If5kL1Jz8ByynFjPVfc
r50D/ypxlfxFKj6ttIGNgwLKppoJIchSdzr/PTmTpGFgZklhJdc+ics7e9VAQpUYEYp0PutIIUJX
nB2KfRRDITXC52aKz2j4omBFhIOYfHQXonPtlCCKzGpwFiHBQ4cOOGVKaxyhk7wutwxEhRGaTS1y
WmNQKZhgzxqj4+m48Q1mn9MJtVR1e5lTZeiyaAZ0CEOuEhrJVpU2OTWdGfvGVrBwg7gL5R3x4pL4
4mwLEdaMWhQ/VoZHdqDTxreWNpd8gy6TZo7/RPzWz5+9g3ezESw0zMlF00LybSUW238UlKNZZGaB
kvxZ1cHZLa4U9y7llr/PZdS7wJNEOx9THDdN2E+MyxO9kYO6wasBlFyi7xVTHPNtWZJxJIRrSTdY
K1PBARKsYdhpMRzlJYPre3W4MtxtfECeW0F1NpUMJ8iXu1y4TDP3YGX8Qe1Sb6hylaV/TACejYUP
TSFewpWSd+XbBReFZe8T2o5RcbC112w20oTAP3ZL8jthNmqqiwyrjr4/qKmQnBtTJ/bQ/uJqGWGR
kahr+jtoyoH0w1SlRZWymLcmhJtWw+lMNtpaVzhJwxAJAlU3Bu9TtgA99B6dVl4Wbud6DiBaKqtM
+CqYQtNocetibth9jR7fwhWHDBbmnSXkoaZ4quhecAKq2yystzJsGB9DernwRrd3h3t7D1LNqr8w
QMWBw8dGRKZDzM2vqy8xys9nfcTOW8HjTpbwlK5kIIvBqwPcR4O+vPfzVBeRL46w+zCRy4/TwVmC
c/oYCQjHiKOmm5bS2c6l6pBzfhdO2z6koJ0+W5K3msNfTSvO+Fz72Y3W754COtPBU8V1G8hpQnOk
88YJWMEq73UjxyKmhR+WK/8T/jcpbw2fUgzvO/mpWciOxC8aMRHW6XAeHXHuk4btOoI/FT1YB5qb
dvMv+rlUJvjywE94lcS9TV6tVWTv0tWtISSBXVNi8Mc8N1tfa6GqQiw3IVta5+d1bUPOS3c8XaV2
Z7eOwVEvNTENncUYYwIsQO75+m4xxXuXdwjwY0v6s3Rdk8nnSJhJpwcAF6zQL+gbAGZUYGvzCp0O
qB9gwkAZcYV9EYG+PJitYOJn+U/5vHX/moXHXw3AG3ktyUm1lkOjFq+0bJiuH/0CFhaiX6dG2R+B
GkWU4Kzwdqwaz1QiPdIEFqJNIZti4+Dk+xgViZwEkmb3DYhfDb/0Yn7UPQXh5Kmb6Rt1osVI7+Z+
L6QUZzG/Tf8IuXtUJ4crZPe0wmSHWlfLtcWl8r86PurRqjdGoWNXYq+U94LfSm0LesjatNMbqWK5
DWpTBP6G/z89uTBArm/eUVw6iQ5gQeCP9g4cmejbqmET52YnsGYl7rAvAsC64CTQroRk54VxcSub
auvqzs+yy5plHPVK0ikWHxS6oM2STQSB6iERhm2nUwHv9vQVP2A+thCY01WkldZ9p127D3eHjrlb
m66ATtoEChCYnSGo0vUgWy3EGcwfw0ri9yM/NBYsU61vK54Ua01wFSYTP0mdRtRb/mbeijmfw8YM
ThvcQ9R1kBQvDdZNGoZ5y/thKJusXrujAWLNKc5BUKRlHtYH8L17ZL3p2OIHHS5NWF4lpNMP1WWk
W54wTFlOtmlX3zprZGMeJqtmel0AlK03fCgAdR5OVKcGs8f5mYihQ3TtqVuEZokXI0o55O8zjHrB
9hC3lFUMgGMO5pWbybA2wwAY4oLJ3vogIDDDKK1IoGVd1tL4EJoFAS8eq9c0UIhKVpJnQiEuAtB5
foCrh8u1lfSm7W7Gxe3k8DWeueKtNhzKMIlDraLJGEK3VuEmAT3gPj4oHDijwWKqxH/6PqC2QQWR
voEaRkv1hPVlByfzBPlzxwcqxJKIjTo0YEVQ6VgMneMFUzwuxpfSS4xkqnUmWudaxHNbwxfHJ11n
PBw+/DSCy0Q3NWOwaaejbIXen4IjGfGUqORHyiuBSaM5GTPWNULEt02EmVcR2S9XggE28ePiwYJ3
EloydeQMTzUrJGPO5n7r2EA4rhBzG+IK/Yzhg90Ofb/W7OpPqIdsXv9hfT+eC2SpQ4ShAi8HOmTh
Ot0uKomfc1kCdQTTl5uPuwDJhvntzFVZLcbgJtzs7E7CgkWcmp2JT6PMi/+6pNHQ/j1GQqWFrhfo
8b2sHeBahfOrvIa/qNObgkK2qV+HUBfiiSswNR5dC8V525U62t3wKrWLln0mNDY2MrsE0XohciQg
nohXqaaogeU7rmrOmXWyzkVPwg/hlmT5+gE85M39FpAn1nsheiVzgiaWHbKXyNy8W0IJNL6lNlAG
DQYqpMA9dZolgc2863u1//3Llnk8oyfMy8TTDTLgT8ejfUhHkSkai1p7ZVX6X7Zzo2OtYS84zzPX
nPN2TduDeI4t8SQhEAf+04q+dROWpJ6L50IaN5H12n9yTgDM3c2/PQ/ZXvDgv9dsG9Q2QiDvGpZT
vDiQTXxd35yKz7ZZ4hq3xKPfeUuHtsh6u55EltWjZghVzejD0crK87Q+XIHMkg3vWkfnX/XsDgYd
9Y/HrDfQJvUCf+LCJZZoFc9e7Gxbjd3eHIN7oDHRh63lkc2DyUba0xc+nYlAyQhCmTSINGOKgUog
pCf3c7HWYUhz7sJpS8NmhDkaBOEx6GfIxeALFANv5jbMJGqGMkswlW+NUxLpUb3NKxLvF9sMShqX
Q+Vf4Kqf/jDv3mLtIXRm3Jex3xK5B7oJF5mDG4ITdoPnV8f/XysYrLHRgWe1XdV2aE4eSMsfLu2Z
oYgcXPx2fTCYzSwFVHchPUGA0yUhcIjjSSZZbDT71Wr4Hn74+7SaAbXENzfLF3Cjenap2UfIB5sK
zlYJy9Bh6NUzk+t7DiSRuKDx++Knjsgzm/GzyGMd+p0K9XlgsTmMKz7EbVawmupYqqXaR4IfcyJc
bhFhhzgGJGnqy8IAZcOKUny07SKBsnlreo4JvSqPv/9HHTrWC1TgFfIE3DXjlwN6wOg7StTKozI8
c6mrwM3s51tfz0whvOPShCO2Q7dUOnG8gaN4IJe09zM56/jQnHoNt7unrWtDyKFMuwj7+CxftlPS
SH2PVCcBIDugZKwh3OIl1WokVfuiRkl1yvER4o39X6koD38QRCdxP6TRkKP2EJYqSL4Rr+ZdTx1O
8qVeby1Oa6yfgjyGNVqZE3WZfHQUalb04pm+N9/J0GXgIIWw/g9O3haxQrliILu3tMI7qjtaNMrG
fbMRO3cI+MpcS2+vYlVUYl4wf8sXByPtPbkVjZdIbbrsyDv3sd6MXX/rTf2UJ8xTSwYEQBm4bhZ6
aKHJPQen2Ou/R/YnKZcOHK1xsjAqoor+BWHlZBtTUYzz4YXITI4tGieJZRpt4LN4SAOelcJCdazj
PCqDC/H6yP+CD40o30BvZHzwc1R0E1l7s9EOZuhy0beesIu33kNP20ALGjKbmUmX/h7RX4JHo3hs
pwGjBRYdlOO/+062iF2/rNBKAssYVzf3jzRYHcIAmNphtxjHlNmI+6LCNvZARjrTi2/+S2sAFeJ8
F1j5RREAeuyL8DNMVHSZMpV2uf2C0V2QacXWqT7PWIWco76HiEt/fWV2iysIjHMO1uYlScbqhDdw
0JAIBvp/wZ7/LBMM339zSvdUygOKzztw1QnOgpYTzEXHqiTB7YZG0iZOAyOZ/GDmI/RhnNwPUHZj
Rvn0Cquh9XqIMZy1A0vvOQx5Hbi54Z50V1U12M+C7SMLm3g7+JsSuOmMAy3sQt/qO/+z9jqC3qLk
mJVnnEv57KoPKr77xktlyJrIx8r33xhGxhvyIzruuUBNdTE+O5liev7Kc9+35CBTKRWC4Tawg7gt
HaRx4R6QN+g6mK0PmOBYTU6ZcAtYTtBlC3FdSvtsAgUnRXp0ChqntDdn88xdgSx1oPO2rxMPmWcv
q2iMSEOmR41iVqGz2l65xYi1IdxHWL1bGYKrR/K2zmq85Czq6+ZxkaUg05OT6riumyiG+r8tYWVp
c+JfhWFtn/6WdK7biHpIizfQgPTISq2DQPmvDuo3eclUixcAG1UsZZgxnRx3mJhriaQWeTcF+Odv
jTofrj43Le6r6fI9fFhncA0o0BNzMxZZB5z5/SLOOk2xU+RynLQckKpSCm98h/D+zPA/LhX+bdj1
n0AhD5MEnAbg4rHqrn8z6bjoFdfWNjBc0MMdXMnXnYPkbNPKMDz/7p5EkRjvaZ3Wgb+kFkfmzEj2
iqoMd4sLvofKCwZH11bij2sTohUXPW0jUKeTKTW0VDYv5KG/wbM9S158m16C60YLem7MHur0r55A
t7xHwJRv0qakWn7muSsnnOnqCtqZoIpWCT+uJlJAus0oYTIK7M84uHv+ymJIdqm7oB8wYgQeiUva
ajnaeZbWqruQ/JKb9AGHpi5pMCH/XoIT2i+KPNJJro6WSji4CMgSywlZC/rkEQ0QjEkADDwNMy1K
CO8kkeaQheKxHYZomE6d3Vp5+cx7+zUzkoI/odpZbX2yfTzPIlTGF5ROGCvhM7YOJdeXniLU0Dtq
UQdO8sGAOPmAY3u67DA6l38CInrC8mPiP92vrbHPdr5Du27OyWPkMNwiDakmiWOfhFED2QW8iW5Z
ivAM/4/FJiKciyaFaRrF5Znvx4Lq9cw7YKgSaR/dEQ8ZqaF0MPfIGfY35ZnplZvUUI8d3ZQ9FPHc
pJ4hZO3jnG40e+7CkLOezTW1xVff3vtHOBq1RVm0SVhoI3x77mdNYe3MxFRSmrHU9LEVxiXyyPMu
paWZ1pi/AocyHbrThalN3eXoZkcJoN8OHDMWQrZYoCkO2/JU3fBkWyYYX12jmBSTZRVAuFMaWAn+
5I1atpkJke7X30teDgt28nFFlzDHbMePaIVfcYNbYnX1EV81+G4fEnDC4oXlg8Xv+8NRllJXtvEr
ZWsa0l22kp1R8zj/o7Bl8Qcj2pS1Re8A9m6Wd00Kkf3AbbqyDpeYNYbv6OI3fVK28oVPj3EXsfqc
Snu5Z9LKVneIrVM4/tc0SRDiMefK+rk0Q+YJnsmNzUsqlO7I5ZblDMzCWTmJkQpeuBEsu4TVQCi6
0SD3MXYjBlRYDVxtEBA0+kYjeaUjdS5mJZPx3pMH+8Max/WTvV+cfkQ4LzNL+7XmAIStcg/6qKoI
Fl6C6M1qV69Re7/LSgVbK0aN9jyEzwR8O/R0cjBqbcVhuMpnnLd3aseOnLeUqp7nCgQHhplSbDg5
TO7P4be2z4rlGkaEJSpipjC6T8I6gowVfSVPiPkPB//cSOe7F+lMHJaQPBkM6BVPPeXcZP5tf/Rw
uh6+7kqcH/XSpq+kxF3GNNkKaL2sflURkyXNoJl/Os1F5yE2PlYy7Sqc4olUAKPdZepjTS8Ba+SY
np1vcaspEKu1d/nSchbiI4r8r4wm0dXoi22fEJX353bOcD0e0h/STU4vGb2VgKsRpLsD4sGb26rS
CyxcPFhwXYRQ0JQal0z2Y2j6JUIGrbZkwducARp0MTq7wL9+CZV9ScStf84EuMRQkJDeU/eq38Nu
sxetaPJxBN/byKSiaCoz0COiRRfEqLLDb3FnQYeSmsnP+W+M10Tvek+Xzsv9IpgxBoyLVKN7Ktsi
FP1Nz7zUy0ppzxmwcezYeUx9IHpCKjn8/k320p9kfPvgQ+UkIWkx/0O5vgbqBxuBPb1GAe5PzhqJ
Iu69gRN/yroNEcs8njN6vGZSqu7DED2O1fBmtFVb5LuuuQHMPhpa21eH6CHoTU6EctGcJz7d4qrR
7reJVCsZL3KxGhq+CM19DQMJMi87FEkSL77OMmcyFn/pO8A/q3ywiARXosd6g+Ooghc/am129mw7
2dDzVmA0PnPAgGZjEZ8TJAPylUOJJYLmbcaNCZvmnILnEs5nrVFhQ8bfZqJzNbDE5uvBbVRk19sg
EpIoZ3aXeujxcRVPLV+bvhO+av5fhBpJ++SgqSVZioMS7HFNZOq+8UdwEXsUjW6Osg/1dA5lHUj4
xWQSPqsNzV/N8A57R7VOa4zwejWRybgRPi+RE36aRxTirtHOMMfAigcz1y0oHoYsR/R4xtOI4IE6
0nrLrpbjHV4E0i4ysJpXL20aRc94w9UFm07RUo6cjrvu+JtR4VwEYKbTmtWFokgwk9qfgr+Ebyzs
0TfMeehY7jiWQxy9OmQ/iASd0uZhdatMdNvmkWVzX3FgrCR3y6tQPSOEcaPhuJoVk3BGcwidTPre
Pd9aSE5Ig6MciqjriLDWsi10pM+jZRe/yxmlC0D/Et852EWk2czwx2X2Ln6lvBD3FC1kkek/Tx9w
AekJVupLZPwPm7GqV0ZoDPrvuskONBhkmpoYm40X+UvdqxMUsI7d3a/YOconO3McIWQ5n/MF+RN0
dcok/LE7m9fmjnvIRBIwtjVRdhnBycSjwpn79tUn7x+sC5qai3qsIDTsN7HQIuT1mJI+syPjSgUs
C49pfU1UvcrnXciHgFIM+cADB/FcgalklgRINMsNnx2+m5+q+ucJPLKvLhcgrpdaW4NvxG258m/x
XIpl8KKU5UL4+4/yDRHx8tV3EcHcFD6IdfXaVqU5UqcF7L21i2iiDzjYk+OjKrxiueITS1THijEe
Q1HpHw9GoccSAxuO2sKhJ1z98XHXy0EnG8cRE/e3AC+JgVIsZq+iXDgDMsZHi3qcixo0TL1pTc0I
znW9dXJrdeMmgmNEdn1OpU5tVZx1GLcfDNLobqbiAuiRXAydfMp7TidcwcFHg/LzRzFsH5r+Uisv
HmD6VRAtS0gCfDDjMojRnnEQwNcVGyGjs3dZ8PbG1RT5tlLqeeSv4D2HHNW0bxePtTbIsLb3+zVO
eqqOYfQ1XlK/9RVGqXsEDuTYbuUTeqfsn6oM4Fdo2y1W2BbabTkemY3M5ZffNBP1Sc86BMTXQNr+
N44fBARpz3quFZysD1UZElLAvZ9aPgn86DsG/URP/yJFqHnfy7/GwwonYDokMA4B6Ns+/ofX5G3k
Pj8dlErvxakkxHxcYkCfflYL+c9XAi8jj+mawaNqGiR+7glRgk2MAUU3N/6c48UZYZ0R8rKW3ZK1
a60iiz/SunVUJzJ0hIQ1f4KHLSPWggtLJ8PQB9cMmTKRRQNRzteI62WBV9I6NhK5Wip4s74BX9b1
/qA6lYaOLxnulmjstP2EJMDZeiMyo/7tkRJafmxFtV3hBJ6EeM3OoffVzBzlMbGZ4mVsa89cjJKk
47qLebJZuKBOLhARbRZP1ZPHsAulx6j6ZYH2n21mLfC0so70qVd+kZQEqp/zcgrh5iXYo3Tyf+7m
K6r6jBGAlmk8lBRPrqnBPbXLtgGf71K/4WmOp5leHdQ689cDsEiD5nJHbpFvrQTTRiptVxiK+mdn
k/2cTyQMZ4CKlnygXmxV/AhkcfBnCv70q2sg/SGib/VnDzSZOJ4btrKsEeUba8wDboz0lZyPF2J+
s5cMC/n6g5oC1bSm21RhBvJzrqw8JeHRjrTr+aw1oVjgDS0UR14nvkTnd1wnv8W5TiGt1qJavExT
+denMkfiZGGFmTN0UyPpqayLTcT0p5G5wLiOLs8iYQZJEI6EFqH3zgVlMPdDwOkAljODtLdAkLS7
BYAc+C4YJs22y9zBxEyorLwiFD9zhIPvg33RXP0+6+ykgewLpwDX8Gqgv33lNY1cc4HWngxPJ8/s
Pdi7WobNjrsNFvIaJRLPWkI3qEgdbiVyB8F2b8AzjuiU1WNcny8MPovaOCc1RJ6UMoRAgyH5BRhC
EpOCuAzqQa+yJPm8fRa2WJUXJ/4n70l25MynTWQap+M+kcwACkbRMopcbkhsMOj/EqtTs80eAQOv
H3Hgtt4C2UUM1n6vugcTcNokIKSQ1AZqFv5yzAROj64F7P18LzUqeeoc87QpiZjU15hE06dAZ07F
k4lT2Th0Xk2eU3VpGBYdys5b/MCZJQ9Qm5p94KhtzoHKnrj/7Uh6RSTN8+YoUXpZmU9DEYuX3IeJ
hRV3sqyrgtNxAv4HbAgl4MgfynWVayZHspHwgx3P/DzP177+gMm6Zp0KO8N8F0Y0N3U21AhkhqnK
+SJLk/5LOPMmnYrBp6q7pgtVoMsq5RaIq9GzjJKXLsFSfXvA/O8R4Cdg+CdVl/noWv1B35okBQtg
kM7JvxYvW3+eNravevQRm6RiNxDXoBiiwwNGRV+MjODdlNwk92R1yW2P/vjp011iXygGDEC51Q/E
VLotMdv32idZOTk5cZ2TKHCJjtQGF4YmwTnU8JIz8/O5lcY2O7ZNgpJ/l3OuBezQ2q2ocpgZDjtC
AxQw1V7TgeVOkhtJPsclwNUfTIviOH8/EWZpmqovmKUTq8lFjvHbpf2EnjdkXk47kxKaRyFrsxdV
s0biYkB8XuvnK6bBLsbeiXCVnEhybLHArTjlIJYCwrGXvX8b7w41W1zhpAXi4ruqm+scihOJ06lW
9JH1o3eObVn7ZGYe4LNb7CEvqKMLa0BBpl+hylvZd7VxTfylTtMEu1/ThKJy8fginGADfAiVeftK
n0hVnsPh5Lmy3h16dliFOCD1Hp/ecQbC97B0JsrZHFgF0MjacTBeEzpduQoVGHuP20VMxUE5cig2
72nyzkCVXTtloT1S8hrhdEsfBe2jO7/bvZCsIjAUCciw+9BM7fCAvC8n85MelAr/5kjSuJtmtq2Z
LP4dm1RPbs8QQH27/oVf0jry+u+/u0Pudermu6htUEpNsa6NicWyuV1kap4Eqn5tlvsWUfi7TOrn
+at2fpajXCjS8gS5DyZ2HVZFaRkGIGQR7XR9PighuFmQurDq7muryjlAZl+/3l4VQyzIKp8Bd9fV
W5Et+n2GMlWOwDvzEtb2t7v96EDBSDHfK/kCTnVwrnOQI0g7zEkIuSlFgyzH4hC1b6rSxEWFUe1T
x8KNIDSl5HCqTOuE/gMPHzkVrmXrCyRINJ0vd4kzOWXAunJdV1gRWB89NPWfPik0lHRozFm6zWUG
jkX5lhhglkVN/QOgKIrkKA1VsF//28emLntXBZeKjfFr06xS9BoMZlD4wQlJM2bwbTcQt56FECFj
KQYofuZ0HPFzOzMRWXgZWHOjDM95knOxLl1lWjTiXHVxsGpIxnm2Au8bHQVh9OXaOiXy+jqnEGws
fktBbWm/DtMpVJuwnOIV9QHpBUetWUFuYb8Byv3OWRAqDqXt2L2yIjKEclmt9a3f/EAfVArv6gE2
QgzNc9vm7ckV/AVVdIYV8FLzIoZZBJJnIV3HMWpgKGifbdIXQ+HXbf6CFEOo87zJvFie8ungc9ok
A4NwRDw4mRsYAvyBX+2G4jsUT20Cu926uf6/GDc29EE8q+cVxztqYkNO87HEL3E/dIkLq7jY4ZvW
8AoIDuV/7tqiy3UwIR3roOBoqNQhzHep9WmitwyChnYvuzF8CBKoDF9FZ3+8t8QsqjrQHxfai4hG
NXudgULLQZmdDdIMDcTOaJnWDeZatb1kkaE/dpxvHcnaNlNl4IBVYLI/UWBjQfugdml34N2pdpCi
Wvi+8xwv54TFDlK2+pKK4xNrqv3wzpFy3a4hYKzjgGiIisbt3tlcWC56bO0vuRG8f4ao4SF0e0wx
uOm4a+4KI5Ka38dqgORsJT2awr5MvJar8BCsi+nOkD0lAYtbIwZHv0tzT4I1A/uAO445Kje/BTr9
aYXOBvtBIOxCDKw0MfyxU/206xkNGjzhFVOm+YxoMHF1xAbfusrHp98hWJbMkODQKMW8uWHEIqks
dRPd6RVgLMb7AQZFOSU5sZObnhIGgzuXTEg130kq5xNKOuv35O2S/fbPw4gW6A28eR8qTOLfm20L
96aS4pk+Utv0sDiNWoX+v7i3Kc8KYLElEl1V8TV3lD3u4QuuE8DxGEIedP71NfetSjAZrnybh0ZD
QdrSKVHAfmUPsGZy6wQTB8PZJvjrE3m2rzwUuGHaxzDEdfDCRTogK95YVWEOR+pUHl5zG5ibRsIA
pvuNARyo8oRHcpFfqSvQHewfQHTl49FTtnhGJ1o6I9YQAFxzjYg3P7B0Fk0tKyvnLqKe/+3d4Q8p
dehcsSw463nNHs6RMhdy8nnKK4UMwFmr4he+x66TMmIFbJfS8NXkZcnwq0szs5EaqqCz5Ra9u+1W
2cCvZrGfljSqJGjYFd16gMZ8fkiOgr2AjQfPGiQioVqr+FNe+nilWrZpbKCt6KWuRcMqvaHRhuS2
F62mztRsH3ZGRshATu8swFbUzJ+w8T/byEKcYZLo05DVSVQ6lkMOJkCMaarVzJEidtxpkIveQoj3
roJOsexbK9ScxuCEANPCaGXHPZCWiWWrfj9Ei8Fzh3cFs+Jc3p11t9JG46NJuqGGDF657YIMmu64
erbGa/qYvTgLKbH123K4Xz/eHFRRheoAoT05aADRZ0dkZ5Ovg/TbyXwr1YeouFsu3jN7pizJ6ED7
NbC/p8ViPW8l+xnLIfEJpN5t6yyh7mXxCVscQ6O424E1ff4ZxgHqeGgxpIBU5qPg449uKa2mFAEW
/2cg4f3aUL00WqhgJYT2bytdXnWPFNNy+GQ2mARtxh0xheVr1RNtag+E0R0bE6IFZB6yjVYsAzZ+
LQ2fztcQzaEHg5laS77EWfAoBDsvOHztzqrfs924tlTroR6aePGyKed1RdzONhGQkG5THTyfq2QO
/PmDqU7QbtzhkF3uNNw7Gn3veru0lPibjb6S7DciUdbnHOPc/HaeRDKmN2oote7shDyzwIqkls1z
mahi3D4tYVlt7EeDAgHJomI3IIRZEWtlPMttzTC45paVmUpqR6wnrFYI3S5r7DEnEvdWik8dOMgj
Y72dyRKXFP7069aBEiNR1ETTWrpPsRkyjVucIROKGL3VrXBgl8RhpWpmv0tzBgwCDy3HOUwaSNy8
1OdFIDGareDMM4pOtD96AI2CQR3ZLPJIcbsvXO3GSxOw15IP3N8T3EZyy8zddSU+ftkgrVgvfqgq
kHjk0jkjKn0jejGFJKb4W7YgMm9YcgSOK/LKa8L7pyMn8yZpc1QImVWR80WuS5+oRUbTj0tvlvEE
nEyKXyegPgwkJ4Lss0rkTyhtV8RMP0vwYYfxoB5vgd6tFJmxjumJdEyTmTUrkqZXzPBMklxwGV9R
rWrDfOAJJroEU5T4MKKrh3GDv5iKjqtUJLPIT2ahPu3fcSolzmrYnBENrUsn/pvSqPlHKC4ipI4n
fbph/5T++saCKx4Vk+QBNLY9hlNx2VsFyzbmVJ6Feon+1/YmYjXYUEFVShv4ElkPWXDHIyJiEK/M
mSur+d6SB023TpqGjFot/QzxbioXih35QbhDy2cMqaggQ89UbG800zYqsAOMeEifKZc4dJ2MuTVc
qhom2pHEBDvSy8zA2nm+8rqpaaDb3eLEhTDxYuuBlMvmApphUcxavy+BHoHq8XD4dHjVtGhBXxwR
Zfeb6mULnMuRrYFk4BXJLUhsM8R5RzawuDFxsRicSPe78SKgbkqOiNW2Ug2A3VigYGpQnRJG0kNj
yfjP6uSXfoF1mHDhOKKDnU5LGU1J5eO3Rh7g72G/wr4nWf8iQfcMdh7ZzRjbMb2iLAMERPDeYjJP
tIvBggO8RG7vqjpapJBE14eo6Fda2kI/8FqqhEK2985JqU43lAJBvmJJ+IOZ9Ba8qDE4pyhnT84f
//ZyCiwZ8b0bgwdDoxjb3dHqRhW9x/GOdmmbiUVoNX5kUeitIV20mfP/w3XLQ6qktXDWOBXrCRBf
JYifTUknPW1j3YW7fEPAOrDZMFL5NvY9vnuxu44+hTWLR1mns0b51xSobeTYMj1pC6gs6LNXVMwP
1TYGLxs9W8dEgGjdY8GOiXSffzk2fWB/CqQDfbXytLxy91M7fIRlM0zxB5w+iPtm5juc2pyj5WbT
3Qy/3XsQxDmVJJXmjIoIAbOr5o4RRK8QmM3u6O5DtkShLg7wCGCotnBt9J1NLypKinzpIR1NRdCJ
IhWeHMBxq4ym19c9RZmAYYGZdK5CTvbClhJN9BRu4JS7+ZrQSkOsHNTpz6O5vQQwudsD3fIEWg9/
uHW8+mYR4tYxheOCVMSXyk3LmHkxKPb71zRT3FCe6Dgtg31q+WA9wWB2I2BeVnxrxmIky0Y7JD3y
IaXLE8peSbKeTPbFI54YitlZ0U2/yhpIF4CgzF+UaPVk4IKK4IZhV/swKNWt+mYz0zjjfZb79PFb
sbDLwjLhNSVYF98henkK/tjyF5ResOZt8kaKTzpFCnN4SfpP2RMiqt5+Yd0qmp+Xh3X+ok1FDnV+
0J4flNEmAaDrJj7e1kEVK21aRC6VqEKqheaDuIlFKtQclikIKzMgbfANZdDYp/q0qpNz5fXWQVoD
YnEX170mf1Ph0bV7Yf4tYWwvw3Ic5J/i9FSdGKnCcCyw+d4fJ9T+vMNBwwn5DKHI9dAfg9XI+ugC
mhGjRcs/XJBF8AtC9Jk8i2qH8gmDuqLhqCzJ/mohQ5et86ZGaAoRktpQBoo8JO0ZpmTFeNmv7tN5
qa8gmdaD1KbZJ6HVwfUxOeUPAXH+ZKzISKkrCGZk5mTgyUeSB+DmzWa43xuSQM5D69b5fU5jXPlj
yXz2DPtNiI3oqpdfa3Pa0qDlP7Lt7Ml/Js7UsOBdYncty82MecgP1J2AgwwGEiPoqEWjDmQPJBfy
Ra1B29h68//WaAQyFGSIjonSwG50rgaCMNNmuy7ZM2Q+JJYCbVamkmhPDnKeNxHlT+7yGZIjVqwn
yoVfXICHCs2N1kgI2ETbUwKcAOtJ1lHQgWg6EEFhH0KF77WINeY+zToeJsYtL7ggYNDJou30uClV
cFhJekyWFKnCKjDwhKGE1pyG6h7+J9A91N0/nBROCxhslLUOQaqbRFZuV7duh52cVqJIUsKHaurr
xC907GRdPPMDh1SerDhaWRIoy34KT16kaSdiBsXjIyUQiaEnpeUi3ZiZAvb74a71JJ7XkQSNxz9O
ZDFS/RAVhGTnwqkXh11/QZpIBZGYZz00gGvXxO7a/8bdak4p+h2K91RjpEugrO2CddfqSe3OnMyo
LtEV6S7qDXMyQRtON0Yy1AuVxve145Xpd9ULEQ8+iVbQcKOocblSTZ8gnlHh5ohJhVP/OlakldV7
k0hGlxsROqy7nrZPYoaCBwRW7h9mE9ZsqSqCqHCm0j8mjdMI+91Xzc9MeLzdURBMLgQedKo2orW7
HFkhBHP6jyONvKNskk63/mz5VekTLPXEl2JhCIw8eQpO7ExsZLIlURz+SPrEqADTyacW3IYWfH5J
UODjoatBy+98hCwvE3L2VcdEtMlfa0hMPzzFiBrpH+x53IFBuK7P6lYRJ0+NrmTx5oN/iSdGKG+x
P4/cdpJU2Ob28UFEdNtW4RrErue3bJqHjEoQsgZTn+ZHVGl17f49A4b71Oo3qBhlBciDyetsiILT
4fIxlN61IWc5aCb8M3ui4H03PNwHqP/ndCbo7VsrE3/m/sL743hv3W0Bdy1L9M+ej4cAPhBd2IL9
DZ750OS7CvqZohYIJGLh/d4auFbmwOD10mdyvkudurbN7GY+o+SifIXArsyIcUZcgPwOQoVOR3rv
QDmAqN6qS6k2mC6z7bInMWDcnlX8e2gyADEodZJfr336LrezMSLrOHv2U0a4ZBGgmkyIL+VGzVwp
cLoiSVxc9Qhd7suhdIuR3LSicyJYpVNuqfore97EguUo4UZf/RY8UtOJ8QOB1rKpHcbipX1yCaVb
+cQFXbFpZH6k2EnKnEaXRZPbzivPFSYleubiuWcgnQs5NOyj2qEH32ccbqnZQc0oAFFd1wVRcM35
lqbSKbS0DkxA/GFPtizI7N9xiOYJVd6vDgPb4KLgJiTkRxlGzXpq46GF0iQ0MhcEkXdQda2OfzjC
75YLr+fFlovLwY8VpXRvGYIYqnRahq1R9QHOCbi2UMJnWwn1IfJGmIL900BuaNxZZJZmdNQ+yZtZ
kYl1WiOFq8p/BW0k9o98k3L0Eao/iOP6dPgNzLnxgVVtF9cjtgZh1Q4DBMhWgl0PVapyEK3QjPIv
UUPb2cmZ+a7ucLPxQ6lB2QZ1b51o3w3u6zjFCB5RWOCurlHNHwWsOgprpbzRA52zCuGsKMzjY7mu
KeRn3e3UoMFbkJ8IdIQDPIuifHCNfedff4TDPYRteNqNfq7mVMzBuDZZ6br7PR7JqjNCG7SaImgY
CCOfTfEISTkr6I0rmgakzoGT3mfaAsbn0AhiAwTtTqM7ul1YyyG58Fy57EIwjykKLS62VtGpbFM0
s742Vj7CSd0qaSsKFgT3IoZ+gEhsHctQ+tzrF5GnHv1JCxZoUTi3sOheUSDVCxnVWPVoMXSYMXQT
lSM3sbCZbUxi1I3bqOYJk0aWFNY3F5CxKPCl4zM0y9bAk/AP5I9wV1MiAqcfZO1gTKhJdaOM1HDZ
CdL0KS7ru99nUZm00EcbwG5HoPbaiLo/kUzU1lmOzaiY0PbcsWL4VP180SuFwFW1WbVvpZhz24hv
iBaJYARsjHh4FAE3yLsBvv5+Mf/QbSrjT5z43m9YnA91FfQoHBSHY5qTzYIl+3UOLQCrcVsCHKlg
db8ZSOnP+AW1RK35+9X1Ue7lWynbJEfnHBkYfDGKDbqyC4Vr2dNP9uholiafV58M0L/ehfHHFLag
ujVeTaqv9J3v7tzEaTy5IcHZHJ0lmmb6LNV+aWI7KspfA9TI+Z/J6z3D3lrMKMUHJG1Fk0Z11MwT
5J4CAOyFvjjhpntXhSk1MthdA8yPcY5d1IFhB+WGRMabCQLo+4U+J7BVXgBAZbrxIISbrsnInPgl
LmUKBfjLguM6/8L+yBolwTLr3tJvCL2KRv3PLRJ4h39O/I2NS4KjxFrVeCXtVpfsIP0vyEzvEYJ8
FVG4/4zMrusSUohQ+QX4YN3O7iyovQnubQeXY0AjdNB9nE6U5LfjrPPuifZJ8GDgwpI9+JUB9YBW
y5qQVxJtLBFr6KLPjpkyc9qu1nwcbsNEaaqUsO6pgeVHsOJPn+IZ1AsfL1FyTDidzczqgRGCDGO3
njzlo+d14h4+WUES2tBPjQHE/IN3XiDePVejTngjNGXjXnH/NosTF2JiERA6CH1WusXIp3sBG3mr
mUxtq/RPtCRBrCKBxKXoUMA6t1oTIfRNxCIZeyvnjnzadpKqXctqv0scpWGVotJ5yhM7IxgcK2K2
fqedGtCKQ/2uf675NI+p3gTG+V6wS9guOFK9hvwSHq4hj2bMEzIWRLGs9fWfuz2jDBLDPowmfKhC
QKurbW4z9se9MksLnIEv1ainuopEYud1uOWiVs7yODGoKoIROMgeUsFeBFrQblDQPtI8kAghDTgq
esQeFqNokM20sJ229PaPGSgzKOc+CB+xN4PgaZMqe5k4tIs71cKglciYhPUfZS+o90AkKc1POXAI
MaQSJ7szpZAYf33SopOGuAuH9MO04Ja7cy2Ryl0Ug0FF18q7/4G8Qa66HSZ1kXcCDhW7gneCn957
Vhfa938jjjhZ9Jy1JiBX+P5IkZy/hLHRWBR4Pfk0vUv4TW8SZDtkuzo8eNu/hyc2q75ZGO4LfuNU
XBSuTBEYbgGKLdXb1asaaynDVIMrok4oFjZff0JIOvilmrWBIg45v/SW3+W4JGC+9pXX47V7ZqS9
ugzfUnzZpBprdUoSlqjUkS+2NoifHjKfFEbVOpDn5Dt8oeP0KbscTsK6LWY0juwxs5Ben1K3XUt0
FpQwCNTsPwu7bce8vdlrNI3LP/Ksxar72uhIkz/cStCP2br7dy8+UV6LUo6XSeA4G1xCmUj53CNW
Pu88YLHfmy4AuJOH6SvuiL3qS6SiHvgUnVBLxFUTh6pLNX4JZfJMNtM55VXZDXLn/1vrXYvEi8c9
za0Cl05uv8lR96Av6kgeC7OxXrlH+RpAfZLcLdzUv+W/ACcPKQJhHOSpkLD6eWH+7K5qB+cyDlqd
ZGVQKlDo5MY81T/9zAS+RrBZn46/Lr+lmHDJ90/9GCDBM4DtPok82VAh100dwGNQmTROOYztDcn2
qQCHPSEXSze53Q9a8a3uBTiRvw9byO3Bco8VWiSe31sLiqHIodpyUoMuR2WuvV8rcPiVyNWKDPaq
JIQH3CwH9NNzqe2QgUUz+8jR+mMompDiFwM55BVWVNyd6tWhodaEZGWrCmBdrWpGV7QIIk1IBpuj
Z1bpWcjM2o4KcEtQ6qnnqH1fqglK5EQ2963/hBjVF83Uh5XPVMvY5asH3K5erB1FuXR8WimTHTfe
PUBaFS8RZeaLVfUCQqKhoxtz+0lLtHk4ffrcjdkh5f6/QA0dyUKzlSof1jDP43HAGjhsYMzKLuLI
EYkTA2gHZdpnLQMRKHPoLBvSbg6H3E18VmmoMIAxh+pDeqeeu5tP6D1ffVpHtREXVd6fyv6sfEhI
xt8brgJrLG2aORFZwHmdSrsHYeG4kbPmudSkrXmT23tTrN8CiPw4/JAWtyDiZWuCtyIH6lluBaMd
krThvxpQwl6KSx9F36+QgXOfZgw8bLKMo7AbPS8tU7mmNi9+ohsDS4Fyi3Uy2/ofB9ZGBySMzPqw
xtmw71QNqrOETwJ2sFDpbdi0w8IB+E+PB2KUMJt8vPxma1QQHUdLqraFz0Ztthxyud8zzVnAzt3M
7fe7lGnQWXim0hicEALoI3uueAk6CKvLB9T38Rc0qNr1xQYQvuPz5GwQgdFinY/4d03kq0SfKjba
UriOalP5/if/j721abCC1p5LGuA6bUyWfuj0Fi/gq8aKRJVPaGo2r5SMrTH1Ga+k5EZBuAJ+hGFX
4hYnoTyVfVp2TGgumJvvIQiE3+0jh0iSqN6TKVeMEKmkh3V963GoMDfdQDtZl5Pu7fZJG0TztS7N
smfdfkiW6GKP4PiecKBnqtClAvge1F8Wisw1yT3D98XzF3pOcjgDVN4h2GHE7VHMeyt6Dm56yaGs
RSdWd1cp6/5AVlsBzVspZnaRtgoQL88npnxtI9llzcjjCwkm787qPMblr+V2EiYtrpceJmWZiSrP
VAa3NvP3SG8xbKGD81/cXeVhKN+YRsXx5zvDnkCwPglkVcZzbBSnfGduCMWrizxJdQRRK0oAHND1
AeQQ3ejc+DbiZBRsL1yTllmpbzv+/w1B8trWmwAvtgb1ApBvMBqg41iOPtcv3HS17md2nB28B2TS
rffcx4a5oTQf/YkexB0wGPGsh0lH25mqkNJ9E76jmjpXJrqISeOF/AQljligjKcN4tJ+NQd7HFfs
P1eVLwy83LUlMxk7bNe8sRpi1zp9VeG8GfNnwVCKGfmczFeYYLKafH6ts7FXWqe1LpJlzKIsxEIK
e5Nn4rPEj03LBcDfM0Q0yQBbRyxKryn5eQWf/YWR7xfyJlpFqE3eOtdBLB1KsoW4KA/pDiZ+1Jk+
woyz8T7dhSgNtvWoYVKpqpFpmSa4SeEo8FsH5J7EmkvI7sy9uz/VyDTOgHyME8Esh+kVaNE6rVK9
2W0Mspbli8NXXGAyuBZtcPAkoV/EbvE0um83mQSdzZHM6lpS7iQpP72uQfdPiuSpToW59+0rOOsg
WZFCFyrL9VGfVL05r9iMoLy5kI6c0n5ix1tnvuITE+JbGFFmF1R2InZlT2a1fwE+MLkgNf4HnNi4
rfOjvlBhMbCEd3dWQYgkXmmrbKHvuZl94PhEBuYiARw9Nw10/qga/15zbwiBRMeRG8xP0cG4NPTl
QkWYI4Ngk3R+fz4xlG7RN/lwRon5Y6S1ardmccsJfN/TulQ7lX9ZGWLvhHLTQ24NnM0RJQplkk90
j6hGqcl1QxmDp07VzOT423GvD98a4TMOaYMee9ptyflMGaLCxuvJyxXj6jhFr6NzEmNQ3RJQgLxn
XWbE8Kdq27xUcy2EL8I/uRof2C8CAOfqvtLPtOSKxvI2cWDnEIOSUpPf2v9NfkDouvaxpuRCxTWE
XzWOAAIRY3R4MEOdAMIZHRlL2GK/YjtTTgBjSFtK1A3sKLF1YYtvA9wh+IZIxYlsYDTvOpD8jc0C
8aKtC5Y49PHczRLWsaQUsYgLQPFfbSW151kH9msmjS2JzSHz1mIrsyjaT0h89/NsB3GzS5W1qgHm
v3iABt2281loeyNp6DNfS4KpVfVmYUxLV8pnusXFFHRig3R54L6DVDN8SXUdaJp0rdLGZ7xLRhY+
k0tcZj77pQpKbMyKOBoZM560ERRMvipQVCM5dwbb8zNHFCZwNzlOqbgTIVglmF222tQpIb2+uRee
a4qrKQFMYg0vfFHfoAlWMD08wuk6Ty3ynP4y0O/C1QBcKuRoC3JydFkmI7Y4A4lgvBzlgILHjF4p
dxEXpofBkeEoPkb+cYhfc5ttrxE155t1SbZ+f/HT/w/bCQynyUqLn+N/SsZQnI54o4HBDHudGlhG
iZ2uGfteNf4DVHXeoOIvEFlZNOmvCV+CEkrGreKjWfsMH99dS5bLhjHp9dWUHaMiGPW/xBqLcIJl
eR3GdPRCfkuALpuUkq/dFZzgWBEP/1bo6IMz+Ww65sgBJ6HMfI2UimIAupmwdFoM7XOOHqLVTKPe
1Y1bPxlgIZRI2ebCec89ZtQki5cw5eiiCBDuRALlBu5vfud8QOUky+EmI3ZUkNTFc6AcA2xBKhGa
oOyz1wSLyASDcWN5uLR0FERo3FS1GnMCmlByo6rFmAxhwLrVxTwy/nvb/XJHW/7E6icNv6vX98+K
QYWqlErtOjiAmNmmjqiy9qfA83RDhByPli6WMuVnvqB7g1PrHnHUYUov0vJ8yGJusonRcLhCHuC/
RzoFALtTOaCzcy+BqIi1sDguFWTK3xk1cfR9pj0UL0gEHXCTwI+4NjYqJ67hoFyWmaUaO4rkQvgc
EimcXkOatKHnS00vsEvWw4krJyEn+o3zEAT89SpD7OyCvxBGhNYt5yrFzu8HUJZRyanmkrXD9ZbE
1YR11KXWlRRIGpcwxDV4OyjQzWKV8xG3qu6pu4nyH0UG/jXe8yLZvnKBOFs8pMZvye/nShw0gUs7
eadAAnL/K56Hdgomjku8W5mSKjBiJ+2BTVkiiwO0j66lD8TOSO5SYJ3JlB04lx09JsBKZa448DeC
04+z7mM9s8AnQ11JAJ776mDz2O6zMoXMbSTrEg2TA4xfMdb/icdrdRFeoDT/ipBa09QxepG+3IZA
BIvkmg9PQGqXrpr0YkBmkyTScm/WFczAFY7n9oUplmepExmqtbfn6CJVKCgkwKUD5j1cKEsV75nw
FdmfCbEiGhEHxnu4K8VQM4ZXD9A1Ln8/C67iMDMk2Ane8BShYT40h6Aul6cbzxu0uHnUfyfDLYBZ
7/izJklMF1y8+uvUj2hOqRrwcOqRBqrcKCQYmMITChqS+LRr7qBMqDiK0Q51yK8C5X0WKOKSCeB7
tcmJQBJzFR1ROkKnitGnbUDFK9BdLYzq7sULYg7Kkc87q3qcw3sKgx4DUcaEPUWG4y0pKeBqjuEp
/uxSq4g7HoBUj9fsX9lXx7D5y20Pn0mYgBDffA5op2GofjLYpDZctoXxeUizufmna1VCxpAdAeDg
8bSxrSnpVDbKGZ+kN2jhrzuVl3anvjVGWx1KY21IL2KlqIt4gxc3gbrXboukii4R9Qm+vI8J1hiP
LPa/zB/AuiBxsyudBfhyqtZh3up/afmMh67VwvPW9LL9T7zNq9psJAFaa7+oZYJzgpvhA5JX0NGb
BDZNT7cGFDuwvyCqQY+KKDlpKybiAtG//bjKlD0dhDXjmCocOV/0+4I7h3e61cn7T+l5eXWiarLM
yyhBFYMDFf0BSPVrnJhR1FIsw6m4usCF7kR2TkVV27LE7bMCSLX6bmpMj5efRUsWmihHMgx6+3HA
+4j56SblOWFzXn3jIIuF0Vf5KTMUMUp9sYQq9Wb1j1aRADj3edHWAm9vULstqPeHLP8+CqT8udix
xsV+N+9JxZ0n3lrz5a6R/9q/gbeawsM/wsbNkQ06HWCpcku+n/9Xp5K6JMihNVBTbTgTPsHGXEes
eds/KovNMSl2SXLaEM59x5LRsnwgFttF7B4nFtSskyYfPHq26L5IQWgAI2r52CgX2I9Cv/oResb6
75SJ5kqbfjWE7ZVgyA+KHyRuULgXzSCqFqLA1KbcSOKr0wfCnA73cGXUvn1FxUYaESiwm9iFx3yT
88xN/gb88KxtCFtC01vhdUXjSkJM4sa/lyDx2hwEUyBTPksb1m44/hmc9y2hXvlQAFOxkiAirLin
D2rhtMTq8wO1QF5x3yBLhpC1I2SIkqEpx5DJa7k7OyL2M38K1Lakjv9KtS2wX23NYqLAHiMvKMuw
2AX+WEvIENr9id5pn7Gr6cX2joQVMQMPYxMXjA1G7B1AI0YmoD9NSbRJA0uM+LEmx2ge4cparsI1
ctEvM9+IKDskz7ZHILk67tHegMxT8Qgp43XoVELnuCCUPirtBuFuD9xGszH1WTv5NxTbmtVem8vC
7GAtf8NGiXs+syf/4OGGPV+RaQ2psp8dh4qmQIl4ilrw1wohxbjdqWtRTSNLwcoPwk4aRoQNFULM
ni/4drf8bcXdSfuskkXGfVEGvSBLqLPOuH/Tid73VPCepq/t239I/fWaSDEqg4OMJigxr2i7n5NY
iHy/6ry+QzHzzN5fzrMO+3lWhfuOXQxzPNehBriuURn0w0DUD/YLJfVBnlX1wU/lI9RWG2HtwccZ
BQj8CxLGZfpKvWGv9+X5WUp0Ify9WMlvX34evWh2VjLvXJn+hwuW8Jd4xhLFYTelr9yeJMYTIlsu
YSyqfWiWWakUsnGL32G3DZSZgVatE7PEGv8TYHTug2zOHlvrzQLBKHpCZ+9g1gDQhkzpYtdrhmob
pQ+WToBEQcJlJf9Imbta7xszP3nTuG5t/pgZF9qj9K1u2Y+eITD0Vl3xyvLXKTcJaste0e3ASWEA
nV4zbc29Zj/I9klMEizbiiRR40sEtZ0PL3OLaIMJwBXvTFwNlK2eK0gNNfcNIJEKAHwEmVITia4C
ub1Lh1L6b8Q6v2HsUeK1CYE449PxPz0ewcCPgtgIUBTVy7tf1e0tsj361xgHrZrwDhHBq9vqJbvU
BIKQxubBDfOBcbjyOXsMSgLZMhuPlNoqshOCRcYlM3KAbNqAc8X19yzs/yEeNFbmNQAs5vapal6k
+xECmiJtWgq4amzf7Q21lbmTjJWl8Ro4UEwXKCO0FwRwjoQui6r45Bt4ffFQL+ULm5xaPtw0eVN5
CqhXNBQHVEdDLkL9o4Pod/hJKKr1GsXklc1N48L7pcEuqk6leeaFP72IbOmqS4g1QUSfweGYI4Ea
Dt/kobUnYIxA2iefFv4kLQOSJPRJuV09sdeIa3TmNRJQwAyCZ4K/Pi0h/czb6gCIuR5Y2V93QE0u
oKOchpl1fQ/tyaYXDK7GXLM8MbDHgVXnBzNxGdZ+sgjk4MIdW4hyfGwelH7KiEIsGPN4biOwyzI7
3QWblNlP0FQUGovtyd5KPd9hGPD0D5oYsmuglyrNOGMuuzWduIGZNVZHFX3vH2fuQk8Br5BEnAWY
BIrcl/FXLxl4qnuvUAQoT7w6WBJAQzEj+5ZE3dMdQHSSHOPJ+Yhb87uYgykr6FlYO15hz392SPK4
roAufrgVMinpYLMY39ozfwaoH0urWve16u4z/5Hicjau257Kofda4wqOJViyATuUa49voYWbAYgl
3f4UhxpQQN4tdWh8nMjdrqycZXaespB8Wsq8aaQFYb/DwUBTDUI+77dCcJ7MnXu60zY6Xyd1Odom
caI1p0WffCgo1fVnX03Bn+iXKWlTwzNIykFwp6HXtY20nOaB6EcshEtpbj5C+RRtHPIiX1fGlfBn
B/xHLAeBwF3SMA0tRxyuXd5XS9S2D6L/FoUK6DgzOJCUmLucOyTl+lbrlormaR7AM3eHjihFUoTU
5fAoCA7k8nHYMuacMMF9YSwyc9gBZ1fpJ9KgOo/LU8+uSYY2AhmvmmIQBp4FyWrzgmvOH3I+eY0l
DGzHJt6z+Ayh+sPujiomS0v8FoEYba2uXm/b7oTeRoODTh3jY/CcDBF4Ov5YVkhnd4yw7IGR4esy
7D9aMfWf1/pyIhpCBp0wMeIW/yuihgpNXksOjExLiHeP7tj9g7IKqAlWPKmXUVheikLMBp0PxWF/
19n4TZ2SnJUTky38K5hPc0V7kIVepHDrrGmLllzxS9vAq/gDO9B/Dryjwa8vlghTGDTy1zcp+r5z
iB6HvYnp2KrYhWWPUrnFSrUjT8hufWF75hJVh1e5z348xwh0s98X8nVuz1NsyQJ/VD5CcMUzeFRV
CRANXT4VzUqx61qZBpO8ClK+YK2ApdKQkKivev7FKwDifSHTyW7TctOlfqSxKDobAudBkmtQWqgQ
pJfCfK349KuyjSbb6XWOd5sxO3DBu8N09YlOFxiQCnYHpoeGdbu81FCn9ob4iRQ680Dff8jVod47
hxgsCJVSgum7/rjXQOlt1jeLOZiT6hsRklv/hVWm9e2gcepjS0Qz48x9SrXtM04iPX7CmYyBQy7x
9sIlHPSKHIxKtZyxn1jbaVMPp86VdPp6t857ocHxXonUa6JUQ/3+9VL9B6EOWwEuhzgNRUwXKgVH
cTyVp4Ueb20XKQqsk0w/WcqQ6MHFqsMlV2qb7O57ZJucZ5PwD91Rd3OL+tuKPMp0ZHXKWtyYN9+u
91kMhN45Y3+4TdMpNfijFRdUA3Ut9vPQWtAmRw7GVWqgsAFX76MkVPpW8UxCioYot3ffYFnH+3T4
EnldTMIRdADzhMzfHKC2DsK8urB/HEU8tfb2Tag3EhruZt7xAKM9qgGpvhXvrXe49CYLiLkVM/2l
Kr9aD6VLEajbGc5wosQ2n7kpvLxhhmb01yFNSCg1qoMi3NLpqYw9ru9jPgyh/T5pDvtOfBZXRS+U
Qzm+JuPiAquDj7y9E679sicD7mNqIW6i0Wu6dFo38c0muVQt4NvZaApqQfIFTLRz1yGK7HpR/XTD
pqbr7JbiB/FGv1KFRmUtNHi6F+PMmbwzKKUx7LDz11gC/8vO6uEC/CsoCB0FFwUjezL/x8JMabKQ
qb/OMIdCyWXPbNHTRq3JDhxR7PhvQLsHgzjqM80pkC8gTCJkkBMhBO+MhAmii46gQBHppKCBwySa
PpDChTwurBYitIIaUgH8oH7audRlQtAKorBwFHVKUyvwthwryH93QFRTjOSN0WUWlELLR5edwzcM
sR2cNQgj+TH9AqgALrhS5Y9S9IYmZNx6w9YW8GLCSxpRNFxOZ6Dxhjf61HPZcBsKmb4m2bLyw7yF
waBEu67BE1Sbyp6p+HiIruamlb6AmKQVs95tXWmbdA+e6/QeMXdwkfGYLf/MH2jQhjsVqWbYvlRD
oLZPZTLS3Y2vgMwRpBc4xl+L5Bg1UoU4kQIKXHNkaOXaBvE/4MkBuNaKt+oKyk3wyLc7y9UUM3DI
wLDECdmhltdo/wm5tI1dAPr15MdM45MPBTjquEy0ZAwfj/5zP9ElGs9c/xYlZ4nr8LpClovnBQbx
z06koQB5nEEeBpandFpxOoIPrdmaKP8cRwWdIsTd9kqETbvolwkIyvDg3acL7F86qSMrABu1QUet
RuZJxdv+p/ZnZQ4qQl4qOwb+iIhlChQNPk5Ctyh2Lved9zb5nX2oMFXl3wP8MD/Edj6DNAK9oAe5
AkytvM4rTtNBHPc2FQJCYBk1MAJFmIGKQbmEiAQ5DF3iHtvGsZZNLwj8Z3xaIL8u+XXo91KGL5pU
cegSY+o801UX1MqVSJy4+OjRGMB8Bcj/BW9HmEi83FD3hQDvsqjjPBDyF4pJiKn6Jc/JOJLHarTf
oUqrhQbSqwxJo6+2KLwnfxfbHQWq5fcQ6UrYWN0ZYLmC3HiAUQO48ZglJd3cBvGC/ku+R+/R6srW
UDUgd0rKC0o+Qe3vKrChMNkaOg0NagyP7wSEoqV+WJVunaXlvXkc76Dyi2h+nE/bp8cAfq3EF/i9
x3Z7ZGaSlVQkUkZI3J8pBlrWSJmldr3ZAZjOtD9NcrhCDDICF+CvXbIZ0kMwAXt19mhJFA9Wu/i7
swunKrrFk350auB/Hyrx3hq2ztsljvIPp01DLN8D3bIXAZycaqPYBMy6pYt5P4n1aXvX/kAk/2wK
ugFALX0frGpgfm4a+J+HXOdutVKVy41ImoUDGU8egXGhJXMcMIlYtxdOu/yeXkuR++UCWqr2a3y0
62se5oa9tpvpUMmpfBPwG539+uK/FhpBjRF1raKNp1eTWDHl/bOpq4EAWMGJMuJVlA5LT+N26r9l
6vQRCNEhBZTIif0r2LusIPuSDoPeYm8+JH9IYmk76vTRr7LWhMH1oHmaS3Ixa8gSEsXB3xp4gPK6
UraKXmqoEnO8NzaHjAPV2g5aceAnnqFe2U2NlyleHz35m2VQxAbiKf4Ra205/xml3CDJWkzuVIo3
dhxEjRuOvZmOZNv2TKIjLamwH7uPFpodP3uzB2Sp0KPnBCB8oVCaLm5/zHTBk/AoobxBa/SsNkZv
wniIRMl+BStXhcCPvdb4SHpt7G3MvPVe6G+weLEEg1M5jAoI/F2l/sA4s8Xp3X8PyL8Gqcs0iNdU
tCe/KIJhoM2woQljBw6TAVpL3dahtmeG7FcnONXpRpLgWaJkwqN0FH8AVw7yraEYmEwrn0TFaCzu
0zTEeytYrhU1gpe02Z5qkWai7YwFzquBeQDg1CYs04WnrBw1nI58eXuzdO7xg6BdFfdAST3W4V2G
1BReopQZxYhkPx3tKs6PBapWiNTx5yVbqYSQFeAhbdDOZqS+ZLY6jZ/jvDrcXi9dAtss83xQVQ6t
Jm/t0LnnXJYCiUazK+HUe5w6MkL92fzf/jeFCdO2L00Ow2p0YTH0ctSMdIn0biayKVEraF3sp0+w
wKQ+tK2OXV9ylH5zJmdPL7VE6JIQM/51jXi4aWnODoIpWUVJiUF3ca7gTgi1Ig8qRHC5zHO63nb/
Cps8odyXYZaS6TRHW2R1hCDACa/Z7OaVipU2XCdfsqQYxWvHXrgiD7qH3P2VAEmUt7QghzJw0NFY
dfF4IZx/r3TrT0TAK/9PwzEEjVYWKnNWKwu677r0cTj1rdESSucJkDytlmtIfyUIds2ifllZshg3
XQlWo8VEBvphN87LWhIfYUAHUzFR8CmKuiO9+BMVAXAEZat+hGzZYppt5dm7jXe7Mk0KQYU748mE
do+bChrah/F1yEzBLWr5fA7MlWHow6CkwAWeqCvnjT0AVBFBi9gqpdwiKnuIrvj3XM+DCkGGcIuV
4+R+SaM7p+pcvHG637ngGzzVbqjdd5C/ms11Xhdm0zhTaYfjC4+W4MrgW7Lo5jP1yfEGtV5Mo89w
Wl1iRgaVM6Syl1CS9gIQUvu6wFfIUqs5O3PrTb7LHUHp5FSpcSJATtKljVhhyZRKC+Ocu4tKqnVN
1T2yquKwWq31TFH7NGQV98QxMnMrhHlpwtc0MGorT/v+v+lGnOwdCOjQt92Fr2YblJ5vMSPLVu/T
tcbh6KtnQsMpd4uOfXY7Y0FkNZKqyHO6Ym8afA+/sayMUWEcYC0BlwKGg3c/wpuJbAMmeVct51KJ
wlB9ynB3OKb+5g5x2g9eRc1fouH0iRoqZo9Ll81T/ErhDx4CLkzwShfxppGrxTi2z7VNkhv9xJwD
3VDtg1YH+O6YmqQCK8fJbyGQzKNockE0z3Uq4gOpkgjtIJPGUHSulZkZomOsjNX/z4tbYShJgQ0d
zW9JuNjHTIbu3DPu89iG3ty+FcNcMYcaaS0k5AyPldS+IQgWV3K/a/9OXq1eDxtxPrvOS9qcEepH
AqmzN5xpRTLk4eM7A0Ooa/xf6yr1MGADXdIpO61iljZh2L2uWMeqGmcXPviHu2+olkiUOzHjkvQW
DWoYeOOyLOA/JBLh2PU8lIk+e1BzmxUYR3UFfWw4xGCu2EupnoUMdJwPzJgzXv+ayY4olnLSTNX+
3NYEgojFPqqvt84pcKLyYFoTDuto7GGr+dfaOTyHQPL8IHRKx5lOZxCkw2/RkcSyRbxZCaxDa096
CxRJzofcBdHw9EuC6eTEeD41g3oJDFRiIi56Z0ceZwF7wmhtI37Npo8qLfsYVB9HGH6KIcFYGJP2
qWgQ/NvCOGr0ixBq5sGwWZXwW6F3c6NkX+OImSWlVp0JEaALZyFqw63x2cbFyn0OdLxb4t2fcRxc
5nQQoJRuVnX9qzOdoBJGllpPo7uuOGaBnDU21o9BQWL1VO6j6uC6pDyFwdDgQ8tEkGZNEAptr1xq
f8WDM5eAjrlwCVoVgr9k8moNxdB+M86oGOs1mYW50dc5/PovqJEWaHTwF1HE3dEImCJDlvU3p4/o
RSwCGZDxoaNNm65We7yON8AoGKXFomArjaP2cpt8UZT9LcaPtb2rwqBcQV1DQV9YYxTD1HMXrwBj
0Fz+X7x8hrM6K23HJEsSPfgUX5c5IxeSdUoBk5srZbBOJLfS2ReTI5OHDD/3mEPUQxzXA10c1YiU
h0JID3iPv+0VoTH38mOUkkpo91nwI7ae4/wOJDMY57BmtxXwksTpQzCCCobpFF2RpK7GH4ROg7Ev
t3CAbKZOqsJO4+hAaDRQL24VmnAf7LbKEwvS7ETHh0CSlAPM4jkwBJ+5oDyJwnUmBQw/VNHVc5X/
FhOBL4mRpJS3jeBGSAPRTurlBmM0J0OojI9cKu9nqG0DHcZp2CQSSACjWWPQDrq3r1qyHf6F20Nx
pGJsA5AU0hh6NqLXq1V6b6XDNYDhINqrvjGvj4NT4tjPJ/09mX+/zDRZ0u18bxU+IdwEwmVWPr6P
k7XAVC71o67EoskbV+2T58lSxMpbIYaeVH3kKY2TTjS5++KO7FxXFp+JCHBwDhoVqrR+pAqweun3
uutuO7XBmulvH/uU8kaIQcjm9desXNG0BU9KlsrpvH5G+h5Hqa+97JAaCdWQYIP5n0m9J00zmhEv
cicfSjdghXJqsaXogjlNRntDjvoPq65ZD8RsZNyxqlAzusSX4MxIrN05u9qJCxgzKnXpPLr0ISBF
Rt0GsnbpXFRRmWW4Yip1GeIyFiV4ixND0CTPDmmaVKHc6muwdiej2mYyTIzgm2NBvwAgDZN5vT5K
shoHSRXhOJ/yW1j/S0H3olxM2F1mJqdYomH1lcU0ygGd1nOqDThQd4y1WYil/rVcHyxFmUa334nc
/7qrK6o32DCUeVGGiKepZeWtL+54nklfU4Unu/IBYqt/CqEVDXG/HSzUTJo7FesxiOJrNEq2MdZQ
MIDpe0h+b49AtIYgAZdYAbJS3M6x9h+NffF/pmnsdP6VM1zlcC0xRC9y+VpTxjTLqnD7POpGqeRs
DiIIVZxGEr7wZhGepKc5tYNBXJRhSHN4qxM/4KnAL0MdG5Ui7FGizl5FFegKZpo+rtP7ciwuXKuW
igHqnbUviSgSFJy83ACKm0juRX/uGvpYC9Ck4WIjnZ06uCwYZtI/hXf+zeAmIBn9Z8c/XIvyiW6C
+fnhlkTnKUJiRH4VhAj0/yrHfF3FVmSBPwuA214kgCuw3oTY4VTYh6FIDbUFr582dav0WGZNNUdE
BWU94WB6sldXUmLDLn3YbVb3JviTyhIaR5Q6Bjr3elPGU2O/P6mRDJIxjs611Raufv36jGATSrLE
VbMHKrJ5Feix8LxP7B0FNHgzCaO0t+UWZlr11krBNk6y9eBC2e4nMSrYd+I8SIo6gXexSW3C5opT
QsC0lxhnzgnuMkDVpjOlH8KI7zV0+90F5c7mQ8Gh1wG410uOSNwFMVcduj1or8Rqz7JdOzscXWpP
CCVma+L//okMqWC3iFoyIKLGrRcwdiFgw+eashklAqJ/wWn1At/HlgYDm0oeonxLTkVClxf9f8Lt
pVBL6ar+vIgYb+kD2ArERL5VdWFk0ESzzskSdJp2HEj3VmZh7EyQkgRgFS9P77dUQXIE8MwhH9y+
erGY2m6B+oblUpvuNIPXjKUcocekhT1zdxSaSx4owBksE5vSES8GzBsN6+XEtaL00SLfLukd2DcA
9cPpsQPxxt34N+cFeR6F/CsRfv7S9cUnHWpH+aFE5EpQfBAhlZdA8g/DqtpMQ6SnDGZIRuJqXZEh
pH92RHHQLMAW7oqeP0B7/uCkU/aKJcA/b0qfXJQSZ9OQ0nKYlj73W5BkShdojuehIYCjY2JbfAri
ek4g8ctciQ585XCK6q0UvEpQqALjsmREvW10pHArmMiD8wK/18AmnrNpopKuiWfuGMz8pItNVJu8
Dk7VWOKY5lcSa3OtVxjgQsR6NB4glIXhO72/L8LUQxJIncaOOnBl9BbzHI1h2HT0bLiFzYvsDX/X
HbE83oHFkG5PnEG5UpAzTfZX1IPPdpSQFQsNx7/HNxayNz93Z6gvJAjwhtyvFvd5dP5LxV3XCZni
vpDTUiUJX6Sv0VYcIa22R+VYn+UMJGEFULln67hUd7LKjgHNLMR0f8D2vghCJy8B23jKRffAcnY3
FPpaIGUzyfrvsNNCMCX4cF3EfD0pIEQHim+xi/fiB4omawZM6KhDNpTg5csjuMEtVfUP2HnpA7Wm
KmDRerhCH7WvyiphJeFtknh1IDRYrcqks7SYT4yC3SfFKvKHq9G94Vu/UDtRqv8rtMKIlcPSGDJs
mJIYKNoeaJrK3J/00rYrdRoZLJn2v6SSlI9yf7eflNPOrYfqjKJynfsrfMzXKiDjWYUluaKl/mT/
WdQjyFWCh/+PLU49h4Q9d86bULS+l/VpqBe8K0aasWv2ozP0eEnCRPr25K7PaZaVAyIBjOODQt+8
NCyP43uKAjQE2WrU7rzWhVcPrC2lrbF2PFaLL/Rs9y+JXlpFS5rMTv8MM5S9uIqd4oIC52lfGq9X
xI8R5DutgXe7h584Oo8kAFqNL2VtxpjxpvcOQ1qKtRuofn6eN+Fx7zWJdFY+A5s3WIkwjpefSk5/
DBIqLZgm4yivOu569QkLiBeWPAlm32KHcmWeP8hKSyAMgD32j2p0X/sLHugruondxnirJJJB8JpN
DCr95RzIqSd/yM1HJvM4Jkhpwq9pDIm3y7fkpZ4Cu9qjFqnHIhTiQHJ39moU6ItWkj4kjCoWlyE+
VO2IKnzBUV6RrX/VrMuPlJSSdPekJJPI+DiLzQq09zYlhAbCii0v8WP+J/gtKDNIGsTy9vwJ/9Cd
KxsrTzV3GucPywppeCHyFapkhkqLfNOJPsDlY3xpXTeFRSKy3haZVw0PQN33LwKbyvgtoNLt70Ye
gF9y+ZGcOVJpDOLslfWk78LjbuI6t4NHCbtZ/jdE3/l/GVWY2z+MHerlj70R/e9orY49DorNPuej
CKYrNN4JDOETuyCJ2fL+QFtmaH15ENQHJXHpLDP2rY5QgcCzgblUK6Nnle6sVwpRoxYlWaFtDKeN
/gm0RRC6+o7SVUtbR+dAS0mT4nYgZm8VEavuc00VcSqYnM4Rfv848meaHftxXrzRjqZR0n5V9ucx
JulXUDsr6l4az0PvB/9R0T90LmDMT5fWQfvVO37yLIev6yN7VQdS4x7TmN5v/DmST8tQFfoLrzQY
L209BCzNEPEfOpv+Fu4BoCgxVZLDdBumTGwFDP9Cp8mdYLAUFnDgRMcihdlfpaYpKcBRLOQiFgXy
IjaFNYJeKclZ5mRsS02WvdLw6ovutBbdMWNWfnfcegkkLbIzhsYBnrkkrUK75Mhelb76rnXW2rW0
OkorFf0KS8eNCWuG8cDGUIFVI56jCSukKb/R6I7XAmBUMDC5Fn3N9ROmVcNWIUcbWEsoP8l4wRU2
VO43KXWlBXVK1a2rfb1973E8rg7hVyogRze+6TLIgkum53j5EruvmlYOt81jlOS8q0ymfsIJaNDu
oo3mHKjTDbNUG5qzoExONrGIiwddA1BlMH5n2v0oapPunkQEALyz/TxZU2iXcZroHiYzFiHQJAvj
1Zd6aL4AAQx2+KZwKIYIv7Ne2glxlyG95fFLMjbc4mBW13SSewQCdSuyR6wfuaYYN6VuJYHHJeAO
BHgrsNDhok3xzx0j6dZVQz5s+54f1mBpVMey3NdWmqmgSgaYNyR33Cnmr/owBNeS5yTG55p5XzSU
IJHx+/F5SCJCeFPF/P8Uo+kdUyjpNI2wDOQ1fI7zd4pdkc5lqKhFtLiPDAYUDivwFLPCGI/IvH7E
YmXwzZ2vJ/XYP+bWZiWeLA7rdSrupZ8yRopX+lWtddzxgMDrtjsI9OeE5Atr6lPYflGNuFnv2NvE
H+EoBVfHVP5O5rgPvKK6TrxUKniPdiTLonOpx17cuE4oL8oG19vUKWTCg7sy2/1z5jbRnN6KGv99
P/CnY1ok75oIZmvkGqseIQHprr9MrcMGJfUpPcA+6mQXA03m0cWa83SxE6VIEBmKReHT3FUqGjg1
pnPfpe0CfaVejj2zmLyZvRDGFV6mfphZY7gDLrKMKNhqP6m4RCmjAyggqJfNQTfMVE43V7CJoN0O
fVn8q7WUoajxyDUOH09cGxW+Sjw+vX4hOnMVrVGKcB+ocGwPWrAyjxPO74lsFK0ZU3QdRIO6YiTF
vllFki969Bd8G/xfqjFZjB/WpZYHvd+SVg6klTXS82zv6HVqr0QCc3fG43EvWKIN/2DemXjGhbNw
YtPo3v2X6ukXLCisg/UwnTEsHryihz8GA20QRXkGfWJwcLQSFu1i0C99stL32EJ9q1kLrX8OcgmH
OiyGqc04oDqdcZArl8JBPltvhfifthPqKfSNdqwzxBzooTRH8StZz28QSKRmk8q4DU2gbI0tWwTq
YqgNo8ZCrEBqIG7yKJcVEFAZaspuIIJVuYCbM6jrfOyiZqHdcv47PyDdseGBgT2uncSqlQMKA2Dd
M2h0NNrpwu0IIBLRXfcRZQcw2oYXJB8w7yF+8PKDeRTT6keOHaYHAw5ONC5yd1JvD8rv0LBzsm4a
9yik21JfFC71gt/wKxsdMGpMby+zpyPX6wxrlPZDy6Bjg0dvTXm+rMCD8NOnmQAOtn5zRzJdQz07
/y5xDLIqPSma4Ge05lGOfC/PZMBABYDdyII7gvgvuAQ3q3jR6q4/9bpDbRwEfqYUGrPsB2GTczKG
2+W3xi1VdLA1TUlbf4OYeVlbg+SS3lUbA43PsoXAaqWZa/xsKKH78FUz5I4ernAleN9eiJoV94kD
5TS8Rnz4FxmAUn66XrALwXlxx4I85+A5lQAbV5NNRO4v+d8GYFSsAEwr7N9rJKocUw6ECCwU3UCF
2ifwN0SpxfbswGKFW9uFzjcur6ab05yCzl6Dbe/7kN4nyCpH+wGsbmaU0CAh1xnLsGBPkhV/RoGG
eh9CxEIBVPTxQMiDuqQhnM5iIcLCi/Dz3iHs7pOPLWqcGj1/VoQeOZHYN1FHxZC4CVQxPAh+Rkmx
ZpdnOQUG85y0B91GZ9q3agZ2nuQbEE2GxmbHoANXqLaApq8Wj/G0Re1EfHh2zqnjHYLGM4WHdtd4
IYPFGqaAowxA5uFu8PnZSqWLLeBiYsEh8CivxVa7C7RxXUcoyp+0Dfdz7FsJOH8tlOTW//DDBEhc
p/y1Oyud0JF0NT1vsK2xYzHt70CTfnNd0o6+Bsc5NAq8pJ7Gv69uZ9NIJE9AnBdKWzpIZmzLe058
l3r9jT6VwYgVpqwElmQpNJR8S+up9AB45wzT//QlGyyKnb4qIRDup8JsMEwHfmBUm87WIObYr4T+
2Gf5k7tpjplqk4vnRmxz7ZSCg4Y5inyKDMpU+8yx3CAT/mPGYPmjUd0GVtbKPo+Be3FKsVitodDH
eYdNvYy4XWkq5crKbtbiRy7pKDFWo/aVCW/Bc+TWOqgh1TZ0fsXRVeDhvHcBY9+EpilzLJ2oOzR4
nd1Xe1IebjSbNfBvUs5NBx5sguCrjuxyI8pcXBsf+mynYplEWfEYljuXopG+xJOpqgvZlxBplohF
YHnZlMy7J430AgciFCnJ9mFkoXfEls2rEhB74NJiQ1mWBSQOaopiaEriGVKDbqMe4B7XrvRtZFJD
s7DDnabx6SxDWntrEu3xn3s+YhbAtpo8SbFGUZuQAveA/zYYWjBhdkDO/aoCMdStghlPygQFc1B2
+00f1qsxg0ExYlr0e6z3/qsItQAVN3QpOKxMG3G9r+sSXIB9Nl4KDxWhWnNHehxS74TCwttJM73w
ez67w9xGINHCahFQuWBJTtaWzm6CwaqrhEsPbxz+GcB3LaH9G/dkz2B0MKJaxHAJ05o7a4Cz2R1S
G5FnNMCuiDalEd+2Jv8DtdwltOJTq1LScLRi465IQdAN0NeL8+XNEHUkbbmckd0tOqOpWEdHTyfP
30FIduCGgLoVIt0JEFsMmZurAD/r0zcnRp4hdk/avruQVKSni1JBzicp8oRyZK/r+cP0dBDQ2dj0
w+esSfdknOIogwxqKxSGHo9qXTHouZOW7a2KooBtkaXiisRN++QUpahWPhlmXiTDJu32y7mabps7
ewziFCem/ocIXwA6hziNMZAMv+JAGUmVaJ4cVcmFgbn5kJt6oofXV9r+Isv+9lwk+b8f5EF0mRwh
96zJ8AoNJLuK6lcK60lTYAVzGY0FFLGiQC/N1Spk538p+THEkGcYzlwIRV/hSvts0Th18HY6FVWi
MkxFs1XyA8OjWVNQ14H/XnuOXJDQBF5pTvHHoVABBl3HmvjYk2XwwLAtNUU4qImUMlKxDSd5y6jx
8SPjdcKlmRMHlEGmmnAAS1BBFhoThAykRLeiaxJNW3gARPnW0aIx2nB9PJOrlw9Dr7n4j2FiGINY
J1Va+aFqmv8Alx4JK/xxTZpiusKM+BdK7qcUpGt/B7v4uPr6DImoR0Io4TUKQgatycWaLe1EdTcN
womyaoYSGDd5TGnU/y+mBmJPqB52dVlHr9NDwWUW8O5Bm7GBeMHbMBJDRqSnvkF8JUqrS0AMCUi8
CVSIHRTsQn+wgobvTbfO/5G+79L4NnhvD1OUQQVDQ61a5tyvPV//WvVrfH+Yky/1dA9lZjnAkTi1
NyCmrSq5LpPvAD809M82AY4fun3ceQTpsc5qEeRrX9PNt1OR4o/6RpZwXq1WlZ4IrRW/eWzNIVPu
WB1Ka5fZA3Cds7SzbZRhycfVV39WNG+iN/VIrTjlKxNq6N4/aGMYu+xxZjFpWDJDCQgiWRaMHu90
SIaEXk8crLbZULjFsKeLxG7lPPV0pj9itm+baAWMXN7kb2c5sCj8a9mqIY3hCbrjJk88JAntlzyr
8Zb3d8GX7uOycswe7iJsKUXl7yp/GebGWb3z1IJxXAKpfa1III+ffSVtAwyUK2ma3mkQVWMvJtPf
rD+xEmwPuVU0aw33WeZyZEhcQiNw89nGH5uy/jprBrA49sRqzRS6sQzgTwDyX0BGQ6HRi7ocxi0g
xsfUXQq+20mZ78U3+Dkm1/krS4wRg0WspE/0qDq50fwpEJJLk6y3A4UtceKvetNM6CNJ3/ZoizUS
sZ9c9PCoSuYQMJq1YjoFAi0BcZ5n4Lbx5J5UUissC2Pg8BMWp+gyJTuJ29fBHIqZ5tOZH++C3vw3
keiGeoeM2+JnsgVEPo23TaqkoKoXgvimlGvTYRYij7pN5B8dZ5MfLQwLqgkBArywdL+PTQIbfBLt
1CkDbjMsezANrHSDujSMTTt5A0LmQF19iojQPclGRqrZwccODt6DxFAeidnnpWgnOdVgJkdom6+n
Xo9wzsQphhW91yPaoR6SBeQ5SCqlBIyWj9dclHw5JsN/MYuHU/DPTv9npCgCMHsJK9aGgB98jldQ
znwvjt5q17DqjBE4NrD7bS0AcIhGWPHe9onzZFwT9CHgQq99JZU6w1BsjbAMUV06cCHQtUTFa/XI
ms06hhcW5fjQZRy/U8VbepSUNoMKhLSSHFQdqOfy5hOS27HxCtX4lJZF4YlwVjsVeEL7AewYJBvu
Fti8Wm4VO4zJvTLvWkih2KPMsK+xo4I6Ib2lH123DnB2iXpYKylQ7E/RdcCXB9EPd1HS/Y/Wj229
XRySTqQhZBpTuPujmRla0xfcM8nUphOITWh6haFBDZakx6ibBkii6a66Hp7Krlqh7FtiOKZR7EzE
Uj0TlbvWU0SvWGV8OlgN44YXRlh+Hir5aIOTHGRl+tzc1XOOL9LtcDKms2kjRoO/gzUanpiV04ot
dzUbAIDN3TSdDI9czgY0MYNZJKj2qncLRl+qL5jLkV+PHR12Hk+ILGgIYfpRD1TptVefYlbRrTi4
JGDK5otQu343rf1jhIlLUI5b2FlLw5t/Mu0dybkkgp2qsCbZARQhM6gIJTMjXpALTxYRC2OQnPgm
mHYdiEyPt88XNQc8w4SHgaa5Oa1AYmdE3zqSNHEaWLpRY6pHgFLmQibPjuwXfiUZO4LFvrQOEBrZ
RLMmEwho5gdtPB+UWMWdTZwN4Ssn5x+xxHdtY14ExBTQQV1hiagQmS4RriFaX4qJofLfsHdMsEQv
TsC75wcyB93TYNe70rwiZpUIzgj8kOXg9yrbETPKuRum0pJvqsQjIRTMOOu1xOlNpbE/IKfZ9SQX
7ONbMLWEcRxH8/77ZWWZjlP6xzYWrShkA2JgVyrgoxbyVpD/IQEDvRbVutehX+CZvMkqToVnRpg1
r6afoNIkrzvK+Imhkj9VqqMxFDgdDbbkVh6edKd8v5mm9+o1rdPUNusGJf2TC6BFsSF4QraI3sh7
qvPZRSeDbYHKawtuVgR8UzW/fDwKErxazkj/k2PA4vfDU8TPkUzC1SuN40AVzlirTlNn2kBYFMNO
zemARB+Ndx7GDRmbPkKFKcCJR0IVHP/VTCEqCYajSOW50bhyjc65W9fq8e5pvjmlm38zxOIFHTx6
+xgKk+PxAAGdWCFC1QBbBq0b8OyZmXjgzOTkkHu6QVDZZYaEzul65WAk8BSctTVJ6gsLGbJpqSV2
1fe206T/iGz1l1pkH/kiDAaYbfC8glUwxNakDqaAWWSnyNCoD0E2DrPZAdeW/WG8/NekNtiUUOL+
eJcACGXBROYHokNfwgGJ9IPn2gOeRdZ6CZqVRf/8RjBqUZfho1kfxgcoR46Iz1xyZRGc7L1imM84
vpa4li5LR5w2cz35IfvKEynOlAxkxjV3v2CHldLPBor+0Y7sz73a9av5i0B7V03tICznJgfWrWAm
TzKsCfY4wRc/qu7sru8AVwpxvoPaYVrC7tFbivYj4UtuHtXUApV6gn3yfCq0dYurdd0g9AYj5kIC
He/MmZnNq6N4Cgo4U4YbzfzeITuaJjMZ2Y0NH/lSsiSL7nQIe6ydta563d+dnDLGKrygLrY/8vxO
rg0svq2klvnmR0gOVao0z5qKSW9nUdi3fmR5w353rT5DM8WUxRce11da1zT6UWYmepHgtkobwiot
oj4DNdMafBBO+tglxYk/NhSmzVxWrrAyQnwo5Im+BYxlAYpRhCUCXWy54TEel3CMS7Lr7t1yYWlW
64+xm8tT+MhGtyzsZA4X0PzDuoStA8rtd7g8MSAWTxL7MSEvOgcyCCN0tR4MoSYulXdYR8RrsFAb
rjh4Wankt7Pm/bKk4Onz1p6LlPvYlaOQPTFW7Tq1HFpksL+XzXKLhSsNb0r/bj4DAFmcWRVOBsd8
V5RuepnXWPf7Drau3jF3w/zT89SYS/vHSelxunqsNS4IjDyDLLuPsk3eIgLYj0fxg+ISBM3siq7n
guSapaFjZD5hxBmlb9Tk4bVbF3N488cRbg/y565lkPITU7Btc55PzXJ+L/yAUJM6aK1VbbTUhBW1
xOv3uj6LYxCl1UUZeAknVeug9gUXHMkAr8+SR8f9t6R6GmsvE9yCjY3X224P6+QXcVMYLinQmpsE
GOctimnWkvI5pMRmtxVaLMKoTt7TuUocfTZfy7EK3bsKPGdarS4ZUDD4qt7WBHPhXu/EpJonE1kh
iy8tY2hcPQyFG62pzi/7lRwEagvl/rqKkjk78Zm3tWhOiYKR1JE84CrH3Ru9Tu6J/26ZyjlVMucz
IlfD6iOKUmrt4OXtZMKMVOS//ucsLRRoVRo9jjq4rU5bANY4hxU6tFxsKTEL7GlzBknjOUP/AWnx
7znWDR00pYN61wl391MY8rAxJs0NN4lVXtSIbWRkuurEd4Npj0kfM4Q8uX0QG+afkToftWND87XP
pxOIdMLsHmK+1cgDYDlvGZSvgRlSeeiUtYUkUqcatEIOB5/jrisBse6fWLiurewDNKAYkmVwBEZl
894j5T8UxR3M1WU7TFzfSGr+k7JSOn5dioREcWsi6rhcAIk0WwZTzZyOMBR0VqUZWcdqy2vNUhO1
u21rDfzVNPgR3GyepeYZ9LonNpg5PjrGfXP6pK/0H8Dz3RqMgup3dQriDXQYJrYRDtw4hA7vmJSL
s1+gex/F8sAJ3RLOCtE+eMf42G04gNDq5bnyQ3FdSG7bYLUTkwvaqagS+hnVui95xgjvMx5V6WwT
3Y66D6FiXL2f5f7nUBW9b373+okUjAR+gRBCWM16aD2Y/BtO6zxMzGCF+ZEfKSdYLl9yYuiXSNiZ
xgKaRv/MtGef086Px1QZ8EFIUzx+BvaI4MBwU46PJS+6zVdf/e/9vJEc0S3dCe5GBQ6cLBpjafUT
C7CB/jr+wV+3d0vKz0Iu9XtEf2pmbwKtRgNYqpapNve2VYF3+ZjvD3Z9NlMkD7mjwTuAs5Qtfjdw
OdTPfgAwLnVawdSVCV3NoRk9+duplZbKVNyJ9gsB3JKNhHw7T0Hxka6oL2PRriVMhJXlOmYdWOpx
InB84AyO4Oxr+dRxYBWT0fHvxk4u1ww3J7cn2yDbO8Y21zFKz2WczKkN/0EycP7OGLcRJ1P3ujA1
Lt0NSsGSk4X/2zg9toCxRSolxbkVh4AAtgpfsVRW05I6N3msH6O7k3KciwtBA0w0azGsJrZLdSPr
LJ2BwKftb2VsGHjksmM8yak0NpliGOx/DGEWZZPk23wGFf0TNfJ6DgMVB6TPTJROtRr4BKYKbmYt
ft59JF+/UhCFwyD0aHpQzjaGn/tcnlWBQoCon83hUPO0vLwqBlraqUwJgC+trDtxd/1U0StE3Nw+
vrLQPohpL7pLEojryYEFmSWG+bXU0XapGPNO8rifa38jFFVlKYiiG3Jfa16RNq2KRHEWX+HytdrV
SYHrvzFjgmuMtIbwaSuJLQtZF5hcMc5u2upa8gww+paQBl8X4J377qL3w188NtgYqQK3Mlwy4WyL
pBIGtWLzgQnLpk/9JRwIrnFY2AeHTAQXJb6CGw0doWxodVMNzPdx65jSPrnFwQon2A+n5tVdNm6l
fJ2jY0WskawfOtGbNZvgHi00uSJgn58qiiwYmjsDoWTwKbqniZQ9SRRXCe+ZC5IyxNOwawvb1Ilb
xGazCqs22gZr/0vNf57GLM7o/3i5A1SWDF/Zzy74Y+F3GMHpFn5KvMEhbBXqYNZTI7L8Yd26TLXy
f3oO0JigH5UjQ46xJkpIJ+siWzls1xXDzRMyTBduCRi7BGh6hp1NoDIG1/szg075THhzOvOa3ed6
UkWwEvLK825QYr2jXxriS5CuK6cvANDaChX7aQIGdhW6W/wJsxsYi8ymnzFYk9OLEthx10FNUkeg
oldvZiaYTvBy4NSk4CNIq1Ib93N7gglZd6nPKeT5oQxRs8evgFrzchgBu3NJmMXNGLaB3Kn/SCPE
KhwiThUwjAgjWiY5v42ZI3bErSRCRbZmpg4ZLxv39CnMOcz9FIAH6g0U3KDUKDmD/3Xl6FmcIUxq
Zbihigp9lCyn4ODMBW5jBR2y/mUop7jeBVcd67cKVsaAJXAdTYqcsS2k42J7jgebB4Cv0TdkcqER
4cxPRv3bLf983NIGxHKX+WdjIGowylHdJz69rU5TaEJZuKQOwf6b/00KASZWXYaaLOyr1NukoQcE
UmOt0DpZtJ1qys++hLXUg9Rt4hW6NPi3yC+IXnKPJe2I7O9EicSS5Lyesm1yr0Off36+kpLAFWPb
5BgOhr3jD2Sj4iblhzFtXxxi/nslKTv3Y0bJHxRqZ1M26q3g3GwJzZoCZW+nOf+VlnL1wKORqfxg
DcQNO58lOfWCNF3v/8lkWbLHcuYR4jiYDElRvCwlQG2h+ZNHD+Y11HVu/j11AkcvkorLW/jpqLvs
kaTdZBnL9eou1wvfl9jPdk4gyFS+dMxhtIsjDVeGERE8mpLwdAExrEgOwk7gKrkEfYcRic46OKEU
dzxDarU58ruvZF9FLqgsKEzXuVaX3pIRonzmZ9UAIoJjthMN1lNU1FCt4mhSMV6XoaNVCCRNv+gJ
zMX6DCfaI2kHHVgSBcCJDrrh7kW3uuMnKJZcafXeVWnn/xmLiCP1gtMEHB7CUIIeAMgXERwTpkhx
sMAi6M5urGTi11M5NqZDf8u1zQeKXz10H7QuzJBa8v/PynjTQ4IibtwzMJtMzYU1DrBR9rw/7shb
YUIyn9ZgyYJQFNE9vvlrCK4SrvxjodinI8ZpKZYSr/jV8i1RrHphUjVYX0//rMUCgz+iPYVLduwR
FrWYdiLNKOogcKuoRrO8i/Y9FOv2YZoYg0bXPqUwebAEWXzeHMzQ6O8/wISMbwcde0Oc2UaH36Ks
M0nUlli0PdpQ74wtQ8rYtlxo0AYmZ1ENE6ei48s4nZ+BNFClhVqcM4abRUOgYz+IfhpFYqbRBcCa
KjZcl16apKx7TGD+ZZxOsy8ZGjsMNOSlsRk8woiskU6VpRk24OsaHs5gowMnDzyJeenNtTC045ym
GqcSF0lf6IJiJw5idUe/UDDfM8WTGzsTXmS99niNQslAi1dXtsqSyM1gCajC9Zw9JCNEB0RZFoNA
Axna1et6dlmP977/K0EAi9ONBxRLKyqHLtbpEi2jj+jevi2pV+jD9b0R5HdIPrVowjqChRqRpCEa
oqP/pqsFiSoMeeYJGLExPyFyGdFH9cdoSj5lmwZaP9etbECD02AkY1UJ3SgnsnZXiWTVbHdqycx5
VQUK67Lx58WzIw5ExpP2MhpI8dg8abYApNOAB1et+D731dxH1kQ/qcV/ycyWAXIjA5syRBEx451e
LZ3Ka9czEWN/wbt2EWpE3PhzXnKeu6XH9YQ4/OFwqD3Q4zN1Kn0fOR4tTo2qwKNxfR0A2cuS1OQG
DWQ605kRxOQX+G9AP0tFO50xzCewy6YtvoTsWk1YlmUS9RMcCdgYnEtWP+XQhyFtFTiQv0R2pW1o
rKsPr3sQnI8OkjCglIZiJzrfWFioNMAiQVnNp6I8aINPYV+UzGnXiFA6fKg3G+EwxY078TeJxtro
Il18IFCVgtPSicWymBlXRa9fmQGQKesXln85z2bJjwb0B+oHdkxfcq/sH58CVQO6mVyVVLsOyH02
EuPWjbpJv2tR6vv3oM8GEn0PMDzU8TU8rClHcxOlOy0TXZ3+ddJ/e9HOX/NgdjW7HFlIjMRkO1s6
k9Qo+DiV2TjWTdXkTrmu/rwjiESy1HsDc/Q76zZBQS2Uhde2hKBsSvWtry1sVviMhpK8jIvxNi36
1T/k/8ww/bm5WCw0pQgUaaEvLNQ9h/LcJ8J/JhN8Bcv4C7rOabuxJRSoGpb4pMtt7/HqT7TzCIsC
tVoBJlRF4o3tuXc3IJB4qGxO4qvSqIfbaZuqQEEEdued1fZv048uDR8lS+hfybngdRd3LUB8UoLn
17US0uLboQlECLiFFVP+4ITm7xtjxOhyvTyyv0tLLFYLAmn+twMCZA5kyCaCJmmAga1o7qMgJB7j
UrMxcaMlmkNLemZC56RuMutHoIdpOPrXoOytu2Sd86nSdmBB3CEE3EPvCpgSM5CktkV0B/+/5NSm
hWVyXqf93JaNsMI+YqTstEVkfZjqBFDx5iaACGF9P5XflZ7ZMVkl+tZp6Chtbo6gBS2AgdYabvuR
GkwKuRFelC4iRMUSargeq5ug2j4GivNXeF6v8tVBzTOVY9TpwLembowhbMF0pLZbeRBVsInrRNc9
Yh2AAUtBYRsVOBLjcJpdIwEqCc5chou7PUpxFBMWomUf75llkrUtKmOkvHUSL/ZSBtz3GIIwgm1J
cKBiSzjiKkeDQul/BxkXoz5Msgxh1bsJ2ZUqlWVeZC8pP18l5/zGCbxi7mWevmIsGpDNQJ2SqdIA
yu2emNfs455lvGIVMcnuItcNYY/DzB+Ww5YubEIRJlSBsSii3QaKOjRPZuOJkFFte6OpOi/3J9d7
ByLADCns52/VacNoqfNGIRq3xEoM0hYhSwuICtsGbEI0Kqw1OTfgUvQczcnZ+aLKl6O5iRhdhCLV
RmFJnZ1eit0t1x/j1ki/bmQ86pv/4m0AiNrAaF6yKvkoKAK8pzbS6maqrcDnrGr5RlFHv16bjwSf
iw5yQjJ+c9J8BT9khxA+OvTeqpFKJQA1BQ3fWGQXAgJTy9US+Xx1dG5JqG89y94q00qh5tuU+KIQ
gpIAhS88BNrGSz9vSozoRUZ4Vxqll89X9ECBbZou8WYKZOL7bJeAf7V7XKU0aogxm7j9ZNakmA46
TdGVIvAc1AOM1MUfR+6yFpaWHlscEeXYleFsudmW25+7L5T9hHJFIQhM58NS7L8vA64EPaXvPm/Y
tac/8jy3TpvUV3e7+76t1h+XWN/mkGNZ3oPw9TQ6Mn2H4x/OrmUt8pvJagqXxBjWEHWFWv2V20cb
onpyqOrItuRmAAXqR37W5Pq48hDQEJtf3GkwOuMAmgZ8lavnRJhh0hlUe7wxmZ6/g/2TaRbViOAn
pmTR1Dmba3ca7iKzx0j5O1I54uPT/C98k1RSb7+l0psICzuifVVLaec1cEtj9kz0Al90b6+29gm7
go0kCHlu4FlSEDteMQ++cx0v7T8KA7EX4ZUkUySW3pm7ItW6FW2/2YcIgWPALm8IZfDhNWmwr93g
vutBbBkryw1NlBcc3Y7fkjW4y6omsC3xcPysVYioOUkzjFkjKS7He14D1miYF69vodonJwpfeywH
G5IqTNCsP7K6vwrVcf/3Dy3+2rJyhF4YLRjIbgRP9q3EVVLY4+bKtpqiJq69hczb40wQh7YmgdTT
Ymgq1yOfU3hwVktqRDEgmPLqlfEXwTbmPERwylHrRhcojxzW5KFH71+XIGEz7cAxkjRHUh+YPNty
JCtR7lHkTOpuN8v4McUot9UBXTNT0c3nGavL7xgc/985clXQAWHKkqNdx4DvRtUK7zL1yJkEy0x0
Xan2uZhEu+/QSYzXWYGLsDBM5kFHBQ2OMQRdixJDPIUtGuhqjXvqLYpAaODzq/a+5/Wa7uVcR8kv
w1unMMJ7dQywJga05VS7G7zc/d8Ew7kqdZhxR7vO2Jue61hNOkjKk085IfZhuCbG7ksiP7pp8aJ5
AT0tJPxajS/6vQQin3qjT63EQRjmuT3csdck4FqkmTp0OV/5/Ge95irlxHC0xNELHAqtWBnhKj5s
wRJQetok5twNhdzjr8961v4hpGchhP6DR7QewcCtAeVvk4O3RGcsKbNuO9S52uxb6vv6Csk+4m75
SKH6UELuuqWrGyF8UWuFBqbER45i5OWFQkmwQU6hwMRKPB0BTRxVwk7PzSn81BtorilywEKReE1K
qcxCEK3AI6WkOXG0qycFJvkDSv4K0HwB1CWXt7tnT4I19NXX7wH1U401bcKvkqrjZ3meBFAhQjly
tq3S31SbchTUj+s9MpGI5YgjU7R48svRqeaDBLKkPowZ76IlmNmZo0yvjRrUEWHfFfhoSAeUu58g
6eKjjZKRLjbe28akITWpKE6mxd4Vq0KdUX+JCwnVl0x/nSA61+8G2FN1nMq1yvxWjL11ff81S83k
9KD4xlftITgfKjLqoWNVRPqA+IIXrwVZXrS5gxa6kd/iLV75lkGp55CWjqMOyqoNmr2nOPNxdqDZ
et6B63sH4t7u0YBpiWpyzBKVhh9BlEt4WLcln6RXJn/jQOYjG7ox2WKFbNuZt+1ScjJx47GI3QHu
Y7t+E2DGLaBGqx+k4HeqceVu46em0wIGJJYyiZsiPsjrBeTjzSGLCtNGsSs2kFHoe4RYqbktl28j
V9FKi7dwD+ltqMnHoliG0Vzi1hKqotq72TR8+Vkdmt/INKnh0n9BtgcTZQu9VP8EXXmHNQFTg8pn
XV3rLb065VfJcFcjqE336ousmqMdX3atF3BuiQYBaMywq3Wky+tYXF2d26h/CnRt2LCpmV700xB2
9VHHNSEcYkisTJFjlhIim8IRPyoXVTcs46PJA693faa462Njnurz3O/BnnTaNKlt34jzZuXwJuzD
ji7sV0uRxKbjsnSaw+DdWRRE/zS/cwD9fSapPr2M3WUDHYXFrLzA61GkhXHr+jdCzx1ag4OIr+Ue
w40mjj1aUNYVZJXG388wFJjhyxVoaU36zzSRpD83xGLSTEUuASIjbZXCBHKekqYI+uLrgtQwSJ5L
kdda48tM8nlq3Vb6nkMJyonbJAv/2j9sUy2mcGhjVjJQBaVJNcRcJbgF0vFcQEC9Vy9UILvdJ3Ri
5ItkvlN3e9z13Rbd4lvJmKKuRHy+O4/fkjt1INIY02z1B+NfVIutR4nvA5qzgSrUkvFGcn/y0zkL
uX1TCZ2wyev8e4Rejknix8ilMRP3GbG9YKfjOPA3jVPpgWhxtgNQNpo8wPDdbzWPX7grtarbpaI3
v71QYiy63pNREGtRc1Ha9bQQ+VdsMDB0CBzREfvsorF4KVmezPYzSon8UYFa6qYr5eDqCCBO4jDb
mIq/slSrzeMXFQ49h2lXz2gsVpkW2zHQyFIxDuYLhWE3WvWvoJ1QBIcKdGmSkM9tl+dwo7+N+0L5
+PZcoA/BHGxl3LY9mguK9/OjEaEtx3k7PK1NuZfbylBfAhyNPvMwuGryU62zIDLarcEKvMq+qEJt
Yf6Tofsh8cfKQCTPcPakUZJB7qD5Ev7/F/0n9OJu85FIhRFatg6CRQxKIp8OtZU2FQO10l5nm8qS
MKg2mW+NSokINy8AsSx5/vmO45+3p4CEHpwA/0cCtQAiCqfhxZvtoprSUdBlOj/B11g2TWtR1B1K
NJLG8eCg7bqnxXSQMCHTG/EfqepMacvy5+49J4Hrucbf+QqS7FVy21pT3MMDw2u9rhNVxPWtUyGl
dmsASaeyEVRCotsoLJCB+DAKWF+3P5AJ6ngDX/KCnCzKlkc7+MbBE6OZKZ4a4OzjCrCcCNF4NU1T
u6iT497U7/3ILopnNW53U+kbO5YfMWdM5TJody4jSQxjrPYbSvFpuwSuHNE6BMjfb+iXaGykxlSJ
1ggkQ47gv9naqYQP+IGfRGSL3F1dQ1lAXryGE2PnbqA6k6qA2UXK2wOLG3Nz1zeGPHAjgk9mrWn/
sIbPBstRB4TqdGokNJ4NuyupUQS0Gs8FrxO7d7surAmO73cIu3m4CeNoLksRvs/Yj7dZTSlfjP+l
dPRNomjLLsSlGK2KNLtW42JfwjsZaUlfIB2tAF/w0j4A8mEgtYBB05PNiAj41H4eq8VOQTuWLByU
ulX31N7Cg4gkT5jAexE4QvrT0dzP3VDPKHnCC0RYU/6W7YXWAx+7/1jJFOAF3DOdc8ChPl25IR9j
EjdzWvXGJTDcAGYLv94Xrv2hcky8o2EgJXdc3qujyzVTbVrDFMGMpW25TTYs7mnFcaYp2pPwRnyv
mcvj0vB8bf0u8qZhhKHhqovn3rH7T0dLl5sY2ypucpa5iUsQyBuX8vUQyYB3w4fAzQKI7oXdT3PM
YrBZzuhBtFRjpKU8s04QsdDkQfRPIZpfdeXKAT7HWu1Gn5aGsOMXvxpdfnck3QbJUQ+tmD34ylMv
BDwiHPV+BPophECw4mfmya7vwWlV6HqayVzt7217uDUT5HwtWP/CsKa/n1VZ7KOVGXnwPGerjsCO
CS5Wsw8ocgWMLj+XV4dXIFsmNs7eK/TkCLtBtCMNpB0gUrkZyztiLZzJ6VkNU8Ahtdvmr4q6rg06
GRf1hZu7dkvRwB8aNM8fXwIdJLybfHWc7X+8UhhIMH8ZS7PXdCCGj0OVJ4zBoreW37cU8yOPcXUI
d6gx7n0j2rfMGdPCWgTktw2jHhwwvuCXTD/fBOZRM+JhBs4ywE9sQfneE9QBXavw4ugxrqpNV/CQ
kIxdJ7xbqBrC1iyHbr9umA7ER7uKFbAiXKkBb8KkZYKNO3rT/eecmOefSvde4CgcR0OI2sUepM7G
h8BSaeYhnH4AqSsJmOGSzgPo9e4RnwZlrFvDYo1bVEK9+ADQtrgFVrw8DWscNcSUFj1rV+KbFrny
8poS6xwAW2LwfAQ2DeACb8vlTijSHnTjT1eRVCfbB2j1yx+V6XYF7173yPkdkmDM3gmskkrKixwG
/hHGlxOwhqW4bctuA0CPin3l8GzpgNf75fHF1VsszU0T+7+nyT14Wikb/HrYwnHCNp9UDOg+meTC
D7yDahqQDBRNNwlVJvUzv15lAhzsKo5G8hyk079qKUTt5hyzZKngOxzMBtAs8S8d+qTYeIjhZi1J
PuTM2Ed4W4w2g/2xpykNn/gvObl8/YUPNdOW8shk/PdV3ompXel/sjNm+QmNZHrHLH0akWLfa8T3
dXa+86uOZp3NVnoMc/ryAD0rgTK7cw4J7M08RSSevPJVf1dgth0/ZVlfx5BvgTipO01WBLjnI5vO
u+x6fwPVDaRUGHpYS1OneIZZAujCWOorbYdTZhgTYkJ01SKoGgm3jVqpkzKqMf5HZsd4XCutLt3K
fVtYUm41csmfxPBDC0eonSAkQtvU+16x97O/cQnkHrVMyOSM6RryZC90rWEls4evHHRn84q8v+Mp
D/L4sQ1JSzMZg3/xIifku5jto3ZeTPd9Kujletl3wWiZRxrylTIXTgU4q1uIkKkePbkx4OKX3qUN
pXQXQcXE2D8bO0hWWM0WICvQqSvEOOJvjwflwmlvY8SndTE9LjYSyjTmtkAHDXgMtsZfrZCLa0bh
GSXtGAnOp8cPGsdFg4z1vxN33RUB/gF5GGbJQpBZ9PkMfSD24G1VY8El9261RPzOksvojibjuj39
x3us/gWJ9MaJ6e6qZfMrJILaVAEcoPCvWFx05Qk4lZBuczpJD0hcDk9feRZgN4Ane1541mA/7skD
Y7YoAVagkhdJTZu8cY/1chXU/3Xf6I8VfOxDnZTjQV6wxJHKq+TebSz1lDUOG1qhk5qiHbWzvLUq
J7OdSFkIBzWM5wcXdsT3YEIGb4eedYTSekAkKd9SVKqVOgdObWbeaKEuQ07RHTzDxH0vyXOsHxMx
AVa2FWDRUEvn8UBJdI8SZeTnVnWcmoMhk1RWf1gM+oKKYaPdJRKsc0OAmbmeHrrxruRyizH6zJxa
OakvHNHzlsUbAt9R/yLawd0yUs/YzWBebu0nIVSlsPfb583LJq7gppFY4ZXiLqraou2jyjFcG18y
PT7jAliW3M1DZPRlAIBjP6z4k28XoIIsFMbRTYuaMy/gGtEvVv0Ce0YnFS2Ax8RbnVwAi7ds2OxF
v4cwF+TH00VjXvh5OGb7ByEjXinYo6VZmyqhrB1KJ7dzt1UFQ28Dq4Ua2K9Y7N2I4rXIGiM7mltV
Wx8VSYaqH7wnv8h1ESD0sMBdo6e2yvz3yXPRyGchaiB1tDLhn7hYt9/UE2SPF0kzfoudriA8UJTL
jSMv9XPvoH4GxUKbger4F8jDXpoI6lRlpQpItDz7Sctyl6wASx8NewldaVAxuE26/ut59erGRqAC
x5XIf1qrGtJm7CBHuMvknzZ78fQpPUuV2CZXuQSnkfJhuLoc1URuhiXVsSr7H3wq73e0GzJr1vQK
pniruxIg7lOfQa5flWXvTpMKBIUSEjIvZEccCdEDGXnkmTy2tyN4EIkbSPFJ5Qe8teMGejtNNNDz
9S6qDF2sLf8lSW6EDCDyJZBnlkY7uU3eZUm/b2wq4JwOs1DWGQJvtWYkhLpD+wp6F5dIVvLR+Uoe
xHdiKGpvH7gVJPOeIp/oEPd2TUlvFrmkZkmscOyZOPDr+Uo3bCgqA591b2qOOLTsGAsuZlTVB1bR
ys9F13nL5fHFW83gjT6eVEpJotrXiGJG4Uof+YDAUzzCbemYtMffL7KYdZkygl4i2kc/wy0s3voC
oSAft8U4bjfgbQod/aHisWzuv2lnkqCrwFxu7Ocm3xAkcWiwSStakt1pxQd0f2zJF9IKWl7YuLDQ
K+WSGCYYv6r4J5ORU4t7KhFX2qh35n+QJZwVhSQts554LvjkX21pDB9e37B6EoxtJ4bgZnYdpH8Z
VnAjMCKf0J0/p3zXCrkPtySqMRB6Z/bJ3B8vwcHEODzD4EyuF7NBmrTHGisUPaCOduNI9gSxu/yp
+lt9cgv3buIq84gnRp+q0H5K4IxV+xMWVLdGCHDyRLcrVgDi+H0Njcn4vL7/Fe6ipoG1aBTymObs
mPlBAkKzIxDA/X/m4PjO/x1yXTdDe/HnvT8bnd3sSzRGgSNAfi2iWABb0s7CS9WHqhVQjqUF3CVc
mxz1WQtoblbyuIjv1SwFkbhSQETPXECT3jczh6Aup36N8BYWgjbHXi11B3AAg8k+AzF9aM3ZikDN
c9IZ5vHe6yQxmwqPCiFc+EEcweK1NbShS3pN0rctY0idbDAYn0vrKkjPcaqi2ysrBpQxTvaXyMOM
7s5A3b8ab3XVvEVx2OKiZXVXLuvkmEMr0dZVIP1gGw+CRnzWUdMxTHdjMkCN3nJAdwHE1Ef1qa/C
b12LeDcEaB5Qi2Dp6lSL1/MWdsfyXJYs9BUewdXcUii2a5Z4cghFWUJ67EIt8oQsOZPblSepwcDv
9o9/wdrbY9kAMrfRaw9yq8vbj44h/p9KOW4t2v2ewP2qN808JG2Wquxmd8MeAFhow9nzxYk1E4vQ
K1ldezsC9cnfpR+R0fOHxq0nXus2C36pKLuPv88BVK9ewGdi8JImEcAQzhRbjLkTVkGCZKdiOJZu
o5tU8kPIY8jL75I6s77wNIxPl69q+IFG8ydNVxcL5CGbigmrH7CNKPbgny186j8FRwEp0zwduYSn
hOF9cfC6vl9bplhdGUcM1Lu258M+CxXdkp/CdaGAFUV7xYUmIeT2ikBrwC4GJuqqziHBaRRuhTYO
yZo8r5EhzmpbmM1j0Qx4WK9beWFkRWkhQ68OHth2vUr1u5E962bLxOSqSwWwgv1VhyxjTqGYfuM3
Dhw6GDdmXK4QsnGa03MaXhdPtrob8HVjoDsT6118dG/1mgqWGUisIbuZf3JpVz8mnRCkXTeknvVT
yL2u890o4P4Q2tC7Kl5CUC+lOEA+6dkSvQ/OsDee06LmZZUf2O/fgFouHnNlpT8p8dNI4J25GStJ
+iLzNrUzg+OyOBMm/Ad+aE2D+UeZ7bpgiQkjypk3BXxirTExhmcbg1xZR5WbuWQ8WuD5scOIo+5b
HADVRZ7XBRaxO0evquQ1HjyAC42ZapwpAspfhlSJi/+AAdmz8zEV6x4x3WTPHKD6jqTr0BS5L3KX
nFI8RAB76JSEWWm14bUgN65+FbATF6ir7pDK+DPQfQ4Oy9sWuNvYAdNBauXd2UM0noevq1+viIbG
HXXEI5n+0P7HeI4C8cf6kkshjLoM6FcNbxRv+KlNbNIKzoN1qBwOIrpEvEtZb69FtnzqsVCkDhM+
zcDMJ2jGQaIOPK+IDTyO0IVdmQUif12eaUxseV5ta27Ld7MfHVFh30nWuLgiUkbpJv7xXlpa8WsO
ndfuD4SikOEN4YKuSnXtwjaexjJppuYeBPkZc0fezklbbzSvl8whgn472XEbwGB/60F8+JWL9dO4
47NYvGzuMH38gD8YtdhUd+2MMaSfXpBptkB5z4Uzkm8j2XqjIy2sz8dT4guY/iGYS8PpLgQceXXo
TSQv/8sNPlMJx6aYleFNMFgD5KprdjR78j7pOE4+8yv0zAFpUcaqLyicQNxXtLetKKUcrUntBm7q
GWk+aiBmRdy2WuJ5f8tiKdoREiNUB2ks2xKrHSEfb2YdmfY6/ufQAK4BZXTTbO+nKPa4bs1wsuMF
F65agLxz55mnoHyceBzMcE+ito80cA2zZnBWPK8ufxpvejfIukFs7WqYj05tQMN+IxEdZPhIkrRh
IM4HXahK8hYDx/c1Ad6t1odxmSJBgKdro8S1lgNl0zf7ZzswfIerpMHD874juKAU+G+Tb7EO1VQa
dyrzq0Ri27cmMzKV0HNRypDtD5nXzz8KkYJBlP6YGjtApoX76STlXhiFSs8khZKgKhBtKw5wUkT1
DP53EcXmk4xZCmKCMD1En34Ac1tfdKhuCE6hUO41Om8I4S6wxhfVek2JX9KTQpeos0CbKbVRPJuO
a4vrRSonVhZQdHCcCDcbCTfp+ddpTYlgE/M0tupKmaulHaFgRD1GQ4ULDpmUTTqoGCeH6jQzNBeT
sQv5dk1fKjnxI+4uvaKBZvR+F7+jY+2i0dZUcMQas4F8KHteKRcCgES6IlszsJ1kJkFEJx40ddZY
j23LorMnB58i8YzZguqxwT29uiouDxT0lCQinQHvbAO/bpTGwtiPAriV/QNJTA4/8DFe1KILLJtC
ESM/AghY49l76Vx0N27IIowg86+04SIxoEvRXDycgiJcurSUd/P8WkBrFmKeCDc2oX30JQoYjZfb
hz0zmfuTCe4eIiWyLoRUk47OgcrrtB84Zb8IMT8OaPcMrXkcFHLAc2u2ruDmj8l/5peVQGEW9am9
42CCKFen8+H3frVcD/dbOUOJtIlxpWEAuMy9HiO/rRipMf4oughArdfSf3Nr8pUfbsOI0xzcoG/I
zY17h/OP5vjNxeBwlJMm/o+CskTh8VsBBZ8HDwLkoSFUDue6u5NGfL7LqEklV2akwdaEJQpTWe61
rZpE6QlqP9Mg/KuZvL70czR5rxRcXqwdD5dM3dXJ5LQJTQa1gO204A1aZyHTbY0r3XleEwsbm12k
ms+AqmKBHuwLpXA/DAMjj8AvPL6MfIOLrjyQsG1UAyFUna9epUx60ajVIu0Q8n2QO7Fbyel+xh6X
kOAEZuESni6xBKcgf2dIL90IJFBq+5LPg8UPz7k4MQLE0flfLV/XVqaDbNnJHVDyESIgVujEvJ+d
N4EkQTBCx4hDsowjj11KwIeR3GR8HAgY6Rgv4OwKATlmUrjmAk6mNysknzxSckdEvMost/8Mj7iO
J08wWw0B+XVSLjIluUl9+Rb5tqwHeznJAJqeAu1UDzx8so01m4uI8OL+eRYNJwCIgx2oOKannZH6
pIpJt+q6tnsYAKQ7CFedGdvZ32AYfr2LK6cT9mBDkAHBAdsETt4D/LTbinmjGKcE8bN1IAbHsdua
+DxWFcZwEbW8aeKWKpLfECPzTJnoYtivS1TdrIND22pIB2ujoG9isUzk0iNggZ61TDkYtHNOlBby
SKDMsBpgoveRw0emtBWiQtzO/gtFn27SYyUUmHQvlFtoahyoU80HEq9c1qdhHTChiVoP8xhf3ahN
AhiIk2nlkduoL/Y1aywwe+3ljqbmn1/1Rchj4vlHYXsd+k7mnTOBD05AD+LuLANKh/U+O5q2JqOi
UG7zHWhkYBuKrPJ8J+ohPCdmJ7WlowpwiyJV2JZevLTLd1z43eqECJPunXK43iBxVuCuSh66038z
NSKhp6nHwvD4AFR+ClNDnqVxSLQEkQTlHlsKdJyjbKmxb86SzomGaa2SG6VwG1Itjt3A9w72pfiG
JpZTOLpKTJxRjMfvr2mqyb87ALakZqNxtLzjTgtZtVgK3WnDPB0FB71MA8QjOXmCc3BpWG4wzUKV
Ra+702aOWR6/H1JNodcBr9fomGZhEZfF1U1xboYzi1pIinlmfZottR076L50MhOrgUHh0Njjlo6W
mCrdQYlEgpvmzRm1NL592NKMP4f6K4tANARdgGOvR6lM8PlAdwtGJER58nSHZ36fKoWnacMN6m4S
CiHPej+/Y9FcKALFZ7CSnPW9Ayupfk5UX3KDwkoH2b6hdywSLeqyJEfrJDU1uoD4CcNQMb6VfxFQ
3dM3XULUodMz5XB9EKp8aCfyTwXdvqx8vCGfr2d9p6z21wPDhucHX7nzFuTc3xSWu0ecIdGR4jBY
lLOXpFCr6dyWmlk4T9Enxi3SJfOMpt/AG6gqZYUoviX0UksosyuNW3oaMUMyoh0eHOAb5Krxym1m
huKbsu6Kzaq1T2EalUefIMNZQqKDUhrX85VwCEsoj2FteOy/x3bd327Pgza+Z9ulOhlrqiEx82vu
ZBcSFLu66tVYJXqFTGz+S+fpPvDN2uRqkUTWPQ+QYiCVmOQNvCAZpDtF2JKl9h5DjiHzMjhtEjwC
8WWkfzgDSQ8WM3yoa9YSDpVPM5f+p0SRtWPjtcddzMfigxi1Vvx7Yu5uMW+HdMUkcl/ZmGoacY2X
tBZUQXk9yk+9Bizh6srrdOU/8lDd6mqgTqN7ot0906zjxc7NJmZLbCriLK/yMNRzgzzl13yTzr50
xTAwdwpTxf9NeIJrP+MO4WNkx26IOQJaZMHSiNWqnYByKm2+f6+eU7TTy2+481sCITmHLb8Vvs9H
4JlrBbJqxQY4VdG0TZAyX79uRXpYJa+puSdkXtnCkRaJFR2KlXD0XqupHHQKoZTlE17XvZ2HMc2i
8thoBdtv7Psp1FF9ltuQiXBsDTfWWJqP6NxhHhikrbwgHIMBLg+o3YdBvR2/t7UN8zVBXwNN2nCa
jYHy9l2zl6Z3kkSCwOdhbc7rS3tUr7R0adZrXWLxOb2FZMf3PuxNKuQxvXFS+jZFNy9PIw4/i8Xo
+HME0S4iiZqDxh7gHh/7wRtrfF4NNNEXaXIvU4Mfjq/OCgqVFjOuQbzJu0lESx4kYKleVjanDZhT
JG7Z64r+h168FnxN1ZCCv1FUD3RleMpCv5USp3wIbt6j8MHeNPlOc6e0HwwGAy3sOBjyuzLzeBFY
LA+5+xErZw9wIqt9bqfNej5121uNITWVivmUjclEwTAcuP+a/anx7P0jwc9DcZ+/i0DSSyZ1/JHr
sHECsXvXDMwDFx50qLRYsKwpNkJ800B0X0R4PcTQeORzbI+Z7WNdnA4Vq0ustJuPh5bCmsL2JfSG
AUXo2F56FECTHb4zZG8CBN3Qx2KcjQgLAxRYSxyRJ5y8sMu1q9VbN/WwYx/2EcN0yNBWbfv4S3VY
tsEwAwtosyoo61r9WMWZsuM0morzFj3kn3kAKo9q9l4zFbNhF+FoZu7rcm9IvEzm5//Nm+n+ePYc
2mgpf4W0sj0P8aUE3eWpz4m9TEHSc+1+G8HkmS3glYokXtRrWqurJ6uicVfD9vv8Y0E/RqyktXdv
93j4acFuUPWmBFzpnL4potuMNZLORAGt8cM53OMJWEgbuCPTw3994VIINyvWQmZ34hFZF+dCWtXc
dpQ2bfA68tPpx/sKUo+N2yavGDEAZK0dfSUTqFW4gbSyzlilv99kJ3jkamRB2ICp6elRbNCdoOdI
LwBsWPCPS9nUtGOX1t7tceACPGU3DjyUXn2pwmAA+ywbH05JdTsHUr28wZrdQSJ4URmeL7DKoGjc
n2OcmQ9hNPpYryL8peMa2eQ6oGgKHbedxatNcy49OevDKKFwx3aD39HOT1oiyG2Ff+ReyqEuW+mv
PALZm1+WE7Hd/FVRBX+jsYjp9JdUozh73zCBLmDWzVqLIJjXYE/vFqgJYRqpQI/34ENT4m7rXMp9
C/K2ElJOp7kJqKNSv0OeRdadjlNkiRe0hVz3u/OhtpIkVODWbfVhYzRbe+wrYw7IS9x15JLPZPqc
yE37mrbxyGNTQ9wNdrfSiDUSfAx8dN//dq9x22dVBjZZzm5Nrml+et+b1nIMpa4GrWxu+s7W1hdI
l/tBYJjkDc9e10IbxPSUmaqTkFdM1pF/ljH/AGGbydcqwR/OZDjhRxmzJRtjZ3dfNLlaJcAZYHxP
bN223dPeDKfaNFa/oHerx3G8mUOT3iDtiAV5eQFPD75bsvIaBkP9yzj1EU8ThrSVOoMKvqJJFCPJ
rBYvMklRJSaOBUCEfkB2dOXoddG4jJpVlz+4AGXavA9XkTAt6JuA7qdMz/r8+rda7H+AXP7lKHWP
0/aCmDeHxlLicmtVbCmCT2zhoaAczJ2LPi8KgiKEpc6oa3yim4TXPIdtSYIKDd/dNjNJwif9t6SI
up0BFCQjqCrTeUJVpY2vUktcVYHADIeoMGaQTJjpJIMgb1Nn0qU0XlUgtn/HY20nW6l5oOrCiR+i
e+fhoQaM7GYSi7pPSw3dhXgv/gbjV+gm0HVMHCBk/2Y5LEjXTEEyOpZ9qr1MhMEkCRv6lyRuuSS8
HMu+ZBBkyywRarVQmCViX2tHhnFM5ETyMYVGnP0Q40NIQEXNkero7rQX6Kt2GDs/a0oyhTDLHatM
y7G4vTDgY6pXY2x5DRzcvooF1ClYYIrXpgYfQhUrF47Fgs/RILECohnjvyBWDkwX8dW4O3JYCJog
iirVS1Pbz76nEfNHdrlVAXUoESZAptqdghmT4p1upMA4Fy1f1UE+DS4nAfTdT7oSWz55gSy9E3ax
YgOgqeVc58JqJSTKspPidkoRwHhL1CETgb2MBxtSd/gxJUi+d4GSrhhsa1TbFEs/RNtlDezKJoX5
LUBSR2VG9a9yVT8juhsLkq/WQVrTozL6VhmvoYDX6Qg5GGkC5k1sZLBqv2eFP3MwLWhBG1Ig7mIB
ViOhD6isIBaMSrRsPfTcoFnT1NPHPt+PbbArIlOppLS9JqbKeQn/F/jBE3Pripda5HNrUKPAMSgZ
sVsxKzwsPVK4MT0ZxUipXBEUUK8KaUdMlx5bofTS4zaed+BGOBxoRd8b12xz1Q0zIRVGsq5qMFqg
FedYK90PfYktuRyikUz3xeiHcTKjaSTntmSEfNY9XmwufkIMXmbyBY0Bv4Nq7UeUpiFOk18IpYeM
R5S2CwuVv9QKeL2oCwta2NyAVogPkhDHTCtzuqyCm3bkI6SNkh+C4ZUhihbuN0x4g4SHUugzPUpq
XlfZdAsfauBcLL282UzDE5223KsBidgiN4PTnk8P1EtHq93jytJi442NjyL+pkKvZDiatkErGscA
faJWAWHyU4jrd9NhKU3DCQgE8tih/YbesGZohrukW69m5pZJ2yxGegf6hIerx62fW2WQ7+CC2nXj
eHDsGAEv1T+oQmZmDxKqBgYspl8tE6UW8rwXXBF4wK8xPMd4nuswJ753fhrYis+4vmBnAv2LiFuA
RMRdvQzIxnVrOLwOvqKx2ilxf0jzYpTSUYrHgwIxfvf1PGS6tJbOdWl/VyPeiav5NjoME2+uwsEu
UWzmTriPfFUhAUFA5n/J2Chxn8GpNi5mzI6wpwfP8WtjpcuNpPPX7N8vS1aGqAuQHcprR4K93WrD
UNZCvvWqMNzYtN3mf2mgWH1c9/cKadDrghOoRfFt26xRNyoOrzOyRYsadDF4vB3HsDD92+rVpG4N
IKZ4X0R+cVH9VN5XP/eQktIosVK9HaUvm6wDeF37wWJsQ7UrFjmrjVQhUSEen/jCO69UKnRxI8ak
Z0WBEjf+XlPTQPtXwyTxANBXXa9kWw9niVGGgMAijOkJBo3UsxK+muLzz5n20Lmrjqsbjkvmu8WF
z4qiiK6vh03nRE1jvQncTVHAcYLQaxK0+akd5lZ14z4IPijwa+K0vV4e7M9Ue9JlIRKYQuSMfjJa
+txCs1qnD8JeLtRtX0k3FZiEKoes2VgUsisvwzz/dCAYOdNWrDphcuGu3OgkxLPw7nnvV+MadVrR
zEDm+P5QF0HBbnGnAsi3n56M2scTdYWyAPrBHVIQ+O/5Z9MfK2m4CZuOIJl8+/IqI+4mpt2UAb13
YJdd90yeUZu34WO53HqEcPxdmvmWZv+IUGU2z7Df4EfzaxQiA6tX8RwyNLIFSn/Yx0nG1Jh2/ENu
ZjrlO2cVz3TG6DTPbIqB53DLliCJ48aSO4WwbAKPx/dU8C4ktn65wN18zyPSHmO5Sudk9DXb+qrP
IPrWDcgoTVMRsDiaMG6S2tT5Ob3okKvesTgE9EAHT9uybs0G4aVt/+o2ru1W5HF3m8J/QCG7c1wY
vnkOYaLPlp+AMKXaqJ+Vr+2M8mnmMxV1wldMy6ZjDrKP4R9UfM1q5ui245DOJTSys1i2hbuJ+ZtY
Tdur9l/fmtt1fxcnhbgh88KFYbhYHno7Tcaz9pxRChiPIGLwvcu/qFCxZbRDFWpY/wdTsAG3nclv
MuxAhYn3Bhr+xrcYBlL6DYt+4cYuckpNRC/khA9Q07rycEJUqiWRh04vieFPmBsu8Rfv4AJCNlvl
B3lVdTvdxYChDTbFsFOim+NOf4KdmbGJJ2aYmB2OwynoTTMl4jMVF7UNddfGoyQyUssp0tt4twB9
2jAtsukNh1Gow3wrINPKnsYGlr+F5jJh16B7/YFTHrXu1NCVO1HVLsqvA/aBUVWh5UatsrD7ZvOR
1xIqwjl1LdnBenwiF06ZSjJH3yUGuCE+xAf41+5NAyCPdQQrS8BTN69+2bd/Z0tClG1EXGoH9Clv
PSF/EN5hOiJO0FTF7UpkgXF0nknBagk7Q9Fii3MgiPr2j0iZgPmdVLh2en/Ck0DI99rkhLxkB2yW
QhdtcRDhm+jGAcEmDhpvSWRkzWZlWJRyU8of/xGyliZ2++wvGi1yHpn1tvoGmp/BFkdCy9cAQiwz
42lw/3QGhRHSG2tdZe0a4ykxfsc6vEHNLi/jw7D4ID3PBBBrWbsWsrT3pxi7qGZSqx3JhZTnWzKz
9rI5lXcx/sgHqIaacqDdmBZJF0ALH2Qo9bVoiPX5YVAAINtoEZ5lW3IbjQPlJ+L9VaSM6mrMrH/1
/+CGt9arqideKYqx/v2hzC/6faM1lEJa7tlO2sz4PfKM4V5TD6RJstAhX7JxY3e2uEZ4rUQrekGG
oCwrf6z0KsLnT9xunT/75gVzd5NzibS/kCoGvDlSuFP2lYRmWJPR1RKtkMmFBIsq4cgN8ngUkscT
6AodkS5/CcC27ZlVKG8C+bGeVVfhNPww+Br8u4fgfSe9S8THm74OB29n1jqME39Fwe93PoKXbWG8
av7lhuinqybkd4BQiTbe+WBW2YZV4bQ9eVRb+Ku5qKVW2kem6dP1rsT+hMovPMtiiLHFsd/X557x
8bLOrziRXNMFXDk5TCGz95+JGcB8dbSTeuUHIddw+RVgbAp1TL6MPkyLevdFYNtCLi05qg2QV5Ik
gwdRPbhAej/AfvI3y4G5ZXS3FgqyIQ/4aeGrArvCIZLbxrk47MWskvM2+l4SXGcN4RkjO2BAKUwz
Dt2v/RBTGVUnWaF0BP3p/PusrzTGvbH59KaM0vttmmisStwaAU88Nr/aZmCNb1yo00gPiAIFE4kX
d+pibmuL7nNIG1DLAa9GtJL3/CkC7I8RhoS+T0kLdm7PWhvTdwwQQUYF51iy+7yQyqIfzUmzi4C6
r4Nb/03gkdXYXd78KD3vO6eWabaAM1jjYhXTRrJGzSbZ4dHo2QGtn919UU9xhF/gpirVlLAQqGmK
QBxjY1BLU23YezomN6hcEzWPhcTtVKzuRZ81NKbBeCnCXZ8PJExFl9+mMsDs2HsrYVIV8TCGA8yx
aBzKBBkHSc42cD+ml/67dvL/KXn5WMFulPcv3ObHvn8OhyyiKQ/T7Vf/vsfPyvikZBGgaHcSJXN0
IzoYH6TexJCJKH3fmfOcvP1baIOr2PpBydCgdI16K+utEu151NTE/AEGFgKBBL0fat8+XcNsOXrg
ExbKslQ4Kme+ZZFU3cmvjEXGdFEhl8E1etcCSViSrfYIp4F0Jebbef3ti6j/2BOdkYosrKCizFSU
V1a2Y0s4zKc+741MKYDpPTfQFVVq0TdqvnAA4zxpEG8O83M9H0czbaQQboyLJMyaEq3q6l53ZrDI
z4qRPkfHIY1H14JiNn2f54LnPjTmPkbodPV/BA5/3wI4XjZ8rxZM9MMy0v51UkjIwA8F8OygEU5O
h9R76jAbAmbw6TU0rvK2xffec7SKPuJ3HpD2W2OGsGiRdQD4aflTUjSFf2dTHYKFjox8meh5figG
tQDIyPT8Z6zXFqdlcahfBw7ynu6hBFuzvMoeZaeWRNNqoQSPAXsgwc21wWaLsMRuO7mplXiSzpBU
n/R7hZEEdbIEcPVslIAoJ4u0/ZTSV+Nc/viPasoNkxn3ejL/S0jft24SLY8WHxUv709GjnF7mKUl
OtFcqz+qQ2L+Iwqw1s2WfSiHr+g5s+7jDWbJG0Z2kUGVhKPn15v/Xdhz3AQwuyM5e2YJvdDvG0CJ
z45w5xdwU1LAs6XklezZ8tvWR5aHZqbbFmCVHCPEr2aHRPOrp065qsQNHErtzMijfK/bacUZDWWx
AWiQVk9zM81M19l1oHeH5PeLNJP+yQ+IjQG5QEaT0eMIiD9S4+UHK8QCB6JHULHhuH+Ir/90GrRg
J9JdwgEPd1zrQ0g+dsAMzUbc4Yep71LTyebjVga1buEEFRHxY26fYAky7T6eMl14UYZgWwRzdoP0
ehMLbuD9piGhxGNFRzdTLSMbaqDU8NaKRpjkaWEp3Re38FO9lDqp1mqmqmv8jtwO/DLKZO22fBmj
t0T3yimASOnivdwCmJFUVube2AcSr7Eo4IpfYmzim7YpYyQv/tzwQUmdDI+bcKcMwirSCSl1NHLL
eOrGZYaK3J2Z/C+hwLjd+vHGHt6B44fKtU15bsbPE5xQbFvVddY9xMQXSvRwSAlpCNBLOjiLxEgI
2P+VJV4hlM9mU7TgELlHgLzEmNd8nF+I8tx1LyEhHsE6VsGm5orvW9tSbriIYmCw22/hhfNzVRol
Fvjeb5O0w2TwW1QHCto0L8Ealjlt+lNnxCEeU0XhB/gr6g/QjDP8SqHkcN/CB0OcwjTRU15KmZ0O
jBkQ5dM7jN+HH2lnAk/K6DuYdPHGb9xzVIPnOcmT/pVbtKkX74UtCK6Hn+ePZiYSLnBF8juGd994
WoFPA97v08j3OW9GdBxOMuPmTUm9xHhc2FytepDlqudZZK40MlrRfPwrEPx/nE3F3Ugd7qoJ0WRq
cGmHjXqFMwaTGWY3Sj+m440VzU7EEdt/ymyDmxDUtp6SWj59cLvJ4Un+xsiGKWyVq1YKWxS+E1gN
qIl5jj1TazCy58XnSNMbnR/cNHVIsDTz+IHdVRPFS3Gz+H1MMPytbj7rY4QlutomttFJRrGAlg4y
YkGrYuxaz8s+Gra2CFUmTcoMdkhxTpZZeHYNbxkPEgEz5OLt7/Pp8NAvrABSLQVSec7OWbdbJBHV
PdzzGZy0qhBHMSprJ/FgzyrBcuNy92VhO/kHOArVLyJgb+NjdgF7GQqGVnCi943ijd9Nzyn7dGRe
vjjnFn1nz6f3FS8tsD2FacQ5TGCfkQqz3SrdcHG0z0MuOvascwjxeAvBugwBYRUgiVhv+/naJfMC
5Ot3LB++zGKxvTHYOSJL4ssfIxpb5JccOy5jW2dtd0nyFHCBagdGZ4v6+8b3tSjo3+qNJf12yE/4
O8EoSG3l/BNVBrsIXphlu3j3ST3aIfU+8ddawuPknifCf4x76kFbApC3okuUPkvT/yv5LAkur+xF
clnfPWnJhFiTV6sMChb0aWbezpKP+rCZ9Ac0wvMPhswRTeeSuLFxjMD3TAedI5eGqpcxQiPUAFH/
IrB/7W9pbJr1Idy9qAEgLQJvZlLzOJd5C6Sz/L4Fg2HKwMonlrTBBHZ8dnsG5PfktO+yw3RXrvhm
71TyiKJbyVYvCC+0+h80sXGlJaeVSq4cSOzAv3Nxi4z91St5znyM3d98FFd/qqu3Gi9+f12L260s
7xHPNGnjaOYX02saEff3sulo/Ru3ob1HEyI1NIvdHVuCUGOA2aevypkgZHse5tVq2yotlHmn5hTg
38CKDYxmGmO3bUBd5bjhi97uJaBODUZ6ADb+Bfvnuf5bdpYWptUJOt14nzwSeBwKEnbUQsN3Nr5I
jLvmH02GcflaOzZgzWIp1XmZrX4Invy0kQG6QrM9KHOFSgF1tLdm6sDxEMv/UggR4thKFQhoPir5
SAnTiFulaUaj4lNNf6ZwLFtagicxqGByLbPqen6O2CouKuXK8xgzZRlq9mLkc4DdDEG5+H0/165A
kbtMu8tWUWnsB3/q7BGZLESv4Oj8Jd40z6XOXcjMpWwYOg5o/BxvmgfIBiHuBF40mvhaj86PDhKi
bBIt8oMtzYyHoEoFcYS+FAwR5i4hKm3U+qwcOHcu25N4n6KYOptiUXUv0HMlxCBZXbjLMv7lVTS9
jPfdMyqGApOeRzNm3rkD6sk5kGwsOKSBn3golzjkEPqrdMa+1Ko+lQMO503DjmIf52mmhW2OI5iL
Clm+2AU2/FBq9u+1OrlmUIMswgj4TsNiLxxawayVMuDTjOsiRFEd3KWjVIYyU4/DC8MbglTB8uBL
pt2biRd/H7WF58Cn1yze5z2pDhEuaNv/tfuZ2aM49Gsxqpr0w+WB0D3sO8NwStJyFFVueU4f771M
HJgs+d282M6lpTCUmqAS/57wIBY6bn4JR+8BE+hz1nGNAaJ+9vzGUzeAqIIfXCAeNgdmKjzLCHg7
k9qPMUcF0Oj2MI7xZLN3IBa5QD70C4RYsJyMi1AqfAht3gsenCwCqmpgm2h89sq7u39L0pq8Eq6V
Uxdskhj13XTBVrOgBjhDnnX+qaTyeIIFZH2bGEsezMuNjMLRb84Ybi0dxG44Og/qLtUGIVp4swXu
50Q6Q8bNhY0TuuqFyQ//dTzWgk2OyYtwygbWbADeSg4NTvFKTy0XLZjLBCp/6aCdylOW88udoU/r
+bZUy/Jvq1EaKh5TFnsM+PPZr7ng6IL/g7ijqtkCHCJZcuGIfddP8HDvs15xr6ccVcgUOzcK/nMd
EQl2fZNFbuvQ6f+NpbdG5ygmMa6f/+hauT5cKqYIEEw6D/OqMSNtZb/uiVc6QAiGzUJ1ZOpYTJcK
dnqqRAaGTqbggXE+ZDrRJ3eJumdnIooxP8gy9rqmio8LM6hV6/xKlJBGTP04yE+Uj7fxma2KVLE0
AcjSVTGbX6Cb3h6+IaOD+4QJKtbPUSlXXy5BM5PvIh9W5Jjut5H2Bp7JWq2LpfKRae9NmqF+AGBw
0vdOALmeqRMWrpsCP2XICPwGNBqdM12JKpVe1yAIoZn3estb6k3JTjT6Om+OhIH/n1nzUSJLopPv
fBCodHedLN5j6dfCc2eWkXs4XbG73do07+R3ctY8c/UHXpVtj6wncBlALfV+s0dCd6ckxx8i4SOJ
Vk9sVKt6aSTVIHnNIJN/DmZGJghQ7NGp8RkHQz6I+PYfiNNWuMy0XYBTL3BUJEQ47wOM6Z/dCrW0
o3UyLf8+3Vl5OF+qGA/BNlpQTREry0HNZ3ZPztkzyyy07IUd0hdBZX2nF4Z1KKEn84wyY4K7Sgtf
o2jWBGQ7ZGbdCdF9DU6EkCUIGsy2Cx7BWHy71vQKBML/vry7sYVMvVkB4Nwhzry919iZaqmCMjSd
GciAKALmELCAbM2dqcReFhNxdpSz7vpB878OBK1JaHFwVRhaIxywNxClziW3WhyzdFpyTE1OkHBu
vLlf2yW1yIuawqk8Z7Pbkp7kRzfzUU0S2xf1X8x9DKsI+NeJ0daCg4KuqsOjFQpkx7hA3jlvQEEm
Jl4Z/sK1eHep3vJLvoW1+gAadl/lifPH8AYYppcGdV7POvETT6fQRG6KORdvXN7y8/Y1QdtHqvbl
PR37EFuoBulGHgOD1e2R/Qdr3RNnbGEJGmkgKDSB/H68VNGLLHeJqVsjdK6AN8Mbndw/YBt5fyf+
nG8HUlQsUrliOBMD2H+cExzoHIryIekjFq2Z+bEEjX/xfkMArorAsxFo9zgyxcEtYdWGo2IO4ZRF
YW0HxXAj04/hMxljgVuJjsjdFdu6Xh+ETSYs4DrBU1AdwEb7G1pkN2dboGm3i1LzSqwO9pR5P84V
4pNL116skTCFYzTLt1tEOJWqYKjrxr+5UO+yZ4wgNkxKDQGa66jOuVeljofavxq0SBgwgMcpHhgz
ZS/U5USLUt6wk7EkSUXjbyn9d3hhWrWOi+OI7jv3dLBff634BOQVOEkKfXTYCCoZ61q8qwXKBRBI
fOFoUJMNUVFP7fbj2VNYLJ4sFGiEJAOm9J9xA0mdZceAsuztVU8ly3+aUTTncfJrNA+7y/w4klG0
dXb6go/lOx8NYufopJAlP/SZSMo1mDNS+6jvgJBRcWqBte2Sdo7NuQG4rGtBYc9bkKIslrwYYvPA
R/hmtdajZXGxqOe+3ZoV32cbFl4SiAQINCXKjSYj+YFBSU2vPEcOuMM7XO4+qFziN/FeJl2BsCa8
UwKTdmCF6sYCJOEp5xu9Oej6SoEpxtV7HVZXk4RWADe2HRjr6Y1UO7Uk3astKAtflbd6Zzn/OSud
Uyog5jtKKj8dzG5l+Zo+qbbPueQ1c0gRX8KNFj0YOOv04UQ/9eobbHQUEkFeGFc2VLdUWR83SUm6
vWkqMSYxTkatQVMp4/b4D3FxfJ5/ij+XOfRFQsl1gFiVDkPGC4Z7z8RJYy43HZgqCpW2ySQUOh9f
vFSUqBijNZleQPxdNDUR/yE7JFYrIBM8zJsWAC0M0Qgugv5ngLNQNI9kuYhcnO/L4LfttVovFw5z
0V1sw9/xzXFSBJXAGUOJNG+zDrGigVIDmjyoa8RPgCP53UEwfWAUf1tcUpCqqYf0rTrSf0wroIhM
p2s/6HQabWAg5hIFyqj/WgwRyK5tDqkMh8BaZAmTpWuE83vb3y0N8zYm+mwczv57UFbMSXxnhz+Y
aWzHD0GwT0kv3h3WgE3JeRvox2+d6zElbDVcSG18RM79QHtoMiU6v3KYqz4Di9PI2Ska7LEcBytE
TBgSXjuVsVrosPop7XBN9ovVlZUeJM7D2pbunxrzsqwK9ylfxXvjbx/tO0H6mSGprvBaeBguLLOH
3iAw6ju0yvlsh+pMOqFrvjiF0B5gYHvKcE127guS/M90FjbKh5d1mOuS4V0e+qN/rlWj3gjE6NxV
KnwvyNOqqS1UKB/vBDpfCM6KlCfyNv4igrwqc3/8z870uUUyblplXyfDBSyQ67yBcN32+8FiJR27
7b9uES27q0zmLSf8shOrSFh8C+Piz0EpEH4pnUV2UJMoVNy8Cr1xCfMUCREFeY5BONzrtqUAybEH
vIULzVnpjuXoFD5Xz40zJVoV6pHZyBe+vvQzlVuXszWXEeNleg1Bd0FkBUoUdlzRgxwyqEnv7KW3
O7N+sIGDEte2jmz4sbFE5WSk6aKeiqmkMSRSUNYjqnvWUiOpTXICVKd/+bWylQna9K27dNA/jMln
t4Du4SIHMeXzg644/WsNCX3oOGnBa6WlYlPHew+X8HotOLHvavf9QZgg+w4w08udWxBd0Ju4Ehc6
7DFONbxRSL2AMtybh/RN3K6UTrKLGbWnPdR8EraGnJdHwl0zvsRubwE1xkGNXqAcFBKnu2rFha1O
MOP++a+17COSlmIL17CjBfvScK4qbr72sb5rJp/i/IVNTy1+RgXNurbAur8jLypMMk8rg8LbRVvi
apaMR0PTDEq0y/lV65hdLoYNOAY1aJ53v93k2+DQ1daFOZ13YhrnFL37Qv4emDF+P2KF/B22uBxo
h7Y0enrNWBiGpM3MxiwOlDXgDfx8EKKvryHzWTp66g7XLMSB09PO3JAejt234uUKf0JxGptXA7BM
w0H5i5jpKi6uF5uUo0LEynb6nD0JZYtgEJRRy4zIXEyL0GmD76s8u/wnjXxEN2Hu6TSOI3VEoVOV
6FdObcXrUxOjjbpw5KYvbotwd+Fc/a9E93ECg7uuJBsGbV0L0CwQ4v9Q2jbCz1fjNgPCv0oSJaLY
hjlgtlrFswl/LpYponttmYuUaUnmzVythu/mIkwVud3pc6NVJuLWJ3VnThJ1b4pYmEpVADCmbI6d
EpH3Ph4PS5iK3UleJV3N5EyrEdZyEqvoFZkPRTCZjxDTSUdC62jBWFEvQ+Ptz6K0zMSh3RWgrEBa
ftZ6u0Ve5gyodqBit0S4Gd4tRLGkzUeD9vnCYctjFud5PbBFspim6mOSoJDGdA2OZqZfkqECU4ww
BQDcQ8u3MFxBvJDvk4Lv0jMS2ofPnrzLiAmdTJv3Kis6gGGCe++bu+8Tznqnp53AeZoSj3Ngkx5n
4Pl0yXDuNwBXCCGo01LPUqZY6651033Xh7DtB2cx/wU+a16o7XbSDHXILhhZm1bEZhdmPxG4/geu
wSiQm3wHpF5kVGC/6JzL5zEEf5GVeCbPlJTXTCJuvO57BYsga3GBGyqn/tuaI37JBuyVoIX4dOC8
YI9NgTgYU/TGfUsRXhEWuvDGAWKQZGJUyXOJA0FMyVneeaNL78XIasrLvN7UCrknV+dVxIAvtvdI
vzgPKsQKe5qwhW1CHN44rFEwrHwDgJwJfeSgP4cL9zVnUk03OTmlV0FqoQW8u16YMYXVWYiv3rvI
qWk1aNyEFbOD/c2Ob108E1TiUNwemzGsGxepoJY9H8xXFuqooC2mmYaU1ujDiLZ/S2xbCD3QO1Lw
1FuxyIAilkIKxEOT3YWYTT/ftNe42CEXmGZFm/bO3cxx+xJQ2khXCfNPvYe3Ac9RIkbqZmYrnXeN
+TZZsaUvp9V1mNJzKmZv7eZQq9aT47dpl2BOPzzh2+g2zjLqLQJTtx/U2uNk4TknXeuqO9+tkzI8
3LJjc/SHsugo9daid3m6tLzxTmxMEAr5CceV+ivIfhAt2uGawUT99G+NCenM640KG0t551jzdiP9
CBqMas+AWUUXd0BnQi2+GlHUU7smm4EMfU3dd+2QD9MTvOsG9/2IzH8qP059B6MJVscELt6izNFQ
79CLPPOpFDltH/i84tL67vWUqFmS/bSXMhCGubKrjzlm0TUes7fw6fGKTqmC+r9sKXyZhDDFZ0FR
3jCX5eNruf+dwzMf1d7igfNyX44tdEyx2nUZyKSvMQiPGM8L48dEe1lp77M9u+vQu9IUAuQpSDnQ
29l4Xp4lEUuCn5XB9PpzALS5jeQvL+LAoxWRBBNYDI1ob1wA3ZD0yFvwXACXG/v7sLmdhCMDLoNg
DAgoXxTX7fFz6vZwcaW4nuDWA+Gqmkv4cHhMvNrprQkjmWX8lRcU877feaIrYc2hgYHgafSVIqxV
Fh4vpVvpJkEaGXvTf6aOeZRDzu0HJtr0QhdDz6ZRDruPFZusvgZEmV7Vr7jghM86IIDUjxMhTxBD
FEzucvqmpiG/GzxiSYADmyd8V/bSFJiF7A5cLl0pvGoqJOKQlFKTdluE8OIJ7c/Usa+469UhaxLD
zcvczdB+kxKDriV1i0lnkZuW/W2rEt8/w/NtFCSu2MCyTbQWXh5NIVUp8tOu+7HqWVuorVzkzC4i
UuIoFSOK9zi2pUPLbIwpr+6bkny2EcVL4hGwl5qOck3CWHbRFc4d1ls9l5jqCkhWQsr67A9kLeRF
S4Mxqq73lTLRUSNmZ5PvHLiyH1aLW497l0jKrs2h+EEXzl1JLzTNjs84pk8VZFaixrEJ+37iN+n2
NezbsOLLgU/66t9p4VxICS4xjD5lLcdBrYApNNA+Wc6uj8L+OLzdJkJaY9Uqoz7AyMJhN2A+uOMq
xx6Bf/bbuBTB+2sBuZsLbCMEQQnLuBEWW/y9cHXy6LdwbQZw6eK7obMNhvbj9hmmIO0LN5wEY2lE
C2n6RNiCqyMQgPVrrMS3R0KHnjDpBslTgoghGAWCHuBoyB9PMj4Vz/zzd41UC2ilbq+69oZuGHRI
OL9/1vLua0yq/9Yuudnw/DpdKEMbuK93HEUhGqq93hOT1qFk8DsTU4s6E8luDOwEWUNXOF20izBe
08D5itE13i2yjhPTTg2kJPwT0NgbUqwbHH5VwYu3qBxz989wnsDDs/lN8VTgC40jQtnXb+AkhyK5
rijsNb6oBSTGgyP7wtys0RQk2NVvbnO8dWRg735GFd9wsFqrdMyMp8H92P6TQps3YBgcZgcbhH9t
oG7kcZOODG0CBz81XPHH/0lNXhNhos5+NzLCLkBsZMWfFpVScm/cAyR/BJaWtjyUpGUkT6ZSWYsk
ZQKi+eobZDUa2mU0Ae+XI1X+So/TF1aQ5Fi43ysWq9yOZ+SGKVOAKG4hRzgtDOGt9R6VmZ4bfKZd
dNPk5y5TT2MOk9XyiRe2Y/BVIF11u38EMFz+RYP5k9nd5eAHkrjRgAKe8UfCGf1CjaZLIyxZO+ks
VGuV6jN3paWATDuvtt0JezNOlJYDLXgWIzPLP3tcDhXCFyUZ5Ioy1RWKtpNiXNJjSTX/qRHEB9T+
hb7zgJiYKbTCotmhlhcqia4/qhx4Fn8ixKW+AXhcfX5l7qJzTLz1Fcr+d+/I4J3L5ljxLkrkpwAj
3YMcYN2i5VtYun4OJQFITQvgFGzmu2Aie/q8J+EL/8BzOd2rRUQJWFh4WKpVUmEfzaJfuGaNtF4V
PkAQW7Lzv0WsJ/Jx47CMPoY54wKf/FqfnoGJyEKuJldgo0k2aWLm2v1zAKwDIsngXl02e2l/065N
5ooyqKhB2fSFdrMRa52KgOWJIq6b/0Bw4X/y1R9sF/sI6hRM5yc5iSIU7ngWK2zv1+xTAGLizr+c
jkWfxNXIqcMUc5WoGhFOCYuCoReoy4SCSGMQBDy0PTpBCbpIF5/ev5nCk1fFxbsjHekF0UgycUL/
6/EuLurx6vnbScQinLaQAnIjcXr7Of+pMG7LOuUYEjgapnDDdfrXH0LA9zg2caE7eGyIfVXe7DDl
aPRysFObmoz0L7AelNjXPI+cdBKMgKm5Q2v/Yq4C8zjAzedbfR9LHaqDU16CnD7IEZeFKYdNHKgV
R3GOm5PLRhzZyWz7b9sbAgROmKrQb8aNcC8tFdj9d8so3gsdxiF9QAi+NdPxakGEHJszZeQdSEM1
JxkfJ3mO+aVvwLUWLSxy/MytYEz3Guf1UWdWgqUOPAQJTmm+3HVh1o5A51dqpIBh+mvmGCBtkg0V
+sTqQ/L9izHQ3tPyYasJBWK4RpY0KymycbzNQA1VMXGKJvHJjxT31QDwaxEtVcvqmfq2aFuUWJ8y
V043yiXk0OZXhCDphGWmFXknvPPdaLKaQyj+sGXCHYe79D06Z1NUUDpboUga0oQXqmESn0XG1A3T
iuSmmxX79/KOng4vzcuJT9jvmFxa7pTXXvfczRs9UPZUZCg84mUJ1G/1XtRJODx6HaxRLjXGSbln
y24E1u/IU3wt661gLe2w2Cqh5YuSUV/AlE03QdTfScdyXzrHslWjaHVRn07OkABFqRTLMHodcZE8
5kUKtPLjiCQRBsT46WEmUw5cBBzFUcaDgRRIY8POG22Yv3fPJw4m/IyyJjjDWb2kRaxJtBUqVFX6
8rexPGSAxyJ8J2w65eZ8Q9i0sR7Rl4M8laCZH2osFm6h9tRGtD6KzDmUFmi6NwU1ER6nThF00DvA
SROCyX51J6ecjjIf0WNztas4u0oRPWL8xGEF8x8P95t7RVqYx5upCn1j+q/K/dM8KERC9GUmZENq
gB0jRvKNle/GC5wbkZpxB4CWy4A5hKks8zoSgvF5FWIWGr6Obt0eulIhvo2iYSL0kPoh13w9QlRK
FT7qnlC7v0jhr/tzZpjDWdBVg2yC31vcfGH2Jcz9MPfWRO9NsruBGDqn/KuYJrzBoNS6kQI97ObL
lOQyX8H5IKPx/0kXr2ZjsImPBmb/HbYI85eU18BPXz3khHVKEsXu/T+g/pGkKZbcxsjvlHQXBFYv
EZS9K+NUp8S+JDxGISldFnxGX8lJ33K8br55Lz6TUD3c9dFXFFLjzI429e4q+dQ0HeJN7UxSkNYT
dphJrur2vaqaIyPzm/g5wCJxDSo2rBBqr+jR1TiGXtfzXUV6MZCC1yKjrKA+duMM9Ym1g/k/K28m
ZX3U7f84/0t3gJCZ0hj3ssvn+avqpZQpy8DXVW3DQUOQwhR6UkGQFbiv52o9NXyY9a6eGis5rsoK
INLAlLeYGzZzadXcQuPo/cIMJeSJ/0iTLV8GD7ukkuFEn221+hIBih6rvM6q/g6G2L0NYbFijedF
q7EnvLa2ybzNGbDoiNHGbPTYaDXQCR5upnmGgnntLMhiN5VTr/fQyLcCw97rGPv8M9Elj6q9kigz
3kjDhYkBFsfCyJfue3mFLKma0bd9RPUXG9MyxVbbv2m6MVd4yC/goysMdXwYnVU9FZq5EM0aR+KW
GZfhcelNkGbPn/7wK+1RRQfDvva7z7sYeNqxrk9bsUSbHig/i7FYI9cGTNyDB5gbfYCKIHSbvXiw
qcQLhXkY6O+OLcWEWLzon1/f8A62zmVGfq9qPaNl6h+9/L5o2YNe7nFUVrgpqD2IEkZQYyadQlcg
fXx/4lnaTJ5345cigd13LPZV3Iu7/B0wJPzOnziE7yOAPerJtqIi5tnFvA1hkkmELvBEBVatLctU
v6pjSV1lOIozZiriefW3mQREFzKyjwybrlXgUtl/Kr4Fyg6mJmE0EDewALoGWpg0ljOniWLq68t5
jzY/FlhnaupxvCQe0Cf+C+CACanfWnEVPmGjgDnPGwlfVdtSelWXFPMyzxSqvuid6h5VRlh0mvxs
67nkpBw3UzT6Hk8WXgFRkMf7zy9W9g5bVKJDaaMkX7ENWT8bWNLGRzBpS8bXnShTaibYWfhT3Ny3
XbB0NH+cvX0V3KHIlZK/RxTYQdokMRtmnjc9mCQ9AVYEuKOIWz6i4Y2UHgzasFDmuP/LDLODulwj
dhNAL5nzsBRtvTcTTTv83noqws3GSlSL2X8f5ehKQ4Oyea0vF17adD5Bb7YJQ7LvBQurUjcYo5am
7/PQTxJVc1Sk5yj8K4DQ7J4FL5YkmvBsV7/oA0lCbsPivENi3rIfarI7XXydSIPbpug6jSJsZkHQ
2YzNVuy/Z2bEatWRyymAcPDldBotDS/CFhMk1P322hzFoQwi4dSD0amGU/4pUmX0kr2NLMqZmrUq
0i+dUrPFvGnl2s7gB0pNPA27MJ0cBEVSWWHWySsZ+SkqDBH61Vm6xN99hebey0csoi5TI81F6F2m
s/6wBx36SKZOVsQSci3YJu2GTFqeW3C9sJbi7h0VSaJCfZe9rS6dVgKCPi9ZrIep4rHMxR+q6OYk
iMWl2o9PMjiLdSn1uLBmtud+2r5YM72pKcRV7kX3/ax7kC5J8maRbozSd1GJqtBRgXW7tiJydcyN
Y+aEe3/1R6gLQEc21yqsQpnXpHGWV/R5qAm+fjiH9eyxVLccgqI9/7I9bSK4nrOUD2N8LOjJzi0k
ZUFH4cS4i8mLK26mt/ERdR1L6KWGOmYu/OEH+fhj04ZIPihtLV9C5GfQaJYCjkeuEoEOJGR5QluH
kvIZ+dGBqh7f7JRXR1vQ8M1iHWl3L0FJRua709ASQ2ZxJ3MipHPPjAXBIzFXh98VZzVBjvyAknhl
Du1b+XYo12TVCPwN9hkAWoz8KsDsZSgNUrSgsclRZrEZ/rWAlg1PaHybzswqPsyO6wEOIQPh/xmT
oSCupO6ih1bm4/Jco1IXzh/7flTPfs2sWtu805HhZ/AwM655gyUaGCHyGRVmNYIizbMBhdHrPjbj
9otzDhxqolZl5duJ2mUWXw/eSSLwNRwHqq9UZQjx6dd0K3VPVZIn5rYcQkzPJrOWa8lbunP8SZU9
xLfL1fPK9Qc2zJbLtM+2tE8+fRQoCKPOYpzr4F/rXY6e3qlXoOcq3zbTv4u1Ah7QWnbdqUAvaGqJ
8WAbiUtpebO4+78SsbFt/mxQPayKXrk/AsSz+HhbGNaSfaqJUmcHLraHjLDqWOLh+4KW0pm9x3L1
thulfH1BTmPqFfHRzoRNWaBK71XgmofCKUXhnVNV1pGgj7+MZEysAKp66c2VeWILkZ0abTsfvBtZ
J+cqLjzwdIvfx/Psiiovk8czGuMoyJEbfTtiFE56G8iLGRwVhGyv7pwo97RdziFEVLo18V941V9G
TR6mdNJiTk5sA07SlARyA7JOZKPPfMnwUld7wgf0aMs2vS+y0NzIUyBoVeE56xSoavdoywxZczvg
6qqbt6R6BQ4U7xA6TbHRjOqUZn8q2qxlWVGsZ0z7pBVgq8jPVgbsdKyzfa9CWlYjhbp1LJXniYxt
ToOGmNSz2UNSKDMHWgB7003LTCmEvKhMNgx23SpCSjXkVY9BEGWMFZooMsazp1q2ZXWMJTITTKjy
kdbh7hYkj1qo6DHetRSvLxL77DCkYq5SwxH2tPULiCxsFQlNtHsZIMTWUjn74J7mo/2EUOwsG5Xu
4hh0xgVYOPrSLEgEBKfjM81yqZ5JZMsShjr4EPi6y2N3uYT11jf2/iB4veYfWTQjCwS/ZOBw+xUQ
e4MJX13p2WSyMPgxTI65U6+fENNCFchuPbNYX7AAD8Hw6ULNwA2lpMm5q+4tKcp8EcrXiBORGpeF
UBESrrz6K4uMUjP0WVPH165a2ZyV++sBYIWxOP8snes/UEiukDRUjZFffnaqyh97OlsL0ykGmddJ
PlE1Ffz7eJPJsCjVE3rDYjd5r3eghbV2VqWzgZny1dfQJObgtdOvxv3Dpmwyhv1YTCGZ8G7wlsiC
MizsAwhssYHAWY6qUPzonRp0ySgxwaBONSN0Wgv4pRs+r9HGaRbSOUPFaexMeyq/IaKW8AJCzQKo
GqYMHb5DhU3guZMjrFKjgzzyTfDBl1B/3qr6o1rjzirnr8r0Z3R9NB7OQLmu6B5tBML0JQSgxfsH
ElGdYBhiGfwp/6bU02uybUJcBiWJ46HhVJGTf2W7qsKBQdwzMx5UUfLUpz12tqpv4e7Rt/QL9xvB
/lBD+9n8GPpcICm3CY70UkCI2gC0rmpmbFnHTR8kuSQBZFj49Ow1Aq5f270wy0b/iOcENzCoHQQ0
rGZ2RLqvONPwp4XSH20j2ONAD2c/8LB+/WHx2CdFXSMXFTeDp7VLFeQxIZv+AdBMaCF6uSS8lYJN
1InD7ttRdlQ4VlxhaOW8vjtLmhgbWTQFHI+j4w0C46pY1shhDgjcFUtCgrew/WsSgdto4xpfs9OV
W+csjCoSt+gFOZ06abc9am0cPdg2BBTB7O8XzmhdJRPC9nuSySFtpYHLCoAjZB8o91XaYgRehHZQ
NvqleUfIt2JDGyNqe2/zKee7Ft2jAZ/NxO0TMfugkeBzRUrlmF/rnoQkRP4EvBxkbkseyTIofbQN
meJNj9fva9PLpr/PjvwX1HeQayue2neCI5FCNwV85yWPQtcdvHbTkVc/7zgoq4OXlY8JHtfjbzlh
gUVsGOZL04KegcBG+JO5xjWoYKMCtZPOKQhcs5axgkyStJa6425iWIeabSNBqg5T3L/J4pEf+1WN
C/k3bDFn8espah973HFLppFEp/SDxnFl4H5cSyYYiLqm8ryDkYavSvEjjl9jeoLAqoGmaeksM0hU
KdSc432/ay5RzGpR8VPhCr902a7C1ECCXzusVHKnnCLvs6Rsq2XbMcH8B/24VHUuEXtDdBgFcTK9
4iionoc62iy9VfjFAyJGgQnnmPl2D8NJMgR7IKhhsJv7LIQxFhstzCN2Cje8bC54ZDgyxb06FFS2
tjKW6HKSntkgGUy4Qenx0hdczWJcQBRgJfcminZKxGfJTRrCaaHcLnFcZmlnd21IjZnG9L70Hel5
X5LuJ0yq0uwj2ei4zrHpdEo668EczJcECPloIp45OQiFLVPKmI8m5rE+Yr9+ODHWkAC9GIZI8crS
/Tkv0Amc0QS39Z7UmGTyYFWmfrXML8YVj/5QLDM8Hi6AOYfxc5XXDiLvEbYukSFy/z+GYnDyGLh5
lPgcN5aD9jhtCCYI3b+idwEkSNeVn9WJyP9OFkUgZY2IaI8P69KTn8bmb0sHyzlP99YqXferdyD7
/f93GRWt8wLc3PsI6odd/QN/lBEHg5zSFTDv9f9Kge9Mdw4tgJf05P7dOrhqO8UUCRKlJZaP5Hkb
qt3xZodIGga7ryOiJRdXuigsW6xsYwWV2I7wxlGgKzJW11Cr/BLmwj62WBeWujWQJvNQrcEpO//9
A4LFtX7ApyBeuQqc2+YbLCq9z0KxgCiUT/8wS+CFaNfmzj8svmxSkxSdNM8H3O3qlCBef7Zev4O3
DkFkhk9wRgls1ghwg4zEEoKgrIE2KkrQS0yPZ7AqHfRvhkY0qPrFCDFrLP95kd4yGTsEhRFigs40
V/FL1CGoJFQXeIsMG4bUezaBb3uYxhuCsb+qX+yZ6MsC93G3z0C9EJsCoLJA9MBK+dzfX20NyCZf
WfNet1Xsq47sj5slGIc97tuU1jPYw3uPuLamrCNK75li08OEZndXbVEp5qIQ95UNn4a8xUsiWOlZ
toKml4eCj0f8JH9EJjDW/ZFGOsySchO2nwqmtaHjboy3LPRUWto2NUZ5ccknBDHUzvzVK1PtoJUQ
rfvomcjsrhc9lB4Id8Zjt8gihuaNp8I9fkUgcQLBWRNzx1lyThvD9Dq/waqJrk7HhZZ7W0VnW4m5
TxsIEGfEURc0zH2qaE7YulDDrETOdtomqirdO1pngkJAA3MdEuX5PebnkkBtE/TwelzZnxgznD1F
lRUyNRsMBrYi/0tL4r7tC2TTpffgDG/Oi3W7usMnEUA9tkn8JqMQP5STjXccyPGHnH/iDjMad19J
HS9cfF+qHFRGUG3GObHrS6EQus5yFqwEsj8aZrGJLGSP5a5SXxTUXylOwaLTeedrrFArv1zqN09p
WBdhUqVVkbfxJHVTn0cZgNXoWbrpg2K3/iArrjY4qvDldtPENW+7/dw6iX806Y1jGzy/GXXIVMdG
bKs/zzW+isTEqbEbYsygVpTXEaPTyvZ/K/As57tcF6B50l5XRzqfxA7jsx0lLwnVko7xV5UuEODG
85IpfbERoN64JWsx8Zot2iqTSWBCUiOEcZ7p+ZcfSUKcPQB6GpYc9rlyqtx9S5naUr/w6kJOv+su
xf9AU14y+uS3WrWpaRfuh09ofGfq3R976qpdPDbUazj7DpfagM0WPct1TGuK1uXOlgwRksUeqaQT
UCXFZnRxcQToUhGtVUCUkeeU9HgsW4B8dMfturH2Gef7E//LYgNPZLOJmAmmSYBmG6ZPGmkirV8F
oicOgC3tbrnz6pMk03dYOe6dbBtm6UGoeabACG6E9obkcpwOhZkZ+htSWb0eEo9Qk9SKlUlywTaM
ydbh6hfOcz7Sekwi7TzQDEM6ZXWfUK2X/W/8/G56ll6HXnprN0t/jU5/Mv5y+geeluAmXVU2u2T+
7466m5dTfUXDpDcDqZVPFNrU/QCFHXhjpM0df1huNVj2kvKlyyGSoqz0ZkuwA4xrTX0Wqg7RqjTp
UR0ufvbw0jt+avb4cWdYvHD9Mzq04Rz+6ApMpxzs/7WDG3hihBXqijce6mNu2nsDJxsazgl9bC5A
GAkYxddLkMaTo6n27lQRBIgBLaFU4ZcrOnTlQzAwVG27vze1GVPRuLk/2hsPtVNrke4vthbGk8BY
UYPY8V+4ocPoZEPYxN517+aq9baFWXi863TqDb1Hhou2muCB0sxfYZWcuAIolOSjp9RGfv0IsQHA
YT6p7W5sfoSrJC/mfwCu0wgAZPVN++2E8jM8u29u3lteK+ZdaEjB9OZzQ4PwFEw4KPcDHmRkO8V6
urZeoZGgOzEO+xLiMXOTE56cxxsTaScbQH1nTLgK3X80xCcYH+YKWUDtyLaMuWCbk5PMFBLMuyCf
tiJnOp+V9tbmvpV+rbujRwTKAQw+gKvPvjcJqXUO0PJPGkKMqDbN7ZotEjqIvx0gS5BLoUTklAGv
SbP5oi4lym+NqtXcvBZy6xZbeVLUGanbjzaAXwbp2laGT6xT2cb+za8My4LWuIHO4Bs0V5Efk2Ur
GZE/73qELp1yVzaTkTgmSj+NeWUH0vxr/Vbh0+TOU1gY8TMqx4MF7Sfo4wXcZW6WXCQHHBQaJ94f
PKqQeeluN1//fWBrekIy++AKMJvRA5odaL29szMUObB8KNW3s2n8RFmw683X4h3naEEMiyemFG0V
jju/yQ6GkBTTWPy2cpVXYlez0HIZKdBHK9E3+mm4hCsFp0GJLkd5Vun//ieUDnxxAX5gvOe/6U4R
iIJjMejiBI9/xUHZmyOhAT/59tmKjxnEnOYi+Y3qUi/5gOJicl6ielOeStquXOL7E3TKSSknZHfy
8Rx4OGOfzoVU9KWz+GkCT3Qv35gHzyGOi5x2ytrgMvD65hpqe1BH12UaoUeIlD+9dLBP7qSRSKbk
C69DkHlIBHgrYZQOIuE5QbYaTS99nDw6mCMvZolkEGt+LTUBiVNnTF5+RsueQqXJ9WhR/KJ05FSG
2bR+Yec9dFrfL0m3IunxGZGYIi7ZTbqinvjTEEjPG2fsDqwyKTQv8BikKwn4Knz135CluzzjUuaT
ekCCfWRSN+A+N2fUnslaFPTkYU8jyhayEHix5DP3vzwyaCPK+X7jEJuQrPhqv42vnszRpwA1gOgs
6PdHNt8/KGJvkg1eN9WW6ZeIbn4JjL/OQh5xH4zTxQsNhEtN5SweNlnIeKBxvVwxhZ6w4AFYg4dc
ehiRqlqIWaOn6NWoh93frAJBfK5SpCO0mINzxsYpr+jyDPpaiwBqohhNT6gQwTkd7/8WbuhALyZ8
x/Swl90aPfPbiQ76BwDr2eaIZ8qciwM33GipBkjt06W+hTNAOiLlGP4qxJpZKCGnGP1cw98dinHr
ayxbzVRVo9yZvvFu9zfLKJe9J88jc/79d9DVs3Psw+E999f04rpZm8OCA2Kvfi23amaW7migqQcH
HIfuMEZyff5jb/ukdusstESJLQlQEICMvFA6nj6VIqYApxiSZpzbSxrfoC6qz6bsW3OxmE3wOZfu
qSGL1Xq8dsQyLvA8tX/0UC2nxQiHAY6okJe3lGCmtP1aQ1q2odN1RyXh/tNazF6wkekDXmw3R8nu
rEs7FzrG+k4XZCWevIBWygV6mbZ7OnMKgA7BpqDmGntWFdsbIgJhR361JmbahHnfa4fcxDUPe0bm
Oikydp128OrqGrEHokvV3rWSMdTLakWsxzKhFSYPmmwJV5oH/HCOfWDkUysIq8QoCG6ZIyazvCYW
0QI7yQ7se9MKMfq4ZSVlJWIWz3iDV7CLpKD9tjSSgAzr888z90gCvAOiA9Y1xGSuFBQ1iSm+7a/U
jiB3YQfEiCcr1N3R7BKMv40MG7lWqtJKucHO041SFmddSHzmxCtEWpoBhwHH70HWA1oQ7Jq+UQkp
x7BpvnhEBfH9eq5QhXEL3e8nCmewraIw0VzszPZxA8sePy5VfYId7G5CeNMCqreqDCmIjdV3RHii
yZqk4YlGsBvLjAKN22FBXJLQLJcDXa2DI3RU7ufBLCeEZ6v7ohhG1dnJbFy6XezTvhtGui21PEjN
mE/oMMP869C1AKMR8egrYWOky+yFLINBsJ0FTVQa/nq5VqcXsQR6h2aWykN+9wmlbBxdePzYfuM7
c+CsLLJvPM2pImVAyrtAxhXUre5jAxcusROgpprpkd0jeM8Xvm9JHApSQEjzQd9Q9VAIqQWsK0eo
fUCKqbK6dJGRDEEdh2hKw1Vohwe3+TyVYj+b6atYRaCpyMKY2+9QIkOINXeU6rjd2gAKkz9RuHhg
wf1JApYw5LFP5+CgfPjo/UAklg/Hft8LdYPyIynrMVYVi187UGdIf/AxMKbfQB08xkvqE7yYBx6N
/zk2QYmjBMgD8j1PAJTSa3/xFXNAemQjltWzDOzjyGEyYbUzwaKSKjBixuGhHET5jEZRnL+MAS3m
De6qj5g4p0OZwJF9/+4udX8vV24JpoyyRieAUWxB2Y7XZj2P9bbQUboQ2qElIDQrWtdl+uCH97vM
ZveGxo/X6EGarS43NETUCbISBpyDOFcVxLWoKSn4xbo4KgX44tWWOOFYSYHspJ++eG4DFLG8w94F
GGW36qOrgT1y0WZBDzqAoC5IZbEVT29DYFiq8APh+FzyVMS4fCrPmHRLvCmogKa7RlIJlEtnpalo
nZi86YtMGMzPEJa8D6zNqhpRlWk/BTUFlGfqtkNN5vxADjPdqKkhr+88pJRnVCMQBF2aYpIjP35Z
9MUCzVnTJ3qB2ewjhE/SDQ2s+D1HCQ7erWIJz/pUlgZBRMTb5rb3L8a5VZPVPnsPt4I1sla/qqLG
H/XurBqHT0FjW+l0U3uC7xXuYm+9XdUN4cptrYU0oTOp/Jm+sHgNSRrFxKqQWu8X1z577ykLFgSF
WGnpwdZ4LFOV1EkPY+vjraYiMV8NNORlaYaeegkb2eUIujLgdOafYf0jE3eCc0UQeqKfXZjISfD0
CEJmawfjB8oc91GRUdhFsM8sSxUGA7BQ1/nVCxdIMqD6EWzdCJIAWBEbYd8l1OgAZWHdiVcLCgv0
BS6RvcBhsrEFXWd1Oo3O4Nf8/pbgsmCxdTUO92ZYPFJLAhUKwRWdMBmyCw7xyrvGLcuTWk8Ln/N9
WX06LaNfKpVdFh9gvkqHhwqJ6zBDqbfnN/9EDfTd2jTDLvNBdth/T/qqvh665PjooasLx7nFukMJ
mvMyfTslNdtIqiGYQZ0HTqwAiK7+zYT7330Um/mHwBPQvVikFa94vIlwwfn06G9V+4I1rz4HXrda
sfs3QWoQtnD7fyWYR/nfPjFYF9sEDMUp2EreW/pFTKSARgE9cgrPVWUxn5uc1QZnFy/Q/Qc9hUsx
v6rdZ4bskXZQIsoqcg6TPBJfwfqaT0EJb3OhskWJY1mLkk/HfawlavIgaHiaN5CsYYY41fkccbny
fdr6TCc1t/Ob6n3F06ZRZ2hwuJv5h2pqgfSKv6CRLsBL6Tx7BL/0yCLqyiA2lTZT5uO9YcKrwRaF
lw+GhSKXrSpJxhQby+UvAeSSDBG2GZUsetQOhmFzl6Dz16pEKIv9APYzm2p3m/OtC45ZQFvMNdof
roj8GyrJb5wkocqMN8B76c7iL4o6cF23nW0+EXWC4h54ejgXC/73XIS9n9om8ir6IKGt+a7xSD7I
NvQOS6rq5UJGohWPzFGWvtnMTHLqEI3cjnORzXnUeUQw8FpWkUICt/uwL65c6RsXrMs/XDSPmhLp
BAxdznvUH9/Tf5yUdKbqnrMkYwk9Q3AaK+JP2DeDuizidQGlnVE8Ymgc5OYgVq48TdiEOKGE5fja
agqGRaPQr9djuUh1JeUOgJmfyeeahct9rKfYMLlvoBAIUXmPjt5va6wJGE69AvNPkTJJwVXsx+J+
KQr4yHg9yxTmDIgd3xAKO70qlfeHrOxvBzAIwH4sNd+rwCJMhr8kgdj2SBwzKBxmDw3Mdmc8na94
p4oteZALQ0ordfb55Yf99lv2cZZe8xknomvcjnpN1oAV2sbvTxfTQWw8vyZwH5LwZifKZLsY04KG
8aOrD8IImn9VAp1S+mSDMX+4Ap+kYqi2COGSlfykgjXhxafmR4S8zXjbIKFKNv/XtYOaSCdar3KH
cjyM1RfUxWQoOzg8GgZQkVwzgVRfvpuYFiKFVugzKwu10LQbQLs87H9+pH022JbMptpGWIq4RUmG
d1bfcI9s5hAs7E3IRTvwkMBEhXQ7sLp6HkJN0gsCc2sgXMJwS1k5myQd88QMGaFIxwbB8Xhk0oEy
qub6CgUYc4Mn7dB/pFJYdvpfD5KpNchDxSkpQT5GCQcAWzBp2K3vGXMTU4zq3syuty9KHZcPYOVu
YYt5r6SYX/ogeyyJ5hol8a6og9mSx1nEa90uqQaI6pZFd36hIAEnaCqQeaB8+jlLZobSL5Do+vE0
So9IGKpu5cOARkjGuf8LGEfibriaOtudmnfwVjg6CZM2B6yL/Pt412v/CaQwtD021TxMn3QDj46o
TzRgNYgoTwAPDwdrihu7oQnWKVsx5kd9CNx/L40oemOuem1IWqbwXZT6WB5C7so2oBFDJnIMMFSk
9zJyKTQfnT8cpRy1a4fMpXxB1Cn8Ec92hqXJMVkakw0B8o9Z6S8ftpcpgssVDnu2WpbLfOENUfEK
/PkGZPj2XYj1XOGgftUL0GPRsb7ovkI6Qkmo66cyU7HIXjcyuMiyWZi7OWebWonyau4Jsw0kUUrX
bt/78UUCy3oxZK/20RW0jC4Ztk6tmaPoqnAhdC8i+S0EBExre7DO7aN75Uzgp0SwKNC2yDEiDLMc
XpSQH+49KNd/Li7IFTdsTY81MzEEcHiiV3ZVI7LHoWWYsRxdEYL7ToOHbW8S9n59epVF722LuJoG
oAu0irVACzbN15Q3AQ+b1X6EZVDogpLaIJLRvztYp5BuS7K6bYleemDEAJJmwpR7SPQJzUJjjb8O
IHmFx7kyJT21NPAkrtHzwxJiDhveNulLAA2Pluoye1mUSqj99d4raGhFLwBjnKFRcpw9hxZxvhI7
4I8VEJzeKHSjWYyjyw3CZCEYV3+2JAFWwEIqpmSckoOCl+75axXXjMXcHnXlcQbuFJB8TVKNzaYr
NVRFo/+Fi/athNCg/DnZ6FiiQM4QuNwfp0cLIzdZavuxhMPvEw3zhL1AODw6jCwgXFKwa7ZLOHul
j8nA3SsNkQC46LOrFdm1nOl1ELk2fTkiMhCU7uKmMcj/E9x5MN4LzyhKmIjQy+BkKfZX2TCCwFXr
hRNNEQFXfJaEx2H0l+xO7GqAzB7OdF/s8TtI5tJLgSuKDnx5XEl4ArdcoX5UlgwJAhmFulCfPZb5
N++nXhHSh26cWGVi1dcVZtf7xPqX9b0qLXfadAbhsDLX2eotF5sibi3rqCXLv9nuTk8J7z+xqbKe
EM+tRjpISnMOoh/xMxAUB+K8ESocFA3kkKOMh8yJN8QUDsAUUa9BwFIoUAnIYep0gx01bYtI08FZ
K4vrQWE6NA7tsXP+OBLR/YB68pQSygWIwhsR4pHRjS8Me8gQFx4rmHbTWMyl3DV9eu1iHm0HjEH8
ZmI9qaZTXfdGDRpdajgtrU3/psE4Z5Q+EAZFW/oaW5pGzVk76wsiYRaA8OIsmtPpHGwVOUxjBDJ+
yflOWCG5lsen8Vykva07Oj9Yt5j7lB4HSGqoUv8ktcmgTXboDMLms0Y7SWNrGUdOUvWi+3ACq14b
HUKHXcAS7LUv/DXCW5BDKiKC0019mPcWeUbDQ1fAjm05WX5H9NgQOHd5R2VU1tazmLlkyMtYcoOe
BolAlN17/e6T8NCFA/pQlfmK8hzvjt/HVUAigzuJbo6AOV1RGUwg8LVbUjVX8f6+fRTXv+HDH8n7
HCBAmp8ZZhcU+4DPFzJtiPnoVzCy4OijU9RKSU5dYlt33ezviyCvzBbreRKVodXX6fnohFBY71ai
3GmWpAwWQtcLTKCd/HAX2KVZtdaxSPNT1lX+tTxxs4ZBtt3qAWzVwfU+O9aal5R9WQQgXEqkQV6C
Ot1l0AMTKTMqMdWC+gKY5ZLOwjPURsbN5P3p9l8mEVJ+RUNXqfmWeCVWI9kcYrtOz3oQvYh4Xmn6
/JF65r/2sxqYec1+vdHxPAuuTgG03Mla5jB7/DQqXTygbW8EXz1EQlmhpj4RfJmfZjJQgBrYwFoO
qK9+BQjhSgujNsjpA3jV2lU/0Jbea6DSHUrdI886yOGl6B/kI6ngsg45u7g5lhmwlK25sqsO/5rp
9BouyiZ7kemHv5FDH2ZZYto9pSDmxg2v+IFagSHV/IhsH6Ms7uCD+7T1U1Cvm9kI95Fa83YCJEln
3ASUufT10dIoIUxfEQ8EGFE9n2mBpy0aWuqhog8AYMfed0n8Tg1FUp1NddiL9/wQ6h8uRsNMpHeQ
WW+64sg+JxDlDA4kfrwjNfmZiMrtv/nece5Sch79bmkQ02TWYEk/f+vuUCtysseiTIvjPYTYGzoK
urLIi8W0NOcFlOA8nPhKSq50IxxRPgPaBzgBg193tW8/3wqlS6TU2ghdLAl2Li/IRA8lJXZDmI1g
IdpvsHUyvzObGUHZpw7KGe8NtUkFgHzQQG0DCVzux9KNiDsdUe03EKyGFcDpHe38klivoy2TQanY
KBe4gTN+1T9c6M4rRdOKCE0z/UARhcj8VfQFQG9d7rzcpfMSYGbBIc86x/wdegWlhdWnKK5RARdk
F/BFqUK9Ghr8dBkL1W/SqQXCArlAOnrKeRqYSIs6M/geR8mlOgf6vubKZbdKYQ3TtcjR8U7e7uNS
z0zZEt2561ofUJdUIodjJaeA2hKaBqttzk132V+DbeDWGgKb9A/SN/5RLMAZ1yn93VCZu8rjSsIE
HbhXApXO+FwE51XOSrNmooUI0PkWEKA68+6+pYGhg4bNoMCFEAK2JbRD/wRp0i4VtZFzNVl6tU6O
Twz3udM4gCA6TWuTcuQ+s1VcGQtr4jDVETqFVtKX902edVVMYC9jtRQSNEM6BukJ81XrN5ViLMt8
tjeMJRSTsuRIsV9ln1DnH5/XKdlpNFwZi0fSqzE1R6ZTWBJYDbJNGVDAH+1yHHlLaeC9UDM9BGoL
GGfivmlIHtLLDUtyfeW2vqXPXB+wDvaxGPfqFMvugMPl/K82xszX8r5FBMl8EylhAyz+F/w1L5YQ
L7SR0pcr2Eqmugu/PlORrQrJN7pwqSMWLUNqfQPy30lYjiPYvVX1IWaTxLxxrwt7VOxxzK0R9nDP
Pg5hKbqhqzjDwPdQxHXvkyDJNJE+snScA/BCyTqOiWus+aibXVo6P17rnZv9o6rmqXoSfFeCSuZ5
Kok/cTfLAN7gdhPvGSqsxKq2Nh6kz1KT3Vjj2V0QN8XGE1ThaXcEGHM+LwZCqpNkyJ6jrBamJwRn
FhpTUZ814pVOIf5N+jTBie9FVj+SggQHNRYbqhC18Mos84fA73MMDJZ0fvMgggVsssujOWSA895a
59ciU1KWe1fd3niftoH3i8ICJruBJk4L8ecFMMvCeHoL3d3Khl7Yuv80pkk2k/gqUqHy+KnpNwG0
2h17CDRLq9dNXFkIm2NdGIySLbgn4Ds0T96QmQhcaKKpG0m6lgrE5mRBCxCGNLR9csCJoSnYBf2b
wgu9LwCRJf6cqeCR37ldGxpsk7XPEjlJgavwHNG+2XBW8YkgOkoTt9nDfmmgPLlGEJlaugaOVpNF
zxMqjyInJJ7B/Yyw0z/YhdfKOiRdKknOAGQUQZ5nFG6+7+XHSdTMkpRP4MkjGwzhD8ydjictppuu
BxmTqlWzdmN2QxLX3rql41cEX9GQ+r2lGCgqdxW2hMgIeeQ8r0WdDo3wN5nXsS9VmIjk7w8K3Y7t
0EOLx3HwZmv9V1rxpEPFyRYUcqxe3bPerCuC5BCvFt1EV+CJoUJk9pFOYKv1bQrFxN5zmnlxh9Uc
B3gGcdMYUiReASR8iGuw8A2/nRbUC0vHo0bq4MFmyHk+DFIpTlpcqFeXJUoowurg2Wwzjxbaj+m9
xV/jeK4PB0Ev/eMdOsT694UaVv1OcEYtylWhoZmUPvj3R7LIxrFDJYV4SuIp5U2QXb5Esqxzw21v
OEyWrQLJHWsWdu8HFJGy238T3VDJkEBQUIx4eo6c/WkCpGsxEn3EqUoN+YP/l11RPzrwx1Ryp4oD
huv4r92WOz80DtEO9qzcSuY4pxpDNPoTyCDvtDM+F0KaY+jMjtRLZInGXYo6/fBfaWc5miwoKQsj
2FQJIlulwC659tq3ehqgrKKp1CG4S7QGCE6Ht1kqdMo3G5NzmnXhXdNVyyvoITBWCsMRnr7OikUl
jD/2jl20KEeGOGJ4ae/URc4qUniLIptQGoEA0mCjQahj9NHmOL/MIjqieoOj+XTq6zUv4KrJ6A0r
QZrA4UGzDSfRi3UkJywhIuXgW6GmbPf6uq3apLNlBz/sPBWbudTKfi3XUI1MFdNgVwEIlFhCSv5s
qPDDxUgcpSbRp+KLZAK3mKusm1smusLIZ4taH3V6mwsoPhN8y0CHyyZwEoCC+2a/HqNA6EcEnoTZ
Noz95RKX9Es+8ThQPKJF23RbPH5Fw4xCUtVnf1J/L2fssIKLq+evTinKjK9fsPsZ8hlpjPoUCjFT
gMejfFTIj3861exD2nOvTZCayesieSx9ki8xE213feXHBpNTytVcmFwl80HrxGRAoM0KoqbiXqcQ
4a8trXyq2pWGY/43Sbtv709RQYjQj0HKRGD7f58MqJy3uWZeKuWyBfZbOr+Gh/aicrt87ByF73Te
1URUWuSn1H3a+sHz2ifjBcLeCMxUGlJU75aSn1CWznaKegektIPnbGedudli56xGbhg7A2TKn9kc
P9AKLYbdNFsZAJqb+gBqiiJiX1MyS4gzoaC4QG3DFVNkuGfkFAF3pIs77JeYudj9cLFqXohZn6uH
ZS5kLXpGBP2wAZJOIWQ8nA1spbCfPR9D7/fZalpUJwuNFVhRFcm6EqrIA1ax/Vk2gyWd3rlEs85O
TpdjC3/ylAUs+celRnPEX/ixovF/tKkHYZnoeYcWwRs9OvVnyYeE7pISSuUvYp04YEAGBxvfKBql
BHEmuHAJRBxjIRkQOmSlWOWIHwJ3SBLMoOCYra62JjJUprWzPo3eBZuNPL4iffZnv1ZgH5U9Q8Oj
vzAc2jRt/S7J+pFe9VJUfBUd07KfRcy9e8K0WhuVYnIkxQrMAaEcEoQ4HxzH9X8EnNZl0KPVnlAP
lSjfdh4SuWFCA+6nHPd0dHsRJLs58Rol3FEj2COL/9Q9rkTv0T7bPBK5qXiw6A5Hm+jytNNcOcfB
o7SL9OcAUcp/F11wpbdd8qEbZjo2IsKgfbUVWx9Myu24DQMgmVfIoNfVb09e32D4TiLcK0g+Kb7/
z4mgsRrHxOnTpb8Gt2b3viKGCeOV9TXxe2FGF2EVKKd6QHFPpaaQvLtlcHoK9weWd0UMAUrCnlLW
vxN4TX8mNvY8upToVDA9/HYogPAmA3V0T/BqWrlY60pTQWKmKS6mIMluEFhxw0SuAtchytjW7C3+
jdbE8pm7R/8+gdRMx0VU/UWZYk1RdYoP5K1BdheLNp645wQI2IirYr8339I+Ji2GSgd/P84Dg7RV
AqwYSvDgcO/SBnd48jvpe6giTP1mw7uGLq1ZVupt2yQrgfJNNUFPBjA8fcDVFqkt+LTNBb/ka5Uk
HAVNIDswRlx0vs2MQubWOgnaNo20JOe9tqgDDYcPrOYcc8b4kT0pnkSFl7+jOgE7QMAX1Vw2mAYE
K5bVEprOxLpr5P2A97QFWzRe9R+c3Wmf0yWt1jCn1vPddjZnR0QvSHP8FYrdcMknHYYgP15p7kvf
aUT6dYNtaFWZekva8gX5Vfl8y+2FJQ157WU0Pg4iBLxTylVVLdP+9ZBNMNlirtabB52xRWk6K5C7
N5XEpUdyLfS64Phroj0K+FUEtunQ4f+kvgAqbbQL1xXIZmcCJB191c2p1REnRdSAOLhKbywGF35l
1fX3JkmgLyRi0k/Xdobp71J5H/TUW8eCS/iGivfw07g58CMEcxF3y+Mf9EzK//297CL/FRJmDuou
eKYDDnhelbo4WKtF3NKz3RRBj5kpv5lAx/GLmGVT4fGoOTi6xqgi0Ne60QaQfiEQ9UeAKBhCFzi+
IX99RZXHXe0+7x1fsScoWw+Wsxcw1So3+FQpCxs7p99Texh9SZdUzGhIFzsv5m/Ijv/bcNEGyLth
UP2bjmnaH8xL5XtnpL9J2/SnCrnPORq0DpZUjbwz6lNVD4oSSrZzGGCz/AFL5bo6NjgigHTePC+n
Jme+N0bYHemMRkCQ17HU6T1mWqlwq2DoaBkSUgjRGFECHgT5KST9UB+DRpir09ITqr9BFjequGit
STmxZftGwe/jcJkU7mS6Tmn9pxdd3+3FgY5EXPMxE0eKBwkeQ3nDSbsmg3DWfmEZiYwnqBUbh27Z
XAfPCyHaWvvIYv04e/0xBZ/8Ml/Z+dhTafz8VIU8tjGIRHZOHD+X8ECJ431erdI+VDYZIg+CsL6g
ac+N7yMNSW8UuF37gweR2jlzB7wjvfMiivzn5f4+NxA28Doav/s7bMZs5IXh7n1IEEugBM30ZgDC
qLhmaJw7B9YdRNsuk5ozW2a/QkX36vnUv/acW2mCTw3zRQnHZ5VbKWWe/eqEF4vZSHQx3z4zHvJW
k/B3cd58ZyuVcv3uJAnA2Wzc4VEnH+SaGvWQ9uVPWqvbWdEZo7zTOt7K+bhi6JHVzwqJ6VfCfy2Z
1wtkCudY4SG3j0JLI7SxaC6KNeUfZLQE9Mj1GU+rBQTUjuRnmIMI/TEMnLPv9m/fQVT49bm3okut
OIe6XSxx7TT44fsfbYInKp7l8rNxiGRzWcHn+mt8KlgPkO4WLCmvnSs6LQZlc8Uk+K7gYVV+Waai
h0TZU1Sj1EuanPJXUtmGcwQr9k+TPEontQcirL/A6CHatJdFCPEgb0T3mM410J3Uj8stq7r5QLTZ
ZaVkJYwVn5/ps81GZOli9UE6CuNe3eYqVHDxq6xZuVQ18cS0zoxIkl3rJ3nos/AEjsT97c7zpoiT
b4ljLVBGxlcpbrfgaSPo4jEHyleLtlnNcyPkCVAALTzpUVzFVTQM15fSJdNEbXuZaVQg3MN6HhxL
5/CdIsIQIrsM8UMwtWyBplJZTFudwuUXnU6BbZLUHL8CyG88nGfnlDs3LXsPTa8hTf6Qx2puQZjJ
/QY9SgPFt5avAotGpdVHfT9spRZGIDUOTGwIwbRXCPCMEnUZ0VJeekB2QrMz34xUjwAKrPvvGK/f
cNAj5yCCPk7CmAsuO7RU7hVoG4EFkQsDRhzKZKJsprPsIw2Zmk4qY7LwnVygKk3ceZO3L8zFqLag
QPGSeL65eqEYhzCZW4ft/Jr9GoVGbvTb3JJqhHRdCMlnBeeBAmMiHjm5P5O20fsJLz7plWc27Yz4
274RVgiwNWuwANdYZI49FU1JtrLYIx5vAsisnrmPisWZwWM7leYPXkNWFX+2Kra+tV7mCz2MswYz
qVqLFb3Gp/jYjJ+TUusrG4Rjp/ul41GyR5fCdbFv5Gpy/qXVZVW9dp1rm5n95Yo/dhGSjHx/QFfG
VaDbkBnu5t0y0NJtqZ0Xf2wqczccdcpVGiJA5RooNTE5pBBnX2T6Us3mvuHJx0a7hE8pmHZ+w5LG
Ysy6D3l0NvUt0AcndcOls8P7AvP95fe2X6W0Ay0xxq364mFbU8EKmtpnHJDCRrktut/u7Qtx40pL
WpIP0+BTAYziaeEOVptpRDu7EvoXxfwZP15ixQkXbcroYwOjH1FHxY4uLdrzv9SFEFDmeqtretqB
Cs1LqyVw/OUbSqiJEXNHB0Q9Z8tfAyMnePipIEBeBggJNpPXWqpUBfYF/MLafidh6jBvuwWFLJx3
MG0SDKm9wGu/jCHV5H2dcjOdfv+J22YGq75UveMwScQtF5zOX5e6HyBP0ogKCGivf7V7V6e0i9I0
DWhvHqOzRwJRTd3hOF3/EZPWwQbQuMtR3HwfLZYHuYLUrp3IS4r1gxiwdDGpIQG4Qbwnmz+XMGkU
PdUgn0V9xubgczwDvhwW5ZXv8hIgdXFAaAikxaJJI3K25QdAeYk/FW20A5kPCzoP/xLfGg/aH+Wh
AKojSxgTrHAq081uRUGH5T6411bCDzasZC8qnjyVi7XS844c+WRxkNxoTDXLATf9mOPVLKNFc07E
b5PRwuQYX78XQEgNoo4cRkMZsjDFLXlJl4xKdpt1NqsMUAF08T/2Frje5hi+XdG2c1W23YD1L0YE
ZUPgy5saYylGD/hWJ2pLuRD1Ei0MtMIe/ejxnOmHdMyBegg8LiQHQa6rlQt/7IcWJ3A1/eUbKW5B
fVwGYc6HIp+vOFbhFsHKGyGFlQoJtOceFRQH4jaSf7ZWCUl5ULEWq7NT9dhkE2OYTCUraNSRuRR0
1uZtEYrOugnJIm1ppMNDjEffAhSlUl2uOOJ2GfHjQAq676pA9qw3ndQMouoSqSnvrBjqhl2JRJnw
5IKelqP0PHG/jPaSUmvIJu7F+4Tv17gcMIIpbS2xL33OEV8DtXJEnrW2ovskXXjofEGogjRNjnB+
cAtvetQZJqyV5AG+j7XxwvbgVnXGnx0Z3gJwRglUVO5VpFq66rOd7sbwEedW06GlCd+cfqpCcVZw
UI0vyKfDk6tBWNrX1Dy2Rb/KywHU34boa1gi4Iibz1btsdMGnhPSUsDNWIjrdxwCgis0El+1NsO/
el+7kBIRtsFXOvgnk4LjKygykA5MuA0uxerjlxRyhX4s+CioKPkZbO/X4EZw4lOFSwr66Glxm/3Q
sZLaEM1wnpNefO5O6HVm4o/Wo2VNBVNkRyhKIxaT1hNV47KXSUv/rOzlQNEJSPA24GtcSxUqxhTr
gH2zcQ4JA3mY+ZntTDchP1GBGb0It23ILJ38cMxhUNfw4EdLVtuN4ZLk8iYaE4qOtTiplxo6rQBu
Ze2BYFvDF1ukl+RTdDt+kH9qS2JiQxJGStiBYCPsulLStKYFoGP8ABc/NdtITv47yt+QdkoKjmCn
HFSCc9Gt3OkuYpXrC2Ybgq/bwFbfwSGd6H5N81W53ELjh9mCD7DUdTq5a9HabWPlaMR05iYXsqQj
sMpivSAFkjyVUfT4/5Oc2FRcWAqA7YiTYLLSVxoKXA2xahdDQ7rQqlWTKCKcwb40QIvTcItY+1nU
jXaenKqUovtTil+nH22Rd28epcJTueVz/aGlAkBhMiAc17qWJMnC3t0TODMbFEANePEXPBRGzRG8
XhSes4AdRiQsxlPmV5VC9dlB0c839ND2sGsJFsFiqJ/mV7dF5wrSJC0HOITQYRGjMPdDHXKDVSWB
bzR8uvOWQNHrxJG064oF5Hd4k/K5hd9QlBduzHF4tmVe60ymdjKZ5m0WDcTu7+6Q1iBp5+Hjh5Cu
6j6iA/zZ8FToIB53A/Oe5K0iTfnlIrRBqN32crAtBRMwZ4ahMTpPrBT3MTGYNyeDvyJCcUhUeqDX
b6WAbinTPm98CVdjusxGHYJcieJ93yi564J9g+vKQCxvxEAGRskt+D/bDMQsU68peV5Ppqhl2KF5
fjs986GWmS5f/U6a6y5hVMf90pxzJac+RfOzGcuO/PMfARu37I45GlWJg0598JUcfILs5zsoLd2t
ZqyxNJN3a8PxraKMtDVHU/TjjX+U2jgFy5DLwg09gOOzkBySK5Z2JL2mfqbYx7eRcqDAZpkosUmo
in3BtUqW0RGxyAea4Deky/XiH6/VrfPhMMK2gF2KZNMSE1gL/dUz2uf8RYCGdOVxwJpEt56Wpift
GHp2IjToc5EHs8RBD1cMyF8fH0EDIcIk/Z3U6yo7MKtQXGLZuWQ6paLYTp3FSLRwW/T8s3cHBRuU
PhJI9Kj/ef9CEjJKMFvXtD7zHSDLkiWvQK/gToB/FqRKXcZn8G3ITGpYIcg4cV0Tq9zB4FKhHnD6
yNAKd/DfMMr2V0iBrWqWmSp8qX0MHdD4VvUxkCcN/VsAS2KSi2RJPLg4hYRIPyGBfSOVtoa6nTAA
hXlEyIRaiW5c7S5+YgioA63QuNdKK9f3TOSlAtRadCkYrk4yWH00+cjii+1ZisPZdIL4hFNtJcpE
+rmwHL8WDylu3cWUd2CSTKjfekfpkzjItpy1AcUmmnNZlrxur0W6u0EQCOVrM5xVGJui8+KqScjC
TF2i/QeM+wUmWElZq0+GD351ue5PZAp7NI2R3oJU29YwqEIJK68VbwQMO8JhcHmhrBbQk7IBeP3Y
lJF9uh2ejW9rn2EJLEKD5/oIZy08JCiNnS6qaf3asSFkE0VUkmC+gKamsu79siSflLFTS+goyCuW
SNSuGQw/mkUaN4RDFsB81ABDpQCcgeb3qqLnAh53ALhXtANIaHEK7htvM/QoyejQaBl3y1ry+hjR
NqvrorAakIDooauLDe7Cs1ps6fBn+gZ7YG4G6OoJro37ZrOVuhfAiKvMajZ582zw/eIyUOyX5WgB
fVn6BWUQJUSNdvIS8AqpNnyC6gBIyUgW3sSwbIy79po6ih2A1ItD3oax1eD3Up6eBMvAFexWQBhU
TgaUriGTvfJGfvU97uIHjJTvKivry24juPLU/oWyYF3KY9UOZ72K6M+zjQSS0c5UeifzYOtSedjM
fJ3A+rH8+0hpPFKTmfThlHMM2JIF51W0Iw0z1aHqkl4E7Qz748WgoVfytsO/LomZOxaq91CH4R16
4uwljLAAJs/uB1xqOQDvD9jXC0cED/xvQjYhR/S7Sp3OCjGoCx9JxIXprcaD9GXbcJuyApPg2si1
15t/N5rHxz7TKPxl6fUy//ZAHn2tNZqjZy2XynoExaEjls+hOLSaCoqlVYTnEdTLz2X+w0+vz6Y7
cCCXrX7YXcuUlAnakq+6SfRU0GIc4uYMuHuQ1WtFtEeDCHi5qXUgBTcYXBSe4sRZHjhgVklbuhWI
QGiLjdTOYcKIesGG3Ivcq3yVgoaplZfJceP20DxL8bJMrbBJVHfNcjimUBS08CjwHqSMkKZiZNAf
mjb3uh1cpo2TQyLU3HD/zUmotdpMUDojdtlQO6Z4qkaiA7CFziXsZDPhYuB6mrdVFvBG6pOEGhwJ
i8HhzbtJp7lbrnGeVAIeZOIYDSTrfckyc52HdOqleiIKgZjsaAr6wKeKdh3eFI8qHbMRikmLMdO4
GvTx97kC+rBC8lE9rcNt/J+6lA+a52i7ZZ76Rq9lH8dKEPT34TH/nR9peg+RzMvJ4cZh5Cr8wlwG
99JPHv51YDbUH6MtogcnGH3PkJPnYg5BPDiTdAtPZunkglwBE1uUHQLX8GdMbcc58VyArj/f71sD
2R1LZnib5z7jPudHStrhhoCkR4wCv1TaSoukETFrZtxkdY+4QPVzlC6+u9kj9xXyScHWervsXnNc
PYvsX5nFNLQbqp4+L389D020pImcWk1IiOA2Vd5bReLt/DTYUimxqgMVTNS62+Nv0X4AWxHBWsZs
zGl+wtEE6UVgkJrnEV3uTrSdT9P71IBXAQw572FZR+DsgynJWxIrhzvu7+830ny6/UhizDNPOmCI
SBoBoqptmNyzfzu2NNguJgvJ/hl0C/5eLcSAGEdnMkinXIhRkPOAkjgFHMWhZAx2j9sYlNYs7E6r
JzlnfzRwbEIbx3NOVWxPEjCs3Zy9j/SkXN8GTbsPmP9qhWN8tzxHAViKoIgvE6/m5+RaE9Fa9KwV
PscC88TTf0CJCiq9ywodLwdzoWLQw4U1e/GtLNh6si9vFDDvZFF5RPnt1wvPDc+50oshOevnV3PP
OBR771sfpJ0W32S4cUcyWLWf1YsBqhjweFn3sAERuM2mnC4+xWKgW3sro2lu0rYxsx692xcgPj2F
IkcyjVuJuucRnsnDdrKGXKqFqbRqyhs9efW5GO79nSUP32mJwx8Cz58GAEa8265u4GHFYqNc2uUc
7yEpS2gfACv3d9p8XBLGyaUc+1Te+qJKwF3QRJAwWQcrKMQXdZAfpPgcQbMR9PMPEJ7QTedNsgSz
xkt5ytF6l8VZjVOogCSbETCrU0ihQmaVGt7OrNmALvn7juy8E5MjWBG/LPjOuC6sGJfpCmG+g7aj
VVGMhdcBgUQvr5UsJyQ9bXm0vxUU41t8WU2OuvcZ2Rg0WC/GeS7BFwLL+paRwGjzD/hsVkTJD/Rs
EfK8NagPObwPfqbyNm/oiR0WGkQiyStvGOsssjzz0yQTpLqmrtUo49AlViAGO4BmNmpdH+NPVcNS
wc5DvHuhH0ti2zMJrCb1tkOcZpKRt+Gz5GRFxxXAC4AopUsucmHLpN5RUmOAbA8ITY/+7nZtNqcV
Q3cSYkNefRxE3rGCQrXJbhMpwihbYaAL80XSJY1lLdHPAmrszOofDbd8d1boceVixktw/IIvWPbZ
fNIbanwwRimdRpcXjegD4GjOFoOKxLx9VutAZg52WKbCiJom5nl7HvfRALn4g9Hq9IjzBFpKvzP6
xJGgq7McWQ7PYaYjpkrq1y1s0/96PZIaG8+rJ1l+uYZZLhKedEoP8AtPAU+VqVfiLoP4YHp0CThE
d+EwnkOayN8G5dguWbNDvwIHkm5RRoWF7543OOkytRgk++tukAWzX8hfBpgLa/ZFg4OjTvifNVhv
F0NOhOpD2AULHS64UvBaCeThToqPRQfvI6798ndZQ9ucon3Y7SaOxXLmejum9NyR8n/jOr6qUucV
A+FqmAB7TLyVkoEEMwmE02GxnILUfHQ2ZtbSDvonr32JHhZe86rTa2e/sC1Wqts/li/1cS+tHIkl
u2k56/wfsyM5rjStuYY0656OWSKjAIA9EzTZ12q5F1nu5TxO3hBj5OfLbp+6mr53x+QtKBSFcRBL
4MFAkO/0j41gsHNiNPqxJ1PVJayCC1M3eC1aMwPj/WvewBQmyikaENVsR0Dh+FJoNI+WOVCBPLB5
tf8e6nPGJGGO8V9E+cy5CGilRH6OU0+MgMV0cuZBIYXXgvEA34fE7IBq4ji0HYSUGsIRFJdaVvhh
SrNYYBVl7nWHQzKBBNolTgcMTOOv5VjXluqiG+2u6O9UPSRU5S2qVEW4X6fyP+gutYJ+zMFaqsNj
IaFsZxjS/nXM8aNrih1OKlM+h8m5Jh+S2WzQco+gfbCCo8mC7hXCi7sbZlRHI79N0IWPwQ6EproD
rewtPD9UDUQo7WnQZpElb0dTzXXV/3k5CJVexnh7ARFt0uQnrRSQxtvwzVJY2fpi31Ev27sgHSDe
1NZcJJQtWL+pHXKO6bCNX3xi59/8qIk7kfnqIt86YfQvpMcsjCFtnYrdGGqcz9ZIouColZ7Nd5bL
l8NMvs3wW4sQ+b+SyRo4/zIrrUYdnQ+1FOhwzdDUBcX/rUKXNvmyE9D0aDHWU6Pt9iCmSq3FlBB/
Xe5HSn+xZFQmxcb102hc+7/aRWXqfcGEx4EJeyVF+HUf2uFXyx5DX4jE/ehSZhSC6xqraKOobjs7
Hx7EU2V2Ing7pauL7E4+PQ04CrRguq0ENSPlWImakg5VlodV29iKUBjAva7dE5bUFCn+StcJRTC3
X99xyP03VsqfzJranAQwbw/FwNNORPN59QPkvqXWEmIVYZYW4R/lEnUzbAAi5gHEy3iCYITOQm3J
HsxGnBGLyGoflwE4m2xNK3+1FZQBcoCxG6SBUnyO7YK5qEwBa3S16PylPR5TA9Nuytz3zQ4WJpi7
XvKjMOPoOCl2jQBu1pBoIyv1x28O/PjRv6zYM+s+dst7idAtQblErLDoSrSIrNJT3RendnQhctUl
LCo/hGK67a36h82Ma06O9HpKT+ubGwym+OIqc+7DYvXRvxTcEBgYNr1mkO6Sgvh2BVZq6eAG0uNV
FKs+Ym7WrO4di3SBFIeRAgH1XZhFE/NleB7EjFUYi/ahmawPS2yInrYoCoiffAyflWLttASDj770
BwvnNWky4o6xRP8Df7rsCRGelsJiDZoJODqmGxxGNfqDmdcwaZ+rrWx0c8IeLopIPLeki2aUPkpc
D+l9dlk+t9ByDqhTXztbFJDkNGcGLS7vNkakK0i8ZKMF8aoe5CSTxxrEuOFxslysDK1l8ks7v+01
qFnWNIcyw2RqBfOEUoLm8GVDiQlTI97jcEU69N2uM2kJ0zYFmnxjtCmQfhHFECBQKbjTYUU5Iwr+
1JijeP9Mt8b1OtpcAF3rMH+lgwnzk4B9BiZAUyUje4a+vXOdwsV53DllZDTG6MfvMONX2O4Ng045
Dk+ZNScIpiF1BKpwuBkZjNKfP8wXBkwFxEygkC9fa1yvtvyWB8KesDqidcvQ/ugJBJ8cmQ9wujU8
cu5DmT9kOlteZW4UDxuWRs1WQNQaoLulCCbbZAZWyy1zZopJXJasAgB9N7SHEvhVTz6i0J5sGqRW
v05+CTo3QURw6h5eIooQyQWQHvjXGaDGjMXVdPaKKmYbJFcjhHYgJXrNhPUo3BeKEFDAXtqv3EPn
0R7KTAFSQjewn4eK1ajdp4wB589uWFMalKf/j1vRKQZL3uXcl8FxjfFuzpO/SJQD/M2ysbFsqGpN
5FxlO3XhIhPiAHXko6yvJNqK3TH2+5/sVm5z3W32Pv6lY5BG/AZtJEkcgpyudI51cj67ppFBTjm2
W+9JIeMbhTjhKQ+3mQuGHeMZqKtIczDgh0lXhgkY955wjJt6z8Njms8M42t+o7JFrj64mcW3BfSA
wHYkqpORswwkLdJ5/WQCWagwAC6SSzYFzsTkvgijmEe4hbje8vJZeGDV+7lIe1H96oOWoYUBiWBW
M0tMNSJiGpFdXEqpZsCB/rQWR4LKB3kt5PzJFjJEziXmG9IbqR3DQ/dh7N4kH2P1Es3jZVh3+x/+
tTfyC4kXukS3awzyzWmLCD9F4TZhMMMfQz9G1SE3InGpbOFE9Im2qAyvudTaMTcFYmt1PGytTQl6
bWw50pF6T7I0PH4YmuKj3QYZipu9ehm+6Y2JBeRh+YS9epyH3t+jiZPxwgjGULw6gLBOZCk1kqc6
MwgkD2Ygf43fsMtECldfv0IVvWlDr8R7RV1MBuenHMTWlk9O4V/1k1mQu/o1a5XOG8el0xWT7JJh
2BZxsgNhoAVVIB7WE07LE672tA/avq22X5qClBTZ4YR9nCLFjsq/5X/fSuYJT1ejVJAvFWFBmEPo
M8Gchm7s/8nnYa9rCW0kg5dWGcNuhdfKaYGCvmjpdrinVgnL0aPJccHR1x4uAmQS0uOf+DAbxxnx
HHgkw2ic9QODK9kKq7Zb0QKZjpBbtG69w0uoeZE7NPxLTnOB5TN4G8bbVVHjbeT+qznl5ON8je9x
7pFO3AvLJNRR9w2ESFgmUfgk6RJmTVrwwpBSzhaGWMfUxSqRihOHVyNpLQeDRmt5NOuESD7JxrP3
SpRu3kIyXI5nCGdD3mwZEplGQV51R/jXq13PCVg/euMvfo0ZJQUBxiDBuy1olivZACtoZyBRk8TK
arE7WzkHzne70Wf3j0lWaoBei5vkxxxiWsZI4NYzdVUMwh4bjeRueUzZIctALPvHlpm3S0W4c2cS
rirpRmIH5D3K7S/yxW/AzrMLXoirJ01hRru/k7rLiALkfpVdJRixoJqOZXtIBHKQahSTns8yNKZi
6jQyX3IMkkJoHFAPcocefMLc2+UqtPLlcosIRc58c2GI2jQEQVqFuEsrK/8k58o2ZB2QO7xhz4GQ
X/gjREpXYRtQ3Z+E1jJNSXoMdh6SBNhuUeH0fh+4PIzo9p5jb3GGWDFgqQa57T2e8hrDzF6MY8Xv
KToDq7XX4uf8zTFLY7/tguVOFuXatdsjtE/WSh9qooaAir4EpGoPWetEMyvmeRe5zl53DfzHCEkS
UGhiMmR5KDPWvCliZLjqoat6L/VnKijsatTTLqM9sgRLCNi9EFURzz56xjQAgLxH/fo/CL7O0Sat
yObPPvz7BbHPRRDxJ1X4gCg6EsWE/P4F1trIEP4L9h7If6crvqUHs5RNeNYUSYa+LuCeT6w0XO9R
hsK4v8/xpjCxnLzrsPvX7Ag8W/vAGYijoFopSRne34WfWYxa/LV5ttNJDYkVIEzVGmLvLMCr9SmD
xS/1TBmOmMPC1H85vsm8Ouiq6hmND5bQBOr5vRH5MxlRLP8XmRs0WgQZv5ItLiEOsD78vsqgDPAA
3SLq/M31mQQaB3DynKoNP2lE8rrW1qfIAvdclEXMm8rCI9MKJLQLhZJ7I/QLuxdI526dxn6FHwx+
dYo3CjmU9B2PA8Awgwq6TzUnWAVFXYXKrrxAbI3deSlr1FUzjSu0PoDWiI3WLsa0jnQlT68ywTjC
OjGCFOk4PlSri5lfPPZmlBnus06VHx5J2ztPWEZ3dL30bjHu2wZqPdN4hR0+htqGelJCUakOOyde
Ji2QHWysh3sGSD9uypjzSQvG5XYC8pNjiv5X6BsWdmH3grpnXKC/Q41diz75l393u0QevulPhhkT
WhlPy2BsDcHnDAOLSi0Uv3w216MjOUMVIELRF4qCsHZdMRcWOqMd2kWrCH1iVCVUf3iWWzWUrG1M
ki0vQRlIeWMAQbIO6iPiNNLLjwBg6fC+YSrzsdwKeNB48CsjHSiZ0BQ/U2UwosXNhdVVyzElnXgz
NBa0RkzMJZjz82j0CqFPLPfKY2pehsWnjZBXlIVyndTCuEjZEE5JCFgmyL5mxBrCoHQ458ZvvuFW
eQ5Ow0rixkHNLjTTDVFfPQOeCwwaDK24VuFtY3/LtncwlPZnECpAXWJFfWWgIiErBex4VZkt3heL
W5iK5T217wDawBXyhe3Ev6+bjJUKzUPlQj4tZFNgI9h29vMwbCf41fFOaAiscZ0ZbP+vI9/f/kah
83EgSIK1+jp4Z3z03gSCkciMHomEPe4fwRDBrifDP3A7L3l8x7SXrJp1sy7oQs2/9/d1XR/Na1lD
kRMqaHY9zzHVKSug9bb8wfEIbUp830jsMXmpr8cvU3e0mS5n0nnv9W1qSmI8A4ETujLo3GpIUoJL
lN19KOczpBjZqvJpTvzlNCarlOKPfRGwZcptbI6iYoeCuUDZNnKfXZU5fpSpH3gFVJvqlKeJ6uCK
CqMXlgDnukLUpI+9x/F2OTx0GnNx2hgCyIr0S+XVvMqTUiMQyR3AncfMSzHbz0+uN5uEVydal83A
ZAWx0h5Vg4h85NxR1Okl4hd9KTKzv25+HGibdV6tQvKYF8sZYA81HHthm6hCbek0md8FHFcRJcne
+x5HqFVPT5zM5HCYIUqygc5+O7URi/iVeS8iUp0zt9ozVIGBtasj9K5NClp+fGNLX8KiuRaWRk+i
F50jQ8B52v6QE0EMbDvoZyu97sLMJ/UC5nlJ0NL9xDC7RGBWxDOA8iYqu7/UwsJso8LGl5FSpArQ
p7tOyKWEEW9mPct2yc0fhqWrWme/iw6qNHyEb2KpSv7yoEiS7YJS854oV8YUvxtcIBVWHtgxmnw7
xLOoN0YTSlVt8FsBAG+PWzHyPKHEgxYCGWDsdMJnOIXRNJdOraQHVJbbd6izoDq1k0rd++o8gkKP
qgI2KNFz9wHypcqOnR2yi610PgZZmOm6ZTVtTRKiCUE8PmYqVsp6w4p1BMWdhW7bNCBQRqSxZNxn
bvtrew4g1JbKXfKdJQoYjU2fmg0PK1woxGlXWVi9h/4OJ6gs7MKct3WgQ7wpHZP+/gmv+j7Mpatv
01jG0KP0niAUzGkN6j35wCHZjbfOj0i/VZnz7S0UcmtckdC4vIKP8NRlYmDDSzfZXEgNuqvT3iRQ
snbtai1ghXYWAejRmw43CEEG9arOXcoCcyg3+xyLEoSI86ngxe69y04gGuE76qa3DgdeZLmlQCv4
vm0MEgVkOn0qUUe3d0a5mcfmPYWLVtbrpFH3w6Sc8FAsLLj1DgNdd2JJUs16f//Y/LsoqOdmtpzl
KFSRldCJM4GtTjxI6DhPezakqHm7Qjlwfi/Kh/t99sSuYA5AVOCMl7vElVPPeMfjh0wNTcPTHrx8
ouQ6cW1+r6yfM8RWhE4SvBRUidJxMUnD+KQxuzvHFrmw55vbF/1KNS2a9mdH6rYbE9ua6xkni4hd
Hlr1HcQmUwScMVW5LVzC8vngKPTcF4Aildxr/5dAA4UFmajzNHdrSBKEUZww0NzPPwfiByfbhzeM
qcIiSyad9hBCYavMOttirCPleJFVLe9GofYcV13fWw3nG8y5YfwK7sDo++7b4ajEHtMXbRA+cKrx
Wgw0vO5kpaj9T8cE2TzhNGs6l1qsrR/1LThCeicMayP9e2Vh6abLVtKdPxpir9PeIV9yMoqBUw62
244tGeNiSzSJhsTS1/+GMPMkCHuG2Tn6tFHYIQAXvyJM7Mkndrl3PKyrtHfGwNcQbxPo8MF8/Lkh
YOn1UYs4VODI7zAEE3pR7sTCuD+cQ3tPt9XsXwb8tiR5VwP56Zp8/Mt63veFjbjHqrW9RdT2yW1l
rVfzOHumR/T5YEUIrps1IyqCr3j1nCN8LqYWofCXXRlwG1EA55au69DZpTrL6Au4+ZfblUx3RE29
XLcPAE7fq/yd9yE7zDo/M574oiyFnQfUrbv8NMu/5W+S3tA4qxE+xxlzGBd7cr3mg6TcOnTruqSM
R2T+rAwPN2L8NhiMZ7sGDO/aFzxOOOrc80Z+Go6MVc9mFj3M2hB6goWxlS7tqW/C2db9ygLuOz3T
GY7K+A6fh6oNsvOJLYwz9gJdsAXQBTv6yqPf/B5NRyrcivfE5IN07UEjREv8369KIOfaUpJJDvGT
LaN7ocQjKC2ReTRscdaWUAP6NlWf4EfvpgLbVSvbNF4rG/2jUMkDcxKWMFB3ek66VEK7W6xYUygQ
I84F4wpgLOAwSW9o3EgKeE9+NFhEWMIjRjH5N34wzRZyg8a7rZg9OMN++onh/sFe+zUyK10U74ty
unIiVoSFx1zeilXPno3j2jiArb094cPaeM5pTcR9bpP219WT8Cnz4MR+xfxMvxwZIvgQi2ZMIXge
PyetqSdZZ9d55Pq3EzkdDf0jLmy/d4bQLIv2pbNN8W5CQGa0JEUnacR25/KsBh6Fc4Esx7M5Q5RU
Pb3B8qjKZlePba7NigtNbrxP9Zt1I/5XJNUShsO64XCkflF2/9g/I6saF/9vyjngq7x2AyK6PtEb
W4sggLwLJ/iFe2temE3FYle4zI4rbehu/9zT44vGXo4djGHz6S41H9QsCbk2AzrR7PhiVGp58uVG
FwkIgd0yZJ44vUUG3u7tqoFfTrY0HTFjDd0W3lCA9U14j23SwQF3hw/a4ZpUW2HbVXGG7NqHhyx6
RT6M5R1B3hPDLvFYd1fXkZDmR7TQXIRGiso2GTPGVcd54B3vrriLDGjRFV8QHkgUfmeDqWgeK3+7
n9USVp+7671R+nUXnzB7cE8NgkYjZsEPYpiWoRh6fIk4f1EhoZXv5omIPC63BQJEm5NW1rXg+4YQ
YJj4R9pMzfclWHmuW8mokmzmAAO/S0wAbJ8mrRBZXeQrFQr9M4UsSc7ToEf38TmoM+TIYHxMlMET
Y5bvIo8VPf2mJkJd47fHqUy4kZfRvCmWTGAG4Na4ZTvoQOhmZ8W8DkOtPIcF9JLOwMQTGMhgdYhg
4b83nkaBLg22WQnBOwM7vCbPHuJ75jFHfUVvNqFGab54mQciOQQ/LJghbDzreyP3LWPZVOlcKmuW
S4UN18fwlszbQVOTNuGlbAeWuOJ/mKC/P0YPh5kbz0RMSVCuxIvgz8rhVpAlJwhC0rWbVHhuCRsj
GQ+p7p0Hk+PUqO4q99Pg9Cqw4fLHJRDvXxkxyggy5ZfoyaxEzCutFCop6kpzzwwI4jYvBnw6otvr
zweWSnTuMcAGG1CTkkWhAC7MC1Vw1xUmJ/r6VcV1NAWvwwJVytlYn9nyERKvVYxRYhaQdNOP1yp8
XyMP6rD29iKY1OV9rkfgIuV7BWCZfmkNmx67FH6VoE56WP5guKs3GMNl2zTInauHiSJxVvEpoL1j
zTCrPcLhZ77FRiWWsV9LijpYN6FCmSYKhVyTmK90PWjHTBfv6PvpF06NXYTf07p+rdVJ5fOHAufk
GEmmy9ZEiKriycTC9V4NAE/pJAPUhatVj9BOt+maFgOHyKiKKGkIopzFgyQ3Y5m1ytaTZrPE2S7K
+BUCI9n/zh3mkvplbkuy2+tK7+0o4f2lNY+YMD0rf7i5M/sE21sJAyyGfcvOHfrLI4nV6KIMAcIT
JPwxdQlaE92QVZeHGAYxeEyietfgIRqyb5JXZGda8DTfrAO3OxMQdgCxa/PAnnGiYqKUBFWzilU9
Y4gEGo9NCttQebDOx6dKcPuqFs3ay7CI/IaZONgK5jWP/IauzYPiWSO7vLR5u6aJ69t/rLs9MUlB
7Qt3ERgIPBoQWCv4SHoYcvmtw+K9X42V9QhuIr/KvuABDnWRjDMMnT0H4PxtLQXU2yCLtZHrCkHC
jA2p8fV2wKuq2sOoBddxV9eYnINR9FhRTE6wDiDQ8WDlQ/TGGnYIGs25agL0I4ezBPjh1Ugp2f4p
vhXit0py4ezvBivHKebfuK+YGVz7XmYY7z9fF3LDxTHyPDvgs4lqqArRN40fBC+t1Iz2pTmYzyIs
9Ca4DiaJGcPepfeU7RMvTFgEo3if7zMYO1F23ZQP8kC3waB5dG6UpsPIddivVPHEC4eMJvWIYg6e
Fz/22whLJZRDYcB14Tu+ZDmbe5zz8YHFMuctHVmb2oq+V5NHySlPBMIETt73ixuPiPLrRIGN+hE2
jvgU5oVVn/VNE1HRGi3dg3UEYipLoajzs31YeJ+jWhdxMBuJntXzdPgPRgQmJWtMnRcHF5WsPWFt
HsLPpNbn3kQ/qJ6NQ4NS1mLhVnmkPw5UE5yHhbP0JwaG2ohaNlCQMJaEWOZamXckk8oYZVu7S3ep
zYBdN4L5m0qO4O8WFB9mssuTGgBNvQ30DmltFm3v4c+hFowJpB5FMxsoFVMXzt7ocLacFQCGrn/u
GVoUU05cAKmaqMq1aUnguvJfs5fjfvqGKT7zS770KMf2WIMosbo8zG5/KsSaljCYU6JFQEkhGtOU
K6OIKOwG/xftiuuni5tLI5VixnXaaQUVxOTYg9+XvO52rgyeHFHZY93DxXXLAecJ+cPvFVwXdD/O
EAklvzLG8jrgvAByuwKqkJVnqGsYmGXNAzaM0oLltH+wo0O+9V7k7bIzOvGLxFGLHdXrViJIBl/R
YkM7xZVTDvlCE+2cQbCbPKVLgtvqcSeHDiE5lZTjNHkAWs339UdUFANrWRrBB2Zu8A/uyv2z6OLY
ZlAsoiCt0fagCFAfUrevpVQJQycK1gVwJFc0cQqj6CNr6f690UJmHY+UyW6dluQxAoM3cKksyR4T
R0LydfyUcOfmX0rYb3eeE1p3XbEJZwUeS5fALVx/H9lHM1nuuHnVmn9YEu9vgilc0k6DlH8VhbD3
ZeTmPbn6kesArPixFCdfc+8IKZa21KyGsTKw8mv0Ho8VK+JnVbG27nxZ1UIUiI0I0b/oq5yBcpAB
HDn+qisyi9byIKQfMTF0XB4ZQZL+FwDPEjkDnLr7cGBTVrHwldUAk6lMnfPQNdilAO2ENxdnanbQ
HOfTi8YWZA956bChvK1nljBLsfqXyx+UaWCVDrqX/3skdArkADLUfuIaoPTgl/Fg42bO4XrVzaPW
TTWd28pxU+ASMmo+GqkfyUepW0Zm5OUbdMRgDL+xv9h+5dFC/qo6MGe55Or1njdiWyvjh2LN1s0c
11EgJG0YvBOXybveZLupLq7VEktr4LtO98LlMT528KIFwGgYWcRZDlYNqO9ACOZCvd2Tr1Hj9lsy
N9OgEB/MWKtgj+Xq6Fom8iSse/WdByr6+zBUEveH2qRV7iUovp2UhHg/ZI1FDKOyedAnEhAzkj/q
I+rykRbXrerN4wJkV0AmJEmjVDy71RggJDVmy5HhVDMvc3wJ3EBT9GhiGGzbyR6RIYtyrxK7zMNw
SJC6I2GbdCGs7VgoLuo5JcEJRokKwym0bsZFpzzejfQv4P/uKcbu65yI1Ufod9FnWRwhW4NTvTN0
JgmlMLo+FIqNzjt/7jsKuMC2OG3P2Cwd5uCm+peGk9p4SvZW/pl0HHco8l3jdTHRWmSd+xBOOAfQ
4cKwUElj+os8BhB2pGBkUAkM+Gs2tpnAJYUzh/NfYoW6QS0dzqcNJjenS9GHJLCqCCLDpJndHou6
i93jeCuzxhevTDxafiTUeORzfZoDR5Yn/gi7MqN5X310S/QdqcPZZ6lxXjd73Xt1m2GglT/sbdY8
qWVb1Ax7aHJhvc5sT9Yshw3Si/SBZBM2GGQt5smvmFCcFcq+hCp/nvxhDwtBEjyvJ0J2zidxW0NK
haGywe+EkUnyscIZUkApJdx6Ku+M1lkg2kEBJpTgqK4IvzhRaceEDO6FsBDksKiynu4QbuLPlvIH
JPvpqo/c8dbXoCqDq+KW83yMMd1OvNIdYjWdGAVBBUaabj93E2E6EhTr7NZlr8mb5bMzSxT1E/Q4
uzCrKRdmo7V6v2/tDKS7D/CfvS/Wl17hB0QJD+nfjMCXTnRsjN50O1gx6uVpnnPlaQa0Tdo45X7R
DpM2KVIislILVwHDqM+W7zkN2N9WqlZKk0Rp/rKbuDOXonsoW2ab4YybxUMPz9fy4K5uZP3eCneL
hKNnwCrtog543cs3/UzmaVlSEgKe1Xnh5Nm882i7lxaxb+dwKdJILDwByapHryKyOrzW3uCNSwGw
042uThYmwKGofwgVzmzOlRiw/7+rycRZADZRQlKJKk95h3spW1mncGPSRrrMiaidrpkp4FS9CU/T
CUoB+hpfBIQo+IRAkkpV2FJcMSghG3fnxSM/WxQOb12I6ky5q6ybe1EkhQbvg5iNygRNxmeU8T7C
0C0bRo+fL4ARw50tFG5VpbQyaGilPM6gGamWAJHMaiI1YEQB57SSpnBYXQDQUskvEwhEdK3qUm+x
pjcnOXSm4c/TRuhjatsmpA3KUhTGN4TthLkx2Fsg/xbzV0vF4Q5456rFX0DQnaVGzVEzChSVT20X
mrXx0rcEYDClVNihVkmxnPD1CHpseatGXfLVRsU5VoBESq3dZtYlXRkjwY01c1UR3IdgisLo5Vpk
KuNB1GjzvGkrylG9OlPd7Rruz8m5OSZXfewP2e1mCQDbwFODU4zLBMHusP+z9tBEXWKqQRYErot4
qqDKwLMTEUIfvEooSaac/VstW1Tucu+WdPs8FSGh2NorAn7j59f59awfJ9Oy4tGRpMihlpKLf1Ln
eSaXC6utjvZjTnLyd3KDWjadI2Hib7IUu1evqwbrVCUXMI+XCDzqVsVZ3UV0nTvJhs3VYgX19/7H
Z/PZERpKbvJ0j49dxjlUz+01R7ftYwlyvO+WGn9rivDgqE4qZI84zAvvy5W16lMXVP9X4vJG/iIQ
3WIg72iH+2t+oy8ITRZrn2OIBWpFTZ4UhwgEO4Ve24vZpyYSc9TFEzvS9aNUFqWNAnXhYRoL4UrJ
v8ecPnec+ahQiW50mP0CruceBh4pOJXX+lE15L/sQtV5oyjN6nW3zSpY+Hk2Ece2nM87vPYyRw/o
dmVe1fm1j+/kRASH28VKguyhxQlzVOWOVwuPz9Mp77+eD8LobZRZpppAUpJUIVuHmQEjphFmtD1O
BCSsTiATA2UQxrHHp6ojZR+J9bA+/jiTgdVX1ALiefBlQvNB7ycx0WAu+QOnBZLHWQtXQDa2Uj5k
af6dI4S8hU5zY7uGp3s5A44HiO5TJVeS1hDEzXYA4sFD9L5ACrrVHmiegWrSYp2i9umTtv6vaRCC
dCLPc9Gdsj6flMnpa5C93WkKnvEwbkGEmrsy+JPHCPUb1lCkgW9jA0QpENXQRjkHYG4MkmSoT8Bl
AYr4NNqpNfxHaw/qw6zQB5i0UQarIJdFLyJGwhLa/zOWkXIsN5BWeA+NmBC5dqBzbsuuzpkfP1Z4
V2DgIDKfAtpJ2szOPCNrMgDcz8Fm9nbhqa3ZRW1JNmjDqN2oDRn/ohbXy/kW3jdzAhZ021dkWnCQ
/kz4l7DHAbyKE0x3nhPK31xIrSyx2DXUraLRyaIb0D3fw2Q72Bz3ni5uUDmEir03ReJ8rX78V/0Y
lky8beg4GbPxLDSVkOVgFYRWDH7ZtXUMVWq2MJwm4wPXSASpa3ZJRBDZ5uAKCsKVPwoiWVjGe5Nd
Kj2tacfaoMXtmScuDb5YTk7BguEZSd2MfRAY6asJ4dA62l98t5QgyonZXlIKCNmsi6DZg+bLH3Tq
uL3oKlgF5cLuUjumMBZI0Y/KVAhZiXuCJUgI10LxMKyBsIA/qX0Dep1EiNFjktnsa4JZ+GuxyGzP
t0SggMaYTJNQ80Wne8CiyTaQLV/liQbI0VBYGHQNrQ81HSn24aydzKHJeKVtKD0feQoD/N1aQ6Wj
UzJlu65zvXLegMzCFe3QBLEGZ0gChgsizv0n/okEAptMA9U+lFJkRu6Wp2PkhWzwcsKC7cTKViik
ky/t7TAmoFGrVaDO/2zbs/HAMiGCVHdzwkwNdyQajAFRMD/KaNXUZ9hxc6kDVaNkwsLaGFzoljP4
F2H46YLQkNNiC0osigxM+q9Mi9lgasysIBhzOosQTNY0q6MmxxNaPmidsXe27qLu9ZGILTzUVEQP
cLHj8hb8x0OabqNunG6U64h2wG0GJ4L5lkMMFyPjLQfFUh3G0iXV0wsCdkinSMW5oAg6hKzKveFF
yL9+BRI8oQNhVFQ9NgEMPtkVdCJpJaRsyx+tvwA59U1a8rnz0wVP2RVbcVyvLq1oJTv0Guy2+qVT
pvAuDMpxrJBaYcTBtMOGnqXYwdnJQu5Sqqm8HcuCKyr3bR7nYdgH+qsrQefYUA3PKHtWeivQYwxK
1ULE6VewIh1TJP5a2zss3Ep++q10LAXMlwPTYgZAlbYb2dMjHF8VhUbf8AcAaBVv2qqQKu48ez3N
TiOVf4LLcgBepFkyVOhHwlLMPjABNmI91HPTZB/6scKj0u9VpPPq7k1is0t3o2vtglbSk1mI8hCV
R/qSV2nRpbFUZ0jriO9j2XutIVn2cd0KOrlfh0MQIxepqvtB3cO2YI1MkTP0vMfhr6kZfMtlTK7G
x340mA1jholBHJroNCHAbhuzzmbf576oQ9MLu55XbyedlsBgZidFZWFyIO/qGSdTuDfgUfK5qED7
nOtkigDlSw8qwEEvy29zVdFqYB0jryopR1fzTB2Lefg5KOJIeU/IJUe08B03NpuKofdQmiLAwljZ
2gQoq2tfUs8kPdOZSTwNpOp7O2Ch2NqrF/HYf/vd0zFvE5vW76sin/t+OY3xOWsO94bIgaRTeeHv
TOpgRnz6c5GHONdbH8a+r9ri5lg88F4OX500ha7vu7VvBiPSDXU+I4eavW0Sjj3NfwNQqaqTux37
cn0IFfIIX27HENa8j2eSBCLfZ/ukY6s5K7Sasin9Y3ISUrkc0dS4vC5Ba9uVA+zIn/F/Yfq4G7xd
sjOnd3bvYIZdnhLw50kevtPWNfaLIhSxuNEQ+M58DnEnO099cwdDznsjj/pZQKW1Imak90Kk9Bj2
GnJpYvnIqmlLxlUThsVD9kEft0HkEmEi9huzac1iMsVOg8SqXVvh1gMDwk+qBJLKn/HtYec+ltJc
olMZ6DHZTpcgSW/v0zKOGirBadVbi8kQw5bxZagPTo5I+jrI0ic4kilMzilS8s2Xm3HXlNzdMije
z0W8GTp9J9fweCKvxJmRSywCwpbTYIAsfXYAPwB5BdW8w2olMs3h+IgRRy17gzNRhEkmalXN+yMk
FOchSk0lgMDwTsJ+OuzHVEsO7buQ6cssoNaJ9MANzm9MrOVsdMeyExu4HccOZX6Q+M4I69dOfTw7
bo9iuj9krlX3MwJmkpOwXlzmxEcRXe8wQ55Km0B3UQAQEkwMS7x1WJDpmXQqY77LELdqn8F1exIN
yQ3A302eaML60hyQgqS7rL9e7WDA6p6iCeBUnX4IvNNOKNHmpxYx1YwmG7qDUGq7haSJQlUBKt9y
lXAMjvq884/Ak9+S0b3U4Xv1QDf+5KFG0IpHYsvT3M6IAGYARcEurpvsEfGV9yTJJgd+soqTnLFx
Qhjgy7tzmMQyV+Wq/JeYpADA4XQBTMsnGG+x8dnif/0iiZh+oRe7aD99cLZRHt4QCCSsVD3kzS1y
A4qNBfcbIuEgcKkaD0MunQHiKd4ZfD9Xl+3IDnPO+RnRfRST9V0TB9ZiTAWIZ1x2ELXSwCLq6MEG
p9Rr0fvjT6oxZhiZvzvqhaSc9nIXdsfq8hbI66cacFe2rlb5jbRYitb6nr4Hue/iMlPEDPyB0PN6
uRjaHaMZnUnHJRC8etJaYX+FNW23D5A26BVNInIaAcn/lCm9jDzzA/e7j9T7hnDQji4V2KdmsmfY
9KanykqVLhl3IsUtDn13L5ElXWgRyPo0X72HJ6x+P1D6APJ8KmY2nKF9wzOq6/lfcvI94hWxroPR
liqpjjSn4m2ndfxUcTiynOIgPZi6tkKQ4TMyx+4NRQk4KzrOx3NaQPWWVWMGY+3t2SgOBinvpgPy
CWiOFOt1FvNPnfRfMhCSYiti/B6b5O0Fe7HREuNan6OzU7DueuBmy5nurZyqqZs8EJpR+0MS4L7j
necLIEit+ohjnVCtrAwjXYUpAedIhxRHkMGHdYJ31Kd9ljYmgZPZfK/woBRpo2dhW09V+YfEiJ81
lPiFzvGS3gvKtpgHKEtKYXrLR2JUu8N6IocwVWdWzS2/KoybV9uWlYX9+MVzxdXhbJgzNj399brU
WfRC8pYFDEUn9Di1d8hueTus5Z0Ial4Wlyuuf1Smotqb93gHSjEaZ2VrEOgpB1a5j3dyu7sFTDpu
pwcIdOLSQOApQLDZW9N1GYXoEDBCze7Pjzb7AIMoGE3TYtjFS84yC5BPwoELA3MHnbCw5nD3uaV8
8oWoaVfo+uGvaN0MgaBbEyhqGoLPoxPFU0BpC/PtPHhoGqH4LJGCDWhKdSpPC3PqAcN67z3fIBAV
eUE+XfPCfbOYSQ4hpcDQKqG0E6DHLP+MB32YNM3TAyFQZyl7PSAupQdm5otrHWXe8IVcRnDR6lDv
sxoLEPdbHA9C8kzzF84zvRYX2hhyQTwGTPm48Pd4xDm7fwCW2QdaiG+AUjhqWOZJk/kczDuu3W3g
PR5YZqGyqv24R8Wl/ufjKGkoEU8RgVn0yjiri1LfjekdQiqVuH1k5JSQgw3s5SpIh5MrvSHtEkEy
fC0YZluDm4qsHubxILQiJy6VtTHcrMC0eouW9caRPuXbhU0G+gYaQxi+N/LHIiqPUoQGblpGVKNp
uTdcVmaQBxHhoKUV77i0AmmENyNDHeps6sQCHtLR+0+wdB+eIK17iKUO6NmLodaHUQy4XxHqOiSZ
WW0q3ayfFgi96pO3w8jA1HMw0ps9hx4TOV4i2kluKH9lHuoMqiVK0QLWTFqhhfB5PRUX7agQWzVK
OHp82+tyjst1O/s5YRDu09A7KQl1XyriKaWHRibODJT88j0sZ8rO2qzIil0FDvcSibfXGpv3rgwx
8k4scXqmJYr+3+KuPmlZWpb4CVkMg/taHmmF/FL5t3NYv8GNVuUrPbUOm4NYpv3AZG9NT+eITpiv
vDETW63l8l2aX3TUxaTx60Hrgd1zuCvRxnjWav41bRO1XRZcTHEpW+WFFfkOYJdxvGz9h1g3C5nj
JTX7uMDRstE1BNrMuh9XVcsT26am27eBTYOaF/BmdpvXLpwNo3YAIHt6Z2/sDlgXAgbTWDnMjwVr
miKtxAg02HAls/XTJ2IycOcyXb/UudByikUbCwJY/f8KZmE+Sc3ruIpwGlwRlyh/AxuezvbZEGx6
+1qSyXWM6nLXOMOjbHPQXAAq1Dv34rq3ficDEvG5NaRCb04tllTaWPVmQ+sNipCWczEw3jAWSJsS
TCQTpZhNi878WjiCoxyMasOufqp61lAj9UbTKmU1whnKcnMFNLwnL+jNtdZqmD1GK9KQ07Jz9/6N
ZvmmLiljvicFCgWS74bzLoGwjN/HaoVaAANdTU8E1oKcsyQyvTzRezTK+C2LYxNHH+M2QOBLkEvd
ZMNX8Is8p7BW0RTQA4w2aP5obVmo7n2Lv4Jlla/73lB+xYQ8/4PUECf9TbAikFl5NjfmEqJeKIcs
xEE/7XOg2SAcEoEw9J85doqbrs4OPjYncAbEZHIsul1Dl4C984FEGjZAuINunrFzGtEYee+JLtOF
9kXViknioWSeYIagZpJUKcWgu4gduPfBjA3KfK/g3ei90dVBzdOpOaPOtntc1qUja67T3sFSF2Qb
InUTQHv8CPJW0V8lXPM++7ipufRFQX9gK1IjSI3KRQ9x9Nn0MQfl5TOfxkiWjGnaD2f/5IA267LG
aPV56tyJlQltrh4udP1yZ2z1qH/EM5sfMRPx/1tn547SH3S7KJHJg675MRZcctyDFG6Y28qbE8RR
+E2FOAn3lLZY2aD27t5i4Hv/LtcOAWUdnapYBmMiwQpEANqXq3PsIqrsh9PYwtGAKRv+gSndwF0Q
q75i1TzV2yfUxp3HFfhbMP+HawNZST7CJbb3VE135wUHVSlVVUqv3rCj52mwS8kFt6S/t3QBznFs
JYX0/ULJcs82Li3ffaG0XNi73t2GyUiun6i5QlUCjN13rrI/lKgK8/RXSOqLZtkByH98l8l+HlzP
8bmgg9J7hllGDs+LVJFwwhhhqUaI426pAggYtLkvEwMVJeB6bJR5skeaucefAsqgtpKj+hcl8KYs
q39TT5uhD7G8dlhWG1DtxVcW4TL/hWhuE9C9if3c6k0i+WbaYlKSrSZ9dhnI9oWTuAjfUDTY6CQP
hmcxZtTF5bVNKwBd8piKIrnxoRbb9drqu8D5q2FTyb/1LmX4kgbnJ1tExd9GaRTYZOnvJEdRJXKi
rm7DRyG36mAFlc4Q57SV3U7WB1UOvywGWRDJoIqMD0R55/wFfF0hFU3MTWyy3K+C9YhU5XkIV4qv
Z0YYH8nSGDY0B2yQMrfA9Y5nfSftIPNc/D9mIuj+2htExBWQ86BUB2peYfidss8ZzMabqSAVx1a8
lax/gLC6CBql4TO9MnO28CA0bIu+OTwDgwR8FaU4SuzmZSYox7orO6WWpGz7u5lqj+0w9Nh7xctP
PehbHQxhzbfhQdJnTpGjI4pVWlYhUuRSpidg6yqw3OyzsXGATHW2Yxe8ECTO6UPZeh01p8KaxHPX
N2N2EwZIfykXoRa3V8GIiL7Mb0Y1YawGtTfIgW1Y2rTzuajzrCD3wonxgpN+ogRhk7yyXY+MChZc
yXBSjgep45vZS7S8MYI6EfBeFwylwwcaUTj2LGA3QlUJxF8p3kJSGLChSyfGiVZEPb9D9GR0YOI+
qnSi6zAq/Do+h0sE+WrBz6xLlZtPXbmL4GuPEgJpOnRbdcImwa828nUxIuv0xNuod3BHeG0pMmB7
ggpEupBH+1Gv0mBvyAqItoA88IiBt6eqYE2GMKcvw41Fc5OHmeapJAXPMraT8DkVtPKgLQ7fxIOE
rkpIdWGNzxc8+AGwfRi7KGhZM3RCYjHT0mA3JBhK60M1BcNQDJ8O36aHooTJuo27UMjY/wVBr/XM
WSTmkAdNfVkyyaQA1EClOgHfoLxtTVBY/ycYX/h6hA7KwCfpwXaydDbKaThhgpO44PI5xJOVk5Xw
Y6zzBpusRadUd63Xf14d5cWFRa7FQdWxFsjStmU3+qOi7h+cSrcwic0+rClHCCv42Sp6OkCh1O21
5MQJcmBoL8Dy4WKb0DA+kxSty5dqYT2e8yat4WVDrPEha1IB868jtFVLK7cvV1GevWAFzDzmYQKo
8OqgOX6/T3oifmEz8VPFtKEzSIc8xuq0w9/I7mDkiVaw2Wi+rFTzZymMt0LuK9TvM1/ewDw740HR
fYY20/YeeeyrwIwaeLn2d1pLp2VlKUVL84ex43Jyf1oct+umSIBIXSigpswpLsWLeYp1b9COCU3T
Nope8KWf9dtORx0o0JnncxRm41jaVLUBDHbeezsI1ZHxB199WG1zuCvL/pDIN+Av7j1hSq9RbFoP
oxTAMun2WTCjQVXag4uwiZFSovyM/Ve8zIzrywBLCVMt9RpbjwMmBQ1ikK1gNSQnap5ka8l4dN7+
046cyhNisteoNVVvlQQYzvB/dDxtrgPRhJc9BTzf2goIxDUOIAOZXzyVkhcUOMb5CseBBe4NuHHr
CuQDgcYT1QBQhTfKF1LX4bWP2lNQER2C8+8ZndmnwRyhmpTNuJzNAZlbpxBsw6VfUWHFzrM8Nj/e
ZIFJZuFJ+9lCzxJG6CKnM8HVFRhmDwiR9nwGdWjhjvzQRfyx4NGaG7MjVUxaVhMhKs+MOwn+EPcH
HYwmxxLPM7C4nYEFFMHUb4X5zR8ZX5kXNNallP4qfvEGHSZEUhTyEUAeKwNZEudusfLop+yLt7sT
k7hMGmBT5zX6ufC4KjKb4Ipe5N2weKRAGqulHfBkgpghdumO805A7LefWnf9IqEIxZaocI5pNzLg
RocefvoFkBkUGJqE/8p/7qCS3Y7OTdFDprxeD37J3iR3IX3Zbh2f8e366q912If+JqE78FO/MfyZ
YITscam/67+QDCuJ5rPSpObdwu5tnZSrSpf454Qu7aUPPohMaS5y7jFDDukipf8CqIkfnfwofFW5
71/b+XBK8h3P7rEVcp5bRumE9y6B0VlZzL4032gjHPxmRtEz35LzCBlf0K1lomTdvWZeMUze1nw0
f+tqu9iQBLUav+CaHAYVabchd++VAIslW30zutEK8hqjpNgbve1Ia30nSjeSw1TzWISQ+8bWywif
fR5QSmjVJjaDjuwqFWf+XXtaTNwPSNfMwI41GPIouBbbLKq1StDbFT77ZMJvvHiuVhh6cjN1SfWr
6qLKpdnzJTFdzy5Kal9e787N8OHLeBOM4CNG1MWADz4N9ytYyf986QVzugs+qLH2Y8dBVnuOI1v9
dIJsARGgG7/Kw46jL4SfIX4DlN70C4fFMSdSmrkcju9R0mWEJpNCvb+C9ggEyY68vTTCan/ERuyV
KucQ8JX2wFU/pBpgH6EGcQSPsiUgo7rOxV+TjrqyddvGqu/r6nfVxU2zSTEnQlDol6nzPZ1up0E2
Gvc6mdUXDPa0GHmVOo8Y8PDhehqX9beunoxTjY5dAVNAakZI/STTPjkVzPYyGDJuzYsktOL5RGx5
byHyS2kkni31zhCdxKtqSdnJKdahujbk6UZJvh32ZzBDq+m8yIvA+ileah1izaL2XEgTj7jjs+u5
aEZXeEF+Js+4jVs58yOOpeG+LENELeCXL2ohWfKknug2UNNWErSPrhbjuWKEu9SuR5x+Op3bfj4f
VIGj1LSAvg3khJqDFRTcfPwmvENOdODLmw8Og6DpW+WV+9gRww/xcH9XCcop6cZCpntrIXpsBvNO
EoaGByqYrK7vV7GIA0weEAmfMvS0A+xpcH3qdef1zVK0jsS2O7XR3xO3Zv/2jNN0+HPEsWGN6HqW
1142aNfrGcV+HZ2l6qWCIHhTjkupOBZ/4scZoZPn7WiOR6hhPLv8qqtHMWfs1/3mtkxewTo6ICM/
f5THnXN8S8dSaC+ivmgOShqbmzQc2R4MSSnbxFhfAxfmRrUIAWrJ+ghCVMKz2Iiilxa6P4MSvDIh
MRTLQFaz/g0UTei9859XohKSFo4fBIG7deciPKUrigU0iK3bdcFSkn1LGPvyKMfhPfECBO8c00IO
KKRD59/F7ybrdJyX7/TVhgRzWWBg81kN5FJFyEwAYtQaHK2xMrURpdaa4DBf9Az2ge2nkjMeqr81
9Uv7ES/ek0J8F5xFthqp+YirlBMqavP6CtM+Z4tAPYmHvs8WoNWb4mUvC/XSK5qrLHcQ4Gfgi38f
TRis6KRsHsH5lBweufkcEYQYbL9AN/rikqMPpsGsMzHCMuco9bZ3+ODSwIideULgfQnmDw/GYuaC
58UsBA5xwj/y7OYUZA6afIGbj9jRth/yZCT4DSATOLaEtYDnFz9vv/ZnuRAPRFemzcWJ0+MBWiub
TeubvYZOcOX9hzjsjFwtiJIPozurdLlO9ZaaHHEsUgXgnEazuqDc61xhLFhmygNqpXSfIoFxMAzl
cMT07w7iztjW/k2HZP3M+BX708yN+sn3oEJ6dDhtyAjrjaJm9CljJfunkvcnBp4sZQn+sTqa/BGC
YtlGyX41SbZ8RKu+z6n9DO+M2ZLURUgvgkC8xJncRT81w2o4WwJM0kQQibOvfq2VlTjFxvlASArR
wySxjPin1Z+gr6T12YlYaCLkoVx973Q9UYqi/ES/mP9atESVLbirYb0lnYz7xLAEiWD2dWwStbxX
kcXQGeLihmNiXAZ8L0CENubRmafuybzpyvpTCsMxZzEM4fz+u+mKXuuGkV3x4neGxoO76Vk4q1SI
pXjIul19TAB/LimZJMC3tQtOL2HJWu93Z6pvn/jSfn5tGfdzt6HrpNdPChiw8YnsL8rKCLK34x27
ac9CJq4pKycvxTJ76SDNmuyzbN1APEc+ISdze3zPVDrsFQCLtwudTP6D3VKo/ml7wzT075HMtRDe
jr+Jrsu1mAIjO/LJHojZOFeJMzzOwlPcr0Z2tRf8Afp4Z2TkneyCcQRUTtOYmUoaKShi2eARsdAM
WwitS0L4v++KjvdnxW2Z5cJkvkB1KspMA66HQAktfhctTKcqaOn+e/SFeW7S/FVh1Mg6E4CqiIBn
kYFhJ0YYElD3ygc6DRGhy2NGW2fzOn6MpjtCZy92F7ErFMLA04/yCe8O0VP+BoaEj8a6PpE02G+8
y0AYJkfT8b/RmEPewodEGi/b1mxtiE+xsKfPp9jc6nDRufrWNmIhk9ZvE+lvU7XW3VY8WD+6ssXF
t/nzPm5RBDHssXk9uB6Ze7wPqIKkHyVLPoC8Ge1g2Q/I2s5n1i4O0WDJL6KgO2WjZzm2p/8+ueGp
xfvHSy4p18+eiSVmkTHli5LDPQ/PlpjJkhIBs8rJ1cEYcFwqaGfjWBgyCdCNs7dQqDS2RdZggEvA
S0712XqKtZuH3uKKT+Bg1zCWHNgGjvUWjkqjX9mHBsnxbaGoQMwURqLRfkw0oUACU6EXjzzGVslG
AEbhT8lracCFzVRxojgMliBLsm7zyoPRYNqiTinlndcRnAeZWpdTi8bm7LquJEvgIASg6qy8zNAJ
I/AbbWTbIvOSqZpkvOA0nYqhkUt62jsBPXuFZ5ZnmG7/jWSpcQTF5oExHYOOYygQBNHathP2pLaK
rSz3FTtDbI6NjOF4oK21WwV6qK/d2pPFElRXCg/hUzDic1B0aQ0Dsph9p4HFA/kxKv6htihMSEUF
wRBouTznkKHqrcdXJAQ4bCOOSzev31BOLUD1YfzySvfu6w5ERTGhy8nPRTbKu3EaoHSFj8Owv7XN
6XSeb0tttIPfz35C8Le9/Pv1XhIFSRYgRwy7fC9De1/HufL+XKBDKTfgcI2EeFyR44Q4KVwIXXy+
7HyLFOcre7fdqL4AWQjPDt3gOiruB6SMxFWakqzbOrx8/0xoj5l8DUGGWFJYZoD/CpW2sHX/YrZU
KU2s1NcOcV3qU1e/ZpdAN80obdv7dJ/mqnWEsCCoPrUaOWvxqEI7ITUGo8MrydgGaTVvmU2C+eMD
c1iMHQhyu5cqLJ1lgNEbV7Km2rWtwYMaycN9vVXghTj+R+BABop+OR9GNB6HfA10gd/Rq+EeVOMg
gYtxOqvMUDWlvthe6oTMJoUwmdjEY53aqvxZsR2TodjRZqS5buWPNmBDHbA/uuO13wZDPfq8OUbs
f1uNJNTJKQrWZljyqM7yQHtqh7NY+8Mx3ZOKAKHIukJ5vb2HWXjzlpLjxFnfb2NjrSC7TCmoOAqF
IvAqgEjKvFN4kn6SzJJmkaAgSU4GXZ4RRzejUDC+dxCauD2CxnQ9n+K6SZbwzLIm9QOf554t5tME
+38aOgQdsWWnGS1w0J5/Tjq6sNPsqKMS/QRYi16oEn8EKIwm/0ksY9cyA5JJkwiUHCJwRvTE9Kk9
nFOJvTi0l2oY74jfvMIGn5DxtP9lgrfncEwJ46q7N1xJlu1Ac6wflFUBaw6GnomATrACklBIFVz7
h6+/Y17V/EAxkZXitoZBmCpL/40cLxXzpg1hOc3iiL6Mbvx7BueDfeH74ReCYe6UEkuA86DTosZN
dq4HfNyezHmsiIVkVphxuragNjbV6XOnN+H1ROi6XxVkyo/nNI3mYX3FDQ9ZPNFD4HjNYzeMMfFZ
NHX+E2sFqiTEkISrIJNPzUseJYcOPsCAlyERPuBojurZUk5RMWWlF9SZtKFPfhPGsoy+0mA3b8F7
k09BEdWiWZ3iQA3obk1DPq6AO1cWfk7Tgpy5KSrqTfdnVO9FRHRECVUV3j0mHc6XQnScqQcHk3OI
QRj+c8IRSAsFa5neCugqILEfMMoONpbIqq8telbthfF912fScg1p2Quyt3aT7RUuGJJz3CZgvmVe
/u0prh3jcTYJOfbiwYqBJjASvMXr4rDzGQxejbCpOAl+hnapQ4Xu/qbkiiYyAidmIj2DEgLNp/PB
rXx+5MZOaYeAVzTOPaSZsdMJkw821YSrkrN2W+tyXZNgZbQDDKXO6T6adAwEaswkoADrpa8Sl0NI
yocmzGIz0RQdhjPOgSaOCtc9UhiLEWeW9pHXfYuVo6suzXPNb5vdu7mk64WBLj/UiqOBEIRwufXq
cn6idWwwdm9kiWa9DAdh9T3bRYSCBVjMJ+s+43REgfbChH3MTHF5aBdLghvohvWOLecCd83EbeSD
vE6scVm2huYiDRVuYzlxe0OOQ7YAlFYaXFMudHdAnfHfwHqBuNlO+niWAQ9HSLLqKoQwSrRYZSrD
4TZ8mYEsop2GGFwQof/xneg33hrjAsl5a2ZQzX4JELpFMajdD+4I+Gbgcl3sSj6z0rg972aECRAf
QRgDf8QVUMdMCJpgwzVg873SkEv0rhpNwD7aLBv1v/Sj7BVo+DMfJS+q+LP2U3aA6ycbTOh4ir8o
2O465GmMu2fRefjoTxVvCLAwK2/JmyxLXKhktEH4SK0TBrCBxtBUUkIoZwfdL4+mnPyEwQro6iW8
8+rLRUF+0dWMyzIa6fPfzYqVXwoUnQ21vp6JYblLw8xDHB2LDRGv/5w85+6+QMAIUGLRjLMjMqxR
6nPF61bU9ze7eRSAzhVUtnMncgXxzD/EdJOMFVX3mBbYRwOyvZoH4HJESmwa6RvqGbyBWNt3v+JO
jyGrpa+HeTWjDSN4ZWwL5ucrIdEl6Pq7l+QLchW1bkKseflylAheFqOPgp398gyNlIsr9HobnaB6
Z67fGD1rBe9manqBYCfxkdEWX2vf6VuDDHKOzrJVUrKHuAy8rM70nCuykEw/uA2tkSXG4n0WTxuV
6UEYpFxoX6EmJn46tYJCMjodz5O5j4jewOYFuRGNzjZmfaLw7LsrWZBc9DnseG/0z3O+PVYiB5tU
YwEngIJhKB8MfRtAJAY8WzQqrOh9mfBWH5GSpyt/yS5ALfnzTVvW6bkn5OlMELc+w0Rzki7yVUBi
3rdtNpVS6o/xJuxeXW7bLgNFbFJG7NzG4S2RcxFehGmQw/GuTPU9Lf72zE56HJFEeqvXLvySi8Ym
5BKy4JcI7NEbE63VN4NtGLEUpp5fbO3pG6LRYMcTezQh3vsVH/RwsO2mdNJ4bWyUz4hkQrwZfWBK
oKTEoFzZzQBWN3jJyOXSrt+jEvWrD0zMiQZkTlpPCarI7KYe8c6QTyN16mwG+aooUk9nPK32/XXI
JnNRT6hyRTpt0+70Q0T/IlCegT+ENVan0wCtygEyRpmFuY9sq4N17QDzkI7jH4/YZceyydMqtokv
eYyuwCA9s4AKosX2ufVoreH52uAE/C/o0YUT+PMjEpt72S9BkzWsxMq7cfnP8lBtazjZmRNkDA/F
ZmSq+d6pSvWUDF2rg6ZC2nlTuO2r9jlJe87RJE2yWRid62X4yc57D58FNJp1JDFxnzzn2UCRW8pe
9PJgpGffWPd1Gm6KRvlc0Z9ST3h2TkJLVr5BKMlZWI8nRkvzqfv8sKM4q1kfZTrmPBq18xGUEuIk
KRY6mQ2D2rutlccWA2VHsIwh8rck8UioD/2Rt+jtDdDVZg5u9oILEebBn5jWscC+Lgh3GPx/+N0H
mQOadR122drXljIkwbz17Ipdw502DcoDxFZw3W03ASNPkw4GExDIwtofx13DOKBdBdeGdDFbHf4H
Vd9wgDJSJQGYW0NBum4Mclr4vgnRFaMQTlipYuwW4kG7zXcOFIB7md0/oslhhDs17ar3p1k1JCWG
oTlhkjg3XzQSlIaX+rkwJscsN/Kt4Wp6toJ9sAQEACdCYgH11mzTRYqohOO2uivWI4HC0wgWMlog
VsVsoS1hrdu4dhdPmKnrTsUNiL+8WcMWJUkMHSozufPqV6h8CjIf8h4eWur9oPkh4MMA/PFzbTV+
qPWL4oo9QayZFhhnkjCUjzqXINt3hynjgDFsXdBq+CzWqhE4oa2lqexxO2ZKua05jCd5ezrCRp4P
XExmsoiXPKDpWOxUZCXl0++ZM3K4oZEV765DVskN+phoL05Olt1gW5rBkavRtyU6LZl4HdkJOAex
G+ewtw6uJRnaSepujoNPqm5XosFzHnICz9xqLaepSKrwrO1JMW75mP08JOZu6cKMYlCbxfN6qB04
H6cirKbXAHIyJerjUw6vD4qmgv9JksNzlSxiY5ifecNmDDrO+1iQnMlVL0zD4VH4iGTAaun5MnBc
jiXzErtJc2gtbhJQVeb8XZ+jVYO2RClcDlCG9az80x92SQ/pNVDuYPduvulfmFKRA2Oj+BDLHan/
vmZjw983kc4jreaAMKtkkAeNOFiLy1DYEaysMUcl51/m1ils5dMErY7YM0Ap/ghmLTe5CiIvqaGP
FVgEiGOeo6DsVsZmUQzjrIW7eqzDp4WefwslRLMkgnl248Z2G7LT5thjSGokWH4ERKiE3XqJmaBX
mcI5TwQatfbWnglEMN5YxXCOPGO6DhGi3jaXWzrLDRhgO8K+E0Yro6hfg8YfNSAgzdOiuMcD6BIz
NrbgCuFItoEOeg3PAKC5YPJMDU8m9T41K72urH+Q2BD5LckSJ3xTnIremZI0N/vx31Mh86yX4zjo
rApn5dh7pumFeDlzAbdB1UgAfhVI2IbYF/ZT2m+//XTnzdwHeOXCFBiBF6Cim77nkFgOP/QtPk22
VdjVWgJYSfVKauWz28UxPX74RsAfmpNXFN68wl+RYKwwyplNcwmYucimnLZbO3kdLC6WjtPU+Wef
S2b/ZkeVEouL75sfuDGLeqaDOOtrnEfq5Baq9h0YB3T6isv4b8TYwZg22ccYoRScRHIVHsEKdLm7
LpTY1YgzJVRj7+B4UieV1AvQ00TwHlxE4xQsyQghMljAFHJraOLktEN8qc7q364Ielp3461n4ggK
Xkxk7hoD17mGr7GfYiabCFt4/BOWYFsV4l5L53ZqtI0z1xfm3lLIEHfZMIcc7IQAqEGf9d8atD3q
enxeVAHOV3eK9wSwfNRG3CHFbPJ+4y6nPlALC2R3qyw5Nlm2IywufQbUwMQqfon8DOLpXvwEqaVv
kjscrRBilzeousPAc7Ewt2EIphoyb/Qh9o/DmK4pd5+vEqRbViuxFKnvtkQzM6lpIMF5Za6J18uX
HjJOi7Fy6EK6m4Wm487vkEN2Twgnthdmr+x0cmWNh2L2HKGOSo7CDaNE7ZHMrKGzYC+pzkOJkDWc
w/ULUB/QBCwptj7ImHgiCImJwItBzUoTIg2pSwi0TcvWLt1UwB09JtX1+S/h50gFxbZgvy8/8xOQ
7+wjVp8HAwqrmOjB8YEF1LHfJB64TYdak+IaOMPHCZG9lrzySAic0nfkQSyktKIQU4O4lV0S4IBi
O38/75CXmuyQkNXA56Z0LgiOUo1VCMgu/oT3p6DnHgLLPRMJPCSqMMlEcSM0ln8HPWqw1luZ8DVy
cIKil91R9i3nrO0WAiq8STJ9Ekik/QOWxoti7FWpxSf0022xpLf72zeLHNbaDe5U3dzMOwMFH25z
/LXGAinpWluamIn+aMtJtkTSeVs5okEqiJxynu1EhxB9G7jYqXlpKi62ZkTgUbtuSyoEDfY2N5gQ
JbNGttSG1KxtgvmBA4SpNkkk2On8wPEqNWPaJNRdWAnw7G/RxauEG794fzxV0bPad5SOup32IKAb
fAPJB5KSTSGKMBTOMHMLfzrX+V6slBewUP8S+1o4Kkf6qAIkTKY2zD/iQsqyzuX0vyzBShilrSrO
XwKyLMfIqFYrjvo/a4veEojHY06U12SAsS3hNiw4Es4xEA1+lV2b5kSjac3MwF46Dmaf5MNrTNiB
lnSettUqo9e0Bhm5DNETl9TvmF9DszFgQNU5sSwRO5jTciEmXlMfvAGOkqplVlxMsrKnDZipkIKO
vrt9OW1N96J4ro0H5slUNHOEs6CJcIHU7g7Behrs9hXCWl2z7iP4BXww93hq97pCHUCRY0Z6d3A0
6ImFxFrVFGAFCGPJyFe0vCaigMaMqDvpdUSoSL4bJRiPl2FLQAzPuMRb35zdue/4uTqhPoVf8dOW
UXj4vsMVpJ6W1zmh1+BPvxGITNRSiHR4afs0U8hrH+IRo3opB8VZBm4LfaTmCj492LMTmTxcFLaZ
5+IumUv9RrYXc3WwchG9qDwALMvD9bfBMuH88Iul62j0g42TeBTKYEJbvICXCMcpuY/g0pnkrEqZ
FpnretNM7nqxqd2SpQtml6f7u4lh1yAZLQxEucUzV2wqsmikgSBOehsHr9G6IqaVW5LQI4nAnsd0
z6k8axcJjHCcXia10QdXVgQsJGVHODQLcN9z0wb008LBdja7wBYuSKtTAyNCzAH8poqrXgYPAclD
/ZexLjASMTJg3VEgxDUC5tJP72QfYXxNKeaQVuG9wj1iQP6jwp9RC//nci0zhLcldkcSPur2dhgW
kJzZ18cgC9lg8syDg92X7ltb5Onc8Hsx83+k6NLsxqJrLufEUBK0IyVAcOoCjBzSphTv+uxn4h30
pCz+ZDX6JidROX3RIZyhWPK+MfrqR8S10RskBtD/odj1tGSXv60ogeE/4DONP1v1wwLdr3ULaJWy
FbA4Fs3YpjsB2CDep/ESkJMGJG7e++e9+vsVt5dPJRrynNuhwMeQ4SLuz91DrdeV816AmoNY8H51
jolyTiJCv/zoSx1D2OOaPIe1Wz30TMIH+GcLo18mH1DNoPMy6nqCkDggZRINgQuN3WJhEx/+WEMh
JZp0QYtW4r92kZ2LsTvqNNmuGV9XZ7b0+7N4kS3elq4FksGj4Ta1c1gfflgGkuoel+nKRUgrmMPS
ooH/VJMgNtPo0wvEYydt6eSfP4M2jonJDTk0Q7mhAMZZKpLIYGwvR2BlVzAjYAo+bjUCOTgKHcMz
LmFsjBW2g71kMwK0ZeNB45Kezu4cr5QPyUuqVwccEHywJJPv5oP6LRIohzJaTvKCkQhEid8xzsKN
Yc1Xvm0p+SDWic9yaW2tmYubz92aKRu8tlrHLuegBZEqUJ0Lp74IJcXMEDnCEotdbgJRnKLHlgZT
jFAZ6pt9dkVEB5VYoSap97sndYRcw0SWD2USwAWNhb7Gv7h5kgztwO0KumGszlRtOwOaO3FLZodJ
Cv+cifh7LR3LNpul1I6UBQKhTB/9W82Lnwx3P2UXPA7mplEn9tO2p0Z1wT0tRdPwrE0U2t6R7epz
C2PeVg4F44lRmGj659Yk8NVTb3UXYHpcv4lje4P9I5FVJxN9B4Rhn6Vu4ZnjCEIlgLqAyWZrNr/Y
O4COtA4WtpJcCn4PW9GaHRAhs6Mn2+1e/httv0mX8sRHyJLH5+NUa0x+mO6k9wfuOIaQwLc87l81
8dGvxj9y1OA8uIy9fQYpZNlMyG2dacJDYPR1WY5ZvKPMjRdlP5jB2vP1TZolIiKipu5Uab1KvtsM
lqiiMvjlIL30O2ST2YJETkfw1hYhq8S2io8ABLyUxpn9M+sq+9HmlRoFCDgzF2rZ/xrU13kD79zl
Np/gDF3bhBgpWOOGlWGjInU1m53HdUUMhrpe574TfM3UetpeXxZMgFlDUzf2z8wLSu+85sSzAzkA
Ng5sCV2Cc0XtL+DK1LPDIxlRdkuo7CBp/d6zwCdd6DDQfM8zYyNTqOd7v/0dSBHY0B4B0c+RlHB1
m8rHiNnEAOOUOQZUocgwsi5IlJtisjqaLBMlKA1ClZ/LVxBjkWov9/FTbzDzFmCuxSauoVrNCS/8
+GXHG8lmR83Qf8qXWXodoVewnqr3iU8sHjP2L9wMeq6EM1ekX+9jhc3n6VwyW04FEVdT5wlY6L1K
Vka1HJ/63UCwLxNdRh86UrZeVLVdbU4PGwQVJg1bvFSfGBzYPyuJK0tFxRJRFOCJXqnDTKx9gIw5
Ev4I4WTQFQiGBOVhh6pxq5Xfq9vnpQ1OH3nJegsLLU0eeF6/97kFE3HfZtRysf+03ZQ+wfiQPzWy
lLGMBaxNw0fEKyogCBFpojjs01aFMkG/a2qBF0MYzAM1Fj2cAFJWSM7v9CIfmz/fFfw95ACSHkGH
kq8CHdFKe61xRDggc+HlBe+9l2IHOQPkZYAROFlHTAjQQslc9PiFnoBVV9C7NSBI4DOPoQceg8mD
hCsXghEtKqMwM2OXxQyz+4Qc5gAIRu5/G0KFeKeWCuE2AR5d0pMHKvumJmJIk3tH8oRZFJO7QXxh
d1YS4BhEidtXm7UtycVIg1JhA6q+Y5mH3qKmeiLPyaptPXbJff1Vv5ViYqQx8Tzu607Rj27VYzyV
8RKOm2d0V6tUiLzG9ZTrLXsU7URsOgJNNZW9We8cgBSTOA6pfxIj/ntw5j/+aRs8na+msSLb7o8V
ElzfgSfVnuJZb9hahPaVL2Ds9LXaMJFrKlpC4rtKWpvsFlTZDdJNdZT3iDNqVs6KWycJ1IGfD6eF
Oct5aXsl1wV7H3AkMzGhc/eySnfrRejdHX1cGviRe8Yi+7/j5/pWChlJgO7TLMZBWw2AX5C5TsZ6
40u1C1HEPnuJyD0fdBL+p3AZyUyyiFLoRKInTsLPtJUvki7w9LCeZSQnX47FUkafog4kz836oajx
HIp5smpy00pRnKm3sLMAtHnXWescP+JD+fo1wKxi/zE7zYlcryCfCo6JNPrbSOKoVjnUwxLOiqFj
OISCbtnwooHbRBmLfN6tqrmnwl6eFBK5rQG+yiPfOXa52pgYxjQUsDjVnozNmb9AlDUF0vb19gSb
SOiitqnvdjsH17PdO5UXylExOg93N1aXnSm2rc73NjSwuHU9rnFx549kUeufNVV46r6LIXSRJvT0
BGXfCV1dY/w2VlmY5+DyhuHonjKWku2Nq3KqYCUXU8CzawU3kmTKCStwUuLk/GV9EYZcFmYBOVy6
bVim5q9X1plg8osyuF256yrU1lBskmJB0b8pVlURA8vqKoegoVbTQSSvAD+hSJUG1mPYnOuFcTpj
uOG48SOHAX5fmWGFvJNXVgIR6eMKJb/Ufwrs3kwacgxC9K7UTBKGRfdCT8UVAGaXjxZej+RfX1/E
mT1i0wnDYIfSAh4UKRM8CUlF2Y17l8ZPHCjjYLQRHkFKtGNwkcAkl6z5LJUB0E3bLy0S/g7+64al
q3QneffJ/nh50hL2qC22YGJVR1nujtRVCi0IFsLnYc3Hnya3qazAhkH9O0OATvZN16+MbuTLQRuU
y8LTqfVhQM1x/qqOfEgP44yDNYcktbFG9o6rmXrdFzTC5VMXNueVf1kmvVhUXoDJavp8y89XM1G0
GeGORuptsQSIXC3LkQRYdDZ9pxDgVDUdDBBCmPfM4Zh5y5JXTqUdiOFynA8pgh8IIkrVMcq/2pSZ
hYP7NF8Rqc8nCHvAZNmrUaRGnzrTS6JANvxM+nu8syTwGAcrBy/02QxXtEdMoUoqgz8kHGm6Puwd
aot3NAFWzfxWQ1OtHa0tsq1l+6TMAduD3T6aI9ds/E8MCbEUdAEmtviHhU8WB+9G+52YXfugoPpL
FEFKUy0XK71gsGMmvtgMCvgVGymx5Ymyk/S9PrtxGWURDGQZQKhgSuTHMlJyZi7WzSuheOW+3VKR
DdLKi9vmuCjR02d10i0c9g7RIJbSH7cqqsSVUP0e+WHEk5pJvbFeDMhJCgeaZEayQSDj67lO4QCk
mLQwKcjpNVObMBM7nPsPgrSohv5TzuCYSGcvv1xHWU5nJ7HUopanEnzXEe/uYX2Ih+OWTPX7Mt0Z
p6HLsP9lY9VZ974OgoaOBnslK69iilgYQSYyshJepo55A+7kk6wqqmQuT0O00slAayEtLroLx5B7
RyxKSJjzlCxk6G8dCVqmam3gldqaErs6Fx4rgDN0dd8KFvHbLjdfX2PMjihIBvj0Sc9jVnUixcNz
i4JrSLEG6FlqUz5xeDu/z+2bLh2IlDkBWJRBoIJcDbKOAJD2NwZVI0coIXaOLfFTvsP0+4eqyk3u
q0fSnG5UeWXE/GC2ikAm7X6ICGQLMsvm7p1NTfPzxoyPGIcZ9W4Zdgf0qP8YffGZGA1xL76jcpJT
LPn5wlINpXJH8kvgOJe6rfe6PcGKJw0/MF7gdjGcJ1AkJm0N0M8EtQYoTwGwThrFTv+qr0dVgauo
bnVetVx97uJqh8902HmkndPDvYZq3P/njvKtWVa/oqrcj1PWKhbQDt2FUlyEaziQUIGEXXZaq7pI
iAXBOqSyJ5oRk2+XOcA0LPy2U+snym0o7FwX2SOOnT+Kxl50fmZ85cGEVHBnMFSNvsciTJ5h0/oi
wXAeug/hZprkZnLjvWd5gQbjVaiPwBA32xE8w1TloWZG4MkE+OysJALDNzHAHPNi90V5Grxbapp3
6aXJpMItJKe/LjzJAp5jOHWCKfTiOK+9zl7Y9EVTRVM4REzO6fG9ZeVzkUByXj90PNLfEFcdTYe5
NKlCu7siH3MsYYwy+QT/zpje4J0Ofx+brXOXZUa26XczeIJK3BN9Kmu/gOS8/XBtECtX0VHD3NpS
711vl+7SvKhS5M+kLwEBVp++bSBK6wpNRN957M0FWI3JfM7K1AhCT1uMl3u0u7JQqOE4xU886VoF
p6lo5i8PgnRNqXXvwzmGYZZ19syspUjfzDYwl9PFvIGM6Pz377qzSYaUIm0i5Op29iwqs60Tba3v
DUHT5JHG3LDzREKzVs0flo+oXd018xfuJY+Xl1shciIjg4xvWae9akzaN8sX4n9F+6btobPPOjpp
7l8Nx0tyR28NCmNCcmQJlLwlWysNcSQlaUZ2hCk1ic3KIyTsif6z5BpkKgY/hW+NCZY4oZ7Bscf4
IZBOPKPfOaTSqV3rw8MM5So8+4avvrnjG11VCggFPpMVxYTSyn4vE0CwMtLStivusBdhOySsX91B
TPJcCigsXZc7yODtm3nU8L/qX6HTUcQvoIl0sL+0AUlvrQvycka9yAWeGX5NkBVG8f6WKefHBgCC
Oe54ga4LQ75AEIFa3MUow+txwmt0+A+H1/F32cAWjJ1lYLmCthotpsrTiD/f8QpKo5N2wZPPTJI8
lbFAWFiEzLmQ6hcEPWH3miU+sFyKVal/+r8dOAjm/lcH7q6E6/Drlqiq4C9XwA39Wby9rfjT5uwl
5EqjSYfQpigz3hgvB5zWJ+5y4STbxh8VX6R5mD3KgS18iSx7uTUuoPykKyu4S6He2947ypEpzYi5
nqZpS2cydKdZ1o1F645TiP02uWvGDiGjrzTZY7sfCaYQ2WAm04/m14jjiOSlGR3Iucv4UWkFYwjB
XUvLV7ZWWxja14Tx+EnDfJk8u/47FVEwDn7uYxXLIgiO6ttDvzvRf8MLYITuVOzs/pjgpOYzCiwo
GNdRb+UnKG8NCcsN44W7qO8BROy6F9tIM8u/txyIuAc1YJApsfZxVDV3EU/r8z9vfi7O4ACBV/CF
yq/+W59CWtWfHMjoNDs+TZnjV8dv0vHTE4tW2Q1eCxUdhK87DiC/HeTdZXYU0ByMi3/SA7zLxzVU
BGRIn/5mApShDtlx4a6KwvkoLAmJF6bWnZ74WFaq9jffbzYbpFwyLL34yH56OvP+SBsySPSh0u3V
1f/JfL+6hG/ZszuwH7Nzvhv4/Fr/3yMMNx5vL0nF/oo+FfG27/6f9oI+Ky82nq90tgJaSX5E95WB
D881k8MjpAa1EJ7UCOlVR2p+tvQQ9QPeYBp6PDdIivuPdvEipDKnaRXNMrVCRvwB7iuLp93enHhh
fmnmqNfk4nrDdYGP63Z6FfV+Ztx/kQT+Wpi0CL2iDDtSZW7W2YR36IqlmwAf9TjYmCyBNkI6bStU
3f8Sec4P8gn4o8vgUIN4xuLfEKCVquW+F0GxhUeK5NtJQDTp7+WFkGKY/6dJ1LCgx+EnMkNt8r1X
++evwzuZOzeZfIN6Pnnc7XUZYOE2i7CweKcQzHO5YNwhzR/K2vqqZJ2djTOS6t54aLBmL+KVA1Ff
2MV1A2D00URjvbXo4F5yVNN2fDpdnLMBDa55b6E4J1EoxF5tHRBD5Em/7qfspfFiPihYPtCVXoYZ
bXhVjLiYyaArSrVSG4TgJzDUu8fg/ngWedpi82vY4rbdpdItU3/SlZJjmI29zlMfeEkBPTdZ6uMG
XDtNUg4lRpCvLwJnGQaiZ+HAZ2IYP41q+wPmPoKUeSNjimNGRCIoxMB9eTJUMUgg2Afv2LcLsF6t
Szbo39wDoRaQQMzM0G+S2B2oijCca2R34wc9lqQqwcbhlvRSjQBmHs+KO0/SQzU3fchpl50XJnCn
515ArepFxmISlvA9UQDxlmCdd6MEtCEPhgqQgiC9Quvbr9NIbFzApud2MU2dHyydddhFkQnHcDUL
waY0aYytCLCC3J4dwWLZsRt/hBB4L7wg8Unuxo9YV9YUxDSpoHJoElvS6HN+/tBQtycQu0ODH/mL
p1NNv8k8RMW1TPlMTVfd6auZ4jBVqItQ8RZjLpcFnr5zMClghrr70EQwlxnSvqu3GS216m7gdMd3
NXCAuDCUrsNSp8sJfEL4pfv8a5lCcSXVPHVvs9aEYmRCg1XbX4jKz7g2tNZcpvMk5cUziMC1ryqi
28Wzb8+gM/U3omwOyCN9KelxB/eY/u4b8h52rIHEsy44LgDnQ7OAVehQXRONUZ5U0mQmgOZAIvwx
zFLJOiziEl3QEAcvgjwjF8maeDEwxWXyrez7u8oJ8bMH89oPJbciwnDRaTfx6Enk9JqUpm5Y8gfc
bJ7URuwLvninC6P22NOUoJE3/Zr+Htjp/wRkBdypCUIYsAdLMW9FNyrZs6Qcm/EI/wpzyUoe70TU
x9fb1R0r7edWFPmMT5U9EgtANZgfmAm69AnGuJhxhMfdQQm72gSCGXx+K3A8zTCCJt57v9Krl1+X
H2xOw/GIdi0M32vO0oA/neHfK/8fLZhkcokdAKQRJFV9HuOnkBDFZWMCsa+k+h8F22CP30sTheYZ
VIfgejoU8xE2prRUsNy/MT/eMW2tZLiL62g468IoB5Uvs74TLf678UadqhRUhtUXHRCNcdcmXrrO
f75d+kie/wMQaher2YSWWAFq0BcxHHiQJ52OY49IQOcSyne0WPxeJzwPpwxqXW45bEE6+i1im/OI
bVT1ZBS1Z3llrqNDdPiH8GJnXe11vnn8w+tmTGsFr60ORoAJsB20RqPxUN96nuKkeqT3MQll4uV/
wNyISvbVFdBY6ZnnvIs+7TokWSn7iybkRDeh7rJEZ32rmbzMKjSgZ3fgn5ibS4HHXCDtdTmTTMKD
+wEG8cTg9Z45OGhBlW7HVu9WEY7mf8SBk8kuKxQiTwWwu/oLeZXDfb/zz+JrbZDiK5a8Ps5sKbqI
XQngp8ym7uQRVqELntTR2titEUlnsitiQHHuz/GbHO7ftOIHPwOCW8dKgl0vJNZuji5J+wJw54bN
7EzjqY1iTfDsr9OgmqZbCH5KUgRVwkjWzqEg2DgdRMvF5WKQSKGkjJb+nXvNZYtkZUzL5clqmLon
YZNBrdbWgWTQsA39IiycPVIWYTCP68e38fYBXg7xlsRwT/W2fJRZENtfoyZswmTKyqmJ7A36jI0/
nilmW2MN4lmVVezyXIHEDMttMagOGPZZlv0Sn/nA7/j6ooaoIapWM7rvNhbb5LFiKit8aM8q+O9h
ICEhZnuMAoBq34jz8FFqBqMbHXF5O7Agz9ecWTNZF5FljZMQgAqFnKQvgAzHV1zWQCISmD9tyVtd
jemwD4E4RJugehMV6Bg2w97kXUbyycE92aXNmHUCX6n/Ys3YjglNU7BUroYldo8aGDaU/F1A5x7u
DbHv08Pxh52TXwZiOD3MR58v01AwhhiysWEfAGvsSNnF0E4Jy3AFCUiyqATZtaiww0yRBebYK2rF
O4BTX6suUkDpfEjCiXcYZN2LvaQn2WUtgl0TybRzl4VI25zm98Kst4jG9w33PaIjeF15MFVvKzbk
JmRX/epsCHGi0bYRAXtHXhTOfwAZyQe3ZJXfdX75caUysV4Ho4hNd0kJu+iMwkEjK7NO32oigdqa
Fv0dhe9qpjLJy40tEL0bfRWIiAtSzFkX/rfxUfvKROyv5fwgxEKarIAOX1LRZvM+T0URwAuftil1
Blux4fbQcjzJytcAe2P9sY3+MjzfQ5r69TmjMObpR5+fF22utDR5+vB/wUvoaLUBZuNr2S64wQ/q
lSvXDE2fIC/mq/hlsrMWmz9CUJWlP0hzzRGXcWTODSbW2ZMxiezuEiFhkmATdjs8fO8hIFyZkkXt
Mmls+DPqsoxgVB3nMqy8bZ/G0SjMFZ2BbNcNAgDNR6fBQeQzc2iNJHG84Niu5a/ejQu+8N/L0UwU
PqSOLnwtVI4ySzxaqgupvfbq20MULEjLXRqy2RGitenQMjZO8lAy9xoMbpaZfV0EQLfjdO56ut9z
foES2Zzx11XYqBDtjyM9PZSigQ6qxsESgXauKpRdsEBHyKmmdvAS8kmwHlhcPY/uPMHS+hJsdJwy
muPekCuNnX30YfWF17NwcP8XQ5wbvIiHGvecPh1gqNMJ3jmRjbT+lGoGlZJ/bx4UHHdMXbGdg2ti
RT929TdpxORhJJs/hyfjGQ0Yx3GYtw9+EPZG/T+AIgeXE7/GKBER5/anmTYITcjFQURylPYsebSp
RJICoVntx2BNftWxn6xTg2gd4P21gg4Q1Ztd8Y13Z5wmyaFoPlyi/6tKfmEAKzN6410Vl/Xh7OQb
QWYmTa4TD4Ih3eoQ2DAato8o0KNsPzR0KjJten8pljy9qdN3l0Wh0i4CTiSn7eKS0oFYAj97jc6n
e8Uw6nFGXN7c1uTF8JOB2XwhmRhL13vc1awufTvn5jQOzcNBob19Dcn/oD73M4pLnJ+JlrK5DEhN
5vboaSv91Lbu3iW3aHxQC7GtaRY5uQZj7UGLs2F9kqAHiNSXDFQj5rQAL9tQa3x1bTv/crIKpfyz
MPvDQ5hZA07oIA8BeWfAINYHmZnb0I/K2B8nQEeTIS63e/NZMOJyiBLzkf9YFxJMdKrPANW2J79/
ZPqhnhoN1lWUt0RYqMco0qw9JWZvUcWecCU4IlXGPN7z9vllx0iygjwfkaAkALO+9z8/d16kKbaL
2keqDH78j7SCgydScgZJc21F8e1pALMPmnBvAxzvIVyDkRKK/6ELA/dv6716Ku2wlkeLBk/24iUU
bQ/t3lGlyN/UwadxKgfl8tRmuJPCYZiawUXsgbWi10DLLQkxguH7NixWQJekGv2hNOktKExP1VPX
Yf3n4DOplpxVFXSP7F2gklR6cJSKk+LlGJBKdpHY4WkaaPXyWIL6Bkbh5F1z6qnt7z8dLizKVXdJ
7SE7hFY90fK/bxP7CDZL97VCo8VMbZdaju7lvwDqEhG1olRVOKm0YQZEk/Ij6EgaEAZCiR/Jm85w
RHKwUS3QQcdfvGKCMcoZiXc47vG1ney6ZIjA0jZEOWdhvKHmmcU5y80Nec2+w4irbny/sIhvNtbP
kL8pQkX5jLOtWEukJxD8c+iHWZqHX6CyUPExGE6YiuvNlNEX2bHX08JQ63z1Upc2vyrVYxrgDLTm
NTHpZp2+cMm8Jtlm8h0JP22QPazXB2/QqD/qjYZnDgMKWDnlPmFXsMsqqt9S976D4yb9S0OA4tF7
vV9L4Bou69UZ01jFD/obgYntpdKj/z0Vvv7tVh9fbOAonQ6wFP8p/t+e4KbFiwzPLXSWoeJrigRA
OJ6vCpDAZDOcw7pQJphA3kSp1S+T8Miud+X+ELfKKbOQ1Wu34vgjCPvoauAzr0cvIntLDnqvqd1m
eq9FtfjOmkTBIx4OWrN0GJWjrt0kr6yxg3oUbsgdtTZz2DZOY6qI8MCMmNpP6a21d8leCFEwrkW8
I3AiLObEM1/opqpSlj/FOtYXLpiLnPHxwG01eDbOIdj0mneTnaqNFJvwdm3SsRsYRva2SJPt56La
NfOqyCuTK9UuKBWE2aXThzNYgNYZLjBdNj1dW7oDAyZ08dcXDQ98GNUs4rDeZunj+zdGUCKN6TDQ
gpGHMNKZuVOw2UxP6NrSW9Zoz4FPdHNQm5iR9XUCcZmYLCgrmbVvowk3opweeFLOwhY3SZVXvkMq
UD7Pb6HlMimXCZhn1QwhvYJOomcMloEMWeAZjyCTar+LVeTTNbyQEAVY08VnFjr/06uYdei5x4q/
IhxcmbxhD7WFdoeWOhbo0c5LQ5VRYk/fXhpU05gYdBZ7Mrl9ZTatqV6mhLZbdTFvQEUafeorDk3G
eRxNRn/XyQwlB36EaytfFMywYaAIJb+pWuRA25LwIibbCvCwFT/X88Wx1tNvZFVWBMyHcaGbRYeg
wqiuHiYLd+TOPDyk/A7ZEEAkre+GNVdN+JJbsRBUCSLFg7aVeL+p4agiC4bddoSRgAWnKX2lqOpm
OaKT2fC2PTI1FekTABI6GwER8EAg1OwCQuuYtFqU7KORnwmdkvbryXXDS0xqQfzgLbqkVxQWQ6Ok
1JbidSe0oWQPdC/d5Nkj6W1T6FRywOW015zhxR2LI7OvtOB8oxTHAoQPCMEO7Yf7JKqusiOhz2FM
RB3ZnUD8+l2MtVfZ+sr8Rm+357QOQeJh26ziBH9qqMvB7ptKvhz5tv9uMrKd1iIdDlWiyhDv/jss
V+9W//Mpr+dluLtm1M+mCT1s16V1HfsbcYUsAaD1z/xs367MxYWDnWkvjTw07l6bNldkxhoJoHOo
6n6voKeZRz3wa9h5Qa1Jt2fmMHoWOFmV9HTFA8GKYOzE5TGHaWsbOxZ5elMttnv395Cy44YWlub8
tluKADqdZ4gBhAD2J7ASStiYUW1SajCtWox3pcEfbU2SWt7UD8s/jCILjCrAGzNsvqtSSPu3D07q
nVdMYgRQbqMt08uEyg871joa0kpLgrj3m0h8imxaXRluSfr9l+ufTeeSxwYPrqiXpka9Z/BZPi1u
GwPZaF4tZefgmF6/509mTMWhWxjPX6oQGxK/1EdAoIUEwlSp0mKRzRL23vbms6oTSamAqjEFaW3Y
VfaN3QDFT7RANMoknCmpJ7RFeKLWd5l7Zbf0IX1d8KI8ohNmLoz9QSNjVtqaPkicT3Gp+UVNQgOv
MV75YOu5ftq3Q9901HPnrYNTbs6OsjCi6YRAglUlIZOAjE0EtUlKsytEcGlybpa+p+chtZfkQKLB
B2MRTkrsUIejZs4xJ60hBShX5TE+tMcvgk++58ceD3pGalf4X80dTKbTKRQilvsz0yBjg7+D2f+F
JoyTc5wtCbYcDmOzW2ALP1ThdGze8BNR4w1C2SWP13nUM1WAJiBMbhM31HlbOIk3UZcfepLrNeVz
wm6eFJU8kx9ZG2aehz7v3awZ9flC4yoXqG0qSQV0+yd0o1+jdKobS7mxE4H+k/gombFeaWNtnQxR
uO+06CE6DRUn35PEdiKAq478ir2Wn58JpZ3KofGGjQ/A+gWkMc4bouKXQ42w6IE7PjKv+g7409Dq
K2oQN4gqXhYBUkvKDLJ6ZA9nWI/WxYjKvAuZHngT5oc5gJOcxYAZzVAGnNELALmzYwkHrvfbWomA
O5Ar8TqIfsoB/IZRkZ5tmP0A3QyMNsIa9ZJ4LOO1RWO8rZjoAl5mHoCr20AyGPDjWaVLZ0o4Uavv
l/kPYSBBuHELi0b/52iCxNGytoK0uXlkjvJzPWDTHK5QgBFyVcQx+JLTICozuVl6QpbnY5fow9J7
gvkkNiQDhqmGhrmbjXhUc7KY8OsOOtk3d0eizNilJnzLaPhGBRAQYLnAv/wBaJDTPi0KKdyJH7rQ
vwEZm+XeKjs6Mzs4Vd+G1WY1cg9f7wIQ4xF7VPsN03qDzHA65l508SbzqAeRTsnZZCBsCHu0xqop
jtp+u78hoJhN75RXmVqWfx5Gn7fIvI3HYIDI0h3aI+uw01MP9yuEZK36mEXU/XvKOxdRHBKC8V/b
NybpWpGh4ot4VJM2/Q4k6QjtvcsDZpdG6E6mMCinr+27a9fflFhiA9+k8RvNIWemeSNoZZrBWOp4
SyfdnlZRFw4Xt5ByFMt3wiuNdV2dHucFhAIIvluezgxXMYLIehMOdj9yYIAQwQBH1Za6cR87vIuz
vXOqY2JX4eGqntkJ1t/nCjYUzFlmXZwrTBlDQmZXIgJE9+LXexJWAoe4G5zsBOQ0gbN6bKunJtc9
vRpXBw/T/OwsXaS5EeUZtg+8CXjzPyvtnwvlOJ78ngPP46D/WUiA3VNSIpT3VvinS/urU+YA41kz
vqvnNnbkfT+eLOglOSgfOKZPGabfkS//IAwK7YHTqZbMvEe9EnMYVa07Eb2r4lbZ8RIC6DHlK+1V
D9A0mUzcGJQ9IqbM26sQyjrnCzEQyqg362K5QBpzVBP0hEBzuGxq4dmmcdCG2OdhCozhi5e95ESr
WKPksoiLKIndLOCzZ7yGI5NyLEanTtVH0COrUXRGOhgDKZbgV/7TE6QEMXBXnfLkw50Culeft0+O
Zr3vD2vZG+b1+cdxLq17BOsAdKOjYvjVHinDfLvPiQXQcI3bP8MzTHBj+PIfbGIfQ2jm/GTmX4lr
vtY9AS/ipp/7i3AdF/Sc5e3sof8QnHNwiAwZ2KQg4n8J++qWqvbRlW6Q3NGWjf5l1qzcXpjR1xr4
v3kJ40J5gEZAHNQwv1L9UlyiUvk2+Hn5FKV8RSJvWPFq1qmfXJ43S7sEpceG24eRx3gwW1HLYp57
IU43Q3WYhQh/HF7tN2+xMrclx65Ip18WQ5UmasSBmuKOFd6vb32nPQU6aV5ZDqFfSiUdr9kg5lu+
SmCtTZdqVPb9DlNTSp+xJo2Gj5/nmuXZbZinXIqHd4yUiENdP7nkrNsGV2gIxA44AHuygD2LFl4m
Sl3YbES+dB1TArsqKMdFbgGTDIV3iqBbDQIPRG8V7eR8yGDlIFSrsYukVOFClDxWfO1h/c/3H9lv
IhVH9yElDP3FLhO/nskbW7e/T6PyJiyklFSALJUbuCQ8q25qnTeixl0w+BB5gjELc+rBdtcMl+/T
Quh2Ls8fIdvqHRT9Xk7ZOdizZo3TdWKl0hgKERUojT6if/msMueFNu/g94OpStGLmGTiIsF2Tm/x
nVq6+eSJVt3G/EmBRFlSHhCjIozPHd/Rvd0oQZPrkuBlB22MGG8HrX6U27+MgZxMH6y0FgiPyTuN
//ErD3ECb3YQ5/vDztJgd6bQRacwA5EBIZSjP2jypRWV25KygSx17vzdkRqG6wr8IycDzO8j733m
XBZlRq3AfiUlhQf5B3e+2rTu28D5cBI3VM5d54KisFZkJbrpYuJAhtjNV6ur5ETQ9uE7wQ2thInh
vH02/qsYAiZBPNwCMKUXqN8CQAPlF33NQ5CguFJsdmSAgvu2iiQ1GNWn5UVHSmFv80BXsM/1NrgY
KJQwonotwZbnkrrrL1Sq35eJ3k4DAK+AQIJlhC1gXh0nChMIJVia0kOQTo4k0qkj6KHrDGJoX2Tr
6E7JxlxIvydN7JDEZ2dNH1npnzObns7iVmNnf7NMygoAmmXt2tQjsspWdD5wB0poVEvZKqTMdCT1
F4ok+6uGoVVwjRJ4/NIU9ijfHLJ6w3VOCEcnISUjtaDHSIuMoCxtvYzIUiNqyt0wHX4TOPFEB9il
yPb8Q/00nnMNwwpeFO9ZY2fvIBcsJprw2licC37mfLnHht4+HYYSIRB9IETTFw2W8aiQ7hfmY+NB
7q9kzeYomGv50WiNN/zy3H+VGnW2Zf8DyYjvsL5UHy9vxSAr2ygrA/NrL+LVzHF/CayAf2FbgR+t
dFlHLzn+W3xNwSYpPF3PZCf3ralWneKypxnbNToXwiRqwK2nBkNRfBO5KRpj6XHChy7QoLpye6fG
eb5c5ZDv4NEZEdxyaPy1AxKOmdeiS8dN85s89eYEQzq0PUKH9rkUZ94PEVFmLzstgCrBbcuzLI2L
zOrJ8y4uAAJb3dAj31csNj3BDyXQMKc/9PJI2mp/u20awNajx/DJfJ6alXdq3IWtvwuKw37VF6V3
10Sz9TKKHuGk/+nTkUrdclvN95pbZvrMLsunuG1XeLgNz298wVV0IbkzBSfWwSIKn3XqXq/dXV+x
fTUwA3Wsnfd1GwZXfsu5LuK/6OoBkbrt9YGfiizwIZMUB3ctQbTkmOddnIkdyZPYwOrUH9YWX1+i
8lGLQ9II7VLr1eKEtnj60KcxIzSiS1MKFRe7uMBaBAzKGxSvg5fynSqfadLe4nL3fuAYwEAo0zhd
OInDzJ0rR4RC0vx/wV9DZh5sYpROI9facaN22nK7qFnwvUA82N4VTHwcKEB/RNUKC/1HVMj9CtZl
GCsI+OMyQoObr4oi4nEVmmW5194r254QV9oF5KN6/xAWN1Kpcp6Yst8+siJKbm8DEQGsetlQ1Y8C
9jSQArSAk4RLWupibIK6u7FiDxDUxouym++S6eRD7MGBKYQdIraR8Bz9npsDAzDo/NkCODCDibW7
f5BEKWdbH5otWZCN2qiwCjaVDeMXTZtktOXf/E0BlVry3i7oq4DzgdqD7z9kOA1BvYf8aDsyiT8z
EOAzW6VgGUqtETZusLFnsQPs2k/hhgb7y2CK4nuJPxyVamIMf1TZl4A2RV+zZrYCk5N5K09vEjJx
6E7svsTZ70BNisHu99csigwkEo0g8slfrgJzVk0jlJC1NPkblusc0LRsUXsUGiwbP6z55yg5j4Lr
phWjxCFxc3xPSTV5U8RGu1Nq8n9pyyY01P6HH8C31FZ6dhKqR7M4+3b1RtPIHEAGFDDped8J/VdM
OPqPUSpVBs0zxVyDi+o+UYJJZ6GGyUieK8REVhiz5hYXw4CpTxtdDXlzuWAcIPAxdIhXzlZ1loBT
dawnKv/c0e5hCOwqalOlVWdc29NOBchTNq0n6sZuHlNs6mcfIDixMQxjKqKuO9mWkrnvnPLSDzc2
0ZFY+xew27r2V5w/H3yG81/RjhZEgGmGlfMIc8mfw2EwyCnHGRx8J3+YBbzl44JbM6mm6zPRE4d8
2rrwXDbhN5PcSIDb+FH+y0f0owy9iXhGSqzRg/oKTslLbp1I9AFu/K/nWqdkejKfcSeGMVcveE/7
VHZynAsv+WqYWcOdCoGSBpY3h0VmYXfeYUIw50u6CzlfRTrv3197Ot7wXwUr5XOPKKoYDErQcaL2
HNb7TSorHdNMieDqNh6fktg7yKrqxbqImTFGq9kXB6+USzcuMpqzC5aPmcszFJq9IK7Y10EUbELM
FAgbeFbtAdRjO0aGVXidak5dEi1WqmzazXv5sutw2CLK83KSjSsrtd1idwxQ/ZODnwajY7GYVAKJ
g9Nxyc+9EtZC+jZMOCWFj1LKFEwYBmtxZG7yN189DQ4zTmJ8F6KyX/SwpSoiVLJNfqVXoFA5pqOd
f1EyljnsjREyjVitBeRbXcC3XzMBqimRVXrMiEjGsaOnBfQ6kr8TmlCK6yZY5o3Vnfb3109cNack
3ujdlrQ7PmbWTiUjht9BAeN0iBPb/Wsp0WRFb8wbo+S/9fkluJRd5iitmGN9eQaEbCpE2FpcLIar
8in221UooQbOXOBjv4SQGkg0IPWOmD1mdj7VUJ1tgBlNUEyZxX7Jy2dF7xikuHXK9sFWqdOwXxpV
AtRsBHBVrKSKuzIX3OQUGi0i9q8C0J3TF9QAXJb6D3+PKWMvWuHlrktp+15FdHI4g6J15ERt5c/5
hlFMOmW3VkV4g1wIIfJU2JS45uHqAv/sWbtLaYeV/nVKg+I3TtOjIwW1baLqPrM3GWk0cuz/B8+I
IpwR538HcolWUpioQcnMY2Cz+Rb99WHiIuMV8KD1VUjXPXJ1BSNbgTYhJmJ0Xu7DzRSp98trx+IU
7/IBq9K9EvNBx3kzCp0/zqtF3F4Rr5ayqTgJD3JzSxGnTlACleS10FAxDifeEODJAPbrVywsIJ8E
CaN4VaIg7S4Br8fAdIsSRvN8vFFK9opKtFW9Uyic0AJsP8C5xx+XHVr+DE5SdLp+kzNR/EQGmcM4
Qf6juIENJ9vLIB9alNikUmos7vPfAcIZ7e8sIOZZH7nCh+KoK7JtmDU2a7DwDsvx/1VkAHrSh/vN
cPppT1BZgaDAHEY8Dbd2m6EARRUU4z7jeHz6S9/dFhIRWTccNaJsIJEJBKhY0ek20vOyznjp1UPu
kcsfQmAj7dZY9vid3q/98vambc2rylJiQvqbitEPs/Qk3J6BfIVH7o+AWp8CssVG8EBgo/+6435P
HNOjro3gFEShmCyXTHrSJPu8Q1SttfiC252sbThEJi95oCBIEgeSfEWzMGwD7evMlSEaaALxak1J
OezbcQU3WBxH/zCfqpUS0fNVNFb8rSEhpOljCRL29l/icOgzaZ287crGN8ZWj6ejc/CIGULFSBK5
ewHoKA1CMCSxN6cIabFzdAAqK8Hmb712opd7tpJkWnp2dnJVp9ESpjrXTwl7PYaj7Wdjx/z0RJBN
QaovyIa8Itn8s3H+rBP25fod2Ag9L6RGSyUc+atnH55R3isOMFxyEVJJvy0dVIPD4tJYxcKEVm6e
y4DyzJk3iSNpivgLPQdStbOjrzePkvuIMFGCNYUi+9YoXEFtXC5DXRk6Nz7W+i3xyjNSzQYg9+e0
0nLalu0K2vpWSp8XurT/H68UlMhrouHezrHOZbL6pIU4ugwoWq3LNlYMD4sWsgq1ORnUxgT0YbJc
lrvxCndbF0kToAeElteNB7tnm79h2meotQvY09NzLPTL0TIHQRUpwO7XW3EQmQneaRbfvZ73Ypka
Rw37J7F+GHTSsRSLATFFU57ivcf5plfoiieCFEZQz3+muDbdI4ZSl4qVK3fBiBJliPfn69MOOKOh
+Ax+K7alFUFUtzMqcu+kPv+L0h/xJFDszIWHKFCKREbvqAY0fehphm051R67CsUCHHtf89wxzbEm
vbTE+vXQE+JkKRLrRm68odYH7rrqF1A7q/rZXoFAjh6B5HgJq9s/bLkJ/gNCM7fCgT2SZ84Y+X2G
K8C0MxjZdlwgrHrCFafGdHo+eaKfpZsgmicVh+oqWrHyISGNLgPhxxuytYmhe5fIdZaWyKrVnghZ
/lu7nKJNzaPSTKDWHw4aGoNSJXieYpP9NqLG4YWISQklNRCk8dZ2olsE2eqnTy94ChLYviuGPjxZ
5ja4xzAJPJzoO8khVX77H4MlEps5fwwFS0hVARrOLEP+Pxjl7pRfDMGW4YGVmyghf0XFHFWXomif
ykA/L/Y4PIhQjoh2q0JE73+KumuB11MCb3UScUbSrvZhgw3968A7l78raBLR/8xkcuDQwTrDmJyO
YUe9QR3Ex+vp4tvu1czhLWTv66z/Kjzz7pVeG3//po9YfFLqrzxgCDHYSg4KQEOM/Zuiw/Of0Bjb
xkSkofdCSaWh3T09P92DrzjCr0C4jw2COJspOYml+wOcWPdAIaYhPe/LCJIgOw/WW14GeA1O5OUY
UMmi9GOCHzTae3Ctqv6E5gZKpuBDsIy32dTsjRP24wUKqQ7Ol5ORwCBPZxNTpKuK4GYFqo3243O2
a6lSjzgDUa0ufBpzdPwIt8fDVgygPoM5A7EMrRSLmggopP0WGT/wqivV8Ak8z0TWlFk7sPvcrhSN
ybZybFiOfU9HpNu4Gb+lv6O5xUqobnPVCly62QYrZl7RKYGnaBGqsCzZQQaKLq+NX/RlvdVNBJw0
PrfPnyM08Lb+Uf+YQHFOTDac5GUcv6adwpDc3QTMYjyEhmoMDF5bFgJ9e/7WBLa/uNl9O+6sMIvs
5/k3/KQPi3fNH7P6FMKx2lQFB/sUSBo1pqxcAReqrT/zbFaD2bfG7QeqvYeDUazzpcsl1oLC0jxU
+iCv7zkPYXlKLVOb1kw+X/tM/4x0WH+LpwL61lQCj54uy+I+j5mb+jSjW6uy6sy79b4rAGDDVbYh
mev8zNq60hgzRAxtHfDcleEoURqhFd45HQcaSMVGu5c1RbiSI8EjfRyZLYd+GVOu0l74Txf+aWnq
427kPj0Brp2IHckEShmgWIK/N5eON399n7C6DsGGNtYzgXEqCGNfA5RhnKGk0p0U2leuGhlMfzY6
9t7pBXMhJz3YdHBUiY4Ikv0xKxECtZ2Q7dwQpvD4bXB2YTc7KzmMJi0eB3nGM98VUirzDr5wFP0z
bukaYIaLAg1FxF9mxnGqGrat3A0fAclwBoyNbXDHAzPVKI9kzik4ruh+BnuUnw6tiQo13FlWZqGw
b9UtWDMyNhdGKc33fsEyWbhXNvC+QUoHteRN2/vc9jZo4JcgpxPXZMS6kAt9DkVBojK+9FFGHx7v
hqLv9Da3quc6yWAHbiMjpg07lqXoYnu9ucvQLc8FGNieWvVLYPxtMHQiTcjA4IsH2KXCWpmjrTrE
t6lH36cskdz+lZvWsElOyyTlkrfvT+h/IqlVme+IZsi3DMs6KoqcpaQit5flCT9D0prJguvJNhP8
gzQ6SEVuXNDd3ywhStZDFKgDVB4+rEPv8irPapuNZ2aD5S/Ti/WsM4oCxwnz//Uo66+3yY46SzqP
fEeZWpkoWtSgxuRZnqIMegXvckIxegp9dn79iaSc4fC95v5NBvhhkVoeUDrVJNn2hTfuxI/RTiCt
Ird+5sPEoNhGnyLQAhMOay8yXeO7prGy2sMrwsiwmfy6U+jRzvCzivnlsy/KUifEfZ3/86fGIarn
MYRDNxMpG/O5ZrHZL9cetvMl5m/q8tf7GB2uBz4D/ZMoUMothWhiK2AE8Rbi+8oL9DefyZBQDLkF
UYn9E2xZ8+hrUKXG7s7sm1CKDdBHYinfguGqJ6yGdbVY73vI/jFl2QBaIBlcVIxnGyagJELHecTZ
f/33kimX3igygFS8smi63RtB49Xsuv0GJfay2bGrWDD2u5Gu/HMwNa0ydhDPMSsjTD1f70iq0Cqa
cItCWltUv1PVyIioIHce5YPH5Zq4Zz64h1+mfO3Vj6GJHze6QB++c0xsQsz9eFZN9xTtLh9K6v2M
jR4rScNOaZB7VRtY78f6VDDG/NgjglenXhT498U1jmRAQbEmo/nja9h4ynjB7KXqlfqqmbIW+93X
LHBdz/cTuYgoNwLoDw+y4Of5FFv+7rsi5/RoivPArCPE1as/QcYLw93cWnDDj1kcFJyoN4R3JsrO
sOV8IUyWWN0x6mBz9K7o8mT01SMu9Wd6zXkrHBgucc9IFKs8QssZFo9WNhPPrQt9NALCsP9QDdGX
V8RB9xEoM7uXfSDVikXCR66Zzp25wuM5FPcayt/vF+Ts+dai4oskNJqRtFAp6BKEgbLobyXhAs3z
rOaHWWz9CgqiP9Hba1hH0FrfcuJxQxL+T+MRs32Yy3Xhe5eEyvALhwsg1Pzvar/1i3NtgwS74grP
tO0Qnq4WGTn3vNZb5+l4iVAkDZTWOwThaGpt1i3pxUzUC5MnKiUmmgvlR48xAPVoyAsw/2CvEvL+
c+mg6d9B+Q3/mKwiiRKWPI/SHY0/OtdFUMhh/l6fbGddpG4/w2AY8UC628zOXE9U6v388gXR/KJd
N8arcWJM+KhwGUMW2xmSELC8kaer45cYqPAJCKo2xIz/dFnFE/qMQG8zIMtOM3Gw5bUcBHWm9ejZ
0pVs+tJi5MIECz2MoeDKVBz/bTamerVqYo+R1469c9YM9yoVvXW4dvK5ugUe9T6dpf2eTisExwYU
TFZh0eT787PdE2TmRIUEKlvgZy8juWWcxwOdoVAyaigqO9lB388liMx7jPdXy1RZck7jI79Bb8yr
wB3DmvTq+BpwKMa8Fzhw5OoBisZco5x26iJTW9OtzPsn4vvV2lbBF4eYMqvQN8IzuoriAIOBMR3Q
o+Z2Gap4dZIXMWUiEofnFWqEXehoGh7+qbx+6bu7iQsiLv9Zp8zmKD5zhPZYqQyBkDBmtJeg1yFC
8aDubXgp23vO8c4uHUudV7ebHVIPuEeSYFeYTS2C6bCMd6hQDAocsHVcVUVnhy4TD2mrXUcLnLdh
Vq4NNxK0pWJQO/QP7VbREJl06LXKhq6Knop+rYml4APc+CPXBMOgeTiJpKA5FAkLQxSI8wmk1B/Q
Tj3apshTInvi1LxAzYccd5+vEIqG18T8MHxTlN+IVBBYkOBcNevbDORy8YGoI7HGv7dtwGP8F2O3
Wj3Ohl+RKehuwoK6KlOTu8GX8TOnrfpgXZxGVjhJJZfYHd5b2p1L6urDECU3hbQ2CRnG9OyzFIrh
TBMYNcMgQRysaEYPo3VqAwnY5y7U2Etnk8BVOo3NVi/K2h+rcFN+AyrVKbxsrNZv15stH61PJ01y
oQx0ffJOO3uhjLrzYt9KRs9ObxlBIo9v5S/D2CQhHwQenSsSW54J/eey7/lavkp+nahD+PD/wt8I
Jfkr+S1UKVC2C2U3gw0W9hx3v+HtWnhcnEQOU35L/NDNRyNLWAICZqVn7ATZlg1Nafwv8Om7do8L
qw1pKMsbWiOMkYmeUxDAfGBXWqUXBzaiCjjR8/OAXEcIlqDcc+8iweHUsATWemKp7LDxpbpcXLj6
RnxkSCSsaaVxteyIroelfADMHa0HHFCmR78boKrbqpZ1ioCiYCYj1R6WDtIE8QXaLCQKFqCKP8va
enPS9e96Xv5I9CaamVFsU/Gag2x2x+IlLpXtfNhDyGga1aMkK1wC98M5DuQN6BlImy3nUProzT1F
VSyIalmOxUw3hc/dGuu2ei9Vnm6iNhSObWn6ek5YTCHcEi5dC4aSLh+Je9SYZymLK8WfztcnjDUa
68X778D8DHGvH7DaQwIJAHwKKbJr0I5dADZpDeAuQpdBmkYvOKlhfB9IxNgiwmP+Tz2TVQtTp7Bi
0hSoVXt9WM273UnJebizdRgKnukTkJEmURoQXHLR9alTu+jDwyMAmd3B/uILEWKTT90z2adE8Hm5
1sMg+TGTeumMrNko4oON4bHufx4RLXBbEpVErZ3V8IUHOvfzyGDAc4fS6nc08Xwym66LFgTDiDL0
crKyP6Zl+3baLTJtVLJReKeWbF7bg1as2blceEdL+1RiwNlB/OKEFmYFlmZkyIJa/n20+rBvd8El
AYaZWi35axwuXp+yUhoYH1Fq2RE1nXjWOIobcf3m8IAQ3M9kpz69ZucMfFfd6ROEY6z38R92Ns+Z
0j2YwkU1UjIbcvJl9iMiz98Qw3mxn3JRdM8QTH8e9Kka4HSgP9mfXfwZPdPfYjP88WxfcbBz2bPZ
tsw6Jt9J5i0hLCRpUnVV1lhApS1BxSnINbrQ0b3KRtQUU7w3ooNghZ/NedI0cNaAuoQViAyui8q8
Ejf8BE13LgsD7bE6g9KyVE5zNYvI0fl8LNdQsL/EmGMWMSyt1f7LTJKCtKmmbgUWqDjFeROpYgdX
GkteWPlJcsEPxgi68o0kp6r4SjA14FiBPWfyDaHJ/SnrgrHYgA5EBYnKNyICcC19e0xDyCGNnTOC
1ez78682/s6X7izF24DwDVYOL8H+uAzjHhfUmktkK9d3gdTdeEBycLeJBRwI/aqVuGiumP5MQi84
/rNdr48Khk2yMhZYtLAMwlFg/5Z6lNA7u3RKbNxuTxvBYTMOaeE/5wKw+qlge4GiVaPb4nikwglB
R45pX/HXOQ1akqRmEyzSKZ/KNn2wYjgETHgVLez+EUG9Yq8ZNn6Wye7sJfBtyiUDcIp5J7ktaZgE
9dh3nzbI/KkW+dsjZgG4EbcDqdNBzHSP9p65vpgbUCg8dmSAkmWQ3jZWIrimvhrulUV24BsZiocc
fRvHK93LzoGKWobTUCmLTbQtIFxgAcN4uL90AjYgwL5sT0IxU08ohO93RTLzjKJLuZeD1Q+wYHQF
bah+ujQkTKe1M2JrmoNuOFH2QOQxzzxfRRbRSHABEwNq8IV1Rd8v3NlRqI8MgCkO/++3YrYfhd/T
HZY6Tswc7bFErWoYKg2n6JDIZuMYdWHipkkTjlaD5BTkl3g2CIgfUY56WeCTQrTgy37826z5yanr
Pa2GZv7oHwABNnUI/PCKNohJxmJjdOPN7T2EdStIEWWBxJCMJZv2SVP+6UuXq3BRgcZFstO7MA1B
16mQ/Prn8nzBfPR0YAzjrPDBdeo3BdTED0zJmnWgos7N7FH0/wAjQpY/aKasycFoh4WTGAuXerJu
ogHcWMATQ0sBpWS15HAtJNlZI1S4fNS43iVvW0xkElnemzsNKTe5tzTXZKydvE23B1KBGWgt/cGD
UE9ZYb4N308tc1yoA9iEbAX/XzEEcebgpTuS8ZmQZU+y3pkiUXmphx4HBdwPB0EZPFLSXuxfanbO
C4PKR1rvD3QzY4BzRUHoeBZvSMSszc03aH6fJ1B2SJkCtTvQs/vgt97Hb1OoMzEQLmo+BOQ7uc8M
GK5Hu3aJdOCjxSh59uvivskdHfFEY2guxuNjtkHbzVCVrRBmcVIk3yeaGbfgs6fKbhejTPuNR1Ch
OEK+sPSjqNSuI8aiTnoD7oJBjYN9hVr3gUzbBDHLks1sqN5nNJfTx5ri8lpPTCboPsXiC42wZ9bN
GJChk+uToCdWT6CManIo7uKfRAO/WC7R7dAVVXf/RWASr9393x+JLyCO+1Hi7q34Ix01Ir05mNI+
HSbGG35stlXaZE6N1RIXL65AYYFAseD9zmJSvt+lxAz03drqDbIvnkFrR77HTn031qIRGZSTJPo1
vpfqEtDgxysjr+U7kqGdD1yVUT8tjqbRP8bxhzkl/ljU1r1T1R6eFIhS5IXcLK+j/ARF9TfpR+XQ
42Pe9sjKve80zNbgSvKLo8flInCpqcd3vX2vt4xm2jDBSD25v+5Q+7oYZi8vnWA6U0ZWEO7SF6qg
PaDU/mMBrqukVU0gA3H3rJwLxiiZSVlsAMrQRrR/JEdK8vDU2xtD102573Tezje7KyldaxSrtb2x
2s5FCfiX8sM5+mVEkWCgtdL6Y7oRLOlgyDgpjGwkNshIrKrbAOZXez2gycS8M7vqHXrtLLYCsAvO
w0e3X7owH2Zomj1WYiNljCDg68+w7TDK9ttVss/AR4r5c9yGzrMdX/4vTTPQR2ZgTWydPB6cncVI
BO1PFsXdfE7szovF6V8OEY3QvsAQCwf5KgPArqFF7SKlkbiu2hN1vkZ1iajr/CXWnw9yljs0EreY
KdzG0Ywd7UDHhA7lmvyVmrPDkwlyY1rV5tcRK2vm1WXd3NGRwa30vydJ8nSptDmmsZUiiSwUdqFC
etb2WwnlddLHTxmteAdF4UBzvUeiU6+/h6EiGtCThXYM3qKh64Uom3tntuqlgY+Ks50ycmEr5Jzj
UHLycLn35kiG+TazmBP1ADqa039TCtnFltwRw9IslvRVYjuAVL4+kDfNXYzyhdzUP2/ep+bWAk3A
Z59Y6LaLGXWjkTxXeOo360WJ2yFirz43BrdLQcXiESHHUQIMceUEvJ2ezU0r6eDklKMITwcyHUTQ
l8lvjwNePqfmi5KdIlAvn9yqAHprSlOZLtOET1/WDMSCQ6EWCXrh4n+13Darp35tzWvtvdCkxO/Q
SzLm8gnj5hzxJwfKdTcSDrnxhRom+867XWy7jkVljTaT5gpY8M+KfUY/M2NBaTds93P7kcs8scZ8
4B3/Aeg5GtpeW7ebX1NvtX4E8ShAySNBF0fri4dtRCMSDqcB1hGrogDHtUqh9JgFh6p5haxmo+Sw
6/gy4sxlLXSI1L9w9N0qwsL6yxmDmgPJK4R/Tr7s0Y03Hc0POqyzyBm8cw0y5+DvipMhDkSMlknG
sQHvLPBWju+K5HNkDJ4T24aKYDhmDoFDMtjTL7A+78MVZ1Qctdzt5vQu7RbDfjdPUg2ZoPzmtQDp
gqwky7zLSRLmnUnalJCzJ1SnramkVpdN0PvufPpF2cZmlflwEQor0EE3NZNLdskWo8T74aPDYJZk
th2ZilFf2U84AFUMMPoBPjdKayY+0IcTAcnEP/CA+e/U2XLlu5b2a4infgAGBMmK/SZkMq3oWO9Y
pGycTcQC4BGvoUgQaWQUCjJSQw5hwZi8q4N4GVu0lvcYUNdWp5xOx9w3M3q69TvmO1ONvOLRJact
cvUuJ+D5SfaIy1QgF6qbo2PZKNrLH5jzm1/seOheUYP22Ob+9mNtdUUHzTsBJWIUGeD0YcAvs6W4
2dWu5lsu9Y1zqZSAfiTVk/z+pKqKi232fGZCN+cOvoog+6f4ow0TQ82EYj4fIiioly1DRDj8jjRI
mnJw8RXdPBjLp7zb1SL8zxOLbro0w1xqMbSFcha+SWw38snixPylYQPbiv/JO/Ci8wqBACWOXxVD
0P0hLe9M6jgdmy8Ngm2SRUJ03R/wIR3vpmaKUeLpDLRnT3qI/HbvdlemcPF0tKw0I1rm4KBoRXOt
TjQBjAV6ih17Z3pJ1eAhp48zEtR9ws/aR/4lvAdYTT2zlg+P+nTDVZKrKAGXo1H0W6isL33hP2Ps
vt0Ns9Mvhz0IcgnJYM99vV6FDlxxhyKRxHhGCWadrJBr5UfwiH/narin7V1Y06z86H3u+xo3RwNu
0MgYHjiG0A0oHW9yOZTzTI4UcB41Jj9xSltWW5cxd9dZ8FzaxfEu5gmAqfcpZSLu6O8NSQLqAGOY
045kDkMSPtxOvH5t6soVk/SNDC4X1laXeCSYOWQoP7HATamZoMD5zisJcAYGYocmQ6HwP+tWSVig
boNq4QHKrEf+Ve50JcG19xZF1A0k6P61YhUTGiUoDe7m98KFvh7T8Ys0xHLUUa0WjP/Xuua5tgle
BGJR5Gs5OgonK1KrkOlte90HjOGVPqOJA5kgIWiYdnGhm56opcmGF/OjumdDjiTiyq4LPW1cwxYD
lf0mCgg4ZAXDAadwI4wuefssjOe17+ZIDXwRnnXogWeuTG1l2GGMLB9EencPuayeesKl9PlLNTeR
I/FckfluUTJ+t3qPV3VMkqfeHi5wlUnEZmMfsR7hbqdAYf+xBeOz5+LbtzgOBsUBo1r72+qUR++p
HFQCrm7yBp/REmDD/D/iUCe2ScNwqxvzxeTNBC9BLE4uMn++mA+CHGuNSmBSuZvGSkNheRmsDaY6
ovL6RY8lzLMYqm8DXxskhkHksc6kxQcrF0BSI8ZzLaQ/JEyL1E/j6MaN9LiDwliX52PMq4pp8ZcB
HeOK+/+0vvj/x+/A5vtrIRaEjOM6PHMkoKg62IZ8geK65fE4kOUfuW7AWBW1JWOvV8PgPfefKoM9
ItxCsiPdCqgVEHr6P6RIWzY/D5rhuR88pj5oXdS9m6d/F2MRbjLWEdQBHy+w9CA9bzactamSmFYv
0MUBvn+cq1zrsaOpDucqe4WvF3Pkbq2ed/mQE+eqqX8DjZeRaDK5T2Q7Wp9rm5oKlSZvBp1ZzqH/
/KBWON4nw2il6dwUFQ61V7PoVW8w4lc8Qyj6GSaRfVLYCMIX+uipKdBXTx2PNJyxcaz7eh0ivksZ
LNqvST2xpJUAXb2KHUB+VMIhnISeWGCoZKkZYlSavfXPRkWhIBi6qoO4Jby6Yanv8WZB0zhpJrt9
dh3gChYU2RvbuYBZXkPA5EL7uadWPcGm5VNOfoDDu6PatrMo3xQNDzgtEdT9orz2lIFAm8jVQMPO
7E6gT/CJVvzaXarvXASVJ3VAKbGxvb01rceGSoQNAiyS4SXAuY9B2k/z1gngLhv/v51Yr2bWNvBD
KiZteRnE6GB03xwo4lfQp9CT8lFvRoBJuskhGdJo3ajdutCA+6DMIsYDlWfAq1SbojeL4LdX/Wbr
XHQY1NKdhyrbUcs2JmXc7OgWUw7CuH8EICOrA/sMeOYR/osPkvI1X7I8Z8n8PrI7jQQEWYKf3WK1
C3QrHG77SBstEsih1GZHhSKRfR+XG3PdI1v4sidsFtsOQ58siRrV4bRKaUx2VvQ6E1VJxzy+dSvn
mt4rqLRwg7gnpHTH0SHwPTEeOLwIDPKkC/2fwbIncKtZAjCmMMbIqZ6eYm0BUPF34YxjHHIQfgm2
bOEhBjUG3MHWzj3MQFiGGx+F+Ey3GgS5YFsDueOJpJLHb5T9oORdNPtiGT9qaCzHartZ40RTgWxJ
10BpMcY54N4BEWkij4QU3mcJzD6Hhe0VqyxUPLXTi7NFdix69qgc5qhaKhzD1kSwLIszYpv1Itbx
xlFabtjOUodikd3jB46UItJe2dCT9z95SEhcZ5tFqe4H7ksU1jtgRmcw+StDvBuTdWIWsufWCtKH
x+ePEAE3eca70XOAw6aeJahgU+FWJeEibwgnp6qQBRgAjX73ZiMFJTUzDjCSgpz7kuLUzhdWwzCt
STK1dbF8b2kSKv/BIs6R7E3gP9lTocdXR9XYw6YycWf7bRb/MuKOdx8v45yQ8qWM99gdQFIrWvxQ
HMnEmv3OdJriWyMQqxEeE5RyIbOaJxXaGq/d6hOYcTN/IP0IlZD+ct/DI0BVldSvBIOs6XYApoLK
rKht0OCflcwJG5R4Ye4f0Sx/zYbdplD/7qkL0ANjqh7GXGmj8frSoKCR2yam9MaajA3rh7VtfRyZ
4TKlHkf2HMTlNZyHjNg1J4T/GIQ9L56Lgbv7NFSJLJuBN11h2pwyk5R7/O0NmYgAy8wzYFn99raE
kUhmSjQ1G9eEFbsrsvG4eSabBvPNsdKJ0oo1O61w3UNxo72n0gmNx9mR3jNNQDjDOrr8+EwFMydR
H9qPRt3Vhrgapmcr/Nx2TbmIyUG8lr/s7R44GW/YDc9itVawtQVPRTuv/vtN9qeZVZZB3RYVldqC
/wFrfRPruP3icp6/JgPfWAcBdJp/RnTEPAVtoGnECT2MUI8//X6qj2xa+MPW779uyX3sowfVvANY
fgfIc+uWeAizPFbDTBtRGsiS8TjRQTyM4rJpZhnWi4sq/05YyrxAF0C+yz3QSwWsujKtwepX/6Nc
KGo4gCGKKtGVS2hfoo+20hYhOKxM6jJI1vU6onD/x0Ujg6KOpIdDCLmsR/1EUbiGuHbNyPwqJHTP
6jxiLAVF0h6+I7GASZNoFnD85ph7GUKvjAuJhLUn8CkigGTwNiWm0pnp7IAkM3DlbmDzUZsWKyh/
IlxoYo3PZmsanz/GER6fZS5AkGQ5QSXhZOOV4gOHG3AwOIpcLV6V2DjNQ4+b14PQm2AiiskO5ifa
Yw6Yy67XzM9ML6q8rJViN4KZ+H9TFFRXjTb5kZIpE4X2JMtfgvFtmXAx+cJ6qtYxK1zUlob7TTRQ
DrD6fzx+K1LG2myglEVYWMhNastmbLPBzn4ion7YaVK0iL7cjX3kyNwgK1ZKIG7gNu81rZkgX39o
8ctxvezuP6ncvJqZBac/t00Mju30nzliNWXJnWdfsPm5U//2aFNaPong5zxIsW9iLMgvxbMdwd1R
EAHqhhGpumtrcZNSZuvJmXvR4Q9C64usCMyj8lp05cptlV2ugl6FP3UBJ7g2MGYYC3m8N++QX0wc
QR5DkvPnFdLeiWh0qNA6276x/hOxVvbMYh4wMmWzZOAxs0vm+m7l9uR1AIr9/GmARx36CX5D+HIt
c72BCFCEUlnmXsXbnM+LYrgUt5+g7a2eMjkrpEgA5PrjOkx35bhXcPOHDuZQ/a2B8Ia1rJ8pCrD8
Gs70y7qo0oWICSiv6LZDpwN4398xCrP/FpG51mKJc2ExuoZBb1xpwK/GM6U+jlt1OLB4Q2Lhjy+U
3K5eXLYYL9m+cq1z7M1MT/eWRJgl6a8y16ATDvCHnx8lif7ksABF+7cw0V/mmrH0BMo5hPX1mtj6
jndK1VrJ387Piou2pMnZ84URDQFwZavD9W9pDLYLXL3dFcD+Vsf8j3ztowJSR7TmPJCyTu6XNn5B
M8PX2arJEeJ4Hz+RR3ldHlGltClj+41w0hG4R6KUzv9e3oGpe8tbn9Szvlax0Xkf6nLSu5Nt50aa
CGwHDHJaAjZhxI9DwI2ajm+YWhElBHgHtAe+AxiTX8mqg0Wt6Al9QBeg5Icxkom9DebdPC/eDXxE
cGigLQpr9wn88cUXHcwBXimGX9Orv9HmmfkrgISliFrPumexdyAatWueQV4qaV/k2Zw5V+RI2u0S
ctJXtVcQIHY+mvLiurgERr7ppx80jWXdZma4HTevQlBMjmICTJv9GcEV3Uh4ps1G60MRikofjbzj
i28fOVTv8sa4dafWyP69cGJk3/XtAUmR7ATz84aBzcBfaMhVsQnepRkXefXKkk98EeTthjwMe4PH
WaQ46Nwk7kjWFeGACb/dyuI/3CpLtXZJbCMg1k7jgzX+HC0Mkq61cE9ZlTSL7rzpiM5GVfH4t9OU
03CNf7ViKKSvJ9Q3nIp6n4dSG0aQCgZD86dfa7zy1S5xBmXgbB1EZzsMoaRDRR2wxL79rfIVsHYY
fZbI13oEabr/EyKSPdcw1VKlUXcdW24TRuNEQvoAApFxc4TCT5gLMTCx9kTWpU7jvO7rx/mGpVEI
yAcqNwNE3yoW0Or/j238VtgXMtpx4gWwev8rC2CvyQ8QN75poTHQW/3/q6kuz1j+uFbxUk/lPVcp
A5yUKTP7s0CA2eS01CL14qPjaO/EDxIlqCSzPGtUhPAAOddK4BZuWlgZrUeRJLKIEV3yYpnzg/95
93820HOnJ997PKwrp934ebLb1L5miKa+qhupdGUJCl3hG4VJ890zk0QGMNGpKi/ZVjnEr6aYPI5M
25YND5XQ7NpelK2qJwTyTEoITR9B535GpmYPbk+ligKDu2N5CAA57P0oS6EqwLz6lrieA9NtoWjW
s1J8qYbCA52UoNyefR16PpCm8Hc8OAX+Qwcr9gziucmuzZ3Ui6SyVIkijV2hg3Ytra1EqsO4I4mo
P32VDRxbzbu1yFyeE7SG/vFiiuQOZmmLqQGGNKLs7wUJAxEwdEEWkiGMIcfaKSQcw1EyKxlVlJjI
DWJzYk40JutD+kzPWkUBjLKsh6ZpWLG4Ou00intNqsqZr4Q+m0dtdgbaUP/3d5BQNxUx9BaX6HF8
vs7vSQ/v0Wxf+Luobeq9R4BY8yDZTl0gfDFXawrXYy4i3ivmxccNkIirwXiWiDbGNdIgMXtQ/phz
DrmhiNqq5MGFC7BZLrh+aTT2OldFKxCm5e9KSzRTe9moQ4M8UQau3vReJKc2IDvkf/mnLj4X2dLK
/Dn9WLugpOWs7uVLGsj/0435FzCqaJBo9l8QmbpRZPE0KtYAKxdETz+rxvHuTJMB7gJojpSH8Cdo
n2iebmmwRrRAa2gl/rn8skwLKnGFU2qllEmXyWi7eaqd7Xt414y/YUDE2BxledAaYLjgJyFncRNc
D2CnmED1DmNLlUwvg2Ro1ZS/mWy1PVEuKpp89D77LGtToRfciFxarsmP1xngRlduanTYZVwpmzuz
uf/zsFwxUJ2KBPMJcmWx/euMOtn+tLpmQ1d5YJeGZUrhHBuZT+6ntEmzNa6c8xffxS9ovCs2AGuQ
cOVJJe1SpO1h4GGylOMN67vXjSMaphkABhivN+wrVRv4opSjoYr5fbrzFZhPgYqRzbDS5QJDXySJ
Z6NWqi3e+NS60UZqiZtC1t6rDnPBZbB0Bsb31ARxMXCxx6NovdD9lvI5lx0wh9Uq4OEnMYuyU/ur
KWbYK/d2CnDAd17xr+VVBfwlZGZnhcY8lwcAgbI3k4GqA2KBMH7TkvcBRRtC7/nwYbBddh53fB7s
YlXSTh2wb901dDTFFmcv0I8+sgXp3zAUW3CxmVs0hc0OKZyR3hpzBcrRG5iHBdvGZEi1dsue+DCE
ccM7K/t6KWn7PVOesqG1E09RrdKW3AVInWfHLQBf7TzRENVbNzJBYHENYQ7K7Av0epoegbexug6c
Hm1+gBk5ckxotInBKuwmUXox4URi5Wq84iclfAWzBsYigDTPcwIe+dlA3c1Q79OJIMLSbnmZQZem
stU/02hstgPBj5IOcfzhLSjcMdh4Frm3APrqlww5/srctGKL1HOoWb6hTcF/h+XG/l8KOMYu02uq
qjU5RwHHVFdj6lpDlebd1Z//czWhWMVxyiz1cgihpqNHxZn3XnwiCvqa/o0LqgJd92OE8H3FnnNM
ZCDFI61AvGHGkHGHOTSVCG5MFZpU6X6beVG25PNVkAHAXOQmAveDsfMve/B//mq4gomJxcX/yRKT
Ko3BTnbD5HK5Cqt32ZpcWKOX6KlF79Y6hG7o2tKBe2PFNrGs3ASVuKi/2g88mVNfxyQ230peL8eV
mnde5AJpAPpWeyAQpd1Rx04WNHXMoOaAk7iWNZ8meF0+FRjp8Dp48XmwNxu+L2tilKRVuiOG7an3
UAXg2OedERCN3n1tixwm50U6jeQP4S+3w4AlLTxD7F598qXL1WesA5zowVD57TvaOJUWULaOIcgK
e9Hkfpp0bN5ZqBdO3GGh8SwsEQiyARFnwg1rBC/TYQt2Eger43S8F44DsMZGD0z2j/scYpwuR+EW
66iTiV8dYlecqpjbgEs7DJqCVSVQlym/hCpB894UGx2Ku6BifRvVi3/yXdDHA7ArXywLNhJwYnCS
XAoyMEd+WEMUo9GZ4zO3FYjBDxIhSrX1E9RwoM2BcCLcK+8h0YgbyGJ93lqmAQwXUs5T0V66ju6s
r0ZfjPH/7VYxmpQGuOA9Hd9qgE2Gy71Mx8ANXthqvw6si2KyID2UZeqE59YN9JJuW0nqIFcesLsS
WwJqoRi4HxSmaWxT9plt0Z8Qo5PSi+fqW/dawRyW95UrwnnTkLW+FuOLvYuIkUFMGOOzEQs7FLB1
qCwVEcvXgylBQvMr/r4oGqqUXy9VkqCvVTulInrBmYD7a/Ttc+4Ed8TCOGAax95FfFBk1uXaKEXb
AALr01XzTyn7ltQdXqQMjqWe1plN8eALTIpb9DyNTLFGRrMvU/DqpaNafkS3lJIZFUITfhLblhXQ
jTTstQR4jIfh0rl/smgXJRZ9Jxp+QlCj8/6O7bUTze1sVDaE+9uj8uO8DOm8EeocE/hJVHv7TtGb
m8iVeJNb1vNWUBKwEPydHcEXGi/nKPe28ZN3mrgEOPk36apClCCbBe7Pe+paxTz5bYlTvx/1yvXZ
Ns1KX1fnecg29iwoIKHRznI+OTBGlNQuJZVsnyH7wkKGEeChjURDarUUV6hVvYCSjrMzAlIBHYAf
nAMoQqMk4M0igm/VBq3MNVyJIu/30o4mPcR2x20jJDJqax6uOF0LhPo+uSnqweM2LS+vjt0KbzXf
uuEL+oCcKH7Zkctf3FQqRKn9DpinosLAsWUByXQ5hBsQNLM3/KETc0J+Ih6ZB/qjHB4D1D5AxnzY
A/UTE2ZUUcLpzxcAIVVfo8/VdnkE6NDkpxyZkEIuVIhWu000Zbr5KQPihMuLBI56moxfxHonENo5
tF8arGWoDqI+GKWHHwAAFqeyPeUdXCLsG+y+BoDzeeFAPfD/dg2M24Xm2OGDcAViVJemlpfAhqBJ
6tmn3rMYA6RJbMzaVW20E1g/JwsCjskSglnxrj5sYxhzmh3FuRfZS3/ScYhEZIrQE83oLFVkUAjz
E3yXHkyThdQpKCG6kf9DHv81Yh8Srer4pwxJwNbdk3978mOWgNIIlXBxJ9I9mbbfrp5PQ8YS0/Le
cHoYpO8sVwIGKW3mY85EOD0ubzUrRLaohjIHNjT1alTxEGTluU6YxtpNCvwjlCMBX35P/DmQrVBl
9dPk2zbB3kXphMsW6YezMxcjSxFWK9HJpXpuBb12AkC+L+2Jnzv0A+64Y6p2En+Y9yzSih1lLGlV
yCMdOq9J3hv+aZDG+mXmNNcNcvodV/RwqpEsOWODLB54kQwsswHShuvzsUcbQjxt5hHyMnbvDFj3
3G1Vq+DV2sbmT3YFNDkEvnR+MVbmO8m321yCB7Qz1noOJABtOptCRxFvFpEYPlZSqxFsxgDpp9te
SySFcE7hgJ/toMt2lca4NPidUEfxAfN48a50pUFDX1R/XpNbnIA7XDKGYVaKnk63nwir1R1Y659B
VgXlR05AYtXSE0W9O6z3iM+PRXoa4y62uN2GqMCRJwku0i7gqoV606bgVRgTXG0DBddK/AuKHRDJ
4JR9r7qAOoxx9K/mCUQxdmQtptVPLXZYlD1AzjAiUPE7au5voExxV5ihU+69Un7fjB64hVj9bgjM
0L+Duq0+jZkXIE67LeAUZQEvZlMHGEOH8UoVivqaKIWYr9mxL+p1/vXjNW4vVyFrR0Wwo+cwafqR
kA5fwagXhppmGb3yUaxVblImjsmwiqlpd6hlLs1YHRyDaoR7u+Ltru1dVTG8VnYbf0MyQs+JfYL0
Jb9RHnKnQp1WeBt9l5JdN0r57QOppX9Lgsy/yQl+lfeziGmTkxwCeDiEBeMnsFkBSP3OVZeqWoj1
y/Uh2951hBcwwg36ACbTfuzjQWCS9q6+9YzRYWNCRcmX2U+KAhDqbsCWp6nQ9D6gSul8SVu5piD1
VEy/d+Q4D8S09BNjJhk8Z4L0yO6yFN0Ig5qIpVXWAS7tl5YASspAAZRPpMlQ+LT99CsYKqcgc60V
aitPshQCvoQXPf3PvhGs4jSXhVlbj0ZBSoCOfnf556VY2AZzQCzVZJaW9ZTiAHSqw06l8vlFysg4
WM2FyznjTaHTmSsi+kBpVnajXYJeaKHFMeMdWy0kK+BY79B1zTsPg+LiNu5fnNwsuvnX9fkGLhGJ
yEEy5pJCU3WaIG5DlcLL4wWvJsbhBlrORYM2dGqLxp2t4T+yBoLj62ZlkafKVzLZHQLCMhhVaHvA
uTMFXywkfrq97KnG5XUJno19Rd+4bVzW0eHKj8UtwfuBcOlDcFHxdoguZIoyzyZsRGBOVOQTIZBz
O/lxui8rAP2Dp6eGMJ+5j0CZFm3D4wWj/nf6XliwrbPLUJwZwGZ81bmJaqDQmIxccPruiFiPL5J1
obdQVyyrei6/tJ4p+4lP87CIHYPbwi/PQRXcqmWZfIaQgAO8GB+ep8+jOVE1PRJhA8wxQ8tS8esf
mJ568UMxWt4dh5mf0jsc2ZsrCbrBPNXZtersnkUqJsRsTLeHrL0wsArQnWlU1zmjAt+A6FqKFJv9
b0FJXXgPMESAIDSAFek1JpLyt7IhPmBXbaNIwKvHHdeCCMWVdvHF0n4fo7kdqEW/fgTazx1cd7sw
Bgrc69UA8Omvd+MVosdxipeX77zLdIgEsMXR/BGCO0LuOZJew/OQlzwLP4erCUGRQxXfogGlV4Vt
00B3PkmyxYkNEKvLsr9Fg8lr68q/U+ztqvOdrtJe3IlI3uRsLBnE9Cvpu5ej+NHH4wmUOhHaW4W4
CX4/7g5bmeJT7LVbt/CYTGYWjKvMCLy2CFFT6fozlNTtK1mkHbbvKuwGmMY7VrZT60alxgYR5Zxn
EUC5KSddND+BcKCvV6raVj08xAQu57s4VzfRAhSSZGHk3j9GyhMdr/6v4zgsf0QDrUVgs5eUDRER
pKEwgI/qO17zEBZhZLy3EcubWKPQbcVO278Rp1YNOuPDVu+G9Tt6qhXZqP+GowX1iLzMzj5hZBZy
9KryLdyMWV/w7m5VjvgBz9gz9Ip64vfj9svBcrWIExStFD8+XAh4jg2Bhvk/Vy2ah+OUfb5tLODn
k7FTw873I36OdxgrJp8Ww5FpeDpIHAAGtxNGfd5gCSQ8qxDdQdZDJ5sXFffRgpCxUBkL3E8UCqH0
rAfiB/fUIOVvGRDipaQkkji4G6inhc10j6y1geoH9bGgSoah9foT/IQ0KTR6NLCeuO3bevQgpraN
WSwAg6NrnX4nonIkV/Gv21gmX5swlos5FRig5jOqN9HWWCHp0TSF/g3y5PuBcxs1boKXu0UT8gze
YY42Be9GEqYBd8SIGvR2flSnv+2B2g5PznCDU87P3icXyn95OYvnSm68A3Sg0Zd8QWl8JLG3TZtu
IZzL914djq/KjAl/3hXp9PCozcKJggCBLinUb9CNOmNQKlIhbDPddkHeTATFL2N1H6X8JVE29P2b
lWw76ngUSHTzzKPkJmWjHxlr2zmV3fXrWNqm+KaL/6cDoGylNd1M9Bu9y9LzQ4nBuix9LKWfOAmX
0lA+TmWPx23ye0+pEHa32hRzvfL7ptPsKk4ehB71Lz+InF97p/KgyOCsBw6nh+yvhqKJSi5xJG04
WqGkqEvZn+sFMmzl4yUo7xDBqBaniGamlW6qAEBdB8rXgMumKFWeToiE1Io2rHbI3ai31quubJn+
t4NG328SVdjDMs80BP1hinTfn7gf5ICLFSQU7OC+TeFs0DtF1mstionT3vyKBXk3e6VXuNGtUsWN
LG1uJGT/cQUEd22BW4KX8SyiVT2D/bZU53civ/uhyZH5JG+e5iUuBs9fR4K8EVgLmmapqnlk53LB
O3h5lbuEsZ1LtFk333NYeO0Ihm49gEEd/GuBBXmm0WCrNjHSeYJaBJP2RO0cqFGerwY+NrJBVJdA
alMsQo3SVYKGspzXjOug3Qy0KDOqfOqxg2diOkcVsI+hKFmUkqMDn7iB1IBxT3vydwerhVht8aQJ
5qfbzmjPHzUEP9OSiYVY0WPxWwqBNYogxTw9St/Cu3VKCz/U0Tcad5gRQjN4vFpktxKrVj0z6wQe
vu6fN77UJvYPLK9a4gUdVTiv4e9d0AN3kZfaNI/Ku+nK9RptAQNbV14npjrxoJURo+xXyl0NPTvb
bDYar8UTUoKURBVH7MnMOJuIGZjqkbyHlhHzU2sKs37oS4JlVNTfwjC0TCvsOUHjc5hg/JVoruRH
uD3/v5Axf7It0wfagxFQgEuzUVfZsB9jnrpIAYPaeKPWOB8gSo8dgOhCgEPflh1cQDBIrXI5vICh
LNfgi1i6BiE7wudK/VVlQQNHIacjAGKoBaOG4aFLOtIO+TznKGSnR+stJg/LpMw52IgExI35MqqM
EAu/2V2fLdsqSw7XCGHigQjRRw0oSL/yu4/E5uv4KD9RrWbS4HDS9/vqTMN71f2n08ZSHO4cNc/i
ofmW2eXCgGksYAjEAcGOKpG/n+1qP+tp2Al53CPK7l92n3TrZMHzo7kuQ8PHElLozhofogq5blI7
8lbtkEutx1S1VIEQNOybjOBmw23a/BVrz9sWaK9HiPOPQQvd24xXm8jyE9fr/2CDZEPVlW7D93rj
Va3+xa29LupVA7+xG2KM6yDBj9q+KMY26bC1niz2FZYNM0fwNTR2SriXaUPFzX/ZloNinCekQDin
9wj951fFI7d0kWpZizDltE68r17mrfRmuZSt1rYWS1/cr/H5FGJ9tIn2qS58hX44xVvcTF6PA73q
c/FP/+J7CKf+/avtMKhO6n7Ovc2uE3WbyIWx/IlB76ClfY26tRvigLvCUwyiyfNZpB3CN2/qfjnr
kQz07UvmDOVPRFF7759+Hkd/iGY5DiGJ/6raHautBHj/BCyLZudQsRacCRoGdpEGjwzSkWdz2Ca0
FtjRWRSe6LZIK8h/vNAhdpoT7COxb2fJBhOT0drOPVTjGWJ0IeXcEFBN+ECfPc5FMnTD+Uu7oays
6WoIY0/mB3J7A0gsa6FED4HXHhxz5O7LC2fVcTREL+I6VoXyxTD61Onup4UucEs1v41wJgMSatXa
wumd0ZPf3VZ7l7lM/SLJLQvO901VUcbFCxVKT24ssHjSH48XQD1LSUtOS3rTX/bPeb37arigMnNP
1mY4Bdxl6+EYMstBhBj6ZW5Ovk3vwqXCTTtjMMomThrdieELDd3lbu4p473vvXyQ7lLLxAgA8xdJ
da8sT+JulF1dOuL5o/5Buxgg7gWa7++V2T4eYL3ib6RKtMl063hxkLO23SeF2xXJDmvVwLV7Jre9
LcXoERuWAPhxqv4XPYlN5yK8V8w6PoeCaW2Z+KU9SllsXxOeN227ocWOND/7ECnj9rgIwBPU7qw6
Eub1Ic522SR9daJap+xV6xo0YVvzNeHE8vnAPCBo85YPuv8D+WPXU9j0IJVK3/ZAu7nOAZFxKjN0
lf1J8ZlGW0Bu6U0bhy+TDMrYHKV45Xjk9esSfHsi2FlfqXUJAhbtwRqfGmn1WQq/gmiTbJJnO/5m
P+HHwX3z7Nn476n/D6O6oBEuh6U03K7IkqrSLsNQhunwkKsL7wkzzHirkxCuqEaLcKegL21fe/Xu
MkYrhQugwoKTbVZ3Yo0v9cvXAh91DD7wRYk+C+uuokh8y9E7liTMJkuITp6LPGyyGtcElCSAYkSQ
Yu/eIElju55bPGTJDAzus9RNPXTZZ7vlsrPCpSWYH3ILUIV7lBgEyfGUBHz4e1GMUJ6pbmZIfugb
HRmGCIaDXlt8Camt5NIl7C34uheR32e0dw6skXDdvCMDSOcRDd+KQYuu912yPk1VMS+8b2CGMe3C
mmgJtJjPhJ9WYFM3nTt554Co3lM87B2KbcZRvMjRANMfPeFUctejMUjHt268y3oMQE933empkqzl
xb0fAssNTBI1pgwziFK/9LJSEj0D/f7DCg01O1pzpzIkMZ6YbClC5hSW+p9mEPAkiSiuyFFzZE1f
gZUJwNvbJG9k4Tdt/fVFCsAT/MF4Azwlp/AcKJitFGcIpe+FeSjX0vKR8BUCfkUEEYKYV+52FpZS
13xB31gpQWBCuAIBfpLCV8zpaWHqLRdaSN+jshI2DWbK72ZqwWSqJHP4NT6YiBGCw4jUiF/VvEDN
7AE+HTcwU6pI4qC/6nOLORjxvkmGvJrpd42PsLXFHTTNcQ/x1G+dctSd6Ilw+ASbs82Nu3oK604g
K3vEhSzszHsjkSeZ7GjVVfEPamhUUFCghkjoC67NdKoGzZv0ImMFwnbqJ/s465rhSWFLExgvZJsy
HiM7sPpBbahWELxZ+lQxUMMcnElb2uoSgR81RXZ/pWokbzms70XX1N2MvmGvitjmdHxMSU/BIAxA
LiQkyib8NzpiTCqAt7xHJcG295N9SRMc/vIyRwbb/SRwhV6+Rh51UOzXfDEY6b+vLeoWHJUp8K74
wHwYpKvOiFcUV21ZGOmS4IqsjNCOR4DEToR9Rwtr8RcFyV/J1d63ovm+XRCEeXSjyn486tP/+qgs
3OlTTdrhiGuia6dM8ybAGktXd63QnaqjKSEx7j8fpZ/H4jC3cSagiLrDKayh+kGbRdndt+LrXm27
TeNz30zrxUXSCOcjLGzdrdC8z5eKGhSqJFMLnUqLKcYVG7Z73DQPbA+t7QHX2S5ZS/TLZDcVO6yv
cXEcpWJPYJ1hkGr//hGYmOGOeAU82nhnDO+qhwCVN6LoxreiKHYnSrMCTH/VVJqxpuX+1wu+AgRM
nHXy6vLvumtCLJZ3E/kGBmNex3ZUrifs7Lax8Bb1USUG0650eGg7WflwJcoj37w+XRTyuumgGObv
u6rx36jw0/7mmY6KP5BqJA7cdoqqfpOeIIsH9W8GVb1TDdyKB9tPmzD2PBMe795279j+z2Yhakor
skL3y61bpYVuG+AB9fr4zcRYQuM/mGlWvI0DJPq6mQjwweKCY4ZGWV1C3RKWOoDn25euuywv9AtN
chHr/s7FBVPZ5o139yVcAJbXjkIRlLU24BBynI+wJ4dRiylQG+A83Ch8PV91udbwwgtChjaOKfuN
4aNMxyNlabeiQVf86wIVYMhVF5Xt01OLPmUEanqS9F586tYojCGzoactYtJBwoZDvGboJITQ9CgV
YxRiVj2gaMQHsRQOFCLxHSxNXw/ebiz6AIDce47vbpzglRSPfj4/o4BtIFl5EoScC+Ap1L48+NDv
E/YTvh8D/bokUFCtFjFc36i8cJAM88DLg49tJXJ1xfyx/iTjXRPxbfmm/xSa+PYvMa6BXiUin199
qXnp/tqiwLwC4ibtTFg/GSRmXbq59UtiwifQO2sS5TMGl1btgtGIgYuRHDB3jAIIXZ3ENvF1q6IA
DwTHfLYahoK/V8FIlylDqg3gi4jGLZr/jrqofiUf6wEpSJmJZ48FZrfLsfRyA0El962yYbh7jCaN
V6F6xTlshwjBkJ1aPHNXQ+fjFYr1Z2eQFaSpZitmYPVjdeERMo9ARDDjX9B03yCSqpAedZkEBc8g
OgifNsDBLTnxSMBzryUoPMrYFpVbez1M/po7Qct2eB+MjtDeeipd+vd0bcp4DSCzlU8stw7CcSdj
UkoOJnbEj/alNDFrrqmfAmusJXB1UEV9671cWNHlG55239S0h7nPyo/hkc9mSbw1FP0TpfqkdkYC
sbsKH9BPjmATeRqFd2BflV54fjyv/iGY5C+5tw75n4DfCMwqExkrLlbr5T6H5Kv5+eUzR0xL13w3
8LJzDKNNGaUAANPvuei3aPDqsaGJuzX6s2cA20BBKbFWcbKob6VnlWTpqC2zQlmNp7Gbu+/CLtJk
SPIF5mT0gs5/zS5LTdvEvJaHXofmdnLHeatJgf0KgC97oWIG0RhxZBLEvZNQaD88dkbyoNXgH9DD
Uj8TcJ9vU4GB92xGkhCn9r08+qiWIL3q1Z0kqbPy7JL/Z0IKsZbr3o5hQzVsykjPnAgsMau67eoT
iXoiNoor3jIuaCPZ8jVpgC0hZm+ea6O+auhfoXn56zYDhqZBpIgt4lZWyasZZyP4iUqdvscpIjks
l2Ca+EPneH8EY5fhky0Wu02QsMhppAk4AAdvJkfJ25NeLhU6QLlAXSx6rxNdoy7PhWKnDFK/qNLi
bt1akDqiiolVH9SebjwlYKsgyveeCVjpAYoEDww9yP7fYcqwqmFaAXN9EQAGwyPx6SwFarv7z35k
94dvz8AdEg3dT2+bVU7VA1LvVpzi5G8MoAUNMFall3CmBbh4XOVhyZjsWHKYyfaP/SZVm+FnKyVo
1oTl+nGcwM8OZyepDFt7t/oU2kdoFOZKqNykwQfgfxWtqQPwrhj5n4M4Dozzp8IiY0y2NTD5iXrF
khb0hsxPDQgRXv+dsvT0YVCAc2zhbxryxL6UD6ewEFrR8gbcSeWrSkToId5c1SGJa1x4qwIcYUdp
/W7saAyzEsVWeUJM7aYGHBtQ8gDBXGveGqA9G/AXYep7syYX6QZsUF9V/wGWOUz1rEWtetz7iA2n
zA+dJQ9zbRYNXUwa+u4/69ZArTs1s3F2CBxw1QFxPEFb/9YjLUCqcn29fJQoyy5sUPrlelCE6KJE
31Sb7MiJto+QLlTiIAyF5AXlO/1Nwo6KstRgz/c8WJB52p0MCQoLhS3okN39WtlQUd8pL64vdvus
IeY3JQ7ptMrkeN85FZ+1V7Mfd57flAutQ+zY6piGWAoLxZhkfcpjiFoJFLWuJoHE0ypO9iKlc9k4
rq5xaiQDQQJ6Ny/RMom6KhDGMHtcCrHqGHs9m/AFvsor/atPKkUTQD7yOXMdPO9CEtDXWJjfOb+s
BXwlLHifTLPjHCh+P8XO0pStnCQnb+x6EhTVgWFZa1WEM2/baWHiRDmLvy5REabyWgRZR/4Q4lwM
pxMTqwvTS7JY3UbmUtfwwPR6wcqYiSr2Yuv59x/PMjjMwg3THmxNZ3e1eG0ASKUZSb4QkUdgt79t
qdAwc9wHbnWmm47TOwKuWIdgIVfoTHeyW6L+ox0i/gW8HW8JSJKpurPYkN2cZ1EMys+H8m3HZPfn
DYJqZCp9iIe/8Sn97oyhdmVjTvk6yP7Zx/kvrfCg1jT65m47hDkI3/TtcTg8v/iFEPpqo/4H/G3s
TXsO8YP9ja7DyVPtkJxp43l7JHAs9u7TLrBHTqedsbbvLleCIn+0ZDGHdBf18BvC8N81RYbWE0j0
FTdC9IXhcJE2bbXF6q5bDpS4UEy73kAvjUzBZ0XCI2gYeVMRp6TNxZMYPU6kYTZjad7b6XnUOYUr
HoGXFl1Xy31yddxB+SzkD8eeh5DjoBWmQJHWaswaAfohMVuyEg4a9Wo1YXBq1B3mnl/uaU5gt87x
pEVTYa1HBdyY5GVKwNIF60OtevyolBR+0CljfPMHWGpI5zOq7I9XdpJDiXYAqw+iljooHRwZK1bb
0qpR5zN2LY2FlmBGhVw5QLJxX0lCojrgQW36YDZde8isJWir+5XLWTh83eRVFMozkZjmlcwq3vBl
J2eaZilBAeKWrQ9bHz9pYTzmizveNv8J6NouwNfdzClWNmGChf1g6hnbdNMnndE2s1z7aHqTtrMn
0kgWDOjS0GNuvBNsCxAjL8SE1flIrt7rWSZS0iQO/s1yqBtEvLAFx/MtirQHK3eO3MT884BbHXc7
ALYkuqggD8LVNS7qt3aHu3mVu8WTLVgAzqu8yree1gMGsbvHcTtd5AoE35z4K8Khsg9jyVDwGtrm
d6FPCUL+2OSc20p2wFgVE/UPeBwX7TyxhNvVvC7bpc0z8dFo7BeEEKh4OzqAQkqqy7VvtXjoiccL
AIMIG8xwufOaqzKLNLJVDiw1sWnt5yBexkFc5JZvLe3gYLnQZHRuEWFiRrF5FQabSOb2cvuT++6K
Wfj11o5c5RCVdxdPo7bkZ8i+gIZMklpmmHzTqE0XA7Aj1Qnzr5rNnITzlnNaXnCOufQNBDKujaNZ
+8wZXu63F3H/VUzlqJaZHbHcFHn7+eT37fIMjCMSiDd4Jl1RVPDcOfWo63joq4z1uIeP2eJhXNZh
hNFNgH+VG3+zZ4qXQ9YUZc4yWSKgr087Q5/ZPaKSxtZaTOHLngXsjfKUEjqVzOetwYVhy4W3RHh9
zU0+PTGUojV2g8zOZqQFfFxoU7n/eaKk2toM1hqNOilD3m2OIyPKvo8UQPYsWu6U3tfaHUkWbCsw
0lMIrQTx1a2CbYqPj8C3lBVO/mdpQhjwVHjRkgLMZHQByAuKH96CRhMf8ZAXEUifgRLeuTchMs5q
hpA3lG2DrBTFlc/LFXmfmEvQRrny3bCcVJWg946y9i7yXwdIDb+r2TznDBAYVe0tj6j0UhFh6s5Q
l5ofLJRwheNEdttXOQ8Q74b/H16jqH8RdGhVgxq0HoZW43BJ1uBLgnI7gyFadyfUlbdR0PlMD0cr
x5DDG7xOXRhCblbwRxOFrtXuOxdtMZv/3uC+6ufEo+3BVWD1L/JiB/QWC4MDesKnKz9oNfwYhTdz
ObFIH+/cz51bdwt4mpYk6l4GwVG+BvtYgiq6gdHpHN/2OifZupbGcgCwIaunraB2MV38CrbFY//Y
pOMCPN465i6KxJv+BDc1iMv1Mp6s6Ay1SBGcoigBD1dYaknsBTciuuyUB4Afi5CicQb1/as7rmKQ
t7QIHL7VU346+2NfUcsn+0zbJrLEFeh+PWz75KducSVjuR5hkSK9qkUOTYKiI6sjG3Kig9rO9CsO
kUuFt6thGlqlepTY6K56Z3sTU4FpWlfBhkOGM/ODRtcOx66em5zQ9/Ji3/7bdVdTcuA5wEB/r1qD
gXPCMSWMcoLhQWD2WQdQsmYNVsYWUrf22qhO9GXvXiD7WgRltr+QnWPfWO62PZfduhmo3F15JSCg
nbyE4rpzTFh3abFdGYBmn/CAgeZSgU/M5Rp8KrWsj8V5paxImY0UyQih/atLkBgCT8CEeUDqv5+M
NBeauUChtj+DY3mdK6egeWL02+AUdksBHa38IZ8njyZAjXLq4Ob7a3HztWnud2hio1e4rBzecfB/
BWLa4OoNwkp9xnEQrM+WXINiGiWqzxjYqbp+CbWip8Ox3X/KyZcLwg9WLHigyfut00cboFpcVvRc
R+wB91nhMUjO+sk60quw/vAiC98cphsdb1HX58Dv+ODtbN36gJvwkqwcBxA+5l8k03nQSQvE9LfC
GGNxyGWbDF38gCmz/LmPyumgzeCpBCXLVt+HCZU1ewADvcMx6bDrIIKsELIlq2QkAImImKCTrA4S
I1gDPoG7goJjC8nl8ogVWEN96ghiHU/oClkJcXcivnPnit1wNm5/A9LXCkkZWOUv5xxaFwKURXQX
MMFvKlg7bTR6StQC3RZ9QwqQj/4zpruFRtou6xz+Z+2lSenz36fPZntuyj9mrsSqTA2KAeLEtY+e
anwdN77TMJYqHxLGkHM6toQCiUbzbPjxxorJZKh1JhFhB8IcZ5ckSbRhx5vCYlb1M+Th4hVdn9qa
5hs/5dUY0TpxaZVKzxAn21F8uI1A1bL7iUkAOzR4KmL+cneE8T27sfSDf6q0Yv8m9ZEDZkxvXbz1
lL1eVMSvdrhxtDs10eQ97VuF6TIuYm+mlUA/8mWrGAm7k2UodsWxEoL14Nz6OPUrDl8eB0rpRSrs
Q0IYKjHCU0oP994XXffVGS/GaczJzdfjCZPdaoWYKSQWE7HYoyzL7mT/OjisNfLqrnuvf9TK+RPu
H5FseoNvtLZRa6ST5SWH8eWJ012tEC1yK/srUdSwkU1YmoIYeKhh9/w9s+tFBUDKu714c9BxP3hu
XxtThBJRH3GGDBYd5fWdF5bgjIacZ2//Hr+UoJU4OWvPtWUJH3+uiVAO6NGf/E2BzmIaZO7/cYv2
DMwCuwhLyXnNgW/uAljFuxNuBh3LPKB4XxrWB8a2jRgFVNZe4byJV085axtyFaZ3pVi3TAlaHTdi
qEYALRHANOUTkC3FIKIciPPfous35wdI9EN80kKAFihwUw36CXCQs2yk9rRPVSC/j0tCCnon6wgp
uOY1hAgWzpTDjVwA85N9G21cFqzF29V3qUUW2cCbFaYikl57aJqz4kyHUoYtZCIIVlZC6dqr4Ato
LgZvJ9T0oj+LPkfyQX1a+FnH6nP7oxBU56QzxX12md+6bLFQHua32pJFe9BZPfWG32A4NTvS0x3o
F4UyS6HHw402wM6EhgMzMn16v8R7CSEDNd/CCbcs7vVBmESQszMyk4njV+HEPdsEukEm1FedlL5k
skv1EPvEfQ1tEKlgiSxo2/u0xIp46voetK6sRD80PSdj1KXI+fBO6+aUnCmNoShFC5IKm7wSMim7
0PvMZepObUkb2v02nD8+wEiUvtwaWPFzwTaO6ftiW1EpdZ0Z8jT5734THwCltHTo5xvWSTChY8b0
9YSmfTh78iMxXCfWua627jtC0xjxgGaoEk59uzCO5B1t5GrEnQoAlLghEui/FkLydqU6C19qhVdp
u0PA/33+nMT9mYfBQFQwwWVdbN2tCVDFJHSw/uXdoYSpHmOWUk3T8UpzhLSdwJwRFu/sLgFCTO9E
mdhENWdWgOH5LKyzBEfyPvUI6N3nYvkOqpEfsrDX4/3cMiykCMR2Ib8ruaP/28jFqXy7KPQ3ZZo1
fQiAjKjN5rqTdes+AWarWXaAB8+EIzJSet3CW+UdW7/jVWgFYEs4pA85vBQ1iOR6cpc9De4ciRJm
WVIUN7YxcuTTCvzr68kfXJQtIFepY2asJdYGetp+9HoPh9WBgeqvxcK1IxjJrwux+qQ8jFtaDSYF
0YrfXqpl5afEOkMEIJDV0mrSJyznAI1yf/ayyeQk7fGf3JykaMDO/tF7vR1VTFmEQdG+riCQlEP/
E8GcnF/RrPbeL0iAgYZDuZ0idw253OSKO2gf9eY/0dkL6ad2dbEB0zQRvbQ9lnfeBsvqdoosqkZv
uHkrwEpGDK3C8ELxttiWe2mcLRUBxhD6j8374wl5OxppZiZzRONW3vShrlNzrIOJsTEaRuXIx0UG
+0xg6jDbe7kkwqcrTNNJmTiaeQHD2EKM2GoCdDYTc2KmRqq+HJY3RlAcbvXI9+DLkPSXkjYGlAqf
aibe+oCYIRGTcLkJJqpcz+sQTw6pt4hslR/8lqVqnoQTVlMa3IPM4sS5PS9VLbk3w6yU1rBuEild
440czLJtvU1eMYTx2OwL/YQJydgKx3yZkyDpqtR+v/4j0sBlgld/GqCqT+QFCH/mMODB+6vxl7rH
EKvLDklQ1twyFWKoEQOkpBYbDJrcxBauVXS0DwT1ll8mcCTBMyfv5B78W3u/4Y/d4pq1hqiPVjQv
rWc6A0n6fW+qA0cc9gSYnNWe9Bj60tf9wH392CUw3UdJY67S6o8rRpl68TWb2umqrLRuWP9NCvWx
2cw1D11b3d4k0ooc9cEP1GJ5SXiBUNJBORBHZZhQiayc2sjhBsaBVZbAlx1CS/G34+UTsi/U5JP6
ZdawJBg84BRbzCJYxI4i0sBQL5IyTMUltI6Ua3rQy7KQyZCe1nNaWhKweDr0yBd95Xm8FPky2yKd
u2UY+okDravG3LT7G+FpWMXUD/kVKKFZoeAUGikkOY9QBzaawlR01qIWJi1Syf85K3xOsU2rZbdS
82l9FgWI1oH4OiiH5IwIgZhtcjdiF/bNIPC9ra9FjnpQ6zjryA4gDEZqbqWdtJmYaTwUU7DtT1vP
1yLayIFc3/bR9awJdYeauaOLg3ugX9sYZ1INXgaiu8LgPzZNNiwYe+Eh3TzLqWjd3+9hxNO7fTEu
SXb3hpJk9y5aINWURvY6Abmyxin9oPUK7AvTlecoIJ9NdbMU1S6T1mGoJyW28kBaPob6MT46ZHke
73LT4CeCMLY1gr+zaTgr5jSNw2U6X4Js6ulVyeL10vcPpNKUc/kB+KXwTUl3oreqvDrooFSm0i8A
w/JlY62+joGWvlGdMrkQtyI7p5CC06MKgx1DyyAwizGq8Fe5fozkaoQ3qJxwhZNYpYlerYDD3s1H
Fiz5rt72Vp4JdlsHshEjqbX9FJFL2m9oL9moRCk6xQ14KDnXGS/Ij7vmx0c6gN73uq1VKKCpMuLc
YdnttcmUzsL4HXhuAoIX0BqJg/s2ShZqYx3wdOUyeBrm4bNqNsqcvtOEtLD83cZkHPC8vI3mlTYY
lC7vV6l3I2ynG2tlIRaH3SMH4zktkfcFsW1sZlZxzyByqbbFzWY2Bw+NG8oK2E1YYusZ14Y6Dyb8
FiuFGuwNM/uvMhVLv81R6SbvHPFf2CzrB5hMwAp/Ctd7ZoX79ev7jVjsDolbp2tzFBvyh0cVEe0V
/KofXEous79jlTlh6LiXbbDoWkDm+qY598ZjrsXaICsIdokUbHbRo8hXwkQS4smhaimRC33/jjbf
ZocjXfZdx7r2V7pPCzjXh13K44mI323ulVcz2AECia5P/R8s7Qxk0O2pNsPcxK6D6pBTkV8bvTM5
k06uVySVXXg8twao1D5M2NaQH1TQfod+BUG9Sye5fsHASvowv3yX8kAuYKopvgDSQ7k4KBcck41O
NxSITKaZMKbRGlhurRo4sRSzHpMymtGPRwe3nJKzJVev3qGjpRfnEv8PfJa9WZdwHIhFXxMHSwoD
8Bvn4MOa6J/Jz1pXdiikyMo46I5mJfrBlbTDwIn+3pC61NJM4SqbKQRwYQcB5wB7642qvyUWENST
IJCWJ7p7cQPO2adN+OTKt1ux9vaNXV4cQlHcMRdUUYQ9edhaO0fiAv5UoIzv2n/pI/MQKqtoGvla
SpflI3D3OJvMM/5cFNRnutdKUCMOWjaN2Bdu/xJHzT4iw4U/PaLK0MNnfd10piZ06Tn9cnUObycc
anBzJb4ra5fuiPsjuSdNNu2Ps2HvV95qlxFXsYyGqxvz51AaboVmxr9ivb+oRwdYhD65wn54oqvw
3CfquJbAoENPaZI6kEE4QFhW46daNSZtRt9DSbMXMJfrWRnx1tF/1KoIzXfUK2hjgxp7bYqah58E
G3+INgo/W8bC3pgIm8GqLQts0JuJ1hWbJMjU8zrpbhZL2PPuxy2aPvXHgEGavpXDpWbrIv20zetW
uSBsly/MTkMjQX0zQ6dWtmorLXnLH4z7w8OTc8dDnqsXlASfrHKd30GlKt0LiGG5Jbs8qDQ5KAj1
8Lr1IZoE5BuTE+KWcgZNmpQmt+n8CzW4qfDo3GTcxlaZhOfnXEwGGq1zCgm2355mW2TN6nvCMBzO
Xgqnbdwpm4xSqx8PNAWPeEqiUNsB4Ju/CDc2RbxGuTa+12mMFCP6+vNdUFx+oTS7ScZlt5K4iqVQ
dkKIo1DdDv8bcdPR6k3UNMyDaIuJRzvvI6YQ2VBDgwbFr5GvFpD/s/118jyCh1wzAObow8d8YWqd
y9KzTk33cbriJ8UqQskTCEwfZclJgEEQB7OUQGFHmGoAiULwp+PLuZ2jJVF5EeDbKXuDfzsG2u3g
Jq2EkUZBbfXbgiy76+T7pxop2UHX3zf1c6h5mtEOR2dxmEOMz+mULGGHbm2y50qP9TB5fGEKy/u7
wuJFaf39QJpgc9N545RMxh6x5EXSeOamCi/Ml4oz77z6qnYJbIS5RKk+AE8e2N9lB91DNglLVSTq
vWys50TrIKk96adO3YVX500dUse7lubk6c58QqK2HsMVNgrABxUG8RZ1PMmD7SqElpal07mjD1dv
xB3dPEXxO1Knr3QazDUJqzN71o/bmvE3crafkidamKPXnvSyO/XbMssLcZmls0QSV3tSzrI1NrB0
RpdGXeFaBtroe0D8O5L1uy/TofeCn5ikFUx3k3fg6S7CEwP2t/f/AT4Ft0pUMY8iHhL/EftNwYt9
+sxFgg4QYLlhVdo87yGnom8qlabABqET66wyhCXSun+u5GFhpj1Q1Oml6acDCo/2FsZzdULF+Wbo
JapXJaRJoA2jZ36GZYFfdshPZFrxGIe/U9+ah1SW85NxRGNLvHkUgEgFKYhGf28y3uQhG4wj28Dg
FPGVN9IhGhxncZmCMeK6E0TPiCyjORikIOAg9AS/dSkl/Uus3g5K2FM540rHjrc7kOK5ZeHRPF0Q
PgKaBX04JQ69/iOqBghHFfTC4LRVcZodN6DwmS5AOqcxmXLYoHGkRFVaiLGXErgYIeok/6JkXCID
ToWSN2GtzdGhrCwZjChor+3CZ97QkflNq1jEOwgvrt2QOURdIdwg3eMGDQ7xXmSvHkPcgPUckEPN
uI4jrmFUF+raNTY+9ZS8ld2wRADnsnINqJZKkjCNRuQsZHKQQtvLtJk1fp6NAlJv0+Kt0NOC2r5z
6xjzGms6vqKjqywMl4CHEUFP515tTVk2mUYhdcCnzvF4rNU9Sq7f+aK6l8zKAgwc036g3MYT23Ab
KJ2hWzWeddaPfcR2M5g5My5CQ74MbUvW33mAivhgVXVHgItb0G7X+0V8MqRkFl47BlCqjFHIf9qR
V4Nomv9C4KYHzcWLJnBHoKiaQWUd1ec3im0lMc3y29VPRq+99Bj01sZxYQv+GutKvaVwNo06cZFT
iqI6dMMNBu5gPQ8s4BujJPKuBY2UGe2OfCQanAbSeqwnKBwEF8jjNYcydE0rM5ZNjZ8GvjK6lsq4
6DdYGgGtbZXCrcU6+0af70o8J34vfulO0STSGG0Y+OvrQQ54QztjhuFAwHFswVpxHaPWCRkqaZKY
1zRPnVj72MQbUU9AbYFL3XDgFx/C1NT1N4cxnyhyoQsaTYU0kM3yqnrr9tMqae5S2Lv0Yf22vH+P
RBCMXsv8FuF8mWVAXZ3NZUES7VEfFlb//SN4oLJ28QYnsurunYncLx5XB7akz9old9QJMUol/AeZ
RmvQ6C+jAUhutLDEiZz7vJjOqZUK2+rJmqRamH+znoazdyGOsGugB4XfGFmUl8qmAiVIGXFrfjQa
6pqiC1M3FL2aBsG7Z4j47wB0qVtrGSCjVgGa+92qsjp5rm5YFUedVvFRfQKsdpqqzezaMI0ddB7H
qTnMF69kdzjHcV8sehLsIx4oqu70sXROyWNK83gqCF90ddNHBz/jzcHVmJS4qEyKVrb+HvRDmfzK
GPnBdhtRX3b3E3XSDP7aGrUuYcY6puKuFaAAW6zqeAehVPF3QNcwNsFzoD8VtQdqLkrqLIySdQ9F
pIn6YSrOwEXFjyR/1kZVTetVdH+6KtbBdN57BMPb5V5cNwiWnCt04usD8YjP+nAS0WaMtvlaI44h
LyU0DN2v0JYDv9d8Lz+jdvzL9ROMwjLeiVa1711mKLtGKLRe0QeVWxahnvUAAjyQxoShbB0vOVvL
hO7S6OlGMvXQBtt3yCX1BIaP9+7aHqARlVJyl+uuOYjjesdjSelXFIhB92ddAHU9vKtRQ436ZnoQ
YM6LIW46ws1m/XW1HOOoJ/KTWvj+90pRfGQ4IS/gSsGmtUh6mRJPQTlE9yJ+632ezaHuSucQw7TA
cDqfJgvMiD+os5OeFsEghOVZQPP4zNydmXm8INxBAOlULBLHDg5Dqmf9Cv8dJA5rR2P8cC6hOAXG
/CZ2nNJAWMRONJEf2OWlicveBe7YGmQItBi6TqaPQehyyUP+wmPu7ah6y9ciEv7Jjoo9NSi2XDdw
oaCPpghjNz7H/3BfHY+XF/FErdP4VoBFktV84L22i/mpYrgLlH27er0lO4wOzsXZ4rpxCTFmpfwn
+PVqnKf6gnACxbAvTxISzXNs+Yd9CO/H835CVjm4nBAYOF+KMnEg/JRxaHLlGWszv/lkCQeY89Iz
nnmfGlvv46oZNVumb4D6vcfinhsPs7OOIcryjE8xxZnNbhfviJ0PDKY211r2OsRSh+RoQZupFimZ
eEvzH6vsAgQDwWslIaCDvyFvv4R89cQQ1Z6WnUw3KvWX09vJ1kIB0rMNJz0dmVfSCJ4nKgmLAscK
cUokzZcXUTlv/DdtyIacL1p5qUDiqOgoOwGCcdHOZurotJSfHfmAaGn58oLgYYiQj41QRdxru83s
DTMRV1wTWTxnCcwoTRGt/Wz02gfmqGZbeHlxteE0qtxThLn4IpKbmf09earmZIQ1Dy1KR2lKh7Bc
OOPwKWyPXgw/G2BXjztJQqDt9/TOS/5aW3+33dGKn8wWL/K8IACtkb+ihMcY2Fvxpm/b2iyXAzON
/bNm0wGe2wVBF68m59u1D67jWmBUnpt/MbsnwhVEm0irjZ7nzMILAlqCpXHn3PviuAH1CJrxTOWW
Br3OoBGKShstNmYr9ilxNdqkHIqIK0N5voBPG8zaG1kL7nfzYugtMpg7y9vZ8Q3YXXEs8UxRNiRI
71rOZhHsC6wDaZb1cY+T9yFrE/A+JCrMWQ7GyPpSIEACmI9F55wrMkUsiZQZDYDpXJqzJwsXvEAS
p5snQumi6ahEZDHaB6BDrmSFBC2+IE4qjDjNdGeqxw/nNhqW8xYgrshkQ4H99w7qNjnSGuQj17E/
An853+UCjtP9M/Zsq9wNzd0DfVj5dBol3IGBA2qGMx/uzMZPPArzqkgH6Ml4huM9kMUWff68nQjd
6x6AvrbUz1LlF2ln1s8BJ6wkrXCiqXT+kboRHznWd1NSXkbBL4Zf6oIS3OM7pbTOAviyIAPJzQNJ
5ecZPb9hXC99a1vZ3mzrYYjPeaqb3kUyvXzJ+p9atqHa8O6YIPYESGseKFiToDdzf3Z73wDQCqsN
NzCq/0VucSwUiKWYWXMUp1YwqIu7q4sLFmLZX1uKcnz0Y5QLl1gJuOp/gcK+L3PE3o1c1/ME/jmx
8jb2WVusMQ7kt2/a/IjxLM4DQqpXR2yKZf6nqNsaSfx740MZepxBvP64b0rzeCpsLqLDmrgmTAIM
DvTkfp4Xk9B9SARJSj8EKVq2XvHj+it0Qal56cdzQ83qBL24bo/4sI6EoFp8A7Lcd+Y09Tki1GEi
CRrFEwKL4qaGLAmuDi63Dn3g6dRbHQ9eQiL642dqSpjsUDdPUynEE8q9UydeQY78c5bT6z4E1aTL
pyD/SRMLrOoj/GSYhoTPir/NE7X77fb3IjnWnCLtD2SA1Sa7uWTFSphGOJyjLbGFjNoKqa+onqVT
p26C+EYzlV3aEuyG1QHjY8IxxS2ArtQktTrMPrUUWiQIIE0K76VNUdExnco82gJEkaU0TkLULwV3
gtrUE3+X8r3pmSaq6nXI+bn1XKVGeECWQ0sDD+O26pdKm1TrTrwQwZZfy2IaLzC1mOSr1UBigoSf
CyZOxuercY87+5Pebn1Ke5SodJaXvwe6KcWIE3wQ3FO+fBmeHYT2Y6Pa/haMkSNFmhwmS4TeNTve
3RvCnQWZjSVGbK2a9tO6RLbcfqd5fODKt7fOAQz5Y4IUU/OBAP4O268C/usp1YEFbQNzOchdR+2E
1T9eSAV9lNP0hZvWmDGEeL29Dg2lvEQreTki3CwcKSv8WuEuJuo793xulvcc34PUtce+S91M85O4
p6qbfd76idvj9XbCqe8+Y1qvkx8FsJGnrj88vl9Ynh5hbsAA/na13zLuhyP1CzUgLxZwztzbdcCN
EQgPHfwYDIpEQBx+wC8vd1ghZVH8N90fhGR55YX+Uv/yeCvjLkG1s3vSOcQJpJlR1TV8Mx7jVPjE
wY86Uoc5M8LgRDXs0+U4LjvhVtxQXCgYU83cbmwzawrMM+dERaxtI6i9v8cvA7eIKWq36q5+l+Hh
CLNStC5/yrBm4AvKzj2TmMI4RjMJ+EbR+D1pruqq1MEhVOt0ow08bHMugBgoT0Dv42JPMM/f++5P
I7u2hG7uvejNmLhSvh/QDSYbAwztMWQbsvQzB390/LO+92+7panqAfYcwVp3L1WP4WCxBPPNqUMu
qVk4UtgTWIXBzX0mwDOqVfxFAIWTjgEwxdbFFclBV0UMzW71GBIs/20+I5XT4CRVACNKBRVkjxBm
1nZjFTm4TZM4mj6ewVlpjRntYpeKKiak4xOuEDaL5nbYI0pekJurV43qJ8r/fEuXr1ziwdcgjhTZ
JJ9R87NwPrem3lUGj1i1+8cCjJFABJJdGKZCpAQ/V0gq8JqP7i5OdVzgGc0z9+NW6N3xu/SuaNKn
1zaHE9z/QLnDALTOQgNrnJlkQHNGEZmNH/r/QjZAvbYj2/KsH71mZzhnxpOFU+gBSk8SaX+oQwXv
pCZavv7SKz/cDl3OFMm/75z5vX1xFydqJZNJwS95jrhQ6uWQ6k+Ivny+h/doLIOdL3yPW7alizPT
sP6TfHy9d9Bd/yHhwKG8P0hXmtBc8NUJjEefvJOF6J0tXPZehgARVbxK0G3650XgLCGiaZql696B
JqqOJSH5X2mnNig2ny5Va59ex4+tICabmskW63lI/nkNhAV3pC5m8dAGAtFFvqMMJzl0fBmDM1J9
Y8vAl8WExqgpnyupM3xpq02lvFWkzTNNCxy47wB3cPmNrWEmPPCWTk22k2apyfVB81WixhwbfwWW
WT+efPDZ1i0zM8SLSk7X3ulgnoALGIqNi7BLF6kezty1imcAH1Djs+Hjm/PNJxsjkJ/kM160QEzI
WAGuiUydglQXbMSktZR8sZuEQn8UGKkvEZqpRQu1f2dmaS8pzUM/imG0wL4d4/1Rsl+MDNVCYtQ2
ITPF4AhzpKruonJSaeBpmguRuJWogXrH0+ocjaT5DnOjVbRJmBhPr246hd1wlZN7Ts/TssdgSrg/
Edft9MyeIQhMGQJjL9gI+VLwcfIgDg48dXi1O2xLo++l6qzh4NG+aH6K0XAj8YS1mitPKV5f18Pi
uJlzqAFVY9N7qZ9BxDSVhSNp9Zz0U/omhxBsd5NGGyTo0OjvrJ1Fhuazw+5X8+IePV2q8yk0N8dT
QoIkLnUtkDBc+c2EjeBnGvjHAH+hq09bAqdw9E2f7qLIYaq7uxg+jRxaMjwA9zAFlJWJNoDIexim
SL+bkvICHNTw4WP7DWcQnCnDHZyGBuo6Ceqx70Aq+wLeH18mC1WbWu5anG56WirYongMVVs7sFfv
vSyX/oIkMVq7JlXxUD/kYik9mwdGk7hCiJ85LHMVgIbGgfLKpxUlWsthFFDilFVOvwbZiFq3mf4Y
H55EnjNCe78XxWWOQUdPby9Zy0zCHGxjsNLOr0357/BoQRMlUq3wWz17vh05/QecZLLjuUScIBfQ
BWmyESYcuR+JB+8Fb4A/10AAlP28oL7F11Opv+SfySGwl4RpKgQ4AYv34D2sB60+TTQ5sVeOgR+g
NIMmMCWz2GNeeY/Z4mY2JNaMjG9wM5F6G5qOCRZuJvI2QoGLjVaFhLEfVvSWWO6S1AgufenicgeL
+fLnWORkVskEPdwQGqQMyfGU72bLsfEgW8stzL3pMo5OtS1Pwa80pjsJkJETp+hGN8vMT7JjSLbD
mQWAw/TNKJvbkhoM0TBgNRpXtI2Gtqad8WSx3fFWepH0Iq6DbrHwd9R6FEwkbc0ewMiEmpb3Sm9W
Okqx+ZzRDihQGrrHWtUfKDSyBfzfa9mz4LzAf6fmGxX9f7+Y4G+sngLUbqBjM0z5EiLz1uijZlBZ
KEzDmVH0DNgXynljt4jpQMsEajYotnF/RSCbf2R/JZTf1pHv7J/KAcFKpPj2lGc6+u0bHAPvQ9Hr
mAxCNI3nIsxPfe6nYXuI1SovuWWwYagD+/1SSvi32djEVRpcBSrR0ft5r6nl4uWBYTaEsdJjqZfD
3zMb6ip+mcUfbjybbZxIg/ZOoOIkoRgPgcuKIhIUKUSi7Vtk0JzfPyhZmcW+LEI1Rpf7f9Rb2MNE
XzAdS/RL9Dv4v6el7LnLSglVTe48WZHnDGplgGJhmjSJ5UUhUez0n5i2G4jh+TE2OGqKhKFAwYQb
XkjlGOjelXHrz85ubup99X2jWydMshy8aExYyDGgpFXKYmmH5rXbKtodimTTwoNHn82Mc5x3ZZMO
SeX81aMk569M3wWotG1Gr6GXgybelpa0oDYS7ND/kux/w1KTWsj3WEwByWW3BB8VB/wtOs4UhG9U
71c2+Qq7c118i1+W8xtbw2eD6O4fGMUIKO3w29dumZpJCqxJG10vn2juX7suFC2wLtkTyMSddGg8
3cZTKePBuKxjnU33Bu8MrmDtslQaXxBBdrt2+7uNy3aAfouQV2VHmo12KenvOo4ri04m9VsHABml
LY6fr1w9EocMTox/MQhGXjlMXJCtuMx8uGqiawmLhHk+N1mXhn97qOdC7k7kBwNvj4/G8wZUFFgN
6y5lHoFPcgHI3nr/XgdovfyTDbX6ctXVxllisT9t4s0nhACq5XH89cyAPrEs+FMbROJnAOE65Y10
cxrT6nhpRLmzFCvjptKIWGQYyKbd/0GwWLcFkzgVnTgxsGGftUo/ua7r6QU5qMYmVwprvGoB8UGp
XGbpLkPbs2kY1SnY3o+IpBImez9GuX3Hp1741gFN0u9HJqblQo/zyEJDVAHtQtECNw0i4z2mQ+7X
2z3gOxQtmF6tApBO1ke5LWXnCjTK73pe+RfEsI5VHKxIrQVJ4vg5OD7LsCqmbi3f2sDjjtz3ORbE
HrNf1cDbayVSob0qYidhwMxPrRRbxOghgBMNapL0tnLtyFKAtX71X2ZWtu0oUWW9kfTtc2gEuVuV
O+Cv06wVnTzF5qHeJIYvviFd4CvniOtkBDiPTyo0OGSwLtevIYx4HtPWq1pjMHjwkz1LBdjZlnCH
Jo5y5cl+RVjtBgfUeSyBvsekm1RcIvkRS1FhmMMN1rGbTxdO/6eN2KgWGm1M3zyvGztqLq1odJ5W
7/inBqsnpeCU+c6TWHsCkWyzt1Qf0eCMIgFSfGI1qjm0u+pQE6vgAJuhIXZ6B2/83bSuKKgpwMSE
UraL4fCUlN/LK+LoeH3D1jUEoaoWUwFsmU/qUCq3I34rqDaq4eLUMXFnNm9ZwRW1dzHjaIVgmnQL
gZ/GdCs/s2uxsF6HLWJI7Yt4NMQCS9jBQw4RWlAvSj95IXg8sLITWnyEMZcNpd2DnbJ0N+2t2dq2
xLOsoIiKZar++MoGN7Xc9ChgYsnwz9LTDubrsDF0On7WCpv42gWKBrPYY1NMKQ/a/CQ7MDBqT+nI
q34G0Znsvv3+hBxi+EWYdZzJYGvMDxbPM9gpBd+/0Al9/oRWxdyTM8lGR0sPlj2ZGjqWijwEdYh3
VBY6m3B/YAGYevAAciq9K/kwLdbfbsNSYTule/uWlRhuH3HP1wlWgLq09204Xbp29WFb6cX88nvC
R0zSOTlugZXbij2prwiDVmHye8/vvxxMyYuswKAVjO9VdogNa0Yu01dbcwJqcjubOZOuQeSPzVRG
5RHTYOIDQByTouWZr6mfy/2Q8TFZ74f3jvaQcbALu/cihYjoMCeHTUjgEwqKazxY5hig1rYwMALu
qTtE9P1FzyGnVEmKwJfKqnSsRyScp/XeDRhVVzkYlIu5+z6D4tUbd1jaWaD0a21PPRA/ixfORg08
ayoVs4iqsGtw6+Hw+xQvNznk+aNdKWffadAOAx1W9XMACUiuQzsdm6BrzYwWVt34Rp05zbGkftMX
uoUiGoBICBeOT5Ej7tEZG9szBZz57ThU/T8BtvgZCAQ4fayvnOcFrppGWrSqBjfwF4vFEruBVQff
ejW9ev6bLvUMgu7Y0dYoPr6H6k2Z6f38G0WtIwHXEyfYeCaWwHLT4miQaNEvCVb15+wL5R/C25fD
LIVlX3G4Asnxif+ieCYFXoSbemZLx+IkcTmUdzIFoH4bsjJZvzlZOBLarTKKG/FhTNjY1ztc2M/Y
7rG8BK+ru/iUWmWrhVv/jCznVCf7T9SyhRFbI1W9NZqiNuPY6WEDjEtGew2IeqcVO2rnYlqBQOXH
glsdK6cFn4y19xSfBZzbpKvZDiesLhGHz7idVf/1XM+90B40VQAo86/T5HFISdIv8J/lXtgPc7bd
LGb/mrVPCo9/Mb3kmVt8RSHrrjswunViX2UorufCvV8c/g/n1lhQFU31iEKLEGAXwYn3z13a+QN1
Ypxj9lehOIeLvWWcaWWnKv7tp4HEov3yvwcC900e340yO70xY3ZOUAB5m0PmH7kkg5NZ4CqFMb4j
5fh96gWWmhxJuCrtQ4Hu21Jql2fAYzO5FFUFRiyNW9GFEXErtipjywV5rCij//rmZ99p1plni43H
ZArZ2LiCd/aDag4CYJyogHhIy36gAfnP7UWNC7qic8rSBwKS49V++ur8iSXJKY9NUFNbPv+gSaRC
ULyXz1+OnUaQFN6eeXhZ110+K6QGrTxUExfu65LeCYAOi60gBhaItxJyHKcVQkYNp70cMOkL+WH2
2JlhrysDbPf2y70/hMRzIRjuQy/VJB0xYmnKuiPDKrp+Y64BOfeqkryxLT7bJP9phTvBdQJw/2O1
ZKpVUjiD64PlV/PPMFJMU6JUaojcInHEpDhHMstui2CxAcSeUmIKOq8krq9dUrV6puUKTeQrGim3
5ulAlspLjTj2yIBcRd1WKhvaleEG+AmqRScdnahkE9XZy2rOfU7nG7ruYwmLdK5ZjZ/SaabTyw0W
Bctbn9YIrjyEryS9Jm5LZ7BR8DdiQo0U7UfMabvm38Impa01YaIEtWtpkOX6cWIJM7qZY/SaT3dk
U3IN4Vm5JfdVnZUuQZDIqcZz837VqZ6RZUZheVd7OYIGjlr9QdWlgdKcjnw+5KLeMt5kHpdkT1Ab
0VavO2ENhD0Chqow44aRM0RqXY3cmuXriiRqxbQu/a4FNQ69D47lKZ2Lu2X2dPRte1PoDW4jTUev
BsFKRDUcgS6sh0/a/lTgn8KVW8MPnn1ciV9IZHoS0dtBorJ08JN1rQ36yaXhxMa3ownNzf8SCs3e
TDKXzIQGfZdckpZ+GJJ2rUC1pSLz3s1cXTzMegRE2sn8cmkLPhRJ6Ows5cGtAeXdrz3/NBeVarD1
MEpnlh+IlwkhiGtDyg2Gn1Sktq8wtevaSRDlK6P6NjeNWx16PIqzGFca5cnwKS3q92TCqP84sw1X
Rx+DLgyFL+iDnbAZSjYU4LUCBnOuD7oKs72qDzYfMkzZJ+i6tLd3jodD309yhCg8xgVhIcstNL8y
hVMzy0NlCCukTsWq4dWyy15Nb/9jxf/bsgyC/KBMJfKCM+QB6ZeNEqdKEtzNHpkIu7tMK21TuPPH
sXILt/YmdaH+hLN0F3g60EjcvFUlHG0PV43X2mtAmLNk6N/8Kn+iUmnMAyxzcCTinEu1pIz3sVhJ
kfHB+2LRNiJimqyl62XJYSOWzUldpBqaByeKOBNhOOk5dNwuhtsWKD45T0RsUSYWZZ9HolVhyeci
0xms5QKfX4wb8jgx+UOj38L8BbbBrR3E14yQeK31gsHoY7n/wdFo8Nhha+uFtHaDFJ/V0Cdg6kwB
Jd7QHFSsLNQlrQ7PrfnmmfLvU4t7mTdNt+WyisOFVW8S48EtPGYaap83eKstZpUjVII743xUONhR
wJBQscFP+/YwIBf3wZnK+iLY4BrPLqgtrKFT5DPWV3SFjDQspFL1rH0UfuWVx+4SVph99O91WXVK
yM5Aeb3t43iM0XFU618hR5N00GMgmgVm0u/5czb2c0A/zPkem6btF05nIYBx0UPWAE9ZD5bXLNRd
mAKm28IYjr0nWa6bgVHfkEO7BFvL5LeWGubpbUuD6WFpZwrYssrf0P88FHlilG3f5TzCYR80InhN
c+9I52/ToCVp3dGNXWsk9l+nCd5q+fqS5pofTAGJkH7Z8OIkVjcVOhi1/EY+CadI0w7cfvvFiBZa
hKjKFP/6K0dkr75y0EtEYPAcq6FlpvdM4BnuTpSkvsXpJyzOGfHeYWX8k2q7Jx+xOkDypIn57dGq
Ho5Br9Vrk/4qshbCWkoKA/cyONku0ec3iTijDr2pHE33PpJqb0w3yr3vdELy7yrQ3QrstwOjq7hv
FdJgvv35GduVUomipZqT4MTDCNjOp7DJ0etl1S6Y/qJg8PKQgP28N+Kog02XTuoW+MFktyRzyvtk
gIM3vLhVNAc15SV3+Lct7bohZ2H8AhvY2fV0KdA3YcklmBF0LE+FIXmS4XyjF9Gw9Law4fQMURoM
XSo+AbFx1nVt3pCz2qUJPSIm5OJPYO/dkpzYUbbxV+rBBKM4iuY87ao2VgkpkjAhLyoKYBcy+FrV
GfQStsZ8mJO/9BMwU634cKbvSrKlRUv9RxrK9vkGhBIgUes8GFpTH0x84oScmrpwd/QVb4EzlGSM
/iyzPRaYJHbHnq0JINJ4FN4C7Yk0hoVlyvIbKRBGYxaSYyTV+sf/fzxKYM6aKpHtq3mC0+UqgHwK
xK6GInxlOKq5QJyjkXfyOlrIuyxcGiDDqhrZMpQiNyfBce4iw4ONM7QpkhxJOJ8uPJ/h+YMLToyG
fLfPIicV0dT/mxeH0s4mR+NKCMczgPXSRBJ4n0KudYNIgexQiIyqjSGp/lbMp4xOsewD0oHlFXK9
9KJAfHUcQ2DjWCIhmTQZ2fU9CQPCbWAyuBnFzv5LLGK03Fk4ZgxJcHOvcXUkqGFk5J+9vUitIMS3
AhEwies3cAchMWNR2oqNhOMI/RbD8/6NH/d8okW5drOR23JMo2BytZs8K4xnGtXstw+NWHV5dVtf
Utr5z5wJbmkpPEsgBTDsZlmdNzaOZyggZxuLXnVkObVhHsJP+eV9g8rdl/2wYNG7Z0ocNUL0aeqa
0k3IC905Mahf1I7Vo/tdHcUozTe9HueugQfYr9q356YVElhgACQE8KCKFrZZ+W/6qkoyVzJBdwFZ
FVh22/aDiCfHdUNafutMKO6EAjqYm0kgtSObvKGxhJTF2KjirDVVcEsiJoeuKvW9UkhJjb7OZETr
A63kCMQ0NDve85OUwYwqbW1EZK3dDqCDS2lWJplsSEmoYcehxvMO69TpVBLp0VrJKezzctl3M/FQ
WExVdJKtN7s/Q7Bbayey7gWklerfSeC5MSqCB+qdO9As6SLo6VNltydWElk1UUq65uj//8NhRcuJ
EbA1I8/by+Gva3qHbE1UBZMPwLGxJ5exNjpC5bAD+KkB7/UPtJ1OAkiRu31DRQT3L9DOPdW8WxKa
pPfdSJnj02V/9KYG6JskaWgQoYRlVoxC2WQaoG3wFs5nXaygvI9zosoYaEG8AzEo5kdIsBWEm4gA
zZB59DakEkeT+Zanrl5vanUghOaAUuSujILSdLQr5TVaEoMte/TLcOWPhYmmzd3H+LgDX/5OevmL
UWBusMhvRNkHl+/sEBXkRNXjmRS7rWGLwqf0YKfwIXWmMa/aekraYLAzbekRcaTNB4ZFPg3+cZfr
sfAJGs+qnyiuEgunwK7CQPDqI1dZPjIldPExKFnill53joWoy8mPULwVTPD11KuWFZvOvqFvaNyx
Xix5oY89itLhUnJTcpcJDoaXQ7pMHZmz2TrQbR1L9YhPFRwxT2YHuzLbTr+uTFdiq8uACtHk7Tsz
mDfcduoz/NpbsIc02hfwvBNH40A9djZ1AVdIsy6yFIYwij9HnSW/ME1zGz6SAgrCe91L+1enCniA
4cPBRsdml2z8aamyDITOEzKjNK2XCGhcNOuiHP97L++dT6wPq9ORb1Tzcjv5Q/XG3gGz1vv4gMtP
uPg6ICgWqdkPZAPpnrVh6N55OPB9hSYe7TVTgPXprY2nJpogqRi93skMn9xJWj+9vZgrgsMxGG35
0IZdGXaCrieaPqXpNEHAryuZGf6RqWv5Mnyod/P8ZDy2mHM68ejvOtAo20WlQZ32Ql/eyW/qibjD
s9aCzqf4CyLhQwMt0R06pPsnxS6hMunJreSn7eCoEYa3wWR6xKlHR5B8XcY9VgOJIjYwUeYWPYAe
J8znHKcJIpq46vG0HpsQr6L3IOBB8hyKi4aiqo0TBbQIVJui4rBuq5f4W2TneLocscQBJDvSxo7/
2WliLShMdw7PY7wpgN/mIzdvsM4sujvQMLTpU7IdZqj2FHmdMnba+wh9AMdRbpSKPYSFV60TOw0j
d54I1231j6PrQh449f9KozOs0czAL/lhsPpdciZcQzqJkFISIb/zajpQzGTZwqDQ7rZbrvqTvwvG
J/gmWjrcvK90r98UmSSTqriaChjppWkzILfD/JuMUmXnqcZBsgHW3gA+YM8UQJmQIa8Nj8IGB+wx
Ls1SSvvkI4S8F8a9gmEi2N0xh6ZvNiVS5OjykG86gA11AIkijay1Pewx/D8vVbjp/WkTycsWZRaH
u9fFbQ9kXbQGjlteCm7mRSmPZ33e1fIah5Fk2x1eLsrLH8ycMEttxRtZNftnZLlRV3EdCFwOnaWd
TdG/uan6n7hSK01zb+o4GCZaM4vn/DuVYE/OkHuZcobJZPpCyswf3j9VPBUjA923Qmc1p5006s2t
Xv5tOV9KsRdbBGB6bUP4gWeUb9kJIC5CRjuUVCa8k6T7CKF4GTKM2xV2alLro1LZk0y6TEJ1K5CR
PdOTuGWq9EnMLgzmK9KAVtpt5TrEE3MV1Qeeor6OM2keOWUO6NMU/EPWPLgUbTTkQVWz/aL4ORA6
dqQAUkx0+9zYXf8rzfrvsyc5bgTG//Ikm/H89nxdBkt7ikmPHPGgCiXqyK4641Ui32G5oFCNlGph
+ZTlympal6eUpVt254Er31mWwCLG6fsHI+V0Q5Qj2SGnc95RDLKSTX95Nd8OgyneSYW3GMKxOXLK
YLp0aH4meRYlOpuH+tfSeVONl0QyvVyFbLGS+LhRzbn5/CzdUw0bFx73CFGH02kbcQzlqoKKwvqv
5k0Hp86YSb+1YpGQ5531U0mYPNGEQ0SxxlvbmPuX+jGdIaUCJ4w06JzvXZQ2mDw95vuGPPlRKgs9
cIoO+801dV3IlNnuQZh1S/eOr3zHMypHUmNIeKS4xa3LB/2tjTqQOQXNCAhlXcbrs2tWTccBO+dQ
yOXpdjUtwvXKRc7gzqPM3JSYv0lNjajbwmPH58sbL2jH3yJOE2vh4qKbiHdtLwRWTI8Oa7eiIVtm
BojROFDhsQv8lfKvHiwyrsX32VfQWRfrbdvVPDEYVjL14DEWwpUoKyKPry+Rr+JD4IJ3nh9OwCiY
sdCc7YA+LUQfFGCdEnp35C5zy0W4zkSPgHORl6ngcNcWd41JQQ64+/8iWUEViAXdSPgZ90d8tgjS
1Cq+FYpDigGGffsQaKnxsuq+CnBTPoyIom70hFAnYw/9N93Zym3VdSUzxTpED35SBtBzRcfdnSLS
EepFPlTyWPM6btYqekj52NzQlLYNk6XOTTcz2r7RTgw8o9gyxvFhXtvQBG7be/kqjOoIv18BU+5V
oketEh6sG4urVNavJKZJc2+Q3e1tNImCj6xP8Df79VCfH6+94Dt+1nqOnL33VX6sEANiTLgizen4
FwA5zc1sNai/6tsiK0yU3vso1on2qxIp9qmydCKJYEJMqqrvrT0WQCUwWOSaSrB3nsU3gh21ksd1
owoRr8uxBe9WimUKnOwUmcCWfaZcC30zEWLjUiC4mzEpK5V1YNe+/X9doPZhLsL0yXWp/vsy/6pb
ZbBYdE8pi574CQ7u/OzvsVg0a3hzWwVLl9/FqojCCrhnc5IgCuOu3X61N7wpQlmxcVbQEtl4vcnF
V9OiVOBgoBPGO7fqeWlBgRQfVEmFqsuk5cjnQz91RhLMoxhUUtO/asEfJX4m0+P37lgnCleLjdE/
mmcllgyveg6B00FN3zjHjiZASmWA/Twegy2Oda0qQiuQUE4fHiL7+KlJ4WostMfJx+HMDu5e/1az
Mf626YHtlrUbjcABsY1LYbNAXUTR6fLneVIR8fIatnX75yIOy5/TUuwIUaAtudPrTow6o8hBRdgs
O3tEEoQC5MlkrMS+ECiKxSOMOUtLTJF1TBDFYtaHI42y2xrlJzYfm3BpJKpbtonmshG+7KM963Bf
NGZpqnUvkb3frzCdegwLE4hZ3O6z578XibJtn7GCk4IUYo9QIS5RSDNv6vRCzgOO8D0dzD7vtfpB
p7Y1duKLpepMiNMhOlAR1Dozn9ki2y9njqkdJdvmhNJlOOZJ8eRZxhYYaiL/t0kUah4ai0p5NVC2
vieYVk906akahCYq/Orbbail0omHcBOKxPMgkj3hzxQTahiR4/rzodMX1yRE/12OkHKDMxnOuBY+
wl3AZDq+hru2dvrYFP74qMJi8G8mexbjZMclk6KPUsukR/frNmauwhke4cMzkohapTbbXWv/kc2v
2hTzjyG/uvPy8bWP56bt5Kn9zD1ovFUe/4I4uY4XUDIfdUCZC+xUz5GuTAksV86ailZAtnA0F0au
sUEp2iN27jXrSWKgevNOge+fBhD3+ZBnTrFq+c1lQaq7JayTotinkt618hS7/KL9IljzP+CvvqT0
1/bUnPOYZH4A2YS+6aT+ai35LjqgvOHIPllWyDGGkZMBPIdPkHqCBl7xLCiKoPvd/GxOx5GE5+0F
jMBGTdvYJr7bYAZY4WFSgtpesiMU/jcqkoumg/eGG6Tz9nfKyvQy9/jaF0OybfXsxb02SraszTfU
U2wU9Ytx8JdsfZcAdA3dPiy+SxJkELB0qKdnrWTsgU/fYsIjajL+u0EKnxBaYjH+m1B8ILa9Eduj
0ajO8XVx52tcAJDC2fW9XTyakm3xNIcA6u7la0nM/zr2uWLiKzdoRAN9gzE+oqgFqWKHiEkeeNq3
IWSQ5nAUgivHsdOnoPvwymihwcCn0OmbZTiEljjNBZZmqOGA6sO5isHsE77rvxoti9KP4oh92b56
ohF0nLVyDkgY1S4oSBHRFYSTzcs8T3YrOBDc102P3gD0P43zSY6mf0fPOSIPUjUYRvvDDayDsy8m
fntJQr6N4j6ZVVrPd+6DlpqT+Av+5GIfolyEj83hcxvT2QTTfZJyEqpjrPIIaHMVZU4blDgM6a+m
WEWlfmctBNhCL0KgnSSiXU7xon8w0t9bKfVp5jOs9JWWnlbQLtQljJjp5IExvSaFzOVSkHB2Bj+p
shBqKM7P9PTPEO7yiWPnEFGhMK8hm6ig0b2bleEJ0MfMCMLglrd/rLVbJbqrKB9A9zA7xkew1KCK
hJoOBt58/jo6rdx0UM69JOqyk5rZAFGrMK6dqPrbTVbnwR3AaQit4C80H1dext5bH3Lc5HxrE5rK
kKtOMZykeHKMTxZUZKvfyZCK75DxEkpVCfUEWCZtBBVdyNo1VvBqDUAowoESUoiVySJTZPEmtxR+
2VkEp02E6Omm9xuKvla/byhM7n70cyCH5ZDJ9C38q9zODNOgSb7yQg84lrfaVZq7c4eQs2AkgN7I
TyRiQRfnq/jjmKVNmSLb82/wTOHa0Blm7A+K7B3gj0ZNXGEgyXIDH3vWq8oIFlpgWjnUzDmJbENE
9ZuJjKjnNaKdWtMr4WV3L5Ckt3HsuuMFfjrHHXYgXs/JbATGlfnZqKbnl6oUKAKVE9tg30+sJhAP
3mLd0hms1HIpgG5LFwyYCazf1D6LwIadt6gjYA6Q8SMw74fdOShRE5AG9lqbYPS0NhcnBbYD58B1
zsYrQWZ/LY0GdbUGYWbED0FGha930cyBsXmBcrTS8MyTDjY1wraLzrLmTKdlt37CVr25GVaoQgBp
gGpWHEkLmwOlCa7IMdAWhHAyFFIoua7LQQ6j8YLplYlka6e+b+nrmQrN6T9ZZ0zlR2TsjPBDEypF
lOKXIwlpMYnuGpD2rcf+iSjt0n6od4310TI0okd+Gg0Hg0NestncQHyCXUMRd3/Ox2T/HoWfudj9
WaGSHklIN93UGoIfOP9ZxOi19hgrFLwq0mPv5fCQGEmQ2iyXWh3ZN+AYOSeJPKuLMOuRqXWRd9gn
uVEoWUkIy+JI7r8BkoVRqKSm9JthbCvt48l425hH1FUi4lGpPY6zAAqxhCyDVbszgSBYdRl9PEtR
7eAxTg1p8AYPvufp+8u7TU94NWwiuPBvJfMGaFpSc7CGc12qVGDDywLyxgesSZK8yulb8jIJEVTF
dYNevKrrQ3qojZJxogaPhASXSmbXepU7GiBRzoV7ItThS+qwE6EDy5lPESqm4lWF3n3yiKa92hbR
5hPIX5ZBYJZ9xhuwXeaWJdkbPqulGLOhZ5BoxWKN35wzYLf97vqO/D7zaFJ3VrErBvCYeGb4x6lj
UOVRj9I05Vd9gbaDVVTzq5+U51JJMIHBt+HaEmjdU+c/xGMBSOVGCEpAstioERvz5uFvyWL97oOK
2J3BPXM5ZuE4DbbhHvlIJ1FVAC/lkWWq+66RFkGE0pAvlAz01+OttydMv32gLfPuwrHA9umndUkE
qScjKfqGFg1Q+LQkhIAOcomd8QjZYb+Q55KIyiYypTDhrMzykAmlJYul915eqjZvYd4M++tkyHjk
LJ/36H1IMVdOvDn4q7rRJCFMK60MUiEbk4iZAO1yL6Ubk1g3y2zrSqpMWegBwqangE8T1G65ZVfQ
UfqJ7aOwMaD8727GqR1F6sfHwaGswGo++IS+EF1in9F4ZxlWR/uz3VYCJ907J6p/BdKZ7hTO4tec
gfIdZLL5LS71sZwDeZ4ddjmPUgcxc2qJ5iEhdL1GTHlh1/dywPDKMOnK8tbIfuW66Wzfjj+3gAf0
Xquqr/sjn39nuRvCFgNayQuKNLTYRSpZIOj0i8UVWLiifiw/2Rmt6sVxfAbIcGOWwUnVWBTKIe0f
cNcKz9bQcsg6251eb85N78ZBTFJjftaD1tUEP+p3ceQbk9XsYHIeYDsf4dF7ztPgSKlba8/FzWhD
A5OXgNZ3U1qr1QnjCi4FNLQAze5cDL7GxkES/UH2/jACNTXgOosAORg8HCYYQy5lAOQiQKw/7CBR
S4zdFhy+l8a0SQi+ucAfWqdERl8HKSKxDzmRQ+OGUPOO3kIomZ7NxnFi00jj/V80X8w2PBeoN7tn
GoTilYDx0IdmNte969ek0TpXeCl5/HB0nmqcosCWV8okSiZaOUo49ecTWJmI0DSjJ6BTDZVZxK1n
Wo0xY91b9ZGxBvkk24ecsE+od8eiAp9ax4RDx7AxgPzGPLDni2XL4Kre6NcBnuPWn0sfCElbbBHo
UmxFt3ax/ND+34pcSPKAwAeY08fwKNJjhHjRUBkLmpgC36KXLmUVErS/awNjnTnH3ujyK6A/L0bB
5szpy07X85R3jpd4fRcstQl98W/z6Zp87FyroUFPnAx6q3GPaF7u1nKvbWpYMNPQjE7DYYbviN1w
gsKFZAUYz6JSsWz6sit88FT/gQdRCACJ/rMNKt7LTvQmsRqPuO5Z6s6ZqI0K2y5p/57xmRBg2Y/w
EpjKObn00x0T1nYeZ58SppJiXRq9TCnkdbNJxz0dfgiyo+8PsluBHwX4kjBknWuR4qcKH7Fe2JYF
MQq4iLq6iQC2+03kEHc8hO7P/7lds3E5QbyGz6nokDC28dHCpNOZL5Joh4zyIp5WI/9zjgMIQu5L
oD0H5eip7ftsdQFjPIfRXLzzUqpRY3Lx1JFlfp1QqVT+8QMDCOt9QkPtLACb6Flf+bMbVaC/P+S+
0akocL1a9UzN0QQ/Mjotaj/M9UxG74NDKPbdjwySYPeIWl6HdvSsGeQuWvEXOulsbwT3JI2QCjxb
2TSYrkP4OlIOjtX1NafmrUCuiTBhJ/Ka+KWO/zxxjLE5cp1636QDRKb9z/fYA+pLEUwGvNLIbEyW
08rAgpCUmyBW040KKZs5s7FPOGcOP0hOMS9o9acQUJqXNLgPY83ZQwwE+OdmLLNu1KvgXp6MtW9a
u6KJmb622SR23qMo/B7lPNtpaRSAvNTdJnuygq/L/LbycpQjrkF5YInJ79e4kDXxgp6n2gxGvhqo
KZXeKFiyKqjtM5UyFeGTARlqr3VYpXrd/dXIrVDiIm0SdpY7guEyxEzd2eDbyBxXXNxcnoq7xJ8E
4TJeENaDGUq/ItnBAwYsjwEMF67thSWCY5I6AB89bHGvP8WDvC66SGWaaqNYCBIO04fsqtD0QsHI
sUiizHWYblaoP/gN22EPmaIWXcWbs0rIjf/r2LNKm5022gBa5Nj5cTyAJElJNfxloXYDBFuNQAdV
onMwYQfqjtTCxGcpZzuhY/m+s40CWbT+OrFxx4/25TaqG/Ql9FtnDNvpscznQuaAryZp9OHnj2QS
gSYVUyaXqA65QfmarffxfBA0pZumQp6+ChuyLTIbzFrxxDEpjDSDBQoyL8wYItPZutf7B9i5B4aQ
tVaLokbzTg80m75xj0ultDiJZFOtr1YhYLAXOqMzAkAcsXMUEKmgFpiaLBPi47PUAoc0gU6PLEat
IwTWXZMoREunZJHdRKrAXso5KwWJAKt1NG41SRnl23VMfcAxd5y8Jl3ppk0cMgZ5xCdJHOXk5Vpv
dKXSEkRQ5icigi+JG0yIdHZqpHmlayn5od9JkiBa5wFCqUJKzdBtyEXEq0PalLtTRwxFK3OwiOcG
nvXlNHdlcozG9JCH7hR0qQ4gSj9H5ppVLur61S/k1UHCNAnRJJIUIt8oTqr1Fozomak+/30jj6ro
07byFCEDAIaN+dwMAlqT6vc/HxZb023iRV8R5aukqddtNYsY/+OXtrrUgsV2Mgd4+dW+qZ712GNG
+RZdxSu49j+1poAuegm5z/fw6YsoJALo3xmA6sPHvON6fB1JNQvuWcEacuf2wUp9fnE8fMpnZa/i
qGjYG/UKVt5lfvB5l0gqIiEpiAr0OG01KZFJVgw49cJMcIjk4JFQaNx5S+QJ98PjOEty+pdUdpQ6
BhKa7sTNXTrs/z/mGNx3bB87HZ/j8MTgAGN5jQP3DqlsgAPNG16krcvA2mRqOyP/V+edKyfsUs5Q
ZBRo7wG6nzC5OI7HO6mxb3hAhueJFvKQrnCvmGq0dFdC+dN0kf/n76rYAxBfRHITxgXp0GSSp0B4
PWtJbNEuif7GeeW+9VkCX01KPcuzjULWHzxBUO4zvvd2gkLSOtF3ScZYjuGjE75XciThtLs3CQrL
zTnPvX6oRlANxFvaJgJynxNFN5YkL+SBwtwtgcPdWi5gO25atanMi/nXarPsXtyHoDP8jHnSG9aj
HGqS1aQXij+LRgE9CCX6BFvSCSPucDUtESz4bzrZvfJBiRzimd7ePCtSZGWLGwFq6p1l5X3phlbw
EjOJhQp/bXyjNLa7d82orOf1tWeTj9JVJTPPmpe1mn6RqBiJogak4U8S4ZQsvzhMonBfTOLWW/LK
7CzWVbxYnZxMrvIVLpgwCs9sPAZOX2xtToOLrzAa2pylLztKtPtH0UMq3WGAOqH9uNQcLshgoraN
NQ05AqL2hv6sscC6v9M3Wc/PV3QiTZRo2pQaCcRiPH9kvZY9hStlaPtH62I5xVhrOub3Dw4DCGbx
rBmVqJamoHDIxodHP5YUp6h07WAhZcPtxqGG2sUNusbCa84Z/y/Dhz2UFUHD/U4F76wQMU0RY3sF
MpE6INJWLeO8PAToMjb9+yDCVAyOBhZqt8nBHA8tTMXpaR+yaWD8nmVW2qJchz6ZkMKXpari22ce
Rujw3cFCQ45CejPd2zkxXRcpPtdWgoBeE/83PNIb8lKZIOu86ao1kcRwLP/6RIF0i4TBHJQPpoJf
au4B8q5ahdZdEZiWREYdlCFc9kKBmAw8NMr+w6fChoPMCeZaLwVRtP4jt6ZkFrOY6QZQhhgZ70ub
KS5XQkDiAXME8F3iIEySXwPBA7yIhE7zhcNpgSdIL3Du866PE5sPpTT5eoG6T8mr5Srpws7TNuRL
xQT0QtpgCeqUXc4c6PRsCRGZVpLmJf5DRzzePqnGNOKo6Bgxrbt95LhbVIbXsEUPViFlkBgg0EW6
3tFRIm55VvIu8ZvMmopK0qKv/Ln10kxcVAwYu3f90JBD26X6HAM9iDeM62XxSfF6+llBp5GeMs/H
2YXm0rNh7NEF4ezp7AegKwTu4PfsuUfwZnWyQzxThBQQSaM3FxqxLpJK6AOaqrAT0Iobu/y0P4IY
GMMQsaJ8Lx8p+ehoaFA/IpajWu2DU7xLWOfKWxYY1SD992hYWp4UbxQEvGLuB7cUqt7f4CtFTf6D
RzHhrxl286KOsUYHLRK+MXxdlBTo3MTKgkQL94UuKZs0KI5Lp7Kh8xGzeDkpYqT//oQqB3Xsu3KS
QicDUIEIzWSfP28T1O8f1WeNl0fKNjsR/0o8RELadvmT+cKyAOkMyUlB48ONG/ngNtv7XizcADlC
WHmwjS1CkqODQfZhah2vrD92KaY8tPmJkWAp1HF4suznALHe1wFRtpxAyW69xVy+uT0wJEdVn81B
D+d42DG0u5MK0PwY1DXCTJ6d0UUz+lV7HiUv82qmV6w43as5DuMPGBairGcIGRRYuFKBOTwruz3T
HQSqIy31/R8DWaNgSyACnbQu4vrzSsMxSQczKuW6b2EmFBqszWthnJLVdc6krt2qrSP35rZK+62d
EXA4OnIQLYyR7XslFYCLtxjNcCmcJOQ6swZAifeu/pWcCQ30dR8mMkUqHpkRW9nN/eNzz/nP+d+1
TgXCl0C7cxUeyJKdzPxESl60AR5YXTUT9BmtoXaXlSXwFJIWWA3JW32wsFcfMl0cbx44Jt9xM5xs
/JCC87odJrkh8k0U14bLWirV2Yn4weYDoqmGw/R4BbcpoxiSKZlRpMy5IMAgRjcoUiAHQImvth4L
TEu+2BvZ59s8roQrBSJmQIXFjM+reyG1WCNJXYxy07X1v8rky6U7bqptohFTvTJNwqP9Qi8+vsEw
yE+rNIXjSWtkjcH0kEB5qQn7j08GTqLUj/q4TSZghTgXWp057X9j5X2J5nTwO2ZmXFOdDaJIsWB0
bMyrfKhETiVMXs5fURs2sEr7ibSqO3cLD876ta681hGaNNmwIdRgg0odh2R123YQqawpqB7lac8n
bZQsNdUaPW+w/N/9irun5Vq7HlXmbOVn1J7DH4/rmvDUZSnSm8izfGYsaTv+X3OgmjeVS9nBT15u
4GjshawE/WlSHUIFP3HRlQ4gu6l6SCKSEE6fJRR2VlZSkhFzkoRb8n3MUbZXZ0SpvAKvyJ7ZwYyh
GnHIt4TxKUCbQCi4aWu5nu5KVOuFQk806uhGDSsL+Vk8Z1y3rCJ8RvThC7RS0XAX1fyK8oquj5I+
Yl0R/rB1IBiWfUiP46wF0FxnFWf7MLDFPWSw6eF65NWTMBqj5ZOOG43MbQwNN0Yi4HoFEJuvvaU1
SclV+3Nh8uxmqtVBupjVmUJeK3OGz7l7sZr/eVlX/w78T40kOIwdx072nRr3ZwSpVP8B/uqciOUa
OALUSJYwo9I29kKEpIqMi70er9aQenxlHwuiPi4rqI7EuUVbUIdUF1fZnhbcvl0uV2eVyMXCdOx5
UbK+aG/VDv/Pu5SuckqCnE/eZ+5Q9jTdJEcZ6fpi0W1OqNjDQbUTsbUyrjsnHVmsWxLywo58Ac60
jZQFIAuPyLkZAQ0MVpmCwuwCKEuf2U95PzckC4TXCWMUoXblM5GXe+xt3r67gSYQj1/EJnDJgs5S
lvJMlOcGgyV8iV/6dQVNdsK/Ttp3l5feds4aVHES9/lt/ggPt6xx2VZFJxLCD46xInImKYgCd1i3
7rwHSYVL/r/MXZ3isi6HppBf3Da90cC9pvXNHs70JT+GO4Xjp7yqcvIwEO4YZkB+yj8tOpTNZqsD
7vuWX26marBxvhX0kREeC5yWvdhOz7voJ64Y1QVDCIEgtJOKixlLMdAbBkxidRzoSZLGZkxXsLsR
MmrkgUeobHWcB6cZoZCiDniV1zouVh6SD6aH74tMiuFvhCbeqw9OrMGDg+jBdX4METJtkH1Q+US8
Vaa0ZM92Hr1wrHsL1CLjYl8kXthuDokgSTeBd68dJ/Bo9c48aSzYiM3hSfadcX7gmi2FZtntQe/K
r6hMIf09EB9IR2muzYPrZv0BYhRxMruYLdrTWL0YyDV1ej221BmYG6Kygbworsg3bzNkJ+XYlQ76
qkAum/KdX4/Y0vFopEXIGeokbPm9M6inK3xUPs2zwul2dfS8AxMpu7qjWV8iSscx1qiNy/0M/+G1
Y01XDRPv/DKBmU7b8bbiPMcPiyYQBZxBg2EkVa7wvkSfR2gxQZvtnngydLjRhlAViMTecf7e3x2N
UD6PkIJYLdjtjamX1pFhURNDtqJHEXDSlD6DpMeDm6tkXB1ux4GoWTzsEAIGvuJo7NcIDs/CJeL6
KWGknHeME/1bAilig45QzQGAj0jhKFiWCfYqyLbah3SW0tiyilDllOtQfArSNOWmtufMT3Qmqt/T
JkEaDOI+Ab1gJEvHCba5XwsjnR+yylwvRBJ0gmvQ/uYjxfkcNl+ZbMQr7PHPTakHKRQWOXTdGT4D
BVjh5bK38svM29GpJIFoo5L20CaJJ4Csft/grxU+hZ7ggxC0wXDqkwNHeZhsP5+alwDg/xjqxAkt
OYbFXCBevFqCkpDiRoHyf+gJJbjH4jdabyHGIApdNvRVscSiAFmyHZZnE+ao1XzVkZy4aNbqJ9F5
/TPxMfHfRWD+xPUaQ2w0X/3kEQZrfcddU/CvuOCeKB3iIoxqAdgwcKEd6KWNN23gkd0Sj54ZNtuG
MWRkyvYo/uatcUPuVpULGYEatRMXrvi0nlPRkzE4/kornr9ichQZHHYHYSCWTNuPMD2LrmygKwg+
y1ETD0wKzJRSDbMCr9vgVm8Ic54xheJMi9X5mu1DHSUaHZItu2RS+J6rA2XLfsDsFKjXftX2fZ9d
ADWnCFhSOIGuQS43RVAMEjaK5fV3WZ+HOcCPIjHZaxCWXV8AIj03sLc5jMkyIvlX3i93uB/FnN+q
mtIly4/d4MomOYpI+MbVJpqMHnVdfAmDlPQfNm4OI+52YRZJufTmV5aJagRREu9nszGnSme1kxuE
d4U+avpCaPWT3F+5REf7/GMfhg0r5zxWE3NY8j6IvzUWpcgeAWHiOAlBC0VhWlX6Vqw7N8Tx5Vud
K7HdcqxEKdBPKG+gm3zjXku010DRiZdJU8Mri83Qfl8zKadqjX1b8GapPT9xLh7wh0UjHbbJantb
JNa7zgcXHnC1pXCO6fkOA0ihLaRvHbWkOwawavYSJXzXzSqnEeUv5hxuvA0sNeOC+5MXlHZLsXq7
nON4CT4ka77KH8+VAbNkysqiXpqMzCklKR9hQCoch6bI6lxURkQcIrgStYTF+cFjJzND3vOtkuKc
d5C6BEnCuIEDJyRywXBlWyDzXMYak+53jqecK7rwxuspfQJZkzzQGAZTHtj/91c2asuSgcmYBF3j
FBaPq0DGopmuYUFmsMJS/lyTrc/oMl1ziquadKuKO7O2bsW70gQGkyd62k1fSoTx6WLIzUudCYMo
mp+MyTlsZ1YEGsY+6H1T8rGAqh34Fh+Z6A6hEDwRDLyCvgHkTp0IUoCmt4gC1NHE3zn5hJdd3y6B
i/COVle1IKObuvtY6Auht7LcgRlrOhQZWNTuLwSrPxvGEaWwo79Yj4G2n5afgh7EK57qvAQCzsAs
XvOMFrAQ7WGE5bH4bR3fGUcUZJpF3F+0Db5qfzDrWqL8uOVpZ7fBWd5XvWqkOAbHh5S4GsyuZ2az
TPFJDs6p5bnQKoAV2BrBUpiKkY85EqeApC2P7zuWcCE55B1yNzHpuIu14KGM/I7JHB092nzc7Z/3
bAaqkkLxD1ZB3gLTDB3u8Sh7SypUPD965uCcg6af+e90FigDv6SWloyCB6vS4xmLFaDBR/4U5slZ
r+1Ba8O4ofClVB6K90x+vdF2UjYvNgYv3bxhQp5/Zbv/uq0FkT5Hf5wRXgPYyArqOWg1P0oMHRy4
DpXaUUSe0QgSL83B0Yxfvd9pjrLNej5QqdZpy/rbXTalLH6AqP76yLlJaiF//QcQ5UzI49MUObvI
u4/+3ZdeXfGycWwHoBxUuBXCe5CU1R45BU2cJFV3jO4fSEBXMEp+bo+jZj6/ZpQN+xA57lNiqXcp
04lrrh770RXJ5tIKnBeyjP58hYpUSQtHqaJJLIEuE9IvccJ375jsu7BppdSPZvyloGZgyQOhOjCN
7pGwlA2oGHtlPts6GwTh2QloQ0ymftmomsZ1kjA6ZcsG5Ylrhv+Qi5YSYtA8RdCo5fjAtKN+5szC
aQMceHRTlEQdbGgQ+Nus/8dJAxeHmGrd7vRph3HcCnvHjhzR80TFQUnBtEWbEoP+HGwLRaX2NihD
FMune6k/ae7kZdI6K7FmB0dG84Z8gKWuK9lAoqPSzvRSgzCPxddH0DopuC1OBWzas+273spUy/Vs
QaBBZcBC3n8//iXvQrA/kjlTqGFf7ipbn4/y7j3Ks0qZC9TEAJzFx5UGQCOThDdvIltfuPuSScxD
ynU0OKGfycLdh6FFE7LQoXPp+XKITv7D8E3IXlkyapImL3yD+Q3/04fdlwOfLoFiEzXU6OG+wH3c
tCsA/zO06AEGCmtL7tdyDEFg8RwwBmPKyHFqGyjwAS7RMmawpWdWs49pJJhviyqpjbAi2X8xW6di
uu7/U64bHQ3Qv6uFSjxR0dJfonghj8e2+KTyDRLuMtEJAaXEEOOR/YmYSzswkZW9ozUZvaZ8UJed
ufKuSGVrFqw6K8oPWm02hJmKsp855VXRf54xbeNHl2V6G8hkepOK4bOhpILLOGhkI+SAY4kFX/KG
7m0gvKjMwFiMw/y0uxn2AUDARYIbJQPsjDduQSzVsNooY/HbhKibCUd1DwI4hVIM6eU4ajoAbnuE
KvayyRhsxVBYsHwiRCiB5vTKm/ili+R/LP8rjWJKJljj+ksGX7HaEzAB2bW1g+mgz3uvc3gbPgx6
qRaEDHgoKcaab6FpMTVLmk0tH2t4cv0m9CQzd0klkilwrmsX/uaVSxT350KKCexlGu57xn103SvB
qouP9IuZVNfeoKYMRSTXJm3ecfqPGS1makTMTXT+F5QQzn3JBOPwtuhiJbSZW6NZmszK2RpwPwVF
rJwOc1BmjdehC17lFGTyk6wU5raBLbEWQIgKseH8L320wjymG8qvoKHhInwOrnpgwaOmbXmdYl8D
U4u/Hrefp05PPVqEO/fMQEv5uV/2e/VJSW9MXk+TKNNTntp6TPf3lIMXh73EnTO1qhw1kph0SQPC
4v4Fm1tMmdCUTggC50GRieQ0msJhiNP2DCZ0Hl6U1IqQHLlp9Y2jLKDVwlNrTHKf1ckDQMiwR/xJ
7Nv9KCHxFkpti1Q1fWkclQcoh6vrLbOjvNM3auTBsTyYyGJEwn7YSRqeOzNfgec3j5RX85eHrrm0
2yXppDlDwbH01wLPIMAM4LZIrKbuiVGS7+hcthCI7cQhYZydh/ewBHFNYR8X9PsY4s47LYE+DknU
8iHsIA0042m5qd26u7EKJy1Vy72I16Wiju0bHz1uMnGQaKQILtWOVsE06dOuuf+15qjwcgZJt6qd
cDjXkxbgLohC0dbaukGEfMZ8OSEA24RozP+Syd4oih2u92s2zcZAhlH4izVQNOpIVSLh5Jp4RENf
t4iPJyEmS/nAaGID2uZAB3UKG7h92w1J6TlTbnJ348YDJPZ141nnq3wTPI8j3HZWpY+eLp++oXl2
bEAmkQF7iY2wFv0L/cAcf+XUpOg3CiTb/a1EhrclfgssATlZtAduza5MIBO93gOoC+swzn4pIHoS
coSR/tFuiXqlFx31G/NUmg5anHQEf1Gbpvq6Bq5TbuwmsIlJPobkv/d0Of5gUqWB79gql16K+J+a
usbJayHvtRAW2wUiPTNGL4GGiOCjklzMSwCyknGKtZzUpJDO3y2W8oskmfKPuomN6RPajB/zrXNO
Is0EhHIzw3weZLDVlO6Txcu6mVaUtBIK1RBmzgqnjrm/VqMFKV67Y7zyAZMk5CLb0YIbDByQZQwL
3oypNFgGho6/lTE99ugszg45u8oWsdIdT2PPhKMQzbzyu95OoFiZhgKnSG3Ao7b2LnXZm5eWMz2a
IjXO9TWqCfh1KgeG+O0Kf45k4syDObm7qxh89iTUA2yJSlmlH4FXhbsp+aIfOMzIFSK+k1O2Lw27
bDpD4STAXpPpavn3RaI7EJp2SIDxbDbMUF/g/y3q2+Ykw4+GnjthxGu1siTjjuM8Fr8cTsX3DvGh
yeWz5Hqr3mjH6a/CgVPbHyFprBh0aG6teY5VCsQx6XM7GW+duNOuZgHwlDbjoPgO+TmXYQWXWzGK
mNEFPAsWeXSFJQdtOtXQsgBR9es8Fx3pzLgAARjMWahr5GBry9c0UHMP+sCsFEhIUfKf/EnOpsx3
0xTM3NZFu4rN6uqL9lZIIbGZQv/VpphGO2byaS1a6lc2V+hh3HMzODyB9+SCFpKLvHgt1ahhL5jS
QMpkxOZrt8738L0YsEk+s3bkM+yQnLahyhmylBkcOYwsRISH3j2q0Q4hJZVzXYHV9D8u1jv5m7p5
D3fdTrMSUBS/UPTiPdU7sI+e26QpKGourzExrEspsEIdCc8neVWi4I/2ZOxEeoUy4EJYbCZWRuld
nZlFjuPFCbT2z91r/ZGpozzOPzD3Z1Y7bysv1woUo/+Hu/AKn/XqcA3rHHR4uzgsRpgf90nByF+D
8zd9NWKQcSuQXweK60jOBEeBXS1qYdClVUtwWI56327SNjxYm0jqDGv0U9c3R29pjXywCDLqpLli
Gp14G2IoFiQT5qn77x9gc/jUW9cgsmgjIadzkq3oPD9ce+xrM06ik9AFfh4usqyvU93yipYRTJIh
M9FXbXQaYEPkTP0xwRSvjARaUgaHsUlbnzum6r6eUU8+QUlnX2NNO4ceQyuSakOXL5ivcs61f5QG
ywffTv/16iS+Gm0rafysITBwS99hLA3UPaXUI8TQYSvzQRBkSCI9+Cj6ZkO3eneilOHRx6LB+Zgg
dWpE/Y23qDDzx6PNc+w6i39ddewrE9aHAIbfbzcb7Ron/vs3KY/VMnJ3FX4Zj+1JNJwQQeMFc5gz
29gf8VpFykxps6dZ9xtcbk59ZRb6Mt6/0A+wrGJ9i2qPHPGQTr8xasH4ECCHHwRfKC3ROuIHsNc7
c/cXH4AWLmbYwMmsDITiHDF3L76NAlzYdNMJKTnqVUO5gt+TRMcp/pFiJ0NLzoPNKb1jURHjSfIH
phS2DvpfuSSFI4wQKwuJUO7zgwq46NRnnCAy+eak3ugnkgGkzMhckw+9y/8PmTeqtwLMmINQFRjX
+QJqc04KB55pgVsvqwO5n0RN5qUXqn2tXO8h0X6HiUc9D2+9YJKm2WliUIB9VC5OQbPGzO2bJqBy
e9uQ7bZx01+H3MGH+8VLzgtdX9utm3FI6shS1+fWf1hqCsDvOH897gkYl8mB7hAEBkIAFKb6HfoQ
ELLyL796qm2tv1RdZEmdBxyTURx5H+bZR/6CdRWPpajkgmUejXNjhEE8MmsGXEDbzbf0GaIGK4Jt
tUf06aYfAKSszNedoMQU+nBzgTTHGogp2ZYEthUCFTG4c00P3TChrqSsgP56GttTMpdSG0k5xMfv
m+s2Rj5hRhdlmll1jzMwus2p/gEqz9hI0E+VZV+5P6xW+JeeVfUx2X01K5u7gF7Wve6ERay7fqLS
iEQBEzNixBIKxQtW3WMulzVVhW5whoTtmrr4ZVDGziDmlnnjEo7fOcfvfeCRS3ieRaTdZBOP6Iei
TB3qBv5Oye1AJ6OBzXARWnHVHyV5ExMF7//kc9XlfO5LWW4akaJXOg6hV7Hxh7y/xXvPGg4qAXmd
nNnA5kptyPeqRiaqhVxM++E0akULMeSqtNG9stnEfi5ImP0KvbIDxp7Nge7iHY+sY3BmVLB7rLa0
Hw1vbfAWrurOazB3L+xGdRLYqqRHk0S1AXKnTq2ZRb66lDVjT7DL8GBgbbwvkmYTYjcw6h1WjwrB
2lRSEhflVbdEQoYWtlZvDPy6GZbuEVL2p6lcEVgbBNZqaniDc7Sjo517CV/Z0yMvR/YivusDIPg/
+AAb0Tn4N6U5h0eKGO7ECmC89K6rcZa6Z6Sx4KDFGf084zSAPK9eXZdz+j3Go1SgSJZJHEwNeq4Z
EB3u5dfXV4kEHsrP9027DH5toyti0qpMPY5IH90s0hjxLQ904KqbU4w3pQdAnH+eocmxj7T4Vp38
mN/bLamPK+0oHjt9iGICU7Qxj0DN7+2pCtxlmSzy2acjrhDckcLN9LqthM9FkuJ0DyO4p4Tfz2Oc
lgt+GDAUmiE50wzYHU40EHW1AGgw1dsbBrqKFXXE2tEYfSSqTAo9r6CudH/HtOBZHnG5Qh7u8PnT
eipSOLpDnaVAFvfUeiRdYJjav6URTbU4xOVa6ahqXdUWewtl2bZxkly7goiDn0+oaEnsOekvhE8t
jJ/XXIzVZyosxNtqTLGPZd4+hQ9tU4jOFtckLygtGMAEX6r7yiEtoViAQjeM/L8224LRa69CPgrw
IQ4sxb8NO22DkNIlWz8UARhKf42xbJoAY+L6O0rChKYK/6ExJuwf1y7Vff8980OIgj6wwWUpLWox
GMAnwtGXr4I+Ve7WUdLyhMjiVHr7uuHVR19yh9QPejvzKblRycs4HNeD4reInzJBqaiBU5ABRYV5
yR4N5uOtV0BhJr2SO14wZDGnk5RzKamFFL+FQitf+NO1SUvY3B1MipIK7hdocOFBnDbAD08S2dxN
TxRWA51pjdC64W1jPi6Ck2sGErTY0NLRihiDtl2ergT3HkVek//kNLtVBJxt6uAs3KgG4Y5f4t2L
ta3xQVDE7n+MeOwQO/jUK8oHkJ2WBhaWCn9gskA5V4VOqA2ApCm1yD0dbFrsxlrfKiDp2swVQXgw
aZSaOkSpeUIVbmViRdBr/aFM2y0XTDF2QVJDSmo4ZPyLugJwiUJS+IikPfbHHCyFnNxblTUQuWZK
j+gnkQXH4DhGwojt4M0VMMXPqj8uc8eoreN1QBdgoGJwBegrtmLRymqzZrOMY+QgjpHrsrL6GV+u
27FkpPWJpE7jRY2kNfw+KnHX0N9ftDUlpLml3tuE/6ijunJN1g6uTK5nrIuO5E2bbwu3/gLzhwKQ
JWTzNmby9QP3uPVHeLWwusFGiasjIvYG3IO5w/ys2naV7RB2HcoHkHzLTJngnOdhKxKCjAmZdXdf
U76G2WYi4qwo6NtakDV1YHoM5h3BMyqGJ32b4Z1AThgL5OOxaKVJsgJHiYWYTc/RVO5op2GkXAOP
xZnEXvoyT+p2I5QSi1yZJjDkFdHmUjvbCsjTC6ti1s8LkqW1SDUbartuHAR8Xcy+aS5XOkaKhKZs
3O7gI26jxWKcOZcVZFtn3Q0yiomaGu1ovlqvP572ag+5Ae55RXETJqUvhd6T5cK9ovOgSk4GEVha
wf/iZV29EI9vYhNQN30EMvRLbmSU8ByIoU7gpp2TgcebXHUvDQ61AmUG2YZ/gJ4PWoT82ps5/MFG
/lxZjUvsK1rT7+8CwllVDDi0j400PrzrigF+Jen04BeEsElk+pVqMcTH+2UqNwCWh3qHlWD7jooe
iwFRrh4+ZgIWXF6dDRmK0ex1tnCe7/rA9ffIp1xduOzL801iWUdjWrisbP5JrEZ3fRWtFIzNSLze
he7dvO5yFJSgWoqbgMfX8K33YxQwtJdVfdz97Ua23MzfjannhDMihDFgOhN7HkMfbR98HoRgoOPp
gkI1jO+R/SXu2l5ZWiB9nRvIpvxIou/fwVr+jwKeHhEhlaHWXutZ92l8IYy81klgDhBrCi2chAgz
cLIhjJmcErp29bVS9unVC/bT8ATRduO9hbUK1BJ0S6493b/T8p8vGFxYwhfwmmj0ElHXpq+NxjUA
arvCpRYz53ZoS1YHGptACzBFSTVRwrT5kagcvPI7cQTuAgoDBR0+Or54NZYQTk4dT3VrpqzZWyN1
6Zj45jGQuv5tztEKtUlbYrnmcGiKmg9lpKunDCvP4lJHGYo+G6MVfqXxowa73mWaoGVOGvmGMtmC
3XIFS9v8oSs0e0R02AYlQeJq6k+DHAcFn0Pq+VKwhpK1zBqKuYYvvQ4v87XnZXfBKKyqPfUf2PoY
t07vKgBKR+Nb8GyendMg17g9o/0cyn6g0Bgw1LUK6JLlhTfa0Si38hSsD6LPHZdatARY8B4UKOVo
WccloIf2I9ikQynJhtjr48xy2wIcfc+ggCzKcta2IKvoDITpUF+d8TPMQwHebD6kLPDpLvFrs8AX
dlUkHXMqvl/IZuG+nYBAbK0TGSPqHxsQz8Iqp3ynDAfPzYRL5lhkdyT/CRVwFw0yQwpu5ejoJXhS
d3EXmDxIPoUOUqORJamQKHczEcpcQGxKP9cKbgUvD7PlbYWIuUmUPCsuzpQj5M7HTbPaoggcjAwr
wEOfktFXSp1H25jyRONHSrzvZgI2ozK6BYnAzHz39TaHFpvdS4f7aqaCpWHxHIoM18lvBmU9+8Pn
J3XMFOIBCZMmM1lpR6WZ4PjwJlyzHnjn+4UgPXSrwG86BVsa0Jgx7+8YDid9C+VvNheDa4N/YJRA
WQV3Jc5gqGiVNhhKHWzaqPpit28itQ1OT1QU5k9Pyre7k1ErpruNbkw/LPt1lVEi2dOqRdMQS35Q
Jwuq5eJN/pqrrG/LYG9pcdBcrIX18nDAVgZA0r8/y/5cEqWuTjRgeONWbeg6Tlvexs3+oNN87ANt
yiHOpIgv/naRjIIQJCdi3B2eFlri461v+8MuLYaDipIslc2eQXHjJg/oDifv4bJdblqBP/8cASon
vCvSGZ8v9DKGggX1DamTqyV/3nq9vy/c+yh7R/A35PnyFTnV6Jjba/nMT5irRirk1TX+23ERnioY
ceyJZNyZFl/OFiocTwhnu1Js6R7njYxvgKe2ja3Y3FQl3d47mtzmdasB3Vo2RpmJe5bv3cojEkuo
2vZQOuZt8AAXLu3M/q41bknb5ymJ6IXdU4IKpmWlWA1Z+I4gLlmOH34/Ty2AvUWDtYwKk3qbzThS
T8gz2OjdrlcuZx0yOpcPSvzxtrUkdmmZ1RNcfD82mrGx7fcpk/8xAzrveRzNBTsT5G3ohV/ZgeE7
D5yN1qQwsPQwMWISq9/56M6B2/Kb9LO3UsifQC5f7CU9G5yl9f2T1HjTvxTrE3ir//wTwCoeAlRt
mlr73Aup6wncUghJdkYWFEVVWv51v3v+7VFMoqcN61gI6oGPrYaagom0xzxTs+lcz+5ZGlkujzIR
X0ryTdnWb5I8nc/KM9XUSkzwbsXA+QkuAl2vyIeIVGhzP5keXQ/aQA6/S7A14BG+kSzQH9vMuzkT
B6dPkPPZp8cfYG3VaT+2RLHsAeXjJXKbOTIEX9PnbXfrGD8PAyEFvSWpXAD55lb+chcl1CNNYy5s
Q3S0ZU0zTx+SI6Pg8pnfzGG3uGSo6lJjk6GRQG4ucRzCPtTb6oeDsmsQvwNs4YMwgOeqicWajuhR
iesHzbvK1t9OlxdDMHc6lkfEWKCk8jZlY78irHDc8XKqrhqdk+GWpZ8Fd1idGtFrEeKHUVoOrhgi
ecdLb1zkbqmipfmqtqkFuQ+70Q1MtKYUyCGzTDfNnbZfHY01x1tHYdsMu3LiQz3Q0WVa5o5ES40c
1RusLhJLX4wiufjl7IX3NzzuPQtd/GoRS8rI1xrJco+yBV0nadP88zh1dPbH2lmuPJetDbcho9vV
HLcj+jqpFZpIz2dLb8iENilHLXJ0oSZNmflSD6Ycvx8E31UpB7y8SPQO8LfI9Z9eIiOCR+40GBiH
neTzrx8r7wsgTUIEpXaUaBRHGIZDP87x2lcVQBA8MpbIDdaOnQRIl/CSA1AEtpJguotEnU8UjNKH
j3nEMqn0tuOXd9DugObN4eltrtih4b2Z25tC0mgK6Q8x2d8Ljsr97AEULeBVB+dx/z7svW+ot7N6
pi0z2auNhC3dKRzos9clMgBaK1K+NXeqS9IB5JMLm1B1xJ7Mpp8OSaahXdxubZGTM8ern7oXp2+x
QPHefuyh8oLOY7ceBsicQ7Gk4m6nhJ+EVCbW1LHiYCLAfBC69igNEAzHSHuOoAFaUTYPkY9HFps5
7DFD6wqZLiQA8DfmJYQtt1M2F9x6lcyh7MdiCfrmfimTs/pyQTrDuXoRJ9KyFNzZ+SLDl6ekvwWM
1NS9Br9EODLuu5SmoN0W2Lfz0Ijb42VsNOJ+U45y1AwRY8AKj7TD9X11C+ivL7086yoqW5ajXlGg
340SXCDE9fvFRd0Vu7k2mqKAAWbeSrpP/koeuN9cvBdHsQpCUqYfbH9MHxzbvJdiK/NgJOWSspu9
qXLD83jLgAwl8pFd3TLsOOBCGGMQGG9HQW5nnhLa9D9/w6ZRLtKvzgQy6RB1lL2aRa3Wq0Pp/GuP
11XqmZo1I9+QJNNH5b5SpFM36FoKYGhkzyVWrNz/KhfJsqx90q3DcSHr9eHiFUIYWvo70MXKveK5
OJH/O+iGGxJ0NExlcM2iM8wQqYp/Gq+G1e8RR7e409N7hnk8dDkKmcgLHYrZyApk4jCndVVyEf6f
VHZozaFGLcIoqMHJuP0yBC23wsnARlnIYEAMU63Fha1rtLT7QqPUylgoRsaapvpY4/0qGpaC1sU/
PIYztmNNrfmX3SiNWtpfD4t0qUVV42ehVq4TrMNeKHgCEroCVuDjMysG9JA95Q/LywjEUl2EMWFI
jPlz5mi00Q35O9zJRqlOCblaxg4fWp4IM3Wjq6LSaf1YxkN0Ay9GErVhHIgb8OdhI5lO+R5gWnly
cVxd2cz4sOMtyr+yAqIcIcQztzP8i5qQN8bSR5jVIVAIyL/oYlbd1FhQZaDbDtrkrafAf+1uDnip
Y7KgiFUBd6Y1cncaiS1zuxlwVhyi/2JrKYMXXfZAb/ZnzqqnquMvxtdqJaHt07xZJkYqy1KLoIcd
xZ66pchGfsI/eO4J88Z8yTgyxDTZMixdkCayhKNicI7xeBt+Hqr36VciugJPd+Spv23FnJUv+bl6
cba1jMExGs+uBQZv3o5QlyBifn7Bzt6uQ0Hvv4Al42PvNfifhbshe2uWloGzW5ox46QT0CGhrS1r
dbZNlrAmGCO2a6pZt7UBbnH5gCZ/U4iHJQqacYd656omcLKCJnXyIMpCCLxjxWf/CTRI0C5NDtak
MOuPdNMUt/90i9Sj7k1pPD02khf13G2qJvhbfOaVIFzgPas5jEdZioO6fPrKlNxSSeFEk5nyWycn
DooSjp64HbRnCc8fTDTkqu4TpOPFDZncLy62kSD6IHtUj0rvO27ZknT7CNyerICpbSF/Jk4phpi4
ZyAEsseXkRQqYgAcmMrt9lafbh5+kgi1IBhKgPUCPJqbJDdVlftePBDnnu4prz5KfZiOLD2L/ony
YASJPYUjSYz68ikgb/Dr62VJBHAU8N1yYV6NmSm+/PFWyKysTCkCJDRLktIvvxAhA2Hei7HKe2aS
gg7c1Jb2VyNqACM2vJG35FpXwWGYx6L3zfJVkTqIkaniC3Htj3kLgD+dzMJnc/v8ZSqzYZpPlF1l
744KE5ciP5910byjUMkZtKX0RxonrRiPqS/BtcOw+VD7gzLaDoCnqJiDqA58s4uMwd/I5ZPW4Ukr
Uh10ezZp9rA8Z9qBoZMQzDBuxYkb1TJx6KfBilaVmVEEv7dA1jiIP1GWCI1Y7AUJ7SBWcKMKaJBK
oIBRIpxjBqC+LHufqINy6muHwLcQ/lPzLeiCTBDAGs7L/MQcEhukuJbbqXzChknM8lhybVlBdI1s
ROVuDAjdSNKqbITvyBkXIAFlHfs0jpGDyu73E97eykIMcHq8EhRYf5V10ymfKZndUz8KGmb5GMx6
x4dZfGvhJATYxeuhG6v1fCZUSwnmFsB7Ar/WsgEAzpmED5omzGzYi9e1FMCnS/Qk41dRu7Caai0I
8U1r9GdeVvd4fzP0tL+E6HWdVlS+b1ZSev7E0Ge6DoKl/lj/2fFrdcl1BjryrDCzmGn8ZI6ignuJ
0TLg9Rw82CPACUfvk/DbGuxsyPJc7AWNKB/iV5Jp9P3SgT2lz1B5DWM93iLB8SW+bkClUs7FeXuO
h8YeFXBi3AaRNVh0yL26IgCPvwpfif7NY2TVGBSHhrZeDunPmeYW+syryh0gGvs8WUET+3Usm754
aszst2GO/RdxFIWBALAKP0qoIB9UVJ5M7Du9I3+PMYRZRbhQq+Fmi9HOIzeodFjFSRAkmfkE2DPl
isPuJua393mqUgSCtmNwlHgFLZXDMgiP/NnHQXT6TYyChMgV8Q9CnU8N/e/RphCuVXvJVYQ91g1Z
ly63pVXfB9XbBlcEcDsiGWCwilQdbJ34vw711xllyLzK1cWHNCKjUlCXMLRH1t1CobrbUG2FEQge
VK9uThiYHiyri3gYYG5wYTmeMSgGPn6wF+Us/rY/IF4+dlVyK5LGftCVW4sLSzmHZQnXMLyElTki
+EcFc5vFHxJXFBjjjv4OoZDQWYMxpxufboLoSFLXH1l6zIhl/1X/RtwFGVDhxR4uvj2jA9GH6dU4
KDQj7gGYleqi4Km9vObx8qBUVXvav3JfmejS5cvGxgEcD+iU1+5Fy4aWXdhNHXbInt4EFrubpfhQ
rqo20OMP0w9+KhkFb+9jzf6KzEBrgjLfmlj+w26Z9Ut5atDYKN7tP3zSUuLQKmTJOevprcsGqkQc
wERcZ//rQHf+662Ppa58BYNjxbeytAPlGXRh5UPLaM6/XZ0ai8vjK6pW1PNFIaVhQFQeOXdEarxK
1nSEWyXBd8O8CSynBxXXaoA/rwf+y5pdiPlXng51d7/6SNvB96rodv6gvaBJTxoafWtjCk/WnQg9
aNgbOdcatCBdImholXThRis/IKZCPGHEzUbF/No3nloTXfebS3Z+xAgg9/CoAgVhAgTEnHO/gMEc
FGnVWBQ0mD0VANwq6xxwoalpx804ReBG28w4lakemT+e72u2UU+IBsS8J1zKteo0dRbWgLNAhZN7
yjEG1imcVt+gEAtNfbeYUPFB9Sv88Y+O6lMvHoPwNIJ4cRtvDCcYGid16GV5Otup1hWqwI3geI7u
Vx8xAVtNoSnjqKZ9z1jCeRtsw/Y0qmpZ9FfUclOvPaqqNARn+dZz4HwL8Y44t767NlnuhZnTVP5N
q/uLAtZiabH2L/AhlliZ7djQ6+d1vPOlcIZQ5xI1axaucGXOJyChcAtDraqwb1ByqXXSyPdbflUJ
U+Prx3/IltP6uI3pmaP+whI7BkWezKgjhUrgjQODdk+eJUYlVu5lhluZn+vTELKvxVVC0Ss8M8Eo
yBhDrNo3gDUQkL/QCw6qtcBu+8Fv3cCzoSZGbUQm63z6DlcV7LvYXiTnnpFa/FMyTkRjOBtUp89S
LJ9AoqL4S3iZlq9uRjTtSy9fr8quhRpnuNfzDCYaboGEV7q0teJTKEshixEETqJJTGdolJDbh+8s
+vSZbkyMwW8gFFb9gqm4I5f2ssXZ2CEZQ5NPVC/uvLMXOB45V1p3pPSYA/vof0kFYNQlNd7FjdGP
jpK0N5VDjAK+KD+skHOF7LLL0R4zijE3W0xDagdqtCyy6OMuMVjp3NN1Rrcrw7Wg3kCUKwRDpqrB
1dhWXKaJWU8hzAGTOZxcxhnzG+ljk0kUZO62GDjzFYOC7i2iOxpX2xRXoORBXV/VYceP6Pz19UhZ
OlWVQJIPdyBQRNoQIogMC8Go2Lqn/L9un8lcvkzp9O2ywb9dKj52qlBLklRxQL1h8eFyAUrsxQMx
6X12YWMS2uFz53nPBz10tyFE+yRtCuqxQnGNjamN+PtGi+mY3ZS5HrFQ2Yu/Vmp1dxSKfT5rilFT
KH3CpraPehCtJZQiAewZGVoY+pyx/wLMqI0aSDShb2V7B1Umg3hP4U6o1fgWOue6Bue8lgybhj72
GDeJbsoNh1J0QROnCPIyAKin6+sLyihiH0KgDkasos9T0Ka2tKqhQHzxPbNqJ8Bj/1Tf9UL1ss0N
BT6M8G08h8WByASOojOCuOTMSalTc0k4qnOILoxPfBAJ+c6roohHKZbXsxy06iMufC0WdvMOK2km
H+vs4NeWJqDN850XLkLm3QQzCAFMgPhUOkXBi8wghnA7Enn7pQVCZI8KBmgdiAx/WQZSqQmnpfqu
wPeaLUMzLdmpqgTRLY6DqTTXTyrV/+5uIFKvM6u69dB3MLtYzI975RgvGWEd1/lresISdDlyE7Ag
4Wwsb31RagvSqnCv1bpyO1MLfzyXqDQJ/+9MRhxza+Kl22VLm0SQgl/C28uI/C0mla4R4Wo2IYTI
YlNgUu+Ben8WJ5GWmuMw9bSzAMHJFXJmj2qQcgbqs5zT7Ir5L9+t+hILKazAUhMlxxRCsnaCPTKM
SbbFQp8JF+765j05ioxpQnKkJxUlJMcMDFP2InaXDRj08J/LnxWcNGaP33ZrDMMz+BryLhIjHdr8
7YzpORTq//E9xkotQPFu1eKLM8UwAXLu03DtDaDIZo4h2r5OM6FVKNF8BA4Sra71C11sIpVuIdHq
WgYkfOs/Rk1AO6XOhs4HGt8ePVgDXYJO2Vs3pmY2zOCXSIkkuzAKiTBrLv2MaEMJ7E1Ia24bSCRj
6a0QXlBOiFrYgNP5OHc9vBqQTuhrX8OdLor1ZMmz61RuOwf6W7oolqgbgNqxcuQyDjr3snOZ+sYb
568imFs4fvwHA3xoVTONL9PFmAW1XSAmfogHjR/QYBw7R3Sn+207URLzoQsfRXoVN0rooW2fk6QM
Pv68GMJ/eOnNUoTW7aXMc75cIUZhEf6ip/NPWeloUPn3u5eiY46nS+ITORYfJtuPivHPjxHtBmml
JRBNVHPdStLMdXp+qExcNpOqALhwaToXMMPDxmcSX6UPeZ+IG/Is8k6HUx1KcKLukdB2xUzHPPYr
pGVVQeP1iMO8lrYA1KuFC8qf8sEGmdQXPoSKcDAYkGEKvSXHGjyt89ubsihGfuzf9Ksgrcn7RDeL
8lnjLGOlr9CMjRq4BsUaJumT7PoW6SdnnpoPlM+p/HAQng2QBiJ8cx5QaKv4FPFVO4rxBae8bCLz
aYtE4a7Lq2NvoPD3qJKIzQ9hQLvLH8codNIKUvbr+qksnZdj2ARHXoq8/zquoFfHSllWhdowaaGn
dOyudhXkW3p21Wi5Icwo9HBOYlp8y+icvXd58i/2o5tCFyGVFCj4j6jEloa5STx3qTpOJxWcLcES
/5+NJcinxxlikhk4R4X4CUsTPCoTbMLoyxjCwdPpKuS1ZEGd3M/LHqiYs/KLCsxpL2FfH2ADleUo
nC5cXjnRB+b33Cb5FMWiYDWUJ2a6YwJ9z9RIutnjUPmf99uZK2US6xLChBH4XjWD7zDWkvY8eMdB
lco9b97rgUq+qxXg8Onjr8YiWw1Dd29+D7QNHQFV6Ui1TFCprKSRMOa3+3CNGOIAf6LE4oF9noNk
Vshpwc51+5kYDJ6911E6z8qinzRI8gJiZUxYfCnYglEvItU/qz+ylmNyB4DVsSa4XIBzuxCRc+hG
ScZV2QdAUW9+YW3Z5IhWDwF0tTNZOoCiL6ATu8iO6E001ZrDwWSAPPeIXvZ/X7Kszb+YqbCgedgA
7iZ7v4MtH7dEGscX8SM1H/mT7ihWwO9ZyROZus8LNGFyDSF90tSbY6S/XLTLfWR8TF7k6EJnFEcK
o7RhbD74/RFCKvAoS4jDqjQOZoMTsH+fOkBJLSVy8Fn3a5HRqz5dO0DQYKKdm6EHDQ5XFmg0M5jN
vCzRCVUg/l8sYy6BePBeMbXj+NrNyYqB2DoX/TkRyzKOD/E3CIOZmcL05+LKtIlOzv+1LkHicUdu
yD0asWc/+S1VWH8GkMeKDLi42IT87DFtQDYSqSMnZE0nmvZ042R1ePEt93W5msWL8k2rkfQ560pC
optd3hOpJM7tCfzXm7yWiHPUKgxSVaqv4WjK4uZF0SfHp0tWQdpqdTVRn0EIfRxNLOAYe+NgIWPx
5BZD3NcQbpjITUFXv8icdeDVphkIZcDI9MQrV1zpm64qvdQnopIXOTuevo4IWIb5ZJ2JFxJT61t6
xMfD7qBVUypoAWhPzDBVmKqJbTgaBs5S5HM43CzxZ2XQe+QObJIxQhLJrrUzY1oXgygIVVVTCa7u
KrU52WlDnb3XY6uu12DrKquY9iwXNGMlzMx6nClllNihQYuKEZn61LcZe1lfczcTVJ01S2kmBM8e
3XXcwZnsu30x+H175dlGd9k3/f8igkHUx5mV7taa1PAKsaOH3BOF7dI6zqzBTY5Af6jKQTGH2EN5
XYumB54+kno0/sWEQDwFr/adFw66/P4ux3vCMIyAeXhcfny00NaRT69uN+pOednY+m7Mh2GHN+xj
vZx5IeZ+D7BIDR6LmPqXISYZiRvfv4NlFHndl5qPDcPRYLe6AHnAMaFWc0o9bnzcnEjs3Z2apwUn
GogluCur4JBFCDeHVZooV5h76eP4Iko2WZpxnj5xuWAdXhJwZ3tbkCg3WNHTO4s6XjCo+cmt2YwF
s+9YBYfE1oujvnsUYMdseYrnBg+G0Y7yT2V1sQNNjygqfvyhGuH7P+QUtp1DAirRcN/5gc/KOlgK
iA9qiRPDd357S9yjAwZoBJaDZ7dFwAtFLU+YxgTN733mFPTmKe4/DBzTD7dgQUSa0icBPnXWh18T
1zYVlR5MqtFgt/rm3IGJVoyfBc7IJkTCeGEbjovxxtnb68/c7wPSj775soU2siLfSdLMLikK9OIm
CSKy+am7w5TCAumYM7HuV/2HafMXGEJCB6tUSvOdZUNOWEngQDC/VRIkK76dt76kFmiQQBWsq7+N
kqruf7DS5z+g+U8bmLPVMv5NgRAE0pTrw+wfj9+7pOiPv2f5PAYPghONrFx4XURtIv9ik3oPA2qV
kOyaJ9a3Aw/QmtMWFBqiR4xXUa4yyGqqf0rD8Y3MFoZskIalulFZEZ+//x5MiLDdvOxSIB35Gk4C
zL4PwQjWFog1P1wyaTQh9qMPln+rCHM0bIqQyBeND9Sl5qaI7Rg0tvnmSzYekSqiyYhMk+9d83TI
fQkudKWniXngzuDk844O3+8xhsstJigzI3bZxuzplFzr3VkWlxkpCZGLojcelnUbroo5EWa8C+zW
CtpZ5pn4Ux3/zy0fbQrz6d5EYatS/tJMbds1VAuotqS0KUt/OxWlWef1fAMXXeHiEPgXsF5ids2P
8i+gHnz3EoiXdgkRDIe2iLJTwvnfQNWV0CT7hS0hSuZfWs1JKCKawbkzIgJMRQv+3mNaCWS0WD9y
01CyYlWezn6cXtVKeexl6oi9ROGICUdYGgWPJ9Xz6qwvwriGGrMjHXWIbLHFAChRw/Pa5qIpTRKG
T69doGfN9st3KLcvYxxRmz0VyUcPzpImD+RBcTOywd/+wTF986HXcabmW4VjhVIxMtTtxtQiIPlL
6d12oOzK6ifKW87M5vJs2m35IroQ2kDh8lpP4GbBOK5H9A05WSybgQHn3QL03oNGquo2HbmzfwdU
rKGCtYf6gEySHWYZfjApyviJD/Wky+Oby/f4SNbwMeFGztoTwbQJ/CoDQEYWFQOrtNoiPVfu1jIW
fm4XWL5FlxVg8tc9PL/JnwHemVML9Q7I2Oi2tZxMAxl5p7hOGV1/gpvtSTrLYGqxR9ht6G/vZIQc
XTvKN5sNRu6xW3BEyHcgekiJNTlKRJDe8O1zy7lzH+DGNLQiZBpVn2EiQtM5yHtegQDP2sPeVjm7
uW6qqb4J+ryjfibqTJBKLnaPJqFTEdzT1c+GB/b5eoW6npWjjhB5AnPLTXUqfZpmJpgYvtLZmXlz
iL481uY3lgUmxk+AE7mYbmlWnmJF3qgaqNWO1a0G+HmaphLkUS7sb9GkjnLDb98U+0qmflAVdwjl
TsfQBf+yTtyxFTKgXsfuoFGPhnuGzQnN+4kQxcBYlM4gBo1dyHbutAxO5Usu673LV5dSNr8LFfFe
ZnaZG2/Vj/JiQShP3IWwn8JORD0I+RGRt1pHZAm6jEVK3Qfg6F/VGs/yNeX9JbLK+DAtKFzHu4vI
58eGEVgAEX0ZixF+a62akYCuXpcs7dnOqoeYzf3RmCRMQ3kodhoDvfhNJCNcLAdfG7h5nR3kpXvD
EY4yrjOO4fcn1hc1YBpMl1rqyaLPC09ZLimAZtI+gKlR/PNMG1FcqPp7sWeV7lmcZ66dkno0DsDX
sycqWihIaeAx9piiFkqXx29nXuwg3II/NQcvTimdZtOciOTnaqhVREE5tD61Jp04V2DaHNtKCCs9
DiUs/L6IRafF2fb81stbjPS0NcsIEQDLOxMypZSEd7kNiQKkVBGe5Xc3DCfEdf1swKNxY2jqnCWE
ICzj1028CWZQ1wQHskOAXbjDdq16XMpJM9E8OoyL0b8SltbCygJD3dV9Q8kMSbwZNBrKa+4UT9Ik
XpcuJ5jf5oKDt0bdejM/RAayQ3JMg/ovlLExMkiHKFa4iuk50mnkz2943h0I3dh8h7VRbLwy4AUc
C/cY4Xratdokkbw+3PekvSh6eH8+3ZtwII0hqS/SGAJjx/Cq/JzZbRL0qD/dWQVmtsYbAvDmAW7B
SKd3izyO9V+1GzjG+Xy0oiKJZrDZB6er1DKTZncZ7WMFbptO2qD6hHD1yNT68VwX++cfbqjeH0H/
K9QqbvVdGnuf2XNj0C1UeDuRbJH0bB6Rkb7DJggc5H2JXO4DxDYFR0x6NDmSsnUyAQ7wQff45oto
PFE1sxLThrPH/mC8kNzBCwbNdiEheWO5lNYnPq2lhwJ/MGKjxtEFBNYN0zcsA13Y5xHIqP9T8fBv
GUwQiFBzf++vhcoi7/0u6dvFZpSSMTZ7uhpwiFVoe6MZ8HWolX8V1Tli1paSomOdUE55D1GOvZlt
CN/qTjDaVA17zNW+Lg9YEH5Dl7bI66qCSAgIYDsNIdPmt22ayJFGmH0w5f+0Ha+vQShzKBMccFn6
We0OzUZk4RmCkEcbYr2HyJQVfmFy2e4yAtADFzb6P/a6u1guz06WceKl9IhBwYj0qQKg3+241l6y
Ix2YFuk88Y8+MKJmPeWSt6v1mNRC4hbHHTfkgiDRHjM/NIMZodxeyfol40IKDVEWpPPEWp56vdy4
4AONDKN8creuw1iFdwCPsEp5+/igGZHQcPLBuPnHd66/yMPwn+AcgOeWG2nuNe4c0DSP74ou65HD
uVHP2Q8DJymwBmBYngLipq+wbQ4Dpq2gFLqXS+pCgAANX1OzHRoYqM+QOq9UI5AMqLHfxMtXi8zE
LC/P4hUwo0t2RZSu59kT43sQIzPiU14jPMZdShvT4aFa9LM3kMCYZPTiFiEZlmBqZpZM48kNPn5A
brFW0pTkZ3rRwCiSphpWDkzXod5YFRkj/5hjmXKjKFGZaCqKNh992WcZWzNRwlPBVwatnv6XlcvM
U6jYaLa8hZ37ejABfL5jofOtFw3s+AQ7Ra3J8XPK0rulIWWt44LMP92GYnFNPenPQp+BgPZ0a4lg
Oqb42o3bn5uuCZ+7nhcMzjPZkYo/9Fb9Vx0reRs9gULNdrKd6bdNdtp34Icp+wPESJQSX7Ah3jsZ
h0Qmm3tR7eAMxdiHk80U9pBH/LfJ3HXvTDr9xuI3PwVJpmPjpJdcAw3oA4hjpyTqlfi/FXjm7Y6S
As0qDbbmVhFnkvBWfyZeObmfib89kGle71luASL0TYBmBHwNg5SHG5KE/eeYPbu8RUsKioDIc0oj
b8ofFfceIxZiekP+rHurBY9YMvhDwWvzQaN38JN2QO+b7U0FuwiWM8FHy0YMOPq+D4Id3Xl3SMdW
WhObJlwoZcWgCp6JEo9Uc8xzfY13tFlpaDjLwu6F+aVGDK2YHiLohY287zPU4hsJn47LXYO3Mgsj
Z95qZBRpjU9LKQ2IxXw9xW489uCoZhjdcj6rafTA+QVrk4BaV/s6xDj5VWTkPAdbU2k/AuqwMK/R
oFjRyM5NNwZCg+3WeAW+9cqKuZ+L/sXYrRRxEQ7HZkGyOZBVwot8RsJQt59dOO93m32lnONXvXqt
99AYjLGwhX/M5ABCOX8nI5mNAbxM3AOOYSbLFBlNCchO/RptkN/ueqgX4Vr/VXEJXIHXQG6tDig3
OG693nrRivTGdthvJuc1SE5yobfI9s9CcuZN8+xK/r1fMK6m1ccG6EBBEH0d1M8J3pJyGg92UGmz
QWwaO/Cva7F/JWtghdRxYB/yKyolffIJc6Wwdw72hpdBYTcsFlqKj42diiNx393QA0l669y8voZy
XQWmxbHW3veUgcPcJmw54jhsDGrnu5N50sk3ep4ZtjAotGBP76xk57MHs+MLtq+k9hS9MarLRhSh
Ky1gN54y5jVI3+ilG38GcVnBN12MM+fiNKHSCe9s71paaqY+b0rjATF2hWOXp75Jn/M4wf3mUxJJ
ScB5vMSjEYbMPb/B/nv4Icsiz+hmuIhPX0ZEHn62NXxFjjF3YIdivxszzYORoAq2vsC1ELEtHnUr
tCPWMyzoMT0AD3FMxyLXNkldd0ZDOoDkL0KUZn+csMWuI2ukw3J/m+CUY5vskaSI5E9J3RJaHylP
i3EiJ2TcQec+O6PPab2Pva71dNQ4FlWiMRnVge0nxHur71OTxbiBJvzAmdK5M5OJGFCmu5UcQ8fS
usPpehXJ8bcHPS6XmXilK5LBq75RYuEzCbWpFnRxbOIXb8tbK+fKlAM+s5097i2abIqFV/kottvd
uONBhjNxU1AuazTvE2VB6M1ujUKfaC4pfGRr6Ue3mVOSpcoUxpyVZefOOaWtddDlGX7F8MKzVvGx
d63d3qeDZs7tIbe5MoSl1oPVwpAsEo0QD3kUKxNYH+KZ+4GVNyUVfYHwuExFTbL73X7Rhhns/xW+
NWBUCp40sy0nDLI0flgBR6geON6KFXrp7CDHX3BQkKiE2wAm1kXUwwCWoTNdqki0TklqNodaRu2N
47YI1hZ+sWsYBTndhpdCXVAI3b7JgfLNZqQEFrSm0aiIt9wZgFKdyEzyPJkKQdvpve4LhgdC5PMX
7XwJcVKcPkoNEbVa9L0MkpvsH0sVtYptVGT/mr+/dQZ9tVFIx+G5bq/5FocEcbi/w+O59TK7uAx+
U/sOBceqe+ll/c+0MFOefjEaTDISWou7kKV9Y3hZu0ujDvkpyKB3oqRsvq9P6yxfLBmcS0kX4TbV
QoC/80SV5UtE9/r/5GBPCgOJa7BUNlHYfH6TIbacHW9as8NsDYeXh98RJW3zc6863/xgz1XolqUw
uoP2Kr497gENR3VSJHr01m7WJkYXiVe0EX9wv+o7gqmOtLLXDVobV9SQluO6Cr8yNNBNVR2yFaVq
mfxSpnA9nMecSRFNqZPXPzdFOChAbpm0ZohPTJHdodMv7hthcUPlDCGNzKVCwjxg/jhk26VbgFC8
B9zdYrB9Gz2ylC1LktX67ismFJQcq7RhUh/s+EH16QGMStorGoWmH71BsJQnQEbHfSTn3flfK8oo
MWgo1CC4ZsHkmcdqBvU6mUZ8KynfDgHV/b5NlioclI39grkJIOdmKNsEofqe9KYE+mSE9pSSF+L4
5iCElYBR28pmBtZBy5TVNwY1Rlf/d3ASIa/aNOBnhWv8otZxJFZyYqHcpc0CT6ridCS72Aejgu3x
rmAHwsz0uSqXPYygoxkSa9pjAutigP7170MN4ME4uDVjspY5mRw4s1AOiVKZbf0scEV/mQfNGSXa
mMhvFz+zFLzmXk11jcBhAheP7wX+VYj3tQteofshbqC2A8T+JwPcV6P1b0Ym+LereSRDLivRzfLL
rpk6FOp21lH/hBXrkeFaVjpcF+T2KyyRfHBdduviDqpZvxhbJVkEilwf+EMXbJTU0h1sDRTurDJ/
pywfybj673Lg1Nq6tpa/GMlQib1BHwjPUBP5RN3mDgCyC2GbFJ/dPXktcVyjO+1O4U8F7mePwWiq
NYwPVgnN865tyaUALTpTvlN4VoDcPZCnCy4yl6eSxbJR/8Y5ePMzQ0oA+VNqFTZZ3mn0MJM6Fo5G
sSJOZ8LWNUxspP8PM3jtpThwTfwdTjsguMX9gbU0bPmH6YjVFo5HnEfyJNlQVzR45aszeAVARAME
+TjLCOc1/5N7tTgeADsDGVXeIrzqTySZMkvpy0TWVvPB5na/gQ3PF8vNzVCvbKSBM9Sqg7RXVKiF
roOLyPiwDDb/84xDRE99XNWmoP/LbhmMdzh9GYfKUu9ugkA5BqWblaJ95+DMrVNm0+mdqOy6CNED
ozFajvPXJEgEYvrpKbNBZ2Bxy3VCR2SKQmX//DV1mNUzj61yX4cXurEaSxbkBZ+sVIJ6tP/YhpW2
5ddmZM8tA8C08zO8ZiZbBARBF1Gbi4fy8TQZ3naxnVzavOrVfQsH25TTyjYMOfp1leYJvz3euq2j
dndsao2DHSZyfsJgQ8ly5L26QybtCAXlPI2MWalsXgTUDvJkaTsPbnVvJsxa20hVLMmCC3amnaLg
kbEM3QxZ4sGgwxvTh+xjQ3+OH5+7d85AUbSuECgPoFj3752HXgCGsvdfp8fnPtt5hXLvx3KB97eh
xLhV6Dk+Zb5fDyEXGLKuOWgOIoDh8+yPFFD0/4813lnjW8cnVrF11nUiOIobORyYnfOwuQa6dueK
ZnSPxTVvKazVijQKWUbFrpAvNE8kPVnJgHVCF7NwMYIu+dSNk3clNFClEq2R0TXaJRaABs/QjVDZ
YupFUNngcCdBr6dqITiRSCzBKrccLM4pa0DuuwlU+CZvxhZpnTk0juoF8HnweJ4NPM6I9WhsseNY
1qYbapIYuL4txktBFWtHhz3rmTqdM5JLAT+Wr7nbWBlh3c8fk89BNlCdoNOLJP1Y4DyZf7il+O5S
4GdYLh+pawhattVKbAy7aBNufpmbzeh0Dq5NgUXot0O1YNuLgo9YxiKX7TiDe9KnvATk8v//jBHN
JyPe3RT2IFsyqY/Q5qwjNwJ6IUUfCluWCsOVFXQAv1bOaTn2Q7QvAWxeFS58inCMdnkhmKNAjr4D
tLDgIQbAoyP1MalMKk3054xKiTGeZjb/jyPxrJKbDBu6edBV1tbsB2RrnQqJrGHnRs+eycZu3P2J
v27dzTmvN+1WzmCeRmWK0Yfm0BgeL0u/OF1FAAgkasuxO9E6eEu3g3arm8lt2VxYbEVeMdHBLFLd
Sw02qvnHdtwyy1qMpOEmuQqvv4cATLIZEd0NFAqBAqvcwHNizQJchbygN72TvFVi1LdZ6WZANJSu
s1q4zKr0esuy3Iu5k67txiDjArK0FxXBpJDbMPIv20H0FxAjFLeJJtqVoM6zJfQSMIKNAKxV0rZj
9gFO0x6/GZ/qY6kKkSe9LBjRUTB+IEq94qQCjp/n+mWfrdmTlgHYvBD9Esrl5yf3hbf/x+FRitnS
Wl+SG6y2xwZue6aXvrFCxLDKMfAnIvhgdYyEC/PQ4ZIFQODkJSRVb31isQXJ0F3yn/byEoFxfIL3
kTpZ3W2MetkUEA7f413tQDA/RF6LDSu8vU1sSgKG2lvkEK1vkhMOc6E/38OlEwCVlyZ9Bqy+vkaM
NVtlvLHnkbEVv15lnLlewJHVdTLq1Di5LgFDIfY+nG5rMAQ/qURSKxkZdD47dHrr80IY6EMxdoSd
WQqDdN1CqhtPR1g+tRC5r9TUqh7eJ2qKNILzK/EJJkX1sR0rnP7N7uHfbHymscVwEcQRfsUYaQNM
kVmyNzXAaioGcA6/MGyrYPLYcmMMmQfl25l7XWWj3N7Fgyfi6uxvIjDmXYrBz234FZ6Em9FaDnoV
nI/bLxZbD6+CTt+Sb33afptQ+qU9oN2rr2y9oZBhYhojrQORx7/wAufKELgiS7Tp/t+aSffrRuNf
1kxRRxSh5V0JpE5oSyKxdNM0B+lnJaX0mYAqnv4KwY1dpUtj2iLQkxHx0u5WRcmyWN33/M29AcdX
Fa58cX17mRAQkGnTA96Q6LjHp9L+CmMgb0IDBc6G0+fe13N1YCOrlnT2cZQTWpnimbZ7ahqMR6e5
ShI2m4Jdc6cV3jo1LZWtH5mHX1CKo8lGGxYJ+WgctK+2aj1ty5p4ncXsc5o273XPC3Yi/mWiYP8s
Hpd9PFnygYxfhbQ+LTRsz49mDFGkCbynVOo8e9iwfvS+46KDfN75pO4WeDeSd/Gf94Z7T3TY9iJD
NUQYCAbq2j5q6/OolX/xmHEeEON399JwFWh054nYfKgO8MFhqC9/T3kYBVf5A/gK2SQIq0unEw7/
zsleg04iP1zrDOeasX19ojUs73w/hJ+SdIe2NZQH9ig7WKpvA+K80CMfQIGYaShASfnfohPv/bck
H/JCid5agSpjZLM+p7HNtX8ULv1JajVCkswwkf4XG/LUk84z1aiO+IViuUJ7x1NYDe+1mXakNjxo
JiEIWTS6K2BaNihYoxUuW+Sd9fxp6soWnlSP0+XO6iVeDjzZiLznyYPeZby07WcWDxY/apnRqrtX
xcWtozuexBsjAA8z6AlHMWDJ+HcpMt9UOuS9aoFadwVtxXSHBXF+3PDhpLMouUJs+Lk/jFiukBpV
xmpqf5fXV1BOMV4rxtO0VvHyWyhfKB/BSlJ+kaF1RGN8gn8vaTXzPLUW2EANcq5ntwhOYz7vMLyn
JShVQT2iR+sUI8HROqSGPOVmrcSbTkTir1XgsJa6471m/0aZNDkRbKVReD+Z2uAB2HinCdrRV+K6
YWScFnITFX7zWtG2cfsZPjmlK64loqnIPMIgtmYqqlP4CnPXDYdlMfrpplJB0WCnHwLDjdBFYIBH
oJ9BgmE6CwTrDPMxTO81Mpb4ypU9hKvaV4Q8ILeU6+KekyxBVIlyglvRquu8zlvQ77liotg7oUtv
KUIcZbh9CIbmdry2G84fUeV8cNM3VlzoBmfG6HqwNPVUlcJPtxUgGXNgSRiW0L80r0NrlRR4Z/hy
MBVjV28oAXeM7ryoz9825dkYRJWlk+uFEnTWbZhW1hSHpriRnaj4m2CEpOVXzX2aemC5qUqssvip
xcwNZhEFleH7XxxU1qu5kBVQiiyPpCM8/CLxZWrzjF0sEJqMQi/shkHbmMl7aZrUjOxGKvSKCdNZ
y4R/kTPhs98g+oS8GXzxzPyg9o1Tw8BPhidck48eaAJbbrlmoQdaQFffCvgKwrtX5cqi6ae/od0i
EGpr+ZKJysaXtgFzAnCcLDUt6EgU3xvgmpCZiEpxsOMUhvaPrxjdHb4qS6l5QcpXERQTPJePKptH
J91rOsU7Y2N8MYG14k/tk67G+3Fqj0E2VKJUsmA9tWj4n+Cvj+2/UrqyBxXQb0euDjDfDPS7PEsA
QGOzLdJh4ZkJFrZRGGVHUVlpjF2JkwTNFRbAsUGCYKq+Dvu0omAqDj/ygY7B0EUv5tPe9aVrz7dU
lWaYbGFQDWen4OeMUUOtCeYfQa0ZhvPQ3qAKy37eC72R6A+Mb26J94rLlTls5IcAVky+2dvm6HHb
hX9tiZLgDw9ExU4GQngzTZjMwl3qe7gtvOlM3AuAPhJzdSTPvLTEn3w1McTmD6KOp+aGmHEeUksb
NVHpD2exVAlqimAZI/7QJAQtMiGmEdIOsEd2S+kjbx3J1LOPt+77BSPF+WbRSyps0I+4rOw8Nx0h
U5qokO1hfI1nS3gfNSuAGlO6QlRaaJP8pdY0akXColHXOu4GZLKHU9mvukVjonMxDV5+6q0loMkE
1eszZHkKipRTjMup9O33YpcOabA3KiomjrbTeULwLORIs03d1CUq1/SnQWP71R5KwykUnUUBhwpW
IC9U29Da20+4m+H+70QTXxl0EcKX/p5U3xIrRRas2z/YA4YkyWV/GByN69sb3wBIAZsSlG8sJYE6
HO8/1PsI3JQaPyNPyEtmUSSXxr9InjfwZ2Fd5lEdBajM1J/SdYZKz4+zhPnlSDQYCgRkG/Uig9ZT
zbvKdpHLYtARVUu8PUgOcGh7Fi9rjdKsoBLc1u42rQqbcinXkN+tKToTP+TF4YtenEMISZpAiJtj
e9TluQXDroCe9fVRbJtgJgtsptAKwOtW4OSSbOKKI7z7tcJHQ1Ms+Ko9Rcp3IcDpCrtQht0FqZSq
EUvC8vqO58ZnQFMOL89n9GCJkxlVVWG0YlIYfMRdDK35FERKrcIc6dKP54C4SQN6u8nETHWGgADX
2LDIVq32UTJvwMGzoOmHYYhOR6oIWTnYouKWXr8yKiAHYgov/JBx8jlPoBNQGT5In41YB64fKIaS
NPvcs1OkkSzQ7FXtTt6N29Wq+J2cTWhkLHAvKHk8gaOXKBDYDDXu8M6PX7CW+40d/MldYxxktTyy
pgZ4sHLctttqY1AjgAyc7F9MvqqxotUFefFiX5iEef8gCtc7EXr9D2Bl7NVcRn36Mr44x7miOEjT
WhZWDcOw7fHtmq3W+SiWeDO+jR7V9NlNLMKkTszyIvrKK1w5MJON0hVYpyXM5NFXm3l53nOhG9T3
AB2cVE5MInKGlRPOgacvEYvHJLByV+aKwtW9yZtzGqtYkVyD+5COvCQFbKHLRjiDU76QB2Tolrab
MbPmqHPNnyBzdZBjd1ZfYTIb7S3xWDLyfM3eNaawZENTzJqQzXM1TpZfNFpAlc7S1IxZ2y2lbJGP
ETBclxVASlX4n4IvZvOKgs6yYYpI3iWJs8y4uZmuMfavZBx525BH1XJO/qLW7xPufsrMyauHZmZk
a2iLwPEjjyKzZiaunAnHuxruWbSfSKEqMIYSWUvF0nu7b5Jl1qGRk0558KMkSPhRHRPKDc+7vjQW
LQC8rXGZqOc1r7ms5pC3D8e8pNi0H0mVB1nnHY05Cs4PrxV4DE2l51lb78+AFjst9FehdjKU2bb+
7WkPdpv92qskKqe5wz2O2pSLDTLvvXacP70LKpzssPOvYINbQqRSAEKgNoem4HurJnDVrSUQHgdl
0mWp4zbAz0BogTt9rQWRfbdj2lIWddD3mx6rsOuRe344tKFEjAQ6wfd6JNMQ1UTJvJsBCvo3atyv
0sOBH/FPiv0Y0P9qUqxXZjmHWj+9ZTMlk7sm9881NQS0zNB8izG/scI4p4bqVXV28E5djzJ0b7a6
Fy+NLo93inxKDM5X22bhdQ00NHIcHyZ8AzK7ym+d3f8DMe7N+BrWbfucs4k78A6oi/S/nhDHnCbX
Qp7xbecDh6O2eW2/Oj+eVW3w7IGDcZevISZ63tBiR6XJCEWe8js3jYdTwj2z9r+AR36EU9+uAju5
ho5u96sNblvIt011PIu/p8YxNhMq064YoGQIjY6EujDJ4gtPRknfsGdVBs03tkad49npvIv767Er
VLcjjWIcNieqjhmASPs/WDmckSWM0UbzrR0DFADULTNAIkDSvFZWOZE4OkL0Cao9wJu19Ca9BOBg
6P2UWYYuTVHNUmuH6g4A9WRXj9ouFiMsulDxTDDNzuOM2Vr3tOjrP9CgVgjsJngaycp6kgVmD8HG
G3vF40FWqHTN1LcftCQDDH7C8x4xnibgFh9r+HeSywitR0fEDj64noMD45WNQsDGAOgIoaDVe7eR
JSSkOEUZAWg1nHtsCxfGQE22HmnXHis2cutxx1ZrR0ZZMCwjRCmP7yTnv347YX1pc/2daJzyWEpq
tUiqMtMArktF1egvBLaI3a7bpxnB36mW5ZimunE9LZOoIq8b7qtv5UGoGCd9nxZ950OZoIbgg4Vn
aUiYJLtOEIhFKqvXp7yj9o1Zyc1dCPvPMK163DOsspcyVAhZPbE61fSwyMWYM+Q/ee73dVg9I9K8
YDfgAYIrZqkDCpxWi8Uh/iOiVavwrIl0AbpwMgC0uDUapNQ9QRVViz4DGp6lO6YGjvFSets/HWBP
ubBZGDaOw7vQ9HsOmxslTk8X448KEUiQ95OEJQkrlUJALxE4+0UBUtCBAwrZIJthVcYpztpdqsJh
C3l6Esucf4jaa2EWL05b2bTAVd9I9cLPIxyvIivf2dI69XeEWlZHyhUeBHL+yxVSfkRV44rmz6Mh
RZ+2QuI55nZARfUrfvQYFkN/NbLbYsQTlnU8xRnCSJ3xL2LWTFplsIRBCfomsF1MTGT62r/QK7dg
PVTosc3KQnoFCnIFY2NGO38tx2Slb4Q8dIWYx+BBs1w6kkWgdJI9qOmhVzFGmxEe7Zwr1o7KQB7r
psUvM6fKlilb2yXOGAsxeTIUaTESDqa6gORo73PH+5lwSjcRayap7G1jRIaAxmAmpb8fzh7Z293r
WfsecXTEFtpXS9y+2oKhBxwSprZoLu0i0aC01nPzs8ALIhZXWt47JOaPZmVbsE7gxWy64V62uNAp
HYDwQJKuUvKmYWJUodJV9fz42mS21CgJhrLnEVQL/sM0rzrcAZNOUPqjszICxe/zIl9W9buckIik
X2KVUs5HvSugMTGlzTnPthiMdc1tS4M+4umzidBP9uciaq/HClCYRfAalzgWqUz0mNwTKcS1L5gW
x9MxnRySX02do5/7zfGs8kqOBEGId5pDQjhDK60mbIaJWWmOYMjWJpJx3Lt5gIHMgttAre2ACy4j
GUCHIp0QbJGHUtREs3lWV65M7pDmEWiZk76QFMTd9zZP3309ePSJ0CNSXVM8p2Wt0z5moKiSKNIS
Bzb4RZx/Q2XJK1SduH6DJ4O42QGzYyBLodBxcp9s05bt03r2x0Q7XRaWEQg1KWXXUX7wEUtO14oG
fSKKZAQPeLGtxKDH0gHl3igpPvhVpQCXPykhP2e6RfzbAcLHFoJ+eYY3vjquxZPtdEOaSjmlXYX6
JwlhYn534KuUZbUanWLeoSKM5i+tzl5D+pXkq08uMSarER75exNLMj6RS18dI0Cge7NQaPgWkd+d
pGOiO14JR1jhHyvTIjnnw2tMOuRQH1GO0m1lFGZP9pSkTxADXF2wsvAePNlXP009R6PriypjFkPW
CPf9I3VNqDtt+0pOCVzq1XjCqiu1XKz73aLhPQ2L/NvQ544Yqw2E/R7sTAbFLJPga5jmvMhXtcCp
nJE1NSr5F+GnpnPbC+9TDqoZbUGdWmC0tY6cQY6CqZ2UAzfMCXyGa3qjWXmaAHkNhPFwzy75Fw7S
e60aZ42nXNwpNPjp1Nz4mRQ5ZycGveo/enarchE6bwwGqUHRgkt0URrutRxfp/c2Y2RnIsp/BZNw
I8zSrWOPwBDnBlv+d7kKtychtpPVv7ndLo2hWIJ11pcLxeur3dSwHYasvldpucIKWvMfu40QapeX
UJFwqxD9rekmkyy8w+avr4OPcbQ3jcqWhn0LZ0CREw/oiCD7f+na6fvPnVehJWP/d8WDAd3wXZ7N
I/DaJbyag7hJNBQjnGJgBbPKf2+HmonKfPrd+19kCy7bBlNztL5adgzTiIL0MFuyIId4pOqownV9
U2zFfF1BKgCEF/utayF1mFIc12OiPbHVBep59XSmv5/tQ55JgwmtusYYNw1HgKyObBbHyaiWZ0p5
i21pqrai6dhO8VEaDdx6sQpDPQZz7p4gzNjTIxKFGtYyJ6zrYsQABrvfzXjPbcwLtgNuZotWgwuA
/EIZnPzya09uEdabEEThBbzE++mAHKnMnWQZ82tHuuLKZvH/voaSzuhM4G6aHtAjb54lCU9haqhG
AnmVDjRog8m42ykfj6xiPVgmplU2kz5KewJQG/04rJorO4MFUqICgxUpPXIFdtv/EBzeEG8bes6h
nSjZE3tgxjwhYKrzh5P9e77X8hbWzPFbbUTDsH7ngn66hxic7Kx0VGqnNIplA2tjM8rrnTgLNADX
o64hdDeOtqDuuENwIX6bvSyAqJ/CbWuOwBUMgLpGfBzNTdsFHaAUtHJNFJpkWtijh1n+YQnOIZZ8
4311cwK/ds0VbIKaHrTIR3dIH7hw+tHZILneowdnn56iQ/wemA8U/JVPLcOc+5wwCSa5kBUPkKyJ
Mrgjx1ZZ530dfVdrOOuYFTk1fUTKPWBFZmVRubpNCBQqyy9brWcP9WCqwvlJiyZdFWJzleYHQ4qT
jlT+m8FDCB/PUxyhl3aHNo82IruaRpWGNA0r8W/jdHYj0U3c91uOtkSVB6lTCmBntUdjmrmpt3Ha
Lm/+xTiO2T//pU0qGNbdVTFyLhJ2FncdacozIorHENLfNfB0cMlR1Lsq6FNb5sNq4JNhJIsFd9zQ
NCLgT26c83eLWlk7RfWmZHqWSsqEJNuwBPGUwjJNHv7+FwgNEoSLHcnYmsYweRErglPTKWfNV1zL
nMRJoMfYM82dZN3lngXEaM8AwOcZaKakHUg85IqETPXHdrV3S+dt8ihcSM68YvBnhhqkOjhHpiWl
FkFMPBBptmzVUOgdfgyV1jY4nhHVORl4rKgCHZjnhkA0Pkx8w/raWUrXGdJ8D6+JQ1VEX50Lbv9b
uzIpkKXoRM1Tx2FuRgaVJjTURa2po8UOnL1b42gULlX75sm9bn2B92tn8B5SC705dlcr2lVEX56Q
XErF/i5nnJqlM0G5ZfBTEHFJkeM7TIHs5zuWpdWwFHbXILCTbCGKOHf7c2qlrHVvHZMWyhdJ9vDa
313vBWQ+4nJQqEfrfp+x0HTQxyJOobxjuLke+Wp7uynP7ly5O6Vf//4qTvDPgdD/uIHp6Fmdo8SZ
Np08Lq7AHpb7xMbq9JbW+iyIpkpq8oF2pKRVbd1HgHp8fht/aEj+EJdLgNvqg6dWEmH3NrC7Joqv
rPwpzqyWueKl0NrYxVrYABQZo9DHEL/b8Pq1CUJ9zpTWXMjsNORa5aH9Mt71gC+KPqaVDIEouvY1
3enGW7M3Abk9LijWVzF7Xom0sRJ1a1ysBhS7HqvE/06eUEYLTs7P2TiSuUnE+kit2ibIBVpipxT/
FZnwrOi2e6kIRLpz6BCycuAr36c7WwgLUgVTxFKjHJ3siqxd5akC5yQ99PRuMrUrUXFe3Bovu2KE
yd/lJzKvbv5FcwVU/1znt4Rj76q3/hZbcA3v4GgYZCrl0SIeG1FhZ6QRAt1Ewxm23awxL3RkbjeQ
FYE6ZwLl3yRS+LYuIbwNq6xeF0wa/aiuxmDqG3yRGl6WuQDBoQl7TxjvZg+mbIDvec4n14JG66gP
Rgdrhy6AMENvUf9daiSxzCa7kb9vRxHW599ss+Iks3bJAApcwaXrU0un/TEvgDnvbdC1Uaow7LHk
nDCYJEphS1rhNy/9jrhqrSyFCFOZve4MIbIXVhRAEqBI3/LVTqZqRRKTqMH+BfGT7slIFIruy8R1
ZQ/2iaXalOCal52DslvmTlKQ5wZSO7ZsMQhpsfo/imACO5OlvjcaIA7qFAXXGQPt567DypQnlZqS
axO0bCp0Fe66FmD12ZPF8UP1O3X05IAcc37n6cpyREabS/D1uLAnr7OXdu8iuuqhk/rhhPNTd297
AnRs37MZzQNSkl0aHcAGPvpKlsDuet+zBcO2VZ6cOagq2TIeoldnbMp0gtropTz71rcQaYtgm+Pq
HZWy0b0jvozbA5KcfcF6YcskVAYMnntZqWY8UO+anvoOOwd8i7fYJsa+fnwFr/tLvjdI9uyssDxL
Na/zT26gykuWl9lIM3BGLYPiqqNz3J447EkrE069XirSMX2sZQP6WNfIhcecyVLJkAlGyedpd4n4
vHZvdH5YjW3zf6tOYpARpp0PLhE1YybZCZladyaqhy6x/jXoE5z2XgfzuvXq8oZYhJUqIYSvr+lZ
a28RZcMWHwTiiWcuN34CtbXcRh/j46d46OHOcSMB2vtMAczm16pHWA+M6OwVT5Rr9myGTcPiN/Ha
8cfa8FsuUo16Q7W2dzC4pBaKme5ETN4rrHa0Uw2J3zJOZJCxW5+Tb+GUiwqpwDDWXvnYmM1Lwcrs
8NkiON+pacnU/M9gIp43TTtT2XDPB/ZOcO2U1hTy3Snf1PR0gbCvzL5pe8kdfvWeJHT4UwU7DyPu
Cyrgw5n00LWN4F+xX2hubEI06A5Jv9NXYFzT4Sl+Oj3SdQG+6uCtcIzN5ZOCLcspWGBVpKBI0aIn
BT+yHACAyBM3nPAHwzgC6oyEXpnRxnNZQ6WkvyyWdLz/jZB0kUXxvUInAR/imnBYAf0PgDNpq5oe
4MycpTdhxpXBO0ZqGOeh7H8gf94TU30hqY/bmkN2bgdu5DfPSck4kolljZS50GRBh5tZGydN08o7
FPiaQwN6kk37tjTX063acbYigxNN1ZdnrkJhO6NO2ICgZm4DNurREnQ5HKp0M125DwHuc801SwzL
SA/EmeKECacapb0heMUPENc3b9RsAkriGbDO36Bl6SaLCktMEMmdcQVtP4BIgVx+nvfEHSZ+7Inf
4zC7kxc1p0FlhFogwzOnCdTJFqp+i5aRzxoBHJEmArR0l7y0CVx9WpTvvQkr1wBoxDnjCE1j6qy3
+m/J6+mx0TclbXx7H4eZWqyGQxalPygfxhuvnz2tfIGy/i6QxigAthz/Bofy/7AAN3VDCTKOQHYR
shXLy2kf6WCFPV2gW6CvtLynMMxqv8N3bLPO4Wz1biOnGU/nU6GJ7toYUVUPyLdhI/U67LxoIoSx
ztU+9iVZZ+DpzAMokVe6JHTzWT1D6tCHG35Mic8YjBvx4lsINRI0EeOFh0HiFu72SHk8stXnsiRj
cA29+06+IOInN5PBD7kZb4QwmkA3lVFIZ4awQTdbgWOpqv+7pAE5M2EeixSwRM/c74Tazv91ZAiV
KUb0U9ux7HzmEC8HnV/6h8quXnL87Jc4FxMF6Z+WEoaZidvWxOztIayN0tssf8fBjq3/k82HNYTT
ejSP7Hi8VrdQzIZHw1hFlEdebywwNO4nOJRPetEUq3dqqPpTbxHBFpQGHO9G3Wmr3tc8n5GGZXSR
cDMU5T5f/fWrSePvD2XUNgjzaigXpJT30w+LpgK+gY+aQff11/kr1+FEl+pMtq4MbgePFGVGTe74
TtS8BGKuTp5i5Rrqn5cgzwVaFmazHt5DnpdDD2fdvbSd1c+P0p+ZRlqnlyEUDWWDndR0SW4V+lz0
3uJt9Q1MzTbB1XQJYq7LSCSHuN6WhqXBJ0TyhrxFBJI1C9svnO4Ec74SXMDMabaACEfNTTAA5OZJ
zHK8LIX0xePlNAhtQDOnSRdL0Tva44sLDN1gj0uM424M9T5cm7B2czO0GM41RjsWDj+vg7Rmmk9R
GO5I7A6AcMf9+dsiy4kWlJ6wX6DIOreLHvzqaA+7qEv/fHdhHmG9bajn8UFihX/VtaI9SJMOhFQD
ztIX8Ow3JRh7s6dbOXUvnGNGuUX5AwFkSDdC8GJzIwH+RvPNPrZdt/8K6RpHmKcxUlUVV4hUw5Qq
UpRprs+M4YJ3sw765LdwCiTw3TjDA6LI8sgsHbfSNFwsAV8BLzYjeQhwxpVziWaik8Ix0Nt1sXOr
torH7H3VIc4wMslOcUA5Nkb3O0F/KFBC+sXGXv62JHoZJJ6lsMOGEz09DQXRDEDJEHSH3DLWJ3H0
AwzDGdqR8qrdbeN0Abk6j2Ykwon+xlQgsMGatDyfjpSP74W4ptK69hg6g/fZWXbKEtCaj3jHcmre
P+wvozngeWOAJEaWdk4LjCHzEGndJsa6C5Ely/0UvYjkZPnqKX/tIzWlsZMPpHApGhzLUSQyNyuY
s483EMw99Jlyq2ZpEu69Dany/M/zao84PNulKb1Mq8SocXLAVQEmC/+TGUMncJKscr5IcerCFso5
H96zKVMF3zEiv2LgTW/HprmquzS09q6+DUKpO/X6PXBYVPoPCbNgxqnlhyDc9ltcSUOtjvIJAUdI
ct/3QoDHLqfGnTLaZi40/wH1CFAOW8KQsiNroDiqTl94xItRjoiUd7sl9Hbc+2a6vvixZYarBLmk
EH0FLa588642s3xUIdIkuS6D/t0RtJMoqsKvCazXxtdj2gMYGOSeJJE7nBwd1ZKvija4nJKUB/p5
+X+ZJHXBmP7h0S8lf+1DJgD+/fYm0WTlROBBO24/iPBBOet6d6o8J/ZWK326xQJv+ixucGQRVv+V
5zi8tcVeBs2zz8L5ixD4IlTj3DsJIirpDroRtWcCzx0s5nzUhMAeXWB2XUhl0C506yQckKPPsIbd
EgeutzCQpVDIijWGFbm8op2gjQjlgt/71wugGciqpYtaZUHMODQ0RBag86APXwEzpmcMnvNs8mkb
ZywKmSGM9odmUy2jdn3wVEW32EEf96dyUVSoULyLvFprIrDpElliyvtphI6jHUYplgWc7lzv0VQE
2A9Pdxi1q7MABDUaGVek/rdih1FwKWHSVLn3yFzn2Ytq1if4m2lfXaSrSPm+MWpElg3hMNSLbbBD
DqmjQsf6F6WKs7lDjaksWvlVVKwxtv7jzkEfphmbXgImvukFYpFqtIUkv/ie5Aw2PDBrahvZ/nM5
rCdZSYVVMBdC460bggeVhLByTd1pJZIRCTnyeSr83IVJ7/2gvRbmwhhJpTotVAtrep9UzAlBSutW
v/V0JMUJPBVymw/dKxekSNrY+G1Dw0s84H+UYQBVetR9XUzeeMJzDRs7T7JAMB27wu5PCnXfBB8T
3vr6q7XwGZCOCmA6axt+/vTVdiBAt6nM+j7qmUrzgLJQtv40Xxq/jdKAIgD/09DYOGQshyAV1ild
mulKZC/o4/z7TulFRglAeicDf2ZlVOIQG2shqXsxPc4fG+WlWlQVCL58UsDiXopFj28rXCePqZbf
ENIIB8ZjLjXT5KQ7OWkCqXNofjwsTMkeFY+dePgZgQaGnzNEqzSNP/ylxhBt9QXmvN7i0UGo0E1E
Y/yjHyQoddQD5GqwIE86v2DcFrjaP/OHnTHTOc4Qi+/UH17rD5IaaofP+N9UU5mEGbDaztKweS57
QX7d70NtNuAxwcbWFmQytG89teP2YfYyND+YT6Krx0nH48ra8e1NB9ZcKoBdJbu8uIU0yrxDx4fW
1ILDPFEaqAZELpg6lcyXPrB7dcB/F0LV7JpxZRLLbohPRyK2y5giRl3ah4ZM3erS3KYGUAozVpxV
E/RtTOPBr0QJ7IvfY+QmmEw7twaTEqlB3lreTQUKwx+fwPj7p3vDuzXagtbgivs/e7/mKwdHt8dL
dMqCo80zpOVS3cEVmVweS2b8x1IkI7ldsvBBhQzMmgFANChY+4j4VPQ9dHLOEfZBH/JJOFJ7lYvz
GDiqFjVFfbBlhbI/x+k/mA8vYC57xfRk0SOAzfpCVSMaIIsMj7Yrn9WjBFKQKrHzTpwVwp1M8ECV
xHcphNlYkTtE9fm7pyvkoj/xukeEhEqq0lxniUm1gWVDEnp2RbfikOWG3TjRlUJhINk1RaNih1g0
EnA3KoMDMZ+nQ34N2oN9yvIkNw1vhtmoZCO8SttTlmp+N01htozSZOE9Obu6k927+PmmUTmJC8nw
6d989BYQFciKTYr6tIxtmqaHE553FQS5p53Lz0UZKdMWle5XwaSI8DfBrSsSLzXOkjdO5WfilHBE
cZs+d2HavJNWB975tQUpRY6zyApwRZCNRWPd5IEMWejyaJeEc8rsMxoIonhgBdmU0PLOczfkHprt
wufo/gYWVPthQe4Vax4cdDapLYiMnFpVAK+BoLR1VNIDX1wXD+lJxUmzHif43do9G1EF5rb7rDSR
WtoBVF3LMaG4/e8xNgfnNH3YupLegtZNtcl0D3w1qGtEN5sZye2P4HvBWmqVW01yKkONhU5Bz8WP
Q7t41o1Vp+RQ4BZerT84XsOyhfsQw3HkUM57EjTBIuAYLSgKqszw1sYz2z00/mS74cbDagpJrpqF
DNAn0KdRVyYtlO1xICFkLdy/i80+OaXmyLlAF/fSnuyX2k/fTh0cvwaPIdzSgJdwGDR4GNm3FBUW
Z6f5ZGTsPXopPhqVHUroEktHbuKOjGrBt7rmtiYdxQZKYf8mgwHJw4uE91i0RhENfGmtgd2YrLmI
YugSKuQbn9zxssA4Yc8Z8xIaz+ReYLBxai3Yc/APhBHrBJeSgcjCnHZHCVBxcuZ5Womsz+5GfA5f
PYx/VSQAIDA/kM/VOsIR5me9WnId+BZq4sZx5g4zrdf3ArrAozSnR2Dl0KQxpHDx/lBvnRCA0MqN
dsIMm2m4Rr2E7JcNFDbaBL/xSehHIJ7GYxourfLSwLXTxYAa5SxQioCUN+KnFY30PKjKsSyxZaS2
teWS120jSwLmnBqLuZmmmP5aNRv3soqUpDgLbnWBDWFfm4gSD7JNRHqFrCRsQAmrYP60eVRVMwBK
VqOyeEDVuVkvyXri6iJk6u1Y/kuMKx1Nl24C7tUJIVEHj9AKDMkt56BeD7oTkU9RlJGczD5T7A0T
95BjSxNmTzSx09ARkhcbmT834uty+VVCHnD4TGwF+LIcuJuqAZnB1fEFtjRAGu4Ff+4ncZLdDl3R
tQB1wOAd7qI2Mtm26Yhbk7ga+Xkr8a7R3liDoKy4mGL9CFaES4+s261T9FqsbyK4CQHOf1iAWtco
d90h3dSvvKtybc3ojtABu8ZViybyWTgymMnpOr7pFe8Q+yhG4lDFDnAcA/Piv+6AlQFWsYUMs7oO
iAYncrX9VPHfASGF6qnqYeZigqNeesMHYNL4NEY0VJk/koYsFhGjKrs1OTMhGQ9/FIEMm43qNKo2
uXc6I38r6oo4zAGBbiMI+D5o/je4tc8yHekR1qCav6PkwF3Smuyv792aNRIFAeQ3Kt2gfC95ifLM
VWuhQA0N4ApKfDDXaedQMQ4YMDSerTZKXwbpyus6ooLnWvPK1XIAWJJq6zVaHsBB/dvrpyTSGul/
9DrDRiEySzZavjyZitrz8orsE6X2xrLAX6liWN31xZUM5ouctqjoLTD3q0LaipmL3sm6wDxTBmUP
ig847+5sS/pc/xOvrAsk8PmbSGZyX7ScxGYpKV0I3omngfPMpZzYtbWq/9Al0JHhCuF6iUp/lw5p
X8voJD+zWkdOcEjhP6XeTAZQzVdf6CC/twQ0onBZtGeYwHYsN2LuNwhAGlwCTM1rM7mJwJ8ZGtKP
9AJYw/mb+laknVIxlqKcM5Hywr7nMl0/SDmEuwzrZIaEdJlWm5Zfeljwps+uFeHoDcu9asPwrcwE
ft0X8n4VYkIzRoqrQ7+F28D0EqPvJpW9LsDnDX8WCkmaHkj8kufR6/00S53u1mO+QtA7XmeV1Pyt
RloOFOJ95GDpDMT9SmfJG5sjy+iAAAQd/ABMybCDbdgUNa7oLOaS1g93d9RiD5BEvEee+E+qWfTg
+ik6RsGMShPY8SS0ab+pnfuegAKN1WnYfuDC7lACIr8CrwHxF+jGHEKHU/Cdmd562lUeITJVLaD6
EWzh9SXLmSB64/6quOlp2ipsisM1hNgrruioUqv68+BU7tVQryhQetVM7fYcCnV0cDEYkMWMjhlG
skyC7XmoelVjd90Uis2pFdBFErXXz02H+nT1gQnGBOqq9I74Ce9uj5JmLt1Um/vPOc/SzuB4yYkW
waqPcWeTjHbNB+WqrDX1LSa1wGt5iSngYhd+rpBrDG7x+TMzIhNPg/G4aZb+EWcomqIwoHILjMBn
LaBnq2W86+Nd2ucgVmSuHyzIZphII0xtW39qacj+6endCaNG5o2h2U7nfxmQ+Rz0cNuAprNC4ei9
2Kfe2dyHKuW09LOokloLvXXGvm6CMXb5w92VTlf5wHinUDOhtAQSJUNsgKcTJJUT0bR3x3uHojn5
dJhLKO/wbI2I9hYyMDTPmcCIFMnixWG8pquYH4hz8TcXFPhX85jmNps25SEfr/XSFzSRMYHwSIal
SCGB17COOAFUnH7QNgAOWFRVJsXPvM4gkfZpasqaJnlM/o1oWpXCB+0H43Bp7RH/Qx8RbQXwx3gW
omm8aPlpTRz0xCpiZ+PeWfEDv7r8Wm1WK7hke4Zpz7WPE0bCtVugymHEg5y1jb5R5uo7bwdn/0+t
ZHtIU0oFwri1zrXkxXgZVZBVyfAqLmYk6BMvSTYOQfet3mxbshTDZp1MDkg3aaRM3zkjrjOvBbvW
bwZaXf8x0VTup5s8hf+pDtPloI5A1iLgb7Won6jDomzTSs9I0/9O07lLLvSjvCqLiZdLWG3hv0u6
KaqgJkKKxxFKpEBIX6BFMAVDmbqvpsqdv3bVNsUM/9paQatXe6audBAKZ65vGpvtol4+/Wx8j8jd
XjwXLmg4hiVizOCGXzbR+bsYpcbfNQviDiceW5xBRuH+3msEXmpfq56xHYL65mRtfIIQhygsSh/9
BKYRxJWc3MKBfUNGDW2z/lV5R0mn2bWFF+u8UUkC9HU2yNSPIEZWcE7Ka9O6dxA8zwhC/85h4iw8
CNxqiKplRONRI/W7CNuMLGDtW27R+o0mADpbTLgHRO5OjlsyC8+HgbT11Mzp21Yby/pWjq30C0Q4
tkWLeor1GuC3Y3Zuqmrlmim6N1xrKQ0VwxP0P00QaG+HUoXZjBPDQJFXmwaCJWVDKyKkVyOUaD1h
ezKnxW02/pXLH/WKka7GnuzOWr8FwxpRrWmm1Layhy/VZV533Q+b7wqOhtpZsv5izLEeIAT3Z1D1
sWnmvzTXDNIFnFr9Ga6R5fwLmufD8C5WPXw3JlLuCz/A9lZDW5v5T22n2cQgF01hxrvyPdxIjKhS
/jk7A8XZApE47VmwPsJ4vEPgawBoiYbGIIY6TEeieuKsZe78DVHuJhRdiK6eNt1OyQhIuMRhwxqY
X8tRtFWPYqUMOwAiBB4eHqKZyYI7a11GLdt+VDncvPjaHKhWwegCaCwCniYMXdouLraGJ4L8C5bW
lOWrEvrhxLc2iBX2no39NxJuDPBPEht0wyVu0HHYLTy1be1HDyPVg2PZyBAH3KaWz+7H5O+EjCRP
fp9VMPbkZraS6npuEqkET4tu+ZMOgZcvleo558PrePJj+9X2vg8YeZER2c6k+ghLDugsIg0nHtcO
E7+8nCYlHboedq/BBhwGC3aEiukcpqMzDP+X3hUyl5ckFCoOqoK29MzWSVzs0HbQB2JuYVAt0wdz
a0U7agVQ8HyTZuils1QGe183XYJqVYwL0zU2a0ggjiahdTz+3JC6JSm3ZA5GO8ATgN/1ViXrGPaD
E849mJJMTJMOJrQQTyL497RYTT0BFiSlZEyQyVaFBqHXjceiJhM6Ok34Ja59yAtMSB7MQ90Tk1+G
g/xL4P8BNv4M3AxmWr7ZhEOe/aLh2Kzt8e00D4g7BLnm0jPowNt6gaAFmn3vEPeqiaRu2LwuHJrH
fGWf8XXxl/EeVNFIrEOKlc/bMph+F/LEISo927pSoATdtTw0yeOC/Qbi7vCGsQ6lR92lRJf8RFgN
bkqV8z5lYWKN/l13apt4EdKYlkb5zJuKOzSQGe1Q+aziZKmaGrj62J+H8I72xyg9pKsUb0K4vbk2
eateQrkS/s+idDOzAPMzUeoD7y01KOHoKPww6/q42ADf5Iggr5itM6Z0OJUpPqsn/+vr5ly4zq+f
1+9ga3mKEB1gvbpu3uN4fxTshDE1vVvfjW4aaOQzzUEFXpnGjsxMh5wO+dori0XzCGvArJlhZ5tv
INuDbNnOy41dMaGeAD4t/vlohj8TcqoprCLo0b/J1VoSPtj72/Bpd2aN63VSGyXF5hLDqea73IkY
986QtWo8TYrhKgXPSIyNA4fkBY1LvXiMYFh+5hUEIxucDehfPss+JYuV84r9CZi+kNc+BZIHjDDt
Q7+UWw1Ru6bzHxH9ZyYFb96MhLYOqA1/8Yem5/CrN0VoznqBqyM2Pc/s1cg3lU027U86d4+uCKdp
+MbTbhRC/r0bMR/q6BOb2YxACW30sxql49irGQ+d8BoTux4tE2jgr/VPmonHH4XCr5IhJF+Wq8Yt
3LTHhK/qhK/D0/JxENw0kpVCULLXSMGzAgNtMq2222Igqll0hq0t6nJ064ktcaVZyhsaiGRI96ww
1uD6UbzpQB+uWk/hTYVuCp9h5sRzRi5deLot5/xyKKNQYeoZT2rZ9qTO4+/0ObjSQOnAZilKBpP6
R/PnKo835diYKPbDfJrXuqbstSJ2R5+PQImP9Eer1/TUWWXFCp43u+xR5VOb8gnEqtiLP2f+gRNg
p4lkNloLir4n/Qw0Nf1UxEpY2wgENfD8LCYf1AEhIgTRKgAT8GSzAKmFjvN8C0wVeI048Wy2gtlv
+MK65cGzBaVjRb1Qgoux5ikWh2B5prGguLO7tW0c2cbRDqND0TzKVxz1C6KzQ+5/tWuLHLwMkHxh
I/CMTeCIjRmBQEEteer0oCrFI10C0XhE7QKhutg1E/XGecKxxLiB0bZpsoF0ifhyWf93Jhx6Ny3Q
2Go4DOfYzAjbINAY+84Skf7P3Xsm1KrYxCwWImiZjbbUd89Fpk7pBE4QCMP3n+MGKXtAzWpra+PS
Df7bOEJvFIO8sLJ0hxw9YbTNUSDCcTvNsr7cDCZRQv7pE5xm0hLXVSJPx5k2iRS2/SL34eyHQkBo
h0SYc3CBx7cUjkKCKaRo81ZN9VOBmy2TErYtAlm3VTlcIuA0qz7xb/gl3y+WKDP2ljyOeNyiDHmP
Ow4gyDwx4cUXEIikWDP2Mptc9KvAURIXizZEMEkV8ZcH9IeODxCpYV6+/mebmrHLP1BwyHpWwhHn
MHmk3/zXUHMF/Cp5olICtNyEBJQZGMbcXnW2+wQu97weubrY+0nzbxT9Oa3bM4W8QLV0jowPrUQ5
GCP4m/ynyo+2tkx1HsjvkZt+yXxqGBVM9YmHurAlaaNJhRrL2hpUmUjsQPdkxZVLfssadKsYXwjA
DozhjtkJy0878MPUe/okUJnLlR1xkFw0idNoDOEnLOXR0azmi2Q+K40sjEeWG5z87mpB25x/xKUU
2YodabvXgCuVOFLLa+ycJ0nkdLdsB6XTCe4PJxUH0nOR/IROtj0FSa25TS/ilnhdE1FJ96Xd1RSj
v4CYxEYYOoO7CJfIm4SFeKS+I7P0mHZFvD0/VyA3fCgrPQy/EK2oDPQv4zb+Y8Bc3Pb0MgD2+Sex
CS3suE0Vo+32UnHtIM8aQrPJy2NgcyItduS4sMjc7wHSwihwbWBeQHkQfogfuPNhDZARrUZdm+jo
xC0eIGhexoaWtcRWoDSZwN0uOgmO9aop7eGbquQPqc/HQI37BebLmKpWhJworDU/2rdapL6uCDeG
jBqX+e6z60Qkb9H47EndBi6hm5YoaVTn3IZn/1mGrabWzKLgrKLYy2IkdXPMUyUDrv0NOYwQ+1Ik
fFe3tyPYAi+g8JUft+Gfc9J5LXxKERW0EDuY9oPdb3BwBZTHpXTUy7j4hxhczq21viWkKCqwMvN/
T8UrFIDzgV4O7Ta7PBh7bG/851aKeWCcv1zUEFLDugDii15qNXgVTRzqzKINLnAoi6l4MiFaPmhB
55Dxm0YJspEYrv6eiOMH+ajzDhKzMuDM9qDIhmfXq6zOejyhQ+UMj1WvtxBL29dXlSGtNJTDw8r0
G8prkpJ6jwIGhL7CJtZzU2h6VbZJlpdeecmtuCzI35FsJ/+Rg8CITSmGwm7L1R+8yws8Rz5hCxsj
d87wVvi1KUirBGzzdyFmlj9L9LOHPHuMGfPi+ZToRq7urJFqfefXyav7wVqBlj1BLFxs7xXTbF2m
J2tGGpqN23v+HzZkROBEEiHJ6gH7DcFyCgJpx03lfT+OpsUAbWPpXt+HoGqSYmBob0CIqs8YC9WM
am749vc5szccmn6gYFVHFsjCHxa9wuBSvzRo6mELnKiVFZaz5bpCDaSyGayOT3GnwMxhNVYXpjZN
aaa3CIDX0mCtZzLX6kTBL7eMk67TRmLRrtN8InG8LLu+gfURwQb63RHl3JjR+E2SnyvT/epdYZTm
j2BM2fjfKmYfP6+45YfH1PdXMw/cN+QBr7foOwlXwHcBcAInsPvn9UJGLF0GfeSZrobsB1wooPGo
cqS6fjcUwzX6JESlnD/gvSrmJiWDi8oJzWCpKGlvoGSNsWHs6LqieX4h0Rma9IqKaA0EoeI+c6Sy
bhtnR526OEziwW63GyLl7rGIH4hTdQ8Ashv7JgTVh8MXyyLXH8LAQj39tVi3iMasIjgDL5ZwhRmb
p4aSYI/lQeJkSg0iE7vbK/FLI9GWh7eiUZnTX0Cz+hAw5ko7hjjU8OPZ3pD6Pyq0kdmir6/f7KH8
dTVOxZk1ms4+V0+cYv3J9Px40L6CdgG7bAdZkyBd4kOoB/PSTgdfQcdWh8uVWG43kIImJJk08FDA
Bwd83SUAuNt6cDW7Uz1zwqT5iAwpOHD0a+F0hvcQn/bS8qi7vXqFoAQxigCB5LK6X+Nc39jPRNiY
DneJfFoAI3JmLjgqGmHMrQ2tiImLpdi3JH8IW0MScpfzy0k9Lx2KGZNKCZQoI+iIgH5JAj+qu7sl
d+17kzfXyDZ5931eguDnf0q+0/7GWLA9R2Rk3bbb2YXGiZ1Dx7nb9r9eF203jyNPgpA8jQNNdcU5
1M0JI3B0/ti0j1KN56b/mYWBSfh7teIZyjfjD5P088lu985M/ATlqU8EVcp7v1WPdVc4h2umeaVt
wjDJofNI62L7vj5yhjU3wU+7umD1q56HR1RCYsoenRoVMNB4nilh+BEKviGoZiR5S0PttcPysvTn
YWncunXnPOWTg8i2HJij/Hq1uy6ybXW5rIvmHDt+XTpDKV3GRVRe1yoggGH2QOy1svnbpcx5YeB9
Q6cqpnRQSrDwWk7PQFn+76z5kWGSrWgUgDDpvA30Q23Fec/0hzUwR8SQ5pqDLiUzqMQotu37qMIc
B0yEwg7BiASU/K7APGOyXWFu81CpN3aCuF2N7z2HLSWqywvpjVRiGDhnVRqdkvA939v0VE+MVMDE
ueKZoLJAJ/+bYik7XncfGDxiaaN5/kAC0kN8wXo1yzNQqyTXCSW7VoRPxxJsGFM71k0OCfA2sogV
OIND85toAsl8tDZWoJzYsyapxk4F9Q+TCeULahCrXqCxNKG3UatAD4Rg30aC9z54IQjBA1cino/t
hrowiBjQKU9WEGylApLlBFCoygtsQeEHRk1SLqDCOc26k00GG0gjCLxhmuD3AJWeOa/BQg4Tl9jO
KApKswY4wYKmPseuk8QpepfDWpXo01UQdOwBh+e6jNTLg/9wRSIff9zies4EpTGP/rLhAWRquyt7
sAo1F7acbXL2qbm4PXVyZdDjEFdTssXBZG7bvyZi135wARBycD4gm1JMEEz/D3028ak5iefPaDRE
CWCkg3G9qj9J9n+AuwhUwDSCmD0RW/Y+fKdANWRh37InxbOVor/ChYbtdoQKR2EWa7QglbIWooEd
CezBAXDo1xzkDJN7B5D/GNgd9pKDA6xYpEKEiV/hMXDlacc0LYJanknYF8nO7KlEI4+0fZWnCEw8
URvyf3R4vFQ/YV9dTwf9ncGPQLCBt726N1uBckasZDTDJteJXfgNqHZjxDh0/sfZC2WHo/uXyEUL
OFASruBh4sInpBp5af4h05EHSRVxGm19jsyrO2tUtlYVy9knj7Z8ETf5V9BbU0f/8TuwwPKYqfr7
NU4v06skoeStlswh9HacemgKev+0KX6pJSGFB9JsfQLnuGV4c+u04C8sMwFP+ZJb4Dc56u9i85MN
1sKtHTw1sjLuGlD1l+stcXfh/ktEqzL6eW9BC+OvueFZsqXIK0yevin64lhpf1bIkWgmk943bqiF
V9IJ/nbF3geZGkJJdMTFc2tXcYlTsutP2DnUAvXopaxOJgkRRMYrDi2UFggIhdoVfjWtxTT8TIce
/40NNhgtyRCIED/7escmEhNizEUCaBBgb1wSVbqrJExNeVBMbnDgpoSlAWft4yRQG/Chg4vD9xub
1otjRfBkgO51IPUmDDHcSvKrdsnQEb+349xQQ+H5n5O91jo8jLBZQiUF21vdMQgOOy1FsU3uylpz
q93lLRlFPTnoxZsqLUn9IWvdGfkuaFNJKCekdJ8GbEOIfWfYlOtm+jpoSy/yEtZWqJvWH2TqEgQa
xyLt35LxTlnT5E0EnXugZ3a++/2ccnocUVoJlNe+Lino2y9G4Rc/xR8/S3gos7a+8IN85yIn1+4V
MxSZG4BN89A+Lgc0PAClWYES65DxbOP3PQscUEO4bJST3q2V2ojXN3MNY2XmzM5MHUtueilA8L8z
bG1S8mdIYsUyUZU41JGTeBRdZYtSUfoMdQ9fFRSHQY07uDNf4Z+9OtI58tR78fOr2/uRUtqeA6wI
CWurJED8T2kNljwQNJ0An7HqjMGPCNUy3NDZmh7QJzkAd1uIXLrF3yAvUKoxMAWa20xHIjDFMJwb
krm04Htc9ctZ5f7DogVydbO2RZzHnw4I7N6BTzuOsHK0XIWx/lFe6Wxx+sdmQ25RsYnmltrA4Je6
EwC909h3ElNhYbiQZuo40XO+IXDyGUnjHXqt8bCwE6JN9TGo3k/F3WUlAChyL9r/QgEybIiUpCu5
fjhKjETO8e0o5MwUMFe92MrOMGuRd4rEb9BOx6p4B4rEMPDvPzf5A/y6B+9vXpo24F+Jn7vRInzv
Em6IZI4c4Jq+SmV/fWHGMOU3FSr0wyOnHmBKEbPN4Nt15eQoJ+3T9b4EZb4i09F9HXlUMcqjisH5
Lkj5zWUOGq9WP3D6cbiurdLkDubjYbr1sraB6OckD2mvP3Kywo3LAK/1Vh0CJjSPg+eVlPW7UKk7
9sh2584uyR7WjoNMlnu8AcICjMr98LIA1Znn4lzYI+j75e94FOcpIKvoLMyWRSANYTyN47BHqLlw
yRI7ZKeOyOuxi67FnHB/UVqS3L8uGGRfeusPyfe1GVjRbhzucToCEsSpVzzwUvF/w9FOtv1R5LsV
+VC4lfk78xIoWmB+Y8S0LB9Gf2aso4WlRVd67i3OEvHs9beITD9qTcuF7uKNY2IyA76mxDUG+9EB
IAYrsixHWXsfnZCgxYbO0Q1HOaXpDdbDJNO7K5gD00uCIexBj9KyFRQ2f0P6Bvw94VR+zAT70zzw
ODn90bYPWdXLL39eKR3oBcp6zsAhnEP200R9IMtveFj1vSwIyBSSxzt3H5kRZ5EX2+PNyI0PhgC/
2rD3+087TMUv9T+O9BaHjmmPmr+DjVBEnzXkzVFF7iAx9r6FOtFiiJbjYzPFqnP2fVa4HBOHVBO0
o3JqQ8vqa4znjVGyq3sWblVR46I6eIN0RGEpos4/JKeEh+ZJtZGajiu0D034dL7Z9p4c2D8KAT6M
LuFOilNbjTjIcdWh7lmilzUmLZo+q1yL7Xy/aH29egelafcY1ISIgIEbFvjAe80OJBNcjOPvoX+8
DwT32NIKsfGglqQmJ0XvgOh8mk3v4Ew76cSQ/ImZSEEFZrv+IzpcTlIhoqifVvKzaJpH99VlYK9B
irR52TZnxVE3uOh8ifXroU8tOEwYonG6iOK4SjflWaIr2rrEV37JVqyLLTfslfS3SZVH3OXYe4Cp
jmvJBDS0XphTXP9lG/uJK9HJeiDiczyKjT6hJ99pm5D+M+Cp051ezh/7Z6mRKGISylp6ZwWGyWT6
GDM8qeJU88NtGuAxAWTLo62OgxKk5OOghP5BvnjZU9idtLmkxQMUvEhi3vQRsnBS+rTO+n6Srd03
M8A/w9G91Ah0qhoK8+YSqmpyYKLMOL3LzAKalMtn0c6n51qKkGbV4DIcAjXEwMwR/P3IF+MrSNO3
0VizDzCP77F8wK/RIEAU0JcwDHZ+WaenV3fSP7wYtLsaBKG4E9MrN84LQ33+/DaJLGxTQBYwbaxN
+FOwC74jhDLbh1YPHj9e5v23LdsV4O0FUMbQtCc3kdYRelk+fsUHK+30LrDHPAZKXnfagEIPJRnZ
pAOVvDVwgaECVrTXj3vmW6Vat4iTwDL7sNjk9FlcZNd6yHMiMgUmVtC9LEz4nmo1VlaB0s2LGsO7
t0r3GhUY2z5qGSs7lDUOkgMf97+Sbd4Tym3WaMH76VPYxfTB7y8k6/y9ubW+PnvUEZDU7zWrME8b
GPP6f8WvElwTEgfl25XA8e2D0mI6F1vPZn+Cagmrew7adruqlYZ3y1SnOjYKynPcvtEGR0XqHWMb
tB9yIu9mInSanyxI4nyHiBPZGy39tZssELEWQ7/D3V9gn65qVz+BUBG9kwbcdvLyfrT78+FA0vRj
zQjW+sKA+pSqjBX/aLk0+rncPggUpWGMWcRBGkR44FTITxToNbX4gu68/xVuoIkIMK5j+NKYa+8M
j844tPWKVjolAfa4gH8NgreqeAUNS8x6Fqx/6+kp+GghiTgKqOM7zvj9zyg9Ud+3LEdXkSoEZzlm
FCdrm5IWmtva7ZVTeCeu9+qTDoOxwDGp96jwRLJx0UY8bjyazo3Imvhk6npNLsUfFjoRgHIRmndG
sEdn+/F32PzG6m2Vpli3KoZDnbfaKIyNDM9aoESjzdGs345XEn09s0+2Wnx8eQm2hfK4PiYnpBDH
gYEgboBHP/H6h8K37jdgloACxK5bInp9nHCcoVopWJjphIi9y/RbmQopFQOGofqRtdRyWANpF9sR
WfRwkiXrtbqlTYHnFBFVe3rC8GHBEzGQOya+Uo8I5qghlTNH4qxCg2kPCjus6aDFfaNeb0GB6n7z
jROv3I+HbgEGq0vbB6PnVgnOxbHXuLYx8sEJ6RpjD9l450aaOZfEQq8keGYAtd3gaxLl80+XsrEn
qIbbhSsHWMI4l38MlTFOTlXhsIRGRfsabnhMXYSebq4YPvABcTdi8VmAoss4/MZ/seAxgJMtoP4p
uACmqx7Hv/5WojGGl5yAo40v4tbBQ8LSIxvUwmx5e+7KSN3AK896iBawlvq/wjp5YT8E9+RRuoq+
zaz5fDczrqAZPQtkxAI0ewuQdEhHKc+SPDVY8tfCS7SeC0cHrIxgYyeWyplNadJRU7ZC1BNgEOhd
e2V6oj33jKFzrx7Up8flxT9ec0latjvpQD4xc9Zvsllk0bFjtcmFLL2P85Qh0kZvt4c3WAANrQBW
uulKABsPyBYpgoOPsGkhVl0q098jDNRiQQvvhkDxRXOkaLt1vXBbko3+YrhzGAX7efDKTTCUM3pe
Cx8GTwu1KmRdZAwc8ePyob/7lxRp0NKHNDQM8lqEfUIR6Uvx8+vUVUHNBIQQ/MC1cFFEEL/L6Kae
acMpDv/rBr+K+iV+/l+EoHzOC3UPQThY+0YVUah4qW4ZE7zJy1M/Cux1DOYeXBy5GqyyzH2NUsa3
ltLvC2H+VBArWW7WuXySFh+yXLXvQ5g/0j8FR4KQ92SJvmp2CVUYpgcSgy7hrhCwrE5EwQWauWHG
hQb8liaCoDsj50LRBQnT5R2J8y4gE8ORCBwHiby0iwPD9nSRqxHe9Kn4hWKM12KbU+nlYj23FMI/
ft+a6rum8G8729ZvuOHcCol44NuCQsCbvDjw846+yvYTvxQIROCRNP/PQS1S4VHzSRM6MOzVxL7p
VTLI9e7j1h1sa2GlT8xS/wJfiXvcNiksnRBv8BOhU56NYYtxbzGG63AhN5zDMGIgp0qcYMZPsP4M
VOztbd0dZ18U6613zTGlJ9hF2YZwz1THfbGFu6jC0xkXDAxVKn1Iw5wGKIB4fRt3CkfjJEc0LMJ9
bDB8DoOBabExvW6jGnqCi3tKMVdbTARxihRiTjF8WxojVAtt30/F3TdQiBOJhR1Jho1G5Gi4Rcas
Gsoem9prOAWt94vqb1soi9ZxnUnaWyNKcdMWPnCsdZZ+SGcOF51t4mWOtEjg3xuoJvMgARmKWRon
3Ib0t3E5BjF5iDCGmkWWGvVxm6PysJneo57H/qLgYRjTA9W9EoA0AiXNQK3gh0QQjrkZfMKlwW4Z
CSTaUlavd0m7iY3UlPoRUScMWPhB91AbuA8/TWuLNvS8LFh1XyJQAM2wF+hrRegJwLaMC5MVlN82
2cjFMv3iS4da8u3S1jfaDluEfZhLSZQ8NT/ApLCUIAlJNaM3wGWT34oaGFlw5Gf5crzfrp2Lgrxn
yFXf9A87uy7yEkHd9gDWbyicLyT2hre/VM0fwjtmVD9PRvY5VcE/HLzC1xLKs6qjB/iCRR29KnKE
lz1o5UBbgxksyNvHyyXoG44oh7yKZLRTkEF8QXZLAl96/3Tq/IqnDtAJVrxQcXpzzQy6+PnzDkbE
Mqe8bEjTomc+GK40rhU+17+c8J0HBj6KVNxRD77+gcmnD3DSp/J7gAKQA2a7PECXQXMEDnXtCmmX
iIGNdlLddFw5aA8beF03kfShw56cuwvT9DTAyseN2rVH0ESOM/Jf+AipwO/vA4tr8l2Ox/Xs7vNI
RmGt1/QIXV8ukiSCcE4tZULPnPMMQY3fT6KOkkezm5CTQyPVO4VaZp7OFnpP2H/iYfkt82+NPYbv
F15RMsn8K055ualoVDUfhlUhXU436et1xtX1H7BRfLIWSa7l0sMGr8xyBZCMqKbHbfFOi4Rd6VMV
3QGmB943zzH0WatZvIXcg5VRsqKWugZ3FDbFyIoTSbf/kIfZy+0U58TKUH2CzMfgCEaHmlxYV/ZB
JkqXm/KqgeU+KrRxKvhsNSwXclS3m/gBnU8JkusjmmCOOA2tylMbaxh+xOkf6roxAWrbz7o/nt7e
yoh8CKHVyJs39kV/kJycSKviW9H3FzSU+zBklvcgZHjWkgTJI/ximVYwqShFcVWYCwXxwtMaNZjs
8OOOY8/2Bw6AOURHm1xNK0sxbp+f4bvD8kgmK714xL+Cuzdeq6NKIs5KgBQthIrH/yto1Ow68WKC
isGXIlPF3jrnsB+IMjGs5KzdmjXXUywgvGLeKf0Xmyc5nASKOegwk7S599GfU05IlOgMJNFr/cTB
joPS0BDdSwjELaHbTq/ZalY5Jg8Fcl7dT0tozzB7qKE6YbHlctsXCr1AjIwjCvI5ivvaCzIQ0ILF
htqRwf8JKyXsvXajSPftR3eDeuj6AdBcqtvklZj+TgGx3T0/m9NG+e0XnxY/ezreZw0xxvJx0lk5
DstBgvh6GAF6f+qiz2Zn4M+Q/gVbHjYTqU0q1Y6D0Lqd4kupCqYzP77rkUNLLpZx7Kh37S83PBZx
mcDlqq1V8Wh8bfHW0m7D8gXUOsi+MZNXKhRar0DqGpkiFnCbBEdusVK17EjXYO2ptU5eVql8wjh3
xyIcwdZvB8wAWlAwfF62A0TZ7fPoHiACTkj9bgBRr2AKn8chnF04cJ3sS7AMF8J8uhuQmyTcByDX
VXgcPSJRbKaAKlPTPDFFQrgmLqMDcDpEL+EgSD655EqNqIa40fJsX67I9B7PvhlsVIHRLMzx5cZ+
iSZPU2meVK3OSgSYq0g/9K5rBNr2za7eb3RSUGHIGr+k9poxh9UJuEeBDTpf1t5CDC+Tg/l8dchW
XlAI88/WETEpwUkpn8uVee8rwabYW3UZ8oAHybyEExuDSAim+uKI445oVobCmNh2A8fyVQh8WvCG
730Ykdb38YNw0Vo3ALwZnoXXZCWAKNSOkcZB9Wn22lbwoyVdYqS17FviMCOWLSA2FL8+BPX0U27E
9kXaeKfYX3thwf2Kt3a8CFziwcDrCoHz5wO5F3SeThwEs90dG2EBXK89/FmDrecCsVIrebecDVra
zHH38yCzCAqCw70Wk6HuCYdZlrI8b1WQLI76l0nYfad+8Ubo96gsX6TD8uYXlq7/efox7xRxwIWP
ZDAAoQrOBXSDjAWfptI+cisPT558cqeergsVJlaYDXt9cK6ELecHmuNQn7XWypb8Oj0ZDkNH0OeN
DJAG4bI8HkSGzguG35vqkQgHRcSMBvwoG23W+Q9beKtawiu1PB4Kw6bSMZqF9RPVPw2+JWx0BJle
Yx3YwWk5W4MTaC/KdI9sL/kuvI4hs6JPlDHQg+WKMdy4WnXx4ZmRNPXpk6KoFBLbGm21vuvW1T9z
lC8oOI9fCcqnFxSR3Z5MtZNTkbH1Eb1Jbbo6CmJXvaBk68yHrULsiGPqN+6NCxOZE+84lyni/I+i
5XBU3pDgz/lFldmwTrGOTwsBAJeYBpPte0fDNuKc0C81fVHiOlw/VwMqDVsGMCSkVdm/aB8jC6tf
p3qmCeD8QE9fvjkbHSdDV3uBYSVHrOrzkXjVv+C8BtRnIFBPvTY9rcYawV8ZnIxcH+FHtsQm9mwF
L3Eifp9COs6VPCFPk63bBJYlLAb7WRIP2U314uugjt7TKJm7Vp9R4IsI0jew2ZwfuaaHXIwF/KXm
3YmaWL3ArRxCgfJuN9PuwHby57HPG8AjHwn/m9vNzUCP+E4Rm6iuRsQP0q5u6hBNFEA7F7mSk0yt
14z5f+A0ApaHMXuA72vGakkEYe4QrPcKyvPhZbQz7pXi1WZGmyy45DIQUlORCU7hwCe/CAW5LauS
LBzEHFkd2OLUOJnphVr62YQgJtshX+0ItkmY+/05EAZDu0CcUgxS6kufTfyua9j59EFPeT5wiBr8
D316e3LLN9THFWWmqajCyc6v7UWhFJyYo+9h+b4FUoPmCdjz8Alto0rURHcJg00yIhBacZNq5npj
+dGs/5Y/K8Vh4fzSaVps6DjlIp7v8fVI+Wi0ojm/aTJwhKDkp9ulQzoP2Das/ictZXbTHPidveEB
SSAmegvg0en3zygYthEbia4hh6VT9L2Ud88/DG8mHuL4fi76fAdRSQTB+rxT2Ez6WkaJd7sBENrn
s/yr9xYexBdhm6BTgfHGwD2v4ARzVGqGYSYSMB7pqjkbS2+O2f9xD4+XN62bY4HKqw11vXCfjZqX
p1txWJY4a28bpID44M17QiVDvezQFKc/xshm2faQbhxYT/JQM/qYSipxTs4seCaU+pgw190U2XMK
L9VXzIkDm0ACrcyyUkgl2oIPWwjiT/4iFtnDluxmrF08Wb9QNwF5uvOjUe1pqWu3Ce87LdMmVOQU
lKMvrVGsXX+PQ98O2m95McvWRh9xFoTTY0XpaYOIDBSz9BxhHvZREAdE7xYuyiI6wywLOuQwNnCP
AgEy46XH5TXAA5OvbqopOlUMCGlsuIM+sajUWpbC44UkRdLUusts3h2TJnAa0rwPpwYFHdseT556
RNXm48VKxL+ZBG67ciglWLFmL4u10rpXH5bALVPsOGtQ0VCQNFAVVyDSWvayNokZFDYasentS98h
9qCGM0Vcg4PCERuTRtGAZKF4twJZPyrRURFAid3p7I8BHudVS1vE51e5fkb8k+zdnGlJvQP66B+G
GtCWbxBioocarR9iu0zCqKEj3vuS7rz494dodQRZd08obWXIvlwM8B3kAWlclzfj1l14K3b3j9Ac
ZvSSNwHY/Hqe8JMlkZ6KaPhqyizGPrQquqj8kw3CC4ODxLm40Mpr61A3DnZjMDknuoVQhiFKymd6
1LklO64OB7CTpFDHUsj04I8Nc6eIEIbioT2jyqheOyRUK+4xPoGuvh8SjyvzLnGgjt7T10pcBDEv
udJJaG/iVBwrequI/2DS218oJqNz8BlcKlZXQkrplZBgtR5ADhzaflg0KHShzZ9O5MK8U1h3gfm4
4F/q/YKX/lR4CSWeqZsYrwfezQUjgOgfQT+epL/EqzFD8wfG49KpXorLFCjje23TD8+hIKiZ3dZS
MLFqlcnNM8dlZ4n2AQNkUZTKSiOYUBvfIBPPimZfKtq5rFfySeuOH2kV4ViIGw4aVHcFTng996YL
nM9vRjbA3vHocgz9FiW547uAC+VGTYlYtmKUi1Xrz3uhv5phA8tFt3diXrqGkBO9HNY3BiMAU0LM
sbBQph/kpuuMUAT5Md7m9NP+ZazSHkOr0OlhdiZHqO5LDy1xUhHkfeikwQG+NCY/vEUq9wS1qvZB
3cb8W36Qu7xCQBxLxEAeMUfFTe9ulZgtymEo916q0RhFPEPNfMDsg8Z+eoi89AScUrDHJ+EhGIHm
TpNxt8X5fdqMAMqunwKLJTgqVgvTUMOisOS2fhvPO5pnmXHvkhKJlRC5DYttwHisgxb6FEWfR4yB
CrSMupP2pNa9ozBZe4RwilWnjVqDC8iIx6/by85NxIm141oESV6mhI2vM3f6jGubeGmnn1tdTkPJ
BUWIIOBOQf6Md41ROnytRCMhg4sH2e7EYIyqN2rvhAmEVPebyOtiFBUOLKMagnSd57bS6UWyqeIK
Kd7NnKVJKdafAsinCrY4KQsQOY+peHK7vFGR8nTXi+1Sq86yaydAS5ftZjlJTGGkZmhRNXQgdD6+
E3IcFBzA0vSYBqHsHJFMNugmOFsIXLOgqr6s6qDtVRc4VHU/Y0llJbghAXRNLzi0kCI7guSbZq5A
sfteUiGQIMODtZHEOoV/rjzKilAOWdDZ7/eQsCTddd8YPIKQbp7A0ToV2PsgWLPdnAKvtNoUX+FV
R/Em7Gavi4nBr39Bw4kSsDhAWWRrNbxwa79wAo0s5RavqCJYuDVEsOBbyFq1N4ddNNA7kIUWbGkW
CZRMITB9yn4w1WRJmtT+AF8SohLVgzOjrAn2EMFcXcXzhfFIXAkEOM7u08h/xeUZx41OxQsZYVUS
md2lwkjRV9w3Q728ZHzmVZrDLQE3pO92GBR1q0qvXBwxcURKzAwvOeJDiTDz5wcyUZMDjpwrzm3h
6CnvMv+7LTR+5N8EXyxAwtPsod2NNLddBwP1tLW2StjSApGce99iPQX4LFcF28O5hQQSC+N+Zlnk
Z64Db7wRigwJVqPZt2UFeozvR7E86rAlY5l+wMCGhp3c6K78/8koXjQyzkHvgRIa7RpCtb10PTbm
JZgrYniRG4+kY3xDFkz//3JijrIzV2mFCvap3QO0q39YH3nao2ftU68BsNtkXcgOfOZrxsQg29bo
jFsC7JcT5ay2ASqP5pczSJ0OdIcw7Gi9ETY/0mdqLmkZ8mxy/9nXeSZ08+BmKrTd86gpPlOX2Yza
41zpdKzy1ZpUY1BGScGzVh4YcSM/B55XoGhT8fS6Zl1fW2RpHnzjIzNmgvDxcYrJ1b8gunLNLgo+
xUhRc6MhfjqygnIgSri+Babb0Tc9VkyOCHbw6NJPOPHKczFCnotBB5EHbfiKzJnFETiFzmEBu5Qc
oEFReMCpMLDVCv8E+MJ5B2XDcTtG+5BPqpLvsYm85ijCqS5dXjE/Lzs9pjIQ2Lj3doRjY+zEJuL2
EJ1Zk0E03W290e+6LjPjmF2BuHjQ61HfVSRVFbIuEwuvpoMzKridRX2gkFIiBndh2ou0l9mK9aWP
NFEubobjHQkJqKXBe1Js8PIwiq6hQ2ceKakIxwciRtzgZfz/Dd3FQl416/0SS9sA0xkHdwljaFuA
RxMC2s69LW9QShiOtRjDjq4udcSl2l134Ojk0LloStYDTg/FzzGPx+OCKiOBK/NN6vZMxnJiYh6d
j8kIJJqTJWwUcmOK1EkzCmz4xz8zIaRXV+9+S9N8OCw+PUolzx/Zo+Qjzi7X/Z0Dm15NjzTfkmu0
+eBijECz7bIDkc0XhgU7Fqetp1jk0iNNNU7t+Zs2kAk2hD/dQE/1yIOukpp9e9E4Lg0/k+GmMNZb
gU+mYnDxRmnDhL/4Yq90DzLxn1918vIM41GL2/KGxekJK1ms+ow8QsWWKlJbCNvAPqf7+hHa8FJl
4lPbUfyLnW7lkKR0rLQ83aUMfWY+Oxh+rjjdeQKZ5KJF20/dhqgvHY0Sn0no0fulES2t696Q4qWT
m1xN6TpL/MxYqMkxfL0dJQHG6TFtTxr2zMx4NI1ASU75Lr3xd7XQoAEqUC/oHSe4gt2fVRSgkBv/
gqhE8dWjMWBaCFHxkFXOXHl3qgKf7snlirf/wHowd/CgpcH0RlW6Sf+GdUOlYdfqowuhT0jlCZ0x
ORIbYLgJQvEQlIIOm0Qc3+EvgJL3x0neJdFWRIyC1En/S6ytufNspvJQymRhtH4m0rDrGwxkxiaU
SKiy2SqXbxDRKHO2cKcHGGUY/WXy3ADY3Bh3BzX3pTITIog47fpmzxayYim/jYlLWborYGpvcm8D
xbQEVevdKlclYAk2C1mUwzSaJFJ134+sUxAKJEX9bADA0QY/PdepIFb17+m4eYNaCJAIUkyQhDyT
7Vi2e2NesCveR7LnPgM06O+L7rBv7EkJehHCkXe4KaDKXw+K8MFKpjknVWqe9oc1Mtz/fgAOL9K4
g2YG1Z10nfzjd385cxU7jb3XgtW87f+YKAirQOe8troj1Isc+oi3WpxG/GM+BvAZxSLwRQ7eyeqp
/j1pk+JABauHamLiN1L1FP8dFSv3JUKZ8OE+ZF3XeCUlNN8of9RqtWRnHbG0GhDLmiAkA5juBdg5
3OdHmTVSp5u2dpQDZNiy0Zpr5dyM+2mKcME4wxKVNzW7tfYDQLzQdlE1THQ7lLT8I1sqy112vkuh
T8r7lmrZ5OFv3iKTFH1abQzhwEocCK8AcT9IKm7jGTNWZc5TdmjZ2GsrR1FbSzvLMgN3W0FEUGVA
6yWiDeqlxNzb4MkpAED05yFnqFkGTSR+6PMP13odZuNVCWzYmc99ZWvhs5l/6Z5I6TI0xOOhwEFv
mQqmGdksKLMMzYeBWZthc/tgIPODMZ+w1MJWDt0qbZhU2S21eNaKUx4nl56bd8tzoNn9s+7QSNEG
OE318V6XmYl77eXPfPgLzn7pzaWhqQCt1npsDZFQFAssQxFjz0hvGDuDI1jWdZOkW0Unv3ngoC72
lR9TDzjIE58U+lEeje/ZdhtUNWVTO+LDzbYC3hDEdTICJ86lb3BtLW5nOVLskcWWWNA05zU+wQja
hc6DbMO1NIYxIahXOpDuv7Bfy+bDlnkLja15TN1wsz/B2OBtDQWOD0AV7xcPm474m5Ey+eRMvBpQ
C8Bu+s5HHGv5B/t+wDedvHpLZjxT53A8sWx51g2xya8a+fJUQ8rUliSyq/+YLUsEx/6NGR1MoQXH
Ob88b7i3iKBTKB7z2V4NRS2rP/oqrKUX38Qp/fUf3qr5rrD6oHg5sKyZ6spajzqe/04zfV9HkFJ4
k6y8E/c4H9B5R/PGTT0c/03NWy72qS9QORxT1EZeFNPqHBCn0FispXik/1biMHiP+LkA7HpSsdT6
WlzpV1twWfsYPCPu13VZaAqUPm4MuAFtNI42hUHxpaTmqjB3MIZaJSzKJXrzPt4ck/Ob+b53xZCk
owKi5uhaH1XHCym6Nqw3ATNVjlR6Gu0tF+0vOTNG8RLDp5MEzihEhnfO6zaqPh5sZ/AupyGgcYYA
XHDlqf8p04/zubT5az3ZyTx0+kXLDnw322XcnNl7mUx3p0qA6NV5jjYhtnqnFeQFlEtuNvinChfH
OydrDzwXxm07ft6cqqUBinPKU3bJIxaDR9H4uxRk/wXssQDTSZCbjDBSuWUv08lmSoQJx06JE9am
As7hVXMnfD0U+Y5WIo2vEVsJO/7cn1r147vzlESePwoB473TIBEFU8hOjG3CU9vqGCbn8nkkT1rw
Q+bgzfByepWdu1uc4GxMNEpJPxcHv3KzZCmnihbLxEHo+qWaPFwnC3VnGn+OTTXWIPm3v2T+E9jA
uLNA1F+Y9m6jrXjO1kUoZozJV1osxzLH58DLvkyecIx2wJiKal/8jvmlfFHhi88DMFdqriTVu5Jk
UmGJ+2CMrZ34JFOk25suJMg4jLedAdw3l0XeJpXzyiy3MzfuHj8BkXov1dYOQdSYW9vKaBFiYN2w
p+gT/922OwEuzpc/NTFs/+U+xcX266UhI9D6wXInx4aWoboCig4Bm0sQNAMjQK3MzPIn5yTQl2Wa
mmrFrBmsgzDyMSHoVW95S05X++MW14JzU4O6cBv8MVC1FKV6xCG32s9zJePZCj/XibLWa5v9LMxv
Lj7LANoJIcLPJrv1Wz6qje1zfPRRZxIwZaMzxcscHL8SCz2QpFn4/6QA6BeS5HZY7g/dcfKUGhT7
HB96+kqfWBEoIZqlrjfjB3xP6XWmaD3rqLPwrl9tFPd5IUi4VKszZpmfVPMzEkP/0H1sYPMEPMN5
NxiF3RBvz+Fl4DKqLcoOQxT7X4UlSAsTtTkhCbFCTWa5UD9IK95jmUO49lNaBqFzYHHhSUMut3dG
o6fx4pz6cdOM+dw8xXupprzwb8rWdIWQkWPGOxODGVdb5P/x/yWyqNW/s6/uB8kmgbsWYvRXXTL4
JaBOdpnb/y5eQTljiipKZ+B7xdq+n7TMmlqUDRJtez4m09DHXB89jr5LcdbgxkBVm3eLY71MJcRU
CIatLWGfBqjCB+oQL37UeTsxzGbDjttrcLKFT3rY1hSMLvuhwA1ycS0NrNQvCDQgFQLwRpTn/bpu
Ujrp+ZowsCWg2NSGQVG2t09eTeifMQoWu6WPWopVig9FAxI+mr+iRecfjFCDPBHi7XmEWSgJZyip
m2NeMbO5Enrq6Nv6dSbMNqaeNqCG8pmQ/DML16jMXetKo7hxJGc0GzVwxPNIEE36CObwtAHVXptc
Xyp5C18vCh3/Le+Xvej20jMwISjxej0G7nHxt9LkftNigSxp3Uj+vRim9xdlYc3zKGzxElpLtaid
WBupBdlBw1LuiyuYE66N4cGBqKLhVwDS+7IFLh3myFocIdhzZJ2iiBB6/n5/WsOzJdGX+tzHfOCd
Rzvag/EYmJONZELrtqXyf8jXozPzHQrHkj8Z2mLy7Ly3DEMxfROXJMxND859yUzw30UD8ADqCaqv
rACmf0RpXNEpDLZePLzo1KnosUKxZolx1/BrFqn034c8L/Gnbinl69odtfh4bntjhd7F+x+J3fqL
JLgXMgHshdg4C0MXjUwE3eQdtaEVHl3n22XY6fUJyJP9K12i1SMksLSP3sKpWRl8CgTDnyxhOAZV
ytvME6m3nXkI5rZnVIobBgtItAeWMT6q757GKnxOzWKlVoetnEYUpTkWYqSo+U0J1JDjlGTsr2sz
BjKndqtftWeYN2IPKzAHqKQ4nvT+O1MnyVjkSbS4amp+lOIpG5nkHhzVfvTmkkDqRVme+AfyW8RO
mK+RpdBXtlW237u3m0rs8Ixu1GQbwV/YeOxfx0jqCgoiJJ+wCARol18dzXaceZKnsRamqlVIwOHf
ZTO6/X1qD+GNK5ojsEMb/PnFUzSYUaXCbqApAe5nR6Fnb1dBSHPfXl6mZps5uf6D4WsY5HHK5Edr
901lEcSQIJJW7muUTTAxK8tZ4GaeFAUMfiXQdtvbji+wlzcRfvU6rZVSGblJwZiSM7mlngAAsU/o
44sgt6dTivN6lfwd2y+Ql8eo8Hxirn5eC3y1k/j7Mx6Q/aKJx0qcjNmexF1AiHjg1Kfce22OLWw0
DnZCaBCbL9NYeWsb48QzEVYxyRXL+yNOYK/x39Afqt8sJvcf3VROpr33P1+JLGlUTffWBIF6Hj0+
qeulqtd+oyhPi0xpqmPiY5Fsdrp9oh9xiHIJCZ0rMydT+pwfJWDRO4xnLbfZZmmFzQr9aRREhNqj
vfU5isTWXsg6c9rAbxS3ALuqLQOk+fbRbjA9UFxJV3KWuy6g1QV7xSEGLa7vj+mNtect1CLkclfV
2p27SQ8l1ByXPkcsvgwjVPmI51UVCzuMToFf5mYv2g9pp8xPIque4fnU2QG4GsEhNFZjBEpvUjKG
sU20c4kviq328xwf91Uqpn9D5kDkQQk2SWVEUku1XFXWyUsPooxxGJnDl0NtQ8BiPhlakYGOqRfw
uBPdO4BPlOf8lNmW4M9y0zUC+S+wa58o7/EIH49LWhKkgFTNAACidicIYd3lgYnvQ6f546vSnfSp
WXLpUC0q7/QO82eLC8aQG/QTmR8ceYpv++n+J2buAiHo0jTuj3luGjo+NBlSairZ2+in/NbZMzyH
ivuMWhGwBbhujqbX93wvVpU3iUJGZgPU8+EUKDP6otFEtdheVhRbOi4atGoygDWFF//SvgygyJqR
nwTwmJGodFReWA2x3iiNewzcxklIY0mFjPxybp5BnNHN62VI2kSJlCAjP1dHh7v9s03bXArggK0o
4W5hg6p8D0k7u1YSeum3vc6sax2ASn/cSA+0Ha2GzUkrX5QYw1rJ2SPcwEYYEgRYXPM+F4Gyvloq
r4VPyJvSqUzoUPasvtW4YHtnheg3BrhtSNJjV6TtkzGQ1glsBQpSfE7O1l0vTgROZfbs+uCNMzh+
y+4CjhjMT+kLeasSWd7nzeqE/UWBwy2JCUBKqF4IAn0mdVkLgBFk/hTv0SFLH/0zqgWoFMWkAaY7
PHAAXbQiRGC+rn4vFWlhE6L4zA+rfeC2lUp5f6pigCPF+42R24nxCAqLYnq0vtTdlBKij88oWTXa
F6Cj0OQ86xYF0ieWu6DBmwtdA8oq87Ux0LDs3nVmRVcbfDJtdGQ+/9rCh5rCjUlML0Tk/RlIJKHv
r8EbwgnDHsm8OYIl4sYog3TSgirk3y3n7FC9VaKAiHqMBtn76mozW3ji4vvFxu/myKRYcPRCccEI
99qwMr7pRfs6Rh0aJ4eTGKsSAgho5DfwQodxM8qAiqYJkgK/mbHA+xzssT9RWjXKZTLWwrsiAOPa
uSYWWgHiLZJf0t0a64WMRaECGotRA4BSRUrqh6X58KnYiQa3rHaqtdYB4GWhhUlOEvHq/NdCn2zK
l2f0/YCCNYP+fk1BEifrdazpL2YH8tEf+QtN6mlL6ecOaSAk/fBfoVQhX25ysa8P8cgq6JGzvBqR
ZG9E/LDG6WF8Ttcu6L0emrRiql6SOuvuJ/OXGuiqQtpYNXmu5DaQMRmwpUsxQCwNPvdnNEMDU839
uhrt1tvmiJ4NQGPHasLJSL389QXFxclXQNYuLRaj2+hYD+r7vJqQXyPs4Z2gBt6AYsvvNKv3D4ll
gXA5/cuatmLDxwJSIpxE2SWLF2Dx3g1ddDCuRLPTxs8wUQ63jczp21XolQUpjBFrrKrSIqJR/u3m
7/USd46QY2xcfMHsFfySzwU8Udql9ACg77PgTPXCToFuUH1jUGBSbadNyBMHIefPozSw1vKg//Ea
5sKinUI6yCQ/t4/mK1r/n53gc8D4UR0walcjXQ/2Ja/04vRnzvF2SFBeoGZo1tzRHAyS+r9WcWMU
8EM14jhUAWj3B5jyIt81Wi9mt5trjUI0ON5oqmox6qm/WzMKg8pJpEXGHwDdJBhwQd4S49kX+Rsy
aYpAf74BUGCH7qHJbqnSVvI1n0mu24jW7gkNfiVuTGzSEFYQCBHsGwDtkRFAjU/5gsLxlzHF6ndv
Td6jWcmJh30k72ORHxOJ12BCGn5vTt4xIG4SIzf1QrmJ5hZPDaUjBUgfL39jQXbyc6/Hmrm+ng8H
rWuU1nMB0ECKdXf0d7S19ev/KKVSfowYIqk3i7N5duErzLzhf5n0dG+8smHd/h9Nn3YIuJyZmjha
1dVCRRp1sBwIGU8ig5axFDTodHd18mmzJWnVWVSVbkHvRlt6ZYYCnYBnSNhwhs91k6olqUMy0JtN
m5ttCytfv/PcRnC309noki7rldZz/bo5kjdjR6rLs0dcuTFN1izvzg/MhxKRBvvqKOeT+0Rahlla
rmX/3s+Eu99B7L4xWhTHVVNpp6oFoTWDcEmH8HhWCGa+eplOqdRnyJ4MDJiExz/7F75GI5aSi7t/
EmeE6hS0D2c0bCP0l/uYU0W1e3rCCNJ7Z816NpzJ42ef4Pp9J8288k3fX/wICmhRfNRmZIs+uWy3
ADmKuGt5CMTEDn1AQYpmQTpb/oasL1xgQeV+GlgYnZRPryc8G+XmcW75mDZK8bIrFl+tYVpNWRX6
Laf54q1YA4MDIcPErt4P76yQGQAvHFQsQZK1vpJ1hIYJJj1c+oieaF6LUJVTO3gC0DHiIGHkEKY5
wzIiy9tyka73ppr9NKqXyhx5qywvhak4QsZKsMtqp6d96QixC6he5VAut006Gr2kqxWd/C/qVRV7
YOvLSdYi4uYqxhrl1unyMO2+46ueNcesyTXdT1WC1fzNj4W9D1YBauYbYutXo8AYRYv0Sue5kK/l
KUG10qxOd/tI/GLHsK+PoVxqSEibksmjl53/mNr3IJgCJoOwYdaFqZtvnXYQBDYemTDVpJkIhJK0
XuemzKO8q7ygAE2SFO9E9vk6dAVVI3j30IkyNRfGlpbaFcbopTLk4LolZ6dWxTp7JDSPUnACBZDm
Cf4/yvZnVBOyZBS9ia8x1PhxAawVz3Rxruwz74R6etoodqGjcaua5CTozJf2W9gMEAtNcVC0ucPN
oMsDRsRqVbEFQ61eN9ij4hWdNf1MhIbxgiQJBAGZNpQSkaoRKIr4thL2i51iLfwbyTQ4ESOvc+cA
DnzpwRzE2Ep/LrXnSm1Mjqmh76ATmpbKtdRBqha0kaDeldRGBCvkJLlU/9yQn+47e7qEVr1zeory
91+2xa58WMhcyXj3IkCy/z1RGTkW2DInz0kSP6HDAcfxwRBwZUOpYEX90DPb6HKl245IevDwHvpD
VXjNaqgjWntD4+oOrluu2zvTPidxxVLAat/iplJyRQxA3XlTNrZDGGPm/NMUyQo2TAL80QXdQ7eT
5oZGIhK5zUyMDRtafShEq0HtH1OH9ZmYNYmV6cnKpV7rq8u2V0BYAyRUf22qwADaodbwCAix7/OU
E/riUFPLoAWyuYdD8NUrEcD4uVfOwQTVpkk6ZOmiFTip6565I7BHvXTfk+xvCAOxKG5K0mK5AnvM
AsUw6+uXAnqTb7XSzziCcv7LDvcZPzMvNusnF/WivGow+RK6wkP8guJVV6DbyKhUBFfzgchJaCQR
2K15etyty/tf4gXTfZMRQSTe1amCTpIUykE4wWTw7yKjC9K4/8dL69syDn6dHQHkSfgLYIMMny1U
TaBgr65f4MY1nm/pVy1EHye/QntofS3X0IM45QmJgySnEwKglRd9Xz6hjTeHiObeQdD5ogzyGHjK
J9BT1REnY7RmDUmncGCT6i6IH6mO6dwwN4EFWtFA5zgirbwPx08EnT660BHJJQm24uZ3hoG+L2uc
P5Ck0VXLNTCUSlmwxkjeHf+9fCyWF4K51XnkslKqAGEIbBo0ESO+Sx/urAYkjJqaeVSZAjes5urk
7kmvA/5Haicv47C/fcHpO9jPB5xMEafU4GFqk+p9WcZVx7GGycGVVGlk5Nro+QWz3Sv9V7vZGuSS
cv8O2cq3VQKN91hsMi24Ovr5I+PCJ4NmyiQ98mP20zjO7fOWPBQpFcwzxOf03+yHLvvy/R0uDWyD
v2Ksol8kgYwUsIuG24Nk0raUjuPMZ+QqLy5rl9kKCAlHsRuJ4NDOzAr4VNjtnlFuqrdmtKV1Jkn9
l5UTsRA49wYqq84PZtHwnglirWWD3thaQYUh74OtSZQs1XQyA+Umo+q96BzU8nhJwV7OrSWek/9V
a7i6ZlItmAQ/gEHKfY3nT8qEChrXxxzH7gehYEy2YjHhaY+CsTSqfD9iNUprVKip84WAl6Zixcka
bXmriLIHXMD4+nEF5dQsdAaq7uVNLfLnvPVVqtuY6arqaZNGuM8iWz/GrhDg+4f+dV6ZRJET3vxl
tO87yxhkj/dhmyqKtwtXbgl8As9/4IDcU1HBQjIkXTWonhQ6kIYQhOzT6AbLwZEERr/RQnChQ1La
+oPLb9yil7m9yh/SCU7v3mOMn3WJg4iljbKztLPrpVsT8OvN4p7ZMW/ByFeImj8vXKomAr9RRT5e
nNkSdn531bPjaLoA7G2bHKIDIyrF2CAQmEUfFtVOE6YRKbkTBod8v+ckcP99tg8+jpJhTBWoxBQd
KvbE9kz5XcSKcNP8VoRPrerjYydCAUznIeB1bemY0D39GyGqlJvh2MYmun8Nks4CPL+7k+rJw0Qa
lIcbKtGSo1mGkbvGUZmbdV5imM13eMdlbhaHEyinDar0bf1QjIp8sTwfGEDR0gyVfHkRpe/0GR7S
Xv9a2oWDDfbJ1jEtWbw2qCG3MdI0I+bxebMp7fPasrP1BKlpYKB5vhdGQkP5A786NxbZD7NYtHAm
LfXx8jpeyS55wNaV4m44EKW0xx+kGaNhPeeIpCrDhFqxJ8m+f17JeBitTPfbJ3qTVkDpRwQeo7Zm
eFKn5yOyWsZ1qGVLQDgqxRY+H8BXls5kpONyWdETqGciKqPKviNIJK2Ukl6EK8pOj7acgfHelU4j
LYW0hjLa09wssM+Wuc5aIPWTgpwf/+Xpn9YJxUu/FB/6MXF7ShRap52WgLOE/zB39w2ZYz7s4wLd
XJ2WAaZpH77hYE8r8IJaMoWkp1LQlodF7ovTHLPVdD4qznWRfsvVZ0sSltiEcTb2wuu3/EA5UX+n
6isHLdp52zs5CV8eX9PxK/wTno1mmuOhMPYlPFN1rjQO3s6MwdGj8eooEDI0Dkp3hMz133ewLVV9
q8pGaUdVxt0L0oZNLYbhizr6Ia0XGn5/F2JrnPHof9J1ek9RQBNypiZhsDE12kguBzDYqrvD4WL6
uLJuQEoZXw36HebjlwTEY4XgG6vB9AMs/XoZbJajMxg3S8Z1+1ai/5ic28rwQ6lhGR2yNKDCnT6J
cYSHTGnnpJlON11zKvGJT+85qnDBLq8j97X6YOkaXDgG0Aiy7Uyj8HG920YP5nCgGclTjJVL5fQW
T3hwLgqsko6mNeaHKy6xTQWRub3IDC5Q/dgbZNj9Z2l82qKZlkpRLKv9EUj1T/eP4sZCHX8VwOaJ
pK3IKYGHt3ama1WPmeF5ddHtAuBhU4mAVj9zlOOaNx7D8z5gz3Ke2PGEUb5H+ReDWhi8OLKLFRE3
upIhbIp2c8yKilgFf1eDFA+/uhcb9qYPCiO5Z1kw8ruukPZDBGdrA7Jgs9ZjpuiD46iI6wbuyVri
96hXfv71yr9wammBwT6YP34VSL0k/fcF5olW5H+Nut0T/MNJBrhdg+BSRhPpy8v7ZnTDtwfS9/l1
1QA5bvQN4587eZn8TY3ZPqOGl/fUNG7TjfrGwoP1I152ZwN1OKS0tpVqB0J389NVdaknYb6Z9Z/3
I6bBrSBN6gbKfloKrzGjIDpjITYZ1rflQxZOqcfDZdeMN18hd9iGHcYbPjrPW4klFjD91aB4rY4d
GjnSqMz1kW/+8JroK5OuupFWXgNfZiu8x9ti+cRi0FwoVqUVP3/SGb59lLY1eqrvFsBS75lnsa+D
DB/J8VBD8O47gmGZXKRmdC0W9m79ivbkU1txIMuyaA+9nXDypPUSy24W0tdOQb+tWe5wMXmPZ3oL
ApqBJE8mSfSAJSlThm3CpC1CyEAxKMcxsNUCWWQx1vtgxYHPCnmWaCRwMh1zXOSq24eweS3XDAG1
zguX1lKYuRT+mrxrnNq/Yh7g8xK4wB696j8FAUphLw5tN7f8/bYrBQ90/gkmHe1YkXZsfmZH2pEd
Ml4TD8gWDprYIfkOPkenpxK+VdBA0AYC7Ggt2i+VHvY/Hp5XQCVLfzoOjD9JOzIW0UFjUaXt9r+V
qncb2cbdUvvjLSLrER7SzT1YRbtl6qq1YpNJ6RCIjM/nafc/SX5nBPY4hINVNBvlmwNlcTl7r452
Ue6EO0FUWQymcWdEYQrAL5oLq72CJYJbsoTIlYlKeHO6NTs4PVRCSgVh2V1+Dwfc1MKfITKtWXGp
V99sv0vh9fU0olyuBGhRA/I6YmKZE4Bq1SbAeRFcqcqhISM7p5iY4z/icKyk02vSY7XVO9yFsWo5
gh+Ya5/GZm5aDSHYeNNdHWD6u56D+gzjEuOAxnimgwB53Jo4xrPWA+w1RGPewPV+p32GwAX6MQw+
xQD5EYeWe78Qez7kqdDNGwsyIItLuo7VnFbUR9hHuD3f7wpJ4ck1WIpo0ieJ7dLuEbkT/b7fALuZ
GQPSvPgUZ+Ctb8BboX0+k+w4vnBfquFDBc3/f+24UGVL4ZnG6v/vtVMoDyPd1nCvBffCeQwb7+Ss
MsBw9N5n9fdE8hIEP4koElcP5IAzTFChcT4zpXSRZsB7scyUvRAH8VbhjuO+BZVC+LrbYygYOIDz
V4w3ib7TTViPgZuTFub5kM7JYFwSfy9V+n6sZqYAZiC3rpXMRJ14xmxlnMKchK1oJB8Y6BzrAg58
6FhIdaMjt1Uzi7SEmqI6d24SFgkKzFJ4CX9+I6oBLkE1z/VqsDj+bfvpDM+ggYjRvGonH0c8HcGC
7fJIuPTi5HO/KSB6mOkJFQGokUxIE6DGpg/DNvqI7LVtPUr2Fqk9vW8ommAVJI7tisuimVjla75g
8ggobNS8b0Deyu7mGWwkI/Ydtt7gDOoVgdx6xItlfkYkc0Aa+P6q6kyTGVsOIi1MJPmXTwqMAXvy
18riS1QUixorcQGt65GBpfStkROW6nRIFu4n9AyvAX+mEhkVEDaoe+esJn3jSu9wrE9SrbfU+nCp
Zw5dfygEQBe5HcpE+ozrULOEgT4+fAORPpLVROCe6EDXEuZ2ZbRAgs4I7GTrJ50b4VHqhgL1n7qs
wLpOnOiTeVp11KfnEt6hhG54+5AGHV5ouI2pLmOeoRD66x6zThsN3In7a7lpbAmhO/m9WrNLR4Nf
Tm/D+Iqv1nHB6pCMNnjkYhlAYnKaX7Mjis2deYGYlTDWVPzuF8Znr6tUeWRnEt9r0+ADTKtJaFUc
8Q2MfU1MPi6v8/kAPuqlEseiGsGQbvEnoIU6y6PgcckcONLgo2m8HV/Afh4mF9LhI+P3qx6cWPLt
mfOWmCxuJDK8qR9aSk4ee4gkNtxGXltxW+gye3lBRk/ltmW38OvsmmsOr4iZ7eEBAZc2m8SYtSwx
vZhT4pLIHMgd6UI8e9xl0uU/CsCxyn7TO32cpWmNX0vjeKfNSpoWlDTlKkdpipqVIHrDtgIBmHDg
XzoAUJwqGqIq5nfLnlrBemj9nYcL/qrzcfhRGOMN2SDUcGUhQprRFix9qs6FQRcVqGpkH9r/jznU
YHHNRGn2q+mEpAmIx9+fFFKYpQfrzoNws502ilgHaUqZv7vRAZGFDob8ya0BbMgpb4MQdJHPaH/C
ivbw+DBWgB1TUBs2CbpYLUnlfpSphdFCp/psh0IVgFMn6Cl6o+92+dfRxk7tugGWrC5ZJcZResjC
sIEswOad40HhroVGT7aBtDNla5/soqrY11MU49cKF04/WFjCVzNUCoegyoItlJreRG8C7XnojIKl
vb6mS+M7hsRgMl5SGefhz64e1/Nk5Pjk+tMq7mhRZ5iwAvZYHoORD6krPDCfb3UnpxK5F8BlEWKL
8MoywrI65GwZPmHDcmbx3BcmPrb8+f4lrRWzNfmk+DFNiVBKSHW6AgkqswHKoCrMs3/pgowF3zTH
96aMF4QX6JZqDdmU/xwSNlJFOX88sNeSOv6MdN8t9t8w1OJe17XiE4rS/jXHUNEbWQcUSt1z0XTn
aDYGpajDgSMhlrIrkzhm2Jq55ctnxVscKAoL+zRsPPegy4MsyGDV6bCG/NHGrZN3KJzN+XWxNW63
9nyN2wed3LaKu1i+bkM3EQkKqN1ua8iqrab/fwA1AbMLq11FOmgDbSuhlxSNGRc/uYR0SzbIxw1r
hK935zABIQCmMNf+NIxlmdoh5Cw0P9rQ0f1/E4iEEpDo2z7mubHfuTfJ03+9kWpDUEw4OAG+V3kX
vMez8Jf4T4ExaUiOBfjIhxBUciW1AunttblAJfFE8o9C3Yfg3yfHZlHpDc/Q4KKsZHFhLf63rPKz
3D6MgOqZZv2dno3SOSZsR7QOOty9YeGY/tGWcIlmvx4wLMHpyt7XZ0kld6nbVhgP5x4fyBkvIp18
kPAjGcQiepoKsNACQ0s6Sm7BAxDH2QWcK3+viNbq4KgSF2S5TCBvoLFnUe3HTHJ2+Z2fHH599JRu
sZ828FDj7kuarD1gEJVhh/IY17+W//7L0vr0z8X/E8L1A8gunhCUMRZmvY3DVvd0WuHxpsbuGOVa
PI/hqzYekgYaeLkCt4AWOMOQIxov5cqz0Zmri0F218hseWqzoY5dMiMLvN8l281JhK5nOQV+6cno
Ym8P+qDw87jr/H9UQvQaD3GTgtX7+BOT8nlGNRkoREpak4iIXN1T+UpJmlHomDJ0ybGqUR1I+MdQ
8kfbYL/wM28He0p6que9nsEb78VoBJZ5elfbt1zxsjAowt3L2oRxqc+EkpZUPjvvfk9Y25ucB55X
jgTiBml/1rc/1UBrnh5boS/6hOS6Wzfpwqh7moaeGSGyjEA9oiSLT2ljruePaXweR4Mr0k3IDglO
F/KqfvVXWbXuovH1we2px6Ohc7aoZPWZDSEhgpfZHE+RxF4p+1kNY9ZHRajq4zabJTLxXAmPlJ4e
vbNgxjI3I1WfXsAZ57ihECtR6Y05k6j1i1IASnJ9jrdQBYe/f1J6sXnBWXAZQIgOHqnNezlHcfCJ
ygwWU8x4aO5bWPrzxIL4jZjgerqRmUnoI2Sb+sZiMvg4hOnYo/rMJYlFp/1bgIMUZZMiCk7c2OEU
mimUwZp9Y1jELIrQcaXSZETAGZaEs/7rJxstxnQygeU7isFTm1aRiqwU+qg9dQOjoKTwneuvQ2jK
qWpDxEYXBd0sgP9mm4bIF+Jz79Y1udph42SO0FNjGRQBh1eL0hb73zwkGWnrtnkuQ55yplok3MhQ
FgKVKVox1pDCxyEUwnAiLNUv8vBE/p/lns57HCBLvCFYnZmUuD2K/Un9TK1RQXGwSGcwc2SLuKra
gztFMtmOeFVxIVNqs8NbNm/i9KY9VOlwPqj+ykiLcpX6p7tSygBowPreu6vhGSSbmrNq8auAMJXJ
Pua+pUZSbYw3peORIYP0TYSf70CL1bLzPIJYV8Bx9M6mLixXbM90iUXs8FlRNRT6JnALEPlVFtk7
hN9O/Pm0aM+h/4u3dwKMAW/MLBkPZ5aHli8D83U+YVUpZKjRNyRoO3MJ2iIQRJqaER4vl/sicbrV
CmFCJtVwIYPt2OFu9jm6ulXPd74E2uQVNYieI+1wFY3ZDke1NIM4mCwE5yErWTqB1cJ5pa4QYbth
G9+MaksLGODAPi8d9R+qGSHGUtgyF0DlHospl9eH6AHIc6dsHTIGz3Jly1sD86mboLomvyLOiHRo
MJ/jHcs7QwENJzx2xlPvKBPFgrnjXwULKgJn++E0JWD4EwoeUl2dGd3dVFDih2BDPpPHWV5+FdZR
51fH40jsQ7UHulMVmp6g+2Vkdqp4Ko4oAkeqg051DA08ifqkftYlwmvlCF0ESIR1Zq1o2ZmDlywZ
G7OZIyq91D8N4aK8jAdHucOW8MrHF6ySXid8EY7FR9eYlhdSiw8PCRs6SXXeY/L4ce79o9ppG3qI
Yl+z7UBq+nbcEtTjd7Y52JpI+rDPTMu2FiAAkuoKKLJbJjeyF0bW30VUVwKznovxd7IE6LpC57Ga
TGOFXIyWOWekmLtn1ym8vj4ge2gIyPixsVsDlpnj778HzksW49TSPkMFExqWd/lNRVRlbYxKWzB/
g+PQc3b3GVaWOmbYOEsf3gZLOrLY7iHpAWzv7wAoCAwQP57QeyKuBDc6WThQw4/J6TlLEa2GTyX9
JaArXrjasZMCeXJYMz6DW2Y2X0/wG47H+2Irle+SSrmH6/+FuEj8xO57y1SXU4/YEaiEnbjJy7n4
NvqVHH1UUO84yd4GsEkYCSc39rUoFZoOORuHabIHGWJ61A0dnflEjD0RhXy31k4RJwLAQ8VkNPSP
/ddAv8wjSgZlg0+ULN/G1qZaa2o1iPM5GeOb8HVNJhuPJMnmL2Ps3RzTju/17NvPoB4LoNvzqCtc
1rPxblY5SQVvRUBu5WOfNto7rEW7Nww/aX1uyfzTQ7HRBuHqib2Po+pw1p1cjjoJTrDODJxs059i
vW/2EcgSn2CghWDuRy1Gnm6vR1Cmj4krUql/i4vf4lBD0YJhuPAPfSSzF212fM4uA1qJQCt4x4Mo
ArYMDgDo0GukUv9dAshnHoC1BcR1X24sP+Ux5Zkd55lRlDGtsrZU7Vjv7g92B3TvTUux75rnXTJW
ggBVv3Owihh8fap9z0i4rGjF9ypYbNU/NcmDN8H0EBesx230b55kMeFhYE/eGI8ctRAB0dEE85z+
4X5Kl569z4+AmTqPWIOxHM9uR/AnorNhIgmdDjfo6JapUwW98b0dVmVUPv1fWQqTy6MS5nxTnTrD
j1KcZq4bdoisp08i5E+x00vxFYlgUKRCx5dR1pXmlB2W5D0h1/lvcU5FET2wbnIRRO33RfahJ6i3
CKuvAAzt7DcDqR744R9YuVVqBnGYnhYWRw6eAa/0+ZIEZrKIRROczQDCIvN9tT1qN3SvkJ+kK/dk
E3Ab5oD6KzfDHswW9k5yRNRyHGdq4kFNSJxi9kBxBOVTNluRRjOJFK0o07RocN45Z5VETpaXeMYd
X4vmsyY6JzEUvnlmJQWktTXrD5qBIMijNHr748UWytm2kD1+MouaaRqQgTHBz87RZdSb0ByeQ6LX
F1/bCA09hywNu0fYSwf/MA7Ae0JTSLCF4+QGA8WqRH2Xx4BgJky/Si0OZie+IUuxsLu8nTfhi9O6
dbidPH76mhvbLIFEcctXPB/yuRW1jifSUvhHjnAF1YaOWHqybehphMCmexkZUWodw/BRA2e01rkz
YJk602+2UsChUcLfGAbFUhqaBBBapxC8zsbgEOnpuwj7x7+3Ufszq9+r3jt0d8J1S1lm9U/xVbgW
oojgpU2AuApm0GuvFSIvonrOZ6J35PqH2lzZ3sPm19pfi5O6oNQNTb3tAVyPPyez6te7wySvyi8q
TaJwY2xvXnLZ3Tf2frbhc80fWApUi+ci/LM6qc65pp6X6JcnHqPhoq6blOrPB6vhFa3/y/S90P+j
EiTzwLyogXC7upeUoodjPvb9Ai6FYQe8wKTLC4d9khvB0+zxyAGCEONJk+yTgnLIr07Smxau+Q3N
AT4tcHhdbTitcMUjH1u5YTAjEovTKsYEfk4YCgylob9Zb37NcPBpVsUzknpaokWOU6/qTZIAPc+A
+kABussSuFf7iyQN68sLAREkT6vVaA0E0F5eADgthB8Iv8Pe+gh0e7NbuC75s2RjnCOhRHvs9dIN
FMGL33g+o6d9fPoPt0IeWhPzOwI19eE1Zsgu0lOunLrNe/Q5hMV7n+0WZD3Pk4fIct/dgTn1u52F
N37CQCNGhBSSx4+7hOk+hI9tbPGxEqj7shhHe/j0IrznMU2/y6LCtOi1Rm+jv5RiOiE/+ctv0rKo
TBHAxKV48MGRcntbhZhWVzePc71g+I5hyx3wZJ6NkF4xEUtOEHBPM+C0CDyRoxqPZZh7XvYafw5U
Zoo9HSc99vE/Fycr6Ue/eOsFj+Yo4QwrNIgjg+UarI8sgk5HcECNtVDFILg1IA3AtSgL9C5y2Q2B
1o57SN5NiJrAe+OomCh0Fd+BuAagrkm7et9fFMvklBKkPmN+qIVEn+LY+EvccXuZ0ITuxTHhAFEf
uWDmi9dAbLiEWOU6OXjrhCW0LSLigId8fRHw87XppKd8vSO2B33q+S21MvH1cw286A8SwYr3GKut
cfgqhIJOYRROgYNzFighfuy9mG7cumOEqjUnN1XJ8plv5TgVuv61giP/E52s61R21XsBHbceKoLq
0wyCs3yq3Pwz8L2JU2Sl5S4wxBOSZPoifQl1K29M8NCEJXTj7dmlNr2JlPlBPV/whtFscxs+OwLi
S+/xFGWCHV+QDNPDzpTEZTrhfJlW+xQHlpICy5/oE4tyGvV6HxCLMaCD0w6OjHAB8INmJKHadAif
vGxGx9CMZqtFtW+H/o2zeGpaxjzNif61MyjHRmv07ha85cyU/WLwpXKxsTVzp28O/Pj7mnYbjN2T
nc0kEPu9Y8rKHkvul9wn7373aCSy5b+EtHWzGuH41dTKv2c2Qv0+uJX9ko/fsgCas4iHUxP3FGcN
g9ZDfpPc8I5RO6Aha/Vc2G0WuHluOYIdLpTCGkld6JBaiM0n7mUhc92ZD3dVcfghboFj7QOZLmqT
NxDJS7iAxqdxMx2hLvTElzid48l59+or6wMx+mRG/rPRfHmMLr6Bp3eUg8PjoRvBNHy83u3N/fIG
8SnrliG1WLMb3FbY/5sYQkqmb2cvQDMhxth6y/wy8E+hImS3jeJQ/cVOOFcW2EftKKmIrYHxREXS
f9cWmQPpdIKijhyEoqHz3pNYss+dfqySAIFYnW1rLLJ33DxBT5ousV+pp4pAMqK8bqFC9vsbfgJm
Bt3xydmQ1Y96xlUXfRZRNPPSC5Momsm0s9Z5UqjED0/23vI003q62GXGcZiHVkZpPFV7/vShAkCc
u627jFoipLUHgWyo2y4FIAbyEOOy06C5YUDqLEWPMV1SmZMRU5D9mf4bjOpISeHpCOBq5mAPfDYS
yJuAe+8YxfUcd4OVp0GYrJix2X1QnwBpTmkLAiD6rA4F9lOYKmqb/Tln+IpP7AcQfZReebkdS2X2
jwQ7Dbbo3z6+s3wFuzJTVkWlAOmtQbMiC721+eKtznMpAtcePnS++3zZ7XZuJIyzblUZQsKnvX7l
r31yTjqSsFD0iESuJAdKsn16eEGBff594Cf1TOtbcmwP3t73XTecFjZjyRZOHdIWOlCovjDPWCHj
4auLObqC2RVxJ3T9Qhd4aA7F8VEMqlrWbFHh778o2rHz7TW/SZmkGIMTUviQVgkL7xYw51p+3jhh
RTwe+ydnCvxXdAEi7VqMp+jLZcxf+XMBHc2c9V6YTv28g8EWXLNwldao/xh6kwV0g6nERj/Ycc2w
za2ClroYr0FAifwnQVHcaycSgVAeL31OYstHkpmMJaWlTQ8ffLiyfaeEZ9dU3Pdpabw9ayPrGgKi
ilBWk9VJb/KjemrNBPT/YEMa/WLHSAa6nDuxO2bYrad0ahtKChUxj2UunPbnx8Hym/8xFyZZvYx4
bmpMB3OYVpvRLkR76Py//CDFkUnyNWvfhS6rg0/FZX9l/bGf9swVwN+XQ+I+THnlffEPvNzeVArT
wf14s8zagavu+s2NU3Y+EBJgUEzbcvrHsRi/yIzWwXSQGfBglDidoL4p0NZYbO+lZQZ/jJYhAuvF
xaEvc8rSwFsMANabQ4Qn+Bx0sTV7bO8xxXEI/cUhAOarCua7a6PislGBTamhs3mdAAaqJDTTsD4V
Ha0NQCoyZ36WJZEi3memVnthfTw/SyWCmPR9W77QJC3IW081KMI1eMRSORNLU3GSeJr2y48/vApG
+LJEfH0PqgC5B0+1BmA2+ukHARfYfJKpCJh1dLQmh1S+CdtwqUjGG/8zqqF24csw4VwiZG2N5Zm5
0IKaAdlLHEdsa1hrAUPQyykzut0DJCs13Gibs8H2xRZcaBMc4mU1MnX698rrS6XeQ3cnPZpQIZ5I
hR6mLHgOfvmOxlODloq1PVE68chkqKN7qKU1ubkVnRu/leo1t9v8lrxCLFtXjBub5XLSGsQ0Oo2a
PTO0eCIbQ3oqf1JLxlM7PYi8IIpU8yEPshZbH4dAaJ2kYS8HW0m1+vFPIA1biZBo+XRRmkO974OK
byQkgpbucZiBSWHUZqaQ8kKzPRPjJcvQ2r3RmeLIS+HCph9hQJV/2k8WGuCipJtk3FUKMjk8l5gX
PZ2M9t+HmQrT/bnTw7pn8kFfCirftokYI+gaSmUocDoKFnfxE9aISiVvoYx1+ONaop/B2NziGsLX
y5R9iyl5HSElr3EqwEKSXOXhhnEUD3lQF2odCnOOQzaCnaV0cvTPt0cJFNQtmSBZKfTiQcs6xWlF
K7vvYPCFMPoZa0j2UGRMqlyGAxdxtMGj1xcPJpyvWE/tW/g1wisvoiW9FL84svaqq5M6J5AAW2RY
8DRQYVj1FQOrrtTPraEAGS5FE/V8CTN+bUoQIITuPFQ7Ne/Y0+KyN8OEx/M4v7xNWrUjk/T6NXA1
PlcTktc4jyUfk7T8z3L0nQfXmGJ952mlbsHLxOjaK2TYPonNkwPcrSvF5ORwmp7IaLcT+V6/U8eS
Byk55WPVQiiptFhLRSufKkedDIhbke3fnrLrUDPGVRvZuoXxbg6dhssludTEerBXtbBO53T0jZGV
IkZYAmGpAsfsvLOJEaFHDdqdlzk9Ow/uFxKhJIEY3U1nzuwMd/+O+xT9aymjffW7sjwoVHaozr2n
KJmrJfA8XV70quukBHN0TqVFh7/XB+kn4RnQI37i3rCkemunvM6gTKDoX6dkHI4DBjQdTtaWFLlq
fN6wj2/1FS2CW1uCeZpCftb146y2Whk6FdTaVJkbGJ0UXQiads+/YAbZMWGZwURqlDsk6WT0+541
7iA8E2FqMDJsa+yS35Jho1aFwq64wCrDJTiDt52O2i+wPBFpet4ZXHpELH3y1LnG5MxpoFlIObcG
FMycy5KTIg0MX4DjaUBV3ojR+wdXNjef1iBY1CypVqjv7jLo8xOpxdSIVHwsmRWkEvKQ4OAxiXqw
U7iSUCbLkMu8hFQ3Q6RIWT+4ryjfSH/3K5YNNcRcoCtalVLZGyx34rEUK7o2Zk8I4Jzlj/a/gRF7
6mF6GB4UB2SSfAPGW3+C4/eU60O8jY1tN8pgPjNa9X+LgmY9r/9J8AH5jEgEdwTLATxtRuOAQI0R
K6oadkco/TkJfCXg0jNJFeh+nNt1B75YTAtDP7IAfF0L/JQ1XFFF6v9uVvZLma0eIhbIb93tKkXn
qBGsxuxqhT6I2OB2fUu1WflC+VN+UeMWgPLQhRVGNvf2wc3NaKTjidNBc+KRdzspKoacbTzY+dq7
ioQxlx3oOxvis4TTGn3gCLEUwfqvokMgHirk1MxcPlwZf7+W97tJyxlmTNfBYDIgIOS4JU34mw4k
tA0Q9ZLZojINNHrL61SJzbulGvbw2stPL+PfquS6ndn3DK3rCLutG1zx+9/lI+r9KnFutId7RX+R
na4YneUFd282gq1lXqd7+mq3vLmq2sHxgahla6sxMxyfSfoHWXyF/4QXMpjHPJblKohRijal+orP
NmbaeiHcuPkNcDAOQzwymsIbYbcxcm/e7P2nr2HqMSK8/aTMg4ZzrVHCEhzWWOQa5FEpyNk7gmqL
uvQRqPKScWZTc9/71ut+stiguAZqgDHLTY6NJpYaDEZ5VUTV48IZRwJM3oVPd/O4h0y8xC6RnPC5
X+byyLE6xAesn8zH8h/faOSCBRJkZHr53/8Jndyuc8nwNT8GaEppDOGea/C3F0RSpXzq5cxUCzPA
aZfTHLB0NqaZ5ViDKTV7nmgh4mBky5sVNEiuXTXk84xaIDYT17DtktWctsF+TJYbBzenaMf/PXtA
DbWky1912DgYD+VrbZdGsQbC5GWZMRyZw+v08SUq6VVBwOy9fLWaBArFcRnsnx5UOY1FCpepnBRE
CtUBrDQYbmRNaMg+8GkjwlYOuqpG/AypAZs+bOrSsYH20esYAnNvpDKxXjDfpbC1CvM9+uSZ6ZuT
W3MsgoIbzyFQu81WZTWEcsw6/5yeNP8aa/XCaZqcf6Mn5hQHZNegmEMYgPe1/xEirXgHhzMWdN/r
C9ob0poCYaifszr8T18JjB5DnK8UHHViBgC3OFZw6Ot7ZIGdbizzvAcJD4zsKqbNUH+Z4zSW5fjl
XBU4zuzObGPAjM+C8Bhhz9/EZQeHuWGMQGRQkQRr3FY/499kBYsFb2chdB8v/kr/Rw9QWfwuZ+hb
dw0McrbYhUELU1dkmUIWE5NV0LRcGiMGTI4XpuhYvsDjRsNaJ76E0Hl7Jm0CPaA32sg0GM0n0ORw
EXTi3mtewswJNa5SW7PO9yhS+GBq1dzzgBXZF9p+8l6oSn/+jISGZ347W+aWa2C8gyAcdMb4fdTs
37bB3J1yHGAVwYCD8v0Obz1jLn6l4Op0Q1S7cxiuBYPZ/UDnsowRK0B1W69y9N4vL+jWnbjWxBjJ
KYGRtrGjWhFFonlIlZZFg3MNVebbFHmxiSBLqcLNKI3vbX67iHMC4dIN7UYh5eJZXrvqrIOUOIhv
TzmTFcyjCb69Q/2k0/Fzzewyg/1oEUfgtvXhsfQffZsVVpjG71DJXMl6cYqxac4U4HWQk73A/KAn
6faYp18tr32on9enZoV1S049bx259Sb5EPGPNjXbPtx+TRKxMwBw8kWFFGB63MlDdwZnUP5Q+W9x
ndIZCN1v1HTQpwM6z8f8uDLtHD0Q72HyzkNhB/pvzWVxdhqrHgYbqHttjZaqikfyYd656YGgMbV7
kSKtrYJOsVaXSczdROcPQg6ynzleQfwMCuKBOSnG0DD0ABKbsRQZSdCJMfSZoa21gyoduWyHVBXB
YS7dPWTiNZI3usZc6zITNAZnge02Oh3FTiXVNtV2XoQPMJNglfvgNBSJhokJ6WdZP+/pYFuBxQ95
8iwPXR9Ngu719ER8hNlf6+aOognqkAxjWhlzAKwP2y+hmp4bj6pKJO3dpgq7JpazgJ0Llm3Rvv29
pOjt22o+kOKd0b48AFiNNKetVCd+DYO8zMKF5jYX90hBO4ksv0fN2qCQqyIkV4A7ym1FyVQDpQ93
YNiXErfeBRkzOJ9jyPcIYYHysawFMHtzuMiL46XGFncezT/Tk8toASTSeh8epRbcbGrTyxLjmEWk
PtsHsj1iY87g4RAVDo7ae/1tKge/6aAcNeUCb7Vc943YgYaZCmtdK1lziDJqSM8hVrHaYSxLD2Pq
PXt1omgcAva50KerA6RKUFNPPzwqJm3KoAVnyOuPbNajQPY/5UZeNa7WqBfuH6i+GrGZuQ3RlSxW
5uhzT2Wxv4MI4Rg0Q1VWCKglXWsNOaSekLxctkSdNq6q6Isv7IQKQX7oCJFMU5FelpoasAj85+YI
aZcZiydcZFv8Rb1l8CSilOChCI/P7hoXKZLr7whpoTR5dYTybAUz2vyQRvUjpxCoL+Oy2ugh0qbI
kKhPgXp8FPWLX+lA7fTKUPJPfYWucFq1KTG1hDKU5EQACM77fsFkSo9LRd+PY9ikd0lC96imIXve
CDI/zImSWJvP3YLLNpG+HhB7sol1yflIOupm4B/MRQZVTEHSWGk79fs4yHarPhyvnH2ByEPgut1n
ck3gMwTPwUEA+sgxpNmidzoIo0Mvms2WESCZDg5mMKezgYIeafL6FguTZAg/rQ+gXs0icxGF3BGq
wpLO5ZksejvtAgm0EB/lMjDAfN47iCj7SgRgK542qynqpv/ts6h9uqaMfuvKFS5eBHhhQe5nXvZB
5GpmPn47sqaBS958rlmMUADbmKwgdxzBQ1KTqpbwpR3LYoIvre1EETlQDep445lkhYw/X0lC10Zr
AZ9JZP/MeSIKJxKmbrvt5NgDfaIkZlvrx8KMYX4OaP77AhKlwBVM7OdNoH0y1Bxg4BM6a57SjapA
pjht/f3IWe/1zt+UqCJdqkc7eNA7DzWBJKKPGmJqTKxclEeTx50xnlHnLnOIinOxFdlMvRoSdqO3
JM8+7wGcL/zUiuMXw8H2q1Vc7Q3BRgVV3dc2fu56Zsfj11/CTJ0Ni2uJNnPHR7roCc2Qn4VtOoQC
R4tTO3j5XG+CfBHEksG8yuHC/BERtuB852uDKB0VTGT/FoXr5tEQU6QrKjeRA75gCqCEH6myMLUF
BrZMR3p9WCX6DhR629fy+rtpuUhbbuMCJTK84rESIG2rseLHFkYYCchfDuc51/lHtGLuP07N2fAI
8lGZE2I9O8bvcrRmW7jU2SeBt8IzpENSNsLjmKhTnRcB0BmwrEFjiGkQ3ntDKLdpRMKmdvLhaUVK
MHqVcg0duwOBWwzL5HSUZqPaZecS1qOFrt4m8P2jpSC2ADpqtROPSz1nCGvZdLV+RxEOPzMQ9dLN
d7E2NP3ONV1nC6oXwi6dagyrv4f4n9AFOrINn4v/fS9QNBvQew5Y2IGPuuuGbyXN3apzpOMr9gGX
/r+jr8Rj9ullgGZflwkVzolO4CqB242D6N36XtgL6SF+uW1y0sYiQzSku9eRVJKpJesXzvi7u30a
ncmj/XfcN+qpxKZu0V1dUUxPaLYtcz7oUTdiVQR58rihiBYscO0F5CNnRaqVzL8K1GoY+ZKAXjn6
ShPguWKX+SMrB3yPMS8xlhsiH28eBZTkEvBHDp3ezPD4rlCIYlcb+thaLCzBvCV/xT2QvywZDUSf
2lLS7PY6rZ07ZbSEAkLKhRpdV1Iru8lC6cobmz5F9G5l0Ou46EdicuFdHKn/vTCG62urzf63uYxr
FZVNuJua5IzrT/kJrQeCgf+WHc17W6mmrQl5/rvQ+EwZcu1A3wWjhmDOyIvL0tP5aCq/oEQubwuQ
ff3hRhZAC2A91s8Uftu/aPdmXx03E93/jN02rLbh/Er/Hk9TSqi1T2b/nSro//vMjqwa1eJ3xDJC
7aPPg7Mmp221gFwvilk6k7peTD7drXnUKKy2+NtOKabVUvbS24IfMqFY5t58CthL5qsiQ/h7+3Wx
OGrxodsfL97hpvbdi2qzwLeLFHF8samfK+m+YuAfe9pW4wl6Vw2+QcdD3eUScxaQ9Q6eLiPEteUW
tuRl+NutTJmEfQ0NBFgNYH1QisgtBc2H3+9pMAOdKruQiqbfU7GiYr6evCtcq6uJZQXLELMNao1E
DBibQCH0tSG6PiQyPcTwiA9osGmszWigtXMymSUEdJERFc4mJtn9IAvezXz7FGKr1ROU7TWHcGTf
1vb00sVNq8NDHV+md9d4+2Ukme//FQYlhnvn+Yw8eVMdlUTgw8bzMsTG27OAlwOTsFW3d3RX7um3
UeXzKIMFOru75919o7iAYkIYHMefVjfWKjUJqwnA1sIRlPm5mIab5h3FDz+wNqPm9P6qANKTk127
4I9pAgTBUhRfx1Ui6C1cmMsviniXz3qeEAJEoLizreMbg086LLa/KoZy0ePsP3rFJa5xDOMFP25y
AiPjKHeyuJsTF2LhztZPrCZfFl6MsPV6hxyBnPoUUkBsriHugq5FtROg8YD0bvtNdNn3T3obxV0g
/56SHy+TOfGgAAaXjZef5RsPLLF1SE7caA+jdGgu2qGOXVD46sYqXRm/IrU0Dt+++YVocZT3oQYZ
ayS2eWYM9lHyvPcuIpY51N6bDcA9Xob1EG3pPF6o34eim1ftfqjbjVQSOH7lCzVnZcGUW4eO1C97
uxhuWUDWAYSraX12MFyUqVBMcQfGPb3ZPXs+0R9QOHK6J2Jx44Wk2pPvfEMxMVCnTpOdLk2yKYAS
QcaJ3C+GCnyl24AiQD8qOsPz6KdDvferkky2f4A3eif+DNhWZ8HJIQmd7dVb1dnc/+UBiHLqsqTS
6BQqPB6h5OelkhFMEBtUoXlFIZ3mXcdNvgglthCxhgAUKkkm4ZY8+zfRhslUD8mHp2OXaYS1BGdG
7QbqC+6sGKFvhx8BfR3Pdz1AbJPP9G/QoMQm7DIXfxzqnWvijKqwGu00VGpnDanQSwjbwNu9sUa4
aDq/Clvq0mUIeXGpWtCjSbN8/KisHxVdoBp5AdKsLZ4odwnGfNgDzDcWN4cq+9ZyqA3bQnxTZ4fy
gP+BZL6IUv+InhX0gm7SErugbnXyH43XfDdUql5M7ETXH+q4xZNEhEyVUnWbGrKOsSLEDTl+N/Ws
DZHxyOgxyIPkbzE9d1+AfDcni8Exq+ctyY0b/mp6b9xkCqT6vej+wwfSjkjuv3VDSOXYHlmFj8xA
hZAp8ygdrD9uen5DJPY0dgHTUlHzEaPZtu02taf3CZKrzZX/PIv+C/VlI5HuS6Muq6Ip2ByZSm3n
lJHhvLOziZko23XwOcUGHGbXNQrDVRqDGyaqgOikem9MRr1T45uBu8deYnf2DaywMUpvwidQsBAt
I+y+C2akC04LK5lr/WnbmXIpEDW+ZvQcjsM7tUfhDdDn1qMCCjV5EtEQAc9IsvvGLiWam1nEW9na
F9Xkxwvxj00glfsp+pWojyz13ofFt8mJYoGdjlXR4OzotII+H1/FwkTucgRqOcVj45DW9d2IXEY+
XrXNh80Wk3urcXS5sz+svLMK4Ck0dSiW9uaH6t2HWoKNYfMBwRa5yEEzrjG0bWLTDRHhbajZ8/9S
TJCiveD1DWjj/4rVYWShLQZX6pUqoSpUPfJ46zr+aSFuVYNL5VWtc4r6VOCjkZBZn0KXsFNL0tr4
TdUXnYc/J0lRcgYh3CuCcxMgust3KoZm+oRfpS4WfMx2gOxHQFdFKaCVEh2iwyzTp4O1jC+XJjWW
RYVtK43cMMx9nB37TJdZhDD5xtplkw8ycBpLwwo6lG58A8bVCrFRSRBwexr9JB0+jG2eXdbd7sf6
4nn2yZuZ14pFjEdeLddFMKvQ+wYxreh1hiaLGGuiqDHUedp6pdzt9kscwKaJUB6VtPX7/Dw1P7Cl
aSInwDdY/DOaVHYhG1zvEpfa3J4+aVW+XAvEnKhAo3Jckb43oWN3Rgc/hDkh6iH8AfJZM+XirPn/
3bt2Cq002vPaR4corfkOdHIave3kYMEs6RD7IRxG4E8OgAS5s/H+KiLzzgg+QPY4MICz/W8g/rxw
5JYs4975dIcYGzl6jmFuk17igMMdCprziJwNK8fafWZIm7LUIg8xap1S1+dF48tY7RrIwRZqniYg
dgGxaQVlo5mgvYhrujPChGi86Gt5Zx22FrW/apwVX9CishTkNDsTgVcnCH4djCFmtHlxJb06HWWP
MPREgHso9JK4A9qr3v+J05LIqqWPbPphsNslOM7BUqoC9HRs96wnM+6GLMakjIkQH8Zomla4Qg7q
3Xph/o5HWmtmbr8RMvw5dFRLq6+6AYj4N38CEKGmhguV03N40PLSzuXohxzPLaOy+fOGey5Ra7lz
pbOOzrV2b88tU2hQ0oGfrbdUt4pig7Ih4YTrPuI7U7qw8XM/rGmDjpMY16tN2nQcStcFBRV0YQxw
8HUh5jQitkrlTUkVX3Ld9IEQfnwN4XtqwwV9Iim7eN8WuW9MiFZ9kSDXo8vHUBeg9vKCZq57ideu
v+/OUIlgD5SqriCVss8VWt3fraIAfI9As2qNd9GYoRo+R0ZiIP16M2fy+J+Iim74XBPd+a/5mWSh
pvXvRSxEkkt0RFsssQ3Y+Ku43945odDaLkVtLuJl3Pabz1LdpU6MLxXEJF6ZO2uIrnIGlSgX2A8C
kkBm8hPBH51KuMUbf3aqcwGci7yy7i5DnN14eAnHyCFGa3Lehl3kfs8ALLV8S0VQrj+bWwnI/wVg
7TU15nZBM21qSEJ58PcZajlT/trEH6sASujFoPMlC/6hjzg9pqFneIUjH/wom2hgmoQ8e/B//0Q/
y57y6U8RAQ7ldfLMdq+60tQu04rM6cM7Ab/htx4QdIy9acRImKzSZNr6/P22ZqfRHDsTcaRjlFM1
4tvRPvlmDdRfHrs+MEMkGW1+UOGyk2gpzffDbgRsRs8rNw+awWUwZQooPWhsq9r5p3e/GvBJBGJO
OCF/TZ0gUtL1y8kcikz5iZG9GhmMr+GiFuTnEy2R56qr/hJB1s8wldZmw0OztYJqpbaUCA/B0EUT
nqG2/Yfrtx9seJ3ov89tcSCu+q6gS3ccR+5FyhxBH3pt1vcMcYXy/Hz+Eff4MpJhAEnok+yefkSl
Mp+7E9xZooN8cWecUGzMvzODv5dbGHLIPHDGEE0B6UwN3IMdlnH9SZKeORu/nQWvzsOc1RoNMOum
5SLZW8uNSYewX+TpTAYiGq4atiWdZfruuCE8+EfDmrpyya49gRqGd68hCfXTPxFgkIticxJvT/N8
AqDlRWoW56Yl8lFExYbKcleVMesSZFxDmcybXfBmOi9O2nzeV8ZNZlWz+vxgS4VZFs8ftA8HmMAb
PrriT63aMafLKuBAU8SVW3c89FjYG9DYf/6kOUq2xJ6kJUXRM6b3fkpkUDbeksQmof4YACYwqFFd
pLW7vqf5YBXTnu/G4NJTR7qmVVyqVlBQdxw2U7/0hpPMvjmkwbNCSyF0PZHVWQ4ncRVU3SPEU/VH
E7c7HLpVfJyZ0DKBScYYUC9yVtwyogjeDmT26VyTbf4XWOvDvAcqKNEG+djZcbyV4+VAd77Xg90s
xk103x+IhuajaBgl/dw7k6IvGyUspRwkn6zCySG8BLXapqCsf5LB1PktHUN9SbJmBtm12FW34sgT
7KCQ2O3lOUMMmoNdxN0/8yIuSFDS4+j7Gds09QT+pdWKHZeXP4A9UrA3LWN/FqJrPvRv3u/dba7p
Ggyf824Wc1bVpYXRpYwLEkdwUz3GE2snD3VtzHrt+pEV/2G6J91o5L1AjuEgAr3WN6lgCUqPucah
UGkD5cUsL1TqoWOgT3H+B+Nmkfv6Pc15HSb0Rlf53JcblK1n2wtU6aZ6KO91+SudhL4slFSK3Wnm
XyhIUUaTYaEdReD3S/EtHcPu36gxs1oj1NymdjiNI6FN00722dSc9G7b2oOHkPgyf0sntU3YuOpr
VBEBU54f1GLIXh7B1sjZg7RVPzghwX4LBYn9nbFGBI5eToaehJ5zhJzpW+2uKlcPrvFFMpwHV3po
lUmLuM/rvXZI9JznXpm4nu4CIMM9XD4J/8hhczbm4Kd5cwBnwjmpRvryY3Us9y5nbTDWmKq8gKfI
V1imFPIGYmDWPquMqfD0WYKKm4WGSwP6fS8lSDbJQ3IOw4tl7x3SH+IqpKwvom6z+3p2YcsuGQaD
bbZXECqzLy6pC/sWliJAilAz9ZL7jOP4pQTJmjjAUIcmEDe2CdAJlnq6e31L2bAFytZinUfZs9sF
zbJgRqH7AOGR7stzsnzcFPOwuX4NyghtvqLHggoA+icvUVdLcB/j0ktumVzYH/9DmlzMmBAHtwLX
AUpmyIsBUvp5Tgbkf1Pv/oZ/RU4mj2RUTBWbVS0RAXa6pfTGcD+xLDjrHhWh29xvGDf3EZ65ydR8
nnf4RAfnTAIGlzWx0N3AhymumDLY7092973GH7jJqVuqwMjP1HQbcZOvV0/LWyj+e3d4Yvnip6/Z
wYYZIpk+AZpNy30yyAIN9bT4jiSHSyCAK1k2je/UP8P51GLbuPyMhDtLiIp4D/nMnTBhBz2+Irou
aD10wKAj5YM9PTD4Drj+wB6tw09Y/wo52izIs3qbZkYY0uI3Q32UpcOOTbyHr8jF0kT2uTNQvEvP
FuwwKbR5X6TP+NbO1vHioVJQpfIwmMg4Zejl4VgJtOJUQsq74GH/SZ1RF3eaD65GB7Yfkcg8uYA4
1gwTPrmMwO9fwy1hEIQwhiHJX0YKNRTIg8oV554gQzqgEWsfQ6hiS8acwKSTC0PfmW4HUT17RJAp
h1qrWhsjxhTb6iFiPm77BN1WqwuIQmM2fF6w++Ntfxlfv9h++2M3uqp9Lj+LU5Otum/8SPzn1h5/
e4ir2xUIldIZ5VROeLCT1aA+rkIKVS7Ud0wsbOVhQIOFcqjFozHVE/m1/xe+xeGK9JPz6FFYjTH3
2npoixfUzmBvCnLUiiCIy9LXW91rtTe5Z/56VyHKCfEZbgtWOqoVuplUu9T1jRElgx5yUGzzXKdm
YHhekBxpxYu/c2LEMmxOLK3EY4zRDciJyZdiUVEk5Ka5fiyCAk4r6m5FpeeJJ2HXIyKDzIYVP4uV
WlPoxqUzovBZ0axCN54+u/OyRl9nS2/1h3Q91h7x+9oDSy+ed8jat3VIAG+zqa2tUnGgV5fITKIU
0pjWdf0oXZH+PQzoDNgGi47/HhouJrk3UoyVGiKnH0vrfqjoT1ver5Kpe3zwvEomSF0SSdheIn+X
6z94SRRDXf/kRL6xw+x2PkaSD/m4KS7AdqKVcn/zD+CDBG0VIsNl7yeZ3Y4k252BgCh6JSRGDIe+
43WpFUlh43JuuRTIoHx1SK4jReqOqmk2p2qh/8esUqBbzFKsFhXyOzvGZV7Q32p/B3UvDvB67qX7
6ABn2K8QkoLqGb6v4zIUkCxQ3zsRou74ZVKJNVobhiX1kgk72ZyOyinQ/NIliuL9RHncuXGW2iM1
M/QeUyZGwa7LSpP1yfveWzScjYPbbOop7+A69jBcZr6dfROjrGUzma9SzFUcrA+pBFqk1XJxIPQC
fbXwBGY5JY6cwMxG5DfeAywmf5BcoUdC++aTweLNot0xmH0jPCIvUmNoh1/4GLelV3eBgDIknV6d
8bR8XGeqKeMYYkxtrQKYw7EN30PVB2TMP3S0PSEegJ574GLsJ3LxIBnWsaWq9CMexCTeQAJ0lJKQ
jLvrqf8L0Fc9S2K+ii+7kJQrBT2M6vyF0+OZLYCodbb9Eg9DzNN+q7cP10Pc0N+FwTLAf7f0Mo48
fwVgkVDiep9Q0/2kellGTWck2ldMrqkIpK4Qf3gK7Ly0Dj2jppy+h4h4LBshnkzo06vawMeCUA44
AuH1rYyXbhWaown8Fi9dMy7fslnFw4DQhPMx5DGHl04cdMcYEXwroxzywttHS+Gk70Gmd5yrfjly
G6HHdxcsxGKhfrEOhi5g1zr730dEZpQTxZIF2ksE1PVPBhOWo/+PTyVrtxK7JtjoWM7ASj5+EK9V
Om7c8H19hpn5K4nMYK620S00SKi4ArJ61nTYsD+iMusiyomFsDiasQLhXmc/7O0hj5K8ySoAYpvx
15AEnMxtXpjm0i3pQ2SlmfozaXYA+IOFaWREjZ8IJpipUM3wwgxyX2/KJoaW1n17+Cz8m4v3yCNR
ZDtvcGkgO0gkhRT5fVES377DnjKQDE3pOgKB60EUOhtBj6Zqd5QE6OfVxOSKDDYuxxbffPlt/LoG
hFNBtzjPeK0W2PVeE7fRXhOhuxWSJzAPV6AWp/tq3ceRLni9qD9UVvBctkbLd54ZghGFFNX3ghcl
BpVqu0kyKkRqIVGu9i3SdfKCBdCJLcaqbRKlpqibcdIdaoWmw32y5mNocMU0BmJzIB/S9C58Grvt
XGYklzs2zWIPhMo8b0RuB6j26bgsHhPOdUHO4jJq6ekYvFY0LFWhvpG3aqic/ZzZSYdj03NeS7R8
/YX18RKQJuQA797iuy0EsAvDHM7Pg26mzsANifcsyhVli61QCc+/7VlB9hiEuimhnQ/vsaAcBMWx
8Wf87mJTAkjkxt4r8EZI4C9Jdqan0ac0VK6vijEqA7v0ABz7Ezb9+zRfW0NgCgkzgog9zkz6T7te
Lxp6g+ivbJ3yLOJIU2mkJ+pdKfAlejH+qWD2xMOh8a+znElD2uzAwmnAH1o+7B6m5gCmJjKlcSc6
sA3wNZKM/Zq25PREalMFQCyU7cnemjH2IcgXLbexrHovlcPgq8G2531WLc8kHHzr0JZleQttGOqT
tvJR2XdyJhOFfkPUsSnMbbutyhq8x89RRSR35UvLnqGaSF5Gi5k4JjOKjw3U4gDr/loCRMLK3acu
Vokk6XU5iyfneiNKf1UGomjG9dBBj1KLtGrn6aZ+sMnE83QiJMCpHOpnbGFPxy/Fih7vQz6eQOPF
LH/FtaBgxuB48sU57dJCBTs0ONxN3LSEz9FrMeD4LRZXeM1dwSD9GjCKxQJ9ihZPpcXeMHNkOyRg
ojub0c6/WjnVxTcaRCKuxqh//ChLMj4clXOdLzSoobLAlyG9oHuRzsE1T2OYidD96nK/TRd+8QpM
ct0BqnCAKReMrq+hqC/OGKLfEmMPF+FrqysLSJL9OjIXduuPE5o2RGBX8GgDFBZ2eVZk/HT1rAyk
Sbzjd/6DZJ9JSSwPcmUQt+BenlDT1gRuOmA0eGQ5mn4OXqkag5g7p7XUmtEYwMcoT3lDwk7yEJTo
lnErWFpMRpJGedlh/tGcBwoF0wxfJJhVy0PLaU3dpO+uw+kQMcJisoj3SlmHda0UTukFrgUh5RcH
Y4vzqlrkETrf8VOBfIATE5LXgzXRHsNvesOKGgKZxKRZzk7wPzAtEpKF0KReQ+SDpZs4WhUZOPlz
5AsdAy+7lkeNN6zmou3lePsG76IqU+wZuFIYN2cx7hSqfcoa+iC2wiBOwkmK/j3D+HGJ8Go30ZRY
3MKoQqCkQTE4LURYj1i7mzs9m0hADTdeelnixzV7S7umueHSWIkm8wSiC+dqYJm0M6B6GOKWx9Pv
E/jiWVh3KrHvNyNVbASGgpOAAm5y3YFPmtWtliPEVkc3BK/2SeJ/MZVkjHsRENCS2rJYDHumwJ8g
1SCZUCo6iqfSEXAT2/cjqze5gjtMSq5taR8ZdA4+yHtJGgVOBUli9VgBhRFeDN5l5ckSXQAGxY1G
9oFDbtHEyHO8v5UWemtrR7iruyFGDZHwMUMN/18kMnAjNDqplLwuA5ie8yi+WXlSwIkrUdwLbsEv
g113jp9S32q+zAs0s2jWn9C9CJx6r+yfpmP6vQVPsMyDOWopJdPD0iCrDcjjnZoxTTF601KcZqAQ
0SVlVt+Jto4ObNxEK3d9wsZ/dEYbLoVp93q25C9Jj03zdgM9WxEeB7/o5Qgf0OskhevkMgVby7+M
c/+Xe9aAmOFWOVpAuS7kbW8n/SoqkyuZh0E7r049c96eTeBRytfP5xB5Zd93efqBosybwof94Zrk
0xweAjZvVPTvnXZFTXIhT9QyzWuCArnznGSFBWWEuiKN41Cn9MrsdkquEfecCdC7q8AwBSQeKQjF
kZd5CQWp6zR3pSwa6Tp1Sm5vRE3sSl9uKoVtK6dXsXM1U/sIAVNJzuvWNaREKyhRKkU0aGzdTxLs
ddR0oY7GaLiJVUHjpHkA/HFLCfam9x+d776p3g3x2vpGlI72T7z/9j8B1wuQnUIcK0GdXwZHqzT5
UQdorycUTc0ihuPAG4UTSjJeGJ8ZM4CeCTpQ7ikhBCrB2ofhnB3gXcdkuF7QDsc/YiNYHHaBuxpA
gVD0c70w9S+FJQQMXkTAPjK6g9wwlUSShKITqiWx7/V31P0YPTFo+sLit0mNEqN11rcXrJTUG56Q
NKhyLQ+Xf8wCXq1X7x43/iFIJPdMRXbyb0RZnV9qz2iOPCFkKSc5h3e9RFyzeZ+3nw4C6zJGAsSz
in+dZfdN7hdce7MKTeSPQKO2+KMCjsSssB1U3rVCF0zlWaoXvRRgAM7zIaOFOa5mW/IYYt6+Sgnz
z4i1o6zxlUFgC8Kt8Q+irqMw7O9OoEfzHtpJYifp/s4zOuyAi5OxM1JvZ88eCHsUaU9zvjqtInEL
pzVtvuMfY3XC8LJ40io/uQxLDHfLijKBmthDXxiWxmzz+IsuY3IeSGaVUh4vkZJOnlLMAZEOJRHH
dRqBbHAvjfoY7iVvlVjjvV2GUmWf5Ty4vLeNUHXAV5Ov9Du6tT2WvLKNsSc/5Tr+UVKpeL8dcobc
cw0miIJLKUg1FSlTDMVGzcy510WmSrhmI0bnjlfxgtKi1pybbopsOaMF79XUwvIThBl9/POeOiG9
idNNWSb3SfkQscRbE9lF0xUBLUqhXBr4tYtSfcJ04CdXyD4i3qdQhHKzFLLKfCva4EVBE77N4B8s
tME2OjlxKkf+OX7PII9JrpszjsNPaDB43nor1kdMZ0MoGF0d4TW7toEHqeGvL0XghmKXG8ar7yN+
gSZCRp6MjOjLRnqGZhih2m9BHfHVYG15hgui/xkyxwAaWSPesZ+4NvcQA9gN97QfmkRKs6wMGFhA
Pvlht7LwmyiQ4zxsaHuafCxpm7tQgLFk3Vl52/Ngtl5+msPJLAdvp/dahof9IlE4NjKDNmrJYE3T
VYav9V9ggsKvxP0jNPgZAmn1GTts/meVxDQcYWHMgk1x+SEqdxPqra6tgllIUvHTa/X8pMwYyyHG
d/qJHJuMNqNLfw3c98MEpshVX7gcJ3PCPUhp4OOaFYSwpvtqBBwe+Sy8/gOradhPH2uugxP+ouet
SSX0h2YfDNoAMWVIO4DYx+URCKVQP7Qcxj+j3JLrji+NuTcdPWMn3VFQMHa148JKAwhftkMi32Jk
VXIWT/S/fVtE2b+SPXP4Uc/qdc8Z7u/sX4nUKot5Ss2vLOsYlPuU+ZaLCkWP1EKF34MXSdozKJZE
luhIZQcvIzoB2cQjIzA+4oyCbARtRzjrnWcRi9t5nW8jH8a8ywzYSOaSfUmTOSOaDWmwNRdcBF51
aesi9CzS0cmV3JZeeUJUuhR2EI+fKSxveUD8XbWIVJ9z81RNB0KnrAsg/NnEeLs09SArMzPUpiKp
3p5vA73FAF8v0fzPGTwT/F/WwL37kdi69dvxeV5ZUCf3y2x5gVhJ5SXlFtFPMaZzxzbPeTDUmxCB
15NblHQnfqZ4lTL8EIywGA6znISiwzK0x7gt3owdMiMRUmC1X8x+T2H/CInH7JJir+tqSVVwwiTz
zTsY8ULuDaWq1yopwGegLai8dEcAjtHomK91qlPdUdCUjf9Y+2r+P9AkyLDSiScKH8GtdiqnUVIJ
ZRD0L133cmBPN3zewmVBgJFYZjVXJH62EQwj/pkR1K3sTTY4nEs73swHyA8j8hLmkzEdJF6k7/MW
X63pKosLXxWZpvgzdzrbKSqrD9iE09l/miTr/4d9cD31bkzmVN0PvMEbm2t6jbAhLcEhG3qXnPvQ
mI2D8uOEfxEIS7mqdYC9MvVhHgYGchknEDxwrhELbiIozDpTBe3RfQ4+jP5XFVWyvECEgTaMFBUa
AdQ2xkLKGlUYx9vTkA0FmNxIETXk1ramMNN9bhnWncMHlZKsRw2i7Bqo2P+GtCvf0s0Y83b4sKwp
T/qngMxTRS1pqNRQ2YxfAt9lNfwJxbzszHyqX2U0mG2hZiqub8lBX3Stmz9NuGQDdvNrYyRk4e+Z
mKD7fn0a+01kEr6IK2fNeC+JIK+15gwc+3gVN1ZBSvcpu9Bdxd3ZfaWfYJkBshLMTkoqx3MUYMKF
UU/OnK3ENXFQdP4Sj7XrHiiBt4S7f/yMRApvEsHR4F82zHVAuGYZwjJ+NrqgvmMlfLk5SOtWcj7M
SD4NwFfJhYQC7Rv7jPwvagdj1sHWzyffQDcQ9uDI+zifppuu9koFwGJFbZIovvK4V0srH16jlgCY
AJ4OWm3fLPfqIIZTbgpn54EPkPjzZHIh6KGJAhT3sOWPkNu/OpZ63lzXd4gUtSaSWaAOoDKpMTIO
U7gTxho/7QI6LhFNCSQrycrQ69ilGCqvD/pAATg4E+eljmvA6jUANV1FmHb+qTLhBRMRr+L0kVpX
Qe79Og0KLQ6TEwquR2XRJxGeXrHnDBTMrw5j5osiMxafGM55ZwD+/O9n/5J9VgsVsQmLrR1YtDSH
cf1f8AWMCy7iAOzuxFHC926k7UmmA0nIwGiUqsctWPvyUNCojVH4Dge7afzgPMi2E4yfZHoDKtlv
YDm3Jz+5GWnor7RcQeZtHt8QBo9s6uKswCdswSnLGRPQGwq8O3f3g+CSNUY+u7W8/VdV7hE5bVp8
UyA5ZvCE+jIAa3+W23tHl3vLAh1BYBID/6lG5JbPbk1h0XFPDJ2BqIlXKgOFgF/JtRq0rLPx8FbI
Mybhxa40z2eeHhDd4nmg0M3CMWWa4nQ4ww9UEXwWgmiig2Bj+UgOKsgcjreHtnQRndCof/H/4U4j
JFQcQoAquyCaRqa8MPP2xxzDeg0oZP6KZJXoVJUUyJe+tbpLe4Q38TYuGVsma0QkvyMNiWW47U6d
7gBKV+fBD3F28lKuq3xmDEkiYXjfpRf71mjpLIhW0hJPyoGYx2kll1rXlVQ7JPbFwjo19XPUlTeD
dwjm1/FsegcQrE+HAK2zO4r7OFBFlo7t6n9bD8o01WegOPUKfT8dl8o1Ab/4QZ11YKVTIK08cC9g
a8GrWlHYOLhESw7upsoNfCTsbKSEvTL7I2tCacLlPiOHTMXxlsQpTxwRrIXaQMv5+h0MDnjQC68k
49CWvKm2dKwxu4/ebPoZoGAjwrdxhp9nm+NjM9ieX+fswl9x9W5CcOo72krJZtUm0yFE5FDswvGg
t+Z4pGpNLilpbKLqhqkQgliiUIEjg6dX2JRTTDNQ8D8QB6C8r067W4/0pSBs31caizRXmT/hk9h8
pXPCIvh5fad5WYN9SiFtKv74w6wQJTrd0OegP7AuUsnm/zC5WAf4ad9vB14TlAvwUcrlppyVaviW
/4EZGbyRqiReG3BWVMhDQjSd+Xs7PqYyNOjND6+sc6PSlYmmDT1KDEt30aBapEbxHLdv02bt0w4c
CyQEl3BH1JyA4TqPUc9O97qlSKDzkQumQLF3sHhtFgJFRYWF3jzoVo5SC71iRxMFy2HFyXvkWxc/
8pXXnqeHPPLq0kSCjQIZES0ljVWCbh30/AKYgFWjyH34X46EE+J0GKDoQZX3E6GKr0rjdFIWoK3O
KN7vPuE488fPI2Qf9/6uMohxZe1c45vWnMqHy+ZU3qVhdYcfD1xJTdYJtwlr5WUhDozFbOCsreBa
hM/OeJBW0avyE4BkhL1UMe9t/4/4OeS7p7LFFaWvc+SfOYg3Mk+GCjcoUxhyO+1kXiJ7tx52TOhD
WSa5fVALKK9JJaAS0Z+5P3bsfCmY/nGQvfpZP7dAWmZbuGqrlbZWFVjn1yYpiUHLwo0qGc7sFXib
FQcSvAWumOltFgP0/6UaZJ86hQ8d3GkW4cN3U41nStMmB5abX0ntDu5k9Cn6nrQdGHkvWmJkOBTY
dJMIFNd8/2ZB8zdsDI+tLAQGdq8divTDu44kJDy7zFexqgsu8ifaZ0Fsbg10ACDLlHgzx40/wSHA
MYsGV9FeYpSv+2cFfTs5Ro5ZlGW3oBobJrkb0/kXgLMy8ZBTGfCHr1ZbeKPtWJL592bmR5LSEQYc
SGyTe6cUrJ8YV7M1tjaxtmvAq8PYXsmir+ciJbwD6A8BEN9kzqq2V5mxpOsS510Z/wVouMZfY+3p
DwAlObu/UcUJ9k0/S4d6gINb6OTYMYWutu4oBglhL2RmB9RVbARRdBzttmN1BFWaCghJTAnGnf6C
TY4TVizOLWJXVJM7ur6Q2W3cLgcBxwH1QCKK7rJsL/+f34ERUx3b3Mwcb89skt+C++cZ9IVBSNJ/
cwAZ16OjnoO9GAelIx6rjUdyPNRbFc5B1Hne5mrNQoTCbTklYSjptHSd+Wnd/ZXUMkMjcBr7ctYF
6xPfgWKSGxDkXtSwxdcTCaYCwzhxHUY5vZgwslmQnARm2tMWUrrU0+cUewDVBHc6anmEVvKLLjrq
uijGj+ItHKlmwZYbrG7DGbwBKVIOoenfzO0rRzkwpX7VL70ymgzjMPvOH2p3E3I15KSKn+2pBFRy
ofa5YdTJG8hmT7mFeE5HcyGYdxvcTcYkhBSO6JFGrG3K3K0rdxiDpZDHi20sDBy3qpuqxMkERIbY
EvKYnX3Vrk1QVS7bMfPXt75DlUz3w8ACaoR8gs5PFMeSpMe+n0RAwkme9etd7ljttr0EvH7fKzmu
4Y158Qmh5asLYTJxLEQR7jldFKbf5HXxcDtoYWa4bK3+CTFFVO1t29mKrdJFYTYyeJAsH9dcJNCw
aeSpC8T7AEy0U1DB+z/qborBmHSobyJXjP1/wQUyt59jrHHYcnRZc3SnyUIaKvwJ/dLtdPotgRSZ
lqxE3y2iYEiG9yDKJtgh8erMOV3Woq/8X9hDg2ccQs+ZEC+YFC5B5K3VNuLTL25lAC2Nz7l+selW
/nFO/yEmdty1cpqVtmwdiwy5VJFEw3EGxQxGGM1VFvo/D4RLUy22hXkx04Ck7+gSqO0WNt9cB5B1
GDYLYPXNAQhN0OBTyuTPqqAUNc/74OMYsiT4MXn+/F5guTFEkkekrXdASahaK7cnvNzphEoSDOgJ
2+B/XRDlbXgUNmkZahRyke0WTTsovXUM/cyGh26uIoHFDIQyxlFh+Ww5pbfJqAIL4oICdTc+8GoT
FHLReSnkaGeHoilt17c7zH1mRzci6Yiliokqz1f0IXhY2qGG1snmUrc5DwJC9TBYQ53Lm/2eTfQz
+8dawTz8lPYygNXJ0St4I8/71/PsAxFJtOhBLML1WsN5tGrrVykafuFkF4wHc56Tp5TMTdUY0UTF
rmhQTKvfbmvKiIv+Uk2VOvu6jHE97gWeAkFOQUVZ13VlwnEYFlUK4gFarsTvXf936r9mKc7dnctR
E88oBBySNto5AKox81R+qiajJQfN39QBgu+B/rft68m5nCQZXP/PM0z22P2RBzuo0FdyQLuQDPz7
XisdZReL5rLDordOlKQpgyzKZBbU80+rFz6unKM0BPWxo1Ey+Dt1KcoJtl3ygXJF4GvpjuVjfav0
V67vAd49ZnYWFtib6pWQ1GZfY0icNh+Cdyu5W2x+O4Dfc2PP3m9nrlHbv+woOUjXz+KXFTYYHDao
2+7SxZvOC/R1zHZC/D6xnh34ejJb8m5VUnz5lP3wgPa9rycsNSQtFZmjHE/ZH8FRhr0ekhlcTVGn
k/lTDoeiUnbMA7rY4o88M30SGgGBKnAUoO6X/U49m/eCk4+Hv83CsDr07TfPeVc6oQEvozDxAnKg
4b051u0D/2wHAXeW/v4swsInmCkwlEXgecqEnnfviA+ypzbUjaqeO38G0P7OZbDxY1hcE7Zq/SeJ
X7hpZZxAc6Hr3u9hdqDHCLZTkMGGeUA98/6lrvv1rYp4N600VRZy4PwH+26ONy1Nvm8Y5ArXQTCc
c6D9ilyM+OyJcI5SBHULP3dy64xobI/Fw+N4fj0DJ4uJIXfb6oNp2vUE8yfcDtA1xM5dyG5Etp4U
Yt+ADORDh1IuhunVMT7n61xhkiUHfNr3ldzyGZGVbS2jf8+dk283FwUX3PVsG0S8x9jkFIv1VzLU
U+ioD+l6PiYi563q195Cu72jO5vnl+f0xXh8viVqmSZYU+9+HhX5I4WkoGmRe4Frp76q+1Ns1R6o
XKkuzb8tbQUbFdkq7LPt+Jg9psY8d8zvK029+LpF+vdB5zD6roNXX6IDu5UwcCzyMJXRG9LlKl7C
gt+TCKPgIz4MVkumVhWlOJHI9g4sMTrl/nd2ef5/TMWbB7ZAk6OHwQ9cSpULyqX3NWOzIcZhT76w
jv2Jjer3phL9PdFix15jibOrA+DiU32dHdoOIRT5wMpVp8iO55pYkGEwtf8MVnBtQK4cuEDSweHR
Ani/KmaVKtGuVqyEG9Ox8xVZUysUVrijLxEBTAVUGuMo2JOepN19bH6mj9rcpYtpZeMSXg92wqNN
nfg4efN9MV8FlwxzNqusJV7MJRkTgklLB0tAfL5web0RngeghkwvWorVezXXRSGvEzGQwHmlZ0aH
mBjxs3DAmctCZrc9/eO2Os7Gp15OqNAsjeRr59SlpExCCw8wzvB2G5VALHoBNndta7S1d4Lpnzub
Jm2qp+/Qr24uDOxuME3uqmYuo5ZRgB6ORqptYssAvYJmAinzUjjSLSyVzjmwgY0Vv9k5ZWTRy708
pJdXyfliufcLkzExvDs5nLfgBt38tOF1aGQzbzp1z5lO8LXKV126b2hTucb5hsqSnF5bdNhqPsK3
6rYOpefOzRqYHuZ0os8HFobNe2kg25rT0XqICdsKzTPX4vHMIUO0SRhOzVu08SH1Ncb2z9JmtqlN
2iDOd9Wwo+CTJ2ZrPhRmXGK8I/2+XGWLSvijwTdy4Csq9JuKcLzSqUgRvGtkILbmLy8XWhiQdpII
v3hRFP6gx+DpaCVU/DwbDsRMepoE5VgwMpKW2HUAEC7MsTIDosz7D+dPK+SfOy0bitlCsf56a7fL
QhUSow/bMfFEqBoCexajygDVzOCSijm705wLJbXndC7CT1ybblsYv0O0kbZoADc5DfVX6N40e1EI
/CjxWV62b2GrN6eNpPbPjgfWjOQDwYsfBMjSfAFHx8rOLDCnAHGGwpkMJVKCotsexeZdsxOgZT+p
F8HoAIPKcwAb11Lz/UOF5qFGvS+hGlzmVYYeVgmxX4pncj/RJB4eYty94w7uZlndTuqA4XBpuFcR
3qG7Adv10t7m7Gzsp9sXyM+2p8nc0yEeEKq01CVJt0s4N2MbKSxD/0U5jv/xCvlKV8i90+ZBvelS
DqO4GC+PNUx8y8jEFzUDXHIz03ECs3zgDxH1UoMBeLnRKSnUxmVRAWgCEhO0Ac+dmR3zre/v1tg8
7qGFRiCFcrwgKCnourFKMrqIBxMGFRJBrG7r50FoI5jcwI49R1qk/6m99hJJrQ51OMdmL0Zv3vzm
Mfhg/WOWsUqCATTz8DZUDL3wUdeUpDlW758Ypc+5lr00icp/bv/YLqJnCiPoJ7KYs1u13QPMzX9w
1Dmj+U5+IoZSz9wVAxcjXrHqZaks0YMnHiD4Z05cHpQJLbBAyguC9NU3XpX+r6RbTX/4HuMPPg2I
n2wApJEu+5CmBdFrjgvxgXsTuS7QAVWdEyseFEIfQ+frVtuRdRh39AoivfdK2VCIvrwTfGqEV54U
GvfsY/8kYJvlSvA7fQjuTpGgDzhjQcbKm/VGQneL+QQVTbbHrNVO9mwiC5fFJEEyt6sBQ9HHJO6q
Mcw6JvNOu6UZ+Tbg7/LGeR70GzD4G7xJOWfJUNUXtYT0/wD6v0Fhr7OjiZV1kP6jn9IDNgfz7gXm
aAJg2NrzE1qQz4k6uLzZgMDWw6qYH1+QIIVtR16tuK+9jwmTyQQp4LtDl+3Ok9+BeV0EZJZeLE4e
3g0SJ3DRDuPHnzqBklcwbQ+A22uFOH0t973b4LOzoVy4i82ZHgcJjkQsYGBFEmMHzQ7IB9EsAExL
IcbyCxZUVKuuF79hHzLKE0cMeKY6YXp4u06OakeRZQ2/5gidJaLa1fo9vR1IuMuzvpdaVcm8W2NI
ybYraDhyd+Wg9q12SVkBT6dSeQCI1tMUINmQqDMnbafjFeaw+Ux6bPRNKf/P5CGlFYmyvvdRWnfe
d04Sq+hpB9ysjmkvofWQwoNJ10fTwMVe7QvBIV4lD6J0BQLweLZGctauPArtOJwP3NN+TGPHRDvH
KDZwi0RvqJo7BjUS3NmvX4fQkLdLZ7gyDJvEk4cur1CNyKqlLn6rligC8qZs0yW52KGMQXIRM4N8
T442Y4MwJYa+T3wJpi1Q+aDw0SsarBnutFcj3bvHTS8aETkLgQVf0fw1WoOlfNiqyAeYkOEIjQA0
aJTVqjMxr6NhU1VZ0fDchCCeSfU0F4NOJyhYx+N/OdNpwqtkgz7zEBvl+Dnx2lLL4GMS8S3bDYZV
r1lYjk1/xt8AOx7mHlX6X0V1lUUfDAEu3DG81qBRn0vxdAG9WoersHREygd7GoCkdSNRwt7s/MBj
YsGGjYHKwIK9+DwmBdQfHl+X1/I9ey7KqKWeN+IKeCBgFE2JKy6j4YjUVBr+uQUdu6+8NHplvtWE
m7XDBbweq20GOIIcHZ2mGbLwIJKi1zucp/QWzA11VT2vEwAFh5G11eGB0Oc1hJDzpJes6SDR7gnT
VnR5tA+HzQk9QqmSMAA13GYYyjc20muXsoundJPmpPjQ5LIT8CPx+WPSI67bfAl5mhnWOXF2SYaC
OdjiZoLDU/ZuY5LuUpF2YOj+X25sqP9Kp1thWlkA4K4wbtRM6rFeEPyQ258if+Xh4y/uKQOQPqEI
aA49HeCczVCYtkdhsZvlbrbBMjQTN5O5VVU6jO7BmSyWovM12tul9/AqgmBfGClbX4U0F6OQ8xyA
B+gL1I6Rli12tnMP+mJ8vcuEFN9XU1gt6muALy0wGgjcn9MUTVYzJ8l1eGNQCjnQ2qrAC7Z2I1Ri
3J31gZqqxgOmamDJmv6+26tOwhVpNeJEPeIp8SHVQGt44s+TfdWuv++v1q/Iod2UNkbWUe0cZHyp
c1A5YpbbqgU4RnUhOjlIvQcXT/0VkNXUZU9GVveIwj1O0Kvp5NLAsPfqproLPq3rG6RvHm8G/cuL
dDMxoQ4j6zT7j9dqxj0YTMGI/AgfsOmlX2loHQYyLdc1FQqlDU1n2wr3hSFy9xsDkYbByOM4fQ8y
TvWdghcbIs2cQ02vArgP9x9N/679/22HSEKByAbuBiss8DcgKedebg1Dt2GMFkM56DeSWQ79idX1
D+u9YjlJGOkuwz4ShR321+T6B3aMKHAe9+ACg1Y01R/b6a05oOV+9qQnoFWz0y/7Lw1NPiBwKGWw
ag3o20oD5J0dM3rRHhFHLqkzmVTOG62tQvOkChBRkh2jh172uWWjteDRS6rjkhsM3jvec9FHZ8ee
ON3OOaocmMpP2SDv++T6O8d3ZJRDwnJZvjKnrkwC0cKqcr1MXfo2/BlW5MGHhT6SxfdJFLSmq1Ti
XLg5NR/6j+yVl8dBxkIXks0tDVNiAjHDUsx+POiwrB72MZg8yiJvaB/FPl65Y0qPeVAxs3mMW5Jc
bp40vSvJSzxQ/VV4tF2Ku1/1TB9KyFlk2jxt0c0rophl19D1AQxJqea0b90tGeX0twLtKxDz5Gb9
nNcM4yRHD964jO11qhLEkPG7bDnDSaVYIaSICKJF5H/CTjiwUgvZp0bv5wZvdB5+3JQej6te23KV
OSWd2/+5ulOMelk1+7uODt4C3Pc2XNc4EI/7vohOZ6PJkKxr1zUuNzBS2iuarQFlwCBT6uGtNj5u
LRznBmNxCKRfwYQoVpJP0PDkXgJUH8CSaWtyThkhpHlggK+dg9AvR6LC0j561Gii4oIuVW23uw8S
BXIRhhYzcabYOHxo+ckajxgvRYFA1owkWFDGluC5/OGXzg0yFmoWN0vIUeUw8CEtelv3DjBW39Eh
v4Smp76iWBmcfs2qkW1JoromvENNeOG/DGTtFx3YKHtzb2bBPQ2qupAHuZb8spH+ffkpq10dYjw9
fV0fF87IgyuaSGV7TFK15v69Ckcgd+1z167aQ1cpky/13OY1vCvaiz9P1Lt8R294g+IDYa4RT6Xh
K/9aULaohm/gKcIb+lVMVrhlLHrLF3NoxcokuzQrRdZknyOHA4iJqI7ujv5FPOgiith6tn5friZa
Lb2LecKxWeSJE5qt6flEPumICudjSKv50cc0OROTCQCuzhI/m/zFNLdxsRM08qyZnkxbY9iUikr5
GPeDuwJoFlW48OSV03bLCZf/v0nO9Lc8WoNbejhOzZevjuUe8sZaZ1im4EtRzY0AGYb8dNvZl8OQ
wKIHojP3pEJsnnnV3uCB5qhCJD/wT0NkhqcwjKACacvUX4hWm/I4U9RBow8qnpkXKCG1dD1ulu8x
Cw1AMiIl8rCugGlSylin/zq5C3ahdcoN1TpEttUaYUw73xQTZyO7gamZyqCPh3fd0CHnEvWSHJqS
PPmg1HMolLq0i+CGzVp+o0HEOxHuHodycGQsT61ua0hTUue9YO/wsrG0nt+YRkrOHlI1oMAuh9za
YB4KzAX18s9a00hDiTs4haD5PqUAM0RMOl9Gd82ZlF+uqv2i+Z+huNmtWDICF8FjDx//x/fVk6+t
7jK+SZqlmiBgMEqy1O1tcUfkNiLfSK3/XQT9vFO6G6/YgiSd652nvBtlixIqHRUq1AKeik9RALW1
VOBYaEA6sTblvuPL+PndKevA+hQjWFeqhucpsydo51VJzP1fOOsvpkKKX/kSOjcfIz0PWE2rqgjI
9tbpev5K6jyFPHXQyH88P+BRPaQd9tUFEQ/7H63oVIaXJ2Of7Xml7gPMAgUeaqRekKKamGfSBPR6
d9+8jB0MWdun6GLm+8sFh+Af1Dw+VR3eXnd8YuegNbHK167uVQFqt294kFUfIxuwE5VLfGcNMli4
57LXxC/LcKxUrdKLSqmOR3pyiQC0f+O6zVSdEtdCgi2UxFp5zF5HNouSY1RSKP9za3NXvejfBbbb
2DiztvYWGYbIddPSUu+tlgibBaS9wMoJBZakQHYEugnZzl1ibKcmZC4bQCdnF6UryYiwysayTmVv
EUYFL2r3DXV8H411BKKREl16nwrBP/Xf1OiAnnQ3Es+vSTBhoadg83um81O8dOlEDtZjMLLmj2mW
Q8yPnxpwpbN9SOGDOEf160Aeqy4yl7QfZhyaDEiuUx06qeXfe6GhwU7oe4jqtNu2u12a+OCSiCSs
HoAVbUMre3HKm2TnPIMmWJIugkrKqb3jXywvj+wyDUXXv6G1Ll54m0i/QQ5rcN68xewfyWiGkH95
SHPSwdlbXXgrIoOHY7297e0cIQVFk2Huuws2UgFb7O+2i8gTBF5YDu3MaiiR91rklgQahCnYIk9U
9bKm/jhCl5StSq/vUvPwr6nU0ZGI7C40LzX/ZZb9ECDzQue3f4tGYc3wUzP4Pz1KhOvgl/+SgmFw
ziJu++pCXVh4hQAxZjkaZ7sHxfJNxX8/5PCC1RLa9LVSOyL/5264vFTB+JGtN5B1js1uJM6tdFpW
JcZ2eDfWZ93+aQ0QF36j17Q37nCMLffGcQTwIb/Krf63MSor3vSXIsMMH4nO09KUhs0M+VlNsOJS
Tq5bPLfQopWOCF7SscwKKjtgfKEHrtMUAFxruGU6y+spkbVmPFyqLjY+qfMOKLZ11v39Go4Ycmb8
xfEZwbSih6MYyP7IUTebmbm1CAHTrUO/4tJYPRrFe+Yr36DrzoOQF5D6GYbJvT8fWdsE+YLo9uCQ
kxzHzehkly6zDHux/MhRMdsZYNscHoYf4Q0Bx3Pz2V0E34bAZITnK4reay6bRYE0lRcn9TGPU4uF
aUpAoraN7tGsx5AhXh5ATJe7wQjTNrotkylxwRqtX6st49lHicl/OTWVO35mJ+dfxO8oJb7K/QoB
0PIrDcPMjxX5r8esKuBxio3nWl5Akq7OL3FbLdqm6ljFwg0MNUKWNwxN4qWdD/IxfTZuiqeolXJ0
AnKZti5gA1lvreewMEiJSKPXmgXQMPTUH6LV2IOqy75zg8TPWHnd5SRO/mOafLNGEFJ++O4x+wUA
4sL+/1xjnEFBZhuJ5u7uYxGBFL+Zm5E0wMgPfpLAf0ao//WbYoWS4pzvgdDii3bcDAYL+7VpCO7U
RrzcZqY57/ahgf7iFknGCgB7cQnmVflMbKQ36s8cxR2ilcYWPP4M5SfcJtsvfK8BvDIaT3Piw01E
FxVITL88ZYo8CnlIZx1ToQ89SQLvLLHJAbX84/Wxr0IiKu3dZFh4+vddRgKpwMwkSri4styX6d83
jnVFWwAcMMokM1ZMEYTUR3rM9l+GRuzelglg9BerSRy9eX6fXib1tCmkGHQmAVAcRSwkh8HmpTG9
N9M9Uv8Vv5vO9pLvJaoj6iY2ikhqIPCeZ0VsVQVIuvbmL2S0t1Qdu5ib3YgJ2uw790PZduMgqT+U
waLiAKsFx6HfCSIqoRzLjBp+bIyvysxBcewjPjz+/cyIz9vQDBLt6nlpp2UiyB+fbAGZ6t5mg6A2
XfFde0Q0BMfW+sZHdhERO5aEM0IfNPJYuPIzjKStp9TR+1TPScQKDYDtjbvYZKvXTnQhgCuSDMHR
zKxfsX6KD5wHXQu2HboF71me7J1OFTfl4ACJy1p/nbkJc73NTKeVpNcDNKXMyR6UrcnN2w/mJ5QY
NN3ILZ1H0n0DkclZxtWbnCZyIU4Yo4B6USN3Zu3NxAebVLV2De+lGtBc4Ujn9KCDS4/2uimSC8Kg
6dOjpmkI7XG443WPdSWsBvuAreqVPKKrMyCRJn75aMFDP4Xymfo+UIczwj4EA29jJUJ+g4SEO+Ep
iHLZaDNRct0LCWvvGfkhCsPrrDToIxlR00iV7OV8e7H3PgIZHLxu9wz2STaHj6HWUTb+tU92tMwX
vP1CRuf60J/WWvYIXDNjDYENYiy5WkC8u/t+WGeoZyv5khrC3F3HSkZkyOvlbQ4AQ2VTnepJ1d8l
ehf0CtBoD86KfGw+vqlQ1EHSdp4cpBv1/YGYCB0JsI7AUzC60w6OG8SCjBaiW24P0G8TtJxTy5Ix
bUDMjXv28mdTBczIr9edCYoxkiI+imbB2vC2h2Ykp0EyciU5LTLiQNSELqCmoyYIHynQcQZZxG5E
sTDMaXD+XCsPsq1RQi9xlWz+XJSJs+OxNJ5j/RxeUKAnoEHUvvJuDNkeg2BWK4SnQBaaME2FgJAf
R3of0N3eQcXj577OPokz+QEMkIV2FWhj8+ONO54oXOtfWBrkGnQAmX8wXBb9hUHFXMdhtB8cRUsE
qT+O6Vd7KFUC1+Lfze98FA2u5Xm3k5O6aLLKsToMxlPzh1n0H2j00nepupGBbTJylXsLi+RcpqAI
L6JUaHAcSsAPb0cYifjIzRPA5anHlog15Lcj0J0MzASiX+/FHKd5enAaEl7/Lnu0eSKqZnkfNjju
Md0lgnKpYnL/sK32oMEm4yUI3yrgG+QANgwiHd2xEcqp/8I+4bXNU+ErCvrcNyOEmv6u8RW47cmD
5c3ReMhiU7r+x+R0GzS5GnXFp97QBBAfSvFyjpMJNy9Jrw+M1g+rhcySDRwTvh4vbJQdi6VHPd5A
BEnUuWXxTa1bCuD8WArjL29v+3J61nIxm/PPsj6NDTEDkhjZygKj6+TxCshGAEktGD2avvRu9Uw0
9gGS8axHVNQ4/DAqwWyhpuuNL7B+odMYGr5ywmSnlzgYAlOZf1ZEJtZbaTibGMAUff/FQT0edr5P
kpIX6iLv1qbZnf/y3ycHbwkX8RpDHeKBqQ233HQM1YHCHv4edOIHIl00m70t9ya72NTJP+dA+Mmx
K910PdLy6vzrANiW601O67ViX7erTDipPquWNnzZ7O2PweSUO6WcgzCioKl1esiLFosOpz6705Ri
7sdOVGPpHZBYTlQ9XzOz8j/ed7AlACdJPUbCBDoKoYUiH7iumFJj2S2rZcHVRquZEvjSP2HmrdBW
zZ5W5lTcXMMc7MBL6/TxbVwNhwN7ZAXpkcUG0jbiNhfrXsGrousDQB7ITRr2ZQa9E8Ky68h1yBsL
JlwSs1LlA+yi78X7LgVZ8NulvTVJeGXYLTzKMg3pmhQMLBLpF4PzEYrlHvDE/uxZgTSm/Z05x8Ka
C+TOxW52aK7Vs8yvsL1MP1xqAs9ieGF18850g9gym1dgDDH7gCEXGSG5M/tNnQrvgSJgh3vmzzdG
wd0IcQqW03mxabTEC9GrQcAe2AI+hmbsBHtdziWSf5XDlb9Qu/MUlNRfFfHL8xhx3a+Tbfzy9k69
TsKeB9D24o1bFCkw8TN/JXbFqAc3kAGUSNJkHMsrXfnssqaqjTQ0VDBs0msO7AalGR8GRCIlgaEW
DgcjyA0tI9xWP8P3oTOTiS8dAwx8ZOme9RTT36P5JXYf+D5QYY6e1Tf6uXfg0x06rzbQqAE4xXAV
LNiAnoTVDB39Gn6ejNCkjnjoa6LIHc9nx/HTbuFnki6nyAVu1oIenVemVQbSg+zQFJ0nb6YxzKpv
5t8UVW8vIUFW/0nrXi74R3hu/o39E5viTcizNL+cScidUVOsyqFeL3JbGeAtf0wdm0kd7ROazwWW
oss08uVHXPW5Jd2e4z/lJkTb3JB2REy3NfKs/iym43bQTJWMeudlbBwOEus2ogC2gt7dOTvcWwOd
xnkWDAx5tK6WcBQf7MimafYdlTM9i7aYfhci0JSe+FK8SJWgUIuKun3GdpV2zs7wPJOmtluimSpK
xCQrOoFt7bbmg/3mkv1Y96fLNVxSlTAtOQl0elwHCe21hbp31K/HoeEkwpRNmU4ff0uZBMSc8/vH
bxQMIliDcUu7CFfv8ehyzo8Ar9s/VHv7Luz05UtPWdVtFXbxpknOEn8sZ6fAlGAGY9a0Hwy66pPd
NPvkFmHQ3iBXOyvcfOl7btWZMS8oMHEBiH3AhdmNe5felu6ehjfvm6/0PZ5yZRu6e/xBwEB93FOz
BtCfw5h8fbHz/T312dvY0ksXLnCtWnLXTKsFHXhin0rh9+EZyR0HYPTWEuuqMvvYTtq4X21w1ewa
U3zyQlc0nYwLWSDxAaP2ZBQChDLof4Htb95cyYk7kLZzoky5QITZBslgtTDNN+cEiTx1Yj5dvEcE
O6g2SpvK826X5/+zHpH166moreet6FE3DneFlJvly2SbB8FkPbCEMOAnwZmkIsZ19FEJKAlyFHMa
9yrMYsi6NBBzNvYfmQzQuknwIvCn3gf4JxdCsyTAHk4JoqwCdG34ijIaAisTsrcHt6UgG9ZtjzbG
W7386LT2QVsVX7sSJzk04JMYBtV2Z5XZtsebMWJk/17pDQfs9EUAUHE+mO3JRRYg3N0S58gCXYQC
3+iElMCpG30L9JlDyX3dIN6XxgYh6N0bSED+sVlo9dFvP2bHJ5MA2q6Dj+9n2ur3cKIfhkAT592L
1Q+SzQEzl1jPopGP34PGOQCJPIoa4FRwQHPeWsvKSRdfqhTjUBg3VC8JXATrPcIvJKpwJaRtdrxL
haGRGvZKSPCO+X5Xo9xGdgFaLghmCxMS6z+iSXT208XOCra+2INS5Je0voZCcVFbYd57X2xEH02d
QIjAQLBUDOwwJJ9kP4chr8mRjISQJBXjDDNt+917GTTcO+7rU+CJWapBGrkjjVYfG6/j9Y2zfDtz
yUlnKE3JRu/NgmlQwN2SQylXGKvd6X5D5p5SBGgawh1Uw+ZYX2dCNWpeU428NYbr/lqTB3JtFM2N
9c/Shz6yS/0qS7cTgz6SQgjCmpHNugeuimBD+T6vzYLphiYwJmqRmQU063QWI4QnVRMLwK5Jd4Zo
gQqmNoGNAPy9klbAb561dR2vNXfYiWcfntuhMqiTrB/UZFH6XC+umUR8cDEnV9N1bD60F9NHiPXy
Puh4jSeJA0926kFRyPfOAj3iT8016FgpC/j0qK8shkXPUkqhh5u5WEF8qjKRQCUaz3CidXDf7k5I
3iU+D2j/WYP+rV7CYpYZ7H3eD1Gvs1JeQlUGiytkb3wnfoVDSFnjT4olnt0dpOX8wcEOMhzFHp6r
Gubx0jdsUIIGGvhUVv8m7+54C5nn/shDWNEImNh0wnigLUbNbG9kpPjVsUYP2luf91LgWNRw7Zrv
NOzIrlSNF4/XvwLUMNMKntviQ+BuJ4Qi3W64aaDSCYk2rq4SXNiNPVHSw0KIBKH64eDg2rJ17BMY
EYHTrAiSvkf3H9jucZti9U1KyrsdeJ1c2jeMmm1kS1RVxefGpHbhxos5FYcKC/Kfm7pYM7Qn1kjU
Yykz9JmYuRsBzCLrFCr11srHVHl/K27FJK+gJ+FlyXxEwdEESFgpp9z608pqE8uEqm3GeJhoqmqd
nTsNR2ltQJqnr9Ew9eyF3zYOlNhabgdrbhIm7oXWk0l2NtyQ89kYNEklJGMqqv3fQceKMRPwjn/r
QRnG8UjoNkzqAtXJn668L9VYYocRQWlRQF+Akshd8sem1mrOmAhuqpKp5XP//BvsRw+WTPjbYJI0
a3PX+BkMBxUzK752HklFOKcFgoj4WKuIn13IzOY2WIaxABwFsPTESg4pMfnuKhxzoz6M2Tg2HUGN
2zVKTWgY9ADInW49VYAYIh9eQkLoNy2NFtuLJBd9l+eMUR4Grvza4n99I3+w8B++vQ5kwK60vSnP
OEsKdTuFAryRd+4YXyqgabDiHjqnYmQ4Kq/o/WUYTcXzkXPLCIda964otVcHiyTDT/9aHU58zpJz
I+hiKdoU47ILL+azXwy5USuh6Do6Jdsam/grK768icP9G23Y6mtpxIBCarjv3MAQMogg8iTPLwHi
62pfxz5UH104JH9nsqSTVf70UiOoP33iCSBnhZTWrKZWjj2WWCAfMFl9IfUcIVsjTlYDDvzuzyyo
ry2y7QEmBZ7FMYJrqzbXtT5lim/JSKZiZcbyYdMoWTJBFinjT5VakqwffWdZTivn0wthiTlqs26P
9ynbximy4lx1F1nlIeNJxp8z5qkKw09RZrj5l+FiG7DsLPApfmV88IQbsrX2GF+CuTTRN1LpMbBG
Dbe3MTpv8iXWJ69Pj6S5FfsfkbqVB31/6xHUm7ANSrwhz67lrO5IkTCVywvn3qsR844/ZQnXPqqC
afEBIClUTmJ4UCrZZjN+4y6aLvhWyh2ig4rgBu+sguByCMFOUZ/MMDnR0kXBUdGL1qYous0LTk15
SHUHuqFS2iFGUKckdJyLeqk+lNI59aNEYXGMjF7F0lOof4AdDJSfgAlWf8z0iPuf9ENtTKsgZV5v
/QCb/BNADEO1I1YolPZpBWsHyyyp0s/bJOxedMUOmTAyux1Wys1q0Fh1mJSMFFPFXvHrDNq65tMF
J/zH0H2s8oSDPgbNr3CYgYzGAHAFNeqTcLJeJc+0ZP+YrpQViFWMGL0s2L3nf2cryTi7lRnQdOHk
Mc9ZSVDWZK21ejYu+8YpY/X/k+M6h2VqEloC7IbU8LKxl+vrNCRLvT6lnPEisQ4K0XGhwuvMK4II
Ef7PzOksEnhcNCEw3Y6T9RaLrgOb/TW/yRloDS5xqu0168CK3Xqfi7Lzw1z+ILphN69oVooCxR7D
Md0qgtJ8irF9DUqI3yohleRTQoBou8F/UOTyhgQdCNpk1eCMWWrgx3ASJNwX+cX6GIB0fQtPigPw
W9V5iKxqf23VN/Tc1G1iTgXVdxw1AHBcCjsH6G1KhV3jIfZ79emnTTuEarV8MzMeQk4+B0mX41cP
LIrKSyC12gkMKumFkj9H9cQZFqrMcbQsakdeveV0o4fy3RzdLGrs4zsX027lnJ1oUeF1tP+MUHDK
euGuOHbsH1/8XMQuQKw2WKZEuT4YeJ4POn2rwRa6qruFs2mZ2/ZgwPh2HO+Vms68MMlnHGs3ZxIp
ZG0nB3w+Eo3x8WEhLNBztSKcPu1b0K9Rzv1wMVnyfez9mrqGb/ZcoXas79cfopFjJQ4tz1Snka8i
29Rc2onGBN7I6cV1BNOOnULH97yuzwYJqkmKA++FSybZa9uBBSXfj9lgXVwTGP4di8ujOEm2QH98
KNELR03HO4lI/kAq8Lpj0IfCU7FDDtvTU4I3moisYNx3m1RAx9lX61V44L8AVHVLyRBBAS1mDuQd
kpleEQ3elUveREUdnClrbW4IIGIK3zTOmCc6bkZipdImO3qc3S0fa3Ay1L7GLHFaevgkqtFJ2BH2
1/NANyDcAmfYymOKpnpHPvs9lzjpUtgQjf0Soacc07LNKW+ZjN7oQeEQYmgtxGuMEdflrryAa1WP
PtuuI2cqZBRK4EAcqinJrQsnKrN2jzlvM6GfuGaZrFdQJo0BFPiof8Rd8mcpLX1SysXhYZED2oH/
1EXnjwQQnQzF2w9+N/w6D8D5oVjsD/Q3TMB+RiqIQnJs46Xm28RPj2jbeegSCTSHYBjkHMKIGB0S
paCi0wxvYyA75s5rv5wezTiGkOuyc73of3BLQEcH4w1G0/4ODMl7ezXM2g76mJESFOQKAo4gDSFu
8jgmeRSwCqFJpKiU5E2YG2He5m/2nlq9ordoNC04s4CHiZWQXvnIeL/dJ7D6FB6POcohaOZwZu5t
clHTdqf86OdmSgo/5xMVeW6Cysx6AJzo8CY5neab9rhnZSITaUDA+KrJpoXUsemTVqrXF7c8A9oE
8WUJH5uSxlghogCjwXucXexxItMjOxi8KjkE5O82RFf5Wv9pic6XhW9tEqwGRgzXrNZWfXknF0q3
YRgTgSrT1gwKLCNvkpI2aqMXROGEsKLp2p4L81etZA5NWet/Kl5jm96z5+7Y+UgrPPl4V6yBQWL9
myGTVf6Zj0BpOEw1xymLjKWrlJnxvo/Ms8L9jcnLQ8SxNgD4Z+aZBnAxYIVYaAwjDWaPXT8/F2MC
x+CMehMViREzpDPRQ+s/8dKM/4HuoRy4l6iyAQBnIs+X2/uOS59YGB1ViswSGQqxYwrv1vIm7/ys
RkMaI1/LbFiCoHWI7ucE9KkkK85/8aDpQFI2GkucuLBiUK7kIIhSJ0aokiXVLrt165W2V/ac1vX0
+KuAuHV+VqpG8hdnyl+M0fPwFIoH+GEIdAChpVqSzEuuY76L79kElkrd9jz787/o+/5AX9U5zgQ5
qapNkjRitcZdD8kgyiyu+p4sDR9PzYhKD9cjRsO9JWfrWmmSQEns0X6Hn1m7qGcbgP7r5eiwifp4
oZTrPB0ZSy6zoLUh3QqzX13CX5OZVR1iqWoExh78Br9IOOYgzzvpM9RX8hf28MsxTOiOh31fH4L2
kXeGfra0KmxHSo55ezLKmKNwyEFbVrDtgViaLcYzpMbwHPx137nUDWVntOQNZi4TC4poDstGCsAs
xrgn4Y1kP1BnK4sD1deJG6LRVp9VFV3MCRWSueHQTvgPzrDtrj088m6OTkycXRJ/U83SFrE5SpTI
OOk7r7L5ZSMlxZU7VMOHjt0xYISAuDi6FFve5rheo6bUWWv2NlSAuRiZHAZgCJK+JTCCeL9Xm3fH
pxsV1BAYfF5pBuFygMIUlpcwqpSMtmXBo4KCRApyjRHThjbWS3KpWkt47GXn5bgTgfjgZr56zY7G
Z4Sieaxw42z4kB5B0injOdJ6EtwpIOr4kSlTrOytCQA9DyjQLXord5NFYPC41a51+WiNVO5yf7R7
N2hzEIzXQ+jUelud4ccofN3bNoIA/TQlAcUWUurpvGPE0DX/QF6Wv8vNzRBrc2gFGYGWfV6N5KYT
mRitKp3uv8d+HLljfnbixB2dP2X499CDfCyunXyZ6DZVUbGJvml4ghbqxkoJvxS45lnec+7tk9eF
wPhlZJkJN/5vb4c/vCndO4D6+Dbnic9KTcDplc86OAaGiDP7uULsMB1vvRs2/B4lr9rsUvz+PCiK
2bMSTi+gXiRSSPvHMpMC7nbTzDz3KUxUOJjrOM6rRDayQOrmXVZv/LCeyRmLeluRloEvJSN19Hm8
Yc5aZNqaDyb2gp8GQYUbmjIFypW1iL6EuS9AelHTAq7K7Szk4sTppOcKH1E5hynzuqhcjVya86ay
LDp8iMgrEkd8vpvs+ebKDdgdCR+1pcndOSNJzIQMAHNyESKqXc9ZE9A2F3+MjekMyRMYb4hE/Zxk
XVou180UHGO8r2xw+wPc0xC+fAQcqoGphrk4sFa+VKwJbylqqwKbr6pTVM3BVzQoxjhDvMgNjh4m
QP9HJMjM0jC03WCbPk348E3IJAO8S4LYR6pDsjWcfx1oly8wdTDW3h1G6OySa+9Q5GNcYR88fcP8
tBgt81VBClYIwsmSmiuDw+C1+hyBQAI67at9I1q7sCJhBd/Sfq1j8oi/WIDjjSnAKlSL9XzkoG1z
l7S49PPj4xmjR5Q+qPbifXLsCoEMjwzSBI/q3VIqdU4m1cGowt1baN2U+mrVydTy4HSkHzlI4fmO
JVwMrD+2FYUUSajZ3v7bur1g256FTAYcsVrkJhwn+QftEKB3Ynkwq2syP/yFw2z8xq22F6y4w9Xs
tDar7sfQp5JQ6TCXOmpBX0G/JugK0k+CemJ6VPMfCNX84vb0o1vRxuE+l/xIWAfV53XKPQ/vBVIw
lfqQlBlCFBvESS/zWSqEwWXQ4oGx74kzko4QkY2QtGSYI7N2Pz20/f9ouGzZYucp1c8egcuG89+2
OPD+STfJR4ZIDNHGX/rUrmpVxt72l/q9BAQb5+aDBAktK5CuoTOBrVdr3cPyINKL4JgTqRqNsmEf
VL8aCMZx1BtV50u607A9iN6DPHY4UlA+Fk324OLgtc7Y4aJhiy3w2cK30rX6+FS6oIpi3kX7uAhl
VXcmfNlZvUeZYevM7zKfQliaZC7bvH8+Dr7TtZNEnij7aOnDBn2xmoSw5EF+n/vPv6YPID0Z6EjN
H1uX49Fr2kN8Fk7yQ9tGOpZpDKAKrvAPq9Al7OPs72oqPnp2Bea7ny0i/6mguMDFh+VvStoM/PL4
Z47TcEb7cltdKeNc3i544IFjS2jdaZ0zLwNbqOMTXJSnnVIEU4wbrrZH0rWEJjRCzW180B3Pw4Wc
GqA71uVTBeOAyCkZBMyNBorChqkVe+4sUzPKuPVDj7b21rC0sEUX83Lm7FcNSSuizOab+ykzUREm
uB4LbVo9pDHuiKBNnUSalboVOYrps1IRisvNJpfWLCFBP9HuWWYDszn/BVsHbpOpBuioDmZ2fiGK
zzEC5gA85BfjPFjdH+4sZBafY/mU+JYdFgrz1htwsLaavEta74a5Ab/ozaiEF1BuAtSFU3RyskS7
PTu0jly69qHXEbX+MDUbAn5CcrL3+jSMCMYyzC5vkUv8M8W54tpc3e+C/VrX2W20d4iSoAFX8hx6
r7pDpjegS0CJu7LWKX5ool1NUs1Qo38s9G1CXcw7gVXP3tBK2ZCMEJDHbBGYTBAWBJBAHTe+xQzI
R20BeG5my/ux0LH/vAoPPS+gzDUEr3ic9H8kbxCIIDiJljMoYz+JDRPuiV8EtDi1ioDjE2zOHSDS
H1nfMCshQmqn7o17e9+a2ZJk7c+WiJhEnQxi1rjv9P6Jnp920dher2oikVBv0jpOfKoxk7rgz1GZ
e1kMkBLPFonNx0G+Hi8KKY3m07ZA9KqR+c/laUWOXgVpjdG8o1/hSdqSzb1LH4BLgoe+h+dSNneg
DjWeBatYXkwhEV0wHZH8hiZ+T2WcetdO1FvroZDH2ffWb2cIcUWGLjqH26Y2MuylfhZUYwvVMXf3
/6DVKqeo7QerKTQS2mARdgzjW3BywdkcArGZwxXqx7/s5HdI1AzVNUsAkj7CHdG5AaySt5FqI6Ea
xos2hOWKteeKSeocY+sNB6kUl2KlSacX21Q0qDR4oacVHt7Se5X27U9cfxGDq7eFlPIKTWOb79ou
ixaD4wbPFxF6qo/Ht5z1tvONiD9Kxj/LYFGrhtW7mHwD3ut2GFeQzGUyRSTgIIsP92ddFjC04Pw4
sg9lgWrEMqagYUM4sLivyEnLSZu1A8geih0xmf44Ou2spn7FgO9LkJU494icNWO2cMK47TXWd5Co
3rDuySgLLk39kFPw9XGAiuzyWq02epPIm5QVzTt5VE/oAFlPyhiIP1dzr7jjJrPLXb9tbiSAa+O/
HbgoFFzaUR6+kNCdNbjnnL6AoG8G/eyFQiz1WRuOlmsFmz9tJH1xU+Xh3iJBhVSRHsUsXwFoOFF7
SUilRmAvG24nHyX6Oqkg/vE7uWyHFV/qLODUNBsbYFj5PlR1/AuoVWvacg5G+dF2mA/nvKtn8sb7
re9a4Rc4rZK5U4UPnGHlLvqx6iuiZLSsLe6eyDfBOuUimYnBECjuvq7IeJImSPeTA3lAsUTl2y0A
p1gtEeIqT0a+36PQPeu+jj8xdehtq1h3WZxVogk8+4N8rOKcR7Bl9H/oqbwzL1f9T6/pk+h0GAnP
Su7ZMs0je5wxllyMifFiT5euKpfo6ld8tbAg5z49FpjUaMN86Ykegn9XbF7oW3/pRrKW6qcc0EUm
ft3EbwLKD6aGVXz+yJ27UaOVFC7k0RRHMUPNTwbm7CRUZ7aIGIVH54S2bMe9+5/cW2KDRZ8o1tw0
wLavRXKlPl/4OrkdHg9pHDAHEW6E9CE4MyfEdmppxj7ejHQ/Xuu1awsXm+i1xCLLc2OGqqP3jpF9
171RrFVkyvUIkqcuT9Ph3A7irhUl9V4kMhZGc6WRLYr0rtE6daJvCRKjPLQNwOuZCJqW5KSvy+u8
0EnCaMzsjc/ePC6jE08CZry+IIINIVnbFmJjiwpcUJDex+ACjbLl3QCYeQZRWjR1curnsWpnmZ5r
6FRFf7kU+5ewkpBBY6B0egBSZaIu/F4fK7ljT74uWRTQSGSLRE+vA4pH+d2emvPcE5miiVU87aAb
9epRZPdu+unxCxd0NV/EUEg9V3avBIFqpgazH4H5r4FNKQI91gtwIMF6c9ZLo7vqBWDreFvqidmx
Qyep1EYta7vwzJoiD6U0X6hNmU5L/PiWNLNY5jSoEWqfzNpR3VTTQHuaxikTHm7yuN1TFhI1/5ZM
ho3+BZ6TqKPBPwZQZCsKOBiBIKLSW3uDQq1HbQWpf0KUqO6/V1M26fPr+Oyf1WmknEnz2MJMx0nf
V4EFpWD1MCWczxKlsGoauvNzzj2ox53URCW7/qWb9lMcjy//Kf6QDZrb3D9C4swxaRp2dmQKzCKM
dWmpCfat+nzYik22/rbDiHksJWvwoEWZl51D/1Sys2t7Riu9XWUoFH+djEXk5JtBatizdQOEyNO/
FHfoxQoFS1NAJHwmDRwDohMOjjV0UknDoC+C86MkjoJteruLK7Rsz+J1PNTIaRhS8GsWvkmfpTFd
xNBjL2QXiyubZIILKwgLOeefmhPIp0i8+O9iukQxlvgjU8bkgH+ZpBuiAoCU8yAmKXaleL1W32rA
M6eV+1xYlVUgpd5BtwdNEZKtVUvGgu5CywiMF11tAvK1lhJDVeMPTtgMgoUg6iwuoc1oMO7sUKMB
uFEmbfCpdtmntJzZJJ1IYFQsDvuvAO16I3AtQ5yRid4MYObq/007JcbZO5qIhQG67GsxIa0d9Xzu
R+txS3X3ZkzMqUVhEZ+63GdnokDxLcq63euqcWQNJe8sksJc9xF9P8NcgKOe2AplxkCZybiS+eeX
bBWCrZQJZOnEcmsaAmc0tpNyq6sgyqYOdEZ7agRHH4tvio7wCBPaLS+CjPcgUtl9VxF+yHX75Klg
8+azHPD9w290ONV+3l6meszFZsfljHPij8XsglsRvVqtjzWKV/sdGit6PwXU4dXA+DDYBLQzoWH9
hNLF1bkJauH4Yv63key+UiFyA5PY9OaVazbuuUgpfe0Q3OYla89ocNx+5McVbeKtfYoeIMq+r496
INz6cQgG393B+DCrfH+HO/a0nBxMNDy1BEjZTEBA9ofbxS32CWcitTDH5oGokYUMeNxy3Nf9BOLS
DE/B+gK2RM2VVFfV3PIyXn3iKsm8lNut0gxiPPA5zPSYkZDbXOARfc56b2/2O/3eQfS+0aw9sEBr
+VsKan1rKb2zuFp22WPeH0OjTGxG7sBTcNES9PtzUqfmnayEWWu/17eiq72z1K1OXk/wc0XWOA2t
iL6YH5PEn1rBLXKf8VzpZ/MVotJvjbG+AMK3l+cpKqJoAdrONIBUTuL7cscgJ9kfJRrFPO558UHR
aGpubCPJwpc1lRf6I/LaZS0Rwf0jtjK540xp/ZigLbNzHmfTtOoffy4qbR76N9WyreAuQIl2Ew9v
iWqBZH3wWAy2u/a5Qitlpwdl06nJ/MtPQy4mqlEwmTfSByOr+J3SLKnt1TD7w4qln2qVfVVltlZw
LzXzBpjDYAnMCgaATishrjhovtKIxHnKIaFnEPg3E0/muEz8YWckAFzirUSTMlHknJcenXxkIg6F
wS6DguM9J0jtatd+hBWijGbNn9+QCTYQU3T7VVnmWqeiVDO2mFR0b2CiVQdQ6YTL5LhfK0CSaW23
6BySe6XlIO01qC5e1aiS+oVsyC28wK4OigPVnjDJfq1JVGKLVN4fSMpNz/D5vdjq8c4W503AVS7t
3p+gQYVcY8kygrr3RM9UCfNB1kL38E0KTd7ZDM31/ecLzKjgxqBNVQbfz4OVeBcxFm/wctPlh3gC
HEH+YCN8kkErGOeNHECSNNysXCgzTPpdCMByK5huENyoNd387t1xM7cj2HKrdsgGYr/1b1O0fNot
U1ptim0bfJQO+B2kFb6vZIqxeb6Gmqt3ffMbUdWoZCxEwqcGctnXSGlR7NlEvuhe4EDk6V+zcoi7
ZfDqqwk9mZGsS1U3SydR5BTqXCMOPMiAD1TYmAlp2pVzMOBSF9Ht/bjj7kiuqU3NXmzfBSB2ST8p
apM9b55WiPg6ZMHrWSExZPS2IN+zRBTZMvM3/fHD28j198yO6m+sy6G9Gc3YmoPUwiB0CDBFjzOq
+tCM15+p9jWRc4u4wEiPohJrT4RUWjpKok6taPSBzBLTg0DfGYDPFAeTNGJq+hgIGvycu2s+N632
lil0Fs9NRY6jRM9uZKmlVVDtPR90aRulsevnvX/ze4sH6VUU6aLyV35iW5gHSXzE5jOikkz1w1ro
AhCVMioZRFT2nAe0ROZJ06DVtmyGOcJo7BzFj3PpIe67oZPqSrQOJ24mDiK7z/BzDMseOSTHtK0U
Da7bnFbM+PUW+xYAYBdXKzn8SGhgGl6O+l9mn74gx0JxvHTow5jfLF0ZKcxh/R/ar37iSagnskR5
+R5TUxTcm8nHKQ1l9NxsLusdv0+ZYYVln+tk6WnTV4fM3LoqpgpE5ENph4de0Im70Ng+ySXGKMFa
okbbAI/wAIWSB1wdSxWe3Aj/aq0FkB0zm1kfQqCOwofiI0YxVArhyFKyxpzSmk0LICBJcEpfnTwt
zrMsMJR/Kjs0X+nDwep5YZfQE3hSv0tg/b9oQf5CJTNdKqbiltSrY7TxQSf2aNrB5FI8ZnYOLo6o
cNuaz78QicZcPWbjeAY/7gb8WuKecAfskaULImS1KsEI3DMR+h3ZYFchNdSB96N8+/STivwtlfiw
/0lpkRIsAB3kPnlcWAs4drCBZLLB0xBmvw0GJgIVTIWFDwWadBbvBARQ8xWbCPgM6ccosBxzBu4l
yo2pg4SCj/oYb+9B2i9WPaQGMiR2UtLRBgB27x/b/Bt6VOA+uNMzu/o72izzrOI1K6Nk6TLVZ3Ad
KR3/6Nv93gbq6YXftIrOPGs+dV3T28BZsJZtVgkP9kfWhaJY/0Ih58+5WJVx+WdU4b1bgRu4Yt5D
I82RPhm8cH75fFf/+kKy5yOrjEbRWYl+3gjS7GqHlvTHusCl1c8JZqNunwkTrtyTs/e+D6UpUg/r
Ih4DS6ioftqPWiAOzOini+s6QyD+5FYJwcjavg/I7XwAnnhsO2ogrv7J/Ib88QKb9+tJWCB0Dao9
KQQ2kh56Cn2zuIS2llfNjdrH6C7KzwOyuISHZaqTtMinvs0gQY4TbksXGBm1j+DuVdLNww3k6pyj
7fXrZj4yqAAiuOLpF9INeWhIoGhITuuYhvz+K8CzFxZeqZ5lTppnHXjzVTh522G6KecPcE4tfg/D
rcEZXbY+H7JYp1jgqt6BXwqo0wlxN5LhUdU2+zexxU8sK7Y8Ffv8j9CMAH8QEmGXok+or6MgKodJ
zqCXuj0aTxHSnEASUG7vlk0YRPOrxzxbZv71Ftx5u9mueBHc4FDSVHOYOOo3m77gD4m4G/3sGRlE
8ov7RG8g6dDrN4IAfAmW9gn5qJtUaJb9swjnDH1Oqznpid1z61ElHKioE1XzVWLfC9JSVaJRab94
JLt+5ZJkFK9rComaIDKrA+voG8qD1/KfYzYPkqczjitT04O5SlR/EsC7nJkWz+yDsp+z+pms6xlY
U14sOz+nHkddbUbzBuoRUocxL1c9Pmi7cNCHzKKd+UJIJKhFlQXtBbZgicOJuWtAT57tceOoMCoi
aFh/De/nPDokTE+DTy90O+qmSDBxNCPIYLtKwRV4uWnhWrv9TYgJVJaQKTuUkmcSYf+kPbepWWjO
uLqgLRtD2nhomqYcvVi6Tqka2ynPwBScwz5xm48ybBKJXvZAegO+fytXJQGcNaJxWLo6jTktuTvL
i/tJkPVWQKkp2iZF3Qc0NOf+xJJv+Mu+U1KZtlSJqnSb3I1lZWGDPYw8nKPqAtQClXZXUxyjs2Ff
WVWVpFGncdAO3/wKZOofISCJnILTGEyYFR1ykZxoGAuB1VX3J9E/TEvOxH2gDnA+dOyGyCmrkEwC
lMP6xwrIskVdmnfv9pVpkmf8HPB1pvnEhIptO/iKQQap01KvC6tVnMCctRcSyIHry3QSM6oR4J/C
c8XMTqITxCC8OnT21ZTu6FJlNb17cI2588Zzn61uCcBQV4K5dtPy3oASIB9v/fUd59YtH/geLRmB
zH9tsr18JU9F5I8gFtucLYOZqUuQ7vZUGgdMTeIDK+kob0SddNmOANfBk3xDJigxSiOwB+rtaxae
SW8Aofm+l1YBShOZBd61Vf+YSAyq/uysq7Gbugyfiv8bTRZIUOLTmtQPPqoZKr9l/7I0UJs2TDN2
zMwmZcBGLW+5czZHwQKX6ZnksjAwxNCySN++z8pKKHcdyHQHTwmLokZ7QVdS2liwQSaGxGWit+0/
0BAsa/7l288JSZZ/3SatR/Y6ccXSkDwvrk8NiNSeYC0xYCJN4xEt45ax0yZOIOS+EoM6UmReFm/F
zns2wM5bKd4mRpGA046I3UrkqEHjuCFN3Uw6I33OLD003Dv8PUFjkUmSY0dP3bik2UOwMaa9x4cH
SHXT+tfYOkWs2oVCdE+Mvo80CPpaiLuoh7zq10a2Oq/YJFSnBK7JC7+KIXNPDEonb/+/h5gsTbLV
KaklYyueTjKqFiWFPDzMehDDjIEMq4ZNiS3x2Ld0gj/ES29qfF39rnaIJxhRlIHWGpx7ApEXGyBn
AslYSn8qStuwx65rprCkrAPIgz9DGSXI6PGfRTWxyzstGqoZE5Ec+jF/LrrIojkINZCS3lyxVsw0
4VvW3f21UAZ8vQrGuQr29IPPDjNvhjqgsFveYABEorbGlYM+QfMqRiqyEZ+bLe9VPE1vEHn8HFji
THEcOimcs81vZXD0xv+quuCZsp9C3v6lQFCXNCgTigSQN9DQDF0WdOSLlhsxRQupTUP4ms9Cgmsh
/+RkVIxQaLuzowWkgQ0kvLx6J9jTZ1ebXaHQeWVmenDLJqNrIz8FDZfFn7L5LQmwC/JhW/C3C89g
7QDzC8RHD4uQAAwSHMIEm0boVJtBumwA9nx8Z4MkLlyKcBbcIRLmSpoFk1oFlUPCd+Q2K4Suzo23
hHmc0k/ux4xZHh8O1F8/Dib9t7xFdk8v/9o9kXaAkbHK2NUH7Ln1nkU1paV76RYBmGUTxMXxxdXT
M1PqQuq+v/wzGNeN3u9Skcn0cYdlkH8ip6qP6RiPVF+7NHiDMKhjPxN48sVsoIqd/4XbDbHsO+AG
8q788uRe14qK25x+pejs2LWX4eYOhqeBtLRRMMRj5bHGeME4M3sc0Fc/gl/9XtD5nb3/+nqqmSPV
BjlUzcskmB/kySDas/cEnmlZUanQ9i4o1vMCKz1O5KPWPdmcMXz57X5uc1NO0Um2Lqv/XkMf4X8B
NSJOSK5zEOb/gdIUWdGXPYQp9/oflFmknDsZ8fvrcnATdP2u3XIynKZkwR1O/Mo+y/BZHL+K2Udx
jZC9EygUdqLm3Q4EViLDvrxpp1XwIuDlXA2ZOBXd/+BM4ucEmGfaR9K7SOa2wyWTX3zOtIMvnRJD
LF8jpp/W7OlLpamo1zaZKCDIVdMNL/Cbn4rjJkKZDXC7fkpVGWIE2ugO4QCRJFV0LW1bOml7kUV+
JvDhScRm40agxu24/AC/CWtrqO84yDDonX2Gg9QRfI4JHj87BWQ3G5bAZtSjncaHR8jre0hhwM/N
Gch7h1QVYX5r879wce+D05m4HTXmvz9Vclw4gh+SfYryccOmQ4f7TNHw+8F0OMG6ahRSJ4Y9cazZ
pKMeDus5EgBySRCJ8ATU4IPwV91B9jw+a7TlnhfBlZ3+Ly1sizaw8VkYqV9tPyGZNeZwn6Jzp1Ul
TLUmZ8Ip39/ZQ5F5ylSVgV8B6WEo0p0WLqNHO8ehqkSPKozKhMe32deNDEZITx9LwvTKZKmVlJaw
IUK2bewe88sWZ2tXn2RSP8Hzb21OE361zsFL4K7sLcMvWLzgKqSjlEWSsT92zvsjXVBu0DXV847C
SFigHq2VaMYKs2VtylVdXSr+IIOj8wAPGb3yTDiz5gPmfv+okXNA/GviC+gJ+rOJVrezWBjTrcIp
ry2WIGjuxG1ilYrHSnbov845RynKdq1InwGI8TTDdruuf4G7m93OvvNptnDTEhAxi+0tr9cGihvM
l3hhzaBN7xt3Rn4ssnDnbuIJ60ZMireuwtwUT5BmLgLdOpt1TaGaFQMWlC2/COXATJW1qmgR0oyx
5UTaSP586pBidfzs1Yhqd5/ceWqVjlnN5+ftNkCPTjcv+IBOyksBD6v5waK1XIQcaER36JuabsOH
/jd1C1Vc2ao/1aqR4pWYQIKSVDvEEuPpwKfPtJHJslcGcA1NAEdJTJ7oAbPcJn7NPNp2ApK0ZOlk
SYNc3FjLdPd8/1zJycm4bzRjwQ1UKz54HBJbUptbBgizeJPaAPOPWhqayQ6TnhI+UfVeIM7nzYMK
zKWVGFgnKYh7iM/3PkLtoQCr9X4XVdiMMaN0ws7+jdRoMo1tDQNCs0BEhsSHayotlGZyQlA+CgPW
llEjnEKPBn87qi+7Va+YvImCFHNgPMeGOLJmYPzvY3+oqGhl43W17JWkWwnfwT3pRNhllftbSOa8
3qrxSpdX9q2P0RJlxPZrVF9D0Sgh8CfACgjrm33zCFEK/+vrnEu2frTz6XL9F1Z52PF264JZNYDT
oe4DcHY0aeKCZZ+purk41wN2h5x4TZhc5SqTqZGXajivwVN9rYv6kf5W33EVQ9FWLNf2dodz9hb7
kFJCdqSSSh5JIxd04zJfTlyznl9mZl4mJ+LBrxUPGFOkkBCGDSFj7Lv5Al4yf6kPZULrW9kVvVyJ
6vx3dvjV43qRzorVwHIvdb9LtZoR8Cp45EAg0x8F8fze3DZYRyE+tWucrXUEBEp9wUYtC203D4M3
xJfQJbWmyAuGdvWFDKqAHLDNmoZkekBr3uN1CJCxymzp/9mcBw/oC1utHHkHFqcMnJk+3pCNHHDx
/Kqf19MnQGiQ142duqTOWs8it4nQSAfNkN9Q8aF/fTKKTjNgL9mnarD6MKJuLJe6OJxHH09HtAzI
g7ZTXCMfVIYphHFkpRK8pjWEwIrEPXlnfUh8n3ca3TzC35M2GGfGj2kkeNNrcXHUn5L1EE4Fzrqn
8XKDnUoqY7tAYsWf/iAeVyeGSduFAjVL2Izqrqtsm66K9gUWRiK0FufH61RINo6tL43jx82aLLuA
7b/76EIZvX948flEtwoCSHWY+z04h1XvucsfIhQNLoQMWt3Joij8HzW1I695IkJOAhfn6p9LneE5
Tje/tMiYYfS0mX+y3+uREAp5lkAdjsMQEND1jbFscBYRTmeaDdRtHY6zyvmY35KX6hyaYW/yVE31
D3OBslpCeEu4a1u5V3WyNuBAWG87lhNsoGEqU7wK4YMX6qRcOl4auMrTnyKyDiiYMrnvk41E71GR
n2N3KZeggF5KMwLZYCZsjSKgIBotF0AWx8H9WTp0Cwh8HxZTpjgKLE/cEHGg7WKa1h/GSz4FQpH+
AaM922/x8OVK6yz68g0O5R4Jc5kIEZZVFuFQxIJl3eVDSn37oXacOpDPRZKTQrbM7ELGoIsPfEsE
dKdOPrS/Q2ptzGGHnEASaAmSL5ntudcB49zZvsGPUs9OAiJAorJlSapM2Oorrh0WQOV3k80AXaVi
YM13O4a2ziK27jxSjVb/HTZjh6DiF8UN2okLruxV8tS81PRi8Cl0m1SpRyZBSolHdLkJRf9qWHXC
luRvz6+zflGiUB93xt0X5wFiL+G7+IYIT1px2/mlamTESB8kr0R06IqmvxwTrzqxDAgsAPaaPMYO
zCHyLNJQSxVfBFC7ZH5tW80guUoe65hy7ZXKGZba3dovnMZA5i/JU5IuCOCEePvMpWDOHOCxLmSP
VUcV169/zpKbPqR7uXQb7rDjOSQhz/yWCsHYzmbyodavGRq+tYbA/EkqhKd9X3rCpiMcwLY1lt63
HPJzLTl+dqWRoUKIHJm+UAF9NKxvA5z6oaRbZDQCDDK7sQlihx+27USY3tXBpQnazCSS48YV5nRU
0HvhPdzvxDSCVaRsuQsSuMkTIT6OXJKhC8AbKMwN/c1Dei2IjgroI0CxlwsjdxPBIj6j5yGOBqUY
PPwbD1r6YtvE2bBTKXgNRai0cTCWs0Wt1XBs5ZllUkK+qn1LMF6KzpjZ5v3NqNvqkLD0x1Yy+RBA
GgWFfsIpzeP6UtM8JxPU1yVXftOuIkyUHMhWFClAHqMURPyczKxuDbDnP9OKNVaHRPanueP2mLDW
BsAA36grmbja+R+zYNGjOw92XJPvF8J8VUM1Lq8HsE3ClUdow/nV/h3p9ARnV+5hRNcXhTZtjM9O
B/f+bTHUmM/irQTdkJ7YMPHTXGitWFgbSnXK19QnSvr5J+2Jm8S9549mluePNIYs7a7QU1mAwbuQ
UGIm7fH9H6HX6WblD+jON1X184luZqY9u8YHug4n2gyVEEHtPiizu/vxbl5YOjp0P2hdzO30DcYp
Cu9M+fNtt5PSeKPma1cxXJEu5Eofq0EecNkNfSQ3ljZWBjTYssSJudvD4qKESxaaZeKmx3HIIDWS
f89BBA0hnoPn52Tw/WZTSUF2/v3XU8ZXzZfhxMelr673KbcmxS8F+9tIkuwdAV+4LjfAhYto1+lm
Nh4vwzLsTb0NZNXffmxJcziQ2cr9lYkjDXlSVsLN2KyXxBkuoQgk+Wrtqym4n7lNOuOmD3UOpIz6
10drJx0iW3qMAf2INEfhYa/BRTcmzmWhN/PVwr7pBJ6lmMZjDZDwrVD1fKFxnpLDUi5RPzuPkHNg
H7aj1i6Rn7w3XZZ7Dva18M/3n4Ph1swZc7lECiatM4727l9zp4F62qGuG8dTd8xhntZrLRITlXBg
QSDjXmYH/MGA1Q28xYJgzIPUSnU0ngbjj6HL5UoMOMv4aMkMJ+rLEBwRBnI/x7GV0wWeNb2EuHx/
3bEg8q9+PiD7kmvEX+++LajgtnPkqqIaz00j2B6DN2yI7nrzFUxf8zEABcoxC2igG9CooAPjmRiK
LyI3wPr/xknsNAfAUdfbKzDBTgTz27qMymuX/78ic711tFMD6r1i7sf/yM9gJpqBSN0/UJHb4mne
uFgGWmhtM26g7abgqRo4/CYrc+Id6hWUabrPy/7ckQSmpstK7KnwByqogQYsrQ4ckSQJj8VHrsub
mKl60XBkC0EZLXyGtRPXSGcXL63CEfKTaQ96zWcg1u+UHCURS2YVzdPKjls6wqoBKuGa0cqpBqZb
tDVnynO/98QdjFR2yfKcusqsxcZAsjmFnWlyfu+2mA4uNU/iJlIYrgb0N/oUFp7gtyPrRgDsCY2b
vZhYcll4tT+eZO8GqubIXuKgSwovnnnOWEbLlIxvGbYDsMYhNBmiTId1feLnor9haeF1LFNOS4M6
hM1R2OPoDncCOg3meRfOLorbuuipfd+l5WrMyE2I2mNeNT4fq9nIOGlZMQKK3xPl5fb8wr+Tq806
5OKFW04U9nwxqWJsWpMetNHhiSrweWLg8cgJFhsna3rwSQluqn5FqVg8IPL14fFyS4H0T6UfZ+A8
nlCzqQb4LseR+MOEWEjrVigQZsw0VaOaq16n/XELc2X7dYRS4kd3UA1Cf/ePUmAzqbVTdcsiCOgB
0o38uBIsPKOFN5138j1pjsNAAe7w0SKdNg0Jm+XeizAXKimsolr2uZylslaJv38VRdf2PXIGYLlK
0+D4UDHbhl/5wjwlMifYbPm6LGiptdYw7n5JaPVtbCA3lXHjfdEf8L/akKgrqBiXVldTXIKeY3xc
nOtQSY4kT1dgmTGeqeNBI8Nb0VP0M5SglUXw1UdhVBdSfS38vlRamOygGDId2EnFsX50/c2i+lQJ
HrDDQ2nNXK5DI4gTu0VESypXT8q/KQ0LhHxvaS1AVSNjT+DLpw4NxpwbgIcen2EVcnE+y86NUgKG
y1zqI7gDjVTmrt+rA+9s3kDjDAal4vwQoLKm9HSI86jGRpUifMeR0fahOyclQoGfhYb3Liww3j8Q
Z5iQtmgELDGxjvo0cPqnffm6qfFRUBn+BSUVIMYlB5WIR54QQRGiwr5up2F2bt3LWkl/UnOIM+4D
c4ZgDV/DyPR/eHtxUvrR/0tpPNBPVay2Wdse+WjkGidn5rSRK66DUBW3+9ciy+wuKwuVjgnENLNS
MRv8CngvC2aiKUL75BkKdQ6g3lSk77vSASZuw+XlE/5cbOAPBHIG9fUGHBbvJwQymqNW+giUQ+Xx
6u5U0eOCXhCwC7ODLTx5LjZU0N1nr44kClEP+OaQXwjRzbSKAmrgnui4qK97ZYKeJxNbn0VhrXQ+
C8l+jHsN3JTERWFZWuesAAjLEmeOyrMMSQ2tnvZ7oT9pxDOSJiJJ/Qwo1ojOa3XteWp8pEDcH7Xi
8S9CaQHt2Pr9jZP0wano/qbmXwsv/+4iXLqCrMUX7zreAwEPROVbX//ILk/KslOZBSPGLEyS1MtG
0swSbxmcUcN8508LL0GPCWuY3nZyaMHSeabEkhGDMLmX5R9tpMFsCJC4qbmt6N8KOcYnhziKznIv
mTxrCkrN6m048uKhJwCoEJqPUcTqNQ81sMCyCA01i1b1XADKOioZ+/WmpJD6KA52OppLmmaMd0e8
sDk7u1U5itdc5Lz5mlDAof2VOVBHyfhezQBNC/r+lD+zHdDNY0FZUU9oIYtUIToMugHGoI46zSkw
NYDtEt1N50PWbuqCSOjY+wUlOGid/Cai45HUGhEZW9hGWf2STcsU7SKCH06SN1KS7w1yFtnigMhL
z34JDtLyL26mICYkjlaOlKbVZE6IiPFHYVbenWX+0CpFyl0hFYOW1Bgd5flnh2Q1fgLfz+MtrnfH
oc1PtDu3YeEtfn+BmxweXGe2/W7h/l1M5KxLYHx1tgJNFhAL882Xp1n3hwr6J8E+qO83KHebWWdy
b2ABhqFmyWbPViOplhmK7KZObEdFJyupuQgMV53mqiFPntSsMvM5NN79uEVc8Hp9py8UvPLH9bxr
SD8UaRoH7VykToyJ1p9Kz2wkbCZoZ4QgPGEaY4HTOkIG1rps0Rt1ixZ1lTJ4KplCy0FFAtTJpk+j
Yurh9F2ofJ4tMm9z5/mQS7WPLVDFEuAFLQ1/jEzZNe2P6bt9JDXQZ6vfY6tk5YbV3nYV7Kpa+laM
6bRAHEYs0KPT7VW6ao6Vi4qrgTvKtwUQSzg1QxKRwc7ynxVZze3+A27STW+VlAw67Nq55McYXOYF
XSkcha4NGaUAuwuW+5Ezpf0qIV94c8pMAtrla5TCHqyPGa3qXuPBy6wdnXuvHh/MWO45m9XDRu5W
uy2e+95128EviurMjXzmlpq5lVtLnJ+7w9hazC0T3sfIQkHRpFo12sp8tpgEihdR6XPm59MFeAag
QE47Wg1LWCcclFxDvcD7I0GlWvlNkFJ7wMCzun1qw0cUiLc+e1DMrzzFU/ClY3m5EqMHzgwUIwTh
ghPGntRdXbjU405hmgL+7Youz3RSvD1hUfnFtFHBgxuJyupIl5IX8WBA/dr4FcvRZjnwhcomUjEO
qQ/JfvooUWVAmRGDt6NaAdxVNGCzy9/wEXorLhNivixn9fFJyw8UU5w3/gOF2V/K1QF3vrh0+tNt
QLTM7JJrhMBuxdkILlQiHyEKVCekA3tOwKFtj12dGeo0kc01DFiT8pYKJb6dPnO/VmnQxAw4we6a
GvrZLzKs07LKzCn3ytvz5/uFvf4vfP7IHSaca9PabsTIwpOXhKXH4+VZEsanHoz5jrcvrs60Jlhr
y5Wdc/0cge2XUaEmp9xRTVQZXp+kg2dRcd4yFUv5EuHvFFWrJPJvo83dKlid/7LkOTh1UsODCKmE
hjONDgOoOzoxG3wWQ8SgcLkC+Po09liYB0UkP9SFO9QtRog/jXtOjb+wj4psQ950Cbgr9c72dFjo
wqzzZxYgcddJcwZ/SORhxiApGvyD3eNQbQHq99uTpSvPoQztdxfOS6QiTOB66LDuT0LU7jCzO2qQ
0tcBaalXTtQ1zZpj5wEIoE6JrGCb64mt2sK+ha9i42fViJg2fKI2g4Emgv369ZiPu4gK0gEV+Iyy
TLKPgGb815GRntm7zWoOeC2gjgTJzxayBelbjz0gD7Ialma/hIXXzzp7ylE46q7sL8/5um5XiBFs
uNYzDV4YUZzLUrfv8gV7srnQoGvZC43xQGOvMyxnNNSSl3BEjhAH5EN0LWCvAhqJ7B4YH0FpA6q+
uApmp/JXxj5S0LgBC2ixXNFN49Pt7Cas/g1fvojv+CKhxoctRRHdvmxqmGSZNuovlLBZhTxJtk+k
h3XJjB/roriF55jkjGFXKYRN5e/8xdlm7grgUL3TfqCeKdDsiKzFxftGUnwQ9d0KmCSfa/giiM5j
r/fHTa8M22d0J35qzr1AYYzwbGC4mbJzV9/nPdX7btpNWDG4NVrpHS9rpQIA9XTzvRpjevkw/W5o
lPTts1F0SJgLHlJlP3ncFXB2nEz2fCZ1y2tbXVZFuqmxsaFkflas9e9xS050vahi3Ood7rIYytM4
of+IjhFAnA6UR0I7g8f7pJE1gZtPdzcOCQdTeE1ZSqC7EJU9TlUi2jn6m34HykB86RB7qZvF85GW
Wadf9tp407Un35tB5f+5PzdL4sBeBm00i+1xYWTFJ0+aNW1avSFYJaPySyCkDDLZfUrlB90Rv6Si
r0y+sQ5gmp2NlfRMsQPHoIxGF7smVhG/NGiknWRrdkWIUWWh5szPS6SAzUr1HVNtgtY9R5daPW3f
8aArv+6j0pdkSR2ZE2xSmfdunoCtujND/xV1bSAD+yvIKTJPxxumutZ3qA2mBIPXNMOB+ZxmgUj6
i7LKPxkyg9JHHQKzxuujRwV9+nfQ97T4wX27s2+zYzFASFxX1Njy5Kh3RiB2B9MMxft3wHDhKzxx
zz19UB318WIuNDXIoRRwlq64u4eWgO1rRFFa0l1/CBlehi1Ga4au8bJcQwH2TjCRNRip2u89mizr
miwA4Pv+bilkZncldVYboh/7nP+7u3wk6FOgivq12SpP6vF1ObvXdGMfdPScfYdLZLpiS7Mwg3JM
4wFtpUb6XdzugXpg9To8uDaTuj0bgbGeKVy5+kmdbIM13BmjbCZgku2cXCdx9BplLMTs8VdYwgyB
XDI/Qh9vhrQNLNK5laZFunVMkVQgLJLTm4sg/wreZn5jO+8zBktOlOxXd5wEmY0SiST91WFUfcER
uzhW5xkgt337KqqDzOn9ryp4EBgye3vkquYKqhMZSbhX7YD29Idyc+2Fhvx6noj4zUHJS9udMmrC
TxBJ7XNHscS4oxIEMMPAfcrs9ZB8ZTu2479c3n3bMNivq2xqUaBgTO9/mhI0vQATYuXZQBtxSWaX
3+z8osTb/N9wUSzigECbkOpORNlCsHG+SvMGTseN1Vn3S4O1vdNdbuxp0ath6t0h1OXrLLH6U5oC
T7NguHFM65vETDRDTNX9MxUHL59g7bwBTpPFW0mC4O+RGDYaXMyUmHlKWlNK/Gwg3LhqMk5aIIE5
clTBg0H2PDXQq6WsnB2CkjanosLfOfCHfqaqebi0wHK4pMQB93H5ZvZeAHoen5Y2P0/U5GFbQMi4
6Q9+qN3IbmIAvZtWr7Aa4955aMEjx0s1v3rPBJNvJI550aY8io7KbAYWspjEKevuthPkz+NzQZFS
fqQJ5oLIQfe1q8LJeGE0+C1m44/wvGVqQ+Rx6CT3C+rCwuua7GWbXAHXcZ4a66hAB7BJroBzubCs
VWNrvfX2xcAZw6hLcmddQXk+KgIkE8XbnkiBdXsJ1y6QAC9AoB+60qV6O/hGk2iPTzeqPPZRK2Oi
pbXdfHnrHmh9IDa3zNdjctBtji7ja2MflM8bNA8kWlgS0E0HG3iteuJoEHUkpEeLz7VUeDDu2q0q
HKpjlAzLX42dtl7drabBsdVayhSNNmNAsCIb4C+lR6u447uSNVUWMCXyXPbMb4r5Io2T6+uhEpnT
B8HtWii6N+t/LZ80FeQ/ySQhqbpCkXjYXzY618Qly54ckqjBq1cRmcI1dHNxw6pwkC52snxdOMab
KNGkz81/o2kzoOTolmORV9Fai3o7Uq+25YKjUOQlD6Zyv9lE/UuEaP7gzGYu+oGd7mb5WAd0jEVG
o/FYcdn3hebkUTRjR9fkq9Svx4bRvyPYla6DU73mAcOKAn1MO7GQXCnG4+4j9Bgma42ePwx8ycDX
UoFWJOsbEG/L0HS3SgT51z7EgnnRQjlPRKxJEK8XYJqGa34ORpnlz9fFp/lXTjGaq+3HVL/hmkmc
1RZo8qWQok9EZ1bxJoAUIW2chP6ROX+GSm2RjB7zRzAqrDwvfaH6zdX5uqR90pnu4OyqHnmJYT/r
HrHTkpIyTnLZ1c4GAmK5oxcYZ9FY9Xv+L5hUK5BuzEam2tCHI40UsaqnGU36CdTLMeEkI/pCTzwQ
n3eg8+BmIjuScPiTv8p8VoEVXtGae7G7Rm8TL+HgkDk9YQqgjQTzx/71Uzl/My7H5sY0dxGfCZ/G
PF9Q9tFgYuY8rkKFGq4pEsEoGp/fZuxutHYiiaDkb5/6RUoyYGg7IP1snT9OfIyUd5VvBXCQdlo4
1HrQg6nUmTp2rLGKThhClQdg2S3JRK/gm57Qcoa5Fe5PJ8AnPBq2g8aKO8p66lO5NzW4I/WASfOJ
Q/Iw1K4PqMP8F1AqpqmwT8ukakEB3STTtJXOmu+ilcHNMfH91vz7mUE0CGcMtM9z+keEbSvGoh+t
OiJs2B5MoE1tQeWHlNpRbdXaNss6dSdaP76p5QuslmY1ksFy1BJUVZzDAlPjJjgMC24Q62TKcjK3
WjtIwmYkV9in0MZjY3Kxpsv6TX0fF4tqY/dCMmcyLo/azhX+DrFUz4+is27axvvJ57A/SW3nz5Dw
zoGXJJ/KbzVIV08k78BChgRuBCdXJ4mphGMjJw8Ot7945jQUCCrz8enMoCyI0lD9ccTbnODF+hLc
rVnpzzlIch6xRseqR23eNFXEh4D0ThLz9urHP7REm5JVHw73ocKzMQmBzrx1fCDEhqRd9QrLYrqu
1Q8Mu9LiwtdP8aQekYTKdpsyPs/vMrPn8+nn/S+xwZr4WOpq1HHi4pD/57K45ceXgKF9UBJe44PH
Agp6vHI21UvHjPepIBuDDlOor1maqPcN4q6RqxNdOxNTNKCmsoX5NXdP0YtxG3l4lEO4TrfI4siG
wb0mfOW4O7MVA7xNGqFEOa7Wnw0VuR1mT1Qv8qwAhyjMwm5HazgUu5j/pOfZptw1qsSvcqNWLvxi
jtkyS8YCqB2d+Mv/gXY0S7Z0+g8D5Zpk9+lN0UDe/3ML+kvCkI/TukW6uu7S+dHN03/8qi90Ne3T
61qzohYQTta9OEaNRviWgtQD2PFyz3fi26feJH6XKddPtl7SMCZ1rKbsWzm9Ni1PYgD6ldwbB4Ky
tb/MxUd4Ktr5X0ExbJPuO0Jam1+HOsOU2dlaKTwCnIHQgTVlkMAlunZE/y0kD/Va4c/RNHyXAHeS
XmuFYZulygEtpvZsmmn1khokE6yrDENsL5wt5qEi2Nhqj/yZ8kmx7v3PrBgFNctkXrP7JvoJibDF
hQRFCxgg2VtmUXbS8FKdAasmzQ7ncoou0cl02l8wdKT+ymB269BTJMOYzd8apC7weqOaa73NCsaP
ws3M4KB0QqBviqsN+klWoze/E2YS/YNBa37FYuRKBHYEax8RaEgqOVnUWKcVJHqM6UVurgeZLeyM
/ZjN/hdK1f1l+luTUf+OYmTM+GZ9OTyrnRdhzTbVe2KpdKVSSRHauh9VbW2jbuyS7jIxteFJI4ng
Pcr+Oa9v7JEOGKEeeM0i5wiBGk+KjoC0B2491Y9t50vYqmKutMF3gUlppgRiKB9Lcy6zcdTKecrv
7ciEeZWmEpcGj2n7uvFOatftrv6iErtfM9u7KYnunR3qpOVut6WqqaZ/nQfo/MPV/LmF9x50nG4V
Rxr45kZJj1+dYcZULae3/LXLFUH9KnZtrd+GnVgyhC+Fz0PxVBLeZnY3MPomI06G9boTaDKrvFIE
PNaqgaXI66kEyRVITSxykm1HHbYQn48lGkjcULu+SJTxjYnT5rj50Im7cWnj7DiGAP5H4ow3i54F
6lLJpLH8Ro7emiOvqRt7BnXvUcngtUJj+43pxBwRBDvz+ii9DVVJLQsjDArFAIEbxrvrMhV963UJ
2F9NNUiBvRtODqme98vYpDK+wVhZ1dRP6AlM9O8AIfEDWiyAmL141T+XhTY5mncstdNdgW4w0oFj
VCmFx7A9co4pNKc+a3oyBalyfIVKbsZrFu1556gGvo9wTdkPrwsMDfVSl3jomli+qfnlWHQqj+5X
ZaaHx8hOx6bF8X0xdvnuCbCV3FE0Ct6fWLLXfL4B424mZT4FAzerq6o1FCvMbWTFvyC50rSo25YP
7TESCNGPjrCxCefyq89/cbptagxHQXe1zmb3doQ8F/xgMXgkall5vWqHpMuXENbCmUD2wK0lAfcR
kHE7hW13Xv83FiNrG2lVTTSDsuvHO61kV8DfSxXwbVJjemjBiZDW5Afauivwgn7VTt/M+k3duXDf
tHMSJPGQ8wKmfcHdy0qdrX6vviXhH2BGNpftoTxg7h9L0FZ1Nx9UU68T+HcfEc6NhJ1NHRaSTG9i
l5EuqaUolypfS5Au4M5S0dYA0TnvaEbo/CnKu4IjTeRrrVkgpy9+cDD3aOz/x876OUk7eE7jEcLi
cmm39b4Ewz2tB5irOaOg4Yf/Gg/FD5RYXkXmc/4o4zV0IP8afuFXsyV+297QSg6XhrJQZgppmTei
KGPxMNzjcrv5BUi6veNgLbewheF8x6gjdZ0IjUhoutTkECNGidIYxvB7lJcx7KTrzbgr0MkoWKAs
XaB2PAqAEWoXm6CuPFcXu+9F6HFNWke4ecNMJl5VhirOQ366D3P7nEmGv4oBqWkd/vV9LdJCxR1P
fKDy7YKu8pQH6SG7cW3OqwtOpV8wa1QKeOY0qCCiI/pG0oFd5eohuoGy30HhMZTNeMtTPQPlsiVp
YAmd5u6DYtGSiTv9h4wV8mpvlL3gUXss98plbEs1zoYFmgXhMdYi+E8jf1N/KxahOB13ImwYOTBy
Qxprlca6ABxDtc+yrLkaW+EmV2jAfjjibeug5v3h6hFpel7kXxI5OfnhIvmlTbwaZi79oTdE2rt1
jNrrBBIcKdPOQUcXVFF4EOlW6YLniSZxcGgwzEyFols9AkvVuKJojL64ZfzBF41bwUXytRDBb3rW
SHkyOVCdlFb9Sk1V6JHBkwyiENykS+Wfo7xZZNUrRYM0MyQXlb6MexIAWvXDQNOvw8gson5hFwSP
rYo0Op17B+y/74ROQVlXSPfsoVgeYk/rYH+RMB5jO976oovxvlRElQxzc1TFGOuk4Rv0H5H/HIsQ
GVvpo8wIAp+xOybgpgaVXDuwQQsVhsW4S9/81AuY4HXlqwV1o63qxU5c9rDdiK0ALp3LCJcfTIif
mrGMCMY7+wTo4j8HoB5d8AKQRvEB6ABgfp7+VOy6UOCYtTHqv1N+ayMeBgPvUV86gf8hLKe280z7
H1xUwnx+hhMEd+KZClq0J7ojxPxflwNNqjkFhzGOCj9xUgY9HSv46VvMU0ne9xaFC+ulfTxNFodH
4d0Ym0NaZLc143b+XBREPZKnVIWF2JQXDv61ns5hhhZZrNenMJzEE6vb7t/pBQE+aG0iplUImkvz
rgeNvPYAddCguqDyXVDMSFO4w8+w7BCK61uEIngW16wXoTt3JKFxdoy2EqPNuBCGcEu4AIeD4vHa
d+POgesoS1d2OouGcsSXRNWK2TZOzCI0tEP5qKKiQHXqJUu7cnBjuv0r6CWbMEKi9bUtftGdVxNw
2hdeI6J7+1q96C3B/8pkyE+o+AMzCY/PP8hRuVC28htt8H5bfh9OhZJn+3TQrRro8B6PJX7vZqwk
I+0oZmLuORO+5HflltPyNu2L7UQs01cOb9MoDKfWEbHP4CRHlkcVyMkpHrHC/vkPHTVKsHv3mgRH
4d4+IdSstOKTsSZA9JI+sc/m+KFAme207RP9UOyprHVC2LlZJp8y2fm5PRXJEHD7aVLfnEwuzcZn
Vov9/XMh9kDhtw2pmrYpen1rgxULy1lc0dF31WF9f4RTDYuXNAfRRtpWTFZjGeYlVNfSwS1eEp8Q
PHdZQWtJ7t2wjsk4UlUSMZoCztf5xvT19z49rk93PMaRofIiLpWpFKPQ1zYzlPWRb3eQdpBzUvQR
c9bP31JONAmqdXoCt7uW+u4MZQTItgi334QCmLaff+gcvXBofa4KvIrkJWD8S1JzVRGuTAz8acH0
7W39vhlOaL2G/7mPKQWaHQpOQslY4lkUQF0kLr9pytMc8Np/zTs51EMrFIL45WubOZRNioDWps6G
hVgYqDBk4rqLHObltVYuT/+ziLr/eS9DwNBvnAZn0l7ZL5/X+rFoe7J8MWbrZk+cn7lzSlhzPEr0
RseaB2GpJsOqqQ01ejr1GJg7E6k0fQGDJj84f5bxe2cW73VRP5L6tVZb9LR8xyNbPpZ2cOM7xcuo
oWgZ/8unXVb0q5OltXG4oqPFDbofCkfgpevUoZdrW6vLjEp/GL3B669zO4AQujVUN72Au0oIyqc/
WzMiFbXeDCj3GX9nGcpRW4NWITSj/OWhicnLx/ORRPvK3FWy1jj2Yws+1MF+EDXsG8eKZzUHyPRZ
9N7t6h7jloXIUXLfojQML4hO6FO60dbLYuwBN2x4nR/2rOxpz69vBPEkBTOq1JERAwsFnIKlp0qN
+qTBLqmlygashzrKqA8OTlCwuieJX1QW0Iwb5h7NQxrnPOAq2tY0ez1TnrxS+Ych21Arc3Jc1StO
kszuKta7eJBVuH5aeXewKunPH838t//IgkXDm2rXLjNAgPzWK7pio8YvDpODHrrhrzCPrNzyVjNl
SnHIb6dNvCo9eQ5VD5xDc4L6irIxzYR34NGoileDgJ0ydGmHedrNXJ+fq5RMcCzeoUP4Acx6HnKH
rcG/rDwSs3uNO49Psn4Z0liM6sr9Eb50741n+BIfoQBw0IhP0amPnqophCoWd6wC5brJ4+APXdkn
rDwDPgyoIc8gtNM3WwPEAEovqk2hX5xpymZeac0jd4yOoKjdCRcbObXkkRkYeN7b67RpW9fjM2yM
Vm7NI87fDeC3iMCzm9JcLFy6R+mOjur3xXnTCDg8P2zPfLT5A5rpXag7FzKa1bVQL2kNafsAN1ce
jIhMcQLrm+oD/ojFeytatch1a0kquA1vhbOrzbOiesquSLY/xx4qolB2qkH/yKS+3awbaNpLhn9A
xXe6tJBDJlWhUlOW/Q23PMQeTQ5mYrpdUqN4TalsKA76sAOEy2f2dA0fHQdT0fV6TkystB75apAX
HXyyFua2n2M8rflJauRzSnH7AfmdVyO7+j6FjTN3/OTiUAeqh/Ppal3/irpfY3Bpz0wHYVsf8tlt
CBNvj6/I9nBRvhmyKzUf9lR3+ORc8bkE0je0ODQyT5CkMIwzQIvpDQq6A65sQXIi1SGCb3AWmblX
AYJ7TMgE2Nt2gmjEX5icl3MHk9vupem4Bdbj7bz8zi9QkoISGZ7CJdBPiDK/PBwSPawCqW5k710P
lEapq5PIE9USMEFFPLVJoBX0Y+LXTkbKXsd8v/Puiuls9TBPBJZ4lllQnWcCHbTaSSSpDuu4JL7a
LUffqmQW1gAk/GO+xT1VIbEeuqOrMVTMrQWYdBk2CP/z0ldeDZmOo/dQx1TQD2BvrL1PTmxxDCmT
cjbZl1aJ6ZCFeVVGd8kHpImFkOcWneQbvgG/6ORSsnYM0Tfv+RpqpCH0sWOe/0AjF64YoI7bN+mC
keGpHbDDNe+o9K1VdSSAKqcpfJJaLdl1gRUeFWuL8V+Uk7DU7T3zANXQPP1jL2mDNsFs36LHaLoF
CGsvyyJn4WFjMRd9iyQmX5d1BIr86c8cmWoAMx2o9q1XUbEGH7TMfo9Hm6P8r+DHp/Zj6R+xtsU5
t+FqLQuxhOSi9nJqqOnv3cdNCJR+oKQX+FBexw+BVtjq2wDUplNunI5JCROOkffS1SpeESKuqXQ4
P0Kgi43o3bB4zaNnG8S5XEAdU11nfIQ3GSMZMNqsM1nxttY4kX/IqI/6RKd/SjfKvYdp3ElWL1/q
QJmLRuZpLwYltLs6RNrVbAByzmeGSFaS4/kci+5gsqBWzXdEjdhn5FqScnxp4FDgQaiHOaiTjcih
Kwv0nbVaZFzbFTZaR8QhFTBfYB+9V9IRUqcyZDB5F8VfmEC5KFAAudEAAg6GMFSVS0XiGBU+Hg01
++x4mhivTIZBufJ0FjuhLMXSC1V5WK3YfrY6s1TrvmBjNMWfhQ3WPQxia+AHTYYjVaWi/YwGE5NH
Sj4KPJODx7A15XZgrFKPlcNo2ffaoHWdbDkFQN+L9K2aqD8aHG+yEcAr7llz5S7U1nb5egwC6FsQ
qrh0Ml/YcLWp+jTnrPtMdreIFkJkN7GBFNQEGpPmsXw8gw/FvIJBIeyyKYB/xceg82Xei7Abg/Sv
O2OWdcZ18WTivoOM83NFa8pr3LMwYDoXW1MKHXwrReu5rmf0ChYCI0QnWFlWew13ZT821bIIoXKQ
y4DjyRmxWjE+druG2gFN4VEzhCyqCBZ6fGvBnJdnBWgQyVvbs8vhvQNH/sH/H+BF7i7QmrIC8N5F
mBNBThWW8p6X45JtCREj+L4CB5SSQWrxZbEgqYYmGrE3vpF64o8TOsK72QPFiQgAKZpTzhD36xrt
LInk5HHyR11nwDv0ZwF1xbCkpt4NzRRQds3RUH8r3MVCK6V5+YkwhrNaMgiVwL/CJ5saNdL5HY2I
eCZt1IYiQ11ifNbdMPeo6imsJWeri3ZGSiMrahuJAOAdL/dVyORdrdrqra1ySN8REbEC9wpOjfFY
WygckMzb0FsAYGtsjHpsh5uzJwQdSZCBj/ammwa4wu7qNzdJBC7HhVgfW+ZLVbvWWHee80mGGhEF
P6s2V5Xh1yTHYBKtgHbscOT+P4r1zNCEnZH3sCNNmKW3a7FFGa0PkZXgdAfxG9R9F63TOgBZ6VmX
5c4vdqINPzPVt6DaOlYuaGV0UsQ02Y5W3j+uBAuHvC+C2y+rGUIH4Ycot5VatF4jCpFWp/sy5YdF
bPhjBjAQQSaxM58OB3AYMGx0+dVetuw6b4ykMexhy9XBVEVJKD4SVXDwE/5YI1jwKDVvGaZHAyZC
9Ap3+yKqTvMzAE6EpH4iy0VxaFhXgypHDTy6Zs7r3DgflGWxf9h7HGAlg/VlDHa2tAVGKs9NlAej
7me3e0kk2FR55BETJQS7k3vl6wqFfZ5p6k0Khgsiukpnm/AC0dxKPQTKLxSws1AGhiAXuS1p0L1k
WnGfR9NKugDE+r2rHrKqi50/9x4ZZGNNvqT+uGk18fa3lNRGJE7qOWKDEKVI8W1rOBxOjdmgnM8n
81pBeW/mq1naf840vE6goF0m4mmJMpRciOepnvnPknby2DmZgE0r/v65f3xALqSqyoGXqLe2Q110
LaezxWNv58X4AgiWSNOuSfFwMz9nDiOfIhA0m+GLs3XOhn+ySbkO7hIkAMIh3eFOya4JtYsHWkMn
dDnpYmq6SCHqwHA0b3LO1vKLLgP7p9xbac0pYQo2DyO9++P9iwULx5P1d0VdYGI6XuPqBmp+ldZt
2OICTV+fbQH4hzs+sZKx8k6MX3t5NFXImizJemUzeD7exHZLx06qVCSfyM32fS0+aqZQbHcSDGvU
58ym7q4tpxsSr71SWZ9Z5rPQ/7hAsdLpUyDasT7L+mt9xiYCA4rsEUKjasOWWqCqBrUwkbP56cuR
jB+Xu/sgG5zAUiXqnJobt32Ltw03vR5v4NrT1+7OsDQcEqBhASISRj3utxe7r5JxcTf4ZWTtKWbZ
PsL2D8UdGziZ7fhcW4gyAntxEcNZPX13vBZU+Qp70qyr47Mx6HE/NYCAfvibSztNvMU0YfhobHLN
ekIO2L6Muh1vnZM9B0eQfHhBJo273J+iWa61usFcTR01e0FPfJf5aTqKgAB8D6ADtI6vKoEj0Hlv
LZiQsJFn87WotXo4ytEsDVivv7iNI0r1385zgip7y7Swk3e8EW6/1T0G2Yn/AgajoJ76UyjNT4XU
AOXFVTaRzWhz60RTO/sakWhJyG2ZG4PKSTKiahoxDBHOD8DtuWOcgFV/HB42MWyBGqy+ZGTxIUNl
66/5LttHgxMCUHuW8OvtkbxvkQqzDS9lw6d1nv3dlaKrwlMIw8CGtA1vKabSe1JLlROHUFNYVnxy
2dp9osHJLyYb5GdP8gnXQjTU0yuQlkRwhP82lcxljv1ClAaWLxHvRbPMOu01+s3xBh5PECMFMdkt
jsAWIkC6TDZWmryeZBzRzMr5mCGoqCyG9EG/YjTrtU062XlnXS38sZOCS/P9JHAxLvwpePU9D6Wi
6ZrdUClpQ4wS5YTeGRYF+CcfIidFkMb2hlshsScWSmaFIrK9p3SasGCH3j48nEz00alqKOoOs2ht
ycfdXTQeDLGyQM+NkD780UsPwzwb24Ir1VQnTtMZVS/6Cs5Qm+tkPtFle5BW7TfPOw+IdiZUSLvf
eUZECT1e+ZKLVZ0d6+SGqEgAaZ+0P57NS+uAWp+d/ySgtCxFOgVQqhDg62/7RtzzNxxB2sDNQB9A
VXK3rMNFYjjNMF9ccb8/UITSAYy/aqZ4s8FT3YIeTzUzct1Bucd2jYn0Pol7Afu37DrpRhmGu1Ox
QuzAI9ffS95cejgXUl0bGQq4KvfMw5NKwTUTeU532rUWWXB1ZN8xkSuOszIHb+icG/cRi7hJB3Co
YjYoMuR0g9HlCxAtFrLM/2v8aOjNHiNnOQWwH9TZ0EjoLz8qCe8ERbkPYeipUuV33LYiTMlvVGUK
e0IdBmEiuOZxzvllO5+7g8yUvs/pOySJ79arVYNZsspDcSKP4gm+hV6DNpritLJxs2XIMp5Z1QoQ
wReJT187fqFvS4PnG20StnRWV3odrUz7YHOoMRGGYmEeonX0Eqs+IGWdwJ5aghwQRZkjM1Ml5G2J
Ae29RPD+gfcAfrKDfx6Vqh0eyO8T7ArWj2E1mnd5J6HTNPehBT3+PcaoUS+cJCt1tFPRQCLUK4Bd
g14jhFNHTyaJ5jQlEbS+xp9pmKdB6ZY8LjtLkT7BZt8e8dVsLo0RcmPUK67ltcqX2iF7EgkBlk1m
6sbIkuqhEByRTsnclj9fKIPY04gIyGNKPyUjwso7EU6OJMF4acIGpB+nSt96cOKhu3S5heuBa9MP
ELMA8P3A6ZFOyjYrMcmk1aejNdpNaYIekg0e4SfzLsJbdbD4pU5fx8xZEljYYnZysWt/FZHosRxB
Z5sldFE85WSnKe1d80UjsZLN+Xdghe19NnFSvPL4gJUnFLTbacJiovCaN0zJVgfkIltqBlT6ya3I
5Znv34X+1xfHwzj9FqPGx6AmdKeWJ0lIVHgvRsvtJSHFlmX/2hyss//DDtaM965Lftkd1hfKRjdH
mP/Yh+Z6GoUKFkAe4238YU0VQq/jRCz4hzKu6H35MgcAU2/xAjfFsksTGv5QDeo/0TJVCmLRmO/w
FuKN2vsizvtruw5J7i7QkaJ4ZCgY86uPWM6GxdUF/YOzqmb2k4hb6GW+yuhyafR10wIhMmlBfKdC
nShAr9JrsoDd6pfrMNIKWYupw0qdir0Zhz7UFdpxn6OF5td0DWk+QZthsW6rxYmVi3yKKXuiaJsj
19ipawodqzgF1gSWLHNYc8AXIWjr+4JXdQFlxRx7armZJzatg4V6Tj5Da39/o563ZQacg9i4xeI/
PN1PgpuzM/m7d95u3U/L28jBAfCNMGBJPqrVt+HpYDPscwVnhG2aFLxuYNqA/gIV89j2aii/WNQl
CAFwjzXgk1Ys9JjI//sJwBlGSm6uVz2BiuuLFzTaMrkiMsX/jSIqTnUtBKeijUjGqJlFXNl2LztK
W7vMKu864otoh89i71CdB31UgqfOC2icLu0Ho8DulVgHQODU5Nt/FLpqjNHI8178284O42zGlmSD
X9K/YiFcYrZ3VEBD1SGZQ96EnbdDIGx/FRExjMpDD2jHDab30ZhcGJFNyNpCb9HNs4U7R+5+pXfS
5uwod+R5fhyDvGUEtqeRCTOK7vdFY2kdVXgzVgp79HULE7+aZlaBr6ANmio68fV0J8eymy/s7o/6
Gfyd+r8G64dh6Ie9gYNxG/HLznjgJFM+R8ZW2PifTi/7HBUNIwLnpVmQ1ZlXaYExxVWTJ/G9HHxM
5aiHvMg4tT1uB2BS+xsvhQPQGSrpmFvl6CSEBm4ME/vivKDIiKgOXWXbN0TNNHK3Yx4g9pUBUzQs
A1PAl5XKCrnnGilS19x8RDuVtw3WL2v6x0GAiZbkoQJHPXE9CejVeJhLVeIDC91pWK1cGBKU2T44
UwGR4FdAhV8AeSEbz18exY4qVU7rF1oVnt45IZir/m4p+vAsBn73W8Mxeyip3p3Ka7PTg5Xeby7y
HRChMK8j4CGKLn+IIcfHz3vNEkjVj9Gd+Tw6kO/zaey1HXN4m7/Ir0DIz+OD87vaMzfmLmOcSGUE
BKOFE6mbYmPW2vxAZTdsL/obiAOa5cT9G19cZ97oBkg+zFzwK/PS7pYKEAfnh4RPdAc2/ZwXuBeF
9Z0KWj9T0MyIiCQOlQhxW81LueF6VcouqB+QeGrx3smwfwPFbVcCE+nZ1/CprwFRMJDBn8n2s+vX
f8DRShJPVxMCvBxl9ecuE5ENVmKLKEZsZ4B4St0WARuPGJ2TygpC3IwHH4JIKpsHwihtsnPa274h
Ypcl9iAmSHcXZzJRXFFFFRAssEmfJAHlbyLS12cgGPMkpwDlVTBUWWWbcSRq+v6TMgzxm8biQYKG
cjGdBbF5uMn+1bQY9szZwxGpfuKIAwxnJLvZx5avScZ+965B1DdkS2myZB+L3YDtde7xP8gyxVCW
b/IeLrogb4kmxBHHvYq2j9iHlM5ZEn24j3pdmuJBzCAAT7p94KQ9Oi2vqd8op5mbQi8YpM9cufqq
Uka8r7XzlNdsIe4MmU9rnSr0OTpKkOzvIWnb2kVBMnEQJ05qOGMaB0nUCv6AX8O4hTrz+mh2hRac
7DQQYSwtdsaCO/zgZxC/E42lYsnh+X0CFCJxLnzcvM2qv9Tp+TfUhDAgc2sEMNIrT2YdeuGGJuOH
8L7dWpCN/nelYM7cDHynVKFxcl8LSF33N9Eli20fnHESLHOcfq2A3V7pdVSAbyxdLu0LAjhPHgLn
q1fPAIhBvCju8bdnPxEnKnTkHck1++dstGSQ2sQ1IToYmEK2/75XEYDY/1rN41PnqU6qkfdf7U2V
PQsw4cJ8n4LZ9F49o+UWdodz46PhlEVWoyflHd4HaljjyHMF2s4pBNTJsV/4wsVWbHVVTdRoUHI7
JIaI5moTF0FySEGeV7bsCc2TIbmvOT6EIcNqsWVHW5VPlRys3VSmFCpSq4jPoOlviPw5zIh5W/Sm
CBv/9oYpc/HqoJkHiPo7yEjUigC1FGsVW/CSF9IdwvlItgWpoL1EUoElsqVjYPXX3ShUDvzQbb0K
Ow+Yle9XTVWlvsM/Ta8PTIjfLdxXvpY+mzsulefHLHCYFNaUCsXExF63j/VC8IkiRNlz+MLUwInm
qdUjVO1rzpQ7yakXY5W21IepoTBmxQa4H8eG7j36FnrUnZ9jUSxSWJ9nxwYXut6IlBaPtkRCRDHP
AGBUOw/QwjtFWJuIgJ7IBTAZ2xYfovxI7z4xYcXXpxUMzyrthdG/PWgb9I+wr6nohL6D6oTJf5ZB
CoP9JfKZBdvZAJ6KTkOWXv4+Ze0gYp/qtu3Z6EKSbTNjaNyxbgvEKJISm0mFaTWqUgK+4UXlGjvl
9StIAxKOfqPjI9EGd3kF7zLv8QTyTsYiSpnFIqVmrCB6AuLY/yxDv/Icy2YRCfonJ7wmjMVYkTOE
oYwLJXOGnkgAVV7V23WDshBSmd7rWRdg5ZDIbWuGFAy5gHJUi4jQubi6nmGVgVTDbUxooRrnzW2W
PnqHyh2ievEWOGlTgUEGlQcJ2w75cl1BJM+cwrSdbXdBHgNgQ4gMcPLLyrI39/it+zjyIkDYVRFq
1CWHDT8jgGN+lDOXPKeKpwxQcsf9yG/GE2f7Qo0VHCauKtAM+ld8C9orwnWO4I8VE/1+V/yCEF0u
l1d9bE4ujRyZBHQ7PLYHA+DjmOvvIbjAhPvMEQKPAFZY602WGnyNd/MswGLVyiBLpD5hduFDG3G8
mR84qg97tHiaG8hXbKoeidmvHMgegu+oN0YmTP5ZILWk+H3O9Fab1HwL2VTIgKXogoxRynsWfmOP
KZnltlImxOMq3ieKomxske83V5f0YZy83abrMllRUaKR9/BIAOT9kEUoyk+XRK1Sx6a1LcjyIBrd
va08DTYb1ikb4RioGoEYuD0/fZAGlDEg10Vxp9o6G7uJRxpEaXJc7isJ6HjyKTS77zvuEGZbw6Sn
MqDIbnWgiuyQIGtSh8TXkcsDB5auTJlTlju9NUKL3n3zXAs0M7UuQSxjU0AHa1Tv3u6fZd/41znO
jEI3HVn5lwFZmurJJ9r6HP34wphbUncDr5ZLekn6A0mM3OQvNAVsMhWGLIy8fWEGVR2UQiMzDH4h
rafnxAoF2ZrvB0UiVDTQKkM/dZH1O/fj9/ga0Hq1b8Juw/pmGJ1+SvN2CKyjoNURlqlCYY+fbf7p
/GJs7ycRZiK9JTT/D0O/yf/2CmQ5qKIA27z4WiWdXRsCMhN6ZxuGBk/sddKB+oCcL6jNh3IvfdLw
afT+DA0jInbZkK+0s39Pm+GmFmP1ka8pmqPUSl3d/hAWwqnCe83o1cXUWTKrK/vVccg8cZNCFllx
wSG9quKqSWQYCAnFPTX5jbmfowpG/A4oMf/LBmufzrCLcZkcfBIa0h0Cav7eogCVp3ZgzLbSw40K
etznx7PT0hkOllsIWyV0iKJN3xxQ5wbaPejSuZVsurybGjq3kQnI/ttEaka4+MrwWXFdROjp/mQw
LpdEK8IuXKWfXe+HhgiTEjS8E1Xc5JMV+kMlwov4wVUyzBpio4kUDJqG4AmiKKLqCyL4fN0VOPTg
UYqXBe4nWR+tMakJ1avuztaRHUGYG8YfkpcNQ+3KojmVNuTT6HZI8OuW0xKCV3Xni1984Met5hhb
QJqb9VFTZjtr7D0GtZcYFoUJvia+nWoUY1qc/KnNTMoy5fVC3xjDrDJ3M+gRzhIcjz7LERcG9q3i
ynktDJSNSiWbOF12xU9qrsqS6GSFQwHDVWyTY+6WnJtdZN88VGukq27WGx9SfghNPQqEfcioMbNT
bzVfuDdAh6jybK5S6k83a/d1cVbIf6KIZmX+R/uRwmRCEH15Zws8a0KZhgv7XMmjRbg14gjitvHK
YVDu7Q7W4J9sFTDESobxnxiRbtSPZ/QPxze1XN9IYwNalkCAM+nlunQhpBqp+fzQdAgs8vga3hY9
BK2zZNuDxwF0AksomV77Ok+yI0s3R8B/fWBhz349IBlBsUBwiFTw7Ql0R61kTvq1xqgT+Pzx4CmE
mgyTPgPOf8qh8pZHfzSzDJfqcD/8zgEVsyTRxhqZIPcAmNK8lXC7SiPnV5o4bDl8g94qCyzVObez
BUT8dNl2+Sq2B41cnZhYGALU400j91RmstLTOt+9YQ3eKboBOUAKlT/PtEBsBI7gdwifL861BmzF
AEHxgwAGARFP+D/8VNKIxpa52IYOHtw7yHf+p6VgEP3uAXDGWm69xzW3lhIusmO9WDNvmhj56La1
31VHEAAzcayQ1GKt7m0HUqLtCltlYUCu8MCGuJuBnclNTu1THtmPemSZRLTU/KyP8PYkzG469ube
9Imv+UW0I5nDqc8ghbbCn6vEYY741AVp19H0rd2XQxV8Zf/ehF//T/sr8Kw/JzdjpQZtMjb84xq2
JbMFSgG6jyClIs4SPZY9vbs65QPBdLJkM2TzxQ/8or2x5+3vPZHAMEVgNz/QtbvNCICzMSZttRXX
EPMxOPdJerUlTnraILiGwbumEkHYZ6qphNudlPkOgQG+72po2lVQIP3rGGww1rBNtTUw6uFrbzBK
wp/qw9E+tSLOfIgYb9O07/lX4GvxRVgI0x7GvsSLWSZVOR7DQ26XQYaNaSgbW0foxC62Du2Ei9rB
WgloOimLnvnmnYjky069EXOGgrBQy4Tx3keLbwAxy695TNge2r7EBKTYRcXrBplp+aJ7BcVXbUMN
ccnNfDvJT8QzZFmFxLE5y1FFS7FcT3X2/+TfOdpYfVsCoOst7qDapblY5z/viquaPB63H/QuxTze
S7kSJehHxgdbXzLwcrmmJudfPDlPr5ioIJkmSDmeyrE1KhJKhwQkDB5mKN2UVCVUSvYUoS5imwIk
naUy+aEYyKQX8rMOCF/m0lwEfR37Uq3/sB6a3ffO2V9pMQt/JIhtrT3YCr+7Q9AGtj1fw54UIAbv
xpTY3c1Tqxnw5Om6obJCY66dJaR++VoJ7oHgfMPkTF5iaZXV8UEVJ+EEldqDE49B/MXIqIqt4Art
6LSCB3gMmMxZF3sSd6VtaJeDiApzoL8vBxkVT9lRYrmLoCWb0YO32YAsHU5NyjHtCZfUnLcr1/zO
fdAUJyYK/zU/PG0EOBgVl0LRfpW6cK/pBy9rFmSEnuhdOebtLCn70eXukDGtVXviaRs2v2jEI7lo
dwOSX404vKtSQ0iuh9etNIWDjQQg4NegTCPEJYu6emN2jpMKSZ4xlz0RXVXBe2LEJgzDaKnwv3e5
wihbZORzSTAW8llISFFglRF6Kho/KTXAc1jfSKQhaWi2yFEY0M4KhWEUMS8y8KPQQ0x8dTXHztJp
YxKRmJ2yPMYzqqJN3zBQ6q5A19/IQbS+k9YkO9WtWBC90UzdBlHx4GwGLeU8MT1RtTPc6Fkvuve+
260j8xB4sAyOoMdtIvfrrhEZaLKd1Xih0TJ/+DwJYxnjMvzm7S8Gfk1fB8Tn3rnbgxUcNFbd5spd
2oUgpw+SM9oG0m5r4ega6j7y94bjCWSw8SMDPo1mZqT577kY51b/Qf887yX5mdsMkrTbRvSjdEXc
zhAK34Wu2iU4Bda1Ts5u4pa91LwWW8wd16oiY1ELa5J+18eHd0/erCBdlhblDO9WEiSqZ5C5QA0m
89rie9wsNDQF08wXlkCUepEr/ps9Ec/HS4vtyutzr1uw+/spZIO03IeLZCM8711Fi2ZwrlWoBBiY
D+f61WkqN0APS5lRUtY/NC82Qf09fQHSk4itpbW/V1LMThlRP05Hk2MELADnMIuE4vFmovphlhfh
znMEEkesB788ycpFtQZFOK4iUTY6WNEAvMg4WBnSVRlu/WV9EDTbbgbCz8cHk1AirVz6lzZRwoqv
NthQG+rSy9iNxvW8iY75NLYwecg/2f38+mXQV8AJQnbINO7CB6yE4g20xEtE4OClmcF9OnIjlpvG
53RxUZr9jhd+b5Ft7XLrq6b2KrMnj26RPTEhz5zN88FqwJ1wgsjo/TEQxBzUjEU9a0zBpQSVleBQ
QK04mJFW3lv2b3GepxKTUEq7EAxU3fcyOp5CcBb+s6es+jVg0F3rJD5p8BxHPggr5P7WFESw3Vnr
NzbwOYB1AKIrl49GFDUdDFnjW3yHEg5UDxALgY3kaDtd1Y1yfh+wgrnvBN2/q2xE2zm+qvCz9Ahu
hHsxgbQwTvV6KIb11MXJZLwzFE9dlsob7pEhvOX8z8qYYYIVGbRo2nt+t8j2vxNo9JQdRBX6F/Uj
As6oC+U1QUAFf0FmADkQBnQp925bQT/kJU9cft99yekSrdG/JqG8hpPoQURyZf/SeODRA7dYpo0o
CXGACUzG2nmhccKxFN9NnT9a+qSpHkMYxi7mIqKt/oV71yIw59hqzBcdKAQwMAKKNhZW5GUfB5jG
Sm/bBNRcoXkJTO3LXBkjV/BzlHDQk6yDj9fGaLL5GvNr3NpZyefjq4BO7ery26FJg5e5rQDVXEFR
YRpFnIAV3wsBYnBhnKAITrBEK24YGTjP31FrG6dpacS+iTkQ/n0E7ore72jna2VEmecClc3Lfbbm
YOejXi0OPUY31JBL0yUJ1N1Lhvcr3+tNay337ktCa0MmFRPvufHtSZk4a6+O3i3JKNqJBVwEHvhQ
GmBlKgAm3wZaxzbPZoL7YxloOGQWclm3uz2Xp2FTvspTfC5mTKOgnmIPZWWcCAyZmMQNU+mFKlUH
pQDh1d8314AntK3pDtDQwJ0ns9FL+x8rRv3KwMBnWd1k1S9XjTOK0945szX0PtloJhRJ0twG+oe6
j5z8tNVDu68dlqAObZOdr8n0xqqOImvj4K5GzSPGmxE/ZqdzO01E6mUjQPJp8qxfoEUGcHRc8eGO
XXnfyBlOgVx+dxqEZNsPrnwdDm/Xbmm9Z/jOiIzoVo58X5QCWySSHy8+chzYc/oLVAx+KVoguoD2
kIOUbOolR2yzb0MPXIfM1ebu46z8HlH7dps3ae+KmvDHoXWtwD1KVqygIrX5p8R4zmDkQdCeB3mR
GK5KGuW8XMU25ay8YfDwefGRRSMpjTfPKwinIu6Gd/53aTTZDh0LoDYGxchr6SskAJGftsdJtGLE
yj5gIuc+vozZw42nsehLNt0Zfvl82zWQFAN/9DOJqFND8OGbL+lpn+4oWoZef4ulTl3ui9Df0wRP
HhFyi039mD/DZJ0tOMdHNwgk2FqfYd9el9Y7EzRvyESeUlLcB9ebU+QtgJaeknEmGvFPFBbyTvAL
fZ8Th5S7qpp2R+p80ygu75rDyU4GrERWnXkAm2o0bI148CBrNgdKE+DQWhWYNmVXu4NWYfdirep/
5un6+fILhE0IJpLoYfcOMDlIxtn5XE08w7N6Y9UZGYEA9wVdKeYiazX2YhEGQA6vkhb4K4lOt0mR
+wYmJic1uOQDTZRQq78QwF0Nigp3uE9svHg2FWjwzbkiMWgdBE4eKXXGnpN1btVy50xNMQQs2tb1
ldK6fltzKroUwXL/8065LX9NM9i5jKZoOd7V2HVvL5Rme79kQ69+to5LYcMoHEvivtYWE6KyN+JI
zFtPGiZ0mJKFU95PhCkRXPcDk+k2gKJLX0dwUz1cPmCy9AO5nAO8gLWcgFU+G6eqIuFQcOjSSDF0
xu82TO9VeNXnPR4bLKyXFaz3gStyJg7GsCesgj+tw90HGQ4QZsst3LbvehziHPdx8fcby0tyiSSy
qLKRRLY1c01mQAsAW8n3Ex4PICnLiu57yDiXnoqQFWxRwdbeha7aJ293kgP4kNqbficiY3037aA0
awpTn78NSkg73IUcr8sj32Pu3q9AJRGJb6Pk2hIemO/21/AT8xCyC6OtrlWvwOI2J+AzOswm25b3
D7hrGrd/UAITkqQYni3PV95Fz/NQ8plmepmVN1kis7rh0C/Y2rbWhKQeVHCGQfd4EkeuO2VFv87t
2MLixYLJu9PJvS/7IFjhG/9sq/uhFPO7ryI6sn/f4cY4Q2CTvqFgHTmB9YTAID/S22IfagZyhSsQ
LxvwcvoJJFFh1r6ZZJSp64wiRtqQNDoSsNqbHfc4gaiUFimWibH7jstJyI5NR3423yjTbP7Yuu+y
yoS+G4e1jUzP7IojIFzZtT3tTbyOdi0ZnfQQidDtrDaHpGVPQr/QAUB3676DsqZhdLeGPSaeejaC
r7fexcsz0mXBZ/6wzXjMYD59APXBlkiVakWAo/U8DxIXRLXXFdGbVoP7/z6xfcfH/YOyyBnICXPc
aI3wViSyfhjg89cgRstEGBjM4C+GOCau7GrxjdkLXhNV9y7FNQxDPGh4j7GWVo4sKp3iQby3NX60
Z0tAs1EThhU/OghgTcTn0gOWccG4adqgNcMFaKg0dok5pYoVUVsCznjT0Pxmq1HB7kvwckzyirTo
h6lfZnpcScFWwUllLRMR3fWlhwRwhlRGik0ZUirJAf8XZ9rvQHNFLJkMl/Ha7C2YizwAyRgmS84K
lBOlIi2/o8gP8OQe6cvHjoj3dYL3kjw5DeImyLDM4mNmZ1RFUpuQXiy21Ea7I2GfJuo5+03+7Brn
nZelgWjB1k7h3+hPWTxtjxubYhW86B8101uUQL5Hs//TeRyvnTzkyPafU0D71bNG3qy/nVx55Ge5
nL+epnfKo8DWeVxzPn/kh+jEscUgwFzPgwVbZ7skBKtKFcAso6VvNt0KLYyllaKBo8QR6UD3OViz
BTlTXh09PrBcopELiZZA/NuJuhL3AFnRsJv2/S+GEZRbYsSfjU2XCR51SgE47nC08OsmhMA4v+of
4k0FS9I2RLrlOeX8xZdp98btoLhedb6F4WoVZoytfwh2DgLKM2rDzouefynnpO715j6tWXH5jhhq
3+YknOXYdr7pg16vbj3KkwIjh4OIPLHOMx/YeKqt/E24Cl5kMQcIq/cu5wf6xWX7j41QSVSuBHa8
5/2rxxBOb54VUkgLeh2u9GSWLVxVIE4/5O1lss/s3drSFtxLwWpbs6FkCdkPD2t/USXmA9nnk42y
PEmwoBkx4w6bH5NOEI4l+lYAzXmtIus8w130y9dfwHLQ2PQpcRQjPjvklePxEskMBcAAAYYPHgQr
0ANtQJMcGcEmeBKHoZt++Jfnb8tgZuodYBHeF57NkVkKHgt8jpv7yWiAB5CxVggaYid5fMy4Jm9N
LRc//jQwBatPX2Yclb5cwCMybL5H3dtkhpNU5jNjHovuMwlJzJyeskU7qmHsYMXjJyPoU9GvvjrL
rfiCTHrbEVQLcK4QMftoaMKLaNVoofBrL3qAqq8c/uetptk/toHW5/65BUQUIn/7KA2C1PNpGoSS
3jnXtrmdeZT7sowzHwUGIp+yPSYR7jK45W9M32/KjSZTke9+3w3APpGg+i/l6gziER6rzVfLClcx
/xGZBEk8frZa27NHDB4Ig56PrV04qXv/weG05uNePc3ngGMjAE7H7CXlbzd0Y+e38oOFsukl8ZMi
B1JEC+FZqzhAmZ+3l3/KMl2FDzgYczfgyHCADk8nmkr4Ilw7QtHend9Bama5tjJlh/DDPxKrqPL7
J43wf5l6H33K4lDSIp4QjSGAYsiY7YAfvtFfwe3usG/b26nZdSF0/3yRchAf6kLSABGSYaOm+Xhe
wbBuxb0GWOfch4Y2khp0Vt3emWozlYv/r5LV2l6NhQvVfBlyi0Lk7dI26E0ywr8iysWe+cpQflHH
QprbxuLNL/12BgujmqmdZuUneQQg0CkugFYcngKGLGbEmPb+zCjCCpHA+vmKQrlPvzoVEph0kIVo
TIdEbKzLQ9otufQ4ZVfuIcTq3yVyzmjSQQRmfbvsfUTjkwE2qKtezbDte92fnmtmkMP1L3esl/Fs
4jkJ0oCcCLdVURm9Gr0DJkAhtKXSQ7Biq6dF4lcbyGRMiW3EP/sCElBjPO4lINbN03fQD9IriX3b
bCPZknbuBiixTdTw87r8lUqSvnm1OsJskZEy1JmXHfswFWC/ZeZPGL4POtFr//FcC6PihvAk6TJa
PxCoNw+qeuBQ+C6Eg6xjCLdUBduC6gHEFLdf9JJtpKYrDcSgbfwkjMW+SgMwLFdJqq8pmY6pnhHJ
qAeh/K0M//FCpRVyqgUo+GAsawtgWKYsr4G2E+GzOXa6c75tprdYbdsTcn1IJlfzqoadXfj64Acl
56bnOMmBUAd5nksCkEOkcf5YhkF6EO4ViPWYLd3LiVtXTg404HzHWxkxXpvKLYxqah8QymIK+azb
g6IYPOB3lI2IN3K9mMn+b9nou4NgB2MrMTDM2tD18+N2+uoEuts3t31XiJID8maTmMkBvWi9ERVp
nAAY3YwJEmfUUg/ikZLlzPmhr0jTwdb9Y2K19mwO7otVyZE3k4gReia5w4MxjdM25QrL3Fz9lPZb
/BKGkVdgYQh6eSw3gvPg9KkEtWQ5cBZ7U1vGH8H/5wC8tbr0vmzcX+UJUFBrL2B23cfj90lmIVSI
j9OysQLQ7tWZD+ij4kGuB+53tugfPM7lH2u7/rgAfF0W/q5+htrSxOG26qaQgKM2VwiBpd4t9bfe
hWog0ARgFMoYaiSl5kHwJr1fyR3tEq1zB7vjoFnQwaRCWUZpnBGpm50aLwj+69W19TEWtrtovW/l
0gdG3ewO1IjAhL25AzLb23wMa/MuLs9rUi2mo91ZclcUxkL66kSQ1vMZsly1oPY2xhCBTC+UbvzD
VCpkMojNOziJ602KalPU+XYa1gEVRcaIDJ4iaS6TV8Het67NFaj6/tsZ0DW2gXy/vs8Q2wC/lUgY
p5pB/9oS5ILYOrgUFD6mAMiweEA2ZpOVEubLEdjINHFRpzmWHPx64uYD8Lx8oYRkh/B5HjFl6M8y
adzJ88iwHijOrwQ1LeLlA5zvJppXMvPlsYDeK/dj/eheBq1Vaj0ZFvU6nXlAFEtwMmAH/uwC9Q3j
djYz5yaIAj8CQf4JJi5LWAa0/L6kupmGdAHcMyg+FfnSBazF3JQjT/68mHdbx3OM645aPqlWji9M
X3cNhCA5ksdIOPLU9PlFEZwxviMBcq/pIN+n1uxR5I+AJwlYHZT7uJF+u04GptygL+HsVuIB+ubm
pgizaXvjXpfqJJEVQ0PE2PxCegJPl9ZKD+GCYvsjw7HeZ1qIEJYU/LYIyxaKAZkLdBdf4sWT4aZl
MD7uSyis07CnULei3oG5ZWT7XLIf1MWqLptoWgTs0erdnHDoC/1MKx5sAI4lbMOSwsvCAjhedGnn
JV2PDV01BNNGwcxhQ8jsM+MJWCjGy8FzrjwFz9o74q/KKDiQywdbKg6Mk3PX/pf1noI9B6qwSLEX
gtjSepLVAXElT/NfksOESumFrSn9mRY+kH3n3Oye1mnRAJA24dO0TR9K4ZofLlHctLvQXCBRxZUz
zkEWbX7d3fYO5yPWLQt1+EuEtE8Ep49Dx/YU+LE/d/FjCUyWQaSrDEfAqUOtgS6tetwFiAl8COUi
VqY2n0N+j6Rr7qnhXGqRR3CjDCgtU99hkTRLdpQ1u0FkejGaslyXoVmJ5+YlizT5XaHmrDQ4IPRb
CZ4mAxS61aFy5Uj65q6eY6+pUWppWR9gY0fh8zgw8MtGjCToMCI63d2FrrcWdUHoeDdA0cAZdN9l
O1pr2b+w738RQ5iNhJN03hsPX3mFve6l6oLF+PxPrV/Tta2pxHr874cf43MI6y+1h0ShAwE2CEtH
xjZkYIJXHAPdXgOTMagD5KeNFGou5M+y6kimScHqKyZjOPG6f2ur14Qd56N3KZnpFbNY7I1z87Ym
8RdOPMY8bVwDAytosM3brKOUJ0RGV16rxDMkWlwq3jbh8VH2dw967v9DZCTWwNdkz1m3x57kQETS
oo8wV0OrowV8rR9AYaIMT0NT4xxUufczB45hx4KX+eKGpz4y0/JE2Q3CmTgFaSTsvN9sCML54IHQ
p4HqGy1GjetDyGiqmBDoh6zyiEeVRrSON4yje1pNjP2SPwTw0/sEJVFiI8aA87jRl9g2MO6uC8UR
VACLoqglivMovwUYH8C0fIQ8Zuv4I1nRtRsxTMUh1gu/GJHfrWebII5SqVyjrU7xJMivCwUZw30h
96ad2LlKf6p6k9ta75jWVQzvI+4WAtmJXbbFCPQr1nBsDcsrKa29VQWW6lPCTEckccjGoyI+mnGX
qbyfnMQrSJxcigAtnImWuMFi1wQoyG6spTxlKF4FwPJ55BVtxSuwiV2LgDnWFHEz6658W6+lf5e7
uFR5s6TW/GGtd5RTKp2Kd4fyArp22e8VshwG2RAAP1rsbKU2DErgK7acsLgQH7DvG6K8r7jwMfCO
Y+SCrtI3lNs3hOn+Vs0Bxd+31ZxyBnDehmGlPMfx0chWViYUC7fuf5OlI5NbMkLPOD4Jv+KAGGsR
6oP5FUTl6OCME0Ozf9uZZtYRB+rKyud81jBeCvtITqvk8UJcsh4aRG/ZjTegmCJysAvUOtlj1Bzj
quSEQRj97ONm/u8EavID/MHVRpwcJwYjktNhAfV9gmK+/pTUwzbUQqt4/fUQ/73PnZ68z/oqJZwT
DHhaxzmr7Kjqa2lS67Rnz/t3zOCquDaZ4PNPEBgT+xwYkBGwAY0paGVCdGJJ4mBOmXWHIGVSIqNj
bF+iy8nONWGY30KIPFnVlrgTheglxg+7L7alLrUjGuyZg+9D6WLkO1js7eCHRNv4okCc+/syXg5I
29/9gnGNLWlL3FTL581BxcQLWQ4D3G88WYTClGf7cZnJ1bwkZqp0scvZ0AHSPDDLor5TEYqcqulh
vxGk3KwcdTB9OLSJzGVHvJ3qBF6Xjz7F/cP976+L+JUuYKHkO8jb678FqzVhNmqZO7/VS9xoXYTy
V18BI5YISRzAMGcJQUnt77iVcqkrYM3aCuguqbAI9UQ9wnJ4p6SUrSPk/DsgHm+/7Lc8KMkeYdTU
dzg+pwbVApw8Tn1KNLvyK0uyoDxuSUaXnAjItUunWIedEnpQtuG5PNbw1GPRDXxSAHC4uA1NFOHz
6AVp6wG1JZadUnMRrkUXgm4gJf4ukiEewEsODX+1iZGUZtarZFbiM5+C8Yc/JOcsxok4KvgFxlaH
KhOSAkyAvWCl8QbhhU9JvCk3h8N7csnnbeiqI8UfY2h7C+RrQC96edriFzDPvfASMpbpu1ETZ6iH
W7nhVChZX/eEQ52jCnxhJ8aOUERnTIm3X/VZa5pXCc60Eys7LdaYYOw3nDzucR2ctPV5jZ6AdLvu
fMYOS2lCA+fIvdVG5Brfo9X2bz5k17QyAhm1IvsknnbYQhCCTUbjobcYQUvCppqmJ2hIhPWLOSen
LJwn7yrN9RX3uoNmIak3nGa+AcF7CnJ0gOzD/uKEjZcLpaonjyJ2Lk7mH5W5+mlyoc0nmAWkbjTP
ls/fCjonb9ceUYpTEfvtI8bm/t1yVRXTTmlDfr0TP6aQx4ol1w0WhF1YLA66kCqifD/WhJfYHK2b
pYZ03Vv59IOJyGBxT/VKHLiGh+kphK1kuD5D4Rhnl+jZrAVoU7Jcj/S57bvnkio6/Fwx2zWKpLQb
07RgKKoxenYvbPyulLntuMh8BElsJwRoBr4VG5Zx+LsZolWZBW319pB1Ibqb04rBb2wwLVuoH9NN
hQ/j2cWLiNBfBL3REoqrorZW/F8ChJAW9TaWz26p7FpAD1prXkP+35SvCkygVgBaqnxMALkdDSWZ
wH7nbJJK3PiAcyvJWmSGQCW/wqyP2OBGXUsyCR4QqljGYbNU54fT78HHtRM0/Z5hlDOmE8ZDRW5u
mCrLVX4ruX4M0IqD1rCQP38MKIgFymNbZaosZOaTdh4cjVtyHlKyfyKhCPM7PNXQTeuiFRy4jHF5
GY+aTOMXufYDMsWzRQ8drdTbXTgR8wiek48eorBA8p4ZlrGa2n8YFelaZUf14uE71ewPlT7uqfZy
yNFz0Ich8YZ9xensdM2troLqKMGlh+xkVqcFoEdhVqH1hyrOH/5aHrofAdv1roViKljM2bAGIk+H
I7cM2lMAnoyCqeyDKlYSMA8PHFZhb4nowQ7jqU4HGKfp5BIbT2yFLGfaoLkrAjzUPW5l6G8YREPp
C/omVz5pTyGwZICP0Ia50o7DQgpWh22Y8OiEGX/OXVSyn8ZSPOAYO2cwuNRp3zGK5OvGaKvLSL+X
NuLY45kziV6aZcYssu1rrmpDOWJYpy/uGihH3K3usVEse1pkxcP+G+er+1zqgCAh+7V7bBVhfYrU
vYnY6GqaAmLsY9rl8Wp8ATLQjmAU6se2uonOMl5sxe0eW53LuSt8nbN+HAp8L1Ag4baNKJqNbBJZ
3iqeq+92iy526QhgBNCty0b982sgQvIzsjLwkLHVmOVBl6LBI7iLRjziVce4v+3DHj2+MrJQ7ddk
NUOf4k0LxKJSWh+jKVTSAUZ0tL9oILmHyax9+XDd4xHY8Dc8AyPzkUGl80f19wXjzOD1GdJgvVUq
DI/apUbf+xGNDyKevVIi36PLBRhRDeQZ5AjHF7DhjxfEZTunPR48OBNmEzruguvPiNT0sCYdklJO
91I7VXOUu+IbomSgl3U7Ilo1D5BGHLl6iexcrcEe5wLxD6/P71Q4cgP0SepwxcA7+lhordz3dRyO
7UnL9DPvsy9IMgECoRFuKgFXyv70nzuqaIeLbbo0p62tf6DcY2cDtk2bu7CThRrFRlgIXNIg1xQi
Q1QiuSngedZTJVAgbVLcAhDvVY3R7vVZIqdJ9CEF1/7rXWWwyv8tn/OVdvGlDxzg+GR/n4VAxlt3
m4Uj7JTzt8CJE3crqOJy/Hq+QV9k4+75sO12haUyH6Awsjy9jU788VioYgay3TIMtdfkOGHOuFyV
6G+Pv/7nJ4mOE/0Q6n5/SEnL25e46hJNpS0+UjSimY/GminAsWF6xb7CZPpeSyOKtNKIhv1UWY3G
AL5e2GnEooFtrofwQL1UKYTrEeJcROkiAn9cu5gs7C9sUPf2ojnZMWlgtj/QASHvZPft1t3fTldP
foDK2CsidEqCHwwwHL0LmfOo4OWojc/852eQatzqwmg+cmzBeFOGpefBg2BPIVpJMI87vqN2uuZs
N1Y1jdZWywcFEOyTV8K35WkLFYPLTo86f/qjogdJKCUEJ34iuxraklvHGqKOpzz19BDolvP5gGLc
JYkTW9DGbqOHmd6g5n522t//4TY5sRw53Sw7aBX0g8hCxDUJkcTBRvNAitCPzytpEtOI8RxdRcbc
yNzBuONsonemoCMvSmy1ZAbxP8YvkbiAR49nz7mCSEmSUjQjf8S8gGDZ90uLffEbyguVxjUmhHSf
b13Yo0z+L+uzLTVpViXrSg/XPVmIZtchRH++PsylZi1h5FWrcpaJDtPd9k0d4LY/5XXFea/+Np7i
8pb/BH6H9/bm7dZS7Atn2mxOTolh8ACWKuKNYHzkjD2brQI44xzBqXD1ofVYPjb+AiyGH9hkXvEu
goolIgjFL4jYl7CzCvqsrsejBSUAVWo0SwTMByS4pDwE3jtGVe4PRAC1O5gCPJTaVldSlVY/CE/a
UsmsFSn4/x+NX9EddELTuuqBHn4aZKuf1K2NFQtR2kPZTIDATj8CNEwZT+8FSResiwbmpBlqLx3D
L3DDAHpMqvPZ90dHlyX2qOPEXnbe9VNHlf+fN5iGfuUqZmGfwvcu/GNa5L+Z7a89xVDU8lcRODiu
dnXMPpIRhzOXeuLO4pdGK4qDcv6XsSfRWnBJt9WMwrDCV16DAR3SH8kZMwhwRjUu2wwXn5LxeHps
A+BjE1wmDVNSIW0asQ3jUl4Nkfl71GflcRhYlInAiOOa4XfNlD6DXIWiQJqgfZgkZPc2mpVxsr2k
bNb5eS0sHfUYKdjGtdQY6WkfwPcF9Kq3z0QdlbiOW7BUUzGoZ6F9dlYRHxbqdNWBIONbumKeJtQE
eHOaFkhesoQ0r61R+KDcV81oh9yAO7yrFWXAO/FEAgpy8m5ykcs5aCKbQ8xzIHY92Se3xzQxgPol
BY7XwrX7dy4SnStAyDtgDPuBwuEdFhvhsclowIqGOw4bv1ZRZ3ZsNayHhBBFrc3FD6kEB16j0mIh
5wE7kpiJPFXclvhGC42Od21CSlSVjGOa//CBPnp7GYSFbk4F8d2KZ7kKUmKmgjziLt0P9CioK46p
yHiLn+CUjYyVY5tfdT2K0alQl2KpOnymEuk+0h2gwuROLxtvtEuHvRzJaheACDj2LqPRHuq9lbv5
AXSZRXjFr6t03EmBk6mqVo+uWqSrGisasKtdwn4plZXDYHphOsPvZZZ+5sp+T8PjXC6nHJa9QQSu
3COjM+QuruSju2zdBMi15hoxTlJ6rTJk9n1zVkkmql9gdkyfGCZq6YaWzyNBzBdWgdAh7Yf67bHS
BMxUhEYf8G7Qp7gzKV9hBC7Y2n30/Hr0GYGnzoAws/9qTOdp2oOgcoXe162fBh6+Y4B6ltPEl3N2
vH3+Cjr72NWmH646RKLiuTvfjn6DUovvPBSlG0sEbGLWciWG1OT3th9y6ZiloMYqGJk00Fkk0NXU
GEwu0Ouk33btnhoWxUr7K7cImuMmq5pgI+1HK2Dye1DJIF+Lrak4Fa20YaGOz1xtvvzrks6boOEE
KGVcSSDKUITBw3rRf8rsgMrqzzDg/qhMEdE+igCIy1eTMvoeafPkFNu9lRYkoIEAv6wT5nbrBD3v
5qrlQwZon+eghJvPNoLOcHNE3M6ggX6W8rmWQcqo1qvQ7X4kqCM4s/n420DUKBUQAwMGafCSj/fe
Np2SpEkqoZ+gAvz1vdiRGQ0DDRBcSw9K0pksCO4LgbkM7/siL9rwBXN1AjqHvt1P3w5Q6w2IX8ms
1U6WBKGx0UBRoQ065GGq4W8A3S0+Jv29OFSom+ysOfS5I/yAdWOhzyhe1QJU7s1L0CGnaBsjNCds
ChSmI69jcTTOMRkfLib1Fwnj/UmGD0kVYpF25JNUo168zvpzITXb34JgITWj2xuK5M5Cdd4tMwVC
dhl4QfQf0Tg217oiVviXY1alAHs1+74KnxoAT1/b1RQOcu9t9ZBTRf2wO5V25886/eZW7MvfNJjJ
Y3/SIW9ka+kWTBJdLDDLklxd+d27nZgEKWulvlEWM+J43khJOETB4Cga79SAk99LzGOmNGrkmvqL
iv7DeQ7FthMcBdMt51wD3xidp14tRKMrFgKVZJNZb7Po9Yo+hSsKVneC014Fmpa4zepORwyq/07V
Wc4wyTuNNtdRkE7nGRFSOgJWx9DJvUppJCGs4BcDESmZkSPewUGajFo70AXeIFWhN51WjBS8EvbP
sxYQ+NbNwkjSl42pWgQlf2biENbbUpj0WhW9Z0Pz2poQyVmqcp9Cqe8amhCa+tclsF9283V1XYrx
qCR700vU2/7lExmuRW0Gfo3zG7FrZsk+FJthaJUm6kn9lQUEkPyxeaHEkC+UC2kOvjUC97wl6vtT
EgSjfT57FglEeM2V9oeYCz5C2MNha/nJb47ItyCQtamLhnj7BgPe5b4LHYpIM2NtDDB+Gpp4af+W
k2sdscA21nMIKhxsqMBB/zr6VRVj2QlTz3hDxvUKyvLBf40k5LbThSFfZgD6urkVHLj8Z1AMlLZr
0Siej/g5qYcaHkIXRxgA7KtP8EYj00chLHoudKMuvOmUSt2o65F8n6Ms2q4SnPoyJmeKmPHMR+wi
tjY8xKz/0yuSVdT6JgNYpVdSRjc2leTZy13pkA4QZi7t2zXB2PNIXKJ+XkvRflxVQiTXATeFhunz
2x620zwt3qeYZOpUyzvYClRASOybdLvTyP+CnulNV2KhZH3ChgG20g+JGjAL/OaILWmp3fyYmLwC
q3pvjiWmtvlqZTCc2QenUp8kmwVBbHeJjqSnfUZZfMbpBo/2USozDcpJBw+VwPMor+PfQsjJWuMv
p5x8KWE0XP/EfY8E7Fx5vpQzriFRvHV0mYh3YDjfWUFUePP756NbERDV58pvGj94QZC0SGo6LKkp
Z7wJuaqvHRGNzFO+YY0wkQzlTaNFtuWJ+gfrWNwBYjEI4279IQ8/I6J7qO5t55EY2qlbvkNyGpSR
t3xx1EMjMZbYfHncaSmO8XmsNTbh17S0lmdBOGKWR5LJlWhtxUe/g1okhYcn7m6tR8nFjSocHfTS
5acUJsnm7ljzSY7N55kE9b0aoiINOS6XPkzFZwZXucm3fjotWTk9Dbbxf3vFTwWhHF1fFZr9I63O
04jxTrZ3njRiWujD7+B80bQaVky3n0ZC0T/m9KVXZwHcrTDWbVrttWyPDK7dE/OzBaFT7IgiFIqH
MdAMiVfOTvsMw9gRl0vuURm5gqM6e4iNX9kiUBjdsm+xTuFbnJrBU9RbGbOnnIlG+9ufoXDdGdJn
cUkMmzrhDglsNKhNrBKTm9FT5ERR5DifVDiNyTmFnAWThkrn9vyDECMOrhPIxTAtl71+B3mpjb7k
V0p9ytrN8fzehs9GupjHc15+G8IivWmkJ8Z3KrXoRf22b+68uOpWPia+hWNpPn6qY+qxfkvAJfe6
UaRIt6mMJ2EfFqe27iJN7bdyn6uAWM13+JDQwp2Inovsq5JDEPaY8vydwEe7peXx6OIEb4QVHIQB
YNMpirdcW1xkP4mF5xYADRKXhRG/4IL4BGWNXo+sp0TTAsaDoAMazaDV6ffojsl9Z5XgxrmCJAlC
yqyI07xUbGDtttnNTso3WzkZJGjt8CpdERWXBZuVcWPNa94RAUzngyf/G3Y6idXMss/krhEHyExr
LCDZgCulqRUSVSWp7XT8aD8GrxK6a14ClapqrqaguHfLqt85e+c+ULmQ05PAIUEdPotv9PW3yn/U
I6TLnUvEZp/K3zT55MQ1ErxpIEP0GVqMDDgDxjxNaHUotLN0RuBh2Oa1mecp67TbObDo/tMjZkpc
IyafrzyBonsOGHA1uJn2UhCIpqxtMhKbumL9pvJsFdkYh/d2P8dwRd5cvQJZFxS0O6YqVAa73ELa
mSbU8QKzwrFYM2ukZQ8p0ZxpFZXQdDql2fUWFzmGImTGCF2MX6g8mpfV+MUwOdA9zZXj8ldqqDSd
tq9J7EC2goAlDHqzQsnyXabfX0z/HIzAEI9xjjDubIMuonWOWi5F4oUWbFhWeOpUCbNDO+lULBMa
pkHtQQT8STr/KLrYjRdWkqANTMylmCK8pXtxFgrL2BKB3GHV031V3q8ayoQrw+UhAVEBTJS7omsB
8TP144viFCg2vYuBo2endWJ0R8ydYYFtM7Vu99YNhx/F7/vUR8mP/HJMmFz9JeC71ZWkXkERKByr
xsY/bFA2Yq8QdLseIfoUi0hL+OKctX5AGkWCOGa1/0i+YmXacjJqBZL4HSu+GVh+8UdlDR+dzQHh
X6yH8Vi0xivPTNnb1FtrR+ubeeVcbZTTnI3Ekc4oFZzxSdyL1is31XGj6P/OX3KAC1tbV0p7f5ig
BzH44vlTPAujdf7tukWgOJxlgX4skJZgqm4h6vGZeG4IKley5Kn8ICMTriIaW5qA2KibdkDGWg2m
WCaE1udHNPXxS7/tYD0mTndPY0Zpf4zPFipFd7onaYZWl0E9Ogo+IgXQdDOi7OFeEMeLT7ReFUN/
flVtVAAydhClHdzIz/c1BkLNlYbKs8kyDOrAMtQMkoc4Y3pGmSuVFpwaRoNCT+WJNZYTqvHUmc7X
0azLXwF1BUFNomx1chnKi9hU31w0jhOs3Uae8Ru2Ujxbtvgr9pXcJa7rsvXltu/Tc9SnV/7bHhcn
rsbtC8sQp0v/7CrDPl82O+rrtkS+upSS8lr1yduAEqJz1jYQ+EUfU/nl82W09HRI6rDZudAKGJBg
FZkEQzAoSXTkV/xv0bNXW8DvECUpjX1bvW62mT66j46etpgpPQtzXGImR0hTTVbimsuBUsUaJcaZ
bqbpefinMhwhc2/Bql0EmiXf+ToB/It0d0hdQYosyZ6X16vG79NMYLh3p7b51ribCZSedwZhUPDu
tlZ8jAy/6C2LuSac2ecE5dENqmM83L4xj/6gzIP5MkwhyYSBD4vCojw4i7xp98/NYRc/S5K1rrLt
qbci5V/KKq0Vw3ZZWOEKtshVgUw8webv0TqzbhtD2xk1VXI0l5Nj9lYUXUZs/kpylSL82hE5zkO5
QaIeNs6nyT11o01fy+JL+0Mx6DSlwhMzuoReioMbLhkU0VLLFVT2y/G8qPwJy89P5a9HnK8fkjTl
hE2Fo4jOeSpZ/9ZpECadbjDWH7pybOTLTOrFrBuZ1kZsK1w6WA1ToPSL6pYMJmej3/DR9TrZYwja
StJMp9Yzpdlg5dVe8uB1bUU2YXPJfvEBkm7F4GBh94XDiX2RRG1aJYfYQBh/5kUn+rvenUJY6LOx
qdUgIBu3X6rlpFnRZcVBPOWNlSm0nrtflPNI5tHsq6LT7Xbl79Wyip2Q1xmdsFNk7IBwpzfxUFXd
JDA+bUUWcBLLRZPgpH1QmWPFc1+5BpS/TARat2LNQKIIL1bg/C6VdZabDHa0o77CGQitCh1DQnd7
IGU/n2kNzBWHlvBxQM+hh9skYjUdav5m6sGWjGP01tA9b34qiwZPAWkA/D2qEdvGqCB7KDj2zn4P
MwwQIJZS6frgOQhhJmN1zdoPilMJXN0TF67NzIphSaBdAau7Gl1O0Fsbupc5uoEihvFCyG5g1Wqe
pYyE2MWSfMo8qYqHCsUHAUSxtoJPG3b599l/Zmd5ITnFHFR67KPdFj+joBv+K9Aa50+P4ZlBNl7G
G01553xlT+1XUzT31ilqjmkJHKrYXRX/d3DMz5kwbutDTO4U1BmYGpu9wFu7tGDwrTn3YRj4PKTu
QG4mOwD4KMlEcKiqf47laZP+iRAK4jwf/wXNWVFCSid9osihB79mwJjhFBv9YTCxQKJnm9lhSfLp
LQ4FJxHfOW/h5vU334T9O8wT+mRN/B9K9FWD+TLEheC07y57NFN3Off+yTPtjYM3BCD3rklZpPol
/FVC/ZOV3g/r9xTDakxbYy1ReL6DDYuxKBgZZy/53ihf6vEJVYWM4V5bZ5G4FYWI6iEDuqxxQSKh
RFWJbXxrHp8P37srKMKZwvLjvDWeE17lEpNLosAAUxd/KS0Sn1uEhYJLYCtgZjkZtwjO4vXvBvgA
KRk5ggZZ7OSHPcm2kVABW9vRSUEQn73OY+dWm79ErLDctv+HPVwnm1C5q14E+hNollrb7gVwlFgS
ehcgqu8I1u8IODY381NpQrTnA3wjfecMmQrcOr9MvKEayKE3kemnRgTUixfGcatMf0KqHHRWLFuJ
oeqEzp+BcGv+T0/9BoGicoezNyYbB06ru+Krciy0l/tUa0k0s8eajdjd8WEKLnwSm0CyWwJRiOKM
J+aj6pxaKL8sswHqF7La3TYJRSsYCVv9IOb2As3GE8+qgVZ7kDrpCgZbQqeo9R9IvqFBHUs+uhO5
rFOaRggWqQ75sy8qI5AMcsI+K3xMju642lmKe7zZ88g2njfog8IzNY1h1Z2A8wuNcbfpttpIl+0t
IkN2T4lo3ZuwZcAa3drbMLJIZkktgs+hlTFTPXFtD/yFbxowQK2lEzojFCu0KYsaIhK/BR2UJB4C
puFqY9/8QQaaEs2ld70iO22eqbkro6CpPUFkPD6jEkkAgK5/pR3IClXTpDCRmTs/TQSn1dZkFRrt
3+ZNm9lSC74aNnmh0+Z5qIsRoKDg3wcaCtghd4bMYjuRMSXN5ku5uwegbzvRUbwz+G9+eUbsFKtS
Mqui429UYAJXG6F9bZWPZR3+av0/mmSgmtOdcYefE+IMVbnIuQzP0GKIPxJGJPMWb+SYsreqWB3z
tRYpkQMavvlqbzurFgLDY1FHoTFqJx8zVllH2sZowUpgtlKf4NRMnCgeM8HxVYBYH5GFe/EWEsCN
2eA2NfJn8qUA7dom+DzCbOwEuJ5icoHDp6LlykSjhmcD0IOXNy/wIxPgioYI3uKNAPsNjRXbdWjz
zS5V2QOS3aqepFeBv1tWHNOMWazJSyAdly5l/2IV8AJAmY1yGOhrKputT8EtoyAfBfwfS2vdyYPC
5icaWBwARsEfteSK5M/7HBp3BmBkLMPrSiaHc1vb1AfBGJdo6G9ygDRNBLzZC6dwvOOe1XkChK9M
oecA70FVV4zZGQwhiVwLK37mbPFSoTyz3Jbn/bscFdcKzeypK+oyqYVGVTNZJ3N5at+66VtY+jU8
PE0ENvb//6mmR4zcBuaufR0lYGhIKtSo4f3Tj0cG6FNRerI59mvl8kgwkzXGZiYoFsSQ4jYLCrrE
6Sb7IJ7hc7+n8yVSQXKgexWhohLak0ejLyL3KtHZZOSlkS5yseAfg3yOfWJHovF2/jb5yVwnMjgc
RhhwfMzqgVbCm/8I/wHlQqoHcMLa4roGT6WIgenx6FPoHeAC+Ts4/z45QfmKizN762+upGaRxvU1
6kRto5X9uHWGv0eeLIZ9DJXx4/8MUGr7hXx1YhDQQZzJucp+1FFYcaRb/BpCw763ISe185YkdPkV
hYxk1Q5Q4IbEkqUv5KdqDba774g50ZGO54Q9PCuzd6jIa2KcPsSbFPrgeJWXPkQoW8kEPU5wRilB
BcSqy9XNO1IHQWcfHNQYGFQ52DvAxoPVetrrZhNyfXGi2Jh5ulUAX8R37htuvTn5oaEfGg/9uOUh
UqPUEz08/59EtMYPgAZE6n+Me/6Dc7GnehfC6v5lOSkA72oahDcgEa1Mv1WQVoMKzNgj7T+hjmJu
mMkXnDECvVuHPZJC1tXg2iEqVWGqOJvwg9JmBUHNL6U26JPZxgMAPwqagX+iflz/HbbAkkGnHIhS
kcPwEYCAKECM7oZ5Up6nUEahgJaBNx1RV6J7bxVJRZr+PMY0Js/uovm+461KtE3+EaXM+8g/yMIx
dSeKDF6zEFYp6E2DudG74DAxgC8SuGiL1x3+0ix7NnaNMqK4cw9WA7snh0Mt+fCACvZMKqMLpftw
eKHgoNj+vi2APHAcJN2R94thEQAQPa9Zakqy4X89nryTB7fsKFBvFhejQXyvFjjL7vyRxBRf49fj
kiccb8WBY38i3wPvv4RzQaxMyBhYDPbsBpJ9N/GP5NpoEXmYkojCRhCYolr+gz6OAUgW5Bw+RH5n
YP1Onxdnwdcnx9+701PUQmZ04tq9GxuExW+1+e9vf4gxZByd5qDj/9OWrJx4ku1uNOap9PhJh1aA
3wRgmmzTr6gr6+dtYcNpfeOQsjokO0HIex7ggreD8imVMCKuDgCzLuJZhto4Zmoy+kGAJpOEIots
r72SHLH2yqPWMIyIfjKXBZ/wbMuu9Vr9gh/0hjpZ/kT1kToTgwXzMGt7AAV4pRK1wabQbnUZLVMT
8a/bt0+W/inBMtv+77QFi2XzjX/Xa+RObliUgfiFtCLuMdFt8rAqU2GdjdtjDF1pelxG1MYkWCeb
4jHSlnBTPQ7h87mxgDyKUAnQ6oK/gsUCK3tSbArSR9Xu5KEulhAUfhmqs5fuAOK2elkAQg5ggVk1
BsUqi12TyRRG9BCOMgGfT9gfpY7Zp7/Ckb7bcpmewkOF8yc7RAixx+yGdULu1z6uO6sESxosrccR
ITSbLvmRIgITzm6V5qRXPdRQyoY+dEQulbF5L1S5SOLo3x+8hfF+Yh7SqmlfNP3jZmT9YLeDVECr
Whj4hiKjz7kbAHDiD1IoJFwBdZ1PYCtdMzX4mlAiLbpWZKsOoih9s5AOMjZ2gm0uWI8M4oShlCXq
/Lyehqs2Ee6EvYeyYPznKnBH4eERBXSKqbhqVuLRz7S/B1xZjdjK2zZl+Z7l3gDY4SHQoIiHjTSW
rwbEbPL7fgjROs0ESp4phoo6k/suu6TgznliG1oAsGswHuLwzO+U3G2eivHL5XQsOrK4eRJMyYhg
jA54Qi/udnS+pzKGCqNelYIoYp4jiJtZz2v/c0LH13SLEpuqhVcdMpVIcWGS4J3x43Df7zPZ2E1o
bfiIGKaiqVobTU3g7yd2kggYAhLP0518UnkSDTJDf4nPULJUv+wiItyiCoiiUwtQjfY2dnASdBfu
raeKLJMoyTJr7sM8QTLvHzUPBR+lP3rBvRBmW8f22sxJmePc7KrmNjzaEc3E++V7kLtzq5+i1Fsh
nAd9LAPpAsD+mCxd6THPI9ViQD2mbbwv8/KM5okCuZsp380qZ42y19ImBVVnLUOnUOcLlxihmJGw
RUrA97uTJeUxlIASkqbf0LztP9Ak/YuKVUdooLeZ2b62pgBZ9S3fyvNLrV65jBM4MVhzNCDjLDDU
bHGzd2emYOmO5M7j+XV+MyfszO2edCMjoVi9Io6gNAWe+NIU2iKL0dasnVamnEPOk/EddERslCIy
dcY9EfdH/sKnuqg+TAlQUYwiDpUnF78cW6swJTusUzxVRfCyh0naT+fjaVx9LGP+p3YT1mQ+UZXF
kCecgYV8GPqboamLtEApzRFW2nXFQem7L7sRichc2h4KCoz+8LRUWY40vlF1ZULfhhMyuEob0IW1
9tY8O1QhC+qeZD6C5nmR0AO/isNerFTowqws+J2+3PS6YJjkDEeoDdx4y2LFv+SvzDBicvs9dECj
Y5ywlY9KUbPRNVc+xtQ88BMOY9C9tHU2hH4zKNsFhykQl0ZpRJ1oJ7zsQFnDco5rtdgET7j9WXK7
PeOmzJX0jpVdJLhA02B0grxmq1mO9EOcPFJEY8/hUG7wO85JGRuiGSBUN2fdTd7XTm1Ckvok3LgF
p/MARjlVuPv1YQIkUZrit2OXmm4h2aUTmTddRqJAieC+J+4b/FyKNVCIKHicH6no9m5N9m5syrRu
fq2Es+1gffxOW46wEtPGoTc8unUZMmjFgiCASYVCWTreWViK9vFMVQeaZfUnIW1nPMeiH5AkvSp0
z89UbkudfsZIC5Vmnv6/K62SJuUk3GM4n8eIVZ0iEEswqOl+eeC3Yd7uki5w4JuLuym153L03bVc
wWACLc1ou2nQtU+kYAUAssTlfw9CPy3dnXW6dsRnp8O+oChufCaThfNWi7k1dDa4DFQx0kYfvr91
OBIumFqXCyhrfS+vHoH+fziP2Kvg96fRH/Irpo+xyI+QGa9q5ne+FYQCPZ79n1snUc7BETIq4kLU
Dsaex3p39ejubfIK5AzP3nUPszrT5YHqLOxOfTxcbW8XQ+Vna3jGyeDsLIzj7My7qcOV/2KeFc03
X7S8fs2N+z3vPv4mYO7XPK3EVPOsbW9vPqo60CnyoWO5NkhrPfZXHRTVwVvC/wr7xABFZlRWP66S
5DGk4qBMvru6hI0jFD13d2NfXGXy8y62Qggjs7jkhvIvWQQRwAuGuj6rUsWRMrj/MiSKR3yFTiSG
AuZI1In9oxGVf9JgpVOyxD++UmVycXZtH8bOmWpFipScfk5fEsMPKmKY8J/fsIPIKNpbsBSlX5BY
d7UJyxfhhyDMrLZJfSk4WNwOCJy1yZxI5wu9ZXY+vY88/+teQ21xKgufjQS9VFoq6Xc75za8uubT
C/HDUjR/8ngc7/sov+ayxow5d+RgUre46g3dff4JRBR5yXotoCGVDOjAKW3PSB/9ysbaD5Y+uoIc
pKG7F/CWivSIXtiHibNuelxtUJnjwP0IfRULOshB/j6me0GRGs6rylF3+yMAJKTsrISNHkPFvAMj
d+A873qax1FgKih1A+kOekSK6afvN6cAMfIMc8v5fevOpWV8Aeqps4Gy1BnDmrtasjRpXT64fg5k
ipQCe9x39ad019ez+4XbQj9UXqJgXVwbAaJYhLSt8qXL1wMA14eAUXObhayRgBA0X/wubeuJhDTX
xyVIwNTfcnnPv5MKTkNZhDnEyny755YkXcBEGIAhBz4f5gyYsEOkHrjcPZzLje8ow/A61WcHoAJV
v3vkmzLFEjNQcszV8ugzy5J+u/AEJlnwIRqkzlvhK2hyCUlRIaTcogQ81f/inKevPlKfG2pTLsr4
zVLp18fh7uiv3zaIiGa1n2HL6uz0bmW7FJwMmBQn9CEsC4VfL7GXjAB2N6dD8xOpCWGOU5GCZrgr
OktFPoIFX1LnLUBrIgwvLBdNXrqeS8QYvQgoAamdf6RRpCSTaBAX8A7M1IbfhQfylRmgPSvULD2K
YghTjFahQSTGSxxPbGctOIKI6dB9F6A6KCSTslHkG+syIHQ9W4iOJSIKDTlHh13UxFxThzypUK/a
nhNaIlacekO5E16zWv2bCC+KNgyD06HEIKGlhRzbVXit1VqzvhWmI/QBeDGkVhMYmZeoJ+n6S6q6
lqY28EyNwkE51d00vmNSKsEvWNnrEg2VNYjl+nwtA1BZzBsOEw8cAFvK2uALdOT6AgO4bmnAVD/L
0cWs9jz/pI0cXnMlXCtWHMogtTmgtfvpfhI1j3rBpUewUVylT9mhUYvDH6krN76bgnk/+SDSlN4P
vjqDjnNNclRFlNQ6L480vqsekm67Z4/DsR5DOUfzrOioOacGSMjQRBq5QXzjSES803xVyXeL+H6k
ZtGU445ViV5PKelgOgOpMxkzZ2tt95qXdLYPLTxIsd+aGgXh4ISPJ9XLIdyk272Gmm0tN5JJdSZ6
Wk9OCPcrPc/TDsQOGYTu971VHdEc7gZWo0hITbmNRuJSnrwPvRTYlcic593dQXTtOO5GU3YoEFcg
hoev5lO1c4zEVoW1DnoL2UhX3NEXNjZN4nuElYMR6jHdRGGRtNktB6t2YDBiH/ctr8dLHULw3Uu2
m6qsv2AQ85/pmUUS0H2psmNHV2ua/cqnbjD8jSV8fLmTolmWhKfQXv1oXg90S6/rh/3hTBYq48ud
7w7NEuEZ083FRSsbywHVmzOqzLO6KZXOJwbFTIl++seDgDjWzhASfVfaXVidgsaejyfRTSvxwUFJ
8AQ+d7vs6XruwIr9MJEA8Y4vAgoQGj/gtcbpSJ9apBoGfBBV++AZv7OIXJX7G/QhqgNPjRl/nor2
4qxTjr7TOQRzalvFBc1XPP/w6t2gyM2ljt+EinDtp9+Hf8ZN5g19E5JrLOHKlLGqSzto3PiQT9x2
mdHBmoaBVNA+l9aIh0O7ERsWduqeU4RtUA6UcA/h/KW2pLo2/3g9Zn6mi/5527bAFOIC6wUM1w5P
3LS1CXpEVwoH9zF+2WO01BboD7P70LULpJTT4+9qPZ/MXEwmt4T+bOkfc39bKJdkRJIZYQUCes/G
f9jumQ4xzkxgFwXdhztqk/BEc92jgKGEWX1pXWbx8dk2vXsb0V/oRLYL4Q2URS4qnLEHTyIY1Dai
JbGKLGSYQo3urkUMdJCa39sH8wsMk0Y8lMCbJofXniGxqbDfyuhTffficmPdow+yehsLVT3P8Gso
d7+3haWbTmGuo2fAi10+3GnujQLn17fqSzFBQTFAHO8FgdWQo2BPB7dAIh53cljq+tEcMcFpNraO
7RVaCet4Gmzigo5wp9X2evinyLvN1ZywEHmi3n4q23kko+UNJhUSn/mJScA2h7a466g6UOyiSU/7
M+9eQSrmLn+R1SC7Q7EFsqIcOpsjla11t9AJ/M70d9Yac093AHnILDmrvF9/RMH8CnhIfAFe3P9f
aqG9Nc7OA0bvawf+7QmWEK0F3cu/7bXNuxdso7KMAWp9tPbqtnbu9GP5bIsFbLju2WyEkcZE4pMl
bMa00gfbJEW5GBJlz4fkVDABPeGTnXGWtZK2jufxl9j0567GOrT9KeY6k1Khl59BfMAn5zXIeCnc
QVRfG+DCQlg6l1JNdEhaxcQU8HRwTGrcF+KFDC/cQ1CrnuiI6LnweWV400BurWYk+u2GeD+/wUPd
2TjEldex1PO/9m0wtDdAAZ4Jhtzdy22OkoEEfkVnCCpFYILttMIeYyRb8kf3SYRYt7TY+mRUgBLw
1ZVf2nkrDpVz8SiOTQCZTRAv0aGQgLbFtyx9CtynphxAjnWL3uihcr5Po8V6EOkyst0RhGK8/2Wv
PVdDEnaRtCEDSzULcXJYr6POph/G5dvNqTpe4FhK6d1qNdvffpLS/sRPSj6nUkGG5xC4VtSTfdb6
GZtCXSwxeZqav+CJTqAHQRbjjR+XxmBVzmWFOMBmxHJ9ssxUOjSpFj63x9AFBzWgJgkuEWOUk3Hy
FJaxgwNO7A9O5YaZd6szsaifI00je/4WDI2s37YBKaFYXaT5wBkcYbcXJ5COJLXD7jNjKTGoW/Fh
pGNTI/vDs/CpSuXFC4pV24FMmBtHyxAD66cmRIojkzV9NKA8MnHjo5A7VjUAwcfx2KsHT1DalNz1
tPyykNXcda7Mbalmt1DnIFBzAOE4hSpE5I5Y6TIEJIibnWFflduQfRpjGlKmwfvMwwhxWzxF583O
18ZyZNA2vHAR1Kl6FLOr9x0CMtKm3/hGg9r5LdfwmuzTxQpGtprP6RqHCfpsm5GK0JF4Sp5yMCup
F3tpSJZ8POjNU7BYhmVXIf8kaTmreEbeuD/MHhh596wsyXbTNPBDvxH/K8R0A5DabQ6WfDoiy1ov
HiA57Ejr0O3imt42sKgkzTflPTHDWC2bB3WcZv/yOnOB4baaAK/8VaADUdnJTe7wH3u4yXhtgG/9
G5BjsatqvWghp6clHE+GZYGDOldyuzded2m6KBwK8QCWZaBMsy986NGVTXbLlL/MaMASuDYJO0iX
kt3ISDRvCCZUalgfqohSVnkthYNpfONMFA9RAPjuZJdOPX686rudv24IZzQRWncsIzvkg3RcRJsW
GiUtogI1knJwvnemf/QRGlpp29TRaZzFZHjL4JC/ECitRUZ5Nw4icMlS737fXpmg7hQosyZFXHDD
i+aDeYWP3b4PLs56fd+9nF61yw+3Y0bQ3P+sA16ij9QQnrzUDl/Tel73m1ryI0J+/A4KPc8jF2Uz
Vl1znxBjq3kuQISHBmzOoElg8cnF449VLEoKh5gCarA5/Fj212ep0KeFX00muJA0OWiA6FUPtytZ
kxv3O7fF8rxajwAt2ET9uVEGHqDCaTLCVKhwTrNa4MYeU6OQo++hDeRngKhJLSP8xxPmPudMp0jd
pJQ3mJ201wjwDp48O9sB5Wr4BO4ZPC4DjdO9BBPIhTwQJ8QZHq1g7GVLbjMJQQtRf0nw6VHMCQne
JU1wkuH2Y98/laWGYMeAhRDD7j/xeHoaii0eCuRnMvA362uULGjCkx988a/lHojve5m5lflrL0kr
P00p+68Kb6miSMW/7E/lpZNb+d2AnN8TpB41Doy2gwqQRm9u2IsGVqPUcQ0JmI3u8CguSj2Qxn47
1W2wuqtBfpV0LN9vj9ou10gB6a0lilaqCmYg16KaxcQwJ6yUM8pWRCnnxxa7XPFJURCx3dizZS9S
MCVTbjoRh0ZzJWu4K5Y/1XIs1dcbLEGpjmByLT//h8NdmjFy5BLdxP8L67y7agSIahosyfI3s5E7
uU1rv9UWwyVnJV2gpbhBt8UX9+MiXthilnrAoAwbMXM53FD/GwHKQC7/0gc8tV/7V7CZQcfIx31v
nac90WgYzRUYbZ4BS8Ksf3bpv3do9utwHK+3PXWKqzXY+6yGB6vBibmO3aG5EXnGhvYAxJSL6liJ
uYcKGRsc9d9F5QXlrMwLd3mQcOVN9pzD2i4BEaX9HwLuRP0fyB9YenLNYdKJrGEjBsZoHCIp8Zd4
An3BUWvWHQ2dYxQ/iU5jxiyQhsLTmhtrXqvbLzk/zw0F3hrpD/dQDIR1/LEMqQcHxsE6aJY61Cdr
CLjF19vADCxStG3eLrUwXqoK90KF09EIWQnMxw39dxR8PRWQglgOLgeBfz1X30lCmK3ilrqnnseU
1+odNllxA6ayujC+EbMxCnW1zQk1uTbMZ83M4m86bpHKEVLaLEjI2SwKHvrA35ohLJbRtqOAnxWZ
lo20TlzY479mD9wF+6RdpE5EVyKeYCEv6sV5B6KtNAzaIDuIosRBTDOPHaysDJOX4/rLjlfnaF6U
aqt+q33JcLo6Dq7GPAVGI2AGNCKR6Xt5q0T6k4gb0OEZYfB+WM66FVG3/xMvkFARt4RWksrXPtny
R7rWJU8yfuco7jepKUGXfxbxWPAw5FHj6PSLeSrfAD42Co+8KMoIOCxAY6QB6loJ93IJKRBJ6pdr
27eZLUWxkkTB4911e+WdP0E5bhasMfZdN6/GQFJujKDSHdmDPH4R8E2aLd9aZUQ6rF1JvOHmMC8h
EPbWa3Epo3Q6aE6/zfDKc5gXCeO13oZTI3dTet+spHJxg8aqad/AcAlt6gYTkSntcXVMtKSKmobJ
WVCztSjQRvMh7rZUh5nDDKWgBgKaLtvovLvMOXSCwHoKVtDVc6tBubLz/vBhHRzc66SwNPGAKrxW
nzFjrkEj6Cz0z4JBoj0FOOnnmph1nrYL5nXV946wQttnaWLw6nnK7pI7pymPgljIZW0JhtFLO3zX
3cVOAiIEUjpHV8LVT6ebGlnh0pA1HgbCfbgSmpukZOE/12b08Xh1p4d1tT1/VDAONcIhrp+C+Rl3
E5jtvKqD7Cx0+DgQv6roZKAi5oBgs963Ra9fjzrCiAcLeDiRDTFX/PTnvVKX2EiU322U/IfOkyTm
ZI1oGhiOdvnYuGjFVjtJO/aHA4PXaFam+2CUqb5fMh1oUlUt9fRy02+u2eo33kXokTwGvZULvbIk
Z8P7f/AeaLHCLfpFMLZGRcshd4dfW/SDmmBgXAjfWVzLp2l2uCXL2hRujLRF3pnecgy5I4kZU9Q0
F04s4fYdLr+gW/bzT0Kt2hMhP9ri3po4t6+7G0jSDxGg0mB8rz37d0cjGIubJT6d2F8CZG9VxPLG
wCV37B0Ns4Uod7LdtJ1pp5xgg4XX5nAJt3ZeHYowNhP92FBI5udhOXqx6eIY3wu8Y0TvBvN0p0Jq
028eOrDEH1J8OoSWS1k1Brp+o/nepWZI8bpu0r3oW11ptNhhgE2N053oxN/3J4qaYW397LBr+6zu
4EX/cMgKWT3iZI4PkRURzWGT1T2obGddXrsvjwL+7J1eZQJfu3LYo526DeT5PMJKt/LSLzL2EEZT
y0p/q/bhQKDTt3hXIwPdEZ4q9HQ/zQowkZBep8Txp88Fg+MxhbopHwoLNq/Vk+57bL5QvLdEfzxb
HpIAxsRvKCPf7fpwJHI8yGMJhjOtP9GJvsDT3tsIRLfPB/MuQIxiaa/LIhAZ6rK88zK80spFlu4+
GLaSQLK9L3PvRE7iJ98XnMwiPsBD0K0y9cdS2f+WmywT3blu/OU0CbMunV5nF5YJWVFLE37a0oZc
jUZAOlmZn7KPOa1s1u80q57XsHIrPHHnA3NZj44a6PmxoQDCcuFm51TaryPV4Bm7DhS59sKA7dC4
LutP+r2Hm1sTJuxILDv9AxhtnJRn4H7kGn8Uv2I0Y7+9fWG+y/D3qha/LSStQwCkth65BIGTWQI3
Wa78vzObIjF4eJe2VBoS47dmQUgnLh7H04S9hmGS5o9Bf75AugQhu3PkLjHSgSpL++ruZqLxpSRI
JBrULo9l6kHb+JuHOzyB8pzYjpxp2ZCS1D7R4TnyOI3kR9chxg5OnueCLGArIIZ2NChWOBvVs5Tj
nNP7sI6M53258bslJU/EmhCSdn7d8XmAelo4+uXPq4bkC9zuQPx7QrGISORKkAEkDtdHzKUwi5nZ
g7Kefq9f0ANjU7B+4C18U3SKu/CnxMXCZURRZMH7x5pxRUUjtnuRFoYoBr4Ona9iobvTxkvIMVD/
CimKB3GpvsdqqEpN+2zG5vHtzf+d5Oa3sz2WMvTmf+yxt+Yzo22lE1143ArnVPB85Chy9yw4Y/Ks
CMpocEy2VJs2GYDMfM5lux7JZ/OIp2zfiLAW9oAiomJd54GIMaD/13yA930PbKSFKH/hgXfVMoxs
VfIt/9IupOsGOzpSHunpeTtc7qQ6Sj7qOE3wnnZKNjFYVe1nrGWT7w9aWFHUs86SfIFUkigP3PKS
djyKKuL582L53UcE5DkLu5OlL5sV4C1YfAM9cpf/R4voTx8XqyLPdTrV/a2QkYYbZlx2FZ4R/dL3
Qo1C9jleRJflBT2zE4xM3oPjDhAkLjcCh2pbKG6jgq8Zycj6JWYn3hSP7DABUuuuF0V6iYrwCq1K
VLWhy3yYZ0JbNXgCtrXAkh9uQ1RNWSFjj5WDL6G/UJmgN9TxH5PPumxPBCrE4d+dBsB28TyEwDix
MP2979bh1sE4TKFAfKsG3dcBY7sqr3QcPIvlBWHUPmsrd/7KjKyONibox5V2cRP1T9a2f/2eFYi4
FUJnLc1S+WXMLFMbHZ+kx1eBM9iX9sSSPGfkKU8gaAPe5W8kUwWjmX7UkuXb8j0mgw/kW/oirM0u
1d4SZrY7Y1HhKDlcQFiIv7yViHigCouPeX+rUv8HL3KpG/qhN2Qj+k+rVp9ZBcM6jrPLCA77PE22
EIubKwLGcmlHKjyxmaUQo8U+NoGPK2+Cz2yRL8bTFtTHRTbPjZy9X2HfTltLvkD2J+6ONS7w0xs4
2B9l+D8mD9jfDoO2FVxXd4vcVzxXvF8vUc1dIcT03W6c2M45iIhrABS2aW3/XH6io0mMagY+C0Ka
Kk2+z1WoSZtdoMQejXHJxuhdldwrWPlmyjkgw5qa1kM1gUR1/Ak+ZQHUxm4oAUUE7dqnWWwPExn/
SWVf//okFhxgXj368syqmWrVYtcfDxGnpbyZFZvD4c4SdQ/Rw8qC8RBRpXG2WwvT7lt2s3j3dCui
F22Oy27SdAb6ktR9HbbOR9YZQABV51j2q7c8E3mOW+hlFfSzW4Zq8/inxLfcnvEYuJmpitF8AtpI
BG9hFVG44jKs0xkAGbtY2FvBwp+fptoNZiBdGoROMISecnM4GnGNeQuR1q9AK/MffxTdrJ2NbyWn
pXnAMeDxjm77ENwgxJoGaovv0+612CMj15o7u0RsWwhCbpJU34HYpEPJktzoU6nkoQKEBWJ5OjH9
kENy6ttTtJp/rfeSMt/7GWfukfAdX7xDnqVDMaMP0/F85iAxDvPFeldjAx+r1WiQHarj3t5wuiz/
OgNIvGYAijoEMPPL1SIc1jHr0XNOUReEtdL07Am+RhV3Ccs4VXGha2mPbR+8K+nmqSct4QSuqrSd
GezQ/wvD8LohzniZfUn0FpBsKHr/koNODVAyjVgBbg4o8+vM/OPysgpem6Qp6AmSKCjPRUIkTD3S
vkAnLCqhU6whKpwoGU5UFFze/8wCMidVUyv7Tov4xTHX5OAtrnbAVlLuomKhvCe3toKT2JYzGYza
4kNMCk+CDOlylboxD+Ssy1W54FgHIjEhLLTOV/8zo22CDzwhYntoIa5GCcTP1bJHGMGjdXVmjffw
rq1/nHGcoEM1RdwFT9NHc38ebxSr3lBqKsnwU3rY9Ar+9SDE7XQZZ+5XD2+/y6ukpvFVHXqDt7Re
fD36rKWMKU33lBRwIyfbIYawIELtsOe3HvONDCQxztV0cSgXf3BDRUp1g93ut5lXsuRhCZ89RmTQ
YvPEE3o8zj9GyOhRG2g3bc8CWDEqVZFfjz6RUSZFgup8YDQa6gTyEr+j8OrMyDFmq5QD66Vi7Rqi
txqxepdk8c5l6YPAEZ6+b/E15TX5RZEBUDlEwsXH8v7RAxkda7cDKXO2IaASe7lcSKdhzpMuaP4F
PVlhL0cQ4G5UNL9HCuzzSIrYLPJgy6MpSfRvdPlqEM7/JeWLElrctI/yuHM6e/HLiRzv1nJdR9LE
fOSt9WPWd+kLmTvY8PjcKqfsoiL5/bwXcNK8WGPxYZggkDJBkDWzCJ7rIwcVj271OGfVhROhK5rU
IpifQafa3U4Mc2QXen3MF+bvhkTy3N7BNpaXwbN/gJKzvVDCINaIFlGYIi097Zm7Nf7s91vVbzUI
M4lT7+tGg2URvn09wD5GGUYyVPEx9TvQ2bz9BfrXkYgKawmdi46rH6nRor2lBRomaodVNjBb9tuF
E9U6HBUCb1nWa8xKbE7CL2ldKxTwhum8fq5NVUB1ZdfA26ZYuU5d/vLR6xVL10xRIgTO/cudE9KR
EHntdsXPRlVGZGWBqEFftYl2UVcZieviyTFF8ByNG0m/a0fy4TJo5G6S4bIX8JzP9d6Ef6fCq9Xa
pWsDWwBWAmwpch56kXP88aJCoKEKemVaF78rq1RThQJJex6LyJU1TInBjpOK3fiskY8/+69rHNd2
4ViVwgJbfu3M9BnSWRFUynBl/0K8efbs65bA/dpmuYldXZ6+xyp1zCAArlDNV2grhgNFzdIHPj4/
1+au3zi7fsIqx9FxkvamSIiCDqnwQ1+k3DF02YF+wFsT7AlVDoB4lH1jNTWdanu8QHwVRTViz1BY
+LxFp4TZki6BBW87OKFaRXygrvhP+ZPFdNkCmkYJfEy37QX58ZvHd4Anc5WUJtUNyeVyuNRrXQDX
O2uAKNMY5BDo9FoyF65k6MbwhUfSA2Mx0GGt9EOXor+sUQwIycXmUJ/mvQrmO4/dLg5jg+H7fntE
qWuHCoxiUZITB7msnLww8I1nzPGUNB8Id/fGKx6Jmj/gB+G7ZpRVcOkFI5ghrPjKog5b007VnKno
rwxkrdWeTM2MfebRdxezGhS5JOXFpf+VGHRwO9eXifvEmfHHpcXGG5lERH3uv8AJnbFJ+pxAF21C
IgmWfIuZXMxhBJaUxyJmylqTYv7P5owl/U5apg8bZ+F4ZTGePcPH//Ux18ieCFbI9Bwf2DFLLOnL
7jTbHXVCVJvXaj9Tgn+YBvFVLSJvsjcdYjsWiQOYnPzKsg5gpGiClHnyZghVpmOlepV5hpbpDVPy
WmkH1G7wlsoTY2UNMmjwAuhSpRHUny315Wqrx6kEiE90Za6kWjqlgdg8ruFXnx1FNh0QLk30mpr8
ozBnTKg0ap/WFKLSPpvXdf1J9RzUi3/Y2iymAVr+unkjdQgVrKQBYZSvTrjbCp6ZaSAElqBA3nUE
AafvXwUdMzqpWw4z76JLZgdDa8r4k590Gy4Z82X54aaJd+sX4Mm0nYx6sduxbSnggHAA7fc3mLSC
C74ySR0FHgHMyjpPQMtrXu0lJZgW/T54lmNotrcjYBN23ePnnlfqVKrQSn9dN9w4jgJVQRCqZOg6
R3z4YBfOl9WTYxxpAAjS9391qGn5GoA1rxUoqQe9H8dzcQdO2HxHM0YlK6cC6OD4WjzWmx3cUdeO
XsohV8tPCWHnP2Q6U6+Pq4ckEtBZ/B1QKz4fU0lGhlU3wyIrcgvXF1J7b2iageUydhmFdgIjAAop
lJbeK0UFQ+W1h5JwNS56ahbtM3l7ipjxtOHj5aMYEzSxaq9jcxj8/FsNzLrax8ISrDWF+0pwv6H0
cktdrDzlhTQhphFg11fBFaTSBLG+Fci5XObUczYL+joyLkvb6L6f7KAoj29FQMbpiqvqNxlo9/Jo
0MOfrEosrso9oOHCE7dYM8SN5PXeywzuwRqygtHtu+5+kgYlyPBO/yI5v3VoYrxwcy7OC1PEPj3k
jdSjUM4DulXnjG8ZcaJkHxSVSn8mbFHKyubtnykIklQtdADPFYyuBpwzz6Bi3L5Q50bWW8mmSjSd
NFGBN0I7+zd7wJ843NA5JnIdgxXId4tyyPz709GKgegiPCuUbU+TjO/ZEXpJEcLeQ19mMpIUaybc
poUk4WJ/mtIX+Gqr3GdGiccycF/3tiQgbiDjtnd4unOg5zRQxl6BggU2CYgoge98KgJ7OqlbOv7Y
3c8qRNBRgbo1F4X12oS6nqnd/e79SSWFwVKEqY55d/nfK5faEPB3Y4ZdSb9N/q/Ua07gUhmCJHUM
woTfN+WNxMw6JVqEjf9VH1YiMewaJIDtwGtVzBTR+yYDqKrqRbtQ0vx2GIGZV5Ul2UzSQOPacks8
qLUREE2m+FdqvVv8sPhcB8tH7i8P6hLs8cLC7+57lStbLLLFcCd+2eZM1sU3RneOPMsk8L4DckEl
VErKYB1DIiNmvJ+eFnoag0HyxfNHorY5DX6n7Ws8ZzzB7l58upx2ETBr/jZ8QredB6mgQKySLU8Z
PvIB6Qx0NZonoHqxvGib1PbJYObm8FUo9xvok0EqfSAQPaJN2Ntjb9mSOBDOuqWhOZIP52/7mIa/
jIZlLGoSW7cJSA+jDc1F94oXpRZriQ2oX7PsGe1srqmJJhe06vZU1RhEm6DrHE/8a81vc9bZPWD/
Le8SWy0E7RYsicKEL6Mqnvr/lWGyb+f0+8Hd4pTTOxVpD76RpJYw+vx8RXY7rtWMq5mHBnt0RK5A
rkaCTr/kzVhleBNrHaD2B5ambyn25hF8jgcT3ndfRlB8givkUzIX8y+1g8z+/Wye454x4HY6m6F0
lj/idc8Q+ZqQZtOqkHCRMSudjWeMZlAm+Sy5W5nO9Cn5RxG5rmms9qoUHOOw8+sTZM1QKb8yjHgu
UTfgxViHTIZqPgzXu8slVpx3Q4snF3iV28fOobGVFSadmEJIhHpEMfkF74XnrhLUi9w+kIe3tXPW
OmPujVU1Mlo9H89cN6iNDAx9vfPo6z77IFnOuH0ge9ZZ4XpO38kx+64+uxdvIOr8PMGzf61x+Ymz
+QkYyamhTiW2V6ngwN7IIJgOXzVO3DLGrRAKU1DC4+ICHE/hnrhdR6oCHIcPFNWo4f+L4A/GBGQ/
bc5a6OIXJKtzsrbHnju3ClQJ+GpRj+H+a+j0KvOJjNYI2xfD87C4g9fa1BY6Spvvwz1npYrXp0fv
v5WJEiKFK5lve919poPa34eRVAk5eTcSWRyuWJiLr49+lYlicUeG5CMxG+E0hyNYVo2Qk+oVVXx5
UNO/CtKFlO74njzuojaq+tOX4WOyjTKHN44msVsMdDpEOiQ/lJ7YksCoo8inBs84GJWI2kzdPIFE
YIHPeePObGGjapQlKFxazLFi36HPUw04mhZRsp+QwpxEjR3tiOI9b8JxeTmQzA5zVYwtyYgOXoVD
fXZ5iEM4pxIyCQmysmfs/IGy6287TgzCdE16QQmzcNFG7VLZhDT/A5F6GpNANrcjAax9njpYoTGC
neInxeHcflC205pEW5/6f/scJu4A5XNFoaN3XdKAtjy9IRctE2ymQI0J+MJnzg2CEMi+dgswABae
/Zujy5sQxBAs7kRcIJc8nGtAmUIbq/VjMKSPYRSkigzhcGsM6YkpDguOrkd0L1rmSuqVdYZPf6tz
bVGdOa44rZiAR1XrkRBVUltZXiSfUWaRt4WVM/l+8N9S33Gg+3PbX/AObOP8NEM3vpBR4M6dzxX5
1Tph3hbKsosTfErcWLvCYGZHfLjJebMEN/8fBt6r1FSiRt7HqUkJRPuBlzqEcB5Y1eUvjArVGSsD
NtqUTbmj+7XxzGqTBFwVk2IX9ToeqHwbX+DIPgAEqqw/TmPE+uvOxPGavOf+6VaOO4KXY2lX9joa
CrDFB/Tc0ETH2QFMxD5AmH+ViO/56jA6PliMJiNNF47Z4WZKtbbFqqJVOvWRHfV880SJuse+b/Y+
NGs+x44SblXE85doYxSBhv7r83fFqLQqw+phNrI92ERtz2loJ4HM8Apx0eIz9JlfSbh+8LLmCIeh
hbxet1sqx6Rmpt/PDJnUYgFQrzUmAsqBp2NBQj7pThrIVC8Fl9WUw1qVMhDCxgM5vDB9fM4dJb2E
SuqvMqo8Aywb6mHO6MS/T8Ob6WGi1X6zHl17UqpNPiQkJqwfVrO0P9BowQ073GQ2eFuzVWtqsWD3
d2rmPuU3zBURUrmv75zBM6J0mE5GPzyhusK22XhET7iFggPo2xQXV1ihnquQt6mkXXVtEWzgmiYt
zMo+wt8rZWviDmkpCJChX7KIuAWn3zRD0YbKPYrxlp4tXRfA4vJAoGXonPsrnDDCB2c7byXRECbm
LAl88ChgeljGrsadYMprGYCPB52iV64evlenXwjwQKri94Ma7xzLQN6Z81SWpHHA9yCPNZHz9PGL
Pm1cg3xt/BYg+PIvzenf6URQM45QhT5JKLJpSlRBWw8Lu0WCHY71uDDkuiRfPIA8GltJbSl64ZVs
sNKKkM+EgGhqtDBYlJsZ4aRME5cWO75d5d/ynPB0Dt866EuTVXqrK4yfiXm694qDJinhIdLhuSxI
dURGgYDbdaKOZFPbF48CR6fnCCbujij96zPlsv1JpTkXGdda7+ZDuDy5Zvpx9Er8YFlfoIWQGut5
/eFEW2PfhTwQe4LDwl2ZmTZkhdsffZCNWVwRR7wnbP1Ta8BYjotgEhelpIPOE66aY21gUoar99Xr
8APuZp3KMZfmogOH7RSbjybIqkwIcSjTMxWg2gGqsyZ1gmHoow+C5zpAzc6AmMCDR3W5lkksJlwd
v4DsX0MkoK6mfE3Q8MsS/6T5vDDHmynDCFKYWB+/e+rqWMgclyROwZBX5Niuq0kCErzYwptIfoxh
CgV3TayBdVYgLJUhPyb95mvSfFd3wIw4MeOEOm0NOIRfBjdErlKoO/tm6HbC4cVAgwWhmwsqX/QF
PAFwBXZFz7SKkXy2GSqmPOLd38vT/YkeaZYK3OTPeaTkJYKl7Hh3jjHfvpOSXZmgcYYn/QiqAHSR
wTMLZO3+RUyDlajjs27To5fC8lEffTKyONBqyyNEAa+Wiyq0DtvgHAxTpKCGzFvydoNYKnQwOUnY
npkauyq5sezNuyLvbw+id+kItB9aQfaYwINuP2l6CRe8J6M3FRd2gBCIO3YqZj2gIce3P2iyHjyG
8n0H6vIipqD6NuLKWG8+f+Hva/FgyYKhyBziT09j0DGpWbMmT61UahP96f8ZMVxXY9l6d79E/4Bq
2dUZuJpnkmiyKOgHn6tyRhMYyPjTYL58GBKU6wtmE54nhktU620+q1YZbTwVTxl9WidQLAOZ5v61
uoRcyBkFbBl2SddEw8ZNV2FN3lleFa6jgZ5ZIxb54VuzMFb5ChcxXDZUEvkgYOoS4gNusuK8Spkl
pCgtXPexkdRuk22FAxMk0Pqy/mdP96Tzr18bHYv4/y9WVZN1Qbk0Sta3WExtGCh0L08lfqVJ9F9t
sAqTE2oVYvDTCASWyxaZnPI/6CG+8dLagRdm5rN/6J8qQisozXbT6ROBnUpgIECTFK32/RM1kKrv
fgcIMc8pm3D+M9rNu5iI+fiqtnEmz4wmnBHTUdLplxGxOGE8xvecfVuKb+Yz1J4YvxGhnk7mLSSz
FLJtjZFZb6dSIdZnzHBQEs6XPJTjPrZA4N/elvEmoycZlf/1iJTyd++U9QMCf40FM1F4+/JEs72J
L66lEZJcM4c+MTXep52BQNyclWUexXMEHA00v518GQbbewEAT+ATwg2sJZO5sB3DsRueJt36Y4BU
a/TtmRZAjs6KGPmkTnxnsus9lcYDGD2uMbUetLEtNnScCZHyISjPmPaMNNdqJGC34vIu9v9x1VTx
9o7sjcQa7/ZW31qjTKyLgj7lxZ3OZnUbn+W1/tCG5HcG3j1KZ4yCvJgivspDQ4PkX7jXyYoipa6m
OaOLghdgU/AFkav6XLyQ2fa+A0LbKT1hOaM6Dftc9kNY2xYmYIFSOQa9qU1CEFRgPyqB036SDeRI
BQRw1P581/yCnE+dAG80XS7oGToicDvYd6lvLaeuOmvPBvLYd9M7EltEsU86M0aAnkNGQnqdl4LN
n3q7apwa9V3G5AIZva+XoTLzmeDC9+Sn7FyMI5CmZD9bUiugkIto+CGF+ZUC1NiyVPW4KZC9mXVd
1wlgF3DKMWeOnDeyG/p+6I//LOBjPNZySK3At0UT0zKw2RR3fAL65zmRo0+2taLzM51K/+bWAfNQ
Sh4u+llZViPJ5Pef52Jtck25iPqLictPRPuSM/qtlBIIwswrj/Lxv5/+CmPg+a9Qz2TeibBhloOt
a3D6wW+vRg6klyqMvTJxB30V+48GtGdLSgBiw1MjEFC/fwL9T/76ipqdDy+l4XppVTDlRO/2NtiE
sO7c9eSl1rmCliB2IOstN2QxAdAJ5Xl5+hgQAzRuSHYHK2KWVaPQnSOhEEbNxNhuDT85ucdJZoyW
6eZV8nmnVv218nYKh4/+G95/iGPp1zihMBrZugYMKpDo1EUBr4zamcVUv0Nr8R0hBb9eQcYfytTR
0LDfmCCpcXWIyjv3BORlBswpSzqlhfdOUU23GDzW45igSeYvkiZkgUnVW8mmWYnxU/ZO94T/dKgp
IuPrWSv8X5VIkX7baaXp4dy+ftUVt/1NXOh7aUXC7ItWTpad4VqQt1jpdEjKS+rUfjp3SzmtOWiI
PPdMYfsqTrQ+a+IfdfwxnoMjvvsWWmBa+rCh+SlclR3sTw687o+ypCNpJcb5mBY09vkxiauCzsnl
Yqz0XFR0Hyq5qPkdGX9JL3Dh+PBdxps6IbJzUKS5SvHVGHBeT8cAwu4d36v2ZZgbcRbFBMO9BTTY
OISV/FOa6rbohKDkXW53soD1a7yc4J79bXy06kn1Wyu0aYTHCZM7SUgvjnzZ7a5vXPxhHkcqavbh
TlWM/cJ1SZL8njnWUhoS6e9jjP3KWcS7KGCVLI6iZViI7gWngRig0y+BSP4s+0szCeYOTSf5jAi6
FYcLvzjYCvfeOMDzurUmv4Y/ajifivixrkV2o6wgZ9eZ5nemaSCSCwI25DUCFUp6Bs4rt9dajxnO
fG4E+vOa1KW2UZp6jSEtKG0j1MWFlOUtiwZd6i9DKX1lpPt8ET7kgXMRVgZFL8OSu3XbFijDej5z
mPyBPXAy/l4sjjHDU6u4Bq6JlAKEQEjoICg9DM+PV3tn8z13e3MSFnldCUk8jDxhWzEUsd4VxSmG
Z+gnoR5Z1Irwl6UlGA6/4qkygmXebA9yZVpS+q/Z8duDLPISCPiJ8x48enbDGWBOjDYAGHu1ntSF
OiZjxvLgsY6RMNl5JgqPSQrUaCBOmQDsMg3z8J2PvKABIe2NGX0q/ESZ6RPC4JJvI7HWUZKEwN+7
OkoBMql5MOhcwD08YGMJtlPcT5jBy93LyjCavvbnopP7xcs5aTrxeMulW9I3SOaj6V+KmMRC3FM/
i6hs8vpsssxRg9PEiXIT3n8lJYIkNp9wLIUR0dffcjZ3DR+aQ2bbGFdB4NbaNGWJG+LP/m447sMl
jakIFBUjfQpKcXkNST8RUVbBipNKPDDjmFKaE9mXTOEj0XWQZPBWUplhAPlaMncfnVkniovGXiDx
6nqDM4lv7edMxi0DIVD0Urkcmo/OMLkN8xJEGlcZEsSWaD1Bg6wJAqCvMm8VFZmzHzlavdipf5cR
o5R2o7ih/xz97iPtqNUxeyGLK/kF4bRgRrXpo+Tw2dxx2aEr8PNRUkaSNobJcay0PBqWCgEAXUed
U0pdKDtQyZaDlFRAcCzkR7V1YepIKqCB9cwaIvlr9KBG9ZGA37lpWYFyN/ETM/pbm73zIc9e4evq
IUblnwqJ0FWBeZ+TbOTn5yQnRpCIHYDWs8AJszPYyqpcXhz7UUq07ZcwHBr2OKhftMX1xINkVr6F
DhqUV1dGxOqkBfD4hFF7synqG6JRQrg5OH9svB3Enoh/+dRmlAV5k7jFeTfybht5CH7jGbLQdQN8
UQvLgm6e66tTlVvk02zgbptNpPz0yBuACgKoQAV4F5W/KzqNqN9E48fdNJ2sDaIL9QIWFoFwR1qi
J2FFYtJg+yp/g4sKRDHGFmmmlGvHKUQb/y/iYosLk9s9Mg1NEjvnTwhoBhRhg9+sEHOwtvAgfq7X
R+bRXyrgFShbCngKCyO9WfGo4kLSwgvfzOTNNrHSqBciB9tCNStYtjTU745LAUTfLyocuwBRFJ4i
5qTPv942n+b0GBu5ql6lxByOYTpomMooOvqzcAjq1XYp8StQNofZ4vBZgMsIaMpkHrPglLSzTkKl
ZZK2/kUBY7qIJbh7OI/PwEVAHyicqP+A/BhCbfN8Di5vs1349IqjbT/52Mm+Oc1O5yA6782kfm+A
Ml+LDRvpu3TpnV0ijrO+5FljHwCapUPB4ALKrVZND1k5ADKD/3C5s+1f/vmP0XCPwEyEPYxwKdjr
HKhVpFnseEhFyweqnENg+3eTgaW7nJTqJ4nRFfD0ODhVt15T76N3zS+t7QDaoWYvakCa+Kix/Yxj
WbzeAlyv5xn8E34ZdgmRpAbMrcFyfNN8PCxzkSTKlORvW9HSMWIDrEeEXoE9dJ5GTkyCk0qMrPKe
N28LVGbJ46zxrEvaLMBUZyu12+/UKR3foAlTBY/6f9SNGsokH29mxR+8ehKGjFrMvRZQOLejRcdh
XCUreRdfhTbeV+ly3v9DHhLgg5Xnaht2mGAhlJU+3fpM+YKILX0MELTTyIHviYf3yzdSPRMCuBLG
gAFjlWlQUiO0di12/fkoN5/a+6gO36R9QFAGXQERPH+ABGsWvdM8hkU9jXU8QtPKfrerTDeqqJM2
twJVC7Dd8uVbfJYH9mblCtzFrdNvyNC56Bfrk0jaFc2CsN4yQwo0Flk0H+lPml5RVH9zvfmp8SaX
wIM212LCI5+e97BXRb5jsUviNDvpG94hAoSRgqt5Qgjt95WGwGKu3AFqN1KSmDd/C142Vm/+e6uY
XOGzmupdBmUfcmZaeIpidyOq1XI1/8WBl9T9Vmkt9akHUQZd0fC/AKYnD+QKj3ZQWLC+4g6aVmrw
z3CrSR3pQHxiWQfCRt7WpegglbJT+yxdDpgZpeU3RZu9nT6x8XU5uESaTgp3CWc4BM/ONn4PzTwa
E5qGQDfAJfFUDsGrMqoWscq7SxTYNMDMp1AET1hJGdOoR/j2lXv3VU670L1PI2mV5VWmrGaWH2i7
8PeBzO/gSgb+HSj2ElPUE81zY2IehrNgbJA7cl4O1ZqSjkOUZhzP05rvFdNyQiqwE1tG+I63fVCN
4ALq8H8Q6TcSkawL/p+1VwhBhyhddyGBHp9BTNR1xBRicBGs88lX3GV0V8IKxRMZIFNLZUPOIrC1
NYI7paIJF8ZQLdKgvUwP+MFapwHxg4gGx5Cr6MY0Kq8O7c6ztEjmnPGjdqbEejRMvtN2s1HPGkam
2SrLTOX9PjPp+0btgtAvKg1OJAdgXQ7BcC2hpW0qquOP8siuuS3n+yTcnk1Ty9kAAntISjnV/3eR
uspMhO7rDBc4olAe/2cOCdzHWOQtGafin9SuaggtIy4gK7FsJBw8LSXCoJMEazZs9lhEb/A1anVn
5weLCFN41GsfM2yovRN87W3hcj59x0E40tX/v6Oupa4dqisOQUBFssX4OYf1biAMk4nHCAtwh0dQ
f2UTNe5WJqHtM5XqWBWMVhEWMUPBAJ22wKVSr2fmj5SgDWXT4X0L6iT6PCs+d4nOAJkkELBRc53N
zvl72qteghvgk2r/ZnUroZNPAbV3y/RffGeZHehjO3zdtowotqx28lLYQ4t6XBWyazep6tSu3JhO
udnKDS/i3Q4Hyca4g8DCGWa/9ueDDGa2/Zlk6ZvQOKsbKI/uCooptwJPjC7hwgTWc0APq6z5XjzY
rWNPoZrf/r0muaT5KgcAq53CLFXkC9w0E/B70qg32xJVp/glUCugi6iUHcWvySIm6roc98P1XTz0
dANXVTBdr9LTWYoSWnKcl38P5veQjZR5kFm+9Husbn76dak7BOkr3o7RpdTeZycS09L+2CKZURC4
NDJy0zyr5BQAuY9uKRxqWm9dTL7z/yjNc/iu6rqevrYjvEi4JP5nbj3eqHWWDi0hy2+/0qGUQIwi
YAQJfuhfUqcg+IPcLULvXkcvIE/kUWhwfskwTXmZt6vVcDraMVTanJYhM0EXiZ+9lwzZUHv/Etdy
koLO2/r6MfMEGP8yjNG2v8O0Azb+6Z5sWq3jjZVNJ1hKr9V48Q0R3PxHesvGFcnC/ih2a/V+IKgj
xYCLTrW9BM6RiXDHgZOWjk2nS1F1ILsYX0m7xHQtEExNtSeXFuKNbNaNNKNioihhejyGZ4hkTEdr
F5Hj63aONDQN1jmrPiHPxq36Kq7/gjM+LpS/zU1fgBUwY+bIrJD0D41LLelKPYP+Ze9vutXO3KuJ
DsVEB5bhRC4VbaW6IyGQ760kGgSJbi+nzSE+6efnPFPRJYrSUHvzWGfC8z8XjuxmLemIoxJ8/rcN
3bbTUxtv68DcSLWpltBj6wmsp23xPDKWwBr8yMywpLhrNVur4zGPJCc7fPZCFP2q+AzbdmSy3Ia6
pQJE864fVDUhfpJdj9sFNKMeDlj4aXW5xEiUHSf/y7JOK91qINkwHqcM9ZP6zfpGO09eo81LNnRh
E4RrJewNh7M/EYKm3OQxWCAsuCXrFwElBRzeUyXegQQ9VRZMk5mNNAk/T/93QQTDwrjYBqcSQo5F
Q5q+Nx4BcnbKlLKdY8+mCpIuMRelpxFglkpCrzK9h7UqGDg3bdUcvQMQWW1X7wx58fEV7bfDX4Oi
OsVlEnhmRcQk2UAJZ9oLkStgvmhARGV3m2cKuC9vxB8aGHcRuvdMespkPiVJyG4na4rVj7/0AnVl
qngnJ6KKTLF/jqV0VGgAidlPIVJsheD+69Huc4cJU4EPZvd6X3rUMD/iVfUMIszV5jicNEmHiVaa
MZEG9hD7tDKXRbsfArLjmzgXAaG2xM4mQB0L3yXkxJeZqqmFO00uE6t0CQL22diFurJqDdNw9b3s
5FRAAcGoBJMRxX0EvtX04LBRdtv1lXzQLlkmgAsxIw7ZMKQbtHEkQFN+tyBukz09uhL/5gn9m8gJ
XtRjApuBAC2BF4xVZxHWpRJoVXAtnm3woPAHm9zPs4dF7ORCMfJc9TojD48JgYGyUkhDpCBAJEdl
2GIv+OPBG0ZwWpUGcL5RQp66CjgLbDGZwNeysUh5hwWiImoTzVNO9BmCXHHAPaNJZrk/gl03Bp0T
DQ9FwT1SM7REe3f7UqVN+ucl8REZeQ499SMA3Dv5ScXkrL6/AlPXo1oWEb/uG6BFiv97JB5zszp+
d1IoIw/y5cqP06dpDgSLSny2VGEuf1oaK5NmZNITfqgJkVojxBZO+eh7onaDrSMYKeLErE06KDYz
2ES/CGR+tvBzTxX29R/6kOoVNcsGNtHBSqs25t3WJIe0KDwX4tjAf5sindtjJ/LN/m9QhOgkBql3
zSZJF7F2OmP4f6iDsq46BsVI/cOLNdGyAYAewtBaZWJqCe1LSvVzruMaSYAh+wkjj2S/4E5x2K7n
YQc7bPHqEbjr1U5ZJgdZqVlNPjP4nnLQbVjd5ShrTK2KBblL9sqRImTkWiw/8WtYlePea9oCeNHv
jVnZbM0QhfCgB+xw4qg9h1XbcrCwc+0wz5y1leqGlvSJCTnh8Y30GhXVg7KZ4mlse4vobj7ZGZYC
w7FShZ5p105MPx4IsgNQN2WjKVnTj4+LRnbT2nxUuvCZCLYR1Bgrj3WnoymWr0SDUWXqwgkuFALT
zorbgOW3vdNTOU+ylF1KclXd57hHx7saff3VBjBMFZecPSL8xU6lz5B8CpDHIo+2H82bEFuQeQ2v
uMx8ZlYWSmsQz7Y489vrBAn6FrKRbQvRxpfcOeoYMIZL9xBqNV2wc87ZQLQ1C5Bbklhni+eZzwbs
gCERr9vrCUjJB+Mk+iSgaWJ0m89rwr0Prf5tW3REYH/WL0k1UiF6YkJc/vG7u0LQmX2GvEgc+uVD
VE9XH1zIQvU3l0fBstNBUqY9NMEkATRupYmc/yFZBMVK0j5TFWcCP3+Q5bVoGhjs5Y+YwFj1RzMU
ItQC1x4fBu8LJZ0H8T7V6joLV7vHrRJiNrQE/sDbCOnbUD6RC92F5Pc6ttsqMbIE8HtgxLzWhSXX
qZF8D2k2ass5b2QlEko5d0h+pVjqLQCx/ZV7PrL3fOvUzAKbqUJmeY/qpxJG/XODArr+gLbn6cgS
h+O/lS6aTLioBTQuTZIQVS1kkMNAukhI1O1R/Uc5sX2oIzAyqGYE31EMbxTs6GIdQd4dcJQ2EoZA
Rk4nAuInTdUFHIm3heVpn9KA4GALDsZFjvDRnJ1+WDl7T/Wl0GKEYd6rFvOrZ6lGYvF+O6Alr6Sb
PirSkiesipbfgc7Ju2waRb+K5mThCAquYXvv2uzUre2doqaMmwws9FzrqDYmIXfRYQov5onGjPP8
Wzkbn0tSAdgPhActTc0DOlVoHIpyKRnFp0dT8WyHlu+lRwTR1WxXCwdtfz8lD7Oe28UqFWOOrVsz
33VlQeB6k3AmJ8H0d12vmhKht2R+cGeVJR4FFDnr1sQZ+jXbb5eDZO84al0R+HGnze1ZLp986G7G
K6DoRwY3Zcx9z+ZOjrcEm8IobeQAdCY/ILVOFK5s4mwTbsOOn6jPmZPqscWwv41+5zWfxnnOp8oj
MHqHgeMPJ4qcEx0Uexm09zPBN++RTYinu7STbxP2qlojWRLxcnDWL4/L+Efv/rpnnQvj1UK/4eXm
CXobh+iqHvZxBjTiqC1L9855lGcEoHUuRO8DS9i/0B9nF7av7+meaJvduSxqDN4c13DZ/VsNKusB
rI35J4MYpFjrL9ut4qDXfeO9CetFR7afJjh9WITx9gieLAtMqFTcnd4NCHOypUl/EGnWnUGGY6Qx
YXmIYWKswyJVRS0/uFJhDRKKXfGM3RHIRAL03cBuIOi1lpgFMaTfq7GgAx9M9BQ34eD4g2DDHu1o
13B39bQURCklthrOG7v93FE25oy1iuNQ+KkNXsFzmuSgXA9nxvqkyQardiHOUVikEAPEFABj3klA
Bs651oqde2KGY0hVl9SJanKV3V1ETLlvNxA9ug99YXpp3U6Jl/In9u/viMzwG2MzSVMITPzirH4u
wiRhiGrR6V7tMZFtRINahJYq5/AZeMjao5nWTSpvGKyKe0sd1GwS39hUX8f88A5fljZliUA+8PvA
2fKci8ySmz29CBQf7m9TwpShHFNUtU7Cbj7W1m8lpPj8HqzWRtotFMbVqSVIzn+W9BsnGCU+R0YU
Y9cMXomwAzGDjBnPGMnJH4YsaCN/59U9BBhYVga9YAS5FCVH4PUJlmmUV7Pxzhg2JJQwC01h2qaD
yDgXAyGSsgPO7ohj3GFED8MGiVC8z1g5iTwPZJkQdYrHtQlDr8wDC6MomGxeCNbch3nsK+1cYXJF
2LB7EKKb4NYa7m4jucvFEnh4O+xGHOlIzZVlPh5KHM0jJgh6CJWU+1D0U30ospS41JZuvvNRph7/
Upz7q3zkheS3lYP98mD6nqaK3/neMGg9fMrpGWzdm+NbUnU2QskYgl0T51RIqGYGIHuQfFlg3PMK
bOidHcqPdH1XL2MnN9E1tR/0MKyhG+eUb2BUl+Ea/t44o0r3eJbbZA610rXyGjPzNQqnJesgBlAV
5FjEhNoK1QIZO6zvsHwX8gLT3efTbODm9ruqXsQjjyjjYh/Z6d7fNo/BH4C2ng1NAVhJdH74Mi4j
VCd3eDIrA4/6QWEMpRuhUwG/o65WwXIeWFOE914z1YxrQIt0Qt9bHz+c66cezqujMWE0CogwTPmc
MItDfkrZAUE9phY2oXBQstqVgd36fLW9lU34SQbEtWI+kT4QlNcjL48cGFFPm+o0PwCJlXBDM1KS
uzHnnDVZ3JJObJyq5o/Dd/LkwCigyG7keDSu6Trf7iaCCcu62ouhUEwKTKAW0+LUBvkZhGyUS1/s
agLEORrAlj1wCRxOI3YeiyD2Pd2t5PS6yiGMuUdL/r5iRXvVCoR1qepTg4ISZ66rw5DhA8KSt5RP
6r0sBReGk3qoVU+0DKwYIe49xGy7GhntTJylvt0LB0SDgmAyrI9OwqP0By4ErwZ+Lv03qDxyHZqB
slFTZRkdcAtBhV02XNplrdK+ttyAzRYNWga7EHTjApk0Wz/dl/RnGDrD7MbS+X/ochcwpD3nMa8G
cbGMDLCdXP9k5gzkcAKKKgbASQmJMC6Af3PdUNmotn3XeoW70Agb8nYjFFkn67tXcAxo0J5v06Cg
gK3QSKtVjZRnDKGbcwIUBFrRTXGMa5smJbIP4a6fqf7f5k0Y5G5B7VHS0exYPR2g7Zeb1LJjCoTT
ZZWgXd8ksVQgWizBCzrZ6FVRAOci2oupWmCEcufv934ZwoYYN8rsJP7pG+FMpQbcdcBvEFMU/CpR
UciKSMroT02d0B8G6qWKsToemV2d79kkxiWfN+JMA+Sfmkd7F1xiihafh0TUzGj9sNkMioA5/sfc
EWYuFVlq29U8j2d0kp5PeOvJC8n6Yx7btrnnnThrbwSt592C0zPAZhTAR7K0gPRrS+GJp8hewn/z
aA9iw27/EXtNh8EYYPYD03KTBeTxtEQIuPBd2lkUr4y4Sm7MQXnwv5pRg1IXegaK0OjdzklehDon
Zx0FrL7Xgwfsr9l78VZNwh5unYeCM2buLsM1tsT8kKSzRcu+pJoIN1Uzf+3waRdU7NZgAUY40W5/
Y5d9DGlEts8vwdbdv0Bi/Fcakl8GyjEuc1XfEE1mO/Trt1mR/viDR6WbsGnZuaYiiJg4oqlt1mRY
d/KJ/h4J5f2gHx0zMN4t4+RYzRvJ1oGJwnWGfPZjuuNkQPfcJzXs8aAMIRY71jhtAPVj7Kkh5LX5
t8H7QCdWAaAwVfcftmOOOuGI46qUsw12/Qvnzq708GUJ+55wDyBzRihNBwQw7gkmEKS4mzD8xkr6
h6WgmWN5Wyc8ntbt3aPADxb3GOJwL+FS0jLWL2l2fwpYBTKPZ/WJFBeQMd1WngHSPzBuWBQXKsO3
EVwvAOLeB2Q+0nz/Md4qY16sNs5UXS99CDOOQxiQWbVHkqsc/Aiy4rOpdllwQFckaQkJZpXG8qkR
1jM2x1a1Z0M2l/PAPp+TY8DJfER3v8kB0t+kbNetWLCz73GDmwS/LCX+E9VF5B4H3WCHx8s4hY3D
I1cV3SaIDG9VCLCEJKflMzEt6/fcmia9UZAbheO0q1ltHOBWy1oqx2319coOxCubBlfi8z8HFlhJ
VefScShQz1TkPC5zKv3tpgg4IAYhVdKBOU6vSkLq6L9DYSbRssyJX3JLIR9fgi0zAX2VmVU6Ce5a
0OAy4vStw8f5ompeYViH6Yp0kFxj+hxaFAEoPYa55Hti4SFZjFcC49C39G0UNJ75d85nBF+jZdHv
66+hiM6GXadaCKGAzium4dgfNUazTb1r3tKOFs5YqcqB+7s1yb4thGrtPCCru8Gl4dNQVWzMHm33
Pm8s0Khhx1NbHtmHheOy5pnMz7rztgfN6RiulKeaVE9MmRcr8HPH3TeNwDaKtuFWbk0RdnY8hSmp
TNLM8O/74mQHNPBLQsc+5VDwfBm/0/lHaB2M9EJ3eR/agDVuem9gXX7eKVEwS8USw1cz0qazaiGE
coqi0qAiHfZDcnahf2ufosBNrnGFMg3RiC2l+nMyTBT0WjjbG7A0IV9CK1sShAmcMn/Qr5tnoJDm
GRESVUaPn4+rUGzWGt7ZFO4p43ciB9nKbHxmVMSD8q67HLd1e8LB+vzI7tJ/g6XLCdNkGHToAsui
HJ9pCszI/NypCagLlrvE1tyr2drme2Z+2hjuOcP1z1KT/t6EazMhn9jYk+rW90JCTyHwOMB4VQlP
0rb2i+xgyGHScMXG8QzYd/bvPLBqNdeT+h9CPas2a00aHMhwuji5bki1gA51yrB/cqk9Nou0AOjO
EznnKGuTKFFlNGX22BpLuZFHYRU6wE8AeYBNv8KVxNolz7av/e2p5bjfZlwflzOBijFrAwnVLZgR
Oeza+cXYoGlwd275nljU+5x4ZAcM8qXdQnTBVmMDc/Z+47b1HcSVij3nPLyT9ix36SJypDbks5tC
AHTyasPJ5nSVPuftFB8GMaN+VgQxHGf3k8GHNyJqcZ3PhMIr8UaMWt5ZfYJvknfxzumgKSp1Fzsy
0VvoleAD/ju84XvzZCD8NpaLwsT04W/1cKxt/pfGkntjZZse2KEs9y0SonX3JxUHNXo6hOvHIg3i
2Wmsx4vYkLXBx2cXYmPJkaQFpdap4fsmRZT1UR3GxYPY1oUbhxvOCgLLAQBGnjDC6WxULc/w/EHX
BSS8nzvF5D0mEGCSVFHf+nj4sqdhdOl0eGGunZYPSLXngQJk1jvGFx3Ef8hXezM6fLCG9CxrmWYO
nKrP8KdLVsE5bKD0sjVfMH17wi695F/kR3oQOCO/xvGPGMeVKp0Q6PKfWnQVdxDokBz6VHaHfofW
KWJge8pTfMiBzLx7TErtbhjMdl9GWhgKMZsuEF19ovsfIoG6C2Es8KyZ6AB22Ktxdz6G8VFd795R
s8H2U5Kx8nYqJGVPDzeOJVVlqTd6w4F3r4WqeDLBYfWSZuO1khzTS2m8uYT2FDZN8PyXU6pbI4ST
FiEhHieSnSM7/NmnmMONb/MGOR2kBgsnX8CjucW3QmjP2pRUuHA4Td6J/zYxEXSUZley8CaqvojW
i53Mr+N+p5o8LGy9zG6w0rgNeMzvOkk9tS2pGhc1kxVQkGU6ogB8Dkzp3aADdfclSVGqvt+GRUFK
/Sp8VluquHxkPSbzwaxDAscTh/u83+PsDCJJDn4FIaUO2NPaeSDZ35QSmI9uATNgHg0dSWon1TKH
uQw/OHSA8zswkHHs8oXqVNj5B0Er/UuKFTuInYwCCuI3QCmiu+4A2z/aGCEzMew9zdyRPrpWLjJz
nbY+gOIdFcvUYQrJmxGVTMjvC0VRjpWxtP9IxqVMYd0AigGuoa16pOHPAgXOrvtX+LX1OxE8UrZD
B0TVddLvT8lulEsBMMs1+W5gtOqBTeesThNo9Ogcn4dxBzQ+gjJdBbkKl5bvWmDysQ4Ex4zVSLsu
KHtFZfMEvwvisOWPznAdAWc5Ud/+jAjLkXFHJmWBg4ZQ4NXh5an8bcwdCHxl0LAmghuxpkujEzD8
iIaZvn9uZKmaEYmbNPKmbBRUe3F0nv7N8StTaxDwmy5lfpJEp6FEB+d8WeuOH7KBAGiLzWTEeWAd
DosNRgwddPebdW3/M7oHdE0mdZogQRvCnB+9Osb98ccDbPzQIyV65+T5B+EpZCe5fQoVQ0xgjMLG
YNTkAx2+qPH89CXVuUo38fQ11LZKFAB2eMOnFdaI2yAGmlfvdutwMI3sV1B7t7iR6uw6cGpSXYG+
ypYCnpti+ZrcrLmy02NGKKuj0ihoymzOHKLy2XKsvpYtxnWC/Uf1R9CNiGGDzu+N5knePq+YqpJ3
ZK+udbWOiqDxypFBnVfv0gReT1eXWSdmXiZJQ3Uo0RDa+POb8sy5p0QPqmbBJsqTClVojbWyarHU
vSOQbc6YqJDTzl1WUHpGOXTaEL/Rui0AVY03hQiNLzcmoqqPv3fNl7hhm5V2EYtqCBQPvblv29qJ
fgptNDY/mjcN6Lg1N7Tlxhf5Ow0HS9Helz4U0X0ZHgzSdLebXIa8Lc58j6gJx/VyZICYNRSISi7f
rLHwHRRC5KWFaJ4+F1ccI29JQWeqY0PYVsC5gReW9cYi9S1Rl4JrycwBaSQs8nuzyg0Xw4GS4J8O
xyzvheySkNQacTr9MmwertuQNdttxV7XUoqvdVpVT3lT3Xqh7PheFCc1fwLJ4uL8Eu83lqvGzHjV
G4zCqCCekKWtWFibZO41uMWevv1/+n91GEH/sqaJ/BQXcSHZwN6UkwkMv9q7EYICsRPpsCp8c5BK
8YVKoYBLvcMVS0QWAil749yeJtYjyWPK27bJIfq84O3oLps/TelPLsyKX5k89rWV89i1dUT2U3ga
Vq6l5ICew9WHYxTz3NIsnoWl4T61Eey7KIydR0auL3CJfOVTpirv6Nposw0xAyyFGmvKbMQEcrNT
YDByQpxWI9oRTGiqfZfIxdaluPldOkvuRFKw8aNt4aBe9+GeW3td0IcyBOaibZ0V4A28PN88j+wf
7yTnsElyg24e1JFShQH1aJCCbqRnEKryaTT0Ho1gjBA6FSnVxTRSglyQfPZPNQMI7AB4jXQml5eT
J3x7BP9kjyi5IkedrctDDvFYgaGBBfF56Y7iGFnReJ+ZJdTXgVx2w5UeXT5Z9EOEYDSgdBAZSBjQ
KscCFZOie3t9fv3CUPi/YYDE6wGO6xuqSfcerk0I/p28bvq0yNLl8HQ+v6CFQVc8vvuA4/4Gq920
YApvedcyaNfcgGL+BRIXG/DDArOwGYet7HMAjwatd07VG/2JdthgD8+SiE3Y5l6i1B/eL03TDvKG
6se4p36fq2PEXilKdUhnikiGBrMa6bOXE2m2/+8Z++cHQ3261OxVq/J7e+XSKWWFW6L6EoFASbI8
hbDCZDrLwdDCOa7sn1S6dpaV4qHl8wr9ZPW3SiGPpZvOvFcNUNa6sEeuAp1gOhZh7rFOqB/0VPpF
5T9ZkzoyJQ12ry4AxNbjPZN0uQyI3uhokr7n2ylRsVe7OYvrSAj4Dw84leXh+Ac+RAjiufQGLHdk
3PiXpRtVOFqcxgI7S6GJk19kghLzHogqUl8vgb+TEe3YhSjHl4POWDjkzL/AWPp4h3NyfH/N7SRr
yFAWCRMAGUTx1kyq/v6d88nV55LDYE/L4tmZLiQFBwQZE83JTDAFLZfnMMJGmm2SmL7kzaa5jdHL
f4uR8ZS+onwZtVqNeqHcZT1NxsuWK0y2hDN6/p1z5xei0pI19iWCDSDdBfuHg/E0vfN+Za6YaqnS
yloBKs/ff7E2uTeOT8uplDrRNdijgt9btL8BY3FgAoKaBCWF+ZwvIIy684U6p3y75CIgA8q0zWeu
F7MDPY3r6+bjNxcEgcpIyrqc1qPO51QsiFufyIsnM33G4FZEH0YVU1ntn8a/4rSL3Ni9wcb7Qvyh
C0l3x1d0bGONwR1FKSosGsr5+ZNq1YAQNaKxHc4/iO22QSYZvy6iCTNPSGHeL92nS2OTgwxfRgby
810cZ0ctfJcuMd6VO1WG/CR6acHgOqhUMn1s9HUicOhyn/oir493r4NrlRTHGemBF3X5eSpnhOOh
9ytvv0Q+7PQNPUVnMVl5aqa+wvzx0CvYyycJks1S6bYE+KmusFBzr0PTyNGfPIS74QxVcWb0e5jz
ngEII3kTvfsQQLlAkFdOf2zS0AasH0I3YbNqcoB+0cmgJj1E5v0XCYNxFc37bvFGXqibPFxc4h+A
o8QyPZ6ija7PL0kAvSV282fwfZXWwY7Ej6+NQcpwjFjpH6fRbM8EUQ7j7H4+9eOOu9zRjdoNDwtH
xSdeP8fd5qFUCVSrMg8wzQoxsLuBLaBxQ003zNqwCrBbyzjsAGGtL0kaZ9aJ1X1UUZ0SV6I0qYLf
M21VZ/OrC3KyvumjMeZ8Qu+Uwldv2m5fEFwuIllWmoSbNoVCh0Oy2+HCcTnDzNrfiywouOSH/EjY
P8KqLarERiMhqlh2GJeQpiB8cDZW25mhj9yNjJL/sRH/fSXcY5G1x3ytIV5rFNGUG8jfq9peAVrx
1+f+zeuzngeL25bifjmHveCTWS0NnIZQWx1qckTkDmhDFJH/x7fRad9chThpIYYCIRAt1FNShY8p
a9SATx/FH8cmQ0FKKNPnYC6BiILEFUCEcRes8ymkINImdqp2KJQ8UJBZfZh4isASdLmbtxJVB0K+
gUFli4Vb+hZpUY0yRXeqRzhIw5TBakCLvk08g0MCpZoEyD3LQ/4RUCuB+QATlRI96aX8ZpwLDFfT
WnUkcT79//1Jwh3TxoLfdxkh0WnyO+LPWJzc5PvzFElad6nxCN1iPRzK1vfWs/+wJz7xs4R1dwzE
5g/Fg5jvKdRLLyBJlzpZPR6k5XquF3OfI03RvevggMPYG/h5bUDaHdS+u1PPHgvBlw/dG9/fNOiE
GEVJcEbrMoryzrbYiDugxZUNJzVe3hGMwScw205Mg7WDN34IPITc7w5mR8RZH9rkvxODUNEdI65u
j4BioSuf2dPe/E0nR8TaGQH8Hc3RhdiIwufHNj81tENeQ3ytZOEL25sOh+MGb2DYMnKy2HBug7rt
3CZHBtYnXLUQt0D+g0laivxyk6TmwvI/JCIs7Up6e7vUW8qiIwWMSYIlWfMDBUh2ayjQmUBd5T5D
3SV5yhzu+FayeSZPyd0G5e4I0GsqVKgkZXsORtisaTVR61Yvwz21PN2T620gvs47urlmvXj9YIS0
lnFyOolan6xc9un3XYt9ZbJWy52PXpmGpxqcAA/zCn6nChveMLkmDqnAfs4w74fs+A4NEXKNc3sF
IYtZLx4M4u35b2XioBOIJX5Y0kjuY/eyfwUE/47l15LaH/kheAEuuNeGk6F47zUE4ZPY5Mz2WDKc
xfYzgdhTbY17nV3HBHEnBdCXrxN0lNX9+EZtFZR71lRgjXsH8gqfw3wDzXwvhjOlXtVfou+VRgdt
+77EQ3VII27JzeIr58JMI148ioKk92jm7PaXDIqZaRn+xLYhNWo+n1fi21AiA1tk/9d6o5KoKQ36
HIBnXpEiMd5TKHfRb/O+sr/H1GbO0WeozpVF6qbPA6h/g1wcrdwSeYJi0A32gwI2BQ9GVzRir6/3
AmAR1pzsZ/Y8zDQFDLMLGH0ZE3ctPD1nGNhEX5Z86sx3Kni8k43ceUid/qPaAwqtR4zA+IIu3O72
8LoMD7rePAhHqRZYvGX5rniU7ZCDSg4t8g6teKjKbsq9QtWK0I53mSRb0dn6rFtotiSr4pmYdjnd
lD7LwbzGIxFEGt+c6yfSF1FN2Yu/kFAaOZPnKJNNLGB3DM5OfXoIcjtOvosyezjSBsIrRQ6ACUqk
8I3s8HtM2ag49K9nkPKKgQ78CfjBiSf/S80+oBC57StqUjAj4d0nZ2/1iDzQQNOErj8SL+7YsM45
xBi1sf7yZRKfqzZukyOogxJB9ZcFUVEbbR1dOhuyorudLd5PQ4qLwxBtMEPZWRKo7VcRWActFhqy
MGbPvHX9SlMvoP/lkmCdgUAs1sXtGK4TtVL9CqwJZh76aF35HwRCTRND1TxRX4Jm4ggqET/1ogbc
iXl2bXqH6wQCv0MwaI9lRQrjqGYqzRC344aM0WyTtXezz3zvwcWyJUnyr1Njiyg1r93cNqNOcCxn
yGggzMvbUc/Rwp7hKnLCyeMxXDkMeck4qGsJVeQp0A5CxKaef/Cgjy2sckqf0rPgbIhubz+pB3ub
af7zra9mL4cXVnp8OHqjRzOb0eQ9966WKYf2K55kZ1PNZVh7tUbFJyA90ymiT43da3vLtB2Mn8tT
gOuF307CfAttlr5dd1JgZkV9UJDpJeGR7zy5ea4wPs4Mdsifljjf3GsZVulSQNV3AbfBuT8BYtuu
LLomAe28AefnBZ4edh7YY9zSjQapMzf5VkRoOApicP5/XXppP07thVrGpV/cyY7H00oP2HL9n9b8
R3Z9sw9qNMs221xONIC/iyc66Mi82A1DeustL3MNJgDAU8C01kUDqnxTksBJaM67Vcj8fxEqbn7K
z6TGEaiUofxWOTwPXwnQxwoFexHy3fy1bxM5mXorvneKN9ykEf6+i7AGVFPFdi7cKtHTp94lxD8d
cTj3OlIvf6/CB/XlcrP2s1RDqKeSYS2fSVpo6e25rTZRnBRaUYqbubyieFxDYFGkHsXTlb3Tzi7M
5mBdQ/L+j0FTJhXswys9HrO5TbE7ggYtt1GbEvD+XG6DZ7R/n8cfcGrV9Ts+T1wFFqkjUGK6BlGO
qHXm3mTJeplaj2nU5EEJRF9+BAqhpOvHutuulJMwNpmqoLz1I+clWlz+3an3sjWSF2Q0P5b59Ppd
0MyQ2gdYnSkjsvKu2xazmXHonuMDYcxR4r7YlnSBzjh4FxoieJND6cAAbwmeRsoiJ+XF08ENeIpu
t/ngJ4I8VZCSRIrJDQzOm/KUbfw8thdilDCGkSIsrzHo4JTf3FN4evLAqDAOj1n4xTtHGdMUjNSN
M0lG3e/OGqv5muQSUVB7rGpmZZIm4/jOSb9Up0IIG6sXj+3h/9meHX/XKXm5VCHim9P4fysmeUD7
1jtIuCN3TU278+Jreu8wliF2uS5t2Ck6KfQUoIKYYEzIt7mRqi1Fyq/t0peqVdJCERBxPjVvNeap
HJ1f1Qtu6jhyKLukPz7CmSviIOKie3ZpO1i9G5g4KP2XqD2FUHDYXhUkG8gc9GMsuThl9o6tDJ6A
ejsx91jcZRr/ErBv4EOw/eCe4zm9nYSzxhJpl5dKJE7k2ZOrmc4ZwUKrajjJBsHpp6/VwzD+eftx
o1tyzd5rGRvAZcB2p6xpBKJ65TE+LQTIGVMWgRSKkoFeYao0bsh3FGPSf7McITuR9SfZYagbl632
vJtT9C7TYxw67YMJK07v220qmkjngEMzsx6zEK0C4c2sF5Gl0NaJ8S1Yy5CjWGGb8THy/Fg23hGK
WnTWKqUTi0aGaC+Pg5GO4ID2yUimkgxJibaFZnHk07zndY1dZPHufvs5oLeY/TyBDBS41FlwSkzN
prmakxryLT0fz284fQdavllcQWFzdbsZ5Q+VWHDY7+jqvC+VA6qDJjWNBMx2Q8ZDiURyULy/v/qB
huoui+MBN1ukornHsUOaW1Yjetg82bfuM5U17LCaQ3HPm6eCDAOqK3lVZx6DsaRc/pMxyrIikKxE
kkLsQP2oCaO3Isf8rfWuS9WwzCiKo97lO9jOA4vNqB4wLUKI+QgHzsQcrEf1HAXst1qKRmCxGEpN
mXkzDxPmrRfxKexYVPuhUAjoAT0BOiR+04F9QY50cqyKEmfonUbCrumqrrNLnsZvZcddeubUjFAb
3IXDPMV5EFVLO347+/XxoQ1FhN8nm1Ls433dJOCnNrMwNSBD4jp8HNTBZKuxSq7uiA5eVS//79xs
jyB+utv5cPI447+QlAfuoQ+zmmkWg+wE2T+YGiOadUEGn1+8Z7hF18bNxl0vGEdm8sGKBG9rUO5b
XsAP3FeaUVInlBRnvAVWuZMgnmTi7qJGkC5HYL9Mt+AYJ6cnxntlBgAU1PhZiQQLxrMRVLUp/7U3
EYCrYPBeAwx7Azj9N3eFqpaBfRnkvxixOq60A99LiyqnIlw1Lkxjzqy0Bd6GhQWJn0NLAV2MiOPy
8ukoIiOMQDsTcWBNVdgkD9czvbEaSdL3clcPDqMU7iYdUCDW8JnQTbASoL8WuYd6gjAAqI51hS4o
IMexi+AV7aYegTOB0uINz4B8IWXwxYHSxFGupkb8hTTtqmK+04q1N9UbraZCEpm5WsDg5JkZS80k
FHhJUqHCDD+C9wSrem2RfecJcUCIiVU4DVN29oUU2wCORI6r13rySVJJjF+/+Kc7WybaiRuhzH84
jTeKR1jR5ETyFYIudY79gzbnr9Eyj1Xi0C98+oxIMqg/bfd5MZ8qDKjeCws/3TaILYLn3cYFkUbY
/S7eKl4fef/yVGKBybDgvCJ8CAa8GAx1dstqvEOz4A/Wrz7ghpg10KsrT4Bx6vHXPOKUMfJxlydf
GR9OnNBD2VOcsCAWgwTMBJCQWVQqfBWp7ZsSa4zVcBIctD27UKRtJjhTDL1zOWTwy48maiNW5X/q
O+EXVWq2Mcna4JQdxmH15SqNpFwdEc9HbqqGdry2C+iKRzQjZc2mncEQUZ8w6m+gC0DDqXmFHFlb
osiwf2Ry+SABcp9deyKpIgZaOGNDZGg7MDijeBKyBB0TRcPVoWEX4w7TYv3RtYxJ+QoV+KicGnps
UlxKvx3uSIS0UPnnOTglE0piEG8UJXYa9YilGOXAQB1sXf6dxAY6Izbm12KwGTf3ETrGr+gbubSd
hkJaX9JAJriJTgFnEAMjNNO5dZuuYWOZ4mAGCtUjEOuvRHN0C1z6ZjaUsQ+8AUSk2d5avSFPqm/7
t299ys8lRsUi2asD90+EnuYWxkcSTPN+250g465JfOyuvByR7nn4L62ywSX62johd2m8zTHUw9GW
evU1jpqP/kuscNnnC4xdJOCsbUXUp7P0Lg3/fbDVV2zl+/rTn7Bdk2rHffDK1gCSiFKWHy3OmqJH
9ya0ldenQ3XI9bbdqP0wKwy8XfqDJvM95YL3IrdNEf02C7FpTJaEgPXxGPjzmJNO1Z4dOnUjXNcM
PTtzbgYk5MPIlSVekCKbchljdSUnY0kRrHxE/i8AVAcQJlcuqRd0EAvDz9W5U1f+ciphWJZ5O5h1
e1N0J4L/jBh14qtKTzvUp1Ci43qju3fOf+DgbKi8bRsDvpVBYiPUSlNC8OKP1EFiPM3tI6L9ISQd
0djTcSNPP2vKFgrFsuU9vVaLZf6rZiJztAum9V5TStIydssdcoEplyT3LbBTJx7EKrHDgGJ1jVR2
KqVPFZTbr9klO4USSTgR5G1DIsAbfYCrpq4EZpnoPDwUFq1xw3P7dHdcXKcg/IvVbeOTn1l8EDvJ
7hGDxSLZGrcZ6YnHOhgWbeemT7DTV1MnbQ6qbRXXcIVr+jJ0otHATKn1YzpVFbmmYPulqdyL34Nk
feX6rKlYPyXdhpRIdtyvb+XoZ/jcwW4zUtFp8iGQGKi2Vk4JFSBCe6Helmr5MHKcuyAhTOCT/sHO
LZEbeyqd6bY6BQ9KMRDQVRYYphpHYtdmZdIH5wMoahOfK8ZBPUie441AeVW1qVgBfu2PAi5chwLe
rDd0hpLbw1oD1g/9JxD6deh7ltULe69xRuvXM2i6GyaKtpa9A1dLcd1+ZI37TNrZDcQDV6tZ5/bL
dgIY2hoDoV761Vl6jfDTuWQnUymKLM/+FuSdMArzgHOEflsq5GRGkVimYt3dd86iFB12QKhz+cBR
LXh8HHkse80qdkUKvzn+y/ozQWe0+L0RzSc7o3QrnptFlVX8fDOo/XAGTSQ66Pep3gf6ccunOgRV
934V06Q6BjIY3jhnq30dX7KKDCrKYAUm+gB5eV5OWDUPZdjVvkNh0s/ZxwhvrMDbwVOiPkS0nDVg
zBmxd+JdLKZ2+67Tl611e95VwrFmkTQYkj7djnN4KYF03BqPqSSx9Bce32IKmRSyPTEWXNR1Y1fh
7xe2x+StM1GzBKoLQKCETMFyhHUV5zhd/slhOVqSDFJ6YHysyTli4pCuB1LUi6LbBP9BVG5kn666
H9dunNr4zbAAnaOQLIDoq3r7b/VAznbXPz+AWGlF1nsZwCIRHX3eoz3aGuciA4jAO9V/tTidJhFr
5GWBnzyqaAXbvhnRlA23G7UAfIGPzcRPR4hEdvppyaqDJ7AUVDP2DIiVEzLQ/mpmSRg0lA+xbUmx
C139FJAXHb0Q0weyffMIp7t7Mc+SmfetKKbsRNPLgL8hcNGihuTD/eJKVfvEL7KA/NLqzGODXhvp
DZGmCWmOdsvyNZc6trcpD5G0wyNE87JOipv/yEHEJWDvc8HcIHjEkyxoQ39IQiqoBYzrYYXLJ4fG
7kLgXoIqeurBgPywS5ptDBMIuFF4DRvCpuml857VvJWBfGPAO6vEwZjTmUKruzlTh3TBKHeP5GCL
fUzr815Yd0eNKV4OZZxkTUUqkgj0oMuX6BJj6Jrf6Gf1XlERQ1ZwbzxZjPy41rxI3P0tG35sC4e7
DPeXKlLMn51ZR9J8rr+CSv/jNZec8W7GQEky09oOiIA4S8TNImSP3+SX22yFQnSsUfT90g3sEUmo
sHfdaankzLPmIJyortfx+fg5DZwXQxjgJxX6HJARAuu8VpaCfYvf554+knm0S0/bnHXxtPPQt/Qh
T1k9mgajF4CKM34eKUWo+UjKIQAE2E2Vzxnbo8cjqG4jyf3NGEtq6RoBmcqAU2EfE0piJl7HFyRA
zJ0ZI9/rWMlRaK9/fQYN3CVoS/SMQ68wYNOpy0bJpkUYvwWnXZ8tEWR93VYdtxf9wFp7nrwCRbA3
4qHbXP/IDuV7ysAL6feNsCHq1aSIwIAFbjpWfHwF/n55A0TP3OsbeXtx5k8U2Z6JuO6PiF+QjgHi
cl7D+xG0x5AZZHPAltUasoRdmmmIj3k2ElCoBwTj4FrOnI8seCr7F7i0TNb7SMLeiEy2RQyNJXem
C4ZdaeVSthRi2kKCDEmdaVRPyHeRAJpkYcCN5FQG496g8yBxAMAaIJQ+G0axAYE2fsBp1tilq14i
TvU1xdD+Bn6NDQhUCuOr8e913NpbdkBnCB5fm35QvjTabJQALJj9c7mUo2TeFSxCK+mvjPUcjnDj
YHYMaWuLJ9jvpVswYxsgOi15RqCCOf2WmXgi8KNIOIrU5EgOd8uE+RZqMjyVLrL62TW88e1yzOEo
Q3jYNKNrDo7Jg1+WFBaizX7ql7JdFZIQopC61FjL0bVEyC42s3c1jsIvhxNSTCze/aQVav/Rw/sx
qyjGF4WFmYxrPTSuOUU2dOUdh0EJLM5M5jWbAhUCOQwGTHXa1FnTot0/vTP+vxYt1esKNHfFjeZs
brna4ca4tKBTm5JAeo6BSbDKZMF1GUQVsoX6HB5y6QuXHDOm7SeYNO27gs0MZWdDR04KJPyEgd67
WK/T2bCjPU71CpZZenNAgXcw6x9MgrIpCFp8vdyehKAsatww6l1Ttau31EL2l1wxFmvfgmBXl+AZ
ZIBW5DGmv8q3IZw0ZV4QKCiZZHgmZOl3B0rTN9uV+I6Qwsy29fEZA8a6W1HPai8ImFqx4wOp1e+t
K+Rio2Ibj1CTF/iajQoW090sY+UnVTds7QYAYGrmdMyj1QtoN4wBQPpMfIyKmeB4beCVtCYcETHF
BJ2Z9RZnBXmlcCCoi65a0KG3WrS4tLRd1AgOL0/SGfAZX+4G2nn06wYWOkrqGoPPo/DLy8mAjaa/
kBGAfiFIAUBmIO29XsKdhbPdXtxrgvYqgOJsPi3l9lgxqfPnn8ZnQ6q5Ta+cFYnj2/nfod5EJUdR
LqvzpnhLw9N0aFpW6jP61585inPklpjeE5+4Q8kfRZ5lNVrQVuMxg50+F2MWDlgR0c2yl51ohY3z
ZIxGNIRujLnamxRfuXeXgeJvcTaf8B+72LdUJHo+OaV558DA6eHhS6u1eXljb7fBrJOlrTEeUWMp
G9G97lmGh/KJ2+L5int80bDGGvHryubrUaaMVLloZLSbrSywK4j+mQ0oWsNQK22wSaIXVxx2gPrQ
TS1Lm5TvuuNva6hr/jB+4MAU5c8DdekjzWno3vgtHgd5jtZNxe++UZUbEk4Zcp9g7Eku7jLwl6Qb
h7FcdkCm2nzb1z4PsdX31whYJUV5weKWGOBJimTkf36/aEun8aGeXqSDcVOieLZRbZObaQroZrIR
mUf3S0zRAZAN4VzTMiC5gxZvT7dcMQb4eafK1rAYhIZ91X77JjOa/xCsYHWbNhTWJ20wq63ajS6A
JOBMK1jrjuhzh7xBoYzemodPK62GX/vvlW6uia2xmEiGqLXZPUEX3J9b6rAbyGZcf5wV4N/NBhD7
4HRVUT3EDhW1LzVJvb7bNa1AusIDE27o+7a+A2Tan2SmfjMmJYs/zN6WaNrBUt1xJlc6Ktba9ite
xe4/LFPJVrUB+81Boq+Xwkze2X4hGEcbbRkyZbC7Ms/C/EJRVTRe5h/3OPevSZXt3KcWZAKfEQN+
oRhLHcVf0pKpXsoCDSqlIaBM3eBApTEX5C7lmNYxUt8Su8FSd1rHVTJTQ6NibYuL87iKPxXww2HN
8SLSItEojdwM8juhadqg/4aLQmHGyJYVt1wxXubLdcj00vuiea0nDhSFfYAVSBSnThyXIR+/l7FE
jqU8IU1O/1ilpxJKrw3TghX+7JCW6PW5lbY+PEGxNguPJuRrT72oc2ryp8niydSPAoZ3a94si2fx
GFipfC+MyCfIec/HhVAjI/I3fYM3O756ww07Ng4RhTiEqGnsDtd0oeO2G+WGWdAEp+c8IR/oKvnI
6osqLmJuqBkS5QKWRA2/U4RnsbKQoBRzS6ykLk9BSVh4x3hj37fOkPtUEgUzA8BafBTJggmJEnXL
t7cttzcCwra/mp0xWDR+EeksghQ/yKYtsLSqQvPLR+5eHnmelrfE08VeieRc8RgueCiMcSeZ36cU
Ibo1KN5mQzUrAYbncR8ltHN7CW6lEUxLtoMPPL1vtA5GdEbS1FtL7kgApIsf+hF4odc245REUZJp
oWg5UBdSAtMq+RJNvV0hoyDIrjApyFYCtsZedgBBc5FrWfJiDjwlq27Lj2vFPMEcq7EFayCi1y56
0Ldg5Yt4lp1woN7FxRXOCPbqyGW3lgbMoyf82WIShE0dF2bm8RzRfX369eHdXVj36a0zVB6c2Sfw
8313648xU5xyl+2x7eWMyEkzcxMOKvzD88J45x/AjcwBtji2jtyxRH1VcUBsjfkZDEBICazp39PP
teCo73wsmgIW48UEL18cYx4DJjd5vrm3YXkuSAVj/C7q9XjoMT0bppFhE2mOgsxJVeJlxJx3C7O9
hzhDWjeBdZ/9/1MGRDeK76FvZFszM5Ip58R8eryg7OBzt74Og197tyJnH6Rxp4J27SzrEBvrrXDr
mwRpgRGvYCti4d4SDNnlRHMMr9gwsxHPTrTPjMM7HxKoTk/6xMWOuAtzpFTPMs1BXf1sOq8/zfOm
49a6Ak+p4Y6nKirvG0KEcpDlAu2vD8Dy7IbX3dL8L3CSQsXT5hBIlVRzgSahZn5ohviS518EqTpV
lMKOLEoONCFKK8pv3RLpYnqAgMlOjc9uGD8mI8uatI+SWNoJ1SSsMy9vrFhfgDCMfXPAMl0YcMyg
Lyz8sd18kD3KfqpMsz+iMaGtsnNMeSoofPPe4phB6ii84o0JCRUIXgZ7/O3RReQE4ceff1F5weGG
c4ocxr+hiEiMkJUsStMqwZCRAn2QftGKEL8d71rRn/GJ1tJ7tSwNjImKbN+JBNePACdFvYjtf1Ii
ZDqa2hhcp4gG0L5CLsPha6CU2mPt//1QyV67LM8uPXUPJw1P4rAjBjt9Y3Jd9VIn+Rc4256DVZ5o
38IRcqnc/3Q0jRb/He9NYdUPXwuyX5trJuxoFSFI+llLtQMR0akcBfn1H0L3liAIT6DfXa+6foFz
uG1PpPcAxK6ypSLOLIGwQ1bdHJvlGHcqninWktFEdXoIA2C4ubnHiuZLje95PuLgFxl6QiYeUEJG
y4cuqWPKjYck/iQj32Br/NRq+ppcG75EZJKVRVKK2zNxy8B8Rv22WCuNmI7vdNDA7qAfkY2o1q1q
QnN9qQ3ZovLjK59zGG1YmCm2gNfmHtsz1qnMXndu5kEsyvqaQxjgsJ4rPDuKPkUJS2DBn84gNVPw
Rf7KeAuSkvtbfXY9sqPk4RIWPmZKwDDuMSzYYvvp21bZup1VEdyC4NswLeRpLEDb1+4k9estGzFP
ovigCxharp1Wz6Xaf2KQ4SJ0IRHZ5uMl1QfRN+rpwzjDvZiDCuAxdASZ9XccHHUoSEaMVXtKZ9Qa
BygCYRNCli2Gz0sY70nFMrTSJXucYTog8finuxcRjKOtRC7RWhSbEzvyyqGdwypb6bGeDlhBH/m4
sf6uk62gu1Iws4Xt2moD7gJQT26sg0xnOxWSjQVuhBG7RVE34sWxALxuS5CgebmNXOvzs8RGPMlv
nVMUoRrJASCX20ga00u0wZ8reuHgGfllEysMgGs1eJLmh9cxQw9e1Jj1rVqAPrYpBYNm9KyAROc1
H8KAwcx3UZW3xPUHONlQUhIYMssaFjUOkK0eIAGvpfazf+iiFl6zhEWHsPpDODZMXyBkIz+bxG+U
IuVXbmCq7rdHkBU1mjSoaPxqd2hj291uziATYxv+D0qakvczYk41zkRtZiNjx83+FQpDtpCOt5TP
asHe+sUgYfbruBm8WA1vFyHKbHXi7G0oFFz8RzJrCZj8cQH3ohfAMz/WkHn/1uvW6z8r5CLSCpP4
FxlRbh4bv2A0KtNXEjVurworAArfMrJjYPGqePWdVpO5wbupX+3C0oFeDafyFbaZQ58FXPgBva/c
zCscTxzH6hnEzM2Kns5yYDQu6cHaDB2ev3pGHS8wbfF3/AZcqIYgNW60uy4giXWcZdOc0Z6HwlUp
1jCZLZ/m9w2lvtSMMHc5N8SKYKHGsSEDCc9Wqu39+rKGrSiVuPVo5aQG2zCI5OVNWqAP3i+azVPB
WPY/T5iH90DMIaZFU9Ed4jZ2T59RS3vfc1sQCKGAq/EYY6XCPcBPp0XofTt/rGpo0NSquvgz/LvW
sJTw6slStxXllEkHfa7yccfwuYaVo+8RAM4w30Gl+5OLdb/nU14HrermuuW4KjU51Exilb5pkyNJ
dJ9LNLnOZwoEjBCFYXolkieWduYvi0NNK9c5APrQggtvJTHUZFlSmpmCBqIE+HzgZggeIi6T9vJ/
cuj4IdY0XTcnunPdOX/5cLi2n7Z+E6xs1vLde/pMUDR6Q2zKHaIrKtNWpBueeEyky9XawlTos1I9
FGwcRQX7UndfsbnkAqBEivgqxeP6ktWSaJuSFYy1AElpd5nuFDyaiRstnK9p7qTkDVZrwNintORU
2q9Nut94DA5rWxuPw3EAdCrmlV8HkBVyq/MQGWEwScy2mYZdBrxO0gqIHUnN5T5q79mP1KhhjRxu
V9o4raWphVgX6soklH1PWAax7bs3j0ikgSNAc+depoDu+vn/qbnUT49HbWRDoLpzKpQMKwp/dwA9
10z0UiikcTiRuVhvd9Rkdg/TMQh0N0n6MxUl5Ait2OSMGkR/v5Nvaau0Y/YFZ7khaLOLlIXX8xCa
CQQ9xMJlX0uUCoP2HxKKl2UCMIhf83nGDvLUwrS7QnYVQEfL6btqgdtYST05MUjABsWT8VNt20yW
YPhU1qraBBhDrW4w6KXWGVDGNfDmkBhKKNMg6EMIPZbT2GDcAE8RRNLuSj9sZWYtZKi2s/yOJYcF
Pd8aU/UL4zO2cjTZJStmpSdkMhLywRzf9mkOGCDG3mAkwq3ipCSXf4yIxGlhdKVOhN4nbGTebk77
pBX/HLMCMLaLvW4qffMgmKdprdNG8A9X8iXjiBPcy9lzB9jfE6OLFPafJN+7mvp/6aWY2vAYVUhU
KuA4hHcE2RyZiZEzaiC017X2CPMhFvFrxfzmjZPCo1cRkK1bcZ2bki2xxNhfnSizEs7BRk8HdXnv
yiAYbjwSRN8/ZcYhEEaxZ67HiDpTuT8l37Mt7seGxZ9RO+H7CwDY+RCWqzi9gxpwsDrVkXr0sWac
RpVU4T82DgT37VDeGY6PzFUbfoikZaOw8pHn2BOCxhRVxMUxX0LF/q6SmovAMZAfSXgI99xMwUt8
TeT5uJ/vpJT0U8gUxI/1mwrcPwin85mwc4XV7dasUdwHmbTKdBtcy9bAadd3TKJIG/MmRVIf/6Mt
oxkbdeMl5JGdohpeoov9kRPxyzbSb+H708+pa865/Ix3ZN/x7wu2AJNwoEG6LUaknHtiPLm/LgQL
v9DaVCQFNSjAHMFS/ZJWyTyFSwxTh4kEHDU//uy9KNabFVxwN75nLmzua1qC//3rrL0KwCvGl9T8
f15pZkfJMHTs3jetKfkzyjt9OZu+Uo/7VdSfwDjplyJ5vn5R23TCJWBYgljX+Gm60/Ely914R0oA
LIFxiYGEnVgZM2AWN6rPu9tVeGWmk590lo3ANZ0wbX+NnkZrsKb+2mFTqqXuMImA0epr93DaKzQA
nuqjNPfNeGoObD7O6TbuwTB3fvd7vtruvmYxWCsbEY5T8MJQvz7VFIe/T0nHDxeNoXhxa2elTwZY
1LOJTcG9l82GERGVNg+XtoaKJdRuSAfLR37GkrEFFolAz4Ev9Y0mSUAoIgiEaJT6mnN7MyuxSdLG
7Y0+IkNX0uSPXdrlMqFDn6BOrSLlyz0yV+HeGsmbQu0b5qQDzjDCAFa/ik2z3P0jQVb2jVtHABfU
pyA+koma28mg3V9oCcCxhE9J1JY5SrGoUp3myyXFuam/3dydd+zIFmwIuYo65ZhX9Q57Zvl6FRCN
0dgY8JnA/074p8Mo6o7g63hBMcsDRJla2sR59K2vhTwutoflpB2N+o7q8Dkwoq/nH6WRtvttODFw
WCO3n4NtsJDCuOpfKTXg1hBRVe9DlIX7hxWOpOMNfAYbJxdQQoJnNizY8ZM0xaQbjROJ8C9Q3bkK
qutfX10Sd+BMZvx4Uy0hqrZdMwMGDkAKq0gWUa+cqlI5lNX7PZi7bsg5yQQK+Lqja47z025OmpUq
y803O8ndvUNaZVzEWlHSRZq0sMyG5qEw/KMaZO2wolPSvKw4Q8pmygBR9nwaZaDBHIElk0Z3gffH
B//HytePlvjCCtIuv50Ha+Bqgnkgxi9P9yOt7i0JAWwpVmxlglG4eCuvN1ulWKDy5jMBShikSD6Y
OGmw4yK18/2g8KfJ3iAPIfuN6Qy0vPXw0z0XP3kCV6o4Ykfn0/yna1qrS67NOLd+hadK0LHmbbRi
+rUv7Afxzr0Z1GZ1/KhNA8V+6uH4L3MeDw6PcfqrJWpBA96ZwgGNmOffRoWHJZNURKwGIMAyWwHU
mddPgnHCEmOxGuiNimhy/GBYy7ChvTa0v/SYFY4lk3EzCwV75aPM2qsdeoZrqlgIQvwkvaBrGgRF
n4q4hrPw53+tH8ryG6tprcQQ1T3uw24bv29hym6bOL1YZJFPI8T0JjYezZQA5gtY+NWUXg+RtPQL
oNVaMFG2Wq/uPljN6cXKUi3RrXFv0A0pno3CLOq8IwuA2Z3gE1FrJl/mg6XoZ5ukQWMsoTg+iJma
ieV3IZC/yEUu7CMOnUmFxIwCHg14PxC9GfhKxApGQWibpC/WjBiriQbQ3QoZNdFecvxbQ8piCneg
2guj3LcFkwd5E3S2QS2PhLsOCkEBP8tfpE4buENY5xWpHJRi6GalVIlMvpI8YHkyp75m/6pX24RY
dMzXn8Y5Vkjmv198jZ4W3qI8sq7ABxzhaCcA+N1RFC7eDXnw2q1OwD8mpTuSj4PV5sTiDEj+33gn
ad4ZrwSuc8itROwSYWqE3462xlff7LDTekqL1Ed+KVwueC+gXn98vnUtYfzLKLpHaibMLp/9GF/Z
hIjSsharvIJpcUGYvGiC30GM3ihzSvBO/DV/UVR31QvX/Tc5YoyaYVn56hcJacweCQhtoAd05gW6
hrEABYrxg7nAltez6v/o7m8Ke2r69qbixh+IV9AnfislEv2qCiFvE4uNkflrX5b5sIZpWSX4zGuB
tDXNu3ZgzDk8pWEyRSFe2l+7be/Z2PdN7f6ay60OxAmGfmvVr+nNLU0b0prUZo/eKo8hIM6CHt3G
sUwHeZH5/Bwxs/LR7+kdtUjhJhgjwsjwlNOutT6XuYP3HJNviotvZUIuCwsgK4wU35fPBb2+lRmF
TfTna8UpnAaNvb8MfGypJWZSqP171K3WbNmug+wLuA+xO8ySO9bOaZ72uPzx+KR7XEIqxJZ5hPrX
8mxJTNBX8lvAVP0giDMOowEZdfHRelx1IK7XgzQSdtIWK8VtMGiUQESBepcEIUPH92vDgyV95vZd
8UQooTkYjGP9Q+Gnch/2ZRuz0odYhKuPH4bpQdfHqM/qXB2NEvg0Jl+qi6QXeVvmeFvxmdXlSREM
IIGK5xV97KvJf793pRUgqxzkeqE2rsgTcPD5IH+YV19KaavMsCiAYy4IQD2N2lpSMkXw8l5eEAob
2Quf/xwBh5eIdaQ7HZ5V5VvqCsMQiK3zLCYOpviwyNbtjGeQJormtpUuRAZh/DVAJJZ07KH4cR5P
/n/b/hFEdngZVXip5jHn9pfF+2jXsvqkhK2k3T3a4NhOzEkJoBkaBebq6V6tDTGJWvs1+vs6LpNa
lqh8YNdOVO2UGH8hIBWzMwaFxipsLEHSeM+fAsLIc9vZ/golJ9YlNqcuO//vRHcxMZNIJpKjF9cL
Ac1NWfjUK2m6D28hzfimXASuTp2hD/3EJOA26/qXrN/k5Zc81HebCxwL3lurINqOwv3QX/yqu2iN
8yVt3EgHTdQWfKjbT0vogpi4Bzw7Kw38kcINgcCMT9ByvTbSKQ3O+A4o751jNgjHA6n39Tj2F804
iqUY+VP+W03J9yN9nsU48XYQvTF9qCqnNQ7A8NHIh08+ll6pWDgKxabbj/wWCpaGVNnca0eVVu2Z
rB5nGK38ckb3piwlHNnNcGkwWulIcFLACUORLyEUORUPDDUu+GBuyZuvpNeCoAZk/dTEBxQKbdCn
Im+SaP/2JZd95kc1g8KTh78njv2pd3evp+61c14XFtAOG1vFJt5cA04C9w0yGhB202Ck5IN7dwP3
75uoYIpz3xZebI8H8GXARV2pAXYgwTt/2jynOjzXXlO/RilUcWUud9tt9C7tgjCvczUEKw+xC9n9
mjFPiDnRg/6TjxzGqQMOqQSP5knBm8gosJh7x0FbPMbXF+3yXttHw4gj/94bv6chJrAmNIvhzxX9
LWyhoIIbBc9nKKd4OT51FYH+ICEqF7YVIsflirFkOzLaKbdnP4rrxc9MJL1Xmj4lPInlOg1p1BUG
J9UDaD5LXAeohyB4b2lZaVAF4vaW20rQKQtv0MuuzRz2s7rqwTdKwpsqUrIHdFTsmS4vyJqWIKZT
MIJooJ3u6TuyZTFTw1Hn2whTLlfbm7MSNBArhMYDzqpxqxLxx48Ptz0nxh4rr5/rnuUOv54U56dd
FYkxOCObt5fmlBW/rtSa/ixtUpLGRomBPRhvmQzWH7mC1VCGZK5v6u1BZMrdwzgURmg2Ow0PsRea
Jmtb+pnGJLwzTykbcrGmSSZ2tj0/4E9ooWe3Im2Mag/HVzZeRCtwisAOtVSjGZ3TOrgmsLGWXAyg
E9NsdUjreZbWqKUvz3idoi4WU6AeVZytAnozlg0oxgTEamZzvrbZrceMfnMxvJ40psxRt4V1PWfk
YQqPvyBjnAPT4yuUBmqkdN01Fb7/jX5rVZBZFp6qwvAIz3sdQQ3a12YoirgOb3uZXsYzETP6GOId
AwRoQ4HhlpraVDvq0x+rKAUgebNF2VELUC/b/tb9KKXSPFDpCQxIwlEnXIRLXogr1Hp//wXUzVt+
sguIzeDZEWSrnEeDK5gPMA2zprPpxY2nZXzD1BzvSNZtYn63ys6XJPbNTQm5QxA78IMq7TMlxBxj
D4PWuK4SyWUap+9YFAjnbnnuFc+1tXILkB98ZU7Uy04nqoOfeUkAedxEaZ2ZxaC6MUbn1UDBwcX8
n1M9F6lAEsAEl9HVA9nTSabFblXuLpWDjOA5EdM40oNJh0bhKwzh5AstuYlz6bdw1TTIf8MYPv55
7Bp5TUw8C7+dvdbOvblJ0jtRVA5+WsXxJJ31ODdmSJnsE+VQleIDks5AJ9tcTGHzWltG0/p7v7H7
TwIFblONaVhnBtN3YthQSwVewdLmXHjryECq40JMVw106QL3ypeSYhyYvNYeJl7mN2lNDA4Zsd5P
S7sQNQZ+Fl7DiUJQmOEtNujjzmNA/CurizUE1bIgrzxVhIn/1hBWL2Jlosy1DlG2cX1n8I5z62pH
sMP47W/4ty91rCLjxiGoj5RLbhz0qx+bml8jQ+ydGSCGXhxpRS3lHWc/nM3IdzvPx1BXP5sN4Vc9
UrOGAn6rxDyacy49cEQOqRmJtDpCf4P6cZPux+SQ4ZuLxEfPyifVjN+JkpQnORpo83656+lZPHqg
ldkyP2tyAn8ex1t9N97QQFlUUSqzCAmb7oK5DLLuZYSJYB+iOOmkrCAPOPOJItlKRSTbd4gknJY5
i0zFkQz7ouIfRzL3Z64OKwjTi9TsqvreCRGEUJr71BvwrFeCgkkoRaW6BfIFOpWL6cUrOjnYnieU
GUAk5V7O+JPP63aH1ojcUwJLNAmnkd3+rdw0WXbuFLKM/Idas5ja/pYxeZ5zxCslQU/KvCSHLIWo
RZjZTEPE//gH9XRyLcgU3HIv+zMaUUNzeZM6E4etuq3DVzHIIPSTSZQcxWP9WUFh2qFvS+Z3Ilfi
zMJznpWi/C/7qC3Qxx1fr/9L3rDz6GiGD9VA7x0Zi9LE2/1qBLo23NsKpthiikSDII+Zfnwq1YiZ
O8eX9T0Jq1GlLWbFJ6MdaBoXhL8bLcCaocI0u0JemKzX+vWqdvQbYGY2nHwRpwbf7nRLR0YWmvIP
lwYz+mx41y3C20hCVKb4RuSq88TFE+qBmxGxL+odh0WF0mzVc4u1TUWx1IspxAZgN0BkMlOHW07E
HS1NKEuQWaIbS77g+aJF2els4XZs5roU7GO4eHj3j+nKs4hqPRG//mAKVjPkKnyrYTV1Hi4ZXOnt
IPcp6mkFmqhtXap9b/Y4f+bqBffp/zux3LWij4TNgwLaSv23C/hoPjRDsCEziHamV/2mvMjlgBEk
XXtBhdAObultrZFqbxnl1JaB5EG+MdYLtog/Jt025jxkj1IBw0sIajVBJKpuLGATxNgw8Ik7fqLH
uv2aUothR7TT4knGKk8P+4nokUdoP3cxuhr6l+FC6QzkHy36YMeNBIgAoEz8UNXZs036IR8NmL0V
ODKfEcE7hilIid3ssSO0pd9H7BCRW+B6QOrqETakGLG4k8/CmxnnZoTer1uHzPCJtII8j1NJGvDi
4P2J4fR0rXK9p44WKgUKFBlp6YXSPWZp8EUd/lFRXyfPhXejGUWGax9cFfMOeJ1G2C3T/VxWX+hE
sAcTwNeZumqDk9oGhovoATzDQtNoYuO789dq67RgyuPDo/ZM7ys3nafC+yyGyymdlVyBN92z1fqy
s+BzM2KLLhqUqI7bODdnQr2zIk5eYDx+ugxFFEw9JFeRvbtZMXysmDCBc/gsbqN2K141G/qyiz45
MfcupTZtvhLZcfVHwlc1A/5cD9aoqnQySZKd50XPrM1ol+mtwRAtxK+lSAv3/7R14xwBQD7lS9A9
A+nILi23v2IaOfpbhOUejcnhxlxMf6ZjJsW5zI1X+yjbExf0TR+N4wDYcZYetPb/Ru1XZo3SLpeQ
TjS6/zB67NqJ2C0VJQefyO2TD7Sv4wjgomUYHO2eGl0itWfnCTSDPFYa9XXuG5On0A3Ov8SgUtbo
ek5fB6Gnve39OjGYB9OO5uzB3uQDMzMobFeD83kqqJUYtE2CwRrIHS1z0tE2MJRqQFnQf7cw0IIQ
VEJqn+6e/mfJUwKl8+8T/YWxrqINtHRINU+OCMOtyx1uY/FY0lOBKGTknIGMglEsFlyBBQmWDUwS
01Z4rumMWGZ30xv7OE1IkrxE5jEGDroQHd7vVwjWhWx9LleUnDWDQQlkDSchPFEKaFe2xGuOp9ww
sd4nYi4jSKjhX2ouCF4JcnWJa29UTGU9LgD3TaBnwhy9Wzh9hWKkWTDOHo6vVJZQ6w0/zdu6lLrF
9zkIo2BppN0yEshN1WrzD8MU4N1cha75uVIdkpS85jwa5FBlUL/vjsb4IVCVRTL4UB4eQgfGrMnK
RHq2euyClnpm+rM71SIxtDnpDAwEAQf/7oHGTh3niLTJVB+1EU17ODYJKwrPnx+VH+T4as2B0HLG
2ypaP1zZWqYjZ4soSKd7iosdtygc79n7FLZpN4tdLTSNgEzlSW+m/BxAv14BhojlTXeMeNCnSNv2
JeYhBkp7H+EBOauRANTIbBZU7ceYnn4L+kxHmnrxN5lsu5utaMwwbkrfqORC3aRIzMJpDrOIbBss
9mPxJcYPUufnOL/AIW6i/UVd0Pd/muHUNNcxyQiueNfTTgVbQ2Vyz6hDHGUySdEa5J0vEVVQia9+
Z0lHKwdTgz61XXUmcIG3GlmVAKGVK33JwNX1L6yV9W1itkOPbKKISUFdQL9HqULYVt8h8tAmRGyi
3COrITvCiTLcPCg13zOxfksABQQub39rVI2w55vJ9Mmvv0kvpkGZ3jtVYsJ1p1zJ/h0It7FtQ+di
iRyVUMqW9x2DTcy3I49QUNniP2E7vqX8gaY15+v8JjXznpwxaCJTm8/k3/sSLt7zE5tDWm2SluFa
/sCpRX+VGsX5CB4JSdcvGjDNDQZrEu15WR5dIa1HS428lTYnGAu5TPSFn+JJ5g/3//fzyIBQPfsG
Q+QxZaAoRi8Uwd6EoR+htUFjA4vwZcl0foZQcsWE5XCIznZk0kkhYTiDnGFa5FG6CYMWikA0fRWC
4cF8Qp/OoOWdVntOR5hpy5U1+RhrfiQOrk5AZNUeQTxD2DKTJGH/Yw39gcgZUKHszIkqIqzaXNPM
UVK9j5lKOWObehkCeyq09jqJM5ooZvERxUXKloZpPuD8lQD8oWvhqbXWpERO8KT47DIJz7WwNxRC
pPhAiouFg8Rezu/pIRq1NE576ZUknkIMFQBrlFdRVUGijKg3e9AoS+qYeNNs8FaZLjZK9ZoDcVK1
JZagZyB8nxJPebXfIRkns4SemtGngLXNDfCNlPDUIKMrejOKofrYB397FJ1whzgKc8xDWuypG5Sw
/o6TLkucs2Kd0/wsm8z56rLzHVzss4+my5d5GEQPAHCp1nm/lcCNubRILnKs7A3cGhafoI1EWt6v
CdtPL0pV8X2JV5RVFvtS/1FjHGOeCiqKYVUTvvGmgSnV5nkagYBVWwrgo9F+NOfvZ735+l5i1P4u
DKEAv3YwPGYU6XtJEHggL5FEftleliwr+WjTn3524SvaffkB+2nPeN+3tRNyRlKWmtv2LhynF4eu
VOLAmim1Pl+2+gU2VEFqJ8Jb629EkCX7HC3CVnLOOmbdc5VLMdGcVQwmQAyET1g989CHtPRzXlx3
kGZHy6VqNEn/tk1gIq6MzrSkhVF+9knhmzVqTiHw51Xj5PvsINmX8Z/0qwv2BQbSztenQCsE7fD4
k9uqokZcIEL+C4nUEXagcclHOC/IpodDW2q1SmpozITSZVBRze2Yk2FislQSOp2rFmWmbeM8FvSs
2foCZsWQL/yVr3gvcXoWCoMdgMaFbjJMgsfJr2dARUJk/jed4YFdKFxT8E6lxQ062pyOyyfhnHyb
bq1mrd1Iuw0viyrGBEiHXyKCnF1Fn8eD//e64JPMyMxruxV/WVNnUsvCy1/mBaX4enm3teypTuSD
19aUjJ18NelJ7gAsRXp0FzBNmK1nIlQk83P6nF29edGR+M2C6y5RhnxdFrDBjyQbLJYfgxguqoW3
O/K+9YIPaaxn00GP2LHCBOn5H33pj7AqGcVNajsOs1Q+7FAIRXnfvE2thkeQvSkVXdbCYN/+4Ql/
fyit623sM6ZTrjAqj6ND+3Z7bdciSR42WY6RF/KzypV0WQgFtRy96HGS+UqOnbUHyf0P5TyYr3Mi
WFp/C1ZPeUq1IFPXie4CchYqV7K4CeMh5P3qnhDOSxtQO113RoR4J9N/ap3RADPH5fERS2lPbcWx
cEs1r6JGmQrAAeNzH55tNM9z9mk5/PqpQeYn+Dte3OThiclRDwd2VFb+00yzqsk0Myge/If+RrMc
M9kSyd2LNi+pcY1DuG0n02YrBVUyIKnJB8CukDisOGIb9VkMNqHkwyeUQWtYj2TaMxxwF9EIAOxK
LjlEhBQXI68AQ7mY7gjX83FXNDj3s79VH6k7m9FQ7jvkznrsXucOKXGIla43mOKrz7yXmr1Gykpv
gL8toC3hdgO6mLxJcflNFqGtF6Ko0HlNecNQ1PBG57TxJiQbYB4K2uDzsHC+0XqxUduCtURM46kh
HeP2ADujDcfC0S3Im+etQOvbJ79UtKpEXSHlmaYfSUsxdvcPmdbC8FyjsX5q+u63HpXwO0wgxVgY
bVvvVLKTwPtUH+wWESRLjsY5WDSiFTXldeBTkh8aoMc0NHcPw4Xh7XDS62bx5Hj+2aqiHDICNwzC
dpfpHWUp+V3/5bXjvMz+w0ZiXeXO0Iky900fggBUXzkoPSatl5Q+7DxrSdd24kbbNHu/gAjFFqz+
Z1vZYuR71FCpIzgXkHp3qT7gsKlfGlcLCpbZ2SY2z/nN+8HyaihIAPWcNSvzIebhDBNQnIGSBXHJ
+sF+xT7B0fz83ExX3DFijvVg7V6tQcnoVkqipIviLgK8QYR+7aWTOgpcq0OQkjjbPEGhzu7LwA7l
6AimE2MYDQrUd+OUGRrI+V1qVXjihpqFpbC+7WSk/eHQj2WE5PA0jZuobsZH+3WXt8dhCCSw+Gk4
6S7uFtHrweLEq71gGwpM637Cv23BQjMjVzK/vjaYMpm8Akc5GRmst0XM/+u7kbp1ODBrs2XKP4xt
Jc2HNlzBRgxRTk0rEcVZjDlGFuWzAAJTb/I36iNeLwH1Cvf4lkQPnlrDXRGjJUurQ6haJ1a3EBiu
JE+H95jkrpYgEtRa+fNYTbcYHvPLA0YQEbX19ib+upcQdZLx+BziHctImD4diNMS0ulMQYB6Xbdp
7oJrp1uX7XrlGeWdc5JetUDOJwptaVmbH10fnNXOtsjS29A3ElbMAV4OUIaJqY4l5lX53WKZiZA4
pwFQpVmxw5h82Ox4jw2RGM1Z7/Jt5VhuYT4Auu9cLHPQ7QQXOwFOQkD7n4f0kHgYc5wzfszQMHoT
9oE5eOVJB8fJokPiizKM3GRHnTbdwNEVAedBmn679GWZWyMFyCYFI08kDfqVbRzTSN5U1rtAeloB
JX9k2RBx02AM9mv3Frm0pK9fx4MQqA3mxUobzjd0ndHdiho8Q99XryQ3YG2odvWz8phxmboUgPCm
eNxiDo4KpKezKt/cEgvFuL7QWDGaDgGxYzIxVZ7/ku3MGy5jU4KCtPx2Y+GnDi9DBkomUSHz3LEb
Yc1uIQ9WfzT1lf10ZzjEWExOOBFEgdpHvOfm9IuRg8ZVqSh5EwZua+/XRze17ubh+AnZZDfOLAVV
gtIdhHhOtelAjHIyu5ewTaKoj+S++sqgmVVzMRZY2w9DjfCQcI+/1GVa9oQK5RG3y2jjgbhpd4YD
SDkyM2DyCE568aoSL5DnbIrUL2LMpPBIkYtKLiCeVEivLrqpNmV/srGs5Ixm2h+r5/uf20Kfb5rl
bGKuHleQdgnc7/38kT01iC7NAaynqldKEazr7K1TyPDboExQnidfpi2RyyoQKMRBkkA8rmdru0k1
fNrZeF3xHSpgLS/FEpr7Z/xmfFXMaJUobY+ByX6CCprci7DZJbW9BqN7apDTbAejJEGUbst00rgt
F+Mw/7CdOXrH7Mm8tcj2cWj3gQp6HD8GKxhLnerxkOqRcmYerKDyCJIOARSYIJEn6kMhN17mRrk4
1nXYhWGgoXNT1EWdCNeNtbkGO9hwr/0vvne79s1MgQPJs9k144HFre2SHagVcU9TnVVd7CvibMab
3t/U9AA8zUQtzLWBbqObfiDWRUtGB8Aa0rr735+Nj9zfZLXokll2XW5r1CmE26ZBZ8OznuIbFPFI
RpZZ5JnR1lReQSzNL7fpPp8Wy+DawU4gTY8DrcMiijW6mPx0EQMogyBjG7pxAPqviRT0lnRgZJJC
MNlGUBb3Bhe4qNtZgoH5IKXzkhnHXKnCmjk3y3inLlHB1C/35FxL8ypPLC5sT87or+QcxakrNtum
EoGCQakpdHJOGLRiJWJ12xgmEJEMkpYif4WC/UqJgYjKfLEYIg5Mbc3tDW/xfdY0eb1f7U3HP6ra
c8mKN2H73UmicgIFDVkTAhJ9ZpYjylL594lF0XMqXGRvhYIzAjrg5nO/T2YdFSdOPmJZmHHR04O3
vzFQo1JFZPXwZm/0ZEsk2babtpwfsS411rg9z1B0tjelS1j7twPSPwlG4m4E0RRi49bSK/23+9md
2Q651sgTVXoLhhjPy2g8SJSGXvjEJkBBmeK5YuPVFbiiOgoXLW+1pnj3YD51lHRL9AcK5hEqUtzG
fBeGwERpr8OrTge1S+CCJ2U/QE70ANRBoHFvCGQhbIbHBARKSXY0eOmFD4IriQGNbMGoPtu6NVdz
erQkhYggdWa1Gj0g1A6kBv77GhbrcgvpPTa6ek2l+nKWK+/FsXFSpNW1AVQaZeo1eAtiMmnMmQAm
QrNhaXanDQgex7ChKsNDjPubxkNHUM8b4u/QRR6sP1xF4BVGQYlZp/FfiU7hHvUrboK2m57mqUmD
W+SlqtnPwu81S9MYhPxuepeuTrBWO65wexbD+SFa2ETiYMX8YdvOus/hZhy6dW9MGrJ2Zz6yUErw
qrdVyCdt6VOjkzaji9z9L56BhBlKYY4NbKVtJGxum5KB3tKJzugCNGikmnLrHASHiUdR+Yqw0v6R
9alUH3kELlcWUAAEJDdfLAW6eB1WE6b6Zcw+w1iRJI0xEbceITUsX2ZDMwQs+FZhK0SqcQb1NOE/
opJgJ2kVoxn8Ay4luUtUhjOrX+A7VgYQ9Z+9dnJzBDL+KRZ+i0bnWb6rQLQc9CG+wmY2EIseZvmC
W4TfDrHzwHizJgmcndF5hOepcGrcDoSYu+UTK71quShIZMr/cd1InPYrJrFDJ21SCznVNF0ctv45
z2iS7O5NTUB0OnlRmz4PLe/ATo3yo0Z0E7vKg0HfYcSh/jQWGiNaIXIIAeGEd8m0k2tFkD+U7BEQ
fDx723IG0w6qygdCUN6gQUjw3vbhqcjEHaIOW0BKnEa2xh5osKNXg05ltFasiomIcvBDnFzLcGTg
Ug0S8IopqfZdFEphKVhJ5QDJPYSDmktzPL2BmpBuC5qzxPcgZwDpMQGHAiinQ4zvgIthrTINAGlK
rwZ0XEqFcwRKFtmlVFl1ACFlqEjFLb9gRujp/cJa/Bvxd/rQxxH5RIRXW0YhbuxFNZ3kg0hKqyK9
Czx9OTBlHmORh3h6lnXApTt6heVa5J3uzZRRRYYcZelYIcROXvLEz6faQlJFqWhZqRsnpmSyb5TG
VEKBLrxjAnXaocCj8aepUpfRmaW2nVTvGW9pLvSNITQx/RQhCZQMt0StZge2UsMXvh+cGjRrqIqU
k6DJ8oNMHwRRpJ77LPzBs9U0CDSrJjxad32ACMU508J1Bsrm5kR6id+69s1xkQ3ti8iJNW5AUTKX
faUuqdTcbDMmT3cmwfcmzNvSybNtWKYA2wdm4CDVbWwVvZAPmO1U81+zFY7wj35/8YAHCI3ZZLyA
LxM/y0IJ/RyfFJ399KzgxJqtRLWyxhVxfqi9pr8Pm9tQhtIqUQne6Jw5q5VflJlY7ccQTDN/Gvg/
7UftzHTDkTr1BSSKvpzxKQkJND1e4hfy1MLknghAdht17JETNBHF2f3XbOPv7sxzaQFFQ6YH6TkJ
doAEoJ2BMGobu5ugws9sHP7MKc71YGmZfZnTPQ3iKJIXeqYNWV6UhLPgsDDysz1uLobBrhcgFUFS
fK3sTSwm9NiVhxhx4IMu0AYqdyTdCnGV+iZKpuuwEVcsD/+Py5QPwtulLi8gBJOKOfHOpebGAeB3
mQTfhXRflMGx7tK6iZmGaRg32x+Zg18eYUqXXeoMrBNUJgK3jtISsE7PHrVdRkWsGiwPbcblbzb2
gcZqZjfzHT4nxnLOZq2iH64a0zr5MSPECPOzHWNI4gdtRcmZI2/oT8H2Thr3u6LOVEK2oiBU/8m5
GIepQsFIk+iUjLu0hJ405j5UiHSawDVElto8NyQ3j/hhYX1XbDJyPiJauEPWphP/2XushWkUeTEC
oS8qgMlK5vQMD8+z8x8Rh5ilMq1ebllZT+cLo2AuTJEPnkSdBQ0O+jI4fdGBmjxx/An5DcvnQQLZ
nqB4soRWcdTWZ1PlasBbSW2/TG9boFdA5A4Swvu5oBEVS2514gLF0suhi8PpMwOoUk/BjJVWCMOL
kQHyZCcJ+G9cmOy/F8iIxLF3h/3CjU8OG5519D36MuzKWVyzXVQY/HdRxcNjgL0DXiy64Yj0UvfY
YmXmDz8Br3KRV+zMOrFNt6zpQB0tZG86s/ruzPOAaAwHaFtLiiuh6Zzn6Gm0If7uXuI7M/M2zjca
eIAsh6DmSXKtea9itoML9ao8gi7MKa+MmFiem0AkSPBNWLQsKomvGtQY8Bt5O68dJ+w32DfHR0j5
8D8ZZBH9EJMJrEbcL8lxfypnls2oFoQhpv826p8zZFCLDiQIObAUBvIp6OEm8CAiT0OU+MANVxxa
f9YZRUXGG5k+qa5Nzu1R8ScSZiT7y04N3edAdHMnYwPjpmLHpS+ctb01ozC3zML0y0qFI1K65Bkz
MQlGaKgZVaoNQRncY/VGjYyO2h/8ctz7GCJKjJ3WyAFASNds2HygYDUqbvpYXH1tkd28f88U6w0r
PiCeZimhyUMelhiKxtWJs5T6INL/BxLGSWFo2Q9SXsxd2oNIOE6VGfKgjJMjbyDRd38R6dXA4oHL
88e+mjAnHhcY7o11GaoYYmyUey5m8t+vlJO7ihfsQ64Hrf6VUcbqaqCozTIYu+OL6wq+ROADo0Hu
paG77uh5rQu3LE4hpas+GfvDAui23hRPlyMtw5xEf0kXoK4t5tXR5zOdNiUt9wB5rQJSkwPTZ9ZJ
yBS3Awg861tR7n7H8lc7oxF1DYRlGM0x624ToCbEijqaX77ATIkLJaEhDA3CYZ/pYXJNWuITdiF+
t+KRA6NGLQaPNsf6jEbmOns0ARh4P9y3dch9PnB9bqWo1FSsb9Ezd5+pvSrv3d62m/EpVCiuh/7+
qRKJadNMhMwy7mg470uSWDmNQwLwWiBrbK4vVr8UfKAuDSjciOniRc5wmK2Ts6HPYE0kZjEzDAkG
9AhJZb8n3w1i3cUyYb6k2MIwKvCkzMnlnG61XB9Hg6Aq2hna5TafJd75loqX/QykYI4xMpFOv0V6
kJKcfrRep/sbXjgzhrSFhVO4fce9E7D9Q+SY9g8gU59EMwzNNuJYo1IXR+KxwO1EodVWxKuDge75
1PCe8fbnAxu8WVCHTfTII9TnhgyQ+b1ADGtx7fwWC/51qlsQ+IBCPecRpaeieHsgxphK0ukMSzvj
jowW56hBVwqHfGSbG+DEWy6S9bkITBXXUSTeVnqea4nHYJlnyl2p99KTs6v//IviBHQAZ9IZPZOV
L7m8Iy89scqDHaArQ9bEveABxiwUA8bo/0RFznTN73WjT0/4RClhc4MSWdQG1A4TlzW0XdjjZ6tA
LrILMgtOyvIaeqqMDt7xBrEuo2L3druqf9FWJBot0K8REzSwhygvvWjhXKMfnyna9o2ATcP92GyV
i+JwpyM3kyQyzOlhrtvmwYh/ugih5JO9iqc44OhFmhxv1UdWNBoFQZAW6mSb0qyZtCbi8aU1pRAJ
TXHW/wCdgDth91XWre0fAHkcJ1TEGoiwywCYA8e0OosQtaBbcAlVGgfFWtbe7oQJLaZkOK0ldpYK
2Y8hE+pAxuPPGApYjcIzTnAQkO3Vo4Lj6A1XK7NBZeRa3alexwu1Cw9uOqdiuMUrwOjkvV5zlaLG
RKuwWm1dECsHYu2o0UiS2Gc8vWBJ9PfybdwnykS5bQN3VNwhc7z/Fq6yxjxGwn84Sv3HIh4Bc0pZ
eTYtP3F5bgwp875LGtt8fwTNapRReflaSJBtGREXdq0QXHvEDUqrUIZkpE6xpcTjVTcOuhNpWgj3
g5ALspnkGfXNhH1KGNXs4Cp/DO3o+/2ON772iWOoZHCarDqPF8ur+lVKHjQL46UeBuH7ecYqrYFm
AruYd+JLdS09re+UrcuNot9HaMBWLtqENg/ivWnyyr/W2CgJyFlb0Pv6DuWNKAQNWd0IiPADgQ4L
h+dJn43FZVqHTZamj+BSPYR7Co6qhP2zYGInqtFS6flhx+XNQhur1MOsXHrs7tG05VyHu/CDXPEu
O4FlMZ9G4vvcvgxBy5uG1LapgB44rV2fMEHwTDfB/86r39VcqfECItgP9IWjtpgHkvt6Z6WpntaK
Y9yTJd3EiOGSJRfg9v6b8m9l0DG0G2AfPM8eP1FSL97hCP4tUstiwvINEKmZ3N00tx5afj/YaTjU
BMxEgt0PF362LKsI+5DXlolZZZcRthmMI2vS3jnc4C25Y14ujTlqGhkkxwJxyKCF7ASpS7UfR7z+
wBpbdojpZBKdd6uni13xbXQqCK2QCL1diczU1IBHzEJjvbbplw4PWQ6Y18pBTUJXzojhNN74glLK
ychSPDYCgoiKFCXixjveDiT6LZDkpSJ6BFJlRj5EZb0oCi15Vu9SuscVWz9x0nATIGVIARa7cY4G
Qn6e1KN+Hy4SBARdmb9AYlB3499izgETCHGTmHqRT3aE2vJP3IPZ6/nJskPWCe8wGprvehyXMo1Z
g9vA6WpdMTDPli1J8g19AVEnC176/5MbNWosebREkWoVu32HX2JedFOSMKRibkiY0SZnoFVrXtfG
YqWjs9w7umYPvCIz4teNRn8BKi6+2506Oad5RHyQpz1O8brL8B8wCS3Al01EeboDfjJucAUq2yld
/fleGdG9hOm3yeFo3aFvs3TXXENdFWt3GJ9Bmh81o8R9oFSF89Chr86tYK2mMVgyQFgFkNbKbvCP
FEWqT/jgLxlk2drWZwh6kG6HLxTbGwqKf5M36HWnfwIJwZTj8xixnsi16fIyXr+gppH+R5psg60x
xcPdP15Nxduoks3J1/tXWih74AxKN7iY+tO+M6SAeeBT2ljlBXT/ZP8fE649TkaKdRgd4og/kYSU
5BIMqiNLfw8+q1kByPbmYHwA6QEq+UW6BgDSHMvp6Zv6PpjrOlHEEYjZUcI92kWRAcYrxmLXycEa
Hm5zfg7HJhW6aK1brB28Ouzl475ieJZLS/jW9ZXmCA/N+9OoE/gbInmdl7L0jjy4SD7lWsxk2gEX
peknloBQc7QRxkkciTzoSUzza6Hu0uSBSq3EIS4iEB2OWipSO+29/XANC0nzlrAlq+THdxKmChuA
xVJte+LGL3BBDWU4JwnYbo45KYIIuRIBnd14kTUf/y3VTdDmmZnBfh4XY/HmeeHNxn1ooSLHqx5c
GrbuzAcqG456Ych9Uq47+0Y/3VLVqULUV6s7XFMgZGdEMUxb3icb7w2V0rjbzZHYPrXtsSl3HsKw
sIq5GsPJEZ0Tgm6d99gHMDnG5HOJkSNvXegWhI2wGYpbNJDWEzA9QO+N1ZR64wbIt0mpbyfY8QRX
nEAKNEleDhnj97uiVzt11oSZPvV8UPilhnfAv3iqNvEhwSgs1KTdYHSzBThurJF12a3xTyBwkh/V
Zkg/oFJEqZ4RRmEQPIGihK9TPqr0Gg0DOIlMd/tr2Hoq3cndsJ/IhZNBK+5EqL53JQETtSINNpfG
Q76jDobUwqVE6gKq7K/mTECefB5wj0ObAkVkEN5ovXZejuis5uzDuu6alCxIWtcOZa8MRGNZBJFq
IWsEnER04SyQ6e8yukNovGWkWx06PgKfUARwe5PBb9b4fNG3IWqbg9u9cD8eV56wKgQJNqWaOUWI
W5CY7Fir8UUvwYwYNCexxIo8YU0oZYh153iP9KicACbuFiQwITc65BPyl3T2hfIvZ9odAN5BNNsb
IkzHN6WmpdqDwZ2mKw/J0AjqlgY+j+knpiBnB8tpLe8bdIg44a7qg6dZ3dqvik/IgX5PrvJZIBBv
fBMNhp/wlpUIV3Czj+HceJ8fXlDeRQ7hvpYqmPIXd5dLcZ+9CDeHdJ0devrBLvxztD0z9gHYksq0
E9v6gU52NVRwdwkmFkzhT+qxANmKUE6AsiPFukUCJmiOGgAg7Yt4htiyE3eTeXDWtm6daVvA0WV/
R865DmxHiDO1j2FjzsPi2A3endeD1DG/JOA6WGmBcvcpIIS63QGm9HY4viMmOjt8zlJl8gnkXgTE
OrQoztfdBm+oHWpINf7xjUOUHIO5xRRX1mYo2UH9NBJUX0ph+pf8IInAjDJBFJcBKyXXgtqO1JrU
78l3tPEZxfvAuJJAy5ySNYeM+xxYosRmAkpfDZV9GLIZyNxbuZJ3AEtdcJZnHWAJH+50OpA3RFPN
9PbhRdAhM8qwrDQhEO4/ygs6RiPj88mY8dL+yvJkxTwDeUYG2W0gadV7piv3+FEbBBU4zpMYS5WI
g3K9u03ZtypwH4A+IRl3QqI+2zJQstzzS647jaWViwYEHwNYkW//iDtP9AmLqgUa00lSetpUpM5/
W0HLKl5UAYO76X3U9WfoWqAjqvjvmIkdl+krIwQcfsvXFUI0PY2DoeC+vhk11Mg66nPB5+ARK/Bb
ONA1l83L+Qw+lChNt9zXayc0Mm3mxg7uVLbWtQk4EV+ORS/qFWwZQcOgqHkU7xW65s6c5gS3jjcF
imJx1v62UgkzTIazLLvBrT0NbO0Hv4CRzFQF0f5EP7AcCJEhxVz3ghXmvu+ha1BrdlXKKW8vO4oW
nYwAD6rCAoKcohZOeJOng+SmYleUDVssgGq1gid9UVBwNO8rxASKm90kx8vqfBezvnXJXiVkAAiy
DlJQBg1ahUc5ppmvkIaCX7DX5WAjQnsOK0OYLXepFInpwNcZuLFsXU/04J7Uu1oVpzhonw++KS3y
kn76aviqb2COg0SE/ObkpGAUDgRm0IGeHwlzN5VFoT/OUPnJR5xVOJ5Yzt43vy/zNS8E1ZlUt1uX
t04nx3jv7Z9y5+j/vOMAFgR2CLfF+QRAsSqrXAkf8vuKNK7JbP23rERTodckDYyv7L5Y8Bd4RdBd
ibZHDWzufZfIRRyYCyP0M6zBDo5lOGPJ2SY7WzPCOzR2rnJFBjKHICgP3GGMwfogNwA74E7V1UAk
O90qCBH43aNAtS6UvGgWhNjY9NmMKUfSj3VXSnDVQRhaGrcPB9K5dKvHsiHePFszuIoBP2OxV7c1
T2mMvFxHBN6Yj2mU6IR4vhWXDQ1uOsqAtkzx3TRudM+k1bayCX1p4sfqLypXYd9yrrkK5/LD+PZ3
h3ObgCmFcwzdPA9pKzmuR4WzIhVP2B+ivHN2x31DDGsnAsVJMkKYH2HbRhBHzX1J+yxNDeVzRAqD
UR6mzm5eTWvK6OvNh0zfoRdk6NI1esCtpqIZJDGcUHKN49Wm0Q6aSV5kmboj3B4vfT0Fjn7GMeJG
+6VMxrKFShpdKkb05+lRVq+QAyYS7n5Q9JfoRe5mmX5N2Ri2DKL+99Ay9yx1Yn3iUl+agYeg97Ne
9fw8sv9o+nQTp7XSaOh0nb92R849DYB7i2SdAgnloJf8Sn0SnrTPNg5xDcjo5iAS86KYb3t77Vpg
jQZXAbx4WIOrarmH7fw0eJCAbfaDaKeXF2qmA6ZStkgqxaNU4tMQwtG6/cxO6FJYSY2B8Wsv6t2T
iMz+GvTyqgS/hGCZ4nr7V4Z9t/9G1z4uWo83SmEe121VIHBU2qerVQ0lhr9pxoslrHfGJ0yo1Q0b
R+uIdMe7QYYB+sgHzmYWPH/QaMRFot4E3fZO4oyKPaptNQ7Y3CyeZaYzkO+o9zS5uiKcUedDfdO2
9/rP6t63Fn3a41Ijs2lMHB/lqjwHw6j3Kd9K6Ow92lyYutOHVH5uJHCYUz4yWI8J3YdpW+OcUnfD
zb1IPCiilps0Y7E3toIJvAziaY/eWWSbUoX/OSSbzN+hupSl+l/tXzbrG+xZHPz8tWO7/vsrxXLW
xREfCJ2PFUPE5ciaPkLnVj3Aay6HBM9J1vXww6IjvvhDky1ayCluvA+N+m1gyPo66P2oMuUB5q7F
gabPngNdzTWZVyAXkqR733egvF+qYCn19Q27OKuXowoxCeR+FaNDGohWVgawkVoDohU1JgZjOn0m
MZbGJy2fZFrofZifRvV5OAeIsZSWNPvVcdNAV3KJiJ22kqwsrzD61d1LvwSeQKhDjl2knmY8Qm7Y
Z04sgsuII1+wyX+0qMD9TgtCaONcy4ZXBN3/fxnA2MLTjNTttDmpYK/H3h7jBWnS15VpumwP/bXp
LED2ef7e7NQ/FicNTczWEZszlmexxH9+1c2ZEHnquk5lE94kpLyYG+D/TZ6oEgHAyGIBXItIVvPi
a0M3+dAtDGgeTQF6uFpBS3G5yY7AqOuKx1/tvNuxnvCYXNwjKuBSJJzNKHFP1yZJrU5YlY/SDWEb
YRHIcOaQnl84/YFoklpHmHjVukP4V0EFlP8SIzhMUCjeu8BAB90uwetxQgDCgr1jDR1pi3yxf9st
JpbSN0FRRrbNY1XgsYPN1cteskFzLIGFW3D9bPFpu/bq7F+XoMlftMAneKjQEqhtss47Wsui4dL0
OQX6GVwFGC08MqoTyjTF2KMTKn6JkYjCjhg0i08WnVHeELSAhYxd/ykKXdpBPQQQ4qeJ8CPc+RjI
vAF3XaWZ6BVV2RICjrHQ+Q+z0yMw1M4zdJZC/2k8tfkzI9n9n92gQNu/gOW3lWlGviq1LQiX9wiS
00dYXvqONWSBOhMwlG7WLjY9RduzRDiHFzSeNgeu4LN3JWPKc34hAO7IbcjewTRSoU74nGe8kOEo
1BzFblazIa7FgxZtfufAt21gOYh4KbBQmIrdRmAOIvLHNZZhzrsgNWTUKrRLcIJbYpJkadllpos2
0CO7/tJrJ1FuwTFkW5o0LzIzw7/mACFmBlRuCjWwE2wH9GiYtP096c49VhV+MAhKCbbaPYNzChRN
leB30MURLCOee/uSSe8/EKh591PLPQo64oEwNYdJ/ygiAYsHF0FQAgpnTRVhNI8DvGybHwOSGSeS
6dmm59XkGI8vcpXHT7HrhsYPg6IAPnXjf5+5juWEYpan47X6YZ6epr8GPOnKFq1b/QFz/nSCMvDV
RaXZHZ5nsr4lbjdp7SsBb91XYYF95In072jBWyFMmaZ1OZsYDm0rCHqUf5JrdE5tqGgfMgkCqQHX
opKT22+gh+Z5FL744vMJfFTFK5oRWa5SX74Azxc1rhQqFWzTQUjmXz5bL7T2a9Ft986hciTrfClm
GuMcyyySmYle7aeb0jdlEVUBL34woz/vgeWciF5n/mDFyk6i8vlNbLzF9Se5Nthf931Y9vkbKrYx
81qrycigM5jB5kiKjijrxt0enJaw6t3WtSg2e9BXBCPRdy07Pt9txgcTba06bVBrEQBY9yVlg51I
O56Ta1+E5picGnZrlCgPWtSErM9HTfHa2gZpMxh+D1z5/rvubFrcnoiVhQrBibmlRLuDXrooQV6N
92ckyQBqwhC5WGhkO5BguWTALmUYMjKpmlIg1D4JokfFTlom6difobBUp2yq2oyuUKVYea6OLQdc
MJTgEanfK5RYXstr4YzKiBwWsxsxOmuztuarUYvVm4Ir2/A2McIWgYC5fDjsbFOEBYZVV5L2p8ID
9f6Je0svA+2jg99Qw7gXKZX2XMChU1hef0/uxMcVtnhTuBnihg/oWcWoWlk6+AIS/rLFCQA9oUWM
pImpgwCgszt1iQJkfu0h+OAc5Zww1he7TSQ2n5s4RCRIXPzURaKlTtUqYWClqyG3YlR7zW9Ik2ZY
RPIbDAL8ZOijnezOy8yPk0nqOgCYg+Uq+w2bBEt6JqhpjigM911YKeLNOOV8LP4qs4IDxphPJ1tI
XZz2KVqtC0mGioyL1PIeC5XXjdWiRMuWLupjS5K3dFp+I3/Y0ujyhx9G5cLGFLQIFmJhzVe5Szkm
OPhyRPLjILjKwTClQ00p26CvjXqgYFuUy982JDBvbpsUyfqs5MawvxkQITeH8xaLQz9eRig3fC2y
vPRj3MYkIzuCwh6m13iyIPkfJE3ymwfXAGMB6YFURV6LKt92D8w4W74SoYMGUWANl9c5PAe1WmVV
KWYYJS8iPDTvLfYLseJ2CuDzbVSDCeO6DZz9uodZrKdaJ3ggi6EFDFnlC76sAg/2pWogwdQzufIL
FG3sz0+sU+CghaOYLdag1bYZBpZ5Io3sEoIFPkPf3dP3ml0Fp9Z8IjMn0fvnhP4eLK5cjWUuMd2Q
iPT07rAhK8iALjd80DlsWmUtA1C3YlJZDUgZyHDrPbDwhWxOOLBXR+9Rr89WRKjjZvXUzWCiaPRI
MENnjDjgIxhMHJNhCqF7dv+TPTYUJYTiCOo0hy7z5n9l1XgXDr7Ge454O8vzdzKeTWiZNW4TzBrt
eB+y0tSaMQ3NNHI8w80a6waqh/4gylkrLduVMAWdrP9NiEcTwsiJO6z6LHYmj+KRhll5t5bLTO1F
ze0B5mWVHJ6L7nDaYkBcyHs32J+LIVLimPaCxRTZPZufxYc9JNKG8Dys9D9cSYCYap5fGM9Hvgp8
t7hSsOP96F/0p9rISVmIJBcryQqVj/dYLNi9Svn2vPJD+r0vHZsSplIeJhK9eE8nfsqxbbYHsRz9
07n6V7LAwAIsOmenj9uCrf79wVNHKkpLXbDYbiE7HezsIUQIKazkrkMyWDwFONAyvIqRLL8hCNRA
anb0nGa4dNOIh5wy830PRNd46zs0p04A0Af7HHgYNxW17gfQ0vuu0ve+NiCKlI6CJVWS3qWVpPtf
7vgc//RkjJOOG37xJ0Qw+itVxcwXjYipXYfuzwOiQZWRhjVBOsdNawwFTt7A2DrZvTs1AeRd+x9W
84m2AnOaHTT7u1+fVw9lw/Guq/eXvjTtZ77WVqa+v1p9HAU85ySIQLPZr/a/ozka9i8N+GkcD2D+
m8+ecvHVw3g/wFfDSrymr1p5vJ7Yox4Id/gQGKELBkE+9yeCQcvMUv2siCbB8OAd4O6qgITq9Yd9
zFRDJs0gqgoA1+Zqky1p73LCQHvUyJu6hO9oYeMMk0DminMv/94OaV26P8nhjc5xY2echs6OMFM/
zS6WaFCKv1Dp58NiWF6M8GSmoCGrIYLg+CII9tkSo6rYQt7xXr3hPxg85E0melWowkj0jhcjxjg0
HxkKGkiAe5lTtbSaLRRcJaYg7M5msXD1XXP4Nv5GQhpKZy7oiesqB6CCyOEomwFxIwoNrNnwRNwD
VyV9prbZb+UQw+ptVJ9Pxa26I9ptIw43X0GF0uQ1aOlJbwMmjEfKyOBqmDdFS86VkwINJkKvk9n8
ORutxc7rujHkvwtQTPC2lKOptL2orky2pvZufWVTyjUbdfJJTfpOGrjUXc695ePGlDksSyrfURVT
glwPt5VGo5hmaUpkQpLQNQZ3xnfJBquYa+R97dhpV87wcCYszhYySRqBBqCjhoM9qQGYUhp5jNxa
/iJBqQA6V4lZYipG8ZzNWgqexwwV5EpgyoxPb9mAq8C3JTeaG6JsXyyagHPd1v97QT1DoVAKAR73
Ngn4BusHkyRJwfGDTroq5qJ/2RHNTIGER9QhJjOc6dcF4l60tlUOgwqz1s/dA9tcTDe2DUXn3yz6
NzYzjAZ7XSZvvZyHO8wuucvJedsOBF1/h9COm+9+GF8MN9OaHi+VuWOVTXXvEDMgwLv8reBXx8km
fet03kqb+A7n9+NwGXtAHJQB5aB7eeq5ZLIEjW6VXo+kLpv/lSlBghWC86lsxgZ+44dgRW+SJXej
kcS0e32TE1qda6jTGwCm2jYAjrv7N1oC25fqjngPrehSv3HBruCeEMxOjSgsBrHnF0OBs3JdvDx5
ZgrH9XLgJSa9gOuuB0TyZ21T+gP7DuOqKCKqmRSd20P7GdH9fjbHN1QxwQ3Szhl4Z5RrK2iCafoI
KMKzpAbHHxJcHtb+vbdsTQkkTs7iWQ4Vieum0IDIgkTptEIIuXnaxQvOn+NEx3FfUT74qWxFckf1
O3AMQdp2f9CDzo1cnaHszLmqmVzjTlTKj6GG4JhsjkM3cg/9E226R5BMIXUVMr2tltXv6IIS3i8B
hpAD0woQKXHwAgqQ31lKr96Xc+wXaX7amvNNR7LI+FCotcItdQuFhPMKKC1n0EjTVGf03Tkp8V/B
XBAaXY+cgPKDJHlvxP3dTOKzYULVoB1wb/eNxC3nN2jxhiCD+yB6AWVpPxBcoIzjo0qoyoA5qsy8
nc+aoJ4qn7zlF5y8yo3r5i+qzF/ASgMW8L0jjciXlLCsJyuUaDtoXtpnWQlJkNOLHgzwwqbma26J
XWWpaRJAKclUJYp+rrolbTv1oquY3joozY+hKafubYFPGnxkdm6QeBV+xkBBPBWzK5zqKxiRnSpp
dBdz1+JXnA1FyyoY5pIs5D4rdEPcE4neSNVo2dUUX7Nu9ZDSOtxZ7PDbupFY5JWucky42SngiUJ9
9E34cLWCiza9pel3MD0MWoDL3t1YUu0VPZhz4TSwlAVghUAfHMfn+hAy81xdhXNnGRfwTz0x7+fv
sC4WcqUZX41k/2DNcxyQqJcWEEvBNTuvM6WcF9cPt4A5dUQ5HeqvKg8Z8aG0DDtH4ZNlxNKf6Eze
uLRE4iKY1R/b3MPXOXRHpBuMW/ugHyM31NMWQm/Kh2NhlnTCjZ27iZpavXUe/Os7yuSMLM4LoHU7
CopaAo1uCYnehpSaItPldazcSSlfrTHc1lC8nn3+voEpBvAe6/LDn+Mf4yjMlsSaMIeNzJDotuwh
Umc/VRl7bLZJwWqGNUWrcMTdVYuNKyt2XpSesNR9LmEQ70JRWyUFWJIHY9WxkcwF2GPr+jb1XQ+q
3dJplkVXPbpnrMJopNTKz3N7fsrr6hV7QdXknt+tur/Iybt5djQN9zKjDb74KXeiLV7yn+UEXMMW
meb1wK+jiAM65KxBVoBSGI8p9Xdr5NLDuBTJrAHDYo9JSiElgaoYqChrXnvQ6wzKKfTyPn5Hct0j
+ocdo6Cgi27Uxj7yeG3O68YibIk8PHauuiDzigGaVDIp8i1whQZ/3iU4rVPPo5RS8t9hUS8xJvJ9
TzbCFjBfFZpdU3D1sDf38XIlVuRSkJVZuUp8wCKGrtAvIiU2FGKWb8A7PUFW6Em44TC8Z4lFuD6B
vmjhs4dETmb58FWi6vLYxgp46QPelG5wEEHH8076/w07XpO4MGrZera3ecL9JpHVxvuFH5Hdes5m
GaS1gP8M/it4t0sTz/832VYX9++C41VdHzKRZC419UB2+LRqGzpr8MuQGjahw01h8w/KavRJHpx8
Bn2Pu6Dft2phxZfWkzLiiDVkWUZvM7dzj+26/FCBzzjNunsKXLymsta0CQMXWaP455ZW5TtQxi7h
pg2rk94nb5ZMur5S8YSyx7gDc/sEb4N/4ltrNNkX1oGU0s3vHa7+J3Qc4ht+V+IAxuI0hlmRgfog
TvhmcyXKhxmTE3Xts75eGlWW0USG09MXN5uOQ0ycg6NoA/gewahNlL+bcJgG7SGUPgz1Wrc4zma+
+v7HcYt8Iau44GxwxnQbIgEsGXefpyl3m35iUUJz8O8dnUBZ8YS3KFyfjpl2eVtZPItvZAJZcv8g
vuis5sEIMpmEbqdycMjALAMo/dnx2JY3Ygr876w0OsWqnBCETAA/jr1KCi6vhGK+XtelJfcMvzEM
BUlEV8/jiWONRx3u5CuX0owJlGkRc1BJn9GOggUx7vFvRNab7sfsIHfwzlAR0HrP3WiGmNoef9Lc
NEG/C4PNuyjhLdwPPdea+DOWYUCoZ3rlP7ekhMFGm8q/pbFwx+vFgTeBA/hzF15uTZSOFylANrzo
CWVOAKZCcYWLQmx63Rwqqn2VnLQRDhyvBKssYY0h7ETnU9HAyNGk+5fD71WWbM+23lZTWGmYC9DU
ZZe4Sl8wWagYOyqLvvhYN2hmvt/N2U20bWFi4vUH3wl9nOIyvt2rSQB69sUOehmeIrRCGSvT8dem
y197vNJmaroe08ksJo2Ekd58QOEGje4faY56YiM0LZ+ZiNpdi/9cGmb6cSNDZdmrImv/0IaJFavT
ZxnE9cBk+MJKD7mWiImGUB5KKPhlspWhsQrVakS6Wp+j+nb3ktv9ddqHADMNTzd03SSOF7L6eGDe
LhGNZyOYNoBENVxd+NZQkWCX0ONZMAjWtjqaGQSHpFuY3FYT4uEvlt7qF5UU8+YmsKv2gBA4XKU4
lXHp4SuGEWH5IzH1qISxlIljJqz4QHIGilFM60ONBPnvAksy/fvOBKGPbAvmtX5VGhAS4lqAS6Jw
XK3ncE7cNTI4qAcr/qJiD/EIDj/NNHpzngV7YOpFR/jgVRouOyGYuW4sOP1l3OpUk5reOroNExHz
KD9draUg37btYxXVZmoyMbNIqkUL4G4UIkQSNpAac1btxUe1k4qM4c7DH26yWCGEfsC+5E5n/tnR
eL+bOEDdj4qIXGWcWHY3Bc7BWCgqD1tW6MowitWcNN5p7j6gILeATNx1+LxkqbKOeMIzWku00koh
ypKdImH6qraANvBVfpwvlyBXBEk94yPsZTjzb6z7Ad4jCVzieAp6szvy5cMYNHPvcyjVZoJF8AfP
+4R9pj3qrWTWh52q86V/STK4FrfKtqSd3mogBYqxQ/dUgI9JxvVMhtqNZQER9owyLEdQxIjL6rgl
KKHVQEDTltKi90QWdAXkOFdPA/N2ERbGTltkqH68wxNLNGZhf3j/NOHtz0R2EEofLmFUDmMcp/Ax
xOYP77Z8/8xnzMm17ruD43GQxA4CppKT90of5liWOZplTqlVX6I8pBnYscto134gytf1VOVj15xO
4PhMva7OkZh584eBW0ayiN3gG4r8rOp8jO8wNLP6B+/7fpYLL/h9yOF4KR2Jqwl8Fi0QsQIChhdS
2V6PS34lw7PApm5GihSv3Wa+B/QJvG1ZjCDpN68tOivWP4itxvzUgKCGA9X0mi2h+8AK8Gefi39g
w7pkqvkfLEo+TrbZIQMoo931XcVfMXDXg6pooUwunVd8SeB+fvxv6AS+dP08118ce4/lMJ8j1vOX
CxHmaD9U2QR8Gjw35ORduLuwsMgIDLKzIausnaujIN9GxQCFlG36UNxqC6lFSpbamM4rb9JL0psn
powtDZrE7qXEWpTTFKJaN/RJE3ILaP2RutsuCvrdf+Z2NFK47Do3nc2exOCvtVn5mKAYRseuywZR
3JRzI9zXciT6byyLffzFDIrn1klwx6Z43gGvZvEn/GnO3yNaFv5XAywVWFG6M4CiAj3Ss3jYWKS4
KWUXhVfXtedVAwJ+yGX0fqNIBIob7ztCWGX1xyZ8rf6micb4pAM2xXHKJv0owRQ9+a6D2yJe64qS
B+s3rx+hDtXCXgGayxc58X+TJDOo58rpXajSc207Smds0/o0miN4mwszyO5hY63/2m1dYxk3dTM0
mKEiX5DyRMLxcpYhGaV3J4/Fs4QE6VLLL8AaFU9TziM/I0EfDD9G2OGQp/5jhfwd7pNjM+XTCap6
fYLrYrmtVpCaXjzQVvt3eovEH/S3ED8JkbT+jq7leG08LDJnw4KH4dqVBkHE3L1QOxDsFXe3TPBJ
TekA5Mp81n7KzPXGGqpGqzcI+GjnnOHDzG6BuufnlAc18CSUzTXhfE7b9EfFx5PGz3axelgPTV8B
CyoT+YL8KMjFC5EFIL0GvYrH/Rskn36Wmx5LClAhDA/PXi3cWnhF8sfeFlVj63Go2+IavpuWY9WH
1okrTjwlN3h0v+OHxupIiHvGNLYUi4otg46Tf/fF/sVghegLGd5kJzwr4WJ59YY2JqZmUs19cO0s
sQmD4kjRSO0xxWkDL7SdG/yv6+4ltZANAYuNMZTZlXl0eM9gMv6AY/zbD3OJtfDh3ef2OMLxUGKJ
jD9gZChWFzX7h58IZZqIADb2qPJ/7TOVpLJ62NkgbHite269Z/3Hj034qfaqvOiPcAKDQE7Mfan9
PEtLeXv2Z/rnOWBV/SUle1ZmhvC3n79cSPirkx0QnAU3JsfLOfbqu+BKS9M1ZtCkbgm1HsFRjW3E
LAIt8FdLDn9/BxnA8o2wqqj4p/2YcbVvmlH1e9wFMNvDb6GCvV4d8y3WhWDfNebBfx42lg2LvXL0
bkW2ZuLE0SVMrnukVsRnwcNpwt07UZEBsTL7ZcL+wENHqdVHWd34BIJTa2dZruNjK8HXHrYyONLW
KwyqiZ0ymMlv6/PqkohY/y/Iy8LptY12P2cWqfkufSoVXbVa1N/dp4euI3BD4UW5HuVJJ2hTHWEf
lsu7ky5HQtBR2y23f3b4DO9pJiiN1wdfmDoTxENPdaBUydJH2Gi+gPYpFYPnhroHf9oY3GtxZUKb
/gI7/xU6ckrCMJF5Q8qHVT6q595M5pLLlTmvAiJAMlCIo8a5az1fEzklq9M6UJ6SPWgfK9DAPTOj
RtF5H/HV0JSZYFz+X6UHr5EVj0aHgRibIAWIfqls6CpQ7UkLGWj7ShAdP23DeKDBZ0hwkqws6IRx
zA+Up31Z3MBJNU4dC65gai5DGGntxMyz+O8YLpoPx7yfn5kh5HrREAFm3oJXjHs92qmwwOPDaC79
TwY6v3RzBXULX3by06yV7mu2N7zPS0bg20ziqHNzL8rpKXLOM3ksGLUPfByD9lltsIo0Xa/QJ4lw
sv0TwRYD5eiRgI4ejYVBge0lZN52wCuceudwQHaS8pb+hfGk6IGZgq8JbBp9omkAvtgG6M64vRC+
xF5POEjjqVRbfUwOZ4omaceM3VGgFiJIFqsb4dUxzLZ9f2F5BOhYRqe+2XIXgccsYg6g0A9s7VRH
OSYviru59fE5uTDGCJP3mIb/VuZVb1M2uX5QgiBYoUearFeDN0H9IshjEM7NKS/vBFNCL2M2WbqC
qdr4d8kfdmrtY63xW58OsAK/LhiOu/j+NvNVSDsDMPYhJUZIAWEr5JCgAEI8sww2dNLJCoVmeF0F
8h6fo8EApGjCkI9GGkv+SzkCRlz2xyxqmhXi7HpmwM6Ka6ovBbM/z2ilxPvTpom2+4sL/pmhKFL2
SaeO/4A7VGRmBCA3X4AoQK3K1Y6VDY/ZBYz8SXVhiiYzml4C+ySDBGi8qrM7yCV19FpiTp6OceBI
obsr2NS/q4cQtb0xd7aqrlASkXNA63hrpY21BMuDiMieIBpH1IhurNALEDkNGoy6VBYnRPJ53ent
jeffB13+s2purR4E0WR6yC5sJQBm4kecaTzdpTSAtHYpK3R08UOMPoiwmRyjLBBkro1tlN8aMtPb
5EZ3MHG2e2pZ3fm17UI9JsbSV2XShTGkO6I9xot4SmbTG/BdCYBeIOXMtXKivZDECs3NhglwR7F4
Vudxq/5nwKztm/hb0sjd4+qZNucxYQ9Zt6fWR2CgC3/qdFPAU9gNT6iGvz4KWBAgO+lNWzb425/6
QRz+vUb7EKOb/tO25bN+EoGy7V+Z5C/2MZE3ek6Dj6locny2EkJyXLyiSpZzvYHFHqdfyN2yOKPK
Tdq7eHLGBYXWGhaoem1oxvD8W1VoLt+q/oqyicHSLZL4B0ZTm5EdQSlEqaoVWjUDB3s68oXzRunL
hHiW4ch7xYm4CeU85ks2ojGznGYUP8NaUAZJU0laA+wvYUhMhV5BbxEbCuPUKwOyqpLWPbTluWBQ
xgvI66XeC/3kGYa2uuRgEp3moMbncqEJbDgEoh2ITPE6sq/vq/9YFD9l5sZXKWW8AtPn4HgjkD49
z3JdtGx1ie/JVaDyyGSmtnPsPUfOnXWJ7rtsQxmcAVj4frA9LiB8ED6B3Bunf9Qa9ev105VJ8NG3
z0BHaTo1iiWywJk9anR20gvP5ws4uX1mgOiOUjz5/Um5wpxqqfw/kzB7qObrw17pkROJHhCWMaZl
XTimY87rVVypuXBSx2Ut+JFKyLE4NvMCvgyNLm2eJvq2UI2mc7QIMCYj/mA15Dw3yOfPFq0ZQKQ4
99PoslQDweJvQMA7e0bwXvmuVl32RWV0+3k4bd6PtzOLZ429kPZuuvzOH1SKf/2sVlEy7nS9b/ay
msO0RIdXpv7o0QQk6ulJKMtvge8XyJNkWN3P2xA4u8K/a8Pk413Q7vWBI07j1gtNUXyGKNa3sEvz
xKgzgULXcJcZUlKU63/+me3dc/APAhyg9lX219Z2eDAq7Ltx7qNsUwSLgb6cj2vWcoX6u/nEvrZF
3jGXPXc6zsOAAcIk0hHzZ4EeSkF6R6kAkVwu+hb8ShFcpSR8/uI8Bwylmod+ImHi1k0jUAwCeVmi
WBZosSj52Cg5B4AjS8h0DJeUPvS9PMLm4W+86xLzQU6yAA0zIzZQIvdhflOy6c0jWiYsq83WPgrj
i4yJVJmo98TdBMEVGEVjGp9QC6YTCqFOBolS+Ps1XWFQW5g9jY49EXyPH5xgfOxnEm6a7+dFbIdC
io7EFzdTWFV5e6qXmqh6hbapNwpShhSeWwCVvmdsusGZS/to/eNtnrq2NB2WiuB5P3uFAGmuBR6p
dOKO3wCaeoQkA6M1JgxuHKqh0OlKi4a2ed+TOjiLM3+au5O5LiuSnDQYBU1RxwPwxVwkxZaa58rv
F8FbSMCHajHKDzKlDxJiavmWDL75PdgtDWa2LN/T5MJFW6G6qirfTZK5ON55za1GchRDj9ScYQ7f
eTMONGdCPdEgKKuo8sLYsLcLTAVsHXiUt3/5+YH96MXJVMRJMIyfHVNxoBYRXPr0aS2OMPFF8gJV
kZPZIu+tqdQEBOPVXnBXFKMydvp7cUIBqhFNgrf7yk5a6FyXQRntfYLAJKgXSqM/UhpmvweM9BmU
BQX87Sq5nYZ4LlQvK0usoRGclfHiUmdwHX4P2XUsp2KoyxuVFCu/Crvsb5OnlaQPIJJDrTBsAKx+
JcjUDYmESw8MnV4kXauEh1R3yZnRfDkEwqTG0BhZ3v9d0YJHAQl9Ax+F3/0PBcmHE4ZgJq3YJJRa
NIID3xFDqT7MQmvTQxjFD5vnIzSKxGAdfaWulUpmO3xoA4I/Zr8g8POFQfGw0+i59GnKw4ICSk9K
+IJly57pMKBy+vI/fhHMc+e6MOqv47Ufwu26Jxx8ZQGJwde25PgF7qeLcgT4NIRTQiIzi9bUNTgL
5bSiVG8HV51iShZhmmc1Gzjhh73sQ7B1rFFtYSZEiqjU3cqB23SIhLpNlq2y1Ewvis5s5rHj/vKW
OI8/hSl9sAV59sr14l9oeErFLBIBlseUFZhYG3n76ZmGp757YFJRzlwGu3iTURxY7M3c/vFAyDVV
mofU36HuulHaz8YOaKWDGx7fC7KDRWLoX9qzngOQHaPlz96DG3T8iL24+/0RhqN9T0wGztVF9aTI
VUs8PMUqD47g097eJpoDQppS3sGoea/DwGsWyDDXcwx/N+OCdWj5wf6IDoaLTQSTvoHp0Z2MbPPV
jxillUOQwOrNZjkW5ocxdRySR4w9tDHTboDLRHWOFHZYpHxBztz0U5Vw/dPZsJvpK0Str3jsJKNt
13kVpOUEplk4jlHM3GWcOGcY7KU9lqvKgSlEtK/ZyKX1iuziVuh7IpUr2ZxOfXDWw/2ANt5jseUz
bn7WsG7iait2MjNx9Hc0vPCdfad6iqPSFMUncJ3siplq8s/3jB5qgXCURb7ANuWBwsoe5mCCPm/Z
nSbDm30a/MY327mujRdWZF4huRhvA6r0u5Ospv18KQ2HAbOB82ODbJ/d3TMFO7sdES1a9HhOlsf+
SKcsf4pxiA8FB702tDuDb//j/oWEi9vIz7sQjbX1lpOyysPB5X5qRYqu7vwgx4Yrq4FkhvE0IIsK
5BmCk1CpATrI0W1iYs5tJtozJP0hroOuOSQggJgiVPzQEdc7OKFxz2/XQ3YEhaY1mv9emMRlPnJ2
fp+FliJh5Y7szLes9YbdWy87yzlzrcSAry644FRQySTtI6l1w28HeCS9nWSWeF0g5mZ28S3+wAp5
rphn10cIQDV7QqVka3959XWQjG4rhcD5HmvQLh0fIQeoDaqglnfsp6UUmQwz4rctkz2bnx7WkoCj
Dqw4ghWzigwHiOp/TK4qGJ78dUtACzhg3zul3jFLPnZTWDMpzfzhs5OuNGSgHYADdjV4g8QqkcQW
Lo4C2G3I8CohxbGDgcOJ0Uahghcksf2e1t0Aq9UZ/KgQto53b2cgyHjsBExqbeQTaq4uhdYbpQxo
Bp8su4MpUQoHoilEHb0tSwW9eq4eObNj8LeobL7IK27P00Hj9M/agOe+VtwpqqYXidHFKYrhqA3+
dxDp+apd9H87bedaj8nuojDS4IdcPRuBWeQGik6Tk3+CjwXzxs3+yN5C6JHXO44aEQuFFCFWqWJu
0l5Xb3nX77LnLAKf81UIwCbmJ6CvuWp4kyff3VEaFcdG+uMRNL7wqH5L/8wAGPRk5LRtSd6SAx5I
SP9QoHqMCTt3S9zbRDSC5/Fawe2d90sHUmK3ufdYWGY33u9f1PigRn4Zy1JPiCIHUFi8g0ZEmaWm
vvGDqXB2fI4hNWi2hL5mkts/HCpNn/Jk81osq6Jgp/+IdnP41z+HUll3BgjP6HHz/YCcO1QJHTZE
puqp845EclMRnqqO0ZXK65ypqS1oBrbFYZYWDwZfWxN6GmjJN19ybBNWQ2QEk2Ry083PAihynF4R
EnG0uN5ka05vd+HGTvXRdQHAPIMEH2EDMaWL9zZXY/fGylfKBrSLn8Vug3w0Pwblx+TxnSrH+vN5
HunMVfwCeWGoyRAQv6sN2M6CJJYj/b93prUao3VIiJKbPlI7uaUBpj/jmS2EmXDsY+T2keL/u4jM
zji768e6X4lUFlkB5GwwoZ3OImAJEC1rWeZjHAkQXbBR1mkDum6YWPnMpj7QYIY0YPXruyv4WMrh
/iq0EIGHmwuYOmhPDHW+6xVnUOz/re86/Z7kw6tC6ABApI/jTTEjNVZLGv4wGKpQLeSJjexl+CY3
n0cM6E5oDDlO71yAXmdkCxiR0X54r6vUsNP1pgZjqFD6W8wCEvfUtGZzxWnMXV3KGKyhStZoa5Np
2zd9qGPqVl8xnQEW87KrYGJ+0NxgPgbJW0XTXqunFPXyu616iNuCPg4TI0T3daZfawrtwz+rQ53N
ye066DzoBPfIW4AA2/zj7YIWCB+f942XEBaSqjXbtynP0p/MFiPkkE1mYa8UOm1rbBxD8LMsA/T1
eHKyk5LWT4JTfIGYXgWh4tGbW7wAi9RYaXBcJTBeP/js1XkeePWQ640zwGHZlpC9jRq3JMrmggQ4
9kRjQMmzH8QI04c2KahTBm0Qbvu0OGrL8aRNCZUQmVj+o/Ttkxi6mx+5P9EKWDO6XR4obkmr0TAe
nAKR+y1BFpaG2D8GorNWHokfMDymAo2uPd+NOIDyKz5pFg7NtYwziSBYliz7sHxr41SLXN9eylEY
fYVaymrCd2fKG/C/2rr/SEeyzjHeh7oxPbciZbkV1a6LNHTNO+usx2qKfL24le2TDbL7bWqrJrpI
/FNZnAQLUYn/kRD+NyZj9MNIhn76l4FI3oqEHfm9z92ik4cNm1RTMVEkL+wuK4K7rkWz6a05Ojjt
jy09PW7dJHYgsUuBnbbRFelYUNdOSTLzaQN3s58rFqdbS0VW7wTzSdeXfvcIBMsHe2fYNFBYOewj
PFZliSIkKivqNbKK3VUg4kgCQHhPMMz9fb6uygCsecIPIOzyFXHe5GpRnpREjTgrPPR3lIzfmP3N
4vZnfqq/8qZtsKPX2lRlCios5UZwIVvkDnGRRqcGkHvEkP8/u5hFT16f+8ylBARoanxEgntuxVMp
UbDSR8kIQVzyyME0MJBWVBx3jnq/ZCe1FtKGPAwLlmw86FDqx2kubiekyZLUwJ4T17k1+RD8uOL8
6wi/sogfY1+TsBeie3J8xMP4dBCdy/5udsz+8OOsrfdDFC+P0s4jiCxnFbJJmR2QSI4TcD01AP6m
dzM7YnlvSeoCkD6ZYjrK9UoFojJT4isJe6OQi5wPLsdMoCeieZRlEXG0EdH4f+W5tx0A0i2POhXx
6+z+A2gqg2LyJjgks7N+itea8l99+kdsTPSL7kGqVFMR5bMOFR77wrJDComicndrNFSDWUIlsmT3
qAAVtrEMc2lbHMSV+6iDxVTy8U8zji2fwlpH2Fh+PkAwTuwzNfGtKuaI318xcDwcvlLx3DQhQ2OC
Uba5U5xUJy0Fgx2Vye5R/otBZyOVMRrkaYLMhe/6ZQFWClsWXLsmd6q9qxEq3hhnOZsgQIWgFyXD
gWUH2KbVM8w64sjjXuxhl1PhwXFWrbCh4q6KDudYzLdyx4B5s+mKvk9Z0W9Jpaf7MH9iPTDQCcTZ
/xA0K3uByLDXRwtwxISW3lQ6A/4oL7KeQX0cnKTjedJh1qY8FmVaoI0VSt5bNLRs8gVhlacUoOwu
IjCIUA3Ebw7Cr1LHWksNtdtQMEatxabqspu2/sIfdBvXg9R9XSubpVT1a7f8UcJFdP4XPkWxH1N3
RTb/mQ/1pON6OIy4w24Fx33O6lkf8nsKqWhye7Hs3Px3v74kZMWptBp17hJGwTlGNudR466jA8Li
TK9l6ih6lXPT0RY413KHeJGIo6q+7/4iyhZoDEH2u3lSDuzS5UXa4tML8mM15UHgFluakfkMY6qV
vAWq0+HCq64dvVYY/z1S02X9TOB5zld0hsjO+awI4YNhL9aigEm/8wot58tv7ooTivJj69c03m0/
bolNlYEJBEg06ZM6Js24UdGL1AAp5hjJpyd6Hvh/2ElMCyjeMvD40+5HmCmuVjL7JhLYec4OpHUy
6YDEWqtTST139IO94AB+xVnyVtaPrb25uxA/hi/MSdvANBw43zerJx5x0QCeR1CcBu08Pr1jRkfs
YloIDUkmbELcvNnuVMCeYRjv63bTJ2K5jswQw4NaeZIdC2DD2OZ8dROBIIoqTgjt7p0v4o8S1+IH
ibj+ZW1AJ2E7RrTybKkWwVHDLyXsxdYgMv3ReJ4u3YSjPBxZwF/CqDZOW8Q8AWqveiEdYJJA4DJ1
Pr6p/W1w8ZfhEaKtGNqjhCpy260GKLJID4qF/qff90DtbnIJmaQGvaLzpOiCuKkP830ysv/j25Fa
+q7+mhJhjpHcD+LTfjAmJ2eAbTJtUx3Y59oXrBT6540O7rmnsJ3/7tIn38TGTneUD4TF3yZE3fYS
C0ei2KTHWjauLmrSeqk4Zp6nn8R6Ummh2cbmwrz+lab/4rX8u4sm0uj0WV8/+Sv78OVVXSSUCbat
J+C0xV4Iioq9ofC7D68tBKlKjhmvqAJ/A2ESCDjmw7ePUl0WsRKR2w7HEwuE++qAN7B1B67YfF/T
AYzdu09WfUCLE8FeE3VLD0HqlGuW+E3T6p3YqSPiGLdQ5Otn8dVvVm7oga5hiu1qxu2ocUVGbuKp
69K5p0oxfB1AS3oGRsjoDXDpjFmopP7FylfobFT5ukUQ3s947RNO3ns1c9J1Rh2L8+WRWprD7r/U
o1bgrEHReXAHDUrWKEESRoflIly2/poO/ULeTLZZFLXRNywaM0jb/aY9PoA8XNQYncfBkS62uYcx
55VJR0KUoYYz19lrPKgoermpssXgJt7YQ+G6k/j9Tw7iDc6DiUlPktJobKX3iGTkVN2ce8hEerdV
IWrG1jwj7T1udLs4QpOpV8mN6/UFt5GdfghsEQGRnxYVPWSOLaPSkhWKY79xJsljyzA+Tb9w4IfJ
EoN4pyoMLvZh5C1a8mgr1p/aJF0KMJv5Ae+/Bchnl65Z0/K/ve4l/W9bjvRNlf97LyHdveq1L70K
7011Xyls/pexfDgCuUDRF8887ULuQ1YwpuE6DUHDCOXJTt7u2SGB6wJEP8rton5WlJnhy8cp6bhF
cd+EuUgL44iW1UEXdECDRV3HU3BDxt5wqRZPic67LyjAxGUVEWjlq8D8AZRgdFUzH/cJhcx+qMPS
yEwUEERGoWJG+U9BkJEhv+BW86jztYKpyYVQYPQdZxD/MvcamZcyaY/oYvAC1PKFnnDxIbhE0nmk
1wGPjmR+JZRSglgM0kHeA91HERqldvrPm2ZzPJst1F6WIxRZCwlg+uRG87fcTf3/puOTGTl4KS2V
zRoJwKpE6kl8s5elWnZM2PAtxvgEY5lEI7+QoySLPUfnI2vh1N6NcAGX9H/oNB1x/RnBfxMOzLTf
iEPdUC6X4PSOUgXk93w3jNKa6e9pVFzi8s72R2L0uZcKaIPEe8ehN8OAcT9TD5u5+nioEE/kr6O2
o7nTIlPI8Tfo3Z3ZcKFiGhmYPwbXRLqGT+8i4YbgJTUJ9ok+ZnHBtowaiZ37KzHGlSJokfsfCNgG
LMoDvu3HuEnq2f+VkEtBcm2ik7y/Ea78XXbEj4EtKxMWBmq+OFPFspHepW6evNQ/A3pJeH8MarI2
lxy6xrUh1YnnJ9zODIC9QhTb3f5vXhCsntQPQ118YawbsVkmwubDZF6QlLPv3KD7ke4y6Q0HC5dg
LvAvzjGO2/sWbDwq5UCUWMsU/ddP/OPkOWg/wABqyuza+9gifoiwTvU8nv5JKxQ2u69rcK36EPZg
l2erAGHXzgFWMuyawy91VF76kgH34kz24u0229nfk7GDgXna3jd6HRHdPD2LqyOl7nclChFZF00j
eJbvxOZ04x5uWU4b5VEK+D3Cc21/pRDkfPduzAvKGW+Z+JNdOEu6GjpopWLpZbVryVdoKV9UDxb7
vvK0PGZv1z5GC9zypnh7yrdTVOfG3s7JZX6UnSBm11dhPSJLMq5XxP4wfB5y/yeXxcQgumNhV2Ak
gr10XLnfV91zmZ7UrOkn+B4BwjVtcVxCnwJsB2sVFxDSKCb2s7ewRYANuyzEyktE1x5uPHJW1g2Q
frljUT1ZIYgrEf/IfS3uu3AOg0JZhfHFlI7U+J9B8q6Xxn4qiUNWyt6d15zJtSK2zIwvdVSo88Jq
KQZMAdmyDpEkwS0Fj/R/MG5y+33EKH0j93rxtzHtEkf8RNptRHC0rWXhwNOCuTxT1W9Cl6q7pLWe
/tMboTHWeht9Ty01Ag/d5oZTKjVmdQRMeB1I5V06kSdMNayhPTZp/aQp6SemG8Mtncsss3vH6suP
Dyd8R167Rs0wp+utFN621b3IuirDfuCfTO9jZQqM4ZjWuYzzx3pnD37eHZe0IGnS6PqsF+8YIzth
PqZAVyioFEWu4xNfeVYtwDkNTRe9obWU36xjegcfI7kOHCeSj1M70z8Y4SJhemt8IwB5To8aoNWr
G/h5P5WIRrGFFlmEn8suLSZm8fzExHiOu3iDCKT12wPg5MJrOpgeRas2TfBm49pjxbqarb/qCBR0
hNAhK4lO1+yIOhbmw37msSXZz666uPrT5q+61C4TbdUzXNFqXQyg2dM0oqmM+eFrswL+pF+rwDL8
eHQahM1fZgnK/Ta5ZNFjdY8LXX6Mi9A7nuu1qBiM9srSDe0Iy2BA16lKLOwokAXsayPbVyPAMxj6
24SkTHJdrU/s6yvhT2QHpBUvXvGV3BtQQ1MbJzzNuwvnFXec2REMYe6/YPwWIixzAHvxPC54hu0x
w4zIarcbFB/Q+VIVfRKZzfwTwmpHtDJSEiQaWwKEMd2k3hYD1PKqafVo2B7whENac80Hq6r0mWYK
SD+tNguRQcNrJwHgq++rKorj1ovjU4w7T3x32VXz32WhdxF6IcNfQSqRxwBHY9mQmoU+6nK+czur
ZzDm0MreoXg7jsy/iEAkLL4LFO4VNJ5nCdH2JcdFokgaiGERjh59KGeIDz3030P/d8QVr12Lv6JX
19oJEc4mVGnNq2a9rHUeACkYxm+V1WAUCLvpXFpoVpks/wTlzp4uqemCxsdjZIhkVaFL4faQo6cI
MkHBxLiVgp0PTV/GEYj5fkv4A1VorWSlb53KirIRhYOKmt9BY5DQiGQh2hP/1fF/n4txbEUvi53/
kFRytK5jVnS2upKNd+ahPYVzNeeblyDUoHrmWkHKrqCznZTinIGB9Ng+LgA8ED3BxPAuqKn8PlDR
xhp1SlW5oiXREBoYYxd1EDFz/HU++2oi5lEqbsVItYiHRJptzNhoQkHCSNfpASiev8KAPJS57uer
pucCnVM6xPp1UvjHgLehAuT4O6NKjE7+NCmhjRsnYkCp3IZ3Pg2b1IzrZ0xU+lpE+6NoPH72z0Ym
ZPwPAtXy/Ny8sKG0vM0tNgGrPt9Zpudy27Q+DgBxkzhb8Gm6vbv/2Qimwjwqb4cKZVHfoFqMndfE
CHRtMUTom3skVhFw+Hw97wXELM73MAGeRNgqM8Ri/op39Zd4k13wJy+KHA4hHPReqeSeRuWmx2aX
yIOa9uhvDSeJVY28iR62+Dlk3OmpyxUcDGZtTuG9NKainMneYUni0+DlbBz7P43gJQwxRHca4ELG
VNjwsMKfqV2QT3fECVOc0rifx3Y/myceyQeQ79X5F9MGlVhHuZw8yc3328E2oqasRvOqfRc/nJPg
+jUFWQ5F/rZqAfutY3L6g1jvd3sSaBcKL+rxkv6yLGnqsJbO8CnJ6px+CHq68g18aGZgb5ghKDW+
UATolj+z2si9EO38fcW7rjk0pJLx+hXim6k9Zobxvj8n2sOKWpOfLbBaNCPgqQewEUtuVx4a3YyZ
OAWcQ+NDTDVR7iSB5txAlfJN9dqlP1Ufg+0TKuqwBkevVP19wW8DU/t3k2+2yBvzTeZAkjC49mS0
tzOIPbI/fyN/auBu6ZIRnbNKp5hoy0B0C0SCsb0/f1+WGAAZRbML9m4OS77TychJzYxnTw9Nfd2T
VNjtQQDN9toxWlxdTB9gQf3JWDIWy3kqTwHpDrHjns3TrCy+K+56tYHvIt0vt/frCW5kKtk6QFLW
OPZJdmWbCjoc0SwJmePVNazh8IwNxKt7SSe460HDOg3eXiJjo+Oa2Wltd64kTYG7+MhyINO7AmlI
6NCsmL/+2MDGV3IfkyLHnKtKiq5TybWjniV8eO7KG9ROJP0VCum66R21GzsqoL8p5pHJ4uVz0Ut4
AGoL4YRmvluweF8NEUj/iJH6HVlKFn5DHIO2OHXIRdyyUxGqXGP459/CaZlfUhbuM8jsqN+7Gki5
drBfqvoiQ/LTh/ZACpv2Q/m8QAs3Dlx/FlE5UCtnMthAPTWldRGZ5ttLXwUIQTzloO/sscN+XK3A
IstQgdj7czyp8mMXPyzTEKRFGgqC31WFmgyZ8hekQPaJjAr6CYbOe1Tn+8f4F9nu7Z0ALWFmDbq9
aId31Akfs20yC+eaM5esOz2D19c9IPCjE3pGtN+G/oiVOegg83M4qxMEnwUoITXMJxtDKxUpCjZD
eBYsZ2D6q7rS/IS2fKIxO79FlHJyQgQdfKGg9YJL1qrydIn/+FZN63yom8PQ79KYi0ljYBUIlkjJ
xvKUAvn5LkmF3a/ngb8tviJ87LOxADsLY8ljqfI2jvrxhew/X7AOxPc111em5i4Nrcjrna0YLsx2
2ib5yLKyV5uVLrJ6IjNJuAdivcgWHd3c3t4Qnv8oWiX6ZI9U30cvQ+CIyCrTXeofb103g2Le16KU
eV0x7xszI8W2iFLS7dM8h8y/i2s+v1OxDcp4+B5lv6Uv6keeLo091rYkPwGcDfsSxctwYoY6IO+O
tJVi1XE7Gu7gvBVqGW8n/Z71niqOD0qyXkI1WxXS+VPI8+/10ORAiHFhlgwlMx8FDR5VrttwfK8d
Y6A/yYKjaYDa7n2m5ub4NI7iL3om/kSDfVETSKVwmufVey/dC1ngM2tqjkylkFWvuC4Yt3wCy6u5
38ZUcWjPo5tZhR7UNLuho4OhdnutojHXbOnnBZOLHpRgW6ojjZazUGmQ8j72oTXKKJty5raMpRXU
L3SnIOxbQOHInkQA7rC4diCpEujS/JCJBCvi78VzYB4gR6+E6IaGSTrTsBbLHrAcwKn29PkgwN6k
uztTO7ISIVjQiAPjS0sxI7EFnfDuyx2aelp0jD/oMt903VrCHjgT5TBZ3MNw7AyXp3xKbBwJ2IBr
cB0n5mdJQODRBsfOGqs+YldRTNddQGtMVj6UEOgbLMO7+W322sLainr2vnxornrgHXKKENS6ca5F
9hoxYriGNCMTZFljUaS5NoafB5/SV4h4gngNvCnIDUAoTQHh6RqXcVxoSqsq/l+vvT6udjtNM1EX
M7NqDNRcs7PrES8iG5H7AK5lAT87X7k/tOoaG/PjUQk1C8bbfcBB7ssP08QYobZ1QjAp0ufGD2d6
XSKrYoEDjVjPWnq+lvXPe3AzTnGtbX1OoBwQ38hWykH6zVmxnBNK1JWdyCTT7QWvoNEb8Hu6ruq5
sVE6HYpeoeRSbRxmJlndG/3IAmF6Fnt8T7hLfEHFqsheh4JRENMcaix5OFDWMDOYUiKMxz11g+fa
gsZKQZrVjtEFe5HMkHzqYCmHHVgI9RehqXpuxj8jaE8eXLTXcp0+1ryzcQbMcgClWG48R1/zY0YG
X2qpyDvO5rQiisTusrm3i1ixnkeKUdufBePAReVQO+ivjWsReNRSQ6QZ4mdWxhgOxWHczbxSGJIX
vd+CxBMD8MjyzQmZ+PiCifOtEkdS/QrcHg1ucYUXZpeAm2mUyIKzR65xOVUDFBrnnLif0Ocbhgls
NOYJAx6KsZxbjIPTbMFW5xJRLl3O8Sx6mewJT+Z3de2Mw1FHG1VIGM2m2uB98Pstv6vW2VVpqsNw
hjDC4I987YKPiF/P8ticoFxRUTrjqBQcGnbmsCl5PDp6LKmDXrXnHr4xLLoR4NdLkr980vBbJ549
/2VYABDeh89AlXUkGSTs5K8Q/6EtmD82zYDE5j0qJjAfrIerSdCpoJOD6hpKpFDaJMuh9V8ceeoc
3HsmBmuu8T9BSepeF+XTyPByz+R5WM1JLiKSYCdT7fTygPBMbMYtKKYbTMCnCJWiA70ba0UzoYtz
OyS/UxbgEa8+irWoUj8WiEa6lzLebN0YDUFe+GPQMdIunKEuYdBRU9cF5jvZVjZfHuCmCSoqv1r/
0qxOazvTez8QvMZZJx+wG6TPRSEntWd1hsDf7NZ295f9mdb+x0QpKhuPGwTB468Q4xCHrm9EUYGZ
k86MSJZbkB5Outqkk240zGz77umhMS85gGvZwUVCEXl4JcRGcU+MtAsCAcf8A51sQ4Ivh1+5ilL6
nWyOZIfB6wyG/ISj6BS8XiBUNpPtnYEseq+J2UM7W9l270k7yKc3GYAFK6JiksAzwdBWnClRY4PF
1RMeu1MziUItEmcH3m6vpMYRADYeS04xxXqMp6ZgdjLYH0ZSpovS1ON+MYkeUgrDCt7QshaKUaiG
8XYIzeooJoiQWchsFm7uN8efgzUPcr8ZEHV2K7309XxFGrryyathF60Q8BYVqZ4bG6OSPPlhsF+5
ZnD1KDreAKA7pwHW7LoYD6uXwCtB1BSNyAA+0yQSInVRuTk39VqRhjuOtK5/bJnRkFP9YMdYEnqF
11LCNcYQfvbxZLA+K0jwedfNjaKcBvxVMvK6645ZFbwmjOPbrUjrduJBJitmYzOsaYU503I2muf9
2WyAaI0UUl6q9LTNGy9vS4Vajh8mJaqPdQOV2pRrSnl/zkr/1+1IuRXhzq355nh1ZB/5Hofhllgf
qxibW29pV0nhUHH7p14gLtxNLcGkbaWNAs+aofFOuXdK2zEJMrdXscd12YH/8JhFmmIhU8BuWJVe
3+tJ/pMFSTRAZ0NFrPNtViOtfyl04U/0a1Arza/Y9JgDeI8Y9sWKxs0WLZZW/aXaR2IXk6UGQsIp
1GSkmOdqisCE6QJiqWtSYUNHs4FW7xD3pmx5W8l53NNcsj2BYLEiXZMsdYY3T+jDsb1gOiSzR+1Z
mie1qQpyQcrqmRFw/UtJkkLJnIfYERtu0ibsHHHZS3zGSEtnCMwYLBZA7hwJuUz//tbdK9Qqc+/L
G7HfoLMZFrsjkgmbRIZFyouf6JDTmN8YJjKGM4DOgJMonYdR4FrngouX3b6PdUJihfCAPmtu9RXx
/nMojyPQZuneMVb/YlKxPRGr7NL4jJ73zuuDOS6ZvtmKbiVKw7lCkMm8kZb8W1x3GCFX4eJ1Tfny
brGm34Co/zEvThse8dh0T95ZvHfZS+5RqGW4gCfkOe10sSTeLBv7SzSxL9CF3xjNiKKbj3zHW8xS
QUAEnCfc4wujWfn87oZXF6sY4HThEMhfOfOMB2r4ZSCBSrvSnXD5rNGkKDgCUlcp+ZnleUABZubk
zdSX9fcRGWir2aNxJfYBZnLJm8TBb86J6wrkxpKaqBJH60l+EXEaRlrNZF5YBFIS623kMSiXN77W
RCVhRcqJwMRb5+hTuk9BGa25SIaTyafqKsfAhBcBIcmWTv+FqbDmu2lL9DlyyzHClV4aoCJHJB3T
MjfQXD06OlCZ5QSdteTMWb35oWm5yrghx/vx2+AZQCLaKpwUv/UVJFy0jky82z+R1hHyiGTjHvXu
APqeMdjHzyGJtZRUHvl1Ze2SlFrQ33BbrCGqWLIUCTVEvmQgGxKsd5UoEMpRVxzdffq2X3nI+4Yx
thJ5KSQr7UqFGsf7+nCQ/AaZsNqCJ+uLgPqzHBNLkdmAAL2oFbmAjfl6G1+gP2tnzHuLHcOmhmxB
pImL/mM/k/hKdm9TI1V5F7/70t95X13ow/GcCL78OxRZwcEF2vTGyIvf5dkgXD+MHO60bqloMEtu
/FOpjz3fLcsJXreVhRywAMw2uW4jAksDaryfgk2elrsmwby4RklVDl8WxG2HHNk2+twFRsX6abMO
J7sMx0Z6bssjb8P+6HtIk3TVqdW4u/dG6jbmy5JGuIhSICive5T+S5eYWBXpD7u2QbT29RpEVjii
lEmK7vVQOsBXnSEE1T84WfQOxNuMDcHHvXu17lZYvfd53GtuJRGwteZQ0Ue2F3CL/UlbJBudE8tn
EizkbqCKVZTFYLRypa115gcfQZ1zdNTsj8bi1f52xmbF1HVD1Vn5maNzKAQIeJhYo7+WR9/hNrum
4DueOGWPoKG7TIPffQOStMtVK2AdJB/jq1oZDAvEvzCeDPkW3On1yI7SDI+++pWzvUZ4rZ5ug38N
teuRxvH420DBzZWeysbXX7YjeBt54cs3uT3xKq4makYqfh6b7CBDEU7cxhqyJF7NknJvjDRURXag
ou7C3Cnftnc9nP9Ehj+zDkTgJEv6GVuGn94koIkDWrhKpqREqAHavxIwdzwCiWCXtdwlWpmTgZ/H
FxD5+Ss4yPv6kqXJyXKvavi4BaERWj92UmIC/gBxOu5sIMWXzWugZFxslAcBYAS6Zvh7RDz1XzxG
q0mf4X4ttIgwukJ8201k7jorzq3jHvRr2DwRq5l7DMfH+5lrnnu3jWb5hoVmCUK6h97VSDBZzi+P
7rLd9wEWz4b5nCP49rjajFgcIpXkl4IJpCEicMTIHNwZpoNmWghb745xteAOIB+/kUFhNb53Ay2a
FA+NGnGzKQi/C3p7HTDE3UbMS4jPdeM8aYUmgMXPKr+yql+gSalzlNcc9ajfesz/WDH+8mXV4Sth
ZBW+4vxe9DhYAQhAg2RM9Y65qBWp5BSQwjaZZtUOYzXBwzVoQ7IMDY5y4NojaXtkrbgufVu+pZ/w
qdPyMuD3XHTyyQlx1y/OtkW7X2NZ0rc4G/5t/nbiDX5QkbDeQJm/KTJ/P+CPEfAkeFK+Hln8IiuV
nmHuOMeqRzQMTTl5zBgSa/iBc9HqYxcpKyirKc0COaEw9hNyDI/iu09G+VTvBbcdYUsYnLL0XQv1
sdbu90dZG9+UdwGv7KYJr66cI/pkBxOpuXtb9Ax6aCU0oqi/s2jCXCtnBgtkriUBaxqxPx8P4Pul
EDLhZ39mlHXyXDBK+NoF+Yyr2gFhN/yAUjXjc4oI/m1DZpV3tJWirvC5wEmxjQniMllM+YGtpX4B
sIBsNMWinC7Cx4zpTkiRcDg4qlgZeSSPjtlnf4pAjIScYzJPj3Y9ykhMMjWAr6yhC4vQsD7jJSDI
RTP93NhAO8WaMryLq1yVHYdARhDfX7wbSfEJDgXT0DvqLQhVSJ0wR6bzd0X9fqKfxCKbjJJk1JQA
uSbuYAijcYamMz6ll0IwkOG5X15HI9ikj2WnbCHyfSE5j0BMjNiLnsrVxIkrRgZEAJI1OZsX1L2w
Vw0r2xEv7Z08cdR9ZQ8dTM/vgGWD3sAM/3J3pNbW+Sg9hATM5ZvhBGRocIvjN5TF0uqqel90bn5W
JcVc08DhZqfliHrdnZgqEJX0OhPONDc5BmAfTilJsHVoQcjVLbDkGjN/GRvee6mHbc0N1TqJwMWq
SGt2NQydabUCScwcWwvFRS0q80yd9rVQFSAIbwzqy2h/e0QL3NsT8gvpMOeujYnEXxgY2fFByNda
MV+WajxJQzkznt5AheXghQE++KZ/+LVO+GvXTFLwP6L4/XwZfsybNOAZ5eo4OKCeBYKKrlg09eZ6
aPU9339QQakCUSXndmQ5G33DD69tt+SLl4P4aRNbVQgIFY7p4LOoKnhCP2aV3u6AUHA4JOFmINFT
Fw3a89CgUhegKYUBw7NEiAkwm4Wjj9brbpUs066L/TgK0+xtv69Q2E1Hy9+pEO4b4shDdJdeX59G
VTyRK7eeHLyNRgQf8WdZNiqMG7sXyYa+KHvNv7i1Zp/OxrJfDpw0HRHbz2ttnNlUS9tsTTXeSdfr
Vgv999cQ7f3PKaoTMzYerbp4e2gtwVlfvFHVSBOeM37MIvLLnZDyMiI57c1eHRPX1uURpKHckVlA
B8oY7m/2tCzNNakwTiy+/YNuSQBh3E0oe69jkR15lqbzWS6K9qugTSqlkdzOIqlbV2S1lnDv1Ry5
fPcGjIQgxAMszHFGwCl5i7KejafnrqAT3ZPfUwzC0/jSDVdp9dRySj96WZaRUMNIM1slq3KnWm+r
CVBT80cJ/4Oa9/eljnWXkg9HhZ7nzZ6/6jk9zdaDCQAoTSe7KauRnoiYIeAuNBl7UrHVBTXfvjQd
vsLlxfHXBSL1sij6saescyLApWmEIGq1PR3fJW210GerqS8uPs9gkUQ1zfeNjIBC9CEpjOV9M/JX
Wr+FKjisXXQsooiRfRyR7Zuo/TcPGUs0manoMvnW6XnJ8AZb0IklwAGmP4NisuS/cXmreKD0UgAn
7MnwOP7O9FGfw6MGppx2FgU0esy1qgW5xzFwLE2QCaYVPHyRVRppC1LovtAagwO/0dZ7O3wF5Hd8
n7nR4Wow+uPazTTcOxKIYGAR+cpH/nNUqh9ZHmrA5LC8k0lj0C/0U0vI+W6Y5eJNvB+nF3DHBMCW
VaBIgVmEzVWc9QYHu3cptaOkWeajJ9xgNjBAn+E0jAUjVpmZWjNXb0De6UredmT2UV53HKSs1/pv
6rSXkQRGrftmM4bdoFnNMLa4AcQYzjNsbu0uM4Ke9yE9Ir/xib4fyKKZPQkE6bBFIXGk/vWPTOvy
+KrL5EU671cxnxNpG8HvApkS7AwxCgfXvbyTxUOrxWqNRHfs4dpDCbo7oSJN6GgxM4CztzLweKlM
6eUq80j5AiQv8Ks7tvQWQFX+XF0U6ZjwVwp1QLAUBBnEExI+iL2zvMhOfbmPGfuLFB5U+EhR5g3T
YjeeWXRGieWOTk4We7PQSqa7q/STwTgAC1QUC1en/zjB3TDCeV217ZRCwBkcy6EBAPCX80o9zp7A
nwysvnKPaTNCnVhrivyjUibo7ZCNlJ1qYEzeEDVG9O5ffuUavAfZn1FDa9MKdeUHJzFtHkGUn07/
/yZOPEW3dLwmHYgy+LUm7KRwWQxbToOn9zjLQdqY8JAkSAROnF1Rphcoo2pPr0CUiSBex68qXGCz
ji5AOb9nyLOq6BAJy0H6ogjNogCN8JON3+y6uLNPUctxfai+GhgcMkZeCDUT3sR178dmhUZamxHf
ef/HqxTpUktrBLAD2NXO40QCs5mmFiMWFAm5CmUTegsAKyNZkrEf96ajrR77C9WKJDtSPGxx7/Ya
/+5ch+Y8SrLlolbu/SZ19HW99D5zV5GyayAhW4d3ZwSoV/6YaVGhkk2ZrhLOlhEB5R5tIejDmzgV
d5rUZb1bxs0tmvV8JDsYBY5hVLTaGqACHcrK8pDyznCmE8I1isA4VGJJLwtZIke0mcvRv8Key1vt
Y99g5uOV8NLkGSMCWyKxcRXmFNjJVM2l9tLqtvWHwTCWB7FbUW+E6NBNebIVg8bSbkh/pdbIwqCc
T1q9weRt6y0GMYDzLD+x1F93rgYI6GLAzHgdyFe8MK+wMlNQ3M0suBX9wHngYpuuVDKEHlPz/Cgd
8TBoJI5uxtcEFK9tnYjAVqeh8cDBYU230FUdqWHV/Hca/A0n7eiYwmTDcg9zzCUG4QCOmZztBQuf
uzRL3PBHkzeHad9kqD7VUykur8DJFJXanFZuQPhhh8LMeLavviRDPRNbhkCkfyV9YXH5je7eEo9w
Og8HbhXJP+On7npWlTHg0FL69V9aB59pFnVzoQqrE0TI47zQx64IH6Ju+9GPmXkwRNX1uZ9vyRYK
VJG4u/g7P72D8d7CkzmHTUHWXX8cedabsqdPfW1zmaAP+dCs7M9YoUC5EE69JlkjXHKpVdaNDeZZ
Bm59PWPwYReqKXGdkR8I22CttrDjbw1+pJz+gniQrKnhW/9WL8rXrKsueYeoGcJqBx3xuKPjtjPt
4LiK2PXNXazwLNvWGowcGfHqd1BXc2QODoY7ORnlivvurO/8spV+0rdoz9EjnpAu7U7buLtMVB37
LiMzNOrbp1YQ+RDQGYeWU/nXRcGlT2lmL4Nr68chU81RnawVhMUcMqxLybqG8eJmRE+PizOX+yBu
6B/u9y3bMfrWg/TUXOLEGStgOO69e2cYQFAIxOSYdER+IwSeIfsqYhD5pK+eEV6IUDSUCNkqFmWt
Cdv3SRI/03e75v+Kmjy53cOet1JJnFs/AZHTLQ305A57egL5oSruXKFrKKPHmXiDsBcIlB1zz0J6
TPjca8LOUZlqLN3xww3VtwX/ivtx0rP/JR3f/sO+rslxv3+8RGVXM2ZLNCtmBmDIH4DjSQaamD5l
wOLeIKrh5YIhuO2qCNKtELBx00yOr9bIcVy009udZktioKkgMNMFevzHpNw0MLluDFmI57cww6Ob
7myhuxi3qaNLdf3ysLzQ1zO4Q6D3U6nES9vkW8r3pFlFGDK6Dsm8/zOqYDSdy6CBrmOyc+RyDQnw
8L3IInxacgO+sCRq8D0MPoGeeYElE07azImXs1UlsA7NpF4nBnj7xhWI9pjWsi3hK/KR+lUdHkRy
6s81mvxdjEjWfjRxfCOLBqmhj6KpzYqsIa9i3AseCGBxRndObg0prrK5YscrLB4YrbZ8rzKkBeDu
YZqLjihlVP/s1V8gmXhboDfjdhkDbF3iDWszwG+JROTKUFF+XECVfG5z+WrROaEIr3JXxYZ/G1qy
OTz2SKt0wKgnc5IXXAgpwpSt8xCGk48C4Pwn4mS8zsIBdprpur/KtPt5Ivzz6fPh/omRa22ErtA2
lIfJOCkskTOx6PQiZdnUV32oqNS4wHIQiIIg7KF7CpGQg+7xUhMdTBe3tX+hUSINFzSZPYtZVNi3
STRjzs9xm2xkGG/UhEfE+hQurgDnAcqHO/X5sipRhS3olVu8U5mclRpCpdC/4BRrsNfNub+R+QxM
Li/qWaNEL8BHVsZ5qbo0D5CRuAF0JufUnG8TdUAkVZ8t7MmBLHbUInSnSnAqAAI2Hss9qJfySPcY
q7aMQ72eNyf+L3Js86S/pDJLOEEbQ0+vpfkS07QriAwp0HHPxLUtxEPy+AhAd1GdvIQZDAU35x9b
mrN8MBJzzvFaKoOLQ/c3b0d0wc0bPZ46pLYNJUjLugtS/WURQCV0m+uyvVQiC6yv7i3VTOUCclyL
e7xkVasRhNBjyD/rP4yaGHdLmzoobhMnd65zOddxcaSI5ut5HT9+TDsF7OcLtF0f6n+JwTs+0ZMU
EB5Ub4Dn0FYrg4C9qi85KUhL65GWABdl/TY82mPD21fFYzZz373r10QtF4ulJ9EV0fBhA7+lIskm
RE8nzVOleeiOJnKIs4rHRfuuYQq0hyReEZiRtMtaYTOiK1c9iGraO3rT+7V9/HQRX5ewTa8xVAnf
ITG0l7acE+osWVKAWseTuwCCNDMkKXIiHTLRwK58+DNSGILYYSmBh85R5oLcLdFmS454V4Y+4uxO
U96T70IPZfl95/le51I2cpsTYGhWBxtp6wzIMDsEXZsK7uBJg48pmyXXiDcAvdHl9/uQ0kvIaIbt
UsvOST+LzXG19B3sHq2ZXQBgA2In05IodyBdAZSH9j3JC0s4QD+wkjUBJP1A/ZeuWJb4pXg33SgU
QYIlbLC3oWaqZzC4cvIg1qm+cQbZdRndPQwtyhCAkwRBHRNXcCJ8yiUro7Pwe+UeTeA5J0PYkr97
fFqJQW/ICcqb1Ix+socMDdkH0YMbNpMaUTV9lKQBxogkVl9W1y4MMJqNJAAd+PpXMepYezlOpSR3
B1EQ/5cyecsBvBh/m2gtbYbwZcE+sUVJQkFL0+RdZGh2hYCSxfw6jacjE4euQK6snfDswmziQD32
NbE+Di3h/pdpUSunkwan/VOiH/2Lg009Dl7iGC08XgNoibuuX7BGeE8NLHhcq6ACa/4eQDb/5xSg
bT1G1OmkulhMO6OEf2rRxGG+hrZp/ZQqBVuNfy6zTsKBBWjcmQnaF7AHuwUbtcD2pAxqIy2bVqOQ
+IyBwjiaPVJv0PccKpmyy3aZuzDoQ6PAL0wNJCRkopZH1sQWjANJKDFkGUKGjokxx3kWcIyf2X5s
N6VwATB5bz2wbnRJfS0GGnzHBrC7aHAxl2+8yX+BZm0fNX4+tK7rNsVrmRt6Sin45kfY1nVS1DUY
I5NUNaCvn0wOlpdsZlgSi9DYv8MJ2yClOf3WKI6/hfAf12s59k5sKapnBK4o4QrnoCuHxEyK3RC6
1yQLSjh7+7WcRSCIlZW/p6uO3/R8GAwC5GZ4n/GkwuY1RreiVJWEs14C+CzwFiPXckL3U1NuX1hs
glkHXowlA+6gs+jJSI5HuZtpxUHp6YQr+kGQLEeNk4dYmuWQmQOuV2T18BF8I4jMvg7d2pNyZ2x4
bvYGacl0BOIjemmbjH5YBNYa7VoglkV5IkpxRer0+n48gi9UEYoaKNchQRzXZr+VE8f7JAtWb09v
JTeVxI+y5tEDXqf7NE1ISj7XHovkSchxWhdljat18XCk1APs4eThHsE57lPG/ghEuw8QC14otJpm
CjMtSgSf9z+YPozO6IJXTClcDZTxdsABqBbAV+8zksQhsNVkQTx5c5mQbyuW/IWS3CcY/zu5Y2A7
XMj3CscdtlAbiuajb8bqHYgdzdO0MeYroC3TEZjmZ3Dxshd5pjwKsCxjkyQCMCp0fIAGonZUY9/p
pzlt3BtEekI4/pDMEEYXpI3atFh7BZ4ubPIKgQ1rQaHq2a7HElkfdjjLFVgv4QPL3pe44gAbaEGO
lYz7HnwyAtakSxRhdNvQIYHSILhlER66aEdS5UFVAzKwOZC6gX87fD1WFoNgNgDCP+OvcLpUWGrZ
6Ddau/qb09JJhgurldBq4B/Q3CVTAtarBYDQARfpiPPyzmRSBI/zBZe17pXacLE0aceFrEI9mV3R
LzGfkTogkJKAcOcMN/Fgoor3PjwcaVaBBgN70dYgW7FOrkrzh732KBZGJT0N5VbRKAkJMZay7M7+
FIhJqOhq23Evyl9XxK2W//TrDlywXGJlrZf9TXAe3mNAztSCxyip8bBcFhszfg0V2Q90e2FxsanU
1UESanw/dV76QbVIaDTKOA39SW5ZTjomuTe0QreDXLteBr6Mx3o3hFs3z/FSwgdrBDBdlnF6Vi0g
NKOhn3Z0ndTtlEArTNOlQwFshe89bQ3GuSL9vpnbZ6vvCv2z/86BcWkRNMRyKCLl2N8P4bc88MlW
HGAZu/jtrk3+cu4NlMLtpgDbDDumGPD80HK6meDIGRcY0csrR7y4AjUZiiqqwqLDi0PkI7bUhSuh
VSRRCl8eT+toD5tszFHxQSlu6mDutz1g79MhvCeVLDvnHB405cfDeS679Cujz9MDKz/lJQ/hC9Ty
Y3M3YNthIjmGQcARHRoOlKhEN5972DucZcWrxG6w2HhkiRxv05yVcswANk4hdhxWknDWDxbF5YQ5
vxdzAMUYkgk77BUVy+E4jmnvNz62+ZQjDJXs4FRj1+g9i+heI9zpVcQQHo+NKZ7qU2bfLhwb86IO
0D1wmXUG9OfGd76pG/Mmpc/p1KwNj0pznJsejDoY6scsoDy5MfIRyQQIl7blpbhtn1V/C4RxLnd4
6ogAOHTIHGM1ihQkmMQG9awDMtrFrVgEYaYIAPbHxXmQ6V5NA0pBiY9jllPToUQ+uHXUnmAiN+eK
Oz9ChoxcwqBBOTCR9txmlLl3sd/r1G6P4iPXXrzb2fzVxRzEI/DEoVmFYKgMnDlRWVrJAlSrDZIx
BcR5wHsw5+S9/L1WWLXdwUPo1YTczbba0Ymzou7tEHVZRzmC7c3lxO7u1yqQ8KnnC8mj8q5frxtp
czt/8cyiZejyCNQDyq1sagyJxckx4cQjkc95CyVE/00BDAFCAFsQQaJsDnp/f95LQ3zu6osr7jOl
JjjJAulmgkD+qhUoLbZDRRlw/5TPU4ROrgYyvLUDdn5zS+98l0OLTJCuvHW3sVh7MQWQ+DI7GOya
Bj0PAz/j718kxSYW0JpgkMEmn/w9EyjaK1RbbgpXLbWhrKZaPjq+XougTwh23y6QDuveclETIloC
vMch/W7MhPPrLvKlKzQ4sDQWVCEIWKiKUQsMOEc+7uVM7wjntnh9pUZmBgFwLh6l0HBkB2HS+VVN
kNt7m53uDRNrquqhQVYo7D4IFdGrzsaGhRQ5J+t3/BJ/vqXGPUwLdBswYR0MKTaTe9N82bEEpEit
PzzU70Dxk4hl2b3PwM59HoCHN8K/snee85neQHsTgLjrTw5Fsbx6fAjDji3dIjfLIIkNPUfDINx0
o0SaLbhVz57P4I2YcCRFkgvpmgCqfHcdIcG/xeFb08nCdjsM/FOEiH1PbAGdn5kzJZHys6PTt2ye
gxcO47sg+VTfq+V9l/HPLl6g5RyrR5xFri2TaJC1PNfAXnlVACbeX90MrDkegluU1SuLa8o0D0Vl
9ZNp0GiVqWLTy3VX5otXJjuefkwIdNDwMBDDA/6r/cMFlrjrUw7xaNKXG2LUVvmgI3mSO+n7avqR
/UpsmW8Oq9IV01PDB9lGKLDKnNU7bKZd8wl+iA6tlQJQkJdKUGtwokDMhi688fmD1YTW/wG9oAZ0
Ez1shnOsIcpEWn84Oh025llqVE86SJaHGjZmHYFlbE/4mAe8X675MsuS0Jv4y22NB6Bb2BiGof9G
hJPQ0uuhgWaHtUpRfpI2OYzEeIJ+4QD3hqcim7TwfvZVC4bKQ6xgjypz0R3n2iVPb+Rt0EL5loDs
lPipbHqjeY5BywlfrpmOucnokd2SRaOZci58G5rL9LaKczzTY5Qo/LJjmxrR2t5JtRy43/H2OSa4
vw9otjKKG0dPxC+ISdP61ykxg+1612gPDjyFBm5NX/RCzXRjpT1MHmAFhsB+ivLdWBpi29Ph5jGh
C/qJVSu8APbhM02k6MUNKYmyJl7eurms4FyUYF3gS8gmd7/hR7HmmcS3ZtL4gkpC4dvB54GrTgvx
cNxV1MbM6sFU0o9W1kNSoCbsjTjNpVx77C5y0lytH5I7snyaA4CR3Xyj2/4ifBJdOCjccEBm/gM/
uRcJZGBrINVIbRiwn616IatM14xsztmvN2MxyWFHcPAB3a657nhJM854mw1uSDQjujmWZ27OG2Oy
tz26yJZa5gxhp4J7mXMfr2Daldfziw6sdC9/gcjkNb+5fxGpJXEihwATqHY1wd3Z6DyqDo8BkZ8X
9wJQTr3mq9BTzLc3uTWKtXS5jLIdIw3TocmwBy1JbTF2gHCYVrOrdmCCGqmnI9j9W0Ps63BHx4qA
arvlduun8jKzwcc3xpZ8bIOYmC7mbKzDQ/tI2gayev6Ul6AZUcBjjbBaorylgdLtsPEjiPRwGqm8
L7FIm9teXSA6E+4cKx5U27E4ysr7/ifQ83efo85pe1GR6oqgC00uLZm/xG+rgJg3EZR+qPoB4H8a
CEmmEgY2/ornqcQmMlESjiSS9YGCrxNtD4TPvrvaNyd0k6nSEC+2VfslVqm77suPtnw2tcnUeLER
yQ5h38uzDUWiFJ0rxfhLfETYPwpMQdXRURb4U8ny6TuBMD9ePPuSEHkdMFot26Ta9i9LL69aTdIg
o7+Y+ERBpKLRZTPsel9e06kurWcCKCGmKLIFbmhlpBhFLZdlJPImcqo6ZGJR3WR3a58+7lPsPY0u
YuAt9MBZcDSXnYtMK/sTJqSm0cwAT8El/gwLdo0wG11Hb1mLB8IwFIoMZtC4aT4flmj6AcLmD/hy
lV2AGX3XTPBRY0+NnZL1Il3bnlg8bpyTTCR8shAGlhvVEBEPxaNMtMJ4vvRFX72hV+uFB1cwWkyA
XdyocaZh7yiBnMSDw806VNADA48tF09N8JTTRRkdEJkFXW6QwNJhqHL+2RKTmNmxGW2VYIBnujRb
PPIkepNh+kL+/t+AGC1mq/YTcelE5usICwDkflTAV++wBvik7HUuhVNbb3POPacNkDo8nFo+WGYe
849Szv5SAbbHdCfr6h/mUVCHqM0Lz2tFYdJRiTGC1Socn9tviByu7cyi31lbqXCouap5NHVgexF9
sSt4enO6iMh8CieNZL41zXcdBP4lKxws3rkCh6Rp5UuPeR4bss0oHAPxNCEG4xPo/S4nUyxeIpEJ
owHiJ9yD8X1xobsWLtXH0erEGfdNyghJCZkS6m5Uok2OzCIaK9MSDSw+0KttFigTpZ2UBqYSbFYb
Z9uFnT/UPWn9+KHwtXE1jeWmj63HzkPucs/IxVtBA9U5yS5wvjXuxPCRlNmNc8j+NHL1zHV60NWg
E4IsY9eeZWj+UwE1cCujzuUHcI3vaJWM3slMe92HDuN5Vej3ZOty1QmdfMpZpkkgYeN8aUzhrasq
CyqACdkDygLDOUFCSfbwjKVM6RNZyVxsegsj+0JQdsBlIenHKg2U5S6qIpbiiZn0KN6WlIwbvHHk
/TE1ukP3Cnzs0oRCYA7dd98XrFHe+5sT6xuAJTQckm5WIGfaQpmXmOVLVXcqn86hB08jLNGWuJT+
vhS9fe+IiAHwNcH4TTRFAVPVDYvbuMtzrZQU/1y/f6xQLMjYjQXt9H7S8TO5jOOTHU97ehAxeW1a
3DTRhrldystCROudJFS5lC7+nGUvomOus+eXkxRx0/NSgak/28uzUDzj1piHXbZuEnL8WS6jKcuA
zsIK8iLaSJ0cN+W2lKfRsSabYN6dkE0J2awKU56PXPQZea5YIoRMzJH1ccqo6mmYuxXwxSSNNBUL
bT6e3nXtpg0YWIZj4PKtYci1ALsKkRpymr0hRurXiZmi26IbRwgPF+SJku9q3RVnNTw5mqbBZf8+
uvkNY6XI/Cd2sY1WK98jsVRwsw7swju+0HrSusoT+gZccSRxaYYJBZ3qomfM9U8CLPhnN+ubkK+L
lbQSgZ9rzEKRpNrBT34qxTOlUKxCPEi4eqcI0TgQEaWGhpjajDxxjBVacIdtEHOuh6Ocat8tx2RY
VntCrH6YPEEDh67vwtWzIyYKPMVzgm1l++tmYkRAMeYGS+HPIBZVVZRwGyesrAzUFLxKUetTruf1
tGN2LawCrAKoJIVb2Im4e12Mx9pVBhyUJtsjAEkPysqOr1pqdC9tN/qPbzVuXAMMGoCMUgMq+lid
101gF9lbqLQrPsiwZN2YG2kXSzpF4p10ALUm81sok6Is9EnNemgl4DiZcTj9jh4aYhibga368Uw6
Tnh5tGFa5Z031uTC6Mqv+qS55n3oqR4I0m0LkTagd2VT3E6Dq4odTVJ5I+fEGWhub5I3ZOrH3RHk
i/Nl/ilrIvqUu58YU9YFW3UxbbBg+GnNDqKUlOX528Hx/kam0s+TZmPCx+CflMMEGefp0NE6Kf3A
10Rcp9V/ctO9kxHU3+TwfSmBvaz9PFPfYFAwi+LvRhFxd3rcxb8X74GN57LzjuoaLqoFLy3dslr1
hOPZvqSv2oBnt/oxPmCqNTA4lM3p3rGPBo9/jBiUPEc4NyyJCCrLiZ2li4Vvx18BV2laDqTLyMvg
VkbJVVT8pNAX0DXk4tE2qI7eF7Ek/MU7fj8lwjg4KnD1bM4ElxT7sbMw2sIDSD7fVIp/WQCE/5Tq
ndYJp5V9mnMCtdcmlzbZ5N31kQyYBGkQeL1i6bojEuBWV4f62wZxpX147mOekXXxSuQrjoLOn5zV
Bz+vPJmckd5yFQ/JarJGf4ecnNkcsdRCOl/6qcN7hHPrQRe1QbrPEfoHLyiElB+xnajdi+kuudgL
Chb1052UxTF1s5VL16E+FkJrhJS0wjCxT178XTmwozJVcq820SlxQMMAAKVzssL1hYRKq5sdq7oN
qqqI4y+co7sTNKH8jbeC7IM4UzHAlNP8h0qN3iSETn+CIpIXSmEIHjTxgX4e6DCFqBteGAEphW45
3BBHkzBxUPaD5G+3gDqQSK0QzP9Djvm+GB2F+FttJyGRL+pra64FBya/wtiFiUYCZoMZXzQ0ufQV
14/QwAfmZW9ddrf7C6m+aNsnj/7aFUsIx5s2BWzoUGYJZsFDEtzLy43R8ZhFoC1zXdyUkVVKefgZ
NgZCBA5ygmm86QV2ykqevB+c7syzursGCi5rz1UQ/0BGdKFFSkXZXjTDhFssAq7XHyhsulgP93AC
EPaOGQL3JkfXtAGvcl8KSgHReB8jmC/olpEYxmtNYkgR72+8RMfy+TrgWelVmc7UUQzLllA73QuI
8+L9rNy4ykcVhBGQIDFwR5DdddL+H2+foKEuRuyafCtDozgR7NOMVIquSc/tmAojCLNnXhB8NjKv
Gqt1L2pf5S2E+kvNK9X9kdDmZry6izd+IiXUEbpDA3dOVHvS+ZMMM5IgqPdoXbEvEu1UskaG316b
59Wp7s5wcOq6eWTpBrMfWcDr547CCTMHoNGMsMru0U//kr4uN5Ujkgk6V3N1gW6/Np0xMeuRk/3D
33lDGsCGoLpae9tkCe8BFXAxdt6BFjionckblcZkIi9TBbVDzgf6jxcKCaVSnHsgrOeCXL9dwc+7
Vi9FP78YBN3KXINrvjRsyoGmqCylmGndA5vo1cxOodsuHmqzXComCFcHChw+LAMWRprtaTcvBNjE
02cKc246VWpw+6SYNK6d+7hvQVTy+MFdNPSz+o2EvnsNW727tBgG0T1GlkXJeW9PRpemikR4mm4D
/Bj/zxK4VrozwmU3R/EekVabilxPPWlShYJ24qa2bn8kd0uwUFv6qOQDIJQnZyHM0CS2fEUidVk2
PjN3/p9V4jjDf10wIixfGGuy7LxjgoCnXWLi/OaFMylnuKb9/7JnN1fAO4cZOZXAB03AtA0qXhHD
VoVXiuhhyPhitinp3qOYov41jgQfEoA8y3oyniTFIPkK4aoBjv8tvQVnbxOk1GDp5PMjNVe+JeRk
IjoD0aJJLXwjbjLwc4qfb9wuEjo6Y9UyfiFhiBUO6tdKIdmBuMT0pCS++qbEi5nYTlNaffNX20Ap
7R/ma0Re3vIAJpRb1mOm0SN15AFbfFdiYIC1+xwyb94iNiHhRQzX6JGXlzoE7/bEaEPEvRclTRVy
N9RWy0pEDi+kqq35qBVqO33k9ErrFXASBZTPiGbGjMBPOPZORXMPQiBDAN4JjLfzTKndg0ccQ1zl
UeBbb+WRET3+sigDoKIXUfnjjt0tPTi6SQUy4qOWvLp776YRIo5Yo1dHs0ac++8sOOTVLx73du5D
oZcnQLyV7EwZVF5LlSblZXkvaX8r4BVlwHPRkbfxEYYTLp7fZ7geQjnMZomMSdKqn8FJ6gNEminU
6NGrdLZGP+YMe/lHDdjicnk9thTEcpMTsaR9i2eB9tNwjXrwFH160bh4p2oJHEdWF5k86gnfkE9a
8HPZigBOdhZUzp8cNVC780q4Aefju/o3nnNMZ4uAQUtZIsxvuLxRPDlkjfd+3i0ga+hQ+KQqaP3R
NcMiCSc5CiXo3vyG5Nr2xQF40MDF0OZHPrDkvLxuCppKucVkHMt5Vzaegwz8qrF2rBdKHnhj8sG0
Y9yzI8OoOQmW1J2OuRAsxWgAWjM4ieDy19EDGhzq5VDA5yfTpWaQrpwWz5644S0AHUnIcH7L/rQe
gX3rzAp0CN05af8FUSSRYkFYlWaPbefZvpvqjpqpQZkbldIiBGN3QwKnL4u7DGkK1HK4MjBU8UBG
752esKrq5CYgGZj3hXcIrAAA82NExrx4w6BFTQyKxEvOhgU8Gxqn4D1HmCJ1nzAS6LchvBN6aveH
Yp9aSWdsBfrj6JUpwhUQRp50RTdfI/3seR43t+388zO5ac88OuPZvb1zVWYD8O3l2IERopxpYvb+
CXTjDoteSIXjylq9KnZC4+B6p50lWJ85pYg/hhqmmpG4WgXMBePXh8z8+VzgXKriR5MKj9gqqvpT
4HrSWosTTnHcycucCOYKMQZjeOm83jB1wGiKjCVdw1XF0AEU1oO+kX4Orr/Dfcpt/XAjN5LjII+7
S7FTaObjoKcGfHKXUHWHo9KkOVQv1yg68S5VR8t8ydf7ZImzffA0fj83CQrKH6HzPDBk75dPBi/F
goR/xuSslnPjgcm7y5bt4xZEJd9ekY1UcRdxWplI/4Lz/e59clqa03OZ0C3BCWUn+FzT/suOUciy
VO5PSy8DdO432YDu2vlE5/CSX5ccFvdGWouGM/+whJ96qrH263FYpov44rl5mEIrclPOEXlMC/gR
oimpdrUhg0nBTnorytS9/uYHkg/6zG4k/mwGSRH2fwnrf71K3uEDM+ExXDqQrpF1EdujLH7bdxW3
wvvlG7V/C/cUDwyP8zpcweagvGwrR1xhz6iW2UIG2GYigyUGNxtwXb65vE//JI2WKWkS0iHyNcL7
AiT8Ic5kgnafwStvnjPZu1hn9JYNFu144iUrhmVhaJsRJxAnlnDH50Hde/y/hsFCW9dzxNJWL756
b2pWwi6c7+rwUI3p9lIpSeDrXR3AITj8Bh+tR/a2d3NZM0Kx00oJ4893LaqBpO0AKAIEAcU7z9z0
ch1k7WPBzMW7zGeBVl1Al27dMmlxER2Vd1/Rm8qIOEE34EFx85lCwpqqvqfS0AEwV2gDj2bLdGMU
YhRjSFO80sH5zWBBmkWvXG9pUw9t33Cku7syGD94dnxr5pi5UvrpZzx8dqDgnS35o9o9HQZnmELq
5TN1Reg6pRMp/UAvK2fxKRQdY8op6EOAesirslDVG0OtsXFJnmjBO4101fD2VZqbblarIFrE0APJ
HUiytJpZpoHIqlESnpJ0hbuTlzBUfRUEjEU0vjj60ieyDEQeE8I2gJFurnZdOI3ucdl5rYaPEOEV
6+/9vOj9IRvMICIVyQUZBAWEopcrYC3/GENu+EHwV9p0lQIC0S9v9i3GGNwuhSb0F2QZVoK51taB
5fsqHPk5xXx/KplGphx3h0VEziwNueOucI65k7oIFEw3PFpt8MpK+0RVlLHRRAhFiWHYUuW7IBrE
xFVAD/LpZvIIl81jOGGWtwcTtyQ4dRNQjD20myYEmM01A6u6eGVTsOahtMvWSL+/WuGLkYo8UmX9
DhFLdKKZP74LQeSmq7LOGK6JcFfGXIimMTcyPFch0Gwwap/M00nFGrnPUJFeW6A4yBnjG63SSLC3
DtWcP8S0E++S5i0dcaCdiCzLH+oUm4iy5W90YULHp3jTn2sQ7d/uXW83/cXIZrAqAxNUWapRRFDf
33qV0OQjalZgOoJolBG56wzql9HEexs3OSA2sx6Viin3JEHaH3LMlwee+STLnS2nG9gKdTwlr6IS
jOk4ksZu9YETdO5h8G0kNIMxuS3QhgW9wKFrVwYxK69nNdUnS2IFahuD2HTRFG7TiAXD4tpmPoM0
/0zMZBZ1lKTeOZlfk6D6lRigQOUggJzZ2VDGK7h7iQpBMJUXkbbunI6BbUz/NPZA2qWsiBVC0JaU
0C+dk04Td3weEkqxrioeAbIb96gxTRHbJZreGPNbmLqcyXUUsFFOZyJwNk9AKYQuZ7XOZoxnjxIC
u2UvKYwfaq1KKjsEEL96lOc8IVvwnn2Dka0yH8AI8L3P2V7fKSJUjDpKHq4r/jb4ToiJ0yfl8yBS
7SDJXAn6WPyj73YLbMqppETkbn1GTOjmZMKZGjUj7EXSEiCUE7ZzT35F1MtRUHkf4bU4g/GzAT9Z
bknBHCSvSYdj/LhOf5YvTHZMaSN6NBaUJ6I2G5ElAuJQpOilR6SDKC8eps7XAdZ/eCJBr+Q06RTC
3X3YY5J4cv+YmuDYEhntATHzcg77I8176k7X9s/XyQ1FltpPd/o9RjD9XljE65rfZEZ6qL7ZgFJc
zgTM9x9Tvb6GlTOAvEiEo4CMAOMt3K69+Oq8780yp7JDh0PjC4hQGgtMJJKOT5tkrEMnYJM6WSlK
jmcjuYCm+jW1afJqCXmQdkgl7bIsZFsnG9XK/2VYIg0d99he10VNdN7zw23fWC8S6bSyfNQ6DYRT
fUt3Ks7IwDlLowRv61IFUnyuBOdlcYTao79f6RymmwXFZZjnZK+PWTJLkdAHYuk948t6mF6gfPYd
b02/6sdljij91J+Rv7qPmiRgmQayvRXdp4DB+YfLvgW2a8vEi4CUn3nfPBKHq/erODe0CRLdT5Kc
DworjA3K2PKNCM2Id4ilbU0iBJPggIc+/rR+nNl+nPo4oLvMxiSFG7ABVTBUXC5RSEtMo9hRQoKs
vFUk8ZlMIkEPG6DJ7gLwMShcTYrHVnkbdh6vu7hFs6aIVGpv8Wl0musbnUv34egBkA3D9Gne2hl+
fvZU54bTABVIEIbw/5jyvpbfHUYY1MijXn3bbIDSgEKb7MDyO4a0Bpjm20zz3hgZ6ncDMWJxwqYx
TvsKJfGUoIKG2wXKleLKWUdi4sF1h+WuiDNNPgNTwiOd5zVkBY7JjJwLqpWH27UC8kSZCWNbGd22
YrlTWa9iiyiT0NtjTNKnfT4etQ5kJFpD2UhVwaOSSdeIXO+eQnqa4MTi9JvS9OiYMt9wquHYbWrR
PpubyMTHW6FCZVtJNVE/WLaytvwegT7v2ouEFCw/TeJdJb716eBnaG6ZqU3PJtLUPalhWxgHACey
3xpOOSm85rhhARHx/Ifcv1lzxoPgaSXwZoiseY9mycqRSw5u3PQYlJ1w4aykMA3atc8dGaK89ECx
LIKzVxYBd0j4eLBnuaM7FKHwhpr/MEWNeGw4a0/1ud/DsCPTenoYKv6LwpwGgV0PjpTfBkBr4dce
Xvul01png2xFPoqg4lP5jqW6nCB0UEWOyokz79rgphzuXPm8YMcOAeptfeOMZk5+r2cWzcVqsg4r
iVGPcaHWiDoSC/D5DwiwDCJ9EnJ2rg3PSrrSfSTDlXtuOoDhVuaaIlHfnc2EbidCgs+Au4aPOKbU
PGu00qsewzwb7aKrwltz+efMtSEGtVp5JJ39x7JWJI0H7QPMk6g377AomB61unfw7oqqvzYvNl0x
RP1tONeHrg4R52u06POa9cOsrcoa7byWP28LRhM/eFK9qMgrZhPMkQTzKdu1Xr1ger4juzqQmz1u
mMbzz1ivFYoZkxQZPAy/x2PAV+s+lfJSx8BHMGboQwgQZ1tsXGyQrNrORj/nnCZZHtaBtV2z/u0J
BvqMfBslEdLHU1SvPq5m0FjTcOVG9PNknltk2LNY7oRZvTJLL0C+iCJ4DFfYpC6IASPST1RXuKxY
O9Qo++JCy22voa7IrLPnAXX8/IdI9p65cTi+puqr7p7gLzPAS/rCnwvCK92E6ChhpVH9X29kZAZX
pIK8+sSza2Fa0Hjh7uu0AVdpAoLnMCvghCfoVlZafDyHJ9QoilY1otPv9zr9uJdCrlMaN0r86vjX
QrkmP/TAy+SUiDawTaDAthE7pzpDdgDO0P1Q26QAE4uxTlNfsunqn+i9ZYXOf648v4SKbrUghiwV
Svvtu+exkFUJhaX4tZy61F0GD8alpUTkPgotCobK8Ul+qsk6417NSXtw/mb3Xh/4OAbwRyLghNL8
wNE9g95St/aWU3E+0RUPHkwzJVZOXJTCyJACVlMItiXHN9PpgZq96C0GPqdqjnaSD6brHggmwsgn
z046NYMtfpxD8Zu/bJfD0JTc1KUEI9XAi709cAC5QIz9XWkUdpg442C2xQBEGIX8zZr04VIKe0wf
9nlTEamP+Zs2bvu4seDNQRpQ2O/B5d1givsI9O18Ee0V7FlRZJWioU6e1SIXZFT9AdPIhdRtcF4Z
TBlBvZNT2q1XVAqTYKGJ+g/IHEMm14pDiTYuF05xF/PkMA5AcviLuDeWqvsJyS1HgTrm5TIwaioV
Yq99U7RyccOTDOUn0gng0moP3sD18CAxQeEjnj2R02/VCdTc/9OVJDCYFvWRg6idJ+6UPup/xFF6
nZgG+Vdhn6eONJLnU/CdrgDcTzkU9YVQ40WOKTSKlpDh1qKvhnDPHzvlMYzo8Ba8EV2fa/VzeYNC
O6RsxP0sNc+9kWFQfnGyPkGF9x8LwbbtLzXjcM6gWdjkejuG0uMACMijPUzrs6FRquuDVB2nRi3u
UhkRhK13rSJfvnCYyyp0nn9hBwkdnGQssxKSL0x+pAjrAo4aDt/quJHzL86WKOA0J6c/B9tdsG4D
+PN4lyQqIs9tZLqBdWTs4Tk0LGc+4R7e+pUJLYAw4epyE/kWfawkYTzr7svDrqYXO5IpT8joDbXO
n8OhXQkKsX0CO9c4RTJn/+5DQqVitOjKfY+LaZncmYZ5buRFFVOTl6GPLI/Qb8vWLbJk/chr7QpA
TJqfWBVC5arycFmiivgGOWsvrwYwzrr3kNr80dDpYGj1GDFMDvWfgs0jYtA636MJEbUk0DP4pfGY
Lz4CvIHAy8jaSlWay46qWhX7cn/8NQzwuLLKkD4HfK7iIns2VKk9wFw1+RvpwAPRvx5GjjQHENuM
JN1eGPgLobF3xM/ZdzPa0hXNQ/eg+IjZfm6iUpBkElpB1h+nc/dFej1+2qQPBt2UbMBu5fBcD7g+
ERsoyJe43SWgWZnzYLU7FxDHxlbqwt8SIXK8Nlofi1jhHXTlBe4AnvcyXDEb+WupvKVI0Se0hAa/
nTOxQ39+3j/+kQL4wvMQLnf12ZKpaPLV6p/zk42UZiGBd3W5u/b1u8CIqS+BdXVOGGNHDFwwjrFe
IQ2K9sKni5NI06kO8AHNXHhGt465EYSZDcrKra2tjjyypV/BhxCJtSb7l0t6tTKsIkTdMrcM1+2k
+QIMss79whrswUv5iOvBIvRdw8FzAO8TX0UsLDs0wBxcyUbW0y/it06GIgdxebXYCy/o1uNYUyCi
Bs9twsVWQYW/XF+yfuFq9r/dtINFC+RhbNCXYEOQ7CUkNaph2h2gJLLVBf/rlVl44Y9ph4xcMcBV
zJfE5/LDnq7FK+6nafq01ctD5VIDk5f0rMsm7IBzvKVZqZhuV2EvWFL19k/GrgywBzOJCgTFQzc5
8JuvUK6dVdvhhFIElttFOS2CGn6z5DqbvtpkBZYhPfy/MTW1sK8d7GBs7TTdJN/XrDmkm1V5V156
u0kIoHH82qcfOTcLcdn35wqYLW/xqfy+NlRmcurpnuFL4l/rhSc+MAx+Pdj4kHrieYLjTNky0QsJ
TrXUggVU4YW0X6vxTGcWsZEPGrZiFnrf2aomDQ542h2X3iWYCGyaG/0CDRQIiNCAsOayKlCm+msH
RQWHYDkTasv+GyUpHzIO8rEabf1th9y9SvjdaWAMujJikqjKhUkVagy/TzQLxMv8e9sbNookLEDC
UOHLNmP28d27oFL+8HUWmdUSNYfhQhA5nvZzaQk02HGWUwtzj1G6T3wQ6+iX117FKe/hWKffMtWw
uDXC7mt/J4pNbydB0i+GrVYMJLICp9kk5J7NgNRbvALfyFDfRS4k8WpZ5MBlLBJs0rN+mU6qcXd7
Ma1KqmzALY0/imxxd7iqfKnwImVVHFJAJ6KuAXr2KHisRxi9n7eWsdrmDXYZBD1/txIaifrybQND
0u40ZgGSmKbSmvVDpijkf0BQjmPDeWxdnWwScGGwGf51/yDRPTHV3b5GJl+iCicxHCwkNzWU8rz9
KTZHF84xkgCQPRxMzZU4aYWFBntZ9Sg17WL4kRKlgGbyghDQN0ImGfN5FoOZGjW7uYyqwuOvyY6V
Idj6AuooPZsn//2XcigE7yN3f/eFfFg955v6WzuwOJFViiQDC0e2j8WqBk4oY4cuqctFvoEI7TKe
z96n68uT24/fbx7+g84qhmV9rIZWZZtB7Uata7AtMd0uYmBRFBfHTlXxzyRTdTj0cWTkRcjMPHTs
qi6ZNtQZg1jzVVuYob5q9kWF8sHfBThHI0m4pmS2JLLKOeU2ApF4LXj8zmR7zjlB6LdA05qhy6rQ
NRaCBOK0abM61kI2VscmCsQgvvBGqD772iTBVECWeoPsty0Xq7IpSjAbIXyZsNG3alPu/04U51aQ
peix5xx3YJSxOGFEsrpdaMhWQ2A6zH88Yqc0hwQZBaFEuhiArpdIa0XvZ973csdE8aJE8TojO/ng
y0q15s/9gGw81XBuHPsOuZR5+gbrEvvnZul28WxkjM7Cc/xh2j4Bx76IPCux31b96rXwNMxqohG8
GqK7zeOHYHbuJsBmrv8iL81cnqfvl6VjAEvGvwlRepEEsWZBN8zLE4Hy+Hsa1LREyxLrPnbbZ8AC
knn/9C9PHMGe1m1lk27qo3hbZ741eYHZz/K+yX6dyGhiEqaYLlhTS3lMGU1t7qYB0TZZql4GFIJH
qEsGv5eAjU3E7zpzQbdadXKVNpuQ7VvsONyDf2MSZb4ecNAWy0zmJGmj5za2VH6GU6Nhvf0jH9lp
bToynZ6TSZN26rCuazhqcVKhR9TDVA2K9Uo6xKVINaqKcjC7bqYMFl3XoYGCCm3mpplmqTHx9jOS
7HmU/gptUUemE2YxsryBauNcxynfurfawbq7iUL9N88Gv+EmZEdSJWLlSW8eM/0rPiSnA72hDKNj
ANagwPwtApOe+wALmz77q/33HamvOaCtjfm0HRVUfx5rGsIu1jgOjUJ9daAoHvZn5gXK8OLnP17v
M8DpejnJuNO/fH5aCDQscYrA+466luwrrR4/V3p59Clia7MjI2DCdn0ZJdrKsO924LkCW2UgafWI
/AcfoSXH0GTM/5plhozRbZGpQjBhy2q3I80xkTKEDAXJSRXHNaygHELIwdhBP2IGlt7GwwfGQqy6
sIYdFoQqmmt5hyGROP1dqR9A1/2zxrNuJC8w97xHBuY9hNkOiCS1mAOahmD8P8KNqsqwkzohtbwQ
LUqg0CmQ+YC/12YAq0rscxRQX/nlMHtXqdYh6h2VjAxnvgeKZaC5f153cU/ikXDlXmTaMClPFmvg
Eynyb+dqtZzey8jqYQIX5azkC2LwR5NZkTdRj/o24ceONOjKXOso4fRYgTx20px27JErXpBKiweY
qXESqAVnB7CckisIh72BWABvV0aYkvZvsE5RITY3l258vi4S63Q0N+Pw/WRZC57PkNsGj53K1TH4
zyGjIvjAx2gQqRaN2YZIscABml+NVUYxqvSztNq3GEGKisSlufO/7TRHz7s5hVjCmupH0ubWNT0+
aUpQEMf+CepC8omDNE7Zza8NiA7rKrFEmGwmB6EtV2t5tcTzQXpU1YKXEU/s7NuHP9DODnC/nb7T
pwadafjtpGu8pdj8WiVj0/Od8oXDjPH8SvzSP8jb+Sa0cLGwxWYrIgxOo54D7HC0SlPWX3gLX+Gv
99EMqxdVFR8wJG6IteDPDTtkds6WwWwTX7osTYmYmCBTGfiDQuS1pKAMWmYTB4aaZoecuj7rwfh6
RjLsJlo1xqbpvIl8yYkS3BZ+l1uTbXFSwY6IP8OOtth4tLZoggJ8FJ+f53r9QpErXqDJUJqEEFKx
34gRN12ux9ds7OkfyS8rGmlE68ax+p/m+X4iBtty/WX4mk5c2OxTg6vP6YpVafVZBZfV6Ko+ALj+
ieklg9K8pB9CPtoQyW/K/f6SPE5L3iBdRssAP6tlKDdD2MzcLUsg9XZiNNjFpYrqcpC3y+mUpx25
YNoqCrtu4Jfcs6X5/27Q983wLjpwR9XD8tZGqh5eCJ4UusPxfBn7ce0OutFdabmOzDTCDz0Av05G
vsZDMXhOgjZBBjTvxiYea42rNRZf26dR29zEK27YCjI52PoyhRO7MvEZlAAIEGY839I+tX2BpaWy
Roof3KtrV0lVWBCo1yJkBTlppfIpIFUAXHWmkL88Ksv6dfvJICTQl3w/OZMXdjMSUIv1npaKStUK
HAwFST8rvsISeIRl8k9t3LTQoZjarfFECRCPvHPXl+0j1WRxTTJUKl+5E7ag0ZWfVfINsIAlZtWl
O6cioQQD7cZnYyXT7lUHmAEfw97RY7KMndhqXD7OG5pVpr9EXZgem5owFOfmpwFL57hgRayjzP+/
3AUBXrcfhv9Ggm/rHHzYq7kIo9IRiCyCk8I66Lqo00u1VImuqfodxSfo8yVh8qspPT2nHme1xbOI
5QIraSg4sZBEpGlaEBw7vj4d7ASX+I5ZrVPP7yS2okUdoGChWF5NQyXiT6mqeX3RmCYqMByU0UyS
QRy6VbLrrvNjaL8sFhzRsCBpypOsT7EtjCVM+/OiUX6BZHUfTydicWSflJ5BHn7eGG5XeDfNMefS
Mj9Wp52bZYQVdm3i3GCEMMRsNL5KH5ZsO17rjkMthl3O75o7+Tikd/W/gzI+Dnawthypv+uJCzl4
zVx5tQ1ElF5L6dEiTCNtIvJ0ame1yN2tk3QSeocgf2KFf1HzYk4KiClHM9v7/mJrVQhAUekhIrKE
cwj12yQ8+k92Pgksdjpe6irxdiDuPsPMnM/fks1KwQ5pN4i8hMZF/LH8KmXSxWP55padHlGzK/pB
p/efXWbFrZ24+vMTRgoWwQ72dA/oC9hWWo/+W3mfDe7nLgvMzR3py+kEHnD6IFeIZP5BEjKBFgpn
KJf/EUh+oy5MfY8euI5tnuIttbjScKqRDt2FZwTEyIv0vYf9x8sc4paD9SRivwbfxD5NSyMO0zPm
HaXF+Lh2bV2GTrJmPZhJC2taEJkgnAOIRGYTvQrYDua8ctug8krUGkNQnrfalk4iZZOiv2OT14vs
8SnrTfyHc6C87k+jsB3IvcS26oUBgDc+JiGl94ISi34dzaEBn07cTWc6wo0s4j15UOLkNMMGOQ+m
ZbQI45scooQWruhwY6N7JW4lrXJkytUJaS5vQIrM/HwbKD7zi+QlyJyeU3z2UWkUEFlRfzUJFoRJ
uTIWn09BCCSPWow+MxDpRj/lo49Bt9+GnC3uERjVOvb7hqhitQkCu69j0k9yV3OGVERwlAAV2DWn
PlJGwJXPQiBYdaBF4QRot1AMas335dnTshVLtsxV9wsFwVtLFhgZn78F6hCXzk8+2f40GLdUrErq
aTUpHBh58XKRIhJdH4EiJ3JRzhMQcu91myM3Utm0RLaOZ2ufEyteCorAHFfuwr30qnPgtRbmk5hF
LpxNXt7NzKe07vxKlwDEkX1dvE0cy87VzILzJeFm3KOzf7dckumTnJVFFOtnNCBq9cmHjSvKPFbP
TmclmROYcKcy/bD+BhZ4RklFqYB7IZ6VF8X+0iJew5xZD3Rtj+YJvNhVJMo22hqFRxJGM/tL19gy
7QBmvJel8oFR9NxmWzpU5pi4ChkLIivtTKrAoJyI7mgLvii13wmpgxVbuYrWH2f5ylHyXNhcHSxQ
b+ED2whzudOb3nJmoX4IiqJEmV7xJKE3enZ8ogrc+byQiQONLXNsBDsLn8XSjeufjVyOrx6O17ZC
jECN8cRqyxAmijmc3ScSZUKRE8E4CU3Iyga6532+TZ5IP5bqmKqYMfLxKry9NOv0PAMmLdXtu1In
nUBstxt655bCygFxT8QbOQNn9a026A7tDjBx8KQFs0I//bN4ez+w52lafU5lpL9jyNJLmPLSVn53
JGq/fMK4bhnOcR6c7ule95E9xueBtxcrnHMLqW4Qj/Ipvo6nipiMywoT0wodtCL86TQ7i/VIm8og
zfRUyctdhpi/bMNngkm1YPZCCT55zL6mCZZ/h7lLJb8gwy7ybYt1pakR9SdDIH6qoZEan6Nl3mcB
Ki3dD0AWJG3ruP2vWdvukVdCe8Dvawu3kpnmBkL0IAfjyYNbm/EpGOUvagBgCEMSrsxjgsIGopm0
lFiLtNElWDRObGbBpWvapkV2wFyX1mFkw09qEVkfHmioy7GLm3rJ1lOjSFGb+/HM/CRAzKHQru6K
i2dqc5DbD7HP3AktjwsGX43APK0oq8zpT5QoAk3ENDX7VfPgUCL0j4IwRb91g3MXs6EhOpyzmrjB
SVH9aBYsYvi3I2GdFdiTgX9TPnlgttzYr4OAZV0ed6wNyH3LMG6Ng9bSIACvJ7D176Cm+rdO11Ks
krcEFvrAqzJNz1bU6RIqfY80Ox1W+bLexzVMk4pXbX9Y06ADtpctk4fk7QVa+gZNW1ac44kt+4vB
6gZFuMzVn5zkLamVvfP4ZdkK0rXqedUSy0lukHzA/1qaWBtxxkVt/ZZqHQuMUwWsDFeAJPisndgJ
IzNYUqAp39RdVCDxdFR8wCx6uTv+5G33V2Rv39LabpbVLM+lOvw2XUUgPYjzlcFvnsNpH7PMqv/q
lXj4TFeO43hn1Cbf71yqdWBTCiGzamLsSko2bPrjbCvv+AQF7+1UCjeAuvgocRj9QxIC9ZFbEaDV
N7SS2AacWWtkz81aJ3kGqTNFNy4EMl5tqpLpRoNA+qABinDXqlbDYyjkmdC6Rqg33jN6P90dCtso
odbmYdfuFpBSTn2n+47lGrm/XLK+88BYT5g+98bjvbCGPFirpnh6FN3QeC7OKtDGVfC2+ht6YV80
dlsx7/fovSWkAjVCODRMtVbqlsbc9LSI/j7xH/om7pZ8S4gMpkB4LFGooU0c2gvTLu9hnAm3kb1l
xSucRFClek3AvxM756r4euQE4GYArFe77t5JcB/tdx6gMU/CDiRSjpOmXyJa5hfdo3H6jsiN7qkQ
s5rtySODaBllVZv5z3++9q9bz2IlGA5MJ/EWSBFzi6qfuvrScHKbRpCNIY3Qhba2LLAqsaRfMe9O
Yx9JMkSMsiQQ6kf9yLHkucloOjCmAMnxIJ7Da8ZOZMwlA7h7nRcD20s7n9hY/usfthTKQAdcPzN7
MroWwSWRyZtS+NLHJtD8rz/iqY8pu6n7Qb+CTirvPDudc0dLV9xpBy6Fz3eAXzEfUk9jW2fv/UaX
b/+VvRKKcvpcN6JThVhU5+i1QczXQ8C0gMgKp4lgMxYRbIPrbmxLADqa0A+zzUVrf+pVJQERd3gS
yx5hy9CiXqaKnFvg1KT3V0+kznjnqpAiDGBxOFwzqt5IGgtYfa2dnnLgranBvO7wiyJFohYlO7pp
xTXGfvja5HiRnCgi0WJ33HLgbI7BCO96n+GwPULR1SGI5WIRgpoJTV8ZyuMVJIwbRhR6QJWO/N0Z
Xv+b77Fagb3Ph4Jq34ID+2Iwg1nCQlp5EFV1FYfGhli+Ew5d1/zP/uafnUVJujoqvZL7y0yZfavw
KlWGQaCvEfMtl6X8soy6K0Qo1v+/DbiGpk8wcntIE3MKuTSUljhVSGSN41pEFvozFV2EPYvoWsMh
ghesnufUVTJ2YSkkVksoa8tZxQnY+Q3uCdGOdCktb2GfMRYIE2yCA75Re7CaDhkZgQIVg/PBiYad
9mrliq2+RPtVcImp0HkXaNzmOLcms3y9JZ1dCrjqa45UcKrTt9PEChsmst2W10XdZ3SoZKg+Vpeo
YdyC4aGUxxGRbJymMXg1zJzxZcC9ti6qjD+4YYHzCrbgMSZj0rAP/z4ecG5GV28cQjZO6OQ3MbW8
pnwtsFfBMmPA+O61N+9ALd8y7y1j1dD7kLQAWdAxtO9tN3Beob5X3fq7eEcI+RdNTMgoFr4t8QBw
CRzfn9B1xA5Q3sQv4QkDOFfiONHh2G4ZvOR8LXhIvtU/325iiEtch/RlSXLY2578GrZkepSDGavb
oOIbpliGMcdwqqYGnKwLlUR5RKfBOcKSq0TlRxs97b8WwSV+IarmE1MoS5ImMbykcjDzD17P0s3P
UFji9E7wfHJ2vKcCig6c9vLGHMkvDSbHXFYc/R0PSIjvONCrqGlYTmBCGgj5DK4268cMR+JL//Uz
MfWyP6SW8GUoidSLeExzdqWOXUViOrWn0pY/c4NbLoPgzNcivWrmdKJr3Z25Z1JCefo6j7rhyM2g
NwGFZomZeUn6wpTlB14xNz1xX4iwf9EOzxpFkdyGxHSnPb6hodb4Pd7f2RxStJjUtJkMHCaLFKv6
vlAvfffeWqIuPgSpkekQfiILnkVwbBTujtKccEwpK6POr5MogDMbLUYSNieme7SFI1SiWdndGv20
QqOuSOexI083V/e9TmuO+Lsl5zK8CPU0o0tS9AjtjCY0vHSJjjl/bckDgkfY1+NqkB44Fu1AVGlh
YheVhIOW+mxFlqBCw6M7sU0vcIq7uXyLb2j99TcPzgqkcLKmcvV5EkD0V/ghcUo4I4urATKKog1a
Lwfxws1adurlhV8H3r0aU8S4QWkcjqKup4/zdPMwZnvx55A99fXZ2KbdeVkmTk6L0y83nG24bs1X
L4nh+3weMZMwpnR7eVx7omFVjP5SzaSuy0NfH19CavlfwV9YMBFz1YfuowF5fxsrt7e6UdLiyO1V
w5iW6BMKNLsgEptqsOUORbxF12aAochzBuHtKp3gShLKDZhMZz1L2iCMkuQSD3abm9kY5jXQZBCE
UxxoNG5R/kak3o6p9dq1EtOOfbuLejyxudW7qfPuSCh3mEgegR95KVTS6R5wqOEWbTxgzpb+Ra10
XAQzqrsNu0Oi1qO//fuoJGjvgHfFjo24Qn0YvMWD8/68Yy1BvbgnMV0Y9S+ub61gMWZ7EEG0QDji
2ociog/P30QsYJsI47gKkQ4+x6jCO7fv6EnfrJsIQF2les61iTESVYRJMhLbytvuH+6UGKNakidF
EsuPqBFinMseNEbRzWJarAOfS7689ze4M6R3VJTUW0/T7SfK36eDOf4vYzk5xX2DbS1M/LLsxj61
10u68NSQJswJjsZEQr7SK+3LbHhUCcyfxdpAinVbAF/IBdAZ2BEah2EFaSOXBSrxGnB+ImQZMP6V
RQRVNzw4kpuWLtv+gjMyYYKgsx66PibIV1UmLPJT0MhhBoP4fmxSjIzdVTIyXQ3RHWOxOEyFN2jf
Q99dRJiabayKW4XIxYrJ2OBerAjEYx2KIvjZgMtd159+GAvc5y0MZSRS9v0zogbznmYsTfNOwW6s
vA9kBvVu+C9mB4Ppfw+Ik5yGfOTNuWz7xKK8TwUrkRyRJk8wpUS6j5lpu6IhMlKh2VpO2mFmjZ6Z
81dkoySBfbGwB22U9rUIfuiaZOLNXM9QTE+Ml2zZojzUIfceuONpk7yTgalQ5u14Tz6SiTIhrQ2Q
LkKourjguUg96nraT7dUQCD/pcBRyN2TEwuayXvSRfgJJSy2hAEIY5IjQXoiyb9svbWgQpx9IKgC
yq3jscqNfRJAjbxlE4lIvGVOTHVFFlTIx//LR+ZxH26dM9HMuqzpqcZyOgyS4TptWnFg6pe0huu9
rw475zlutih4MyuiGUVrqA6SaPxiuXLBtimbBiih/4WpnvjpD7dsmaxDd3tQX73UnjwF3b+Pzyhq
A/2hdQ7ianCoxr13zPhJ3ZBs9J9f3UqFcl15hGEI4SqVHvPm6wzf1Wru5gu/O+qFvjw2bxPCKjpB
EUPsdy57DGe0LvgdWGFrsmICh574CUYGZcbN0A2jI6et3NqR/o2V4Koln6D42rxeHqcUPTurpc7P
UU76A+uJD+xXs00q0UnacKdTMPoOD7HdPsqbElPU/nJ7G0BkGISy9h//+mVWbV+dywXG6i0ZZCO0
QObS3ESQ0CwACa/W5vMb1ind2k3osYLOAdKF2RCNdrYaqsXj27mA1GAZNQxiZG40qASpva2TIpyh
qO9CjVqYRvMHhtx+tkDU4ttOVs6+w8PSprRHhE4PehkmktIqOIVgZiEFj6ba1H4RLfd9EAmlIyPx
NC1YvNCedWBRvERNbTYLDMfjqwW7QozEP2WeSSweJhH5WtWpdcECDqS/PXPrstehLukHQFi9Mi47
QQMq9oGNXPXcufWE/kZ806wbCulveJK24FK/BTf/Qq/3P9yh24ERZuOI+KGoDILIkTI8R0DtkSsK
qcS7+eZAKeS5Z5KYrYIZ3T4DpCKtBZdUpBph+BgDt0bbQIewY3JzaKkbsHycbuEmDLCDHRG0CH2R
Ln3SrV2SUFimG4Z/3Unrf35eCAMg+6BF/m+KdxlNp0RNvY3xIbiZXFX45MEp8y1Pl/MqC8a7WPDv
tgG3bK+Lhd1UVly9EUEhUgKzJYIDpBAXs7loY6zsUw9C0/r4WUjwOfCq+Va7v6kDT9k18dkG1h2a
xa+8DOMr4QqvmtoET1gkHfA8v/16iIewnSw7HOmK+fDuL0bJt7RNv+uG/U2FpfUe/G/KrjkGja4C
sF1J2ydpa0ZrtbSw8qNZMoZwHD5exssG0FjV9XM+No/+A74jNZK3Q6N49ejoAKHUnWMUdAt5bNT3
IBgMZ6H6uxFB9SLNR+/AYOyUpRZivW19PZFhMul+QeQYrNnM9CjesrbpcKdeHpR/e7kfCGXjj7r4
qA8kUeM2ObVhwqnxNQkDNcKKIdYZwMttlPnz1LwYmNu0El1UpgMK8svxn03ASYaISftTwe7WM9Sa
XlEZjWc2kCJBnm8htq/HBgDZN2wKaIstPhw53KuojMoQ1I1/QRH8gCe0HPmjeyC6DjGH6NK3rgI6
zuawqnEK68i2XCFC+6NlSuMHPKzQQrc39dBYEQFePR9nItiEbWWV7afqChubnWchTmeZErFi6zZ1
xpV4OMhdj76bWdYUb3AuCq7lf7OFPEKxJkfkisGLLCx8RVbjBLxqCY2yduSbS/qzctqFIvqbqgaf
gciu/D6Xzs1tMn1IKDp6AqEJvNSyrMCRyosnpJJtZkXH/l6/n93CTqLu52mshIUNpug53080qC9n
rSw/ZiThOjFmOS5IIqejFN8yUrQwLDcBL5umPm8mUUwMRocmjxQC2CHeCddlATAP8q1lJ86ROguK
YSbhC9epUvE0XnYewe0Gl86hxUJTc7/2CFEeNp2kvRwOdq5HUPATNlJj4nY9oly5UO9A6xhknkCn
3EGD0yTHVjONG955SWmTzknJDHhQCtipGOA14koQNUAfW7qHpc8T/SvytpWYKttyW1OmuK+wMDRm
baBuR0vfnVDreRFOJKgg1ANnYg6xX25Y1q+nMukSaZrYTDKP4WeolJnBCtDZwoId2uMWGwd3V3+9
+waFFiQqiCYG/Q5nMgEMr5TGq8OpEMVWaGUewIO7Uzs9qHsxlUD/WBJSVny4HpnrcIyPhT9wC4EM
8xhf7i1lAzyRsEa9bFQCrJ3mbPF42RogQIT6KLMWqkbGzkMu3YHn/ZEAIZ9QrRuiuNvfxEg9SsxJ
CykzW6pLGs6xXTHdE4hBWgR9Lu9LxDpSRL0gzzlWwoTXllHxGAicbJPaa1k1Ka8qmxZVInFtfJfo
9dZnvsaFQGWpWlnXwhEmWf5CtEnIhVz2rQZdqmSdwf2F4GqNfJxxTS4RsUTNcAMspGRMyOHXdcwd
1R5cRS/HQKcQK7dYZ24rDasU++dGf1kcnfKQOGZ64VUPqTez/bzIZJbLG/V2cEX+CJ5k/X4Z4GXT
z5gdAzE6/rklbQvYzCylC+8mwfiUs4dvN7WteQOsDQesEevrzCH36oun8O1LapKSTYTBUH29uErQ
p6usJ8WD1MQXk8UAknZzGYdB3D++r1rUfwUOqV7XGQE9hJyV3ngVfUVOxJPmFA+cI2E1n+HPqVqu
4nkuOwLh8Oc2x82QF0ny11gIA7nS5DO80g8CpfzmSwG/3oBnMyBk8yO9aRpaYsfCshI0iEiswuy2
wEwvYy6N79SiAv5HWLU2Ikq1ARaQ86lyqBTiZGPRZ0DQny+yCOpQWZjnijxefB7rpu0fvFzntKAt
3LlEzPwPKCgAbRlA+fq5Vo6sSE4eU1AfIknXfxxAD4WBRo8EqO4UdXljRbovWGA1Z93V+M/H1x1K
Tlg0J9m84Mo0LoHBl/DOW1xc29GnKOONhYtX4zg6xKfKeZS/XHaAAUwQPhDq9LPzNRlSSGX1G4cC
/Mg8RsDU8jUenChPmNQoesXtx/FeABOXY8DUajMyZDl+BtBe01Dy3MZd1GShhE8ULKB30lw0ZSAa
T18oTkH9HBf4lLAxVEXgEfZT6UknLQgrngNyVD2NpwXoD93QvlvNtz/53S3CpySsqHwMVWA3kFSv
rJ4sLigBGX81/8989kcDiWBWFoxqQOvD04fR1fkWVmVorrti2Mp9eytGY8SvDOl5V8BRra981WRc
czOM1oyBVVOF+DiL370elUYGzTWmKBF7ckYuiedaPg2MCF11WrxuC0ZptIPeMcXDua4sueq/CrQp
YDVZ/pRukCenXQxxB1/MmnRl2TN1TCgAT/KdQ87KS6cXggwJ/QqEg66DjW+XGaYVVZBeQ/nlITLR
bR8u9nVEgzx+1NcqF9GY37R6SfcqUYvcNS+svcP+fPtTXJXOPzx/e8tlXFxlGWzmRdLMjT5PMPrp
NY5jE+4gNxPijKajpYo5+sUyTihxIP0YtUmoh4SQkl7A5v1ocOy5ZdWri+gx+dNXKyb6rOU2+rcC
J2kdtxyaj7ALpNoND1Vm9EGdvSF/Dw6oAy74T+wjV9GjaaCnv8IcECHAErQDvfYJ/Yes5sEmyjr1
dN/+x9zGLSiBoVourV2osGpA9hnC47g1eLA4GrBfSryhxsFwtwcEr4lZNIngYgF7VVTSrqjqDxeQ
N7Qi3L+kNA3MBpHfcr87KEtppSmlqC9/12gpTzt6CJK1hKiVYMENkLbMxptSH2gOFWSB2FXIxmPN
QcPg4fhiQKf1p7Ms66f0yfUdCphgee62ffMaeA6bGYnt1m3e8EA18UBp5wK47V16194tJe4c1ajA
l5Ivv8g8FMFWNIaxC3tOsHvidJ9+WHZ9tzCn1PJ8cBDDPxuQ2lLQdPmWm7MVN9dko7QqiVCYoPUr
jvuWghIHzGpORorYc+xfNCl0A7Ciqh+fmRrA0wSlaD9aHPOsJvXTinV+wJDeZLNu/NN7H40IdOOe
yNVxNXZVpXR0dCnORQkGXB/cY+PHIDJsW76ms0jGvPrH6+dcUJPwQK+YshmMD1DMdCXhbScyeZ+3
2bRDV/n1brq+twTPy+YDh2Gl9CvdUvH4L4Jtq6VzDwyYfdRFPOz10yRlfAidKqGxpsuEZi9aUyXb
66GZ1L20WH5uKy7QXrBhnjH/UYAR2gJu6kQ+PVNlCCxubv6Iy7y5byCT6XyOemZ9eFrdirKmK3ax
C70GZZXaDNEmGloe1K2sHun4RA/ivz1eC7a8+gRD3Djjpbk8efGB+/Wu6AwTizfR6v0VphayO8So
8zxpyVJ1Eluz/3aWr5BBboar+cOaAbOlkdATnvt0D4KFoda44IN5IVRulSbX+uwsQwNliRlJ+hcN
Axh1M2uZXZRIgZyCakRzGk0Pb+3w1PkAA4ArzGQMtX3nEr9rDO7t/zRLEebJ0oO5HC0Qc2YXt8Wr
6Uz+sOcl2+onuO1yRCbDk5r9zCVObJdg/6cx8eJxLffvlCrNJCIDJisN5KV1Yck86mdCAd4MCPSW
DcsCCuDPTKwzrdBGXSzLuG5syAV4WVW7Y+bwU7LlSDnr6w2Ahxf/i44017n81psdgzlkiURIZ+rW
jhJRAqFOyDPhGIHVYqRqFgc8DmedqphaXbpse+Vn1GOgBKc8AkqeNjEkNz4ZtJb5QN+CRs+jLDAR
PGSuOEff3Q4S6MAPMOIgW99+KyWzDR/OZSapbkgktJvqJZtu0AEZDznV9dNZFGNGlbe+6EF7/EB4
QA5wS/NJJxfIdAA8MOoCPq54rxoT5zOKE1ssbWXnKVfnGCArRnQS8WMfT4KT+49Ccuv7KypfMKlk
GdmXkvnVWnXwIvkKfjLhXUsVbV+Jr1RNoBJggDvU4L/uNKBJse2l1gwhYdtBlUurXanaDZIIGL20
6VwEtCJElhPd42+ho4iMfmtw6GrTni90D7lpACMw/5qsDwTPyjjA7qpTTv9al6MtWETScLblOG+B
wuxhCQvFzU5yV7Ri0Hc9SrrCFYIlddurAHEHgwx/g0WLfdhp1zYII+9yuB6PZgPsBnIfORfOrT59
tQw16x+90KfNfoT83le76ZRbH0y3uAD9VeefzbPG213HUEkA8SgWmdZhKh6cnC58g4rmJXIbklzm
D4hYaUTLT9ZKGsCb2ToB6t85wYjyaODRJ4TvwzsDYbcfkwpLcZCsV4qEW4TDllHSv4+Tlz0AWJnH
irnU15Qv4BzqIX1ZHN2gKl4oWz2jZkdB2kvpTL8YRfTvNbpJoWs5y9nrgNfuioEwjlP2SBceXRMA
hv415/TMY5MNvTUQ3OuXICchXswATUWYBFio6qd+1EIRZZ6xXocgQK/Pu77K+g4My36JkgsO41qW
21sAPgPoFA9nazv2ReHRj+snb3J3LIEK/XPI1ehSpccWqSCyRe9bOKb6TOi/+CgFDlll1Tm7Xb6f
AMZBx3h9D9LvrNMaBoCfYfZHIcx2j/sMJqCP3X2IWLrUQDvppLZ9BYLlFhONSunbpK2Mjcuf8Rxd
f0iS3pX66/X7wFFWAI8XpNTWIm+/e/jocr4y9wNTr8aKASdpbgx+WbBatplzj/fe7fv7KnazpQHA
bXGzFaXChNU6/4CBJoo3rn7zvEn81ZS9X02AtWvaqiZ34JxwY/Sv1gBd2ndHQrFv/KNqBoV0FNNR
PIlq48xwVmub4+F1TMY6S6BfKzzjSVGIfMW4cGQHVNoDazrcWK8Nvy9I/wLtTkumctTUj+yocJr8
8n2dzWs4GzDIB6ZVzKl8oMxlME32V+zkGhs3eJfd34asaAtQAEiF1+e1HNuP+b+VCMZ0L15pGnMT
5IelyaQxiFfgsG6le8dSQ7AYR4iCJOIJqLp8aSM+CByfoNvLI8f8IGmB26uJs0Vg+WRfWTzvV0fq
ghYbPBus+DJZE76vijuwPKveZOJ552/4NzhdFI2NZLw4oa3GkTVjcYqw8fxcALMJnNGNUdwX2skq
rcR1+9m5+6CjojSmfNv+0IhMjGY0jUe6E43zeaEi/4d2nN98KyREoca0MlmOsxe2htohG1ubwFuP
/TuRbOsQscJTj8bybLR90kwuFAsSGnRQPE2PJArMUFF+zogkXlAPoeOez9WHc+Xe1nDgTOf/hz5w
vC7Kf8OEmsb8rraRHWhmNIZzE/YMWQ6s/5qOcpOu+UlXVuBc3YMmZu21QraLTmufxullBNz3o9lA
NTmh6QOxOQXYnKrkvolI1JXFd1ca4rJpQl9kXOTrMkj6H8WARgV3pj9tc+yEj4koYJVx7HN5pkrV
xyAwbHqSK+hFHLA6B015NZddnA1gYdoTVXAJJ0sw9yv1EGHcaLv43NzAjo87r3+w8RKd6NMWSHBf
Chbay/mw/TaFkYcMGIdEqtJO0E/wDqTA1iVkfJIb7sujGQSh6uuBntn+F1e4nDw4PJqix9LFxE2C
5btpPJXLqqEmd2bZffdtSLd2fwL8KVkW4fp0K7qN3dWM2r0RWSku+dudwa0uhxvCu6PPQZuF8LYy
H4wPgAChzMUyWdwCr/7Czfq+jnzgTpPjXXIb3LfodSTXHfuach0y8KbTUc6NauU6pj+wDKxRvMOM
MU8qDrWvjnPVQrIQSShzL1Q0x/xMfd2Ar3N3P9HBOZ/19czHY9k8hrIM6+u/FnB9BCywtACxuKA2
JeDArYkOHwokmbfjKc1XI61dy+UmZ08zdaEthWhAyHykfaSKgLDJh9qJFtr8bB0mxQPiq6z9G9N8
nqVhinAjxZPNa8P4hXX/ljJpL/NIMDmrRjd9sNPe0QXymAXrPsSnoF/XlSGJGeNlSVTT3ugNmf33
tEy0LYUBTwu/L8/v4V1eBXu60gtRtYCc+n7qoxPxESrvr2muXX4Wu/H2HV6UfL8cTBLmmC0YueEQ
BR7VzjE6chipK5pE3YvTXPTUZ00onmRrd2ccgseXRlxPJjSnsWWcHqDEDT8IL4JtEH/YTpNMHfxT
2V6QxwD7yy2TE8qS6VHTARKPv2lcqLh6XaGhHLPtX9WZT5R2hqUfb/Silysb3n4FKh7LR/Sdd4UJ
FDfzBBZKZ3TtiDPocDlOs8MCPcb1GEAmy6zbbTziBscSwR3TlC0Z+QUe/qognufArPxJWOWChBVs
qFq+rQqI7LVISjKcSuETYz9jKuiyiOxAagfGV35cRwmBU/RhBuqg30PtPjCGb8FcsPCxdOIG0knY
goE3hEX3riN/LhuFccEq5V1qI1JCNbtq06zwpLFiH2vTGbJkaFraPQNe7Q5eq9AcSZl3+hJCSZmu
mvpao8b6x1m7jb+mhMSmgBfg6u1PgQoNXJ3fsfh+KA9SRd5fZvIv4mt9iYW/I3Sxizb//7P4FISx
id2lsp6fCQ7WjURZnIhRiQi18hVYpKLVfJBRGOtA3Q7xJOOi6g1zhWV/UUbt56rsUp47Nc+GAZ+y
XVALBOvrDtn7+wuHjX4zA9wJMU6AgffyPNvFFUER8VB9SUmuaLSXqyTV97NhQ05PirVE7LhY2oJz
GwsLXQR8bPnVjSBWJyX673j+ODk1rFPptyH8rD1mtVL3EOBreqHflzEWpgSlYjFsMPnV2fdpHDc2
VjyvudZ+8GFWkKF1pICvI9/B14KASKweQJQmdTvzzSUS4k48U9bkHHkYAxAW34594QeokxyRPVV+
nFYfBaWGrDQ7LXeiN869ZXfaKam1zY1jREIsLSmQx7DgJ2c3D2ov3pKmDNWyuGWi7pfX+y4eCRv+
kCUsfWgg0m0+wGsaFZsTi8Ski1feTWoOBYOK/e5+EtFNNuwvvhxY1kW1zpDzSt8X52kMolG5k4yq
dZPrtO9fkoW1lZFSntVrxs0X+AxahQPMK5rh2COlUgdkc7b1HPWTEPHMozJlXyzP2yoxaAh5HcRA
95ihKBhMV2wqxXJLBm2e7/gteMdWK3WXQcKJs1JTNIPQI+yk2R0vUKdbKreCRPoyrobt8q1XUX1z
T1c8jfUXjsG0HNvw7/2ArW1KFun/mzrGiuR/fnCRtJioS/bT8JYvaLchKUD7j9nLXVnuq89FAXcZ
AGhCK1Qmwh1DDii5L03hYXuvfiZDaLtTFTqxWH9Ioj4hllIZjH6Qjb0Joi7/4MKPD3kkNSxujD6F
3CbH4EzZwi/K27oN/LllC9oW6F+TDQ/M15rkd6r8+mEhvTlwG67jW5v0vY/ZHPCB2DEhy67AgTWT
VQp5evg7Nu21DztPkyRnZvxtgfz69lszjUeHNK+PN5N3kHf+SaRjtQXpTikuJcnGgzKoBOjqdVu/
tFMkQp2AkME/5+eta+f7k5j/9VoN+dEr42cuOcxZAQhIUWXTAOcQNwtrScvUVFsWBb20fbAvJFFB
qDuKQYDjjG79PWe4eYE+RTA3kRrR2ZZvw6GilV7abU2oD2zzrZT06E1KmfTIjyr5nmgfLKlwQaNQ
rX+gQqXIXU36XBIgCHuFkCxnerhhFxqOb774jVX4iITsHnXTvD6OIkvYHXfFWjwYmztxxWGoXSsN
Kz80x6FVp16wJtfGzHfKXg6Ir8GBzNCSmf/C5cG3uribKTKfyvAG3gwCnY6ilDvE0DyDz/5ZoAAi
dSqXjDIIZ51cjCmIY72Kb0kvd8OzunQ1LcoK9UFaU5FzbpqZ/IlUF02+JK4ZMAUvuAAW4PXZleCj
11i3aXRMiiR4mEpX+xsxpJqO5O7iyJceXwQuV8lHrv87vcGPHQ723MftixKhuxhuXGXrDX67SQLu
nlUkWf1PFUH3YLgEucdkDw5/UjPzFHVp1rhiqPwP1ohj15lw2EFTyLL6qC3bBw6Vn1td6pmmlvpM
C7eh2gUW/etOyaGqXe/DmqTMky+wkiGVXTY7uDbRa5DejtyXY+PvcsrJDzAggiiji8ZF6c0CV7P/
je7MnH8pQ0RM6j794xd0euSQVG6ibLymqjrp4eyiia6eCBWDY8Q/l62bjeYqjvfYDuyhZZOCkRDu
N06+PKyA+7FQLAcRu8g06g9CiVYrD/iPp16dJm7rSubwIKoASny5reeqMvNpsLHKDvG3cM7G6pKg
K3xPpLVB8krQHMx2SXwUyb8Nb1CeRjponz/Sb2aHW2TvbBt5OF8v/1Zeu2wCwd+0nknZHlHmYyNB
kiNXu3Dk/h6KSLEBcxR83BdjAq4qGmUYWVdGDlVDRgU6v4nQm/Zu9z3hgjFPMZI02xOpz6Rit6S8
Z10viLIt7cUlhUjjK4xv8I/ysvCSivCQewsJzFms0I2tnyn/us+2rYRKDY2lBS2KEJc17CjcsUk3
wqZ/m0diVY1y23NIEgyiKq07dy0ENOnnaEqGCMQzDnZJgWuinx1/sTGXWEevJDTHHrdZ8yplSwTq
yy3I0uOFS+EPUCQMGZFH9aGzLG5SgITR3rAYuvKDH/nIWbwELMIXCn4Pir1d3XptyFty9KS0mvYc
i7GUePOu0Mk8xEikq6hXEEBPlG4iRCivXNv4CtvtSNh4Y7lrnLoykqeMKTWgiRjg8yuoxXEpWpeO
WwlrKcyPnbs32blvKVDjA07QphC3KCbjyUkAsyMZwcTkggBHvvb/ewGhITzai/ORlq17rBoNJSgm
Fu3k9YxxElcHxMaC+Fi243JIHnwkf/oPzdrmh5HjQYcu/RY8GSVGJTq+8kCCaCao0PbX32zZQz32
WH2j7mcb04RpSYFLHENGiPknANxRgutWyB6Oe9SUOXzsDR+oJb5O5IiTiT3QW+t+SE/3++5qNAuy
vsSsZo+M2tGTL+nNu83TI5IEaA2vslOZMFrR3pHchR6NbX9l/WTiFYSHxiJ1w89qb2GPCQguoKVh
+EShndLRH2fEe1a0hgXXX6Cfc8p9F7pDcLc+1oGg8nz55KhsbVjTcUwinHwcEnbaHQWdWJvT86Cp
h9G46EHEA0l4Emel1rKcqWNFlhgXMw7J9PeX/CvXxrU9zIxKk3KFD+a5rCKMlljD0FekZsc4MQVV
9JvaMH6U5AIB2bdxJzIQ9Wt+khW+sexz21Iwfs7xa7SfPTjYSD0ERVOjLRmTsN7M7/r64jrbHb50
AppBNuNW1i9wr4GsVwkFms6bkPqkFwS/hDHUHi2+/Sqz5VdifQ62k67QpQbY7KyO/r0WRey2fwzA
BQAe+BbIBbubpAsTru0go+Mcj1C+zgojLeIrr0G5OO/o6OpsIIDUc/TYoSRwSeYduZifQ7J72LQr
KSveD1gNr/sOvO3ZXWkGbytPd6HIjBV+CdzWWQytorN9pIPvZablw5OkcC2sdbAxzpMoDbJQL81r
RmnLWMCDX10FHTrqfS1z0CBaJTJc3yflj7OV1/so0fdoOk4dbCTbtT3Nqh6X1dJvLRo6IB7d7No3
FtxOmEuokCP0aN86+PLe2+LQp6hJqFH0jxpR+Jm7EWfPkJtUGTeggUDl0jhPzDRYwdj56GMGXH+R
81PUAoj8TC8S4AqyFrcNu/4W80UtAtNgqoYs/ZM5hZNX1oROFGsb8/un2KPvOLtId9ugqn60Shmr
6Xl6RpV+b79kosgaAaQ94s9rvbID5uBJSGUWi8VZWlcGhW6WvlYX8Yu0ppLdWDMPZKa1hsDPaoVi
0E9klSSIkmqRPzjnABDSaZnOfiYxyuK69suy4aY4zB8/sR9wFK2BJ8eINFiZt1Pk5e4WTIzt+zoP
tUxLc5X9RApCImyIC6leHTATyFOJBLrO0B2j+f4lwCIyWVp09vf3MGTsRGB7oH69Nj9UaRdAHbDx
vB/jXRWFieOa51E1SgrBNQ4b0ffC1aXszPFTKc44+tLGEg46yZK5Uq6ZsyFpa5zPdeN0r0tWSR+H
h+VAHW746FmCa9HNmJURX9U01uXskJZ/hxV4z//Y0Iv7SnnODLjvpDdvOrLh35wJNxkkElM4FLl2
MWe2s6S2dfwVs9Wqa0YCrSxfM158K2y54qobgUW4eDVhFUFlpZydKSegQSmRNHrYleftCYwfId7u
2RxrB+A4//eVtXBU/PgUlIEYYZ/dKi+S7Q4MGt1iHo85DzCVaUnPwUkeL+u8tMtw3GQzrLI8Tz9e
0D9et+W8WlF3dn7qNMBms+PTruSF0Wpd0DEw7gkNpgcW9kPaufCCR1IOcZ0OuB1V2gEX6FjGU+07
DlRXposH3K2fVsP9xhep1VTf9/LeSeujosJ4g/cfR9P7inH9fHUALtx+d81XhX71aUCmlQvxXW+s
+1VlgljgkpmHI0j/8ccWa44OrrCELUiJx8HB4O2pXNhCpI88AkK/mi4sXRboj8gMV+oAgE359HKQ
vzZbzVh2cteMCb/i7IDaBU5NR3ZJxHGHg16M+RD2Tb2GSJ/v1CJNcgpjd8BLDkpkUbm4wXaX3fNs
XTe7Wr+P2kohKkQVgi+1DaPBc97HOK98iHFUet7g2j/GMBTUD82ZaSZpzVJyzSp48+CuoOzPP40J
WzMCc+iXsyq2N7Er6e+/OQq6Jzg/ZrYP3OG23A5ekpAs/xW0DpMvxfAid+tCB4JesUcJiX+ommLB
Z0DQ8tFT3rsQOcFN8fCqrJv6wICLBIiIumPWst1qNIUzlmFxOooRTjEg/MmjroPoc6MNFqQ2pwJA
sDjxo6AfQeQDZjOeZVgzajgtXDRN2hsmtCW84zDnvrcJke770AUkxyZA7UfMiEquuIaNE9o5HYoE
v5vYf5Uof4Lv5yDkDfzmItF6cyPBSnY/yj62UebuMk+Dde4bj0fTRWkB8Uz9o5P2JXlpHgwFKtzP
ef76sQe+WsNEjcmcjqKqmuOz4UC18JJXkS8aIlRjppCkZ479USADYhoc8bzGvXJVs39D4qPVc6lu
kc9FbBinApJ11AvniIEwbyPEjcZgOOQFFBmaqqKaaV2msbhBC7Va9hsqGoqfRAosy9DRLAEUO/av
ae58Mikh810jZ96ez+ItweS6iFMN4p29zp8owASc7GdOM0isX2/6Ts2tUKJpG/LXzFU3r1J3GNde
JR4IUdvSdZlgSS63/yPeKrYY58stOlBNFkY30LtXodCTcaTtThrBEI68+/LpdCY1csS3Odtk7DwA
mZrQdc0oH4OXiALf3OKPHirgVcpwhLHrO+8m/C4A4Avm4J79wH8T0C62AFTkvYfQiNJD5KlEplN6
TweSUBBK95eM46poMOpS40pQH8xQbxXJ+LaGTKG0oyFvNiyRgYl3kQ/H679FjA/z2V//235Je6F1
z5kWBr/ce6NIqHqdNsNzZeA8fdjw2Y3301uTTvVvfvI017ufygivhg37EHGpJR0M8uyeSoTd1N0i
8kkIPB5f7bySL5BSPDml1fCMwUt+MCUOd8pa+gz0Tal1giCSsjbVuUuateSyYbpYKPo1ziPkEXP5
g/sc+I2S3aFTft6Q95VUBv3oA9m1D4MxR7uK4plrEj0Du2CCkssotko2OJjGYwHMLLeJh0ksuh5Q
+bf0m+/ceMBSHd3LjZMezg05TebFn/9eNG+7LyzIooQlU/53Zaf4fqEmFJaagtBL4pVPIBhpSiZn
mj2xEN8WO3hJ+w5rmRKvs182KW+1uVLdQOgCI+aqhNXICN8WlPTeXkvw3v10ZpCpJ8J3n2ShVJAV
hII2qyy+UvNCRkPxCacvMCZR3p0GM9FW90CdI13k3tr0A8Ca3bIbrkRJ4cMYYl032cgrx9tyYTk9
r7kcdiiQhYT0D7gSsLWp/ir7CzH9T/yDvbuZ5v/Yg79yIyFfPnOO2u/pYMTLhdpsHinmIMt1Oh1M
0W0c5HcPL9zLzeLcxnJBuulRx9i1fIcCnFwi1VP0tvsF0bgdJtxcMGfRK3ELBIucCctcR0l6miFD
GOTgWUjaHeW/zjcTcvL7LYOay2YMIRhzve9M0gdEJPyS3Kw5OjDpBghfkpQNXVnMdprs3KjH+MWx
mGQflSodjVjEDYo+/qh897mBzMmUfEPib6lbfRJmogYv4evOB84E5mQEj2eVajFWSZyYRcumjb6v
f4BK5wO0AHSZg3cR3pbQMOYx0kr/XjdYvSdAMYx1zwIdeMMTLLRUAkyVT05DvVBh2YmV45UKIUVg
MZyHxDAsrj70CRhJqo1G62+HZ17FMV/KmGOhogs74RIshGBc55WnhWPr8pPrCBXWWITCFEKpnujU
KfiNqudLjPA2N5bV1NYMjKuLcGbUaEJEA/4T+te3pxfShDPzdUWUqVhg37p8+FOgWdclwxL+5G5l
mVtEnss3WNDrdeF9QSn95vElLK+NI89GCsyqJLbg18rgPQiHk8EulHWzMxCOiF6UOJ7a6o3vWjrX
+aiPeBan1yFf6eJehzqTUj4nVN9Qb+3MhDHLSHUTv8hkwryUzknY0Lq89Shg+W5zGasqkI19Jjd6
LFFC9C5j3aG65LgfeKnuQ33UE5/u8RYyTu7fv4wLWIztuM1+u4RYfWaIErnWf0NkwXxQW1k4e+re
bA2P8e/P8dTpnIxKEynYftaXqdH7wd+ViY7TrHRJoEE+YjJr6JyeP1zrROdegsrQUpLRl2mt/lKD
VRyabCRFxwE8/NQn9wZ7mqbY9f+/L+LzrvYCBf2I+ixnbGt/0ibs5ZKxbmjbt0SDNVMaXrkGO37X
bB2P77GafV4Gy4N35Yb+KMYFNQE1BnfllhWOkxycKVn2FTW4D4g9mE18IiLW7SAdHYIMsq4X11qK
1cFAZOtKjPmoM5wspZPLEJJ2I3qoeCfw/Vpjv4TLi0pXh7MpvOZOJmDY268MvWZrC98POAiD6M0m
UHveskvsyNNQ7nkkmarPBlyKQv93YCHqEbZmfzDMt+XkkCOniryfUtHp8XpQ4gKsO6ZdU4ZSALFo
vAhNcEpoDSibUfPD05/Xcz+10bV5GfqcUTvYqra30NHLJlYiKQsswC8+4AyQKaahfaj8fZX5fUdc
RpcgUEFzcpfQ628XR4tqyChGXhuXWcuBZJdQko9q1Y0NwMudfXFojIny+hvfDvjdLGBvvmaGeZbR
JN301Dtx7tkLCMPhjl/Pe49m+2O7oDgLuenjxJb2i3HoCClLwGB6+tzaIFc9ksRvOLpVd3kENRHn
Z0cOiwHe/YHdPSld/TcUQD2RbKL2WQf7zbK+EAUjVJ9bEOsBEMP0nKKwfuldU0zn4Rzn3zOixbPy
Dq/61vii52dBS7qBGaDsiXeocQHZpCKWwdqEaq61j8UYedr0YgHp2V+F/yNMvgBhcyioXj+Qx0tV
BRoxfN+xOhsYByBQ6DRPgwyDpMm8vPJ3H6hE8Abau4bFCeRxeL6FErRJY9p/AUa+YR7NqSX1EvYr
GIFKWd8hpZG3d9Ej0U/I4UFQISqXeY6b7PcL/hRuGDEHJLtgTtLG+yhPWEdFTG82StshhmCJDEAz
mstT0wpa7z/2E82o4hmDgAl7+QH2bsNjtbhuQOzEoR/4lGTaUnp5KEiv8I88IjL3pKQT3TKssvaz
PX718Iw38YlZHf+xXWYkSJYqwnni2glVNWdDTIcLaZ7lowq3pudYMAQQlaUj+SSmikBGNpzEJfTA
oDMiUc38MsqAtr1CrxKbKkZmU1ohgRFRPY/LCBh1nIB/wOAbQ37zgIhIHaMKMuB/xlk+wNC+98hG
h6WsNy64Dt2NjioxgvjRm61D418OGQ+t7g8Wfnpi+7xX1p/dxOFWs/gpV422TpF4rsvNeDHXhQFp
fC9MvZ37ZSTHH9TIOXLHTiG4JHXXhqAPB3PvenGVeDVY/hYfMYB3fd6jEDdCrCKZC1VgYrOpC7Xg
iJ9h+nNdvZ2V753Xid40lcL0Vfh3/JcYx2YQeU1dTByjsh5wRC1alti2mRnDESXelqEQLsor+JD9
Ne4jhemZbIjuy9f8VtpsHhhcnJDTuX+kQDTpUxE98muNdeVYfGtyiOSAJjq5hJ6FyjvZLftwryv2
VbLSqFuxAM18leN9eu8d2+qPa0D/TyqmUkKZ3rQXdo4TtIUiHrPi5974tvRdJmBhOS1XTe+z54KC
uEOd+c1wdjdz4D9OZjvbZU+tudp08tULK5Bw4PVMFbJOskUCSr8QC/zLZrHUexGMLyvLpy/JKLnf
X93PhH6xDDW631NxXYXZFX3X96Z/+zB6656IEYDe+25UNkhekJBvPMHcMUtXKO8hUK3oQ4OjRwE2
/1WKIrbGE6M8uE/bi3xxvmNU8mbFNEXIcIFa0DuQt4dZVKKPANg66PsDDZ10rUP5gZYsW52hbpoZ
nm2dixcXY10cz9MRORgeLp7D17dYwPxuuMb+tdpCwGWCh1BQZleoQ8HoY2lqGtsRrz7Cn/ceuTSa
jHqY/oMqEyeGBW6wDW8x2YDnV+ZA52Squsdh7XVstRfNF/MLBlOc9XUKDbxohcx3RbM1pF4AfjeY
n2PbmmVVA9dw2Gjc74oIkKKSIxaAZ5BOp6911NQ5SLkBMgCyGErF2A+0yh79Dq9b1Z1GMGbOXw/d
GzWbm0MglD9fUQP66BsNtJDuHplWolGBONA9OjhvM7JsT+V/ofjuLDZAkh4FW5tKtPNeI8U+jGc3
Q7s1W510ftYpSrVsY+T0YvJT2HjwrI/e1xOohRVdvbP48nazCoAykFWsVA+bIG5YBxxUBTVwzGBB
hKxP5dS0vEYtD46rhcCUg0ZNb8ZzUC7lA/kprYsYjizwodiMyHL57ZO7xADHyuQgOGJ6h8vob6rI
4g0rxezcTfeFrLadnTA7B+jOvgZvbd/5sDvh5wJobVf9FplQZnYCDvkXGWZp6SfSIUgMLVWyE+wx
0hr6R7dCZTzBVKDEeknXGekhjWA4SWv6eRu8f26aM0huhu3kwyacFE3Py+Pr5nRJCuTBycCIV221
MKDplRlLwQ/WvJKeKSL3Vi5W2e6fDUKoKwAHGQl39NuWaYkB4C39Hp1pjgTIo12jDW/TyJrErqFl
nIxXfRPtAPLbNpCk85ZK22drmWXyuLFT06HCvPwOs53q0VqdLIo3B545n2N4Ddddsvaas6xqUxxm
z7WNQyvO+9yseL9GovHkaKl7VFFGmENrxpbyeFqrAuvyXA7coXcJHsF09gn8b41H+GS25XwvXhSx
/JbrM6iepDp5rbSe8t3qT3/AMYpDys5tQojDdmVtk+J6UWXtYCsKSQXU2OqRr+l1wNFwsD2xRTgw
NkSAZz9bMpl/SjGGshUmsLM6a8/+7TNkfqN1HPAkYDUUUU6dkckaN6ZK5/Gx7ert3OkDuLy5fB7H
EqbNvUU2KiNf/0GYQyPzRBXtztqvYHBTqVEmZb9fgEVSG2hAKxmSnC5plK9LEefvSIgMZ7G1o5iw
4g7TTW9JJte6EqzSJ0ahfbru/UZk1cOwASM1yPsa4FJeCvOZgs83/J2Bzfb8jSkMcRt1TyRi1h4l
ddjmsq2+1lvfSNEBhGzevpTXo4CDNTyDqESnfXeoga9Mge8fbgJQpIUpjT0EQ6m2wF0dr3Ho2lp2
3CaGEPkQm1MQdN6Daj5BPsnYckUoYXbw9ykvpqf5awjGHFqu6Ey1ZEddVDV+q1xYXxwIkyCfoTyt
KVBWO2CGkX2iPV+t2vw7B9DncS3Mn2yJQ8NzWJIBpQOaLhXh0lHwIQK703mRHBbx5dTk2FGz+Ukh
Cxgmr3Og97Ak/k8v20N1f0wUac2CKxSOLx69msnUFMyXe7KDx+2DpoHD7QAYanfDV6n/MlS5D6px
8Yxz1RsW5uppAEpHS0UIRBdXXzSubr6rd27Tx7//uC7XWGFdJNMX6dISM3tWmcQ1FXto3h4I9MFM
FKDCz53kiyF7FZgNaMCUNOzuBAoasThIMMlc1M3NLHDGBi5jb6go7LDeLwPkBJExg7G4viE2DFhd
6zDgc6F1LY1KsLzBv/+PMJY+JN7cCCisPyXtaohfwdoZf75U6u+6ZYXh4dEW7c2Qqbd8xXZXov1J
f5L/mF+rSpXSAjEaEsxwdjulT5hBst4wGOVfipeGzmYSWwfBOUERlZG8f0ZIK+nCyvE9I+fypXno
Iv1wkwo3wHsnzpD/+hrEww1CcdWymru79DPEY0Tkw3yysyKVJFPpu6MQPn2RqBvhYYbYF1unob52
ZnfXdn/Iz/7G6KnidQw7xwBalhMDn8hGr2k39GqbDcTIqe1uWFUFNtDksOKNvivjtIKndwyGXvM8
FjWQeZ0rVJMhKV7V44/x+449q4NESOGSy8cghUkYgglvEbfr0e8DyFpFrzQIX5frwjwAlO45mLzv
tJO2faSS12Uct41sE8ef6Adc6aT6xNdCpvQRgPaZ7LHZpcrua5n2v6z1iJUJDFDUjYSG8tihGrVY
CPXB7sV7UPA2JFOC8iB4Hb7nIV5lVLM6X5xuhPgkkqcwvDk2Ja+uV/U6hMIeR5K6mwyoKcVznV1c
gMKLPCGsI+yQkaVMl3spVRPmhJDqkJP01JOdIn2EeyXloqkVGC1ARKV5+fKVnHXEfoh4PVzP9KOr
WpiP7MsXVNzHJE0dKV175r65HesCpb0kjEI8n6B9fqr2Ju7TIgJpp/WZLorgHBX1c2hYVbyD/b0g
iQmtFVF3dXTabpv0obfi6kKJXZUXlHRWBtJCaumrifVMSWhAOQbrOa2Dqw0gojua7pDQPPoRhtqp
HRZaV1NqqKi03CjRrwU5am/U5qsRYIJWyLNdbAZ/Jthzagal3z6LtqHZPEsOZhDiOGc+bYMFhUz0
Pi+z5WJflhQXdpvO7RlJPRVo1tUabHRVsQrq593IpuXBMfhwJttc+DOsYL/Q2auKuXguajqwU5Tu
BB8WBSb4AuKc9NetZZrSfaR/cl2btPRD6Eie5W1md0QbjSeERxlq6IPl9YzleTzZ3jW0ct/lnJSg
+HUBWGdt+1edVUq2plwPA11iF3NSPBIOk0wwplequUG4E705yt7lmW7xpN3ihHn10N8wEKf3Hg/8
MEVYNPgd9u3M6Lj0dQEYw4HQg33zaBt3HAicb53hOEeamqgws2j1/ue42ZTWHrFyOxUR1XxpqcAA
jyjl4FY4rnKdKxhXqAqW+UWdcF2t6l8x40OL/BRqetvqycMBLIQjFwEyAGIZvTSzc7iquKe7ZtUt
sEEKQH11ndjSfS7LEQVdupi1NcNaKJjdwwAf3N9SIqhXFo1ID46m5Am2YXnlZanx2Xk3J2JWOZiA
SQ/DFdOZyGiXBBVg+EgKV72mieFqZMedRRvSHxVQ+Q66+L0qD+mFTWsxxYvc5U4wz0hIYyIVk8Z+
QyhLssbjT/TBrDFMfpwhkiQtilmm6St2L7hpTUSlWZ3dmb5wWk2gtSGOWj1pIJ756ui5LfvZpFfH
TMi+B4lWZG485fN2TW0a7d6EZcdRsLoebav4S5RZOzcLADWATcSzkd5gV6h2ekFWYee3FxqpvBOL
aHovBOLReIuwBA5wW5T8M2ZRDdcUHFec8zeKJNMqxhu35FeKdHdSB68wqHXzhdr4ZDs6x8F1iryT
09dsyGFdWSyQPKa6e3B5SDiViFSSmG3ilUhbe0o3Qc5IShbKbqpYknMncwDgXnfVhgMjvQGdQS6Y
2A6J0zyIuyBEsUxPfYJWRrXodJlr7u8AZ1TQF49OX+UfZq67J3gUdUDIecRc8+b1iMN7lgYCXp5H
vpGf7w5pP80imTSRZoSqv2FdtUBUeqOTfknhBomIjHwDa2YzZNO8Q9tN9j1NRnw2LKwBxXg/EBQC
MbfE/yxtmF9YGlFEze2sQzrOCp4cUUAMhQn6uCmOip0N/6ITkbSqTp0n+QLIpaX2QeF3cb75F9Rf
23AiFLrXuIa371co+4o3n30JSK1qmBjiiER6kfnRc+etFxwPxWKXXXKm+gU+XYdoxuv5I/B+mldA
1TZu4EDPZq+UuPH6TQnLyWnC2/CBR2hF3o8FPoMekaJz6d1GqhPPrDlTE3bWZ8F+XfCaDXalBXdC
RyVmWCEMKLpeWe8vJJkOTjqeM/A0lRGQ2GpB+kng6KcfTpidnaN6sJ5L33XXAb/9mmZ1l8K9Q/3j
qLwa4zjkiwUZ8xD7zq2/wdMkwnHSAdCb9a3dLyAdMtj5z+GOGbbLCCVLYBMXNTPDojUSLkUeIw5D
Qar1FPX+KrSAuTLdpyQvcOsj1Q2Y2nzc6zdTrP21bs0psA5BTgW5vNCJZeWvxhoWrxIoB0/5f3s4
f8OA58rh2Gjevnp2w6QGnN780mDg/uUo/nH5KnenWARfvUDbhiVRSWw32i+TR2Ti4/vEaL7JB+Mq
on8cWgPo0pVlD3Kujix8ywxzk3nE8MF58rdLvETcfVFB1Prm4xOyES+ZjWgeLa/d0fHAa9/l9ezM
AgRlib3IrWPP/dU4ONkeSq/sKoJ0EzQ071LKI0VGJonVEPdOHDPcGqAsFRaNdOJCTJrh/1f8JM5o
rsn5Z/r+U9wP821+EeZgoqzfND1P8mKqdBat8TR7dUNIUnfRGUL/nUJPc9sphe+U4Ogm61DFQc01
OVTeg+Y+xUxJpzHWDa/g2FaB35n4Vb7nC/oySbPKe1ODegLnBx6UV0Q5MjZDVoa9fhvEnDS89m3+
k+L1gg6+G7+oeYM2Ao+2giQzW2r0+sNdZAa+oO6XGshPaqVNjy9lHCZISC4tssTzo5D/oYslDMsk
yn4Bs0/GBeCkUQ3um0uYGjUaV0xnnwrs8oEa2fTUivRddxvwUj6GFssuKwV46XNiCspScl1+4tJk
rEXkuuPJXzYSQkeDq4F+xLpJRzvXCyViIb08KjuBJkd+/kDwVaW9pdm1obw/z1mD6/v9umsYZZ0n
beDujwIbQhxi/1eAEIHeGYF/DJtoPJ7o7B6aHO+7xJuO3syDloog2BLNCmkTMlsUyFfN8SFSM8OC
Gygo88p1HUxr3VByjjLhw5sOo/GZbXp+eqXc3mcB0IkmhoydU9qCF4RW9Agar30ZgAoqWwlXni6K
XnrtQe2bUlAndlGifYQELbNeeBIx2saH4652FJWBJfe/M+fzzQgUHKcIXnt/YmUTRfryfR2heCM5
oEFiWMXZtUfR23RA37XCYF577OMsnWjH2hEipof4ZHfnvE6BPi2EBvC4gUPrrnB513cpt4bRzx7q
GS318e/k3QrufQIJ/kPauTJwT5phZHsmaMST+r0GvpyKt5Gv+wGMxKqXV+uPNtYEbB8VJYQWdPjf
66Q9eGnbnbMmF0hjh+0vRPHj6HUxHY0h34FMNv5baf7qWRjqK96mVMJDeeS7wrDPP7b+gS98Rahj
rj8xbU1gQ7WqfXKctJ/qo+P/FKN0MLjT1LCKQPee+0mFrceh67qclTg4YSQl0rafuHQXS5GGyUW1
REy/zke+791cijU5gDcTz2Hn9D5qBsGSIi/zCdBjiav54OPdbcnXouD9E+8lAcKXBVENRxD2Ao5X
izuqAJC8P/3hI3fxFERG6Kkie9Lb+mKbcqEbmpyaCSqSwCCrEGORS4fcqmmkrDxawzANHSc8yKmW
PeC0YzPyPjnz5fdz7bjrq6LdMb65pvVTpPlQIHp1o/EhEcLN9k6B1fXqHeZoHPM7M5MKhA5iM7Uk
laevR2KHuOouk5XEeULymVU/0XDX3k9frCQjPsSMhR91E+v6u0NqaDTwc4q6YFLYNePEl9BsC0Qj
kMQTfreB2ZHP8aS0NM5tm1ZmSOXblyG5hpONda1dwRYQtYsuXN0YcMe+m2w0tAU4MTMu67jc4oTK
44gyRvow4hgCXm12Tc7kc6LUlDv133kjWQmwIWueBf/Ii15veh+RP0Xj4qaV7g3+pd3wKCwDeGol
CjDf4S0HVYvfdIYAPWj30fQ2u+psbu/5sFMyR9X6b8D58UX1k2Y/xxH9u0CNjxGAIREjGA6wufmy
f09bNoe9u77X7x+wMX7HlZsH9U7tYqyXaO3uew/cPV56569g6Td32jECVzW0VLKLLJY0zKkV3xGQ
wvI9DWVzGBHxgZlOit/r8wG6mw0epGnYBUYQu4YR4vtyQv4osQ+pENtCY3Z6XJLQeoUx/XHCf7Mr
Cmp28P/G9KB+1Hk0I4woh2yzIX8NEh7fhzad9lhL5ZuLuJs7qQvCXwcGovox/rpo0mDwsCwRH2eM
cR1L3w4hDUFdmNuDaNVcaodVcrICFyvAJMZanj+K5VNpwCUK10bHWYZD+tHrNCeHAjuDfKnB4JpJ
QFxPFxBqZ3sqrOFPcqw1W/z537WTqduq3W34y0VWIm0bMeDE+T2wYWTi5Wnzj1BGuyaBZYngYMMT
4Zn2SNaPEhSICHUBCb3FwKg0v4v4dAmHuGWmxgOzESCLZPWCeCjlt0MdiM1Px3hvQjHHepuRDN2F
bjmiiMtRllBhyQAKHTqzz2p83jAw8Fq4dsqowNR4Zqe4LWsFwl+Y+lnvvyEyDIQJXKnCLJoIu9/P
g1OAUnShzw4OlxN+HmXIf+v2AhO3JbI0GbPyBFql2/hLzsLxl3lwX5wmPKrqfklzw8hd0Pv+H2S2
9db+6mv1t00MBQsR9YMNBL0z1m/poI1tXl8P/skztv9knj97w9v8UxvdO0Ts2hbJEpXnnGwVrB9t
QFZA8m8Cri/dphzwZsJxy04ZYGV78gxc8J6VgnF+Lukd0iZ6GXogTDUUeOMkgBmlAEyTywFP1D8U
GhJ3p5mVyZBAJxjWIQKxeFpniALHLrmhzC2/jXRTdeAaO5+pcUfgeYYwn9Mb83Cyp2L68rZW+FwB
zN9ym+OsDYd5UMZPAIgHv7KOXKH34qQKvd4ZRhmePeljSqB/bCfhwUNz/68maaKZBmwJDaZlNUsv
5WtlEEbPQFiavqQ5Z8PQFKl+aOEhsN3RT4l/I4yxFRYwbwL5l3Tqp8yut0spFzeHUEsWL7bhDBhh
7RRF004AluUMILCs4u9l/4LhjH54J7IHi5+j0sA0UtOyHM/3aW83U4dzuZ9qH0YUNmw0dLeCCD+C
Z/hCGjLBxGYBVQoF/fyqAj1SuGJ1Jm4B49smJo63zCY+fTNa3R7IUFufnSUEarMfV39BJ+ZyiEJ2
XFnoI4mq3/T8RHbFG7jD5gbRkY9YgcBLz1gY3SIn2NFct0ncRXAnCRIjBwYbMl9fIfbM2feykivV
B119k5gb8y+Oa0QMQP0dzGqlS0N0zVriZzX8Ok1Vj9z28viGg2rm8H7ayRKqyoLkWj5H6j6vAoDW
MPIGy+5aRCrpvv5Ag+Vxx/hN4LdWapXGb6KuumvvttiJkyy6OoKzwsg2NO0AKQ2bImNwiu7vy34T
Xiwd85JchNvQUKK23sIShnlnGny+jmjNa+7/csYe8tc9UGju0dS1aYdT14CYYdTHZgJsvciJ0V5d
hIAUwXzj6SNy2SgJDWxVF/RzZF2kyxL1yzooyev5gpfBV7iOfZm4j4SufHfw/K1eBxX+/b+H8GD3
s/wiLp6Gl6d5WOVpPD+8a+aZCorxpTu3nErYVhsGjwJjqt0sVqyf7evTUwKn21Hu5RutNy6y/Xal
jP/SLKoJNG9VnaAcxaUtNKY8T6ra2k/qHvhJw1OIjIUj9BaMrNti4Meo1o0eRzZmK7DQBmrcw/h/
TpMcdaXkAOtK4+TTsCliZx10EO1O2T5Y/FosvMJ2gosytk60/aLAr/li7bvnlYV4JUQTbBASOt5X
Xo5YJN0cExaScJb/IfD60vxs/F2w9YmZWMxD74N++0x89ucUBH0A9RbjuwkhBCQfbxp/ViB0ss9B
oTmFyVcU7XCdInyjcoNcij4r+nluYcUf7TqishB/ddOrGrj0h7JOGXLEQwsHs8hjR3DZsac2AlAE
Vl4o9vylEJqjB0Hr44olM2B8vSZnFUpSMzJbVT759sUvGFVe5kJuzOjxWXM6NNjtrtCBfcIg3iD8
RjKL66W4cZdZqB+w2uxtn9kNivN3hbYIks1HBtr6RDAbYyheOALPpYlfWCdMsv6na+qkqMpYM2oR
tAm3q6BnTwgEyysFG3tpyK8g8LIc1HLMCZjc1HWlureULdJYTHXQ+/q8JmuBS3j6lWcZ7Okd/V9r
6/OGCfk4Bl5Tjcn+RuL5GMfebG/3v4aml5mRd1yqkqQbyyZE41Q1iStFBEuwMoMi/3+FT8/fczzy
bYrqWJy10FaymkE5t3l+H9mwU0C+ElguYdA5E41xei6ojq/EseHabNoizXKw8Fv54L/3Qey0AZHZ
luf3X4Z829dXRfGQw5zG286m8I6oluRCfggPkG2goUDeE+DuxnvAQub2dca8CVWa7JyUigzydiwb
wYdD1alwpEHb8r0zOUiRO9yeZMuZKnJQJnpZBYD+drhz8e4OEXQBSMhbfcKe1dOA5EvkQg7viK02
3+cNJ7jY656Wzhqv5+2sF8sJAZLc0ZJfQeUAheCUpzxctVmQo4rrDDjk/Bs81Cjd2hLxvhs8+/7S
+OENa2H+VAcevn886KmT664wa6UkiV2r9jnyCntCCPCspDjABFjGNZvdSDxKhwkR1ZxMUi9MEYo8
iPjCeyA6CeOZpvUPwv3nIINOqo0UM0waCvWdY+W4I56PoIWKi/omtbPcP9V/pNY3jGSSFJL0pJAU
SXjtShVoJ5k3BVk7lmTUcA4Sgo7sf/+R0fa/3UWjQkaSxA8wmBdkA9kAxSlVfN2GL8iLVGmA/k+V
zrnkL7/uIFSw8X8tptEb9TLwNWmh+H1RTVyeuqSaWewwx6N5YuXdT2A5HZju3T/aS/4NdY0Rh2Vy
IzrvFnim1UO8EQ9SQTBNhlPYUIo4im0rKQN6EJNiUC3WybKxPQ/MCaIJS2tOFx9ET20sn2JzjWcS
x/ewaUAx+cdnwh0G8IusHcFTlwhxHCs0ktEH7TEx6nPnqHoNTflmuue1mPHF5zYLWNyHvrnhxx8M
t7dR7h+D02J2ydFWNrdDSmY8nPPy6ByvuCGDz/HvRxc9ZPeOukq18AZWkfmZL6dSkN9UIgSZzeFi
xrKybc/IKgpbZVJa8tRtVJNGEa04sVArQSjx3XE+ZtgAZh4B4QGgHq2BhLGOYv7mAfQRQPtOX/JQ
0Ms7F3be5O1blJZpMlSliTGmCoVFyyRo/k8UsGUUEjy4ypIkE2CaEbd6xn6dZFky6oddomyfV5On
TON2CogRlT+Na+WB9HoMwlFCzUIf6hmjCcnCDw345sApj1KG1PwNXsqGOguJq/A9Uu8cso107zxp
haoh/Fv/NY3p6dBFQ7dxvSfEzdPYZOzsyHIafeTDDLnCFXZ46lvxEGImGFQA3Lcv+JucSJcZseIH
6KUDiAvaPibN+o+OPuKP9Lw1vcLiC/yhX3vL62/VfurFoTu3qa4xmNZoy8NHjVG8XT6qc9dquRcB
RYyo1CINyb6TmN0014yRhIrFZA0IC/BxlbJLLiq7qUxiooAScRtksDtN5w2l6B/IT3wvfp8aIS3W
u+PYmy3MZRw5YCPRZHU+he6oUiZjQX9Mq03lEFhsZMyAVxsUopsrfIZZ2SKqC/1dFwRClJjxfN76
qu+5MtkqMLgG2ShUUcmP/kwuHTxGLG/uXIxsqlZOoLUlYAIOq8ugpKfRmbYbv5wreBfwIJfn9b3r
CcXyJqawOJsHYKtM7YABZ7n96bx/hmDYca9rzFQ0p4a2h2+b0QJ+NaQj6zZYF9veyd2GRYumbhqp
dWmAkW+LMvoUUS4XkFqqq0Cne/dTE3Pu2Ga2kEOc1Uu5tDa9krUDF5JZk+z2rei78VXE6UkHHHiR
i8N7/1omzHJDHzqjLKxBc11tKo5E1NLpXmy6G1/5zDGr6+C6TmUninQiKtkyoxQC8SZr3qpj6SKH
vOPDEm1KRLxxVbuetmQ1rHr98glZYfB0r1YFbePuc7wvJ8qdd2XmzeR1QXM/utUalINXtGDzO0y0
GNn776msS/9BoUPfRKuDuMiG66hYY8x7+P/8dXdmoa3mHuTHt4GuNVhObeHPRB9K+ECfhkp66vae
f+Smn6PtCJTkEAhd+r+0jmhvBb4c0hBoD0GwQPJg3ibuAcCt/LwKpxgsYkt0s77tORMMfI6ZEX8F
w8RIC8vQl/2JZy4YD8uBL5OKnOipce6jz1+HNbAzNFYP9AgGrB1ruMU/U+ZXEzOcfaGhLy82M6l/
cIkiFl3gM8OoW8mu3L8YlrMusXQzvGrW1OJf3WELaws3bT7jeZvUjDflxZdJYEjQnVjk8sevbn/5
cWou3MMFja3oQP+MdpAbf1E/wrpClnsFiJhU6IMGnrmust+CISPcM3X0+CbDdyMcs/lPr/c+WXYV
56Cb1vgVRzGn7dF/BYGQG36IwvLTyDf4g09XZZItA5Bv6u1inFIv71c31wrOCrsDqtitNw6PE97v
FnFGj/KSp4U9x4rnkq2ptXX5RBqRriEQHPPtY8rRW022y8PRtFA+xtTjRAPGD0A5Mbf7d9tizmSu
W9VsIiYR3rY40FzA133xIXa1wqBGdNNu9l/63XlvfgnUlNsUolTAXsOCwwvy2P1PYleTid/q84ed
lJO2M9hBEUWSFH6S9z2hy3I8tztztErwiKN3svRen5BlAnX7Mdyo8Txrb5Xzkld65CVGNv96N084
NGgb39qtmeFNCny1Algsla9oA1UNgn6bcv2OuuGDZIkEEDvayAu92c67TJb3+bumj4qs2HEDMTXb
G6aNFjeo/YSgcbjNhDAwR8eqV4WU89xxrFEeHy/f83rHZ9EtQrrDjc2/g5rm9DUFP6xEMcUibK++
Ac2AWekfaRsowZ7GITHs04tIyl5WknpThwuV6Dqui0B9VQAAOp6/eHnHjOlfzXc8yRtAajMcHsTY
6WPGh1itB/fTBrFZcQqMdRM17C5K5d0PpMD5XMiKru5MuM1GRxwH8LULxjAMqwNxXsRvCVZPguVI
UCWgo0ioFNcX3ndlpZZ/2BC18ASWg9nXgJtwz8U4E01jX8+2ZnwxThWGn4zOUCEcVRO5dsAhZa29
FlbhVWDXJMK8q2791LC29g63bm9wfQS6lRdXKPodrfuvz0VaM1BH7Zfq0OrlH1VJt5i9YMaMHEmc
MwyZkSRiut87DHZMREGlzP1q7H25p3NHjnjUwee3UvW4fTBnq8fLFZ0j59fGHgVSjoNS6KpkuFdW
ebVgqB2rpGt53ia+dv0YgW9s0ABRBfp3ob0bD93cUcz+JAY/4MyiFysETa6/Xxqbtpm/VV8YXGIV
StP5gMsLBQOkRtiGLMbMBguANCiWeAYZecguSXhrv+FVfH6fELyvrzXWtx3hb9Zt2kkLBWwhoTbQ
76HqgDKFfx/WwFAVjwbbz5OjIwQmw3GMUzvbQ8gMPi16KX4sNqG1hxZp+btDK7rxYcoJmQEu1y0p
RdNDjQw/xStfXB40qljTjdDMmKxQL/8sw+4pX2Po5i+cYHnng4fdNYXBOra6LAW9cf8Vz1EyLZV0
qgtNBym/ZDXHva0RCm3AHObbJKyw7RekCA8rXsZJ9CAI5PBQMHZaqx+esMs9LfXm2+7mhY7DnGIO
oK4eNZ7nwUm9ro2UApzzG/OYyhLL64lZT1uV1O4t0QMM+FMNPZxwI87/e5RhXdWawirXMy6bTbNf
LWn5PFyPAiRrWffaZUieWBBu8KerPtPMod1bSB///89DcmD4t4nB5y8lN7lvZwzMq278gqeahPxg
O92Yh114q5TrXLv6E6dx79TM6paPxsXIjpqQB3rDbqbL/+3P9mJ9T/wpgKdaCmMaXCzQ42yXQjHz
EFF8uMwa+RT3Ldios9/opVy3+1Og0oxCPG+oycrm3Q51MW8StH3FFtKNvb4W/65v//w5I8dMLTEh
08EpUfeI2S99kmHq7CKaZ4vymJV5wAkU8cbPYIExf4ZMg3THOhVoy9PY2MXXwGaQRMdMEIUgzaXM
zaSkQOOe/iskuXfIfaZgl/r+hZePVrKvKu/TNv2lI56Qm/+/dUbkT2A6NeglSB/WokmxngBwsfB4
JP8VA8mD9a6I3q306DpToTXNKL5CNW9cKFr727GPDqdo0uahYG10Hn59gtg1+ISTNcVdwwUidEya
dHZEM+gdJtr2SWzRTR61xNo+ncfJT8qu8uUYJ2IhS6x4Pf24hZojHIktEPlRS+C0ptMY+6nyfEyQ
kOEiTBsDuObYxEZz/r3BXMCAB/Ea7VBDyM182aB1MDgc13zBWP/EMQ2ig8Kn6igcWE/zCOIY9PtL
m2zU/OkY9jrIF3JL0A02ohZDM/Pv4HhijT62mkmkKSEhPlkIICwed8jTCFIzUClM5v5+M783LnSq
ULDeyd9tx5L8xCSwyL4Zky8Y4Seuz8y5kiGyZbUuGhh+te1Y0AW1MUxwLMUBw+ytfluWp+qqV7lq
hFax2s2PVcGtGxORDSHCnWbA9mRwy+mNRX2oRqdn4FL16cWp9TM/Vu6JQPn8C+w6uANDP58m2OCS
kjXxmIEK8wXau2v2hYp1wWKw11wZ1t1zuK4wIf2itd1jnAMgvs0Dv9thp2JJvKH5bPebqRO9QkL8
GiKk+owfUO2msuxlNde8xP6R3HUxFf6i7kEPwOPEb/iXCHcNOMeKKoy9+DXuYlun2Am0HqgyWxR3
YmMvLdIaCt5SNIDnfall3Z/9jQrcFzwvNRSV2xaszJyGA5+o022tnXfXHjvMQprKjO1mqNMT52eo
IEJkxzCFodpX33FTzi513UVWH1u2JLsHORAmonvhstJ30rrbBVK7uznailWWQc8E2YHd+eG46eoU
lqxxF2LXbiYAZ3Ivkqu/nQJXkxXarPoOruHhi06cyw4d4Z9dwq/QiYDSClMsVGJtauhqoBLGPZ4s
3fuzyFZmoI5KvfJ/8TvLXwaZio7rW0QkrvTh8MOjbd4YgkoELo+e1cdzASQvb1M7NJyrLurRS17n
41G5xWi0WPv0vbaCXQArZ0HFLnbH9fSBinEakOEKuF/PmUssz+LyshdY7BdJEA2Mhja2Q2AYD1qL
FYmGzvxCC/CMkbe3WYLhJbLJv98ONMktrKOVspcLngJTCLQSCaMZW9b77bo2dT/cBxFMnSRqna1u
Xr2l0hgPop43VcG8O+6YXRd1LtFaOLC2jnDLFsbuz+ynRdOVVrSdBmlsQ8LEYhnPJUXITc8qpmeR
GJSD2kUhnCwW6aezLDkVJZqqBKBObXCHShOmRS/AP4DdbKfoQEFY0+5dZbM58E/SpLQfxZMdzlAB
JbjVlQpw1UnqOi5NzPhgfkRiGRlO8hHaOAmaTHAr/6hasHkCGAJ2QzaVUxBlLUFU+gWBu3BkVhJa
jP8aDBvrIiDhngX3QXteDbx8wDI1wuzNlRDuS33e1W5H8I1wTXAtB5cv93TxzD2cMuo34PyUI4dF
Veamn/enmsZ5335GYCrN0kUTRg46qDD19gCE3vGepkz7/UI366+59p95/yAfpZblpOiQFJtBPGPa
ScoQO+/qKkEIOqhY6GVS7bReFx1PxNa0mO3CBt/TZ164XhhQPJZBRBEhGbXXy3xrT0C/RFEsnkMZ
lVQAHs+Gpf5fnUZSvwni4aUfW8W29F7mJZnnRy1uEVAHUFpCaSA5R7IQ39s8kaXdVAdm9QwmOnWO
jGke8Nxqo13yNMXeLlpvB7jNeddMSCd/HHy8CyBl2jSRkcJ0fXNFRhLHoX96s5WqrjiZLgWZvfK1
kejL2u3i0QaaXIb5hxMqVjjD20zu/EtEGmdTI8lBKdO3u4bz+w9cVo++KZdrUfAi4wQ2nrReS0c0
euBP071PfNplLPwsGy6wk0aXp0b+O1a4s3LoJdoL8pUL84BqP2lOh6js+FiRB6778wxBn0d0f4xd
vemhYvQirBnnW0Tjpa8aG7gGytWPGx8VKYI1hNkuLg6OwOYdfLKmCt8JXnG7VX0autrFbeOrFrgy
S+gwHkMxqjKswiQfwoy15L4Nfuan0OFyg6xrGD8NjYaNjBKXUFzZ0HdN/fa9FsF7xdeNBIF913dh
QoV0BVevaLE9jdEZLZ48DdWiZwgC+tXgVMVhyUjW/4JU8lgHIzoumlhIF1wh1HsWDDqJaK6djHZd
3tDtTZOe7TieEru4XIZfT4rkqOHFC1eRJXNms30hjiWq3tbB61lW5Ls8UVH9eb3VF0UhZdYFPPoU
ZRD8/PPZ7j3pWiIqLYkawRG9oiqgPJwCsEJ/SxWLaGOJpTpTu64I1J6PFLnZFg7Szi2X/80xw+6e
smlDqo2I+J1w5MYBvxkcGnYkwri5jhNGmwyUD+b7lONfArLBuf+QyHJq9Nvu4/frBzKwcdkznaMh
ghBU5RiQ++FfBoOoLKAmXRgHJVm+rwdf5cXuFCZ1eryxglkB37ZAModKTgjc4SzUTj7u3Cc2oqsk
WPk5NO7pliCnKNN3KurR7BplMciNWNkTJzAuxz2GJWqd+JG8URbpV2kdYA9tNf7/f1DmPi3eXyXQ
d4YkgNt0lM+se1EdaUleIuDA4oAA9eUkgWMPlfjhfqQmiVZCpwxafEnEcGPMpgBTVkUIL1WpA/7o
mQ0HxX+iUA/MDhMJKi2Kq77b/5SXbVIvK6ZWUZBUxG5rqHVg3MiHbbaV7QXNtVg2fDl+EJSxK6d5
Lanlwlp4uVbXNZhMlq5PfC2dR6WGtg/w0LD2htIJcsvm4tk3lGzcnbxsI/AVhsh1Qrbgxy9t4pQd
J70SIBDbfZYfOnCBxjTpjDP0vBRsuIZ+ZVtnHduTD55GwPvUg/8eooAoqGrG1LlO7eJ4CpC2dniL
N6nerClE2l8g4NpNk4jizYV6KT7Av4vkqLgodIsD7BXuyVgVbZ0MfdmHtTNcS7Gq7TCshv+PZWvV
8ufKCuhNaLW4EGCqARmhrMVRUpmcNBtTC6939IqCZo+T6PddrWjrnf8TPnWO+dXAnwE+R2F1R1cV
vDf7QB7w26gvBMdvMTap7otYL9xg9VWpeY3EftMd0gcGJn+jl7PSOZKU0yRdKsWTGD6QW4byTu28
ihrV6rXr41fpgSoqT75JXlRMXha1qBxMbMcfK53WybSFY37Dg+dEdYFVnfQqJfy8s689WosOZ/Qo
fC9tGZM1vvON8fOt6y7ZUzDzr38jaml9jqSou+8pwdw1aLPtcdCNvUPQbHq3qH+upkqJYsmQqc0t
joi3H8LZL0lp1GVhBry+0xJyvFYlM9OWJQB0ekX8qINuQaqia1vFxgQopOuJHoTXh9Ulq0GbkEhq
Y4Q6m6DfBUtMQMd2n39HFglf/wVWdwSi9AiFexp5smR3DOuQe1/muWPqEn0uHr76Uw3KZBooLGPW
OladX/boFq6inB2W12bN5RyosobeT3cZrnKFXuv5NGiCqg4BizyupGYbn6WcogT71Fxo3fWElBNd
Ce72PS3lmPeLrMM42fyi/Y12Os64mZkI10/r0pd9BDNRpw9Qq1GVaZON+DANo4oPA3yNlvZUAxoY
JeHXBqNVVlLScTCFjejLJxdCFTtKCmOJjkj8Hl9BxGFAeMTR//WlOAq5gK3B6xKI1zh0nUuu9fgU
6veMNieHG5MrfRYVzpqMIWl/Tv4mh7zdfObRzpzScM/AWYAW3TK/yoCj57gVZPvVYCiok3PX8qnQ
qPXrCSvOkEcmEc1JmaWPBTpJLGT6+8oLTPahieXB6OyIExJLhLkCoXTfUB5oOy3xk9EK7b+KWJyA
I9jQcIjpVylupRiGUIcedQ+weAZl4M40Lx6nBOyk5pw08MjhawSH9ZrJUJCl4mA18FRxscC6nLrH
FMOWNhUobnuFCoOzTetDh5PSi6rcUx29Vvl8UoHwZQ9y/N+OUBc+y5X8nYM7Wr54Jv9mRB2Stn0v
T+ouQldbZyHW8QW8RbD9I9IhcII3YOAq/2s/spiCknAolgx2vyzfrSEsuyQlnD6KKdBnqiITkUHj
y85vIfzXTkqvknP9MnXnNVxOdJmMlQXzegfAZvkhre1hVCa+LoBasefvXkbredv0UnMJJ28nLera
/e8zDS5Rf2v1BZfIhQh+Z+2PT64nb4DOATsnJaCnjXXhK9n5rj8GHIybazM8Joecw6NhUyXSXxLL
qQ3eAcBZHCgGvuE3RX+mYZ/bklBtRDvbSt84e+TsvfMKrLo+cu8+hlUGBXmsxs6U6vUl0t6x3n2e
r72ZlGXUlOuIFbjYFS87+wf/QWCyQNdrZ3cZtqJ1JDYf8YUuVzPaLL5ZSc+aozsAGKiQ3PBq0GJd
29OYl39SDsZYTnf8jJDi9b01bztYjtn0yOP1avJ7eKHbvk8MxT7ISkVxcWe4Wny/VEVJL7W+fmhg
ct2WBxXL+WwkANNzs8yYbhvS4prZMllBS5ppivDegV1B9oxnRhce+Cu0GFyBGI3K3tw7NOKi+QtI
w0227GYTJVUnLFFkOvdr4WZxQm1Dkw5GF7KB73NKlbXL21FdK7TPw5po9NBcuEv0vZycNBuOkKK4
uK1MGBEqcXPPaEefQPU/e4vOUGDLMn/36Xqjqo9rKhBncrtWqe9sq9OgH6OZkWEIDRs1n4zOEhoL
4lX9bbCGaFaSjZrzyna+ajeJVsuX6odicJLASilJqycAAtjaXt4p2ZLdhyh//GPSeOYESSfrCqqT
36NJFN7nA/zhMlNYkArucNIpX3y21BKaxqiej8D6c/DiUXaBS29TtWcvdoQiuM8jwBW7dawsuX7T
Xub5MYOEL6R86UXr4ZLrhNi9KMJ8IQvIS8vtvXED9+6nQkusm6Xba5baXkIVIgEG50f7pG0fhPV8
Sf2X/o3tgNn1Irv8Oy2Na3Rk4mUjdjvTDRkTKeLrXOW0JJjDoeyf+WEk69bXs5KFQeO1rB85CZZu
QSKnN2Eh4xc7qDw+r1KgAap3O05Uh/0XmqvRvR14RKkoz7v9w5lDoiRYTfKfkdP1trvYg7qD7bQ0
4ukStruHY2J3jpCTuPxkkFu9A4aGKE6t12YKF9ELxUpeU+I4DArmjVRwDqNC1yyTtQ1e/OjxGl4G
MBykKaEZt03A3Yk60gUsyd6xb57CM/G95FiEq7SLpXQBndnWhuwJOg3YdAbv+6GyX0iZCmo+ksjW
VlgScVE6UalnOIsnINL02Ki5WOo6kdVv07++sZ5V/qstEele189MaPD5phLO2QYZfadcsirwXcgd
8GhvkwwEOLkb17FIOxtsvQN/hbFGAYRXxDhjOOsEzVfwAqLnn6zFxYQyxa48p8UP+Jw7Lbh4X0Mz
OkhgOZy70/JI6XHQVBvDEhaCXqPOxSTpoJonlCaBec/C10uqoSkZEBRg0ZWGXLrIebl0/39GfwnW
/04yUa9OB3QLv4Lu8Z7Z5sb80ofKbmeP3qM/P3nCBcKFaN6w2kKsjF5fsMMn7mBByateIZ9HXY6R
VS0E5GOCBg5bBd3rTDX7ShzS+pZP9Gw+5RAWd6sP8kJzBLJWPRuxOIPLwbwOZKFHgRtTsUv4k4jX
++u4MD4DiOe3hdMEtemkYdH5/3rVvJW329ADn5tPdV1bIZKmsuN6gWtkCeD0dPYHmZq5tlTcyB7r
YYTgW4j1nWV7hkXSDn/Ub9yCfNQtApvb3d8pgUlidl1Zsu3nO003G19yaCC4WpvnbIsAS4H4BlE4
exAaU28JE85Hc6/EVgVhetbr0ES+HThEh8b4IK5AQVDY+6mx2w9py+qb84qwqlR30AyT10+RgsQ6
J5k3khULGBRVMBtN0qgyh0bF19tRhKnYkhXJL1+Qq6UXDrMlBGni9cGDO4+tu9gGWVRBIJbIsNty
EwKHNWCiiKBhTmwwx3hqJm5Kzouoi7X6Bt0XZPSWoUprZ1ZUsKON/nMs+szNlEm7GEN38gr0LEI4
J5ZILdkRrNEJaAFukA/29xohDzUL5+kY/sP94+mUExsWJT/efRReG0ct12fVtQB5gAN6Lm+QbtSV
SZvyX33DZwzXw4sA4+FKxkH9gem8ZHgEvtvvpH38f44+4Et4eMc5CZFK+PXxrDWlwXUjHAv9R66R
u/pYQ5ZtbzCCS9MrbLxVHR7iPVczR30YBTbhZ3YlY7H+ORzMfFg4NALVXWFfppYBKCif4/MGExkm
eNV8HClH6AHeRa3mU81Ah8YhdmpoLg/w1Uswy0TxXcaDkYCS/DFnc9puZtFRvkibWCpfEcxW+5Wi
AuQ4nJFxpZgxhmbYWejYMtUhI68yfq3e1vIaCC+fRxLYE/IMB1/DKhio53Eym2f02J9mvwAsCO5N
1FXs6iiLvPtBNSKkXcpENsfgS4xyhfDsSfMfHTPfDQuQ640yKG25oWiQO8ePeQAQRXhkPiYrxkvT
PElmUCeL08GOTE/uzRTRwyoyDetrpy4WJiE9rz7qZul+2hbZ2n46tkHbO/A1YehuSKWy3dfgpoJC
7F2auHsSXGmJ3n7QtGX7HyNPIH/kCyuX4AY7uaM7PtmCiAvI1/hfAVV9UMH8VyFTuanRfLnNattu
tmxZALPMsmkQ1eYEi7G9PTpoP9iyngfN9p+u0qDeRj0bW7f69HKXt2+OPCpq+RLkZUvyv+xHG+BP
BbCGKddSrTCVN/MvbbaAyUl1bec8256aXoJ6TchxVCGbWvOTBajdYcGr9OIftVHBtYW6Whj+oTw1
K6dXFLhBAGWdBWTGbtnULG/a4faiXQIs/RDmBT2sDELqwWB0oKd+jBzVjOf66La7JG5lPfv0IDai
Za1+EKDdLfNV19VJUP+q7zhHXwxMrsH6tiv7Zx/DlOlDpgj4k9FgusgL9FXNNhPR1NqKXyy5wdun
wroojzpiWjwz79EaghBPxVhWB2kbFftpAnqgS0RWERoNPAAf0W6LbehudNb7/1GvtmRbcEQgSLYR
1BuZDcXf+d8W1B4NkX96fLI/9Ixah0bLw2e2J7HpoH/j/BMGvH5mt2AO49lQLXPMPclMQep56BNJ
jQSk1/Fu1zElM7nVwIjnzrWJVUGD1gng/u1cD4ksfbZjFQ463UpJIC2ZdDz+Q2HjmG/sTsmPdscQ
5ucHfhnVgfJONJL3tP6+sQoJDcnOjVuC34J7epcOIwq9w2odNbyZpTBQ69C5Nlv55s2XWgDn9qvU
h7p5HVdvNrQpYNPifJR2EaO9tu1BmzbRyVOIbd6JWfEoIWXWW94yrOwQCvgJ2cARzLiDQvEGGnI0
X5yk92gQudxNFCInIbr27dbE+Isu234mKdW4bGmbPDCQy7VqCVAJIDBt1izjG9dUaMVPIOT4zJWq
sEWS0OAM1FJl8RCh/zv1hEPkpaYOzWYgkTeweC6RvQiT08hzrUyxAdOtqQQWEhVss74qZVNr5cuN
MsGiVPAadhGnfx4XPeopFR4pA6kt8Bx4bvplPXRAoOrgGX9mbhitzUz2R+8cpj8FctcHRJ0NZKZp
81bcabMmFFKiQgTrN4Q4jmNuOQ15cDGJB1KEDrUbNV5nbLUxQyd5nKIYy31MqTbAa5uNKgOCawjf
7Bhqg2j2HRbUdsY6WJmv5f/U4WEfaI2TWwYHvPT8mZV59Vk7XjOcHeSPpGmKo6VQoASTJzJtJYH8
BfoY3Px7ktp0bxroJfUf9aE683TbThSxVlJsxuwANR8q8Uzdm92v0HQE82TYYQjK1jzVxsaAhptu
Yy6NDTg7j2RmdJgCsBml/Nh7h6TvpPtD+qtyALjKoHF2kwX/0R1Q/lZdgmOaLdMUGayBeK6xKZjZ
qb0qtTs8pOUD0X+i/HWH0tZsABRH+vbIgBg3OR0Ukiwyan5juvgD+czFVpCnB3e9IDKPHEYzzTE6
IEZ4paAp5jsaONJ8xuiStBoWHM1oxxMTy/KzSq/K2/qNSbVQTz361+fsZO+73D+NTfWbga61XzMF
sIkVY8IJVJIVoS+cDgDrzOxOFQj+bl7aGaFAP5FEpPPdPCqh2Y1JdYV7CaLOnusa4Xu0zzzf+BWo
7GImfMqR7d6hLQ5ZRr15KvFTXPmDvgetk+bkhKOZsR/1A8jCLmwN4oybnUog5TWBWH+61uMHH4eC
W9LtkjkHP6UFVeZv5i03oMhFxnx87bKb6wFUw9MXBUixUriRSnzl0OlLidGanCIciw7SeSU8zYGS
9LESHIb3FC3j7OG168Jlt93t1P6yVFy8UEHAbGm06uFaTmHSK2VTIIdWHExdN/ZA2QircIeDPEA1
skJoD5YcbHdU8En+G6Usgkar+bTfZqEM8gOaHdm2WbP8u62k+kYgkQMnwtl41k4W5fIQw+89iXP+
28ssJJrzyNGorHtxIEPcNCmq7P0aNUr9AOrHq+z7kWcKV5T9CvakyLAb0YtfBnqvjkBX4PWvuBLc
mFkCyHwQgexyezhWA9AtiBGmb8+aw7Q/Plw0aWo6Aji3h1pIm5inEUJQottlwjcvoY+ohAACpJ3f
qVvtHxFoGMUh1hrzIXlrbg7KHp4PZpbmBxwJ57p2MXfQDpBM8MqjKHimT5hn9hrGYVyF5H1SB3lk
HKpEuanuMnwlDGYnPW/0GAsD93zI8gDzVuGuc19uL3x7RsvXZSWbJZFoUutl0SHV1kioeYh/Uwxx
g+Mn1Z7aVOhjv/4LcxWfI6ubleCDQyXVtyBHdebcrOPXpYerC7Yr/ncGpCrPCN1xOVy6r9tydFnS
Q+805gwKYtuPuKekQsaTWFGiJQ1QGHMuUcr0DMJ5aeTn/40IVEQ2MUJrduLznpCauiinAmReFGwB
1exEsdjmMF6K0vTcmh4usqe91Ram+v1MftMrgTUejl/QgLvO7Nv8Kd1FTBfQjwJntFdJ+/ucuY2D
ZErjk/L3TMtwp2k/tmnSg65h1XA93UOz0087rf2cAkZFdIt4eM6vjfcYcqEt2olWUpU5QxOjWNpC
413NMih01Au341n/+yc3CQLxYPfWJlDRkPdnqOBike0pJCdvHvA8crJvBT6Qm1nrcsRVwgXgvwVR
rOL8/rpoPyl6CdA/LS+/Y/1wwnHWB8sn3yjIW1y4F8h5WFlltq236FkgvTfDmFONpzC2coiFo2dz
NQCg7FT3SL9QQmrcguJP4kw7ky/xvRyvBW9dob5NgOnIQnV7sPIOEs9tBZrk9HEkaUeoD5RW25jG
Uw9tGz8quQXc4LgBmt4OBvWkKCYd7j+iloWbM/C5Pc8BzO6OETgkYk3Imd8+uE2HOZSO1NUmAncW
OgBo3fOUnWF/MsPNva/lImGsDqKPoVSqHfisqhtqGrWj12Mgl+X1GOBZoud+fwp1NctnF+FlqAJg
esCSAn2hu+SF2mprhVxS3HMRbkNiApQ5fcm9kMqwpwAOrpIgQG9FAzI05NtM73swqJkjNGQuLbMQ
p70dfkqnb8yHJRWebv52u8LZW/cBpr2RsckUGLLQDQ3l7oADXOW0uQa/a2cONiKbHqezcQetdLPR
nyYRMjP/0qH+EAX7gbczzQ7G9kuSgf3bwgPe6CvqGmETOLJTQnsC0THJlvDZKFAx22piyhkdFh8d
1XWbJeri+ReQ51CtfLf2GWudZyLy2iC7qCu4afTyh1wBiOc5l9Bq45u+eP675Y/JTPU5b4xdvIfA
uo3Nyf+AZP44OPXBREr21GRFUb0gtVD0AYK8oUHenyW4ro8nrFeNSgw/5EGVYh+716zOFAAXqjJR
+ZjJ8J0sqT6FMepHN0Hg79lEtv0xkaEH6T6jpx113gqEmLCQuOTZd5s0WQbmcUghXIKTeP9bkxPf
aPM4dDTBvDtg9flsfCQt+Wi2KI+E4lTqcTygVFXjnQcXriGrRfBLENEiGdDhVv8dctbwSiQDA8e9
5fXcOKjwShHvrLfNZi2E8xzn4vVWuGaHtNZca/OYsZV9vmdGLateCorA5mIyXFObMz03rlV3oEC4
XWbhFv7dJ0HPHIv8mjo68uMVAd2chl+jXXf+7chs6E9QaIXvEDhP8jF7hUCG0EiM+/7MEfmY+C0f
GO6j8nHA3t29ROtNYTqT8HzH/bFUJZnPEc/e0Ue5sHfVi55nhCeF2VWB4j57sQalprS206rU+CKD
Tp963q5KPrFV2jqu25FHG1IP3GJV/3ci+wPj2i4RnF8Lmment3b4huSoWtn+0OLP+LLxg8+tW9uv
NopznEFNR/EeOH/9BNw5aoZNqyl+urxxHCt79Ezru/5ywNe3uTg5N7lW1S8oHhjb3FrPUd/3fCV+
NNYq1QKs3oaIOhbzeQXlL9XDU/ih55+Ia2guFLDy+0e57iX9ZjXwHVXUJNYgC9gUn8XLKe4Kfodd
oYDLRkekLnYjrSoI2d63fRJtfBtGBsJRKJ9RH/cDP+zEHRZXZwJ4kgajv4jQywaI7NHkpJInIu7z
GFiW4LImWWjzTpzMEnUkMAk8+SIZfWE8Bg30MCX3oj9VkVjgvtkbifl3AMzp4J+smvik9ab7+aOY
Bwv1/dx2Kw6AxXKdLQqUtb8X6QQmdEF44GWXDoETCs4zLgsi6Fqqo1AgChHF+wIgaVzLp2lzGjw9
hvLtQ/GYAowr4XsO7dL1macNlaF3jZDn9n4jDH+wRX0+MsXiG4d8eD/b98Sol3c77zaI1CmDyqPE
UREkhtfTuPnFIDmFcciJbSdVM6qzzMRFOdyIKmAFvYX3/MnE4/B7OtGx7/R7afWmy3Nm7TQEhdP5
oNo5AuEdLceMixXt5whgbQzm9u0EO+9LTrpR1Ns8etk/8WyrWjdZhmzFUGlY3HRuvJ7swMgpVIw2
KoT87zrXACtt3KD3FBu9VBy5ThER8C89/6KHrB3AnWlq/TbjgWapxSl3s1gIKh8tZhGupi4ou8IM
vFVmar1NZCYt7cD1U31wzUf7Y8QQL6d7QiKygdCLVKDMkfhuPQmc6WweVMSHcyO0zIsYnfxS7VET
XNk/UpEpEqM7H60eT1RxF+BAwJm5W6S8Wq5iewSkKly8pbaWPkwxLCtoX9CpY2KYMV50dtw9q4Ru
USw3X1wDTh4U4ebe1Ss44PyspVw8EyQuzfKo/oX3IbIWiUYO9JJNwVJda05W7NkBQo7ygla5LbhS
cCwebCVGu1AhVdE7s1nRJMo6YaOlEWz1HXXyePmmMFHd2cN/drMThzeVKwA1O01GYX98OFKBlefB
PYXy/GXVbI0YT7JkobQTKVqocmkutUhBg09Dyg+2k1HDga+v/JCHG6F78CBzBp9RFbkJfCNWmaxf
tcd8GO1LbS+RfKbROBbMyua7loT3ICbQduFwjPLVP92Zcyq6d8S2ILiYR1WQ38pMk7/4fIeK1JLl
M8t5Zt0ed1njcrNO9gYnLHxCgHhLCoNSHHCuX4S0BNjhGEvCMUiGJd5wKmM3oz+lFVN9D1oQNevI
kJ7wyPbOFLYBi39W38E3lfo6bb032eWfjDiTbbnbq33U+9pVv4KYgrGDp8oKZ7zRW1S1yrlzBYLt
wQt8YF6vsoBgUomufE5pO6FP/w38kQCwnehhgICpntmgxRzeeUtjMyESpYLlpRSBavjVj2BR8aIz
/3aSxBX/VN4qOE3118qssTRfAw4+PUtMbOsiUT8O2IZ2ltd2/SZ6PiO49p6eVDxS9YrK6OiwEfmP
TEBIJKgsgpISElSeWfdfnqVB+98M4SQprF/ax23FODpu95vMhjp18g26abhpGw/SOXyP34XTVW7H
CgbRFgPR4TcdtWVHem4kzeOxRyB6jwU8FL7Ys1C7B5hHR+GHZxnWOMrSsVde9IHi+G1vC9AYAq4K
y7kb2zhbpXEQhKablyo6KQC3pUFBf6ehbk2fbhk8ZoFe8KwOu8DmDcPAdONG7OdPhSam43djsoYZ
WfRx87gkhHVAIUFxtratyn59kqcejTvmkE2y8ZVjF6so8QrHUd+zEMktA4YUYuHxUBAoaOwU7DvW
Mf5toW8v+WTlqrXOggWsiZMDAEwVE6GOQJl7urD3Hrr2M0XH8P9bsU8cWFKiHwThwKF9hklF2wBp
W60QnpKG3mV8CLPv9v2xM83FI7uMmzLdWPw1OiBhyuYdjiUOs0qYuz34CeyErxpXf5tlz6xxN5vD
yGY4vIV1rk3/t2ofBXHkA3T4m6eYy0tnIGokMT8+mUZEWzeMiuAAwFgv/ad6B0GZG8W54AgeBBfD
dvce/czJQNiYmB4bj4jMV/+ppXEtrq7Qn42Sl2CkceNU6hlL+phnJYRDL668t/+rAwtUkH3Jomi2
T3qVhI1P0ErCnvHJJ2NFXWisAE+CvV6NEhduf4HPi1h9r2S1x5N9nOoYaxMySP0go5tY+tZ7p4cP
W04J3WnaYahDTgK7trynk5BatLk/HOzC/x75L96DhfkxTjwKkM471iQ4OuvkvCn1xoZKch76mnn1
OhUigluqqfJ5lBfeatBDn6hlKpawnXx5USnN3a2/GUQMsHXV9fRQbewzrfVa29QADjwsXQDmWLXG
cBqkKU2psfFmvIZ98KxXgAtUgH1ZGlXfHug3uTh6uBascmwnIDRi8ShEm4dmHoe8G1QnO7ySBdXT
O4wAEYTjnsp1YetHGQ69cuazK+oXwacuSlgMEwkr7MlK5my/iis5behTRR9VA8MozYcKBVT43D5B
EBXcx9mNIn2JP8Mmbr0jTrjAIE6N14uCRPrvJYxcx6ApB9UcxZqu3lNI4dxzmhcoYj5BN91dfGDr
/7RXXXCNIytKP29VtzqvL/jECM6ok2n2qZRhmEJT8ngoIYe8Jsigolu29I4kBe0UdaHS3LHBEwJK
LV/colQ+myQA8X8C5Y38t5cyxtW1L5VtFPaUkCMMgoowDfP6h0hN2UWn6QnCskuyx2Pc9+PkSp/k
uGpgfgnB92gNoeCcRT227O8uaEvOrSt3OpUJ7ciu3abd8XZ7dSlPdrdK/uxhAZQGXd/R52Zuku0p
ccEgJTPg9mIogbtVBuuJDL+op8TBlMroe49yEeYx+497fbwdYg/iI8xrArAokfwWejvV5S9CePVz
U8+Z3NRIAl1FKZMc6AraSnS4i5lOHKKqy5Js32rm8j1jpncjjUJVEfGC/7+C11VqZBtilEYDId+8
EoqCC45Sz3Bw3fsGWykhZkf81sVV0dyi8hsT1Cw3Dzk8uWU9KbBdM8glek1yn/uNVTDTRPrFYSyu
4cQW/v+DwUB5be6+B8XSNRqZdmvIalGERafFN4JYGM2w6nxeeuOGZHNieB+/ouy4y9crUfjmzuHU
fci57hVr4Sc5m9ekLiCtuz7fF6B2az8yb5U/rLJM3Jbq5pGT9G64TzTnHAYZDT8uQG81WZuT9SFV
ZxrBKng0VQ/dT1KSV9dRf4ozoUrCPUpUYXs5B3naNpWfcsvcm1qjmknAbGpyfOv3GOrThyybUjKP
Tsm0yYrDKwt/kAst1qSn5Bw1z23QTtn2azlHEClq7EnUN4+g4+G3hSMymwlWzetGuYICQwJCoRxk
BHV1cYLX5ogKvRVCSQtG7l+Qful7hcmvQ08YSMNmCJnnrV7fSn0glWS2ixvZVfJEpmhx83vumYr6
eBM771I/QjVp6atsxyVePpWZZzR64RAkAAmACcg7th8+KFJDyICCdYO4oFzLPBgBhJukHjQNNZbs
uQ34+LKjY0MbHcmpDxy9DHqwopUwmajyDPjDXIABzpHc1DA3f8zXxvBFKpGTjjC6BrS4wWjVWmO+
LDPTwtXkOoRbx5XdiUgsgyELuCWRm0UYwWYcImAFkAceLcCSJfl4kmsOHty4mhIaxFaz5mq8IhkX
oGPB+LvUqy5mCOdDBK7ci5syF/zrUfSuCiv9+jnwPvvMFDR0JaCxtHj+VjY2llD/zlydFO8dx2NB
my7X/tVtKh4u6bPVfqqs94jSK5dWjCvRlezkSkQ00mzmut3sNi5MWU0AV/2+3LABl57J1YRumawr
HFE3H96Q3L4BlvawzpP6S/8wjQAkfLs30HI1H7pGSzOIGcJypWWuFvkm6JYy5TDK2GwT2onQmjtF
Xo0ab7LQQ3i7EUCoKS4ZwEQu/hKZA2Wfp++gsGsGMnT38vyDVvdNE/qc30gU8ur5UFKAcRHfaSZJ
ZoP7dQar3Vr6IblVAKv60dO3j9VwvQmnxc4MS9/h9WdPzAgv3bCTpxDhZqJ+PoemP79gNj9WjJo0
OImTvvrzJtyyNDfQeq8k1IniR+e/ZhSnmKzd6T5qIaYjxk4cDWFAAmRGsEEVIgbKm5jcNg48g8HS
5u4dBSDvd3566yFJ4mE5tEUiHGuY4WJtyzIPOKbz8itzbMfdQHPZsJ7DJMTrZZesH9a+joTdKpJb
D4h2yIGfRgGIw3p/+TsicgHR5nIwy95cO9ft9F0GTydtY+kYRlQVB04BMp9MOLevf/k4YqPMflIT
jIz++MPrTrMvd0UuAUaxVQY8/MY2CrlMSR4YkzR5t+/5sRMMuBNs9oLQtetaEGmrv5SS8hLuF5gv
Zux4vFban+SFvbxm4yDC95bUIupQ0bIlUSKfgHiDeayT5GWoAD8T17MzhAbh9NRj9wgzkIKamR05
cVP0j0a9y/dvOCS3T+8LCnMBE7DjQr18cqLTgc0KngYDO8WzkY0x2WYNEi0PdrJGbCHLbNZO4NzL
UeZYpdiEj4hD9CFPLJRk+jfHFtdejYKuM05OqMgqmrxNwjpj+VfErt04Msx/sPnaD5Zx1OUxnw98
GJUa/0MHPZE/E8Qz64tPSg4DssvbKKGZqmbi5U1phcMaOfn2OPePoiE61euwo7KWgoykNxxhaReU
QtYHFo7c+a5urzAdxDsDY8JwB2I4WHobpa24aoWy441Nc6gLbgqJwGWenpxBLtUSdgumZmpa29WY
AU+j1vhCrJCHg1aJZoI5gx5mYDeQck5yjJbPQa+rqp4Q/AKeCnyKc16kiJhmbT3wtrtcCm6CTlU6
/7u4+dWfOZuEXFKHBmklhKAsV34IggAGwN+JH0xk5qbAHvctJ4L6/h+wcNAhdCn1ieGm83LTBGgU
C+1D2+oNmLVDh3r3DSPwmkxngyfjkK2RNt+wMH8L/2h6Z8+AFgVL1+owAaSdohf0b6Pc+TI+rAdX
vEY/Foy5iavAzQt8UemyYw5/mheSeWw5sFsbsVMP3c+AsoHc5jkp3X4Cg7BYktPz8bc3tUMsdies
KoKZAsreJhCO/amDv3gDpRyM6YpN/XPxdOlh/z1Z96qT/o9S8iMrBcRPusWRKEJFV2D9/FaosamQ
hp6PGaseAk6NBecFokYtsKd4e7Vii+0nPZiAJU14Fn/g2zJ6nCBKrCg2Bh7/kz7eCc6hEVv/5m93
HM3ZTFxs+QyHg17N6YL0y6JBK1a6IucmltFV/Cgk80HShqXVB0qp6m+jyqRCbTyE4xVyCZTM0bUM
O1sKyD1g8yXjx0cQNUprI9Y2HVADLLk3OpX6AiOBqO57nkb5iYTi1kXWu7jcT4t6mJeu5bCmE9vb
GIH7e/ayHNt0Qp60KdS62J0CmwFZzpUO3eHiMXhOlF7uI9f4WAnsyyxU6fgYMmV3Ut3clHwUCum/
xktbKW+Cds38TCadrLREBHW+BfKLmjlOvIglE0S+UcVSu1TZAkRsf77Ci9aQ67B8EAN81gmg+84B
yQm5e5aGjrNbhfu9L6k+3+zHaKIbs42zE1VTTmSnCgOiyWPHh0g8gG6nk4TrtaFFV2Ls43zps61b
dpIsn6AoB8agDhzl2O9CqIG7JGAzVTd0A6A269NQuYyy+jvusIsJ9sVYW7lslhM79pWoaZezqJne
Ip8AqcfOkGg5IfuvVGhCODuz6aFRX7RNt4WfWC9zh9qswfNCIoU4QZcyETHKrx/4DGqCtfliTQEI
UwCH+h5GRsZs/cyoABNYn0a7GAU2NYy69Sx7oWjr4XgKiP+wvWn+0QUK9ypxXAzaR2aPWnA0WXdo
jxdZYlm9V/hxKfI53PPr+jMU2AgEh/3h2eIopbqdF1m9yKAI2fjKTC590TEtDflPwPORSXERYV8+
T2LHogbDqYQExVzts5maYyoKPcpujUgMk7jMsFoQ2p3pQeZYOIoAf5g3G3OdHPMDabL9B5wfTXqj
owB3EimRZMC5RR0SIAsR9b6gQ+mRGsZP5M/UEIa7B/CZrXoiaMdsTwT7kNB6js1HrEz7GnwdzlG0
+V4nn2GkU63zhUUU+t7/JPCbdIswl5OwvnpLPHJaIdAyh6CrQK1LDyC2czUjX2WznYf7uT3b1zv6
NmsK5t71ZRxQYFHt21QCGVjczAP792lv0K0JU0l/SBymLgdvaOcRz3AekC0l7TF+zkK/FAiOkjmv
PZYGh7mgdpRoXengLjmYOCRfX/EBGKg2oWq35bI31Gb9uUpVD5JVVVdZNH6fe9lqUIwHvU/gjkg9
5QCtxV8ypCUw8/via32YcQMTTfc0OUKggYbAiz7pxdZBpUeHER0XwmwkrZHhaFGAr9lhRcQQ3Grk
PxbRjWIJn4ZbvWtkhfsme7wgUV77nLc+zfa4cDiPZ86q2QcfAwv6s2EMH546EK4yWxc4yhry5Arp
VOSe90rvO4cM6Z+FpnajAyZV8VjrrHGxMXenNnuh5VcY8VqtTN+aW5EgOhFGDhwOS2UraoDCzOc5
syg3dQ7Z9iNSxLStKjBnmTR3+W34Y0OEnLDayCFJALRdfI/+b0OMRYrFvC9SZS53AdbMTg59PiDM
h+olNsq0G8JDycOO6e5HxzjbDerOPaK12aRF71awmzO1l1e9Rft1xiacdM3/XPzHYPJ7zvy/Rx4l
VYsJwVhkMVU6TXd1Wl/Vm62sXL62Sz4qZcg/975ptwaxW0r6XukHy6pEEfpEXPqn6917rK5uGQ0u
K5WrDbmNKWKJisqxm0tSfkgjId0Ju7RQkBvOtcY35vUVQKV6QTMLV5eAFKWzX6ht6Ked5/ipd/eH
rHHLBNuYD35bCwx+DY6Z1xnn4+zTAA1qeY/YXn+z/AYIZM6YjmWqsz9n+QRU1oJ+dJrIJD+l0BH1
u/GeRk69el11Nh7x8V4IJKCnN58GReJ+Xw7yB2ifuB2lFuAcQmmhwkvy9TfZDRsRcfZIq3MLamZ7
rI8Cq7f68BUFyg2+PK+uRTVIuCo2Xjb1gTI9wi+i7w3SFkkw0ajS/jn2gy/Xnko8b25h17Yj936g
CvNWthA9COMRQKVapKvjz+Fr0ZmpQHo13p5OUy9vE/7CnalqzQdRFwZ+4Sp3WeWVJ7uJYu+B49sw
/wfu4WINo/7p6YskfAbQbn4JQNRGW7dD84dVfMxoYKXb0Bb6h3Xi2ZD0vxBIPzTvnI/wDEf94HQg
K8YZo7Jqm0HTNim3yzyVOlw+UW3/h9COeTTo5D3s9TXNTJ5GRSPg7oUE8b/RptaeNMAAnFRA7SnQ
Q3ZkPlKMMT6vAmBwkp8LRKoNESuozNJR8XYg2KU4MdxZuEc0b/kIbKkBp+5kMZ/LxkdzB0rj+2R8
AeiOk7+ZrGI2RqD54xzA1PsTnDCyBtQUubdKfnMuQ8axjXRC1Y+l+QP6kZBfiFBGHf8F751QOS7c
0kZvgreFylW3Zq8RIBoXDVrqMMRF07MJUpmTWKD3JX7dLJXFGs65neJAu8DIIU38wqquPvGnF54c
hAr/0Kaq297DH3/rDGID3MjGRZ8uK/WEocRKrRpgGJ5gvtufemG2cJt1NKNW7WYVdDGmfJityteN
2+3Cqhxr5DAEZULW5PNRKCm2pCRQDv6O73x3HSILPrYNEGrIbj+6GwKNtvq3OFrXfzSUXp941mGB
3NVULzIHktw9TkOJKI3bfeFwoxm6VvuD9MvAFklH6BHp5uSw+RA+yCNJ4He44em+j6uZo4nr7u77
uq87cvOjweEz7Yl+JZOnAZatAGQAzm14SJ9pAKjC6+U3guPn1TdtjkI1H5/2TqwEmTd5RBJ1W+4+
XVEhkRRNGU2EPiiGv6dhFM5FgwWOhAwrGoSIO89oecnvQ0aiY0Lllh+IzwNMm6lq2Dnywa7ApLfs
BVt+JjHvSA4Ag3Q004VBrnDHeuRwtAWoSwwdHQhJgaxf2Cdgd3ug9RjFVMZeE3g7iXe7Lu/cG/OA
WjAztgVRgE/iwbZghAySqH53HjgrLKRyzc47OlXDrh0bLRnroRAW2sdDpRilA1Lbv5VopxDEUWe0
a0XSeWpZFOXONrXA2x5kX4GEvkuBmj6H2IPpRVLHyP6q9sMBSyBuD9P/lzZDArFXhuEFnXXhS9yS
asNijOf4uasS2ET4VpdnnrH8eAibWzlYglPD94GaqhRBerGuiDB3JoI69fWB0dlYgJiJUHeIFPYZ
JgV6WbwJ6r/NnyYggfj9BkCfk4HAmXs+ndSK+8/2NezqxmxqpU5ex7ZT6His+jM1EwNuBQRXil+4
jhJYWKrCEaNwblvNzKwcj1LRnRY9IrqEPwx4icA97B5IomjkFDUEz0Dd1iXUn8W+c3TZaDPTYCuL
miMiI0kZOocWRg+Pkqq/c0EAx2XGa9XQdHci7rjPkowcKB9tqPMes80Cy3Tg8Z1esS/Svgmfds/+
KhlxhRMVvDcv3WIVOJZc97U8nU6YelPItWSbXxdEqVesL4VQc8k7qGMukaD3aHZsRR8IwpnU6uv/
tj10tVBMmX0fbuLZ84vBim2LFzJOh3ScpDh2DAWZ84STeXbkKQ4Q0do4z7V98j/yQAiHYlMtLkbW
b1xgVl8+vEQeYmPDJHq6xK8u+dO3g9tYXTSl2ZwR5vb7oGwySU9+yNMS+c7920fvokA1G1pzPj7M
XZIYRo0vSOT8BdnMTGTKMgHeNG60V0FZGeT5Xro+l0/g80Mza/ZExAQMmld5Bxe0SPWbShoiX+XE
ZOPzl0uv6ts8uV2IUzAg2EVP6IOXZZV9+eX2otoTqNpgmeWmRjyz6134hPbXmBb9rwP5Xu82QHS4
wAR6whbCEBNEjIqhVstQO5+0FnukQPsY34Q1gCOas0o8mF6H1a318yvSqkjgaAG61ZuXBR9LgPj8
GYxONmiBDDAi0nMmNd5fQ3n7tB0lqaFHhNjpOCzi9o4apiXhs6q5M9VcTpFjY+HjTxerqNwvXSrX
Bp5aH0j04fL6QPrhahRm4xsxSFcbLF+ECCTDnfdTE17fzZnW+ilkNLN52oql6FRLxKDrSOcPcPK1
hID8Q1iUcd6U/zs5j9BEFkiqj436MlxnXTfC8IoAvHSsaTDDlVaHfRv3XSN6LuoB6pe/wigbnxht
I6GOV7pT1gjyLOuJtJiR7euteKSXnAojJnFLb55qYwuhaE4dmS3KlP0BXIazfk9MN20ROum+cmIP
eLPGY9YC5+ioj8ZsUyISd14mbB8JZ/uioHQnjPqorqRwSpCQ+N9W2f4RS5Y8qtPWD0J+uWWESupM
x9jokITthwPxXWcnXWKgdt4lL1HwDrkelfo5MmXJVu9FXqnoyY1wBRPcu46YVbU2w7cgp4uSQSaS
GTqQw5dlb5NYrPnNXxWirMsgPiOqYLJIBNcMyuMZD1lxYd27rQhKHL1vUrvtRN8gGM8Vpt+Wbaj4
TLkPO9l5BG9/VAPDnp47z/uNGO5WhwTGYKb7AKDAJdhD8XEumS8meWBnpGZ3c/14cAA/R4F66HMs
YBWB8sKRQDsYh5xZXXjg6WOgkGDK0idKHcDiE8DiH58egz7AJYv6R09xsxB2RWQ+YW1Dw704V6k7
gD81NzByaMEU+YUCkmCtfYUk7ZBuiKBtuVxrg6esbD1Fjf3gLNEW0+xQgoumKYuDzJ2iZ8s9ZZnf
Se7h/FgQAo1J69oOwi4mhBmjq9pYQO9GQdvq/6yRYoBdxDuaEa+X/JEJ+JxszONLd/f7hlOFYR+4
61xmuDidby2JEbjCv5vEUKxMYeWesJuCekIT35U8FgeutXD+dbr7+pbdnfYzb/VMtvgvESuVCFhK
OZswy/hTXdTiQZDMukVHj3mk78KArX5tE0WInAIRVoX8ZpUkNlEh7otA1jYZRMqV4nUURI/XlSye
UFlIvqNSQYV9Svi5Vmbx9V6DyAqekj+yBFKH+dstRelU8bjBWKQPcdkioct+Xmp+cO9jVnAIKd9M
TIn8dF8AFn3cRkuecIP0BpI//m9T0QRdl5PyHAMh74lgJqvXoNV5YejyI+FLRjf4AHdJcEkoGGVq
6CEqVRphIp1/af7Oe5G/PBtlOj0m/irBqPZVfS43lyHcEfyEAgpxkXIbUAYfEyS/X+T9MUSYNZzO
PHLGlRqURrs0ITHMFS6iTQbLo/1yj2pDwlqYc5E144t1MDo5wq0CVdhEID7Ujord4OY/5lOnJiLx
prvpK9NhB17olmeYRJPT+RbsX8iBgfi0uqZq6fEG8sje597wW0QCcR8IWaeoARkvrAooRhvTsVJy
U+m847uqRg/SNrg7E7XVN7tvl53JqxOGiZGeRsSTvnGQRwulv4ig2YcE1GmyqZUHm0WGNcKeG9X+
XatGlOMrfPX/e1jx/qajXIS7DLLS5IHdZLz0QfTE32bDMqwxJce2kFMFhIHHS0SAeOvL6atREAqe
79rQExupw+EuRdhqyioPTRvoxh8th0MHUa9Z7Smk23YMdqmt1HrteeKv6+X+zlMt653ug5rkDLQb
RINM9sGo8cnXJ+EIumj/Y/yyB11SI3DRiHrI3FUQJ1gyLzxRj+UuqLzNavgiaAAtvcdDXft6Utd3
JlPvs2cu+7pc48RTUG5EJ8aQqQ8R1ct5HYgGqtSNs6yGaHC5dz+yQA8QKvwuHvoYoQN7ang70a02
xGbeOx5HxWAA5EJeQ8LwrhxHMMQJrOD7KhpVAEI4y1mIxR1Tcvy+cH/JwTMU3zOPkWDqSclWPh/i
zAkhcYn3yDdf2SaKIuC6Y3qWl1GQvMUcG9Rb6AGodm1ZEaYdapicz9Xr66B+fkJr7ytw8ZXwbL5e
U5B6GdhLtharItqUXxpIatS9S91ML2Na/jJ8JKrcsLb2x0XD1cMk5IZUQOtOPEKS0PR8MI5xDqiM
shoUDxGkeaQanbI/GETwCVtwhH2TtuQpSXqZ8RqRvZpnzr6hfvPTTToCTqdSIDhpQn+ruzZ/vggQ
DG6YJgSwpfnwjqacgACl3XS6kyDpTXe7PB72wcOvKqp71F309D3b7054vQZMhk6hXpEEubRIlHms
KIFz4xrDzNNklk1U0uJysrJs6Evu2sWsLhTi/YJaywDnQUHYEjW1cAKUT4/RZ6hZFhzJZ8Yw1PU3
Us+LIqp57AUMWQ93imumQCGGmrha0gY9jbiGt5ed4OJol6wWH5i2V7dmy0xKv5mOL6CgGe4sMAWc
CVBPu1XgHgzuxASPYsin/Gq6zFXEkYrlj+jog3DLfUW1ohtiCkDGAgYiyJXklBqPI/5oz03c5mDj
PE2lnI1m4eCMmKE7HtFsEzkevzaMiax00yPRy1QCrRd3hdrg2VF85YHAnu3kRBWmLaigrbodXXPq
b8ty6E1n/J8xonnStQxFUowBsjTskFDm2eO+Oxy+72c/Ztlphr0ujTRRp5G3HzL1Lk4vrrosqo88
yeze2OC82lfnszNAlJcKL2jmRzbwEVVKiIIuDOk0UmaLZ5QPpjppgCWbhXwaMs351Wnws9MvVwxh
aSo89VF2MpTs6ns717+IFNXSlYYZ4Ci2zkv5iM4GrG5+1lfNdon9EWi3ygtNSnwNo+Jb+RxFHUx3
9/FMgNDFkkRqtgO/cSbP9dLM00O1iTVXexRk2a7r3oUq1y7/nBpDLDLdygrhzqd+Ie/Hh//cdjGu
z1pKNrJ82FE70S3p1TL5mHEyqAWQoN1aYnpe6IrFJ7Cybif+BJqN8OVyD9vP71EFuqUzsRyU7P26
zCaA10+Xna68cueil953/sPxWQbPkH6sclPsq6jR1YYiPAFY1z61B9gGJVL4aq0N9VhbL/dFFHsC
WDLOtgejteEsCZl2+NCHLxA+DV6T5Zbj8BADvF3YNyIX5DQnX3a2lr/iFQg71VPOiNKULLEFB4gB
TmN+uwKmrzE7USqczIbUl4KK6kJtSOjR0qoFWL2AHeylmIl67lSJ7OKOw5wLjMYizc9nfryfc22c
L3q7uNMKRFCuQpH7tLWk2VD3Yq7wcY5t4k5GjrxfINKXRmRpUlQjUsEyrg2CQH/PzmzLrPcj0Y7d
jcAu9+olI38XNo8Yx6cCx6sAiKaZhhtEt7Ii/RLOUK0Y0715RURDCryrZ3EUSA8yuR7QfvfGWKqR
aOHsGYDZS0euE2I8F6UdMms06TNUZDLoKYmEEvzs7azPezYdXfU1mbDu+9211oU6wnYMC3d6Q5UP
Lb6c1h5VN2YcU3jXXFuWIrWqInURRPYepLklit8suGZn1ITfegozlOgw0R5RdEnm8ZHTpG8/a4rh
WskZyC/CuNLKnl5EIXdulYbhgaT2RLZ/+tr1FWGkcbs1PIqjbXYqLpExYpQ6e1OszC8zYO8w5nDf
qpcL6ciw5HeMhSkw1TumS2KmNb7In0LrqBIfZgLtDRvWjgGLT7TEQstFyyAnfZ2q99LsJx6dhACC
RtBLFvWGyuWYn49uzbrgjulF7pPTSL9JWC4SyDSbEwmytAByL4EMfgTkiJ6KKc4fC8KNuRkqUk0d
cK4OK+MFmxx4gO/YGybMLdGcnxQSV4yDLtWQnnU3C3kf1j7hVPbb3GlOuoDI/X37lEejjaoBMdBC
1NaOdqmaac/BzPci17IpHzPNQJMriIfeCLkfBuIigQzZXahJfQkPPeSMm7YBH2O87jKaLJyPfVzW
Cb0fiOQVXuwznNdYC9nTU+alF1bsIqqBlqs0EBcydrMHwxS8Lh7r+jqKvIX32NSYuPhO9F7RojTT
YSeHj9oWtjLLMqO5xcxezqM77t0fKuKIgX4oDnQG06RGNiiRLi3MrslQ+1nnwRw7CcS484K1XlyZ
JfG6gWC1cXE12h4RtcE3SokTF2/G0Ccvt0+I+hzntx3UBOSnOWh2fDO8zMLx7lMcjY/PNf63BoyQ
cMmlcjlyLVIKkaEMIA5v+xWhaA058wenzFsu1Fa5VbFdwRnKKZe1lShiOgXemh/qCfWpM3KM2b+p
3SKiAfP6XEs/FfX6HIL1Hln0PyxvMJ6mORZk8TVX5Eo5X3P94ZQt2sGKa2sp/8bFYYVK/11viK9/
eZcee/1dd62xiBW8ZAlhqHTK6gJnuICxDYWscFnJeqqQletub5pWktUr3/wnpzo1VBWyVkrIF5T+
GSwQuT8Md1kOt6BqxqlwSCJIRpuLrlSct0ag1lZxFM0dMJmdIH7c8kRye7VxaNKEvAx2W1OBF/QD
VGycwuT++DWkTZJ4DfL4eCE2KsezCWlC+K4GS5qet/WhDN6th3l4Z1ulYG5f9HT2wBAW/tSN7oAI
DDpZ0t6hY0wfcIGEmF6wYjb94VTsENsGVHjjkRXPM92ok/9R2wUgqcs1aJ3xDClcI74DuekdsH4y
hvdIqPYtvdpP+o7tRUjpHMwCribBfEnIAkU73D1TipAHQas5zjH3Z0iwThKQqlBBq935Y4D43m+N
wZ1smP1gUpertJkQA5yR1cPdASaCMpwvhb2cvilFVyP2iplMy3Zra/v12QJhCzS5uZgm+fS6wEdh
cQXH1Wr6cYtA/B7W4Tyg1t0S/An1Zzou0LMVXBiaUHO4WdUOsi2H7L+U+GtrwOEjxZx9zzyC0cj+
BMCl4a4djqFBlSd16bVzjq8q0ebwye1jt0e3yCBJ/LOUKmHL0CaAv084/cAzvJ5YdPMikDu3/F1w
1b2vR9EDFMhn4tbqAQzVj34/hixDpxAvLxXHgwEW8/h2QayKShMli5GA+d6VU1KdB15m14y5u1jI
OTwA8kc/qeEL/qRqSVIzgjiotJAxLuqPElzmuomI2agD5uspOR2TCQldCF+PK1DxSsUMnzruBAxI
F2ASb3/3lgaOXXRjiXKBYodF3MZ9LVFh+NhVTXGxTUcyUv8ue2njGZYubOFwXkm8tj3dGCVlm7BB
NKlx10+8t9sW9jZ/KHOG9fkX+/bW2ovnx111qwZ9XoP/6QNbkmCoP7+lc20qsI65Fjt0+omzR5DT
lGEo59qsCB2XxwC95d8qUrXWYkicdbhAHf1yeYGXA6F40Y9J6mrTJpGNrXaT4sCehSpX8q6UD9NG
f+znFRtrSLr7ste+0KdIHXtIl7OERyrAmreMG7yfm/mc5yIh5lF9+kNEg88VKauxDQhPZkH2Pvgt
oaF0AdPHEr1fwDfRfcwJ4wLHS+Ov9xxSE1LBkKzG7lqMs1+iidnrwPyimW/zx3DrVn/K3a15Mh5F
+UPu6uStOD858Fo+1cARwextcAL8OBrEGfBRVJLRS8UDh1M8kDm/W0fdYzYz/TSgbZOdQRRZ7RoG
amMm68hCU9ySYEFGxuV+TD6JP9gCJGzlbjVIaImlONATZhzWEErP2O8W48jx0SJ0z1gAOAnd2H4X
lPCjNzc0N+ku+yvwt15akUD0+vC7BRmIF5eBgoE07tpesWONtwQhdigd/OPiBOvYkWFP4wus8e/u
u0mO1Z7cl+L3OStHmOgA9JHIHHNvJEPoyGAsdC6uRuvpMB9TeGRbcIqI0ByeGmJhHrOpNC6PMOIv
wWAyLVWx9Qvjvu9rpQDKnhM5y9MEw/XRfsuFgV/BRKL88//8MPpzIMwicEvHyCkXr2G+iuRZyta3
mjQoUaBQGc3cOygjEpNf5ATG5m2xz9z+pTQTS7BPre1n4TfHkOrkCg1sYQ1M2AKtdbz+9dtlL9+B
1q6oh3Eo87Rw5ijUCsSyix0ELqEIH1xRP7kNDkIC6HUoJ5fqA4ErfUKjlP9JCWjF0HGnd+HsipDW
FMdE5dpGh4g89DP/TpVV2u6/he9G0PBpkt2lnqO5UZKQYaq58TRseVBZoWTszzYXqa/soB/9FwGF
6E68JQFpUlh0VUqLRMd44PldLe4unFZaqQVXsv/kgd80SW7qbzPDR7ZUj/P8OwYnFh1upNNnuSTA
dmXs/A+I+k+evwVxjLe/CTKuhGEQ4+Rk0ZSumqVmwZd19zeKhBl9j/RI2yjZs50ahsT7sAa/pkk/
dU6sdlz3cWwuFwZkkVoA8P/SBskup+IRlFNiBGzy8peaRms1XHIWt7Z0EW1RQvvMf0RxDdxc6GKP
2+RLOTP27XgSwUvyPp3nt2EN7e0yiX8NtHbwR+QBHK94xTDKuPxaWa/lCAO2vctHoEWXFqxiQVVj
9uLklYNDTKvby6ZZRHuakOoHcmBvO7nazzfbRd6UOfXjPXzWqpI7Xa0laqNX0geJDMIgPwHc/Sa6
gLcF27ltgxljZKtGYs6wz5zdM5L3HL+BdSTF6HduzAbpmrUSDZLUiZ+SZh/W0oDcPd7bDfvRdGIh
AncEhCi/UjYClLx1DeG9yi6NflvPao4B8Ge5SkmqomWEQMLOz1a0FoH5I6qLwUyyJgWkQRU5PYde
KhaOf31bM3K1hazLRUDgfcZOUbAv8/AdrvSAblPsgRU//UkzvlG0WdVLhcRQr7ppeMZjigW+sXhq
efLEdmy5CwB+QUPU/SxN77S6rDZfOUx5jdMWyhava39EnGeoCIUJBIMuHj8uL4onmvCEgfxDx3FH
PetQ2me1bD5OH+k0E0qdKih2QRokX0BrrF7jUQ64YUPCT4tL+IgF7ZqhF57SVaTYXlUQ+25jNGG1
4TsSkzi+8808IGucOcDEAgxSAobXRQoEplK+cFr1ZpdxA9DRKT5jpB0x8UJwWNEvjtAT0BDvtK1N
bkb5DN+MT0k9+kveolk/tvujGw659HanJ2Ovt35WfyTJM0NfaJArdj0qYoLBTzjAQtRjnga5tjjC
v9GCFYpALrFlFvUx+xcd9DaeiHtmx8hUZ8uVOKhzrwfSuy7wUnDFNCw6u8+7vwvM8UzhxrcvGzB5
P1JeRArRsDkixCvUD1WjQhqqu+S30w3l04vo4EmVV5QvrS/w7GZMYxQ1u8crUPq8Wr3ChhMxLW1p
p97z/EwCAjBq4szOGBmuD4nVRmSdNVW48ldvyNKAoGgRdZm0LL6jQr2UHfUa7aKRzbDDDloWY1Th
5Xm9+N3cHL+lm2K7gSHi5u1av+jt4ehXqW4Ta+AYYS6gDFvDUql6wi0G56t+2zw+SzRuQy3lc1wo
44CWII2+8V9tvirEXuzP0IBQI87V9uArj5/httK3p7rBfK6cBksSV9tJnj3v+1i5CE+ZGEl6XdHI
VsXdHVTuCallqAp4Sz7cBVSR9+HzBc2djj5Oe7l6lI1+UgEhbgQGj2spRztt47d0UU5JdbUHiKjn
jtaB21pE6NFH/v3lYCiIle8uPJe+0dccFeHN0+7aBArHgwmhIrf45CvHw6CY8A5y3hKbybPRFbLM
DSK7WFQwSXOv3cIaCP0y2OHstIvCYoOkaLliZHNy8JPV+5YlmVI3xbWobo8EEEDW6sc7Xzfm31zx
Srhx06MY9ELw42G1bSYpGWRqbNXsTAquG6YeqHjQaseMevtXPKBeGHlpm9Iw3gdxVMz+tYOyyevS
iWe78HiwUiWQ+4rThdJc7hu2OuTwcwzqP4VlMXaaHYqOQm65x9RSQbcIaKK5qIoA3CN1lMvCXuyg
ge5xhtxAskeH/j4m1ADz/pWB2ygS4zZlSoJTIUWI31MLI0SWXUpmX728lAo5EzE5nsC8D+qILRrL
dj1bB7kXsAw0z8JYlMnzbjYvo9Mqf3wnTtViSZvL1KxSRZK86TPNguh295J/TXEDLiqxnLA3ZDiw
7jTDUn/KcLZylXi+Ou+aAXrJ9CwrMW6wSIcMCMPog+5uPpHEV9i5gixndQByu60payR03414aCXJ
u3GhvqMlDNV+gPkCUxDzYt+zdreHNPhHv4uuCnlEp+BloBZVHgc89P2q9cumpaMvOOMmVDZGgDPF
OLwj4p1vKKIVWHAxODFV90fEr/oHmQ0Bxyv5CNM3vH4+L8JiTEFDvQFGJeejAiBnToLYKUbW4TWM
i7W1XhU++SZ0WIP1LK6zEZwGEzEunGQ1Xe9JbFEQxMcu2rtR0Uu4kYF4ugjt8ke+6QblLAWMLwMH
ae4AZnVaIMTJon0MET/mysT+odsRXC9qYgUYGFlzPlqOceBxipjO7Sa9LAIlUfRVUJcRsncYz7zT
qJGU6hgb3KQ2GLsRazVXKn1rd2le2KO4UWRxMrU6xPfqT43ca7MF/KRJtVcLFnCUWymCHe8GTe7W
cLfvdRS8EcM1gbWnHfHARWjXLEitGGS+IfWWr5yHodNBmwX33m3+3rdbDkvcbhP3J31l3H6Mwfka
OkN/rl6DvhK7k1/vWhptokoa3Gv7Pt5yBg0JwQ3bOL08Mq+ZLf2P3xIbYZ1gCm1a+Ggbg2CYcrVa
i8r0y61FIbR3L/a7zeSUsj8BRZLFvZ2dEwN/SBAP2eZoetQUjrK3zZa2t2NNnVCIdolFB3kXms62
w9Wh0dbNOnkfUinUV2iP1rR5VPvr2Bewd+HVfGImIQXrh4tI431GP4ztB60OadYLp1+zpRtMuxKB
Oe+j8kyVj49ztlXUSqUVzKX4KQoZL3JpTTUYS4xlWo5NrY1JXPGWeczjx6nXexeCxDGNfaUCGMee
mUBqhLPzrEoFbTEzMv63CSwec4U0A0ooif5vMxqpJjU5L5tGeFKYpyFzNaFXcLR9P5emYydFBeCs
wzhgk4D4J6KBXfUO5+yyeBjfibVxQdfep/j4RO7wHf4QtLpNUK2U9goyJwq7SnSakQudaH4hB8pA
rI+zeXoSsk2MeQSHSnwQDw+BL8GtP54GQQkPDKwTfD6+xe3SP/0IOTA2ZwPRrvLrf49DDGunfK4Y
uGB1uLh7j2flB+EtKE/rZuBd4QXU6xMRTUW73uuXl/eX5fqljhlSgWRw309yRxOGdgQJUG7FNNkF
wKszGnGWfighVzmRTiIlPqdvRE7ksLSjjzLFE/UVUiMSabAx7hAcEGOplndigl0XYVDy0GGUNftE
CxJfxdff9kLUP90RZCudQckdQyaDrJp/XmqaR8swUbItbE12wdmtK/C+bYe5JNFSWliW9Iu5OCdx
IIFdVWJHe0XV693Pccg6gOVoCVtMj76RMjCMQnay4dtgXVEiOv+WT8Jl58t9bJhpBTYYThdSZnxH
xGFQWpO+eE+xi79cfs0wfne1NsRLk/jqitA7gIo01vO54AsamZVz1qr/9oDeedMgoghkW+DkCusb
7iW03z78TygULGUhP6R5Ezyhf5iKIqtTNNiDiEv9BcihNbWkV+NHl3fNQtDg/VSB2DoycOyvURj5
wUB+Ij/NBFTJcFmDVE9dF3+CG5nF+IQve9Wq8uaaeDs2onu1d6BMSJ31ijmpgu2itR9fft1pRfVT
97NFRQzlX8zeDvV64mEzGRTkMzaDqAQ/hRdZrC9OiNFuAoAKMMOqJmjmMzr7yseW/r+PMZRh//Qw
PhGNkDx3RYJQUPMGOy2wgPdnZYl4dRUwCBEsRa6xBxRmVJqxTqJsxd+XTMT+ff/Vfhkw69eKDVcN
rf+JYzwcy56WHwruzyH4MKMzsNj+Nc07hJuTzvP0wvI5HWvgli6sUllS7ZUUOK7l+1Fys1rYpytq
dYcxWE1fofH8DAAzeG46fUO3x3wLWA0+xw3r8hFys3ftOjtBqea+QdlJ4b3ReOv7+3aIc86bHXDH
bJSn6b6cDvpXwx8R3dn75JbGF2kB2UjQ/OGQesxaEKZaViu1Atrw3I+bBIUPcy+264l4qfu93s0G
W4c/dMQyvyG+sSJE0yNrf8ipIi4NqHbxg2ASWaSPs0kyrCtwCkFYvIjRqPG+ib9YkSFtu6UR2qJg
u/2ifH75ccRUWbFqFbwwzB5PonUM8BdGwHsJ6B2UMm6Od2ujOedSO//Kdo6PvxhNnTWaUut9NA74
bm0yUR4n0rj27dbFg59wzjzdBySHyD+QSntK4pB2e3Qo/MnXGKprD40qRzN9zHeWuaN6MtMzsH7q
VxFQ/mcnb5lbpmrd36bcobFzyJaADq/1VyjVAsO56YEf8GZVP5WMAAee5Y2H7E1ACcnmZtsvQmsq
HCakp2Z4gzCUNgMXFQzqF6ab8eaJ6SfIDEf1liYm+In+nbmAq7x+hoabxyDntUwVZ6Y5A8ZDtpFx
bj7//MHtiqyEKuI16zFLhBeGZaFuWQdEG3VQlOddPTi8aGJ2SeKItyGHqQk+sgnJYh6UpBXNXudI
OMuOaA7BU/hBnTv1CoWRGO/FyWkms5e0vziqOM+YEVVPw144waXiUksB0o2ywMrD/RIYfVxLTnY8
kGdp4X7z8QDeoxrmzUYZJsfwBY/GdyBjc6FFFBCd8K2vsIOrLtRmWE4i9p1OTKukIaVPv37xqgPc
F/7aKMZhdhfcBthLHw0hP6FAm0dyJRkvvVcjvFLQqfIHW7vYnPm1g42TjO8XgmQostB2AeooFonr
qWhf1SK62ltVrXqlfkQpQHpMWHG07Hw77y8vFVTmerhwjVHRqnKMZJRHzVxinNZ+5jN3ILxFVN6A
ZZxd2t0AKDmYh+WgpZ8VPsB1gD6CXU/WSgN8EylFe379xRZRMLkxtJlugySBcSpJHrijR9tfCey7
lGisyLmL5FRxcuVDpDwp3T+z4DYuH9Nz4OXUF5Fxf4aZZEXufSh8jK3ylh46UJO30g8Y4MR6XJ73
uRIx5HFJk8w8ya334PYByQVChQdrv0aa6uZO3wHEy6NwEgUtLA+ulgRRuVjka2WF+8QG8tzKKo49
d4hrDIjJ4Ci4GW1AQnzMjqiNYKTa3y+J3kUOUT4o2vhlFZZL8ejT9Df3Q9NRElzqfGL5YyQFbLsT
FGCFuDVBAM4N1ron8Cdg7tpJE7VoRFcOLw+FXOb3MbhJ5X3VWFYaOSvhIAMorqAQ/o8SjnyVac7H
8/iP0OxjY1pMsT92dvPfX/ECqTIdGhmFBVcb3GY81UHpogoa/RE/EGrIgE9r9cGIj+/zX3ZkEoor
lYtkkYfIVTm8Bn2mb9sMOF0/EF6tXuHdNdWBanMOsf2Z3e619k+ZlFG1Mt3owvto5ADPhzziNBne
3iyfEt4LY/hA9/gE8hfHYM8B1Baw8Ny5KvSNX27HUfjwBjTTAOB18v3Q3ezaIpxRXu0vrdnoR+I6
QJoLZplTA8RKBAg4pSrLKcgrwG/3M+pYAC4q0V5/Tc90CVl/u8fJYaDsc6NZRpxd0pmsxlOklSXg
MVLogtNhOo3kiguwOQXbY33PgJ2lc/XTYXVHe9eQCXuTyWZN88mvCie3bSGSWlrJvvBBWdNnGe7D
zyffzq9TIcje7HQxPrBxQPOdYmncNCyNzxScsPDzCkzCrt2fYnLh9ztRRpr6Lt82Oru33c8pyYS6
q1FxQeUvUNc2C1GIjC9Nuz53Vb2C2EFVEzB+dv+lYYDr4MBGSZEcT23UU8DXq20WmPqc3cBNocXT
9npRaqK0P9d11e2cn03cc8TVwNeTnDDFm4HE2bbrC942M4J7X2gD8PR8CTMV92MCDWT9DZ9HBrIk
cfDc0I9d4LgqPc3yU4A52qyLEvLZPmyJguj2WzY+iJp+9KEmLz0Cxa5c0yCoQrISd4lowGI16cwC
LV75lLaonTrbobwbCyuZhmSaix/Jqv/6VMccldSY3XUuass6AjmhDUrLhWNsAZT710L+5gBRTBTL
FK+Q+IWulbHuJeD5Ey4LwVZiwn8odrawLTQN7FUCYYQnAvCklNgfapddEiquZL+kBF5YTPN8l3Yh
JnNU32b00V/N5TqR95UTijHyTjDZs4m9s7KGHbutAsmORiFy+PVg1YYCO5/qX7md4fQBWSwNjXfY
mWU6u7rnyLKIsICohS6f3lULmPXJ4pTSorn6AvMCYL920d7vY9FWj4S2IZhAuL6JfZapm/eX/u5x
DNRVnyJUWEh3DiMYkpKYNaJ5oGZPGh9la0gIROOSmDgzJPu1BQcxf25j+7uMggBOUgJ0wPJTz+cy
DuJElT8RbXW4Y4pJvYQrRh/0yMmOl4NLABHRu/l5YF7nrjfKOc01RcZq3sqKigezKLKQdgfl+hL4
C+S67Rf4BAdXRSWFscwUPr6ILQLEJ1KflhwHM80k6y8umJ4X6caRCiLX0USb43HuSC3qhs96unV9
5GfDv34Q2p+o2dL/yo9oGOh3+h1+N1OKXNKMhTwjZqu94PjOjrwrDYk1/2M82ezbyHWqRJH/IasR
fBaB/LLUvrV2SHSmNgceBi5WcwO06DFpUNDTdLRPe9OfFizwAYILBKZXtpfxA+97/h7uWqYiJlcV
xNcZbtfSztDeXqxRxE+PgGzj58VByZs53aW7LjklLAQPF697g4Ek1gdNpDxJVxKGLhs3P7PxUtXh
G7SuX2mFqpnuOt2fCNQvVb13+VGbfl4Q19aJXVwOOkwnv1O2zqd61g4rWiZeszEipe70GItaMNml
Xp+TMg6/CzXFWn/+NZnigJb3GkhyhBcT5TuQLTd86TBohWRBKixhtjxyMizlqtxdwkFYxxTwzPiu
06Ecmleyp/RmXSvTjXE1Q1mNBcLazcJgMZytxOktgao0KNHBqjvTFD1vtBNmcpo+bYLrG6d7D5pe
Q5iPdA3XWtLe07cj744alihdNewD4qezUX4sL6QzNpkBXw+UAdfCjTybPjRB9bppE+f5GSgVW2ng
1YtxE8Azav5rrlyxvQVOfxdFc6qC5Xk4QOIWQtHDWqrX/187IXRkwwLMjsbWSBMqeZ1O0TT9THbE
rLX4dXgmrnbRt2/EKlts8sNrxsdLPETlkpB9+qqgbEo16oIxBdGL5RlVxKqNSLqPZUFLf0Kn9m/M
NRg0i9Y541XmM9gnFbegqU2qPS1jUdkKjjkfH3w3dWiN56n0NHdm8bsB6m74hE9qVURf0DIK8uAw
oWcHX5An1FXX91K3PJlVn/0FnWwSR1YWCxfGqLLtGG8oXOP8rPFZYGawpdK0fbmpVRlavXybESwv
k+GO7KyOafs9tAWmh97mmZ9uFCnKE4YPAPHu+hceGYTlTvZrkD7JC2wyShYLYUZECoe2peh2eIiR
YrETaiLOFTlQdahHuSF0+lzz8FED6aU/f5Mplw9zQ4vqKzJn9lJv/dBlmfJtLLec+nEXJgUdz9CZ
xbFj1UjuhIOQ3xvcJ77+BHD2UPwE8isqWNBZ0cRCvMdQFUZOFcCBgZxUC572pft+mFN2zCOLCSbl
6f8jPjzZPKaj5Plgzc3Raer00s7UOaxdKnBY5GgYvPRZab3meK/xFlj4sw3Z+1/cIZMz6wK2iRuc
CqR2lHoNh6i/ybMn0QEBh++6U8LBmJeZ2hl0XHqAYmlBfKca63P+L8FC0VbXbu7hsIiOMoRTrJgi
Zm6cUOBGCIMy0rHuKaXew+JEeYbcKwEZIikGDUbjPrvQhI2BDHFxHMmTjZnWK2KoeIHqdl2w6H1E
yJEdgxjyFu4DTY3f39XOZQXKFFNduvXoqheF70of2Fs6MSCsXnFiGMS5HEhIXpgYZi/hSf6GKLCj
G9Qc/Pkcexj92R//QBZwNrWIHk7jOqdKsqvK3o4DyEDrLWMK0U8UWUtzDEKAaoFYFJDIBIZ+U4/C
6jx0KVIOOedYnJNOui11bZaT/u+VqCWk5pVAFbiq2gspbg9YZEEvK0+QaD6ktVGU1PK/kuB7T38z
ehq4fWt3mjrBO4EbwuTSddSPjafBDoLOFWNM1C6hJcctUzYx4ozMhr4G1wqbA1mGBrBT+JD8LhUQ
OCLEkxpfuQngmduaehIZXrIQQ/yon8F5yl4hDCHOWEULjTVdPjBVQLtKxiQyW/DPSsu8y4JpmctS
/1cPERPH7IfJz1ukyVxAMC4orr01cf1hI/Jb6QS8Uu68YxAykO4Bh6UoP3NcLtvyhWaKwJO08jJr
C4/m+XdXOBEp07tbgFCUOkSjISTaycZgNoedb5J/UIVw9fMr+Ngd0bL6miu3syMf68rVj9B37r47
/pkGEpH8bly3syq284LhXIYMVQIyrhw3YaaNFTVi1BLYG9ls5mdkfETZFZ1GrgKCqrY4chu9viun
Izh7mek8O7gyhpSJGHPtV8WEca6GwtDZGRT+F9Er9E1TfTKTd7wLCzcA1zi5qGHT/wwabw8qKNK9
qYHl3h0XAaSL+BIczxqETkwL+lQ+xIgHeHTUKw3ZpwNHJ/7iKjMGFfDuSP4wHcz9LB/Z2MOQ1OrO
xo4rt72hisx6mTMPoDODzuFTADNiP9noFxHku+51ghP2yC/vfRK56yLCAQ3NmSNg2MbKDQHqWOuq
jGmE/yPZULoTwtVQlAt/r3o+dWzYhFcMT9HNqJ0+uEHUiksfEL94Nd5OfXnLLQTPSUfBtK7fDipe
NU0Bh8D8s8yuAP8+itDxT32t8TqU0ZfooKbrDNLY+jIZTkLkhzm+iXzwpDBWzpfP/xuPexwuHd/E
yi4QNvTzpOhLgi5dOG8tHwokPxuEYNF3A3mfXRy0BvYfszbJf2umOFK7ohWM886lAoxvZ+uoz9Aw
oOjRE+bi8bbpQTzrpsehZPo6EGunkwFAB2oCgt1b1QQfiUuzbEruYBwf9cgWtfLO09SA9vxXQcOf
IQDRR+wXviVH9rMHNrPgjcs7T3v93zbtOvFmsWkeMqAbuAXz2cYtJlIxnsez4SMJEcmc8IZt5usA
z8ZxDIIBdN0gsWBxp2hjOsphWDnHm0qlTzD4hqA0ezZvbitxKQU3BGZwKOe97XHQs3SI92pk/EUI
X+0L+RfWmIuL8cACMWFKazoS3wkS/GlmeFDhlrnNU0bmwd5ftE/XbDLA6S+0oIiMTfMW1k8KNepn
v+G5l0RGX8Cwo6Obs25d4NqNGvWmh7gfYQwOaEjRSTWdadyA0L712mYfSJwUdqfZh5vERyAasbvH
YMgnV6GFH+atOClEq3+liiw4H3jtsJU5oV2ibJJNSXuQ9ZNLM6trq/NCp3QjPuYZZXDGLZRb5i7p
Apb7KfwXXmLmmN2FRr9zbKtDm9PY/xUEMuRFh1+KQVcCqrR8/ybJmz0s9/MI3qpsaIZNtBiqHFLb
E+v+Yd9OPS4k+cGdmfo9yXqgYblB5RGV9kLQyjFB2b5lGRnZCvm3nqmbgmc1WqasEhtk9+7VmXei
2D7HS4vzkS26aKgbmTDSmjSNzj1i6qrcSfOx5eoWscmkFs7hv7UpLNmiR/079DspH9XTH9/a3uDx
cN7mUAhNrCDl5R1UopmnAgmQyIFkyQ8ZLlxJ2YUHWVTBue6xJAWMi2H7pCENLofIua8RBTSQZd/l
2q2s5xr97eKyR3aR/Ap3OAGMGsqamH4rHi5VPMpQdo2qrwTt50SPodaHDFrHpMQEjYbttnNaia2m
dHw3yNCLzb9FZHCyiHideyw3sXrODnrnPwGfWpOqh1obWMNBSN42YFTr+DzZhpkpSf1udUBfUXmK
j3Xa4QA8WPsAtvEO5gYf+DW+icMyQpqHmKwrDQDU52fda/nd4L16tyomjudwxMd3p1X076J90aan
8CXfj1A7n5RLk3chhSR2Sl1U1qSarX035WegHBQAUDGHwzCwLwRSzPY2R2jYJoGccTpsWskIGgiY
02Xx0bLYk4lgeli5gYbyB1Dfex4XikiEe/XH+cXSk3r+J7p1TcsGh8TGd3jSnFZSbFqW7u0O+Fn2
fagAEEv3IGxFUIaM7FT6+a0hQxad6KsIK9NaHQmjRtp4wnxFrUEIAN3En/ZeH/bSOt3x1xBTsis+
Qz1me8sZxggeldV3dY5+046wUBDTLfMLWW70Icx0GfPxL6H6UOOQvH5+wEOU4gfacuYrVyehYenm
la+b4G+2sYVuwvKHbindc4IgyZunJcF8PFfItqwhx1xvjmRWIUMq2hUGZENRajxWd+g0YAbyfBzC
57oJdHkg8ut0Egw8ZCuitWiFsr6IFBOpKcXzkL+y9s8JglWQPtP0q8iikbP4mhn6sXIH0QC2KeeW
unk/G2SvzD0oYmeiE6BpAgJ/KJOm1b/deh50zTKEoKerWlrUNiv4I2n+cTmhI/Sn4PvfifiD+Rf/
7MzpuCc6ePFudwjt/KLu42xWIBO/MRH77q/IvuohqOTO/lvKwyd7ipCWKo2EDnwqgu+TT/VNDLZ3
yEg/ViZyafsUX4h7uxsMAltMKB6yBO5sDrEYK+UAFUTHuMaWaP1I8drIxSwTSSax9peS2J+BvYwa
IETwDJqxMuwefDvVdOpLjzpxU+1axL5uSzlGurvKEX1ejzVbmQxQDWsjNUHjW741BCRFP0PqAt3R
3S/z9mVakeiOAcuXug3SduCjg5ddlzd4BKQvMSXg4NE24Z6cmX8UJ/CGYT2t8ougijLgkRN3dqSK
M2w6brx0hzenqAqPwjmXO+w709sEx7jsMHypmAKE6ZSQ5XKvGh65HZ4s5Eg7grDgdL+Nfi8sg6Uv
10PvVHr2xqnFUBApQUD3QhAmlo4GlUl8q0BkYqDLkEpqZ/BMSxA86HxG/y+sDYMf/4kJCVnUXwkL
qhn39eLycCsv6RLC6RrIBNiiiE63RGOlC7lhdujp8az+3eVV75/ov2hl8UI7v1IDPdab8F2TELa5
L9BgKed1n6UpzX3y6qDX1fTaOGWpJh6UWwqoLDVEA20aEH0msf9S50ytnjJ2rxXRm+MDtBgx6ixe
Lsc5kIy7YTslwEXV2G4t8+bUbTk593E6ws+7Lw8jumNi+lQakggy2y7hev8CAdx8Rm3T3P92rVg0
wSwmwrotwL99pTloqt2gXyur2E+KJzR10nqXBkNVYiuzae9Ogyum5eeTnlcQV1wZmndx3WLulHgI
dUwFpCf76K7TjsmSWtSRsJDHgd1LM1s7qgxLUrKb7dKmurQcmhoQqGxkEatXuvGgL+ddRhIm2SIC
C78aqiUa5r29vaF7FUPeOQ0+RXIb1sOTTFvZ12kbxXaTsG37zLAK/g0xTwAgwaJSmp1IxuppDYxE
fEUOBJd/DsXKOCHQSEu8LjOH9OfOb3y8ELDJ3iRpE8Q2SeQ+uUDjdYP1HwZuLCWBo3rU6sRb+KUb
oHm3N/5L3xcl5a/++2WE5GQIfbT+cTiVWuiAxtIOd4cmCe/54ziP6hRbVlxJcD3/fVK+3uA/xYgC
DmRlXO3GzJfoTfRWl5vMJH0nfEXWeFYWuN6MfZG5/xQHI2odkL38ViCX3SQ3dRQMTz+H7hrdaAcv
GG6mVEVZyW0n7WG/C91U9SXiuYj6o/4p/s/sNq+000+e8PqzdEzQ2XOg8NQ+ep/yUN8aTQz0aOVM
bAT1hX+ZcWXqMoWkFN57List1cQSMAE7TLDyPogMz1cq8u3guA221cANsvVqgY5c42xfNU49dWtk
/mOGxOf00BQyraRdZt1Ve9t9hKZXR3M/OYan+GCQawf+xQ0S4bQk9GxZxrATmbvVhBuMfDOZcV+Z
4BP19U8Gv4k5o0rtWZg0SATpA/WWg5viKPkOQ9xHuOZfUevmol+CQHYac+VqrgpymJvouPhQ2NNI
NexVvy2oiEWXVdfXLryaeWSMuXe659+tGSouznhX8afnR66oLSKkBPSc7L9t3NaRIcTMiYc94BPq
gNk0Y348UBNh8ETiTziSWMovvEnTYEK70sbAirpRFlp+G+oBdJ03D3dSKHvx1ZxzJS0tWvrNr2LN
EBQyLjnrI+uq3kCA30O1uAPS6v5x5Yd75pHWP4lq637E7oEuuho0qjeFbFWirKf0XT7uisLzIQqM
E9xhssgqxpbhDo7SSYAd+sMvBPH1TFFPaUoqer0GGQ4LKbSwD5vg4shpf7fTLqcqds4Zw192iKg1
PhXNOvvjgHY0mOOITQAPyj37CJx9aw/tkyTkWPQYME4svrV9X3Qrpcvgq4+DlOn78guD2ZMTrS5Q
2FIy2Po4cQUlZ5jQiDb2hsSeHKfH6Atz32yb+k4/VF0GEkbGmhRoaI8lvqlddYCaftHBjq/Hk3oE
yZjpubQiK+Lj/bnhd8vj3GrzgJ8JJ+x/C9ths0PmpKeqKIGT+lQxm0SEGxYyVOYmciJmaD/4TMEs
JcXMG5z4E708CZKuZTpVS56waKmRB6SjDm/umG9wxt//joGdrpX2PTR8NOviqBfayT5HTHWWxEix
HKDDiim3ibc+A1aEibKuMky2Ac/MyFwjbf4izxm8JT2MI2fbFQz9FSpyVvkRAK4FCMOI7YZPXEJs
yIY8EXw0DXHK0IlQs5V9VQ0n8fu3A7Zwg2IkKm6VHz1lTdvxq1lZn9B41b4OzOFU7nKcarg1FbU6
8z3J+XYmFGEE1TxBV0iWoy8qgDZ2uQHrWwFKQ7sE6btBrKpdWiITj0COj91EhKXSXUH1aq9zQAD6
cSnfMQHI2RbpibWbNbrtRv45sEpyL6udRrFG89Nj6T0t5lBlA0eU5HOKBEJWpBMHBHyz7p29oelw
EAoJzJlFMf/x2DYphKtSaNXqOX208ImZYT0xyr4XdUNY1LDn4VwyyLvpIfTOqerqAI7OJvj76qCG
7ovw89QE3cDaiKxfh+NbWzJ6Bz11Ureb7P0QYvnrS7q1wODexGhv5ExeRwXmz2EtsXbb2VtZDnpT
fe74ETgFunT58pUhxnSKJkpiamRoI69zf5gbVp8MhozQpCMEQUUM0vjmQGKreSXA1WEQ2prX1UqY
Vbvo7tjcyijeWg7Sn/K/2GxVY+BgBodj/IR4NJV3DSfyTrtBBdwEMPSkuUS8y+kvdPXIvq+r2YDQ
tLJE+6FF0vbFYfCxekozyY9vyBzsgplvh+/4HqmsUkVFzQhxDev+pII3y/2dkt9+/4FLOL+dpxyb
YRCccstv8z4ZvZZpXs7miOyA/8u5YA8U5b+BZqkdvj5RJ8S5m3815vc/KengtuCw5lQgUQhhXALz
Osc4oMmHTNJDK1PkaJzHNXAY/lASDd4x3pSM9d8mLJM1coNKrZ667xiqBJEIRJeeFibQiWIbGhBi
394VoQ0iwv9lhM/jFmyFCawFAetBvyZetGHBlCZ8DR7+9QXexMd5DfGBSZlpQMD+B5nOJBzVmh1Z
j+R1Jlyg5IbPvEFqA8joFfxl4sW1QnfYtHIbh2NUnFSRFKrSf0IT7KTs6g1D/z9nNBZGv9dXBXeZ
fdvwinRWwvnoAgfprvrtVq72B1jWrRUIMxxWU1sQW+Uw2t9HUFOTyvaiilov2GoKtRjZZGiUzIF5
+8yJQpX3TmOvhigv9C4oiDL3st0LarZen51TAX468rQ0fhukniuzUyfHIrN0SHK+WPdUmDXk9172
ZBJYdQoLG2TYG6SDrsEjWx5fmFZSFYxagAdL9DjS1g2BjCAipr71iOnmpgzkA41QLNtKIvWoVkks
UWVsJerDkdpsTWAE9af7q7sAqoK+7Fe5Y/uxjubq4+hydgxsFhiLmFZFRCF7sWVZMU8K6TuzIbcD
KMjnS194bGJmjDX7eu62/I4rGvXdh4tP6olNIzTjqAyHwRQUOsqvL4pgr2kfhNLxYB67hh2+L73p
yvNn5gNq4LRDiYil6m6u74IW15Kzyl/hLPT82epzxkzHN8TMh/0odQ1rd5Uj9TYNTVW9QYltSeK1
kSrKJcPXBYZ0X2YjxR3B6Jrf4n+7e2EWUu0OxTe6baa3QEQZ8+GTBPhLrKEBz9Ps02eCALjbi8kh
ntbZybsbCI0fa8a/GH3oT1OislMZhr3wrbyl9TQ9+QXqk+cGS94AUObjIuaRr7GlUjp3GMeZ3fW0
GyZtkx1QAzkSM6ItioTJDISn1Xt1vaHoPcdvTg1Lg2lWSEOmKXd2esuYrsstccQf8ckpO/b/ZRjT
P8vmqCP9vMOkSjmBZNDr9A+tpv6Uk900piEVYfEtX9g+d9cUrrb641hCIpBHQSZ+jaK2/Tzq1QAd
3a6zbvMoS8xw3E0reaxr9oxnSLUILfvFe4YMEhucRgf6m2mBG5NiYUagDxBk9yLDv1KNWo7PR0Oe
Ul0p+gDKBlSyGddT6Fnad7R4OGlMLeh7x89NbZNT3EVy+JdqTj7XqS6BVN0Ef1oojH0jQG4jRVPO
5t1rv7SCtS7YKb5+htEJPsfo8rVN0SLA12440bhIJfb6/DdH75BErlx4E4iOZwer+dthnjhDxePv
rzYF6vEl3IWmCeI/Fl/zn6vIgqIydiFi+3W1OumSp8czR2/vx07FAPdBBx7GhWVnSMTQo3x2JaV2
QK1U5qyuStAqC/G1qMPyeLyEskBpVtUA0oJwLBag5MuP9VFUT/k3vXL+C0Fs1OP0/s2glnIaVQXl
JXHOG39/rq7itLfp5JHHzIt1TPmwO0DQ3nEy/ek3RKKM/PY2G0CdKr1ek/Oa92aa6DKAsQkfWzQg
X3iNw4d6z9kTQ6aZj4fyZRqY7bIw3Yy/CaJvlEDi2UiIpdZPEIBaKw8h6UB0vpDrtFzz4kH/XK69
VAg/JJ5svuRAszXxUel3sDQ+GMbqBDIUZUHOvaRq/FfIOuYIlHDvjUdg5+NuIQHteYPNnXLGP51t
cEzhSKDo+G4lGvB41vc2wqH+8gDc9ZhQUvoiKnYFlZ5RkDft5tTFuywp/5zLVM37OuFaUs8uj5pd
QF3KognqJ0dyfC6zWNjkOorLOD3Na+SySCDqqNG8AMoKObX/0VHl+nhjhEdmX6ZpjHTsQm3L2BfA
50gTJTW9wnbyvZfiEpt8YSYOzRq081jdQ6YzF7RSTtKsyVb2wyNqgCV8TCr517hzdaGkKsY2rces
1HEx888AFGf0fPcBNuArvZZEgmyWxkMqkXnRNgSaD1s5dGe90qkck697UIcPKAaWK+V0daYLgDKr
ogEZ6bszgk97ZmKsFLrxCqLDSqRdUOn0rh9lofeQGKyend1pvnEFdizYFSLWgHDAJWOWU4XRbzZY
rk+w2fc8yr2Xqgiw8moKDJtY6poiHzkjt0kDn9SZtIeWmA/GwxPB06xuDos0Xk8+Uy1RHuyzaYzO
3Ur2uPT9jubmybPDA9eRLbEvzn6LxyxI5jO71RYJMvj+G5yvuWTowtQVDZUTj7AnjNSAVRmnAOGX
/KVdiuFZZIxHkPlvWvCcbITRdizS3KuJcaWtCDoUibXZkSLQ36v0ajwsSIX0/b7QRCM1ZgFO+KgD
i/77qtcaYbYMLgyEjoQsnT/9phRGrPip0is8Yft5e/9pRO1n2YQTeNwOXWq9cF07k00ShQ21BRiL
+y7vOJLDj63dk6k5ZoeLBCOrXClkiWdIY5FKE6Ai19PeYrqyQIfr6v72G1h+GQfPPEFc5N3Ieq1N
8/gmPJxLqHzQpAfGp1ahZJiszXJYyACGca14fuDTE+mX0hkYkZU1H+2rHc/5CBC28X0MsjqbEB1v
txsPUOoBb7acUNMMEvd1Z+qnu4pPVXHXjssgDQPMFdWPCtNa1M09TXgbCT+IVtyE79NRKzHJyuXq
YfuVR5dlXuGdtmAuaEkJfso7tHr/98x1Jks5SU/gqDAqphs0LOPLMPVC0mMu5maDeRZu1YvwNVsq
bG6bvtT21tPkKysKPelY//jF+btE3h4d+5nRO93xplkXjJx3TyS9WIT6UxzXuoNp0fX6iIMMCke2
KlYTyak9p/rRpElnHgA7Cjm+JPgUL3Wa++1+vKHxVP81trT+TosHIehyeBSa+MXOMkjZjQvBkjJO
HQ5szsPFg7okYu07mjSPDuykOF73yaCDeJHCBO8S6/rPLi/szXr0aNqHDQLEkgypHwNdQ5MMEbkJ
+msD7u2VRJLEYINw0WS8k4e6ROXBC/IRGE90Tt047QaZBm/AGYQPTvfphAj1NAveAB27RnbwxPZo
hC/PvARxL1Int7/6CnKR8UjYv8UW07BlyZ9NcJhLtNBc957ADS5hpC2hCEw0m34lOfmhvPzMAZla
UnFx7LOO2fMCRxpNPK7thpEGf+PJpP/pSWIWSJsE0IHdpFBTemz4hhpSEKD5qdjHhabDMCd3dWqM
GIReCbonEt0TqfVsl+YHYUDWHn9aomkc4DwUh1qPqDgvWnvRSfVAg18DeY8GLKQ7YLRHAmN/ThJm
tUuW3aJsjTguF06cTLqFL8mAlz2mjg44yl7ZIh8KDCS84hTfuo8RiVy5nU7YkIrnMCCcZesnWggc
AGwpV3GpwCxEqA3MyIacBhRlMjVkVCXgYCv13nag3AJ7fSaeT3nfNfuDQ6+9k/6E8xl/W38k6IH6
DprJ7yk0ipnpMpm2bIRjz+veW3XaD9IxXKQZE8MiD311q7tioAsTXnbq8Kdch7+9c4D/N3PDYo0r
3nlCbAzXCUBss4HEZLBk9WLKAJeLXMCNyMnTU682dGNyZdZIxOGsCCU1Aoi6IlZecLfXbUJKwK6N
uI28epzsUOgRMDnCDlN9Czb5LC5nN8h3Ju7RSkVWa2o2Ded8kXFGZPS8N/C0pOfgAcdPwfcSJiEY
aDf4ezeRjqKwDCWx8oPHAJdPY3LmVu0IbBxckvAU8czKy2Zzpx98dOXO9eFe3Wq8gSEIagHksXry
x4PvfkXtZokJAtkcOM+J4b6hmbUuUi1fsU0jwjoA1zSMPu2B1ZYjFmuhovYmlBmFUpujvKPRmzVa
4cnQUia5snMpG9HsqenQ9pzUAhHUfUORIUTWYjypiCUpVs0NNimbSC0zSRk/mmYgyLAJ0NVvTldb
+STGqQPsPTwHhbTDi0LCn73DTui15bLhw1mVYKe5oFalYIlme6Z3SKGnikH5PmPUo4uMTPFLvppn
miI9RdQQhAcLMbZvrk6YHPQu9KkQgUlLYqFW4feHkZC3ZfDIW5jMa6RT4gywvEPBaPZKPy1c2xxW
rNszbqclt5m7BklyTWpGpAIVVx9EoiaDE0FToLXXoChV+LigxL0lzqeD4AWmOKwdbkTUCbm2RGKs
XTEiyXf/Ygm5xpr+WevazvI12LDLpqJAEqwvwvsTsmcTPnn85vQMxRwoIhBb9tbW3rFljl1g/N1w
cBveapwmP9OnuBgPTmfZypd7+fRQkTnvf9OVIUi74MYlJU0JMDLb0lc5Z6Z6Axqcvvb9Oap0cQwU
bs7JyJIYp4AftEqWFFKyDlV+hNzpbUPgOiCHkLgRbCkqiGTtfA9hyJPQPEIVQOmXQgkror2ChmFn
RDKKtokUSSsQnl7yecVFGNNsCGEuBAQ9MuKedWWB1Q/TSyyNrYXoROWDLgP/9DV8JZruOA2dkjZg
Mb5gvD66I33mXOPRjb2+YRq3Diwa4vCzTfEJZg5NYqeE0YRGwYxTtXLU1cgY2umyD67WwN2A/hqm
bHiMDFhvNDIelDnieE2tJ6V4dPw+qlaJSzh70yWd/e38sESaElBSGIWCpat59SaHWXrpKh2o4LOk
Tjn661xvALrABSFOAZyYR+8L9Jh0e5UoQzNnXLwfGRcy6fV4mmZnfClmaIqiBIRs7zoU75qZX5Qt
c3lI0/0kyWhDa2cfDxSQk1HoUd5d2IDR+2c/Vj5YF7ybiYVgq6WeO/UztWWSkqZunLyQqw1ayNip
kDeUagXwRXgbe515iEJ8Jx9pyktUm6gifAN4kx0uKvuQkz7mF9Go5sXgjKSwz8Vv59GhvBVFORQG
fRAOfQZ0x35UGe27wSiaLUfDdxwy0K2M31ZsI4O5JTOU3ebJJqDm2ZkQpT9dDYuVRKuRpPNzXaqR
3Ps9WYnQ4PxhmGyVzUNSlJAfyeCgkN+xkePwmF5TmN8dJrOXa41W/mfdQAkMCufsW1mClanO8ycp
vIuLMyFK+4QMtACI5lW3/6SrY1IHHw6BrbEaN7vXyq7y2c4spOPtnE+Bhurs0Y3q71HLEk4sOsqC
GulQRD1NiMcsXrEoVovrdirkXAuD/hKZNEBus74I2gy8uod3Ej5uLr8TbnTyk/sjw0z+vWGLfnM0
VOK+WHLUhmYzEV8bZwPzSBn0dM7L+tDskq11e9XPXZ3eHSksmwKlRZOm8WU1p7cOqnNgvzavrr4z
U4HSVqoT2wLZjA37I0tHxFJtPDRFulAwi/aws7oHMpkEUQq8sNWx+c6Pwb20rO0Vxiw8p0f8/5gH
t3jlwcKpDHRUqEFsmth+Kkqf/LeOLcw8gReFZgb3IZ0XipqhMhAuQg6J66t89+XmpPIFrq1FbgNR
rB64v7IKp/QGNejoQHmHRguEN5H08enLvc9OupoWh112dbdqbaYbWOetRvcOQuEK2C3zqN9oB74y
YGpSlvE4E2AERwV1BM82khVVDwya4Yb1nwmUIE80sTP4gD/87/0MZqQDzSmwoqA4katfbXOp3DpN
Aaqszwf7U2IxoDiWvo705oLOESd4z2f69zE9jgpVWHRYceX4L667k3BG7KBvDRFOHhwSap5rsRn2
+5/WxemkQwLFMpoy/N35JYdyP25LTuRSfxtEE/zL10ueMyWsHEs3iaU9lE13+t3NN6OjuhuiS3pN
ZSOd9t+F+2h2ZTiI8vfME4Lp+zZNxgogOpHUVNjXyf6A2mNQa4BHtWtqW85foOhKw4hoIQAafi4S
GhZXR4eLHAdUL+wPdSjphcB6ZvG1QAWHR1kXJycp9+JJqaAyx13prjCQrPARxLOe679EznjY7sNS
hY3wauITOhIE8dIAbCAkU8j02FNXq7j5nE0m+qVkQdgDSohv9tjAscAo7+vMrjBLwUjEdds8eimH
Md8ycfKR52aSTSeKFJx41OMOST1dyHHdeMbp+ka3Oi8nxtfJrCryVcHEkrfILX9YBeuvE2/t710r
E+PTV4t5o37jyXJkxa66dlZCziilPprSwqcywcGNFKHpfqCkLWBO6CLIj/fogccyfMTtsw1lqNJd
G0mbKbAhHtoaLLSCk98lrZ/oOQZ+5J5Q9NeTTOEvD/n23HV8IOH9U7KCFD/3KfBohr+Ec3bniUCw
Y9rPy1DmIbjeBYAkZpXQeBDDPVZEvWbgfgDWDpQHt/mRhf+bFWNUnxozBcYe2usN1a+4ewdsMm2c
IJVy+277TstI2Joa0fLS8jcwsf0tviut9oH1mBK1hd3MsKHHbFgHKn2/gChLcE/OvtQjKJKN3Yn2
OcR6gdMLTwrJw4vKxzqdqYWRZwT7teDGbkwh1repPkMyGFakUGokEqxXkeMxBUYDqVUKg8RY8jnB
x6IJuPV6pU987QXlIfAMT35fgW35E/ODVCR7jsoptAp5i1wkTNdghij74VVphi2tImvUdzVLPcyO
HwJl1eE4hGtggIs1xQpn8eoDImNl4BkxPQMrZ+PtYeMri36yCE1HI21mgEClT9dc0/SSr9WggMoI
PduOY/sxdvB3l8Q7FJ2fcv0edugzSDA7yxcpH8f2oIJaRFJM7qS0yHR63zlA8VCND62agfZs3tQp
/RSvCSy04i+cmnJ4J00YJ7VXLJlDkxIDk5cUVHkdoD8rDZvGg3PMz8MRXe3HcIhyqypWc2PG73Ke
TFKn3J311PxSKvsz9hzd7q89S5nojrBtYiy5hDQoZPxn8qdsPVWtItoTd9YVDnpGHTp6vgsRuwtr
4aNDAr4eRXlzXEWDheBjJri7qxSZA2/7ylj9Ink18gtLfKeMkikH5RiuJGJkDtpqIgDtnqEa1C0h
MY22cii5nNO/rVkt91H3P/d+Xi9ycJ8WuOwqfgyClDPZ0fuLYJR8j5wayEmFBtU4UA1wJlrWdQQn
E2/FpBaQvw2AbYEh1I1K4jvR0Sflqr0gi+kIQIKaeUyY4R0CjUEiVkYwOJkhbvHgA9uuSWDcrIJa
AOhuR99ISyy6R0+a1VBdARWQjqW9HQqyYU2C0Dc+D+jf9BKOVLilIjTpcbYebb7LrabtnwPEdxbE
WiioSO9Z5kEU0NackWiL8LNT+Fcy5lJyGtVzGE3ARbj2AaOzo1CbMB38ijmT6BvG63g1u4PkgQ7n
Yu7O9Iqj+z3ApVRar7GX26/dnsWXKapPQ4CsR4MIVcySjt73K2fzrKUUMJnfxYFoMX2deZ5k5eIw
Q/DxRSDqohekMfDvXJL8hFTlpdkW8+vWQ3fSdE5+R0WriJIFFBZDclO+Mpjd0mSgVuxnFQZjzda+
dGGJQ1UBNodzFP/VqRZvmFEL5YtCWQQ0vEBmGRLyuZNcdsBHyvN7jPLIep6gr8gvR2M2KB7/ms8F
rHSGccqH2JX6wf1/KL1bNqpXL4tH24VodaZz897vMoGtcsZ8KDFmw2bfNen7M39kKxN79MZUskEw
USAvt3cel6q3B221/dFUPrnBO0FC4iTYodTeTQg/COJEktanPNWtQcC5gMxYbzdw9e/PS4K/2St5
gYNir+diaLmsOs+2oeWFgebpKxXplriKWbFPHZYHM5DBruX14YsqO13vAR1yTdhW/Nwz0ffbxX9h
XYISbZz6RK/z9/lYDj8tPL8wz7pWSscfy8HeA+4a/tOcPtjGC8HizLTm6RA4lsfEn4qcbYP3yY+e
oe4YyLJ8XTjxa/RMDzg+3zklFOIrRJ0v7iiMEgACBKbbQ8Ndrfb2p928l3CDsUzIbP5+fyzaJsgG
i3c67N3viJhTEco+zrqf2OAWah99Y6wxxsGY7dCOfvkVcANHcKH4lq4gCfRGLIic4gtK6XrSvl5y
kX5aYI8cXiS+uGTnr5+yfF1iiTmU79hVXams3Tty540V/NxTKefi3OiC+7oZJRlY0/Gm0kHAqPct
uGHxWOd1nvuI1Fm+8tztb+IF3BaF/OBctWKXwBf6/siTfSDu8/Kn1N74frDZFuJa4KiGjoExyYxP
btVdkvW90yUx31/5Es9YySCO5YbKclyaCYo2V/SI4eE/9Cr2lf4IO76v3xGAX7C+0/yTZZ0fJWJ/
RCwDpke2pimlTzQkg8k0rcp1JRczmc07Bxmv+GHpfXeige5nkhK8jn4gcVNdk275DpNQI8R6pyNQ
vVQS8x9NjmuHEQvzD7V+yN3ZHeOVHO/zleK7P6SFUuKO2Yys/+9A8JDAI1hIPIehYD7MO9Yq73fI
EHwqfoa+jrj1iNsBjoXWHkky5cEwiWP88z+gfJoJOdt4heHSTr7jEJTcGhLiS+8w34zpKELb2eMH
JA/ziJN22zykXX+LklnqskqbwPK1sO3+zmIbiwKXd1iYh6Ctzcn4qJ5x352KfW5HHQmJ3HEJT/yH
cCIHUo38JNjP3mOCui/ncEFRkqjIaVBEEWSctxhRdzK131uMHaXCx+ZR9UppkA0ysyjgee+t4N78
SWLJKjI0b+/XgD3iYw6NAsbYda8RJzP9G3YaL2U+f/+ReMW22GNJH63kUQCJ8NIKiiL/Pd8rqefy
bnrVPmvqjIupF472of72LzY7syTq8gqhsWLuMKEZVaEb2ByIjcYVsIKFgVlJdHk3slv7+TK6TQuU
w9HDs8+9TNNbcKa+RKJTAJiBDnr8f9EykbDl/zdJsBa5UnjBeAQ1PIe9HP8pMQ7T2mU+wHsTGdtm
aksNWeRQOfG0uap/rfml43kkDhAaY+lG/mW8J0ebSp3YJnUp9FnFgYi0S73WhQHjdUAIeM4WpKlR
Do6nbYMynaDRm7+ZfcA4JBswHe6ire3ekMjEkLOPjrCXITaC2cuVDgunWXB1hFeOu4L4qZ9mttaM
xsF786Do+nIbiZuihVBoSOgL9L1it5QGv9NM3gaNyQwU3pOzEWxq9RvVLRrQ2HimBiilzuyDFDD8
XWiKNFTodu/PDwKZShyWFS+nbcrQFNdEK8zaGibw8N08ASF0hMeIkdjzgX5ycXklt8FK1bnyhD/h
mUVXDkKeHz/IDQAhAevJ3nIb1kqkbcw+P0LUUHjucTGZa3QHN4XOTjDQZ/HUhzi3AuXUAd7oyi2B
xan4Bi9KG02kRzW2cm2aQaDwh56lkPVwxh0CKAGwbcG/BiGwpAQbrRP4PLDNExW/H54l0onC0wpV
0B4+/pB59o3HgfidWQiGzSACNMdk969KJalbIV4bVCuaRavv8fGE92/bl3iHDGOZaJcLA0TGIZv/
qIXG8hNlGuIzljLBlrblow9GpchryCw3AU465oLQaLIWQruesyNBqatlgwerCLVDKcy23SCUPjcN
NsMN8XI35ZRkzWM58ntwvlFqPDzaONlNZw7XRRCxvEq8mf8K8PflY4jl44DQoq4kzSYSdm/6SgFI
g84IfQAPFbYxRYJ52Gy/YFM8qRAcbA8oOBZWrWtvdeLd9bKCcg/+b2Ki9TlkozbHCXk6Kf4rgL7s
b1zZ1p4CSIHDtui3EGWhtiCWnFKA7Nl9NGUt0n8yDTix5u4fLGBA5XZbRKkKVUXAmGkOEzFT5kmv
PD8u8cqG7XblejrXr2Q+qxslafrQgP1ZpT7RN6oXaMVS6r1HZi03zNAtecc81Kn9ir4fusXU6Nvm
AN6pXbF/Q/5w41MwSeQXZJ4QglY61bKpe6Zr3LZ+Y3aM3DDUDke2HZ+oPAfhvQuQv8uL1lHMMVrq
oT2Y2k5eeMcxLUokxcat22cwUf2N8+raka2As/KZ3pOCzakKqoNTs7Jo/PhfWDYBoiC5hK1SKV3d
6BmXSiDCK/Ju2Gpmne/Mj6Koyz/KSpD2UtrV/+hHDcAHk31F6uSJmwQjiyaZrYD1h/mj4YTX0rvF
GUkwvJ2IM4TmyhRq+7oBdOwRJys8iSig+ZBe8ej5mun30HeHkr403HilCrre9I1F8mggQgOQAlLx
1YXK+v+I4RU28WLF29N77W24XUAOltb1BheLAVUaWCB3wzVzecEkqm+UpkgXoZiccEM2u0L6+nPk
SPktJ0PrzLpue8sxev+VULQjHWL5cbRzzNzJbLE4mQbZ68QXfE3WIt3DUfx30fX9DfVkD3qHjPr3
kqDyg8hooNEC1QfhUpouTMTu9/j6M32OWdkVxWEj/ZgHJXnr6bRlax9N9n7u+EMvcsSvOlhR2Vn8
v0xOmeBuvvBmsHDY34RSLV0tN5M1jKA4+gMx4WKleifVwdldgICVrcrASv/+YM/jWL3yQy6IxBSA
rQuW485bDZogESpkqzZYveRPMHCLKGYEWFYF8WQ1p3ZwRv2UU3zk54jMSV5nJokVoR+Pc7qwNg+r
1XIl87QLBL2me5jzWFRscQhF05NVsz7o1+Cvv2iwZWWiCP7umqlPJVTf192diwbb4O9xiU3nw4cj
+JPKBTssrWp66HdH9p5KR4ybK3Ajenk7MvQqRa0phI1jUongBPhSQwa86kW+A3Mo3IKbsmwB+D8a
5gEzuM5EJRlvN1Mj/Ht4sfNCjDhPVKMvF5PxpCklPe11WdP2iDmjcC7kGN6jSkU8otqAIGWCNkBF
E8SeIWVQDkFNYXtA6pdW/HpNQQT+QoKfooxR7M4mPg4C23as33hfv16Nk/4wJGVzjHkv7QgqWjvC
6HmtbCFiSO18YIyaL9N2eeWA8nbLCmy803r7boMb72bP0qTKNMArXgL5wpm1zqDginifzLIvqyQ0
PrFVG+lRthweLjcnEN8JQy2F8q/ihidJTaXByhFp9vBIOLCCnlsMaxC4uy/ozyjyEFAH61XEyj/H
yVD2eLhNpeUU52uL74Q2JYuwVsPlE5VolJf+VvoKGmKHA5lTOk6hRu/14F6PtwLkbYPH/u1p/G40
HZ9w/RezVDOl6fY57vuomEeLCEwYqGZaiMDVsUsvQ/ZZa/QMHXh+BLLdcXdJ/Ee8HCUJwcmyn0nV
IMYlp8wu4f3u6uMKqzVPikqjxw2a7PW6ZfhDSvhVjTIYQ5H4egxTJ0OyCKEFmv98BJRNONrQZq7E
BbPq2F6UoGRXQA2rqOjZfHby16DBkBNIwrtRtfL6h64oDqz/Zg4kWjEcDwRRmzla02VNBiPUWCC3
GF6szcf8cb64Y97l4mImhqWjZYctRVMqFNfSMVwRnnI60E/GH8VXae89dLTv12dJGrJnK/NTbuqh
NxVg+ZfFHE+6xFoh+s4Dn27taMq4CNqhSqjDWTOzKG1RTw1dzFGbyGqyvlXL926T+ADWMa5g/bM2
zGhJtfq80mob5K/cEy74PeD1S8EGDAFR0JlnipWA51VMTnue1JfLxMSYtzI1HzMct78IlM9paDst
vXdVu5obYZNabbk0MWGPqofBPwJ7VlcArJZ2kYD/djuwSg6JUf062e/qGwBlVYeBOvt8YXCPVMZS
ouq6zEGQSszu8W8arrS+x6cAucWOJQZWv0Wv06eNtqRD8W7fMOVJ8QQ5dQfwEVPPBoS+rWOZfLWW
1T8ZFFXjkpJSkGhhZWx6zBVALIrHcNznejuZgcDVMExYO9FvMz0p+yCcodja0ss8kt53TLX4/0jp
APLHeqPkpB18sbPkprU0rToCWrJAeI1k3KsnqIndWZUllPNZ5hnBLjK15ab/dT000wDWLyulSNJP
63ozQdbcdTD/RNSOD1+ZyFjOqavZA2fm1emTZBAnLv//Def99DQ90wI4nhHGtZdnRGgE8hIykOhz
JrwRqgR8Suo/Z3z7YH4YvgKHbEy9qdh/5Rw//KGXY08PRwcSO4olVtP5mK+6y2VfT6hwKbNhA9GK
iWmJfaQ+STwXOjFmH1vLn8kfANb2etQbGyXxttKefhMH5ojkvWZLcOtKs86yzT0CObBAef3cXapE
ZVHf2lC0XTJo6W1vndheGMY/AbfD3xijD7aVWvbVbtWejC5zVKR5DQRKTEi45qojjo4rzZc63nKQ
Qxig0TFk4M9NLm64Bp00EwkxQm+kKM31IwY387GxRtNxz7gs/8I31CaM3Tv/89ZKZhwkuNCwmpWk
w665xDHWFClM5ri4kaTRy99aNnK5kJKYhDbmULVyVuez4kJE3S94NMQhHO6O33MQpde2x351g+xW
Zs3p15P8Ww2jvKibXmuxI45irEwxHeeZ0tO4cjYrEQlEY8i+E6ETFPHzw0zgqdII+UQeoqNIRDUp
jPYBCCS8WepduCPqeXQnh4c46bXO5KnbDuG25tgBQ0JCbt6cvNOn6aAsS0TSTnpW3OGzL7CrsYpD
IRLt7pbqBeYTOmtK6q+Tn9+e3887YLC90ZHgJpecTYPr79gqp1HQGbL1jtX92C3lAb7OLgvU/Ojf
QR6B/Hal5e5Nviwb4Kq2hKgL7Tr2/+jsP73hZNhmwWwzV+64XFtouLteIahzYARCx00pKz8JmD1w
fzmceOeLuVvgZ+f+x0hfgqutbC6Xo6kK4giBTy6J9DwtTNGDDDqRkAygoHhGk+fZRpSbZx8fiQ1F
de/aaKIujoytSjzaBHdZbudtMw1KmINMdWUCfP5aYK5wUxtCaV3GL1TA94lJiPmRaZJFA6At/VPC
fbTf8SviIslxH6MlCOsTSkolW+r9kwavbC3IbSwLBT0jMGXU+oK+EOGozfnVF/klcO9zmcmJYsve
LsEIHvYODb3nq6FLiDDlw/JJriY/MQcpc4cWrTskLRoT+D7zvaKnmClRWJ8dj4HuBhGypr9y4b9E
aKhMz9qfkF2hhkttRFFCtB9KhsUvv+FxKgwzqza09019BdfOSmr+n6r5Cn/Z0C2f9hJPLtwsq5yb
9zC+OIjPoFnxEQj2fwLNbUTwgGDJ82WZLvc534FpzIAdOVkPxgzhy7AeYL4vpgaqO1C3NoDXefs/
CNoUHaa/cgVSHO/TRekiomr0ShU98OcY3S/X1Q9SSboOLWArRVPq3985QtmzR6L5wHQGu3QFnSMu
M4THzvl50db7ZE0agdSVWZb0/veze8br1T46+X+UgMD7EB3X6mWekkl8HbjaGwt9AfnBRXn3glCe
HiiGA2kG6LuttubzeGO+w3ONPvYqu/g54aodRegUN9BgI4f40B2glh2piojqXobyF6+QJzk0UNGI
TMn21eeHibWE+Os9sYr5uUeRaHEpzXLkiIyvHIFTQriWnwa+RSv3327i5zJ9bkWvkitHwBfvcZls
60JRDMtRH6d0HTwwW0+92VJmw9NW5yq5khq+2B0z20X8buSLINjcUBUCK9XQ//wN8SsEEyye8nHF
YcHPSBZ6Qr/83894auf+E67PjkSRpVXjhyg86fZXuhdcxgwvkMnCuJZiqYhX5wH1DNBoo6cEbctD
j7uJtiDvp3mQ7/YXiGR3NVKAj6032wHPClJO1nXg0Q+NW171gpYF9AcHIqd2k8nsCMDNYiKQLk1P
IxMQ2hpprN2a6jEhY9bZDmV9b+YcnEZWidbpTKIXgsVXUiS440zjV4VSm5g1Rrp3pYjt2R5tAdLj
GLJgwtVSDCLi8VN6hL6miIyXHgTJoqaEZJUJ/NXXZvZf447lfbFw2F88lcwBlrs7Hx44+kLwIgy4
UbD490TrSxS+Er5mV+/GkGfPzx2gybU4J52AkI/Arx3aadGbv+tPKNbE/bbwLSXwCRrFTiJYFeZo
/HmhWTdVfABeAk/hh1o4iOCWd+JYn7j8MeVaE15zl8WJ8ZOfeu3/6fKdb6HxT0gkf2DSxtF9LBtt
tWnv77gGBN3zGFiCYVH9uOz0Gl6cb1YMQDoSvTiPiYr+0wRv9uY8+2AaspO8IZGnMTKoPw+MQn1n
m8RC43hUew4PHPf4mmQjV0z2bKCswiXBsoF6jO/qfBsl3pmmOpWA/Q98eZsjYnTrdbjYBzuCwjJ3
EHaCiHAyDdplJ3Hp2IWvzLARZWfUd55Jz1xyqDB8RaHLuqn8fhjeHEMeV2hhPO5SWvUCH8bLXgOK
yyD/9HXbCCdmJP46tJtxPAt/W7waXa1mhA17GCFbes6sP1lt4AJT4zwEcnQh84wZfeWy6jDOyuyi
HSJ9h0//9aylQ47s0ozmtOE7e+Gn1pnXIyJqlt5VczJwsMeQYrlSe7QTphDO9YoMncz3KkoASkqz
U5xfZ2AyCiEIdHsVdMrTj2+3JT4ItKSge8pGkGwz8KBPs9yq4BqmPxZiZ2YQzIGg5+C+GsHMjBoA
3sa6z1EagcnW1aRa7cpqU/h860IEEK3BdPlJqy9YpA1EXqdNF+UEAgw5/jJlV5+LNrJVhzhbyDE1
RaIPeN9LrzIc2Z1LOTqHskYcWzwPt8sfQTZ8y4AWTDHXQLRjglEJLPNeVtutEhMn8jS4jpH5zBvK
CrtBN8OIjsaUubq2e8D/I76buzpiAOP6QJLna2IA8qPu1LGwaL9t+4mgNwOSl8F1d5sYRfUkNv2C
3Yl9MEBKOvr3gATsiBQAw7+jxVMZY/+i5CCsX9YE70dWodgb45n93+IZSrzr5i54n3q2pVv58+i2
IyR1MlaU0lHBAaLK/AT+qUXaxm+JeYeaJee4XTMEIbe6StRiPASYO6eydCitfV+OhgHSti5M42RK
N8K2PZdP/etwt8BubNoDb5PKma2GJChgct5GE642jnkq2NEDWKJKUssQC605I/mlxGQFnHxqmM2W
FDIk0aOz42pzVd5SNKtPWW/q0sxUtWJGTe87mwImz9MBYv4gqc3dASuf3yP0b/FvWQvJeScHH38C
HPoSOxQARuIx9hbPAmrUgoM3dh9GkMdLxZcwRn3LVyCWP2NjLY61bHyex91/VEnRbSEEVgXc3GkC
jJqol5yOVk0B+Slbe72DMwuacfaCv7axQ9h0N0v0VjZUiYogffJd6dpMIT9LZZRTP+YXgd2fhIyI
4m4A4N/whQHg2YpMQQE/Xwlj/O1QkkLedCMH7LCQmRH8rjoqo982/Adohg4uEdDhAovBchfZVF/m
45okWE3EZdyKg9dlNXG/Pto9RXnvlinrL/DM5XLBIrhBoe9fbt0/lLYo0nb7DZSNiBALG1dz8yly
grAUwm2fipbJyRQLjR411O0k1ukYfo6A7J6glfPupi0wkO6ZQRNZlem9cu3bXl88RBO3zVaR05ax
X7sFTj20zMMox8cG/VBRfwGj4Gcm3gijG0rYwUeHfnNFaXPWn1RU90wZHB2TERIUrDZX8nH47J6e
CEAGrNNRhO71/PAHvxNb2I9zLHa+fU9or9NO/f9pP28J8tqE2ecAZqiKFFCB5YFD+EwTx7KHiHl6
Ccl0Px3VV369HzGOAx8xSuYelukGssSOV5Q6CGXNtk2qjd/gKhwl/NEnvEtsvQ8IE0cfG05gtZVg
rY6VLWBETsOEaFQHCJD8jo7HwoxMNjAff5Kf81aE4eeizgMDOHhKtcqVELqsIOmBbcx+WS4UXYYU
QjiF1ywY6nO3vXFgsS3MmAT0clqpPnrhwnnV7PbcLRojRJeuQvB+GApmsNg10nIybtP4VbcMDPz3
Juf+QaAX9jPQB1dBgGibs90phob5Gylu620RyjBqi7x/Q/nYM6aWIKmCHweN9oCpzJl1tbjY5AyA
bWHDF/e5YckhGrVqEFwquhmZPPoSTpLrHKrsm+gzGHurg1zQuk/wbXt7aiK7uzvHTKgoGY00obkK
gLr8sz+TDToC6n107mRP6SrZLap31jCFVkdwlFiY7pK1YDisloJVf3/5DT/NMnvnrweaGW8l6frN
DYXBM32Hy9uUr9zclGyo9jfYnveIu7gGTaT3r+38K+vRrJNLYfQNIlXbiKa1kgEj6gOLAdgYeY5n
+wN++xNTfkztocmfm7xaHgocUUOi5hES9nKqsdCnuCe9iNc8N2BB9XRrvgQodnSJM3q2bqvbMNlP
EPlNpkTpj2Fa1vIyCtCQUhxfAX3YN5ytoIgZI/v60BaHxomfJcd6577luhN547GidArnz1G8vymQ
1Ju9Glzq0F9Ppr6GL1llOb+t7XwzLFWEnNAxeLzRY+lwMpMESjNEfvTE39dIDAXKY2MKYLbDevQr
IhcTzEotk/KP4TQD7zGRReKGn4SMKL1OqJyeZYwiOMWoYntTy329zUb957CZDjQjfSezXRki62DL
CvxW5T3xIolci0nvL6ztMku+QSBKa2kg48j82yXMqpSoJwdDHSfpomOXEVkucG89mwIQQa2lTABc
vcjupVI0yfhrg5rT+WXuACQXO8MK20/l2g7FSVDpUaEFfL1q+vaWaRCJtZf9zRpHjrGmi5a9OGNb
CmDFcLHCx/XPYny2MqsJvInyeKpIrXnqq568u6HQhyZMdHapjU5kdvGSsT86srRwJ5O9Kw2RIFjS
UdA7QY65nSza5QTn8gJK1nVo7QXg9g/Ex20CBD8WzlYywXqXjP6/fSmJHjN95cDnlRScZw2GRLfP
txioEgwjMSILugnxAU0lx5Stppc2cJrgi/mKWGwdq0BurbZK0bhp9I+sJQ7QVxLv27J95QxURdu6
S+wVtgIFGDNj9+dR/CVVNI7SxNsRzQxc1cMw2EjX3Rhu7PzYlTeq2kMyuyZqJHX6yxSKAr99o6cm
SBJJ37EMlqsqCGenpktuTK72bIGElzVSQg17Q1nCQEsy9zszrOTjLxX3qzLCOkRzjAnTx8mzYS78
Iw5a/pwHoJbU1IzPtlgbKDPWOa/MST1nyA5j50rEYY++tytg3Uxi823MvLQ/lulxaX4oYNXnqrFI
00fVgPgHkMVzeNw/94EEsfEqEnijb4hFNCCjgsntwarMdfJnqJSlrAEGxhwr7HMZge+vtTwyhEbg
95/cPRNZIT+3fp58UB5YvlI6BhroGxbv4+P8WgjUbtdTjIMN+UAmZH21xnkwq2RDF2u02O0Mtwzn
ttj4HfmQDalrAWJiHCcA+Dz4M5l2oLhgvG9P5UWMczX4SYxB8uQp5VXqHM/YXYntZMvjm4BeMZdf
SRkbbAWLpyNMliZceTz14QAn2qUq9f0YFcKfJFk4BlumhZn5c0YH4XawTGIzlxqsl+pgTnKOSa/W
CU71rZzsnaGaFyW0kYkltdHPQNpC9a5MT1mNd+cHi+Hh+PxL1GiQhLootvoer5oahv6xJpVIdamU
iHphMUSNLdhIazUF830h35yMwehr1lDFW733l9GbQl8KnxkfXDiFm1hmc8WkrBfJgRSrz1SWTjzk
CGMfoajvz5l4MFZt3H46KrHRti0Pv9AnuoK/VCWVF6pOQdTiu97e7MdT4MDWGeBaSXrC7N9eRCQ9
OKIEf8o1DaTjSD1vkUwpPvBGVn1rRCTgr9KUz7CZIT6v60z/JToFsG4whUfIR45cgtKG/ybLPU3B
YrMxqqyHp9I+VHfdKDYGWvWK7a5vcZ0Um17b4uY/sk3m+dMijH7dATNGdYbIookbjf/24qxj+XiY
JShXxNJ91K2255hDkBJSoJcxBqSH0V+q7vbT64OINV8Y1TQ0xRG2273VESNIMdGLD7EAJeowp3RB
mVfUxviw6ZADsJsTg0ol738izDDaV6nkLe7jKpoxcotvPf1QbRM/2X0rfvcnkzlVPOPOIik4Wlq1
VKtJa6iUQ5aG8Zvd+5sU1DnVpjVwx2d0jRmGWH4H6e5lHyxAgkyNmwIpehfgdJgoViA2R29ca6Q9
0QWLQhZVnox8bCUqCzrjA2AH4mP4Q5/SBB8evlC2d4FYKNkNdTbnghcCsS3r51HzIIDGailDG2gg
ci7EwinZSvXe474zkoTtaj7AjwKO/VM/l1PSSRL4rRRZHjsDKUByA83ukFVhM1vVyL0mE4UW40xl
AjgF0ZGAkDKvXoU6Lm8adDy8hZzGt4kKpeJObsLt+qorUhTA8uzGlwl/SHc/TOtRWXCW4F5WhNHL
3Hst5aRqfpiVWEkTLHWEdZOnbGeAmpkz88akdyUu3ZO4oTzLUJnWcrUyMqaLZ2Lm0eByb0wAiwZ1
qT9HMJIdHZy7wpEZuI6ZHKlEYxiDVOtZDbtzlIf0z1ivB/TZu2hPcBaw9PY5ngZCorAXnzcx9Hca
o+pCJdTSyM45/vle7GjuaqVJPVS1dy7S8lclTYPIVhUztrlG5kmwLjzja2jSxoQVXUCGh4rt0v/I
LfozatxHL2bq03b9fhHXtlN00eXv6Yei3rgwV66GhlpgnlWAxLAhge/LNbkbYuW+KoZWcfJ6eEVm
gg49HRVSHH0IFLHe2IuLVfcYVwnx0fBCxcvMQQP0zv96YoaO7VWY7kBmz65hgBC6AnS7bZkiwYz7
a9noXnFKrZU+lD98TUeNlSZe9cU41bgaoZ1kgLoKRTs8CYcd2hMMCJZnNhFPTQfWLQny5zglL0fa
i/MgXe0PmmiJa+B0LuqvlcbzYdLGIyx1+PT2qTJDo0CnezZka0xHLzeVeUvyR0QGYuir72tbJy46
Y0lXpdCjkiqsWIPCRrDGWe9nau6OSwSFqqpqmIqIqRAghEtfis5hMXrI7hvc+Zclj2RM4mcygRjA
dnGHaExxoXGpysre0VRrUn2CJWanYFnd/6gWDow6aaqxvr65SAF6T1fowlIJPt2Pe8wqWd2JGt5+
bMdgm4H7n+ivpOKenCIg2bqfvBGUbNfSZ6QOvWUZiJf9Z2SbLvYiydcCSYnvMugSFbxCoJX+u1Cj
O7ndNH6YYfDQO1OAbS4o8JLG3zwlYaJ8kDu87KZ4xhzbYEtbYIEMiQJEuxhwR6uxEPlBSiQMqwT3
ImYHMvBJQydVRl/n1soj/PEmU5bwTxtMvK7pMjoY7kl7xFjqOco0DaEKD3i07AmhCVm1Kg3dFWUf
CNwR49WlBHyQNDbgCCfh+YnsfRM7dapRRG0w3+pBZWsu2EKjGZWugeVgKZeDMiCoX4Nn1DVe4WVw
bzxhJnCnTJEfqpC1dmhmh3Q/TsgAywmGmgBmzckDtJgFXRgrAYLPEN+o2bISVsdjMfWfQk9nl1w/
GzwmfOQauzi4EbLsew0X54MobEbOeHSihf8AYwJbFP63ZeTqAMtGDdLawfHxcYyzx9h1PNZ7EJa3
Q4bdNTltfmpIqYZGa6HbKIReERKrJJ3Wm3t8O2kgRbZTrFHO/6XOFH9oSAyDiBTnW9It0RxbLext
SSQjR7n3F5S3hQRzadKES5rFR+zoqX3OT7hkTLTXoJSWrcWG/dB5mLXxSl4INZGiC3QX7UICC/M2
hKsNB2AwKNEMoE10AmhU8wmpk+hT3Zi0MaQJXUU5bndpUB6forgAxu0OmdrCd210xg4UIWapShsr
W4QmCB4yN0CBp7gK2k/d8ax1+uPj5Ibk8h3UJ5efRzsSDLhzPxYSICHUOn9acNGDAA4aGg7kx1O+
eP4XiAOVmcARgTtNOf10wlFTXa46eR1wqPPt0degwp96V78BDEwhMprfb34v1SSHMw2VWyGaJT8h
jUQfhB43WbYfpGZzDVddaByVxWrQkrCEFswW9TutEGEXlE3lHWJKEGli5Rwbqc9sIBz6Q6nklxMm
ZBxwHFsLfRF1vdnJhR1YtkJTYKzyXXvLCMezjMkwH0764PbPh89B8txoSjkevB5COCREQGZXndBm
lH4/xZLWdhky12qw2FpAgA4An5CBcFmbTwKU5+sRow0hdEIPLAGSSQFcBojMWLEeYplXKcDL4USz
s9wacxWJY39Q94G34eZHtcOF3u1pWnPPv1kNM2YPnix7MClI9rJtZVSMBr4BdYoFAdiIZ7esftAn
q7wOXPaVs01F1tUt6sD5xz49c+umyqbGvd57o04Yjfj8oPwb+Hg+2T6QzEWGCrag0WCd/rCavOWy
MEuE0dSTCvq9VJitRaKMYJFbJ8t/Xc+XBSEBs50hAGkYRBUSEdG1FWBehPmS29t8sVnvvffB7AY8
uMPB6Kp83/TfF4lsMZpzOfp/Mler1AHO0EZwCRDreMT2lE9tOHqqYa3ESbqfnVUbwg/oHCyE/5r8
Labf5bjGPC7YNwfPHQ8XG4Hf0t5MKi+OmoOrKDP2BZOaqcn9vH61YslPFecmhwsyJtjzCXFPmY/Q
TRCvJHyqECsEZA7BeUZtIuUCjigAgExMxy/mCIzC98kWFwku3UHWTNPhhbZTJdkjXng+shVME+fy
KE7iVa94fR28HDEX26GBt5YZ4eZNcD045Ppb+GxxPn0xh79MJEql0eMgjffjuxz+oCqKTYPQuPlf
C4J9LYSB9tlaWLQ8tXow2X+CWXXFkmBfjI46CsmFXTVBhNVdFRhDcGWONGveDI9QCLxxwIXz9XYL
VlVXLxc5TV9HaLDk1NbUa9WYiIf3R6lUdFxi8dmQxAAZuxqY1H6YbyZhs0UvaSpnAQPvtSTXZeIq
ybQNC00+znmEhYT6Xl5Sic3hGmSwY+0pc6uPkaYO2uNY8z6ayI5d/4JVj+kC7JSSOHbugHWl0as0
SS7rFcueO28txZ6ppsU+sRDhAGNFVOT0uZBkyPhfY0MeJ/M2ADYlJjmRjlcU0vVfvpfQYU9xVGpe
RVfbmllEdEP+8uZdx23fO9o6dnzgE2ciexz6NjiSEDgrOXudYOhSERLl3M4oZJC7BeUoZ8ScELij
DeRCbKcjaX6C+1yMZFrsn01jwyAoheRIoHckk3PZHbylpcsZYnB0vWJytV454rLYKdOD78BCLcmo
kDEMp5udhvu2Fv13uJprzHBLASTZgCeZp3+rul0+siW3cRhj9CDhMS2KOBS2ARvxSKRIgkdDT22Z
5tk8ueaNxRja93Vr4lxG8H7vOzcpEeFaCKYM5fM24sa/mB2kxEdNp6SbXbqEeFLWRumK81xBYZ8x
vp2fVM3j3gXQ8lYa2N7kx+gCGtQAhSFm7LuadvT1ncDQHx3a//T8B8/feE2J2ZAMMfM3B4/grH7q
GZpMdFuGEZ4o25s3uBBB7S6JKMO5lWKagtW8HfFd+NCfwR0U48pOLK58UpRnajOCVPmnd7Lu2B88
KMNRwH9ritm+qfrWccNey7VRlNinkU0SwZsQFZgYlFUMEFbHWeqyr6voiFqq0q5bOyB2rWxVF3Yg
E8Z3kRLdqsMuOOSfjgSNgL1BvI0TPgwpCTsA1rEGI2Gw2Hu9dz5pp2IJ+PzWqZ6Zdg7j+yxlP2JA
mhOLY6fD4qog7viAl92t9Px/j6SPc66OV8BBxOfWQNbv/REbTwdg3KwE4au7hHOjVbZQEeRFbH0I
QNk7uqTJmUZQDR88VGVgNVmx0WtCtEY3Zc1YEM/3l5JgZWnOyXmz8raKj0e+0WN1BsFkul68+LmH
CWTYZcj5Jq5RKKmfhrw0K3Qsz7BFkmobsICZ8kyU+l2U9xVAcZCwgZSmmDUIeVlcZ7AkSM2ANyZv
/yL9ubxtFOVKrPGRJ3Vtov+gN/CZdO5xDKI1PkbRU7YX5b2AaAYTFfm3KA6rU2w2T6G4QR8ouKf9
SAmagksSMA20El2OKqzAQWe0ojqn9asRaL3wglL60TzX4mi5kPI6kaIMwUnGt5irqRGWMYv6IABo
WcGBgVQ35j05bvSsq6GlkCVHlcccBdmxZ8cjmzYfBKNpD+VnWXWpiUmcK0boAvGdhCG/mWc4XQl/
P0xSToXppd5LGbkYARSI/P2vKrGtLlFvyMywGu996tZxGePaH2iUz2Z1fOknEHZ4MN3ycKdRCJS9
QiNXdxnuuqXbDR8LV4wOITce0b2NqY8B298F6oNNMF1+Jni+dLkckbZfYPUoqFXgSZgm5+mPgSnU
Zf/ZjPPICLE4+mao+h7ApEn+AX1tjPxtULdhFlz7nFjrRgFrVYWz3CVik3fljj5p2rb63Qb6gM6W
/0yeno70OIXWwVSmZEsOCj0n89usXHR9KEKYwJ4aScGMYi8P66jLdyh0EzOSwo95wIFf61YZPpNB
4a1xE2OoI+U3qnej1SU3eZJS/RpmrjTIII9KkiADxBsVokpGDEEWj19kH9npF6cFpTgXvEGogG9l
df4lOOhKKIIhyShPzkqM+0+nbCpuuIZCN1fhMm6xeV+zU3nRDPzsqtcDaXDVGYmNZV9a0CBKe/Xo
boUJUT8puuKtqhzkV14DDlUhA53aAah4k8Jdp/Nwdghwfpmif8hJJoyPI4yGNjcBY4jPBUjtap0i
jKNaWRGXU/mMQZCDxAjuYChzEC+yUuWos3veHo6XgVGsRqcBwlJTPVMSbcE69FyyWeuNrxtumyvN
iEMj3dQl5XM+gEcxbkxUZWt5wxd4mudPG6aG7ovmkqHX75NqoloGF0jZTn1ntUtyboEYcYbLAj89
iI5/GHhpwDw7FGxUKJ/Elb9MRneUNT1gBfPA6RDlvGBdW/6Kt+XYVTD6av333oTt/S3CxSgeHHAr
pUTZS6hkfs1hJodY6nF+oDfH0meP83DEWc7z+r5xFOWeH1j+VnDBfY9CAd2oJMdgdLGKMk4eTsXN
WYk/1KT7nvLdAvxePrNhM7Z0WyMgiZ00EVVnGw0eHo1qyK6cRuxat4DMlYRqQTK6ETtc3hkDKI4X
gd/p3M8Z9ZRnhdUwSEKsnxo/KfnJemvPj7RrXS5XtCLArpGhobATvLbuj2IciOkOB6MtGw/XDVtQ
tOAMKAAMw0N43pLIjA4eg58NoIgKObQKcIsY5LAwSU0jgVbl77h3PV3407B1x6PEPPpzj4CiomPe
VjPAN3kPyXPULVDEVEk2L3Szoj27uRGhuydvsmI0iGpxv4OXy0IxMUsWITnik0lKSgQ7cd2Yilly
q76whKrompclHBExjuRmscewQoad9iOXWNxxuhu7IYxdc07+vVObHoWQfK+zrNsGxt/Y7LZ0wEYM
FvzHlUdzFTingnkXUCMEaxI/kEOq8+JcWcZOuRZK3VVGxCDCFVaKYNbQ3zOegV6yNEy3lpfRpbbN
v3b/dLEv/VUNv29ff6RjmW4t90SbJCNfvqDsUBkGtOmo75m3kva8NS/rwu1EQRHZGoTqGiHxx41I
LXyHXfuSgpab8nVGrQNPG2UqCiMnCnBINNZxIJfgHnPkJuR84GMkN7SFPfxFxiu3B44SDf2Q82u1
lJdkMc+Ft9YLKM9snfwc1YEqjLIUsyP4DaqPvXSqYPXzVSEqpT9CFyJpL8t0dITqbEgY2o2GDrdR
2BSfMWY42fiCw+OvMK8rqlxiNVlubSmgsodAo1kZDM+wmnjPOZbq888d7zLbYdxlwU4Wqoya2Gsi
s5Byx65DZz8vg301Po3j8PA2/2uzTqT/JVTKI9JB/4JRlqm3c4iexo8p1Y4pqb3K9zk944cz3ouj
FlWNdvgVoODUfoHV5iD23FNohV/HTTLXrZYk9fujSc7WdHs7Y48nz8HAaVz12HBXe/PZR5wlh/sA
a1AmOhkgsvoAyBq0YpNCvcTirk0zKQdkCtK1ujkGfZ7c+QGvrL0ZLtcpluy/WLFzjZt+1Ii9IfvE
sMdt6XBG88MP54mOWN1hOKnLHoVtdQSsrm6qvCrUR/ALTI01QVQLC8yZec7o5IyNjm30HL+v3GNe
yJMifthJrnCVYV3KjmPVEW0666LHxTswRax5k6otazZMhxn8rNJbkvT+TjlUSa9KDEiwb/opln6f
9DHgp62b3vDbDkWTSa9D9s49qTr37yB1PQYltAcqlQhjFGdOQTLuHv0K7ak80M6S+bghAbkYGubp
Wa74cHm+Ib/Ju3RnjDrKNS5eG8kwlDyetLEbqwo79E4pNfxn0ph+9x1vE198Vo5YKYqD4Kb5HgsF
jTdOm4evjariZ+4qFSiQRCC+mgXexLWdufeRXvQBAz5T1BeAwf2RWXQ8Eh6sYLN+v5uQBo99DKfI
ftxEl/4dxiA6e6HNcVtHuG5UpxiTOM2q5uJA19O6dN//868k1IO1ljszOsyWohGSJmM6ZvJx7jbH
s9dV33ycHMUIJ4hifSJmJNtP/yhQrJG8QB5rT6mse6rppndjzmT5cbo1ELKH3x1IV5RJJjVO6CGe
OtgU/SjYiQvvr0JC6ArAjXgspRqSMOIUqLpidBnxdnnjl0QCTS5mw9otCAZ5Q7bafx93OFlFy31I
sDWvXHpHkQnIk1V7vCurDJi4P+o5Wx+Yb1VOwVKmKLPo1nb0EG/kCmrQU5G3Gm4IZFG0eX7D1+fh
e1cqi23byrLn8b6ry9vq99FHB2PsW4noJJQ3PMMQnMy1ZBzeZoknTRfl1+IQP16nPDJNB43VuMoB
Fpew9wsyiGolraS5e0lPn5F0JCspkmBx/54GCS2+wMfnbKpVBvIntTy0cg2aJuWURWoBnfxVTUd4
mTsAcJUXkQQkt0fDYB8QPpRZ3b+e7zQUgK3X/H8jdvXy20Fn5+PE8wpKBjAr+JpT/737fw7uOoVx
/bXrqgtAMFzs1flDiqbq8NBrF2p/MjbRkKL5TL5v/8r2kcrCFrLVamTLwBszUvfINbUp8MYh/aSc
KyOQmbY3KeyjyFv5sxG61vcHeAxG8XXvfv3hCTeFaGjRf6nFgblGmrUXi1eLC0KU8SZ4bXF6i+ci
FENkcZw9N8T0MU/+6gNqm2JV8GDhpepVaXkU/WI7f1p0DCbsvc+rdEYxZXewdRVDRzvNNOmxRgcU
bcPJ5EbDOJpia3t8zndiaGe3Z7FHtS/w4KxbMZOOTxZt8Rnj4qu8gdZxmKmX9+BQK5Ts1VA2jx/t
kRF1iqfzT1jAG8YwR7Dbd6pNu6DF3iZk7PRe3up9EpZ+K0100qKZgKL2fGY0+GDjb0Ar9j6nKp9W
GCLoh2pGo+tzdug/Yv8k7YW06Oe9dt0LWoG8SGBiXyLiae4Vy9nrOg7cGfZrI8fpkgHGKXewwyuA
GN3epuLd7a9mo7TODboO4I3mcl0FCdz5fakvQlty2NDcMJig76ZVifrjMC2TwuvHEfbvYXHBSVwa
TeLwOt01mWG2bkBEfJBnKn6Hvlp3bbqFiPREpoBfaF4f6kxhPQjTQ4BE9mXCgLwJ/mOkcg0Ix1L0
5kq81heZL9VBGA2a0+S/Qu0JachJHVS8IPd/fhLmDi1ltK4UgCcbS3OoDiqawHXiUht8DfkT9iT/
59Vgf9+AIFY5veazbrNS3oClN8ABXVhZhnUAYvNjfI4tElNaMwPMLNsLkooK8aOXl5fvJWwhSZNV
Z437jcc7DpG4o72hQowBHQ1ICR6t8fPgSuMRifKWHkolhLcSGnF8fY46aY6v5LUS/H/Mp+OHnEbL
pxn86quNbYYpyJsbfByRIk9Z5Fdb5fBdIB3NNZXr12bfZQ9jKg46JNCqWSg/195/dUY3u+6QQPLB
z6imr2ApdN6u3N523HaR/YYJTXupuR5dSTnrnlbwFpBAbLXrEQcz70PJNeYtz5vXN9z2z2kQkRvD
SkEP+SnmYSKuR/8XDLv6QPhzCwn5WmfQv5myTTOvGLt7KrZeaQyDJrgdCZ2eWg88moqEToR/9KnB
DssblfPE6pq7EAEpKmfYlV09/ye3dqJ5RdPHBcWumFuEJ7kMtCEWw27l3DQXjwh1sKPJ25G6mYGb
699XExoC4JFriaFvkELrgRKVMAzRY+9OIK4Y0bxrmq1JAL8PjXueLbdw8TiRZYdoeXAzutU337SL
MzmnBUFUwlDVjd1LCopP4LlyZcZOHbmyQY8H0zIzZRUNPLOZlzoUskjceBTYdpWD9yC6xlA5zUVY
U+ufIbI2JyWSiCiFFS/1LOolxuCuCGZkSnIOTl28CgJeAPbZQ0z0cMWHhe/abtn3IP79voTneAo0
XjC5PECwx6oGWO67ZKkuk0CpzFW3RxC/DG6yfHAsbZqYsaZgdOXI3kN+mEwUpmI60xnEpkm0h/+h
1uBIt5egC4iMLyfjk6OO4Or683JJGGhYybphuylq4C1V2FDavffjyod/ZB65Qe9W44DMsvd66beI
SP7GbVu0OLGNgHdrpAybf2iNxh4EjFVdIQIs0L58fPDdeLzBBJ8EWnkfFRh4RwwgX3vac5cJPCnB
tJMOrcZkkg0mVF24AM6SdkuV/yR1uYUptdRcXWp+vUF5FMcu0PJS9SqIgIWzYWAAO7JmHz7MP+HW
3DlcX2b++AE2e/usAbCPURZ0F66stYQ4woVKCeNMqGZLyIj1R1yMuc2WzFLPy3K9ZAWUeg2+HhWn
hD53wSthGvE4mjNwLKjcAQCx9gbNimyjUYMbP4HnaR2Sk1ZjH8XnQX+hSkYC472Nn7xwaDfcLoOg
VlqUJyoB+pJHrh8Exfkpn6bxE3/YXaSoqUlBQgzsTaPMv5vJtGEsBjXx4KmYs5syAw/Ju5STkv4J
CFJOwRfZ0m1vSo7LAyR7OwOkGCrfToLM6gv1ye9BgXvhzIYKPHrdJIVpVUxNs4Wac0jUaTZBLSmS
b/rZUASJkLzGpcgwlu8BIJcYNuSjSyLLEmdXt+LYxNkTzup7i8NUlsGnrPUovewHCYlm5OosDHVI
dFOxMsxD9xZ32sQN1Mi0OsAQn0JAFsOOdJf3eV7rXxNAvDNIfCnHQYAu60r/XbcC9F7Los5URiyO
+rMIgfifaeRnOMVOGbb0ELsHoyNCI0rkggrRS5MDPjjSxymhNwqrzk8Obq/7y/3k+98W/FCv+rHZ
9WuB0L0KTdbrtjjjj6oXoXg1lfY5cp3tjOMD3e4S6aTMTcDtc9x0+0LVaYs/Wtxq2JfdGXxn8lbC
LmPSWPPwPYf/xW8gR2mEhm/fqjusalzVMBfHXhUVdODHO47MKxGMsn7n2DCpZIkikebByCOrn9WO
PYlXhp9aFER9n+9AECmWzUpoVRlZc7GwSlXf8t+X7UlZodKN6M3/EIq3GDIBovbaYPNoc6P/Pbrn
dp9hCi1eDvfSGpuctflyWVbUykzJwGjDglTMVQQ6OaRVeXRRmMUu+TJrbhkQnJLkPZNJR3OtNOLD
JxlnSQ66tgi/qM/fqioSQ+J15rpk6b2Ap7ALarzeYFRNf/rkr/Ry052AkkTNZONu9mRX3Shhr6H2
03q7+S6OBN0jWQTXFW261Oje3VdN6Qeclms/NCTfnOt35qE1nfJKH/zMA3tfx3b3MnUi5zzSsKVU
3e9hcTZUwmU04IW6a0ZHX1xv8IRV4e9WZwfmnaS+oK67b7DBgDUJXfWlIiwKsCRaf3Xo+S+/PEP6
OJGqsRiY44cKqPcZZcIWVMTQTCSfic4kR1vRFqa4WsI+y7uJvnBFDQRQ9UaO7qzzOVFTWPS1UvRa
2Jkm8JQaDE+G+n4DGTTUXR/ipreP9LsFX177LR8Z4oLpa9oFifKnRVD8dqyb6LFKn7bkE43fP0RN
ahZhmhKl5ZkuF5+ExyU98/mU58vDAIjc/i06JqMZFepRWBI2hPgM1G62vXYT0YH+j+4Y7whraEy/
RvvwAI8FgxMCKcBD2SEEecNbaz7uxmYY5IoFUQqibCol9XW2fkTgke5xxeOaNQ7vOG8kj0jImqP6
wFiANNJEzvD2tT8iQSjUFZ4HdZ2x2VciuXLsagsgnHqYBuuv0f23wpXbUBxZH/9Kb3gqvRV79xgH
KHJvttv7bB8ZJHQFxqMQKDEeZSrYvFfv4Xqidz5nY135oZHbHDFeez8QD1tNHjtgK/IH0jVbuwJu
Zz0PTIFeQ+igDYwBMG1l2O8Fo4/cZcupqXGbkIGma8vMd5bUnlWz54t8DaC2Q0lV2cyVUqAMFCpd
/VGbjl6u65TSlr3p0aIVQSIhj0OtOtPlm5tcX1V8x7vly8TvX1Nf5SXRVXRCSC7FQmYF75C/zBqq
i0doUYU2NKpXd/i2x0d5YBU0SsEPSXgBNFM588bhTawOaxT1BT8jRq7c09i7WoSKY+QvJBrfencx
y68L/sTIzKPUAh9badQcsYUvZ+gE8y33kxgXsVdSbpU+JT/B5YgUJiUYM4JLmYwA3n1OwLlWwt1M
DGv6NvboiZc3khYWgcRJQdwNLUVLrQSAMEnARnire6ldfsOoxXC1utOHqzvrxZ2d2uskZoE4x6ls
aHb9j6egKPz40AfB8AsrpmYaWDwvxfLQcJstU1W9u/whoZIx9f4QHmeGC7Irm4qxXEcViLXIapy/
uTB/ZA8iaCXsKKa/2fcb62rdRUUmvsRPmODNi8C562IeN0ONpzx9/WtJZ5b+49MOsoX/nEXnJlEQ
WyHzPNFPXtxTm51Rw+T5VksWQ+8RdjvOvARYUpafVrfZALUvIhdANNkaUEwqoTzKU34HB257TboQ
1Ok4Fl/4YMVCnYGeTx80zTeS9dvw3UAfdf8mQNHmOodEbwV6AAlXRL2N/crWSiUrG2lVQckOezib
KnYvkTO/KmMFTXQ7kOdYbD0SIkfW2KDVNFcVdpVsZFuMkhL8oTf5R2tVN1O/nmZe8L0s/GGP+jra
3yqcnDmwLBtOnjBvPkDJQAI8azoR1GRySnGggaToke1hBKppJHFnqd3JPj8DuXG85X5J/C8iSRJX
jGaruIjTcqQpTF8yR6pVPoCgHVpON0pHZD8oWk70Yw0paDsOYJmh8ses6ooxkGwWTQ2CDhz89m+6
VeyyWjUzwAkhI8Mq2CDKg68RgXE8sO9AxiYqGRR0jV+VipQPX4YQ29nYAcifMewrhZSyWIcEX6xM
qAsMu30AuqppIOvOwmdjOMOALFveTqvTWFHYywZ8MZ4DrME75oJwI5aV3c9FVOsdRUrmj+w8mKt+
x87PPx6Ik8V4fbh2aVEFI5eCYxUy+UjMoMtPWdp7tV3+iQDVWrYwhicVO9enKrpaTPozLGaIFg2H
nq8ArpuqPYJAVclL1okO7Pitm/ImraLCrqe/xo3OWprrhe3W8LEezbp3M/873PmeKjGa/cPLJ3Sk
N3VrRNO+AXmLq/f/aj+S70noLdtfT9T3JGNALJvwHZ8FOSfONHNTsV3NULDjnjoE66HArYTFJVnW
SXyCT0sIqbmp6sKKiuPPqDXMGIPzaCuV8wJDU9fWg2oHSCQGrcAYHViSLLlxVWj5T04vY/eCm/hm
Fuwjn+mK6RTAMem/IqJwzK0vu5CeO7BC6W7HSB/8lTo9l5TEVGkSuyeGVyyMOCffu7LmmvHSG0i0
KYwp/dknA21trA4EO9pGZc12+oDTD29JqPjkaE8aVfCF4PKpRIJy1btF7njzR4P4SxWB+lliHR0a
i6+q9CvSJgYtuUgUwV1EmxGl/jTwNBsq8btn2f4gMiLIOnVI+EJWv0KFvgjUvkzk8DPGJ8NWStpl
zR1ifM/45IqY1sDbCj8GP7LAphH2gsT68Gu7/gDvU1JjgDFBq9vsg9/gkgTWSpVz49vLAtgU3Eyo
jSxH6ihIWvK8s3knaogj37r3Tld/2/hs/LwWrNYFLrOfiIcodBDtlARsYMiilJkW+G4VO2jYuVCv
qY0V/uE5nVEa3Oifsy1RhwXxZHlF1ddmzvxXUMNwyLtz6yiCXu4Rnuusn30WWM3tOiPLQa0ax23w
OJ4aF3PCQA2rzGkvnJYIRDKp6/b7HOvn+p8scUf06YsU53NcIwBIqQ4eenFHImvfEWhW1MH4BHeA
/1YgUJtfA8akHyjpC4GfMY/9KnA7G0w66xSB/qnnFk7eGVG51cz6KmcQ0irWJMCPliGnMI+8aiOD
/xRG4m1hEXTe5kaXt7GLISXSONVlhbDiLrnEddA1Y4mKQ/7QH5U9QX3drBWKxS1R2BJFx1CFjpuu
P+qvewSecUhb9L15bNrKTG5HUaQVIosHDnXJ4HPGyoPYRC9cYBLOItJQTpm1g/zEn4+8lRFV91z/
x2RbLcBZCVNnGJUn0w7sHR9B2pq+HwQHHpjo+fPk1daWyXLWUNOKVPoKT5oZG2E/kVfXglzcQp8G
/GhT9foGpkkyGgOJQRJF6+3/UlLVkA2kQ7yyLTWldVEFUS06u5Ywpifgj5uXB98LOiD+s6t2wCXa
PrgZd1Aux1CoIwtEANczukECUcqkc5OXnFDjakCqlt36UJj28CrNCghfPwpzUjPf6UahVQsBfWQc
dEXa5QuldL70luYVVSzI6fTh4KnNi/BHIQ24MvOLLZBN3iqQ3hfdG6po6YAMver1LyawrffEUYDN
ubNYKSry8E6RxWXVebSVUIdWa8pqkD00Jwjgk0Hli8dhJxTVGtFwqVDn7zfqNqfu/W04vSPsHtrr
YbfwddBjpxf0c0qKad6qeeyT6svRlxt/m0FSxGitdI3eoCPVy3FY9KhVEvlB5MlNsg6FCuqZUN9W
Vz7vzKn3OMeA+x7yc2TH98a4LV3x6gkfCNmhcUFOseDC4EFx3suIQvpvxP37inEb1h954g6i9qyI
mYsJHdLkfXWblaULnI3HuoBbncesmiH8icRLzqcDg4GWkpFQ5sMbwSwmqodMftmMQyx0t9NBCddD
xCEsRIrMQBpUUJO/tWqXBPXCnEThwGLBN5IU/u4i7TscdGdWKVdYYaLKIEY5pbxxEkU5n22AOEE1
GutmMp2jiWZYD72gWq1YiaqDjt1wU8KvOX47tG7l7Hca53+ijNsGRp5CVYG7TxAvvtCHGlDLe9jX
PAIUEjtrwhCVm0uQarvSc6VGwTwKvpAcW7M2Xy6pX5Le5/MhENywDIlrFV/BskW2oBV4RTTr1OVk
w03s/EQFAH+dFgCMAJkTCFCgiicn15VYE1MOhmPAU22hW2jgOGBBmjKLBrB98kV/VKf2rXLwfCUX
eRkrvgdudWO6/5p3pTDjRrn2w73qDBsJ/26qRwKgPdRWzvEpe/HpLj3Tf2s0rL0lHbTSYFFJ4lgS
HpebUG6TFQb6IY3kg7Txeb81D4zm9SiJAFeu6Cx4Bb+l0EjF3kpuvGc/T7Q+ukVKwsSUcXbtiVQ/
EUMu35wKKBq0lE2Fkj/su4uY863IDAfPmrE5fFdS0+SEwt7gW1qjQKELBg2XpnNnkdgVGex9zCyY
7rrEvhvGr4fPkYowmvf1B6/M2d7KoRgocfOdaI/M0p+cHYH+I1sErxfh6gcO0yCq8Y4/esAiniCN
FzbVX9F/7YGG5yjTr/95sHI46WqILaye24wFxbm99cYB9A6xwn/27dck1FaFEIK2KjA/iZQrs2/8
WCuQeelpKus3b9nfO3Z0pxwFnetjzjLnFAPgHvq4jqvaX+Q3SvlZ5LR0VnwCS04mM958mDi2ogiX
sta2vlJC5qSwMs9oG5qVLpm1xl/gIxDlGVrgO02JEGlNZKafy5UCIliDjsiB/+iSNdv0yrU07tRy
D+tuxmcTGnsTI23uImvGCPjYNInNhtEqgpoWEcKWw8sM4u3msZzciDuM0q7yi1zuek1p5PsM+gBs
CyMA5aW/I3KZSBqWNfDkLz8a44omMLHlykV1S04tmhbE2O0Vj5pLLQurP3hH+pOorXQuIUkLvI3A
mJ/SR/F9/1aMMqEeT5X5dlUUQBvx/4ac1psKIMcSEw4k+HBlzMsQwWbTBjZySpTDfABV1fjiofUf
bVDyV7cQToV2PWe18py7ODOD6vbN01Fk7X0xlHDtzrS6MXitsa0J0gD8T4V8oQSqEe3NpI4aW5DS
vpmpoahKb/nxNfMh+gpnPuCy38V4jY70tMo+yBrWkKCaMj5exmCMJV/TxXZTmlLeotBQ2EqGVUq+
shDoRwWU0UjAxqKMePmsIvp6vJy6DTKBcC36LWG7TULaWTlxGNYYXpBvBdwcRm6p1U8gTMWZLNgD
Y3pvR4hoFfZhMoEBx2yBpG6GnKA11NYlhZrCBrj37cFEZsNO7japLUNJD+j4lqhtauLBxYpSrZZA
45jYWrZCaL1F/XdpvMoMopSURQwZx0mP1OqYG4PJMLHnn6No2zEOwKQS/X7XL1e2jOVodXJSwEQe
+TXBieqrl+goPkKB0oMJJ90CBHtt6PvBHdEX3lNnJb32yKGejjbUd/cTz5LoyOK4osh5MHvhqyop
piGDxZ1qH7jgh67pw8pdQ7pkvkuxSDmhCSaBkAnhE3G9TcvFBz6BpVX5d/H6HFgj77A8qJNqidHK
B7YvuLympPiQ+ipgeuqw9/3r9ETvJdi5fK9uVQtb3mB67fQ66R8dsiUg3FcgSxfZYMQg178mVo15
D8UgnYxypZWEbI3Skp8H/3SgJFGtcXguNiJ0ioagWccv9ZCq+I/Mmvu+vQ9jUOPDqU+Q0lip5HLb
qJuxRkEYYQFZoeAnfavKg87YvakZJvrXavxae6i3yGmOb5vpALSUXORk0j5BVjaBa/QwMqNZC3py
bNsJ4cOZ7Tllv8Kw3/3AkrQxTPsxg0cQf/glwUSi+Dr7llPIH1JtXozQ9WrCZy+X5blhhCFa5nDe
EIRRGcyRJtjuf1pT48TMEIep90+ePZc4t2FT7HaiTntfM7O3OeXfk1sNUjb4gbYWPD7OvZJb8nyG
xovTREroOTWO46/0Sv51Vug4z9PLwNtIXAxclM6b5nitGft1GOCKaFq8DSeqptZ7UmhQuV0oeEgm
sDs4Knr6YFuXTUWcjkNm93Fqiqftcqvcii/zlRWZ2cLM+543ZJPwfAchPDimb3HgNpacgpFSaJuz
5+gdNTv/hzjvY3oSHZ6bZ5Z6Sn5rSj5GQNU1qu8fPfRF7K9XpsRfWHChnzf7bFrvduk/1elozwCR
QVU79+Joyn8ManrS+FZxjOpcKvRjEw9wAikerkcJJcZ1lup2cvXGx3s3H1vBjckwDb0Pzw2WP1sn
SI1jtYouXVLrVxxdXwg+KxZlcsBgSJBnIROahb0sI/zu8PonVX+XIUbIV2BmModAd54LmY12Ky/t
hoS+ESibQVeVldWJbH6myrBEe9N09lzFPq1zWFMB00y36eFpJe95UrAFkwGkGoarSqSH+YiHO+1W
/e9KL84uNYZFXirmPHDcpytzlu0akkIXoJo30WC7sIfhkMPCOT6SogDOCvHE1UXkYnkkhdBmsk3x
7pp9SyTkGTouK0WHRm3RJBZMsKohobnEsnCBHSHnqmoLmz68HUzsw98pffcYE69uT88hpWwJ5vFW
Ar4cVRczV0BEAfNPNEqh2CMGxtO4t66MgYMPAguMdvA6T0yQMW5QhkrWduv5MAUFu1gfbQMhpLoT
YyyprSl5P6fS2ec05khIOtVB5P4K7+CwUjAxxGG7ngKlrNnWB0Hh6hxJorvaIA9ZxbsezsSndGCe
kufrZXyHVsOneDzTEfRab0rwgM/iBhLdvd13BSEm401Seba+luSuEjk0AvkUyMzoBIH7/D0SrO1R
0medECCOJU6ydraZkp6UINdQhXGSopSde1tK0UPCMdz3a/ldf/wUYBJdZnccxRM21UA215GobS5V
YtKy+XMr4hAx8AvGJcAoD9V9vELWRvkSQOmE2oWh8SV0SEapuOqpkWwYRwLQLwXbyv9erCL849y5
n5VebA7OznjLCW7BJ9i2wEgfwPapbLyxys85Bg6dm5HiFgiBxn0RH+S3z3meLF+Ovozz4NDexzsn
/jwrB5Q+Io4L/TG3PgJga0khXME2SZ9ZMQDMTezkB2a8UAZkz7fNRpw1CMrU/GnR7N+QT5V5E461
M/IC1rUfdBod5luLLX3paikyD2S0CZG5fnEyYmOP03dBsVEIc/vLGfcX7wjgcu5dzgJ+oNjALoNI
e4Am34O3wwaI3+Y03psL52monoa2XiWEAQbjN1cZl08ZeetFDiYjaTeq3Ga7LSsprB/y7841FUOI
9yco/xvQAnTEwqSxYgjDVspBO3FRTmQbkVSIW9g2PwhSx57uoXymbE8gxEYLbLEH0QSYG0NXwuoR
JgX01IOIjVgOsAmoiPKKgte61t9KA4VVHuU1DBGlBclfcMFL83nEiFpOhCyZhs3AZfqC+7NRcEK7
q+f9MVOE2ytbXKmBesT9Ylvlm0hMFSJ/LSEj1wgQsZxIS9zO68W0X+dGiEXK61pMfWvPnQlKnJXn
fVFlnYsl0Sy8c75yz+BH0XbttXhWj1ICGzsINYGP4lgzHd8uUjN34OiTu+fNxDi5gd6q/gz+jxNE
Lz+O9sayq5ruOy0bMLyZnLK3KzZHEfPSYnwgrfn3plVEuLoEdhZ2NUZRy0QUYntlw0mW9hE3E1qB
1HG4CJ8D2LfAElUcGjfQGp5w7DYgLiIJ3LWsh5ROJg419LQONT0QWVRsn5QrW2KUwna2OZ5/G48V
7V5jxuJKKjvnx+k+geA9tDlNKo/nrYNeRk7p3+TGKzaRYoKYJ9e8ZtrsHBXGm79Rhz8komL6p2DX
xWJLp9AjNVq3ekcJUA/jetcJJFe/lMYBQU+5HWy0/pVxsAjo8zKvjYcx6xRBxiOzGfMGyI8H2AW1
HrjhcLKDw0WMCkQbu8rcInJOeKG/YCChR9WiBZXOC3t5KPVZM4dGh9l8tIQm51D3k8dOLp3lWbfA
AXecqt3U94Ntc/MZuA/4QqAe+6IeY5FwymBKIVfgLGIeXX/YBhnMgpB0yGEAVnTlJgrC6vQTig/9
i3GSVcG5U2Oxsg+JpE3PguVSL7nekZVF5Clmq0Xx0aJgC/YWF8w5zeh5Th7vhUvQgReNrKHxxn9+
5vpw7T6TqYP/I5Up/MVt+MEah+b8JgsHn2W+wj+LgakLvzcTJGiyIKBU4xDCURIbermAwNLyB61I
L2hHTLrk/ty+T5F2wASgH81TVC+U+Yy8MeFmtZ28wSZ3zHZT42XUh72LRAY1XIaK+Vmj1+TE8ql7
4Amg8uJUxnyEiRNtYPDIT1VpCvVTefHaEpKy+Rik8ksnO0Gk5JT+SdlL3iwcenVz3BEB6M4aovbS
uBvTFOtMKbSD5QZVosTGITwPXzxe1J+0p9v7vSeoDRbtXAusPlhv4Vtn0bu/tgU3hDbj6RqksQhx
9eaINObc6ExS3Y7bezbOCS27xBpRoxICdmcA0+AuHx6/lyUqkEC3Is5kktDu3Ru7uvJi1eiuJpee
VOCima7JpqiiXwRwMY/mWQURJTcE/bY7HJu0FcEXQgjjNfFIC8RxfbBVUeCM2+/s05YLH5ki0JjC
Di4JhYmPVPpCdWGKMPZ/u9LW28Xru9T9KVx9lRfsJvTy8lNlYiNbMI2h/wQh+x0cRYHeTg4sGOPG
+ZWkAKEe5/m9cS39/5J+bFkgpc6nMYB0xLrUarehq69ewyEYgl3rNAx1W+QSd0ekEZmj8kNQWXnG
x6k5JHjpyaeAg91xq6TtWrs/38T/s7GK6R+AzqZa7D50m8nwxKnMH20QoNYpkE6FSirJqUkv7PuK
KMAUsjKdcG6q/tvVPQw+L8lEuvNUeI2jh0YA4ZHC1qEFP9lbpH+KbZeDHOre2xYxiJIjSQPq0fH0
uK9uvRLN10kPuWLAboNKLAyq9tptf8yxXv9qxJzBoFUavkF9MiL0eVkDLwL8R9dzCRaogXmOFPlO
2Z0p3tsGXp0bZoGdJA5u4yOw+GZVJLkQOvE28I/UaOdQrIjSFHJ34g9TdZpF3ToA//i8gEySJdqt
uvBI0xlF1nKxldoUSLDqgsHq8AzJGX+VbDWRww4HzZoNMNLI6VMTZoZkxuZCaXbe9Tnaqu6ohA2N
qCLs8sejCPNnw7y1dELfBt8MloFib3kAhKEylZk47wwOLn/CUmGScklDHKfeauQvF9WCWJDHmsgM
pVas20l/h0Kmded6Rwb3p0Pt4P2fmgfnvwnrvoia67cmRKZqESmnhsiAvzHfFQQeBQG3aYyfwCgj
7cMotx60mXR/8LU9KL5LOxMu1dBZefJCqjua38FTxKxBOhdBn+KcPYZH0RNS71lKi/FksNP2Erly
xgOBKXKEF7IyGvbWsrgipfZKun5SinIk5gZ7+XND2ymGqpGlX2hjAfg5XM7BH5hrfpIQu8g79Om+
VrwE7MUkZF5HGWvo3V9+bXinFJ3e/6FDf0yCJW3sHoszuEJaDIeFEfqXZC7sMvs/pWtIEd3Gkzrs
3dQ02e6yd5uqvHVmnL5D0ur2XQhsIZrp08Bws1/Mkzv7hNc5Q6ZUoQR3CcmdIM+vNgW2EKM3JKsF
D8TuWdtybAICxj5Eu0rH/BWNRiLS9OvHE0W/+vzN+Kuumlsq2fR4GlaywTX8RMGlzQKQ2S4BGCeO
dAIM+ZywB1xSKJe5hK78CK/l68+lEkOsAHvn/Xf7eQVZC+N5poPzbYK4bEh2rIXyFa5pTyQeiYxH
3NsrJQkfB4eAujTO/4C2JcHykhoJ1FybQ5k8wYzsmtWIcONLL69XKiHZDK2gd7f6gr3PeqvgG92a
tCulXm54KuLKCJVu0I3jrDv4xEGZOADK+NX10c7dU7UkL2ZjmLX3H51rU1rILljHS3chkjfbYpl+
hEWV8BmqBY9tArwpB92G6dlPmMMA3sacZ0dMmeXyn9LQaPK50h/ZwziNsumCLUwVrVUO0vXUfuGy
1Ea9L38YBBa/EBIZvHk/Rn8tIB1GyFYBkKGQ7rAqoiiJI2ndeCz4KwNa7oEnf07G8AtJeSSjgnFr
qNWuLb/rAqNkmpSNF6dwP/mwHYRyt0KN7f5q3clK93DwJy0ngx00x+w4BOLiqG0bOf1set6XSsDv
PicpgubI2X0LPCxifvZrNsfLrFNA5WNB82AUCpVUdcQa9OPiUUBsrQvBZtFdT5T1FcKfnDfhMJWN
hfNBFN8eGZv8XCbvHSPCdp4XaFAV+V1M0jBYAHBmSvtPs6Oe+HkbSn49p0fkj29hOdgPiMeucswm
94cJJO6+v9fgy9za1dLwd8j9v9EAGKIFU9AB0xgettIUb3hEZjBu86g6Ao6HrjzRa2utSNFsfb+t
Mu0WIEHymRir+PgHy1iua4ROR72t+FGwzWhpN040+rFg0nzn8/tdhxS0FBYey34jQFtTHPk7HS26
3Yfp8NSXQEauC90JzdXKn4eI6zDw4eXf9ZFmV8zWzl1TdasMQCfLieCuk1DwhYqzTfaUJD1t0XQ7
f8OGx/HmBUvWLZnByypuwDWzWwCzw8pX34ozhPAZp0ZDiZeW/1LWza4rQJGhognh6vORpONXg/xU
BC/m8inM8fbjvYV26k6Wg1/Gz/SSluLtyt89y7GW2y/6WiUbhsfF1xRkWCVntzRjLgMhFewWzVOS
8pFg9MhfJ5/7RlayA7uZQcajw1MX5aKk75OkCrhD6o+OcyUJbm4VCd343HbMPjPFiAHbtDSlR2Ew
a5bSljEnMbcoGWD2HnJiBNTobh7+AMSh1XSuSgGrGS1tCEIl2ePBd8QuPZmzPn+bbe/syff6fvfI
+l1cnyefEQ70ZvFKQdFpCUEUe89bf8hvFbx6Wj3gerisjjFzDVXy+1sHNgrzIFEA0TbFD7tGf3aI
iJ3l01RJjcoumXwVlF1gLYVusWRsoi/gdQVJ5G0RUPqza3ImsHeV+saHo2HfT8uHRO2P9GlWIzIU
DkrHqUv62JJsw4WMKdK5qjaMP+jPZTyhzNIzpYTcKdguc+awYHSFsd/Bl5yIVVnMOKxhBm09egR0
EyipfOpEa6SPkp1kos0jtjXJumXpDHBew9cEWhnigJoUwTq5WBT4UMo+KMoweFOwLh3B8L/9wkXO
00VvEoA7vynpcd8W6W/PW59GzL1yp7YGf5E8B9NsYSYHpbDh6Au4eG+Kfv7rKNE/o3OV87j1HAgB
jPX8eZDzz2B/LKSKSx233E8N4sYtlgrRnWwZD/UqkOujhTnsI13pFjVpDfk9Hif0xuT/OsAs8GsZ
lTKuoPCwZwavyolevqM6IrNi2EnoHhRV4gXb15QV0SWWVJu4L1z/e5rilr/bnRQQQ3ComzMHm/U9
U961Zr4RWbY8tYzID26rgFexM9K12rvW83+2bZh9FAMUU4VtQ9PJB5dT2P2I0x+6YiS4ZLoqdfvA
LQEp9iuSl1Qb1cs7WO5rf37FOucLzM+vRV3Sb9xtu5NSLFdblA7CB9zy5pXlCPpGXr54K3ZydTf8
MFCsMdyj8kukGOYl0EpzUYA12/HCOFzphMV9r6SpOysleMVkRbgPHpoS0se3LztBmZ/zJqLBC4wU
TX2b39z/Gr7MM8FP3l0Geuwy9ornG+bPbNiRVD9EKC6dwzCDptpz/HDDE5nIt8SvGb4THD06cxMT
98so08k41txMiXvBd7wdYZS4mijs7dpvwYQFjqwfOPk/HMC1peM8Y50amQwN+BCR7pMRqqoao72C
+g8n5fN30EA05bx9jcr4BEvQadZuj1OxYO9w9JiKbYkS3apaxqhFM9kKyCekWVZ08vYbBQ1JOhkS
NaqdJXl8AD1vANETh6ijryjdTi+clcw/wj3jUQodvhMbHDsAs0pFyeKgtEodizkCO0IOPWW0BTY4
UfR+pYcvXyQJShpLpJeNldGPMb6VAU5+A7cdwg/3XQDzFH/bQQny5Ftd8zR9+/zre6unb5zna5DQ
36TCqG3x+RitbuBnVpetEBtlwKhmZOMA7KMsnvL5LCC7rVJwpovKBy/G/KzWqSJ/TWh4GGr2F1i1
Vj9FnKCn/Jt87jOgdBkr+JohdpFWq173bPX9R9VlKh94rJWGyVY7zo0Ca9MYZXlxlcKUzGp5JS3f
4CXdvuvB3KvU06T+0fxfNqISLLf2T1T6yEB0zQBiWtKOqscpmc6D3Hgqi/FaUtVRiQB7xIbjMeOV
fAQBKLmSjgVWKamFfeOxObc1e0D+cUf4+vbU0BqQTA3sJ1TD2K53LMj/oJb0pMx+T1cviICD8PS1
ZrgJtErz5L0G+udUT7N2K4Y+Fe34tfwdB7gtxC2h7p+bRqWcxV97dB2QI9U2kSi6luGIXmHKJGxg
zp8ywzbNa6Hx09ARYWqfzCu8yUUVWJsUPNBOsZJToFpBHEB7SvYx+16tkub6CQQ0JqQMuIA47Gw8
q7COo6+EhDhRZP6bXVLHD43pU4xgwVlSebmSUGvPOEghTGPbZyMYV3PPaEmrwkv+V03xDJdX6+lc
nHwoxH1Y7RN94kNSj4wH2n920eOjgQZSppMksGgDAI8wWIAQEyxsOC78Gxrqb0d80iJzAb2wT09l
ftigz8Zo9sD6VDdbDcYRVCXBB/hZ3Ar+ZTZm9CqpmIJTA6h97hP7+PnhMFcqTDBCW3mxtL2JINTJ
5fzIEY+rA8UsaNAvyoPneex9Td3ZgiRDIkHmVqQEGYyFNmgV6YrYg6J/NUTyhZS2FqTsGnxgawbp
3eADnNMr+BqPOLDJ2k4u5G2fCaOMN/xtGql5B9CGreZlS3LVYFQfFrUP6rZB+z9cQx29ddikAqpJ
4SWa0b2Q3stKte2xxkC7AAo8c3rtT3JI0uakzll85dxg25rx8wESfuzFQCqCy3P+EF7Ep1zmVbIK
B4DaVT5YskX0NsZkh5ebfTosfXHLFbGvLk7D62argp9hBn8i8PLvHT7NOZun3bs76/KeCI++FZBv
n71zbMaXiNL3s2StQFor2/0xQ0azaw0JQmxrFyp2Vd1qcVQaUCPICzTBrUzqIDXfS/7AVYTpT25W
5rtnm2PRG0iwSJpqY+Oi+gBoFW8dKu66TPdVJYcd8ZzXxZF3PlXXGdqsCjH0LpKRaUCcYHTN4v6o
/wFfWXle9p7+3NBYDekqXrRsVH8Z6soYqcRi61ktNoKT6aDSgD/zulKyeFWLES75WbXyVA5WgeFe
nA1sjx+6gHCQuSUHqwWolkOcM+s1QgpyTerNqVOFldnIBgS672aY3pgJvMgAW+UUtB8O/SExYJrx
59978NwJMNUYCGXzyh+U+cofdNcD5XVqSCfT0nxTwRMsvk9EjCOWZHU0RYQMuYori1bAtDf8CIkR
i8j1txe7C7UaXHOeJpGE7DgDoP6+Z8u1KO/NPpmNOVQNSqvTdKVEmDZbvIaR8LF8folE14iH8SzX
CweqeSbSy1bMwdDFghfprEw2J+epMrpKXN+oa9FwOD1+QAe148Nvx0+4A/vX7hM5fOWe9/6tFjVE
bg1/LY6OosUxmYHz0l5LvvJo91CGCV68DBIN3cgwn2FarP9DgZasd2tjXqneZAx4l1vnjGzXWdSn
CVWQNZJ0VpfY043cisVJqHuKv+C2mrV+HV/HiKmyE2rotHRuif5DH0eSh2uaA688ZvwMN1yvc1XU
waRLksEWVH6hUlzuAUwO8vZgsGG5QdGCjdaJtz3rROtzKRwghd2uYVGBKk9LiWEFUmoG3Ra/20YV
lHiBR9OnjALYhOFxTZoK1XYlNT+gdpJ9CqWEYNUZCbgdAk0SPgaFVB1nsvJvrftdad1dKRxqYLzr
Z1gqt28LqSLStd/ZzYIoL5BTp5yI0dV6+XH9LgqPCYJF8ux8HqBhAFNKKF9EzXvesM67DgkADybY
G1EX+4kffrSUlzWgkBGVEXSMqNTU8aT1Os2eOfbzMFLDYrhnexr3dHplPqnd6/bKbQtKXkwEfE07
TcNkJrp2egQ1I7WQNEcaIBHHyC6HM9ps7+xXXT5cxsotqsPTWvERzAigk3i0s7NVsUU+69R2Pqxw
mGYrSRi92kfA9XTQEUVdHTy9Nbs5LoVfVrCEcJT4gEP/9KjiM3aO3B91K13PxN/s2MOhCSw2WxyF
iZoYtgEor/36NKXK+sOfzOE/+wnMi483UNXMTbd+/ayalRcGGxjNTGeDaAE6bL+zLonGTka+ZmOZ
Z1oG03qy15IO72VAeVcC7YociCV/nNrOLOf71o1NySFMlLW5GhDpFWN8Tez+Kg2fmH2XfkrouRlB
RWZVZb7YRUAnI6tHRiz91bJ3YILC5YWvSgiHf5+gKT4TF5ue8qAARIQrEX57AP1iW1WhtpeJ51cq
la5EjcYTki+52QwaC2UsUjnuVxjVGsH+jJodsTJa/yOwodSEva58dKy3nfL3Av+5gDYBe+toCUHh
/T0rx7eoXd2W2tEus/9tD6LErXfiXhyTTPY8Mc37dOZ+DucdcKJe2S21+YmuHRyrKc0PfYYbufAf
QQ24OV3N0tOvRy8+PakkhKaQZUad/4S0q9qAQSQuvVrewogdoOumGed7h1dyMo7GqbIZnaDhAfAO
nwLxIxjqHlX0kp9tUuF6+RM6NlJOEysjvSO2TWe7oFYs5pGTeI0oLuSdFZGrkE/l6cXgrIewGmDW
WNpXKaRHpAtJkldinyNNwveiPcKzL3V+m3Zg7js3WT2ntC2v0Ic0ABK3Hsg1MkwkJ1OHJpLDTbbK
Kk6kDRCoGYOkm+wmffl4j/P5rvD6QAsqLBblf3VPBH04NWD1frPS1bRUCbKcExuO+iqlQEiqrYle
m3I/7p7A5wG2TFgq54W52/lJftZTh7V3SDJeYctpBWCkpqOByLXoofPnlpC+daa3jCcvFcjENY61
JufPgngZ/rHIJOl/DsErB3C+mZM1FEisU4QY+UdH82RqsW0PX5jhGmwMITQNF/wHArCu21iPIsjl
ZkxRQf4y6CPeQpK0oT0iwuhI2JIcITMNbP5GamyvoNMJwMj/+qW5jzZIOxEAD9Sg8pXwio9tAGkK
MjuwTHvUhvO9g29vJeTTrsDqPvDR6HNUsmDq7n7LMWt8fCOPwaSsKSxQ3/Y1mqHpNgqc+KeFKbhG
rrdqN88hv/FtTOH2do8083rqq4RqsnzhfdqLr1+sJ99I0VMAj6AxXPqj3RSDUm4Yhy3S73ZKdyLz
Ja2dqU8Y5PyQ9DM3UzQy9pWtFvDd8+7mTEBXKyjskl/TEZHqAIwJ6PQVUFsIOCWOL6SHEG9RNyXY
nqfXQmRVaJR7hBZDNmRV3RjbxjcUudUOv3njCEbHjXKyDCZBaPz9CRuOh9OShAxRmMQDTm8OnBeS
rmT1AfPtkK4fTNp6KMa7uvKN2WSJlkVC/VGyvFKdRaZS8PlnsXdPYszrAxkHlTqwyV0eANgbJJpC
beiyFPUgBavI5/U7UoWszFuVj+rdvj65bOrxN/HFX3nEkdVVnCoudrVPJngafGVfdu6Evmxv7za8
MEPOx3kK4w/n5QtnjZ7MPCd6RS4XUgXKNiUj67SrcCJDAzdq0VCeGa8FkF7qNymH+LqKr4ahPjtz
AVXT4RJnlVToIZbLwHTfxRDE9nR4H8EmzjeGL8p+hnRvmQLO9/f3BxHpMABSGo6UWTlFr64ctDda
ass38HaFapWV5zeTi2IiqSBgNFG2maC84EAd6Y3nDNIfFpWUTLWAT0MNUqs+7t92iuGwomOD8WjX
7ZWq0WjVAIDqUS8VJ02hGByEMZ5qRmaTr/VFFhIyt87utUdrgNUG1MIsRuNOzrM52f0uOi0Iqntf
LgIeooDxqRzP9zix6j4U3N/U//JSK1rlopNqySWwW4GJlEHOht4QcBn4JltSNbK4wtdRYxkBg6z8
b8mx4jIyHLBc2kNGI0I04INKgpaNNgcPG524cIA9Dk7mxObvhmRT14DEfVy+arUFFGyfoTwcbhfh
0XzpEvh0VdAsvOiXDY0jL9Yf1bHzGV7ThJYcJdAriYbe/PEKEeUZSUcU55ga5k3kdhkeqFHABBmV
GdXo/46kIQYiI7TeDkaJw4ODUMO8qXhX0baf5OR1jeZN8x1+TPcM5lmpqpmfNme72MetfELP9d37
ob4mZxqvB3WsaWHdmSZxtDhYR5o1tTsdrDJ6jzKupLXb7y2N1um+k+W+mDroHY2kMZyIKeUtCozb
oIpI+WlyLyb/+GWnviP9nJDgnhjU/bqujgWhL0VxlstTMw5rTcKBnM2MiESgP301ElMMbJ+9gzXf
4W7eL5//uqpfyg3QuUs7XBUeDkjcllOXHV0WaKQyj99GAinilZuiXn8bQTYKLhNhQAV4A+O8lTyA
w2Rquug+Jtq3EMncPc9JOxzGWN7OzYt9eN7Ct8eQ8bm0ACHKr0+jkq/69suW8NFv29B9kgLHjCNq
PKvN+dCf5P/ZfgrRjAZQSmVQjtu/vMIFNiM8uEQRap4tcockOWFmDhGNID6H3Ey5glCpyAlyVjo+
WUOS5WoADClQ98WYIfN7ZvFWrA2cUuVEFH8uwofXkIE0I8PxFTBI/WhgxpgV7M17fpMJIfAFzIaO
2hM+X8b53MO/MfEPbr2o9OKhkQA5rucUv3FH2LquyaCzEJf7kNsG+udN9wF61MLAFBfaJ2gp7D2D
YLCn6sRwT5e7gApB2n6dSheETfx8jKkTmgAYpXUqO6c0aoLtgTIcS4zcSh1kaKfKp6ysnu/ihDns
6n6GGWsRF5o+RQaea7cu+b/1CSLKrT6vJ1HpBGLvQ6C3qsNrgbxhZPUzAmV0HyUrexajtm6Y2chd
CwDKJ/ImOF8GFiQlL/6zrBUJcJK/qTieLlCp8TjyJ1Wmk2bxkrkQeLmcTTRUoYoxIrbHBnNL+AZA
9/a+optylCissQlaqpjGcgZFsHuMdgRZ20WNQnrIRkHVRJgH1x+noAUgZdJpDJyJrz9Ld6rU7xzu
4SrXQsPmMBMHfXFzOKa+i8e7Y6GNqXx5rzk7VzJcXpIQ2Q6GVwC/TqoNdhhoFD8RCxpEmCBOPZNt
pPF+w09U+96qipUljLjy8GaERXCIrjTlv0+xpSAaB2VhPSAVNjfSVWgQ98XHVKdcSf7Ipk13jqaL
1aw/ZFSvVRiCMBjjXk2zC6oay+LrpwGWVjRxec1UNgfYvSpYOkByzUiP0MIZxOaZ19Px4qV4T/tg
xy+Zr1k2vPnqhdbcY9gsbdUmdOiYzV2+WaLEGuSKf/KO/I02MT/kPZthC0VI7EMdIf3ARqomE88X
CrRm1ZD3WF0w4VbShbQO+7IGenNv1aCzpkTQzcax8fL6uPeK/l+rwIwBlF+Fe7rIypQrRjzNuneC
DQhtvipBvmiSLauS/wzTF+1Z5FApygFSQ4oe7SCKgq7Ijgq7dPjdMVwa7a+j/De2Gkgq8I5HRu0E
bGaFQ73uOTDJSLK1A52s1UR1n7FyqRdt2tXn9Kw+N90SuulEWVEABhAZG3yomT/+uof1d3P2o8AP
09N5rxQByPwnERjcgTbCAZ4MZqxB9HcxFUDv4YIElKwbRoxsx7WdRcb68UH3pY4ceocX4rK7WT2R
f96AIe0yG0rsIT//2C/9eHB+5+BadYE/LuaGrxSPjOf+kZzOyPI3k52/NnSh5Kw+AUq9MSuEClhj
IiLo8R2Cc2naoaxHdzopNulJumRl7Nb8DD0RXNUxqtjpnZ5zI49NHZN+hXfhGena8GSfJU2Cjhqn
1gG3nRjeFEv9tQiRhZotEr7BSNiK31e5U7pqAmv+sPcgKhiz8y3wj2ma1+Z0OPDE5wCo3A/z4wfU
QJsXvVKMmGXugrVSBzpxNLd5HprytiuCwPvDCGD6VBAgIh69pHWc4OSmvLx9LfKW1zq8diItIkVf
iEXdwv0tFmKOXwfFMjiFz/4dMgjnG7Q5jGqvcsftAEo20d/XA2+LVE2ieatg0DxSPLjxkGG4za+8
Z/U3lFnynstfQnOZKgyIg1vAxxFJz/VCZIob+hhNGPSjVHVYmFBWYi8dI+HsifpUxP8WC5TwXeVJ
HFfM2zOsBSskyVtGy8lC7dDUv6JX0YRZo35bw8Sdh4DnSP3P1qtV646fgyX7Gyoh+U+ZAZ5KK1t/
WBLeGT7qQk7ajeIa3Y+h805gTXORUO2VKM4rrYUZFDQABuGyIOzTfSBvE2dUeL6Ixx6MAgG4+eMv
zwTDQqUYf+GJCxoyXEQjkUo635sC/ErTfboSb+UXJwxp78/lRlqywnrJE5+M23Y2+Pkpk7qBXNPv
e8wb+ZehyUQ6r+AbHzcEHD9Qqnvo3vHgD4SEWpqrzGbrgnu3biMuI3aJbHvq3fKNj1k3UYYYSvo7
Olv1fhp/q7xFq9/WXgSJOEMnQKqHz/26OAPnFURMwOesY9KtHA73JZ25nwu2Sola3cvTuv8/XzwZ
TGeNDPJwqh6pGkuegnBc5J6XwChdE2u/6QUj+wid9BaVoFnYo5PWfa7uj40M0WJ9EiSbRlhHYhg+
Gm3Ze4Q22x6uhciEQf7qGDEmQbmEyGa2BFdRvrr+fgaxUZFKU9ur/lmyZJkHraBumQHb1OG7Tnck
cRtnfwpHUsSM6rYU+0ab+LGOBeElFXlWMVwt27mbwAXXzUeAAahA6egS+nSnzy5JHnc0Ecw5oxpr
OH16yEQpsI70osLBovMI8R6GGurDg8Sefkii6uHX+/tt7l4NavCCykmdKWgxIZbpfoY1LsMCBFlt
D4iO3rExEMeoMWrjHs77YFo1tMwwwQE7POe41GKv/RZ+uZ6X8pdsFOzjrSRM+uVmJBMRKfr+UAr5
2I03zKFK8i0ikH5XHwe7vAsHfQDf/YYti1bxgVt6x+cHDTCaBtLoZnX5nBA5qYT3fyq3DWaikSf7
cMk8xU4cZdjyemfxcuMI4JtNw/aC4GNxZ4FlRXFsspAzM/xIrsnYDgjHIAr6yofFHojJW4Dx1XmY
xLjxSWd2mHmKOT6rTa+Skna9TYTTxLuQNzXaZzKcmk/4MbBTrpAjvKqwnUUY+MoLB6uNYAZTDKz8
r9RvsbEqnTHUtrJdHkDBvUOeaixgQrpjJNG+dwukoxQFZWmi5MlNoLj1UwKqpm6cJ8r9T4BJki8g
zZe4QhBSf5trezyoMeI1NCO6LuFkZooHAPZipPv8X8oULFJaHvvObGGI5PjVghKlR9/vIw6jyN/s
XuuJGy6sQblVFs3h/rhgvVyYshgpbI3JEaUIov6iSDfpnxBF1Hgjsng9KoX1JpCWCPpvpizb6liw
pP2Zf3Yxzmq1+/Jls1527yGxbPw9xQWzYT6H6mPOrN4TA/9yjKRXbV+hpqlE0a3yGork/Kw0c414
+L82aVi64WjRygZISVEvRQy8YzBpLjXqC48t9VAdqry2Ircye7v7LNmRCEEh7fb/rSjKmDojxQVG
ua7soHz+Ns0ROSboT1cb5H98K5Y/L5Ki/e/fDb2dYtr5TMW+qN4FfoY7081EyUh6zcmrKkX7IuoA
gTIXFA+9KzykAmAPbpwmLn25LRJJ93klFsUD4vp1YlqC1kEh6oTB38maM7aXLHIIcNVs/ezUJ4Uf
/foSTSZmMhDzCtGiedUoCzhKau/cOw/+/8HMSMgIExojsEzhuaHvXxV/Yr+JTivKGR9NLIRPDZdl
Ts0YnLNGnrpvpI/ZOqdAoCNB413GbSBeq23Hdm/BdakFjTyZE3q8ix+QFwBff6QIH9U8xeZpFGS0
gmPvOueuDOBXQPAr0G2PTjnyEVJV+dFRPCJnz6J9jrgflPwjbxg1CF2JDRTA4jvi2Am24Dtw+OZ2
lOpaTotrw6eIekaGx4C0R7DfzANzQcTY+d0u+DXX2Hp4G/oGsLj2ijGdv1nJlsxQeI41jbRLEM/t
gDwd1nXDqrl4OTHT2GkcCZpvuyX6EbPoht2TAZb6L5nmI1eOIzHYZnobTSj0D5k7nKb9Wm632L8o
A7rwYuQ+m+11r2Ytj9yA0u9JCpLpJA0BFNHZ4ziH9GVXwkWnSfSqDfrJ/I9s9qR/OjhaD5fxQRVf
5Xz8k7r/2KgD1Fthb+hb3H+yxrH5gBuBvB9Q18KS4PlhenBDRdHFo6WWrn4ICpKAsNhjMnhQ+hBU
NVWVgIEVpZD4bjRK46UjiYa5qhY3eKb6xr/Idb2I7zFpIvXSEXGGY1/ilg/JbrMxfNh/tKsFxvQK
t1PRF3MnMccbBar8xjtEbbEblZvq8MAcrL+WUqlpd/jup8WSZy4ioEjDyyRZvJ7YSAg+3wMLHZ9c
1OZoJ77NZ3lCU+XOYBCc/ApP6NwBFjWd+mbjMeNZeTmBwkaEdF8S1ptuxlDc8lFQZZZwMZtTrkqm
761z+VDVsbZLAcTm7KsehXpt2YC5CKSZuKHf0dO+QpKnlwtZrqkPn+ijbfCZG3d0l8fAJrpTZlrN
946nQd9b1abozPU5q30RVfn1Ygql3Y6reG+JNGQFhQU3CwONHS3ORuz5DHhjkVRJW+H9NzNs8IGq
7i7BpSiniRM3+jva53dYw9JnO2JiRPXroeLW8JqtvOZiOowDCaJ8lwfGSe524rpiwqtWh3ybeanQ
xvVKJkV/iSGO++SLB1sFaRshBRcyQE57Bh7p0st2GD5WhdjIr3lkqfxv8Hsj1C0FUP7owa1yLa8u
iu/PJT8Eftz9bMcCLRTEeWRmlesg5QDhg9Q+XoWsDml9qj6Jt7AjrIWNHGvQC6bNizef82h+Em7R
JGW8nYDpZQgrk9Shz4Wna1KQxXB5YZxjnY2G2+AQZHNLBPuAtJkD0Qj3yL0nBQyBH+49rEClNt5g
yU2Rpmoaz3sDnZZs+9DIFVvcCNel3VbB/XmFrpnyyiP20ncDKwgL6TbpKxhoM7qK1rd9PJBVQ2gj
H4d7iXwy1/jPyHkVcidqA1HxFtTHGxpxon1NmD6bJHOgM9pR2IxmP7RpU3jjjABq8nWbxhTg0S2K
4SxXg2/D2opo30zeLI6v3h0CdGp6t4qLhVACJcnqRec/814hAVhIy6zZHi0jUPgnA2V9mvRupQ3t
JLrWCv/6WCjbL604iOXzexWTuiqzMzvJk+n4h0pk3qcD5scZ9J489fW++/HbK2LL2nt2M2NeByBl
GnN/yaOkq4i1Z3+SVG7Bw7NL5z3xbA25n5TYSxAt3td4IQDpgW6POWCim6Ez3okSEm/xpjKtBHv0
+zqCTcJekdS0iM1M+znhISDgxODskU55gR3SML5xVoxhgN7LpSCzUiy0hhcIV26a8YPpO3z4RBlk
qRIFt2V4hcvcyuz58Tg4rRDlJfCsVc4tbMFNk/6ZuavtGys9JtKBpxT/5qve+5NtVIVkqmd2JJeO
zYiCQ/E9e23YJ1sNOYVuuBloMmvJIvMFu4rDxiQLWp8qd17VlMRHXd6g2jNsKccRevdAuQw71T7/
DYmIovpQi56hv5Sdk+RX9tLYZufpvRk/QXrVqmarsiZhlpK3bJBsxjyLODzZBPZoeeHE4yoHgGyc
YcudZv8b2DQdFQa6umdIF8Um7wEFUA9FQBCaKs8j1xvqJNpWB8C3CsHvlB23N28cHUoKITtstzRB
n9pXCJ4ex0Wuj/iNkelJ7wBR/7wiCingt5mOmbDnQ9hjrKviK9/a84hzHorrBH4hsJT5NPrkaqx7
ku3MVyMTelvyQS8L75CDUdR3PXA/jm+nrroijOUbTCsrAhO0ZuwmMjCl3WRHrDeI9dZq8c3QyWM7
1vfoPWfF5LTL86kuAFDVyNpDQ/XKIvVRhq+xYK9H+d7OHsd71UBDI6GiiKRNT9tiWOa/RF5CD7y/
Rt1T6nMbw2L8uyMEL/siG2zRB702zMQdC3+Js51EJLHJU5IdaZY3QUG6icYTW/W6Iljib4yHC9o7
W0cBzMok0JFEV0M8y+x1zofA4kD13mMskZfWkKA011hXOdbsTU1QBTl7VxJHdL6igAu+MGot1jJR
hiRXI49wTimqQybziyI2fMELocTC5Tg/qYs2cwWRWvWTOX/PK4uq3mnFrI67szGThew5VYZJPGAh
rNeR6jEDnyMEfYF7Q8+QOB3s707oZJkcm6oTjLh9wjuJ00oOSvgFzQ8WjOh62VYEgPCPlEPMn9Bi
gr5+rWHPv/Ap5BOXf0CsUhIzIVO1MAW7yvesuqJMsm2+NjGTcX47hEz6xzl7zSwgfSEhaRF6jedv
T+TSPtJ21BmnXKzkIPq4ulVpizCilWsPhPRH8ukBqwrA80Nxr7zm9wvNHtTzRwXgL7nZ0rcftrqU
ps3OwB9nbHeyJ7hE091F2mg/7XgTuJDshVvw3VVmLqp5cEAd/MD4/EJ1cHAI+RIBJLjUUAT0jpE8
z5WkA0aWmYZVrTg63G9ySO42nSobvWadvS7WNmS8qVVHAECfccrxXTDjGXBNeAOXNgLvRa1V8dYs
6083MZpK9bHlIPcCe6gqmD0bwG6Ufd0xvnK5hoWPIJsAdaPxgsmF+K8lqGz28z/JFApa86hyn/V0
BMgr1u5m0HaVgMtYTtPv/WYk6PRi8cX/QKPmK+E1l87xuNb10Kz1LySIwVS1JvmqC4ohlXE5VyL0
sbCkzEwIj5mHY71wvXgepUITBXzPiULw0cN+rm/i7uDNAte7mMLgNaIkjpHOPe1P5QLyehuLam/T
sqnh7fbEQSBA7K2s8Upuy2QyaHNbDV1CnrwOibs5PfiSkAOtOhTjrldUtMTMHgfIYaqwgns4aX++
Fq+B+era1f3KzvH6aeQxQfxgnxwAg6syGYEFd8Kfp3B4U9adu/UEKvug+Bgm0UaFhtdio5C1E/N3
37rY+7AcihUAe9dKVmYzuxvKRBTRVxE/FrDzJPB3uRHLFILG8bRnGiJjGFyITxCfw+byAVhKMVCk
4IVB26lSSz6XA+qy0CrHrZIqWhvIZmr58fXDkE32rhkA300Gy6F9i4vzNvQvzJD6wYrqM7nn1cro
BzbqKi1TtOT1QnOTR3MVSX70sUqxlx39bm1U42ds6CUpOeQO95bBLwHxw2TzdWwzx0UPVw/4xiSz
pMiD3rfc4vaaT84OPfGvNQqGm4xiZb+qTdkfyUq4ML3PVDWy07eYKIAUO1+zHQ8kyySQC7glCJ09
dJQqmFGB5nJkzHguc2yaIK8PXuiBQSozwTyyGOAROm/cwLOFCk9tk+pWLnvYQTwW59O7wLZ3V9m/
Vt2BGA03YdarWJYtlOkSNH13qadArwQFHMyQ6jDJhAbTGFCZYWSi9jNXJH8dBOvk36aHhAdwrqMV
vnB8YfYaCfAdqhSKRTY0mM9L1k0G5OE/+Ztku8LD6AAz+qo0cmrbhmWe4oLpjQMya2JTpGg4ULTV
3bKkivHcGPEwXrAGQV0fZZOR7Hi5wi6nkPn5SR8U1Ra5F3uuHwWNWEAW0ogHY/VlXEFj815DniHH
eYZhzpp2DKMkuhyHaCz47tu6tkfZIjBBruxzWROHxmg+i5NoNnzAs7k3K+wegpI1FJ4shkQN16k7
Oj5sxGyleRGNePndS8WStfegMlmjwMwEDeUmf8vNJRKPs52/Jb4jqHIMCRTbNxl2PUlIoV2BjPf7
gbKFhf1qjGwegeoJvbip1555Myui4VuXpOC+tYjmns0WXd5dDzH0LBIot1hjSarthanSAOndwwi+
QR5xPOhMLXa8N0LNB2+MecrE92gm/fpkID945fuon5yowK/U+94+a1N9o788U0oqPBrxnqH+tAsX
LaBHsAtpEf0o09KpfsqdNOGo8xXgBckxMtB5RFliG2mFzfnCWEOt9mGLL4L2GhdoLs4lD1+NLIjz
q9/y6jXkGcIhxDEemMbMHe8J8Pc/VPpAZuIpSXosBg9b1CWzevZSY9vkknlA2tNWDG4FTTXw6H1Y
bVdZQPBgKxmoNVlDOaZws65MKXNyO4VieXQszPUWGjLrlfiNXeCpajAoaNDkD0czSXHfKMXsx/I6
XqajENl+qJA8Y+LpiRhEPOPMKnwJV/ytnsQmjDAVQL1KxLiZACtac0WJMm0Qywam/1BQM6Mt1ICz
dbOdTl3aRxXPMLvGFvm3jc3f8wHT72jYgvjouqHAtXYaT8NESJAuXxJm2Y+vLM9XHqJZDz45osOe
oM9G9Bnm0XozqkLRCU013XIQ+VQnC8vvEi+clLq2IXH4EP0ssI+UHzPst1qveDEMc4GKPeaTaK8a
gii51S9PZUk5qa+jV1up9cXpXDiQ++AmNsfWZFIjgMLC5XWNpgvpZfAql3jGz57xsxvvDrqBhjVr
hQZ2WIoy0RRqzVsFcXMx+/1Rdpxl0XcG0L0ehOV+oYo6dXputMQ6+5AmC3cxSoWDk2VeTVyWAg3F
vSBfd/UXLqIGp5VQ4QBVWPbibtddtTBzIFiuvboFOyYSupRdjJLUdU+MqulUZCJ1KE/NZaSX/zbU
spm5Zss4/JZYColQj36VtMxHifw7kyGDYZx0E1w9Q6AL7X9aXek/4arfGY3MrWsdmRh2Dlr70zH7
FnZWMIJThQlkgFQzDCCZqoIe/WMFAXdioZ+sqSeaUnxEmlOGUFYbiJUAiYG0dftzE1aPZs3VpPmm
DGkRWNay4DxrxE6ujx3zLdDseaBYrXaH4uefvQaMs249VT2CFL6nxXFjIz99wh1QiQGwgZ1Dnt1C
pQgVaBJ9PprIPy+TlriBKj7zcqLDKOqXUfu7wypCqgnbwrUK5s/uTjNSMLkR+PTibAA723Tf1Gg5
75yvnZSY8okCx9EPF1xbboho2hT+/BcNN0vNeqEyV1NyZtgSpqqAih0lDyy++B66JgYSnw1JliVn
P95I0lkbVymn9d+nuFH63OgTVcPGONj+0fiiCelsINxDgPV7IQqit6GA/jz4tk6Hbf67JP02RjYM
Ovfk0LUlw1FEaf7ktzXPXUSP9L7kQQOMURcxggBtfhh46KzS+Mb+3vjP3RY5QuVSmMA4ItkeYh5d
ieDOHDf86qqlrKYX6MGS9/YHd8M113d0MbrfitBfThIvr1dtvg/MQtoSiISU+/FaBryRyzEu1oUT
oCRr2y1jNtc1AgeXSYH12Xm/Wzi7XEJ82zJizjGsWI7fB9TGxgIzgFBykG0ZajPXM+FSvWeFEzKA
GiBrvjHcSyYLUy/0yHmbf7639kJ8Ve0Ji7LFzcPp4neqvG3SDvFJNOPkLkieZYHNEORqElmMxoAW
aKNAf7j33LeSEn2bCfmo2gRwOVs1KMqgLdEN+AnqI9rxClW5EeqVLnQ0HsFYuvMg6LMKF+LVQrh1
gN0Z15VNHJyUfVmxxeWppsiunlNS/2aBeG8F4P/WpQgNlbMQUptGpJ6s3/7eHLU1oBO6D7iRXsSb
L5CJ4kRK+vSruW+dtuuyxgyOkRDoxG9pbSNLKxQLrTe4sge7++BUDbWrR4Go7Nyt1n7Ni6EBRnWw
FIpPp6ZhEjNLTDHkRJ7MyXhrJ/PxUSAyBjLz/99yQn/SjZ4/jzQct2aBdaqLl32DkyXtyN58+dOe
IFtlODdpAqPZqQvepBPk4kCtAtzahbEF1o9tYhQOF4XRDJ5uc8V7056Urgc2K+CFeJeU0BeiA4nx
hDUrUWIVW8tQahrxnU/Bw9q/N/XuBtte40ic7fikUnQSZxVQMLh2pMsXeOZZk6u7R2MCx8MHS9ru
XNtrZGSo9KbjgXAItOtsd0bnoWrn42t7q7ub7mbsUCNnIQRh+fMVk2Ep8xT0Ifb8xYl04ZA/f0Zt
+JWKnZueZ8SxBRqJng7WMBkLmq8BnCBXSnYt5bEXT1SD9GYvN2EdKr0OwzO1CHwidUCGGSQKjrDh
RAqA5zdULUSq2TTHnMi3ePXx6smEesONxm4vDr8KkIymdFn344I3knvfapukL0T6GWO5BlUtFA6E
1fbI7MRsTYTWYtrGKfUxfn2toO/9agf9t5pkcJndd4Bcx/MF7blNOqu3/U/PSbAbhRVsOgl8xUSb
Ki2Aj8iEfuSppyr71Ska3JhET9xaww3UiZwPKkJsfzlQUmynhEctqjuSJHMeQAr/xqdcBtIcc4nR
m1907P8ioIg9q9+6Gsqi7XC+srE15jYI84ziTodIOcim3r/GGLMIrca18mWftiGDGpeKpJto2y+R
FhBHMZCm9WVRT6Y4GOqzhy2j5rl6kuMStxp9mv1yw8yIKShNZxzY+y4jopChCjsXWudvdXWch99r
VtQ/A2Zdtc+3OKz3vm3CtYLVLQRJ2sUa0RxM16IE4zE/ZP0m4dDWPH8cY6rcqa7WzjRT072aJW2X
x4guczlYZgsrPVVhnLiPjdKwIVDP+Xxj3eZM9BvmSTgmh48ApUAgvESJy98uQFFbt1lBCjcpzpSb
RLIs+d/dPR1fRAA64XLR6DFHcqtEDn57VJRc0CB/4+q+VBkXaN2Ng72/+eVLY6dBZo23ebbhFuWv
kpo6k0e4t9PpQVWz4ic4nQzlgQEL53aKGXOY5FUYB/H6izdASBoijjqT2vCDJo4w+Z4riay9g2EI
ufYntBfLaLJWgUlxqx3bOw0slja8ojFo4b0vap0XT6srOKj9cCmNjcpNk6xf7Vj3l15rKCufPS0i
7nweUi8InSogsC3dWq5GHatT/IHrfkg9aMcNuh8roQNOfaOcrpA3qpvlGZJ9EwQvgP1Dp8RzAiR0
GF9nSqBXNvuSowngc+x4PQJDs2bTVZYUiKTwyrIHJ9ww2UYtvMQLl3mauQcntanvEDQzDmLCEaH8
GEV+tnuY9KdW2/1wzs/a7ccZjjITN3vlbo3olfEXmzOHlGgCPmSF0oTy9VP1TElhBr9JkXGrIrd0
XkZSpHSBA51o3XW2O5Tjic9RdSHRj6IhTrgty4SIP7v7jgmO1Uj1nTHccq3fPVde5VA7fg+Hfle+
r16bWESIDOfTxMWIPStZ+4Zj+2v5cPV3EpWl1lYDoF8N0xOT/YCcg7Jxok+udNVZc8onedeIJD89
78AJaLJ66tnZWlsdbVrXmqqY63B4UhnXzjPxLb1+pdHmoBg0IClWM4WSMNKlnAmvBAfA/dmnd1cF
Av2axT+r2u7MKQZMfjSMw7wUGI4lyFrNgPFYJDX1IcqepUh+CyrkbeMjKIkZBwGTaQHV1v4pv2dN
/v6scwcwbr5sMfPxUa+B8psb/1p/WObiUnLHrB1dwATEGFD6zRzWMDhbBWmdTsqYSooFVqLeBqHQ
98cBYTSbn1EqwYnoBCOndCsrGRzFjjZLfSObIj/6GYV/Fayfw76gAMPbeCNnexR61o247DyeXtqp
9J6ErzwaAkqfJbtKR13rwT67nlhypxwlhAUawYvAk6bnMVY4OKRq1eUi5BELkfXt/RW2Bmnq9Ix8
gfyU0YMOocL9TU0njkSyLLnKwS2P+YbUecoLO2HNBbkVv3zBdCb+k18siXHCUfbsowQyj4/2u8gc
c9RYrJqERvWpbz4TolsTXz+22nDiDv6t9A65e86wUOxoqS9FkGxPzCMoOOam1K4CoZUZeF8KfYhO
UkcVSPN3yFXFJv2cv7Nje75C9d1H9JJ7WBGJeSHEVXJNGzU2Q7dt8iAg37hB/bb0S5lv4yYTLxum
KQVoj+Rtb8gytwu2xYO2F4l5rxOSHHlgfMnJTCONl2b7/UG7DE9/gvGWct/coGrN5iG8moVmCx5e
HUReFFo+PJRSrt5XalYI98fqyGmCA9O5ix/pz6o4uz/sOINzmfr4VrqJhKkDmdujUA1IWpAxpdVd
dZWPVN/m5QHm/mJKq+BlaPqthIw1b6BnMGN9sogHdzXIX1uJDiW/C1VMx5SiV+6nuW0eX8hzN7I0
vTw6RR2Hp4UICABdXzpG1egE26fCz16pW2zcCRCy4B5qJ1Ieg06dVedN+e3VQqYtPrYEkpqQTG5B
9TyDbNHLwjXBoL/cEosevWvJwHKcSWMZLb74b2bqjWmgmT2quCKh5qdIDTCM8ibUlKDRM9UZki9i
tqsSW5i3vvlbUDmbTJBfwWaQ6R4kWlcNT/iWNyCsBE0dNYN652Rkb4F8M27MyhCToLmnI8d5AcHs
805oe+Cd7ZH9OMru1ctiK8kUIbeAW6U3XfP7EhWKNEnJtA/POiBLAt8jk6Q1hwJX3M59kjzi8Mf2
e7pgePA4UzW51fSIkixt6yi6VGRN/mvAIdBabdkkNxs9crMZLoH8VjamSZy2+kC0tOnTk+ZZDAHv
53w8hWHwufiPpwNrYeDf6ac67f7cmGhLVJiTzRzYo6YQbDMTqd7MlbO5X70krFeHDzRcm6g/qhSK
Ov+vzu7/GOOD/rhvvA0bjB9p5uFexniP/N8jWOdnJoSABUNOF1EGY4lDcutn+X/spJDnHnRFnzPg
dtjbArfPdzdPtqADG7Uc79bB+A1d2+3e3Ce5FTT9TgzqhxAAxeE186ryDVHwZQfwf9MP9UVJ8XRb
F9dIMa02vRrXxcXC+9sEO4FfCzffJhKhRplJKjK5AsJukKeg7hxaCQE2+/64LJMriGUPW6QxHc0U
vTNvPbtmstkw+VsQZKYhUjTuZ0BJLuxaAXUtV0WXRb4xv0IGjY8JoNYE6XP6aS4jtch+HsZTDTw0
oDKOUyuSIqWa4SMT4Ppa/a2/OuOBA5o0DCjzbLL6g+r/KiMXe2VnZ+Okyx90gIlVs4mcJyi8wCkA
lLijMrHNbnmZ80ODhmBHiOtF7oQvBriTnaxqMiXh1ElV8cRZIOalRoBK1EvJjCe4MJ8wHV04ihd0
fXQxq1XPjQE92BtktySwcmGRitkhftAUCbAKXPS5JKnc9Q9c4NJVNQK7RKMNTcw3FR4Wrv53cdOR
AB4Wq6IDzZthzf9+9RA+1IgybvLyX19a/jgkWVMjuf4qvkr+RoJOUA03AU5KiA8hyFSVTWeWIITg
HAdzgujw1tarVPVc2yJ8/QGe0DQh3KOEdo/ePwlSc4Krzg6ZtsxTrIW+ukVtxe6zL3bvlU+7ki7/
RQ+hbxK3ruVX4xTArkm+y1e9+0eE9mkl5IaEiqeEpRetTpOVMqsr4z8R9Heap3OATLC6JoSYWyTC
/AuKPoJbBcy7dDAnpLPOCeek0pmDVs6YCy/Dqf07W/TbigvoSTToIzKXrVgg7CXQA2e97plLuJc2
H1kEelt1ffO30ktpjw5UNuFLYxd2KKFbl23F0Dl3jOJ0orJyzgnzxYkhI2eMTq/L++tYWxWKAVTX
GU3WZhFDZuUijQQHuhMxL+DW5aDBQVTZQZQzrVzXbfYuLCf1YGefstfjkVdl2JwxebAP/tcGNyou
BEpTb68n8udaxU2Ilkot9dDaVm/myJLvdRZo+VxOR2nCnblADT9Agh+feJDkLSBMJvPDZO/yTeJ+
/bG7fMvBdXy9VP212XJRPA3KFrnedjCW6rod/KNGR8vtippGAlzmiQ0t1rZj/W4R32XESXUXR/2H
rDZgh+FO7EH0RuRLzhxVUXXVTu81mJQNP2nQuNwhya9QBOOdFQ35FM9Hwy9fO4PoUHD8OSknF6UU
V6b33/NVXORl8huEy2Xwhk2yU+ppJtJtJwbo7mnXdEPSifnVoOcA9QnIlV7HZ7KaM5OAdVzcKVSI
XeNs1qkWqJUDzR4mX6g+vdzyfcCsUylG6DoxRFXT0Bj0/Y95ZUhzwP7HXasy4H5NIPyvsSyIyWvB
yiqqHH9XSVrN/S3YxVd5d1+MoLHMZE0O3nx3GNs37rVfXhkaNA6JIDYMNud9u47Cpp0vkoCxRpEM
Qxie3bp/ZrJPy8Go+wo7tkrpd5ZqPPinnS0hvXBz0golcBeB+Aljs/EhOgN3MV/wb/a8VNRO78Ex
+M9A3To/MbJMq1plaLeSo5icOCOtNN5flQMKf/HtUvnImDbbkPMXdtOsniVAG3lcjiju209yUOM/
eaK5NvnlDZnLAizQTFstf3+31vCs4cEvEWgR3Vrblzeh+jFvSXoQZkTHabtTJMMf3wEkTD8+3lhu
zpmvQhLeVWME5UPW+aq8a2yTPXhWUBfIg3dGemhoDsYD+NtYqabURM/vOIiyQEuVs6gkJ2JjqIkq
/UT7KZK15g+mf6u07CzgkO2q0R3o5mXj5xILKRoIHyotnyX4sb7SYtSXvOdWEyo0sE6EHOIHSxfo
/ZqpOKY5vx0HmuZqkGrBNInBSCYZ8O0eyHr7FWXGLZTJsPWl4bBrJBqJnUnuD6gqGYLufcuFWZqq
WE4siWCQFn+Za6ZtoDH8ZoZGbzSce2f4Xfm+ByFg3O1V05rn2MYgyZxq1B1yCtC4HaWv95U6LpQL
+bJQa0gwn17SokK76AvQnI/CenhkwKO6jvw9pk/yuk6cmwn018/CTPlhKUKgapDkAk1JzlUM5jpk
OddEZiGVYRa0cGBXGsHLRvJBuMq5oMH6pSCcrbFZytrw3DxpN6ysK/fTQ1BaHI63PcyV0u066C0w
Fp5HDoox3h4nn6jldfe1kXL8HJIlVPRmul7RQMzPzCYZdQhdB8ZOqL9z5H09vE20RWUJW+ZUODHL
zlttDgwdcZXDo9QR1S9UL8jQ2r/hXUl0xzSbe/+NpT4TA16JZQuQQx1UxPXIm9PA94ivE0XplE09
2e3YXc9wbKQIHIZeaWC4CA2gw62S5rgft2K7Xl6Ov3ZjefcB0MQMJFxy9y/By+1sJD2wrbILB80w
HRCmuUQjtWJ4DfPv2Sr6tART9jVxUPby59eAAQAdP0EJQkpmCYcOj5XpVnQ388OL9ZYTt43I+ASg
c9CihOfB5dq0Suzy98rYq2RW+cqq4CNxq8UsU7lryEgEY8kumsUkD40j8s6CLUw7TyBGx0hUuN3e
E4vVURCE4lZH4xi/0ZVD0HNpyzs0N6D3k2SvYtWF+VKH0SwH7F82thmFuiXMum3kkAi51AayEZSv
WFkFw21v+5TfImWh6b/gh1ETNOIAqJYkjPGluuB27hrKn+V/zm5dpB5pSBBt0iXkx/p8zUgHDxsm
3v52cN+kKG23EcC98SfC9AxU9bXaPu2A83PpZ3SfmW7ah/1NvQpDPDVC5LiondRom9sNM5s+NhSl
vRAfxn5jWcrMhpY/PCrMUa8fzVHm41tZ129FD4x9kcQEQYawpIzzGRVaMB/xXwoy3M7iTvydOkPi
BXoBtuCpnUOFUqCNPxgCsLJ6I7joFlq37IdUEcC+A1GOZa/2UnryFzN2pIgg51RTu2kCty8/i6rZ
ac/KEYiHOYC25M7+beGaC4zeVzFShlqdpwZ5bkO6niq1AZmb7GOpdFzhnnPowIhBzwetG7a4pTF+
IB8B4Mk1S3F/n9n1mAPpQbuE1QDwdgQL3i97TjcUhtWGZu1PJgb2TW6iO6zbeQ4z62djD2eq/Kx3
Ol24mev7mVe78Nt3t48GFap4Sw49rQ1quLIBlVeQar7moUUz+WEqqzwKcm/vLdjPAMWcZ4ZnkD5l
USgqfcO5wawIjFO2ydggxAg+BDEQE6i7Xer+Zr0Fi3uxAqST6kETYxC/2mhPZb97FJ6RBkIo7Kti
L3XHagt4wl2m+KjjlshlQuHJMxGYvVe2K/MrpBRwVIu0x52ItA/wNBGwgwv33Byh4bG0UhnRw1GW
43hrJQYOJKu1h0FrlVbj2sMW3Usomri6GdgBtec7dwxgfeZ1qmuqYRdY7i+avgkifxU6ZGcUFh2K
0mQ6C97hATFGWKRsoK4KmPPXQI6E11CIkMDgUybSHjmio+TvKZDQGv37v/xczCQHGVXsAY2diI6b
7AU4foBR432vfbxDtMg6lMXO+x29dFlecucmurcjIz0UXBlqJxy8tn6HovSEQ2oyOzf2bbDH9930
OMniX2cqnWbsB/944/9HJ4xErQgasjxybYXLXyHXByBIjzCnImVvvEnTDxsCXezHGbo12M9wPH6/
b66ozT6Kg5IALBkGuJtz5H6a7DsijtpLEixtFcE4KsPDsI5LFi1FjXmvHH3xwCR15L5ouKdsO1EO
hwgZIlY5k1wOGGS2y+s+NoQ5sk9HzlLsndGkSf9a6ELroZKRIsUAvRUvxfPKMcyX1a1v++4cFWyY
D811Tftm6+23Ho0JBDjb4jknb2cIWGE8smqb4Xy67utc1OfoqVYYAR9Erdz5MmHUJRl5CPgCeUlm
5v8q3w6Nl4c3+8zdVM3xFh/NpwtdfY9ZqrrL7KVYQk/N/iN0PAHTcOn78pVmceI74LW9r9VbeUrK
kZB4Ze3kxMCgmmTYAM3/11kxemeTngmE3ws8GkjOw+NjizBlIlHVKffdNPP0d0nVG/l0CpSHPzJE
bMG6eMJCOi5uCyFiFqiqZM3dK88MrVeW+y0IFZ8mRYNfw+dXD+MPw7bIq+25was6KvYUz2Luap3I
59FPJvcktlLZ05xQRUFsQVfgY+MNrPR0XRf5c2m6HaPOukHsZgIj21AQT9YOwlrKmSKM0I1oy0Pz
9MBSu4xaM+JM3lU/ZfiK1NBa7/YYLTzjOfHfVqgam9Yf8FhixY8XoKZ7+XBhFB+5qFHNbxm/lPpH
Pr3Os80lez7RPHZtaCJKVSZn6yViwEP3ACvaW3JXPRn0ej1xxfrYMklCBkIdj4dfBcPWlJu+phpv
x3zEF8I3iVSTzLBnHpeiDw0y4UaVdp60xUWrggbnAht3mUbr2tnmULjvZqLs5WtbY+vrJ3gadYSV
1TQSOhX68g9gqM8/JbdSoBhpfTjeg50am70Lv5phIyuaAGh5ojkE0X/TbgyanaBj6v35cbrtDjsA
iBj3gVsY6nI5rGiqbnQzeOO4N+vjlFPN4xtxV3iEcclUDztmHem16gfq4HK10WQpI9sReJH1MUBn
2iqVfOkALq0uRfy9ukf5nsqyNBmMPEAjrYebDomiMAYfYl2r5pJc/Qr94OtU6F17IkLbD+5KMz5k
edljmi6n/8p4hV/CAlWhr5PSbMYAosJY5wC2vpNsABs2FgvXHJp8f5evUsmnkaGsWWrmwumJ+rSy
2xia6Q4tWNtS99N30+kcNbOSYKHbL9vwmAQO+i8iMXy6CUkEIbMqVTnlOSHnzTleSu93JpaMw1R3
HNp4i8HzqNHWn6ZFYEyME2HLyO/Txgj/oBohSbWBzsl0IoblrCT5hZT7scAMXWzBHaEYgBKV1ziK
UvI1cUbJXfovitigVTB34HpTrltK4WW0Rawd5/hlV/yLiGw3Zoa+0pTqlVjBNl4ykZLre4Xbxph4
+t32LPSFL/3Za1854MNRaKhPSVuA2UN29ekbaNX5Tv95rxVAkebFDJiCwKBxTlvRDmB4N+hQhefv
BcXtHab2Bwzy3SWwmDmgbnAck6TcPT8Hi14ls72cPWtVqnXjMlGVapWa/jI5acrYktr/LEmywq75
FJ/0vYWUXnmyH+Pm0CHzZv8dJLX8+ls8zoSzomF8ylhd9aItToh09WzahpeVpYbFBWGixdWrje3x
HqVvJCmXpXfyn1mXVz6ioU4amEuuS4X1iJhVhFzbzEGVGUvXbJW+qQ6smKneWbvW8wArS6Uv/acY
1UTEmh+IOGF/uLrnH84RtE3qskaZtU9eOUod38CFnmw3PKoexN7FaXGERfqbP2j3vOKadGyJbmR1
fS1I8utmFcuCLFNFCWskHnc/DihLCUhbRhrYHoLAOMXjDcPkTtYYqep4Adt4Vri0XpOq2+8O5bSu
uZe3BusONB2oz3UCUk5pG3szamU1oeiOPk+oJjCrLL0CqptzZ3DfJUHlTzRz8nLwYugBwMbieVQB
5LQlCWo+95I/V5m4FwOlPuCqb2pq7TwUOu9LiEt14aZImuv6H2Jy2RJjPzVxisXdAayOQLmwd6Gn
lhrAuoEMxiqyQ04/BSF4bJTBLlkvH4RHS5UBWEDIEISRTq7P1/vf4g/mLh8zlhEpxzfso9oO8fX6
UiH3Y6Nef8/IC6o5399+dhajtyh7Gim4EOmN6FCIxlEhq8U9CSEVW4axU2FjyAlBbCCzikcpAScv
T+yXGyavVvq9LvKTYUSqf6ncEbsoCImbIg0QFDpGPy/BR82IwkO9w6GL4uoeE5l15Q31fmYnVeFv
wD8Yveu8XsPZSihnu7viZvxdyNfU1r/uKmByhHcIfk+Ra0+T7fLuvkBE0ZAlKyVdgZ/4AlhpuCX/
Udc0+3iDQYjrR6qMzOXjDSmpNc1oVrahOWDDCdyGFV4c1dTPHW/gXBAXfSWH+2WAIHvUv4mcGABd
w4rHor3c2KiVGN/MnXyjv6J48KBfwZLcq6he0f5Kou5gTBrnoGP+lMQT3y7A2fxrreQUKJmAAp/A
J0uhXe1flVBNqaCd9CySSoIZQ4nUP2ZPxzc3U/IscGQ++D4RPXELNfyD7T+6py8xrNWrXISl11EK
kGFOUmd8Nab1v9elJTtQr14gUfMG1NYEPwSeIwjAloVogrbc4Mxy2yHnCcOYhTwD0kUY4OlcbSWn
cvKcg8+XsGqaIFQVXXt7d8pBKDVPG235K6kvYvAtCSDWf8/0WETNWZ9OZ1MdRIUF8qOhtqmiVzof
zE7AD264GIl5Lg5I9fCtmZ/FLdwoCb85NxGc7/HMKSgiZ3cZ0sngxMA9AJ1TPspSAHMsv2ZVIgEe
EiOl4QEGOcma/oZtoBsXGpcOsUmz6NejSuu2yJAH/sasP05cuVgOn/t2otmbl8d6QHiCoYCYC8AN
h7qrMOc8Jzx9mwJ8qg1G8nO27Urqr7yJE92P/cpbgluZB9Y+tmOztGa1tA9lFBduv8V8nse4GCC9
xfeJiD7nn5ICc1ZxXPAOACe2TYtrZ73oNhayn8WSsCCndUc97tKI0Hnza1TzUC+9e5FfKpiQFsjb
Bg/mE7utlV0Xu1vk0jKYAWcrUWx92s/Ui1FH4rS5X7xWAsWdXMjhZdi9EyKo0JDHLtpD18u89Kcl
7WPaXbe4SfH5dRQuBL/PMyl8e9UY9Id41o6BxiCk90dmc2JAEBQiJpMl1FZxWgTKpQ1AT7ozBScU
TSY99zRB4ITzXO5nxWCw0J3ZKAO+RVvatFkE3FXd9+Dgt1krdAsATN1o90+rZaE3YOXuRiXPjLnD
BQa2xsYLsk+WvZyUnU3djerB7dybE//t7oIN9ZyMsUhWlKXYZsoWcaWswWcvq+9m2DJ8dDoEuNh5
4j880ZvrzzdY4tsYkwMGhtosKdEBrMCFF+2vPlT+zoocAs/TmCd7aim8IK2BGsQVHy1T7B3ZS+mL
ZZMQayZA2WZKjVXkI5vr+mgVrim2nw3d9SoHEvl4w8A7B5N0ufV0rKZKOSvgVjXHlvUtxV+Y8o0g
2XszNWhzqxnFedjXtcQeHS49AoBa6OZwr6vEAAzTfVEU13/ErD419oRFpLo6aX+TPGeoZpGOkLLy
4nRg49bLiIy1KZkIxNUpv2L+J0ek08dkjvGVVy7kMeTQcaXIoBEkcTUz1rbHra/U8k4M3JehNVWP
UY6r1DS8pJlcBi6D8uswXe3swNLut94loIH6JoH9cCqE+vafloN5KEl4vHpFGQtVOz9r1R++0XFz
wEIqkerU8VJ4KRXZL9UAOiCIbE8gubtbyPXLuadpdAxkFxPQ9eGeMaWe76KZ5RwsaIrWoEMZ7Qj3
vjZv/uF/00qqNoODg/+Obd9uEsVyzL6avxjgLLUPS8+zcgfvZ4jCdBtBleD4TsX0qjwVM5vi+sNH
o2qydqEH92ZlA5U+lRYkUlCZSHhOl/lA7qeXm2FpUxReexjO4U3kHzIx8CH0qTIBUk5+B4YnY41G
5RAhJpiSrWO0dcGI3OAlpQuCrxziP6pj6R6oFSTD6ZqEfpNCIdudixfPUwM0jcyYZhbd0CuVpYC5
xCkYusfjDCI2DHis/BHVN2SjxSA2QEYIc3wZcRtIX/Pa//ZZeg//rgIzK2GnAHyTpeBH9I6e9x72
8FBvjMcNWMLOWjFXXiUz9x1fL0TKKdfy65cYQ5h2iw1EiUTQiNPKTItboS1I6oJDmTXU6rluPCFb
Eeyd0IsFOBLjmUqptRSVc5SxbPYcVjB8ML6sxd9vWtpjAvTANu7N4CcFLCJNTUTyQBTftwJCSHDY
vYxgdEEMUseGbUKQV5tD/uuDNp0o5/vNuCTnh+0n3jCnyQALb47fP7/4qd9xncUZ01SeOprC4YuZ
Ww2hGWRo9r/Y/3Fn0GXuXEQo108b61kK6nOfMlE8Xhi2zbqyHmVVfEDj4iuEEqZiXHEaxI372FQr
paDSiL3v0LAktNHXn67/Vbs2+aDAOOCOrDdI/FBXVDKYMAdctCbjPty7F5uH/cDtK5P6LK8YKOdX
eD4k6uhxOMJYRg6ku9076G85okVeMUvint3uyreFhng+c1maPdcby6F6Q7e9eOvLzUw1z2ImF/YZ
DvetBSuZk2yF2mIqq5zm4Aet3kwgnloeBeZVfRJ8xXIQBL5sIYgVjh3sOfmVhrNKo27mjn3vxR/o
1Zknp+ljC3p1Eke5R1gPgTOK+pih6rF9m20Rjek1KBBehuK6cfjWQWamZwRWB1GgbY/11gqpuPBE
ttiCKwiyE0sHgxvPAszh1Hz2eP3QklsnA2l953IAej2hrCa45VFrfrz3HQvXq8Gu9fmjHPhkdtZQ
HbVxeoxnIMB9nRReqOrT8r3F1wEdQsT8bOvLHQv2eAhS8aTixg5ZMXqYh2+1FuYk34k8N2yQxlrg
qg8qn1mlDQ0LFx6bcWq+ySuppQ3gehTwrErE7QWTfwtxVCfGI/0+Uw8AI8eL8Jzu5aNvxofmBC6l
TqXJI3Kz3tdCFWYzxHahmG0lo7nmTzGD4vT0roDUYA+JyihOClsAButffB3JLAXf5u4IaILM2+13
S4OGWyeOIisPSSYPfRhzDiGQpLr4Hs01viAngBI3idySEemPA7nToYwm/1iX3MN/+pHJja1WaJ0J
f8VNg5i+4WqU6t5LfZu63AICsel9pSgchHzHUn+5b59sHxdF6iF/Hv0WkDvvabWgCNkz+ymy8v55
sga9omavjlPKlBFeg2p13aNkvwL0Dxu+JDkCSGiZ7BYEYKtpCo0tjd0cKIELq7hXh/iELv8lwq9N
ar3l+g3qoPCYW9F/TLoIN7/DdrL1EoK8Z8BaEe3Oy15Quun0OdNF84EaGVRQiFaLbFPAWaf2BlyR
ofDOeniLsLEWfRJMiWcbQnYTjvDrlhSgqRuDZFF9HXgGFgL8mOHm0i+cR+chdWoKypS0zKL5S6Xi
vL1XF5PlYGEsu3sg95iL9bbyo9GlEwX3tfGoImAR+brL/A+IX+3fB6TfWMHLnw2vzH3KyEZ1rpXF
lL1KEZRK+nIpS8Ata+pYeJPpr0EuerZ7Ksft2zkowZbj2aGT5tuNiRMG0b3jhAjAlEy96J9FVVSn
O2ah8L3kN07XhGURyT7DK0ZqU+ZdHhmDZ8q//4pkcbSU+nZdiGIppCyWDYWa70H15RPSC+EncJwu
Mv5a8cpUIHvSJMajfp0ZSdIMmfBnoakJZGKWpfeqqKpkkcLc72YWnYhRWCQkqRYdIIoqO3QOoubC
F3Ecszfp/Rf9pQdyAOWZrfHEGiWNcQ9zJD9xKMCtWFZbU0LrbTdvmNpdCpd8LsWbFVr/xkJJG2N4
4z0NdVREJtOHEHzp3dzQGTmi25biH2sWyDV2ZYgS4hyHfKfTRKrvn836FO8zgGx2ZEqbRaf8wkM1
WjLI6ToY5lE4f4jtC67vewPcfiaUH59sXsyWISNfx4Y0ZegLy45GL36bXysNGm6DHBXmMN+/tUKq
ixRZsU+FpoaUpupMXtLXY3aSHGLGcb6QLehBU70CMrgGozu8juDYpI6YcCxpH0LUR+6kijEVsnjm
NJN49RQkNjBy/p9OccNjin+k0XUi5tLiUrieDu235g+mvPJUxY095uaoNx4Av79vV3g5IRCwEury
E3AsCJPeh0sPyhrSUxTp959Bhlgdx/dTGg7nqwe0fDz1wpffDtGdmhTHN2fbCuyuBcWmkZ3ig7nS
6w8rF+OrDnbXx5pF7CiVt03uibeSvwFO5llTXlzd67Bh8xpedvrjA2m0Gz8nlYISniJOAHZMG0ZY
PpC60StZM0sGRK6HGy8peVBBsZa079CnOIJdmU6wfM2hQV81hohQPeFNt8nRAovoeXAZAy4RFgHv
3KKHITjKcxIhbe5AyXeysn743StR1fG+fJNlQ9uCVaZ4PObN/ykaSNYfof5PjR02QN/qlqtbAGY5
DB7dU2+OS9kuOMgidxRGTZBxUCwILmw8heQi7yRzBf8rGfBbudUOzYts7xUEkrAcJDcY6UhZmEpN
5V3FYWTQj0mimMWIxXZQpleqFGOSSbeu7FFVH074otTp2Mh8j/Vryv5VsJhitVM4jkfITpElsWe3
CZHmUhPLAcaYqLWztNtyXIdz3n4cwfmVyVYkj2vt3TpNPGyHlvSBK2mE0dIBH5x7OXGMJ8fyR4qp
1EsjcY4KofqLycj5AYZ2qWWqje8glfYMv4USsKcSkYOlXa//Weg+NkOg9Nf1v99ANG448nrzG5to
vp4uR4F03JTyzlQlnBYFH4RXFapOLPD9JU7LeKnS259Yy5A6C6Dfb8P6jwaNrALI8Ia9NXdOceeC
27m4iAYg7fBQb2VE9dLPGkR2QyZ/g5uZbJiu8LuDL2Fulya477AgtbhSAM1Ji+uC9FoaNcxxreMZ
Xl7x/TzDCKngmE+Gpvt6zRBAyyohbee/IilsWYKEmgY3D4M5VIhEOSGAQfKt730s4ZkSvbnlCUd6
y1rT0tBB45Pmg0ZqbLzWAYEAb8Sz1EbMLia8ybFuMwqHzOZhDBsAh6RP9NJdAuD9aXNmk73ngF0d
8hZrUYmd6kriRFEye0TWmvKqBcna8018xP7MWlJYQTZvjbElSkhUFqCAcjxrxh9SOYrSVhei2X2V
MYB2sexvUrvY/sIbAtCqQBe9GhianwNPHdPsoh6WpfsHfFlKeNVy8huN01heHayiRTe1CSzdtywa
6pfBWr7+NekTZBX7oehgC2lDZOwMYj7qu35UzxcKp7PbXxylpmnYnukkYoqfrkbp5wBI6bX/tMXQ
VOm1v9Eot+wkBDIzHZVUW3Jk+WznhAnzjRvKI4NBTNNnoz1gIUYbnTk9LFsO6KKG2RR7Vue6NXUz
IJMxdl7aR/QdaWkWueggKc0g6UvXK32nt+Z2Q3dcck+ut24N5H4fD9EQhwBZEXAcBZxhwK+yLsGw
7GieqF0ipLNe3cSzlUSAKL6YqmCSXRzR5U0zXPHQR7FnfMq3ylaaQrk9HOlbD1jjQqrW52tTnfuH
QiOTl9cAlG1BFR2BHpPTTGUJj+Ig/+vcuV6RgyVAxkDSNbm3x8O9gj/ebiLGIcQXxi8cFtz+Tk3J
1bgTzMgDraNAHQY6eVRQCqfQXuCmLe5vD2ZlE4cLdXg2JNlciLtC3XYv0z4JDwqy+xz16BSs3Yw7
ty2NUDoJK24tjk33jiwa0aPlCF1W1dRNrZv+lltdt6eU/9+HFPdXk5qOKV3BxraSSiGX2v2uy9dm
+XtSLgesIBXN0p/9dgKlckaBqeRlvwAWB5B96DagYgMz9KnxWbiL1CcDeBbbWZWt3WVTHnbsi0ed
rH7OIZZqHP8OSMzSRyExmSnaCskgK6P/+CRfolitk/1ebZMU8qhAJdkwiidsfC88/BXGORUEK60z
bn/I0fmcJBD7DqvgAVWKltQj3Y4YspJUaYo7H2KqyF19X1AjyikKvwRSNgeeGyz7jko9E6YTPfT5
1J6ecUoCdMdJl/uKr3Pi8iJNJ6lZnjUpLvna3gpxARgj4Pcmsepuad8jfK5Kj5vSC/9+O/igqPvY
+8MzItLn0R2hm7C0LPTZf17JKH4j3o2S0o5C7GOKQFaA3dl8663kr6FzvpqYZndKjtMcRkN8E7Hh
ggLoaAHcPj3eEdkFCQoZGhDCBSENTx5LOTO/jP6EDN9i9w4BNciFE/u7VSQZGVcv3DY5KGCyyOzE
9Wat13lxgZIy0d45VQGvNWWpYGTjX1dlEqBFDjihEgeY5AxK45c1Jz1Qe9A8e1InoUoVbxswC+vI
QKxNBfm3fx2L3CgBiPxrlelGUcgx5oYnNWC/IoUZF5IFhy1Y/RyxNaAuSNuJq5HPpo4qDUFe6yD1
8TlajvIKteiYW163vmgyu7pNFtg2TiYufp+UIfyVQx/z+7u8Mx7OdrabEg8vCtL+/TiHsY8RYNNl
X0gHZHQ2isVkw41YKAbcoPefhYjCcc1th4VD0dY0xTFc+iBlbudcu8JuJR790ZX9JEqfIjEKEENS
sr2+yNktfU8Wq3tphiXcxISQ6nUv/836u2AEW0idWrv4kEFj41V+ZS8CvlSYje6BK20llvqQ1Brz
rMpK6whhooV6pNqExqub8IFxMOIJ89+GliFu7XteRypuRj6FRQvkCJP8cWyu4m9b0H7vAbxUO7BT
EIqquR0VUJ46aRTgoIxsnGnxSW0jxH4tLLDJuUlg4Ceh8cR1l2PYEmg93BjkV8WXNAYXZZ6eWmgD
hFFATEgqkn2OrYdvyST9g9xhNVRwIBoefWZIjHUaG1sVM+JQg9HkFtQpE4OrURrVPyZkR8RDWIYF
p3GZxaQ78LqCcQgaWxIQGNVHWGyE6RnI6BpDnKG+q37ICyqTX5YQGVxTzyyhhtzTaNBd72tpE3Pu
hpJ5smnfiBeL83yCk93YQY0lh7tMhjBwn0BxlrtRnN+bqyEKQeF1UVxeAfc2k/RDKU58pbHyydX9
1402hvtqWQVVwnHmGGZOCRmSXLFIaYijrVC93F5A1JZhXGE37lE7dlX9N8rnkMttFrAU9TgEHiJB
FxciyepggzJw6ygRsd0Z/3AQ/tcPVxW1wszT6b2cnngTURhNegZWi5ECyFpijEdVuAnw8Aqdlg90
Yj/rRrvcwH3UltBo04qK6OSQkjO6pMUfiEiQGP5FUKw36XB3gNEE0IpuSHinbr8nupy3CVGeSn0F
MDSm7LziJV43yMckVYlJK7vQCa01Rnsi4QVu8zmI/2fOxYUn5o2GCwzM3JaPYc0u7/aKBEmT1nnM
wf+E3WU+USrTWakgD8b+lNjiH35qEsW3g4E/hWHEAbHkImE0tnQLPtN/uAcCxuNWJ/RsBJ8xhJb9
O836PUksdCBtqLL23qeZ4ioati2+lpjypSt37nAyf4Q1nOQgLyU5WUiUlp9iM3EsFAO8qj8eUUqr
+OhilS+mNoPpNRR9Eocr66CJxn6luzeeJfjflOIm/nbv9KFC4LzL+2DWP70yiVlj09jypnC+fk8J
9BWFDvCUx/7uUbLVeDRuEiRX4c44zolV0Vzicq+NiztKz/GS5B6FyeaV1AN75/Z++WoZRG6AWbAD
8fWjTFU3GM8MxiUPUWAuXljZOb9b/pacyV0b/jTFGkxPxogRAJb5le68AEL/lqv3x6auRpI7b+hP
z+koE8Wv05C8dopac8ID/JJP47ymmM9cNhDcxslymiK5aQZ9f10GGc3oat2uYLfUdtgRt7vnBxXK
F0y29GvEtN8tC6E4Gv/VwSAhP8aDSQVinwHgMbU2fNCzHVfr+h9IXYdNkY1Jd4yIjQWm8CYcFvEW
8OjfeQ2rSqdoNujnvLvUdsY9vc90Yr8rUFprcDlt3GIxjaUE2ITv125oGaXfH8iyPXIx2W2MIiRa
chL57iy0CBoUU+yLwQMrOsrom71wXfi4I244JLkyKMH47swBQqEKQF/RzLpO14XsXO4ligmNh3CQ
cYtXfRioVWfPzXSTVpjO6VjxyqTa8ooroWDI1tb55VJ3x1MqUk8SINuVxQvY6fD8not2aXZM1hVu
/UmOLO7Y19Pgc5QhqSBh4I6Im5TbGBkOCKTCG8XU1U1AFxXItaPBRF24HDgelWnXzVbReC64xwJB
+2joKSWvNseWY1Cx2gSEnqH7bWTSz2lYKbaHQkJr6jb4tRWD5YAi2ajrTDB254ulELV/i0lGd7sm
i7kePWTW2zZuALJtVyBuuZE2L4md7tUp5inwYLLCKqyixuz16oPSVOjaK4qUGWlwQ+OrpY2ijN9V
abGd9h0pqNVIgCLrvaWmOYOx+5HrV+IFNWbLre5zHo0esoRqtiKHKAvGGsmiNzwfeNzUZ+ogC49g
qCJmn5+lFCWynVNbsUwo6OWcPpUMCKBCLVlQc0YLtjY1bQnTvC4Jij8reHV27cs4o0WZ2/hAXsx8
6KKH0PQwq6UqL4d+qZe6WDylAWUan3tzz24QQbqQMwYE9hUqaI6U+m3RaNBRTv+7ZcL7+ulxT65x
qEC0xiWxuVfpHy5VRft7NIsHwzzvsCZOSD2c2iIgUs6ltn2JB6RJi6qWr2i6nCtJlpr+RzNbR3uj
RACI0eC37j5SecTEJ8C20IjQjBLi1jde6lljhsaEay3K1aDbnvkusYbAn1IUGRAEXy6lCBkFT1yC
V1FVgXZF3ySOvG/uEQrTAR59pLIBnKKUFL+/9kHymQ3m5DOBBnqaw/gActYPLqXGKrV53bW9ti0K
HMLcDcnrW5MXdiOMXo13/HABADJpHaZdhoPoJZIdfnsHpay/o9Mo+2TZAfH3VuWhRjSFIJdI7J03
AlirS5f6dyiJ3jdIVojXoIXv95G9xbRBJksI607zyVQ+GNrcYvncclN2qhBqxGex6SPC8cqrPXiD
omP3He9ymY/x4eGl8zgCnQj/QF+83gFAj+BIcT6m+OEQNQmLVVqpsyv4WbiB6QxMhIGBlQUJrxuS
lW6bAsrTGTHLN6RUxATRtu/OrraMc5S1wx1RzOW6+vnzjyd7IgMkd9JNBeTMLs6DjhSrFgirGS0z
2v4RdruWNLvt9kIfc6HvaP8KWwBS4ZsC5YBQuQOqG3XWEtm2IgFC029oG2zGDR/ZwzDIfsvNuYcv
sJliRWjjVq9Z4x2SutcmONmfmRQgDXEH53gywEX0ADNyTnNDZArO6dqzYKrrITx5OKZfQrHUhMtD
bsjxXiRQ4fv+2ZqUuGFz6q1364PRJTgIscfRlqQD/kneIh+4Q3V+kDpfUR/la7FBfLe2y2DY03g9
T5sv7cODwLeIiC2ITD44aF6xKhUXh20UqD8YSJcgmAamBhf69f62iB5PVe1ACA8pTxFXpiIhdVsZ
EJq99xcWm2ALsdfzmsFbY/LAYnPXXp2gEGTeMFeG6hJLqciHP7Wzmr6KTUd8NmBInwarfUCHARF+
uKSFy8bDygCwz5rpFPq2brhrkZ2PyunPyEARrEWnk5jNtXc9vFbpxiEtBHP2fJnAO1h1W4wd0k2i
CIrIq8j76jPEdZQrqrfZwcwm8b9BTtYOvbrGoi3T0yn1qsPqGaK8412I0f+Uzrid8Xrnp7elH1fi
Lb37YLQOOKg4ezsp9tHqpubeFt+xHw5Km2B9u7xAuRtgkemfTqhAZzQqOHsfkjqYvMa6R15i9VdA
a2b3qd3jWjOb3hkP3hJwu8xz8rAEKcXiRAA7VsWG3RGGzqKj3ZqHtKshLCJ5/kFSxQIUbAsgnDtT
yknDE8fbbvu+SJjOEUAd9/TZ0dcevXEyp/M5A2n9pLwqNXRQEdjJXjxC0HG04Q60t+2DD+VHN+Q4
/p6pSM0xkSZqYUbtCi73C+vLhABAEbxL9NX1MZd1ESHFYKuz3jvjKIbeLq1HzKtFgkBeR94bvSfB
14i2IKLq2CK8J6wBKu0OrdvttyP+I6MTJGL1EEFdU3pdmkIShSGZ4neZz2gFSoJxEnpR9xnxdkoQ
ebZ4Bdna8TLSEOq7AGTWRwnK31/QJjtq6QL8V6f9JbypT7t5Hl/VCUxre0hMFrSSTIqMUYlPXrI8
tJD0trBfBuDImd242VqVI7sOnAe0sOoAl810ev6wKbDRKzCV5+ARmAQaUmb8QJmeYyybYzuii90g
4a0JZXcGt/x0BTEQbYY7+6+GqQMKiDSdxclGNknXOhE2M/cWH4uF5dPx0nWL16yNUSOa6fEVF8Mh
eEW81bZ3D6sHUej96JBLSfSCeG7YTPRrvHdu6GVsIcOUZjbBwUOguBoaDAeKF3YzzQy/+UgcUlzc
fpClSlOPhPqM6kPEa6bQl1w7xT+XKLZDtvRsWVwPSH8KEkN84VkXBKgt6LBdEJvB6gcKMedqIEp0
FzNeLZjB7klGSfRYxdRwMUJswcvUaOtku9j7n+bfhsZktuMbjPp8wc96VGun+GDmpzhIAioeNuXn
GnVmL6Hrl2wE1xo2hkMCV4giHGwEYkyMZpZ6gKqIubbDSSZDbeVrKBHjbQ1opHqMCQt+eCKBhDGO
qXMlNX1ZZsZIsQrWqp3jXl73JRotQxhwVM0uENA7TlNAA53ACL8KKSlE6dBtTEHCziD4s21/FSGP
qcFKuGAn8r5691F/hgsuHbb3nQxMT2quiNpeGfyNS9iDuYVI7HHTgVxJf3MHKh9IGzZcNfozEIj8
rdV8KQU5HNf2yIPshwiKqvZ7vGR+s8EnmFW8bTfgzjF5uifCjTPkaihjb9P/gLPv4I8BWjbS0cTN
LyrlifHo8Otv/aGECLiNaE2B7qVz7/O1zsZM6Jz5oeCezqoPZMBTnduQtu6COgaXsHDGRQ3ABx8T
9lYNwZpS/CcemHeXvHLajYNzvtaeM2tvU/Mf1kscb6cyLQTNqtPSbPtIn93oS542yJ3jo05cY0+y
8cXBCen7JhaV+thod9jeOJVILN+NG+nZYV9D+IWPfiy8d4jDLCR3kY4w8MrfdaOMguFqpgFuPjnI
TOh0MEqHc43P4ullfC2Fj6UjOhRM4+Lso2XzXb8l7TpVqIeCgro0WZkbOlcmXRY2ohphna+nWQ3K
mOXgIvpyZvebOjU9rtL2iaRwz+5QbEdnHtWfor1KvFcTJ8Rc5f4QFnzoiXksdf3MU0LN81r6WApC
ARWEse9rXrvWhxRh/SLZlhWuOoMTPOGKGdzdvKW9UJYEytyrEkwGiGo+OOABp3EEjlq1y35Tg1w8
RuOe2pqRNVcl3PV9mQjOMLEDaxHKDsbgct4Vvg4vqBOi40f8eF/ScnpBbWwDm5soquSNzeaNSYjj
SyNC5KpBdG2OdILCvznKn5uQ/5uSjFY7/S47lTe+vIo9uSpJ/XqS2vCDzwTtx3N+cbu/lUz6+6l6
hSs73EE+0cSQYf++2JhY8w0OEqpieNaL/4Oc/KututNEJbdYWV2I//nj0QSFMdEGZIeXE+p3q4vg
LayF/cCGaZmmxdz38g9B/5SnyPoFG8jrTBNH1uCdzKqjyjYAHBP42ZUd+vJ9aO6zCT0dr02m+u/o
Hwqrf0rml0n8a/FtEZP3ImmqxbHII75KVrIe4qwMvf8uJMRrbJsUvNKEaigFLwl7lHo1elOd6gCK
sKvPe6egwM20k+toI9sHEWkySbG3AaJTrSOFwTMTBftdml0DlvwKoEoYc8kSnL973oK38p6th1mp
abIuM1Y5gND20qFFXJwyYOZz52kPKMrFGbj7h54nKPGl1AkMYMukMBEticvNSRYKBzw6ZTgLCz0K
cKpQV5m3kEKUB5IC7AQsTgkXTvXyL/e2DvWXD1rK2yiUl9GRc6HHfwtqVtkk5B4oV5kIJ4eUeWv3
rB95XLqdXtwla4csFGrOYmt9UP6mrHqflNc1SF9smhOp4GFqfSiusQDp8DaDABx+xJ102052BVnD
GpsNFQuaP3+65FOt10hkKTIBUZPh237K/qXowAKhwxWRsGxlfuRLgFmQchaw5apHwM/omWdY45T7
ha5HzoZcpgXVNM9M+qDPoRG89Kwb7sItFW0FbjO3u8tjt0+7l/p+jSkAye+Aj6thie1Va92vUZEn
PfybMPeD/rjteBzvU5ofmIWCN4Moo7rIebcuOEyABYscTm65pKhcX2sT++9S9Ol8XCDnKr5NGgg4
36RAQYxdSslqA4hb+4ZZy4ckFODL4nTKw/T5r1mz9vhkSunM9OQY/xtSWLU4DrC3QOJLfhg53GrQ
fnu/055vZBavqK8ajLFzKJR41TE/tfmRdyz+9sRlpqemXI12yn+6m/pmqNWK+Iw8CMGcRUTWfiag
Ne+lVsNx4XUIyBef0GQU8+ZhzcVhJW3v/rCWVMysBUhhoof3vjj8Iw3x6wt6fons/nn6D8ARsyer
UGhKAY2bQn23w8oE+sooa7nWr8UC8ShrUVJuzd4h/A1aslYiuaAprrWZJtn57KexSrk0X6BmW5kc
kj8uF+Y+3X6zou9EU/s33JaCLDGURjSofNvcrp9R14x7dIj4fY9mltFqGrAL9v8clqYAFtdI2D6p
Hf7feelbwGXcWla6D7QF7kZNAc4irVbnqJ3wtjadFTfCvLngzjSfphLvhONunmYxuzhLh0wtCVez
p0MXOzvkr9dCgjG0eFwVW5BDj3ZAKjAWrWjXMWkr9V2Z4T+jkKrh3RA0yIqzCc3tiHVdbnwEqTEE
8AslYUTZorkf8BN3LGmsbg72VOonjxDYyJRCQExb0QkoDmh0GpU8lIA2cDMaPmXgA8TIVjq2owYM
WUxYyrBmqhfabc76FPTfcISqwp4n5IOO7m/pH5gpRYCij+ba5Why8y6e/t/ggny+AYBrbiX9q/ob
JEwBK7d4ynaGKgiBiNz3AqyIEGnKY1/uaKwWJBnCGgbl1pu5N7YTcaHCLj3etI5cML5lRGSdiw/B
VXpZE2DwcsolNThBRqINMrgaKomhSFbaJshtvZEY7U6G0aLhM75lnJtJv3ow1tyE5EBy7VcvcYv5
bvI1MXoTZ81TiIksur8ABiCykIlaXOadNCjnZhT40vBb48EDfx+7lcavLS3o7foc2/0NH26MeLHk
8gqv5pCNm+SSu1KUyEbJGfbdS6IvC92L1DnThhyCcbeMJv8ecdeLTNk6DcW3ve9OJ7U19Y10tWRg
VghjhmxFVpRVMcP2MM6jbmk3V2PwvOFAvBPPlc/wS7RH23yxdM0CiJ0QiMlW0MiCUns76B6vb8Fc
3hfEZf6ayrBA5ZwHtGloBZcgNNhCLGCqs/qAA7Gq6mlrJQwrQR2nciDpcMksTsCx/B9A3486+6k2
qR1jSN/BAcKnOOEHtob0k+Wxllt4T3R+oe+fku8HwOFuTW6TUrMJ75TFsYpJn2kOhtv8o3LMPMCz
k11waXqw6SbX/6xh3aFdo97j29u7zgw4LwT8U3n/Ln0VlEzUw8//iw6f66NfRrIJlPr625si5A7g
iE08nZM0/7M89HQWNC6FuaJXm+WEMtMen+4CVsJyn64RCVIi5AFX8sYO4wTo8XclNCu8ljf7U8gp
Xgn/s6IWT7whaOPn1rvqjGaNmrmVw+022vsaThHjCY4rGioqwSE1YnheYyVD9fjSV/wRgLTcAkZG
cl+ymu5Sk9zc5XNXnwH+Rjh4opd+u12MZXgr+T4K8rUExMp36p5mVzpRgZdO2CHF1ZaXkwwGTmc8
0XmPpMbRUARETYOJxeNrMgJzC0pNmKGuWjeizzC14KTa6pAswR7gmZC9Z9s7E5RZoeakULXKpIXR
K40s7MpDzpZEKY7nP42pRCVLQYfHxyxapizFCKtKuUx9Dams/Emntl5NrCgYRnEWNvLlHNpGilta
YhB5+X+ga8Tn0o2vTOO1NFO2tkazEdl6oEU7OD3AQZaarNjLNB35A5zxWjpmdfKkeEhbB/LNgTAy
eCRO33Gmo05aYgJ0H4nRyC9smhyucs5NkW2KX2RI7t03aMel3SAhlDpZWZf4vHaHcD02NnuDT6X6
56lACPzB5wlR1p98Mu9rNNwgBwFDvPLfEKdf0+XhmmU0HdBkSmKN3NYbr1ozg0sqyHk5s0wrL3ND
wF7JL755tkSlfV9wHmkC2VmTuSv8cqiY7UARjkh0JUWITibythzAad9x9EH+7Ap4n/anTYDxEjjz
TJxT5jU3sPHy0O+tBTmHsfcbkx3V95dE5/ULE1gfUXrTaTcI06c33wnhll4vJCfgEsHW+eeJQWnI
K7yJMATvCbGbnKX7Ie2qu3s0WeXMSzrmKEhQIjAy8BvjdxMPCkcI9s0fzqCm+5kRo03LfNYQUxrK
IU2xPV2Yz4GRzzG7wrZv5wiiEsPl4P9rWOtYudtZ3OngKTFuqU5d0CeFUjJH8RJJhyB5NUJtXvwi
XYrHRdemR8rvb1Y5Cqg33m+Si3V/m6DId/tVkecdS/f8GeIUvuD6u0OAaOXhIwiG9YmQS71jZAnn
e3S/jMwDqP1hiQprZzV1eZCCUdgW4fEfUkW72D5cMymJleI6IK1miHqWAVhaJvQuziuuyNjlLbWk
Vveo4C4Wi1Q/2oiUJ5T/AsIl7/25jmQsKPYBqKxgZuxYvaSedj1zj5i6rmgzkr1dulZO1Z1hylqX
ao44YVOaHrIASvDpUhqempEsqkx3TTtG7MwjDljzNpLeOL/wBer1v7s27EYREr9qUSJMU9BO/4+z
409NEEbqadZfkhlPc+EC0C7FiL/MZ2TkKELPhIK/nXsl2KJP7thmyBkgX9MKl261zVYKBVKUGnuP
JdNeW1tZRf7ibF7zwNiddpaQ5OSiEKgsrdquHXINOH/e0Tyvzntjlk82gNB/PJPNGOEM2aDkdvuV
nvRRYUk1aLjayOgMXzNy80t9nVSqncWnFDSxvm3HIOMYIMCG0++iflx8Sw+/9IVK+ld8ATMxBIKb
Tbb6PB+gSYGcZbGWEmOeGovSlLT0yM8x93ycpagQqcXaNNi4FbwKagf3xt+wlGmfNCYzWbBmlO8r
gm8j3ac9H6569dvhb72z3+v5wvLdYLR0YTmreOyxDJ6npCNmaXhb4bGj2KXI+GClt3U5ZfYGjrHA
xvy6yRQqAnUMRltQ4OL56OszihEQXXJqbo2a58Ddck5kqeUQKipFmm7lDLL7Nz16jf2D4zKAlOJ0
gG9AnjbxXwdxw6ZDF1P77E+K+999WLE8GeMNuwOPbahtMohr2qxKhB8PHSZwv8ffb7AMzCcU160V
EC9peAD6PhXQHYUt3bkqtzxy4BCPe5lXAzd+kobm+lLjE2gGJmJIjooECDgQg793VnLFcRgxC7Qo
zpKBorqPBqWGiEycVw0vbNJSPmP6hSKFceSPZvyuDQ3dit+QspJptO9xl4OIG8urXnBCz4FN8PPt
Svnnt8tOsGZ27HMnh7EKsWZ74DQ6MG5MMlXrReSqab5VRjYAR+WpYM9daTusVPaXfisqJ21x3YAs
tFSHHKlcrxJcZXpCMocwYvPfAsoTjQajKocNcQb7ylNjvEbtPF+l7+dOFtkQYSDJq8h8mguMy/hm
1NtbjQew9inIph9ZWiNFMv5O4kYfwVoId0FLHBlYYkseYbYlDM3ffo6B+E+TUPtXs7LAFCiRQuwF
GijpIb1o8/B7FxvxNQdC7VAO15onx1iISqHI/UgtdWIy1bknLVfZFh/cRuIaovwiaCNR5ExlFJcB
iP9+ImPRb9k+2TLZrSxBwrLP9NH4Jlqtsu/cyVwXIuvkM8rzMjDAp77GPz2Scdp5jJKWuHkIwcH2
d/We3b8juZpgm+6KaDWK2z0lcsmS3ib6SjeRBHhyUileq4R1W1WmBFdoHXt7Rt1l/0AtYaKVySkK
c57T7lT2RHb7NJWCHt7Fd1RdmcRSk3QpE/Ah4I590hDOcpRfhBj7nuf306rUqnyuPouD931Rm69j
0Co5YwtyW2W37AGeG2MpsWZdM8T5DjAOEoe/WD4JG5xur+aVZL7citUbg4ak7UdmIA+3qKWjl8jo
AjZTNbXBcqDYzPhFN4w5CexnoSLAU2ocKcmsmDn/cgpGK/gI/hyfiXoqd4p1gCc8SiP7j0zIPGLL
8Pm3mxCYJiVYms3OnxzTUs0IPx/HuIfUUlQyz2fvOmOSRbe+1BXSSWcY2SbH5RgNJ4ojzOE+T8Wr
KNtkoKzND7Af6sqc04ZBuDuXkpzxebiNieLUHSimXc0B1tox+El5l2+cvLiSVaosksmw5IIy1y99
euIyDXVCurhtJs1bEmD3CEUXoF5sB9TezjHFDg3bTiXePB7cCu1/GO6Af8nHsptFz6wfoW9FEfr4
PemLfbHBnWHV+FQ90bwQ0sNlZgXYu1VzMPZ87U4Atn17+jYWkOsBbGAC6tG/dP8QQiukFaG9R+vK
KVWLAzOnGrLoHgppkRnBFzt4KkdYDstkd0fmfG2U/T8lus6YKo542eY3XvZy/B5wC1HzYbcshFz+
INNKNh0MHdqk/7qn4WfLblAZ2WUTkf4bEqlyCM/L+RFdBcXFDpC+wH7KIRi613ExoYVKjLVhx39O
lWpR03sa7OxOUaI+BBBmRn0JKESF3K+ftYCWFIP49DR4UCMyTKwHludjnVnYqE8klDg+pbu6ukcX
JG4KKbjVo4Nn8PHteHpZbdOX8lzSUF9SBjlM5LmJH6ABG9t4pY7h6HMO0B2jfU6NPE+KkltFRq3o
h0zgv9UmCPIQt6gQOjHzGwYdVG7+CE/XU2cuS4tVLjQpDsuNCEc/J3kge3eI2m8oWukJ/3fIlRtZ
+cv+GKMXC2yQBTN02PSGF1c6ZDfeeb5iSyR1+phdhDBzg/GoyprI8RGGJlKSXVbpGoe/CFAujBg/
XWefff6kDhe6vf7WtWk5XN6hd3sZ/L9yoDHpedUw90uW3p9kUl/5xFKYOW0FxLM+I8XgHa3Cg3vj
FUTwavW+6+1/Isk/4yjA+mQmvIPhehSGeMjVFoksY2yLOVuFNDdY/prLFANrBjpZ3m88koErzH/u
D9uR4jMLrQo+wRSAL7X8KtdNLkXqkNk+Oc+roCiPWqALXF5Hpm8XjWP8tSBTUKMqnHK1PyBnMsnd
BaMqk7QyNoWH997DPoCKBf9qwtA07YErZadP5R1vESyF8LwCHmzgH/rXH3bdrJNFOTv0RcwBbzkz
VyfQSxcXJb8gDHHAvUHjRiosM0cBetu0s3Q1WW451yw0av1Ok5vb/h0aFGS3Z9/xpkmY71p2U9yM
Ks+G+YkPuoQcyzZ8ykqnaZlvDfd2bry/c7zY/0u5npIsP4oYO6c+ot5Gt9IMTGBBNqyLu85gqXJp
fn07xLzRYcibPpShixdMlkm1ca0YM/CNUXS5oB8Bmh6CYmT8ePgfxOHLOXjsAgPXHZGmiINorzJ9
m9dtrTTaqDDd6ubD0c5SHbv9Hq7ScUsnxsrKTD03dJsy5GhbXvJmLJ3Aj/f16NFp/14a4O7nEQTM
XEFKF+AGojfF3dbjIcXOHpilEVH8bNNWiYsWOb2ylzvVG/ubQlDjgKBfFwNS50p9JetNtW0Ly6WK
SEEdHBGLr6cnBRZ3t1aZbqz049NMkcCfmJ3wpDjJCLAU1KoK5SHov0hJgT5XDSNkeYN9hH+FwYkU
oI/173ZCyp+lwT79CLGm+Xvu3IiL6SLTSz1iA9YAMXJQvghi8E1iFI8Rx4bfJA69Pgzva6WiDXUx
YXgHMcjJpsNtUeNo7ROU9cnhzmyRPubKcSFCVnbLAbklUbOFmoR2Cf0ihxu1oFawSa68qv728uBz
qUyVN6x8cmIul1cIPguhFbsY9CELIzgOaWDjuNsx6116+EPgU+E7Do1GYRBqKIywg0tzPMMywEQN
QEVPHMKLX8SXx5Ruy08hpVUBWIwG7Y7GqggOJ5kAgXi8g6RXsH7rHdqxiQwEedffyGA+0EfHKC+v
7H0g8fFO6e/2ozRr3zWTcC5vNb65Z5H07mXC5xzcIDAjMIuGGR/FP13pwyNRrq5PaNblcZhfpnfg
KJQyZIbCzGzWSDR8zmWttX26Vt2brHO2aJ7VHTiCZNWieWrTBKoxCJDNC1rwJ1MxqR4+vlFck3Te
0yrifSmRcMPoEEzEIHQZf2Tdqbs5DK3Dzum0V/WNc4Ji1e1AEhVe/OFal5+KDD0GjKA6+Oa2j5Ds
hAjr3WUXM24820lZtZQ0wRM8wCZ7UztXW1dapErzW1+/s718oscP7Btl25jPvrbfScQraKguUG5Y
TxLHdTQLg1cb+aIouC1AMU022NOqddDisqkNK5KXAV977ICilPXwH+yvJOl6DsnaunCCDM0nsQ0K
q4yKDKooBEVVesy9SEMfPmxGpG0K47XzLR2YqQKJl4xMvrEwjF5NzM6wy+VaOPsREx/F5/2SCr08
g5Uq78HX2yOyXz4C4wxYKTROxlwHAQFfNI5P4uFeas6/KEy+EqwUwIFIRSII388ZRZA1O+1tXPow
yNku1Ss37hNsdjz9z+jJUuD5xn32cZKw2+0aOQkYw6wQzCLXcZQonko8hdDOLYO2fPWQXDm7DFrs
KxVShQEUCpSseQZWCCkjarcQg87Z1CECw1szYD7ldu2OTCGLq+ODIQsbuT1pChup4sg3rD5VE4m3
pPWuMAlMAEf74Js7NJLZLZdZ3f3JS8C3aAmjb7SLE7r2G2igjXncP+8Ic3ZqnTKbRSQrTmQIplgA
xenm2dWjc02TShR3jhz7TDFwDHkvMaQEtGr5uPrup6YhxOvrJkHm/wGKLSslmwgJJcoOlDOg7mHv
dCX2eskh3A57toYn5t1et5lbcr91NmJERbAxs7dyDMOnuk+bQmGIc5pwr4D+POA4A+spTFQyWHhw
8PPtWA1NjSRDHpZmgWUUBL4IWCDYF7OkUKe9SI5qGFiOgmrlK6brBgI3n7L93PxYneXijT6Lpzfr
f219VpUGv+cFYjl/nZpIzgpu7VQ4ZE1ro0WT62mOU2Rrn02fjt06ljh2+guTeSuQ+wxmmE4tm5se
XqZEWWVTcQ/xNLBM05NRF6Zup0Dy5VnOPL/bSUYsTc1iWMPIdnR/iKKzVDtips79G3be4LmCIxQO
RzqMJTXddDj52dC5ogYhVW04l9p3aqH7CUTWeOU8Xpmdkxhem17LbF4nRQzbrYNVUt7sCFNQgSni
jbWEsK8kRBaMeVFx7GDbQDmq/MCWO3khsOWSTUuU9UnGaXMj8Z6Z9owVwNOxBjiLOt8dzpdXRtvX
YCJrv+O83ur4tNOVSqsgRxw6D2CSoFqymtxhh8LzgHSFvyv04I+pRFUulA6XKIjSeEu2aOYJETZQ
Xj4kl/VGWMu9ChGQwGTvkp8AT57GlXaTGobm2xw5XS1/4bB0A2FOR4P+SKXGP1oeCo+lFsvVDCpD
xxjJFkh8Fti9o5soyqS7AJ+BEmNwJ8uhp8RebJARxStqZnzPWBGJz84vSmjxH7YG6AT2HOX7MM2P
bfpktK4USgtAYsxBK+eyFVX1LfZbzrpjBrofSfgGBQujru8OkpTtmeILxQ3GpUw6TYgAgM0LpNFB
nZDopv2X0dECvocJE+EfvEFXIGngxHmQq0TW4Rsb+KvX5yVK77Eom6i9JyShXdLRyENRpkQEdT7n
U4i1M2XCl82VC6fFFDtNwdI4bNs8dGckYLbtwXW9JYn4Pnh/A3mS+5s0cqdYn2jP6v9dainJbxRV
xn65Ez3zRAGX0w87SI5g2GbuK8Kyigv7aicY0zEkDmB0nUtCLv7AMh0d6kPyQf7ke5GJ8gkB1ovj
BDzBquy1PIZH/SS6ggM/qp4AdENk9d7NFGSRZSi+WDLe+f4xqqU0BSpT/EsY6LnPdPJ5ol2fQxS4
diFsSWTQWWtMdoj50Fj/UlOtXhtGRJBFm8FKjdKXj8yREqomm2rdBfDi+w3+JiTPpkU5YQFjy3y5
MafTsS25UbkrM61DTu8yR4FycOZbIK77L866+ApYSU8GdCWsQQMZ2sVEchtknOKU5st6DwB3/sOq
3RmLjtv9qHYDyWzMwTBgwrhkVnmD8FV6KlxRhySzkE8qmvp5WMacvXad+orrp4GfVpWcoZWIu34e
M5nziZSVow2cu3Q7rIRn8phRMIkHby9U9BnGh1LxzcverXSpfr9/2UxjV0lKL2xa9Jk0eCMZFcKd
XIIdouuKovN5JhxtHQwUZUi+FPvQxBrfVd/IrF3eLcNK1uMz2+w4heR8g8Td2W2IB6ePae081D5Q
fVfrHoEyikWMsqojJA2WXbXTF4CwxiuSEbnR9NjTr6CbJaXZGXWW2R4WWQkLpedLcpHHYGKMV5kx
Dd38wVaFGjf1SFlxdK4Vw1fkK6yd6SS/Nn+9bSr8GutxfAgQ606DcRUi1KSU9H6utySFL+qgJ1OG
pegI8bO0RyBgAFZCTiU9OEgRif9OWAD9Uu3MIbVvGAoagqnvrcdsH7sSCJahkEj1+sMke90sTrYt
w2zmqt5/q/KMsmyDE2eKFDnWemprPV0m9TjuiLbfXB4IfHgUWUtecUTWwJPPeW6g0zN4kOGF7pz4
0j6kp2D7XHEf9BEmgPU+iFsR0rUiGuQmRrBPKIBGaNie9s7UNAqfLRr/M50Pw6AhxFe7kCCfBc3g
xM8je54FNkVUw0OUspLWGudQpfmcJfgt3bSwI0N/p9q2lA5QRLy2iiU8V0+wYb7uNseQ8JEUW74z
lTm1exkoNxE8HoIGViGmGdkZXRELRIADE/0d5YLOfJh2fBiEIxbUNYYnIC0FiVjOQgScpIM6Njft
2De72JrARFyUMOEjqjpv1CyihOEaL78xTE8zmsJ2e1XG1jWHngtpFV9cHdJm9/4ZFWjCF9cqBrme
9bBZ/k0KNwTJYXh0A5tqscx5Rb29RFzlgcQi0jpN3m4nQvwN4kpiKyeu4qPFA7GAMLr7PU9WzGyj
nwUojEM9d7n9C3i0FteWltly9iXjTG4K5GDbBGR8adFqXmCfiPfFag92NQZ6zvizUiIlZfnORIrL
7jUnnXo901GuNirYxXtRGxEBj8bWg4v3gdOqz7wQ+wiZ3AAEhfEEdtigjW282iBnL8oY+Muu4ArE
aESg9LyR+obuIRQKLPHTPWaIK/JC90b/UauxprJoNc5x0MDI45eTxiZ6JQhVA5AQdTG2tFsk3NM6
cqbkioaUKLtWdD30+sj6q9AkTU3RSPoQ0rfwMmTbnmoFGX306uQlAhq7VBvWhNYzSQApcQgSEk1H
0/HCqqemm8QDMjPX3hlCNaJtCs+SYC3Tpu2SuM449YhRhIT1WP2BjuIncpRkwVH0YZwLxIglRqbj
gMfq0Wb877K/qdObsyBY6jiCVwEZd5DTY0VtB0iXJGXdhfhr/ZQoKlOuMdwX0nmHJngIoj/w1zVZ
Y/2KMYbSVfLQIMqeWrhukyyNcZbQEhK5b07cSpPfuVotNatG9UpfjS3ToxUyGmQdf9N5BpNK1Bnf
G52tt/96xfOkn5OqCiSpM/EDSjmPeRwmIEKwIBfa3Mn/JZbk/mihzNSUj323MfRVB8ErvZ3IJvhN
FzRak/74YtTPLnsAlEZheLokadq6Ht9IqfyRdWUI6RYmQat8hU+9emmHN5OMb4zD0Ez42fx/zy2V
4L/Y2wem7zszmYMbqOf4VbyT2zxgX8CaqXtI7PAsPtg8fFNjeV+PDj5KzMtQ3nJX+Wlgq6XF28dZ
/WzaNz7yRjQEN2VlCfZARiBpRp6KDFGRSLN660ECNUT9OnsaeXLbEm9AuQhjGM4Xv8+up3Pf7JM7
pMT+bunAOxCuO1N9BJaoPzBrX+10++kB7nDVyZO3RNGupI8uCgsq1+TUEUNWRLNNhJMq5y5TiCfX
e1MZDweuzGWYdpAo+DZHoDnCyzXN5bUhTdt0eAsKeG8GFNtLNKQmLjmUN4SSaEUOOpiUT2b+6oKU
HdU3ggaJNxjItzGFyQqqUIjWWkqCmoLPJ2HZMyg1EuQASg2LZdLKiWTXyPppOlRQtv3zMot5T2u0
b5Ak/iIPXnNbDOBFC/L2mmAtSfIHdGeRP6nQaF87JCE9ztk0rXoQr0Wx/DZ824fMGyWvSYWukqAf
DAXtAxfjmLVx3spWZ242qJyzP5PQ+LZXkT+utCCy8LqWlCD96OKtWxUzP7n3c/M6unX2t9pi0qCG
7KDrS1yLs0UQjQL8p4sMArAicPmtC2FX4uLlIcXDxelsFU0IX618QB/525yyF3Q2YcAm1vokSX9O
zuiBZG5yx/Y/T/WxKxUCHhMRH3eChUcsOS8uYAOfYH1AqpmzsL+FZgcFb6MWc42fsDg3skZWVcph
omOb7CjVzJfFOeWlbImDq//UL9+1+WJj+X9Uv45FRj5gWpQLY8CllmKyH5VO6QEu+KBCO0/VOQQH
qljEfyqhNJ1Je7vSrLfbFDORGwWFHlDaXpdj1jji6UhfkFzCc4CckG0uzNkJ2yeZA9oBhMT+7kjX
rHFWatnXCfSPAQmrDdSOEMZzaT/TTsU8EVuRr5TxTDVeEJKZUwT+nOCiLkTt/Uen+8+88vkK8qwU
5iFGl6EVeFPsJuu9OAok8FkhPOVgG/ogkA0zKnhERZDS7YCy1EwfTrJBDs8C/dsahFU7hlFEYmJQ
jJB5XC8EACTrlP5vob1eOTgIGkXliQpJlIOf7Cs8jVbRfEAPh3Vy1yOhXMn4pe/JDCnAziwlurRB
2FCnXPBrs4YPLrcMyJuozAnvrSz5JYwlg3Tl+cgApGpba7Da6dnOMRXQpzFXOd177QjOeOTYBtJn
kLk4SJZVHgxrRfqM+yPRLEaik1c9xFg2blACXC+IItSERQ2/hD7MoBNXomIAdQSYJ3XCOq6ki55v
XGcdcvlM9HJSu644Re95BHsLmTc/RJt1w5B4qbeMPzYBQH2i5Cafj6STucotXiJTdm+lzyf3nViW
16+jVl6OcE+p8ln6l847VdTnC/TBOd4S1BnUeXhW8UYMVk6X22a1zR+DEtmfFCzaF2kC392TZ92M
YDu8Tf5TEhk0JTKELoon7HWHXcWZw3GeBF3qUuMxUju7Anc4fFlc9YEf7yu3dLshcO7TJHZCwWhN
pi3qyZD91Oh+1DF6YdiVrqiJDETeHfZerf7+GkILhNmO0tRboov/hfxHHKwBcJbJCvrdu6MphhHn
T9mEXb4HrJhJLIgBhz1h9CUdgZe5YZEbiym0yWjD4LoioqoPJ9JGd4ESXnLsQ6vM/fUm4jYEqhlh
jtvgABZ2ARSN5qhxLe5aMvNt37ZB+6s9rufwSuDaSKDwFyeSlMTJUcTmjiGRt2w4AWvTJDw9KVNU
8OXeRruLaXlPe39/wbtV2KMC4P8VAsByM0Q0sTQwI5u5bjO8N1u+B0iuVXIir4Q8+5TvawVrx5ZR
SquzxW/64SHQSVwsRL3R0s0UxdUlUkPAxs9+1EJWvrkL1tF2gYwRKrWmqo5w9iqAE2D/oxyw6AMm
AQSqcsBQvWUKEMraLRT8YfRThRwUBLL8XZD8ZgPD1WzQol+WTQX/E+YrtV66AMQJP7dEo6zxx6t6
SgHPH82/L03SFxO3j8N8FqbRNjz1mt4C1yww3J89Uo5buv4TcLLsi6duIeSq98f4b8BO55wgs7QZ
VdX0tMyWb8r6QmywTRAsFB8Paj0Sy6MJRuWzfYR00vaBM5yZKPiCKL927yVCYjlZPk5vntkuuvp+
xfI30q2scUteOr7Gg91IRusO0K7TTTH5cj47ksLATNoHsiXtlyMkq6HBJ+IHmV6M4YcqvlP5mmBa
WIZCFZsDU5Qa/Pd7J6Zz5dSuCTjznWTukYSGNGYPpZ2woPeOWpDIj8rscG2UVsU1O2pQ3VaA4ojq
a8O1hGaMe/CW25BLq9msIxTijAODNIxBH2ahk9iDpGpAStfUcT1jla6WLcn3fyeQO2708goW1ve2
mjGA9Sr5cgePaZhhBbf1uPVk/F3mww5fhOVKAHHXoriiXcuRu1xYG6fnFuAujTPFjnaNCMOP/shD
V7kybNNcqAjsn8Zak0oNXHlTx8l49crzrqZ8RXKix5njrTIfWr3HWdIvvl2qfk/Y+2XLNjDY0RnO
HIQ80gfwKd1TEqt0s9YVIkFVe7hATjK1BoAc2GddI2iEYhWZhFI7SsTcy7lS1g+TMABmgxRRrmCm
ZlfC/gw60nyg+d1pGt9VKtQMvuE2VpZmUfQriDqQBSyaYy79NwYpZ8VuK63BL3vmCfcJrYjsGAng
5WCbh651B+jQ2gh7zBp9j+9Ca1Q2mdwrCMT1o+LQ9K5jBRteg2anSWlLROUSLluDimq6Zgq8GJgz
TAm11uW+jVJl29a8RP5m2Iyv6RI9O/Itfv4gX2C6Jt4ET5pN7UgL0vCGE0VzAKHpX6RdaETuIjFZ
r2YYynsoLtahCHplL5omLeZG67Gdmzb5VHbWL4LRhNGehKQxw8aplQJutZLr4w2IUUsoTURioZUY
8Jt/VEw/fycLGpm9M218fBnDICPixUdPjCO2JNdjEezMTWkgfE0Mc/IF408zZ3Gv+CvU1dH1tG8a
cLOHRNxZ6zIpfiz6djm9THiHGlnZ4zeqd4IZ16v2gJmrs5Jz1S9JHsgJXNHkMcw8GLIksX1xY+Nk
R2a3NtkuWh89AsSIGIhU7NDRItpIoHTZKXrdsg0++Yx5a2F40k7RzypE3JpnQsCwY7i6M9bkbhZX
Lb72U9oUFFSZfjAmtQ5lGrmrFi37sN9FA2kC8bz7Ye9JBCnxALSiLGFZfP8Z7BTa7Iepa4PjlGHb
O7ILGemskC/XrwvvCzxq4XZmtUEn8CpIQC7zk2JXdevSpz57+paQTXl1hKrvQnESBv0/h9GpslYf
oApZApWE0MKaYKgbLCC69uf/OrldaBv6RQYoxmMFYfEp834p/GxDBZZ8zdfvQQPr//d4FdnwoW8+
fg27QVKWYOMnZtjmga8rK9jGl8NqV7m5t2ol3X1x4v0lsbRo239Fp/iVv+LQrBWPJwBoyEvNWdjH
2C1MgyKrbcRn9FVN3HJrgbwK/P345IY1sMMdDddubQp4Kx+jH1bI58rA4cHojCiq92AvI30JHlUv
vQe1I2Wse5+Qbv/6sELr/AxQ29Z2/rnjP59DTheNhZhmO1Zqv4Noar7UtNchtaawCoOUUpb8AXAq
G8WHqBKuR76OKTUz82oCEIzUcgP6chK3bSrW1LISttoOHfqkGGvxgmjuLlHktAZ2bEe2Q4E90JGg
qJgPjhabtz+gEObUe3iVVJ7a2OH3rxKmuVUMcH3vkU2dj6YRFKcJc3EC8BtCBHMxMqFrIP66sRpP
HPhYatX0sQJhBzU1joZToXKY46OFyPSBib4na4CxOZLOzLGLKbKjrKtEdJCePjKILToevRlY81sd
L2A/r3/sM+p44eSNsPC3qrNd3cOoIMTvJ4+jS1x+16CIB6vCwyMpljUkh3Gy1kuUeS60sv27zrPw
j0YPujq3XD1VYjYbfVHghhqQRNRVv3+e10BNuIQ9MnccXRvMHtixrDEvjsIYWDnhgmq2qfXpVi+E
o2AMM5gSdj7L0WBvld/vNw6Ilj93+a8D6IZVPiLZvxtdHMRq3s7jtzVKVIqS/XtAG08xmrSamOUQ
/FMopfkJ6r8dyObnW/CGPvrsUUwQ9abjPzxNs2M4elGrEnYZZdbaewdrkTPs5VpYK5STNiWLCda1
IHACvKclyZ/uA8v6jdnoqXI4P5b9KokZDGeZHN6CHWby11jW54WcFAppfRjLrnGoQLYnh4BkSbFX
K1b/eYtCh4VUr0hAW+wyC4B17S9BxAiOnD5x+80fH3LimF+Re7j7sbRsrWOdY2fEZcjB9alU6Gon
y+grygggx5NkyD02CBhMtaGZwpWeQNHnD0jUR3srYiGsZ1Y8WYNgSB8JGl5toeQB39R+N6q8fW99
hkdeOnpGXvxMwiH401V2BJGlNTTxS3S0uPBhl18gjmz7AakKpHsWsnqM6AARWpW4qRbpZ5En+WaH
QwBHbwyjlVorj1pXc074Vg2HEaa9EmlVYYv9oAj3Ms8I6jliBeACFSJ6XUeR94EimXxTec98MJQy
6bKUtQoP2Ym9Hve7WvENtMjkj4zZqKZ5c0yB9zRSv8EAl1Z4/Ivm5eNhMU1z+vvcOeKliq/mSZEE
C+LJ+HU0OkC7FXJ82n7btytac0fGV8CqZDb+2zDYXdULbu7nFj3a0qPcd1oP4zMJj3LyRV53WFCD
Ya2eCiNJ4GEfbd7OYLQ9/Twae8kswLDiTzgfVCSCcbR9CsKC7hjUTEBnpp9+cwjkm/b6Q/ypRy/s
K0DLYn3s81b6pT1CeQFAAiGKbCvTbfHkFmtR14rztDlXBMkYmGlpH+S3ygYDTmCE9QovGitQh/Ee
uiktG9eMqv9sX0/CzxpI4XxkqzVIfDks2yzRmgPRIL/5Je+r1sJJrQ3Dslua+imh7W3AgXUjGm02
XgzbWsI4CkJbvQv7gKVW2pBYFYxbnixlFTBiYKzCSKD0W1Mau7cqffx7Nov3cYdp8vMwxQPx1GYg
A/RAyvbfAGjrnS92bTTstQkbOvjYkZucLSSDNSOX8hc0xbNl+dMXu69q4QMsoWmJYgG4Wf/Y8Bu7
fUbPW8ifGU7jaMuvxkX2ZyIhM8DgVd1KlTun0z9ihEDl8pXQ/C2aiLxGHRzM8yCf4tJ9V6KuwGTU
I2Ty5v7vYMrkaJh4DzjklrNhZ9g1WsvNEZ9ezE+gshv1jjSugq2Kwwt+xm/803ow5uk2YtXJGOte
c5jq5HDwKWNSx4vh8CKK/BAtkPLNHyR9oD7x88fexoXJ5ZE3t2PTl1uj5lqEvkV2c2U8WSztWVHR
1jqdgUavJWKSl1tYIbGNiQdj4VhCNgf8FP9aeZm3zXzhBne3yRYq82zhJFZGn70AmbzWSfGY/kpa
dIs0S/75tOai7ejn+Kr1ANPQCD80T6IWX/bglkhR/uKXtWEqFf8jkVLfU4ZfhbtpVN/hBMXgQiyr
E65Q9q20z58t/m+g6FF3rKk/K3SxxeJ7PcmQEW/ZMNa0mZN80qp1VupWXTT7OmqZyiX8Ppup4fhY
cXk6W4FF072qdbq4g0wvSyRSV1w/Y+M0igeKhhi/PqnbjEE1w43zeWh9GVS5yV3lbN8gg/hK6DTN
LzQHeDVIoC1jsNuRo/QXZA2P+BVM4jlG3gj149L96dY242EzPQH3CVmjzTBAmrTfKj97ZY5EIY/b
WwYk52ajB7Pd2H+ZeERIpscDd/ora4MHSbY9fs5MiXYQn6nu3M43vPDE/dc3zy7W/WUup5xGrs7g
TMq8uyDgIqz5WyPeaOs5elyuvVJBREO15BgbJKA36/m1O73v/zKEsgiTE4DnHouOpKyAnJaFSPER
HF2NsXqUEjQGkQoni0z6fNhWi5XoJ0Kd+dKp1Dz5dExcLWMswxTRdjtk8Snv5x7cVF1AkaBRMbjn
YXj1WWutOXqah7iIbOjPQbVuCSdbtyXHTRVh0KaWcEMbZm8X5EQMGYSnwZMtOihgaeMyFNUWD5DK
PGi2vGYQxxSDBhS1u/z43Mak3KmuyBR1IbU22LIK33nG0F0ipYsMi/GuPMWfcR4aZfmWAeocdjml
yCjQqjl9PwT+FtkNnZl+j5y0Zsk1ZJmvomiqtTk+g8R0BF685Y6x8stY80v7QdTEbd1pmCLXMUzv
D9NKkC3hdhA0j9mVK/fE41RfKb/NHlxSK8uryRTfJMiFlLco6O10hEvphHhGwR1GWhFMlpAWgkSQ
TuzLJl/gDCtSKhHHeYjKTg2H0V13nvH4HKGNKOZXFC8m0YZpCdl1uq89OQIT5kK2Y4/uzuFowNRs
OtccPRRQ+SUe5QdXx86htTsn+iuWe+KFlNkEbLJ+EoKxKYeq6HoB/Y3HOdavuHzDFc4q78zmc+5u
elPkyqpkiFmHjA+bHjGjqhlZOFWMQ3XHzRxqJtuqZIMVxKBtSNxi2ZCfYNaXGUnI9SMYoggvjPrT
DCQqHX9x/RJVSTd8ZNfKqenAHyLV3XKoxLiCm2kIp51m6d+dKgmkX1RQcDoOsKmZmEEI/zO2lsds
Q98A0lC18PjT49PdOm68EAuAecGzZqgEtQ749AOmfI23ghBMTDgT7K9ghOt7BMwHogwUnJaK2kWH
HNgwMaMWpnEfPe9bjiFgkkosutzXqiAGhT1FKYftdiBIT0rdMVPV806mLMSlEwqxxax8Fc6Rtam3
FEl6lJOw9IGbQ0yEv0RZxXOH10MfyRt61JTDpHNMJDmZA5YD+SVSIrdvKgQ3F16k6Nv7ugk5ID3m
U1oEgWUb5zRjh+XUuG+wqA7vY+GOYkQW8ION+S+AxRuDBW75S4wovq6VmHdb6JykEeVW7wU0CdbD
dZCd9M+xojWDKTMXKuXY2Ont6gKxLWBaXA3L2gPeb1CxaCcmWJNj3i30mJugAQG9lJi1cP2AaKe9
dUnn7Mudc3nyep6bKPwkABrjrT0J70x1jVuZY8Taac4tcBUtbm2kYzFof/TP36nFk4CnbZ62iRHe
RLhDdaywX305VhPCMjho5RNlQkJu+LFxPA8jaqp8gp9tqo32cH1B+ZVyiB3hTf+X0dKMmVCz60al
tefYbeFRDzYsq6CXQkvVS0/YNAM/fZHO4+vHK4BfoTsD3alWHF2PXKdEOoKtMjJA/U8CouvJxTu7
IxkEJNMCVOL7M3Z34QdLy8EDJhCDEAhjCU6zy5zR3H7nUYvtYmBCng4nhN+oZKEBKZn5iEqmH5bu
BTen58j6W99+ooqRKFBsCz/LNeapHSDJqtXdu3Yi3zGKvPMKeR9kLDP2N7VByAapba7kSf5gUXma
jFc1A9gpYW3Vf5McroATVHXgepxFitNjYC8slhlcyXl/l2o2PpYp/QNhwD2PfQHgoMzwYJNhu30c
Flenl2mydfmYaFkm4UuAtWUjiLy6hCGKPCtRwANUxXHyvVDEsLbtj8qj6oDuvhtwNJkwwQGBPsXN
hIDxwiavLuU9aLjSq9vFK6xlxEw1CMZFGdk51cDc93QapM+8bcC+yNtEA4M8Qn2+XTwKoMan15m1
dyB8/OHzcV1oVPOEJtu+tednh+mE/Lg9O3v4xup9B/Ss+3wsGSEGOtKWy+590hGvHFi8JbeD3MX/
C5YI1sKhgBB5OfmRgv7CdM/fcpP8IJY81H1Lqsjsu+ePKKUoAUqaPOy32e6R9p4VIsZdFl8/YVy+
Q1af9m+kWU13CB+/BwEBIxBVGu4l2n1oNTsPF0NBEchoBCh55Ku8es8ENL3sgD/Ec7ZM70TjBE54
T09rG6X7TtMMAsvQY0dwIT+fVkTv8i5QxJMLD3sWSwiJkVFtPCp5brSy2OWFROEHVSN9rkUkTQIE
5TE1dOWm0nTgV77sjw3QEJBDfouv6HJ7uAO9A6iguM44ogzP9AmBd6v86e+Z2DnXOXbvoTcNnGk5
2qWDXytL0KiNl/eCSxgfD+fw7SxHZgRjBaInRTcXJ6umDoDF24htJk3pEmxmeBVHIMAFAtbS9/nO
PpqSOjnkVpL29dIQLbuWt/lJ6Zg6neRo/fnG5I5LtJOm8l7DV3zXtn3Ok6/HqDVWmbMELf9RirRW
/bxBt3RcTroIxhta3dQ4Iya9l+1RyqVgUniCID9cVsc3aaJpeTxa8o1E7fxYVgohZsAuW3dwHSdm
6flvKIkqQwzFTdAmTDbNDVMzXSjaFHMn0iO2A6zoiUvFlFvnaoDNvyDY9zjk9hx7pNPyJc45q3sn
myzck0LGaABs9tsovPQd8AJu2TgTn9oQx5CGnsZ/d3kgHtXV3ISHFGPMEpN822PUhWD3X857ufFp
a93Sa8BioT9JJjZBme4qvYs57/oV+RGzpY8N98VREYc8wqs9fnuf+8JKJUMQ6SB+XkmYHD+ru/WF
W8LtK2FnaQTjDUgx2lm0F+QcJJkWmciwkpeQ4CtDhUuyiaMBMagFIwdH67VhPeskW7AOubS2Qpyr
KOj6ume+CqSzydkIEuYpVbnkeJeCapzBFpeKM2zYt1izRvpIYI/QDQUfcAVTtkUtW1I3GsR3RrXd
Y1/pgn0g6mOogGOUiXcSjeR8FsyehmbeUz0qKHzme9+zBEGgJoUeigSsSBE8ohfI+plf1Empvz5l
NPsjAiic1y8VqQffiTd3ybGDc3xL566U6PbXxl2K7yqYz7nOoMWmcUdncbSJqQucmgsZrp/O5y/K
hgexAA8Uece7WYxXt83E48elmSOYhrDxQbaIsKi3zEIS2GBVTSvgTlt/PTQOcSQri2F1Col/HEDM
NhRZP/p1RWQNQpADvjtbAdm1b25Vj3VfwftXblyTGl2rEga48DYSCtYplkP/TxAysNiYCMqF4gMF
1RQ1IyBahkAH+aMQtlnxrcMJqdlovNevq63os4Lkb3HLdfc7Y0C2SGwHUL0iuJmNQDgHyd9M9nPQ
j83owkjphZ/+3rDiQcZp3Vrk1gnjzIK5UnO2/ziP0LG2Ym+5PEp4Wk/9Rbn+ZG60g1drJEI0ACg7
WWhxCUE9AOIrBDBhvIKrhtS78nOQ27a42YV76Tkfeno0A5EDANAjS3gPRqTwIAL9bNSIoBfIgIXY
qZ1qz6rq6irS30MLEQub6k/dxJsvSpCm1GwDK1hLfPm3kDUlHyRFY0SLQQyih7260Km69s9rA2c3
jt4dWLTaTdCwsH3Eyz8eHwukIM55qe3OJ8G/7qPkx/7BtaSP9a+5ZUspayk3lnMwRYHAWomxT+1x
p+8YtrxTyZZ/z8aMM/xmcwIsHsRe+znfKdTGYaYlIftfESfIg/lsKw0xgQHloZh7ydFQl14ypeen
SucsajpJ45Tcfx83GlHm3seDIJwrGl7ko6c0uiA+DvJEBaaPTI0s6B3eyPZcM22ZFTeqvBUGFa0U
tpv4tdiBLGqpc+ldq/t478+s96bwJod9h/cVpexzgfdjqbJhF568y65TfDmlvwT1kLtKDgVU8Ixj
z7hRWd5Z/B4G2Kxr6zUNE63jp3wxiwou3ola7umoNfv6KF+1ijK/aAvqJINkHG+BCYXArQLq7gLX
gS1Yl5X7Y7I6HlHu1LCzvgWkrj+pst2P5RmbynjZAnfo+too/3ew7YAVwyUWCPT9L6o2e7aAdIxw
D/5SB/Dfan63hOUYJFnj6jCMxNThaYTBAK1L2eoyfaUCDXFji6vgHVIEywejVWgnqHCMSzEh1ftc
opZqX6ndMYji2N5ZcgdEOUuhxlofgRzybzn0cN9AVpsW3D/XyPDUb5vO3rHeNLhMPFKuCe6Lds85
caAa9463KDC9kRkoSbst5kF50OiXwvx3+tBOSJirlvFOVXH/29jHSXZTMhx1LWLYZzqck1FUXcfb
DlxayIwFswHAfCN4u6lG7CLdFax4PmWVC4DK4SSEqadG9gdBqk3D/yMDbtlD3xvLLxVvuOSakv0G
jGp0LtSkIq51u2YHKqM2vGoVxZrMhKui0DXA8Im4FDtfPpUWN6pJai+YB0p1cDjI0ag7vLqsaSdw
SXWbszMtSyDLkXM/i37pZMQrTB/npPlpvV1UFiXSESyUT0aK2O0GA+7dPQivEqxm2YLx8PpJ6nM5
wSn4P/4ZzCY+TefPOrsEE28xunuQ0tlmUawmT9Ov/4HahnmfYoWv+TPd8AMF+agvVDFpwR1cqmn6
eSuTpsGe8FtrZ55WJarZaQ/eaJABrjMuc7+J6GALe/KXwKQBBE2wrSFjwFFBMnG4GTJKL3utr0/U
aNkHNazi2EgHJDzUqkQq0P5spN825/iVzO8LHLc4YkhVILR0MoCkRF91TZVCQAPPqLSsLCa8kYiA
4aO9QyU8TSjUD0VhqytG2COe1vwGSb3I7GcrmuwGt7cY3frPC1an480/HfQ3TtYQ55CD/gJ91WLK
s9l8Er+mK1lXUrFRfuj0gJg2n9xkWyHspa5UWJLIFGj9+nJIzIuHnYtD+8BrMWhxiq5Pve5nfWYc
RU6+md9zH3NQVPr39E6OMPpAXzpSYIst0HQegNqDzI9hAFIs2zYwVvrWRTMreU1GdMZdmohMFD5G
g+zx125PnKM4/5OOL+O4BGUbsFPAh/j2m8RZjWnA1QdIzNCCnZCIaRjch/FzuDXyTBBHWSB8duVC
87LtJrSByxkaUQgIPlozUzRaOgp/PK9YdHcLMaaGBQ70YdyqpY/+j2UdsWuS43wExwjRjoicRhDK
Fn6nYeryWOmpos5kjiCknV31wTDBRuz8tNzNQiqloPTh4hfJIPstg0ZQtDs7pWuxVxVDhKj2b1f9
iSTSjh5Fy1dTJ33viMGM712xmmAQl+kngtBGUibhs07O9fDi2iNhCXhF+/t5PIsGThTP0wbTLk2z
IQyIPda1ISM50GOfPPf493yrKImWLl7NYZvyo6NaClCAg2JsUVIjDiL0n27qZDHBGm1U1PTwhHok
SRM8/7G4tmBwr1c2ilPB8hx8TSO/O4n1ANRls0r7gBg3vn59qe6fvjvDf0AfRWzlM7T5WkESHl9v
heKFyWa4R2zMm+Mnr8iHx9j05pilPVZjKy+7mb6jg/5orvzSFqs+OtwwgnBwWRuHQ/mNvC+C7nIy
ZJbdCSGLL9iuesCBmjQsW1B3yLTY+94Dh2fvu3SBKGccN4cw8Nq4qA1CtOLrsq2Ab7SvFgpmh4L8
Gl7+E3ELJhOaZPJNQk4w2O6EigYaM+dZW15Uc4NfDOBHbnGeRCfCP9/a1/E5lHuaaOxT7uG01Pql
erC+1M+ou0TYDyNAGOMVpm/ZkrTB6H0V3Lq8vj0PsVrvQPhHAJAgyqEdYPP7hgkK26mYt0iopUca
Z+E7t2oSCOtU8vrkLgKGUePZZYZREocmdRNvHZww6LkjNQsr9+T65GuXOUsuea91TFjD7BeXsaLK
5JvB7LT+mnL4v6LS/jpv2Fwk5IbsfAaGUlWj8JnaU1Yea/Gx8F3yxOMt2M7qhzdOJ2ve9xy3+RyD
g/H7kYvi2HvCenmfBMkPECtD56Osge23Ewt01ZqvxGxIxHVnv4LcFVX0iolLVQ3D4IXwrFjrhemU
KlDo5pP8ollaocIFgyGuXy20FLJeJ/lY1vxP+mJPrJSWTgc9ifytC2zaLDRYJlLqghVqYJLddz7n
t64aDIwhsME0GnWpqfj4vv7vawi75+NReraiuKlad0Iwhd/Ff8QYkEnP1bRXd5LwIlf6Y1cQkd1c
C1BnNAGuxi/lXKnTntfLmxu2aDm1GIaqBvrsmqn47cr2lB3gjAWQRZmIy2X7Mc0TKcpHw46VXoga
oeAda5PkCFgXwtjLmQGEds1YlczEGMQdMLVyjZwdkKLZmXqZio8zcZsTF+oAr3P2I1qLhbvJmloM
kimInDEGRAJrSwOw9/XECcLcFuyhOs5v5WvoZaYDYNCq+ZFFzZ0P8lSorEMU0Xarw6oum/KRbdKy
7mdXta9eDyuarLbUM8MCHLA5Qn43O/vhBSPXpq7bIzREHHXEBowIoutaKtde+pTkdC5DPbJDC8Bp
upR99ClWCdDF0dR6hhyVdB4yfyc9H9BYac3cZqTtrfCa+yn0rPp9ItI1GCihgv7Gecu5RkUfl/2e
BMqkQZGAcyJQfSf1mZjaNcCqTxJV9x87J3xfy/+bmezPjxEkruhqHUqeHCA1TpbKoIB1Ai5bccMS
gETDXQR3x8dBeKL0BIP6eReDfqjomIefEbd5JvufcwnTnvDv0tR570fYVUNoJHD64xp/BL+/j975
wmbYKv2YFhAfPMMcg1sX1JN7kqMtpDz+ko68LSKdxB7SAh8vcQP4GRn4ZnGYlH800jb5/bxPmtH6
ASnequ3TRwqQpSDUFPE7U4zW9uoA0ojlNCw6kHGQyrj8MQAFP1coIGjxHcqKPRLb7J9dgxoOaQvl
/4bBLpgg4QVCSMNY9TM2U+HXUq5Sa8bT9YaLCzsjeFfH7udctaADeha8OdhGNANYfadOgPs5vDBg
dqosWGbQhbMBJKrfbvIOjE4aXvwVxxCesX9WW4m2xruRU9jrxlqG8htsaG9blL4Y+wBQoKnFhGQZ
dwHGMXnMBid+8VKleyLiTKKXEW9gNV2jcvShGkPj/Fv+bh0nXzf68qpYYPyOBCn7TWa2tQCK7hNT
l5riWpBVT0tn6W97HskkHEjgDBxxDLMqTMbkwRLZ+uuE5lmKa6oQyuAIpU4PyErP+gAihWW6qNCJ
lzFm1X3kRyI6vXDuQ92NRtPOzEHWY636D3e7lNJgvX7JmbtcEufRsU9ZRijCwm/YOXV4kahb4Wzp
hHNMx2EN7pLpsMtStunMZzQzdF7FmSzkOdos7yBeG8aTi4o8sF0RMuC/4MQEQBM+pVITOxgYZo3V
LLkW2570A2/lHNd7JgNni+0BCvubmpG6QSLO8/WbQbhAltB8s42Gc6w9CM9aLXETPIULsjwTGXMO
oLafKM31a8AZc2mpYM88emLdFHeRM4S+Rbu7dsAfBV0pFuksTIf87sw6CgLyWbJdlniR7FHqfn+v
Mx64ycTNWLI8ZesKsb7gWvGBeEYXCVpmcejVKl7pFok5NvF04E1sKvTJPaNUSVms6MyQd0Q4gr+h
3adb8x956eUyeDPbT4Zfxz3PIneo/75CBXJuAY9Qgq7khDf3ARQ2quDnUnnPwuDwQ+sgYb3bJu/X
alji7YykxDA2tioR7vqj13NsQeYlTyU6BfOBMWFWwEdA66ysMDH5A005/3YqvNkiewl0iUrEhJ2a
/0lgLNJcq402BjXvQiKtOLsvkwzjoGu8xC/YXtAnaFDJR7pCscUySD+uoO1Z4n3hSa0xF5Hc+Lz1
yE3bznfEdxTJuw8EFVL7Y21CV8BCcynlEttXFjd37fvVJ7JyBrkgF6lvxh0LyBAE2pk6BGOc/cM6
nQ/IRG7TNYJIQWiv91KjEzQDkCjQwIXbF3a5cwaygbfyeuz+lL30mgWBXsj5qKnCF4abO3vy5xAX
CsqBm06Rnblsz9/a8LywtqFrBS3zCRlXgCptVBbwaQ4zCToGxiyTFCm0ezIG/GUfsoX2gvNaDz3U
ZFrsTH60KwJ4xPCsYU8MOCL7ecKRBBwG/lPfcnL1JP3/6PElU2lDC7wexHDo2n07zdkh+u5D99CS
QI2uq6dq8rrOkf8xX4TJM1DNG6vGKU+2eSiJnlCoCOdmmt7x6ipPaSox6jXoO538PDfBk8vgzSt9
kCK4XRPFGdBnw6DaZPBbwi8jc4/XFkLh1ZefM3TA7VilrU3P+9Q5aRRd4gShI41wUSy2U+jT794i
ojV7co6kZENIJL847KjZAGPQfiW0YQAzDJ7NnTIPDUcMKZWhsbLL9yFifKK870FYNM+Q3S4kgguz
fDWzuuep8Md0pD9Y996xfiogQj7bAlFqBasp6ztVCOqg522ntQwHSViE3tIimEXLzczq5/wu/phd
ubVNB72h7n8UazF3Mf1xKj+KrifQmc8vQ6SMcgQM007Wbz4wycL3paabCfsmbbnwJ95u/Hn+heeg
nWCiKYIs8QCqWKjNZCHPlBNDTh2kx9R2bPmfaFlWUMTTHbIpNCJH3Oho8v+Z+NOBoyaJYdpC+Cls
XFl2bu4+R6dT3WaiwXcbFME77pDQhK9J1u6cHSprBNkGnLMjQ1Cjxwgttw6aLzCcpCtHUt52xv0z
vHS90C2+pLW4+ITwu5ncHROa2qIgjRLCkiyi7E0l4BqsnFO4hqWI/kRmJBmzI9IicQicwvG/Qaq+
yy8C53Hm9YACihgCY6hpINnSKVFntnAozvKVqrw5iQS84hhvXbPOCuf4guQL6R6l/g5Rl7pMEGbP
ml75tdlZ9+cC/Ais6QlpjeU3loT6zbgohaUnFP9y9jz2RDN2AnUeWq2knVv+O48a+grJJwT5eULz
o5t7knPKBGMH4Tp9zP6kADraZpr93s+TtueHg2lS8Ce3zBNZtOfaXRp/rM13YSehiOiq6oPVMOO2
+9WHxdMC4LwK0TfLcmD3GEz67swRVJqBqDA6XKB+WOsJV9MJ7oMWJjqHwXMljCKxrLLL1B30Qu8A
tdUhy/mzbKTsl/kABrU9Fu8INKREn9Fv7FSbTqcKc9Dnux47NBXoTkYeFJV+3/+2hvL9+ZM82gVj
yM1xPlv12ENO/lI+Px7Mmdbp8L+ejyknZKIKLlDeD1/C05cHP/AQP1IdZioHromjiBZwsxXPWGbo
/HNTmfB6+jiWMJ5OmCN7JLSxpi3rFiIfTCqlxfcAoMf2gJkbliGE6owxWQBBuyle1fmaThzXLUx0
o9jJProbXkjCC8zSyyo7sb9bucCkOuARM+lt/jnF+E7Lxw9+3nnChQVriLxXBROQYovHnZlAiImJ
wQfk3yLbw6RYZJF7es4uAqMxrGJtb4jtvGSZFRadyx4jQ3A48P5DQNLrj8SCx5oV2wMD/5qbg4u2
+fa596Skf1GiIf4tQiMqBhHQcmZ4Xmm025QNnwG7EENJ0bDyw2tBOZEnp7ezRyixRKg/+KLKmtQv
qgqm9RRRbGjjGcbjU0eYnMOwNyXW2IEq3RoIwnd3VWrrxU2oW+dG3imngyDEwvFIFxjz7dagL6o2
duX53OJUn94XW5llwsFeBCLqqD8pSskTLzfI79FWmW+5qbjS1Nhdylx7nPWfpAB3Z7DLjF2R1F+M
EQ3h/01qb9QDm3miRKQ2Nt52uk3jGhC+VsHOLmy/At8JEzOz21V/qHCzYkK54hGwuYTzxsi7sXyl
6WO4svZ0PgzUh3ewWYxPT1VihN6LSTsHKB/Fr9Of0K4QJF2M0WAEJAsN/XOYJlz3Cs3jpPJ+LdHS
6YoAtxv8tE9u56mUNTBTGhV53v61LoPHVD6I25prlT4oEbqJfjHz/RriHNDyFId6WxaXi7SR2cRo
lAaw0Ec5V3MEAQSSOSUMkb4uKjQ43XpHzgYEeJwoNm0vpXw3b6JdCTL6X/2vnWh7/cGbonyQJNXj
BcJ0O2yghEs7ftKRFOZ8tgSclfubLa5bFTe6TVdXuHq3w8/hUWq27M8uoxo3gTCs9vGlhCj+CXa6
SDo6NY6Oh2GXLGhwHHaxXsE0eHAJ32Yy0s08lQzT7pg9WZbcEdzGsKB4m3CAtOMRc1Wj2H6vAla7
wR4lHpriOSMWHAGBhnUS4YN3b3DY9gOpdY2L+KSY/h+jI87Q4JgVShR6Xk73B8fcbNpRDa42rZDw
qzzcnziYQv9iRhsltlNFz+UFPmX/wm7cE1tQ8NjnAJvHHxzfZDxtygGnreBy5jr9tCDQlN56VaNm
4QgZGnKwcwQjdqahWk2bbZBljbl90wr9PgEV4pkbrdRDoGWu7YPVBrXxpDqC0/czb5I8Ie+1k9u1
dBCFQu83pcvjuewdHWgoshqJs+xc6GyoEOQQmuX/Jtr9dOZWRo7pvIOyPfpBuptWnPhhiHpLkiaC
5bou7NZ3AeYgNqnYnWpEiF8v77j5B72Tzg6hvcss+A1Aj/m34R/7rtvBqu+uSDnV02w5YBmEMhUg
p7rMZ0GEsfZefXCu4lvU8Ld4w5nUrAqFViLahAQ8LPNMXiXuvv/iqCyKDSmjufvmk1QvM/IjPuEL
GycX1YCdI+XeXFabi0LC3mIkuDTgGTflx7/nNVWiBWZ/ncKKglkd+Kch4/diqEYARKnbh6cG35NN
gkKN1mkGzZfasjgHdXrqZKM7jcz3N1PxxhAF1sr8lG9MehcVTi5hmvETupi9wyF30pfHk6d0O5N2
aHLAwIN2A9Fc8NFdB5vfJHYIW4Ce7THlstJKPksFR9BI5Z5mPUWmjvZHTDSg3lXsb4a641HO8T6E
YSYLnRESU9TZdwOnAgrZsjtjt+CfuOYeDlLfrx1Xt2NIEZpHYkzCCnJNnNnWucL2Ke/Hi/Z8B8pz
LXORh3/FNkZWQ2YQDA+0GzS9+zppfB3Zrx6ILZTnf8DtBHZNzdB71pucnrlDXVm+Kr3/RSpJQXTH
1sRrwDgfkjx0Of6mQfZVE+emNk+VNkIzFyw2UIW7+O9NpCuBUzYDGzEGLfTZIuxGbj5kvBmGZU9b
FZAQQqK7LXSel6Mw8VeJkqsOFNQ3xJ9pm1DsGtJSsJHDa5gWNa5hjkMmmNOJ763smCAtV5QS07Lq
DOtjSJpCsCpwcR5OFFwUE3q/2tyF4L5qXKUEMCJgl57wdu9VKRlYYrOkG+v05nz5lptIMLE3YqHo
1jyUljfFvxmWoBOn5jgijYLX4/v9xsWMNSyisJyj0WvGkTvKEEXtNzi8ehqQ3HAfPbhy0qeGSHHL
tzC0NVImH5RrNaQf5oq+JNZjv0ZWT6Bkkk8Uq4l/Hbzs8S5s71V2Nl4deQlnG35TBNqc/RG2EnTU
3qoaq5eVZK1+Ey+pXHhpZ/Dv6mS4+9WYhjd6LZ/N7OCzlq1Yiil9HllkThN51pwSfPSzGDWXGN27
YGaCTkwtspdgO2XubIXjkXM2axBTMV97jj+GTRHH4riagv8fDesxzMI0Uz4dl7zzC3fqIwx0gym2
ze8cOLOBFz2qq7/CKleowrQ1XPTdEdt9wDf6tsN6pymuwGDekP6+VCel8B4oKaa+TPlktEjvXQhS
aA7TV7Ga/ObyLIxFwYtTyZ75mXGWZmhQoSFXsJfpMQlfZkAmJLVtorc3oriT7r7weLGz95pmRsPG
5nw43iUOCVlEhF8gbCj5V0U+Nu9BeL4oQZgDcbTE2TtcE6FQ64OuH/LS4NFZoqXAIuIXNVVLlKQr
DnV+v4x5tbcMtwEgGry1acofRj1083Hs35XH0yjTDkC9jJXdf6n4VpiTlfFDV46DwwdUxyyYWs1S
SQkiWIAVG90r8p+iioSe/dpXXsp15ds735lQ1FdyCpjeSSIDiTi7xh0LXM7lqfn8uB4aeIt516d+
MMsLKduIFDd1C8qcC7VkC8cpz3lazoJ4bfZGQ3oqwW6OdWbAIegpWtozz8hAjEtTeVCc7T848/r7
QW91Q1eX64qNPaot8R9UC32FQrUSzrJVFM/Ss9capNZ0soATYqxszy8L6TYy0oX9qJfJDYvtHf20
wQq+c0Tt8f1RW4FWLx+Zk/PWHI7v7DRwwwsu7k1LPy3t2oga/UsLWNV3gKb7jOhk3jzk1UUF1TPH
zrG1nI+c/Xw/nYHvKf43xHXgpbZ3GGvDunLJ8G/RLXuPAplct2iZgk8/4DmuWYCFN5OHrTyt2CIg
JZwVjr5Z71+G4PJNjIoOdh+Z15xJT/fbO44fJKXRzcsRFeerWIJqaLUhhTfLkbqDbu8Q8ukL4np3
nlY8PdSA1zKjQc9uZvdD7eWn46nhylC3jKjPZu2deWjZA37g0ToGmSFYsI2VspUU3Tgs6KEJtfhv
qf0TWLWwGTjA6NI1AxKGA4WfW9sISPnmnGjwKGlWNk3Mg7I+SGsXZxSUxjbCwzVYfoBeRqPCFNiC
Eq/iTHp9JR+a6ax6TeKJnPidwpE+iHBR6it0cHw5oBDb9HuyWsxSxCn2iR9XNvkz++MFMsRhAsQn
lcH8Tcv9lAH2n1+jqlKIvp2DCTamv31IYUj9eRiVcyN1I6q7rvdf9LrF4Y3UBQtu3h4mCRQ0IH5I
T4Y5TCjHA83vMkTA7zPN1wRNxSBaLbisuFnUTkO+ngIrhJ9/aShm5faFcpOxqpK/lY3xTKhP73g2
JHXk+GNINy6M0/1jUJajkESC/lRLPxa8oFjWst3SzkdB/CBG0r3e9HxFo5GDCWXrky8gMsR3iDCX
e7NicQNQOVtBJDTH+FQ3y77fCD7AJ5tqMZ7MA8G5RL+Sjk6ldPUCuDykePUozaNOMcpcmX9IDJGl
ZlUnzLoh0o8EeHdtc6zNkuRXgBY2z3winS5hbDYI9Vq1QXtHzZZxMEh4rIBFh4YIqeawwzX5lSmA
6iHDza32JPH3DOAArZ/QPLWrXgfMVz22jdAqr5N3jqGEGqfvZQJDr2rzrMZi2raeZnuTyOJNA7zR
gxMxm63s09c0wZLZC7P29HZuATOw/W97XW6iaQ6A6IkHIlPV2iygtqu7D2Q+Zs8L0w1GVq+ADAhv
DWv7JWzELsrZ4xexXC52a5UoKtcSubPt+fPLETqRQEdA+zbiu67ASBuCE5Hs2DCKPfp8Q4iq3uA9
IngSSg4Hbworjq4H1eea/zl8OyQkmXVOsx499dUb2QTH08B24l5dgzkV/V7ILd3Vyzq9YvqPWkTX
9fzNZvQ93jZHGcbtZPw+/ruvV9gkw6sDqYIZQB/DCxYIy0CQB1bPQHMI8GQg9i3WdzbtD9yp081Z
gHy40NLSUTQ5KLaf700VAyHzXaVOKwsSOPhlxpQPeSTWYgI3lrRsIvly2i5hPVZokScOnKXv4XB3
aYO5BAHSY9QzWMaAJO3wORycj85TX9ZxqjkEkJnCPJhANKKQfQmVXwU61dyDddE1+odob33Sm/k9
Ka+DszhmOKuX+xOoYumroiFD1bWtW3lcJ/F3TQUt3sgEKt5yTUsJhr6hW+wY9CtjUDFXsGLQy9ni
dJgp3itN0L+Fj7N8buzqCWG5Z7tN1ELWc9OXRtVxVB2NrpKIFpgUOjvKjySVcLkImJjtnvMbdxA0
O97jzWzii5G2+zx2mcaAZ1pFGbfdKGfCmPEtUH68dx1sqX6WkfeVKQ4PtLrqa4U5oAIsqBni/Alm
2YEg56r0rBhpe71u2G9isK5U1XvjoT9lSYdjcVP2AH4JCMpxgfSKjYSn+u1lBM34PLA7ufs39458
wp6d+pOns7unjU6bAFO5aca7X/gG/75IGqCUWOeI0tzoHCy+Fy+k0aqNzc8OOIBcFckHgXsmCT7W
pR02F4Ki7hT8AxcQi37UmVYUY2ICbS+sBvq9a2DZVJGMXJgpZvaof8/ERlhOQPqQAGGcYieEKG+A
kvgS2WJDN/FtMVW1qEekcSHeyVyY+RdmcnTyHTeYGJfeV0QcG3ip1sdDQYgr6gbv/g1UqahHXixT
ceJ0Xdusm++2dytgzkDxbgzFkNYjdcP+qrrz0xXhnjcur6B/W+Y2gcXlvMf+Ckz9Il9SiFkgJYq6
n9qocdvCgxvFYQR+3zs8qJrSxsBl+8juK0CZ/mHxDDQ1tl2XhOpn9u76PSnF4wIwPytGj14PcOV1
bFu4b7Jt71nmMTcJOLoo6yL0FMTyeJBM+Rp8+uVK7pKFXAEJ5vwN6zNdnz1AnC21kf40IRC9gp/k
XLTi8Cp7sWZSGgyoABdfSj5wacw20dr0iSxyqL+XYKuDewlTq/sYNvqeVAOyPrMoDQZ+SHmeSs/v
uAPERi626oSn9wswc+jx7ovNU/bCZBJT5XIux4t0D+GrhdZjHPe+dC04JLKtA3eXfzvfN/T/Ml4x
Lq7OdtuZy+hZZAmIW2FM5i0Q2rhI8k9dBX2x1vqE7h6B8z8hLhAuaqd/rnHF9YczmJBvCgoikNL+
ziXDGyUMcoEgB0b3Fc+ZilLsMzJ5zxiIeUaoRSrS2BByLsxed3hX6upcGBka1fP8M742QRRfySr6
RgpkmRIRjdhQNuNjkyfghc2TzlhGOYQBkybMS5gEPV3XqtqgTBWjiu2XgexJ6UpMrsG8W1oOxVfl
96KV0isW9wxs3sxMVSCVHJYTcIdRqfDqxYFbpD5HyjcLAgRI+6ujNIHJIxc7nRRHHlyILETz9nyC
JMhruZxDNzfUp/0pZnfHIARaE/JHn47GUa0l1GpBflx+5ErX4fnCRKuYyjiuQdEpY2QxUBEuM21a
P+brwVkbvgTOkYosKridEulx/jtWlLeyL31iun0moSRzZiAyKl/7Pstm1i+VMoqK9L5zvx5gIgES
cy+yJUps6tZLsX0M7f+O+9Dm2MdRyGcHuAFHaW+yYn1ZTScnS9L4uBHFLhbColU2OBCy52zHW57R
TbYx5CD0FjLrYqcGNA/Mzn1Uu7qAwkMcxXmlwn0GeU20fVZLYdTQHfcnb4DKBQKZVysioOeWx6RU
25CZuw5CmJQPlsDN91Rq2EFGgceonbqqzZgU2Oln47O3zn2P2lBhpZOUr9JJmIogENXvncE/j2gR
sKpLMq0bhoFXNJnLIje4LINffRHN0y6u8a5lWgUrjyv9CD1ovdd2JE7sv5jI3sTYqr+K0wJFzlEb
vvlaZDFV6H4GcDLW/DnC89UeMelHvIQdo0iV7cR3zRH7cjTI91Y4HvzMYFw0eT9QM9xvARZOz+U+
zGDEqPaHS82arwi6YCL1mlCxEbsON8OVqH1Up9BN2T/5/iTs20eSy0kXydABXLnYWwLqa3CiDVbd
L3EFb50Tvj6q6fWCg4gxKebmf5qUDxc0k43K1NkzaUZhSECE+W4quldmpMAzmja+yW5Sucv/Sqxz
6YjhidN0BDWzJqjDZmMbYoPyjM7o8UR1TcGe8EN6dWfiiaeMZCaaViVsOSvBkaz8XzPDdX9FbsbX
zsXv59qQxS/2l/9J99uBooGf2Smo9M3VWmWlr4VHQf+nexW6t3zFTfNMwkKOeUvhRsufYAN3pxm7
pjxeKOq8A0h26sDnUbzuzYHHqRlIXMTZNqw9GN+p/jWleSblpH/Vdxhllz3yHfQewTRvbviUex3O
yVa6LcHoo8/5r+UO2puxnSriWnHsmHAjDw016SniZn29vk6AjBtFp5YxJg8RSTRRV0Uyfa6NzNuK
WU4VFTY6dZ24qRYDT9jvy0NjdGcwTEDCM/GOgvU1u9VTtwaOCR5DUuT/VGJQ2FliifpmBtBSQ0of
vxAaXhNsNkHJjaK5WTLOMGrExgrLVu/BfG8+A6Gk8XsxPMLW0ructjyqVpQ71tcGFyBh4jKp2jlN
jDZMg8vcUwgudDpc3Nph9bTvjaCZITOOR0QEyT2R6TRkZeOmgUo+Ehxkgmk3TWCwmL1RMsYMAjE8
xVadw5gsS602ALdhTcafQIgXpYl0mfe8v4YSosr0Lad+4ZQ4VJaoewCtevKMgv4nerx0IHzNXGYe
w9dW9r3eJd1lTSTX2yaBboZWpZjhZdzr7hUMy5A6XY26JjqNInatjWcCMARBhRWcXIYJGzv2fLBD
7tISUz4IEok2P+tuIDTh8PmGXo3twt69VQRErsDMQyGphm/QqICykuA8uJ/GGFKJrif+DpugbyDm
tOiqDXDwQEjEgAUIkkh7OJfntPKnN6314D9/11NLWA+kzEh7jk6nSe/8kVwvUJXdO33Sdq64rKA8
cFcErkOqXdXiECy23JTV9GzL9L2FSv5Kt5h/uuLwAj30M1urcBE/Yik/P/4sAFDRulHD+MiWMW40
+I7R2ol1wb7oCmDE7z6d2whJu9iD/Yzis6AQuZz10P/2idNCV1V8dyicHnhB/iXOpPj4+7BZGrJc
9yjVeqqQAA+EYpA2XcSEu11eJ31uhKbFVzSjEk2zQvASbb0RZzQAAEf4h7VvUlDCgYb0miV8hUL0
qtWDoMgBex9WpCch14d6P2tI7URkMW7SCNUD+EDqtl2f5z1GYQjJY98v8be87ZHwvRNpurLnKYZE
R3AIwzgs8PGYxgQQAUys81RVd3Qn1pNKUv570/7/ctB74jZ98VIKcOoz3xcOz/2Nn6f66M77D+Vt
mlmZ8kXWzhKpl/xdShU8GbAc+lkdI7fCIsXeopxf7exXFHSqNs60ig82y9IKrh0RVHiTtBmQZL/M
ArZvryuhella7kMw6x4xGwtklYcjNmUS4J7cXafPQba2sg5LD6DiQDiS2YungvIsga/kfiNAc1hP
kcMX/OB2Qjer/1zv18gx8mqgCv284Pet8ew13VIcxeeGepFOfPQesNd3amPmIFoL6oXFyaaqVcOl
cZCY57euH2VGVgVcqeelsjrfeIGwLDHCtkrtmW8yjiUUYXsgwEtTjSfDiW6fM4+5Ku/z3NTLldSS
lam3PE2JlnP9NY9ao96YtjHd9BXueGKRRXUMzztwjBa1HMfgSdzPHZZY2WYbdS4vYhPq58EUtSf3
MJ3NIVUB6d/7wA6188DJHBnjBnEiuI2cpQzJdtofRH+KvrqCrE070NaJycY7MLxUw6WLPjiFH6r8
hqGRbvZod0e9Qc4JWFrU/HEkl7Ycv2TTDmBQwjcMc8Oe6+mVc7gdbdO1vch7fnGFfbviuyVP+wzm
M+4RfKemsOa5NHJ3QK7C8yYQk5U4JKHKwP5dajIzF1Bw2D9No6TLuDryGWEe0Gu71PH3kKMHZ71P
ZyA5etnR+QjTWj1tLQDySyt/Aoo3Wekp2G16cZZ4cGZvCAY/9vAISbTTELuN7/CgT9Ba5E0nWHuX
AffpNwQ5C2QS5uxmwvJ9VOFmz0p/rgBUV4b25VR0M6Pbt8n8mnpM5khbh5kgLXPCP2FSBcXuPBHD
9Yi8wlVsE2eFXwcx88GHkZHbX7VE7/2HIsvk8+cA812EwIFtXqQVnNSzV75cBCLksP0miDMludGJ
tduepDplKd3n+L8ztRwuz7zHDrwabxSIHFSNEfzTlVu8JWhdtw9tWT6ZFCFeDMHa7bLD7GleoSW5
9jV+kim2xbyjU+iSAjr2wRJp1FcpukSgeZTg252fw1lATtmcTskkf2m/dXOoGh/JufhyerSjhjCT
4uv1Fy8N6izHxO+Yn0Tq4A23KWXmVtTewF9jmPnHMEYd4be8Fhg9X7AYSKH4sEIsKVAQ9vOULDkg
dcczcKh/o6GR9l9m0yKHoy1wQ4XKeno4jdZ8YoZwkC9QhapIsNbPzGWPIk0PIErCg1bek3YrfFDS
QNB1nLwVwYt2Q884/XCasmAtHPqa7Mc1hWqqbXURJKGOIzzG/PQW3lxZGOUpnuDt3xyUSY1G0kTF
u1MxrfHLmdrsEHaALWJ7zYdRNZMgjCmd55CImGug39DmsxM541nvAcgw+DxZC2dl4o54IVG0MOQA
Ddi4FUpVZSq++DRK3aSweXrV3YVzXM2s+mdqKiIqDc4IkCuYWjsA610X8SKgnnYFU8OetcdTzqn9
TaPmLdj9je26FmWrpw1/0lW8ZAdVGNfHS8c9LrwemD9qGbqM31BEKLrrMJFvWnXz6Jqi35o+JniN
WOl7v+TdvBHMBN9WIGZPaec5VN5eiZMWni3xtusgNKffEaScVUkSyQ13z2zJLFNs5mp7N15g5sYC
I/ALauEvCNiY58+c+bN/snscPZ6HPB3YxFJckEyJxvCC4zhRkoRvBXaQoKCDsQ3+6wg2C+21oDnn
DYPRa19pzTGa4yxT6U/EGzWZQdEn9wQqQU5eJnFch85zG7zwXMYCZd9Ht69hOpH+kiB2yAkM1BGC
SojcxOsXCVsUK8JezeieGosz74ZVg+LBvQv4bWVw3f76z/BtRmVerXnLimgN8BQcxFRPVqDS2HeD
Ysy+R5yq4vaiGf2E8XLjeqPcJCJsNzBdqzIqgAYtwtYzBnwLJx7MDQtHXBHLNdRP+OTAj0/g3R5Z
PEzXqEqq2VQDhYZQQXVWpZXnc/Ls+95/D7ebuBkKxcvs25zYbPWrzlNbTa2HE3WMGeV9RmnfvL4G
jBWE9VbeH4FR8B5YHwUPNgIfrR3KzgdQDXhbH/O3C/H9DHxEUUFvl3enItW5Q7Yw39+JIgjI0rG4
MC5aUvJtUm2fgJxwJ+KZY1Sy0il1jdFvCQ9GCo48wmXyXeF2TJYKmB1F5CmG0/qf4f8WX9z6QOLx
eIQzkM32xr/y3ilMskCBe7ggd2BXBBnjVQEBsDu4IVu9zzy5VlAgBRgzgSfzSnDHbTjSdgSsTvh2
bPX+g2y5XHHjH/igDYQnlrSCV9dEl3a/kysCwlCYa7YyOH4bsdGvRbANrR1bujvWd8pxYdz/f3BQ
1RpvW70se04l8FjoenViBJLIH1RtS2D992qEQ+oVlVgSxy87k5Nb3MUMHtzCVyqxseI7Nsi8sivX
zxMhCiehBJUFDRPSGr74FzYqqT1r+vQPJZarSI68Fov07vUWxQlQhzTMeAY63UG2R3QNq/C62IgS
hweHOwpwGM99esVXDMMRD1oqVMfg2RPW+epy5V+UrwD6UbqB0VzWueO6lUA7d+HKPwSuxJIGXRav
5V59JwHJSmr7KWchNZJRR1DvIDNJ+wEMd/joAxJiy9pQaDP4mbR5zmllFecEa1vBcGZ4/nClIGI9
gXIiFcVQrDQvfNH5TuzJsLiQG7jeWcXJIWg2S5wSH5PKK0Dcc2OIxJ4BUizrKigwndXOz+xzAXGh
b2baOskByp/hpdw4ItFxa/dLhfmLCHyASGs1sYfQ39cjU9wlK5gf11nUmoeLgQW45btZHdX+Tkm1
29q9xaW92y/Fr1CH5r1fygZiQSHSiHub5IN/I9OJEmBTqbfnBlx0uJGpU11XZT5BTvvSII8djZ+K
V9nJbZgYdonXIORStMzRdDdmSM+xQIhzjAIsaBvMwC5sbcx2xSFCaUH9/lTdkXLwU7Opc9WFdHVU
wZMdC80bCZoIam+NmG1AaRYyzgh5ChDUVDUoYeYZi4u0eAZ4YIiJTHrUdwQ9r5h+lynL+namobAX
t6Fn0uqQGkTlQXkgwGiGgQ/o717NG42px7EQ5BwgUwi7HQLvpHwWwPFc0Bu6bzkczgXjks8KR6fi
EDIYLRwXTvlv3zmGP3kuTeTbFKP+gkMa74hjG5iTlLyuFR2U4VrxEHBfYUVorZlzNqoe4JKnnrYZ
Ijw/dSht9ri21fj3OF2bkWMSYsfn9PcGZQHCy7gzOYRo2QqK06Fn1/sTPgfSqRH/AMG8zE8zutYa
W8y7oewN0MV6r6QC+yot8NAxq/pF4KqhqeEFTws49IUBY80QXnpCdXlULFvHHvN64pnLL3YHqlo4
P8x+Q2hRvKHOVeq6pE39Ef1SmJqnAiat9hRMJmLuVwf2FOgTeyEf+n9yMMlQBFwXa3blflkl/lWL
Yv2lDlhBp72oM89q8SVRxK0jrvgeUChFCVdZVMmS2UbWjamF6Er7GMvKqXmErzeCYoec7DNn99ni
7VxwUT93LX3vAzDfktZ+1jwKrk6X77IhUIt/WZ6oumoCtcys59AzPtZ/tVZQGRqFfKVFWtXvv3Di
JT9Jl/daPgy+8wi6YD43I3Ofw4PkxHnkK7hXaRvMJySJPnM+WaPpMB2tGURLDMW5I4nUPtoKmy6w
FpP8RCzWqszMJPDn2KYuCcCZT6J8x5NlgYusIQAxDbx9bSIrR9sz8+LTxrn5rA0qB4qvGC8UwEoE
Pg4HmvE6UI3nAnDa/5ntlzEZV+nPPu6JSRETb6ThhOXikaE+JTiPl5IwKozcpWsYNCjMVSsVJynh
G70IpJrBhiQWlrfdwT+Eljl654I0aEMdDK3LgH8zRoLInH4fA4Vb53kSS0sSxKlhS+KRWh9VR7g2
htxs6FS8fjnJ3kf3m4UpEZjXieLyERc50tflr6EKqvAYqaDZz8cBnNfBpk46YKzhmujSHo6zTBD3
91P4SHJvrk6EjbTvrToEoYe4DgIbNg5FBjzf1IVTby8FJSxZlI9iqd3hPB9+6XaWiXIr4UBsQFku
0ht5RsMrGPlUBt+CK1mALVgTvkXFrpEOpqW4ywXwR8i4ID9hwwjgaosbSarLHkbrjjypCmOtOQsO
mTSTeGIB2cbGXKg7BDNospMPuiGTVumQ3GVESQnUT1Jo6Me534X6TPKc3czGbnP7hz1PLmBbmOBx
ZZ2sEAqosgk+qXYj7O6EW4QMSkawEv1gzb1tkSBul6pFbeiIPy9cKpVJXTKHdmLYj1E1C/FB7AWz
OYgvwz1HMP0J6aRlwJ79jYZsw1dlO4GHPVRhVHd42Yli4k5S0i9qIlcKhVMekLN/qU4sdJ2oRg8k
ZCyt4TfvpHHnhF3PEoa1hWLZtJ9nU51IOJx5LoMibsWJNna14ClQ8XcZRMXvKbDK/E2U5iLBANPn
hS9fXmI3ZyBamplKsr0m97QoNRPlM1vZrlIjFIvuVCAnJVtiavEytdzkZkNAqbEqV5MtbV1EwKYu
orghflRFxK2Z/R3CJM2qid8qJ07Qi8NNGDyt97A5ABqbyON6TgmN75GTt+bL8vHyzap+hvQl2g2e
1+QaxFo1DLJLQH5KwjwHK8ijZYIAJUttLPZor3DEurizr1jSR0gfg4zT2b8ARs1iYYysWh+UZAfp
GWGW18ehjY2YKjdmqlslkXX9jcZYwYF+Cxzb3ReJGgIQwOjgL6HWRj2GM1XjjFCihvaKPB2X+xe2
niJyc2sZatzsjQ7cpryR/I2oyg5wBmc3Au8oKqypNPnSxmUHGM753ZWAB6vjBF+t08/3CpafK+6h
VaS/I4uIyxeH3UeNz/hswPvMXSzSVUaMzaHvih3ncWxZ3X9Qwknlq86+J49X28Zg6whKEkslQOai
DK+4hg48wHBWsSZSzjmn1zE7DD2jK2UrCjHFReN1cAWvn44xfTvmfOUCYIWM8LtyoQOJvoUdGVPD
ArC8r9dJ/n8xACpEoho9HLib3kU0nMDx3xI6LO4kKCdR8npYePMlbZ8yOpzw9joxVr4X/JAxGGE0
VHMcV1gVONpOw9WqDBg3pcTljO34VfR/KfVR8qViVMeogz+ZLCNesFADOYLzV7uOeJbsBrOwIU8R
ooDYlL1RLZLGRF1Mp8i9cBqR16aZXdVfPfmNuWODsP0rjz/vlO44CwlqP4RDNSW2iJL4qeQlqrwp
QDtnd/CeVPgZAcTE8trFu38VqpDlh1Y4hezHU9O161TxTdQsfl6FH4wNBvBj4QW7SEhw5in8ad4y
RxKaOOW5QFGQnqx+dMiC7GsOiTE+KAhrkvKGjGYIlr/zQGuX/xHMpE6WlIHiLa7lE70djbuX2YOe
WDH2si95ka61sm2/c6UZOGtI8NtUMUFfEmSfJVL5babppCM8fLwKdOlqGFBtBKZp18ZHZUsjNbWc
yds1fot5tDha7mYFPB8sVvxXZBVl7wjx5XSSVWKhIxN+iGhT1Zs4Yngz8JajaOFUJSuLcxuSanDh
xM+fgkVKeL+2nDtn2Yq5P2gfI/7VXPa+U9kNSAUqbMdn88dkXCVg5FayB3mX8k8oRJUWlMJR33to
XnzFlMx0pEPw9U8qXRIX8GhSD5ipveB1XUdkPtksn7SY9z0MUCOCTV3rchYJa7Sgtjbsz/khr9nI
9uePZk3jXfATdSqyKmnD88PeH1jrxbW1Xw4kxJckIo/so0zEtCx/1udOyVkXWMMDSwptakyKmUYq
0owi3PHtCsEXutpJxLK28JE5G+CJbIm78pFpFfPxeaGwWs+s84X6k9iBOolK6A9JhegW57hpanlj
9mFvmbb7qSvLuSB48AOkioa109lwjwe1R+sx7yUnR3qaElshL9mV75t7phrDBLbostU5d1bQZhmU
pidblqRWiU3IeKQM40cruZ/Lil32jpF7+2vRLDRGkTBi+josauBuyDt29l5kMncZg8wETrTdUg3A
EE8nBeAknkXBgZedFInuZiGptctuAaPYDaqMhib2nm/rnaEJElpaX4UoRK++UASG+9Cnze0qTkL5
YBS79lFKLvnRqfbu1kUtXgSzD8srugSiXUjxJdJTCjvIoPXEZJ2hoFsbQ4CpytP92HA0C8asLqJE
VGZXWY6uKQDsmlnscgJE5FEOmNf8UvYkO85Mzsm1ag+5eMAVLzlGIfQahI5yWHovywDdKr5Az1K7
wTC/vd2qe6jW6vmnBlcXnkWPl0J1m1xrtN6tJHpkIU9zE7lFga0m9NaumkSVjdlX9qbaf8FRAm51
dCm6mdHbV/+j9/H7U89pLhTHW/3bZdSTS+V+oKC8N67Y6GFs4NvYkh8C3W3h2g6UNDaVIC7Vt/uZ
007Mc2IdUF5tUlYk8AZFXob/vBCOFX1i26gVtUyismmr04fiR2KYgUHiUygk0+bvrH+ydGCYN1em
Z0tYJ1Y6mUl8aulXcnDWwD5zR7cAhCQOcXxu24seWJNfQELzr+K0IrmxHaiJnZM9nIYpDxF5hK3w
V7YPdSrq/WFlpbwTnayp38r1RwzusafcCDt8y11xgzXMSIoKqpnerq57ce4VtRn6bB2zbDbbvgNW
GxKT8Wk2Rt1aG127SxQUdh1TdTZ2ilP2WhLgizffpf30oqDIQrezaORKiTP0JmKS1yVzJC7hn8UR
QY8W3WKP5GDuJcORESrIlF1zmoCl6KFNYI1P/jIAbkXccC9p10ZtQZlDcLyQMTZviyKgmc9ITO96
PDuLDWHSouB3ghZHkPBFRAb3AegrlEG0q3wBAhRoZjWmq241lZaFgDwXv61teNeARm4MZ8/tIKea
68YSfkcPXWcpbfg2MWapJcVK72NlbURIAaLo9Q7AcVP93yRPPf3unQCMaqAVceO1Gd46L+gfO4Sn
3Da7bBQNWESplpEAwogZ4qG4z2l+Kn/SEocEFOOmfnyLwXpShEQI1w3UQdJASBz0ROz52nSyWhCG
hV9pzcBgKu+5+uzHRsUyAL21g+aIKhiEJXy+MzXeE8T+OArS5R9rABYjC+N/XdGEJzRfEXgc7qa8
TOnAA/Oeq05DQXT7DXZlC7phzr+g9reQALymXkZ9CYP10lhe5zl7n6GhqaidDIqCOllU8Dvl4ATp
lgH1MKGIe6a7/CLbU7Ko1nLXWgnhbcaOcbFytY4IdaBrbefSb7aqWQOJnxziH5EcavXa/mxfEksw
Fjh5usJJYlR1yG7KWoj4Ag7q/MWupP5k3zjKROIAj5Xpf443rq8XdjVhpPK04ZFEVwHrLjHicVUh
zP4lP5mf2aWj4M5nJ7VWRzh05LrSfrN4E1DQ49nJAkWkHo/cJYkXghX560E4ERNCvDSV4H11Spnr
v3od4yqHpL0oViyu0tjVVDjMgdjsbJUwkAk6IkrB0XwDOHpB340AKllbmJB9LtwRGY1FmmOD/L75
KaGACPLD3SGVb8dT/8nIGiXG/B5VUQlNcW++cauBwNa1E6enLNN2agYcmmNemqhww5UAiAvhGTVE
AkthxQCQNL2mHE7+4W2MQ7k3di5CN+nSMY4GZ7uOIg4QAELjQTDURAa2UELC27jXG6HRdbq81kO1
HiQYBATaZDvZZ+SefEDxE4OCVUJCK5Ys7+ptEwrzngsMQt20CS81jwpKVJ1U116tGuMWns32y7CQ
zt0erUAqmYkLBVcVpHXx7ql+A6U3VMdwzgca8l5oFqstVQaM9xd1n4OYo+E/p78ezsX8tfPGiGLt
eflQkDC6JbI5EnUq6v73tgr2H30UpzcTHd9Cx2craWifNWcmn4cxgfrwoADyi4PSDewUNWdXXqhD
OyJfufA9aSqQextbpMD96gu/DonWw/wcU5BDgbp8Md9gnS9zlx0lZN5m4SW1FM2mntR4B8WNWisf
mXIwOiqrxa+OZCwEbCszRkr1B4COMCGDp5SCoCG98u/JHM8eBcy2stty4givtYaXY+wSeAgGosZN
Q8lDFjdDXjTYido3NHz7KAJromM4zHZsJ9gbYg9tTquGguXvahilt9Uv2UUQ4N0r3o9GBvEItWZD
MrnxmQQYwmsBu1U2Q3GLMDeed1ACzHmpXh1zs+eQWywNS/Ww9kCuhoz8F9wCRSJLq8QAhL14IFOy
kYp+pwLn8zOPF6UYnlnFmQ3bxRQ21QEjZejSY1DFe5xpjCcvSunrY0IRB5bl4Fk5zLn48LjzziSX
erHRSFvykDdNHExzaNuQVycScbYhurvN/Hrk5zDQROCAjqTDYkkXxiHekSnArtuE/W1nUrHbOPtj
/N1qvkUpMxk5+miO7ojeDJ3a8aaZMrecULKNI9rEks1TgJdG9eSmGyZcCveJcX+gRJkkgyIsgMGa
dNlYzxOzm5+TVucNA5oJeCgao/NCcyMzjg1GHrBr4RH06Q6sbGkkN0lZG7y2sPeERtY9EAuXCSAw
kWkrSCZYOk5KgTiVowlXtBgII7810mNTMEj2L5gAWU03m2QV40QS8qtcvkg6kHsX0qE+GOua1s7h
x2ijlMLYhHdhCgFhCgNexWrT0JB0PD5U0ve5Y3fnV4iv0IW+iy6l6hgHpQl9UTH8IUXhOqxFiHl5
Ge2OxmnIPvM1nwn+kjY3eW2d+/3e98Y3RMJkp4J8VsabBpjNCq+ugKjhnFizW9KNHm90gf659L0+
16gcM/51sIP3A1sjUlvMBphi4fb+YqGAdXaDq6pOTQ2W+SzXViCBuwtZcPd0u91j7eO9IhW/rECn
0zfE3j29K/j2/YZGHd8i6H5F0n4vcP/6k6amafpWPKB3fKhO+5+BcYOC7JDRo3QehzVZKzBZyOq3
wa+qzRnrrrgPRvrrc5FLB0w9clR/U+qT4/F1H9+dx84i4ELRY7hCDCIm1aNp8D+5XN8BkgYmf6CV
v50C4BRibQfvNeeFMuHvr7rX8M9mYpvPjiX26QZeGPikkyDv9/UEhET0JtcA7gaygKH30I4ptbw4
aY+Zzqh0kXsrU1TkjfybOjR7Tm33PSZO1gCw8br2kif8E2krgspbb1d4+BRxwppPl042d4zY3mR0
qXGX0QloLG75OaDHPkHC0zVBs7GSXFwZFd4EpA+fgKb9X+enjN33CGunatlufxd67nAk9EUm4SwG
wldEjNYgo0X305SQvqzVo4lFaNmphPrf0cCmbLnjInD9+wr4/c8Pg2cX9XnIMVWmMQru/vn1Nb2i
F8shD3ZTXUgbbOPvW7sIodg/C8rPOSDzuCeUcH8SNPbKUqOQalT5ibF4oZ3vLAfPMGOJ/4dlungb
OCevLsiDfVSk2SaWoFSJnSCJltM0w+BWKdtPdgnV6aamVwU/Wmsx0QQkOKeMTIc/ZXn5XjdGPOpH
G0MIynXfYP40B31aRvNtdKpiQ1eK5f74uIqUK+fFQ+jDhcKwZSTpNCW65RDVi4X1HqexaLOWEh99
IdneEdamYsaSHGj4l5Akk5ecdzTy+gCbPgWqRt+pnC8ic4pSE+Ese6QHU4nn3UFcHiFE5epKPAjo
zdHxiPmGraM4wV27RnikgD+BZwChqdcGDPxWV9zJkjSYzftPTZ4E/gGSbUGE4/c7ndiecSICEOmU
MC2L1hDT8kJZFGjBkwXjmvwDyWanT7yUJstMGG/qAX/Y2cadgy851uuF8nI5UMFb786qYFdYyPAQ
nvYAjqsavAF2m9R03jsGZT0DChZkz/qu4MDLGUDX60aNHfDF1KBTJtcmbnVRvJl6sRRPuNDLE07V
VvyH8rjrggaiKYXAkyvWRbyhuVgGbTK3O1eFL+ilZkWXYf6Z8RgDi9onXaUm3DagvHsEKU4VPLiH
NsFcKrRqz4YM4sVLpeKPKOS5QVsdWC0d0+BZtN2iUfU4rMYl/56YOUACw2VqtY6dCqkdSCnm5DG+
41bS5MgtY6x7HIEinvpUlsTkzB60aU/fMZlS3c8kFzfEZ0ECJMGi0ZkBki0ZHtMt8M34SET4tfJB
0PZ+6jgdoAe791BF0thlIjKg8MUsboAqroigeR1DxUZdVqA4zpp/zqQG2O53F5WTOR57Nwri7mIG
xGPBtm+AJaQRT5+HjKmx1JGNTZdmEfihtXqmn1t2Ae0n6TK4rvVZBG+wpqti5brI4EJdNQGNz8Kr
vK1dVMR4I/q7TlhVk4hpq8Q31ilPKftsKEwbc7b2uPw+Y9sLeYRqIjaBsViJ35pCgs3Ubn/tv4/Q
7P1OdlKFoBep0ZA+p5dq3tU3rlqQD59/sw38XZvPCjDNL22qQi21e4dAB9ij+uzxNSlZdANNVhox
jbRssVHsRKjWznQsDNVz7LvtmB/8+ddh4CCyEQ47UHGPv7k1SupRsHIgD16KZ+1q7QIRzMNB/kML
ndEEfqZYN+x/zvzb7NUHtbsZGxdv+buV6UP7WJa5EWWZKNWXdRaWMK+CBzp2zw+v2s7rLt2Sg7Va
RO45/DsKQIUSB3w/14eX15YSmWm/ERWE4EpBJc0iVLWE1w5Dfg54HjFU11xj6uFQcvp6VXsm4T/F
dEXyp3xnFQYeLkmy418qZvB5Iu0T7nAx3cw0pxfJ6EPf/aUZHW61Jh2eD+6Kbnp1v0XCTIclFNOH
XdbG/NWqjb86L4pgvpOvSga+BcpqNI55Ugp0nvXfxllFDGcV72G0I2qYqAngIq13FfER942K+5Kt
mFIkBKpyHnwwZXsStcytwcob1KBmxWiipsiH463WkP97FTJDS0bQsDSfRb1ijv3JAWN+wAN5hC4A
lr2FXnTlJJmOy6ruVUQ9NinHWxyZUdhKixDOwWezTC30OEfWgn+mSQUa69/VamAUSv/BUz6vTW0Q
tSPQRH6HPXj3ikl/Fs+zjV7zo8L4QkIXdB5MpgmBt3fCTbp+DP41FJMTejn2lqyzbpiptW2qI4SX
IW03TbDIqcH8AI/+6ysoxfZUU+1KnODJC90MektGyeCoV8sorM7Fn8N6jED1TegGHLdYgxx1xQR9
rYCV2BUk5vyEYnOEsyGmdbmEc31xsFCtsWU/W800XfNWl7rH4BhSC78ARjZ3RG/oMra9VqEr04Xq
7qVxMZMKa+7XrHmyzX/ZmT2nFjXCNOet1878uzxXC4NMix29jyuP0MZGCcL5zOQg6JRbNOP5oUlf
mjLnOHI7eRvb3v8GOKNhBEwFxTWKKwNlwJd+Obj/thrg9yNAy8tjqaOrZKzDNxqCGeIy7WQft6/u
JHygFBXX9b0LvPSg20z0jrFqW20rN6M8sMhZGeFl8MNMAKuZR5+FAaPFd6Sx8uK77FwJR0lmWgiP
gNwOulV/FcprlmUlOlta98ItI3xD1yr25PrggRtpi359FWruPc53FQoIoqWtpeFn/QWbI7RUifji
SvGtwO0g3+16EhwjWutnWLlQFwXYQZSRlVjBfL0ikrIIrLLCIpRQsShWdFg2herYCyRy4K+BP/LZ
PcewqX/uM5L5XcQdjW2dA/eGil2ySFAzn0YOmEhem7trP6EFxdC1VnF57yxyIwWLC/AKPdfuJPm3
FGm9XRqQRAp773ruG3SbvKV2wGHC67GdErsP4C9m6GWbB8WGfxkMu8o8fUwiViUiiZgQuF1852u4
H5RVzmyIr24LhwWbhMJMPNjcg3pgt4OOs9gPADOYxDx/p1Ze300P6angUNzW9jCGMxj9UObwxPzW
nnbK96VRg0MlbVfOOhlf1ax4S0wgbxKD1bVuPE157rkBylumVmAtmz/Jk+ZojKNB9ASPRUbnymLf
jsuJFyHRUWhnjf+mvYjUjWkgD24cgrvgDVhmJhScQRwQ+ZjmSnSvuIbK+Q2GsehAaAfs62w21AJD
xXcootMN7GIfdFCzS7cicAbbe9GdNmc03OVczeMcWnwDrsZDq8z+0YZUzNJeLKKhPME8i1TVMkRE
B1PGuGrNjAA9+BEQfFrz+KNFo/RQ1bfQJ2iHn+3JzW6EUdgvdgaBreNQ44vdDbDPNABPVm85A/F1
UOJIKM4Btc29tmh6wpOa3EjhdgR4YceLBBEg3l42GbIsK5kSwVHSqDRSboBrGbKpYxmiLqDA/It1
dTVCfPQcvn8CvW8rfXs/zrnD6qu9JkhMZ7/Z2kvj0Y+kXxpLrqikoztrOF33KaIFNfH3ehVhTpTK
dynIq/VV5AqpP9Nrq0AruizIfPAuTd4Aem38D1N0Mry+Ey9thMzcetlEmFKZw6xtY/TuX9uY69V7
Un7TqZJbrOXp7Xbu8akLdozdyX7hG4P9vw4c1OPWByDou8PsF85lFXl8kiSVCkBtY2tU59ASUV0g
yw0CcGlQW+/VLxVT7Un1mu58Rxt2anyx59xd1wbLGe4D8jQWQ1FvuAi08XlSrAwtIgr8Ayvwnba6
CI9NwqOUE8xF7YxU4w6BpkGkiJO179VjKkbFDwQacfxRp6OgKaRfJfFkYdLFwPV6cM2lNrtrZfH7
UbzQe2yEeTBfhPWPCcYRdkpbINQ2zQqxUnK8m7cvBzV+mPVMhFypTg6Oz8lxspU2dGRCsFjNtptb
nvxhHMIujnnq0CGLjBknbnOdDJ5YwTjYuv2tI4RzvRMHrSO6psFfirvj5U/S4u6gQo+8zv8TutUc
cY20+uLG+iAwuEpwQzobb8r9ulHeeEt0rXaEbG2stAJExd6+JpNf381drh3ieZ+VlIbfu8lVOGmC
6sBO82UkrxZ3wqUitzFZ1PEYSCe3xuCjGQctieKD0fW/sA+mJPTJ+QDhPSc9E9J1j+3HU2a+DiRT
+HnVz9OfLwNqbtPoTi1b2bc2gRa149sGpX8YaKbkKwhqqFhz01iJ8bislFZXbXrdRqXxxCGuMxNk
YZfuC70H8UV5WQSHpzvj262CUAOQzvB7l3vUl3IJRSyhRIbIVnrExmsQxiMIYsx8SVzIz6/TNLeY
r9XgY6qqaDsc+lUt5X8NNeAeyr94wv7zNs67n+VFMZXd3j74ZiHxtFP5mBLOpYn0d+wz/OyjzWUq
DkGBN2RYeXsaJE/QufkbQZ3S5Y5/mxUXjzmGpy4vhk6fZiKi9buxvTu8PG/y5RVi7YippXov3hbl
miJYy25k8WgF44N6qHegri40nHutM8mIPdcTVNHzVbbfg3m41r3po+P57IvOX4/A5uKsYF+c+Yne
g7RgGE0h5RUIUI4Mb5xAh7xrb7MQLfCimZKY/PwI4kvOWLRW/o22o0kw3Hd3XkNkci/8oe8woOvQ
R2PG5AmMnq99YxM4jkvDbvG6EAZXVgPD5CDZYJOhb9m6suzBkYW4JCHUql83tvreQxpc6Qt4ID7h
A57aL2bgS+tQUp/CSym0x3egaZHRBKDY/c4StumoDIGnr+3pbqAGUpEgr+ijuoIpOQb9GIU1C8na
Sd52cpXA7j4LJtOB0W+pjmbOlaL/2G0vHr1FAUg57lE0sSfm01NajKqn9Eol5Wh8EvKjWqADk2mZ
p5S7h511JLmFqt8KixCed6+YV6yH9dZ6qqrvZ9rxDZakOPKsstlN1Yz1zFRXUmUOQKYywUa6dpim
EmHfUtVxGUYDoWytMXFB34pZzUyUyjnxb5VftQAnU9Dnw20JkzaeNv5VfFPLt0Ky0Ye2hT2Mm/Wb
gkBFy/mVmawdtcKvAY+zKx55SPJ3LlMDOcl5Xh69zN7lPf90tnscUGYlfHwDusX5NOEWYj6qh8//
nB+MGxnvMNcXb5/CT4q3NH+bAWodaeitfoVy3U0b5fB4cx5AKTdDXvgB+8qAGqg3cyaENPJvjoSD
DFYa/MBK+jWrgGFQJPy4cqgzw5had7vX870IDCQFJ6teB82teyYuokCCVCMCssMMltYqBCST8ZXD
2EthM8qAxvTq1btNBnE4OpEmFcDfQwD46hxNF8y2ilpMQm8Tt9FLkXpCdULnrmDRLc4Yn5F9cJnx
KxMiHMQ22gMLODbfubu9k12rPYQfsVfFAN+mtvZ5URsAl43iuAZ4zUAcM6oMO2sUIztAQFMvFZIH
MdIHvuRSgGpCfdXZtb/aPbucNSLSTlP8b5DvC10kzfDTd0ANVCleNKNzhJZOnljzPPBjlA7kFTg4
UdxSwe687hdJI60XY3Y/xXlOxSnJXxM/C2ufc3pHFlRoXpbcSsZiM52NTFdmPc/8GVwHLRyU8a5I
MQoOyDdhxaED3BO9r7nzNXK5Rprh/XofIm1z6SXMqv8gnzpRMm7qDz1RTyhR5ThYR31YVEmIqLp7
vUgoZESviSHDrOLezRgJ4RA/DCwpaaYapP3Ly4xu+oLjYMVxm9umdiXorLHyqDZ1EC8BHYvbLHRe
PsvGfYF22TeKOyQw2Zwvm8Pm4YgR2CGAveO9Etyk6d1/ouUcyj81gNiSofwkXv6R/81kKUqBKvLf
OPkMdYdUL0C/Lt0yZLikWoQy10n2+TyvsZtoYbU9C/cAXJ6t4PlE7oXZ3CyeMo4ZfTeUdZXCUAIr
ug9MLoAPHOf9nsRUrp4rGbZ5zGz4JSHQrwPaHk9RnTAKYhVSAj41ItaDmmAfLSrsLTs15QhVFK38
ix4+ACN0eXg2wCg/SShaKHku4vzHd0Jrmjl4hwSPVgse8qSf0YiUdIIX0FTeD64e4akddpnP90M1
e9qI6NJm4UJQEi96S/0t95dNqT88p0Lhc3VJ8R35iAPWztPKaPRt3myk0wa5YL7rqVvo5A0DlE7g
J0G3+Sx9hHCRCg/SxNBQa7xdFt3bIJSkqZuSLHABFKzMumDIp6W316ELy7XAWQko04jSu1dYXdCx
uIq9tXPF1pAnk4w+GUpOEc29zJSkisMbr4t24zeZlg+vuLkFM/ogz8By/RBGe+WyTVHsJGozKjtc
qm44yADAD96Rr6Il31lgaWLYlv0l4F8tGwUXC8GHYQgqbIVgRnxK8K8MiDG7SMoHfamm7H+AlcAt
0Ff4g9CkYCn/AvERS+iy0QOLY0wzXLpBOcA+xamBAHwgXZ2y1e9pFba9A0QJwZ5P78na4b8kdSPc
DZir1vphi9KcFacvavKlO8i2udNwVPFLt6veATcO6SzXa48BX1sm1cXNaZyXAz2IXY6WF4qVWiKZ
/LANjMpBbGdLQbTHp7dPio7r2kouHtBn+k5Uh0wc8VNVZaxxHHfVu9btyTv7pWO7ayYOGB2/dy2k
gJAcJYRrOBiTWKNgApCr9W/ogZDr9FMn6X0Otlnv5Aru/1iS4UGzwReZwsvF9VQz5UK7Gf1Jy6Vf
AfQaz0NNwfcE7bAbiPV0PyCYMyGkKMPctQUHzHxZn0qOI+IO4+SSND/mmI0OmHoL+cPpShR2jwWF
Wdk/is8GoG5lTxTuofMs5E2U9ITZTWhCNMLSn9m54R0KbxihTzmG4BXlJchUram1DJSGqcdFBBFy
YZ++J2vUI4G5nvaIH0ZBhrlIH4Nd4YXZgei9zor4Im5fslnrim+YhyLUgysJmTxQcX/Mip1a5Hnz
9NN4ne49KHSxMGtJt86aFWHhpLDPWJl9JkWrCTTXg0lAes1UDqoshKvwSq7yRNAW9aZpYfjAziJB
Jn449kGoLpXMPg2xd01ZpTdeylsv8mZK+AqCXq6f988OEiQu1GpaiZfKt5WSHbt01qmCSFf3QZL/
aZAckTpOy5SHh+wjsD16Z0a+SSEENl5aLGb1ngrMtVBitV+NkOiKTf+gJuIZ7Ql+o2jwZvNZq79G
5M4AwvOmsgqHUq7tlE9kZeb2qyWwuMw0kpdIKDOgCHvEr6o5H/L+VNJe1jkXR6fT1EvUBcMsQ3ZJ
I3bnrfbcsK8ZKTcwk12AscLpbG506FM0hqMfB9ilEQJcsc/H58PzUkU3sepygqE6e3kqndLDGFaR
NgsfI8B1bubDgwAs/nGvy69XdQHhUcL/B+94s04zrB3zu9qL3EmCs9sa6r6UH4G6ycowdP9oeN+R
f8oBe0z9hNZJ1eO3/c+s/Rk4+4VRajaB0MlJIpDkS2VmWM4V6o/k+GT4bnhUU96EuBDjLKGmLBVo
ixhcQrULSX85jYqnjA3qa05sEG4B706/36wKaDAEWPyQahKSUR1uj0+XKY+w8EkNBSdIg2lVjK6V
6Uy+AKHNY8oDL9W2X3RGZM4Wyc/8y9H1AbDdsnxcxrDXjcZzn5+bQU/8LAhApIAkSmeZg3ASu1vM
mRFhHDBvhNBQ5Da7dSe4QurMQeZeizbkRAWxFp7X9LIJeEmSJABo3LIOe8MleWpIsjArh6TjnEDU
KYgMBEzuZNNk7qlCb2IAyhBpmPqwj5BGzJ+Wfu6xiK0mNCORO6Oaneu5qtY1NtGgacfLvzWUS84g
dj8aNRRx96wsIZQS9/vk2xSapFDOEqNBT8jmgL2T05e5BGX9f1EkLyFBIODIATaxSQOsgw0aZ9w2
Hs8h2Ogwd+EyTtP8q/UUUF+ba7pbFfT7AetK0N7IdWehV11LHQGVDlXZ/tKhRCR0kyHhPetiEO/M
/JMuhDP6mwCICWx9TYKg66HKB7UpE0cPHtHA8ib+qxtGg0416eZ13TMDHKz5qdS27CgivUgnmow7
PX2lAtfD9viT3+T4APCj9B0qW6Na4omyR1qzE7kRe2l+b2lnJNE38ZS2sPuil04pd5wJVSJ/rP7u
hMDwHND3V9gWgEy1yhj8Yxhx0qVmnKZD2ON3JHRjqb/VKAXNROZMdg/LC3KE9BsA7GsNoShicGM2
wObDyDi0KtHYcC2bg5iKkKmpvqC+9lwPJbWI+xrhr3O/1rI+xevBe+u3z/+J1+swHVEJKRJhY81x
12S+gQbBrn9ih564ejqb0QM+zLT9MfKV8wI7beJxQXnvoB1CLqlQmzFleBAd8jB1Il7WboUYJQiz
AzLwBeB2uMMFUYgdYxZeevnP8LMbZwJYmM2iW6RAdBpvvwN08/89j/I9sGsiGXyEYXBICkpkeB1v
x6vqntuL8LB88HF9tCW92baAnX1vXsOyfI3Iod5SXeYGOwoicG//96JwZB8PWWtBehsWNX50m2Rq
Bj+Ew59R4zc7FpFMkebsZCDRflImJx5uPMs3t0MDwC2Z0zOVdzB3B0JnUZOzvExkvyNI4oTEagE6
iITjI9FZGPOckquyMNZsUD8C8K4XnsJXJ9ww8u83T7JTEmnAdoEhLSI4rWMfmX4DgDKR34oZ2xgJ
W6yxqN+n6DhujEmaQ6YOT8rgzkzjIvl5DX334L8N8EKF6AR9Tn5nT0rkTSw0RgfjjxOuBMrfAkcc
iswBk5SysP/egGwyqmcedawAkFl7xSPEJpDlt0z4iBMRzozM/VAK5w8dbfyKdxlsto7GJ0/Ati8V
/q5hUQDIcOTP86H1K8D+/d4zAgIjPp++/zhH7N0fFmFutjH+dAcGqlcOSprlGNNba++wlkxHoVu0
/rw/Vv01qdaKdi8JYDC2XuwDX9ZhbGtwFcCHALpK7pSTjWw7G/lc+wLnKcCaMDq97r4pP8oAvHiM
cVk/mMKTK4AOtjCKTy/n7RgM8ATD7hNL6PgUIfpXsgBIdL92+hSuhb2MnsRd5+ZJiq6Q/qHbv2Ow
0iXmqDGtwIY+rWu+S/5DHty/uSAoG81PTc+UxnLOmQSfnQSta9aYANRzzL1jwpAHVKjdZVCRXilm
2A4MDLDc1tGWNOIyn+Krw7f+H9Cyjf3RSQNX0grxeS7/8rQYq0yiBP5u3F4zPPe36OCxBYvFel0w
369L2fRC3y9n++hovpfxzpsQw1lUf2cSejGA0zBGPaiZFfoMKA4ItWE+Rf0tMemOie+x+mhV6dIk
mKwRQbce5F51VWdr3lyLdp51PG/0CICgHbmGKa26YPbPOYF8yCRyT9YCO6I07cftOgpN1tBqY3pL
9UDdE5Cnv/Rw/Zpioh6V3TIHeZNQQnnpxIPLCuTJCLrhQiVkU278o+j8wCBM9cyTm+MRVyWRyG0Y
FiL+I0RAHrybO8yOz/xZKHBXSpGI2WisOSRcZFHObxo9O8t+6Fu0i6ixCE6hhI5uX1Jx/nyTudss
yF0WNWsSs0CVBYHiGWlzpcindW7G7jpFNGonBOh0wpfpSElbdxn6fCb+hGvDvT9xhy+bnU01BRQp
N3nj3Q1PQdUmC0/ysUgZ1wL3C1QwZE5/VSEjHF0/itBEUGRkWqtE+wdLEFFQLN1AsD8LQpg6xcEP
5A7OpupQU+ffPzsRsx7K4vh1MKwLOEprN7uy1du5mWZMKvjsiLerY5qtwwxJQDFZMTE74t6xBLd8
RY4Dzyvs1fl98i7pavfOeQOIfqO39Yz782u20ZL87LApQ8h14kS1bo7uEddZxVtMiutSZumMEMnX
t3kQuflMP/wT0/0Aj9cyjwvhfTKg//7ZQkyAVSMdt0tRzdrTxZh8BmvI2JbG9eqydYXG0E0dr3Jt
BCd6Pxv/ZIfOrv564P4r2ET/ERapQz2bFOfW2SntbHVf3Z+Rrh0BspHe5skTfQhw0+yKHLV5MkpQ
axwGhkBkRoQkfvHDC68Xv0SuKFrUSVsD97mBjNpFV/lFxhxdlkVayAkxHWKaP7+zI9+FjxUB2vMe
jD0WvoppQJGBtjopY5u70xSk5ke69gQopWiN1MtXRZVhxnZ4+MZOyIgO162z/17duQE7miY0+Haw
OcTNBQ6z4pP0D2ph7k+Y6WhPw76wADRGppXS43jRljF4zMKdK+uF8s+r371r2CQ24QqAIf2+fzxD
i7ZkQev4118n/p8UwKTSJsxJHvuH8O8s2BeEhrM7zdzgQUZ53ANlrJdcnodPUZYlotMTcNgaPwcq
kTfo9emFev+GKikNa3veaJYnTeS6IOIPwIEtmhXZCGSj9fvWpIl43vvynfWo7GOg3C6bz3j726j/
dOdz6PNbwlT8GAtkPp52006mPVg+k7Y3suA+syQCfJPrp/R4fAdj5dbexNkAuPa34343T2Wwsl3V
za54N4ml66NiNt7VRc0vlIBegqWfCkRjw73It8x5HfROq1njgV1mWdtadmeBmxuCbXJw8wgig/ht
L1KRSgewIq4YLun1YZI0tGzbj8G3rt6/BANTrCWD+ASqoDZktX3TYFbzeamSuDagAJ9RAaXosmgy
mds97uetqOxm3I92cLZStEg0d3K+TdbfVlHd6fzHW/Ec6XF9w89BPwwLEVZ1+BMc/ndUG3K51FUv
jaE4/cOKQI7DWRV0Y4avJU2wtzgmYy4mJOU+PldMIrugbTAqwlHt3dGbSg+Z0oGExOZ6ehXtWwgZ
WsxhkXv4/LFy6EahxkGp5QvJ9AWEOyzU7Mi2vnh4KV4kV76Tt2z4hwCEzyjei5U770qcMH+BH4Qu
JBQR1gFYYO9hRs3Xm7/Pt8ONndgXjq7kWQpuZSMn/FvwihkZdbbddRUXfKW5lPmRbRXn6kKRZWNN
EBcy7FqCKmquoxGGFu9NiOFOmmgThonFiAX4e/XmwPBqM5sHrBwJO7cnZtH7Fn4XswyXlaoKb4sN
44NRCfMOD7oTlYGSzw1j4SXLkiofMEEzQZ5hUoMhdLYwUn61bDI002PkqV3FjOlqyfKp28TnlEso
FpizYv0UEA0XQZ9zIVQFUDCjwiRN8aHhBmv2gTL26N0FnVRZPhssvpDIZD5bY/2wU6jLCbncc37A
/b4yvR8UwQTK7GQQ/QhGKIxU5GTB0i0GJqhr8Qoq7uOyYujWaE8IiHaMgH7A8H/5aEZ3zSce6n5v
5vNhQNg4jnbmY1ZnR3HyAYAF0eB/OPK2i/hSrp/wSlDw2i3jde8GMdFKQUVwPpUBSfTOZZGn/5DP
UzRyecYIZsPQCSOAiwYw3Hfs4nEEHqOiW93M1rRXlPJbPidh6oKduknPxVAXOJi3pz8xFmrVwOhO
Lx309/8Po4t5Cb9taTtk0dV5ECa/bpBDlZF52EJA0NI9EQZPDW2lVXa3v9LTjLVmajWgbELD5Spf
CdPrK4JWnamTW8z1yoX1fBsEW7ZISQoUd4FXjr9bsqOlusfFeq129LkoMPjlBHt9HJFqE2dESz5t
KDG68oTiDlglHL2WawwE2rIpKmi4SuPOdGZPeJk8VQHP2uDV+2lWgxd+j2k0/2TyVRqcAXPoSufs
RTyA2JvCuERftjSoengDePYfdexHLnq9xcKEruwxWycRTy2hGdFcXJk4I97y0SuwQuRR74zbEzr9
a1BVBN4jPr/q64zAziWsVKFmvNjNhsUwRi2JiisR1StnlB07pdkoVKAwcFMePL4aIMJ89aUvVLpd
7vN1mEzJpQfTZSkRGUtuCkL8MtyS9LLRMJmbqB+LYe4nQT4jrlNFsOEuZtYCdqaZ6d8PoyPaBsqj
CpQWrEM5FOez9izi8B9vxR96HSvdj6upN8q9aOreI3pC4+MUPksAjM/mmxBJ9h6Levh4PYNC6xMs
R99I3vBZU4Uy+VCqq94zecB7+6mFhaxbwQjVX/vf+ylWFq8L/mYc8pytPArZt/of5O8umGLLEI6f
OgdChyfr3kl7gZeo9IPKysbAWIg+PMB76UJV+y1ZCa6oYFxug3wH4NCpFGELqVaoXzhpz3Z6UDFP
VEcS317u3KVgb3uowuCXlawXYHKBfuGaPjLBvVbUos6zbpwPIkbImXduCoZbkTPhbg0XuNhmrEa/
kTm+0VBlLMfAvSgKdVfIcL7Z3enilBDystg8nSNtQ1FRA05GA22Ma4nhOuOW+B4FelD4MjxbultH
iGGXvcomeWZSq9E14bG4Gn3WL1TsOfwybTrm2tgjurPMa8zJpFgKaBznLY1qQ4QWlSbJ38BFQURG
2zNZVQ7ebgW6qkW851jOS3i/cB98sWqjfpmPivN2zIfpZgi+BVuGoy58QJL2OGpzB99kjdhy5l4i
E+NkLMnBgLYgPP4Xsw6RHr01DgAb+bt8gxNu63oZTQexIrxXux/MqEphRcGmHdl4SGbmfNcnMRVd
Ge5pbqA4PfNP4hQtIcrK93YzdHqhrXeZyLV1wInxUQLT39oGlbzQtu2We9/KCYxclqibdXrOcUkf
TT9aOpTObToxDaFMwlZuo5MFVxgC7w2dbr/SY10tIRB+tN9qivHpBz7zbVP2BIZ46W18U8MIOx/b
R/T4Yq+BsIoqAUCw2mJuDw9DAqnG8Bln2A93Ep+O9VLlsL8/TIuUc4Q6LlW8ffZMhZeDznHIKrbI
a30tY0j5bX5hGJBmfyRRpJ9MbvJ1g5kRzRFyi/CoW8iwJwG1YvBfJCm4eGDRYbXrdLBiQ1qWUsFv
Ka8MriQUPpXqx0/wgGC6KhyjzK6Wzi7wYetqOKqrW+QNB2T0ui4OAi5cl9Jdz2x8iM7rI8V1Enf1
HIxQ/5PCZ6kyYx48SZNtYsEF7h3TSW435poxXnWKCiaa/+PxpaEpsJnSEGtsrgdFXX3ZoFKkp7Ss
xuOSXnxXn3+lEMwLPagd//bDOD0VwA51u2oRnwt0rElWvHTFkWhTSheyxU2RAJuZ10yKNp1XLu67
Ey2OPfU06q9muOdSvQzNqcJyWZJEIer1yr6qs4rIV8/aECtOGDoZuyM1frQ+yASwDM8RDEMqOKIF
g1wYRk1pmDAzecd2kEMbxC4ArwsfFV9QwSJo8E2rknzCnISA1ttHTv4/4awGNLSdjpTw0zLd15Dl
DlGWY2UbXQxr8yrMwDik/0AVK+uCQVObyFNRoH58YR6QyKEaWDz2jLFNToTeo7uO04iANFfFjAAo
sssWF7fBu+rIBCdtESqzX7sHVL98nV7J7MJ17pehbIhOvlOc/koF7y7Q1JHz4NOTKeD7YDms05Hl
AC7n5RnK3q3c+4fnxQv1JM3vKyiGvekTfZhEKNMrQs1s3Y/GotOT4OUc7m3NglDj7ededZ4DV+iQ
pWESwweetzbTUVSncxL7Q19K6U4/Qm3/myYtdLfMYg+j+9Wk7vO4mhfqcW7UIbyj54l8UF49NrAO
dJ4UONyb2iCywJrJ740lQ5RaurzV9xsgsuMsf9uzlM1691rCUpZgU7IOGpCDWbMHdFjfzsNVQfDr
FHPZdsmpjDKatDV2RS0vkG3HV2emUOEP0t8Pxyq8Ow75D/HzOm4c3gkzlnr+ZDCy7n9paw296L9W
7AAyiIjRpbPshQ1kTEdAApQ+TsvuNfoqbdIa07CZQlpzQ0LeSC768fG/zFeFNj8SrVzgccXExF1N
1yg36cneZ71Bdbvk8FhtaFjFQrzq6/K79KnYMKtT1SnyJ3UBBacahpHmxcEcUVsYPC27saonLwPW
cLzENafkKWyEJaw5KNBoJ7krX7wuaOMdW1VKtZFC51xPHIKRD85HoL7VxaeCTAT0zYbLkjStTHAG
ryqzGjlsohZFgZVwj6UVHdpuFc5fDSdZ/jnJ0pGzpDoaKodMpaoXTHtT1py2cKTYy10E4dSe25VF
EHfsdFrarmOTv55Prb4iR8mSjGr+u/KQpLC8o2Ujc9gvQyHaRnGY9yAxHTLECh3LdOqvns0GK5e+
meVVM8pXsQygj18lnGPP7C6D9Qe9gSQFlBIKwgswR1g9DbP6NP32cZNPo7gfZJCkQw2mokQsWnVB
axBcBf3hm4zPHCkzh9HxNz4cjx+OSzF07/Wcad0pJ311WSyHwkaSc4t0VQDSJkGetSn9tb4f2j1G
IafhgxWfC8ff7zRPrixSmQSzhMKmfasSBYtHHctl25T+pMEgzEdJno2BeOap/pcASS8NFBJN/d5q
R0cQqaLmLcTtK3c2OICBKyfkaYQ39lVcY1czA99O/uQQCR4/g0ig91f90eGXjVbF4oCrWeBljBfJ
XDH5LFnZG+3iDDbPThc0RJMHO+Fi9ZP/iF41l4nWFCCiekljiE0x/p48oIAbaTh2RNQw57ZEiVXC
6qKvYtxS+Pffh/RJTPzry3Ki8cz3shZsTjZ6Mfj2JA0e/cmmSBnIvtksOy4e3PXpvl+idKEBBOEp
UcHZMOZdirPZKv5H1avYCKKcvJsXHNraC9GdtmM+UsQgD0O6Xt/IQax+tleoM8W837LVfmsPdy3D
Tx8hqdvUA5HqO3HNxr43H4odgRb9uTuy5ZHL2IYu9YuZArGG0oJ5mbPDMR0P/7Xt6zCtwvzWca95
qlea2kxw/8/8le0ouL5aL0Wh1k1wtVs/GVQOzkcMFiSMHONgvDwZb8JFOhiQrHyOv1q1Tbb2vw5D
1lDs6gIor5qqKpyODvY/TAdXwm98vYOT0Tw2Yk1pD3Kk9bswElfvXGxcMk0J4DC6hAepMVH7sHSr
bHxhxLWIKYwwen5kJXZhz7q2CbZ3x1vBsAr6UTQJNP1bb/JVBgeNcbRf8TSNWwD+k6IZgrJje/Zw
Ft5e8P4KJZ31e++LAMRqWqPm9nFGDMjtFK0yg5KfZeN1LG5dJsZeQ49uzQhUK0zlkdtq450pJ2ZQ
eHXLxffYmQqexY3Ke7eRrGhXWVbHSAE4GrAyQclCQvK9tM3+swWKXK34Dsxma7/29FdULikTZg7W
dJygpE416mCnNE6/91Nn5cqOSRUUqztjR1+eeRMLhc/+7ccDfB3MMI0jb1K/gm5dGArMlJkkle+Y
wz0qebwXeN1VSqxy0a1YrEp5JUnHnRLjjF1wqyBrNmThqBSw4s/H9ZJawxO9pcmrzAaS8e82PcrP
AGW4cjl8+gCQKZSL38+rR4S2ZB3FLm7miuJkJhRDdCgR71j2tuZOg+hmUhMAQjzXLiriLNtv3OCk
By6Taj08wE0XsWskLOz9t69ld79wTOvPYcHRQWLQ1wHm57pgcpEA9f2NMhkc+e194b6WBOQg9Wah
44JNdartknamxSlrTxE4k0goEDTDfORP8BflSzBM1nAOU6YsI6ttMuuZGKFNmE/n2Ca6CFn95d6e
pz3jB1IBKr31w4KiNRMRYOkdb7jAablHyZFg/Vwv7gbYFK9ysUVzE4jvXr7P/cTgV+RY+lkIDGQK
7jnoyMMnfnSShS0uWyDNyLLIsbRPIAD8FhHHurPcZkuFNHRKvN94p3ZG2X1REdlOfjQi/CoJ2FSw
egr6bX3gpe6+2ab8tOsaO3aaY3EwvTrX45ceeSyzR8IOGjDbFmhJEw5pdu7a7cZmvLvjmCD82PUB
ieTA1uw+cbLuHLtTXpHcThObAXzVs+34uFTX6OTYNhlxmhvgT0hgpG63PsUPacQj0WIKzR88ouXB
hY/u1SnSSOH8Jt8n+Q1Ml5tQhRGyQoYtJK6YxOlsRTZMV1nKNDKJv7Upmg+6yLYTThoQa7ojWLDA
33L8Z2F3O143D/JkC3p7Z1HAXT4d/0LtV5ffjdyy7VBS4LRwR5BtEXFA9sATBBjulMuaPJLtDHkR
gfH/nqhBgkev/h/+a4r4zm7ozEqNuo2FMvEbFwM7YuwrTyH5g7ijFfrq99Gm00/NNMjPC84DdfnA
BnoFRryiqPVJgf1DQ+4vDHoHdz9PsBPTTnyDAFLR6Pwrjbv/lDDbLpqHdBNKLqJfD3zUQ+RwzlUH
oR1GIRhRsCxNMNOzSx1HfVyxhHPyIfYg28X03VrbzQCx8faOJUF0IV8hjvaK+P9JNC8N5suS6zV/
VyQEa71ipiFHzS4vogxdXHsQLRpzw05XZbS4h6esOMgnQveX4Qc4yhyJjDS0aduq532V1NDm2NC8
bdEC6R0Dd+CUrg24nNnctcLbd8zYt0g5tG1ZQRjt1i0Eo/rIDsPXtmZZCMWOBKjAXSkC1LYYuI//
1MQ1KCfJbgXe0b//ddEMSX9krVD+G2lGjS85ZoJydoOsiAI7H1f+gEKFC6ZpZ1RVlLe9DqeJguZv
HHNmR+7DFX5OQ3XwO8BsQti7nXVX4HWAf5Nms/fjuFcVsScz8j4mn/gNkuIKXwTLyOKWgRWKfbUw
QYWMumbBAbpy5aYi3HKgio3etnxSop7ECHCqas4m5hisnxRWzW66ZiEhJ+glHZmjoYYLsc0euXnQ
wflJQU+4rAKhKSIpWiovPsEliBpe2v359KB1IGJE1np+tYGsMLvauS6MSUNB8oFT+bQ3VWz7BQfU
cy11OOtno2mv7wFOgksy6mVWdXwbEbhT8T36dACk5j5VDM7UgMQFDrwcu/yhjy+3DgrsgSUM5VJj
tZKEsIltRPtcYhI5egVrq0K236sh+ejGFjdUS/BAtfiPFW67+ocsswHemZlU2rOLS71rFPjZzt8j
mt72CZtLfm0/StG40ioWii4QSaoHze78AGI65LvCVP5fcMNWK5RbhRofEskY+Iv9N4pvk1g/v6iR
prrAwYDzO+kHWnXA/AVznsW3Pb0QpD7Mc7mtK9ckwIEWk/vH+r3Kjc2sF2H0WF4oOCcROPws+Dp4
xo6/ORclhfEzILJl2JZH4UR2WWgb1mJpPUIOuqSapsCl8bUi+X0PMeGZQSuYz4ZCPiqUsFVFAj/s
xrwGgD0CFaS2KdjnGxt3Embix2Ys7N13V836cRmPKEupuVBRXQb/EM4Z5xw82BNYZB6qx6iKlq9C
bLbIW8L51B82JHM6HPQHyqU2NIIlivIFwmlPtJjK8YlvddFPV3cL+h8ARj6OCRIEX/sYYSrJc+a9
zhyfDYO+JMGXCepcZBz3/1ODgr9wmXoBh0nwHW23l+T496WiWJa2w8nHT4S4QjBXU13z0o2TDeyJ
ZUyNCnVCKfe2dSS4dZy4Bf+MphIMSn/TRIhMONdLeB7hqtthKGrY924wW5bxCcBqt/HITQ/jcTCO
pZQfG4dyPsXOi0uk+/XmEVLlTl3DNBRzLKoVtxZdYmaG9gRC8QO4pjqTD29w1HfLUkA5L4uYzDe1
7G6fLSyXXwO6GzKHJW4Iz/mztsQgLfZ64L/z1tkjPKYwMrQGaWQchVgT3SGN1YLI5KfqxHGmOC2g
GWmg/nZE8mzYyXu0Dl/grXo4eo0QN9PjfwPn34Gk+E5aOwExROLFjarkSb4gM2azO5kijnc+rq32
zhPucDsou+mHQ04NfKO33XnK9XGBCGvYokdcxP63YSk+P+4GrF2KnaTiNtTYqsNFZUsJA5BxvOl8
/Zv8cdxDlTWzyr4ObfeBFn1FNODsd9cgA5ItuIPjjrpg3Qyf9rx0Z3FOVPzYlJId7ERop8Dfg8x2
nlp7+kbAXxnpafYdpAVLy733x2RvE2rwydFVJ0pJaoO8cC9ezH0AAMllgLWEhRXXPeQV4pxwT4ab
hgzf1+x0w7ONi3tFwltNbNw/MezoGce59dVH/xiQt6i681W9BoJx9rVhe6aD9LXu3rW3HTYi3aqY
LzkVWpjNE8y5RjvVvs55Hd8sSqxAzu/DBr5pvpSHlhcM8U9M73mAE5mS/bAo8cGSfe+h4JVnjPl7
sI7jKptTUeGENO05tG7ehhTqLyz3hC7uTNdyEas91uQcuYac8QOA6bqbu+9bAYQxqZ/04mVzzFLn
FUUPGAb8VHTyfgGMaJOG7ioY442TYgbA3rJ71PjQKJos7NSfEQ50xnlH8ZZ0Uw7UZIW4tzaVNpJ9
bJ/mgp0K+BHNspsanQUsrCnJNcH75rGrxNVMQWlVWBwlqfBB2WELPU0s8+r7zLdp1sRNxRibmeg7
h30gK8rehzihFfEQ+4WJxWuwRftvo+X9WQ2C9wES94w26P6rhfyEw/u3eg5RbyESwsM7ICmaXBzJ
vsFIgKTxHbXVoXeKajEoBYDhrnjHCDB5HObhaL6ISVOJRkBNQlPAjD4/Sx7NuiyzEju9pPUkZiOC
OgX72vFoLAkjuhMX5gtNBj/DF2dLo7Hxc2NSOD3cm/eO+GBuFqQnxYDaKKwavxRHhC5XfSMoF135
+O/wwn/Ybgiaw8S3XNygDDNH+Pz1joTxuvUFgFb7SeDFkFH5DHu+TlGCap0tctkIUUniw13CIxY/
jjv7mEM5SvKjukMtFEpUlIYKGk2FMRr0H4gluzs4L+nOpjrLiUgvRMqGxgst/WBe54XLOiFZ5YSh
UTsuqNc2N9/WsH/iJWMroJmoEWC0DsOVog+65r6U7rfx/L0SJ66bAcAEE45TTZ9eJt2gk/fjqiQJ
E4Zf2yAt/DYCpPxFaY1gGRFGB1UOcdDZyLPwA8LV8/73xtTbbEZ2yy5bnwkA5UbLGddq6bpE8/ps
3FasTXXnZp7UeFjs2bPdxBvoR+hZarNERW/aXQpLpUQ3wQY2awV76YgN1rQqHBva+LDhRxk+etAY
nukFuDKVqCQF5TrODi06fftrZsDT0Iu8a5SAeNQEC5CZys7lIIfxUGurCF0pZ1Uo2sMdgrnJZMTC
qPXwHZ7oAfrwUJL4rGGLEWnKPNkMBQhK/z1Nt5Dg9peoDAJK1sr8W9suZOvkXJTi+mg4DGbqidhN
rXKXfWgHjQtn04eNrNCu8sSPBKCEk4sLhYpVgScAaDj309oYmFuqMhKn/uJ2VHCn3O8spMWCXz2T
xGGk1ovdXpsJ5FloVYXfJsw8/fnIU8P3gTRcIpxExNRA5X2WT+OUVBiW1G4Du4jgFHsKlNJgFGvZ
XKAMsbs2Y8Zqtm4DO4A24iChCAqTm3drtpPYltB+X2mt6TwDule45I/2NjoqEij/S5EWXS85npUg
eAWTXAd7U7jR4QP6LV0lAGmihziIKXkjFi1SntaLXWTvuvyMJVQvkzDnnW/jNRbPUAFusUxnHfyo
mfgL5BgOr3WpPink07I0Gl/HI8rng7KMTywuaOgEEXaC93FcHIMm9i8RaXnmh5zWtKmufnmNphzl
ukZBMEIrPeHDXxFr9CNTT7YzZ4Vd3mWLzMXnYHAzAZAKKLiOFCYDH2x8Jhmj0L+mQybTwOjZbTXz
kcl8wR7FiQ4nacf8ls2ygELMgiSxIAMZcItvx453trR0AZiAKegVdWRJsu2nRnkwzZn3cK1AUxQ4
rA4T9fspAao217RurnUGbO7QU/Axqbzr3XNqjEZ93IkyEhonKSOjPvF6FeCW3kZakb+g1KTVYj7s
FN84K3LQZHv8k/UOq8C4TpGFgB329xbHOgUBgVMyvSEq0szqd0ypQTGtVMqVR0okKCYPYvWDQAB8
zIPUVM6hRQf/8Arq6h1VIhnce9U4b8djIcjck5bTJzkL7f1gzqctnkEqFC6a3+hNhplN7Rvwt1fB
4HdF9L1LLtpOWELlM27N02ufNrYhPCUV85W3MUYYIONgBXN08X/A8mNnvtFOoU1u4ierX5lyXZCS
Ekz43jy17izTzZmOz0oMmIDuMNhydWIAiBx0ajkvJ99fvNh+X/kEMBKcWZulTJLWjdV7jEZAHbb5
eC/Rmzi4qipBEPjqJhePwwvFlSwdTdIZHKcoMT321UgruLcTWlpWLWXllELa4iHMsCmYWcd4/2Uv
tECtcODANu/T4t8mz7T0RjEWOndo0pFmAoW2UMyWrl5qeJIa6Sqt9sBn4V9qZm7KlOw6l1VXsqVm
imjAZmvRUdZOWbQt+0o0YF+9AXLyInlfCQwW/J0Z9qbwzcc7dyWhkE949QDqaobQz+nMfYt3E7Dv
5pnyiXekXE5jwxgVfnR4kB3fHYeM1WTpBJhfBsWR2ZbtibOPxnmoDQZ8T4TxNbZNSlqqOiSxQVXw
V0L74TUzGKmnwx0RkCxyqE3XjypGPe9qS0Na7wYumRoa7K56WeM9RqLqy41HYdL9WAgMh17hNsUu
MucMKYvz/eKcVkvZJTFL9RTIp3jmE2mQiUM5u8GTv55d4FGlM7I99wc7eHL4oxDkDviS20aPfx4X
v69ZeFYRj9eILy66FTOGSAqQ7c+KmvQrOJE3wKiwIpMruUTatJ76adzeVXXIi9cob6nbdBgBXmF+
dL6uuAnmvG488fdix8axq1cnWjoM0Wwg4ta4NoXO/rVLr08IJL/fvjqwQfuXQ3t+lbs6CsFXmSr5
Kco9iA/lgN390HHofTnjym1mpIgPHbIhtGKff0Tp1vtEsmVMqajh6mKKMhDNhG4btWuP5LXZKp7z
wewsLo2/j56gHu2xUbM2Gasg4+n9SgZWYGv3JCKcv0ZvTdmlA1xTXi0g8dPMYRjveIVr0lescz+6
GHxVGUQ9u0QtlExSADbqLmo9zA3/n84Y3fI80lID+FmQQR+BjguTYfx2irK6U4j4klwn7TlgpsmT
xMjeqKE0NhDoH+jTkH3RvXDHXeu1tjGePqurMNkjzmZkqLm259+Fh5awW3rwygXzZauYcn6s3eOo
zriBgosmXiat5cf6cdiDsNjmzsGV2dneVW8wv1ns1zPXO20KA1UPk+/cUs2v5e+9F6X398qZE1Af
8Qacg1e58VSEVvZzLe1JQvI/J2OfAdvZWd4mMaw/ejEZxALJq9Ce8Ilx53r1qm/wnvSAypLOuPP5
q/QtDFEaUkOkrZz1//gRzXEdEluEs15YMuvz/Ti+HYPCbKkDwUfvrWVWVWJTFAyq5UzCXlCNqpWa
PtCGUoMG4bH37R0Kd4pyP9F837nTNFzr6UeyC5xARtDSEaVb5XQbokRBbhX8gaFXv7zdYFxblFD9
HELkJ1LsRb6Rt2JeLtnzePmzoa23HCaAKBkNY36Uqj0Ialq3tyyJ7221+GWq63txjjKkDXD2curB
H3ooru9z06xKvDEV9TgmSd97aQavRcNicASs7XJAOjVg3q6LEP6tGHSeYMd70EL6Jk/SktjEI/cF
XAB5KWiQRCHJPfTrBNao5d5DS4AP59bJVyt0E7eL2Mom+w0/mxFtoefgi7G5HoG3qeQh7Xx9DUWe
LSEazWuCtaV0r+SpfOyqiDCQaPtjl0w5pTJuyMrk58Brr4hDlIhityJXiWwrxWFBWUBlLb5ONDQu
cK6GHomM0UK36/Bm/L2g1V/8EXnB6S/8nQHpVZEv0Z2OkV1ga8hk88ENxZ2/gS+uyLNqlw+39dzJ
PDeeSfXOZ4TRakfuWYoN/vPP2EUaoLfbU3Cjl/rwTzfOMXVkZGVo/tR+SZEdKJkbXoaJdNw5rEUM
NTttQmtPrLJXpG1LJJECllWrpnV3OvAyiVJF38+LRowKOh9p3UCEd0pteWfcD61HDCv+DdwkCMax
fJ5P2FQOSKiEIakYvjnIAnBbK5oP4c02Hm8arDDZY/jln9kaf1GYILG8YrrcAtG2ps7yqOD6CB4K
EYK8zz4kYZ7zaOhluSxSGMWF24IjnPUUCjhgn3fwqIK/W/tvyyzPyLaPzj8dWyY7cXXyOW+UGoVM
GIHMXXDGfBd3Q742RRMFH3OCG1iU4SdvE4qNwkNk+/u4E5brUydUASyKuExgbVc5bTbA8ILrSy77
zXRC1u705XbgCD6tiMON8Oxbe0d4DqEN/VNLBDpq41IWeFbw1Na9JYseZwubL2sI6QYEphvm8hua
PCEtnnm5/LzDfRi7uIb4mmkeHvA/cZvvWHkDY6RtUnfwEUPLE1C3w6dqdZkCJon+t+rJyhAcC4Ez
pOcR/J9KBhIPYLQEr3Yl9KhMWkoqAJMZidtN4MXoYK7P2z382pPSX1CzF11dmDiGtchNbJOhqYZn
CivbnjYd0VCRIyM7Z3zKm38xsnLoBKgotV/kOERn8wp8FeinfFrJSpU6azTDpUPQIPM0sVXJzf6x
Yb4nBvbrcS77tBPfd2jjnAEwB5ZpFjYuAM12gro+JZTeL0sjUQSDGsSi1Pz/anO5tItVzoANiTI6
ym1djhg/UOsN5gEicJd9vPASWUVEKMrzgftPmYq9jQWNkNK6+W3Mrh/8l55iJBlRz9O0ycXqpdla
qPoyyPp4dAcNiqJU/0es9yE9K0bdp2oGLWH+G9OzJboyitOe5Vee18kEmpaAf+tCNy1LhA8Xk4JU
eodnpF5q4WlTjApG5IicZI+JYjZfBCx//ebe77XmvTQJMlWc9sJaTjRpG2QrOLjCUhX/gcdfkphS
4ZGuFWDJN7lAgGI0XF8u1t3TbsizXtNx5sHC1qnClZScfbMeuRtxMfxZTLuTjzbNbu+X93ni6TdQ
EwVmLRTrV4lRbsKcn4xeQzC36RpDv1KFco9/z1L4htmVv0TUplGe4atgZqucpgwqrmE0MsutJeJJ
pLfHpbxgQWWnWtaZXHgtjIqax6LHB/wxKnYiJHny81hFsW69PL+N/WiAgWN22H+bKIPeXoh54gap
umlo6biIOZ18Fib0GJQf+bweDyHkdu5SSTZHC8u3HM1pu9Atbmy9nDj9figScJyowB6WwSgwyyFp
T1fSh6D3gR4aQHx7ACXtVxkBAxADjd0jhmyMGDPW2f4WqpYKdDVNTeUZGPCI+IvtPTNQIomcy2sx
Ge41znwu91O5vPxVEedBKaTjNFp0eGWrRSH2gRWis7+GdXRORRxIHZtRcv4YnagL/ClAPlR/i1oo
FrXMM5y3VGSB7LCVt/hKrOx62DSQ43Mk1gh9QRnCigbNywoJvOgtSnBOBAbbNLAcU2DzNrMG71yA
TTEvZ9Mm94jTeAp2v/0UT4XcIdji8FOHIG7S1PsFv+6j3zfrJiJMW5ht/F3zIUtNTUkCTkuLZifN
Yb+ijpCXoazYET3+Cars0ZM0ekr+NbMia1eRq1Nfs34TlEhfaUvESwrezRogCxZyKc6hIjdP4thS
y5WJVM3xqQSfmzSHsOakoC7VxfadFqLtgEgUAs6hyThzoEnTn1Xcz0K7o9pU8MAGn1uQksY3UGQb
UBM0djFt3gkeZxDdtXUJKewGaC3rS/zICOjB0vwJVek4bYzPvsdLLn2jkS+OPTB0FIZydxrfa+n8
OXmyZKvQB4GWH8B4YIk7fY9qBUCMyGGyDkQpIRaFD5EjcT1XwkZ+at8GJEhmxqdVJLQCOjR1Cs0e
8zHpNzc4/Dc4qUbax44xJUrom2r3pgX+uYcGyUkdgvJN5chb3bofD1783dtjOVrzjfRyS9RPbxHS
jdgoDk7Kc5pgJFBfXIpi9/zvu3M1/Q5+xzUv1Exd05Q7Ns7DxBmBuozerX91Git7kB7HHTehCbxy
TJkBT3qs0rabpPII6LNN3VVMnVcokxrFbKwCHWtQA+U+5hMYEx6r0kCzuQfY76ST5EWX5LryXrow
Vp5SkS7tAmqYXA6aoFC8xhI2jXY7pFl6F8jrMTe94hlRh8PbLWDdwhMnRHQQJorTBtzwRHeyF7Bh
O8dy3PAI0dr/xPjTAHHnJ6y6gr24iAZs6cTeAnyPbiLmJLfGtfVijX45bdyKoldtHA4aBnpZBAbz
h4Xcjou3xqgvlQgvs4g//Hi9H77PJCJKdmVqyfZpUTSKAaMX9EntaQoVhhdxitFxs6sxB6xsIDJP
T531ocuciFhdNCBWzCJbXG2zg/CIE6SRVOwGNN5xOijBtqoozrIJFfltyqMiwtFeF8S8Gn5VLO9a
WQxfTaW0RQ1FywjmPrU/vYrwHmicY0IW/vGXnrpFDSqGEXQMMIr6Ex46nDMxZIPdd+Jj4smUQn6k
bzb8a5HaTwLHp45RbFTFKnVRt8WNkkUZwQAlswJCqYxZcnvWQ0/wVOQfQEFdtBnPeM4vLhkv4lt4
sdvcS9amhJICRUMa049AetEhIiEvVslKl6lHfjyGfxzWAiSGE2O9sgMuzSinYyHjfIMj9T3phIBy
nLMWsZi5S5lnii/89qHCNcwTA3RwIw+HtTFE6zG4NcaPRtgq0Y+tZNLo120QVQVnl1jGDLjbTWDg
aKhveNXwZ6wndfwTyS8MxCxM2JZD3FzbIErqMdm2FQCW6eykzDzPBmv0zoQaq6FAcWy8uRNfAo2t
cCDlhWVZ+Fa8yrjoLPuiJe/R2Kf6Y8GZj5eSxvaC7m4MAXItC6RS8e+vqpHRKfNiLj6FU6ct7es1
QTMCbGANFzNxlDNo0iIpUsa7Je2N4qyx7pFO3FRHXh/jpgudkg2XIBAahOI0MksT5fdjeg20lHfH
lED95R7GXgN01XXW2b47SBEefNb7OVJ5Fevyx6DIjjwu9VZQa+h/HEZ+W11BEysadELftGicT5GS
XZ+a5Zwuw9MUd9kWs0aK/4XEUfoVqvacobfftY/saZhO5to27yLPISuwvx5Rf0iHKD11vWMdU4GU
ghrFmXHE9NWASWZVQYdi8jLq4b4/d5chiyCMd7HU4MTAJ00S3Xw/Ep1O4OgRFzQ0HjrIGSYAvtbT
6gtt7dpg94K83xOxdCY2UL7FU+blc/+I1TgjaGQEZ9lficNRohqAzI/M1oij/R78UptR6GAoNkec
V0LrjIPftCKi8tY/xZ4XNE34Jwxq+dAme73PvXp8ljXDTbzj7rf2ymt4WX1oRO+smbMyL//1QqC6
0Wc0UtSaOmarINy80/SsKFaOd4nGQqwXMnLz4+3ioUiVEzilugxLjT1jihkqODJ0tIzOTEdxWp1t
E/LCzqaiMmjyQAF88yiHbJrMu6TkatYosTbFOHAVUQ3Iri4rf5zlyDZbz2f21ZK6FPgBI8/1Xs0t
mUAp4LKCTQa8xTnEYOu/DToL9DgycHGpLB2bZFIhZFokuxuSNwTGD/oHAvNf6t1qbocOMDU6Kjz6
rsGmJvAZtGoYLD0tOOPcAY7ON55Fc3VO+EGHCFOCyLvSWN7WnMgDPEzXO670UVP+LwOf0YHmgKQW
GJ4ukXj0/9UE4zhIifZtrWMWPkiSxnxXu7C1SXjd5hsP4z5Hul2vDYxuVJhWC/dy76OLSEI8jBsG
+bonRX0+jsNOJzp1wjbziC72a3hCeuEA9YesH5W9T4Y+bqNPM0fq0gsz20KQTuHUGWBqINC5v0+I
qQuiT8qPkibntbqtllYiz0JfkALou/eLOY/7uqngSFZ2RmmkHaqzqyYA3s8cnG7sdRx8yBu8F4/v
N513zhIX/v4Jnx4ozQ0gBXUe72IGCHS22pEEmiX7wQL6ahFoooyduDAu9sZvJsaqIIxe5PUK6Iil
/bRDxoPizPc+S+CTxtw7Ihmzq4d1MyZj/HHOEoJ8YsqKqoqrAC1KYBErKpKbxKyXMnG5QYEYdHOs
CWg1PnAqRJBLLC5Cs3adHPdDo80HQiK6GFc1XMxvY4HAAegXQX23nfsGoQCCktOq9anLHT2t1sGM
4ifV/zyn/gnWqSp6hPh91zcRur5fVaKAFob5cHdfPaO+E+2tsWfK0p8THXJlOv4FIWndmATrSh4N
JvcNzLXE29NcC1HcdD6d98Cz8z5c5RvsjGg5fnJTeS4DZRXhM78ogDP6cIzEsacAHA7+5RU72Kd4
OMx3pkTPUytwmb884Hybr6DYLJc66aezLbloPjjWjcwOS/iPl3tNjn+/w70ZD/Go2fnjueX4N3N+
kNAarLFIXvhL7G2WPa1Ri1h/rBAYLWWsRC1iDuanb7u0W5WG4jBdMbQXD1kQucyDrxcGkcGAqNVW
ZTcjFjvvj8CASV9GnrrtXJb/wTM4iATJTRO5fwrQH6G9/J8heTiQHonYBBhZ++gijmtZGwuAgjPt
MCIuH4uM7lZeyKTS04f71WPBe9ryTekXARzTh5SUNbPqI+OQV7YCXb+L4aA2/gvA+ARlNTW6rI8B
xquUlPfRhSvLaOcU0I2QEauhSqTjjjh6izn83nkUYRsDTFsEhz+ZCTfyx8Ui0BSqX0qOp81FynXg
buBfIYb5aiYC/BCk96iyQovCAMlpvDfnrfCAb29qh9KTeEjxQUWvlU4uVn38Yj3KtxFwZ5ZRZWnV
jQNUhY1GEmhQIvKUXzWH4OHuAxHxVeTP3nHVU6fU6ae/L8pgIQXpRCIvmbdjoZDWk2pMe9QhDUwP
cRv1YTjJBKNn+1Y+GR2E+sk2UHz0cnx7OpUVMe//fx1PL2UWhpgBhBCiJZXCGrbRmI42T1p846l0
zIfg0kGhjdSIeKrE4weSxfSPt6tVwqbnCyVLmAJ+PBBzdYaO3wFLIPqR8cvH+/+n+apu0bDrtzeW
UhUFJ7ufoiYfOGeCKOeD84xi1vBPfT0zmacPFEQVx03G/jL4er7XYxHtIJCbmYPPqx676wzkriYf
SLJgboREmzE4l3K003rLBIU4zQlKoj+E8oBjwKY/vtuRXfPGjCEGRHK1B4F33IilBKbFnrojSi3K
lSgNsW52D+wK91e2YjattX7u7f0OZ1s5mk8GsBetB+I73lWQNpPaL4U+715FrUsBEjymy4//MycW
OpPA8njFOEINkb0rZaS9k2Wt7tT3B+MuNo8BS0kDdC1gsar6putimvwjhXUQAO/8wfaqzXSaGtGK
WHk4u2kG0UBdjkWXT2ddynYaI2qkwrFzbZcWL3QbQXPS0ZRPIT55ic8Cj3Y8kJR0NdbVLfxmDZL/
Wn//EeZCfgMQJsMieQXvgWZyGVQcFLIJ2DAKNIAhmn+BrB5EU1sG4O1xNVsOPXv1LUWM2JuY9mVv
pwy2eHUR9wSoSZSOiYAGbpRcCsGze+o1w75KxZRNYTKEKnGOH3BbcqCV91Qu9i/GdNmKo8KhXc4x
XftSZnrPbQTYd6xUJgiEO4oD4BKrE05w3tSIMDXCEVXGHogRQXSPS4mCKz9MBBYZCIugzSXCKYIr
Ey0vFY4U8MG3Ac90YyozTDaIZgDidINdzq8ZMYqlQTLEXjSjJ93BiKoJahNiAMrk85kMyDQm+TX2
967At7eMUnD0TP+5CEZ6/PaezVx1aqimsQVNOJotYmGR0mr9Gm9e9+nToR4vPdYTJeSfwGXieZfh
ac0rVyyEJ7OR30pLH2yZm0JjYUeiiPSUI1tKn3EcSg8JUJOpl7N3HZ1WvEAoNnCpBOPvMT65uwg8
ijbihP3VXtT4AsNHo0vNwbEhiznO8FabW+rdfYW9/Ye44smiCKFVuipWkoCOXrtUYu53yhg3c4vQ
+97uN+B3YvExB5fxHZRyGdvvxw972Y83q570KyebclTWxl0drg8hZFGWhnwoOjX9h08SuKZwcrMN
BipHVKbuLpIIbs6JlTZNNxxkdmoYvZmpg0QdDZo/uc041Lsw06kX9dsgDyCN+4ZlVyQTcj8ui5Te
vdOFvMlYvXyxh2oJU2ayqdqECXgGXCgVdTslTOVDr3idCXGaGVEyesYM9PBgI/kiRav8ETXAmQyX
MyhUBXKODqhye4UmAJwP1gssz6wON0xh/F27kTcnQLLaeg8adR/LNM4oDVfALYQ7KUowd7MR4hiX
/3HxNVxav1NqKqj+AOe0448rL5rjLcxgDCsNDhy4CHVLKFFxrTXPtG8aQllETLfPSZr8dnzh0o+a
75Vc1lknIlI9PLqC++K4LmPntJfXdjfHoGFeTad+gsexeR9Q7oP2ei0ubvenyEs+Icz3NHUXcoxx
njwbVBnwQK4cFgiEm0Q19XOVDzFgd6W8tvuwOa4RaQMUJVcN8jJBKl0828WaFHIT1VsjP0gg0ucv
W3H92G09JRqTemEfFs9SoHjq7PYMfEzUL/w4FuflXejB0oBVimctbzo1bwZ0NihB0ZF/yevIxRTZ
gR7mItDgc2cU8MsI9wOLI9wthggoo/lu/DyjuCSgSHnXsrLrBELPV5HrXlYoqUc2Fxpp9JVHQsLk
1zGHzg88Sy0OGkoEPaCBFIAn0rWOr+SouLEDt0OxsOQ49pzPhrF3jd0CFgtRNEx1SxROxH97PABn
WQ5oU9nrOWyIBAH6LdtVIxRyR6D1kA6bJiVPpevHLXR69E9lGQi+OfCmknZjh9MkwYWTXvJyLE7o
rnknpa19iDidiCzTYTdY9JMAVTomUPCU0pp37rPDA5V/xd2fr9M9iDZ32FQ9yBw6ZQgh0QI8BoN0
6iE5Zo0PWqNlDnow24iBtE+/BppNXU1oHOIgsbPhzFUiwEHJsZbNFKqwWqyZFOx74bDW9W/fqzdP
crNtjGDGsKCi6TjzZb4kVlXvXl02tgGQB8QdwUUayRbMj6Vl0Z6ZZlcjwwvJuhfWcCN6YHt5Wu7F
lUqVCBO4ZrtO4B37/j1qBESGQMazB0Fqu4OlQ8w1m1H6amfDmxjAijenp0Ph8s7vM6L0rT+n5/dW
Ysa1Vrv+EQ2Vwium+86WDmCUZWW+qkWOO/Z8410FMiwvnemNXkwC/BEGu6KWjrpKwl5smuCeTw6G
AfZto02WkI6sjPQAud0Hn0UTZ4klAeuVCQJNqttOYy6UCXTcTBGJIbe0QNgaFXRbk1tDJU/6QSaB
Z54eejBAOksvOH8w8Tr5b2kTHwVICsEHAYwiZjZSL+0Xl10Op+CZEdZA3ZuoTU1QYEsaKyBSXxNM
3Z4PmYMz2GLdtKg3YL7PpvGrBO9RHIqiBVoyzkj76BzROaovg1BmsGLZrFgNcgVuyCRk2AYJ18vP
n766bFUoBxGfvGs1dEmQ9DNiLdfoE4Pq/USfslXwFV/sZfYhp7kF5NaONC3tKXMbvDSXVcou7Qts
PYlaCkd/oXdkOgnyGX5SpYXKsNcg1CNkDGMRENtg5SLkIex8nwKr0CD/nw7pGeStXKQnzSMakSAe
guQj+0KYaXWJ1eq2i5iYtoYEuxrxPQAbyVhM0RBJGfnCQl77es6OWJ0fXzx4s0abo0X3/7B2HVbi
9ZcjyLNmNuZqm2DtBHjzj1wl0GdAVVUyy5Rqe4XxXgSq/nsrGeyaeTxaByTmPbJtQ0ZENyLrOb/H
+Z71NGyIJVkxjGDHj7yrFR1jDJIWG8mgTKFXHQEBgwHnWaEJf7jVEvP9/JdGCBtzBkP3h4/QKQAt
eVf0QkhSvbb3XxvP4f4PBqLNN7kRLswyoVXjnoLm6wyc9VI7P7A+dja9SVvNWb5VsYTYrkGa7Zy9
7lFx7RmNI08zeY5SBm9l9jEzjXe6rc+fL2Enaaj1ZHECEDweFOoVYBmm87rKmTNpgnzgnxxJmOaX
BYKc4+7amnpnTwaO7f+cKIyZiOdcZFgAWZRr+oQl543PmM/B0jyZ4vtll6zBb9nLNtJYwcK3aG1c
zEXRP17BA+oYNV9sAVQKqULpnZHpQbqnPm+7nupj+4GARHFcrmbsBCprWC+76HXssziTQ2djm6Et
83Ln4xfJ5HGzPBJ7fBRqPvs14JpjtAto3ISetthawJM5NSDHFztZgGu4L5aU1+OK0NIU8doAjKss
6z2M1MW5Hcks3yJpMyXiSyddja8kdmCIchGC3Bp+RD+ui5h5U9kQX/zZXH6rCRkNao/C9adQkFqY
+dkjj+gHx9G5uI30+78sMCaC5lCtjcp5AxpffJe6kkihnZcXKKahdtAIvfVTqe959Nl7RqKKB68Y
nS0/Bv2Lvgo+7oe1LhLS/KUkhJoD67XFqE/nWO73uEVTlbKjxDfo6ejsEA/LHdosSbOe6gbGLUIM
Szgmgijiz1DVtSas1joMTC/+1HyOrmrpp8Qfe2E+LWEbAG0M08XezA0fTs1OW2xDY0D6jG/4xaSt
X+LjiEk/da2OOWc3nX4pLzB6h85teNMt/cXEWPTw/p0lu5Cv7J9znTvk0ONW0fxkWvJixblzcnx6
PplEFa5NrR3BbbFPe4I9P/KEp/7QAmIO5foNzdw6RrIgT4NPraXOl7Uq6plmwqTwTo+qgIc9EIE2
77js8z7HZ6Y0xpZP5TH3SadHnPx7Pzg09yx96Ntnm36Qu+w0/xZifIU0BDnC2z1TfKzd1xGzr2oD
dHALItX43d7vLRARI10qIuuCffBZOcZtX8r5F1Owb2o0t3eefeXIC9qKlc1Hd0MidcFgOxndwla8
BObHZBvwsVRa0IY7WqpFep31HhKoXkd1nJKEOgDySE/5lEMyhw0foUSBhDcvDZYaDRVrdm4TyjEv
O+lJlAFMMFIGjsNAicTQw3vmi/SUgW1IrHUxSyJlIMTzxCL4hno2p6DoTZf8QHKnhbixQJ/LdbXk
gnIA3tE+HS5Hj1ABdQOKkz0j64ffKrT8b6PUxdd1002cSmyyQg1z6pwkkXfbGR3HmxMeLzvDxhDb
Ea3tps54bGhDWWXqswWgIxNYMGx4BgCKg3QjTIPd+68O3HKzx6tdym1WOazofvkBm2gJ22JrDLc5
31axla6vfuGXc0rJ7OCqF7Am884q2cG6Kkej47yXMAsu0gKOwtmI7z2Ddj1aHErsWGNNmpkCxaaT
nA3GEwgFhCatX+cl2klRBIyPkjVBKmqYpvBtOEwaQttJ7Nbz29YcSED8Tqmsbqz0kZTvYUkNZ6/L
CUod+pc7CVhdDOjy6T3WS/zKe6uziTcYXZqSzMylOppQRK2At6RgCJAsWuB+0nIqzcP7D5+WyOYg
i+8fsmRV98Vu3h9KK+yNa9VWK2gIvFjMP8VbTCuLiFREUPEDeHt5TDoDkrbyDT4uN2ui3ZN1UxVX
1tp1O3s3VvoGGn4lFS3FxOSanz7B8ZAdFNzaHh8XpRrtKw6G4w7+Fp5ncR1AGjpOy4t+TtLe4wf0
VDvjqVIJKhcNz2zFaMdY/UM+91ZXaulgr52PmwE8rlKwd8yuD6VCefMGq8VyIdWSj08P6Yd6T5Te
G2AwobDpZR7YVW0iPvwK47wATiW2Q7abcFiLt/irBbCXRF9I5fQJ8MipjoA5qITEAh/OFvReZEBj
r3bWuKqk7I1we/PLcsdZHTapKnwXV1zdaowRics1BJPcumprY+GmYawdVrR1XG5Mj1m3wLnLuMwN
GSjInJXkPRAfBCgmHg/7qBxX/Zi8vTtTtTO8wnTc/BvaftFL2yBBnORNH2c5B+G55kr0t3N0EFmb
BHdauV3sfVpuqgX41BGAKTmRuL0e9qRkmZpRyLlG5ADv3EDO/duCopqxJn6VGV9bhwVbfNQb7VPj
QHJOlqz72eOiGb8IAiLM2RTzw8eHoMTIYNz+B+pnNJ/ZxWaHaMd7ZnGDWReSBt3O3OAPr/HpBn3M
KYHQXk1Fq/Dcl7o4Wuyv5yRlzCRzd6I28aHT3QdgGQeIxOS0d983EuzfqBuEJYAWBzcWzBFYZgT6
d4X+3L6IbFu6rLE/vsqCKZlTnvmvXdr+nmTNvW+f2c6oF9AM5xP6DR5srmdor0UYwzkNe92bMVm/
NKu0hXGTln302Cd45VZ5X41bqFsq/L7uSMHIRg8ob1hMCd5dxxtxrLHwZUq0sRodhpzvk5ccmwcL
xv35IqkNR1s6shstTxkNECN7HRNt5/Dgys2t5WkZf27BU7Hw2vLIS2OY7o0B7vK2zNjlcHmiY92T
PlljJxQQrlPxWxe3og8o7FDRVBMdHvxvvK/GJggvfYj9FWbdR+QPnUvqBUCQ4QgBzDB1Muu4KWnJ
6Yn23hO7AGEJDWhFLdqStEGSr1otGFcNLiztF4+7EyxHisoOOfF+R+YAv7Pq7xctqD/ZccuHXpGG
YhSgiJ69oJ+XiaMyVVPrUjc9tF8d12ModdvxsV3MhcYysgHdXWT3lBKD1NH/+kz8ZDJ++dAt6aFO
Ql8QHDVsi2yK/N7+VvcMjwobeNb7W3g2tFSaTWxOaDn+MtaSWrYEyg0UTjRSGcv1QteuG6jQjFQ0
BWpfT2HUJ4cfzUVNm3wDTJua3v7ItENeRpGDwtjytJta/hbE20VEa9QM/2HshsyJhG19TS0xuXSb
RhH68mt52LZ7/ybWgzfDDLU55FV3RgtAyb7Bvs3BcfHDTXoY3us9yGMMjlWT2FNThnXQzWId0X61
UconWtcvxlRitNIb6NpOV3RBieWGzIJs9L66K2gVR5+RlKkFA9wk/pas5tnp0FAGWcEj7bQwvmA5
tFWW4j8sMeqiNpgNbC83PoClPunfxexA7Lf7+ZUfg2ZgZmIb7Cqksdl8fs7R/HwPXwiwcR2ZHjtj
BytgacQgVF+L7GhPNKI6dlJytPc0OU6ffIZU9spSU/yJkOmAp8WW2zixAGmGgeObhTNWYL9dYBW0
grcKUlGq86C7l+Ms1Nb1B4LllGRBWyXICUO1KCkSAaNksMDDFkTuxOks3ytiVzkOzflidJFQH3NP
PBLwqY0nr1bXbyWVdqGlGl1/nfH04J7rrKkryQWq0TEmSl5BWdbjjSX81kL5JYJ4pcHD69Meif0I
8GwUINz2gq/WSmbVQ7bh0WmI0xWRZuK1+p4WHsS9T16YqqC4qZKImxiKrsH4wIhUafSLpZREVVEy
D9umU0HzT95S0FTSOTWPu1Z3E7QQAXrvbi0nErNyT8UMu5BMDdETms6RPafT8AnB/z8ndY+BhvCD
PrkVYZIhvlwwJ8uPfhhx8FvEBse/2XaLlCR6NxdXGexvtf+LdmgqaPL3BM0t1OKum4jMPLWAHIwP
sJR0ZjchooJ/UZHRTqf3RPygsKgOz8dnodGiuPAh/sXBDBF7q9agFfS4YwnnGgTvY17LrieKL004
Mb3DK1BMJgKDPfCHXB+bZiFeVAj5NJ/weGEGl4gvqRv1kb0mEXlujTif9dd1xeFvymyjClJ9ESnL
D0OycsseEtolYogYst6v9+lx+3s0zVj7u/V1cdpZIeFEHeu4xS/EiIJ3i3hXYuu6tuSGINx6rQC1
c5UueoiyQyS8O1fHd3pwOW2xqUUiOYXQ4pGM8rrXPWQD2Ojf24sx4jw2MxsZEgvl6i8Huk4JuqfA
4rsySU9ISdAoSLzuS405s04iWXKE8DMjeXJxd6DkajxJZHKcqoI7GcnwDKDIwEGNfmp+WzwL1bfQ
sG8m0dasZmZQOGCJRZGX6fLqz/9pGpFoojGFQIpCIl89PkrjB0++z074HFA3l4/j8jd7v9km5YvU
nC25hbKXs9Vo+ZXUQ+LNhUirPi5fMsBNnSoJdTIa4zITEpm+B6Tq6aG0MjnHfxi7md5dMt+Q7uc3
dWlWzpRj79gYjkesUmX96E9pF5XO3ydf5kjDMxnDRsj2BFTqsXT2Wjqz+lNKa9rVjIirEJpUa3r7
IQiuL4+J3o3v9Uleiypyr/9kjSGar0D58WaIrNgME1WEsWHvqRBJvzWDbEq/PQawe7dyWKPJKaeA
qVmO9ZQ6PkFYNHD4OI4Ray3SYIDt9sq9gySwklIQXdGGr+akFeBapXCz99YIB/g5HD+V0VaLg5FM
dg0nUTKRE1qR9HiGDDMaYefvs1jd8wuxkyGNLV576jQj8q/PjZd0sjMtdjaHy1kKqK99U/1eo6Pr
xqNZIaoaqMbcT3YuhLsc0SwkLiJKyH6zA5O86VmBuB+b2oDH/aa6kBB5Iiw9A5rlxm5bDB9f9d+R
Pc8YvRNAvgd+XvYEDKRkMBHZSPLZeuCGZVX5Q8NepLHFWv4RVesLraGKoXDb68K8oLVz/hbIAqQ/
aOL6FFM8SSdglaEXOC/xFveqLU3dH5VMf4aB5EhMhum7jNXsEmabFZgGY6c4HDxOQQHn0/9GiULZ
UyYE3JFbWmeFvyaFLHvO+NjVrTBZB1camhbOZJMVvnfz7oIFLpsJdSRjuvRjBTxjjQ9sb14LOfIJ
vyrn7QGSDjj5SRGBn7t8r+6v2kfYV6An6IrmN5Egk0yTvCiXha+Jit593x+B5e/TopPHIhIJazje
/kmKd86Dqz/Hf92AtZRco+likEAmDaWIK4DdOWIn06air6PNjEmuZ3jg/k7SGRQ7RwfJussIsWyw
m8WlIs2vlP+Ibhu+gCnB9D6M7yIfx2Aj9moVD44YWdg18PtcWldpxwcxLa9VkT+YcRoWskYXfTCw
uWIfbs5s1p+bRJPCY/BPaHQ8NibA7v9S9x6vj9HxTn9TUDQEkXBz7/L5D47eH5oO+XvkLsgns5za
LC2DNlpX4CFrD29ar0Vy+OuadzlJQDE4IL/3gKxCC51O4XaxStTrHqQGMC9n6iiS1qRau35O3hbJ
V6WWqrklt6zZOGWiZnUiIN3WlY+JlTCu335hUCE+GKvhdCClJy8L7GR5O2tABSl81kY4GvAOP5Y8
5XTKZdgEdabdqbLOoAWUgcyQ4aCWLqLxL3UOCRQ/tZLPEBhpEzHFbJhyVJapwnXorqSFknlBrArv
55Rdni1BXqXuQInXVt+H+oppf79/3kHP6LhldSY67pTAWYulxLdutr6AaLhJ/VGsfXv8WhZpz3qo
x1qfyf73C3MdrtIanoZTZct6Rx5gqlgV65eCBMG8BPtum11DbXlZUED5Gy/462tMLLW85JtbHRPf
IdInVlVNFokweWmVmJVDH7UTZyplD2J/r4k7vb+UsDhwwgLxDLuASw/GDFreP/PNFJzdtjc9QaSs
8dstfqsGcXWoDWO5pNn0p2m4ggfI3Xg37wLPKPoOAUsMRH6soMBb3wt+bj8RCGWMTAVUolEMJUvX
D2AuEvDhOlp9b6k+QQXDW3DCZzXRg3JHZUb1Sfiv0hhIIfMTZBt9L6v7ScE4KKcfCQPhqvIKcEuf
rkU8SvYX1fuF0pl01z0lf1yboxuD//X78rh1n9SN1zRJWE3CBwA4R+fFav/d84ds2GdhrY6gunPj
JLkwivqpsAONuIDGRhJHX+IXn+ciD2tGLd4tyAQ/znth9FA7RHvXkCOacF80IVp92p7AB0yQ/0aM
GJDufdZPgv0NwOpKqy9MwocqP+GDIsSigI8E4yeMJ3SllpkNeG+28ti75i+l1QzzeDOiA6DtFi/Q
cD+RVFe1vZo0q5LuboWupGsxHZCFUd5YblRucvtvL4+2xtqaTFn0LspeFqDKmp8qxv5mi8owOdjV
q7CEPzkThadlLKswpms44LXYnCLA630sWDqHOqQVV4LzNMt19CXsDBhYVL+ST3lZD8XPIrxYQmu+
foQP89nQeFzl2ZNIPRJG/E4uDj7LdMOUPLx+E31HTyR3CskktGXBGf12wHtDkfGlzVETKaL75YAq
a1RDfgbX+IiX1E+hOU1nG2kPkMFZNvsFt9KkHQhfXY/FtYga0EjuQjTQmPH0drJXIqf427DbQq4g
/WePVVr8QYrPMzkWJrofGHHrrvRhooTDKGgEO1MbcW91f/bJwXIurjs6D/flRTCxiAAP2pEwmHQA
pD6SDu36T6vH9Nfw2xYzQlCV9y5pyk2Kva8oarp8Rte3CkUQJM803iRuy9Yw7pphTjvXPIc0V722
nDNag2NZe5JCN+H5ImPsABZALiOGgtjb+kUouH2UPVoPu1Bf+3/sc/MlyjoPIIo9Vcq6d47OXQbT
yIyO4qzEm0hy4OYc/noK8YZJjq+FmPjJ+tEKOXmfiS2TNTzATT3r0TOVbNbV3jqzgdPclLL33Kqj
sMIsddH/vHV2I2kDTV8yfdzGPMRszioYUbXIXsQ2v0uSr0iWKjYn1iHOg7//Nt14XcxCoRDWDkEQ
XTcIDLyy9UPGpWLKrGcL+GMhAVLUPznoN3rc4u/AMeW52yvyYcxx0cV5DNmEmcfCgejXoo/NTYXT
ovw/wdE47SldDD0lmHpsBQGWw6QBAaSQ9usl8hsWNGL/xZxD4nqDEtDKQUwVtcZI0jp/h9W/Osfr
AaRlf8rAoNEL7gqd6jw/VQBpG3yvGuypmaZMoyuDZNvHLJNGL/e2nASl+iV0fSqyaH4t2+5aOG8L
csKyi1umqE+/dygeYq5JyKmt59y2V3hCFlZY0cfNWBW5M8EozuQ0riFZoQ+T9GnzBAbNYM7Att4g
UyGPlgdwr9SAp4AJG+dv34ZfIyzMsDujb5bYsjcWa9LsmNpAGPiiguyBYoxOmcdG4pIrt5NQKkvq
k1o5hv7bMx97uOOv5TfVu4s+eaXFAioGI8ASWM3p3MV9I0uZkw0TtYala/avZ1Jh/Cg5DpCwMTBx
MYNNSMEIwPzc5C2GxPvrCFYkv0oK36ExpZpqIakjQFl1d/uTJ5nZupDLDhCDYRfb9OPUmZ6OqxSB
FctHlw4uyoS1+K/9R7L7xldpf2pn0t/l2KCh6eDB1VpgSWG0OxmXwlhSUMgfGVX15/tU1rqRaod4
Xi2fTZvhnwlYzO6pW1B9l1ZzSJlaqCBPhsIHLuRfd70dNvOEeFOdavsN6RGp+fcauL+q4YgPjgVp
h0Y2X/XKzFshwKlw8DmDt7p9GeCJa1KaRkb/1lIZynWdOKdzEKDipFBKf1q8bU8192EIshYQ7zZv
Oz+Q6lBppUdf9M3wQ2qHXawdiXXE95idSdLzuYRl7jOInbyAJ9uSssNe71wpJ85zkxOymyg0tCsc
LbO3pmgBESV1YBHm5eQhKMgkQ4gKj6QqWM2FcigO5xQXMPIdmwuUfxzzCc/vIlYKuTEtRXlgUDLb
BrhORBy4rqTu7E8ZU3S3OllHoe8QEOrskrUBdT6y2ogMhOd9E0FybIg+MCmnUPMzlx47IQrXRZj7
4lLRrUHtMwFcUDN5PUx/hQzMeqBnTcevReZz/rPzeedTe66G0QBKmvKwSMe0dWFRnDxme54/attQ
yCA+K7cA4pyuQiOm6GKFax7KSTQ1MrjaBwJkGEzb8icZNGjWPRTsN3u9+CRwzKp7/Vsp+of8Femr
CNsqhWOAelbFwB/Vjh/sEbncHaqHatrOzQne6uiUPK2lYt/svtc8vgv1BltzhMlk3V2GZm+xXAaL
gnz1cMChka7Rs3v/spLgVeZ9rIEMkrC8sa56jcQqtVihftt3/YLr9SgFFTj9Pyi/50eqhpBP7smg
50VKa01VM0K1mJAWt48rJoAlBg2WKNZoTtysINapA64Q6IRXmRfZt0TJCimqVMp69xBx4vBKrXVV
s3p/itqY8ILVvRWXre7xGD4X1AIXBeQ2PUTPYI5rv/yF6fIhKSASP8pP6nLhvD3L9TdegzjY6a0i
yoLx68T2B93WgLgtN6d/NoHcPn4E5/emGzE3Zw09dnGroyerwvg1MKFD67hJkgXmZoqk7yTYpByX
vKrNv6vEEfqMQWVSCLUjHmq2aR2D4EOOIj4gcimEqruT+JVV8Piu9Su+QoFAYZI6oUiPY0rPdWOz
2Pt+Bm8hr+cWm4L3T/y0Cco7k4BfC+igzbpfBUVNh/TgWTXRfWfBvFXuepebCIVjnsIt94xjBpkk
C+xWnGcSwUVsJc/hCgM4aFF1ZhNqZUFla76NSBlNhzJfMIeqS1ow2d6ThJ0oXX+CEgDBEl7k4iUj
BMTVgDojJVPQvIXQ8jNGDK52u3pd+R8kq+pIgh+HDSdymvO9XEaIAwOLy8gZSJC/6b+kSIk3f/qm
XIaxHAl8EltixHdB/3pZAjOlJXD81+x8cYdf/D+ppRzqaZtOdw3vk793+p9CWaV5chqr8WtwN7Tr
dVY6zs73k9iSy6enREGBrHxHJQkG/gV2Wwf2YaBCyU77Qfvr9DSz5ri2VnerRDiKBBw2JeG4HTJU
n1YmpRL578VM+epOV5125nXDxduGbD3pO3a//p6BoGiW1UpG3K4+N3QSP3wL3K9rJibbfOzE60UY
msbHjzCuZCJmJvn4mzCfL7i5tWioFZqPGAUjQSDhWcdjfQxqiQ59s0Arkow6XsSkL3u0Ix9lGlKw
/Tdx7GaunxAIESK1Kh9Z0B45x5Argw4fqMa6p40QdjLgfko+O3q83tdEEHP1PKvIse/VLbuFb3gC
6Pma0Wto0QmNwgSHJ+XfT/8JT5ACTPbLq1qE+l80Yac/QuJRu4Y6fFpsAORKved6nzrGDbV+dPfk
Zcl0lkgQK8p6UWwrFVOYddfLbwOnWnYIE14XQyW/3v1OAWvBYlqqLGCvjXNbNE/vd+MLCoZbXyHo
v/419zepr4PYEwqzYCcQdEU3s+EXWQxyy/LmyLOnDDIkuwmaHD7BATiVD7co2wFobOG+OlVU0iq+
uE+fl/Nrkj1yLyuucI6eo0lJs9SFma46Lt1e1meoUeynFVtHMSm6cepsgmB1ujoiB9UEQDVvBB89
dDIjrl3RbZ0uc37NnDoKP1/mgRPJFzru1/5jyhmpEfaoQJ9aoyYEmT8gm8ia4jRblXZ4BFdW59sO
9LnO57a/Ft5iTN6xTv65rUCJMsBxusTKbdYwAMkOkseB6i1fTlqD8uHcs/5l0cZXxAzJ4r6B4Euj
cq6P4PFvaydVBPR2YG2kLogZbwdEZZG2WQFua7JZr1R7D7xeacoyYZFqJedGe08fV7vz5lF17ikX
zNOM0ynoEzmpDw/SwBb4cylF4UwdTRJBLuQXyGnQV+WMvzHypWTKvvFg1S23uoqBiEJA1fNab5Ru
Mcq8CGADgrMlBaZOI6GK4nrcJoFS/a/ADS033+NLw72pcAOKaRY+uaV3zadtsrFkJYf6mXCgyzSX
XQONuO1eUXx/oh2o9n9kYfIW3t7vyi33DiBCTWkMYvwH1FHa6W5O+k9n1idWcRmrnYCBRTOkc/1Q
xPv9sDfbiAePXxqHpKmztsD+8JX03ncJQZzS6Nt+2iv2YckOzkRKH8HWCl9lGSAr5bi+TV4yvuUh
KoUPnpP2nGgKKRwwJRLmLHgS/Xs8dcdt+K/3Kjrn99D71eDghxGO3TgsxO9QzuANI5ZiherG50Wl
67tYdfi/IQ1RXZpyYfPzpCX4mQWUKvFR+9gXeIvmLoVQqHP9kszM2PmrNdggZ9c11RQTEpWl7D+z
ScWOC7TpV40o4VIyd4ipmyCj7GOq7OwYklgy2gtclty4h56dkamtlYxYkhwf9daBhIerPtaXn/Qg
vgsjxIHRSldT1hJ4U/VF1YbW7gTdBKzIW6otT1Hgxs0h0cLDXT5cA/l7ltKiHLYtgHBjk8UlyVVd
z0AZMsE7ezz9lw67bCEmH3QWB4FmehTdLIhd/hh0dpXd5JHaBW19ptt3DrvvTQikLdacey3AsX/W
tojKIuXYrweCKvFSLOTmFTq6PNfU3aiI8acVxOOIH0WYVycMlmkFpT8Amd8csKeB5fqLdKI38qR0
Z+w2U+xRifSwdY0mpGktT2zB/CewDLg/QnRaqTSxXzP5Na0+OU4m3g9NQPbNeyyZ8UDzg3QzygL0
2pyGk1wPWEbN2M+Cz4eRWCzRblCFfVTKRTdEan2YjrWC0Z4oo3au1r6bDrn4laww5VRIqOuv+KQr
I7DzlF/3HkOMuo2VWxADJK0SVxX5+EBo52Gs+sXgxzZt4+sYdoY9s1Pve2788nD8yCqpQ/h2koAX
wOcRmwUOsUD3gj/qEk4Mentv+xAI6DR371j/OcLPZuYC8cJUs5FmtQrWIsSghKXCNyGfhw2lZ9Dx
1vTm2gaa0Dc8mwGrqJOhv0DUZzzlz5C5uv0UYuZ8wsR1DYIc4AG3S+ZYnQMBZbNOeNYlPiUHgX9s
wqjysd3Asfd/c9n4WkWZewv/MXzpBKFx1l0imr/QKf7UV3kYoAZaL3WtAlixdiebfJECp864hJtE
lnaJe95PojHzmDeZ3dKBDsA1d2A6T1/wqPOpee2NZpoNfKYEWvIgPU+R6cjiesSDeNQUzpVlbozE
OpInjfQZ6LPP+ApXxadWm/6+/8lvgmS5paBTk7SVuAOkEi9gjwJfZBBB5v3/3WZL1YAAaw3rhq/Y
XC1r5OO+T516/Kp4d1Zk956MEP85q5K058g/16cHFboXXap7TnlgRVuqnoKKhS8R4AJ/7cxqnj9T
cK7HdRvf4vWAzH+rof86SdtGObtHZj8PS2EOE1V8nGQQY/EEPk38hjXeQg4SLxaiIxrXo/uqO9xv
lTpw+CUmOTv7N92nYv19ffQrLXIbiH05USziiAC9MwDPoVA/LHCRwwUqmcB/6uxUc9Htr9nHNjJy
FQqJZsWGP/P+8h5+PzBvuPe41MYnodyY3wNe3/KzMp+7wBkRlwqUY2MMgwqPSMygfFPWhj/vQ9Vd
KYdhglAqNXHbyEt3Fe8GTI3f2IKwlXsspN/fxN0svcatA9o5SRKirFdo8vT9oQtHGLFwYcIL0CcE
Uc8hKwXWghQKIT6IwajmljVsP5J4ihE99I2p3mqDWK3Ry71gi2vwHEgrGRp7DDHb1yBaNUZ+JoZs
QlNwAaaYhDIFX5FKPC1Tl2Cd4YfM1UCAlCVHDEuo63dEhbodd/UC3yjplb11iBBM5suK5aiN/qNd
RW/xVwHtKDBgvbBfYYfdAE0ubvX+THk50w+TZFnTGMqJbWUZoHtDO28uDzT/vL0JKBkV+D2MviOY
mD/rMyLo4VEY+7oppS192njIWFMHPFQ4Vu9wl8D0HZ8nT72F//42nUWghr9zehoIVZIBZRxtdsD9
de2u/fOoskN+MgyLfRwn8mdrT4Kl8dh7OsYjCeE1zaBwgmevmAf/p6yKKoQSmPgD60W6tW05yxHW
QfScc7m2G7fCd7ucjM26Gm08bBUOz3n5hU94V7shHZ4XurHGoizRz1RNJEj4sFk1KsFaGVtcYVHg
H4YtIRmtxgXEr3/qkMR1qjatwYA/JTRy17/PD9FDVaLX4UyPrQVxTjA+HMa35ycsi3P2fNz69Lnj
u/aFw521bM7iyLWck3nIIHsgIwm5MlkomCFr8K+0Pm4AX/qNn3GvUIJFz3ynarE1lG8gRzCJce0l
As1lsTN4no4Y/bcMTMg71eH8snYvs9/Z/Z45FFfQ1aD5k5O77rMh5J5rFBbzqOgItZWhcxKm6ely
vYZJhunha1Gvdbr3UZfspxJ7XeUqJ0BcJh1kF6zNxdOYxPqCYcz5aGsi29EznxXF6QozvRegQFEF
9IKtYFHIVHWUIIl5Z7SpXd8a5phyOAObVlr6t+14SXnidJ8TfXbiNjmebpO2abC24vBBc3gLIqvU
XVxw/+Bde08jZ70rbIc1JZKwT7eVELuHwbWGzPihQQD/Hf6sSvStZiOqPKsN2GEF9/IN6gHqlyEr
s0eQOismvhGRWtKzDUb/EysUdHWqtNZ/l26u99k0vulltQknjI8I8nnz4daDzCfCKWZsdnNnYIPE
ulFhlO7DwtZh1A6j//q+HTKQ2JY/A7D1Agt8T9KUy9Mx3FIE2CutSrsds3CXwzS3oNYg3PA8bEjd
PTqIFVZeu7DTG5aYxuBmw4qv8hb6NvhTAWvoE/s/CJoAY8JPvxk+wKH8blKR0KsMmtBbVyGfGaej
GDWNTzlBN0U6cUmW0ZpvDUa0Du3kz6MU6bshR2KO4Mbz0wur0ypZeXy5b6Rtsyq99d63ow4ejPAF
mrd+ToEqwGDoXrIKgsrwtow1pv7MHWccLQkMinjnasWWdiduYeUvSLMsQtowkn0CO7FAB5la3TTt
c4q2Pog9t2vV0mf12HNASy/UjGuuLLrSxeFPg+uhYpEjFgCkoNxj3q0DHWRLuy5onS99YVpZ82fb
8k4qOXzicWZqC//551bJDw09c9oFiIRQWEn3MgwANns9sgoNyV6JAAl7LI4vx0Ku90+ywKkuEOCH
TW5OFxIGdfklVIA3yH+QQQtzNS0xhhb6YvJ4ZuL4kvG01Rtd9h3PLs2tj9zURTDgMFTxugXvwoQS
9vg58javro1eN9vBPdMA5WNprLwxCs8+DcvNb2xPoiXedcvLFqUR1FJMpX2geJCWr0tD0HU7RcUD
1FKrFvM0PGCVe3EHdH99o2bYubVzpQoXuensLYHgtWgYw9O7lO+wRliba8lN5sMUv9M2mUHak58U
LRo2/T6eZWMvMCDR6qGDDA7X3s/8SwgjcxEq1vB7SLjmd/Jik2nOgzlCEeYcWNcXwySI8yShjk/S
pSHNHI55xeMw/U2qDhWHYkw+kk6aFsJtp0y3afzGN6qlG74+0KoLXg5uqQp8EwF6w/T7PWOYmr2w
TJoTOeIGA4NsChC6Wa0EIzt/3AK1zCs22HNuvRIiWd0B9l+GqzkzkNQHjlEDs2/aSdcRsE6Wpifx
LNPbWqD/seQ3OmTVSCMSO4pkZ/rx6bGX69xV5srPSQB8VFzTTCQq9s6cFqHISnYvPVH1chzzJgbO
CLQrSxwKhOA6xrz9ZZusOGLV0cvTjgemkXw/jVdjbJneYMb4gflMqJFFaUYL7eBN8asMUoanuhdE
j2wM4IlS0zgNzFzOatL1L0/Jlp09FAIVUHyr/wGDgpOrkHdVGHNIwjpOWQ1ywHZsZpr9gGofWDI7
FQ0bhObpjzty3PRUrQeHOsnggitYjqOYFfkaInlYa34qcVzjX9lcCRPUceX+tj/Rf3l0tu7Q//w7
U63MKKdqI1AIs1hJDUIjEN67g79wNUr+8dOu2yF31k8Njbu7IZIADFcXqdPjldjloRK8r6+daPCp
GM7vaID2rxj8hiCdQQIqKUyjXw/GYV1EE56i6PWilzZ9iMLKKcI7viJGA+y+KLnjFhmVXRSWLjMS
uVmDSBJc2JBHwJVJOPhguje28t20Gdw9khNe01IbxTRfBYAD4dcXHjAu8DpuRP4rrwiD2ElL3bdL
qBGywtxw9nwQPPukUwMUviIEkczOnfA1lu5M4uYqZ0VpohIFmcQtdZLRFUQbe0wFPQ/K5nEoN/tj
Irt0RfCoMbxwoqdNxq3gAurqkzxpbvCWlSWqmbgeixyZB5D+PHox0AFs7hUnL7fop0QL1R0VH1WG
0Z3RF3m3T/itMJ26Ubj8GtGNHMHdRBPjqk5n76HJyOBte7I6+qzNrLKqCf9iQtgg014J9wdNyyMe
PJCe48y3c0viXzQsuAXp9J9b4ZATs8mwxjP3nQvrk9AxV1pP9Ik9mDF5TrEYTV6Pdx3tKToNSnWZ
5ff91roaeSoM/F8YoQ6NgOjKofbvf8n5rgrho5IVuhW2VoBDivcQ5sOTlX/+s1/kymg76L+I5RaZ
D69qLA2nU4h6eSrnBBxnpQEaxwlcJncwBfOGsPtuS61bu5JzL+KN7LWqbCS2xChKuI5BAYgmx5KQ
Kn3vVbCi12oorLlB/DXy45C2R5prpXmgY0t2GOr6aXHx+GcTfcZay56G03wL+D42Eja/WZqcnwDe
cf/XJqWdXwe89f7LnHyG75NSumy3S7ntp6Lq4mnwrH47MHl86dWXd27ZIPlEw/zE9dE7tZBzR6Mq
JDsrScIAw9AjU1IORXJheK/Lj2TG0mZlQG7wHab5LCjurS6NkLkn1boRC8Di524fJ9W7pkF3IX6+
3M8XJRd83bbkNt3NLW9izbTKShnsUY3QGnKTZPa/hQEvHDVogDxlnpVqPhOueDZ3Cpu8Z2uVKauZ
MGnpC5CPuWJqQVRWoL+Q+TG8k6QyMv36Q7VbCxtzMaNm0dY8hUPQTHFsJYbyq6/d821IqKOQCO22
n1XKsH6ohFphLti6XczfGE0A2TJLCq3rBxzTTBThq4hMh0xGKc3HkeNYNJX6tAvdguG8O/LaVvLl
9mbuf+7pSb41vFffzuSC4n9utKPSIqF3APGurzOPt1cjiEqW/LgLmagSI4CRioOPBaLsWZEcIDia
y9RvNW93g6VoWvS0m18UaayMALrwGMQo7/ZmHqGkqogR6IL3HeFU4juZW0P2mfBVsrk/ZgkfLRWk
+4rGfdOa2hCYtj6NhgGZ6wCsyGuXRTUybKcE/cyVZDZO4Q/BF44IOc02mBZVuKtSBXn3owdmds/3
kaCC6W8AKUYR2wxfeKt92TIOUqr15OSlEVG8vJyzAtxZXHujsgGhpduqeqPT4RLtvmCJ0B83ugkk
6Lg+mYPpfRjOudtAGr5D86NMoJ9n5dl2k10TvVZCCMa80qHeb0fX13aen2Nqy9c50+aP1anH7lTU
ddsJ7z6dAJmzSAZpRC1Bgie99/ruZjnHDERgH8EyGWiB5CohPWHNNEYM2GvnXa3yv0YVP0liVPow
xN1qztmGpyT4G8w7IiNjEbmMTHMRxfV+GC99RwWxxbPt3FjGpF2CnfEPmR4op08HpZfJr8wTIw1n
T99+gNfs542lAa/yGwQI+Wx7PPQQ6y5FZFOGEe3bcQ4rZwxjAUkGVInB9h9ZLFXaKutqMIqya9VT
s7uLqonNVPMofvnwdYcik0XDQHyWbGRtZZs0XtO2oUeeR5vC9709tt1yXaSDEqvCirm2rgTIp2ts
PnysFtuFRyOsB1LFuiRNKgTusAjBlpMdNL+TT+1bh/rQnIcBcqu2Aec0GfiDVOBGd7vUoyeeYIro
mBsXCe0p9bLRVtWIdVCoxfOwr6Q1iiaF1lvku5AfjfPlNjXucgH87SPCIkj0xxxYUZ81XZ/OXaRz
Mgx5PJRuxhtIy2zwN8oyuLRTHCGFhdnuDOcVBQX2JM1Z1/bpv0BbA7UBsF+E/X94TP4euKl3unRr
p5xSvVslrBX5U1i0dMvYVXDqhyd/dLXTrV2v2KPLHbnb2nJhQSCLMQYeEoaaOeeUTfve03xV7bf4
O8HU3wkE+qMsXjs5KYRJNqp0Z8ByDqkLzs/Z+DvAJZJE+naaYc5Xy9WVb7tzIaKOzpENcuckqQCd
SGd25HbNl8wMG2hxS/2AU9Af5cUFV85Pq7VLTEHO13t3+ai3Dc22nXjE8FvwLi9GdR2gh6L9cM6K
f5rz8fdFC/wakLSDoYT9/N0qRfVtV+DA0giEygP/CVQ/yOSYYQVzbgxtElQlvEPO0lhVs2KQIrrJ
Qww3KPhv/+z0BE05aXhSyIGjhq2aaSwOPy4P03bZgZIGA/wdiFXNnLISeP2D14Ge9h4XD9m78Vm+
Ea3DtCOGmQxq41h6cC0QCiKvaRYOZhaKfoMST7mD+/IHu0Ft/HaBktugWex0tTzozcwe+A9UvPsP
UtrblZwRzP4BcNShFpzumM62GsFrBIkauA9g5EpZOSBFVrRSi6uKV4x1wj3ZOA1ASwGzzWJN4S/Q
SkdJRAit4HwpwImC1+ZJyRz/g3y1Bi1KEYje2KAClTRHGXWqSeQaM04Hpwod9ElcjHP6tLSOiH1R
em6U6a+aLkBZ9s7MxkoCKob8De16lZA2JhsE5ajnnfTMv+0I4duhZyPECd22KOc6UT0r0w8fHIIx
xQjCsRmlolGskJ6uCv0sUVoPbDwhXxylJkEhjuz49iNfQhUQpw89D1k0DN8DOhANWO+OWhWxuQs2
9ipKa4tqs/1gCsipsanaPYNJT2RC1x0F9GVWaS+NIkDk0c5DXa8zT7y9LOsPsfk4+QxJe7SDXIX2
jt9ZCXf/A7m1UT2n32D0LWxXxl205aP5iFkhk2d2VwFc4CArN3EWInnr67GKPYzFil+Ic1z8GQcf
X3x/1eaXmHKMARdjAE0N5xRXo8e8xXfAIPmth8mUi20hPOV1ohTEuFu7uk74NA9EKKTQZmOWuQoW
kD6FmqeglWX8c57bSKIm7Y1H32T/pTTWcSS2jbN0Td35a2bXK9vKrlE2l4oA33iDNeLByWVGihSo
1GJ7qzdJ4Hm0jpuXllYJfF62Of+kJhPoovVXE7LV59DS1rwEReWjJd3F40LwwViXo9MT3684t1rV
8WXJ3Jq4OmfTvmSo1Cl20FoxmVPkxP6w74VicZwQxc57U15km5Qz2qAg3iaQD/CQ7XkcDHl6ZNoi
7Md+ukKLz4Z+JDbAYrbbYHeyD71LSTSpYvDQ8bwDjeTG/IoNTS/VelaDWa/s9Mis/gPTUv+19por
ekvCnXtS+ApLIDQ8YxOEJvYMoekfbB8luZ7PT5dy6y+ddKhgmU0bZpiyzxdDWdaGKa3Qdl+gDzmw
N5mha5hZ7BmebvKSpOVcRNNBE+CTWS8zkdAWwdY6icAjZMX9yqQyQE6clNSmnLrFjdWzYthdLmYm
RZLNMpzzl3htEnTLnuoaqDQdHlZEEo2CxbnYGLXVJmiC3YALMqEcmmcleg4VDXNnqupdZ0y8b2JW
pv1t7vyD+WDxaQ8Hvqkwjj6YMAKfGEku414E+g39GvTqumYSKCcidrTFTxBcclEZj23tvfdZz1Bg
KO4pkAlZWukPJDypb8xWNrQERBAWaX5JbbgnF5pdJ9FgSjVd/d+kVmeMjorDSgL2oXsWDwkrxYMY
gFYtXpdxOaP5JkzzRFvRdP9S3sld+QVOQpn+PDZwzlvErR6yrESUVq0H4k1ee786BSDAqVBxaMaH
6mTcBF6YIDMu+gVhi0CBkytki4h6W1uK6qC/aRlVuRiHUDrOyM0WflRBlH5NlCzCrusbmrBPhB23
DLOL5m8MHoUrkTEN/3eKXnu6z6UZCD5UV8gkAyxI0vb/ibXcmGynpELEQYUCIAY0aN+PtS+KuPQV
FnrSOlwT06ztrYvLa4ea++TM5wSzpx7Q07tmQaiK8Grc4ZX28Xal7TgTxeWbMRsI1IJkkJlKNR9C
LUIJPyaLfgJupQKLjNkB5fWWUtGF6qMQwQRO+URqw57RCKcTpAXzdA0+378vbw+anTL/OsIu1zvJ
6uI/tx4hV3R0o7zhH4mc8EQbQvvxYTTBrf68grpAbd2t1kO4vZ50h/FQtg3BBzJIRuuF4gInS08P
xTHdkzXZ7CUDbVkmP1GidXLnn+OF9dWxK2dcaiz9LdNJydkg1nxt6hkclYDD9QX2sBmPW/CpPflY
ku56s3DyXOEOoMivhsvciEMFhIPnOEchlt+UU6eloNpiS2FxXf5ddzN/BTOU1SQDx3f5dCwiXz7Y
KaZQEQUezo3AosK6OnAYYr/RZ1wzlizfZo+rFYZAmcCDUSdTyM5+qAS/VKz/4ozl2jRgfhp0l0Xn
v6X7GDgMpdfr6IoTxZPowOmmOU5KvNIaDnIZVHSONQUoA5RyWLypbEmGtvk3EqIpNll5D78G+Zsg
OhpwbZK0gRtAlfx4oKEQ66dirbTJxVzX3YdUu3dDye1XKNFKjj5Na64Nx5gjX/oSsRdKOK+gZ8xD
VG1wqdOBzNY7JtH30WGhlvNnnTI63FfHPlFNRKc/HcV2SrYUWlCjE9sdd+uyUbyrsctAt2FOpmnW
7uc7H2xYfSSJhSv4VCyF1MjUqhuoHHV0A/XZVrz8H+lobgbKZuEt+U4Fwm2Te9ik9iTZUnHNfv3p
SGH05St029/2VCIviWsfCqnXxrssEshogX50WKwMvoQOyqWZySEacRzYjQQ5a84ROFdIG/kfGaHy
GwhYldphEW5y3R1xcFBX8jGkHrFuGOZ559ld3ySqFx5m2/O6VtIwouq7lSE8jAJGzEJ9Udaq/mFN
OU1RVjZuFwd0uViKOfirt21ObbB2tvMhCBPp7vp0ae5vZa1dZykVfN5pd0aHEELwfgCt0EGBA9cU
jBvz5hKFTtiBl0P3xQTDN7YQ3qqpU2sbcHUBKQf+aliW1Oepvt0VBtEJJcSS49wXHUyDM2KJVTob
W2yLlJG8/n9777QI4/GZJc/pz3iHfiatxQDfoxOVeoW1xzBfVb1xwe5xjBuf6lLnj27TDSs0DnqE
69RbeDDE+wQO8XatJRDVy51FdaDvFdENWHYzDp9/vT09JlmdNqa8nKUdXBpzv9JAL4HTPTncwcdF
UvB9zZnTMi6QPv+NZF+SMzuLL46IkALbIEUsUKgFp4MXNEy/Bm4Jmfz0fOtOWyemLmBicA8bLWef
4I9Xmcg6GJ6GTHIKvwadjfd0zyoLGUT9CPGdx47K56if8S3GyDOhh4h37SsvBzV7EHIWWRIVPnj+
+LIcc7YcUAPYVwaQIbkeoEnxbUViPrIY2DbM4OM0051BP6ddI6ZIinbqzePpLpzFgkfZWtDSc75U
ygLs87wo9T+38L3Gzg/Gy0no2/lwSH16JA33SLRoy20Pq40/e7mU8HOciAnpMCIhPeMKbnxC1Exn
uLFbgm74iFQBhtmchzB7bRLFo8D65PBr+cdNDWvrLdgKQvhRbakSg6eBO4La5Oy+Abk0aGcvkGxH
LXNRwy6WfEgQoOJFHx5ixph45fqYqT1hD8PCaCSHMLfHgEkBP7JO9khNvAvxD9lHvBuDO+o2Nccg
C43JtoY2zPCaFaqB0gihyzFJZO2kj/49fWL/4gV4sdMBqqGjTbx15HpqjmsKF+Gid8atjvZ0r3o+
OxWTfGDScf0wTEZI7pAYuPsi74GaXk25+He1ErSP7uKs0feXqCNr36gAAUbi7m36vOlOPBhKhCOM
2qymScJsBTUfc/7TqvDrHhogmc+fjMQC8E/b6ZUC+PCJlGASAzesFHWCz3lXhyrzBrXCZEXbGK+G
uaJwvf0pEEfmuV1d3i17pM8fo7ub+vbsZ2sb5RvYTfqm1Atbs/rxX5cwadPvJczSe0iyTw2nr5xK
m6DS59zyFd14DxxysEoxYzBLU6s7Tl0x1Ooc5wX9w80x3Cxx4/bNa4Dn9RNTWJf9LXGPt+m8iCuP
ynk1c9CyflK4EjEnJmNTcedhva308WEPYBqX/ztpKwMeK+YShIaAtxUBgKDXgCV1LpRmNQ6saz3M
fng27AP+gzVAq/4czcVpddHcJCgp5ls9Nr8xRN274lHz9Wq81SYGe7nDx9+xwqoVpLJk7GD9X6VD
t1UFyU6H8ga3UtqZfdeEJ8QjBXA9cmDRKpa7nxKX7dCdiv+7KXmgU7HFS7LFiyn4LzRJJghC6tNh
qfvvxwe08guGSLrBuy6fa6Ix2E/cLreEwyPxF7FSpaki9PPrztsJw1dPTjo1lhG6Rq4qPSusVPXU
iSWPynv6Xw4w3KcxSH7c4zc+Vlm0MeydTunHiturtfQ6uBtYRPpNQYPEnfJaniKIkEDnunBOGrFj
LARvI0ddWBRLaSTW8b7KKpW8EYInUTTI13fNgZuU2YbJZqSr8sY2vb+oLXj8P7GOnZsBpcwjJZN0
4mEBcIiC5EIDjO07yYBACY/QRlkVYmI4AEMe8ekbFyBC8bdXT0/O+kRtiOOoOCIhbcsyg/pTuq5Z
Uo82SgCVoAwbrcCA5u52iBwCRvRmR4gWme1nsrQ8FCyjEOqWK7Zpn1f/yqUGwkdYZUvPzirHYcm+
LEsYKJkLcR+jtuXJKrMF9tYeFT8ctFILOx8BquMNy9Bgn8xBLS1Zl0G84RjiKK58uyAMT51sdytj
770pZEFSgkXlNYUFNe5QJG3P5eNB2ZRjfJF7HeJ4iJS1PeUl5bLyJITSIeNTGEG4LLlfHYe2wPoF
fmLLLBA/tXzelnO9SS4SnVxTZWcGFUpI5caNDxfhJ62itojIuhv/gIUABBlk3vBHLBMDDuKccQuQ
Xhx3Sh6L6IanjMp77Gb/Yk/UCQ+3STZOweFVgV+JQO4uDPp6v2T1VYFDqu7AsOF7LeGOsV0FVjzC
UwTZQnDebWliJXg5Lv+xEyhsM1QnaramDp2oX90J3K6vYZmf1EDkclYN4EXW4UlB2b38HkoKXv7C
8c9gYoaFCcaqxinhmARK9yKwIwAFS/F+zdsbsD5Gq9kVLjmz39f+0jfkIyXdXrxlCtUyiHCpDScQ
KnAPiyX4l0xXTdXq8qnVQ4URZ6iyVeo2M41talXkjkdU4zqGA5xo3NfLF5jz554o25r7GF7dbIMD
VcRlpHH8mInQowwhHcLl41iSVQuyP9FTngLMVCiHhFG6ATwyZzoljOdL9eGlek7/IjRe8uUyh42j
BTHm7CpmuvPOmGd37hRqWIWORKslK+zDvD5faAHliYT1cw2QE1HQRRqAcwgQEdkTQBR1UhXGSTdY
UkBDX852MN5I+M2eEZ6hS4q7rFpezP8gnu1tnSVm0DMAvC9Toc8vpmVSsD6cL6HCtQeluftH3vDd
m8f9VpRoy1VmICtugfCYEyth655c2w7IxYgk5tcFOMzKYbJ/Q3gTwCINW9QPziBqsQIJhd3XDaRz
JvyYgH5iG9akYZq8kMq4U4cDNAOR7FF2vpGoK+DtwPS109UddNH+scTJoRgLRhQWnO+KXaDvhaKP
wbjpH4RHMBDybxlmqfw4VO4Dn4EfwEgfaVoFyTxnxQl9BUrg/b84sfUqF/WrXcHhHhImQL8Z2i5T
1Nil6Pa7z4IrxkkdZzJkuqnQuRv2/f0688Hh9MN9bTLL8DmaDXJmPsGZMYNExfg9iw4vC4Hai+qj
HVCpI+k7oRWQUGUGaV96dxWK6TsWp4lmFymlJ2+okZwQE0WTAge/CstdspRpRqTnzlp4wIMe8+Ns
rqJoImYWYmLDfBMpXxIENYAYohlMQDamfgNl0xTXnZm3UoonS82EUqOja3STmFbHqWKmoG934vtX
Cogh74lVPJ9pxqH5axxXT6+l7Q4bDoMiBC1d+J3MSjpEqdHONKugeI0ao7w0xgyT5mVQoX2p8rDx
rX5mcEOXGj3JC5z13wAJDX0sNbc+M/Y5jKgZ8FE+zWjOwGPeyLgsnXVi3aYf1TEoLC+I4V4iiVoq
c5rnRF+uGq14tRcgzoVD3qdIWTYTGfXN9FyRhngaJEQuMIwA5iBgEWCtElPvUUZGCfBB1clb4Lpq
uWNK+1eEeLLQm/2pmItBxCDmmlebR7jNI3WN0mpzO77v4GXTGnGl786H5WBlvyuAiDUJ2Jdp4vnS
m4AzlqjGsw8MKwzCxrWMvIngreIPqMb7/MV6NOxNuNo7t95Dx04ydObsrAZO0iGYOHuKsbGyqFX4
2vuINJXtDO688JEteuOcYm+MK97J/V1aKzjCnsUP6IqrVd7sPtFO6HVDOz4tXiHlO5sh1vGhFs3l
uc+/m8jJbSqFQ6odwkqYi+TU11SJvZNd7DZh5k+6FrAPHPoH+Cu/6A7KJnCDouKjtrwxlYVk1780
S2IrelJuFJPDxoAVYZMkfHHiVYDlaUBlQ374tFKhSIrrO0nekWvtXu2V1JNlaXY73D5kvkG57o8X
ECykYxnOOcaPHnjYM/olTxwyhVFQcJ25fAQsZ0ftw1omnf7o7TuRWeXtzY3rigFrTTayzoT7VjkI
o3JJHVdvQkEQDYDxOgSuUbVNUtlt0tJsERYWkC7D4vanlAdCNRj6o93UB2uvqmZboaeoFQgxEV5o
DX0/w86aGcT9C5siehxWyvyJqY0g7xtcJ+BbTGFGK3H2/9azki0AOlBd+jFebIgeYFoafCSnasYc
4aglPefh75gOM+Bl47+IAJUo+grpauLXpqxrZdqDunqYDD4L9QEPNANK+ET0AwQmkkG4kc14os3V
oDnbIdxcJsYvTp60v2oqaR9QqGh6mW0Wg6aQSrh1Wfi7EcFANLn81VP0awZKCuGCuvPmil6VLKvA
E0tMZeupCA0KdE+yZMcDgxBWq2Cm28FnRQ173dbuOZpIFfXiybq8gyuanDqGWXF3G7OE4PA+b7Zp
Gg+iwWc7BAhS9McFkiHnvjwr1KjD5vK9H2tZz/AI52X3Si1t3Vmn2gRgg9Z91a0n8HOfIFGPXSeL
gPJ0MO+4UfDboq1rjhko101O7IWfg8cnK4Vtb28hTHvc0LlGMhEpp/zlKAe86QzC8FtusoNF1ZoC
OFMxT65BOo/mFu2e/z/ux1yW7TaZogBJmOxrI+5129pn6MKuFvbUE9bRSwgAz76/pEWYwbhk0r5G
fZ8YlNkk6hHXbBPr42G42wDfPMLSkaZ4wFNrrlVLUVwkBz/U1YJotzAay8ql0Y8W+BorLRrG0p/w
a8M9724+lUzmIkGwJ09e65GUTM2wbAWeOG0VKGgm78YuxDzZWpdrnPghCqrBHBQukoJ8MyCLtBwr
gK6RgR0b/TytCtniO37ymanLvtkl1BL7jYtdVkI2XmCWsIEcaUjcdwaHJn8Nm4INssUPqK2SmBA8
v3sgKxgARd2bjM/mAeEoFBviEl7ugCVfi0iEGqWgmreFiqNZT93naUltBGUEiupUIUfR5SwiJ1iR
eB0p4jiJbKyAgtkpE5mfasNUGi83vES9M/ZmjGegTXhaOuiNlkh2Fy3v2WML4sy8VmgG/XGkOFEP
HLoQQdoAfVGgAIw7SOcCGtLYOPlztcOUDDbQeYUkRBbAmsdMbi2qCpZJs615jhLD6aWiELbJ7PXi
6VBDzrJnF03T86vwsYjzI+w/Wdlj/c9hp23r2wbINeIgX1Tq2o3GpOTj+Ln39jGio+BazKGt3lbT
vcY79s5IHOoNbt0vfuqSA5MUL+xQoDABAp8/bySomymWlDs7/sv7xf/7lhx8OqDqtGAJ/qVspiJs
Sp/zoA4m1xKmg0fn5GY0jQXLwnBZa2rAB91u8fi+ndjIntlYM85L3RqLil5kSv4WoLoal648bwo2
BXvcB3dNwTsUWkYeirLgYG9eCEKihNFCHRKjEPYQKFCgzU02Cy6m+vcLTECrrQQ58xXi3A38o3lo
Jrrrh/aQz1l2rTe1/4G6WNAaYFSr5Hq69Vk0EnR2eC9IwheMWQo6RtNuBFqnvm5R8eCwVvErHIL+
JcMlULyZF44LMGpAkTdGUHqqVGACEMC/RxjqOwyNMDT23HF4P5EW2MN/g87Xa3QABr30jT+4o4qi
5AXWk8YxcVVpf0cw5mimLkQ3ZvNGtH5SYVLfCawcURmRa/pznHTUM+oe+xWH9KlDbkRDuVrrJJHA
REizOmKPUsIje5lnguw9rLPGoS80u6kRrZM9e0RaxtzazyS77VY2rwuk7zJO15Hn6TfqpRS2OOk/
4PpWz6T70gbhjr3erLP520Qwd4j0Oh+dCVCfQ2NhnkSbNzrfXfAL8OgJ2UVeEC4ZbB6ESxl/LxTd
sDdkSkISJCKV5zvmAZia3aNav5NNtqMgZFq1UrkoCXdKlsByTov15OMmZycoYCVHbwgy0yTKrZ8t
aK3uty51do861ZSaYYdVh6yFsZomt6l3Z+UCldycZiHzzx5Dmoq8nae1wmBKcMviBMurueoAQsl9
paHFXyMJNRrJJf1Wws51U17yERCUFpXrnNplVL0e8CE2io0eBU1fbYt6VSAJJFc/Hpvd+K8u8vBC
nH0AHsIgfpVtSC/2s43ugUenWTyujgz0XboMDse+lcvb1o7v1ahin86NV/0epjFUpVU9RHKJ1T54
VW9ctxmnOCYrwredNgZmHTK/UOlvtM0WRiTqmfeHdiO5gWBMsRtgxDRh8IfLTYdogsRPrPI6lYrN
mi3RUF/kS85IJXYeve9G5FhW3lTWEL+LgRq/tGpyqlyHpTudHg0jztqYbRWQJdJPtuNAfNHYHqQ1
ejV+HX0XsrLNAScwEUbetHuww2xcrYlUn/LENxBExnvPtA6NoA5EkbiqpBkRc7S/tqAX1uamZcxX
eE3uZbh5Lor/cWtYqJRvi39eaaY445uZTHCAxwxCxPP7ZarGlnkG1xKubUHrfBD9GP2mfsngERyp
owIMSLQvdFzXWqHEW/SwO6TqC0fx7vCjJf3L0xPk7PSGKpNeoW4GZ7St7N4xF4ySvCIYlSIZaDmb
uUdHvd82SwBJf4rGjZwrt6FD17mU9JogCgGQn4L0ifVg5HkgbdUODB8gHROufArPz/kqxALKbuav
nSqLbUGXq/D4wWg/YGnpgnXx7OdLOu9cu03jRfHo3YHnLLn9oVL0VclKT6mTW9iIB8k3IhOyAz8/
dKT10CuMk16e6C0/DlGyUlT1NLygjnJ4WD7tw+xd3dZiDeSq20dH14DO9j1LW45h5A+Atmn3eRRw
DdbyTNNdpBZAzeHmNtQtm7tNDIlRoi7UfQ1L/PdEFUVwKFNttdqDFza282zteHvbgKSwk9t3yyH0
jQX0Xek7xlTiZpIGTZ9kQltKhNNweyj12sSHs1cMaz44qyhDAG0eUDxzze/3Gxa3K3f4SkB/iwnI
4KbU1ZWI6NRcGaeFOdq5OTfYcjHlI88eM388qQ25+rZP29cVtPgyUqhzZqjAhYfcphFYI0zNThNb
IC5esDaLdXU4FsoCL1jX5ZANB+31Jz732AEyEMMl5DJCkJhLGcb9n/cqRLgq6YsXR3b+twdMI9oo
X/rwi/28H9UKIFElnEHbMnxnNMDPLK8KxxWWbfRRUoaIVmEmJylXKOzw7QtB78xY25PUNPkOyObW
7TC4WoFFBMSxL6jl8MTnnOwmTzSWQ8qV/GdVbDqIWHChxOxRQo8QFgo30XmEPMNLQZn+ydj+WRVy
CRuebb52MEBhV2C+wRbA+WqoqsCU7b8ZQFIEkU+qbP/AKnbTu6uStvQWLMC9TUo168jL858hIJXj
EnXgPOF11ofyckzs3wF+uOiJ03fB3uu5DwQVdvkcYAq68A1rOHH7Gl0j/Y8yVBW34qL+IAF7hq1s
jN811ZdOHMbM14/nBKk9GWoA2vXKyAr1B7FQTQKb16qzdEJg8694ePVKRPB1n6Z/4UU/vXWdBTV2
cFLprlaO1osStoUULEC6Ngvx7GoE64LB7+Oze/x7ncCHhtP/afYkPPTlMBsmQmJ/oMy6pkdBKD+u
+27zfH3IHevZg5CMGYw9qagqYm11u4wEWxVMBoBQGaRS6i3ZF4MVQJByUvkKKJEToY+tYDPlXr0l
h989Xf/iRfVdj145xMIbkbJMS0UKFru0HTkdqdtClgh6RXyyO4uEsjMaKs2Qd4vrQh1y+O7dBWOo
GbxrhnZfLOkKx74PrNlBmDN65jFiqZ1qRU5WhTMnGqLTOneTQD6paGWOPn9Zj+faF1Ao7xq7BgsU
Fs5ju0TaaFxrsYc+N+l3nfb8F7q04jD0W5lPhxrcRE3xmZe6B2GbL6p+yDU4hJ+rORpxlcZewmqB
qULxW4MS6dtb9PRB66QM5Jci4mCD9kp1+jCdKYiMvDmICOsQ4oj0QgcVyZfiidIOdZKs7fZSBHJA
KTr6sJV2KVx55cQBlNXTVoVeXeXK9YKq87SvWXYEnaSRyg/4c/cCacYOChI7w4tPkQNLJ9Zg5qjN
gJlv7FwbjwElil0NCa+DvBJ1G6dkhUJxtAFOg74QpVyA/jcCfx5hXoHeoP5lPPy6oRMyx6+V5NQC
WADNVZPE0x0cs4XbT8dIH9vtnDqLiXvqXC+xTa35cJV/CNHGEjh8TUoYXbky6lC5pvjI57kZXuho
Gm2PSc2Pzpx/l6Y2gUP1PicfIZVYR5AuBIAcDwfjm3nKTxmh8JWwmUK3jWTyXYEoa7zRhdK49UfH
oYdsHV5+oKLnchbOiZQDj2NrIETlo3oCxJkBrFXAdQgAGHmnfXfNimXFs1oZsaFLLW5FuGkeoRCt
00WPCG2yaQGhwbkoeHCEe/XvkVUibjIxl2rwNtSXkG+Spq6+SW4Qx4NOsFTmHp14Br0KewznCBgv
PlomyqZ1nNqik2JvNskvCMfc7MKUd6NvXf5jKApqmZp3pk7Du4Exv0pg1uNrCfj2cobLUYUFmKQP
j9LXHOgFngGKfx+tbJdK6TqZlfugrYLurO0GQyB7JPF4VEYz+PI9eYr9YnyEIQNSBlyuaHrYfTUF
AbpbukqnWGjjkh3YAnZtoHevNp42C99fJa6z8F67fAf47aconoPYDHy5kbY21ahaBnbRWAvVhi+Z
7FFFRf7XWxL02IPm/D+vYy+GA7Rnz2o2szKjP4Hcr3FDiiByYSNAHzEL3gKN5VdRygKINWPNpj8k
ErBbDTs79gW7lm+lWHanwLRNLWJBh1evGWR8reGWBz1rqwoi00AHeCXdpulaBWoXgKlJ5ggMpIhx
D1xpl7gcumGT/xVqQuti+6sC2tajWd8DNOgFjrcHtVQty/0Awub+Lxjd5ld/69z/YTuu14WLaP77
/lFiP/PtgZ5Oa64rVONZ5crNlB+AY3A1T0CKH/IEPILtAcJrWT7v34KcrIArKNj/LSaaCe6FDBe3
zlwjc7Ekblo+rxyfBbSJK/AIuCYsr20YC2TkmuEXF4s89Hl2cbbQzx5VS1FozviviwX8X2tpddUk
Hs6kKb3L1QH3/aAtxSf+otm9wugAUKJQ+wCnc4arnZRVn9FWEV75PJ3lS2xO54RI/Lm67P5ojlBl
sBtSPzY4W8p8PLCaUspHDFaq6OM7Zw+E8ReNKY5Y0cfws9PSJpCD7WXg0LRp8087AM6avQJ7YYgm
BEwgRNIZvI7lCgpAZdVUTD+vUWuKjqX45iXocxuwb3OKWCPNcgdxcXWOdyByV95KXrGwttSCeEvq
J2q4YXFSk+0qN3tDGpNGaAl/7r4NEqCbcBHaZRpcJH8+lK4JOO3RoPm6OqzWmTz/yEfGpt2wbqr4
6jmv9JiI46CJpLrUDdR1uwOrn7h3PFIWE6WzvjFKCoNjYGDuo36cg/SpCCWtH0OiknEKwbA8K4+S
sCapXNNDbPBTW9rJrnJixZW1xY7vYeueg403YcLCznLwyu17eTHC5IGqDvYEOyRQ53ef5sJtP8C3
blbbiHRCihAwVAQa2p2CW+Q88RUPAYMRLfcRE2i2kleZG4JnmagdDu5X7Tt6otBWaFMCT0f621jJ
e4Ap68C4hS/pMGz/yFM6Bm8U/tzgAiyS+8BY72VYG8ILEwWOzdOCC25NHweO3RGs8u33jKucBzuz
rk5sbD331n51rlKKs7dZdU++++c4RLngtKrkXmlWNigpxe/0KHJsqops3lGTybQFnWg0q8F+nsKs
bVV3/zmcr+WUWjsEPt5U7SQ9sJFke1wAQDovvhppQxhd7QLE5ZtsgiKIBxxTyLA8Y0qvnIjt+4Ym
x6eYX2FarCM1hXChuu5+d5Nds3vqG8s51y5eX8I/mqJhRmNILnUyUrXHPVJ4xOyOfKDPLmfYiGuQ
UwTHopqWaV5Kv3G79161EnxX9XXR4ADJ3imwDDDwemagOH92bsbWZIW/gFNsLpV6PDocKRQ8bBPx
4sWiIyU9e10c0FZrxUu8FrWH2ZMaqoGRIa0J8sq2UUr2db11W9mfkD5t8z6egNNZXwpm7O3jQBJv
Oom6gs9apbWzFnn8sgFidvhPtBISzGsbnqslzJlNLlg9lHUuigFi1s0Tam/SQLOvEbEpyEa0FJ7U
CyeIetjGXKN+cFnfs2r1Oa1m2h7KdUFvZgcZ+Mjc17Ox2nOCNBZe7uNOnFzadDHtFbH1S0Waez1n
NwzYywk/RV9ig4eEuDSUi8doXSccbLn11DaZBmEM/CdwsLhoPrtKCiqJRTk9wGmveBHUmj6qJyG2
SsiHRKn+Yn5dXHpqGEgHnIXKgMNQyfmRtyvUZMj+JzAb2sbHo1YdKNzPj/uwcu8w3Cgbz2fLKz/B
Sf01p4+zI8LLPxS0Nh/WbD2l5+PvXHc7tcg5q9o9nQaHruxci/GJZqoJbudszLUmD+vPLX9nVzfE
Slid9V3CjmXhmIzPlmRuFyu4SCqoMy3wV0vtFA5oKK4gfJf++WhJt1KkdsZy/IqD7SVS24r2N56W
AVl9cj+YrUg+3MAVSv/9MPkHzqUBlzezolghOn7ZALGvVVmzGfVv5EYp228iEE2IR8sYoqx+29Ke
bYz9RYo378FYP0uTWasDdiFhh+i+v056j6kKF5DcnXKQje4FfrpCF0zKNEOLxQUUEChOBTMKXAZh
FTMOFnCCGiQdRQrhNZBPt/IjpAf0h8Qjw9a2FlRujftBYIvL9AL+OWLvgbRusyfCvvplyh7z8MyI
vxIKPMlqjzkFNvwg+RFVfigqKVfZbQXJNjAqOjzqwKww3fw83SOBn/Cq54ldfHSXkKbbQH65OZL9
ajYGBXYb3aU6INq6FNgGu0sHm8N+nPSoFM0q3oKC0xuqk7XK41Ufm3cB1lAeDjjXwutL1qyVPLid
StLi4igt7WUoIwmS7nuN9XmsOeKLzvC/Vpebx4dlBbL3MwPnltlElY42mmd6gYweO54KhFVP71QX
f+OdNw/JL9SldggCjnmBoZyXVPSrFQH2RnAzAtc5KznK/y7umhK3cjZ/awStU7sTYCpkKU6Lxe3x
a1ryLdGGjAu0eYG9MfYA7Ns9tfq0W+9iJYIv/zJpoUt6AT51yC09YJHm4ZDrILL4xDP4GfIpY2YA
pyO8p9ItApJzUTUOqHriDOv6YoFnjfP6cJQwreiQBonwMGZ+FN+rEUo7bP/SA0Jl2uieEpeyak7p
TxdgmnHXeROmuJfMOyEl/Zawb8qC94ZbaT0pPx/XQIo96tJTGkKK14q/8QTAOH9CDX3/Ht/8x2Iq
MrK07Cu2EuGhqKQ00MneLbURJC42zEEsWtE0a/AVv4x/kp1f+Itug4A2PCerVc6z85ABh6uYZY/Z
AeK3qQntFakaRyLYf7EqxVrRhHl+TEKD4GCuZccV4s1G3oFCH44zhZb7fpBivPpes21OaidOBLSQ
sgYCYmB7UpLt56h6SR0yGO78DidFjXNyOHLZRBY1nyUaVYv35uFc1Pbvv6zs+rqiL6lmT+VfVEBu
IhLsR2NA6Bo0X0T9JBrc4pqADeviDghWBLulXDt9zOlXGRyaapJDIKwP4+wEl24Y6D01arCXPbim
kl9JVnyxGK+7qL2iU1D+RI8mY+s7+8PgqUk5lr1dt5KY//SMYf8qpXaDTrHIftV0nwNYu5U5kc+i
ghF6z3FbvsGXX+6SaKpFTS3I7629SdFSplDZS9n6rxf7GJKCLrffxvZ1Wgwq4bxUD/TQABWcV1Vs
igYkg9X5viG2bZni4ZvZkUeWKKuh45QXRox7ljr1O8mOMsO+uqgI7gQEMIM2J5A+eclkT9Y4fEfQ
264d3ViFpCxoMNeBZKQJ9ZsX1DlQHnvgpZJkWRQwpK3RmX4F/R87/R1vV/8RL2SApVqi6y/4vvO/
qSGzlwojCzY59Dx4e5za7vDxiYE9JzcVJPEE4upR7e2rEwgqj+G9A/OZS0YFCisMxXXk0DeP1TP9
TLbtXg45GIC1UyDir0G5Y2u/xVAEDjqsTSGvwFuD0JLVgFKwRPn/tY6L4AidOgliPumMWJqvixEp
O+JluvYe7snbJPUaTof0CnAFKPOIX75WiZE/q9hpyd9ojxU0wD7MhmU5X4hKUB9UT5f2RJSqQni8
07GNnu6h2U6YJn7oZDuyfZGxN9vZatJ5aP5H55d98Hpdp57+xnTiBF6NoOcmLCGCWCVmSUx2YHbk
BVZh/qeMLRSzCKrd4IdwzEXqiDEBIlO6WA0Lvg6R12Fb4bEID3V0F0mmE/CNgcm31RRxkC0awcOY
+HCaqIYD0ToKuPVDNKtQ8OK2YXVmNwVqQ0i4FL9FHNJ77uio55ipfTsSMDaSBVJE69BDPwZJ1plR
6lWIulzEcUklm6s2sRS1DrOFrP08p9wXUm3Nu6uFqQPAcCqsElNQAQElw62JOLv+La/FqX93Ys0Y
gsiUu33hRF6xU1cehQc+QlxzRdqdnRiWYeXq0+3q+BZGniga748Tq+CbEKObk6i7ITePRVJHfCn0
RR9gxSjFxBXE2AfWiCfnN/Xehv594CZ9VYq29UPpWyoT+SEuJ9T7ps9c4GswIOUdQsNaWC/4ZtUl
ez73Y69Ko5DYEoLwKQhrAmCJPsLYtvNUeszwn3R7a+DRHEVDnajFwHwp+8eaXZxCKOohd5ZcSRZ1
n2LdC7BHvweWRI5LgDYBnCkX9oyzQHCKht9MFPWEdnfmScC4NzInQvfS3prODtmjtbex74OCY4dC
Tv/CsATExXROn49Z2sqgVpTmbs7Mg39FjHwREPmMrCTLSJdGdi3yV2zhcWhiIrt509rQZv+tmV2w
oiAcFWPa+fv0eMvcywV5f2jVjxn9Q8Bjk63JlETouf8p7KZnQJ3HQs/+ULx/yy8B4yywXfRRKYlE
TPWEOw34fsVcyfEhWb7ri7oesd53ZBLE5X8j722XzmAXw1wZOCe5d7xYvCPjDXKlMka8yzXhgobA
BnPt4zKlANareKBqGyym3zX8cBvTiJ0SbmYIs3BOsZL08/fEE9ud4rjIua1MM2KD+cnprQQnG99S
17pDzXT5rrOybMs/zQDcglrgqCm4ySylY3GPeZjwrndCHLj7iPUg0iC0CH82H7nmsXQNOQ2y6AQM
g0vGpXC1ewu9x3MTLgAwugQ3DoVGmSxLF0RNo7hT37XtWJZfBw9mFrd1jAsk42xhq6VmGK9B5ZQD
LBf3g/dehKnZnrHk9VFg8K28tC3exXJo+POiFmmlZYcULk1cilqqrDi4tTskH/yKFFfkxOst8vfx
r8sLaP9rxGLbAtsuVHadPm1+GHyAyRXU5iNj9Y1uBn5W3qlvWjFwAEk3AHd/GCNsyMN0gYSmMKvn
0yf5pQQLdMbSUz0jngitA9i1TGNSR8iJxtMHR9f/2xgIjKYFXPidukx6EY/k7PLueNF1hwCBbpTx
+W5g4aLRVPRoxuEyczJsF67J7JmJQ6B3ucUdF3Bfyep0u2Qe50b3kiBzfNsJHboPrnaJcTmV2dVd
MYwETdMg+bGRERV8u9OuS/zIDAuoA9V3Z5Jpgm8B+rvyAGhQlhybwEe6ZL8uLkmuvxafjzOjlqZM
j+lz7cw1yWgGixLskKGeu6U3NSQ48ITMTo1ZWnmFW3lJK64RVadHDJSMG26049JUEPY3Ut2B7oGE
D9O/M/xWHmDKeoIdgRsrWyBtH8bcaP8bA8fDGU22y+h3N8W+gLiBhk7dBwWXx1HbysZldeejEYzP
t//0UR5gzAKXHaycXNt3RSsynXHcpW7lWXj6n3xuRl2xY0flgbzG8RmoWB/ZbZXknvz2l5zyAsKi
MrNlQBHWm4b74h00eDq4laNl1hBA7MDRgfImmsO5D9O1fnV3jpzbtAr/0v2bVdHiyIMSJjkTmHGe
7hdOMxEoRzT8JW5VJ2CfTgw6sZAYLzeaAJ19nJTjsCx14fgDJLEI9VOqvZ2eM+/zxZaQy03V7V77
gWj5aRb9Y4e0uwFdRJupUC/4phwNMf1uWXqYtRW80BSslQaK08bROTKgOgRdRXDaosPb45hvp9Pj
YIlzcwt6bvAKqnUoxQL/GTwRD3tBZQgL7FzBKMbqD7ciYe1q9na0ohy2lPuVK9WVzn2NAc73LnBb
FxkE2dLJut2QNQL7KoKs++Hux8gWRntLOlKlfwPrCCG3HFF7iuiriOk/AlvKpLzFXGxNFRztAmjf
XtbCBFrtzuwCknnB3bgbf4qh/5jhLHzOSkc68uU253k210BlBtwkTuzRdc+6CAxRUN5LS826Hr6l
dXiGdFWLjoqofls1c6opnFoYYp/8fkPW7OaD47ryx5N9vsSJVbOToLf80LaX42vuOYc0I5gcqil9
hEyi4EbttoyWc/wZrvjyOQ6jqX7bD3mAXP65VgJPbrGlvtYmGCkeFBtgyO0g8avyJSNTLovshPKi
yJJq2zadIDnIQCJezkSgTieypEDSoWedI7Q+ylJ8aB5DynkvlpL3nUxhGqVHgcRjHt+zBQM7+jhT
ep11OXQ/7XCETro0aG8DEJpPOCv110i+932cr9nKFn1hKSO0IJYjlP2D7vPpYKXg6hbkICaTOdpl
uV2ii30xoLjqHEVLcxoCqUqV+AU6Udue32RQYAXDJkbmdH0St/kAgS8ORTuS3eObU9bagmyAUuCq
TNboOJkP7zGyAf05QfZOye0PqQygTcHLdCXLO4u69G9iUeLtoPbDPaFL3zkSvRTDem+WsU2Ctz/g
0zblaF360U3wdi7u8clrnf85loP5JGd3Vm4VULwc4jpQXfM0i1SeEinPZ9fYh43c/BbeJ9cxTIE5
meajJhIQ4kDx3LT26lPxPM8D+Bq8HIYh/dVwlb8wiyS2NwheNZhWlDFt9964yt36nIWJO3FTMCD/
3htjfXupICk1MbFdOsEfGzfzaCtgIGeMojX+cxw9K4uiChYabI7kxvr8IWGUc2PZxuMtRsbtkMNm
pCzomIm8KdoMTuZ3XAay8sDGUnuDwssWST0sWBbEjg0QpdI4r59TIEPzIMBVS4KOrlwTYheSG0QN
/J/dTrU187nP1Kqq9w6NlmYidv5bd+UwTX9si1Q5BXoeXCjIB3SlQNnDpJ7ewNZ+OgcBGX8mJ6Dn
Ipi8l8wKyMY6SVTrU4L7J0QEbQCoh2gweZ6K/dY3PSf/JjkpFa3a1P+7kgmnrj4QQ0po1XozoT3o
i0rJnP65oibdke8kedGwMKzZYiGC6uSSftAhRlsEDQjFsKGoC7cFTUo5ilWc9ciDOJfYWp4IMUym
K8HbKxjrklv93zN5Zovl0dfkcvYUAffPTMlgH6RncLuWM3Nf24VvbF6H40kE4jXJbtpTNOa9+bvo
L317h43OL2uVMl2nA8QeJth47RzBPiZzyfixoNriId19Ag3cA9jx65WCCeZvaa3uZDFS+pjeYG+K
to9sbN3cmqTurhOQBXBqeYSMzYa4kl+pvy6wW9nS2l0AvZyZFyrV3wj31RT5tmfQyu7C66KO/Azt
GAKgWuudjfi4R2YMQjlaq26tb0ei/qkEBbf4fW5q5d2Nlq3oeXFxw7pPON2obzSKe2Zb4t7thBSG
xHaTUOVf8U8vn0v0bI+ZLLVHvqcLAMos/Gs/u5C6wDFHG2D81sMtE/b5mRZJ+iUIceGputO7oC+/
rr2ts3ngrtVDyz9JBX5oCEawXknpjoytuGA7EAayyIv+L+6Sypavqoip3qi+6uPFmCXpQP0ySyl0
ZR3DPuWsAaG2Zx5ibJ7xrGV2K8aHrF8M0iUWkQUeIvVH5Tvb5F2UXiL1vXdvWBa0Dm0CpnxFTiYk
goekjlJXXr2/2hxEP7IzqVFM1vh3IayZf8pQvCJmFEZ+/GogIsdNkls7ws7niHcf1ePFuKm4IJxw
87c1PsodXt0wSdhVwuC7JOd9VwJ16XXG6i3wl0VdbGqlqHah9NUYBAh2Jlkoa9U1XXdIJkDMVev3
nWr+P7YLqqSMl2hVLyrO+Q/mbgjL5GKzG0meyBFdz6bKttuTw6KP+0RpoRh5mnpc8M4Rs8D9W5vu
zX5wAUFWiGGg9s/f2i7g+/s2TzWl+oICOkB4FeGLy+5e1PQvua2KFhWVHLysuVSU8R2tS5UDMyrs
MO8MmZDsBVKuDW6WVAJdC4vD9qhCPlnXyQbLwlzkeaJ8yQUB3zl1mu/LEgJW9XQWub2LV30ouxcS
rHNqAUPiqG51FGhPMIJtVgyvZoafm7irgarcBmcV987KaLzoYdxMhu7zQNgtaK4oiYihW9BhfanZ
wvAl3ZLNbXZ8A7sBIPIOSkqOD8rBvrVFD4TcIZqG33Ds6CQebrvmNTv4hswipBGnNf1vVwTp7Xyg
gfQd+LzxftlXWLfeNKTmR56p7mwFK6ZEQxWoNv2mOH0RVidV4l7AAdp9sZj4RVyxILQLztb3deyn
3Ai9z/6w0SSV3QqI484i+p5prB9G6TBic54ppxO6lVjTO5PMAZHuEaiKEswZWqxlLT6MeburjCxX
OR+KUdchZ1oWL+/W9nQ3lQ8tqa0NoosodQziK30g9VuIjG4K44Rxkkpol7ABv2/2VyTLn44n1Yvk
iKl9Qx9zeQ86RJZC4CM3gGxMZyw2nSJxiGUPSDirusujqmw7s322oWfl4RQYbXAlMvsiVMfVHSqK
UxRHSUL6FNJWHjZdq+DXWdXrUBo6Q/inktPED7JQLR/L35L27WoJhlEoV+NuUQUcN3wRfbxXZlIW
OFwZYH8RORR96qmy5PfKsy/vBO9Ry5p/7FaSbTISKkODjjAOviYfmqipEusmts48zOKZEKpYwr1P
f+cHBCKmKralbm5HdRsxYwdzW389NLhvkxEU93esoAubOVG0M3+ytY44JPWsU/pTTQ1RYXlZiEkM
4EJvGYViWtnhfc5AuCamPxOjjJ7XGhYgDtG93iHFgokGopVUV3zYNpok0rpb0iPBiA8AYK88FMD+
vNyZEA2HMWNisKrYn/V+e88Ihu7z8+ynWCEIfMBOGA1qfbNuNC+g6FwcX6KYI9US68kSC6FTZTh/
JKrKSN2A7XE/DVh7Mb2pjszNPnshZ5+0S18yESjqWyFXHeBQvCjC6yl7x/1Iz4cOuKuJm2Ev5YIV
y1xRPoVWDaim+Xu6QFwMGHE1k7YnncA4ZA8gxtKfMWpeoJ4Xb1SH2oFVVK8MynkpTwq4PpWwA77n
LVSMRd14wJ7vi1NIkDrpq8592utwX6ygy5ZOCLETkWGG8wZRQfTyXndKqizowZOel2fVZpijhnZU
n4Ii4gGdu/suWCQOuL6uTaVWhshUj8/1E/jWE4wy0c+DqzyGBGLCHygy2saXuFiFN5O2RrOawzAF
5gi0CmD2xjeWrYjdgFuKmjUZESt04YaaVUSLokEIDJA9Del2ZIhWG5F7Zi8COMcvp2mc3AZvCcLx
JM6jPiczv1Gb8cD2szKmsOSz7+UhFzDdcBqwhrExs/Vewo13AOcVzv0Wu9mhmGwz7nFSzWsi6k8i
Db8CkaQiTtYY2Rey0yOriQvknUXd81oIzGn1BoT1gTwV8/offqBG5Hu3sRbJQ6+4ntT789O61By4
EaL9n15Lo/fUEd3sR1ISzEUPKbJKJji9jm/hej5Kg0/4+wZMc6/NZ6zFQcwOfaJEQEDPOLTG3NdL
mKOdJC2WBBtK7TvTq1fE0crv0+v49MUx/6koP5SWtrU3e8+N6DM1CyMyoRZItwsb67kXXN1RYprS
D1xFBpLfFaIDvnYPFJup4/GqwOJmHGBkiAwoNFxWqQQsvwcOe+snzMbmbEa+NxKRUEFj2IM+GWAA
DGn+EvIJnFH3qjjKnpznJtr8MHlV6XbnOemlR0NgUZ7WWo41Y5O3evUjOgK7CBG1pFbssunktxmR
YddBJU2mjefe0ekwUxvTqs8Cn8xO6g/kkWGlrKsNiAuIpuYSrVL+Unt8hwmOYzBAl6cPdhIkND92
KlK3n8uRNEytsEbN7NU53EYNgWwXRjKwhUmD4vfOrp6CvjkM2MzEBUpS2XBsvHoMU750Ewu1FoXX
62q3+IEnSh/jw8HePO016nGC9fYcziKOCUivjyrZHZ4gZ0KeSB+grdiFGhZRupxXReExVKGC/ocY
FLMDxK65dZMZLbmT5D6gtg+tgOkWKC9TfvroYbj5viRaw9y9xvREJ3Atk8lD+94X+QZEShdNAXft
ii7n35UQOuWJMGKETx/IW3R3rTs+kgzW0vKIYlcy9cVf0WrV7cwQh77NKwW2LWeD00AwqekIIwiG
Tsem/i/FSvA2D7JRNRzz8H2wKkCRp+0M4AfU2r0KIf2G+uyW2rmU8cZxPKULErKf5je23hwgQgZM
8mflkStSuMFoHlBYZ/7CDSyBDS6a77M01/fOiOqjXwhnflXEFO/szEnJIRhfC3HzXiHyp45CLrkZ
rfCOKpGJ7aRXKKwAmZZ9+rIWhZH6/3CIAJxuy9pzsRTjgZp6j+l8iAN620O/ldtFl5dM/d3/Sy2k
dyPOjxKw4CsMe2QSjLI8Vk7Zb+0r7tIi2bfmUBNTzz8dpSVJtWyOxuM0fMTcKEPadI50BhDxRSrm
Lq/VLiM0x9byYak7v63FQELz1/b+CyjrweiOra25RWRBqOG7cqRyAcIBrLcwJrK8waHm7mMO3IyZ
6ZO1p1qzdp5KsOwJl5VHRZ5IJYhdgCGz+U5K4v/wPdZDk50jvZvSVpHuYoX9ggpjf80snET0ydK6
kZERhNfN09+jqleQfeJLOQYJIrdZSeGRIayF5L+p0guSSJItsoH8C6I9L3Mpx4UFVcVUBSiXz0SE
QHGGHeGzf6X2NjxMGpT+S8pe9sghKzrsFNZbTduFzPzEvClyvpcm0dy+rNKakNpxkyEl9EONcn9P
gS6tL4cqdeKRFCfJO4aCEownuYIH2jc9W4YLTck/ImlapElnjHxSoX5CG+KiCZGjh6CTCaot4RU2
tm55KA/BXIw8YgWNJd0YmiKV7Yorc23Fd+3X0B1oHUZAGOIymaKSwCleBTEDw17778pHR5paByxn
fOHvCmuY0ubYo3L0yclsC5KcPx/KhBdJlsqVN69C/IK0oIv0TvczPUR94QDXU34X/IXU8pbFpWdy
LPrhNB/LYTiJUmL/sYKL4L+FLmupUpRWVGLE7HBilvicQQjE+1GDVH0QRj3mNJbZvSxfdFvdBKxh
FNfZkcfXbVJFRu9NNQqBhYqeThEe4hYPAGdf6JcmIINZOig1TPA+q3uilUDrLomCrZ0tM8gFckMD
PfWo+sgXDVSWQI+41lPwAHCuc90bOG+aygNo+aSNIRDCDle+Xz9fUxSIQNzzM7zC3y7/K9JYC9vd
qTUPny0DqKA7CluU90sLHQH4Z8TPwf0JUOnUphYgVWJltsHlcPt5DRAsdxawmV16c4hjsUi/5EzG
chLT8M4gqw7dTHQsKzmpH2HWJQ9jsIXOKvb1ABKzVhr6uvt35YQ46o8GoqUC9Q1kdV7tehXwdAxm
JKxKA7WrIIzUKm9FslgeMdO5eSwSXhoiqnTLv32KJ5qUzWfgpgLb9I28t59DXYzJMjYwF5a1k5Jf
jjDFzGVetjJrUkUe53YTzcjXjQCRhb9of73b2O2htfuVVBgn3527OdWsqC6IyAN5pGQADCNR8eKA
LWVEX6LhQP9d+Vnhb1irGSA3OX7/XvxOnKevnsDptK7IH/I/RhZ2RyeNF5ZsRx0nWnrRD789LiCa
oKJTtaGZQ2394MpIrsx1piyGaQ3GkCDgTBUndK8t1QO02CVeIzDoZgViQfI74VYPoteiePw/Vi6E
vXzrhdKdi6sW++1hLBtIM4aXDWAJzelEQALUVAN1kQEFwvH/ktFpf9Wi3MJ393MxjzmaRK3+Ytq6
ONcFnznLeq8rn319fxS9yzaF1cQ9H1bc9pGK+vCZ+t1aplx2mWxyYfgLNxAU5yapbSXP62p7cOCu
Qjnqx0Pb6bU3DyOuzccDrW8DtzzOGjTVeuktLjFQ/8xb3hSBlIbKOaai01AkXVo7drzMiGaZDmX5
lGjsS2MTsFcVgxE4FmsVK+l7v3LddYG7+za9OMhm5EH++PRRDAnt/aNlCoWfv6x1aa77uv7wS5qk
A7sPI/AKM6THUjk8CD6DWBX+GfMYhguHBY8wTWlw7LzkKy1eHjN+NbxAvc6ZpuaVlFy2vihmeEc8
f/Y4Grzt/cpWAwFkQ+STmEv0ZuXm1gIagMCIq/F4QWHn0sT7LYAzJGRiUf2KK6xm0V9wqoB0nto1
+/WP1DK/UWNZvZ/BuINeOQuoLjYAmdJdTKWFxqwOjH7ekT+CIX5/EM4YtFaZ9+pu+hFCzm71aPjc
v7QfBPc/HvuOKJLLrGyo7LMZUGMBReaXdHYJgss9X+NNTZZVWmVzUtMV3uoPMrTqnmz2om5OJ3BG
BHULvHY9AJ86uJeOBXaiiARsXsRfX1tMLs8pJ/jZ4nwm6NPflHo2zxI1TIwHkhwWob1EOD8fRiK2
57Y1zHAUALhhWq/AIWivajYVF724ss7dLY32Yv6NoiRRyGWkSPQpkkYTbRYSNFwFhXEDQdEMJq4X
thtx+4E65/jo16wSw3vG8beqq4eRzfJRzYx7otaVD7giWzz51eicH0E7iFgYBxS9VO7GlnAmk0Xb
SzI0WCzMeJUH/An7tCgMG+CGDweeqHUtT8pZMp/dG/FRLrlvyIx574i0wEsBLD2ZFz5JYLPQT6N+
gjFWwGEJTbg5xTXkC9+bnhNlmZnFReBGYrgUSsurhpyRGDVMySyc3/WC75ninqTotmwE8LPc2KPH
h0bo4+QGkdCUtuQHWHiHzCLjXmA0WSmJoQU0PGR1sJziWcBXsF7rKswlqE31jZx2kkHNl5VBc7Td
ZC/L6FY8AtdIkms1rXsPAXoAG5vUNePpgF/1xvjEG5bhLLMGNSTx0M97Wog3gt6sNyjFhNCoQyud
Y8vRHPHsP72QTYLrEdoxiEWflRSSFO1Q1DMVJQAMaKldlwKt0TPLS9aJ7LS/xdk9W/ndOtVIruo4
RE1I8fzIApv3fMzye/f//H+y6zLZWUF3RMs//j5VfFr9WnnnuK/5i9FxfBdq9Bo2RHN9xCNcQs44
K03TgieWHBEioN1Futaz5vZ9H9lMOzOxc2xq+snG6oFVfOqQn8hRYFkx+ielRLoozImJWzh83ooX
cW4w2dQr73TM7gs7rriFKRU0GpZ8rK7jCj4/lPvJYDCOxWQUYhlru8L3XO3bpWIR2/pwTgnvzVdv
kLjX/rxL5TfWWw+VKzSsQnZ1TbXTmTpo6rlLl2wx0TNR/5ZBuSubWj6XHi3LYEG8bwWCj5aI2gKr
yqB30JcSjs+xr7fAGemZ9ILFYUXRwMW7+e1ia7JWv4MRKLdy18FmqMSOVrwHrUKEWy9DrsrsVbsK
lz+iRBc4mgxZSKwXa/pZbfEa2pYr1+Z3MdW8ZfHWMPtdVi5khPnEIyCyMoBn/WhAAYGeQRyJQhPh
386rhIKkz7OJwrDY/z89x5E8FC+YaCXD+bvTYhm5405LZYoL1ujsks1TtQ3NY3T2PebsRtSR4aIW
HnqGLXznjXOQrUC4hL4pdBOXrnA2BNh9IdwmN/b7Op4jReBXpyy52JNWkjBZB1W8KEGFukj5KrAs
PbEjzX+SBX/hvVAs8mtspzlBA0Tvfb1vetNfzcDYYbLFEy+HdpDQuxGkmYZ5D+N158TlK7qXTuy7
TjfjqSEwcfr2qvVyk6AuWGGs1hLg2f1sP9DmjwQpdSnaVnOUlrpHGy7oA8yMYG4dIFCP4eEObpIc
CKgI/DuW2sLWidzmK6kd6RFzVjlnzB+BizFWqJgwJmoo7ZputJi+0+SJ+ggcGNujVGHx/CAYx5U/
yF2Ol2BWyfFT2iYY86UNCl48YJQPn3rPIdluTOBjflCpxlruQxy9JDASuQuT3yzAevyS0AXE774f
G4mi9J04fGkB5q/iWgC4/nxtLAyX6wMwgp5plHgnejAPOvL+bjDgVlP85j7HAnqhmyk9o5NM7wsk
zHy1Ado3HANm8ONNNV5zivTEpgh0ZbBOFxqVTpgm4Qrv5ikg6huz39BfAHwB1aXSJS7STQJ06Ox6
+J21b4HExDf6ydnYyMXp0Js9GWTc9ewOKIpyqKTtXAr80ATuyjH5RlvZHTmGaYdUL+M9t++1Yzuc
6/VK/rInVRBrPdb71c6e0/pA8dennWltUENnXLozqDS2UplGvwtwynvIL8+qN+juU+bKoe4EIMF0
GDeZm2nCsr50DclUiVzPIrJXzcYLUSxcWKfiWNCbawILDq2oII5sJnkzsKwgj2etmpzTfkou8EW7
NDQDBZNuQ6/FuBC8EZHt0hwCLs/Jqup/qWfl3mtlQ/Vi5HjJDqIkCl+6Ub2LDrHdNDAKOTm3tiLG
hR0z5BTCts1jLLB3bQ7vtH7W3ZyklwNMA9rmXBoana3lMCJXB+Fs1Rncxu34phe/KP/pstY7lO6u
dl0hN9HksGAF7kCK9bM14yeTANMNEh5AbC+cFkAlDskE+Xo0HLF3wVCxj5U0IjQ0GDZ49XkWhM92
tuwkXwxybF1vowtn0E1FgE2v45hOZYHKN5il1WmkKfIA+hYwCNZzu9CWipEyJafCDBPbxxUsY59s
JEadxeWkvjioNL9sbM/uFG2zFTF9W3L0BBQDmQUdpyviuMHJjAhkkHQjPoCXHOb0xKUpUAfBinhr
SNqfXYj0lCMJO1mP3V/3iSlOYKrF+PpDDG7Jeh5cEJJ/niLVwDLmcYMOCMRXxA57Iy2wCyUmOoA9
xC3kLLfH6vzC8ayeV5vaHpLnjnydY1R/pfyHlkS0bGCPmumldEyEH5DCPlBnw7QTAxgsS9ICtkVS
Pudl0VbDxFdCgoa2us/s1+NIG3h0kfOiNKvJIBINIeH6fWzPPhB5UXW4XA0hF4ZDRF+kB5L6ZGzo
ZHJRGVeKVmSB1+hpAd/CizT3OPzAVnZ8wbcBzY7+CSeb+MoSI2RTk/uhI6sWFL/Www1Sws5I14K0
phlZjCnZH31Hh/sRGM4RYZinYzpJql3KvpIvDEuVMha/HyNKKXZJ1xYH5heT51xrdKnhw8K+zy/X
5j/jFcpGFs3vFrr1cpBJ6T1Zispt912ArmbOEv75UjjVlNMJLx4QHf7BvO8xjiu/SHc5A6EbwBg5
ji4r59ItHb/BqQVqtVctS1zlgbmeYBLgKKu1c7PA2MXAjo1fk6gD02ZDX/7U5Jf1+uVwiiVcZ1N2
y7YXk8eL4rpwRy3cvXe1+TCqvg4p0cNJFCKE+e5JA71SlnxM9DHhebBzfZ4pJPtacsWo4Djupl0O
Jy82TBkZLLeqvtLZ+D20AH5Ne3lmzJzuUHRgJhf8rQWfVu9lIonvbwN1hwvgfpx4oJygt6eryphG
OU32zrrUMe08L7c9cdlx00i+9x9o8Vg/M+X5qqGl6myuHAK11dEjM7YWuNAfW4I8KV+xOuHCFzIm
GRcoaGhwIsWYEn/YT9YIB1kJXddisM0QNu6x1DmVngQ2Xl7uVMhzSVbhUvp/0viMJ2fpd8Jb4M3U
0tAZ9UEAzvXH5dPwY6I29+17ae0VUKPMMT4OwhnEJcdxBmsh1Nr6I9UIjSDXNABMdj1E6wNcTZB9
Rva8HXjvG8ZEvjiMJk94I8YuW+9xT/RvTLdwuQ5GUmsUjLSiG2QagjZvCGUawdcCr+8Xol3qrq7S
ExdWTyOn0RiUTFJ+Z9d8GxQSZQpZJitWleynzr4Zr0anl4R/ubpWaAa+X/h0UGE1ZuUhhw8E4NoR
p8vm1MiMGqftDM+N11cPgq5B+SpkD5CcEFcfaiZ7gcAiFgM3LM+C0I2/aQZZjBz2i64w+7WmT6f8
Z7jMPToco2a9HEXqBTMxMmqtUMD54eXV5+fFIzXxeQ1ATUBrAK8cF/b3QsNqT3K1F9v1BjllfHjt
uV66bNPf5KYs4hDh28XaNPrNNYvJ0XCyxy9W2eMJj+XUEMahuTR3t+FDLKLHSTEu17rtOTD79ozX
ACdFqiMgni9YEdIjBkRV0AAd6pR1I5+PdwP4ew5Vq25Nz25jTFz7KLe3ztyALOr8VBbwC7vwYm5C
FV8Zw1/Se5/B/Q+J32N3jb6FGx9M5yA4oQakK9DDWR0iyTRdDvTzhNXUm8L7viLXLFSr2NrxSII5
QxWWTfzEiYUrw9jHgLJiozZ5qTLwwvDhYO1m6V3jJ8rXzYYwoCHsJ+GzFqYsE8KprVgCp8pntspD
CXgiVScpDcpSvIE9W1W7bnWCr+v6RDhk2Si1/EgSMk+AcXVyE8ZbgXdz9LXbLFPzlb5ATDIVr9lK
Fhothbp4JfhbFtd1fmvlBJ/nhFhUbCXGOlCScE+ODojipvbgjjXv9GwlPgvWtrzNNpbYHgU1UDDf
Ef1iUIykqxTopIEY02kcxL2r0deZV7QBNwNe2gUpaUepRAbtexNraVlkoeOpbEuxe6nyFpRT3ftk
Qd9J+bi5lDt7AvwaSdWP88dV2mDDFk3Qazn4/GAETm6ads5aodRCgK4Dwb3AnxawpxHaXMQK3N9M
+2e2Wqk6dkVILNc53eWn+ECMcEL03YWy6Js6v9hFcS/gp0LlwdjqhufVGL3OYq7s6IdgmC/0bnU/
lT5Wo2xB9LdxtXJkOvmbdzPJe5iAD+d6UglEGkCiv7gVAkb8UkNqIlBtokzi9ewfYVSu4EzsvXjg
sUTquL3bLbTxeogYW0P7ZYFAMURSjHzSlxz+ZFalSOxq0Ae9X3iPWdIewtdfbF1EEAiju7CxQ3i0
ZDz+zh0p8mFY6MlFXF1dio6dVBu5yfH96oa0O59X5G2roY97BtAvDacj63CtuiO07OZZMSaye4Qo
kSwn4XD58CU2Vcs7bucDsfkBPFz/3zT4sc8aExh6nSpM1xvYBUrsKLPbA4mGUC6J2rrMcg98Ol2b
MV0q1ucr2kqQKavM0fUwyoTrFFelCK/M0ZFGKgqksngPnvHOo+6j4y4r6vcgcMZDTCmwdbfqu6mw
mW6hVzujT5elKfiK3uAU7ST6uMHZ4iRu98cfH6pZeBwvhJZdBNn9UN7gKOoPJ5czD6B+Pa1basMv
SQdbRikFWln8QGqwzqDVyVzt5xTQQw+F7qGYERtiB76/8VhCwepvoFlrnX7yN9tXs2Cpg4zNZPta
+vOmv1xAiiyq7HRCSL49m+9BHDRjBDysH/cC0179YTypI6KbhxY8wbcU0Zr/JeS7KBrh1SJSoElS
rFQ/bUQVVvwvQutw94BCi7oJz/nqPs0/ym6ZJB1MQB1R0JKOozbk7Bkz61tZxkc9lx7jKHyj5kEy
PvqjQd528kPrFPhJtMFiYMIur9MDp2Wc2Fxrhf01DyzhUq7OesJebgKgtCGchBvI/7Mf3YbpeswM
ZXsHft7PcNJb3wU+mGOvDV/vQsEjEizKVOK4Dq6l+u6/vEIEAFbOor/944ypoqUQEBe2YzoJHTws
+WYthPfT5A2iYJIqTsuNHm6pT1yE1mmnoRga2EB32jUT0lUM0EcqH/DWhNOcW8RS/+LKVS9SwAdc
MueXbGQ9M7MKD2HI/9CGwP591JLExK63NgEI030rtIC8O1bRkDh0m1UnFmSLNTxx0n0ppO6etiAc
rMuQeP52sdpWLeTlfxeuCBxVNvwuIuUnCfEnB5oDN4U2ZOCTMjt4zrhGFEbJxb9hbxt1uzu50pLX
FmP3xFL7oq40iR4hee4v7ihmEdeT8jSCuasbaJJdkZdNJ0h3YBqxKYbLwDkzmrrt9pDQC6lSjdCP
hddrK++6B8KPLvnzttqZ99Xc1DDv4s/Cs0kAOH6VkuA0RtzOBMwNOB1RREaTTGKrd/2EkTDmwOMe
C18hh1XAhvkIjQjgi38Rv9DRZxdCrV9/HdLlzZiiCD3gP1i3I6mBcK6fD+VNBnG24VoXfdY7F6v4
A+zm9Srs0hxPfSMOKukPL6WcPaRG52mk3I+fB8oECkYoMs09l+pdbcplVUO/XunETkr5o4d5DfQ4
o4dfy6qFyeK2gE6eZJcKM6X6H6OQLEf/1v88w292Tq2h6S5hbG2ILDAn7GI1sMLWtcazUFlqH3R2
L/7300lO7iXXw6Q0Pw/IAiGUmKBhLeE2dHlCbYNouWTVpmRPKFfj5JvE2Sff2M6gblOwhU0DLBwP
0Gon4EU49DKmy9hQ7DAIYxAFpGCAUkbOrUFY6hYvrFYDHDReJMPE9jXFtwhDdYczwotUFidwozP6
S6iqS+oDei2KVT05OpXu8Cm0z0/XrAWTEeAWFVxI485aKexPaPg5sbtaCShwbuJRPxAFRHujrLBB
ooJrkJ/kptCp+lA0wIzjnzCw0psneGA4dZ0tCUC5tZG6r88vvWFdli6hOOVuyNVCJCf8osyz/vQq
l++oBnuG0gIbqs8MWFaqNKpmoISeDlsYkh4zJKCDfYFByUDFB56NE39dZcVhhLaxxl2wWHvKgkx8
vP8X9kIUMhqrbTS0eFp0CuDH3iPp8GOeFfHMvO5aKd+yogJmBtO6C0yejglR/JKi1swKWpwzfTJ3
gTCusgW/8RVZ4ht2dCTt9ZOEFQnQNSVR9Al91qMuSosxqC8Bua6SkaPFwPnwUs89L8AlRSTDN3YF
pYIReX3U9xBOUmuL16VIiHUNePOKs8b9HYM0s6XSoF4E9UNLmkv3f4TnR4oQMSe7U03Ehxw5xmOl
tGTaFB8UpAJVmRFo/7rXzDM+7iR+Ey3zW5BbEzjVK6MuLSjK/9G95dm2ujWY0mVF2SxTsZHuR/ae
Jm1Je277Vpddkdq/oyf1pK2Iq3Aqb/gi93rgHBgQ/W+1BmMwtoiU8Pliyaj+FnNC3qvn534IjvlZ
i89ZHOSEBLNgzFAivuErfE6ZSW+c1kX9KxNoeNqObVKHefpOJJPpstKLraKjWnSOlWZ/k9WONgnj
jMzQOCxIUEpk2NqR0jsxta1j07wviCbCyfjfV/79Ib66umjsbMnB2v/ip7SVMXVPAQsmWxri1ZlJ
6Gg5PfPLoGpBjYlww785Kz+gSiP96J/ReEB3kdOD3TKW3IZB/PMWBqDZYW6S493GnOdBWHfaXXoA
SaaItNHtRu/HtDttmOL6C4H7wQEIgc2psHus2ZTdpGnIQpmEKaEv9yDduvOdhZlo+Oe/yfPg/yFJ
CqoBFxPsDfS5iCXFkcz3uQXUmF+9SqMPEXhy0VQ3g+vXB0/8i3RSuWkluumJZRWagGeBL9tCdS/Y
p9x9oI2Yf8uJ6RlUDcGtleHIAMH/pB6Q/7ImmZcjjKO3W5mR0ZgPe3Ra/bToKi3yCp/b51z1MIDx
CmuIOSfEY5OlpqFipwq+mzDUwA2Ytg1hoJf6mwDqZo5ovdKubjjlefyouJfcFUF9KDDhJ/stydKG
8s6YvJP0nCLxc9Cst3SPmSnnRO49PoH/lLpSd1mQav6HnYGELyp724g7sCz6U/I7a+WTr0lb19FE
9Y9V2P8aOLaLnXMMC8RmBGCgpvZ+XIYAwKiUcuZM9PEglr/+HFeIjIxrzthaCWBS0J6AcsaNBRzi
xm4M92BRUtvdUi0z8/jeG3Ygg+I5lWJMJ6b5GlPv3DQBBBt1u8lDUukO383646WaxA3SQHCzvMAU
Q2ArXVYxTzP+7NoTV2SzoSR1bNpoI6VoWDjjMqVYQ06tdl4IWhSTi7D9WGowzYwjJLjkXRF/FZ1t
b3QQ4SqxYrsws03e9t3w/2bTpzxM9ZDK/3sTDtqWGwC/nF4+O6M1IlcoA4yUev9BXeuRHieF9I2S
8DGBCF5MJqfTZpdF9R0uElxVsx6zaAkthV7qpCXQN7OxPBF0oP/W4ffwT4RRhdNLRbpXt1upH5sM
YQeIS4dRXYSYiK/dQHo9eg5zX8Zd++313k03RbGNCYgPFXJSXVleju4R3WwLQOFfuaSfQptGvrgn
fOy7uIBOQJzX7juVfhu9sR8ITtnr3laVpUaoECQU9o12Fsla2qr/TlitDo51mizbs3k8eqzIL59C
GjMSOGJrth7Vfl0+ajCDr4BRt+3Q7KcoTVzcgMac+xg8qRbeYmRBcXARK+CgHHfNJXz4OPlup7os
sSRIBAcGl6yM+OZGAr7E4zHu+NtPCcK5dHbsojETgU3yJKnIP6XBpKL/hntryAkz8m2Y7owy93x4
D3iRu1ZUTaqtXnGyq9N1m0xsmDKqARRP7d+Xlv6NSOopNML4KYvTk4bpYB/V4EMIWMono6TXVYy9
ewHSVy2/eIjmjDZRrHgFUA86xFCkiPezDn3KG0h5Rx5c4k1z1pENbKL3FWB7RmPRikxuzSjX++gM
jSu5M4Qsm3h3vJ77lfuownucFIFGcDDq8dfmAuy3bKHRvW8SMW2Sr1Uu/yNRAkUceGGlqBHu02Ij
ZY/7DcrJvDn+vS7Y/TAJlvOjWINa+f5txE2CNSHC/inLxtN/Tq2bkv6VYsJceim3WnJbtKO60qRj
6OB0MI6XoWPn3hIa+uo6+Pi92X2qgXUxoSJkEj/ulEJb1neGPk7V+j9TxdyAGkPBfWNWdYK/NFk3
y2fFrbd0WxFWUvu7vR3JeXpy7S5fFeMSoSNZAtOoLQykKkkt5sNFXexPa6kPgnw8SDqCTvhiD+K6
OJkYXeypS+mr2OgPYWv0bJtnidvDpIZ2JfOvKum4r9FoA6o2Dy4WGfw6i53GpIyaH6l8IXCinLJd
7WKau939L4Iaa6OBrb8vMxfdcFzxhGxHuVlTEs3AWQu6qbNw4rSL/OpcUfu99fdkxj29GXwtX4Sw
e1/YJeFJ4puQv5tfAaJRe+H0Bt6Dc+wUbBGeQX9cZigL5wQveJ3kII1Y9uwmNZuFYr1rmxjopvaw
dl7TLr7CCvUKBoxZE+WXRpwsoQFk6BnrEb1GKvE5UZDbPQxmsz3T9cBYTP5jq1tCRYjkDw8NP6no
f+1qAUM6DY0f97Fl53yKL2TBXIhmeDjLWd2ceO6TtKI4EV9DKLXUQfS0WezYuwo0WfrOJ5CG8b/o
W9GmmQTk5tSRWeN/dGVoN5hC/3l7R4+9V71zVOoqjstfoXt06nuI6kZD5wO5fX42jyz8aaEv1Qks
xvqcNhYMzVCANuutvgmV/6Rlw3VozM3L5Ipi1TzVI4GcF5fXtzleZGj2K+wgv2cM/wJKhI2VmcQc
1ciBhHVsErkMAKV3R8GscIXKBQwgt2gjWtb+ZWQfOeGboWKXGk88HCIaCAV7J0/7Bo/toxdI8XFG
YJzFA7rEKG/pQX5Y3Fkmj5p6Rpb0zLuzOiuW0sz6zrYB58KprC4mKWfwqkzyhncO+5JPsFXU8CKY
vd9pb6875ReN7gb3P1+mrSbSAkvTqLiZmFaEVjnsptKxPUvPHCS14e6GCHd+elUNWjdLjTunMOd/
juLo4tGCBdeOG7XSj1p9QhM2DkXXym2w8iEiiWyk+t5P3LJP1p2/ABt+vzCLa0wcwZP0G2YoAme/
7U3+vz0a1zyRXfCaCFiQJnAR8qc7zZqjqgidaHZtvwUzFIW/0zcGOlSN9qNDDYNRQIpuuTdXfOA0
9mtWoN282ZaX9I6JvnZSNzzbk56jUyoc7ktB3AeQa/4vaToNNVMHf/1poyIQGAMUwlQFEeCWRmb8
ZObmHa6JAbxT3r49hNiirdpVc+nGI/jat++8id/cp+doALHW/9FP28ojuhPU7/WOEOTUIK2mz+Xl
I8u6LrIDNpj+r4asMRMsnu9wB9ziwum4LlXm3j0j/4Okbrzq5o4qVYHugHo5r65Zf9gs+7+YYgF5
nZfRkyN47U9cfu7NyM0AsWt3TPoYZLKfdYcsu7YJjGdCiCsBTsh3pC8rOHj4Qqhtz2rfAYTP2Mdd
13jWh/j1bE5VU7iURB0ASresObck8LdXccDZXfDdCYVCI2NoTnUKn35QixOEqT2PWGgulos2UA/y
xITBkKB/AZbeVfVA3J36KqFYNzrGd2eaPfDkoBfB/GqbmE+xXX2bWHk+cdHWJ1io2jReHEkddiQC
sEAnOP5uzfBSFn6Bu9/R+E0fA9nxYznEGyl39BzlYDDrxzeHDOEQL56RXXvGilZ8FK8aqQeFyV60
fYMw9EBjbivw/PkNM6AYCRDWioowwjzzWKLCtA/lyMJjRZzmbcPigWe4IaPigQM/LL1DcKgF2wbY
nByb7RGe0B0NTwGMFylQzE7/A8+ji+pb7Q3qHJlMe0iXT2pA/+pV+2s7G2C+SYL3LBGjcVGyFSby
ABBSyCnym4ObasJcGeeyqaqVYvsFWtHeDjj0oZREh7dGjBNaezRZ1rcfvn+dYb10pTxIQmxCkAhA
4qSP8kWO2m8O0r5lUC7IwX5YHGrOgTjy0LoJ9Tx9SBNrSSSDOrWuNMZfghXGOo4tGDKPoY32aIFS
FKqaQxuA+MRMBCMvI48SD/gRegy1ax2UUhqz0G8l3AhudUhEahrFikXcs4EGSEgsbDzst9oajmpj
RWi0HRxwqyW7wHmQOTzqMe9zPQmM3r/GAVUNkykGEEq/AUJJRMNA2y2H6Si5fnIa/yY7RDno7W2l
h0kdCCg9fw/38esAvXrC+RsSb41rwvjcbFQPsBH31oIAHMB6mlLO1O+J2EWzc0SXIEhZq5cv0OlY
p7MlqNal9odazdOK2nOIkTzWngk2FlempncVAZqaC0Upe53LOdBWZG28hawh84XW9ZV+qM6lsbAx
IBP7y4DCLBRp1QUo2hpKLX0jjXiVGqdOSDwDdd8Fn91c7tt0+xvXbj0lAfax4tV68vrcorDTUazr
vyZQnUiD8ZUXnvu1rvxdrK7kbB8J2UGDvMxh1OH5Hu1vnBHKcLDDbTe8GQfv4sXGyJQWg2DrtYhR
Vi0fLt6L+4reKW0OgPBO7IMIa7RI5dOOYvGzyq2JI+jpaIqkikd/oHyxknWbz1/IlKfTXqIL6Fdt
a8EjS9AHCyDds/zjrFn+6UWCL+Fld2M4EsI6e3fS6A2nvmG+yX3/vj13fQ7Nq5ZwMJ9QfKAVJxo+
NjcOyAs1Qa8UIKbw51g66ki4AR2VdnaFp09OW/a6D0b0JTqXbuVcqm5L4zNsLAXtF+xCxL07h+N8
qAQoJxJai7rSDSg9XNKKcVLc4TxFZnVjcHM4eQwQRIHrQzzq4Sr+/9OZWIhg4p3W8f9BObcMm7Wg
3FoaNWI7QnX4o0AFGlBQzxgINSLma7kXO0mYlvOL6GZk4/1Ws2QbFLAY4/uOMbcHWRIT4V6edhKN
seXslHKfykav9eX9qHYdqLCo34RDJUcYq6Vr7x7B+JpCUQeCKt/o94nxAi81SISbITSVS8pJiAYA
VpkmQ57UMfxcmrn7gyu79peiRUdWXkFCEjBjzqOdm2x9aHj4ATSKrhK8NDu/vz9ihFIMyhOBOcTD
oOC2lNLuoO8+FFPLJmhKdiwEn195NIVH4kiq/iKYB5OvgzM5UKcpCDs5PV+0FuhKjPe6Wx3/g8fh
IxBLiMSk89Bo+7zXME2Cho7jWaA86dqJnuD5YUkESfLrn9azxH+iVBx2s4pqNEmwANA79GcitqIe
7r5DqZN1pnOxkxRx2uEWHvsF8eu5sw/A5via6AwmfBW5zPL93C156VOdKS05Km0ribXDPDlUJa1x
HAbPWox0ehVxIi92l9+byX+YEMlzbw1/sGMwEF13Qpy2ydkBxhEVZq4OgLlleRN6SGQvx6VIefrc
jpuEHeJ1XnkgzoYzcV7bz21IT39amUmr/VJcZLSaeTEuaHrjBN4e/YLO+35y+aVdcXGktKFAV6wn
L1AUk2d7LkvDT5BR1FOHvZxQHPDVQ73jT1RqgpNEucfZZcfYBoUziscflUJ/eaCu0LqynITc8QkU
KieTQqXFlMfAXtM1zUkTRbnd7wCOgEdrF1+U0fJV5zqAPgepue4IZ2dvMexpZ/kQc8eb2dbI2eqa
AYNTK89xGG8Iy8vBLKKK+j9a3PZnWLixzmsEDeIRPvV7sWJSwiuLADAAZ+HzlIqVDl3yv7cFn+ro
NZI8qRYE7SezniLsePH569KNj1fCua96dTXP6BHGF/lfcP+9x0JzfRqkUL3aQT/LCM2/tK/bObdF
ShN4TaKBUJ1WJRyOyh+bmebKOS7k4bAFEdgG3mO/ORMAFVEL0mJQ5Cx9GaSB47m0Yf/4BIQnTEoI
WVuNK3JfYTlnVtPS0Cd8L99IW5eVp83be/QNDOvgv5EB67BrGAl+YCtjcpQuuoRDMJJ2tu3YDNUI
feQ7D6yuP9UjMNCBPxJIE3dEEn5QX0xKtpbosXfJlGUB3CxMe1wxHbQoX+p2sTOo2S/OdcJnYyM3
lseAPMlVyJ2oOgBM85XNswZAypsM9tNKY7FOIcJ0zDmASC00Bl/vZbM+2BMhMfKhqcG0VnRu6+Iw
pLqs86gybwwX3KM1cHxJPVwcvKubWJNW3YAZ0yHG5Ug4HP6fK8P8UJefzeEbBxe2zKgShLJFmfA1
5o63rb7gcq3MdmeXoZtcd/Ccpf+G0AbT45gLIpiqD9R0iqwwTvQL8JQnxaBAHqSdC3DAS+sFvDu1
xrF43PHLTPpU0s4ooFJTFM752F/Jn9fJ5PUovVAY3w5+LOlACsHgpeU+SlBbj5nqAJzdR+7Pieyu
6ajxdTxkXOaRpid8DyuWhQ9OEyeuijAySOAvHoIj79oWG3vQgcS6IPgyXdHEZTERoQlgnEwKnyiB
6oTaFvUuNBF/6le6Onw2lEq5zla7HQDm09RJ4NG/aY0ss8VXwNqYI8NCgMB8kRy4prnlu3FYDET9
lkBTKWtPDSqjazf9hZZzJO+0HDtyS72V85gOEPgLUqEtqUad0i5FETzSwwejr5xsSZZ+P5FsI0wa
taJ6Rgnx7UBcgoAHlvyx5mlMdeCOionDJfAYuFoCB0oEqXVtlx+I3EBFj8ZRbFVtCEInxQhxuqJe
G9Nx1NJ67ezhar60xo659erAB6XEzfcp95FNxCPy/Ay9yeHw5U5BPvZ/NYevHEZRP/IokdEfUc9T
hfylhIh+xSdgHe4+teUT3UUJKhd/wzqhkgoHCThO2ivW0u6TmUzuFxZNEjPxGudL1fAaR81Z/JHh
dXNyAT3ROsPE2Q2VaKrpg2tgCZMScMtRU2zcK+sztVUf4epITvbfU6i/HRAd+LWeu2Z77BaTi9lZ
U37TPFsayaTHQgK61FksOALPT+7SZL5WFa8dOaTH36VAQ7/G6xsI/MoYOmbL9Hac1uMIgHbp4Mo3
Vmuu86J7bF3YRbq57G6MMzVztV2i3WWu1J2399hWukolrlcgl37xa8d4FRZEoXeNB9b8PvMezvNM
1QDNEB3lK1cP3Mm39vRkPYE8X/U+ZQsrbtWmDq0rZafeYPAs036hVp3CAzlC+t1Nt90rZcAZvUmD
S2lyRKj451pOl5nNRlhtVdn1rsfNwl++Nq11vp9RlruhL6VyIlSOtak8XPV9rZLlWaGcrKq7YYu3
B4quiA2JF6haIWefazKKJDSuoVD9aHs44bQQWIMxUp8GpsUlCkFdKYdz8AI9xuS2d+Zv4pVuPGou
vNBEutBy8rAs2tWInObJq8Zkey+KwZn1uZTiZ+/HIKmaJga9S9A1nm2/S19GWF5lqHF2p2/IBJpW
6hFrcMgAI+w48IRUelaQaXNzRJc6ceaT3g66I1hz3eRRtwSBZpKx7rRAxGk++U/0S4OwWkEaAxOm
qvn85WN11rkopDeZNCIskzcDFotw2fpDyqvGxd6cwskosQSwtv78wVetEKaenHDYfu9/XffJbvqN
G0VAEEWuwrqPyCy4yh4HbMHKi17SkpKfCMAguwansaoaEhPrYUjcO4W3pdakEIfcKHg2YxtUkCn5
QE0hJmhFDKZ7IyyrQcxXAfPkT1z5xfMU5jAXWxM2ixer0Hr+0Vtociw9d1MKV8ZZIKA4Xkscp9wi
lgrbpUVpaSaSdsH5SnmXwE1fqKPLy2tmaedadmlosIwiH1JIAbZKXIoBEHTkcSFXl8wcM8fbK6TH
2rqpwVrXATeMonw4ccMkmFfZ3j8Ba01Fqgs5XA3ZxPboAvxifmA7WXR9w0eKUf87Hryb9gjiAOmu
Xgxd+Fh9LCRKdNiWMcyhUwL30iF4hn+kBDD7mAEv1x7SpRD8TEU2DkUMrxfFkMB2tbCCvx7SlG7e
Qkd8deB6DdLfpASPZPDkhf+i/WwymaZWvI1E08M1UTfqehftwIaR9tF0asIAjoBYI/bon+flrLYG
8lfXXb+0jck3r/lOe7CY1ljNCQIVeqstZ2sF4ES0fOa4qrd4tPYD73NvfoxqwOWb15rLo+14CIc/
Pvx9YSPHnYKccxcr6MTocilbRT0sN2kxXpDhMlkS7stj18ftk2LQM3NI3dCKXsFRsRPzbLs0qkCV
z4kUO++0zdk3QOI/mh1lQlYvLD68HicUy8NH3s1JjZkum0AxoPdm7C3QHzXAcas62x36Zl9HgV/Q
kusSokm5+P/mWZJvDFl1ao9gTN9wTHt2koQt0+VlucsSrKEQcfrHWyu212uKWRI/fq8tjIx/038T
fbeAO1hP1rEsL7BBR6et/BhTnKpGcbpa4nzB62lI3cTAmOBacxqrGx7x6auY8fZsQdup3Zt6DCQ5
cC1oMj9zCeUQDOKAy/cYbRrCMqvo6CiFIL7sOXxuti+nX0snsbw+2mi3ianfALlkuxSuN9uKWCwM
ckiZOdwGwgh2gnPdL2V6x+d7btC9rsUzRwC3/OKiExIFAO5KTm4FJNSMXQhunRlEXSFx8XOFHCUl
pzMFhnk0x41+SIhCEWZbiPE90Jk8Lm8NJQ8HMIkeHYGQtzNnDkERrrqbuIwOBeGkkI/7xIbBXk+A
2omUcLd6NThtuWaXWgqxfmyADRrCbSORbENP0MhmMUrA8/qcKhjSca+biEZHBwCNBArEOkljuH+G
mLi+MAaaaQvcA3Se5dQDmytZbcRPtXbaez4ifm1OLQye8a9tXtwZH7iLCCtyaEFu91XBQRCnF4bG
bvLQtHPvf5W3Wcq3Jt5HHiDbD2z9Aby8f7sVrl8mzDbi9pmkCV2hHyv75nQRj7p2Xdu2sylRUj20
4zHVMp0k34KbJv2di4lZE26YdHlvZ/ve9dOEMwKzeB59nuktNMmT0QTvscK5J6BQ6aKGRiJVocB2
+Odv38bfQVf8/MrffrHDUQ9riHq7k3dbDJKxYJagVfyNnl0nROEQL99YgXlSI91b/24Lcc56DxJQ
SOAuTajMZJ6gAPrnkp4rve5aDELX70VO9CqOMToGdQG5EHQsBDlR6dV3Nta6uwCTFFiTG8c08nj9
zBDFDHYCwRGgTLJP9jq5UqPxf0fyV4m97mJUeLe9zKw6tFj9qbsv4UQud79e8feLZz8gWshJ2IHM
UA/ER9CrRX7usej7J/D4glOKF1gAjEgHKcj48KqSRnpIFYMpU9XcvvQVdXgotV4/gvHNIa/jYb6C
uNFoZiaoFCzCf2OR/TOD5A+iuF8odMG0ucyi/MxyGoGalzG+b9btkvnehMnHk56B6zC4sKEBEFS1
UB7C5tccpe29JrDHgC3FENcFPzlNUa0vvgLRRrBHHFvuMDzcotQB6S3MXO8Gm5pdSDf1byqdzj58
ef5ft59nbu+j2I7f9lQFPtg2sHY+OUplsJuJ9LN3fXXVf6f7WUSa2/n6f/AIuXsR0SwXGiEWuR5d
DiImc1BMesmGYQH8l9uTyNxVs00h/7m/eY93pOttZTB/ySQYa+zuM3wApX6Fj5/QOI6wAbx8hcis
v18l4GHvIGti/vlDN9Fv9a/elPgakju2xfBm+w24tMjoCIPpGVDi4iOWsxa6hRrsaFTdgfAnIhu+
RwEfXjex13MwR5bnGgWprQQGggpu5Y6XaHV86DgFLgTU/XZlKV8GMu6hN/VqL3TZ0agR+Gjl854e
Qad+30SWuWZqmasILS/RdHsWS1MfA6XuHZ30h9h4ZJiGtpFYjqsr3TDY/m/KoEgCM+262cGZnp7K
SvQxvzrUFXCQJ2rSibp/f4MmM4f+xIHO30BH5Q6K6MVidFSumnJx2B9B6TF6xIwW1KLiJC1jFTe4
j2oXPlhcOp8BGxo3UNfs9dlq4szghtahzTxi77nSvr0LRgjSJy8gCSUWhsW06Cn5l5vRjbWfC+gH
HHUyNX6GcjR+FnvXg2PyjDBy3NfVZatf5LkKwOOINp2NY5ssasH4mRDiTC2MFhOF7uXqe44LAyt9
ikAqTXbgktv2wnxfudEiwla8mT2Cz2OpU4AgK2Eq2OrSFMD0Y10fTsb2ctiZRIFvIOEyOpkwRF3T
4U94JttLPSt76A3xdPPG0YQZm5gvUz83+PxAL412qhaoUHCt32aolCkc1YUJUhWk2+fJ4ljneMtD
U4hoPfGZ87s9MaY5oYpCRj47R6wPw0GHVmOZN5bCZ1ftCdkANo/QKpIOMwvRBbGFxWeEkWORqOTU
x05QCveBCInpz8Rqr30TmVdQzsF7DLDnXpEsp/0ApjGzKG4iW/otfS0tjJRl//n7NPD5vTRRB/lg
LSyn933oi5qrh7wq0fEXUfXPNHSF/pfa7jWzDPYmDd9Z3mRK4zbsKcYBudEhIlub9w3t0q0qbci+
N6Qdx9bXKa2CwB/aBhKJvqZYelH3YeMFj4tL5YCDW1aj9jM6Wp4CWs0Y+Hxs0xZ3CQKNczZibG/l
zzFV3RmctwmCye38JOJT5MfsIpAIkqcyN2fZw1Ff7Atyu/jsbdqrvi2TyVQqw0lwbCU4kRp8t2uP
VjwwuZB50zMRdKbNrS1an3LbNhUTGrPBsb53WeYsOEL7sy3FyCC5FPkoauJzhuwGMJ47GAFf2tEk
aKd3ZKe9IJ6WTTgWbIJjW9nd3sGnq4jtTTqiEPrny8BhFpbAS5WmnaCXYzYxfp9I0dWlDwo3acXF
JJlPrqxgVKzguSi4hqa0Vl0h7N//E/uDJYZJ8ZC9yoTOhHEw8Zjy6BgV72K5GAh0PCO8jeCeDrB6
6jgMaKCUQ9O9AdLTxOIy+AVSaOpkARaJbjdfwdCCknYrtNtpcKfHb29qVcQUeqse8jzz3jaUdLJI
FGDL97q3tP947LZbg/a2vedLbXwFgYYpD2mg/549P3H1gvBxH8HL5bDB8Dh6YC+Yh5I/p2pjqGMw
kZ42gjuTAqmlw3lcN4jGaU2TtsQ4haaxgxoixETKmBq5SrXONBsjgzNgfk2WsyMRpwqG+xKeXz/z
ubcE5uW2d92bj20wDrOUAHMaXKNvY2+6iw3hKhL49ELq5C+SuVOl1Y9JXLsCBDTIjR8ST+skuvBb
Sowt5j/7vUW/2yW6P7wMX08h1eiOqTDMO7dDyFm0bp3tMk48B5UIhQ7/vriAovxeH5Bplki4i8he
cpJQz8W+NQVEdp+8++uQCubxsW2jWdsvl6aseHbRU4fas9YbVTW3hi2XdcgQXd3sal1FaqIi3Cl3
2XsOLIJGz9cQqLtXJdxxhrYd2H1fTtqREsPKCdzT4StMqV5NMtz+6svZ4R06nj+fZNXkoQ0TvE6A
ApPrXWYnPyl7Pzra14HeiMtlxs3Hfs9QA6EmKi3UezdZQO5CxmaN1EqavikUpu6n2dVqAHTVaDif
OlaxWf8o2u8QLxBv7xyygnB6ZCG7i9bcc+7yDKGzRbdylO4XkhrmuR0UzdIPr5eYe44tQN4ZZeGq
9KFTTLrqaj9pL2SBRtzEtu8N4risWwk4RBKii2qY8kR6n2NLJQr5mrdbtY8mQHaqjY6fbd+ExKI1
0vwbhKRojTuPU/REMIkW66PPpEJzgVNnWCqDnzhj/lkciu9eeKjvVjfR+G+hdjCHvksvIWPvTYZu
ogvsVU+seeOMdCyGLGVnYXQP/PoA14TzOkZTdCB+Bt48CK5Xq/xGXC5z7wxhcHEkYHNnFu/Zhj0H
Xd8ufRVB1Wh0BHUrRZm5kka2tHAF0IbOiIl6v1nrzKho/VW3pSMFYBZw+sIe4D+fPvyx4kPrDVTN
KLZMxpgHU3gdVfufDKQMCDO4NBRi5nzrA1u1EjcdkF54FiPccTaTBPffjUEwN3wZnzq7n0mPcFI1
9iFBp1mIHN4cTRuKQyV90+AvXAzwMNxOFGuXZnpn2F2WEXKsq7Lfmvi7+Um77w3r/1BeuULK0max
xXNKd+KpkIsujRXZxpWqKhO7/AzfQyQd5oS+JzAahvBANSe28QpXcOQjU5W7QXfZhoqLD93/XWuz
cuDeQ9npbMvinQnH41y+mDo8UFhNttyVIMzXm2nuR7dS+99Eu/QJTykjyzOgx99yjumNflHL0mh9
wVMPjZrVLk8fKVE59l4+hCX0iYiYf/TT7rIKV1HA6AxfqnWpLbs6+U3r423vHI1wDycwAxEbTwb8
e9zBrEP0QBa1ET7QHxzg0xEFqyOn0K89kGCjjTLz0AL+lEIfICEs6AibI5HcCXtaPszExmfBdCIH
k9qsY8BJKvYCaGxY/4AbeacFSCBHtlKdu+nRrrkFE38H7EUUmVEYQSZDik1BqOJXXG4OPS23XYx0
godYfEvYHNV0TUhvz+76ggLARPkKk8wpEp9FxxEhIwNqHLUQoSQUx+PY0Ky8SOS69JvQVvQcYGSi
JHy9X5rbRWRu3heJXWNn730mxLhEhGlKYN9A7TH4CGtflntIoaHUGOxIdTuFBU7t5Iwx+HJt+UW2
jaq0UM7hyzC8oPW8Nr3BDpPmyqwhukLaPWFv5aT2JHbLwugnCKEGs5d5OQuSXaE9YG/PzxycvW/C
ulKB0qv8qJ41xVF3YrIX1Yd6RErCnAOl0HF+l7UlyojTLxWKcI5NmpSNU3dtYaEXU7fTMsDSeE14
+e9A2zcO3+rjdJONCS3fXTqL2SEMa+1471ZNz3iCm6rNgWbabe5r1AC9IWi3dxmV3+02BK0XtqQQ
8QXMHvY7YMxLkZRVpSOSU1CaXrx+bw0o1GNnLetd7MrDzbV/o20jhaxxV9GE9eFlneVB+DLMHD/A
H59QPqewQ67+Vl4kA5mInUkDuRAVUPDSK8BQ+WYkMgCeUlEQKmpTPTAbQx4fEX+YfxQ2Dfi9DVt5
PtfL9kpW5lAwL+IunlJnX99cKvwhiplVIbamkU6K+avCM0AAKMCb6o1W4J8RFO3PoXf92RxBSkBe
u/BOHbBYIcYPsU0RfesuYWVgn0nxe67vueVpZuuhkWfMhAwDAu2VCAtCadGQFAeMC3QPRGEB3/Pd
6JlN5qA4IooKc4Z0rbgSXD52y4GVrWXV3T3gOIZEremcohiynawVSyMuTK3Qr/AD21NlISKig2lq
Wj60Yr/NlyN/20tRg3ge/Lq6pgKDZilCLsH0KKkh9JqD6TGNUC9DXWLm49J8hKcoKeNlZrGDTciu
piN+y2/d1PDqoeua3MVfswJJRXrrwemG6BIR3YA0Q/FGcQHcEGzpI4p3b23vs5g5A1n9u455Kws+
1RFBXl4OSjkZV/ZH1pYxCzUSF8U/wO67Yrw67ymbZ1lAxAduxvIh3imb54a5kgudYSrHdYzXWO2d
V5HbEcLuEYDVlVJ36g8n+yZQEZNUErbggaM6Mjc2fOCJNog0K8e0hyp4bEKbhQu3qOJTIjFxmPJ5
ksLRhDZqLeWAPpN5xrHJIUknHK9pVFd2aNgrX1f7kQuNb5WXy1UIZt+ZQgQJMuZVcfI3yUtmIGBG
d/s6ueUJdgFyA7izY7lSmE3qRkB1OoROC3ULjaBiTjvqMRlZ61Rh8iND19Myx7as3IFBpYfUILNG
rUvs9Q7/KKidKdfSJTmGSyh/kDeM4H+wrCUiVq83ldmZv2VhZt/NWJdTnHrCuY2EOzdZvgbbAczc
kOz9Jhqqsn3ii4o6aPLlOl0uL5H0XydhJ5cVa/o53TwttouhK8pkOBFry73JVKjFaYPPodZMrtxL
bjkjN4+5JwZgNOZqxEZPM3W+lq957BRqyOLMBw+jdFLwTvRSBOXHsXjHX+Wgn8XvqdSC+OItwL+d
jljsLs4FwPBvDk20gPZQf+dv2wZ6RVjL9eGWmmFeOH3G0jplHkL1z4WX/UgOz2vC7o/ShUaaWqEV
d5ASjkhe8ZdIrCDDAWoTLDCGYnWWF79M+AdFYUjdUxt4EBg0KrwyIewtqDGMRQ8EFXnECDPNvxcw
MELMcaWg55Xh4f4O1fbNTzCopuSB3MGB8wZrmHPvtJwPFidjmjTYcwC4VN+CSDXxGQ3E4jp4q/av
K9mYKsxfaS+9G5EIXdUipcrGflTd9uaHeLeDldDdeAznRJQ79lFSYzTGmjtVRdSIDtMYFMYnu94e
tLVE2p6Z3N19xW0QO/+Uy2PxaE5L+LyBeFRxX1ZRhUOIYWAJbDUkFoOkamYKpXocOeaZhX70J8Ck
/GBPEV6+QVFrYFMKyZ7q3JHSSX3Db9uvBUWLG1nbIsqNoxiw3AXgN3tTmrKy8AG5EWq0u5a3P5uA
lIPjTaPl4yKZ8qfXqqcFgAPNI0CHjyBvWUEDdB7YvcxS7DrHOhY9xojRsoJWpBDAeEUq+mMd4qYu
wlcnyFM0AHmgEEd4DOpceOj1LDDSt2XFYSz2UtRg+l/KP8I11ZI3oWlKtQCW68Lg9N0WYwld5Yxa
pjFEvMiCh1kDrboig2ySvC7dJzhtr5a25LktdFU50gGUVLAgBRov7s4vHL4Bg2nEk63nd/hnQ48b
XW7p9afR89ac5Kdeop1aw7OA8QXpyTcD90Xo3G6FPT/PGb08rccfq2tCsgJk/GMiN2o2rzUrEEzj
Im8OVmo/HL7N84fqkddUs90wpiUKmPwWSHxKGM6aohHJXvpS5oHloVpRPgRhiImvWGOx7fRW9MGF
871TfPIeBNVx9+gohUSE3ewvUL2uR9CruJXWP2DwrKPnkKZrPmJ4stl9944yNiql1n5Xg3audCti
sqyloAPPjK2Gtu81mDTZAL1et0F4UVk1WJJtxmzYijurc3Jc6SUA8+uvEhFH1bxDG4W7M7pKApsM
IeYpuphPf2tvdyMWzAaSc3PMToPr28d7q096UgH3SzEX9nv82ZaMKr6T2fGuR4fvIvVFCY44zlRV
ejTfqfagzDyFq6J6deLYh5t2hPnkqTUwFh5uF01HWyJxfZnwPtu4AXt73Psvj/r2+IgIVlU1E2mO
X6hpad3aZ3CJh8uGLEs0f1B/QefaaUjJ/t8QpIAjp7SeW4Ad4VdsEYc2sTXJwiff4J2HNaLpopPl
HLAs14tPt5HApF9BeDdZyneOijADY3zBwXiwVsBRD6RGGYSPRgwrTYBCHzRBIOICxun1XVlrdvIm
ARDAydm6NMHDVNMC5p9fMnISPkPL29lTmRz0DVHLgY+jL7iVsPEg6TjvIQsUXZUujHWoss30suUS
IyuX2rI55byZJuT6VjRnDpyY7GRSZ3IPKSRtuU2pmLGykvkYpTcKq15ORBdKNBkhPMN6QdlB3ho/
/LJj92DeS2YbssSmQqS6iaOLrq1DEoOBgdmtBoVGQrZqh0FIWUOj2DWmDXTo3VdZCzbpx2xr6BOR
i2kx3I05c0pHl2W4iIxU2hH3tE/aBdD56FYrihhTPa62YlbMCtT2O7UyjyxkYLg4HLS3BrtArfLy
avGJZJaIMag+YOLCWtTqyicA606n4tjM5x79bqJDCCriccIeDaE8u4QDMXk5l3fjodKhzY65J8kM
nwrMvpvxo0isbc2AkngjUV+Mi/tVqD5Saq8Qyvq8yNX1tpzGOgYAS5nz77Hueu4iW2DRfiHdKY8+
4Ri4HrrV5RtqsHF/44gPuUg0jPhb6miyIEx7iA2DFRjnY4HmO+iT7iSwuuJHNa7xGtz2Ee8iiEXl
VZmSCSwi3hLkmMIZkR2KyyFVmUj2Q2PlKxGXj3N2fPrKFHVrG5FIsmw/dq9WHessSMH4xnWagEdI
L+NdPdWo2MO++k9Fm8qe8Of8pJ407TKRdCmbPstYouJMIWfgxB7hvFMks1nFdqodfu6epeM4F2Rx
PnutGo5miovf8ij3r9dA2SZCdTPUCByZFnDTA/AxSydStnsYIBHbQMcwt0VeVn98DieiWH3fBjvE
0Ij7LLMwd0Ehp2h22tnEnH5CLuK1tJYUFIKJJqXDHvJF8VRJYbO3yDGQ2j+tq5KxWXHih/1b0yED
9j2y8D3CZegdCqI4oNOydcpU6JK1uC/lUBAJP8R3MlX+zq0lS+TNmLsXFigiPZSSov7rye8zuLTI
5cYoAeMQl1pIhBtzxTdT5lw9ZRyeeUaW6eeFli6YZ8sKNXlZzZ9lK735FpojdfZjhe3b7VmJ7CBF
AK5IFD6faJzOYLmTIEYUPWu+JRNEaDyv61kuZxNr4waLvFeIPrTBE50F7iGaET2Ehp8Z6i4wHi9c
O7rq+j9E0BgzsWzB1hztNNhKS3KwZh5PUkYvzFjWsbFkIB3nm+JRDqrenzazC4oHGIpwqXSuQFrg
rPG0pYKvnf3/VhFYk9wpyhktIVFucMZSAu07S8BqwEbWjA07YQOk2E9WzyqraDnvdGTGBE3rW0fS
v5OJvFK/Va3nxR3BiBynHxUKDKp0xucpscCWVgZBEmr5yGlDSVqmblKEHYdPPg6CvsVH9tHmnRMy
CueJ4FvdIluwaodn9HF6sH1MVcQYgWuQiRUI1J9ATQiQrbWjWg3VXdr3GKBvshIRRqYYYy+NJ289
AHbTtplyI4LJWucj1TRqk6ouNiP7PPW0SGwduCbZKXQhy8BqtKdWMy6rs2cHMHxSCMfGkidg3kO9
2QNpXTXpm9+m9H6bJdE9xKiiOvZuk6prVEQ7dsqo4bqu9jT9/p25eX+A2BSQoUeT7bx8wBLePGV+
DVFry+Lq/cIlTHQaLu++8f4Oa4gu+8eBlGO7ZYj34Q6TiGQ0hy+cFXP7nzcRLdCxT5plCZTkz4r9
jAkqspX4PQDTSu8mOTBN674o8uBjO47GIbsjQ6jIStELeKCx57CvU/VUqRs3ZmpVkiIWyKc9+tKM
sRNC59sgyMYzrYIIIQ5Fru2WCgpW4ISRJd6owV6qmq8wln+U55oZ8m+WdGsmrmp2NV5EZFrR0AkP
6ejTEf0h1S6/SCJ48zzVEETtVI+6eDJQ09d2X5MIjdZNqwswbZqycDsZ5cgnzpjqqXf82lM7TL3H
4j+s9ghFzTcErG/+EsoooSf85gkP2RIUnVWWxOLXEvONIGtKD2p6VYZM5iaKfP9U5nj9amH+ccSP
/5PUVnZo4WAH6PPMcan2NtyyxZ+igxV1/4UuSAmCBLFjN9UZKYR9vBmuc+GMuXqtMtJIkpP4A92r
ClaPeFVIVHsRaT6xewPlOXEiscmEgLpLnpV1/fCe7X+h84CLS0pUwkTzqwIf0VUfuIv0k0+Da+6o
8qmHzZVFO3yvkDzQi73dQscQz1tDbiUCB0pPKAgatTFOJ+5RXb8bMvbuIj3Cr4Ns7Mw4mFH0BCmd
q6rcnetoGoi0p5SICVk0nbLC/bVo8S+J4/B9iFnsFABQFWVBgsJsC+JnzFlK55ISXf9WlpJ+1AJn
8Y/n2BSiejdPhzixKlQOl3wrBz9T7PefxhMk18VLx0eU8VvQYomah3uD1wat2JlNjRPrEwIkq3hN
+nJsAyqoXOgGGd/r9ZiUuM5KErrWNk8ifrP5X/mZ2skGhkzvSZN/eCFHiRRzig18c55TXzkcE52f
B6X73k7z7WrJgwSWw9osQY4RGb3z4PGZgPwJLK3CpvT/Ma5XrKnlmde/Az8h0tYT1na1+7PTdZW9
1/IPPNSu1IaREXytOk0ZOERYdo9ReilMlKDk7sjpAHtoS+FDYcUpbDVL+4QipgREv1l6vR5L/1/F
bZ0qAuZ2oI6M19gsa73s04lKlMUN0UVr2iPFzdM5sJAV38eW3a+bKoDkbZSCSMRTUEtD4jImcnwY
kCLi6GkQvB593DaA/gwUkp81IhMmGaFOuXcJJJbyMCodft7CcVnbbBgMuWukb498g1U+0xeclPYK
AMsZe48iht8kdjyGE4xC9ZUdECNwSqcoV9EK36KrjDDyIiyUR9MebVpi0OiV1j/hqT2wVmHpRBJV
GTvoVjL2RYpLXUkD99Kv8ydz3JXFkb7Ooxdsd5sKut8ASq8hgHUgA+iMIwR1UaYZpi093AsMbqP1
YVC7jeK+22aEhOEWX6Q743xS0C3ySSm8op143X2KD9TFDSWg0/8cbDi/CPRX8HEDmaoMCyb0Swxs
/hTxseE30hlKQNp4/SYQnhdl7FwCXdM6QBFk86MZmec3iffXRVSqBvywTkz0vVSzsD2vHM6ZxLtD
7GGmqafrV3cvne0cog7rmRmAO9F1OA7aZybIIo7RVaVSySSSP8NzukNoqNhqleDnL/ZDVXMPV6zt
svsJHUY4ho949ePgsLvJmYEjsQoMZi72JMlPOA+WcKSrQx0+cwPAl9RsTC9lovkRmdKVwtjvQnwS
+5BL5DQgiM9sVzehbNHN5ppqtF7up2VK69AWr/f0UC8KnNT1Mc8yC9X1tFoGSCu+iWIuYirtRuyq
SKgW/QYo0S+uIQM0cVJgKZfdG5T/o1HGHwcB4dAseSxNfbBQMW24NGIcifnS+10jGWPdjpU2tYnc
GoYEkVgnO2i5sVHTCZ/1NoExLwNq4kkSAMAYMdC5sXA+Ch8sukhW5qOwqbvUMajtLOPIH50Gfr4c
8ZBozQRHCV0U9Aa/Y6nwqclipY+u0BUr/mqHGs7LZ0eWYAxHcdSeyhKP7tuc6l8buHcnXhX4G+6T
buT5WI0eBa09q8piXRlVd6hl3KpeJ70mrPyiu6vI5ZRp869F3io8XmIsVqOigOxHVImQR/RTrs0C
Fx8/oSDRjGfbS5qE5cbRUH2azAjDKio7gAu/xeryXU8EQhkfA6IPdfvY5nN77QIwMS9ganNma/80
EJD31ysKOxWTlTzHIJQmk2i8a3DlgCM+/EnaQZe5yJvauySOTE7uHp30032uROR0mfqKdIheTiEU
MoW5RoKjUWBTOmDRNE8NZbJcy3HqL0mf8dejO4kF6av5lVI3oM8i97qfQO9mjZVE1/tb49u/GPmA
pECR8yC75CzE2VGlrnNydVQD5VwIXxW5QGpKyD4wZstN8MN+ABrs3rkYTOINMSyCwGIB03S+6Xg4
UxfrkP/vrHHNx2qRHV1nXPxAfeFu8WM4SJManuTWEo2GcAbEqfwa0AlX6A7zOO4g159BnbXOQEdf
yRKeSUEAzI6GlXtFl6ZMv5aTRt+wEX/zV6JbM0yGzXwBX/uoYrQ8ETxnO8uNP0MAOwoV7NhFjrdz
nqfQw2wSWpU3F9cs27JJ7qcr9dWd2VuXbQOo+2p8n25m79Y2eMI1RI5f+inRBV9MXpdZCe24qv7a
jAPuA8QVUOPv5WzDVRufp1m+/YaV4rzEQPDNbZwOiykEvmalqN1A5OlNX0l3KelXRPxY4695COAs
xkxjXNO2CSU5OAXgRvRkU/ybDNXu+BYiMPh++LPeQEfOfG/fp8aofgxgQWL8yyIZ0xmWYfMo50SZ
PYnB0SnKaaAvTcD+St3SKMNxQZiEN+5DGSCXO7RBNlRRFf1IePK5OVM6jlekZtz7/s+Xz6MqOQNU
3fOBNo+at+m+oZcnBKoZ8RaBTLWcm8cguuh4CzjTzgBXNZENSGt7eVfbg5uJErNclqBw8ybkU+WT
XbLRT8sI+oMw+iMQxm9KyyYL/KbEmfnJa5sHG/dxeQMhtHkSr+e3mwHpc1CIvZoA2g4OJr3aVxUt
+vW45FeU49jWhdXbJn5nq6dFaMtoEkCYeeWhwE3qaXZoBl45LuGoa2M+v5Xgy5ysM7gJU3xBvXdT
RVZxwxF39NYY9dqDoyVXMxDXCeP8Nn7lMM3jEo6bzfkfnnxYQWujv85ZQbbhIkcRegHufb3hnWzM
+tlNT/Z3pJMw36R42g9UUEHSxrwgkWi6Vc/AdM8V1dlhR24P6sxqZZdvF66TdF2b9gLQ+tSr/xjF
0Tm1w60bKHW4YM1uUXHYbWuLbxwAip1B+cppwjL11k4NQG3Gh3jV+tTzFJOJt3Ywo2ZmWcWv309x
Han6YyItgYhsThwyEMHVyaVNWz8lIEj/9lpqIHODXTdQN2GaQoCfcrNaFdxspGnNwOUC6X7R2V4q
xdNflryZlxukdNwfFA663hh2xeM2/VNfEO26/d0o07q8mLYLLJtDFiNis/HbNg78LM0rg/PYPk+R
OL++doLjHHEXv/TEHXPtf5iU10uhCHXZFBFz7jqS5NtlMRaWg21ahZjkI/3lR9oouusogTAMF198
NZ5Ebf+sUhDuF3RPuPYdFTKMH//vuhV5TBt6tJpeW98F0yguTMwBzsd56JyXS86PbWS79b0Wns+w
IXFbtD8sT/m3En0aZ+Az2f+Yd9rMjYW4MssHkkS3Lfdd6Ia4hAZZdt0IpdgbY9+Z5t8cgUEwfdK3
p5cVzejVNC6UBPj3gQ3w6ontVhpWlTTu9FJSioLnrQcPfr8leBSuYM/mvsMiddz5ySejooFCK8IM
etAKUwf498VivUz9qs3jn9n+keZlVsxuP8whK4kUhYU/q61U0RQIRoR2y4wyZuZh2coFLyWbk65U
s2pFq1pOjCz1iabWuoYWE6Uydt4HAV7juprHJKigVcjUAegsIQApJla8D8uEzGqC5qwAhQaHAf8A
lByC7Q4oDc3l2WQleXobg7J4Ff8yspxhIGzFXHAH2jxAmL2bHYVMLIAYA+Yqq4IW4UegxZi3LZNN
EuQDVDqhyW/R0IU9SIw2cznXJh7FW/3qob9e2SBMlmqSpo4owduWgeP8qyvPZ2Zv/gYMByPZb3FC
oVMu4yAjBxTYKuk+2mXbxMok7RyuKxKUsI0BqW7+Q8LSlDzx7YZfiAanw1DNQBVPABS0J3z8qRFf
MDH2BPLFHTPs6Rws3JOD1Cme7aDE8ZYlIOFFlMvexqlgU6WRVf8mkzLkGeizVEqvYpvV5ci+3rJF
p7DIPTohfGbuhevxoYCOOlNfZID6o5YbC44i9Hl3H6JoSQX8glYNPGDwMvk7xRz7eaUvx45NtScO
YCUuXd1aEJGsQsk7Pd0+0C7jYim/wnIgK+HQfskSOKv/u0lMP8mBhhOihUS1z9GnmCwkec4fiSFp
R2urvRK1gcZPu6naU2ZZreU7CfTwTFBf4BV/P4l/6BiQ+M2V/re/hza+RlITDx7buXp6gtr+YbTg
D3Sf7qNkMU11Otm5CP3R3lZHCOTCaERCBv0z5I0UZa6JmMItEc+O75jR+eO4A4rd0hKObLMxK7Rb
S80W4ojCCSYl+TBmRmtw6FnSnxmzENQAXZgq5YwFExJf3PguFwdCOqEgL0BBy6+B8Eo7dZP4QAma
iktYjjuznbfT4XLyYU1gP0bw6QxdUCtuvfDPy/Xn2K0n2JTZw2lHUHKUJ3yJvMdgVHzmFhMczAwf
Dtya8sCU4F5w5Rum0H1djaTDk9EF9gXcOLEowjx6O6xCoO17k/5O7Dce6B0McZ6TAl/gdEwtkScg
Br2yMaHuorx9FJzBM4vQNyNmXXzmR1IARzLI8PtWPe621FexvPWHyTOPjkRVK/iuca4TgBUcKaU/
7cmsKH7qRz860CSTe+UcNclRDaCLpqNTJblgCInGeqDdkcaTErvcMsSeIEfrTs8NLCcVoZIggjq6
6hR5K6MTgN8zDYZt5Srf3rLFmnKHqNE0kCSKZ4i1df4vDzictzFKruggHeZlxOdw7k6GTOPMMQRK
oyvI57df7pNmELJqqgaO2FuX++wDpzQa2VCMv2efYDfv07p53nep3KbqVd+pXlje6HXWd/u2pxN3
Arf6TMrc8s8G8b+xLd5KX+3NmaDzR4yX6cDwhjVWIlSFGydpqK/umc9G569E0GQkzrMQzQY1sc4a
86Zl4T0FS4KpkaCK1Vn3uDSeYQhOqjF7KyjkMl88olT4LWpBUJ8orcZucXn/vp+z0o1cDV6KJs6d
y4CnmHkZnRWBCxw9NWxpbV0es6VCdXgomPvstpZorF9ogvWFxVuR6M6y8dLV8Z9SPPDlAXsEqwuj
H+TeX/6tXidTZdIMQpNT545uPKUEsrpeegrN99DHHpzoI9tayoD7NGZ3WN4yBsIKess/eWyLawll
TbuX7u2FJTdZNjuTWVg7BWOBxXr6/wzzJa02pwgzvG5qJSstJYC5OBlk6aABFKCAvOTiqypodA2J
WzKcBM+ucXWQ8idj1OwRLx0yMCGruxFcGTOYT0SJwn4alp76WKJRpzQD4EJl1P0f69qe8OhwiZfv
/donYg2Cy4KwPHYMQUdPthbRKHMQ00atFVcVuyP7T76Ls5knYMQq4J64NoRegnL/nNjzZC3Y6oZq
/qVOPE4NN6r06vPtGx/vHkqgQprEAKmKL9J5sPmF0RsOEX8ToU9HpfaB2urlddTILTnPFKIViEwS
49h8+Dfen6nA9I+prTm7XbV7HwWKyoogCr08NXu9BDstiOK+DoclySZC79WD9WXohLI1svDcT6il
WqDO5T3V1vUhfqOax2yxqhNAAqJ0WZrue8J5N+f4dOCufSZgr2VT5ztiZqGtSkok3F3mXTOUBPqz
o4dNlEo6dCfV/ILXtj4ClumjzWzEt9XOK7IHuZ3rf55mCds267xLiW3l+VA7SuvNg5NTSKGD3whK
2c3KIzJ3eKEV5KdQ/tM69RFUg8JNXhcGArOsNQkLCgDzLaaJfsBzQwfQ1NNwz1bTM3FnzP6OVHcl
0CXnye/aFzLohM+zJrSXWXmcNFpBgJtY1vTEhf3keIAsM2X4kRVfXkrcl85pncFxhz7DELVzi5kz
YmH2qMzxNQoBzQWGQdBzTJdl22APoX5VEb+VibRfqQUKhm6mO8z1yMDtLbIg0YnHOMTKUaUYu0EH
Xs82+6oAIEc4XGRSwVHC0ARfh4l4WMymLh9Hz5K7kP6IAnpVcT2tPSdWSKrLNdCPw7au1+yEVIcy
0nqEGu8ERr/DorazOJ+ZMObgfIeAIJOmSYuwh26chTfgVc+ddwwGYQeRP6a27BCPqlEUJqbgRkLL
fuiDf7yL0ovK4hYvxTRq80GRZReGLD36yKPyuiQllqtQMJSr7gSeuxoLxzrWUGEEMPGS7NZlzbXp
FWSht1gtzfVkN8z2genSn+dDvaHs3rYurM9/9xGbp5M15amjWAWu0s8deubS63gYl9FK4nDceFXZ
n0FGGWvUewpM2VcphkmdAsqujEMPeQHgu1Y0NegSXb6qYO5ATKc99IZGmDQ7UVQ1r/7H1/HMsc5f
lKbV5UYfkQSu3EmOvm0E3UmquWK59IbS0LFtVdi8We3TpAjGguyngpGfG7d9Ge1VNYh2EODwgajZ
lh4W5KlOX7g2+Cp5ss8zmzDfQdoWrCr+LGUk2bzVEUaKNuk7IUa/OD5P0u83d2aKXoBm7IW/TjD7
PxNQHpS/rd/FHz78eFUPu0DTH+XdiCmShiwIAY4QvnJLucRVQUh+K8KCp9+4k6lTPq6ys+vIlxcM
8NmsnaC3dUkDXgMuVWB5P+5TJ9sYj7vDp0CSRoATWnkcC5oM4O2OZnp3QlHTWR0dW92ByjsK6QGO
VwDcUAyWFMV6cqBNt4YvVaYLt8aw4qz0AGcG6Jswxy7Zir/D1cGrXJZwzPXA8SDFEXNhT3UFzVt+
z/SouLpx0OaKykFd1czWVKE70AhDmNl3J1VkAOndBnCHjOEozfWOcJDnMZDjibHdd6+WMPAjdpp3
zdECmaP2YbfQjv755DNRgOdg6RGZBFVbBMpJcthU8kdvRhRpMA2bJq6VhNh0l+/GOKjeN78Q9tF6
dW9Ov0BN7NVzzoPDyAiR2Jjhm1pjBeGJ97Op1/OOw+1VMi8bVgiTDTcb2gS8iwPlfoUdU/tu8/gc
PTxZjIFdstCzdBoul8/ehgsY7UsPqdP2CuEIUY4eZtR6PaFO0WUH0aQXixqhe93V+4sL7mTyTL36
kDrK2Zn2XUz12CCnwUZ0v5tKaDqfska9OlOmGis8ZdDxI6kMkyvZP8r1OckQWwBRLUYRfFqifABM
5qjPnL1rFQfyTgWksqwhOvYwBPc1WKpPR7qciGIzOv7zJJgChn1dpxO6GUDbIUxjlxc09QCnTAyF
vAJYEz0oK+9Ud+/8bwsWQWBNKxkUyf8FqO9EocdPRygrN8GUrucVuO+jS+gmYpb0h3rScuIoihd6
DucEoIaHGvzOqD/aesunnYYRKPkNzth2ekDqxK425aOsoh8KB4d29eNU24eN8VhnfvpnQnHAH6Eq
5IgsDVovHS9cgWLkd9yFlxhRvT1T6Gqv9FYURDRK6As//7HjL8ehZWGbbcpm90qtfI/gFc0WKfm9
/SXMCcxsaSYO6wnuMWD6TMf59vI5RDM0HyYdpY1mLR1N5qILwa/3tw8iJ7vuTaSJNnol8GHITh/T
rXJVapqw5xBM9B7WPCCWRZRMqF9maNyg673+98RTOxI7rG9m5bwuy8YOlFmx8IoVqtLSsq8Yab6n
9oMsluCfajQr9LpnGbtqeM7FVVkSGmIaWbUgI64ZSZrFbgxHJHBGn81F6dU5bE5piGUb2eXuOO8X
abeYgWknaBbq9VlDUs0igWrlxX4rWftzhMWckRzaxm0ju9kNg3zz2ufw9bHosHIgDmnclalUubxC
EIWJ+10ohRnSBjcDeUPWQGMPXq3XoRmqU5VYeZ6ANpYgg3VCcpQJEviOlL6ndbFJrHcDJCb66BiQ
5poQanzwawfeXJlpcGuhTATkmMCs1anLi+OUhmmNYGqhydjND3gzyRa2f/s/PYBeMXfWBkrb1nO0
/oVTHObyBVcjbl451XiXmI+Qf5P5sEj/eBd8JWCM4yvYY4zNiHMTsRvwOAKXHCerjtIInPF1DyNB
sKn+d2Iajuy6suCN4y/cdt/LDzbMWbGOXP9pYU34kYfL0Juq0qw7cZptyGlxTOnmdPluFhuQ9DJT
FwKyFo7G51DtxdDEwMJ/+HU8YxiyZWgT6upndeF3S0i3tbb0IdRWtie2dG5Aw5o78muoZRVkXYTE
UwJGrSHiGdgaqywVI2kfG77rI4/yUCZ7rD4y46VGK0r6ztRT0yqgQPQ4n7wgEZlJ1HKiGQuE2mJ6
1SHp4tkYYxbSXw2q1GGuLmLip3Ej8aYHDeqh1KBQd5dikBf6NkHnZy+peVUB0w1lbyNJ+5J4oAQ4
4EuZChse/lgs/R/PWOb+ieywULIqM3VPOcmqJ+njvnd08zDVozT+4uRyBTTmWoEp3Gl6hyQckYn1
hhWACpQFz1avdRvqXmizV020k89yfG4oauY7oj5d5qhh3hlIyYvf5AZ/Wiy6qpHoqbZfx662G/Oe
qA/gjcWQYSlYX3xcoOjacOS8Y6i9k8i+Ew25AlusLLFlKzZEoiIdzyAI5gzdG+n8hAhCbHYVGSAk
5F1PNdoy3fO029AJUR3Jd9MOmg8C9o9Ak7Br/N0Cf9qAYqJgfmVa47Dh78xlGUuxIh3749kSTQ5d
5tmHcFJ502BwcF5Hw1uod39S9S05k8xpSQt4aW33dpL84PayhvFTDmoZP1XHsKw7Y700gNUhZaK4
DXfD5gjoa2UcIe7C2/wUalGa1Fmp38M3e5K3N5yvykQovyLbZryvLaD6jW8QFKMBtKMqZ7vmklEY
2FdL1ISJLDkpcAXZwgFlenPt4rLoi4MoLetjolB3tDO4KYEuIahj0nveTbK5siZcyavJfYNg73Ai
uIA0kzWpAKn5+w7EeK83zB/4Y6rHDNTmNIj1qTFgDMqe13TMQkb5ZEP3xqxKoPceD7sn4G48FjFH
3cHctd+4+Mwb+0hdqbFjUdPP4+TOlCwo539kKqRJKT9Tr3VXJpSQQeVKL/jlEp/7oCyBaMV++PFp
OxI1xfDQa7x2qaTOLAVbVSzfv5XrPBZXGXWE1LPt7hQXDFJlooU0O17PauiTm/2s3JVGbIG3kNhf
gCRiQlV6VucaiVmL0UNc/JISJPXlQOmV9lVNDbwSg7GklPXASvq2xpYaGVPFPWyrajgm1RodcdT6
01lj6tlIvrQQ9Kw7yCD8fz0JPiQFpx4e2r8ZFdDKnPKITecu5ysbNYRWG9fXLIM3MJCzp7x4Y+ae
e65lt+8ffdd3QMBpGjn8LYTXXLzW9JyWmQPCH2s21qTejkzpAVvmo3ypccxsmtd7rIqUnTOX617t
a7E9iKero5GBrlL5MzhbfGKlxkY6fhEffHQvQA5CYY1ug648tXUiS+QKDluq/3bIonluKCAD/RmQ
hOVRk3eu6eeTxMRLnbEyehpY+R3FwGqSEHBrTjekP+O+C/ciOsBAd0lGEu2fgi7l9hy1T1pi+HDv
DuYTPCTOZdEWGSNo43eHk6mYO3ZgcLMy9F21vdNKLMVksGm2Ak8kHoagXrnQEHc9SyEzBpqxlKt/
Yk82lofoCZ7rHs/t86QP24A3cM7glqYW2OSg9AKxplHhvPNm8tNYiDh3dDo2EKQbYrivw0q1rs33
nNX2o5kYxCqU4ul5RLFfTJkNIEJpvtwxF28GUmadGKCz00nlVwBPHxSlvLJnxbVgJT77tp8R1G6d
PlGQP/OAivb5lnpA7EjKcXkiJEVLwwUeFdBDQauZr95q975/z3wtnruUCi5R3wIPTrTK9oAQx3CQ
QDiiNCKetbcjDrY/p2uKx65gMQNZ90ZJM7SAK7igrdkkvoBjFUgTpvn53/OmMHEv7o3jVcGvdUM/
61Ozeq1vtqBwXEzI+4mNnJe9plphyNX9pu0Zv/LtnUWOI+X4nBW58w30lIiOm6UdTxcFR2+1HqY7
xs4CaNmnqq9fPTfVDhWl3i+a2JdmMFBACp/pOTp/9Wuy+kXLZ+WGlbsQlrgtA8bBtG++JZIYVzPW
SttdXI/XTRW4i6TXdo3S8hAya+878UlWdRMpNYX/mnno5WQQRZqg+JCZUI+UX+CRQHUm8V0WG3pf
SujArWCQG9U1NfGWK3agJu9+92iFmiENFkWEZfWaSeCnQTf4QaJ1qYOA59Br40xCkFDvg1NWQ4Ew
hqkEyKeMKEnMlJ1G0/NTTu0xg6yflrV8o1UWZxHKFZw9miRzXinuO/5Ah8OclZHFPeCRa0JghSpQ
tHtM6e0bXhZhJm2VKk2VrDnihRns08XV2vOBBn+U9SM+/qx5Cl1b63phdtu+yt6UvmzKkGj6IVER
FT3A9n/GQaPLw0b6a83PEU+5+6A6YhLVbU20tjipbcQUsOFMxqCCdIWelh8M0OKk1F5ipWz07F6L
Jt2De6rDxkvFav+pKdSNAQmqmnAHnHlL6ayVx/IIkAgWqUfQvO2MtfTCDICh/dTlwIlUqWdcY1AQ
ZjkoL/Hq++uj70IU+iEKqDFAoW1X7cGAOvih5dxGoHzoOhLsLIbvZnABo3iGh/amGfYBHkwbbhFd
UL5dhKHZyLhQayQXeB2/++8LfHpboNadRxAzY/W5bA03FhYopPx8qmOrfv6Kv1QHfZH06ovtxvae
2Z3KFifMlfuEbBtF/ORce3uoVD9toBtyiYyBPVO/B1YfeoksjO/zLdaf2/ugDT64nOLOfewLglf1
JQCHHB+aTbXYeRuI9JknkM4jXv/fWZlSeYj2KGRi2cTv9+l7vG7s+FRw9lJLhFpWx1clBgwbI9B4
w7pclPB6aixM+F8lsuTZSBdmCPbdaVYUf2TACjX3exq4nHYkC/Epf7TgRMBcnn+itIcc+O2v7XIh
8BNSS+qyyIqjfNveRYZqD3Kzvhp39FQyCQnVETacbiHCpxfn3dTJtic9FLb/X9Sn+VMD2TSrt6Z+
whQuPFMaUY9Ycqmvbp1fQ2pclwCaz1oxwiVqEEY4JvFgLt5K8iDqcecRcM1uP6xQrgUGMLamDwwh
IQf63+yy18sNshaNhq/7S9XHJZDxrEJvMn1rKavlanbXfoNOgR963Lf+CmEkMzpTGXKlyZkwLjjT
zImQ4eb1wlNbrCafeWhpaWxPdczxezUt2fNrXRfjIopZ6u88ScVZrkRIG2nhytkiW2XkxwwgJqvj
m3cGqg6x5CJQoZhUcrFLLw+rNG6Kkk+GKukVNeSufPWvZxPzC010V9BNv5jRDjy70erLmuKSwKD/
C52Qco/Rpw4r5q+IFKY7BEhp8mVL1pF3PefvorD31ogBzxgB4In2EftqFyuFyDYw4bMF+fFZRUqF
Jj6rETJdN5uke/8afIJhSdmnjXPFycUcy3yMfyqiL5HtxHxHu1YUuqFQp2gkB6+Py8cyDkbjy2sg
DqEgFPLDCRYH5yvSZdUx0DTyBWdxnSd2ID63klO+LaDRFR4WMH0jVuYHJmE1opdkzT49xAVtewZ1
WU2RLnQBwOYrZDCA/CPrK5/tEaMe7y3cILfgAd/ZXTCJ2zIGs4GOBBWHr7bmfXtU2+kWgp4BuKVt
1hG8+1/Me2XGQBTfBttRHhOy+0Lx2Uxmm2daiedtMGOI0LxNSnxePwg2dWidZCBo9xSRERCtAyp0
YEF4bnKk/w9aiOIFaYgoIaap6Zej5i+x+/GozVYSwIgijF5dmmgi7WYLf/QomoFTd6PM5+DB+vgr
3dOFD89zAb/mStTXpkHLbONKoI8sJ1eo9kTpo4O0G8ra0Kj8GrGMwgvlJWjJRcyyS0SY4hDK5Wfi
EAJp2Pv86RzwnozCthnFlHTVJtURb1DJyLaGumZog/SvRKq2xyvM74IxJGMTWVHxXaq96hLVSwCW
ef5nv16gc2ZWUoF+tTG+gzG8n0TAM1/u3opkyhB1OcLAVAAcTZxFAQ3iRPWJS30l08wrhXULd10g
xABsFBvEF5Yo697YW57CmLPXl+XHOZyws0JUGb5uSUMNBReMIuJ0LGhAV7WOn3p526M7YNc5TAig
6FaXDqPOCSgxGy2MtCW39wuUJ2+dBLaHciao0pSJR7TlvahgkYw8XYGpYizEKJ522Xj0R8BcxuIr
s9XzEb3NTmgv/CZcUAJM24e5MZrjzrzbJNxoCa7P3SqgwPk+8Ic6f8SclOT4CdwnGN+DWGbvnhes
HxF+/FL9/CujjxIZ2MxjqeW2mf85M6DMg7TsmjM8zgxqJf2pZtzrbO1A+Y7oPsts6FP6DQmhGT1B
AdJvQXvNqD7D6f9D/i4IdgVcBpvTXc3y3y5PGKb5CMIGDPQ3GpwJMddIUWZOqTESQXl4h72mHL7M
cx3EgdX1QgI8aN8vjUZorzkBglAv6yqNd0SpnoMTcj6tjZWD7cMJV1z/4SHgLUKFsKrx6Tu2QNpt
jzCgU2wFhZX+HeX31mFUgd8W29XVQhthuSE0MhaPzqzcCCRF5DX6MCjoqiCJSgHDREJMN1pgOt3u
PayKmLm1hpV/DJom+C/tIwX9yv1MPx9u8cfEqMVDqafatNAuoAnV5fnPJSLzYgU+t3GwwhYtR/eB
W3hQLa3U+4HX+JhNos15BT76eaid6gBSxAUoAS1OLAlmhtFQxfgqNcD2JI3h9yu5z3ArMahLadIF
oBbnwo8+PZfIweJyw8EqnXI3048LqumJZD1ILiotxx6w6oKDlmrrWLN15bIfuvMtzKkucEqvb5yr
PuVjXcnFUe1qGPsxdsBQvIniGwLcgPatNMcFNkkidOuOvZEDzsO5FGMGQnpGgNO5SNm+erq2AL03
ir86fPyQNfVZaZ3QYWwKKprqdhMPsRofRxwKxl6uoT/N2KGTfNNw1kPWrxPafEnqsxd/Vzgc379r
2lWv/6bFx5shDPWpctqYo95/dxk8boBrhv3ko/PWp6D7yqQEFgByEGQBnTTI0jmnEo4f5EEeVEq6
+gIwv/QNEBG4V/gCQmKji/YFQR5k+N1XjUL3opd7fhKfqLepxqSxyYm2XNb/a+Z3jVk8TTZF6Gtx
Vnmdrw1k9DM2HQErSGextch2br0bNlp4pkmJD+ifK/iUAXd5nc7CkHTacKUJMc1eD2qwLeL8u7HX
W3dyBTH3pQSTPQSVhY1EPGTiiWdfugSSOQpL+whjKbPjzjLdj5QQaqK+EaRY9mM3NBF9UMNq4qVJ
9wlXjXn84GbkhTEtQAgH/n464+dfoAaWk39h9774bsmMoMuQnMOQoiSu1KJiI8/U3JhIRiGuSx4T
a73Tj9cIq69F2UnUiF+oo8HhUrOVcTOgZIkyylf9bdCRUIug2SnNl7YK2wyyXNe6RAe8HTs1pyRq
I9fSAg2NNFF+AU8axjwdtv2pn+SgjqYCpgqAVVm/UPqCgphUGjgwpViNYtzoXRlIVXl7fnUoHO2i
4kIsIfahCYZHnMiVqt5UaviBDeE66MDApClwkERNcUMXnRFw6LJBDJa9UXJwFAqRwItXsCit7kRF
ysbxug3ozW8Kvap7txmV+SDzCU6h//O+TkU4WhmndRlTK2uNWmO5aO/zCvIiEEADNTeopd/IZRMJ
NuMksMt42K/lqs94Vn9i6wBJ+NvAll9TR74jlKayqdfXOQBzwEMVgvrj6nXzmQdUc0czFHHm8et9
O9tGawVHF9jNE/dS/3D5ye0XJSTb66ctyWDtdu//bk54Gsxai8asd4385KH0GABu/EyPsZu/CGHV
3CDcI4CZvhsn8uFWYx2xPhjOWn+FxUeuk26kY+i+Ver2eP58eCyoDlQyhgydn+HyaEXRhbJ+zp6V
ATDig+l5JD46YkqqM67nimvDmjLPx0L6XCQmHJydMYKNEcsQneyz5+6S/VFlgn1Fc4bNCDQDdXw2
lYpRUx92zsuVM1N25e4pWvziTz4Vd/HKq1zqb0RnR15Y8eATenajjXOkhad0KDkRV9sN2KALJV/g
ZjWL2QfB8aqmYv2SqBSW03wEJhhusa7WKKm4LmslDXfR4TB/Xei3oYNkawgrUof2/Kxvf1EPFybD
ngq3W+Lc/pZX6QJpX8b+6+TtAy+vzzdIUbKfWXqT/2+h4auqd6+hrEuLlLU+SKqEmLPZLHziPXow
c5t0zP18LUhwhhg+g7221m4spbtwDktcYCBW+S+DFQMM1dhzCJVchRjunMwPhTwaDkfbggvucjIm
cnBoTox8XiQvWKEY2uIMcyKO1Q1ezEClxyAV/5AQmT529RZu4PZXIZ0XSmMGc74K1SuECvtVDYL9
RUDjPGQG3yzpWTElNBteTwgCsXl3EZDthKXNYnwBHWI6tVZmz4mkHY4kOl4OC9JpDeZKH6gRaOxU
SDsyAY4fs0VU2y3z8kn33l+kIB6aLEX3TjEpofNGQB+3upytvKnr9gBnwmGUgur7QQvEG4sxL7zD
WIeVlG7P+fAsN/l03sBIG2mu/njPKo5vAbI/8z4ZGTCDvfo7nNOBaCIcck5nR4gYD+TlawbDax/O
3iwh7KU6rfOW2wQbaXfgp8eokrRyu3oBTrxiYQgtqeTRE7lrkxN601E3HEGxWNln+fUOho43bAW0
cnyAWyEo79ofLi2LqfclflZM00+PfXtfHR7Cj+pNFh1gIrza3yr/+U73HJQDjD1l+Yx+arOHWJRM
a/ME7ZhAw+fckWl4jsRmUB28tO+IZunjO0nwrT5juSEUWtfccCqg/hzY+Lz/lUu65nFHsaSf/QRF
ejDRw9BBMPo0kghhz8LNmU1LqKXpkA/58/3ohPUM/ISqbdb+JSRC2MHkvoXm4eoOZIA+hu5xX0SC
8AEQSzO2kg5Gbk46QrsG1Oin4beJBcOvH7r1wwy8SRhk0Pg1xtNPaPfyMfL53NDAI9gkLTG5132+
wcQFA3QgcscrLOKIuhko7x2bBbSE0fyLM05nKz+ftD5/aTGJxbr0edBUYcieyM9ECZ2cfRYNiV/x
Eg7YqmQx47/cKtniPGCytESL7Dpi28uIJMGSJ2qusy1WAz5Y9bgxiDE0I3V2hsECtAaNOms/M0jK
REehGxnC6T/MbsHO3agA9n2JLMhw5Kc8e7ZRB2FG7HCkKW5UxVO/28nGGtE5Qzu/oqBnONr3MdQ9
F4ktG/wfcOBsLG8zGs1sN7LBdg+vDzcORf9oBTAZcJr3tgmE3agfyWg9DeTzlPReh4GPJ8RCmB9C
6+lhGhZQu8/1je49sWsSYyrSUP0ZYopzGXPSsHporxQMJBctmu/k628mHGOFLL+Ch2XRQgCs90ZS
pNK0zlM74o9z12fpsX+HUPvBmW/WhV60gMFIa7raf2U+KCzqtUUuHYIcV3yQ6KxbqcGHBJDu46+X
+Jg3yx+zrMtpg10qVja5KkoXpa2svV4ycG/3g4jJzSfXoXTzxpM4EB9XaBnGWkyJD6YRPIYFvxm9
quLVVQNdAcGChYPIu+FLzdBfKwO8e7/bu7UUOMGNFMxQ0rskEGceTR7jO/2gGrN1fDcYf8q4UI9G
D7r2Es89RPQwFM4zOoE4xiqyRmKvdnFMNUdnf9I5JgBI5+TsDtDSjxR99cWjcoPzsosN/DdX0NQe
FTS6lrm1MEHub0TQ95hiyJ63iq49ZXwsXg6q0K4IhYlFmXTz4uK7522luHhqrfuJ7/XF/lus0tpM
MpZU2031kBrfGu9Mqgv+1UenTsh4WM98Se0TdUm5p9Bn5ibFTcdK794v1BgBOqijTPEto+OA0122
+jkUu0OpFpPjDAbyQD35nxX9hgMGvcatnvtCwKYmSbk9kSMKUZVogSlMFqxUe75UFMuWYNdg48QI
Szgvar+QVteoPAhywO/LXxRxrWiQHyeahALxUXGqXpDsHZCZUBVGyOMMg9agkGU1MWsfX+50NF+n
GOmTnW1i5yd/E74dphAOvPJaQQKUqOFPDo1Ku3GrN9Dz9tMbS4sCH8LiAhz6umjnQUHA2e5MDoSW
aF0FFJ50UfCl7fzoPKiEVkcYuEseBrBy9J3RgEVdOCyioHAaxdN9LzWaKqx/GtGHzQB3toKJgeNO
lwTlGMS0Ba4GQs1PuoegmxfaJglJVdTi3mN/yMJUdItD6hDI2OHGTf5k6aEKgLj7YxRGXl/uwULw
38T2QCSckomVrCmy6EZMMZfcYReHf13Comr9YDjwUkFxBBVB1ExXCasSl+7sfG5zXzOAwSrLBrwW
1yz+dpp3XS/jVvI06bDkV72FYCdHhm0iOgd7fqbGjwCKCyJX3F7YLXPXCHA19vATKV3p6StoAUrI
IX3Zmep6stA7oPxZ3l+OJX1+wKDrUAUG1zz9DwMQ/ONrFXg4fXoYILIVaRgG38BPN5j1OqlWp1qZ
K6CqdWU0bLKn3Be9Ir9hyBmljpgYCk2+cinx2D8dZIRYnv1sPRddLE4cUJobTvswOP2adZABC1O4
zz6P6L8LVWuRzxqC40myE5V9ycLhYgiLOo1GBmX0dn0JmkXuwIelDmmqO22vEK+X9mKiVuUAJECf
rIzk8JlPTmX86hsjdAJ76lpMKCG953q79fqGI5zm6HFv6uqLfG93fYimDzvtEZSoPzX/txwXd95H
D99Q+VSxt7jzpKzQSPrfRyaZeAE9rE/BnJ2LkJ2ddqJuUHVaHhot11cZ9QxCKam5Tlk3FK4dul3h
y+E2eMrd+UWrP66LxCB6thKxVITb50YJ8zjz8IKF7gVuzgejAKZAjH7BbQiaKPDUuBPKukPwH3Mu
x/0TaQvwZvsMTBXNVFYFsF5fFdDEhqlwOijnQBrJDR9MgOFHKs1klzlfkR6MX5+lmnNK7WnTqByn
3vNcV6yKcT/bkukxCnIphxr+NQ0ZpsNiTYX1q6b+WdMYxkABnPsdoZofTCe58YWyc0ZZD2ucYBnf
ovwtPQlTB1DATpb+gvs8MFPoh+O/IQMJXPNqguIcT1lg2e6X9qNH21FmdHab2n4sAi0UjisxqzgN
FXb4PI+Wmw3ajAjRoXZwtO5+B86ibqh0vJX+VW7Fq1NsYNudbEWVoTMir9dSvHBJapufvb8VNgr9
p9wwY48EAkpfHzrHG/jR1X3WqKg9q0oftzEDgWRFk23KP2qzK882MudORCjrV8PEJkunBLjQ8+xX
h4Ud9hkkYCN+O7DgmxOYx61RiFyVl+SbtjzMFKTGtz01H4Rtpb2oWbK0SdvnEny2wbBrmz/7jFKx
ptmL0S4x9RJJncEcXxO4L7P8kPe+dC36HexJk09dGIUo3aVHeg3V+JQfo6PZlfJTnDL2n9Gyssx8
r23KXX7yKiDJ8n1qdzOxKXuL69zlnWuq+JJD/SV7OkdJAg+spR3FYKIOWeJ2+6s9gJPDorw2xWm5
CCd6DeKNrabgJdLKhy6LTNEs2cyKqO6BgUjuoQ9b1EZY/n39MBK+h9GGdIM19AXYFHWvLGpc9tbh
L1QbxJoXsSwspGfruFXnyNKFrsmyzgynKmfztn4tSFJMXYKcy2WAiqS0Fl2xUljK62w0fOT1gZ+0
D2N+fhhXm5eRAdfe6B/gcLs3YvHWgLHc8YyTrlUu6APABMER6PCJmO5EuGmXYpkswbP637I9ExnI
I46OYcPHmna33RcOl+vA4DXvO4+SZCxYyxCpnlHkwbQPE+apoQu7ZyTW9ksDOJW4UHwRgQ/TT6g4
VN2Bxm11pQWeTIOpHAdMzE1IyKRCg1i6h0IgNvqztAlKOHakN5k/TqCYK66/+0ZvKW94du9gi6fR
kgnNziZbZ9/547wmGlpHlfcONB8hq6BtpxVaKfRbS45Ohajt7SbICPVJp+rxNg3PzpE/mXjiIG/Z
50NlJ9zAw030O0+75Ozwh4Wq14Mlf5T/9vdFEbUzjbd/mD7e8zL+l1/g2QCh984nviQ9WadgPvP8
Mw8mOGVD3ALQL9yOjJPoASvWLUiSCFM+jINeIWlaN2Ez6/rWh3Qpqqh3Jzog4LbdL5kqStKt1Ae9
fg1a63DCreMe0+2TK8uU5ZDpIrc5rbUoTn/5pyOymNTXmI7EZRYSfTeFXg2BSLYlaKXkZPp2B27G
sf4VvGrXKy/OX48nKyNwuu1R6sknyIo26T7ewwBVzmPFTuSOKyhljExNegwbmgON9LnX/UXfFou8
wT/tvX9YW7BQzWawjul2h2g1sUfgKpSDQtOyjA4bKlLesHYPwjK/JjH1rQPsjgQ42YNrQOHy/6GD
FQK8df6obfA5FRr5VYR6TQFlrvtW9H48PHMTYhvsg9x+f7DC2Od05MtOfsUZ5rPPgOBrtQlRjCg+
RpxBDOFvLFINBL67j24tXeVCH5D+Yh3e4bk5c8yopSotADpcwvPZc2rf3tkMykRbllAoduh1J4eF
NtOpiDEfhuMfXu88qIPS7oSiRqJ/Sgek9/sLiC3L9fs/KWt5VC2mLh47TbDlsrkFpHPsaB/PYi2V
Ve1PNyYAo8oZTDbaHJaSowx41OAWJoFo2CdxFWfZstOcHjs3p6FPcz/Yn8Eu+LvzdesaOwuzAHGv
LKaZruCt04G5NJMbWAQobo3L6AUMcqw9gaBkwUHZNlrHdalEmi9NJrpQuxDhvW1jr8sSMBqa1LEa
teEN/JWn8qAYxmA58S8pp8aqC/cVMyqBnmZr7FUIk3cjnlzhN2U8xWgYNfWed95exLeIoojRuQtx
ECMI/nYHIzJFT/QqkCk9m9WGKTLRTnIFk5OwRC+YMt+hIoOLZzYlIu8V80ocMHed5OKREwbp0ArD
jCt2yW6zFbYOyq9abkV7XRbCivSKdhmahB8cDBJg2bfWiA8sj6J+IFQdSNVy2/znggu/g5VmF6tJ
iBTKpUUopeFLmeSwE7137USUuMGkCsgiRnOPPZ316VSL1K79fnHavJZceUJ2azHp1mX261UwOSzL
wafV5SCfz+dFSMb1IvoF+T5iym8sSVQJLzNFwPoyLFKjXUB9HmGg8Bkm3r1SPZ1upzqiFFynqfL4
UlaC8ECmdNcxV6Nphy8mD7XXAjpDVE70OenVE/L+mGmdZEoBw6z4wkcYFGLfIXWqFKLb2UKvcGX9
0CunCc5QxOWs7d1+xyQshEgLl3RaS5Mhih9Gy9x+PY6CJqEsc2Vvw2ZcWGafsl83Tdog0EDV+S1x
Donthj1RwyabWro8+LZjEqlXfmoAjxkn0YGutyVBmsSt/vgxJUNGchVFmOMIf9wtwQj2PDtbxPFJ
a//VjbImMq7UcFy1zF3obodenT4b9BM7beiaghv2DIHMQIHq6XsNRtyD6jr+s+0DGgL8T0DRkEiN
oNpFmnF+5z0IbrwdRZ/7zJjDhv3Sxn1r01+TZOLr/Td7v+xCZeAnDfOW8mVrb13yPwHrFDhIlTMF
XSnZ9V36srWiDcWVOvFfZfHbtBhSS9J7202eGquCEz7FRs1OQs2RdYtgzxLyEiSj/iA4QKMD8KSf
NXynjrvFcjL2xi1O5yX/4eFRujeCbvTXksV0Q2Nc0LgI3NUU+dxqfJRxmPyQXi6PbYgxHyu+31dB
M+e2ZngHaxYip2xM7xWoZgBS8qnHx1Kp9H5aHV40KEB4n1DqUebppghjJKUEFLiyUkzd685D+xfX
RnryxQvub3MhCXrYQRTqp4t5+TvbOeKKuZolrN0QerfTctzttc7j0o9dVsUWeEtbOKED9dEqTM4d
PBh1rKtdZdZMX8XfmChx4VdQA7XpphbG0YQ+9ArRi8ELiR1g4j512Vho2EUDweaYMw1SooOr+I7x
iFcPCyxAReXChKYbTZ38D4V1BnoXFEgcINclUmC2h70pdECufUOcGNm2AKMkcGJqUm0p3/BarYbt
ZUKjHuS8ROe8doVYeB4FZlfKV1k5bSweJOgieAJCoDZr419HyGmQxIW/V+ikbllG1JY7f16GwhoC
yIIDMWndzOOctpAP/6XePXTH28LPbMOWSPX+ewPWDTqNo2CwbbAdqYWpswf0jBjyXUGXZAkaA6cf
/hHU8Z8LQN8na04ocNFx9suKaGmCprJcXgD2Klk3ULobma+MovCUahA9yNViFOfAYt9UbWe/PBeR
IMTlibMRCjzu27HrlHttHBGeK1E6vpRMK81HS9+angfInFUanLB1lwmT1lXjEqSyWaYV/AwLkpPf
RGSHZj4u5V4MoXPipyy5bj3d3itPNl0i0ViRRh4xKnjNHTcLx1Z5f3tQoO6C3IH4DgVqgTpAZFSZ
rhb/AARfndqHSGs5Gvsev+dvWpAaas8NV2Bn81d8QK+weL8sMbc+tqLogn/XftkQZijFX42V53Gz
4LPtpW/OhCYr2LFBY293An3OORes3kvLSkjQG1PfNgZHcS4eH5ivz/y5WcjW138EZmFeS/jsJV1d
VzAC/sHfANSLauJ5VAhvwtgrngnqn9XhdNbdvjdogMkTiPEMQnu6FAFpVHYmRKbwaD1R/H8O2S+9
hf9ELx1Zuy5ti01k2UCuUXZKeYlu0G4qaK8baHP+pGUdc0oeYYzj0b9qDzPOyGGOnyOUoMGOVUkg
to1u7Pn2J4iGy+3DfK7H9xFOLhTMcXz2X7frWUZvWaQJHZZxDU3/oGxktnfyBe2UvpEs+Rypeht3
9AFa4Wks78hRabd7eev/2q/NsTA5/xao06wZ+DMPVCJfd85UirpGSUYqtUJvNaiSDGhX1QgP5QjA
LmHkdDrlrPwuYXpbsuyLcXdsNN6LOvQqXQ6cm+0/4Sc4Nmpa03T3Et98zPW1KJvUbWWB01bPW885
TLeNfM3v0z21kyQ79T7pjxnRU04ayaTBPg8JVgZlQRSCDmSLYduHV5QYoeuAYjj7o7TYLrT19onV
49JJEmzg5XbsJy3hvCPWRcpDbKwop8hKAl1l7n3m/3FR2wExuxbFlHmc/SRQGKt7J2r4tihRpOYe
JPsJurb+mjLqwm1asjykBdXlNvn8gt2PalxGJrSZrcJurcRzsct0Hd3mSxGPaHG0w3mvAjnaMk/i
GhxyCFLgr/RgZ3VkryI/Q+Gakvt8hDcyBwVFf+WVdAUU585Qr/DkmXSevjWbYlgN5Ls30kCCcSuS
OWECEnrHqzUWFVBBLiaw2K116oJ2EPxSu+C2UdffHTu85yiExh7lNeoJDKCE/0ZWC9uorcfXNkfO
NiyCAZFFIGmf6ERyeqp5VVmTwyBjPNf6SK+wka+r1pEQqVNUSxWzMQPE9TaR8MKwn6aZAPa69GCD
9Ivs0VeqKVKXOdAGgjhp3VZRH3gCt+Yx3U7PL2wMd5zVstckcyeDcAZzyu7GwXbByua1BXn8UHWL
33k9kx6V24MMR8zJy0wvSnrS8SODZZdaIYqFElqmpr4g7RTV1Nx08WDibXm1LHaXhmg4uZpJT4R/
8+Hmlr2pwVjz122x1Ij2jL/zys1qHHPnom/AQepzZ1jgKcclksYLe0JEnAgln0I4zE+V3ev00LSj
BAfwH852FkUyQSSrZvdObbRyHjX7sqEYg4MzDbTCV2UgF9l0Plk+6BzQD/NUv5G8WVzTbhrUdjpK
s6ZC5BbwkNmlL1ue9u7D4DJwvz3yndo4nhbr2dltNFC3GwrH4pVDdWmXHSLRvBrD5TzW3P04hujM
6hlxFkkSVm0h5t7zAnXlBuCbUn1ApepCga1QP6QmAs/2elAipt49HAyxFQqQVYXkkGA196aQ4pVw
GuOShLM7bYO7mTbBdtDQGCMST23dE3gjaJhMl7gU2PK4wu1fMkQgIn4aq5RHptqC2Z9TUICdw1u9
JzlajzoglHe/xer2fM8zZn7nDmUBr16zo3rA4S96l/SNdLAvHJZCTmuROGG4600cIiNB2udzvsZv
IK6K71a4QbwlnofsaU9yMMxnZKoG1PeZkk2xSBWymzQBKtuZ+/RjZddo5hjRQ1a0uxYMcOScQbgm
PK37dTJXJ5o5B6ytH1oK092321wTeoavbhjj/HOmh1tsi/NPPutX4Sx5471mQqN568AKx8hez43r
B/BkXxZjLmLPE5YTclusiNMHZEbxT4gm73g3pd/wZuft3st9/B80zMCnVwmNQi7bw5Dgvf9tvqrW
UwrSUQT+1mBulYUJ9/nUIGFZkmKrEpqM8oup1vmFDUnfhLVvtu7WZyfPB6SXPV76lKkf+6Mht1JP
sliIDQGFexp+QVKMwiVedl6SqTTc23Ze5+cA4H5rl5PQaKSzZz/VykkNPaNsjobwBSSxsGPI7zIS
qQlm53iXQFP+gmgdeXEo4MzNbv5aXtCxzwe5/LnKQuXY0w9xIFirpPgn5Ey/gx6bgXRxx90Qey99
fJnD4UY8wmUuK5VhV4gtWLSyOmf1Sk2xcPCMScY/fL9ghC8N08HjBrBLL4DYmU1q3Lo92aiE3vJ5
w76/4fJZZja4klHCDdqDXaqJr7mmjeTV76/QDoxiKw/SZ7WzDJn2XAYH1CzzIzSxpEk1uMPu3aGM
plt8aeMz7mBq4p8euNiM0GuLn3fsvZCsuP4FOZUCN4r1prrakVtiA6zCDGDydCxUQUXkvPtKBXJR
Sbl35wo5GoQVHqqpCZt7Uw5JLCbHSNbN/xTDg3BI901zZxAFY/qK3p2/YkWLBrA0Ojd8HDZVboKL
31+mIHDq5GNy33ovfL9/wDdQQE9SDIGkNawItIDvs4qg1bYwMKQQFC5Ol1GjZDxXPKu80DgOcm0o
pv+raGzmGOnJcd7M9DqlyJaoT4W6GTgvPXVcQwaxc6FYcb7ZHhsV76Mead36DRlb9R/gQsd2UZv6
583WpFgPEnPAtVfikiGQvX49RKEmeY2ZUXNBdwBe/vLxh46jro/l7w6TPWW9X4F/w61cVjD8GLAT
YIHfmgmYhFZkWGcIfIdmGQKsMM8TxhBDh9u9IS0Ri1sW+4XodSs23txqpzyOHluLpO0jMlQrNeGe
/5hUPF837Llu6N132j0DhZDOwB+2/m7B942v87cew3iAKQnVer8vP+NvsiSOHiay18O3cWrP/dXO
T1aS23SL193mYgkDXThz+M6wZDbx7po7gkjs9EfghDgtXDe3ahBMGEG+hwhwFBh+D4TFA8OYYGnx
uVuuz+DnpNPUx7DAl8jglPCY+yi8bvp/ELK/D8J2rVE7GHGoRtFXEh5eFzeapMPeZm33AERPGFnR
2lqkZKiqZy3k8Wm2+Mzi7miKjZuq0YrsSxhr3vlYWOuqUYfVsSBcOZ86GYwy92IzXjVGmCCcT+9+
hqQvgz6/CZe9mcwzZpee9b0n0y0RaVY/ZbPc/XFxNcOIYGE0vAMEHHCkDrQUhG9j0TINzYcLxHtL
ExrFFbmYukB793HctyKaxfTglSH9nwB3n/wrDPgDDqfNEGltaWKqzwM9L6pcCGeQZVqYmKPmzh2V
oRltnqOJQ/Ta9ZRO3P0KV2PbcqKHK8GcIQ4aouy9jBBmliUaX0yjWYCQJz4fECN1dSoFBOOyO2nN
+qDdumlLt4YMQZUNBvN37uLplf0wT6chpyuQGqDOrw+5A3Y/HqItZIpr9iGxbdLm+dchyYGYnEO1
vi5V7SpoKn6iQNA41tY3/wcpHxcSWQPah0cENWstuWm39y22nZ/2i4P0ihxhyCeG/Ttl2YogATYo
Gl4slDKDa2GuhMbXIZZI53PYw9+gkWcGLroFxYM6pCcvEJmamYxZHf4mtRvIsbNDZaVrwxX1XwKi
NVNU1HtNLwRp/GVTqVZGWRtmL/D6/HpylA7Z+R689akgwAkeGnJn62YB1B90S0E9MsnLLnNy9ebD
v2Ug8TnAeiDYbhywmEESBfkTrbaM6NhmLQoCMHkEhVgO+jZZPks7JdovXIEX2SocnTCLWTB1ZRy/
9vokoVfg+RJ4RHFQxH8jPZWjvwCJXP9PtW3pmxNDQ63B3uH2ykMRogLDS7VMk/Yf9aHjOcX0MVRj
jx5ySr+/WTXfO98vrJPvwxxTlSdpLeS4HVxzanywIpmCBYk7nuoDxmYOqvlfEFYiKhlJ5hWt3tUc
TQnlFWYWZAkhevvF51yIKI7QHU2GjhS1Yz9eSlagffggSEDaAkYmXwq2ZKy2zQI7ifpW6w9eJFki
v7S1/hbA/y36LM7wmK0dxEtm884mtftv5vB4D882rVupTDCrx43Ys9NW4o5ywcjcEvqSa7LblSxF
TUHxD50bU7WLrwUE2NaCVAe3U97iZirjHlrlqWdFhPfKk7N2bMdhf2/bZeay8Vvm9UdvXcH33IkY
WJvpZlcxyrurrNJ9yf0cNUdptuH57QM0whd79dBhDXaK5HVw6GP16DdfiI0CLDGhmcT+WprJJPns
IDmOj8dCtWnzWqX2fwdiPNVydtO5mcx7lDBAbPIvO0H5s9NhRtmQSiCzXp4Lb/CMRJuiD4JJ9RD3
tecD+iH93zIYRv7JsabhHUikHiN88eRjzhzuG9wbvYQuWcwVLdU3kUjYUdcRsb7CBE9FSQi+Lo2N
XNYq0Qcj0ZWHMoPhczL7It7BNTR+UmW+5AAxfB5us3SYwRxasTGu2TIU+wANlLgMNkO+/EBB6sW9
IxUaq5w3jv9oA53FQs3xDXZ7AEiT4TGkZc7zTRzayO+Lo2hNWISgN7JU+AzsE5a7pELLUFx82mBb
MWCBRIriD+xtCPDX+pA9OMBkDf6uT0fErzqzXOJaFRZ1ZnN1ZXdFSpkMDzpFi46LDHAsbYvTQESv
B5Z+aiJSpmItY4eDATS+BrsXK+v1ZCO5J8ihcIQl99x9dVCWDfqsJ1MPgRmYRYKseXT7qzVDtfdl
UQi+j9ckoIej3YnrSHVVri+qzISm9H8IzL1Jea/cTg/9UVSkk4iFHApvCNYHjNsWV27Bs63HEh7W
fNaHHe0ke5NV1KGN8su7CPscSLMGyCJLorQmHiSOj742qvkUxt9sM/jDOCYspxr1PVnXuQvDFXER
jzgg0AFK8CHRNNzuiYfimtj8l5ONnqsS6GL+CcWzerRCkpdtUt8ZGdVg01ExNaBJWVCZjZi653c8
ukNXiANF6tzxQfU5zPgmHbvCUBxUIyRvQ47Q4aMzFCa/gS6O+I7w3kxHBAPu792/DV13YCRIUFIy
i/LWBnDs54eVr9VkUMnN/fv0cEduxAcZf8zGO/ukFAPxgrUzWesNbYUs3m+EaTFf5TN3YyN5qVtA
Z/MT3z+naQyG5B5Uy4mtw+KN1gSL/Jz7NtjXi7CspId+19mVbb5NDDp+pe531YLl2Hz0breXEtUy
DhWZ8XPqqV+1MgygmMxq0F9SMkh0AVmvQ+BrUx9MH3eEu/7DdvWZpJQIVYKBauBL0B0dInC5JBoA
/V3R1u4zxj+Ru3pMvTd/wRXR8OkmqJ61FOkUXAcdy8FB1azoZJOWwtA73EsynWDv/5tI1TSfLLDm
+KAG0c+xUlrCSOf1aXd0U5n9tVPK8km1qzzPe32swODton6jG9/4OZGOoxRI5sAzpx1CjXOOEhpP
aOGwwKyqqTqJ3di2rJKFUK/77//zI/cexRtDZLu1mg17TTmbwaDAfNIHG3j9JLDVzLfqMiDTtiPT
yjjjkN2pXpcYvEObD2AbO8lCYtKeVkRYVD2dMkg0S8HaAIrzyRsJAuM1m2g8Y0a0+WaxrIn3SiIR
Mk4leSFRWCg85kdGOHqQHkzM8cZNxTwsueKtZv1xHrpOryMgx213JLi2JgRdtneFvyGdfiCTPYXn
ZDua26h5YrfycJ0BnIpH0MvcY0WjWtX8pTro4E2o5dpKG4YNFZXCtQxUI4JTq2+bRcLU11idQ1wh
rciO/lb5Uff3xazzrfRpE9tlPtoazMmZD5gFTrhIGPp5fCroOGvPCwm0YtS+fiwhZWHEK3bCdUx+
svWNbXlpcKSw1N5cWxkn7EueEf0WBDxCmPc6LjL1eqhSromqxHc7yFNAmi43/BnJZQ5GUVV8u3bK
FPEKDwdWVL0LTLaE8OHiyMn8WqZkW1nyQjF14SSHSkEHlwaUZMjwBvPncPMUgftf5LBL6jVLxGta
yptIkQhSj5+5MFkqw5zBthnGqmiBM/M3RTaEuevF4rn1aCh1tmGW6N7HaQX00PumsOZJIeWKh8f4
zvcTXgEAm8MYxXVFD27Knt1M0Vr1kZeh9N3FFh1M08M4gYcaBoN5jgrv9Xy3iGAjAU2OFA8ZBigt
i765BXhUiJvE/ux9c58Rr/5ZyKM8kMlCqbtjm80EuKok9vK0dyUWSvc4rKLxU2hw1GeUnr5k/Qen
yUbFBz5WtQYkEg+jjWOkXe/tKGoYj3UmymViwdENi+L4kbbpwIxko5ZR6zr9tg7Xq9q93n88xYpR
2Buo30IT9iBtsssv6VzS1a0EMyaWKj8FMTdMRuiVG66CpNdYD5QVRbQ1ZOxYd8AAv6zwoCljTuCn
AuXbbSVu2/3Bf+PMpksWsP59/nQG8I3KKCBVhgBBtmyP4f4g7ZJBVl5U21MDof85EcZc3GGTOBRj
JsE2KKMPfKP3olmXf5ll6sApFEghgqOCC3Dt+JGxbX2n4pLtu5Nogpocqg2PkDt0oH6pKFObKM9H
6DQbN8/PXi5dMypG2PeSGHj3s2dkRso4395NMpQXUqWhaPg65ZgiIXGnsP+cV+NKpGNtaPQT53Sw
f/KiqQyVph1pdJte465yoVz+MGraywXjTVYMpcmH2pWn9xtzaN90Fllbi9Z05tNbFBKl8+DoEA8H
YC0peuH4tY7AymjVmuVzJOICNCCjvI1JavrVXqpX49TNPLUbihknwSzwJmE6Ho2oLB/LPrmTc+A/
/sCxtrw37Umh5iZD+WN1cOOFMedC5TfOtypRhcdlAVa0aJM9ESVp0PWmgvn6IOTD2c0VTbKxq7hB
QGaWQB9pSrTaZgt1p/sw6GTQo85jqJE562YOPXpAxLWUqRRTeZYECOazeQ7I+fVWegvWYZ0urpge
MsB/xMAfzI/FeqnO5Enr5ovhdXnVAyrh5M2C/5n0Y7ZurFPVClUJ9lc8C6/cYdvCqdv+K24zY4p0
ikSAe9aaeQ7xj4RcSd7fKSEdC//jLeVsgssSNQtylHtGdRkigPlyiVgvTX8NTNvRNbfWzQtX1PFD
E2IcG18Zf5dlo/0yXr8N2bK0+5X7RqOjZVwVIG76fB/lP+G72qwuu09rgJBXAHtakDJYp3mGUjCV
GnXbhAZLJzMpmQsQaaDDm17ivnAG9pSadelTMxDc7hSSsMiaS0RaVMdtd4V81bBcJafP6tdkujou
9rq0txTQqh/RzSWce25QwiIA2/lwgh3o1VZTx+/dMySsZ7K3tBEhSYMNZhQgmibv7z0t+gjT0mQ4
VNzSbc8tM22eOacz0+0YOYxCFdEkuej4Jmuy/P48JDVcc6uUvf/+b4w537CD9mNfrtD2sFHNOmlD
HifemI880+CpXaocOyPQ9OLqBcZcM9c6udTON4iYDg6FFqPWUlTAiST8I01eofYloJGATCCuT+cc
8uJfMG6ibp+mTlYanjtaXM/hXftp88GWOY0Z0CZ61DpnOLw4Hk5+4M1OXruHLEIKxsLCiuY8+yOv
1NaBNCHHDybPXFpORO/dSRm9adyxAjFnBU6EgNCoTuF4xziSJZ8IQkQjbD3Lqi6Lie1uE+jXLwo/
TrzOIDgSNVyeoevxnQbVpi3AxecV1QYSQD0aK71yEeSx6tn/g+Swsw7HkutfqLxq6TQGrFOyoco3
sL4TPU1oOPUAqZ2M20GaEFzCvOMPfowix4NervAycSkAZKFIEA8l6WBZlyXkNgATGNGsXCbrOxho
CU9ZG9xmBnXyZJHIisgFNuq8U3nUnbyZjMzo0XE4KcofNucTTvgn1rmjhX6y3JuQAhcdzzOtehqv
9RaW8JaQl08YPoHJzfOH6eGmLH7FQTO5Lz8cHkc7r7SwMibkbeXARq+G0xE+HzuKS9MZ6wrqWxcl
KBg+muL3G8EISlMz76wCPp21jDSV/ww8hl0HbKgihECcM83dLmiUwla/2aww44EMU0rhK8fmx/rc
Koj5AIxJ0L62DGj2M30/iAFDcdnfNrscyWS4TvxXkjdnWILBzIOhGxxyTGcm2K3uz9tXpuAt3Z8g
ckAY89M2SFbmyIgUaU1OLt3HeBbLLqf8vvhnaAc/vVY696IeR0/HG9OPcY8iA4rCBzemIaSn00Am
mj2bwvOnfiSoXcSc5+D9fYhea+MUCBYpXFlcLhi1aQgFEYtcD0cdUVaX/TtRWBuP0fPQ2jnyKHsL
WWzLOHDlF8tBb6+RWIJqlnUSFGyKup2DHZf+i2Go9HefrpOhZ6U2pJrX+YoilPjGRMGz37WwSPHS
HeRzvpVO8Yu7DK8olhgEG2X/E8rB5+cnALUKaIF/mq5k1H/ByW/Iubt0M/OH/Zlob3NHD9bToswK
qJvMpPbIo//qEhtjTFNNx3XL6+D+d48bqdgaZcULThEYPcViVdcYyXuyECQ89LkuSdBdYFZl2R18
HRtqKu3j+OZ3O9JFC+s6weB6dtKUDxgxVnQXFWq3Po+KT/XeudPCe+eZzuzwSGo7FEDMFqO0nbBx
KNv8WdezQpV0FxG4BeXiD9zImL7xIQ5AN+RRXol2LaFbNzENVIwHaEp1Z+xdu/qYOJl77GzHzunv
UNFZrde0+8KJCTFErsmigIP/mntTPHM8EEvQ2XRFdY5Hzt7FK/4jsculCG7L+sWQYqKf2/7Wy+tt
pmskJ3R8Qt0WA7Q9uIodIdVHEp0JoJD4AkiXr4T3CeQp4EH4fn+oOyNXT+5tEjpXZ/8BE4w6zjgU
JfFIjKZ6iDmRzUsmsHcfiGSYQu1cr8kv8XoAz1c/4k3ukl+AHME22zLaCdrsvvkpwy2LPkFUWI9P
Zyf/bPjrEZRLClgF3E0027uiMy03EqWIVX5sLAirIsgKDiqM8ow6hAYcD5P9MPPPVKBu4AFkkG1j
nI8wTqsB6+3hb0fi3o/PZgcDl0M5yMA8GvprB2w0/y7E5l49+0Ydsi4CVc4tgqx9H5Xpd/VIhatP
YsPYo10h8QVKfhimoHDMt2M2143afdk9R+CuXLB7ztxTy0KKafVmPNC072v/lnmXO62lgqTY42m/
8QmQ/yZC7+OMFfxAqI9ye0mfq6vIH6Vb1poPuWGzB8r8QZRsPzGS6txsK7eMoBxlu64OIOZfVRLm
oCFLe9tjEDRjV/1zanS1LcN+z43Pz6nDc/sVpYcCSB5g3gPXb388cGK1mFKlPmxAuV/aB3dSj0Ot
u/osOl64WnlaYwHb1XiaS3OtcDF/YvjMdudSJlq8OK8ORNpvwKD+CMFm9/RmJgKI14nOlIVhr3QN
QsErlZFcUfZ3zaLvF7pNCNV2fSUvTi3yX3acvrkRgfI+cIu+xfZ5aSfwWS/NV0+uwreY4bHic0EH
ZfXzhEuEtx3jh2Vm/TIUwb2GVCsTfhwww60sL8fg+yMH+Lhy+Hp+dFJHT0E13cSXYb/7ptStPzCY
+EonL825Kugkh55FEY76XR+urFAGYoKxxtEyrQXF0qs9YG87Ico4Rm27cvHN3lTMJiX7ZJSznAMM
yGdr2B637pzVjektjfUKbG6MgExBo5wtpME7xGaWobl/vRFRrcHx9nep6Lsi/pm6sLgy6QIV70xI
0QoD4J74+RsdcNkOPkX1R+QvScGGL9Lx7oH+tLBt7tqIqfLWjUIMqMXR6QVpfL16b9Rh9YQmzzoo
93vT6Ofzl/kpswIHl42PDMRyYjDYABNONAQbuxsBE0QWUyMuVvL7y3LUp9LGHCnYN8TIwwF5tp5h
2LCNzqV3gRdD1wlZFQ9Rs+Jkhrox1QwK5ejnKghLXGXQjGqgKKV10WfEhixkyEwsXSWE8jLB0hM3
l6qKx0CaUBwHmwqk6pfbeVuqx5MCKi0MBxCo1LisFlONrfuBIaa9ekKBPf//kt0ErzD0DMRlJ3bn
X7rgtfAxpMgrHmlO1t/LiSDKpWAxFq5OMYxA393S5I+QojSZHuEETds6d7lnTxrzPFY5/CvxlhZj
UrP+D+RwhW/a98699IPAGWNu4pT9z/U0VzR1vwHEruhMt40jM/m4wZKYwu05X4Q92eWZCYsqY8zp
ifwk/iQW0+5S3R5Sf7dUqFGw2S6ksnNIXtxRmdOGRLWgLGqaXGjpW2Zw6YhjSnDuEYABSp0ytmp5
Rx9QmlRLmwCZCyzN668TGBeCjnaljon5F7ykESVG++ct3Tu9hi/DsKzZzcN0U5AZm5PNpluz3s2W
9ePzmcTpbmVsPeg9DkDIP0Yf8AQ4r/eSn5lb58T4FPjg6VIPwRUHqoWPRa7Xw+6QALT5Pl6qKBuC
pWeKULZ6m6wZJytc/CdzrEc/swwBBZdna1ungo2wv7FWinOWGv4a0YQgTh/t6HWA6tB0wdaGT1P3
tkhzvfd7KHalLWzz5k593rjvPjcGA/MGn5nYwFSnLC1ES6rzwIZg6j0DJ+H+LWojyXAmefkpX75w
C/zJS6GanlstJfJO2JxOKgQGramVCX5dySqnrAzQ+yY0niojY+cTRmFMHkURNTYuiPTWX8KpQXH8
k0wkCGRa0oNocQLUnAAmOZ+RobXoupN3YuBu8fqNEpwLUEfmmcfUOz/Fa3O0wo0e26Sj9OQTA358
VNPeGi78l5jFPE5HxJsa+m8PGiu/RvdUQOfM/jBoFkFx/yltcU3RZVKGXMxxe5Er7uEyH83k2nML
U+OHDX4QfBHIt6L+LvEsFKmWvZU6W0bmQclwbodbpOuX17y67ZcBgQtBDN8CrkmjGvx52MECh5Ue
5H+7W/+vfEIN4cdYdW9mjVBm5MkQnejteVJKaLTGeUrHlLfbNcv+Zm7eWW9A/+/XO1ry9+fPor1j
jauh6bZ1xrIzYAg7s0cNqsc+yUezO1XxI1d//+MkFPC+4q3OcHkJIaQ9/hST+CrRFoj5I2K+9M69
+jy5IF5gwIluaJH1VtVO9Ki4z5BKaY0QXS45FumYilxs2bzNbOJP60797Vt5w6lJJOLJnwFjYohh
dc2Mh7OCheo+RisAuaxfDiQ18AgDq8dAP9t+FxTj2AYD9yAF0a5ot+6IpJ0n7OfE13nlkXHpvNZS
sF3HlvArFpC2ZgMzohN8r9LfucNaCgwVCNiJVKdTYiPCoXMCyN7QVj90NVBth93xivR/T4hHlHwt
SzGiS1R/QTY7/4sG71jLTbBOnXI0NHD6IlitRfB4olbzAdrZ0ubqxaE7pZUY1/5NJsNqFbanF0KC
wrQJotK6pOmHswg32skffRELhe0dxQJUtRj5l0FVeZ5BmsrYYeRPXqGd8Gsyaq7Tp/1S9GvJT5K4
4C5GWOceqkvduxOdE5EAN+rRSKUXIaU0Jxl2+erQLR5uIPtr1YwFhHiSjI9mosSJT6485UEPCadj
3BwzL9o/qakL8iJy2u6gVYUgVwh/KbBpLpX9rP7RKkbgw1B+RjRz2g6N6hzfhEgte/ARFA48yU1N
20ih551uLD0TEbvwHmK886dYsR1o9hvpSsEth9gNgEiDUfExM+51SiN20qKVDo9v7mM8nsRBoYQd
ViuM3wGke9eL+Y4XH1Y3eXS4ZhlorPalBQNtfGueFJdSUZoCiRGwwvZboTbX2cFFt3HzzaXFIhvo
uUZpqfE3Qw/c8Er3GC7ivpo47gZIXJPKuQhbHR46Pp+lGuLvaxNAIpTeiJNr9n2pZGr4BQ9NZ552
EPcawml2IoJh6o/cQTuQEysoULzdjZCydHG2gLYWrxIt7BPBiHfKMfBEF+7Sc7RcwfN97Rmdwl+E
uo0BtCRyVF/L1MAFe8n1K91uB1T1Qg7CebB5SoBlSZ+1WHTFtLz7g5OqwUJ4SKdlqwWdr9i2SPj+
LJ6/aVkgURwJFmWO7Q+WXRXEPk0EfGEp5hifwIKNMaeFroSlMM8ZhJyTJoKy55Z+tFSZ+yVqXjmU
kvG432fkosaIUJSNTHUuEjZCCa4VKM/YitHrRg/X+KSjGq6DR3naJQckFNRMEYbvKfuB/4SLPzev
dSr4knx0wI/V8mllBLVPyhwDVj1e9fPjfQEXDl+FCMryENyoeLyKD4edhYmwgPfPq2PrFH9yPMDF
EgVgqSnlmXOA6elqB/N6jgZRKoJS7TJqBCAsXA0+k7nAXN61taNJEWNOgfryyW/yW1+8UBD6kPYp
Omyhdcnk4MfePRL/yiyztOssHGI80wwqtYVVXIrcGW278lMqrwkUMUgFsV2x1mXmtJCyF4ILBvwC
YTMHlApBwv2af9DIcb9gxi6XaL1tCJLeJytMX6zqw5NMTmyuoA6jBRZs3QlzJunFf3/NsBa8VPSP
qjQczJFUkGTaP7RNdLxer1D+uQvnJHIBytE0GdrONb1YCVN68HIiwBcQjtL7r4kpGsec1qdpOCpv
CO0xOdU4MHUXOWHzxCI531FXc94ObQfMRKIlPP4lY6m7j0z7tM+XLiXkBItA6wkt0cMNeXBF7rgq
gQ/KQwtVoZmqE5sk0HENT2dz8jX7osfUJOBkYtxFzWBb7iyTQOAITiVxtccOLFxZdxbakeUriVi0
FuR9c4GTF6QRCOsc3o4wM9z8gnJNyso7l33CgkEB/TOHZCaCOqny8lyvkAcMgvAvN/fZNcp+lsFz
orJ7JwiXueZtzS975+FW2Gtj2OmFvGzY3qcjVvR3bx81L/KXnCR0uNP/DegyqG8cq41m/YjQKOaV
h3A1jwN0qgO6RIRxnLq0dlFyoTkXHOfQaL0gN68JzRxP/1AjQsdHSb6/G1EH+26oUZotGXTlpfX1
nj0QbbGleR/DJN0vO3Zjuo9D1KtJmbfvr8JSP/FVPvtFzwk/r9HH75F4pWQ+Xz/PJqu5duQ8DNTP
sklLwY4cop/wDf3+qu0BGIv/Pr8ZAIghCGpLWO//LIk0IjjULT7dlvosCqroO9gIokeJB5PvJ7+r
iB9ACYkaf37euzFDE1+xtdiSavgqwTcv+0qpoDcRWEIjlRWRmSNuAzNeiACoaU0I1AZweaJQizxW
bPhhKL8tRVhFScw22sZjDSHoA5CGshOfq24rAtgmrdVwTwH7+bxFkXMPv53D2pEGnlqqmoLSrkn/
mgXS1/oOCNokg15Uokq0Uei3VB+GeE6eloekZtEnzi7FvaEVc+JfDx7AUM1/rxOcoR6vZB/DFTVW
ErwY+Dtr1TaQupu1bdCgrNX5WVICzPZ7RmZ1T9DwgH8AecKkBVxIDNyVR1HIgY2WgQ6IBDmnCwto
7JfamLbKmqYE2b/4DWwVXD2YO7v8L0aiCPJFplspdE/liYYGUMUEQj0klmaF666fIgc6Oh/3FOs5
Qm7D6XzFMHIeUe5pLt5oGmk7+7sDUSVFo3TDlILDHeVZZz8U7RWQB9/ZRFM0qmE77vcXxdiNEXqh
YFxc4pZTjqt1sHuch2GKxUmobQ2UZpjaZyJIrQLxgX9bxTJdKf8S1GvMSzhY+xzBrC2S1JxtrwVw
iuBlbMDT1owqT6FdBwcbIDK9ikGzOfyitXctAY3k8XKnwCzQDpLk7M+WPdMQP9sWaFMgeqTnmwq3
4IXjz3lflNFflQhc/GUheqZ/FebLdKM4oB6Jup3vWGgqBO6i1ICdIfAnoNjWAiKyWTVZcXLoEX3c
sPCdq/L5USd0iQvKo83vicTo3OvvElpJ+MqIEslAU5KnJCTG5FbAKZJob3USU01hnsGLEBpCMthr
aKMoMCZNvG0X1k69rxmKW5aVfiXZIsLy/cOwWKLlhSNAKom+eC1wF/6oNjdulwczxMf4JCjVhlUX
cg9FCETOSRwgcTO6cYQoXfkANe7gkUC5+ovX5xlbl6tRRBIyu7amHXQbH3JGuk/9vqskjn2A1Ffp
WE1CLYvOyj5eGPXl5VJ1Hj+kg7gg0fGsdyzZLFVdT+1B12DmI9tsnZeZ2KqAAp/lGfgiP74h751+
JdW/JDWF4dfOxoQ00giTszAyFHobjvoSLwIcrqtEyxmZeJQVuCtjXbtVW2xr/w6ifnCb+XBPx8+h
vKtW1b1himbgnyktiLbSosJZ+NZmLRu7UihTiyky4iB+vC7QLYgTBUL9125LqNoSR5MkBz5F/JSw
X6iDjdIO2+QAtWrBqr7fMiXJ/wX4UzZA3ITpGI2AyQg2YoXHjzGWo9vUc7po4x6ZgXtXIUr2a9P7
kfWCFnanZl1Lq+b92H57+qX+ESGQDVT7E7PbrXKv9v37AskPQwW0OlC2EdNb4FUb1fLX1RtHXtRz
lOvcweQdDf3MHLPRKX4hlSXlEUE0KeesoOPtfQxpA6mbLsRKM2qwTyVWuYAd3BZh3yZm8mIZ6WJS
iUX2sogrMjC8I9FaHv4aFAl9E8W8y+JA191bp+D/F2hb70IIs5kS5rJKarlCkHWaLV8NcxQ+b3YA
B6FoLnsrr/hb/HDnqqbkR415q6wc0mGsoY0jkb6H6qurETRssSrgz2D8tiDrortDw9StVp03s9Wk
1wdiZgDQUwrrNywqoQIZJ+0H8qSusq11XTxEzrDzFTJTKnNgkZ9bs1E63hryT3DLvkyBlELLE3Dj
UHDmzL4peWaXCuFrvOixYJpmMB48fQSi8tN9QHQOYpcE6HEbUF7/7AEf5FS1pMnTgkPIB5nskv/I
m9z2pE6e/wn7OluuS2pefnij7ST/uaZkpO4BPluMmeYvoh2lp/b29mito9J3rWvAW2PH7JEB6PxN
oZpLyvIH7QwON7irhfeiyEzE09jbuZG0gYLB5odiFtLt/t+LrC6W/ecA4G9Pc3DM41zpZk/HAzgr
ye8BYwn/pZ+j8Zhbh7iRr6V/lVgSLkesS7yGkqC/OWVb5dPYhEL6EzizwXtpcB854fqqiYpaO9Nw
1I3XFsxJnalGMxXB2hjFI6873veGyqcY4JvKxm4gcwMFEIHy838ewWQUhw4YX9zGkZCa4fTgTC1z
6FjJq+qb4Ioccfwp1//ps0sk2cqe6wdvKFV+4mRNHTvs5METzj7K+DucxGiA/69AbzfRVb8tG3Cg
EadqCcoT1MCMgXY15Pnmy/m+Dmqt3u0qUyDOxSczPZqXMQC5sFup2HlbuAuzgUOgn7aPhrvr09Rk
xMlY80px0Ozf/QizP0OffQs8DGvz9kkMnsSxz+6Yrmjhkx7TgakDJrMBcqn3TvXY4pI97XJegQGn
algE6+OOLUWGli5wOgvSAK7tde1CbqP0lsPLUz6fp4UlmID/bBQeOhWPR2mGW/QmZ/y/X8W5ezqW
Bct4uyJQ/nBtaqxqzZ2A6yYkxGtwjYsLeSt1ShMs6QQ0v14WfOZ4E2JWX3ZDHT7AgP/Xy5WMdtkv
rqzUTjY/ksPFmOuAEGAGC98OBRpRFu+5JpWIlDqXXRpYq8MXEc5fy+nPXrA5+dK1ratDlc7wvjfi
QnBN+A8Pk7hH31/XQZ1wGk5yw6mzhM/w8tS3TP7pu/kwndnYyi2KadEI/qoSE2CAbxzoMgnDEVws
P/faNowyh94bqxl9OaKdwNWiwAvNXBugyhj14waghINS5bprMdaNqD7bCbWk4t7eYG4maaIT0GEf
4Z/nUJ2k15DDRavVVtWMAkAxpKMIId6IKUOLKwYIyH2atQKAxiS/Uzg7vfIy1Aky4O9VEy3v0J8e
hIxiLmM6CTtpzNAcoDORnRC7fcPPchjvG3QATPqucEHI40YnamF9ziIK29U+iuxoUHzyaICQbmKB
8qmQk+kfbYsQWa2pODeipA0+l0OsryDf2e1m0Di5YohKBT10ytD4n5JT7gX+Y5Sp7fJWlObBJcIm
NPoGQ7OPaJFJyBQH2OWv5fO8tVTZEn6wwLwAQSwZk3U846y2D7POCeMzJ6maXJevtQoPVpqN8TLb
ogDJMX60cui7hmWScZKgRdd9ZsBy88QI1OtxuV1iK1ofJlVMbCVwH2vejPRZmytrxQN+QSdtFws8
GdDjFycyQqtbAdbi0QpluuMoXpWP5NJZYruk2ALXrH5W66ExWKBDI2xep37xm9HvzWUv+i6gailD
tenw4yuaAvaCzcSrIYaj6nZRcItetdc/RmvX/TBC0CKhNU+ddGuozOxHPwfX+UOpP4/3LF4gKbBj
EQG/XQumjzvUKWEd4pKao7uodIwr3kqR1hZQ58QNGzytkmkQvRcoqjccWWOVUSwzoag9F1jhGyOo
6dqrtHYk3FwnKmsaGRbI9vSaGVM1ZnCwxXvcsvPdcATAqjZN+8fzRtDSQtYg+sQ7fyj0egpPCvKq
wVU7ACH8IXBV+WGb4qf0dNoPgBt2hnREGCXrQYIkjS6CwaWZE2dtJRgRLO3v/sYf2AstUEJXDTfH
5E9WUpY354oAbDP7KQ6gSlkGwI1P8VXJm8FzIAVa+QZEM2AkXrjzXk9Q7DLLDvWwiGpwq50arYlk
BAyJEr/AumyYMs3NDXCcdsXRt/AUNhfPjtRAAjB+LrbqjbFX1o0gTJVNmY+Vzc9fuX4mX4VoDkiq
BkB9WxAfAXXwvulvdI35mcSlDw8az1lJ6Rv2CZj/n3Ff1+35UvFgyRwS5DXjAvzbgpxOuY7QhlI2
83JIjkyGqJLVculFw1Z8odjFzAT80p+aNG9lVTTpi9gYefimQ1vnSfbyRCzmMKgJgxMkMocXm3Bs
hMii4jKooDKJvM2CjCUocruqy1QvlTh2TKcuPGRAz6nR0rYEcR2yZhdLXubNjInAsB/mjSF24E/9
frnqbTXLYZsyXWH8AaHHxIQdj/Ga1ulFLS4I5NpiNF0nGJihIw2RuV3sxAMh20x227tvU0jzzAOP
C3Q09q5MFBl99GzhxNMIrl99fRtZo7V8yAlxk0CmrpTjdrWEV1DKztJEYEAGwoUYR9I2MSIScTDV
ypzgoJx0jI9pqvh41yVi9SUlgyKFi0r0Vyu9sg8S1QWIaYZ1i0RwvQD0xsM9ab+r+NMTFBAu3MKg
+bhB0gOk3skU46dunPMRcxEV9zJHRxD++HpeEHcyuwVTRobmsqTTuDv21nzlUUzqg58VjEiRbhuV
ds3ofo39xeheqCR3zX80V0ws6jlatMrO9vxIuaLHcqGwtsl+CmE9OqwKtTTQk/XGv9xEFItSJw0T
sYaQImouh3xU1Z06k0gjN4Lisvfw0Rv0RKkEwpUi3XwwwT5tkPkYRAHMizr6DRcS5PyRbgDCnX3O
d6LyIxPI0shWBPxtbkZkiu60ASFwlDi9V422QoOivaJ2RAnxo+byFCZKP21XxK8mhHorfNPfZWyH
Fue5R8q0W6wSyUG06AV79CkGoYDNfx4gs+U1WguFiwJ8r7lFkVdsjZMXdHdAavCOl9F3+gDmSmA2
0pmpkBgv4gb33uKfy8Hztv2bdN6l4dhPS2W7TM+/Gplq+i610qqUIwb6R/WaPT8Ht/kD1XSz0vGS
shVyA4fFQDXd7xh4GkqPO4ajaR82mJ6vVsjVNhX7Pjqn1mRv8rv2kSdWzrpuLF3XhvAjKS+jGKfB
X6yYbrblC8skvf38wrGNVs+0KxuQ7ppqcAvof0sUZRcbIncuV3osQgeggUZRhTW7iXY1Q0SEs3Bx
W70Gg33Zfqad6/yTCQnVgyq9fROURcHhviT/XCdj3vM4J6SQ/5ohaLJM+Do7cin3wsTf6qxDK8p2
a2i2tyucGvr4DEPb4wRYe+E4HqDCtxUc5IB8oXmDCfACb48aKnu+CM692TmbrKzNkvU8XPYlQ+3P
3BDxZAnswmmL1Xtba4xke1IeULZkETiZC/3ijGX7qO5cL7ZtEbuFvSGMIoLImJpWsp+ZPh3ZxSOs
2OFFTgJkJZnhCSn5VlAEPy9kao9UrkR7l59db/+Y5paShXEO3253PtLopL7lylGARL3F1knqFQsX
GzGvNpdsOyAVmpkItPj4MQQmg7RWjpVXeiXhM4kUshT7IqDUX+Gf4UyXidKaXLm6toBJ92zFMRc9
lpP76yB5hhKF2N2AJp1tTXn701qMBjrmkMsbTXLtkI0H1NapoFUFXNdym7X6Ku9U+eZL+d7dUr/W
eRnE+HK9ZVebSM2aJ4z/F7HiKhhRKkqGIZl5YSPrCZve9xIJpi0LiM5TFyx1Xd8KzcLzt9TZtwA0
UYuG/0Qc213HsjlAVluRzJngSzC8DIZNTR27LK2ydHTpfhnEA/N8xYTAtQzl9NejxsY4J24wMvzb
auFL+W0Hq/yUwdIuIXFVMbDbzZiOhcHkribPegMCr6IulHYJ7jypb5oLutTAc4vqetWSi6/3Nb/b
fT1DQ4d5KrCkb35NS2yVBdYh+v0dNsqXkSWasZvGpqCdc6SVokQB4HxSevWqamxpN1QXgGsesTTC
d69eFBtHskzonRORaGTjjYIS0vtTTiQRWtsFtl/php6ECU7t5rDdUdPCveXI3DxpLW4h6803ZHA5
TgbK7dtlI2r+h6QZy790NGLEF/fhhZ1N/1HYKkdV+CyS0MmkwWA0TqWtSuZUHP0fiGOM1ruAJ92D
ldjc+vksy3qzc3y+sDLiYq3ykFFRJQZiVrhrqgxP7X+zpTvHjdaaIoeMiUh8zcSNmYWgGRREmgu0
7e5LRqeb+Aks0lOg2wQpPB52dttRqiesdIQX5bhxGcqE4DOlkj7UljanDRSyhL6a+vw+RK5k7C8P
xp55GU7VMxgRyrIm+GwiI3bHdbk+7apzZnpnBikZmPSy+hRkX/J/+XJ3c37LD2GOOIri+Z9Ahqoq
iX86l7Zib4j/DnROOUurlbWUbH86u705PR8hHt9jfc8NZ+hH2Wqu70s8+XANsgmKiZPx5/Dpqj6A
e/HeVQ/W4GNCzvRWO2HRHyD8iopLABvUR6p1lccNzlphhJZDck1kY0LwkXxBEh7p+PuSH5r7q1xW
jO7ZkEqQt87jC8uXz/g3/Gik4d9lnhBW7nJSc+oSDxJA0hQqprMFv8HTCVaa0JVTBBzFjdVQAShQ
PVkBzRsof10YHn1bz+syoSgsYwPbSKzDdJSJkmlTcX8owJUCYx3x4fFOEarDshbg2WiZP3+8686a
0/sdYma0QsDFLobJRRyrHC3ZV5YxYtsxolFbhjhfCMT7FMTUvauC7dB06dYt6LULX/oABdcEDnbw
0ky700kxpM+M7c4H747ryvcDhCUxmrxqqOJsUgv3MiMGG/t7VZoIY2cKoXgXoMWnbw/4P7SN89Uc
2P/vZhmA3NoJNwJNbAhU0h8CmOG/KaUEZdYig22b6qHJtLWuwEVugFNzMkETrW67t3aYn01V9Wse
EvmSiMQ24d3DcHGBWgTQ+CpgfWnXcmX+ht0px9YGM2fqFccb0xFOwM9ItilLDzLu9ekxLN5ZQ3Cl
+OR/Y1aQaoZ0/GtiWH0xp8obghda3Zu5kiQuskWQB0poa6vokcMQ9e1WNyPKf9CJFZZNPNhtPH1d
T03/ahWIxkKoNxRQWRywLMhiyA8L+wVhqrQBRENM8fq4Q+nDZJz+usa6nlEtBiq49iIM05w2/XmK
LjDhVkkSkvpCqbEnBGFweTb4jbufL3csgzHd/dzUymG0ZMkYhCnCnv/0i34zZPEZPs8VMlqfGXGV
37295hQeIiW+pcfclp/i6oE5kUA9RIvs9S98tZK56eck3nR4VdrzwfWHfhFg3cENR8yPYgKFY1aF
0Ou3FEDmDtg00Jasi7vZ4nykjUfCMceDZx/qtRv1NhiC4YSMC7DNaeetlkWGhZxy0SxSOpE0won6
DCoSZ5nmfkiWJUqeDui9arZOBqSnpKx9LwfpudGC9IJKN7sn8eTOA0pYPA82QEz+hymeXYCNxrUn
cSbRRBh6a6kJOiFTO7GgIoAEiGn/RGsgadmE3qnORu0glzBlTsh3gke/1KblpfCf6cd1wTRxdMSq
eBEcssZ+L3W763nGWmWDSlndH2b4B/d/VRLV16Oj1ZpcsiSjwd0How2/MkTkCD6/YntCseGEIvdI
L74PjvW0HeTmSmZ7qJdovMx/ZJONtwv0NuKrMnEqzDwugHFqQd+W5Wm7YBCIYCHzNDq+oKnY8sJE
VdmsNUBj72oab1DZmuD+w/tdjMYiIVsGeDIM9FbnJPXqX5k49/0VuKbbk7FuoKhNT+osBOsHTYRC
Bnt70EhXcSVYcz0pedo+Nwryf/6jKoXVm5rbyCH2sf5TzeOEpf3g0Hn0UjtDeWXjhO48b5QPeRfB
2VMqG3Yk9Pr/toVzfIq5LUe9gdP3vRkpSwW4m01nmmlhIV+gu9f5ZDR3kvXWGHCZMPoda0WuXCqH
ElB+hBVZlOEdUjpGTLRg4QSgjxwMZ9jfkhmjfsSUlxwOFWPW2GTx3J0a+Jyads4Fa8TFac4xgAWX
J+NZEA0SJ16Venbiaxms1TBL+UvO6AKMAy6n24bfpc1y0SRGHeVCK0gDNqrIfC0QlUit4wyfgiIr
ESjRHdNf5TKmUNglGDfiEQwgFMBDmPm+BCS4jA8F5+hcWNoE7GkjLrtHKEHyLp2gp9Kzx5Ard0on
lhWnplcS23YTbKNjI2d/B3+Ry4tl2XnmQVV68W/c5b34Z5cFQoFZAggLu8t/0m2LCjfXzK1Hmcz+
IQGnSxhxre4kJn3sgPObnBVE+qhOyEGWR6KudX6O2U+kZpIlzbIMfXfM/0En0XgwS8UARLDFF/0A
Npm2K5xLDRcg7wyO4thWM4663Kaf7XBK6MFnSLCiov4b1C0MzWz67QvZEcLeqSgGQYf9KJPgV4Qu
w1vYtb/Lxl76FPYNLpcdWRxPsZ8nCmA2Vva3nLxIt8upGHa0+DhnWQ1xvx2i04jtQcyhVWCNI0Po
edTsG9+tD0psFeD+inDpLAhNQhS9zk4nqfFupGAqVqKlivGU3jyjxszkPkaOIGI5C6kvqoD2wgsQ
LFF+p7CpquQrdlBU7spGy/sMJM6kmaiy6vebIcnjcIRq3m8uxf9UyOTPmT1B5YIW8aUHl9GfGLtE
pGP2ccLD0XqKb7Mmk1hBaiBhuKkY0o7u/FbflAUdNoMbwnv8dpvBiEztLYKskQIGSh/+wrqEvTM+
0BZXRthPYypLI+/lygUQQdVK8xa4ysxZZYAG5E09vOZ6Xx2Muuf27BRcbM0JJRx3jUFcQ4wUF+7K
uVs1YTA2eHWOD4wJosbiIU2chxUuhzyfPGmBbnp125Ef5dAyiOaGutTaLwef8+2nCoHg1G7o2i2n
eMBG9h/hwFtkNet/ykml/kJbA564hESvDRvDxMRnHounB5kqezBCEa7wh39mCC3HeNcJbBLETjvm
q6xRDqIDjrn72DLeILsav5j58Gn1hxvs9Wz0YdmM4d74A7SO8xDWjdccXe9BYMVOWWDze34cwj6b
BRlmFqqJtPrXZxRkjwidqPDYAT/tiBKHdbA2OdnVXYXZwYY5l1KUxLybDermtkXqKh0vjOENPjW1
2Fgk5Vw6D/9wqEUUcpBb9bOwXKJm40EEEXjbWBS1b9bc4+fhnY3I8X+snyZVbL6YVz28oatx4z9F
aDgiNxKTPjMZ8v4dVuzPoZpVwW0KWcCrpA3iQpq8PuE5+UehhLjMrwyN1kSELCYXSZb9D3oHQZv7
SNJORg3QEdKSq+yV3aIBXYcjJgxcfJp2SHM/1Ohwf5IFY0MUt/f5GN8P9mnXiagwQCe6LMyDccxL
rO7X7xvcfce3b2elgsekbZQz12e54wuJl/vs5MMSE3f9s3lTz5ejYR73e6vzZhHfXyDlCIdVsSHV
s4K5qCKxWS2kiAKE+dMIfIpthD23mTEVGV7fGBPoMNJ6KyHQmc6Svn1KkCj3Ol/lEONZJoiip0w2
dDLfHflLA0XozgJI8o1C4Ztt0/i/8jJb7Iyks7ZMys1n/m6Z5EUQsIpxaYNQBox2xvEOJZe09WlV
dQgQc5GC3a7O6EfGdR/yxxkpiqgYmezqql7o89Fpq1lL0tqGoOxNe7KI29dJ87ppJ03HqBXO0r/r
gasZmo+0fdvqa7/KVvtb2s7zaz20iehVgq0qXOkCriP6MN9qsmD24GhKaXezljqiOw54hDdwkkOQ
ZAal6rBlSb3dPl5+lfdvFabxXfFd7EQ69BMSh+GHQoE/4IqV9vKfOpDexMqNv6K+iXWprULQvalz
QcmL4Y1Nn9cLvA33QrvF1ngOY+G8yxW+C8um4+ojHtFr1yjRLewC8V6GmoOLWiKwxvk5KpzIZd5O
ztKbssJ7h4qnJZbvDnDzJcPU4ddaz40Ncmbsk015H6HWZ1kqx5ZfnhsAIIpnHKgaSE3vlfdVhi55
acyoVj5yvORUd2UVZdDSaY8qzG8bixHXk205/UKP9+XRTLkVM1Gm5v9r01zFtMpYR5ZS8eW9bA2s
R2thKAoi45ZJpHDRdoMpqU3R/4c0hw6stvQuowxz+KVy12oQpaqNWueK/0uv85B45lrHsES3MLSu
hb2yJWIQ6vC3PlM0jCSSwKUOjVcLvsXyIix8vnSqQwgpOAOeWYx/tJIdd6EqcayGVUuLxhYUsX/a
v4kgf07OSXF/AywkKLkZz1D7FZGq83PCkI5IAUHLiCGKcHWXvfQBdH1/+4o3mxf6UVw6P8vtQ5RI
AdQcquom9nnLv7+zY19O0TpyUs0SS/7baQ24my8WYypjPslg7OrEDPjKm4lnTmUYmAeJkWay/KR9
8Z77BP+4u8pH7AiswTySSUTPceKg5R7yTIj2HC43oMQ2KqYyJx2sYUcef3oszCbXIJgdb3li36BK
DjOntmNBZt9hdM71s9k9WHw4DYNAAj5uOB/hg1YT2OZwBSugvIB/Bgrub+H10nIJN6r0L9UbgEFU
MWBmyHUanFJr9KVuSDUK0L4dMBj1XNgEdm13oN+QqaFObGQexS8I31J0+s9WNyKwoM7NPbGR7W05
ro5+TIUD42UeyCdMlSFkpmyuptpEbUeTdztB2WaEFRKjB6Cqhq2BQiQvqHnjfHgrQZgGI4176IGm
2ur3W/80Eo59N1zDm2um8kiw2QNvul/jgy6ZvcDVOZhuMB80fYIG251FxBz73c0nByIpSvzQydbf
soiNXiXxTaeYkxE69yaho+jnmmrAZyG5ocCKqou/Vsq9kOVoQ+M9xuVA6es4556j/m2abZOWkofB
c6UrXWqc6/Y6ojugvq/y13V1OeiOwywRrABpqvvvSnAKXO4QlXm6d27SopepeShWAq04D8YCU/BL
Qp50/8aMu2gXev3ST4P+m1klaXsq43sCla87xRzEY+JOFHYD0jaV24V2+I2IuyPRP2w5Llbrk3wl
OWQN/hEZTVM/duHwRAiPlTBqvNQsK6xuXGb7y/p7ZB2IzlDBrpvPBqt+qtttUVWtsgnmtB41Ajty
9i2xQI9ODKh8tlZW3wV9qEluoldd8kgFTAORlA/iDrmkpIGZW1ruuruYwrKXcje4foUjKEgqqJFW
8Bn6/IgNjdLabJ1cZhStwybNyxSCktsvl2gHEI6lgLcMzFCnuGisQK22xdz0Y3oqlpjEtA7puilp
4DWHScHPFP5R1jT4AGLDG/OZS/hyPcMN6045k0SxBj/7oCA2mFeUW2PgeMv69AwdGJt2d2CZoMav
ogYmRkaWfEnYyr4uZztMqBuGERzuFnftwc5Vu7jbFwT3zbmPACycdNWjbXdGhwHwMTG5MzurIRNe
bEbT3iA7VEVePqqkaQQ3qmshnLbiAsRvEGKch/9818zAc58RhBz0TlgaYZzGHdJgnD84By7MNsLQ
jI/JJ444Vs9705cVX5cM1WNm+pRu548xQe5YELn5jf23uPjWAlGoN5e7vi41VGKPEEcTH8K4pRLe
RgUp8JFzCeYR/R4ZSkNRRb1ndtb2Nh68EB6wVafIc/7B5MNVa8VELM69XJUUL1lgIsJmIDBSc7Er
6i7/tDDWDCtfU1k71WUe/ePBu/namsT9l2Hoo7QFCrUIAipL9kFJ1hu8Cq1AJYEhEh7YWtRk/Jqm
edDWclUMzCZ0MOdniSk2xjb6mY6abIYqEKrJ8WJAZ7lJ7rgl8c/Y+xTRz2Cx+7hRGNKVrRcU9Em3
HC+LAR2N4ef813xdp50ZiQkWpFPmT+kcXXGiiNtb+4z/ah6NsHOo7B6EYTvRJ19gimUOGlcA94rx
aGDPnqGm1MMw6PKp3rEF6PYJl68DSq1LcVIeboPqUuaOr04WDAdy52007++wQ9Nbj3OtAYJwVzBa
PbntAUz1j3iUhB/NssBz97xjSELmHrpO4pPlS3m8Wng4GaS+j3BiiCMr99VoxV9c0TUaEDrqlLRf
yTdl/rIhCvc2psiyBUG06xOji/Z3gOk/Vt7oD9dZnZgRqLe0JSHTrOpsq4Crxa6fGICEYVIBNJoW
qS0JR2YCbnwgxI6p8aYQ1khlj5/qj0EQRXMdViF/bGzIRbNGrnuF1uA7Ss0DkV0eDkkMFJrb+t0z
0gMDHRYTXstAsp0U99AUVJk32pjsjAWEyT/sQvXC/rPPBTiq4Om1KzjgKM8R0lMPlC9IzJRjzKBj
WFH4PysqodPDzJz7lrh2pqnaA4oPDkYc1+bqOt+NdiP/8OZDS6svUHmMpj7lt2xhKtALe7w6PG6e
hEd50q+ff3Vc+54mDdYCkMBQM7vEI3o8IB1d3X97VlXEeBYgg9m6X/4d5hddjrCDslBL5b1d/pqF
GfGYOAPo8ypAYofNUf4TFMfLQarCTvleZsrTt5O9EDcK+1YrcWMtDzT1A7EB+aavxOj+Pq7cppVg
ylUAH6hrxS2SzKnPkGUpewXZE7Ql3CUGvRPAJbRq5HFvnNhfctEmuUAvmJeiWRhiW5hG5bURdz+z
guWIirBOVbiTmN44qFKFys2J6IN5VAyzLCJipxN8SQoF0BIOf1xnj54oVXY63L3VeL/xnhX5H4aq
aCl6Iu6XqXOxUp0BiaDYkupc3PpheAr3r/BD4vmq/tOWO0mPivpf+dRuB0q80rN5Oe8wDQdn9wHo
TQSdti91emVgpD6UM1N/JTV5iAbJFCfwx+XuPDg4q4oyCuzpAF5BLBzjmH35rsF1iIiDkW197jyP
5ck+BEqNWJii1HzS/gZmsHi8mvLaKIvi4u/+ilQPa7RauFvUl+HiWLdWMtB9ChM9rUSST2HWUAaD
BckJEdsMFf2b81ngDF0eXxHecC8/7xewOiWFSVpCDJlx0dVpMNmlc/s3pEdRnPslhooAUs1nU0W0
m/MxrATkMHbXATSjD0Ew/gEe6cyIk7OxiiTU0hfNi80lEqkTcpwYXf0xCoy2BT0ZSs+KQ1UNBvrH
x2hPQYAVoziGVLck3an6y4UfBaBp1btVa+hQ+tyAupbGdfXYxz+VHgNc3QbUKSTZ68wTYdMEw+vX
Zy47ZRQQuxaLs0GqmSVRNxNZhpm3GnWcyK0DU1WGclBAQPoz4uCE6PTd5WN/uURhbbUP8HsMCnwH
tj35+ZaJ4sTYc2iOeHzdoMq2oT+VbDZOPrRG3wcGHn+8N6yU358I0Ce77LxcLIxPJoLcvWykCLtX
FA4iF+H0ti+PFu6vdneMPQCg0ysJMsyRoL4695qsL5yv8pc1KLalhQuNVP9V2fgwjJ/xvWDCF1mn
4VmgToSuNuxvwdhmjnJ+5pPLEvlikyCb8QriaxdOwnTPFoYsIRD54zQ8gUrYdCDpFAIXzAGuv1/P
JSNg4BWXARSBw75L4iGpKI1KE7LRklF9djTDxDhrQ7NiUeJoV7d0sQ25XBELmbx740r8dGneMBjH
lEGul3eC403aQMy1ylwqMB6rXCO6TH3HtZqXfiQ7IuyPcUG6dWgk9SYo66cml5laklexuHKriK+i
dJRqbafqaSdm5+YHFyXpPYVnfie8C/sfbxiGDQjGctXFf9RSbZaOqppeRI1RSS6GKCH+rAPi+RiT
rSfdUkuSkwCJrjoAc5sJ6znTMVwDkxefRvt4bKIwE1xwLlQGD1S1eqNbZltzqa00T87Q6sWeiFFu
OTvCyEOxSZCX4enjrGpulpl/f5lQ+av/JxOxYUdqon3HLqH0s1o8Umr6yfxo4eTmUOuGdI0nUWBJ
ojpWP1243cYrW+t0zMGziQorv1IjbeLPKM3ky9lkYFI1pG8MCnjvG9itC/nBy7k0Kd1JbXP8Sl9j
LZz0Taolu5awO7ecnmxekbibim90YAIORig/803aiL8ErEAVLMPOCSvOG0xjOG+sMTgdeZh1X3F2
bBVbq/cDIIvn13eriOTWM1XQzVdEhj5mP5XL8+uHbQ69vPdPCJd1ZQ0m0ycdH9SGmTtBM5o97pC5
SeWo75E6FV8XUcGa46bYHLveOTCgvX0WAWrphN3WsPcBjTXjObBWD8m/JIVTJs2WwHIBrYKs+gkW
2lslgzI4e9GfrHIrVdDTMdsBYuU3OPQ+R0C1I6iWaMJnrYQFoPG7OcehqDwDmKTyC8Yakfl4HJOG
i5X7WKEZtTQtEljwvlbnTI30ymGOjbw84GkfVg6nvi6etgnhogzR9K/vIDthq41NTW22dGKYiTZe
/dUqIBG7MHz9ucN8RjeHLEF24FAXVyUPMIlRs3MPO0Rd1eA+bsrefj8sQjykHI+X5xdI6qW+bgGS
wzijg64V9i59evPzYNlMm7oP/depbEqt4Pt8qovWp1JZh0eUpCNAKN1TfQa3lCN9ZXMmsuCCNmMF
lV7f/eZMaQMvUfw4wT4APWJr7t82SOq5PhwJd6eDmBkeLALGKVQKoPbzn3pfAsuQ8fPK0FoqIspd
MlfFxiE9RKnis4U9OeIWCWe+XIVFz/Zq70gHY/A2yShJGuZwkiB7o9xPQ58FjzaoUSLB6PBumU8p
LPmMcdFpjjel1bUNkAPUjWP9YDZGarrlMNRbEgALJ6HfgJQ1/asQSBD35Rx4so76fQATLKuu0+TV
kTaSblDItZU6Zq4TobyQaRbcFvhtqyzfBqtzR6Je1FimZjJw/Ws7CNjpvIvMrPZNFl4deh6Ce8SJ
ddHJeL7I0JwyIMmw2rKC9oSdFETLW7OQHF7OScAPQV/rjpcdzoc9KLfl9VgLr+RQT6HT67YRV6Mx
+2GNhJ1wH3D1d6bwfv5j5lrWyLb6uyYq9igmYAhMnUY7PKsxn/vmhaxEvj/eKHR2aSZWQrwGozSO
Ery/yDKQDjmt9VJ4e8lol4V3rEA8f3LXN30j5tEw/h9yIpxsUCtg98l7Cw3lQEutXqqGmSmijBrO
yUDBDCyEF+G9XamJovLm2Xu/+Zxo9Iv7q1Jorjavmm0R5qCMcyCOIIf6ja0IvmFX0m/UPmgMABai
PQktwaJ3PWjx2xwyhkhZUMwpXWDsrUo7B5DuYE/DCYaOubGkg1cFeychr2Q1gO/PQAr+2K/PvcfY
Cy4yrhKq5ZsUXCcZmhrOozh8BHOrG7Oqt2zbo0wfguwXS7u6tKlhwWKi76Raz/VDojVhLZrJnerp
3QBqBVuM6eGhBv7jgJ6Z7opJ8LbOr1s+DhOu0t2L7X9xNGSd9M+pAYGYFhgxea8KIcWSR90SDBzu
GUxJkfK9db5BhQavQos9ZkS13tLCp+f1/rwOFBvPiSIzbJP0y5lQKxbczot+DjzPjFaPcyC8E4RA
YCMW2Hmfgf6HMnEDxU0QboXih7jk5UGtEXZZ1nPd+SKmbebp09KeH1wc4xwh9Sdk8mZSfo0w9/bx
WXx1ATcKf35tiYNN98NQRr3vfT67WuxuGvKoGstJNoSyXJRp9ANEezkwzNMvGRtQjbDu2Cj55bTS
mB4tZJx0OuvdBw9CmMHDpaWg+RjII1v0wpIQfad7MqRNzRFhtZoO5q0kNHK9qCUxYSqhH68tybAh
B/R7ATaRGQQ77ML1yoiqUphfkbcrslN1vOhqk00OlBnP8W4+jxpRsL3Wox6Oqm0gxsR/ZoMYb6Ch
z+oqsG4T8WXYnMCSBB2fkv0ITj7C4foiPhCGT0pCUUStZjXha9eWqCDbPPPq6ag3SNEgeYRDclPc
G5KZz3paQaN7KLA3+MnofJ9nPtBNr3zNuOHLb14S2y5FShcUt+Yzy2LeNNdkxUVMM6DpoxXN0UUS
Ke6IkbF8fAXLdfVTuQ1ipEwuT8YeBct00Ay59QXuWuhSegMCSPPIVb2utlzsuA5WEHIP78b6cfiO
P0wo4rrF7hryRA8zLlIeUSORdbojDi079quMXqkAS0GNuit/mJZegienEjYDkNhToOEMySG63Kme
4an5HhBGswZBUGPY0Cd2uqEBTki9xU49lQm4WUCFRG4jsXazRGcm27br8Hot5pnxXIvjB8A0wtZZ
thUecZ0qpNHJXe4km7Kb+3dY8G8rvFPNrKQM2w5nm4wc4S9wrnzJQhgkAdXRQpUdRTiME0x4LJoG
WxjZnTt0fxmFuVpNbiQf6t2Pal/utrJJXm+2W0L3y/1i5dZxDHuCJsdkSgwxuGddSp8WlvfjTeBy
hpjOdLmltRFsXuODpb2YbJ+VWWyJSny+e6U7GZ5bJ/vnDG5Bf4CTgb7TnVYBdwRzi8qqGSm05CS4
f7AJaPJ7gA//68m7EtaVqt26ga4Ss7Ba4A8972GHwsj/qAgmaii4Eu4ca6y88uL2odU+bI6IVR0v
vF2bIJOj3Eiu6ArtxGRhp8GT6+efvj4QLyoXN9XSI6RKFO3Y5FbnFmnqZ5E+We2TBiWNGB1yVxGi
GPe1KPRk6DxNNz1bBmWIMsFIDYMpmOqregchtfHkr1m6QNYrliDetbo80DPWxInOk1O9AETozsvP
dRWCER++45oTvuUPjreHWaUFVurtmAICPQQQcYGDEYJ6oLTHeD6W5nnQWtDBXQ7F+QTb1/XZ4WHQ
72r+UAfN0+dLLZASfgpR0QutJadQYmBMRqt0b+tZMjmXVB1AyBKtFdBU873J9d+abcA5J3j4gJOL
CDcPlxxOUk8uQczKrShvCozv/uBkyNt/1tsRkpGyXzyyJCu32PdMedn8sidy+2f6YjDMbR4F8pHn
U5oJtG08mqUji+fhUBmwvSWTyX9gkMyZWARBPTZHL/Ax6b9WlDVP22DkOcaB8zCwCW7STuDDTIIl
/0C/6bg625dgRCSNJziIR84RI+3F/FcgrXesOj9ny10BpCpcRvjKoKkBPhu12h01s0Er6z99Hpv5
hcv+q9NFn5VD1CV3FgHOzVQj11kDfFRh+5LLlPU6BLQQK9xWVJnBFH9nCDppBZyL1DctQg0mC7c9
6NFUqGnJzuN+ZshPAwhQpchMwAH/fKapjD7epwqpP5DTzEkYZID0eQvhYH4tU7UxWtj3VLPBlEZa
P3vIyoHXIqBRmmmZbOZu7Q05Kki1rToUDEPfKsSf3Iw74iErerEatPQRU7EjQ6maJeW/teuClLnM
8gAeikcXMqmCWWWAw2UuJunWor7BVcW7f4rlELFDpsJ+1BqDR42TOK7cyaz04koOVbrLvsHtmZgP
5oR5UPNi7Jk0PIqk3YYDjHiyth8DnYIfiHphf8Lod2ZhipSGu0Ki2NlV5y4qZBB/wnM658Rd3dDm
zbEa7ireTtRBHNPgqLN0IwHvmA6NrTMW3dCv7/LxguGM+vYFw+y74YKcTaMc7Zs5iDIY2G2AT1PL
V71oR8eAVU6SxDbv84QH15mg75zcrEEO3fSoGqlhG8jQKToo/9D43xBsiB5FUHKs6oMooWBiFb9O
sEERnLYQHM7rKq6f2BdftAh4YkCTM1E0zJrloUO+Kwrjuo+c7Cme7rt5ri4PlM1nhXiIPhELb6TV
W2LLrjFnIkv+kDby0eS6E+vjXCRcxfVyWavIJPCDXvjkIgU52/H5WmzEUOCgWb+NiMiz/urAZrsA
U5QW7rVuLNipm9yMgE6w1ZJyrkhINqysYZIdY9+20RUZikZ0blsaQiJVDu69AmEMbQR3sc+0fSP1
/3i6gK/EdjBGlM5F7vkR1ghCVTRJPSPCUTjiTPYNVoAxQt69TLZvl9sKLh8ZfleyouPTkG7PbZcX
OprvQaELD51QGya5x+evXF+b98DGf/4SVv1fgVVcbtqFQFJ7NEvpXo4iLKi3YjnWL52hThWCyuBL
oXs4xUTtfO3Hu4HhvBqgg3ze06LJ3kObw84mtSZOb0Zp8NkPBEv/IKqhU5Mt/qA8qce64nk00CQ2
4T6ZJ2IruCBUe4fSoN5gbi3z6vuiWK2SPzNlcFswCxF2z6jw+rYE0ECpeXuTJYi8iH0PRk0B/JSn
XDH/C6QCVQNDY9oPYENnMr3buvLUqE6NJZdV+r6zhDRxj61jakuJcgOTgMpdqUg/f+ZC9Vf2sTS7
d8+duRaBIFu042vLI4uFqECWSDFtF6eeIm3rNsu1mVv74D7eghdCN14S3Tb03+/N8Ss4dTFiJgAv
qv9HVarzMnBB6KF2TXDU99VAfApvDn/Cp9KChwIWnGuay3ZcN3Wuergf6En2TdyjUWFp/r54rYBS
Iw98dxQcgjpi1nlI5SbHZayO+J8EsvbFVpvhw2DsnSnoMjPtDG5xzBwojgtSOGCZqG/EmA6UTSx5
FPXgcjN/CKdeaCNCX8VZW5wpVsNLVQPww8TtKgil+7MpJHxCg+7xcQu70YZ5uXf87Z8wqDf5pKVi
79DTtw2s2HM0x7W2txguhp2yJFeYTiCKk5fGMREXhS4Qj08pCfTVtKI9xZWPpcDKV+SWvC9BbyVz
PpsCdour1KYNwBOEmUSUDHoB91G5lokyuGuhoabP/iYpcWWmhsN/B6HkeyZuD11rJ0JPXM+7Qmdt
DL5yIkmGyhYmY7rrcNtjZwG88gKzaL0KCkWikeq65aOcLpmPTG+Rz9b9kp8alRVPUB2cC8JRXJtp
dmFV8OPnPuZOTwWhzPqc/1Lpg1vBjGl1j9LIrEyCPnkSPZ9YOera7WeySQTt5s874ZBWTos54Dmh
4qcziYq1Gzm+o6Ur0zMuhgoxL9eykjhu+dmWqTXZKp+L4lEOSagLueC2NDF8pm+CfHvq89xKFqMl
+g/urB1hXmCwJLqO94SLm3grDmuvdfoui0BeiYHd/uTt2VNV3VnXaLMSlrYnuqF1BiAGN7uujVPD
GWLS66ttbdHzCtVhtw1saNRhgYr3f1jwYQHXll4hPGXMHRdMHR6MMekpdL2R5F5a5T7d/vggFlAL
PNTjssq0stl0PvnFl7kqg//33filVCOV95H217etvPRFdl9VnUmh7KOT4c5P+bFNoU2HX7RLJNJN
b5aINf0Tw6WXBrFiuAhNs8EXfIBGNtfx6aHb4NZXCoSNZ5aqNj4rx1Hdd9ZGjyDUItv0g1n1HCAw
oYPPJDQmMi56oRJj8+IMNvfM5q1jgIrPbIc4xDP951mg0KOpea0REvvYIxuAfo/eq5dD+tqDtn5H
t+5003cJnSCpQlT05ZyYRnqFSUJCiTrkmfy4u/Ik332yvuU3Rr83UUAi0u5APuzKhmTdazEUIpFv
hv72STHWETRJ7LEAKYzsFuHR5WfueFTl6UHoATkHMeXy7+65ufK/SV3ASLUKEjFSTkfArNnlQKEa
kGPJcdeW0OEKkmspFfgRGDo18/5B8WnjyZTrK1/ya1xBRkA76EvFt3qQUGaRUw3kNBdc2wdM7tV4
Fmrvax8bUOgdRawKwH3kPZEfK0irXyUp1+UhXyUB5uAHDOThqyy3ADXxXs/kgULbgYI8w2BGCMXI
GeEcorTQ3Er5O9a9L1VjcpNIg5fmxS6Zy55/yXC0ORmV3LjRL/Z9Cc+M9zR6xkiqEy6nS/ikG7yk
PMczwkfuvGOs+EQAeho4SLqLeMVe/eFS2s9uNaS5ec966NH+3gKcw4HNQGGAcsTW6U4b5cgFxzGZ
cX91+ldbKvxehXReaM9xg8feFuYGn1eopDrNfOfTynjXvP0Jerd+xXFzZjkPVcJDSlWTMpnrha6L
O0u4rIAi3xSKDYPVRBMWfDbEPr4GEdMu3+qh2cZhtRMdXzma2VuLoSGyLIthWpHfYy2fXZ1Zsleu
XJD8kyJUEX1CLuJ7ESaYrRNZCsLAR+/8hi8w/PTCqYIFDo+uAGZD8ZUCfiCz+2YHOChk/QE1C/7B
6/V/W4JlGwDinMhCXkA1P10u7gS0Nl8FmgMvZvh+fSk48is8Jn640uipxQkJ+8RLO6H6oGOSawOv
QEB2upKW5JqHdZ0tXdwGP0IX55eKVI9Wum4FgihgVSJEeJeF7I+6QSiUBrnZgONTPL1WpWZ+8lo9
Gzh+lcyLG0V/c2z74moDR70cUUwy3SrBEj+0aKOrgnP55cc9d84mKZ8cs3/o7WRijwsUVHHj8glj
MQZaW60xAvOtcM9/jlIIbK0fyFRptInYegswXXD/pFDMUZJamqWurPY/SMpeHgl/7V/lCj/gViBE
8RLTs2u2TJb2vIgjUQDx1rnRXjzadl9cDhIdn9TG1b9Jx/Cre2yHUrVI49YpAPzLtxcVorg9TsVH
tTl3XbsYBLN6RPKzvuwHxJJQqAUqXvlG8rVklvQGqFEhXmf3Iz+YgsXYUItoYHBFrYzgOyhEhcRt
z78Uez2EOFil4A62YW/E2q0KE9HcNkMlbKqwmYj78VUbXirz9+EBelzcoPFIunxJym/QFRSCYClv
uZkFHbwn+0Q/F2wRSBxhR99WzjspKbj82YslyccnyNWEp3Ql6R5gfWPIeXFZLP1C32653FPTXVVj
u9eIztpWXtlv4vedkbUwKMGIwpi9O2no9dXfb8O+wAkaub5/dIsRsJb+RxUnJfE2nBmEAl5KhLyQ
Tki4C4nzSncgeJP1gRWZF4yEb/hGmvqyBMN14gUXESfSaP9quP+BRrOcrrTdXn/b7qlw1hxhvYve
rsbwWgnukjsGd6X4xpWXVzFHhW9LpWizm7oQDILMxraAaJM1q1Arr0cO+z7zseQzHNkYtUNfDRMU
hoAUHAW+0Qxd5h3lQhelPUTdkhLQHwQKFmEfftLnwhO7eJgG6ONhg6stbUj5lqBcgujY2nkTchzG
gIYtj22zsPL9pLSgEApNcpAZqyzFyXtk1mPE0RyIcc9daXaO/BmNcpGpVHgKslXm0JtozJcM94rt
doaJxfcGyQnp+3J1aDm/bmGsfrlqSSOx44BGm0MsfsQ82FIFM41j/qyzvTRc5btc0z8N+Dy3NMwn
q773JU0+2tXkA8WWfU9ASEUV+4ok5wSr3QvGE5wGXrnPNUa9+B+jv5X0LwjhOWcUVhZ7bPD7wRsy
OV8c+YUjlbcw/nF8TDLU1KojNzWJJYH7rA4Obdoa1joY0/H+F8xRSCqp2MS2Bq7Afolct6ypQWos
frZ2PEv0Mx5jESyJ8fkbxiBg5Le6qalkv4+dQpZfUfe+F7Mo+2mSX+NaKWUPk5pnBCwOu3QBn+O/
vKJnNk0CaLp5e0IEcRg5Vr1ECVTkXitJKg+0m4OXv/aTqnV2e7dgVqQ0k5+Bh2kT0UDv8LluAZMh
BaxWA97aIfV3ZgeIazdlBhU9gDwU3cH7le65pLYNglhGe1eEelPBfpklscdfqWDfqeULEGrZoqhC
8Xg09ivyxxxnSu08dSXIPYDKMiYOiXyMkCbsnJCPtOzunklBgSz04RwV23uxBCOEuQFoY0zFkbLo
K18mTwywInEC3fgDjVFVwn170GQ250IgMCokUwHNUCaBapQtWwMmZDTJYTF8EHe5eyWArXKdFAVo
RWrAKbslNzKbDxetiQIMA4e6ADEmIvIAufuuXYUqbCPMedkLLgByFWcszbDwso//0w4a3K6Jq7bk
ThPgTEKrSOweZNVdsavQwVGrqo8VUKMlNNuoJIpCylygH+uYMdsoToMop6pSV3LFsm5fhIB+6jFB
KqDil67m4eVMuVsF61m4guvgDQb16J9ELSlmSeBkslrlAYJceV8ymcpIMYWPezMBFKY+UdhTT/67
zwf0xKl2NkDPaj3lwo1RJLgeEVuG6GTGb6qNAqosQUF7dY6lk5WilQCC92sAlJaLCZwgkgdYSp8T
21zaEfHQBl9nCShXdRZDPpjv282uB4vSIJiyvW4zr60UJyjHWee/x+jKF2Njqd/16tNEea9FlyFZ
TQKrOoeVOsp38R0Sl6WMt3DGJe89PAA6BnIjj9NbY+e32UKAR61TuuoStD2DKU57/BSyMMTDAPsf
gc4urNADcmocpKU6YdYtYGWjjbHKhkz6ATNrtGYoqbnO2ibyjrlOsc9NPz3aGtqPfLN+/oFh55/B
Fr7xhK+fp7DphvwXlCq/DV4AsCDBdauD4PWJHlC0sK4fMxXzjYaxNaRAl9yyZUVLmgryNqU71fTe
Cyq33XmXq2zFgw0gpnAEpduNLWZ9kcZqevyorBqrNLeKPvwhuKEBOdH0GaIM28yC4nixVxT7+qu9
jyz3QWjkpVT0CNApQdhvcfr+OWT1o/R5HKShOWX/7nx7kAX1wXDPnCvkvchb3Spf+nSMkhHLQfGi
PcjBrBfiaeRIzCEJCzpHg3r3zr6hVnMRNMrzrJwoAEQqWozHFp8JhTPLo/A8jGB0FSbzwPiEjvMg
3cWzPckZ8thcfeuICDtzXMBaabhL8IV/vTjpf9ew6ZYCSMV8pcP3aXVIK1/geLga6mvPF1injwS3
s/V5Mytss8EWUC7eLllQMHYpWKEFEekva/3+LhFCJ/buctgOXqFI2UFsvEpzHtkFTVmWIX9QTKvz
WatLF+mlB3BFKMWmSfFZqF3DKmD4KwX68ACGBpFZcKaLvpCgr2tIqPOWFmanxQv9VFDO4/zHik/a
BJk1FQL7v1sjfswo30o4UZY+lJMvTsWaXAm4FTtFVIxWRmHtlVgNi8gYTlXXFMpAjPBcyx1ojG8M
gm0aZTpC8JkZimSjwrtneuQulqGjKqkbAMzznoyn15+pyOPa4J3Lng1hvaDqCrFT7k7rSpDO41U0
oiYeWwGYDVeGo7fZXC8chBvCy+nUDRUgd9DdzhquNWxak8zC/BZxL6i60lTReIlAVrM91HTB5WI1
atsgAxrzwBlQE1E07gNcch+UY30h+rKjhWraw16QJF+e7k8ZLFi3iq331srIZ9XPwdxZyxGstF8Z
i+CeY9AgiyGPQDVBZn8KZa4BQ2I+bC4fO/WfZTrf9JSojOTJZ8T96U/jbg/oAViw4AQKwJZPmfgM
UTa84m+Pa9E6p3iNmkJhM+/gJBJiXA2IYyfuzBP5AebOeiqNHgfUvh6toup18UG/5gLBjMmAfMNI
X1GkYXBeZ6qsFfimw9wd9xlYTHHMbpRaaR3PxERg18t5LjdVs227/EY4lvFzmA4PyyDuWd98jZS0
FY6iktQyGsglD0DJ0oAZ0EhoolnuGMWDgiLwjLm6KX/1002J/ewbCkZCbbGXZi3it/rGpDEIGZQu
dXyRYUn3GmKPZ/DBcvIvoQ17GnllIWwliWAugS9ZwQoG1jgizYHuiloxWidrCiHxe5IbjTf1XZP7
JWSp/MmDR2L89XcpP9XItXvlkNq9gQXnJqS3QoXUXacbHXTT46TC/xymswRjTPEBdC5iMcl+xMo6
hHjCot8Cno9TnzskYoFhD48r0mPeGw26u9D0Jkni6tiuT5vIsarevk5oKK/H2kGoMcotkM2Lbtkz
L9chj2zZl/uz6BFtsZWHmmJWRQsB5MWBU0PlR59Wx2XAmB686c9iC1d9DnaiEp/TNq5qT1CIj6dN
eXebQhciY40iodmjWrCXGvVRyRaVdpPyu4pepzyQ8actMz/rzB1o4jBleOZo6BeOX1Sn8DJhKfk2
vrUQN7bJo+NhqxRvMfHEW6+0L4+hRJCrZUwjl1OLtm/BB26tnvfzSrbt6GM71+/GxJI9tY/I7hs7
IWoE1+RpRvfMSaSIqO+IBSxCKPr8B0Mg4qtKByineAP5+uFMdy6hpj5nSv3eEbRJysi2AjTmGZKR
juE3tzW8Dcc1Z9Zs5XtIraMOlX+V7Z/Ls15cG2uC/EtsICMNUVb6S+3Em+erbSPRBOjLJjqKY38d
s/91+qZG6kiGxgalNaQk/Jf5XJj7lr/tzgGDl3BAmmmNeB+ov2VJlQ15JoiBwc0X/p2aDKf/TzhF
+LwzRZlOewz1D4H/APbGmdMdZtY4V36Avn/PJm/xPNARNXgfg3HnEtHY4jbLbjhCAkqSlgOgXhQA
FAE8O3tDEs8Fk27f8uItESABnGGdSI+/+kU5iCLnkArOYy8r/m3tgtTUHDyN8K16OnJietQ4HbDQ
t8NF0IADqzkiPc45z1HGPtciKeBhb0B0Pes8iYrLrS2qEi8/E+QVXVef6f4Zb9KQkyIOE4BV6B9F
IgmTHWj30D/oJZNni47wvxuPjd9mW6vN8vTs4zUKpT1tizUo7dRhqbm3zPxd+lylMx4rJe3MZo5R
eQOZdugbMYeYCIyPhBd2diGrfZ3rUPptt4R73DHsKKZeNqS1Jb0xj8+TucBgfCCwN26cs2YC+Xov
QSoyUv7hCUSPJ2VFaekWLfockSTXFXA8kz9VomT3mMOGFzPUNGY+5SncNZvJ7BfFkLZBQQWDwrJi
S1xBuLp3PxyM9OIDNBITms3+ssZygFMZMtqpINFLambtK0dAOHAvT6WVnWPyv97oqNoDglrTAtTk
085O18XPPIKy5gv3ANwzWpyAXBNwKpu0abwWJc/HRo8G2h2YeN1w287LknQ28ZDUeD8J8H3cDbaP
Lf8hiUDKoXQdiLpkAeAI4ytYVsGpbgRRq7Kb/+vXtSoyN6LCXjxE+4WEi0AMjANiT0ZtslWbHIsj
l0KFEsGn9tNTGfCO650/dbs3qH42Bx0iavExQgv4cLwnYOm0D9TiSxe2pXtzsicPYtiHEI0aX8xl
wpa/N6/UI3zwFFcDygSTkZLwkmUT34vjingyElHjgnPmI6x50lM9S+Mgk1QC0oS4p2vGilSg8wlh
6Z0nsIUsSM/3bgwQK9k7XuTjfdrDIM8SFhqKoCGBTWV7jO+Go3gcQh0w01YU5G4xnJg21JHtVz0E
m/bxGCMQXXnmhYakOLgx+N5iNXVXjcFq4f6WHWx+WFkBsRvScQos2O4CqD3JQP6VtgWiZpri9Jda
DE18H6MDAkC8lbTo2n5CXTZ9k2uBuWv7cOjbfCsEJBjW+4xMW7MFbnf49+qPLLt3z7BSQQYxtEC/
5HbnuaxqhQ3a+cHxTpuV/p+UTjg5e0mE8MtEEW8CHeVCHovvk0RDoHSKMUcOXiwqOcA7GUBrpfvm
ZYU6H/x96VPmi7y7L9DqZVmQu12KA14BAC/nekkLa+xP9lM7IrWfNNjOM7U5PL7lceR7ADaw7XtK
jxQGSFvz/dRkoZ4N6tx29vECR91tkNPvV/HqaBcE0K4hDXPMKmqfT6xfAjRU5jcdStP1HraGxw5V
7Pt9qtQRJrItZl8O0dHy8sQ5rNof3XC/7twIb6KprNv6uaiUm2BHoysnu0GHRk23xVsHMcGe00Q8
tZOyXfWbpUQstD6UhnMQFYSIA/xjtC5FbUomrnw3EP8WWgzAzn/EF90HHY56KvGNbh1FrrSySbkw
FHtmWRGI1w9ezYnvO77SDbHGn2VOsC9BexfdP8qr1tPv0dNWddiVPJhHLX8CyUxhM+ljtQtBPzCy
XrcSZqlzsXJh8Ppog7sGWSvwcNsFWff6sA1h+3d+RbufGGJx5SaOIvV8FfOLKKGi16+/qFD4Addo
gtXZrk3r6SRwSgAGXGz/5/ZIbz3W48kkSTO5C5TgvzLvmIg/JqagKuiH3wjr2Mkzilg+xfId6T0a
dN2H9Xx2VpvzId4nt5DIzcK754wIa+ibTXkEMbH5sjKndUzjXoXY94lrROg+tmO3CDQj1e0pYg22
1uZ2+GtfEyaBzMDaSKu7QSYXoh405tJM/hkOAGUeB545iC1Aghgve83w0mqbrinAoGbb8k4Ym6F7
ZbbmgI79iiIre0ORnORKrUgOZ8kAOx6TDuMS5p9/50ec610+JyNd7zj8clc2eYiQVjvc3jIrJOSO
Fse0MkSBJaxUozpZGBX3fyQzI3gsRPsCi1N86bHVmUT/H+IGuyBmDoX8uMJJjXbrE8FRndy5WiGF
Imz5FCcbLceOF8O8RlZAJJKwubC96L8Pw/SU6ZEJOGSvyYDc1nV0Aso2CTTWw61xgIykUdB6N/I7
Nw7psbFghu6r2hbN2dBTli0mCShbXwos110bAly86QziZfiS1zFHqWQQk4vE+6D63C/aQfY7x0fP
EejnjyPdZYrTeQZVpVQ1RRBY7oSDXynoy7PKwwk8s8mvRy+ywGigB7xc+vhItdfmk9i0r6lOnKbB
qoswNyXii647IzrLUmlvnb9rJ5MhZGPEnh8Z+y/pldVgC7m3Z+OH9TpnuufvoBvM3wq1JlNGdKmf
UA7UVI+STjiOfDGT+ZO0YPkGLdBhfwmX/TQPITIFhe983IvofTZznBwPu5YI78SMkPyTXGgqn92z
Mz4DYC4P9QYAhh+iDF1VBpoOMrdQfDk/jBqXd5VgCdXA0UxmHnEzTr2pufk7uaRMTUR0F/xSXoNk
p2telPfzPiPUvT7WEOBUx02K9xikk2i9g7lxToP105scgggYXz2iduqqLC1Mw5fQZ6tU7yIsBWYv
I04pE0s6ekq+DTY3EF22BPXrdFjSBnHk8gaVw2UG0AF8YO36md03gker3r6+4rdKwwGT/j/HzCE7
N0pYHlUlqKDhRVjJXLh8T3vdP7ZVXbFLl1VKgFnkDKmGTtFPI6EJ7XpJIHr397WJv/1hNkJlbuRD
Zqc5GY+U6baf815EC8PIhB5nW3Z77IxLIe9okSBOH16tbid7KiB5NqLTP+wcbqe5VS1eQgL1eEnu
7Ec7jG2c/86uir4yyIk0b2QzBnqiGP96m9iSKeR5Cob/pmmT0myLgQi5prVZ/RE7cYToNZUVqW+p
XS406LDDR12sWWkFfnoE4oK9IaemZpDzMMBpca+ad2pPK0DmNvTRcfRHThBADMY7gt61lJtXIhjr
4ZUZWqlYrz00nQIvXEhmzvz6YRPVeJN7ZlUHD5ThieTdrWI0h4A3V74/ryLhxO3CgGGsowquxCI/
enRqmn7LoUmZt3GemapQtaPoXzQ5wdCryciTH2s7vaqH8bqn/Xi0m1IJhgmwwfgpB/gKqxzblB4y
8gNsxpNQYaOgcbZnTqPjXfz8PWwsRTfCQpfPXNIxlyqBzQZwOkON9S1Uni9d9ZnlVIUG0qtknko5
oK2t4bD++rWCh7s1fSimGoPGt71tWtwrmIzFL3Uum4gkv+4pfazowucwos15LWpdiJTA9Ffg1EdA
ZtAQV6nOnfCyz54Zonom3+B2ivgWvoBT6YcTcGrVuUzA7pxi5Bm7oF0ssSmlprfysiIhm6kQVeg5
TCXj+QYc8BkVYpHy9wzZupEqXIwjj5GnIG7FUdBZ4BqmIQISazhqB8kNUvmsTjvkQoyBKeU6LzMJ
FrLGoumgSClpO5s2c5Sz+CWF4tnTMaTVT2b8QqJZa8mFZ2iiS8gCsH+RooBqYwRmgMMnou53R1vp
pwnxwTmBFCuY8wWa/3ULHGkSFR+LW6UBp7OCqG1ti3JKox+bQcOc2Mg2FBGpuFu7pPdY7pOSnGvl
w7iAG5rUDj9IvZfeuJDgQ+iq1UnzbB0q+0/35iiobxlVes2hoYqWAyxPwC5PctcilBP6OJreGRoi
N3VqN4ofjRJtWJllvruOIgSBZCnDbiWdc44CF9hYMJq3iXXTQAZvSHREm1ICiMkOZDbV4OixT7Qm
d+v3JRpYzrONmNhpW4uddwvxGMfnlR+VxjumteCBSLileL2ZycgzA9GsQDo+Ug4HILj1X34xMt3V
MXjP3jKShYqxmqHYK1MI/BIayzFwudHSOetkbjqSG5SaTnP3s0EvKt1jMl6Mo1IP7sHC+1GIkIzQ
VNX9F8Z8eGr3Pa5mFn+fHUR0ybGbeL2cDR4RyUdwVEPU+JT+x0bgBwfu1Z6skT3+cd99JuPTVbur
UZqrYG0J9Q/JQ+9VoLpjnATWda56oxEEdzD9un/KL4vyV+65/NkPjwDCIaqMJXRoUbTqSGagAYWG
8iiGEhErGbGfv9nWoFVtkqfhqqwaSldTF6FDOBchOWg4Ztg2Bl5YRtH4/L9oI1T7BGmk5166yng5
u3kpqg6LP7Kiajy0ymNw+zAZK0pm6lUyF5LoaGogAbQ1bHNsRYJNCwcFO3dL3yLZCGwqb/Ig4cdL
1gqQUpyp4eoXm7HlB1sXWGLFANe2teEw58ZUcF4MCWIUlpSTd+8cfi8wmpv444OJQ112eFjviOYz
mhmoas8Lv1RokEfEvAbCO80qh35/lmJUg8KTV9bTEOWPlNQ0613bFDEBKSK+ji7Fqm8MDRv+6Ftp
XnjuzNLstr0lXdxKugs+CIe7grZNmz9dV3r5T/F/ST0ucQuek4/LyZmy2WK686NyYk3IzLAhp3Q5
IlPVtl3k1o6aTRBTbiD/MuUq4t1sSVVNs66BEm5uOsHconS9TrSIRmvUctLkUjtJkpzzxo8cI4O5
/dG8MecEyWXplkSDCe7QBMEXw2+Pb266u50CJEhsubF6gnpEdDX1/4hCghiNwHfxDazCc7Y9VDGp
P+0GrR2KEIx4ixfALz0HTkkp3ZhUeVZiCPSmt5z7HWA2I7/JK4BQcbXfqI/ycbIYiF5MrW1m2nMm
INsyetbH9Z9vzzu+7icN1PoUq0qa94zOWmtjTWTuytydJx2Vpd3Bd+26HrkU+6YQrQRJ7SphlY0a
C+YNvodRYPSrMHbyW2NXdXlWhlInK0R4NQRAv++SyY5Mqc5iMs7v4rVFh5nzoPHMYrgHI8Js1yN7
+nO3+Tsr1bOZRKuEnk5ME7rbKKOjPcUIqPcFiRmfNzctJ2/n2nuE+KL1uFnaN4sI2koHzcO2XxAr
8Y2BfK/6d8UsW3lJyLlx8XLZ1JFE9UQ2YHm+ANqWavYet2In7MlbNAX/Zf3fUF/rz+EGsWmy1PsY
i+HtWKmyT+J5B0tOpv4+V+9GJd3ELZ/cv7+U9jpFNybtL90jGATXcLtf+xZjEPZn66ezoGScOGGr
asSNVJbiBJCVBuI15b8E/WuM/zqZAgJtUszju039ODC5Uetznx0R0oaCiJDD742+Cun1t72V4ZJV
er56Q9tPj6p5iD8FUxP3OIisf/aVt954qHe8/z0dxkCegw7HBf04e7x6feW/0kAVDUn4lhGNzAnj
ZaXWyAlHmSfE7rgZUNh554Cd2jXjrZA/mvO6TP3XuT2i/s6Yl6wZs9WEGfzJztN3TtP19gf9Pr+U
Hj2jsn9wNajV0quht5ihe8D+yTGD8YTJdNFuc5usGpEEXqLilu/2ti12NZ+CUgZObZwD29RpsNNr
fBQ8LL6tHUVVbJzrUe3aYzppHDrLeHb+2EN+kxduMSkITNL+05l3srr59+LISF0WOD1scH0HN1oh
VTAvcL9kOeAs9QbaG7pAHUSuPJiUVyiNPpIv8uDs6DiurawiALF1dUrDatAJD+MlJEfR3mH+GJiY
E6YAOubHnijCPeqMEUNpy9hwbp8FM/I0S+lIZ0Z7ERYVpsSqQHY4wi5/CqrFWmxu/9EqLYQDfW20
tE8EWOU27Fdk2+u3e4WTkJQ/EC/0ckahbMp0cr+rzvoL8g74PWoz/oguyv6PHJWTIqQ8DMzL57Sb
LDGpJwygwn5b/unamr2JMkTQhiUAxc2R2pluxGu8oBofx/wHowcDRzX+/Lb4YYbn5fSs5UwScUwd
dcJXGerpiP2eqM5rlGg30VeZDzeZlnFtyLrTa3Tdj5TZh1xK6lmhYY5CZk0NsHwDEper6uwwW92j
10ffS0NBqMhcauHImcYM5DPpwClgCCz4nrUYzwihuCMkbr2aUQFSfzcgddnO3htdonGi/XjyHqIo
hRhLdUsq9fmTBNDBinTgkwY06AApfpm4fzUQaWwX0MbNQsQ4441yD9+WLVkHmkWIzO/RdS63Ju5A
neoH0IGe9WTyyg9RPeG9IuNFsty5uYOgvqrrenc1NZATMCnmF8ZEknNld3MlHvipKPtZMJCEoPFh
+Q8yestU7ebPM/W1dQ0n+Tcs0HrDVdQKYTt2LAmm5kAgaiKtFfoHOiWSjK3GOQ7RC+yVTf/8vC/g
rretEKt6oUjv9hKRdiKJhL45/LDJXyc05ViXGQ8y7gQf612d1UXXuremuZbwXKDryhOEW8Ukc4Ir
snTnsl/Z+7LeY8f8vgn1mrCiOHKhqb+cKj0P4/L2HGZImCy66o7rx99jK5AKfLOY09kddayHYPNn
KfnXyB7v/9fXLr7AkWqEHnyX2PqYR+UY2UkcO/JNq90OvyNYY/iD46UJeQh+pqi+vvgNi95hHZnF
m/vyIbYV+JNsODQgnkZDUye2R4mhuwNkmX9tzxJMdy0k9b9VL46v48a9iL+9z53rc4rqxGfxR5xB
zfItBG2KfwLOVIR9Yy14VIubgw8imb2d5j9GMun1fGgBDgNthZjKqQnfoe5jWrwtiM1oGtPn5zkj
pyG2C+NQuHSYw8wlp5Iy6PVyleOa491SH+Em77ZWH3SXSedkFQqKeTi43g9lsvqqNBDz65CKeSTU
7bxBtpeVjqvwI0ILgDYQn9tYnlb2E9nzLGByRhVNF69bEGyf2d2c6WtlBRd27tugVE2LSxKpqdMq
DQwSzBTQEWTnReQ6ECyNo0e3GX+5hs5573wW044LYMkiq29ueh8AC8Wo85SjclPK6U8cCCXhwBVD
Z94nJ7vsHSLloU+ekgGJ2nlkmOURdBI72ZJjwD9k3Z7Uaz2AvCM5WGHgkF9w37NiZSwmPqHfxIMT
jv0L8eaZ+Y3UDz7efmK4O9h2MafkVJSjPfeZeir8Zxjaa6QuIOi4nH0Rl2uC3KXEFwt867oEnnd9
dQ9Puxy1yfebXYjikYgV9XIkq58t3hGo02T8CIOGyVP+Az8H1DYFu+QCrcYQhWulyqL8SF2aYm/Y
vANpTozjq92olTD7pQ1IU9LDhiAdG8PHX8eEDYnzcfXcwYwX2k/7BYmtJV8RriFOxEQy79hi8C9Y
JrpUheWJpJD+eOsi0YsLjdRrHdz5VOpXIN+HIRwh/REm/wjCjxZRIbqLTRZV5o0lb7yGqOWMmFkr
OHf7II0bvL2nyQGlir8Xvdsz1fXVnmWikXDYlngcDt9Dnm9qU/gZmWIKA5U10qMl0gbXHlzaWjga
/PwBh/BK22CLArXuVJvPMx0TrSDvWKWDu/AToJp5lizGyqjT2p2zdlqWua9DPvGi3sH9sys+rzWj
glbzfNEFp6JeGuVlmxX4OECVGUT9L+n6U08Zq/7bQCuvy7zfnG0TzU+bR8tyevr7vAC1QJU0HWTJ
bhjxTzaBYv96y/FNljcunE9vZkIVMOPlm2eMEH90sNSkGgj0TsJ8RuK/Cc3QkZydJgWdq5segXIC
NeeOAbeNuX/VYkVHOAWV9KDgWa9jTKYiUGKXj6bU03L+kgoyckMyhhH+VM8X9HQKt+3lmBbNzZWy
rZrrxBtcvNIjVz3i5lNzQjG15RvMMFAPE6wVsjqpkSVcaLiMUN8DAnS7Csvjd/8mffJiANuhtQR2
H8vWJZ4YJCHti+skt1attYxEkXpLH+gBLxBpwCMHmv03A39li1g8OIU2eWaKWNRbK/cFWdaaGVI8
DLDyVyWOGYu+a66/Wbi0ZjHw9KzEvvS4viW7tT8iwErw3wyBcYbwIGmb8/SlbMFjw7ca8s/O41wY
xijjSnmQZ3TJ87nQXCRrDgcpOXnjH8/lYV/plENUkMxxddfRs+/WkHvaPIoGnhz+GjCUFOfm1HZi
klS2E++i09yyc7a7IijXjM2NzjJHzg3q966wEjLOKICkMH9B/Ru+/DPuYg8VyE+huN8JAU/UFU+Y
7hreAMwo4Lx0zNDLLimoxhuKsP1z4H+eMawBA20qx0Gcpa6l1vjEEjoWhWI2DI6GI+XmdpzvZWlN
xCEa/LaJdvHeCXeSMXkAFhPwKDu8TnXt+N9JcIqZfPNKjIvfeo8cNIhbfgJl0IKbVvPEyJktagOB
miU2nCsmFiDm6gCdbY7SpNPEvcB/EWVOSq9qTU2wteuvHumau6t0J/3Zpd/ewE3Z5qd6YhVF/mC8
hI8L+9EJy9OaFcMMSUSCv8m91tqmow+YxE+gknt1AtdzGhLwyPtRSXOnKo3WM5FiLXa7yVRc14rs
UK5WdYQG0IpeduWpv3HJTLeNhtORQ8qMB5PprSwjBNL9dvE3vEBc7ZItJySPHIkyKl/3IdvfmP3w
tdX40E8y74ukZi0x0zH2YHYJOj5JeREaa7kEb+bJ/nuhFWcDF/RTytCKr+QdCpgzhSalNMw1v806
1S5+jz6ii5H6KKm5FkpltE8sPpE0lMiuAcTfBBBJc9NsnpjE7TdSSsb0J0hIPIxLmMZS6vm1VYJr
7dEk8ePvzzO6E93nZQRwDg3jfSEsr962rC9ANApApUH84EmCq726oHSohwzHsJLPwbajEAP8omz7
lbbCHlYQFpdPo/0Bp68Y0NiVEDusPrkj/nlxANRcENyhhMOW/jNotJ8jlw+aSdwD9g5y3Sh9cIWJ
ElYYnfwNzlgHIF0Bl8cvMfwxSPRk7EwEDJ0Jj+xsDabNjBS7z8NEUGG3dEr8GRkYP1zBJ/wATNYg
O8LRsYmApJcEKKbIFI9Ng+ZPdfuLUvBsJlPIVlvFJwiUvpXXjarzue3HcahRfwJZfI7g5r/aKx7J
FbE3eiz6NjsxQJZj8VG1pn/SrKiw5w0ZSIgeFYQ6The6Aqctk9mZjHBO1YNVHm+6R33ypiz74U6Z
1ezHaJA2IVkAJbmoWDAG29i5kuuDqLcGzlne9xeCo7Y+RJCTsYDgnfqx3sOWNZyjZVwXOu+fI34d
fyBUR7RojJq6S0Q9hVsPD6v99gmZsoAHEXHumgI1yUxsLHdwnPNHiVPXTJ2IkXFM49ZMGMCTgWvh
dfoTIV+Q7IsY7b2hl02zL1GVGeybRFWq6lJvLEm80SPGukQhSAPSXxNMVeyf0cPoI4PdRuj+G7E9
27XM90tnosemPd0FIHhb9136jKjmSxlcS/ns280BvB5jHYEufwRvz3U8NXhpvz6KdBYjdwdWRk+Z
7HPgzVRpazwnmURmnFszk5r4mLmkX0wmS82dNXBWjKD8zGxZ9aq77rLJIrtDkcPAwrWkBUnd0L25
+n4Hzt+WXKqG1VJswu++CuYMOlVUabBoUHnGguTTv2jdZoWSUsPZJCN58U5ucnCBEBnHTUXoUXk/
8ETxsikr788f7pQ3y2+Segq+WZLiuRrM3l4pERsNIbLfYIyd9WXtNeaXurNLaH2+4KfoUbDs+XH+
VVKoplyoyu2MQ1HP59redmlFR6n2Ozv+PaXyjxiNtl3fzTYKKLu5slUWNYTXgGQjIHFWXo4yfFeL
fqOGwTukLj2J70/z9yfqxOR1tmMN4M9AA7ILwNvzNONcVDYCjQTfFN+Tm6tLhLS4txm341U7G7NE
9PoBuSMPT6zW4LKBv+KJtHK5LGx6vM4NsLb8R1oI6cb5IEoLFXJYcjNqosRTcd2FuLWVrEntVWMh
Bl8X0tX64gthl2jED0uKMq5nOTaVNDPuLhlkRt84zaoM0avAeqoyb5x2OhD0dXk+icKKZS2SwHMd
StmHgYTwkZ93UseR/SpBTypokCEJ1b2FxuzHK/COiX4khw6fXq9lfqUlSm0HxbznZ3HcsogbKR6U
1viMzlpCJrSUJyqWwBFMyaxdYOzYXODGIt4V1wqA04Xv9P5Es2CIyxCxG/s2A5W7KjNMw5FRrmPj
19bHxJoWKv3jYUn+j67jx9OL3zexq19+iSUJzOs8I7Q777uiMb25TuviqZc+hm0ceJJP8g9OSPf9
X6TNnqJZHVVGe7xT1Gjr1eHJt1Oagif83+ZfpEFmg+0UwOCoxnZ7LNYmCkmbtwk2OsuDhfCWB48C
2VOSolaMOS/a5PpjnycKn1qI9NRKivNoYfSDzEcpvf1E+YW6P50rPFTdRDqmX5OZUt/xnCvKCKGU
9RVoLQ5yaq/5sJDDExpg3GDdFpeq6KdYjO/f0srO/lMIgMQz/llTc8tgSmcldGaqhbGUwLGzs8qz
rEUnbPlA3YlCAbnfkeggcl/Iin5ZhyQRwNf6uc+LqDHYGMI37wXIqKcpDZ3RXPdKq0ilj4C/n3hu
D/kQjVxVevHk3K6vRKgIP02X4Ow1SB2XSiQ+1p7l2QeFl7MXqSX4pV6i7cI9MSmiZ5zyPK8nS7OY
zWitKEHY/w2EkspY4qDhFsbSNnX4M4S2wVHngO4zW+pdEOMHImOsrRdct92chpJ85aVz3FnVmAH4
+RnO3m+sCijWwsASlFiqKltq+u7gE672PgEcaSawEcR7zQwzy0Lp/KSTXTuaTNX8Tfw7SU1XDLEX
QRBRcLfM9BaZsOloyG6S7r4vXzAqcTpdvSzVMUp6RPnjoPuePjASri7OMWxuOutd0kQfPkKZ5OFB
4lPGlqx/c6sdysa0MyQpHLi8rj9K/AVAHgpZhmseDWPaqQpxZuMRSIJRdwQV4X6UIge+Z6Gk8Pwo
DBLv9I2xoPvbR6TclsAX/kLXmkoXuoK6VjD8YzNdZkNJ8QIYYxlUEZZclN8DmBdw4nx6qMK2y2CU
MKJ+aPgvBRsw5Wis1Yv6A7wKhTQFsLR+86eym5lZ9mgGaC1myic52ceC6p4E25WSSzpwLt/kqhV5
pFsGgu+GJHgBJdbbufjBM4Jqwl6BrkUzZDXlDrnGPjcy05j1rQQGBmvYWx3V4xrmZ0Bk69NmwXn4
1E8e8V1771hx5vTcE4IzyXxy+g6xXzC24x8gdcLZ/mYzEUYjUS1g34YYbAmrHIzOierXNx1esVQb
z+OQ9igQtlhVCw2iHO7jASnmxTfPL6pHAE2tOsmqstVMaJPs+Rz8e6W0H98rNPaHCBj/g12DM2rm
XeZX/oI2NysTZxGFxJv0QVb7xC4qcNRMuF8OtFJrQ7tp8sYDNSX0m07ZD3ChL/ItRsGUXjGDfsVy
xj3SmhMFutSOAf5FiiAwTjMe5rGKQN9KGFsHUuMqbuhLc//jp/tA0fRUWNKAc3h6G8Ts5ueuOZ4l
w0b5+mF/qJLZOw3q+k9Mj8vAHP53qMNEiZF7AQsF2nDL2V9I+mxqmLFFRT2E9e+VyUNRgSEiPdpw
ZJnNhlr4wZrp8YzPWceoXPMF5tLj/7VaNB79i093fbf5oUZCEZFyzqphT+B3jKn6hCwO+deZe1bc
CD25bb8gHcZmdIOoYIC4jpryosBFLxg/o9epq0lO7U4k5NRx/MjG3VXv7Bt44U9ElM4BLFqd0ZK2
OPDTX31ABg7+1/o2PQjuJzVKxMeDA/5Xm+VC3lT7Lt6Xmv88BIXmQGnluvHBJ8yPbKddLVGHUlpu
SemCNW48ZuZlSZObjTfGJXSX4oWAzVoyRHggNqydG2kc//GS3xweyb3NmY5ORjoTbbTLSAh1Kox9
nHaACejnNFfjByJl+RJLOu5SfiVh1H4OAmCs+eh6e0rNWEK9IAcdZM99/kIWRrZ/ZRI6W+lV+/T/
HVSBpX1YRUE6RLiC7JaJTFJDnqUb6tTu+4olzEcp/bmPUkeachOJn78vlWj04n2C9TKJWudUYMGX
kHNR+NrMuF1XyyoP981FC6YVCO5sUh9f6ai1Wtr2Znj61f3/chb8CixMaFgnRaMZnT3u34oL2cd1
fzqcUwkJMSpyGkYxpneoFyd59LiMrYNwUdLMVIJFAL7Pe205yqx0KRdO87JuXMlpF1FeW98LW96i
umAZucF2ANuH99rVmPGIQh2J9uIQa2zVNcMHHZTgNX1dokdLwW79pNWf3ZekzD9QA+1z8YC+3k5v
Do2G49NwCmZ83oOzcPSMjczl9Mx4BaftALDpgFXMLYFf5OHOE3La1uoMXa7Doitx6tJLB60x/tte
DD8Jq+SdsGgwBBAC7XwzImQANJQ911IkOFeOHe1yRQEYte6oaFeOYy/Ke2gSM9rDopkjzGGr3gOv
pcXsevIdhDyFzCpui8gKunUxzangmn6wTNJbtjHImtqeUYCvZTg6tVcntf5UaZsAeID6M5/mwPEt
etKaYSr0wOSSv6KrvqhzpSZJwIrZd7ZqH+QZwRMt0bQ2678F7hD5q9hqqMce/OvCcgjIwKA8nHQJ
62izAAAJPw/ElqNODf5eJG6eWPEBKeCQNEaHnz2lge5H/fXr6YNlkNfBJHsfsVUMAwOnQYhtet8g
a4xfF03OXTlb10FqTnVfCTM/JjUqNjU86fpeOZsyTaEiFi14XegyzzQNIN0FsFEYP4qZNCu1l42Z
4ipTbXaE4AC11Q9aXRg9hITMWW0aNiqzGPaIP84q+Mbyz0rwkpoD+pJdjI48gwTm/PRFr/jLemhm
aDjSZvEvYvF8YCTHf+TM43aNiGLV6Ei6eLEPNQDUK+Om+7xdF4AvK8USHCNkwD5Nb+hizIV9zUT5
uH6P1Dhyxb42rWRDXvAW+De5vd+L2cDfAUarDI8RHwbNb/RG6oq2xDej/8EyoHQc1/pAU2BpchB6
9ta6Bk8YWUm84i9Z9gIb2jWoEZJVVYS/PU/in2fcxu79QLdsRJSpRpBLjk3exUs5Tz+3RGH+Q9dT
JOzJb9dNpi0u11vV1DkrQCtfmyqO31asyBUcson4NI33iRWX3xoJkBM17plmfM90eo4sFZQgKL2+
qiVGqy9jKT7EBa5cLDdPeA6svegh/WkEHMSPsTC1QP+cdOoU/EHrqLP7ORcgXtr6PywTAoGD9u/z
dT67L4mXAkM3gUx6SamJzlmrZDclvmV5yDI7TOCHqKijEm7pD9YIQX6FuLGhmNJR0JNcTvpofoJb
2oYobZRVr6X+ynB5qT8d+mMGNix56daAcCuqTPTt3jiurN0NxPNRFGn97GUTD6oj7XQRIrbXd40H
xjH6ntZ5A6K6dBGaSXM6tCSSKcJpzuIxKYaSXxuxzZN3OX0jqFXjboqSekDCVxT/2LgBo4A+3McE
T11aIMQWC+svVIjSzrCQnsR905V2oBKiiD+QLnUInkjb0b61XJ+EZcV+TkuGEotODhMvX5Ch2Mid
MGa04U0DxbspAxPQxVQ6x8ZxHeTS9EBzngM+f1vntjMklLxbivrRcLLOhZg4NurV6vbG9AVDMqPg
2QG6wHEMqPg5PS8ZHqJ2sffj7fsF60Uc9elQF/Fube/Z+TQoVbQvmffGcttEzS05/Gbngp0Bi0Ne
xUurp1vU15oNmFPEzRL03yaZedNPyM/5MYmTjclVjuaGORZ1x3fAaBr2MKWZkuU9iw/Lrzqj+T2e
xT26WWBKc7w6T0zj8SBxNajzgmcHYSw7BTj5mgdE/D8SJZNIjAzMB2EH51xPdTKBq6JntzWv+7jX
V+kgfGfPHYT+n8B55lJ+L0EuxAsL+SideGuiacb2Qzsve2tlwBASOIDNscMP1MS6zPydkbe+eZb/
0667iD/UuNEB95rKh7JLLMUPJpn58480at8wgLIk3JJrxTBnlsocurCGwG65U/4XiB77z9s63lAf
Mq9Aq2WrLBbtXT3a7i46MklHsNvLslUUmKYFkyf+mPz+InWjaFfvSZWkP60TC1nazGTtVpVh1Tx1
6IkXXHtnVdfJGYMC+zl41ppWgbtWw/RXDNVW2ZTXjwuJZvKwxXteepzgT+4GeGimunqvDkQl6Nrh
v4N0aoWJJkMtcW2oMezOi+eIGBdCNKgsP01z//OWeUmtZ3Qz3pMkMxKdKGMd0cbEMEWbBxQAtwSH
7gABjrlNZlO3lTzxrD1K0S4gYLf2lYrdjWFH2q9QXtZ1Barwmvv/sVSzOTyag16P3CZdH6+zGo8Q
4+9Y1qNdV5dEE8OU1t3qbWAj62L3441uHvkWgLrqhy/P+vzLMgDJySvmENuMn/vyrXCXRbAFGls/
VsAl37PKi67eGfm8wsPBrbv+U3t0UPZThl0E80xXmRAQXhtQ0T2FmlVGFdvOTbP5Bv1KoUK6cRBh
hEcwjtUNOHFBvlPhpWKbU7sbyb1F8pY+3L+zDHA50663Z7Z6Fq5/IX3pYrgI76NMpWYM1+2EciRE
FlXz2TuEKiFqlVvn2IAq/xd3v2uvre0LiEjZ0pjSpYUSyRBGcMn/E3NpfodFaK1TuFESu+BVzZyT
C4QfPrUryzhEUoHFhxHR50vtjY1LZD/Lelml657cD5q6MT2IScRp0VLgTt9fwL713+OAiTjiw7BT
C2YiT7sxAyMB46namZt9Qgin1xvPoySpVwqXI31BmBJNIo7gEKk/Neo8QhcZytslK36I77uBJmwJ
1Zv1ywQPyJuTerbs3l5Z0IYwif6BYwdGSnsuU4qgCyB9O5qzlM+bucnoKQIY04By3F0RPX3y8Mn1
EGoLIA+ZS3xZWczkCajRTfXPd4uMhpia7VBFhMUh/NPAMdG2yUXVLd1oh9RRtcp7H06hJ77/2x6W
h56Kmh2u5YMg1YINhUvbYKNwTP64f6ZIEMvLvVAd9Uxd6QPH5jCGcgLCB+hk7tKhsVqteAXv8eo3
cU6soHO6OLn7hgz22a8JxmMWL91F/tOO904ehtEOElhi0Ss81ptWVsCAtlgtuuLyjGTc8jqgxyDj
7ZzRT8vPN2VdjvpgsnwRVPPz3kxhrsmEgSjLclPUtKgHGf7EZIhAgpPHFat+fBKz9pT868UOD1VK
5Q5k2ldsavetpQkrV5RCOk2g7Cw7couIhSA7jXcP6g1ZImyTsmEypLI3/zYfywpJIAWYmhsllFj0
a8vEnr/0acR8H/UrQRi/nxa7f8RRlutnxtXzk1uj0WQYybyOR9QE6aE255jVGNfYSWrBTPoJVPV2
Ee90ry+p2Kfrgk02ewIqDhdFJRkgsAw88iDvK2/KS+WZYWhLJKh7AdFsJJNyaXv/589pKULWqlxf
HM0Ds55Du3IyG0m9Ii7cMkxqoxW6Nzq7f2cqKUI3NmGZcPWPOM0h04Day/+VND8xS6w17XI47xAO
N8tP2sigAE5J7FFMUJWhDxaBIN5dXxkqjpYYxerByIJx0VfoEbhFHLniFOA+321tUGkfjJoj2Xdj
LSK9GyRh3lFaawai2/c8R/zWwx39UzwHR27bZnZIxMqXKHpeodce+LZzHQSgipEgyyk7A7t/G8PY
Nmh558twOVGiQHkBbW77/VtQAJsWbidijAtFEgrK3Qwt0UdS9QtLclN4nAJNtRUMRDxBzqSL7tCp
52kgA9Gb/nyzy+sRTo6JfBZsiRNguGBgVo2gT2UJXs5uHI0m8V5ZsI5yfO+bSdzcgxsJHJjxSfKu
3d6ex82n2k9okIkhS13DEQlbDgBR+rMfkBucfODe3uyFNOUgqeiwzHtff+uxTthw/f/k3igeC/R7
fzzQ0nLdWNlwlHR4wsrAZ7GkJWr+t9Q74AaLXospdXthXnDzg3ynIKFsewmW9vO2yzRUTpY0dmEx
DusoE20l9wNy4EasQDcXKlvcDBYyEGI2bKw/QDCX2U5XvUp+bhEcqYwgO03gVbK6f1fcJavQttrt
FsYk4Xk/7J0MtxOF3gj8BuuMcmupaEMkJDw4e+R3mlbt5tvkZaPSAYqQA5R/+X7X8cQPp5lPQ/CM
NVW9KpUr8LJlLIuNvCEd3LSje4ozkxWorrf8ZtngexokD57FS3T/chbW62m35I/7beNN/Mq1bQ1r
AaNj+2bxlpevWaGt7as/gPpA620bJe9WiYxB9AYXdoGnVL6Vepdm6CZx5OpNKGLulkPT+cDUb3lf
HvPU8tGxocWMIdSYojf5NgGpOgiiaWI4qCBEQkJjmM/1iwyOLk5vYowD7n2T2TSMWJ3s1XtCk7+E
HIQsg0iec7WZru41YwzvGhqM6YyHRSQt9uDPFuwTDduNDI5hFbtD1D7Z5Lfyn8VVWmfZIQb+uMps
8Euh+j1rfigasg3xskAwKSUAq5RMVHlHJCSHsLbPuPY7hjGQDNZYfE2kxls1c5HBx1SwHEJGNaeA
mKnagyj+E4CdGhiSiYImN5gKtPchXE+G0mTOAs1JLC0wEb9x4mXSYwyA7H03O+UnI7xEnGbuhDTk
iTUeJfJkaMIHCRhT5YW2uvPi2luDGd7I3lrIQHsoWtUiZ5h+7a1n/XXXThXTYcxuEBZDCwRSFavq
9DulJGiz1piLjOQSLvCbn6OMMvF/Q92uAGXdzpn0JVHtnq5GwoO5jIfubGk62th13vsFF/1Oo2Lp
dxVP95csFWNZjcnNefFM42mgAzFMgk/XkJW+rBogyEUOTxcK+IyvzFCJyiYXc3rNAGrmYOuLGm8i
lcXvzUhtVwTgmw/1zzIQ0bTWRRga5eIUqVuSCI7YNLLJpZygnHieEVY8jkUlL+SRxZPJQmzs0Q38
AfDwr0Fm5R1zNMNQ4+h1Sq+GT/7YSsJiD2H8h2aulkVmbeUm+O2kv9N12Lw3cmrOOMPI8fsEtzoC
1TPbM/qU6pWXF0Ky5BAl4txkUvUtO70mGXTc2BeP2lsgpGBnxwYt+z5V+kEkKkuqRkzIsbMycIwk
IPnXQEPRF8ILzm8CiK4u95lHj4uqFGic+XXmcq+RmXZzHwmIdbBvjfQ6N+HiSYqEFhuO7OF+jjpo
MWE0gK55miEfQRVpiRDhNBRzteOF8wbZtqTQqq/aDVY1x/qMnO0g7/dnTsUDmN0YDLHCyoFEmOcJ
5YfSYi+LxI144NdvdsDl/gOrWWp4a3bbT//23X6dhozO3yGaBIrPxxAvZTGEn/HvLA7AG1e1MlF5
4zaLLzqkWIFuuY0cGKAQT2Ce7pSwAfrYpPxaggR+lwN2G02kvLtkzv8Opfw3JORCmBVEVDja3za8
hFGC0Na1zjrGqQZZBqraZY27w4LMwt4g90xiIeStIMU+WB4zHJApKFy0cBIcV76Z8Dqwd5tpZEFp
bSMUTA7FQ1K6u6H/ncC0DfjW75RWI8Bt4UHksUlM5A+BdikeagEtqbFvWRv/LRd5BuCK2l1vThvS
VCgHs9B2qmfZHJvjdlRGv6g+rVvnxMd1I+gpB24XBSHPGgGZYozpnOl1kmwwQ4eP4PFOX3Y/ga2e
ORl21mrPvKFAtwrEJ4QS6HwT8WYykeSf+oZuuxSGyu8zDjYMFlH+xdYfSrE6cDZ4fiVzLdRrgV04
O5IjmdHT7M8Fj1SLbhK17tmclZ+j7DvuuDpwTlQfPi0ftLl5vHqipvTnf9+54eg50Jz1M7JrP7Sq
aLzUyUHlF+wEi8NFyywdcxo81qDJ2anqvm9Y/w0KVVknts5UHJK44yfayOpjCUCjjBX6BpDcn+Q7
MIoeBBj2Q/rIeOPNEYItr8BRsnEzGki/HQlwVVm7U1t/sPG3FKHIfiJkEoMZ5Sl9AnPt6kCnQBvy
NtmivnjXv8aYcSN3uyox5ektxyHQnED6erG/vR77gy+tc29mGlhE836lPLiOTs20kCeVmxGa4Dwv
Zz7XB4Ee876wxDHV4XdVJ6f01l69eh6h0OZBSr3vQa+DfQZTpOmzP77TjcqzCJYArjgk46OpaEIo
2BysaIrgflt5laUJSKa11hSai5SxF54brLqlZlB8VCau/4LzO5r+biTm4X+z69et65eRyy9Qqpcc
1HgvHy9koJtLS1DFRtHEBJRJo+wPUgvZkUWTtJ+ET0BJjk2Bn2KwI9noGk9FjtY2SrOF9A129SQR
60iYh57lQmbjpSM2LIhH+N6iHPVoZSXFLc0XA9Y4M7H0eZy6ffObo4jPKHnOMrTUeBKADdGKhIXe
TN1JyIarTNt5wl6VEEv3zMJuj6Svhi/tL/EhoCxxSHaIAnt3qyiKW8SRljj5pcW2tw7yIjMD3RW0
E1drzH9GYGTwy52KgCnzYAXbi1s8Pg4vCCn5wSY8e4Am12srag3/9yChmscVbaV8R/KXWeQwAooX
ylnYQ5lsnl93WTqXR0MnBot3Q8U+aib7Xt/Xv1x4Ar7WLJuHMkoZ7b3FVnC+4d83TWqvvWDLpDQb
/1I9r6Ii1fjvi7Qu4MZrOxrUoN9KETe4Yr7yOyTpr6MnqFScUP34FteYb4aU2KqoDwfjdkZc1pa6
UlhQLlhw/Hf7EP2T8u1r5gVGJZnlgRXDojeSqRuLh9oqQhdyEFdXJQv6Vehhw0sUi+xTqCpoZOqx
9wBR0ZbyNW8gpip33sDXDRpWqYNmiyw83v/irhtqAdSDxZtxMilkWc+qOxGp3DdY2MhCKVgVYITv
YfaGTzHAKeUgqdkbYyoFfEuEmrDhV1G/g0rMFJLp4wiQnxGREE1tq3hNQmSsc1Qk75WQqYivfl0S
cPLg8UkzTTascaymZleIc+KSq81oWvcIysZ1O6yB7EllcKvbPp0HOLIyF0FjTEAnroEg7W7g//ZG
nb6vzlblGinoWrjvjBkY3TkQEok03i8AoWTx/TIQhnLdK6pHf+ckCHy1erH5i23Z6A88ecgWbolY
8e1Zd6v87vCAS9XOtd9Tcu0mQ+N1OfhZo1op4Y8BXMFJO5X32Jtwa+o8vQC1Iyt2//6cZzqN1wyW
SradikiYfSmbRbU+HnWbsfydNcW/UlhW19Ez/3Aqf03zoqYEuFWOpp6eaoGWcsxxdst6uNuAulPE
XOk/8EZEmroYcb0sFUqYu5v8IiaW8ZTB9Llb7zGtIV0Jvslht3Nne7AaYgJxxY1jtPWlTNIGSIBy
mZxGMG++N8+kPyE5AMZOwdvB9b3gqbRTsKKc5FUWhbKW16gp+s+rM1V5H54f4i3aX3XlkyGLGJCR
xtKSBRDgd/Q7glNYBaohaDEIZubi06kr0RmaUmGvVPM/cAdWb32gvubxSZnCkB2KJaolr7O6q5HZ
VwaEoM25aOEoh+xMBUqtbvv4C/wly/UPRN1NdHX9howAuO+Z8OQceikTocDumRj/gEg7226xP12Q
QregpXcG19DFrm/bmQl5BKwtoCPmuQfoMA68W5Cfy2tim0TMkKxw0DRCNNiSdqRzVdgXegXo8X+8
Swgb5yCw24XwXNZ69SE23lcjv5qHX6gh9Ef49/td3bWMGqvMzHNLEdeP1pJbzslAv4v8JLddH0VU
6RUpy8V1jvaoeh8Whz2TSfFbkPsy+inGdLfrGQOxL7UlhelUbzTQfa32dnznH1CKElUxDF2IdCwV
zlGVGLlv2VnFfMkv9KJRuc9mdhtl6sW5NmSEj1nKRT7xxdal5WrSMpPc34cv0+WP9J/yvwjvLH6L
JnvzIc8AKBi8ZirY8oZqDYGFpH3EPsJyT3pYi6x7ATHN0zhcZ8DOgwou+aIiHKBM1ZccJqCRqByL
84fB2I3UMYI9ZJ2tGnNz4Asj4qCMWwZfZ24xO/uJre/ieLl87BCpIPjzo2vYag6qQLNn4yn6WHxj
x0s9JI7gCE8Bv0idptTG9gurBt4oGcmHkQ+BeDM6C5yc/TU5LODnw56pVb2pxh19c2oXQ/Jxluxx
Tsi+U+ETtcLKUdQiHEYN9dDiEEK7jXr33K+XzXuju8+HuH/0Ra5uEzM9EfIDpdXiKxe9v3s+p/Xd
TG1Fg+PVdLFhyJyd+MUrqk3N4MZyjeQBIiVrKW767lEtJJUx7lwCTueE/SuB9sxp60PnPd/tNC28
ZLszAzHInfV+ng7ibl1DTfSolXS4Q3sqHeLCtXmV/97H42zLbbBJO5GCMmEgskBBK1n7kgKqt1J0
LdGbCCirjJFFSvsqutBA2RkwKkfneluykfeNRCYP1o01gDF4HRS396vd76ZDbitzV2vmoLYfKzE5
02tyQrRHCLgg9n1RSQDjtJYWNXN4Zfdw4az11fBRNiSPU+RutuKDAz8Ucff6ASqqe9eHsUD+R7WL
ruMKBTcysG0xZqxUIWBsxLmU12dCrWMJWeevEYuJq42YYfR91bG2Mn4gIRT1VS08bhREHu/z2KBO
5Z7ywCO0qyG8YDMVxYIfeM1mYEHotOCE/D3h7Mybv9tT8xMB8L6LKDH/hrSwmKC/JH5R6mynlkxL
Q2EKJL+X9ov4wJPH2p4AcnrVK/oRgbf+6ZnbQ1TFjBkLmYmNwSB68/WxxHIa1GAziYSjNLimtAZh
JM1ptYVRfMnzf+xnUdx1mrcC/MZtTOP+wfXR9iTOxWNoqDkGfoaF75Q5aiyIHHKqUJ7zMmzXg2xV
SF47/cLPVgB+2pm02Alwr4c/udv9TGfyddGhScRJokohZbpguVKzDvHNXMMLxjBtqOCtWdBJdApE
WLOQgw9u7z2EGmHbRvnFW4M+OYxNHjA3kyQp6qhM9yYpt5ne60s2q/Gkjik7lgCkDozNuEQFKP3e
gk6Mnh18TL9ZZxNc3Lb4ryt0PpT6WvjK2FpaDMuG8/2ZmtvJf7SbYsssYi5em/vqUN9b9M9HWffY
l0vok81P9V5EVMfYoz5hKBmciwq0Y33rMKhdc0MHWq3O9U7xYICX4I9k87W6OtAx66fNZCAjRh21
1vMlkaiAyfxA2XbPSgYXg7HjCeOO90TNTg8D61bqEecKZT/lVFdn5a4ZzOjwFvm9aPEvZUcn736G
t/BIhuqgcLthGWfDG9NfrJxkZfAaVSnS6dvic8DZHjTjGDaOJww+x0He+qX2nv+TBMG9oGSDgpLG
HpEkpRPtd6f2huFTs7NslNnduwTYgK+Bjhk6G5dT6qraYVsTOjmkE4njQWlYgjQ44OA+XWOzXVaW
6U7h/nwrlkNRIGLuuj/vooyI+ZxHf2kgT5dnSd3W3aylpPXAX++sLcIQq8U87+QBe6lmtLlM6tt+
f42YRVSnQAisRaMXv1J/rgFnf/4L38D+eF+9X+itC1PVpN2fzcAaATJBXkXvhuxELiwt7njvW7jI
jN9dNNVXF8MLXc2ED4uOw+5flaQXh68ffvNQcHxN1yQtbCKP1lI3z9vTrQ7+K7mbt3Dg8krF92Un
99T55XsTTkFmrkMs8vE1Fczqi4DlpiNWG/scQ18xf1N5pYGntNw9m2fLInLp10X0bJL9Ye8l4EzE
OSwFQ/qQk8HmV2Apgbg14fvoEJK4KEk7/70b53+vS3WYj0z/8P3764nGVTVop1+MdOFYJuVf0npo
kPpdo0FkNO049fzBEhbCEa55DFFciqIc09O+KC+KymbgLCJcEWfeJjwCmuvKTD4tADrBFzpchEKi
aSJeNAFbKAORXrcXqrdjZvGRjhmo4OpF3vPw94O3REGSkg9SC1wV2IIsAf4szd0rgHSi9tpNVVf1
3kfLNJmnSEuax+GXmlPXJCE0kJcG5zS85X8nujakhXKdWPdcnklCU/A/DXDLXuW1CQumhrGHdqQq
M8QI8Dlm5wkAKbMYrzmExYxiWxteX7RrWqxuNWPOTto5cqCwfYuSN3HRNLIul66cU9bMRSJUTLmT
4O2nRbp8UbnwAnL8AF4pSoEZ3A9p2Sb5B249NzeUCRv/eTQOXkeDn79m1QNM2LfUVP/x4waoQnH9
IocoHh3JYmNcsPV+mVkKnkRTaTLE2fUpdxnJqnWVCXGtrsu5xY/sWNx3xoK4mzFYy8dVAYicdAjl
GphY9GmnuTZ+9cOLeuFQHGLML/jJGdQ+b7unGykbjXiwOp0tLf2rgLsGKL2eXTJAc2kLDSrVfgVc
ksZEHISZfTWO42fXOPxLfL+QnDWfDBXLG+cYQH/rdiGi1Q9s/JMhu7gAVpIO7RrxA5rAEHB8Jwue
8FZzN4KOMJVBo8LuaSYxPJn2CyQWTYu93/UM4tFPjl6hcDwAqyY4z88p9/BZuIEa1MMiy0SehD/t
JzR13ZsP82ddm0UYCaaaZYWU4SFghb1ijNL1iFAxvU26asXUlyyQWNvC+juD5KPYlL1mlRXDEhSN
G2upjZq5ZPwE1qcXyvJESu8CdFb+Xv+7KU5RCvss8c3IHpOrNyJwMhvcch3PXDH5AsuQX5XUsRNA
45KqFnfT96kFfN4479MJcIHAvOAu4uuNNF/Bth4KDQvMABzBjs0BX133uvVRvnmiLOhRBJ24EBMH
4veT1h6RG/j1DjAu5D7TCb9hPsXhjpnYal8QvEMAL+NhEDpAesUXC5Hi+7CGHJE1/Ckx0Z0Q+h/N
TfsCJPodVlBU2SAMTLCihm+QzZnySRHhp/dzAirWt2A7mAR7mrNjt/QEIHv/yNM1NAEOEAI6j0f5
fDzz5NjlviixmDyoLILQjmK/t0Ho6AEhN08/HNkfwOUQgVf7HTA/C5vZmeCfvG2qSjbcoN/T9n3X
GYAw3/HSt/SRRnkdh3q9pUjfWRRnCS4VCWoXKnq1ZVtQ35Syk2WJES2hF0nRuO2Er/bRod+9ZX1H
4MWvZX2kB2vAMU9UKDoA98KNoPz5ShbsHQjvh9Njdyec+21cF/z0daUFX6ImVyVtmluFSQQisnqY
ZnlNoXueD+q+IW5x9IiMqzbxe5OZWNC4AHSYK7ub64nAwKf+zm/8RryIwjkSYUwkO3S2dz09Xsai
n1GXQ12RAqiVXKxS4XCvcaOZ2kPSy2oZIAmVviC7d+gz4xKKQwHBU1RHOdjEUZqpbfjFJ9rGv9s2
7kmkaZcqAZNHbsaCBAVY4Mtl4tsB22G0d8+ZPzQnare/gFRY0deiaw0LcIm8M2UZbRsxSfxrxj0r
nrB7lUD3nSkmhJ2z3TxqrZqJIN+AnWNXHKKvQEQREm7uSORLeyXYV738MLy3IZj5uy7BTqOh/yGu
izHPabcrNa+Egg7R4bq+22Qh57z5lQFqDVmbSKv4FqPCy9jZYsO6qts4R9bIQHAPDWQFzxLa40Ux
1CEyzff1ZHAqCEUGTFUaJaY3CdR3VVCVnqaNQqGH4NsThltb2TR64ZFujfdkb6+wggPlOvYIsXKQ
46D3ZdL6qVQsyfIxJfu9S3YThwJ8aw+CDU8N+HyJKsWD5EB/L5jHQP43cDRyTMjfmbGaRHPhkexF
C7vavq2ljQuEihdw7wVspteO9sHVVA5zHXJTwO4r9nhm/A2hTlo5Oy/sDrY4pHCH15osAFNgSwnE
PtL6HOfYxh8NZ25knZXQ6vT1m1UFHgffsPBeZ5q4wK9/2Fpej/2aRhGHwdnLUOtKsGUinKty2Zlv
MfokUl4IJfx29yyAwXl42LPBlgtxeeZeGUc3GWjkCk75mCGrX1Jc//GEFamY47vqwm4cZOojYTnR
8iW1sQ3eQLt03xevkLYB5aGmCPTU8VMsJrEuEC3rca5sVjakzL2sdfdQcwkEjNtc8XIyGpfdSG/J
KD6e4ED39uBAUO+ovu5qAThbg6bCHaKAPIkJ9xMMd7P+Q40W5tsb3QAYuAS1xx8lbiNYWPdCTnEk
/13U6xk92ApJoyxDEjT2tIH716upIpgtEBcwtf25308VjbppfKdYiftPHaeuGj+dX6cQ+4ldt7dL
ZSFstBJrRGkVqAzsVCy5izRVkhKj7yx/wIHS8YWIG8MKIFH6nFTP5GbtxxVSRHlvD1tipSBdYzWf
SM7yGkr7QjEbCdX88giFyyAzhd+tCblefwJXDjdzjk1/DcVSKZBF/AAfaFFyCZ4GPL1WCHofaMDv
LASkEUtQEvDtWI0/C6lfkxHPzrvGia/rLHBPiatjljqmy2J6mpdEVmWKHmBipL5txej7KiMyK6Q0
tVILIhl2CEqUeHe5+4J7tcRQ8xDA3ZzGnI2xWZ1X5DHcQ1AWCKjd9B5vuRA17gopku91oXuldDPg
AZ1Rmbq3gqLHntrfYZqU7avoF68LBZ54NFglqr0Iu/kkLekNe9jcX/naymEx1E/WGNIFiCSsscUc
QjVPFdc49p3MWH+DjaWgOAou3GQCD2k/ifPW39s7pFUnZB7AisS7Q5dv0D21/vNif0o2kJfifW6c
AJnqJ0MAFCQDzN4L/oyHB1pwLIzw4Fc8yEbWtmLz0XJokbpYkstVNqfmrEL/n5u9MtogcFDI4nDS
TRTqxxaek8k2XvNV0Laaisxq5fm4Lba6LEWO8v7Sz62zPEldBDdf0EkN3Q02yGmi43LzXc9HNbwn
0g82gyT0mU0BzXeWrFRGr0IrPXrO5/toVYiKKI+sQmp9LrYPOuZkLd7Gmo+63EXapaPE5evYgUEh
ZDfwPjYqcR3qVmGU1cykHj0sj6kdhcGF7gcY+v8s+J5o7fkgEvfbNDOonpb0by6QXga5f1Gx0Tym
l/DCkJ0QwCF5K3taqzC2QkLbF+fsW4WhLhk4aKUfPluuS1XuwjBdIAC1k/5YFOF//7N59tPDDlWn
k0Nr/EGr8VXdqQ29iV/EwTh5ikjVTLQf9rAs/t3sUTo8DMLadeybp7Jkzq1qhEOTm3zwupc4LZtS
wzIFSrxmB5wYd7GLohU7dPucQqWuXTvadrYOzwKTNjBfQNADuEcGlCsCcp7Oyu3bPPhdjLUMvPls
GOFHe/NctlKficK206LmselPRKBkqKe++ZLBYGmK/gzNy+0KKHZSW6ZGf+JovEwCx83Sk8utaHEU
lOOCDjMnUQ4KazpZE1/r969cduqRhfIgAoRCT03TvePGPAM2DP2g5r6yQcRQb+JSdDBAZyez2bEZ
GMwKm/SdJqBH0UTK3XC9qP+aGH5calb6aHOjhrSwiyXbyerfMnJvtGaJfUQqBaRmwOU7AaDAlPsn
mPbOSAFXAaD8LQd11h5SgHasrP4X57JNs2goLjDXRWEIYUe33CVzMe7CErsS+dWAbO6Ec+EF9KFF
lrNlTSDgi2tXHRHpQjqLVwANbFm4rpKES4N3vkzfG5VMJfN91W0ETSTZK4jTR6DmBPB4dTJzZDDQ
kez6LI1z3kBADOKJOPFA54+dtGyzzK5/HWJgc81+rtV7ZBTaJw6ItPTZXdzXD688hIS8bi88byAN
RBImJDHnvs6SkQlXjZQmmVi9+9Yf8CDsBxJ472WahADAzx95Au2ykXIm9Cqv9AHJsBrcNf6QpOBW
g1JesHrtyLayLj081xssvlyHAP7qvDucvJa7QWFQQOCpEJ3Moa93uAlZ++WHtj+Wly70xvmoVHne
Afu45dR0pBv6JbNnZEHVjdbZ0Q2fNfKojmrkcKPjzN0Xf0f+JiBAx+BUHogGA4YCXHGS16PZuBRV
4k+CnWg6ODPcLRQWKRomOQAb2JZs568xd21QgXjReEhOts+9wmzAZtSg4ynR5fKueplTPofSo38A
l3/23kxTlt51y4UgCUBNODTvXhUFCgEOYrJFJSyeykztpQXD3WvTc0xTf9MHwFtmRQMwnQ+98qsi
TAg1YXdykzxymAnXMMmo5Y3pHgtEkQj+/aCj7xU0iwP+pf+lZBw8H6ilW0EqZfPG4Owinm5Uh96K
OlyK0Gmr6TkXw9N/zphfcArvQ2RuSXHMeLWomyim1viQvVr1PxLFbgMTza/d5+UdZCQnEIfTD9x1
sNrbFvtmQxbFSG+F181/CdEhcym2dqx/5A8OPZS6ctJeEBF1B8LBOO0dRj6pvbZ9dAfbM1b8BBiT
kHIF3vSKpDgtYPZdrW/OAehc7hEAemIfSMb5feO2dPyCGztJM3hWmiwXQr20VAVLc/XOSc3YJgOc
IPWjmos2fSC/N9FLlr6fy5nf0VEAXCGMZXDEloZzpte7U+SmimZxJAkM4pwsZWzioY0FSxt4iqYQ
UxBs6ENHNwER9pNnWrOccNMdyVI1+LPoKApt6qPpHqmV4FM1KFou7cx9ESUJpwxDUDQ5MOU7fVpF
etq9Ok1LwbVo1jJ9LIShoGmsmPSF35pMvxGAIp6Dxj+Jr0hrqI84hDCzqR1/IK4//5z5mE7+gHaS
Dm/Lyrz4ATdWfm6PB/lfJb9lbOYWyBxvYdLIC5vp+QNWg7c9odf5nlUQ0FuoXOGHa+LRTDOAawkn
GhMKn4WyUjvnW6RYKgIul1Uuldid+g9NYzSZKfI9RPotvpTSn9Cdi3iKDicQ19hNPQxj1YLlqokj
6jJlX1boqMjSSaJlIiGAywA8CBpNDY+1eFL07sq6T9fk7Y8Tcf/e2i3LTJe9KooOE5PXyncOWAMp
uE4NJcXEJ3yGSsm0uiaGnJv+m/zOv6gKiI5ZGuWDWqWQR7exnZ30iUl5r8ik9jxbIcn0lC8LnXKE
QOVFPQh+KXOPUc/+gNL8M7h//6s2E310oyAGfeqHU1EosS/4PRwbkbtPlN8BH4UKr9nQ+dvLPeYO
HFAmxvMkPw9Gg7zX9jYoRhcoSl4Hb9kuKh79jfXc0bI4Bt3RrJWBRglOB3VPMi9P9JjcvhgoluaM
HAXzWfiyurrZnmLO1IgA3vMKFiXMfkROrV+vjDjZ2/10q7pGpvm5D88j+VHpDMcptsiOznfetzlE
SFcGaBgVduXsZkAlqIifC0aDJoeBlVgMRtGqowh8Q7jooipOXtTz+Ml0Lf7zwVnfszPmXsVBP4Ry
gWqPiYrcq0cpiGfNb2dLp3CRK2SL2fKLqnT6vEyU49+0DbK2YY7pkVI10BlujFm1iuwQdpw6wOUS
wE0cQXvnlWuw68vAGYkpvAtlqz8waidIU+8NCwt6x8aO3kS/ewVceYyNG9lW2WZcaI/50BR8sV5u
R5RmDJcDcN9Ss7wQP8KeUuOU2jYunOlZNqrseg4GusXX+9kQzHaCNOevxzvyuqEVAYcvMhMQuk/1
BEk48h0K4pGcjNBoAZPR6gY8dhjr4LY/wHs52Mkn3G3yC7H/YYobJmFPTI1+3WlcDslO8jtxuTdZ
LB16WmiufdFJEVVs7+9ERu0+h+4eF6K3LSqh1g/oFzQZ6NZa4O+5Yt8Lw6RCNkSN1+TXGIIpJ6h5
mKrNFVPtT0nubMU1Du4M3VF7r3OqFXs3/9HFmnJeXUGa+pqUIIvVWwKaQymR/TmRtkVqSLrvrU29
+dH+nEoe4veMMKPAAs7XGd4LrRvjHPE82a85R5SbVyfy0Y3Ba2Lj0Z81VlCRAAy2ONe5hQiAXd4g
SCnjvA249gitoLHOTxVvDu1blF5yR1bQnsvLil/TUw7a1BPs43FlyahDFdpenC4ZxYSVfKxOO0Q7
eAhHZfp27RiRdlBVRdwF/r9Ge/nyVVGZlQZpOk2z4mJbsF1R9C/yYoQ8IWUSzfHlDZOkTzUkVtLD
3zRZlJsfYcGx66m+3dFe7JMfdqRVo4ZHnxhWXrGC9D59WutVS/kkPwtV3k0Y1j2NumHPCfWzvaf6
4d6w5rhQuXYg5581kBeBEs68Br447weBWJlw0O/Pvprmzo/2rymt+VmVrCY7S9DKM6D3n2c45Sfd
UpOEukZEd6b9OO0cHVYdFNT2mfkq7JUYh4PmJKp0519h3qPags5sWRm06/sKEneHNxrWBGECosLE
Z9V/oaHgTULTonK7RFTC78nqNv7tJ+tUpgHJramDHXrqQdKDAd95dzAnsFXDdi++vkz7pyKrj/E3
hST/ciIuZv3ee9xn0MQMZB0k91Z0X3/0qwuhwd/86fPHNC6ehMsxXlQ23ZqkShw29EOX5T7z84pq
FjpdWUro8xOjviooF6EWbclgrv9/PZZL/WdKCqrKxayiOybEDAvHbV23kQc8O8VYxHfnNx+G+nVh
sx7LhkLy8XEPF3aYjfjOYGC50dC4y38xxMUMMaK+ADt70+VDQLeclfU9zMXye7jWQkMLeQGZLVy3
u6h18LVz68oBitbyXGQIWdMnTnoS/o6QT579DXyyoVMBaqj8vOm8X83KxAibNI6d3K/oUexFpH1e
EKh4m8otxRDzNTiwnJUMnFJ/sMc6h2G3S7mG0wprhRlfKvTabKSy2Zz/ZcC5U3kBQ4+VDKPS/EwU
xguMOi/SpZTeSV6c8QI91/ouRBhd9wzDTFzW49nSW2Wj5ZpiDz9NgmnjX4Hwf5jHYllsf1vQwCPC
8ETPRNO7FTQL3gu4FUXdutW1nJrv+fGCwfnQt09QfnjwtFQ+VFbspvRWoGCwTBUa3CdVkx8JuEgA
ka+KwmyQC8knbn4QGSCLNRbV9n9VyEoYuTMsMhtebFrBagTdPEfklakoMs3oWiKUjTkVieQw7ild
CZmV7agUF4kKcZ48S5IXaidPHfIB2Y+/oLmASYY2ZNP9xfb2zpPaJWgdyYfS3zo0IlWwCDXO54hW
4u7go0/4we+IBm9bBCVce3VuX33HHOdBsRVZrhMsNjces1ZcT2Nuhf96oOnFzGaxwZyoulWimncC
H4Gys1ywQjiHChaY1L1dLX+/FjEZTAcPUQ6VE3J6c/JGSAzYJ7AyT4PP7DYa/weIAHQHo5gCj9a2
CG/hxqYI/LkFX0/QSau/vvZ+dxenxxYAlg8+ubUtM1KQcr0twYIDXkbI+Jzi+tsRdRK8Ci377FOz
UWcF04LhQ0+H9V2xhjxJls29Mjr/f3VPWu5IQircEeuvPPmy3mTBC2rpj8sZm6w7sF944ze7147n
8gKe9v/oVu6TZkCwwfuebwmwZjhgPY2IAXzjz/lewo1Bev/4a7jWKgktmOWoRbZYXxdhKFPziXJp
dY30U6gatIt/yUOkbFE+DuguHaut8DX/7+p7XcqoYPDIaBPAH1pNtwpwG13fOHbisLLimtmQvIh7
B18dv3hWNT4Hbkp8FG/tSEoPZgvxLqKCFw7AfPZ7T9xreCQJ4zvrDAi0ahKS8lC15mPvXdqm1uOi
H7bCwYRHdqy84eM5XLhgYKnQlWrFl2VQE0s0T5sDEGmASTJgqjGl7/anPS0k3IC/5K+Egf1roKEb
mHKRcPfbK02KuW6LxHieu+uglcVQYS3QPi7o2rMzMPRNIw5te0A5XKioGhQ8vWYPNi9OKn1RBXyK
adFGWZu9ZnKh3dMWTrMtTd9wCs8RI6k3DNXcsE0ZZNimXHghWkBFCtTno/lXKmegJSO7A4/6L3Td
LO6XH6bCHN0+TasQ0G7I9aDOGGtwQ6tvbtIndN9he3Tt8pXbX4rjvDQ1ebqn6+3p2649Derz+NNL
ND90RExv9Q9LwM7A7Nsxlb5Kpb7OBS/kizREVsGGz+0uwgYBi7LPblfv5++DOdKbTg8UElSVlmTw
JBupt6U2MsaQBeRY3nL+irtwo4tcR3h++osFwabJ7+tVRW5XndSDzs5bga3u5KkxSrDdnpumDpUZ
3RXHix3PtP4TkyCGXITE4m8MPJsmrsMiip6XCN7oKf04kO44PGrNgYxU/w0Ljb9az43OTd+8xAOQ
sJ+N3Tsr7bzUTPKRIgwU+F2fjj3t3x5pFbTYDvZBcQQZ++oyaOwwQ7V0XNDZeJrkwbiRCA5jRK2E
FDqEU/0PNz0MJYb68zP21qAntd+hNqkeX+c9qVx3hhNTQnAMxvbD2njoaUIIGx9flSfBf4I1NuR2
QZU9P7Al8J2OXhPdBOkdMDFN1JUXGZg+w30ylwzrDCOdRl3qAqgQRtiDVQF7a1fr9kXI9XdCkOQM
HWebUb7KXLloIkP/LnY7MvyRokEGfxlKq6skcUf5hck22V8waEUpODW83pnxsZ9V2wBpeZDMwPfl
Ur8w3gqAo4Fz5ncAgkgWFa8FFJaGjFgcKKx8H5FVFTAQUQGhaDHhp864ymoliSex9rSqDsX35ilq
368/SwCXbcXYlZn1sqJIkOLHOWjxkHIg4A9qmY+A+Si0L1nwSVu9V3fm5orTlphnpXaPNAUcdEsU
uKwNdbvmC50Wxh9E3oPYRgxxtnttAgjYWayMUMITmFT9otAqTG4talzDN++XaDRNFwsepqE44wYH
gmENbEH/pCaIWiZ4zbObGeUefTw+XXJxVSmhUpN/qVjUi2Oe68re3LlME1LHZDAe/iqdEF/Pa4v/
RgDWSDmyUOtvo9h6fwtRAStgjPWyoz58v0nvBBjgG7vQRB/SQC8BvwqIAmlyMhNNU+b2fm0a8K98
SPBS9E34asYLCK9vXeFqeJB0/8nlTC3F86CU00MtcL2C/Cf/YIvaqycbkWlkf3zeorSi0b86RtgS
3uYpIc2J6imU0o7aLnJZVUl38PE32/rr2+YKXbt/TIGm0Y3py/D5xreKt6W79McrJkJmxquCiuaD
9mhJa+5b0gXh7rfXD9zomW84yx9qKft+WXeiiljzrYWzDXPiDDoOJuc4o9ZCxSiVjnu6hieuQlk0
qmh+k9cPRijyNX8IodUOur8hlRae9dIIDAJK5T021yIXp2RGw8mqcyQJmyII/C45wcpB2yQTHJ9D
4bGUU7NqfSL7w+4UFgb/QPRwi4KTRdr+/LA8f3xgNSYn/9slMJfX6ZriNvqVxmTq2/5jEuzSPTA7
Z9NvaJTBem4GeoHkngWA/uYv9bktPdkcyV9Tg1K+XeTTgGRCP2yWJzNuZDTSnLWsCjf6AIYGsPAz
iYP6erZob1xg9i0KhUrVOHL4vExC7KHqfH62gO2Yd6da4eWDsUUE4oPqena00LbHGZvo4Nfrm/Qx
6i9Xae+903JFyqTfdAJSaM5wSVGwpGE2zFEVb45GIR1e80rfPSYB52rHlPa2s9fOxuHSfkxgiLrU
6/U5AfdrVooK6qqwC/xhfk5MWlUR5HGRCDYnF4HKCJ/TzqNvjmtPiXTanU72jo4zhM+uVIUWMIGB
FH05Fhw5LQF5MC9MyTgy2Bpn3AO0A5DZnPmM2jW7XQf1xy0a1KWoqUcZTZf1kbGdeI6poyqqqzc8
hFBnroovIU+A+Eo0jJhWKo/DNgyFtYOHc+4casFrfuWirKE+O5j5C0HDOlSnPyPkxcT+uAHLq5NK
V+LH7G751s0mthgPHKZdOjintv8YmGo2e+2c4WMIjyc5jq7NbKH6vQhuo1gBhIebKYYbrR07Lv4f
A1fzmvKWpYXwaYrAa+yJBBZ1VUnC3PamNJIQAVBBRqAQc+ZQDPI35SYKj7ebV1CymvXRsyPpD/PS
rA/pZP5p46rUAtLWPnFH7/3kVq8NiG+7JBwkASbqd35U4cRpPBNFMMu8OSZHJA6c81tBUhtJkgdu
O3sUnxwG6JbGsUlLsalPSwde0f0Gro9VDr98yT+k2I0T9cD1eAXSHrXzb4xlL13a7PEwIpViaaiD
GIqQSfbI9w1NffL0+60my538kBVJPL0nba7udjIXHVSE7e3++gi+gf+RVkV1Fs1aIj5bIWXHmmLV
HCmsxwiG3jsqJswLj/nFn8szA0pYVwAGzNMqW1TJA20/Dos48RS98ghVF2XWsQnAPSE25ObN2igI
DREPu3lAGD12CJU7YfgQMaM+FSu+0PEoxBkAaMkHvLg6BQWDAqLRDjvT9wcOTR5QRXDble4BfMWe
bdBIO9Eev3kdPYhcODjAomemt05VlTg6XVdEWMwkOHV+UAi8/nBOXIbB/eZNVLtMEcTxTAbAkNqI
VjLRs9uD2iJm58omNhjb+Tl3JT3OUoEUbrghOvtJ5lXU1lBL6kmSAxvFhUkhJCRyo/sH0jPdjj2z
0qw4fOXHDxVVwsCO4pcJXlzwcVHJHaW3IgXf0w+CcZkNaISluDe5iYtj9UaH8zKGq9MffrAYy4Sf
19K9nC/3Xl9xZu/z0ScZQvS0etzQRe8pUVG97YSXQ/mDox201iMezYb8bvXCvdRkV2UAY+DqFN+f
UYaweLFns4fPQqJXGTH/JwpgGSrl3rCuehpWmFnl/ldloyxw/k7dF2MUOEmXaCPzWCtZMkh4df/F
GMqHisMQh20qZcaq//Gcjk4M+IzjkDDo6cmiDl9GrULjgmjUrKTeE6JHp81ySLH3o228yq2wmL37
15NIPUtwcjIwLpoFfU1EMKAqV8RpOZQC8kj89QxyrmOXWwLPHeoojzKjG0tDGFJgnacUEhFX4ZKn
JUPtnxiw+e6VB3FGFRV+ftdTf9UvajcTibTUrsDrB2PbMkTLOtMNGVqEmvssFIpZjx8bN+EuEkf2
DCuRUU2nO6mT7bzqMMlUGI0vL3fMETtZzoj7Xbh87krH7DciOXot0ggOuGLkzc3TzUMHAfj7fis8
PyqJejsyox6qmUlAvc2In4B1Z/qZSu/5MYLIdhKoAutKPS6Vib5H36T03NN7Wy/qummrmGUrYc3n
PJmz2wRHkj0tuY7TJE3dXGzcVhybR7oewsI2t61wsf76bORzk+W6Xcz8TGuD4Bq/Ea4fkteq95CK
twXKq37nbYC6bBxi7EIISRIZmxYO42BXZKGxt0TASfEmRLkLJlHRNjUsmk/WBvsk4Tavw67m2jHt
lmzBcoKThJDLg7kpmVonCxn/ThBwJhTs/EeavvbzZMtYsgKepmu/ayBL41j8RSOZEianm4f3EWXl
oUSq/aHKLAkS3JhC4exqcrKnmaPVsU/h8p1G54yvM78DTPXnnUwkhKk2QolgcD5+OqkvktQ5Rg3Z
aUk80feoBNdJyjJB74prkin7baSTXxo15rMW0Cfrmv8kI1ljhI6vQ3ypfIPToKRxg2X9AnBdtkk+
EBWKE1tVHVcvebGN/dF0HSIJqThudli8OMlK6LIbHByowuS7YCC0Sw4J7uXCwnG/YKh1iVv07s2b
gOqCSa1c7fHoqZ22eqhXp1VvIEpm1dx8wNjBasEnuUdxC1issE6Z3E7kNfRnWSXd4Xz0qF6UVH9C
YmIbaKyR4+q8W+UkRE78afdLQXXNSxOXZJe1Ed5IDpIga1M0rOF5YhtIjVGZafaR0tCjpaK2WJRe
WxdDV9fjTo4DjxXrnGrXgNqsrTOnQHu+DRoyFiiIsBihXuaj6ly6EnLOgJ0ah0XXKvkvkcnsRXbI
I7GYCkA6dVAyExff5pTzN33NxaMS8TZNOhLqThUYq83C08qcCKKvG+KT9zdrmU4k+AeeGsfuHe02
sN4kRTvQz9XJkdS3ef2T40EnSXEnL8KsATBnsYE7YZXI596r73m5Gp710YvbNIY+iQCNsREY6Sl/
K7/hUAGSeb4FbOyhxmVxUJYHFpjTymcM2qc6DrEiPABX7eNDhek8EaScc1lK5Z3mS/8a+qdZ1Z3X
0fY0WZH8VX7mTWqHSKO23p5lmgr+muL4KSa8gWJ9lzCISqDWjULC8OqPMJJDyyv975VWWeUNZuH3
zCyBV6euWmDvf8nYqzvK0mCNk8vf2wg7qmN9V6QkCBOdTImL9e2+eS4PgS4ALRQOXqgcKxk+e8Lt
UPyPhHEANGOIEI8vCsqAydAE1GIuXCeq8TnQAnvkPKd43hWpb1DqyJgMo1K+/dlzAAyOdxvMtTQ0
t7FX/YsgujZ4gvPfWjIAfGzH2Z25jZKmbZxUUKSOsW+t9lxlPD2Z2MKF+SUoWVOZzmKpMdlw4CU/
yBRngKdJpMJYtP0BepSBvBPdZuYbJxEgm0EEs3e3FSenCiZj2/nw4FXqBIGrHNU1jMeQNOwps5Y9
ewqUdD9r5LqIiMnsBNyTCxdPDditiz3JcCLSLnaDaU6p/pQ/eJIc4KQw0fE033Q5Nl2uva+OUuoK
GgDVdwXjmmJYJeEa/L/szf8I2sVGOQvHw0aSFQxt6u4XXtovrm6/EKdbMO98L8WNoz2LWcngFmJh
+3aoy+VwPJqW5llni9zXTcYGO/+x8GCVr1CVsLbw0CIysA6ZkyLyEOK4Kq2EQwbSLXnUtRnnASjv
m9yKc35jmwbGEI5IaZJvhkvXJ1qa2bBfrettZxueYhKvGmFO3Ea5o3zHuEktquwy7y3SIhu/pRiR
LM6ZCAJUDbyhZSeQE4177A5V/lSXWwjTh//185hVBrKKd4Fv5XVULBoubFIdobtXQbI2NgF++TEm
vqJ2FyZkaToQeQznTjSzwaisAfvPP+uZMwPLyqQRM2+95IEeApeL4jPq+nv1HoAaC61gUaWfQeci
hPDPzNa690oU7tqAtYB+y7vnCO4kL73lxObUSA15zMXK2ksruQtd2m6nTT+vot+qoBDZF/hIwnqY
pSL6pf0RJGf5uOMxKf8suFTcMLjkaM9/hFbQ51RMnITs3ieYJ1zGbvas0fVwO+vYn022TK8A0C1r
mDWNWJTvMeEMij8+qXGkZ6uGKrQ5ZnIBGX3eUCEkK1LGRqmMQ2cC2ZJln0zctz59U/miEJGn7acr
vJc4f1ASkGrvE0bw5NRNxYMn1HZjtQDT8wGCX2zl/vG/Kc9Q578HlIMvgSysknY3+8pkr6FZCJUB
IbvkBKEdLK/EsD5iNHze+OPHAix1Sm+KkXkKXOcWo83T+NnXAYXLwq7OjdyUBGxJm4Hba/3Sh6Se
4EiN3Ak1BMOeoy1/vmQWMYRJ0yLKSgYespTC6oiR5qRHQ2n3w1UUl2BRsy9P1d8ifTNb1Pk6Pc8u
fAqea8bbDi3ApeG+FpVMoIBW4cUOdYo01fLDBEQdHXGGDQi6prUaFCRb6MSICj4QBGzX1opJOzXj
lIrfQLr4qtwjF8ip79psRvhI8Oy64Ez1/mChMtRB1doKNvU4cxc8rNqvs44//t+ITlw7qNa6IM6K
SozjTYDRloZ8C5UkFOd6nGSxD/oXyxfA2w2gT5pKB5VCp7+KKRffEHAiK3L2Qy51MrYmAI+Js6cL
GUdFUTCkf+ef26jeIrxHen4qxCDr2Xc8L5YYz8kGFO4OOZHECvkHR54muSydCJ98PBcFDQqViisR
78rMK9JasiEVVqWdezrrM4ybKi7HMkI+Hgvcl/tsC5ZQB87AkGX4iQdNPNoP74qFmY5RHI5AHU0G
b8JtxWv3Q8b7aqug+KsshoHaYsaU+5CnIMBkraSEukFqsBmxIo95HMfH0msKf9nbKl+1KCE1Vlww
Mt0O48utkvtLe46eYQiTmr10DrxHS+mmVaStXxSQyIHohBV9XMJrYjIyKHxNFGKt4mMoqb2LSM7y
uOnYE2nNNfWvm3Qxy0PBWwo/3pfGpnL552ICgRFufFqc/bRB5dciS5TkTbZ3txVncK1mWz7wkv4+
PzwzoWL9k+JPsjVMmPvsUrOHlHRTjPZ4dkCfhE13id/Mb7AmjS9uNNAN/G/x66Wr2HW9vVRbylmQ
oGBcSNOcYpF7lu7hVlL0AoaQdjhnqyW6cRayjOTOx6tlG17hnUmMtnn/L0Vz8YLOKwNcMd5GaEAa
6lbmVGwEAsLarfEHiJytgU099ys57ZCD91YqRYvJIBFRyJnfSwd4RnGWQmlrdFBQKsBlqkMHMCfn
pVyOcWNRqNh2/wypTHwr91HwMDZcikGoJkT9J8tgKv+3wLoj+4GP/dz/oiIXCbH0BexQ0YSSluu/
hjzOLgYuJqf1QAl4Pc4LtrbSJUtRCnNIB7rnJjlddWYnUVKHnJcjTpjn1a96f0HEMle+lc+fCvD5
mVQdrZa2zeoedVn8hjTchi1kLrIBG0zNN7RUqIXwaNBOCKMhS7umAXzzIyCqPosBEP0G34pUtkq0
3uXK707o4o8lkfKwlMaOnuLmcADZLggS853KQGVkn8+YUibrqmH4BKS+AFs94y8m2x5AXruK4rEF
vL/7rXdAzy3KRzB+11n5IJUIafAJPicHGSmB4uBHjY1jwlgiZTL6waLMT9ss0SoTQDlX0OhBFpoC
vEqN6JCNV/xVkEhXmrxbE23VlZ7HlP1pexTSa3e4NOj51xkwN6iRHPPhCaJKRG3FB8ZyYrS/xRc9
0lUUXv/6whiGU9VxEgiyjSlNsulhbLi8jJKo/IS4p/rtNLOHwb/eapbHEQ2cmylOpnRgXiHk+q+M
cmqUeHuhD3xTegoCx5TOPlCkrqhMgaPUdBQDLvngim/Rn6Eljo2+yozb2yazNOM9pYNyIcz62r45
khMZ+w2i1k/cvX7IVG0+ZfN5J0f+TGqXXwSFFKjckw3jWsLP4ZJbYKFMcMKdK6xQ0Eob9Pw4vQt3
soD/wlvTeHv4Bl1PtX0DQNHK16+DkVX1olnz/BR/0GD7HZcvXReK15ykK+JDra4xf37iJCEKR+Co
FQHWIFyTbjQZRQAIqjAis1sx8H41GDBPaauFtR6nKz/ydPMYVoWjetnVsbJ5wKA6exHiE+fOV41j
D2SDJ7NVLQwGjIsdx9ZPoLdegySUqfjMfYBAYDqSYuVbOPnGptbTLBtOpbe74wKDbAhCOSyiiPzx
aEN3MucP7SSNVT/FDBWIsEJOZVx3rC8s0t9shmJspwrfyFX5uSOnxBfYNKKaDszwBafzSQfbD1kL
OEfFZOhudUVHEmKKi9YZpq4jCT68NLPc/haLJydGF2wVjlrTkzBva264GHqhzxo+9wWnt7LzHDzw
V77RPt82OZModow6/VAbr4I0gz9zG/04HSsFOJ7nUbuPjRP3Pa3TOkNl3yv7nM+B14L4QGVkRaDq
6eyTtgd+8gzIMscZDsJrNDRx9u65oNPnDXkghnkvj/wZcPh++eXNssHOETszrjlbNBg5/xTCdaZY
IKQA2pnkU3BgaFjOOuainXHk7qaQYzkU3qJdgPA4WzFAAVosc2cnmfdBrDpY5HIuWW9FhPAJfE8v
OR1JKHXj3HM46PEYo1oLmeDCQrMA9q3I7GR8dY8NN9QoBMbmVM9Vi39yCvrDlMtvK+75GImPzG2U
JVzAWyOXmj1cGW6hkl8RKJuoxEAE4Ytg8Py7pSiF2WUo6zu3EZFxxuRUF2gHymNhXJGMj/RCG6YH
9KaofSgsMK10lUrKXTewFjXnuVfnp4fX074euGcM7dVwFP8KR1x2VO119WDU7h0+eUQgeIzY6YSY
XJoY8vykYJJbzq5eVl1Ex28BdNVQM0lqFv4C9VRMag0vHTukj9gC+XQqGWW72sbzm9+Ed3lR23DG
T06I/vssBUFFvw8gahfvmuAxusPUTm4kKK/iSASTVI5wJOXXe5cLpv9fDQ3aVs3eRz45hbWfWJJ4
R8cTV81s0dIUKCJYCye3kZNLLwTJYjnPhZLtVvQR+NUNhKwQZDVfQa4dQveiGKXRYQ4MIDdv2xcv
1KCp26hh1aQhKIfSvr7ll6/1F1KWnp0TgL124yR+mrE14eNYO4mLLauaCTg1O1+BxaLXKgN1uTdG
xQOWeJ3u14AnEfUDIaVC5sZRKp/Gcb4yARMPzzchKaSRoN+Pso0HPbmd7G6tqfSNf8fbPbFrmyXg
8h2q7fFKzF8HCEoHoGr+iIStOfOLuzqdP624R4CPhU1PoNq0w4uruIhpf8yg4ecX1ECVn2CfDeib
aTzDBLS98GyAhHdV5dl4rjVqsVvzSgCWOMgYWR1gHIf7MHogTLgP7ZsM/Iux4dcDzdVoP9EkLSt1
OHKdmRkoSMdddvI9U0oz19/4V11opTeOx5Vanpndd8RKZThI0oO5P1Xk6KeiE1vU1UhkT98pFDwR
r3Ii+m69EKgEFlMBuIgNgUF2NVugGMu+RDA1xQ2KJXahdy+C1ODBLf50YvI95eCBCcMoYd1bNzdd
mV1rDcqJqdQOk9IR3yVv7KtucRSk5Devb2vD3oWZKQuU0l7izmZriX6oxbPblI9+a44nmqZdcvqn
6oWlsPqcdvulKAl0OKpqZ8kPCQejBhO7GYKlSIJ5xIpMTHw5F72pyQx952TGyPJWLroAB+PWLi1n
0wdnSowQjNUPZoPwRRdF5Ar7g1HpWHJ55qdLYId53/TLCKPvCgdQSPXnJiIkE6nruGPg7QxFD7p/
Sp0yPQS9/bL0YhZDyNKvFX6b6n36GDwNkTZA+Bfw6eFyZFCw1IR4MQI+rCz9qLVUE6U7pgc4OqFj
JYIPtc9zhNPZsdthz6lrfc9pzYOtDhxX/WIcT2VDdBv43oiI/+InQnmoNVJrcEVy/V8nBHjlQM84
KNmgtky712P9MtDR2U9bDZ9r06M0u9QVU0NHg4ZpHqFNoEiULttfcng+21PwaRmty50RF9wcjWzQ
wTzk+++KOmHVA8zbn555QzZl87/gYkLg9lDUhlpy8ie/RkGo4P8TQlq2H0iaQTy/ObmYpsASBYEU
jEXfvBjqVLClFi3Nlhvx4fdUks88bVw0yseqpaU944Qx/BUnljJztVD2p1Zk2al4TLITORIiGjoQ
CxTffTVhTC7HUlXf/+iZJi+xMTt/ZADTDn4akZU/A9yE4qJ/GQXsaLhUAIK3I5fQvGD2XL+uCDlU
I3AE2Vqb9R7pR021TChNGcJ77TyLJoEBZatru4QNP0Fz1ICrFSBDjvyDi0aBKPRSR1FrugSSfC2r
m2KepqwF0MTmSX/sImq4VbvzpGGi5aiYStBiAK2AgCWCPNAG+Ut8nmyvnIA/fKrX97Wb7jz7JS1Y
tU/HqFkEA5Va7kG2HL82hibut0nuSTZsfLg17P8QXHEEgM0BQGcNMTwfJnXcHPOe43ettZUo/3zT
j4xkkAL6DThpiXQoMsPfK4sUuibgNCLqveoonjafYp6fX3ceCJJYKte2PboAqArMS/f2Qw7KKe3E
SSMRAE+SIg1nxbihZhi7pTXm+KTeiEYlgNkIJVWyF3iY+JYqKCu5aPHn4m0F+1N/FVfavAa9ZMQm
WLEmBdRJ1K5vMSb/JQb2GtLAPVLJGTna7JTxrfTdZ3h4L4ExrywdhYp8NwU8ObTQvzQbjKgpS5Sg
ZPWKAmTUfS+N6xKarrVfrFX3RFu7KT9+REtedMheu0pc5I7UAtxJp+6lhceXPy2ileg/BDm+i0un
PEvn6KfOlQCHjDy+njUcrO6MteL/oNXSQ2ACJ0madu7pLOZZ/IEV+6Q1fBRsuNvDe8k1QPMPtIx4
qAcN6wsSyhsfKCAVS5E/hQhGsEQYPo2e+9INHKrCQZ39oADSiBMZXOV73pQ4zdehfGdkAYKmEgjW
amCBjEkEQLE3pSMctGyfIsDPmQVmMozXTKQe+/iZkRWCHwE3twt4mlTKXIYbMXf1egR7yNA8P+Mh
0ZS5dtsDdbqVLzQsm8TH9b7lP9i2R2dozvnJtHp5BW2wOZOZ8sgJQcX/V+VaCy4GWBm04b7n0KsO
UIWhau3dfwznoFLOM/zdDjrAc5OvYjj5v1KzIYZevAJHDlwtftIF4v2PducoXq5ehEiWx/CRu/C5
McDuWaqQC1sMc2jHttCAeffDeNqWi2SGxMMtur3SpG3+n9LlLZzn7wWUynDRg6shzmJsrp74jTxQ
xzca3nl109bEXncuKn+g42ObQf9wp0nvdxwDLwm31h3DHL/eDjArcO5Uw3fMXLds7aT+nxXtfbw9
QCTusx1kE8xQUoWuQWL9cdZrVVwEdvgJ2UjHHYgbMCs9/GTkonirqSfl126h9Eml6nv1XSQtSfB7
jCF+wWKTHzrfhgsZxMKwLbpmGtOOqzMuiUAzP+ES/7DIKUZeic2fE0TxgCEzbGsg2iuu+YHdnY3S
VTWsayLepJ80wfEL7SxjtbvgSRR7JHLQw/E+nFv05Nm5ARY7nlVJ1ycHOpt1VyN+7p+uPKHBLAYo
9cis3bItDBK66CwwW2kxN/EBW+wLuaxIkfOR9QXMsF+G95s3bhXX0T8LWdzx6Kp4liislIVw11zU
uzUkXjWnmv3BDKO2Js64JclUnQmMADklJaDDvEMfS8lafv/IpedIGKLyidCMl974PpGxjVmhNPFk
MjHAoTU+nCVpfXNM11FtE2CR7RjVAbN4X3s99O6MGOqf3Y2OPVAWThFEfdFyfQaQM463LRLJk5wC
oc9pr8iYQx/9BEX1W5ep7naAWnbBioMNp5h2Csixf7mEiMuQk0qnKeayvrUPB8Z+8/sk4iFq2dow
uYXpey+XxHI50OKkf2XywTwsab3wvWc2DzAWiPnIQwr7V9hO9E8usCraRIe5CORfjQEoHHJlRClZ
syiq97XIE/WxVAiJUQqY3jb5LpgjPJVPFwfn2WK6550xmmDUd/hYrNlwOkEKYD5U/FeI7YC4h/1v
UQES62BWKFU3Fx7bKyL1FawBPCrT0Ui6vUtphHTiOQU4LrgLb60kiiFgohfmW06u9gmb/dllALNF
LWE5Oq7WN2QQ4zO9z2scWOxqgy0r0Z8g24kghxI75S4NAGutkcjiSchdIAGuRtHpHQ9213MyBBI1
o+8m6E8d15yvF9DTxJZfkE/BBrN8Nezoy8x1ngFXWmAJCH4Pp7eHtuxnTVtNblMojhz/2RqFDlSC
RT/YLupqB9y3ks1d48X5h/vqicQYvAGgjWTAZIUSd1Qoc2sg/4CHmcL57QKVBP+6S/C3FjOjh0cx
9bmkiI+BsuyYFUSQ1bwqQoIH0y7G5oFoDhfmSx0iQ0BK3n2dThjFE9ZjG1enIMMQ3yQudvI7SyO3
zp6qCztu7aN/dxh6hp0QL5IsYOeu2sXnfXzQtjSsdW2k2/HBzLhX0j5n6cLvsrauf9Bv78/naL+4
n4Ai/jL7IGFgqyf4i4p8NwCXD0yOsshkYsvvEomTQhhGv9BwyX6VHQ7Afy1TWRs3WufTKH7zBbAX
t2pw5BCMwvPKJSN3L3bXN6jaOY4xHBRJ4cA5HB+e3y9RBhZmbXpz02FhrQAp+mof1XK6keH7MXee
Ngafg+ZDnDiqzS/aL5ODErQ1JO+s7oN6SumXsKff4fnAn6p+j9rcBCsr4IfURDnU3+6mY5u6VW2p
pEyqQPEFN0BOm7aBT7P/y+bMLCoT9ZAJfqXOE3V16YHz/Mwkb90munx/jqWJ1kFyXFZKcL0dTMaF
nTCD/aM6Y1YsmvcJIvchCXq3uHJeZI+lwxMrJvYRIFhg+k633/gf8yR1SDGfpczxxwYSvbxUSJ2E
Ui3T2yuHO92fsb34psoeBs/+sWSCs94qrWloemdrill3UfNPRrNF4tzyy/yuqFD4rS2SNu9/7YNZ
/348E+nrWhIxcwffw2mXkqG2WLOhTvncsMxQAjcJqkZVzBrfL/4bJmvDOlsaC3RC1q4VTJ7e0TNz
5oMwpjLZOv/C5MB8banHevfJPEn6rDEhj/mSJPaHFlKEY+Ybp9wJ2+bXgnpjnz8C9GeiSd0glrQF
uGTE/A2n2qKjHxU9vL9TzbOSvWgmYKfq+Ui13K5arh6fMlPic76Sd9WjHdauTg40z24e5jGZeJ7Q
Tq29HDhpgyDeIbL1UUXHvWyCIpfJCjBZElOYuLd2l5JKR2d5jWnhYET8QdHJRHS3ecA54vLFqpPJ
pvRa72Ymcq2ZGMj5ps4lCtJQGqKqX6oEt/Jk4R8Lmixv9S7MLzJlsSTstNkLdaJIMjo11H/pznd5
qTyq62yl37QbAvH4DebxZ7HJ/ArH3I8m4UADC1WyrDuDgcr+7QdJQ6a61oo2apFZTmTVRsbc0mAw
UC7HD+k8PnfVV0187/bxP9i+MwMiQxiVkV0/RJBp3X7FJJBbVYyOdP/9mWKastW87YyMHn+QdxPE
PFdSY16EvOm+cPq4cACt2eMyLLOAaJk0y2kqLdndQ99Tzbq3zlYbLhAP7DgNGvTvxJCin1AdR20e
ZamqTd12zpWAH1FmjGODMcfIb5+GpWxYb89p4YNrVWPJwfZIATOBM7Tv5sEmvc3jukarxb0QiqzP
FjbXNM5OA5InDNFulVv71SxBaeQwRrIYJ+F3zrAFAXqS4XSags+pbTAowgm7qTzIzLEmp+PJow1z
3iE4JF+nTekJAsw0weo6vys8dkZC4mHbg1Nc1kfBk+H2c+B9TGC7w5HNi6BQ5RqEtBKSxQFAtZ9Y
t+agnPJslstTDF5cMHCacgaLtS8JEPnnaVvQQXiHX9K7KiN5ok/wI/cI/uYzx8K4sLaGVugAVbha
mYm2PkJ0E6Sg/HCKQedYveBaDSH8Amk6ohzDaGid7m+Z2UxlpJeMVaNgpkPmRH4AjM1BEs+mfIm+
w88Ju8S0skvXscVdQuCSVaS334WyS0Es5ZEBXb6nDw3w9xQQAU5AcSOxN8ukykD+Idk/7UsWvlLq
VAzsGHimVpeks+y+nN6m+EizzA1G73oFo0znRSB0UT8AkNm9kJXYga3EkYT20fBq/sPQ7iKmQoPw
5K/9CzSFFXLVY6SlKGqVxEd03OuinV3NESeQkrfOpmjVsqoiFU0TELF5StecvG3tAffX6bWnqQ5c
O/WqH0hjZGsNr0j9A0a19U3+oMTk5M4qFHFroDjPKHHXlfOzKrBuxg9qQCIeooq5wHcn3xsqn/XH
FTmTpL/qMgtgaZVFxqnRwUxf7J0EftxizufeXKGAzS41lZF++FN0hV6dJemc40jLiGQH6m0JyIte
DSQ9hgnSg2oP1c4Q+Szpr1FUINfIw5WogZnzzFQtpqVVcN6uSRAej140lYbr4Sx8HTzMe+s/a8d2
eB1SSSk04DQ99CwCRoyDyYelg+hqprm0YDzLd7vLlEDqCoptkADHs43GnlYtyhZOzzPGojtSEKXt
JQSncV7KS4ZxxmqI8QUaiQTu0suxQUg0awI5N55u2p5y/22cKXI41gMPvnK9dToxwVUTCaE3nv1Q
E0etiWFzGTn3q8kYC+vEZrYgVEvbKHIHONFfsKVwLjBwv5BamtczV0KPm/tklxFTrIpZvMdQpt+2
WvwxuDp0YshuZ+pjYFu2dMAO3iNxBBlDVyJaqw/YXgfSjXHn5p+re1SaB7QCGDyuhLCpJI5arkYf
Lqo1g/w1fnO//YGt3uxDAIOBYdqr5sXkoYnBcYGRH52IpkjBiBFF4aH/jOQxeFBL2R0XeldAz2he
sGMgOeFMvPnkPaMoq5lLsNvsXAkbxPStJL5R1xaIuIxe0vT+VwABSLiffdjyly3WnYCG09fsJOUj
RGqV9XGQbDMfAdZmVw0c33A0YbZbXRuz821FU4gqFHCeV+TE7WZYmHgUY9PwCwuzZtIhw4QSw3pt
IZ/VOiarxFJXbVbxyC/kT9tiWjMUIfQV3o82baqUdD8NQOudAYueunNFvUOK3W8gEsNRfyK+LyLw
Qte+uUpW870Ea0UHAPEpnyDuozTWdPDnk97XinskboKSpnqnk3t/CPXvgUz/4etcKiXeFkJjwYc0
OPTXwKis3i7gnyIARo2ON4izTmLBjkhvlLmHvZEo+8i4nR0aZd8LYesvdBXk4CeN8nfFbs39HSJI
MbhuhI3bCIjgD9AjCGXgsd5djC3VOM0MytVG/t13HF4LxmXG4O6qPDLIImZBlvSpBrZWy7FFRTjt
NmBgFRA1yh5EUOdUIGV3mx69TCdw6R9ID1HlHTSuZIbinMK6rGCbd+aNA4NHrIVV02po8ZnPeDOS
jg2ByCW9KHS07uhdMuxULJUYLzEsBxNP8h7x0q/3SbIyipj4Nd8w+s/O49i80HiALQGzGZjnXbZI
o3h+ASfugOTnUDmC3nKVgq6R8Z/ZdjTZZas2oOZtte1R4Alqzo77SEa9c7HVJJYhgTXbZ5M1GTQ4
YMIVpVA20+n9bzBzY3w+KeQKJeXWrLDQaPyK4HXPK1mVC8T94kQ/2MTw8mBCbDSX/42L+lAmmcHB
7VuSucGrg+r7pSlgg9XcvR1AM9Qq6sw1XKkZ4fbKLANG52UF6VW0ZPkqiYKK77ltNZKZnBb2LIyw
aNoumy3SiCZwYvu3tlQX3HRpwnZyQbSKVoYKgRvYZFN/DYBwBRSxfDUL6luu0B9KbxHVfRB0OzQB
g4jmGGMfv7Rr0dLi3dxAH8Zx8Ixqa9myvQn10OHb1VVn243cCkYWdf7kaNC97IzBdw4V/umHDmKZ
YsohY4hvIt3MHzFW7M5XHj4/Zg0GhVRx1KkgJLY24Yhi9B/BGJbzSkUeaPH0yAbSuEy09OMxsx9r
1a05zTljCQquYiDeJwonVKF1ZXgdJgJofpacwhMSlopjjLFz9hmP9w7zu3fN9bSrNiBfzslM2VyK
MfeU+4LgojyF0PBZjTtbrjZjXCK5sSPrExua7v9Oyjw4R0ZIYKgkXwJ7Z4G2xHTN+cAAhNO6OAwJ
+4OJEIh3syAZG1Mw/d9984A+rrAbXWDlIWnFw5iPL9U4XWZ7F7eIiwr7H98h+XhFCJheY5GbInG/
BvIDhu/SViqkwGgv2qV45hujU9UEuFiJvh2ICDMlzfkCjW7JVQgO8SUZnBhpbRVjwNDAaI+AKfBA
6cM0zhtUTedpPDjiV7SQfQjB6ziemPd5TzewVN67F0eIbgSAQcsI1E667+iC6h/Nf1tKYS2XUBM7
/ydhe9Be/iHhg/NrtpAENr3e5go59UojJ+JkbjOe8281MvLGWvWAaVfilh53IGKN5CpRGMo4d/dV
6yNHY36UdUaDhQB6AM/siafLZyamM6KclrR/b8AsejmnUQrCkcSWz3gkwGNA1Vt39bjwL2Sn3rmS
AMoLnDeFRaZGu88jcA65L/+qQGLkpf56bphDtgsgBYhkWPAxpNwni8L+PkefN1XgMChQtTfXeeCb
CqqoRZu72eKjudK9arbDXN3DwWlRrMDj7HsNSkFnDSxp1Kd1db8jxtzk/d2E0UZuVVFvh1OPLQVU
VlS4erSQtRgrU6B4ykPIEde848L5El4DWDlZkUIEjVG59dRPHoHCCguC0qoxGtMtu75gyZ4gWh6F
SDRUyLXmXkqbMruS/YSXiFv9MUufMGjRTXP/iHYXKDrRszbxPzZWKUgZzMIfOMec1CGXVvVKNhXy
z4Yl+Ze3cKh5Aex6zoCRivtOTjH6rfk3x+oda61OF7+18OBEiyrh6UVJwKRBVU1yQPDLQ+VBHQIN
JqYlldzY/fReq3Hlk36Eao7PHZUjx6vh/NCxlKZbFdsFK9jzg0MoctKxI4ezuEmU4ei6zxpJK5Yy
icJbJaf2aCSgrGzfG88WkVlcr0iRvE6RMldgREbeQZjVxjrgRldpIIlnrAl4NUgG9xjeUEPDU4jD
ZbfTH9o2HLbNncg80Id8ytdYq1D6KXa4VMxblCra3/T0IsqJOVO7wKX4MJW7JU0Ehh+M9be6Fc0J
hv1QwjWuE0+2tm4rfFLDol1ivSDVZuBke2PmHmBkLc+oEp99I2HpQCrbytpJ0GOOKA4jwT6Q9y60
OiGxTbax12ijRuFEF+cBGtOtS7z9/DmSXjFBvNPx39P5Y0qq60zNsZgCa+fIukrETW+sg9MCvkp/
h3/t0zo4zbNxTkyueLUZ86WUAuH+7lVWr2vtAST5CW1J0ZQdAol4Vlw6r464bromduMRKDs0ktW0
KUyRDWrdRav2pMKhbczXWUDh8/k+B8cGdluEMcJ4UNHQzt1vs1ZphtgGc+EgJJge074d9QlcGnRn
UluJrh93JeKNxu/49sguubRixbYfpiSSX3TvlfcFmWC60+YDXfJNwlRDranqoFuOzpwFv7x0/MpQ
3sd+bcmmYeznKINquiaTJojYeQ4zAvq+CfHBg7y2cD6WZi5oV0AmTppIpdEPS7s7EAhDT+ifosM0
KxedPheVZqh4acEr8Yg5loC5M1P1EO/TJOmchOQcZSubPaBsz1EJzsjufvuupYWrtLLkrCka2CXF
1Zpg01bICRnNKE6LnvMHXAOUNZusmelEfFjtr97tljtGu+LgFQsNDAM8NHVU/UNJrr/KwhZvYmY+
ekADiPA8pTjdnzMhJeuvJILzJ2ruxtxgFjTUsA0KWcK0v6/4tv9DcgN4En8tHFgevdRC/V06txId
6R8oEHkhVdVAVNVtw7hsG96OvMtyyyWIOVPAt0sDL0QQnSjU5nwmCppVN+1ZJvpKc7/RBdCqD/WK
c5+Y0+KpbpPA3uvfmTMYm3XUguUIjlrb1bsERkVV8piZbOWEv08c7iM0gZlG7vb/0t0Y81fw9IIo
eG8ddVVgq/AMmnX9OGbGPG8wKQzjk0AR5ZFXW2SmH0ECJLYFSGjT09J7CSXSENEDZIz1m0H2eoIo
QBwZUtNRG/mJQ0YfwfmN1TrXkSp54KX21da1QVh7WtYnGGVOKAalXYye7jVbupBIjqLDeThnCqu7
vFc7/GUv9xZH4+wPWQfxha/iIFP8GVCmhGhNAYQv7OrRDs4j8cEJ0r6ormZqHBm7XbllqY/PrzFc
E4pKgOaOU3ApgQ7dMdExXOjBaUfsogqm3PPb0sGuoMkglivs8lxbXa0QStaidin5Ll4LPY50yWdl
Yc4QUWODMuri8o6ss/dNZxlwihpQIM3MVOQEUZOcCNUD5ejVl4Vf/uTJVMtngf2QlUlk0qP1HZKP
nwtUQTr6MzJ2zTmxPW8Xb5P5/e35P2iS6byXJqdjKSmljLiI8A/Xz3LF0mi2ThaZg36Pte/Or+H5
QYEryZ1+6/gPgNcsOo+ji0vwsHt40pYUk2EAaBf0UF1YUqXEEtpqsmoKqTmPmHEGDJEZSKrjaM0q
3L++lKDjPOuIxiLaD6Q4kYzc3CUM/YH4/1UM7dxlK100Vk5SR4zIS6xOt3Cw4TUBQ+N5cEz80LP5
U+1CDiEAhTRbpuzZ+6Klftb8BXT0kKGTBMO0S3W0lYFFnXMp5JP56DKwhDqd4lnQhflZ2lnz96Zb
c8XXxnzHj2fKptKMGQi6lVGB/zO7e0qNfgqmrkTNh/WefnYf2yD59gDKpwnWihRYnYlq/1Qv1htL
psGijBeBY2QF0Hb0Ar68C/fRrF3IxdXVAMJplPsoXCV3wdHiN35fU4lNZPT0zs87nEBt5dNBZta8
DxVmLEmW703ptdAohAsvbRMvOfVZrVO3XXdUha0EL49U/tVAa4NQ/wMBqlpp+IMidw/VKkYX0RtR
6HR4gdqQZT/qruyREZ4Z6EolMhq1mfjLzURbK6AQQoQ/TlJnPxWGAjuJZed6ubhTkSqqhrgXkKj4
sLteG+RHoSULHjz5dITrHkxwcsh6t1QPLVKMwzwIbBA+CfD9501z4d2+eOAmG0t10hp7UGaZOJ1T
nPsxuo8fVWiIzffxC2IeofdwTtgdTipUeUbTJs+2ClUOoYQQsarkP3YV+C4AeDbcmRCxXBhtCz7I
vrfz54B1NebVc7rcVLmopLIEUx/iOcaxKkfvahUlpXz6eKSZ3bW7wApZ5jgbrbptxl9rPvO0FEsr
LaHRVyVcIY2F4jSNac8PfbRnw8pN41MrW1WZUmO7+lN0p4khlSn/mADsa5IDpHIT7IBR8MmfPQiX
OtVzgSy2GjBXBcgUkaFJNgEyJW/+jhOgoq+F1BH5EoQPfiryPX0oLGVsYKHQF5nMlG3rBhvBFnzf
XsGSNFmo57YL7IZjzxgQ/Kb6O9Lr1MuH4YyGz2wf8eW0INQdMk0aOl9FYhD5eXly5jS+EBFR9eyp
zwHEcGC+k3JsaMnvAil9NYlv1zyw4cN2zbPQIkcG3TOvIp9ehp30EwK4KeuynfnJvec6WCEaCjkC
qs6f/uHYbknJLpriHNx6QdszJAPQGDTR1syCEjCykrJxAOrP+FlUWNLqOtmI1I1N/do0h9y1E3on
Ln2c7avu7Ulg+ltyjJJcE2X3Ctu2f4mfbtzSlMhHPPE8myhzcMUmFmPzCMHEupYaKcCS3AAnnHTv
yRGd637jhhe4ngTns9UGICW0+NPL/nZrhLWxJD3B4nIKgnHG7vQvd150W0lyjE9t4jGVxJXsnSMF
0xYgr3r4cHc2dSssJTU69wmdUx1TGZHGL8HP4kgnFN9gMEVaDSUOnbQT7YkJXI8rczS4dYQyzjpy
uguV0P8uiPdRHgECkNizaw3zcE2WBoXCquihT1xue21791v8KLgdXZy5FfLGgwFGDbsuWZnwDO7U
tj/57lbMgpIVLqkeuu6ZPFLFJZyRZtgRKy5XXPQg5H0wgxluZKujIdOWzBD7hkrEyOAL2rZwxo/R
re4pMO7L4oWGNG49q8D71ghRLheBBEL/5oXf6+NyCrow0a354SY1Y6DrJXITBuAjDRdK1C1tW7ik
1CZTfVzfQ2nobXRatlm3fmtKdEtB/r1I8cz2rbCbiL/U1WDfC0R8KfP7h3Er8oSgjplels1Vjxr2
L7EDtJgmWQe06F9OH3ds+p5XO8FsqNii0rm3ZwhYDUNMOD0kCdt5rkDqavh9AMudePYig5yF45i5
BezSACpQcuOuBkdNNYOjX8xGqMHJvLJ2DUU/e2rWRzc5RfDQTA8ej/P4DAdE0g+KmVjfb2zaghGS
RiIjI0yzn7HxEinwpRvWUJpPIl9RTzZICcXB94bnTA+QJrcHR/Jkt+m4Qod+aqKfTSNAhOyXPpz5
tjV5BZd/6/0BLgEVECyKMNe59Dv2+WH/8YcxSng1RiWs/RxqEV1xjj0PeMau5YDWkq15L7a04EUG
ARrsktOdsVAValeSxVewINGzmyLTo9aVx0VcpFNuhDUyYXbG2k7asjihzKHiKnPmlL/P+iqb118n
JUd0UpgLGDwAxU6l4NqOl3auoFVYmXl0txo93Y27hT4BHJjdQadEvTAPBL9Z29+Msyx0lvLvBqN6
nGD7HQeKzAhmZFhgpZlR2Hku6Lib3G+5CE0oJIuPmslB4k+3NSccmzuOYw2GukO++GyGHR0BVK/Z
I3Xqq0lrxAR/9gdmX2a2mOZVvSxNAhGAT0Ou64b6tWqCEtQcP+7aU8eB8tJU0gVkc01O6z8f4El6
yOtyFDbwZClqoOdDsO3XYYbOJPa7cCQCz67Nj7HFr5zMvqvKnxLFWmJn3/Cbd7p7E/BSMPsueZN3
DT3p6fgDs22DDNSyraUgI9+hGvdwUtoUqjvdS/HSGK5gtcOINxjcWvn8bR1cZ24BKQeGN/MMM1gs
ZMAq7TPiWdb6KG6uhj4BePMI3tqpcUu1SVhNE/SSy6CSPEXK/MYCK0qngVPzZ572AeBdl7AtYUP1
kqOtl50oBrdP4niy+VI+zYub7DBWrQaAxV9V8/Ev5DgQhULc72C0BnlOdZbG5PUEO7+rXL+sEnx2
F/mDc3oj1O8pRCeo5TzCDA2W4KcslSOHy+oDcoiEDdCi92poujSPJAAAw52h7/wwVBSyWbGcKvZr
WBr0HjKHroAcY4pCU8BkMve5efz5UeQ9oN5wUf9JBdvaYdHrVwOi0TdfShUO1rfIAQBf8BuuaoL1
3r4kIpnwSobWZEIOK91FOY0j2EL3Rckn0yzEgTDZLX1G6eXZSGKrL/Zk1IVTocbIYxFeeewjUdP+
ijsszjeMedCc9rXHmlyuYUYvpJTaH7CcTfAQvMF6rHr4i4AJf+tL4cTjoSqKcuRWyxj+oTA/6scS
ArUCLDsKaa2lvdF1slcqzbnZJE8Z1qfeuDlibM2lHLI1YCNHsVrYLNJ56lLrmHFrjgNeJds3tS97
lvVvjmAOBRDmisXH01qJ5yhYOfZzVg+dOiThjQlMBDyWMNvKFOs0aSZ5JTu6ZtKKVh23nOeLiyjA
fYgMMb9ONq3syrD2g+KcYvWsyKZg+LWACeHcqJOXyHlJLOkGsvY/pKUcpvvkOBgt6c3y2lkQw/Vm
AsbwfK/m4A+0Dt8iMXH4Fz9zJE1+ELb4+DZTLtU7JDSr5wrgkJ+oECa2RK7NxvaMMV+zAbXVS1sG
pmfL8EjR5zQS2JzT4ewZyAMIUWN+w7rQIC8LMdXUHWQOZ5wwbaJmVz6FSoiSwwmn9roI26NqgwS+
EWBNPIJ0SIbdOlJ5rg6sA2wcSFw/4N5JUa+ilxOfRxI53Obsmg16SJYCC7yg61YC3SYniktJ+sJ+
7v0PUnU4Eb7i54C8HhfJFTx4ZSD3FCL8niCwlxY//bHHVLGvgeLrTDaDaknKzWcI7Y+ESSFimnI8
MVAkMQ9RWDC/qhAX4+K5q98SCXkdKt9vGz0bXxgYSGIrzeZfvFPh5rFOEZEV31ZivREN7rp21n4e
fsYfIsqAzy2QHqs3f+CN2DJPuJedll2pIP3a2zcRw1laFUMQHQCYUempL5Y6hvz2wqQeDGjCyrWa
Z382xrMe+w7iwehyZ0Y7mdxVmzfU+cMgiAg9wImibsQZn11C6Q7XXPtp5R95Hg4ErBI/wViRYceI
QYdhg7oZgUdGBKsSkZPAAekCTjAplIv7J+BrblnobrJlNNGn0RkAwhk0bsMOwGpDSVqVYlB6srWx
3X53Zkz+shsx7p7HGpl7jPGzEVuwuexqB05STD+I9De6651aSTbySqoBGYBFBRvP91/0CcfR0kil
HiktlG26KftA+ipWk8DwFfxodKH28R+NNuQ32HVr7IzDG4Ols0a/lU8eqeGO0eYqxAQkLm7doKJR
He7SnyK+9OiIxZfhUbGWOlHQhFz5+hreUGEBnkpVSRePbq6pjEaUChSpFtgvbBATv+kqVjjaYOv6
cMRQ2XQPejGt2wQrDp3s+c5nzV4Qa2efeXxqkXH8WQmt3U2BlzmIT2Ra9zJV1rzoU/AjRO4tnpVM
3Hrq6mfeSd6wIUm39zEgnBlCNb9a5BTr+vn7YdrYn7mCNbIuqJd/lBV4ysKVc3I//qYA2Vs4Xlby
w3DvxaCXFowt6vuvzwnTKqGRFgBZRjIPbHFvr0QsMmHL3aE94f4wWQcUOGR5OssllLF4lXV+e3rl
aPvKzWIAoYjQZ7zxsTsbkAiaEdrEnAVF9ajmAae9wwaO/BnyhDEMGToDbcAazSvLFBT3T9c/c+Uu
d6rHL7PvbjQ9vixLB6kC/ozLZCyWM4kA/aZKxbKxH3Mejf10veu75keR7Zd+ut/7zjecK+Ww2DVv
bOYsyO3WaQQl/GZ3A0zJw0AvJSxhyMpZSJP7wvkr76TgYzr5eE2dKmdBZ2AKNONjbzwh7XDqYy38
O9eUNhZtbVa0n0H2Caafc2G4WsbZ/at81VRyYuBtByPJRP1/c4Fr8TRkLR84SL/5WjUSdkB/HAjV
mKYJazDIXtoKeuQOTG+lbzWXh7cjkzyYXKSAC0h/8BUZrUFHQ86bl9MpvTMu1YDpaAoyXszUEV7d
3BlKEw8IKCmFWirwgZk1hJzUYhW/oSZiffJitR8RMkZKUdDnpMfkDOVScbBFgz8NiXMuwolE/Ymu
7GHBbpknqRqsFXvcQiuUk2UIW2+yoE5umHi3pUwri0zQvBEm+pJ6fOBmlPW7KCpbF3+ypNZnZmK9
mc/dcRmsx1BuL0Cjt0X7tYjSxgS67RBXr/P+GaYXd41ogfP+Im3anNvndVUttKYO6rAUq8QXq+dE
G54sLJ1Vfmdk24/Mq67LEFCz9CQ3fBiyrnSG6IDSP/Ngz0U7v4VHomZsyXCCDnRejmz95jvshRW8
EWV9rjwQ1CZIIzEf+BtoZG3V4uhfw52NVTLrz1o3y4zQJvJULy+/lKz+/MhN8z1TJIHrAzw2KIGo
dT93GV3w10O5uRmRAo1Tih2d4+FMOqEI/niUrnmrKr3IS1yQLNlNGZ0jPQSPlH35Mb5Ixh31F4Sh
XMhbLmoo9FtgDrcjti7N9XSdqPZYYR/3PD7i1NNgyWFC683qSchfGUMI23wecDzYudc/j/1TSgxu
x+Vu/uiPhY9OsgKGAvkWi5vpgFMjdxIKImooH3TS9qbWosMmVvTf51Vgyfo8jgp5c7XaBDkytyKf
z5VYITb33pvvKSN4s1jD7Bri9b17s3TXA34u6qK/Bw6igYcJInwYh5ANi2pTWfrtxq2ZjBhxvoX6
EaqBAjdBaaEpSAykwyxIfLuYWzb4XaJxEUEJrln5PRqDcvkeVRvYeZwKsJilygj/VN37cXkVdA/z
ZIAd+qlvPfxre8DcVYYukXtw0MQvVHMGHyeB+PJTY5qrqJIKAJOEBfSE0zyM6n8WPzu7K/9/Riiw
t8nG9LaCEMYOKx9gH8oOXc+UxnFQrouAnmpLlHi3ZE30oHuEtkWUt5G4ObQBZT4W1a5LmCzlPWhN
Tz2i3kRd1ReFrUikCE/bSIAJnP4cq+HS8zx45N+1/siLT+tOuX1XArkZtk+V+bcTzPPyMnHp4/UH
Q2rQx3w/Z4dllDtnqnxgJ66J0At7bfoiRS3aDE91OJwXPmCl3eJhMpvhbSJdF37R+HrfOisUeXE6
GtS+ebpIwBfNiA4b7pwSFB/NUTh/AhCNVxyj6qoh3wpAyuaZKEcP4y3LhchUYdx0JHxjCzSWOn1e
0wtkswTkpitlZMyR334zPP7oCZdsAi3z2jfNa/8WmbGdAJwQtvu245oxuHJkm2t8k1xtccXESOGU
rpveEbAgsO+J1f87TgDn5V8sGUx+W8G14+XiY7iaK8FFxT4x96OEgtPjF/Vqq40VUcbr3CHgfGrL
8tFX5BFsoMdyCeDxjODov4WOEq6NkzBacWQn3DLR9H5VNyzMLAV3pV+8nHGARpvI+MtGjvwGZhKE
9w71pfxo5zzzyX9SOaX3gnWFe4pLozeEwLpge6h5sIJIMKRcaXr25kPzBU57ynPrROvVPK4lbWVH
JjU+U26C8bPHMY6bBLu2Hs8arVS1tyLk4Z7pQsI25l8SLebqmE9BsGKxjFmwohMzUF60vn3g/R7M
SH8sBYBoQNxC2GdCjWGJa6dv8pmzNAXHj5blUL/yNbAOWyLE/T3H3taaWO82p4qYfBqoTFBQGeQD
xXlR2xlDNpj3u5i4roVV4JrNPqtNYRxNa5pxFCnoK4MgfcspNsUPjdIrw5+xg5+M7BtH9AxWrHmw
lBPpa48qAl5oS6z1LSgu7tS6f6ODJE5tfb9bW3rGzMxLbKlBqBaSKtkciZRwAHWgYJIhSOxIznZ2
BAFNg6CWNq97vq0PsnwErfKycRKC5H8cy4uS+hpV+wnSFrav84NV0QBQZrrG1RvSDAcEErIUqkQm
e3old5xhNL6broDBHjNpZ1tgCeqVOaYz2J+U5EO+ElF1GKjLCxyxYuGC1M6QxyK46DXWoRUGlwfj
z179tVzpxWbl81prlWdJ+V9h/wgPG2VE2+0LlnKqJi4k7S6XnpFtQKtH5gOd35ekY2fbhXzL23Db
03kzk7z8MwfCTixiAtgfu0bxnp3ICBEOjZOGVvgXCKUQvIjaJeyznU2FcW1fTOQ1SG/iixF0Nr/p
k8Yg74WuZLeFy+9OVGZntoTu0F/4O0sIo1d23L+rjuLumEx633gAFpe2IMc5KQXDrW/O9OwB/lcO
4L3RjPfcdq5OPk6a3ZZZnYyN1bKQJoPo0FpnsayZGR1cJeFDgttoDd1ezqwEv+pRH6vyCnaDu8xR
jWN/Ey4J1Fg/ViSH1SgNpL2JPCAzr9B/2Si1KBb40e7SBZaugmp8WZ0JaTAsIfSQ/mmVNeLaadrQ
v3ZAlBk16qtF4eyUI1k/PCE/GBxBDSaGbj4RwIXbUaXQArXLhK4/SI297keBm+v0CPH+D7WMN9Lg
QNdPB3dmOvOgWoR4Y28A/MeeCIiASykbj3X4abYeIY5N/1hny2ipfTxil3LkG3557HKzu4jFDLCd
8EWJK0CKCLnTh6lOqUipfsgknBv9hjn17o074OsibkNOOMJ16ol3eDcAfWxbLDV8OjrokPXDyfA7
JVOn8y01EzVcRdJLQYBOWOUE1PdCjmvSlYpqKjm9SAqVz0YNaaX3S1leWm6cnjabdqxsDWZPTWyA
xhw9SaAUtzyx0UXQ64VFwbC0pP1SXIBVmTGEI8/WjSFLsnEIEzHJ/shtIoB7k6NI/5fZ5T7vPKTb
eiqBW9WQb4oFHZP4tFIAle2xp+MkiIsIe1dkZVSbZSJHoLk/fQSh+NQjKg7XF5J0jTkP/EBf3uAB
noObr07dLMYipFkDxDdCnHUh54Zmpfu6UINdXegGGvA4POhmv/JxMMD32FpQ2QuwXGZLIY48N1kZ
cr7mftUN3jD+04fsSyU+KwgscSxI+sm3oHoIh1iccgl6drDsiDG9kv8x+cYNE3cIpgGXUPGjDamn
rFWFeEU7nyz1bOPldt/TS8coRPeK1As9quB3GBVjgpr0KeUFuligLZ0mhe5b2ELwv9FN49f9u1tg
xDToUWwN+rKpvBJ5p4orBdU0zYbdFA2IqC40RWtliUJSX6ehNEda+f/2laZJ7tsZXSXe8ZrLZLso
0YhGc0LlxjNcn7fsc2LfeITx1H/fp0ikar9JcxmRdyFKGsrTVfsGnKn6ue9A+QsDc0c4u4xfrwhe
haGB68KCCXj1ytpssCeGOA06OHuUlRyjpgkG4t8RM75YIVSTPTmVC7GsLK49wHtQ+9qkFIxo4Yz0
eqJX61LPSfYWtmFUz6WcAsQ9lm3rNFn9vAaIdCK2yusdZr7BU43XWh26f/8f2uhb/9DsCh3DIYUw
T7XljNnDhXLjS13TR75NARK9iW4CDj6lB1hmgjVXS9EDX527qOYD1od0ZfX1Qq+wLg0M3M16NKgh
QwRJ3e7EwdyliBChwr2OD+OSyjXBeBEOrY4pkW5B5Ej+9AeppQGvI1W/hifZ3ARucTeMiNMfzEFx
BMHNaQBCHvz/yv9fy9f5ReWu+qOAXYFe02qacRYDwvPFNvuxCrQGXgAMkecDBkaEg+xmZV/nzGWc
+R+allVUA+2SjGk4iOCM35XjoH9W9xpURDYV1UUsS4FGYC/oE3+9niB3eTxS+H8MbFANOZezm3Wh
txING6T1Q5TvVHz1fu1d6ZehM4SE4KT9SYNlChOdoW1W9DD/nFXx8gWt3xw37rkB7OXOmFVxAB61
DmGGiih1bLRGPpgjl4H0V6rKEg+ECDVVhp6cKWBOY3WaJSGtmcwWOTUc5ShdMOLUdAX29j0VcrDt
IqMWjpdUSqtiuPQmL463okwIikouyoz4AxfBVzRSg/+y6LfseggxqrPNPFaKP22q0hPC2v8eSixG
2IGdS8ZMZlaxqSsN8b8aOG7GvLmTx3cp96mf567I+bCd1HgX8tmQ9H8c+6bkfP1KmmpsTyez5S3M
AG4h/WZvNy2RlUY0A6XaqXfo7ul6+RMfG1gOaTYxLJ68Ej3Qbt2cgVr1a89JB4qaroS0fe4wi5Zt
e4tqN7Og8ZvRSofED2f0SuOw2FxgmwDMbgG8eKBoHQMy3MrHZF9d+kUlk7oVUkMNWDYDy977OnDd
NuOTdYWEu4JE/VnWt+iLPujkXI/xGPtNbHn2r8Ifv6exkZNGXl1NYfMrEaFCzZ/Caqh4G1Y5QcZy
niqNrzarz8rajPMDEMZA2Svi3Ts3w6sRql3Xn3cDC/DHcFV5LI4m9+5lG1noD1dIMzC7Z+D8u5NI
kYJILjNTjx6HwbbCUnD2Aewj5oCEZgCsSwK9t5c5kE65iQX0F1Baw/1yutFOZYDZuZKYN/Vw31ZI
QrJrowx260nW9WsoSAmzclnfgncc69pXM1T6aZGq9WSfQnQwstYt9kGxeuVCLSYJHNepbzIKE9L4
7X3t5PnH50CTI/gAaa42eXnyPS6CKEG782b2JjYbVMQZJDysBt7+bwpdevKxy6GQHP1q73XH6ia7
hBHA+AcPpWsWihaXpuEmLZMNjatsnufY1m75yqQGf2TYkIeeT0gpgYWwrcRGDpCmrE5NfWFKFAaG
mNweSGkC26+S60xt6HiKYsDdFZfjhxus++nziFkz0oocmmUXcExtDlt4O+YfAao/BqB2abJv7u8A
Xlaq2amICpYsiNVQ8QRlDQh1ILn8wJqwPxdojylKo7Kq4KhBKiRPRy5rTMBzK+49eDs86ui7ZVB9
wHCLv6cfN3+9UTXPp43OLEa93rKTu6sTmExihjslcjrHwmzxQZ04cMDUdLZ9vr/Fp9H0ZyAi1Rel
oaRHsRJxCFpv/fmSVj5ivrwNvbA91NUHMDst84+SKP9mE4eR4YRvaM/FfqPtE+ZdSf6+Xo6bwRUr
N9J+oTsIE+4YdDmbyVCmlCz2OQ6RLfgQuVqsUE6BoiC9hK5UD/aISRmukkaiwvDtg1Ioskex8qL0
0PmB8hhzfqH70Pt9F1MuhqkGw6Z2JcJafwHwUTzuYeFNvDnjuFJwLuAkGHr49ZgbumYwLLfq8bDp
hLnA2jpiaYw4uFJm0yZpxLA5H8OgeGO3lsVyOjK1RYBE5KyrjpOiVCiY6fYgy/7YBRvriYrj2TAm
p/gM5dJKRcvqk1qEUCRlYePvnaTaIC2GQPocrzA5uakVUYOvKBmvdKp92PsahvrTosVxrgo2AGWU
wrVrzxHQlg+Hdm1Px1VemliUJefoJVbD7+4cQhwaxk2XE2MYnptJXD/YLpMryIc21LNgMKzEdSyC
vq/H78EIMRhrLCCOqiKoAvpk/Vjt3qVeSPOQmbzbmDKN7UTRv0+VCCAgC0uPMzK5KDjiN42IW6Gc
qeU1oiDeMs5Z+qtEFFlkpx5XbYcYDPZ87iA/GhFIx892NCLMie2drMhB7MzruVypP/4OyhzfUBm5
PZA6dRCok+WnHEcKTu4Ji+RcLY6HlCOc6K4Tw8M9dSC0JA4yLNXzeqH6RB91sajdnpYswEPQqInU
UqtsBi7Pv1Kv5Gf8y3rILK8s1xQz94mmmhtHFV7kAc3Zre/ozggif7EtDG/WzcEcEInWi2x/P9xD
t0w8tDCkHuO9f9S9A4ns9rXCUUK2Nd6IxjYSDSuFiTBz84ihxwYdWm+Qk846Tg+ZTwWVDCL65d2l
CpRvsQyUq1jLtMxETBqppxROtoar4dJ6pzzrydHzkT0/wGn5s2QdyqFH50Evjb4oAJOceUKILpWA
HJv6ea/q4ZLRnxhbPZxnT8g8YW+x0R/0dUqHffurFtO3wzXm+PkcuTPNC8dIYdOPaeuqT7mn/9D+
k3ww0owUl8UPecqZmLVYu6Bd4mpIQLGuOelL1ogTHOzw3G1cY9sIz+EWFryUufLuuYPkrhMOszXM
eH8sB3ka8G90fWkn96VYSdHjVQpQ3WfqhPMkMHq+pzPz7YzMNBrFqpsdy79JBaMpnXv/ShM26lZG
Po3DoGbFLCvISOG3lQEHfPPaIHszuecvT6KtyfXxS+KsSWh0lKq/NPoC/s3ailVoph/+OiIDwD9/
HghfQrS7RcpFhciXUVrsUbMTlTk3UDmAq/9dvJ8br9LHavA7bVZg2cobk7K3YKv+aJjenADWMZvl
NK8sKtX9/0Z5u1z2Ydl+GxFd41rQ5ZHdk2KXcHzD0a1jYjqqYwGxEDz5BoiRiBBNIOBcqrJWuwmr
Y454VRKVQdJpJe/HoBjJ31wkXKhReXncNusH33Y7uN7Dhmv6+iXBMOYd98vvKqXYJoQDQlYDQZlr
lAOGk7itwzavxDCeQuJs7xzZVnsxU4SKU5Wijp7y9NaCTu83gSStbdUtvLNbPIj3duwvC9hu1SgI
YSz40K4pOL9+lqGSh64rhOcNQPA78Y+A+GLFPrSO8hHkKSLvJQdGzk8NNuBVbFII9q1bI4XSm2CI
xfe+/V2CC7lyUbud/72wwmTckMV+Rb1eVKULA+odcbDoqt673jnSiOdDdRFnqUXhmjZesRWtQHBO
EHHBaZlwkLo8kMLiqOCisDvD688eB28JBFaCRdo5cwkXUdrwIyQyJNZeRWZGfGPg9QB1WYozXpBw
CDhO8QOFHJtGZSNfNGSGUoKYaHYPrT4DtcvQj9T1FwU256WkzDcb/Wd8is59IyNxvnjBXhkG21Ba
bpbuiWrqpCS4fd8FvCwGp3HoRrfGlPzP/dVCvN8Kj6DxyTivC3wWrUZA6+ebTeE1jWrnnJ/sibfs
dhvmjBi10+C3QhTugNMla2K6TwK7nYpN7l5PxeIGSbEkabr+0BJgJgiiWFtFnsiAeqAvf1Y+eusS
c9f7Vg4+bZpL8HCJtYrYz0mf/m9Tako8Z6wZdiMwo/BHMVvYQYK463yh2Uudmg3l1C67qSQHl27g
5YreMO/NwpvcH7BysqIRNJWpgNvPu+5B3Ye/lyQU33X9NXnnmm+smuy8B6vdaGfzGJSw2uktyQAc
JWgmTQZsvNYhPCLDBlDnxcbcQXVXL2HVkTtOnwsTuq0QOpbLqKVsDJDfFwijZ0ojoKGbJibWMmaZ
hEMj+kIgAxLSXAX6+rZxzw1zo2uMrUDyMAkouuU4+V0FeMQFLjwIEa4WqQdJ6eT4/NidpzixF1MN
tguinaVyBEbZyW6WnTxIhzQHqZlAA2LM6hlQep+qPZdVTn50DgVHElycTALtIARaAWLG0ex6KXbK
OTqzmZ/1U0qD4VlClLbmBysIHlI4t/3B+VwOc9NbBYVz7zezMbhwoBeotQJ9a0uRP+DpGG0n6LfH
6WxL58dSHte+r0H5yfhBdM2H+VvaJ37LZKfjX6gGF1ZXE9nF69VzZmLmLs6RMoDXdxHyGZweFoq4
1zVaZDFIV9Oezlbj45QRv5fxap9FkGS7PJmHXMVGfEC0z1deTUl05RgcQoNp+VpKU0ooyNrV8BJs
jvhJdJrAq16fZgUpMSN++R4g0RN9XxMYOuCimkY6pQZorsreykyCXmkFRTFMbNnD156i9sprDf8T
jUsCLacl0Wa34spXKcwvyP9oyFj6OmcHGPgDmeHFYopTw1YM7F6L1vP45Mpc+J8loGHtDAx1bKXi
6Kr+LpMfJL6eqKF98ZqwfwRhUaXuD7mgUnbj9X0Xu52rmbbNPm9XYY/eqeHwTpARV+aHoMyQvVSF
cAPrH8C6i+T1wbwVs3ofXQoxhCMYQVUxW0SMmSLA4js6ft/2T8dwV+vEg9RaaJBF8Z+tzi8++R+S
dLFDAvXbv+QnkgIQRrMuV5uWwEaJHojRjrpKpNDDK4f3pnkO8H2a98IvP/1MBSLnBoi/qoXcIJWI
sFseCyzsorj4G3dSB0DHc7DeiKdtt+YAyp7HZeVRQx25oTJO2PeD3fATUAX/cX+LjSiD44LRf7qI
4vMwL7nXWVtUe59ZwFKkZlivZixc7oJV5X3ZGLcwLqmIiUzBWAMM/k/fYAbD9rWKNSQDeO9GA1MJ
62E+TC1CvXHBts24/EF6mJlrxIB0QqjF2/WP6/B95Fp6Ao4IyrLqc0BOiDy47vw55210zxLkeqAR
jypUTgQnRIzXVCY0CQXrd2oFSx75PXSdcoFBAHP1w4yFy1rNTmNzfGxQmrWvfAxsJJ480gLMtPNY
HsfW3twsLKDoX5hoSIDZ+OicQWrAMWu/DKhwcvaTpxNSaTOoN2SjUmM622TEeahMDh7XUaJPQsM8
rvQ09Hp5O341pbZq4vocRQ4vyvcU0H4sbxQQTDmeY7SClT9g3rTqHBVYTJ6UBRRgGZtAvLWZFLzb
zRdxFYqloMm7yMejjAFz9zUlVk6lZW+Ukuvi5zGggpl1kE9BGZEGnDrTA4H/ANSQLzP4Zx5R5zBN
3gopr4CJWr6e2eIC6bqiJtKs9iqjKMTvUxR++/2X1tgDS2CanlqH/Djz3eWux4KyDkkfq+2WlEuv
PU5uxh6u5OneFzKsf3qhokbllMawrguwJpA4AAmRIk2K/ga18cQ5C5+aW33FPH+cwADWPqNM64Sj
DWoTNHe5qbt1zPi3kovZx2NSUDQtFXfqIlGaS/rEWJym+yXfYjPAn+1yyPmdAofSfL4ZyzR7x2BR
8JEUCXmULAX+UD2QMJxsaKcDK8JYEXj/LShHNz/OmKsFWZkDiuve7sstjDak6fuUJcjfFdhY6+1m
/FlDW05E4xyIlIBlaYZnJc6d21sQBl+7RSBtLlgGSg1nTfw3AAbtLMJ844oWwVKYW4hg87xCXDzk
JnSk650ZnYasOgXxdw2r7zmycTGeY6pgoDXyd1/vRswgmiVTFYz1VsXhH/kdXT3f9Z85HlBzxPGO
DXmJh27hcuTdoeAvABDZOkkXdCIdpsPg67KxaGXYMoCm/2TxtoPj6vWm1nBisngxan9TyXBtLZb2
tH9r67xsH4kj3nTtcTFcVtF3aM3eFSFJ6L6YKLvIjiHQm/9HICS+kkQvUYqJsM/RAyKBGyNZTwww
IzOGD6n+SqtYld7WdwyRqBzfrGJVbu1n3c2TXKTfzlexoU3Agphi1ztNjrnLNVUibNxLRWNEU647
bDZ0q/ludM5k9MBAW0bzH5tu5sL6s9fKr+SjpmAPgzDj9z9E2x/2JblPT5/JjPwJKOvscCUpO6lI
GH6i+fnEpl6R6yaPFvBET8IDRLH4ubVgEFM1RDedpJ853KVLx4SAdT39nr7GSAn1c8pD+9Db5shE
4wBquqzrgo+DXNG4T1PgHZ88h2yW1kKO7VRCgBrud6co0IEs/CdtOo8rYG6S7rxRJk17I/dEvkjY
tb/jAbzdwyWfv58A7iqWlZm2xf1R9++3Gy3V1UkcJW6R5O2FFGaoE8AW0s7jJ23abHhYv54dI37o
/EVXh/p8JDuY/y8fmHhIir69S2QzYMfXt41q3Jiaf8eEuo2VvDNhhJRse4DMWFWJGpoZPEQVn0Ai
yynQrR7HndQZXOYbdHrvrHehvcU0LVaN0bQQsGiRoooECiiCtbE8W718WNX3BZKB46pk8J77v5OI
HH0wA+TB4BIosz8KuPF7Kvbs6TGvzevEf5csOx/UEpZMGIuT9jbqZQvabhB1mwGr8YoS94XlYXtu
wpNRxtUXTsbXC/i5l5JV1eNufmhDmSHqAqO7/sHWumoBxrwbbGXBoDNXvqKXZrFiL116COgFQ6Eg
AXr5/pQjEMuUUk1aVkHJcN8ePXMxs3bvUEjpAAQcjAoYvKuG6GytdRHoTHMs2mR9HSwczdPxo3QR
QEuUTOJv6jqVcsf3s3QgV+cL5t4TFjxBZ+fw4GX3eVd1WU2sPTQ/kM0ekoR3mc0hkkoN4ltVxt6q
KrrgnQQq4MDRQpp9Z9/mHJHDrbyGFb0kCNDtpHXpZijq1wlMKF7rIEuVBxBchQiYyXsueEWAzH6T
LuVLIKG84oFvK3eMoqrpPXhhQipYHRmm0nl7KTxHnNavy/o1FkrtX31lc1mj9IZqmsJmBTVuACPR
xsnQrwvhV91wU61mOkUknFw0DAFKhLBlV+X29zkhwkVmhT2R0q+cRgrbWQchlC6P1tG2upV1/wKK
D5spQGUAZo+7k0U8bkhjME46PKIJ45zbpyp54NuHXaVT54ZczQOQQpWNTzdIBW/+2UJduO9BtsG8
MxH1pjE/j1x7gCMTM0t+s9Kis4KKOnFZSn6pxuRW3P+/oWdhG7fNsGq7cTOf8lyWcA3N+RKk5/Bp
RVfYbEmPq3CqRRT4BViHVkJZl9AD9o+lXRiOwdS83R9Z5WoSlvhuJ4VtKUgHt00wX6tFj/I/jqDJ
V8/IMXsMjz3goHwTiIUWxrJkQt9eYs4usFZavSpFjv1RANZUGnkD/6Xqm+lqBFSq65WXsb+SceNx
DuZ4tI9gZxZ/R+bosyS17YWrm6NUclMYUwmlmmtQmOyMfqisnsiCyXQ+H/ECHZf84mnw6QAG5SIq
uepdgCC1im//hIbsE+pvRMVghqUWiMSrDFp9fo0LKDIB9BpM0NtQsfnQtZ7e7lAeOikWd+KoUCTt
R+/MxSMc+NZorrAdXGWNrpjCZEAMAPwF7GYfsruGJ3C62fmryhmLznzNgSxGyQ1cURY11+XjTrPr
DXDY63hFscBAVaJt4zQOCCG8wxRNiB+KPrsB3sdA+ASd2l8lIKPHSvSeMBqS0cgcrrMWbXlu7K2Y
gwGGOsG0ve2q1b+T39fRDHtTQXnk4JPJqL8CIm0lcjPZ1MIy//oVA77gkGj2OaiVDDylf5KFC5sl
bV2pHOHVgvBZhNi95kTuIy6rSfEIBoeIGKO/HRpNYpzir63uJjoaN0xu2DEmIUG6q4eDSmomviQ0
nmbJf6nq6KciCTNM4KrMK7mdScXGgs2g/kxafz2rKiKj2UVVMQ/GqbeXTL/jcLCmrYdRGZJhiZfE
/lQZxA1LFXL9gJwIyrsUG7UMQd+9FVfmaUKTP0ms+uPNc3OCEjFXbFSgQnyepUjDQdMnZTNz6Qjc
NLbMVe7C1UI5kQ9MGarsVxVsXTCQ//VqB9sczM3YHDPoB5cSPLW6ESwDEUlAeOFRUtGduSD/u99K
4yL3cYQKdLL7YI21LaTcA9M0RJHzWCl7HLmzaqS5ILSDNPEaQsxF+wSThRnkIw8GElhdCV1DcY96
18ti5LAXPb6eh/gkeyv3k1VKouwl8B1l4HeVlYb99m0ZLDHvdcgPbADipHtKqQCJfi/cvj1D5HB3
DVcWjayIT8189DCNagmHKFjGMWcjcPkm3Ot4tCUmIy0TEU9jQXz2ghUVdgJsa9p3MgFKkDaRnIlI
H8E8465YH904b9iptvht4EBFaALCY49lHnG/K/TmuBIb6K9GFNWpsaT4R5Z+j9a2a/XI0BXGn7Qj
j0C5fXMb66+VXz7rKP1PpMyZIb1MUbcRKo7DpU+vfpf5MokNSlkD7Yv7y2BQhog6hD3M/SoBt9LG
VqLklYYNUNlF+zgJJFinggeTALktR1JUxUE9FPNUeTBxlsuINxaLoIWyVygPW26M0AyeUT8ljmIO
HTDZpTp1N35rv+WgDC0CxqwuwgsvB+w37jKOWcG8qzqKVDIU1Wyx2ZOE/+wCQxTUT/hqAkj/yoGy
v/HPdZIQaNxY+9LI+9PkEYaN3PPL+xevOGe5swOfEGWAIGxSKF1qkQpD4AqSooGRXZqPa8j62nGL
tOfzrAoWEjqbyx6loMNM6PkV+u7eeZcEqOQtRT0rfsnjHk49wH1dSmIeQ1HlKkcPT3Yl/niH+Jqy
nX5TRwAauqNJrjtIsGqNJvCDmhvUfUSdmGsppOOWxdBqIoDD3JE+Jt2hsw3Jt1A9qdxCbSORaEMf
TWibZsYV//3K9q1yDJXf8RrIatEhOHdB7xfaE1XquaPzHnPKUsVGlVSlVCp6afuya2x7OgwYhLkx
rjPcRypSPBS8PMvTQ39Kr3Af6ECKmgg5VtlOuwkFDkybEFCNyC1wpYcseuLAuSbDrdJaFu+RErlG
ttFDryJchd70S1iI11foJ+0DIyv4XELUzF1GBCleEWlTTMaTSgwyX7VdSaMh/BI2nZRlzuduR5A1
waZ8wmwx7yy3R1ikgoGR/66XE7C1jkt1KLh+MvstveT1akbap0sDmegUlub8mDE/xzaBkyquKybE
ZRBKjc1ciGrSyC8Vm2DWdjDYQII2IilZVaHFs6SvHjYm2Eyk/v7643BgoyHaRU/DPVpsuNmH5dgR
0H/v5AkTmQM/DTHdlBi8THUMvVxWwe3TJAUwFaZO8SpHquMzXA9ITC1vC5yd0fgw5mvUJiKuOs18
MDNpjql0fiM/BAmVgFhCHR7LJQ4LC72RVi9oKE0e801TjsFbmjB35gpi5w2jhEQt8V70mOrGkywG
MA8MSalXT0gtYj+rzm44Lra2bfTk3c/gOTBLviIL9szNe9IE9zn78n1KLUWvO9RI0qspTyT1jZzE
0blIEX8dD+gyyIfJiMDaZf2iaSS/MP3TJPLb0B19k7M9AN2wGY/t0PrbpIYjbthZj+qKw1JxLU/Q
5VQgwAszqoqFQ0vFQi3Gq91vsf5xYux1i904I99cKB2jkYNYE1Krq0cf3MrVuLXd7MqPeelP0csV
0jh9SyY2E3Sp52Gdb5VQGTfvMVQ0IpVXHANwv2mZSuPhkrYRPb5pUibuyvhCRMBYUTsSXDfcUlva
8dx5q6hgtn8FV5J3sfgk/7JzCdzI29UvFPub2PSFAzbayYX0j+GMJKBGq1qaMQZQUBz4xMRCqWMc
aQZSMYM9jotnC8Nav3Af7mAUeTC/emUMp8Vzk2DdXX+XcRlAQNH2B/tA7t3H+Fd/ColIs2Lu4aTD
3EEIM1YCy7M42JRWkb9ryH2GbUI8sNKBVtRGW5AAKJWYhfhLOyyFVtidEsfs5+AQOFP+VymndPVF
9bpX/n/FXmoSaPPJtXb5dzXfrsbL/cXuGhQFIHtMn7hFsia0pBMeuIpR7wjE58zftK3kbOO0CZ/e
aJqli9r9qzemKvllEwqwPwcp6H9rOjscQXXaNxHRShZDjcUH0eN+MVDFTJagO8nte1W38/UaNvSr
weEMwjxmMidpL/X3FZAp3NbS3hOAMAbK9L5yojMc9aFC3ojwCOqW9BY/f5oHfPSub9V4mfny9SE8
nIghtMscCa5HKxIx+E4yH63J80qkE+bSKlVxBHDWe6Amud3O12wNGpW2LaQ4W5L4gvT6E47YE9HJ
C9x7lfSjKGXRp2NW3mmuK8XrIwxcgs/1n5lCFS+uSnHFFJlP1CnuLNECRJhkefgxVCfn1NcPQ2Zg
u6BQ5aT2rz4DEVjUPGBmXg4EG2OlvZY3pkzL1w6ulcx3BWwZKHmUra8EOzc9wKPmgCvR/KNKWB6w
4XOw91XfS/JtCnDZmOTLqx49BeRFeNO4tA+nQJa66BBwfSGDqlvv1bxtrO9V8ambnbbOWVtVWhg5
fBq0Jn+nUFQ2WZhTxcIizBg6iX88ttUOhsIXURGxC+SoBdKlEy/hEGnMG/Eft+glB6rrCvmVFbIT
t4MA6gMjgJonMQkeCZhAD4KUjmMeWYQArycOPz/yx+rcGr48xrYOkXPriaRq7pKLDrJRTj/3giV9
b9JjfRhoXY+6S/qpo4dIFb+uO/obJ8ruTnkTJDUGcZ4R/CLJMQ3+UwR9oLTylMimcwO+jrLPMUVQ
UUWuQhpSZDDy3Lx7UCtgLzo+FWXDuedE06BSCHjxE1K/DHfEiYK4ynGX7TmUe5YWRbr1E0Ws4Qc1
4a+TUnZiWqDpAHKZU43s94pPJnXgqTVabIxBRrRfnMtL2X4qGnkqHNxYDPFs2qPWCQxaXw4oXM7s
Q++8P9onasHAGkZvC7zQeAzPFUvMUWR5O8IS6xhwYnDF2Jy3XUqctlzeUmYXEr5V4NPj0LSyMKW9
uNCl5Ya4ziR8q+OexJgTtXhIKp9M1kH2YWkcHr0Wl71WiwKJJDvOOvLZMEeXPXPQ32pMn3dMToyG
7XFeVdv43tPvearwXUxg53rpFQ0MjIKnbAxA8y5vOlMXo4+IKH8r/3xadHblNcSVxSZbzQacMDAp
oI1urpqNdvMaqX8KkqjJNRw88dyZYRWfDqtuAVXE6SyCBxX1c7+ficUIG7hzkx5GhwJ9TTZ65GXF
bn/OfhcJvu8+qijtQC6PFmU2FD209ZWRO0vno9e7DodDxgN3dgMRAK4WBZgW7jxNru8gZoRO1u6S
AUx+WrL2Q9wI8Q61LjXy44ba8KZfDiLgAY0Y2ERE9abcJgnAmtTQTa3Qi1z3P4vOMEZqw+gbYy3N
76QAi8P0eLS/qK5Fm61q/lcATk/r2vmCT2leK8YxNHGO3WOHseaFpRgO5fKsz3q6NW1e//gc3F5n
ASVNFdjQUsu8OQB+wm4kLZmtzMoc/vhAFeps6CVapYRaQsRxdZT85TD1p1DPQ7oDRDBJhlrCoCpT
YStCY3AuVoZmlytGAfuvduwkY99TZsb2l9oYIyEpQ9m094qPn6r9V/KZKogkIlbrY0IFuXq2ktVy
lkuKSIM9pHalCdaqoTG8tViBd0FVqX47e6OSyLSUFte+Tem3GZbuLr8txlrgsAlRqpBJn3lpgvZz
cdPuLzgwAiWVEsrGWFW/sK/obKUZoFObvmvMSQn3xleETMX7wn8qEKyTKXqlbyzJhrnZcoNWxSxQ
P+g7YtBQkVfcsdZcsmLzyDHFDBVfyoluQfg8hu7rd+frpU0+lyKuErljvcfWXpMOfOIv9aj8wPhA
ndFut17AP1f/Npar2Zg6imnjI8xckENlb7VbX4BLK/Mljr1h5tfWgNJKLNcCKLyxnQ8HwvwP83Mi
rUAegHPpU+nS10LRjPDoEwoEsaE9Goo5X1gzXRWLk0qfkk+hbx3+gRsi2+NP0XFD8g9n8S7FxPgA
IoKyhbGJLN3lC5C0eaBd5iDEWZUKgX8WdHm1DPS8DdzqrjepsCJWT4R6FtLYw4wmfUsg6fPMUY6E
caSfgF/s/gyFosfmkJ25A5d0JMp8qPk3RgLprAfI3i8j3QZUG8gpcCRN+TCMxHvP7Ogpz4APdL/u
k2T8vR4mc4nLi540AGaCJ4piQhkt10SX+N8SAcFGIu0QYNsT7oPrK1A91/f0+diUB8jTMJFKU4m+
jEHCa5K8YEf9dpQm8r13QWhAmWFCWvMNW0NRIofiQ3gLcaOS5FCWdiHnE3yoik7ajG1106OhlFpF
o5nB0QYEgxaQ9fFeWwLtU5V5PRnS9s1Bq2QTdW40EO1yod685g16pgaSMVZUMOHV4csKf+8A3HO7
Jtt62+FvKuwPuoA7cxOUhRNKY+m8VkhmiS/y32bgnzBVLlAhOPcHkULlKEdJgAZx2YjhcJ/v9PQr
QqCvWE40HsGy6eWFTZpB7s8eOeMd0IRiP141aQdJdVOa8v27r4Bu94aOeq+sdhw5nCeD7KRHD0e+
aVk9q/o7EAz7F25hhpety568yM1vIRxPPQHiEolWDfqu8w7OveIgaIXWHAqen2vmYFCSmL0LYODh
wSK6Aqs2pHzGp+B483KhlvhzYe5zTokVnIriACzQMRcg5mm1Evft+Qahg2ebtBvO8Q1/ehHkMzx/
2rEVpfBO32sjsJpzE6bUgf7W58p58B1hkTb8rcAnY60Y1CeGYqa7DbLJwWSfAw8YlFq82Xnyi0VE
cvRFPBHLFcHe6aRBwXfQNytj2Cg1bAY41JG2kcEeO39sFY2lvlcTjCAxuZgrPiWZuuPQK9Dw3HeC
v06ZF/10JhnXhzrulimVj+tamg3Lv1duI3ZDM73nzaYi/Y4LRpXfAYnaoh4RqEDa3k4TAZp17oMa
GANKfpHwrShcGxV7vXAPAy0kWBbQOQtmloAbDWj6GKOu5rL1lknAilX8PzJCnCisribyZ9SmAeIG
N8qvKmIAAo73lMeWNUG4gK3OzVmS1w7W3ArGx8UuduPsCOYPLMcVKXbW3KmE4jmNHtNtITKBdtgy
uuM42Q0xqmwTkiKuy67yqKQ0T12jnLOLVglFpUeZYCgtYS8v+JM8+Crnmek826P33WpaDpoZ1cfE
p1GFgAaO0BSLTGk2X6sdKEykauBGdkEheIAc6T8dbKaVlCIBh22WYziHu/JbkiELHJlgZ4hzD3oo
cTbtfwlOx9whRrSjoXWhQx/sko8bHYLBkZI+uZnpl4RwIjzeh/bdzkaKkEX2BGX3p7uaIVQU7NXu
8o+tr0ICSrKcQhVFaEEdUatZvJJEXsITkBYpjF5gXihGLIkET3ECcmhPXjskbkm05nuayRdr+k1H
2oO2qEjVrF/SBxDAnNo2gkCJUfpqS5Qzn6GdA/RHvIxdLVh7STRHQpYjD3/m+eOx5C+C72/JuoKX
T3lWNkL1gbAtmxtTLWxQD+DKz+KSyfSC0ApMWc5TM2jGHEMLCh6NtZvW+A+HbJUF2E9Riy1+63Fq
Zk7buRXGA+7w0HseJSjl7QRXJbc201qyR7DDS/hhMTwWwRYOZ6dGpo/QoRMV+V5t8fG5oexPvrkI
OB4Dh86FOxyGVQ3vx59r2CV1Bklfztrk8+LwgmvuzpDG09fd1FY0UTFwxePYXvwjOnaKCknanL3j
lc4BBnzcWa3f+UvRsHJ8/kCJlWY8/iblpsHfS7QhuTZgd5kfziT3IV2iL6h/vbml3CsAXJ8e7Yty
oayTCWgmIB7mDVv/g1McioPM8kBIRrKf0W6OMyUrTAwQ8bHHkRDOc38WkFv46dSZ0v2i/K5uXi11
O+FyqOBAYpyDdHKR+BRSCR9aJepCOjjNxwOmhnosFP6K4dWZeL+r+Wuuo9qwge1cqOy6rB8nXYNV
9hTZvwNbzSc/1nN3r+2CU4ipxe7/mg8bw7wuLs0hBZb+KnWB15RK6FjfEm1sfEw6xQujws1Oicys
vrKoJ3CmMBYNhA+mTxD1XI0++AjkL6QRJUqMNdKjcKNJwifsPer4UEVxkpIcnGRifPfNABgYzxzt
7oERZY/FQgYY4jLICyxncS47ucSlOpxc9jNIse7dfxnoUJ2VQtUUeEQ50d7FFWn3kIiqiwDsO3MK
ycJ2rcWJQIGCE7MIB4lSeD4tdYrf8svo+BgUC46MRdg9ee2gegz3mpzZfD7i19eMMnJBgtumcFz3
1xNo+MvSd3/f2pQ4j1Zo8s8ND5JEFSaUcD1RrQZr4vpoVIkjZ7CuexfgfjfF0uxYJnFBSQt1kGZd
MHSlhes9T5/feiVxk4mDbvlFWV+Ps/SV40EJQGgZdkyNA/GXxkwQMp2RAdAiulR9SMvYcpjRqgyU
9FnkZZIOBxpHh6tLc49HJxZW9byiCisyxcWg1OgfBgc+EK78/gpDgBiaBZvtftNeX32RLthFiBDi
unXFWqpXcnswX7Sz1Km1MhidsoU4xGik12KrXmdnd89vBlpU2RrIrZVUKj//HYXzJcN8i1J40C46
CfCD4zmOMb0tfGMAxIgHtLxjkCryk8Rg4mL0oTHeKDrvUn+CpldJFfQueNcqvTYv54FJYuveUWfT
HC9WPulnecI6vwYtJasWSDCpYYYkujifMr/O50r7/ydZFEWXisguCSnNaLMwBm7+Td8/Qk2QB9aJ
BXqdyiM5vM9Oroc+SMBgiRhwOWO8xeqe9rQe0hKfh90OVCha2Tcn6Nm99ZfYsK9yJqRKE6tcNjsK
nI8WAD+qXNfIpDJF8LNQ0wBdt7YrJV4XZX1/NyER12cpo0dx3ROz4/YZBPI/HQjflFEqQcBloF4e
FpMIct38FBefhC+CPtDK9pp/DZGkPZ5l/mLYhgNHhXMK3FQCGN+Xf15HEVOXgZMf02Guid65C5H8
szxh8V/cQHAOVkvwLghmhxD1AWxSZ1CrfrEEL2oLzpKC2cETOqaZVo/O5NTEPRDfn4AqkldKyOYw
7G+PkA6L+hmrQwP9ckbTXEx183mT/cZx4K1JocxqlY8lLtiewJyHgXBW41xC7q2G5z/kGQ17BDPz
fk5/O37M/4uZwYTsCKp1PRHHIi0kG06bzv+qbhj5NAkQmELa8WKnYqGThI44QQ0SMvfOKomtYg1I
UHLlYXIoUav4ycCV6yAjG4YBUgVP0Cvze4tK0PwxNdHv3od/ldfAItSgv7zfVEbfFXQXUBt6PrVS
Rdp0UtcNG+5yKwqT7kQddNcxB1cIFRgwEYi0T/0//aYB9oLT5umW7VrGC1ehmO18L4EHJ+/Cm7yk
79FKi8zcjSwva6MC6+m4p6UkeVGD63Z7eXHdGkQRWepmuIE7Qou1wAE983GADJGQ467P6C2btard
vTMC23N89muAMnRuuUl7+NZe0CvXLe7+xKU5mHlY7uAtJ8xippCqLKXelNcJrU6IMGm3ayzM9Q/1
l2FacROWRzWN+0uGkoS2+GVoilGBtPD/AuAV0d2rkbp3qW10HxaU4pl8R3aFCzzyo1OWsIX+ypaS
q2jF8MUjvo62zRL/Mpm5d4Y12LnvknMHgnjID34CoMiaec2Z1cv6bXCd+FV1TNKR9y+Xp0igRGPO
0mCXFlS055bOI1bvmquX1edfZWNT9yERT9sNDJLgTw2qXF0oBqpo/HKcwc/cCpB/ISvzJ65/Nd7s
tJdcaNCRTL8XcDvVpC68d5bm6fPyoQzQKiDpXBGnz0kTliLZFKAE3vbBrs9aMiqQIxBin0ohaRtR
HOSX/npRgMgjM9rRio9EOg2EpF9jNmKw9VGBw/uLU2vV38JKZbEIcP2NT/HagwDxCzmQ3PmOl3/u
6+AvoOkNf+VyhjzCrH1I49zousF4L6B8qPGFViAMGOjqMiLf3eKy+KBvuks0/jcQ5d9IQr5aAAp6
GwXBkWbBFhSwHtxLznwoXaOFpbYjZYyiQtLNrXK8vgFyo+cPsPGKAku3nzIhJojyVViLRbtCHQAi
M8wBfvj6Bh6F6XVSQO/8d1PdsEyoPWy2avR51ERD30I/mNfr4uAy7WmVZM/Vk9T49ZYwIIQw5Ctk
/Srm2XJnTTxQCqwgbRsQaYGgW0JwTeMgKt5pgfHvTR17i39SOmW8+MJpYd3PGXhbDA9JME5HuFit
3Y9FmWBIrNcif3LSSvsulhNYJr/EiJoYHpuA4ndX2/BYGHlsKeHJviGJOm5EGsSxqjVxp9/e7Unf
FCp7PkrYrs6enuzxOoxZ3JrZPv0QXUWi2GDhsVc5362MG4taT17uhtGhilbSsfMxGk6dSH1tFO0u
WE8RyVeQE8qbXtJo9+YN5pLNAvIePHn4FBcbMXzhd5vX1QxaHNKpYXPsAJgJ/64cMzpXUfY69c6K
QU308rnE+Sn5MXrk/Q/gnI19PgUJn+8e1iZ+Uos1TF8aFW5rvQ4tBY7f47dglfPZT8DOSqvx26Jm
1FFGSsd0SC+Dmw+hqJYFLCC+jZeXgDafXGmG70/unf4uVj26bFLlHhTMeVbgQw0pnVBCTePVONdP
07gofAp5sRZe0+cA01JjGKlhHd1ZJx4dXwPaZmKE4tE4DvI92xEVPQ9DcV1IiEWqiRdk4pqBiBqc
P7iftBtzXN/rGiilItAk6RHTG3RQBr/ePw9djnh3gKdGEVeZ9/1qL2otSuwsBG1br/KdWPa1AgC1
evkLvLJyi7MEmPLpb0U8aORLzejUdVPD6BqWmCSpGmWCBh6nLSAu/cPAE7VB+B7MrWkvfPqYwru2
b7+LmED1o5Y/n6+0Sns1q2gEgPrfRQPuRbe0QUzgdyu3Hj4IJTXYMOFVpn/UZ9ab7lOsJIl9VgAI
G0mO9oEQwkkNNvCjgAnSb0BNn5A0NNlvbA8hY+xHEx7V3iYGNK3KcpEcmD+ajHmPBx9gOPl/cZb0
B7c0+CUPgpeRSurELMnsuITVEYIqsZrQ0g0WLgupwFO6d1zLfeELRNiK3k37mRzS7QaH4hkmCFO2
/cSKpWkVp5B/nQwscS2eyo9SNRtaQrMAUd+s02eyX5OJQxPVf7uTHbwNrbPyIORwpvZTp06JyX1D
i4gr6XpeYwEodn3nz4mt5JHrFkBsdyJFPEOua3DV/2CxIGt1m7el5g97olY35JWDYovgOAlgdMYp
04Dj/gQneEX+vWBKFcptIU282XJUXYXf2TXAd0r+3X3PzGl6KKW22c53ZQpGpPEqQDkXPce0F7oF
XjqDcvP9xOTGrYebVxMQfsoNPzmsCm7a0cn8ImJaEl4CLy1+e+70uDcrZdBeaG5anHdl5PkqRWuE
RIg4d0fNv8y4glgic3Bn7Rau3CzxC3+x3eyySop2ltWdehiv9sg66zrB9k5VODnoXsYkSGzOeVPc
1+KdIr1JxnvNLKoTt11Uqtg66fP0AHShctFZyCYZhwvdxfGTlxNuoDqH0mUOqkjFx0VY/lN33IsA
3rzmLpHCQPyUp6oNuVARCb+3fONqqrxboSlzJ3yfbR/EcEjzFt0R4r27juic8XDA5PTNPEn9sWGB
cQiy4w4t62iNbsa2BJTmrSvFRPB6UWRl9ffE93Iy+qaSN/f85sbxEqWMQSj75PZixPqsfKT/HDo0
ScWrje3DGhQqW+wxTNqiEhOVINp96ExYz/VLi+YtlgMQQ/5ls0REqci1rkbDIj8KzpOOvf+GBX+Y
eHF/Wo9s9etyn4X/3Qw0oCKcmveVGZH5KG6SMDnVNwcj6VhFmqXahUtmnvEFB0ocXC/0+tlyCu7u
dJtmHvyC0P79Ckb8l+xeHhzgS9sRD+qNg9/CLvZ3RqBVwESQvHHaC/YfzVxIYpEWMtBngDeqjJp6
Gm7PGU1+XhUFPPBAjJ0v9QnZaLBFNWc+hNqUf9Sl1wWFEfep66uuY+qkf0CH5qexP6Sisjvfe/L/
rDGWq2nuVHr+ic3ThfTEg0PLkWue7La3baIXd6zka6nHuIEVlM3zZMTga2WV7BGp1LYdoyFedHip
Q7Ecv+HZ3onGoCGG7N72LTIQlVvAu7mwml2gxru/9GcJHYNxerQRWZyM2Z6YixU4UaAhIq+F9ty1
xoJTLSDINTxyL5avoPyyMGOdQL3ZWu2QnY7xO+CIvMd8TtJ9qQT1nC2G56lHvEAJj+Vi5gvaRKeG
O8zm5f2Y2d6jP/ITuTUp6nlwWY4JI0Dlep7AaOJ9qhykcbeO1ky3GbNuAowb0+5mtZXiJwKZs2Og
o7mmfD0MC1Y8HpZ4FkuRK33JKK/8WJ+bKAHMwLJlOEj7ycuaLfcLfUvEcUXtsSnz1ESi1srRcORj
JiYs6f6xX4J34bxGzBE0U41jBWYfu+dEQOCMInK69lyGmAn5od6o07zJZ1y0UoPOcrael1C2989B
+txUf/2dWsPKeA/R1r1sS/OdwpXJawXE6V9X8aaoqtnsZJdhnXJwctTH+V7yn/ot6sCI4cbl2Ofx
4eQwUapnCdBqgENQr4TqXYGarLUgqZ4DnK5D4nvQ8fGwrrZGwzEccd0XIcB1RTyaxvPPZjLtzmBf
/8N9K1Q8Mg86dzyBoJM2lE0k+R23I9dpTrXMx6PvifEBmHFZln7tQsHJ2RBu5i3JFXA6oWt6xG1z
tgpthBAXX8LhbNJU0lhh37NjV1guupjUKO2BM0rBRnImQNnzt+rJorCeHNhn3Utun9XV2YjCLAYv
/nOQ974wIknAau3kDAMjkt/N8aIx/kBotHgTdPawGw8qmn6/fI22/066PJNEcqoFKvheNJPZrYy+
t9hVUcC+G7luuhjdReT5OvxcuLFqqeKWdltUa7wgwinvEiW0+QXm3hM6FCGlW0VWj2I6f6BDbXIR
LcXs5dbQ10MaWbY8DIZUd/FQv6j86FIhfYhNzRChCnzdEg92I/9FR7bm5j8QTHP19SoC/iKH1u+L
fIk7R3thWdhh0My2YYWiRLEVj4Noy+Q4gCanI2SUUrJFK/0gtoUAS2g8x/6trfiob+xLV2v4Udcm
JlnDBJNruta7WQVUwOx7/jHqtLqq1r1eq+79IgcfZQy5+a3eek6VaEaKyECGPiwmJM6fyIp2px5i
ZMqTN786UN/Mv5AttLb+UQh9UzMJ7ArEheJ0DED31x8nOkiDili6ntmV7vXXKBYfmqB09EfCGL3m
1T+9L4DgtjpTvcuPiabiWSS7HFXXl+y6smtOzZNYMWBqaKzr/FHFYj6KoiB2TPPdxFwc5hU+1vw9
Jvg0zA0+4ukN8sN7y/sLaSD4IqBYEk96IBS8OkQWFBdEUceXvGXjbeg2Rc4v1o1McIZRk9aZoeHE
TwznuCf5a/grKdC8oZjiV9Imn3KTppWqeYtUK4z4wjU3sAtT7tqLWVwT6EKd6b8mKHpZrKYP9rLh
FNzWqwW5pgFmEocGwYdfDnvgCCl8AIoHMvCzuwnZOX0bkrOlBz9KXKter3JFSWiTCJYozkh/2pN8
8XWlkw3Uc1Ia+vX9bs011Gvf3uF2gLV7lX8DL2A9qfwitV069czOi21n9rlSjC6JJve8HO2YID0C
1U0JGtw5Tl63iALqDjI/WkUqR9GhWJYv66Ecyu312oXFx/K9pBlw6rqJ8ujJw6vFn93+ruEdfA8X
cQ17bRRZcC/CH+6zGZDb4TGy0UMM/c1l2/YVDYgLtfnLBo0Z9vbb6RtHQl6HuCR3DAf6WXRaf0vL
HXS8Pfp4yLrq2c+FJYBfPU7INnfuyKlzDRGWWxYVDBfSbUG/8uIjMFOagxRUlIQUYA/TrbAaUwS8
9nZUoYJgDskkHp3ma4ba4OalRIeOq+UI8DkJmhlDqKx7UC+Gd01I/wURosO4Vk6ivjvl+6ww9nyX
mD4/uhITM3JrFsDohP6dOuJ38qD2fNVL9YJXymMh4SZC5oHAc+QaFD/9nlf5fy4r6pXq42NST6qE
tLrsq3PrtaynPKct3t84rxLNbZTKYa7kae4z3RvvBaZa3AJDVK2Jm8KTjWVYClNwKhelOCiMJgsW
6T1jzWf48FFG1zL9z0pLXEdSesWZMZCp4oydu/yHrp8UkAG7tPDJWznkW2Cljs7YfFB7uZBBB3lA
Mltgp8H+7ClGfXKKYYcyYBmlF8lskI6A9APyHVFy1rDRygKlCFcHNr5AYukimxAAWNarDHZl69f6
XxiOoqWRZFejzGp5itdIjOkF2FuhUqNj6cTNeAb7yACXARqE/rV1yZEt/jwa0SAyhxeP8xhUV85o
NHpMDifgEX3vi7sRe+jJRjQA0gBJrfAaFVJbiCgEGxzVRRt5iu2SFuLQe4os5MLhpcU6Vh2xz+fB
wAibhhI3qpDNNMxAE/utQbjYOLaiMHShO/RtHSUMxPxQXWtf2CeZ4GOcXnfBDKB8OE9UNHFrw0K7
NK0nAGAQZJ0c3+GobAhJpt1URnZUaM5FjDV7mPinrH/HuHbBfyZDxt6a2pjTToVkfW6BdwXUK7/3
j1VyVwmdpmqwqxnN9yzxeYmFJWlnlfOAbj/AHXp1DApdncWbl1CQ8jTm/BNoMXS07O0QNtf3Th7L
7SUmNZsd+QgvefZCa8mDbHn6McyGWn5Y0t6WJkKfd/ha6ufnbM78KEGG6P/TQT9CfejS+yzg7aXF
WdR9oZMa0nFezXeqxB/esr9zzhtYQE6ieIk0S1rc9CjgOuhqIFgUd1cF06FDy7EZ5MXAhwoFejdq
ub21dGnhNnA64F7s4qfwyaesrrklPuztNvWU/qqtx4FX4kvMM1DgJb825/1mt6WoKGz9A+V7+dVM
7l5QkcHGiZInrqY5GQ1wCjtvtGBhB2MDEtIvJQ0Fofbd96pdEmX58hnE8AxV9ae6IyLrKVPj3Swq
l9VT8ZvWZsg/7I9Fb5XveR0DjY7jdQFoROvvEFoNTYgD+OVVjPFXvGMYkXQekGm32JpjDicxocdT
wQO9ErWaDhJXWqs1LLSrFhOj6YwDouU1PKk98J/BUwQKBYpF1Tlx5u20MdMNbfwlkOHK8SmOUm9L
z6dQzLaG+tm0O1YhA698l/wYU2B3TJ106TBGPn69VjqshuituT9koFcDxFC+8qG8DHnZD5Sx37mX
SGdBnoLxgR1ACHkfWfWRc1FVZwZP6v/CfUeJEjhGfNIHNjYEdlLSoK4DZtyGdHYik95/4TVdqFem
KWdM0cJh92LJPaRs7d75itT2Dur5OU/xR3mq5MUGj8fptlQIqMUUvKQj5KzCHGPOwx/b4qsPqLzE
eUD66qHkKQ1MQa2fLpaWocM/oz2sYyy4f9A7slDMFwfGP6XosKDIDU/WRhzFZCaVQq9CpmrxKZ8z
X9IyEfjcxKMoCtNSir6M0VvASH/IfrBgwHTjDsoIWXe4PWmzxiz5n5O5KkHMLno278dsMs0oTdLH
mO9JE4HS3XE5yeV11iLN+2cCyq/ZwME5QFukURlhF+g4idcsRx2JJA9/FkFM+YGZ/Wnfh1VJFSlr
fKjBHXL5JYzfz9WDz6wSOXz79U1ujPG+Sq+OibZT2THTsBbP21Tld+zXXvLfYf/ncMesW/6D1dNd
UTM1Dya0pJve97zxO162HBCZ/go7uRiOJqRgn+TSX7171F5Pz42cC0yA3ZnLQrLaYIhwkqEtnONJ
xBYuFzb70CZ5+gIdF+TLU2GMQABdzGHPvogb12sAMJv9jP+ovwj28ZWQZ3y54gKcz5N01n2wbPIT
sH1S352XIIf6eFy9G7OEXdmANAkqugSI1IeXOv1IKo1nrIz4lMn2oEIFkrrbRMGYc7ojpZdSNWpa
lPv9aIui+XY0wAz1GpNfqBvDZSZwj+zDgcG8iOSsRr8J4hhQPuG54X5hIJ+Tr9BH/p7qKbmTvfiI
C7ByGpEoXEAcsbQQEdarvHvVJPcy0oP7mkCH3gF8TUSrzZgB/pN5Ftpx066fA9I3v8or4XfTQZHP
TERpNtyaPfVaSUPcZg33AFPcpJdO6snankyuO/osnMI7D8LOmpd6bzNPtqqbMxUCzMDQJ9G3jL+f
Tce+wpM1zGJDr3gROfgxi8knXNq2jE18HaFqVU9FSg8aPj6x5ldbIyKXgxygFAg+y47tsszFSqQv
ijDQDdzvAQDv4M/LtcLlAU9ZiG20C0Scns6qslf5OnsPb9uUqc4gMXuEUFXxTjS3e80dq8Ixurcw
RaYx4HwbxSu0COgR9fObVD6kHdR8uZ9TPSQVr60BHSDk6MRqU11/63RZV2rxYy9nGY643Dn+tZz7
XZU/o5gKtdttuMrzNDcH9Xfv7gxx+CRWHtqreZ1fv63buGgt+N5VjnwPzUrchUwra+IRaDLbcu1s
zHw8WFj+YPpqP4e5CFVV7J9dkPiTkO+K+TRRaB8+aBtOsQHtof8E23k4+Ig7E8k9VeKC2ASI+/MH
sDpIJ7F7TbKno+IcRgfwGkpYHBpdEXUmylDakKy0IrQCNH7Ub5rwgJOJplCVoS9bkypzcon8O33J
KUZnEYYJ33OM/zOuyvsBbYrrKppbOCQW33YxG2owyMLUlPTe7o2JIKIVf5LxhEgozWYMWmJ2Yr8J
skr1tlqovJXmWwdLdiRU6KFs++2RXyIFtNXeoIK7fYSjOYO9VbQ83dh3vt3oaOgxCG9FzjJEpG4E
A9WYFgfRjntPndhFjkzoPMeniYu3dlbrQHWGfR53wkEAcOXhSWjTHF479lIe77z8IjROvHKc8eDj
t4Y/haArohh8Kfoaz9uzbVc9y8sx9odXQeLhyEC97MU6V71wNTjIj/QTZlmb4xhjrY8tFWzfbjwU
H9YxGMU6qdEQOH2Wacym/RtGvPp3tCPiBENzs1HD7UHBfpH2EBzB7g/81HZp7bo+gQpGWkydSkQM
ruA/wcfd6Rxh2gZ6yFHO6wTVxXfNgII5Qknn1uf1DlM2tRna+pFKvUnNjlgn8Ko53yVZhcwMZRQQ
32scdiFHRhts2Io/dq3DApVbmbjs5w8h/KiCselDr93+0SfZKT+kujet1MNkdMrjFk9fBsThLhv+
K2By53OTkj4ge8ebcRUDZeZZz8LVrZxs6rkyvI+sRMIJXKu79Wv9F2qoWJIHQ+Di896wpFuIigpi
evXSeKMtXB2p/uQSidkjTkxi1t3WJZN/qe6VdzKaIlCHHxYdVqrLe3BlmTEP8O5c1wyONUlcnkuZ
BSr/KFbXb6f3jnqSyu8ZC0zaBx3/BQZ3nl+vZYtNW9QqKkuncaqgBuyEfDbNsJgS6Uw0hcwxqXWj
/Qhuv7Bmk9xP9gtNONIMFik00HbIwxYlquxJ22TyhLybyOWvRfuhOaxenLPm6tv9Ynw5DH2vUU+m
IYZ4zIuY1aS66TacYSCbfFZ/xjdAC4MN6+nNZZic4OLSywkt0seqp7uQZEL2cLmBtwctarfXeMFE
Q1pUHSmxl7bgrJkVazFFROhlff4j3A8TvhInrf7kDITzBlMzebdcM54roLsV3X6Csy8ZDWABOZzO
bHRjGFqF6mq0LH0/+uAOHSxIE4UYZ3LfbTalaP/4AhD8kcEdNhnJe80hbyZVJTg3olZSvTJAugWd
JaaPByWgvZptZJd5q3H09yy6i4o3yg/GwkaX4OGjEZ9Dpsixh1LR7+Kg9Jk/qyQyO6Id5zh20vHI
v3klMu7YGJ2ttp3m3XwFkK9Iyb7RwXs5MaQaRVwfjxXjxcjwzlZTuDsDBZFjPOehsiFTYYtrgkhm
qCTC3cguF86u2SfyJvxU7W3jDeVAtVo4YyUMHjSapPXZIZUrejhkczCu1h4SQFgbdmVcbrn84et/
LKzjUBHtEjsW+0RgeZVHz4LkaromFjL6R6uhh0U+mGjTtXpFEfycMQfaHUC5qJ/JsS3mM05PW/AR
7NEUUm6otraE2fKYm+zDEd8Eus8kt4yL/k6BT8aLsC45fmjns0vP8m8VZrPn3Y1nsiTR3PEUvkpx
Di+xBnwRdnXBbRmEDcpzM6GNXhy7CWwYqqC6U1PHIMSfxs7AEh3tVda/uAcAdC7S7+bXdEgOPCdL
8n2LFbg5hHfNW4wlR/WCF9fyODBK8LwFyw/nDk+t7TRaKluWiAY/RhiV66geuB585cHlvAAdJ8aZ
V+oH3vNVqk99sWXuleNPeQQ1o/w8pu6s9I6GewPkYUcrTL8w74CySj4d00TZDo1+0+MC/oz7XhCL
Sq7TujCJUN+Ld3y/dh70m+oZlwpoOwz3BX+m85cyfvZMxAZ2lzaS9sI3miyL77Z1DmXuOUOiSKB4
dJm97n3jNYOggYrrcRQQL1IVxyl7SW+Qp/77Bek1RtDbKk5jwD0IIYMCawU6mjkr3bxUiuTMMBTg
uWwlPNP8OrVUS60VzkQACaP3qRXWZSPKsbexsuV6B+nA2rcyjN2NZ0UCU1Vk9lLkEaDRoMhaLzQo
vOXvAIkPzCu+SDeSqwei7w1P6buzB/er4NIx/JyY0P4FN4vZeXaLUFNFagXseY01sKpVVya2JWDO
oENV81IfxsreC3QG5cEQJMHLvZIFEWa3rI+f4hH6+VUF6OuUV2DydZlP2mpkGDJe71fYaEsrHuwu
1A0Tt5fiCg6IDZKKTrtb7FzRouvpXYANylBxqNDnLiB3X5WW5L6pwKdTemPdTa8oGGF1y3peRbdt
t+zkycVrnIpJrs+QlsIFqPFncJH6OQJaakdavVSmBhOKgtDWoXPQAMHTJLaVDJuT8qKeBdweFCD2
89fH/m8E4sf7H0/Q5mR2PkeQlGxpzFU+oWxHc09gfW87GEBUj3TrCoGQCWudwipBxnzWFNuFZo/Y
0fBnI+ant8OOj47HlhNaK31hp/vt3BZkymzyRZTs7/CS0tWR8aTv7HroSzxI9+C86eTBWHGoT2Eo
pnEMA7i9I7QTNQoedRYXhICFzpYnqh8RU53xnDpgkwiVfGBjNuBrAywsn9gKzfFH5TTTCcF51/Sj
X1l8ABfWvw8TlOPsIWvWPvs1o+5oYa+Qbn3A7ZiHEdjXSImvVMBjvWq2HYrY+qFwTnPWcKrHOzt4
zjsAI9BtB65vLh3fay7SJ7LeLZ9ml+wfA1NTj64aKBXOqnyVvedbr8h4fNMj8q2BSk39B1/15dnY
sktwQnnVkcCOyghp6pJt8pwMyXc/0Rs1QPgSFsZD6YWTor1TbJusIk05Zi864oANiiQYhprHWtrj
Y0hLdyRw5tF66zxLNhsT32lDRzz9ERq6OdH7BHHvK3fb2KHqDEje2oM+B6TApg2+CQ6YKmYtL3IY
VkEpXwDQiuwg6gIZkfwH5NdgXXFYUU+oHz6BJvQK4nAHAXAmzyTmZvmLB+ySs17X8NICZdfmFh4a
O6kvAGRuZa6JCoUcs291uNjMbjCRUrDoiKmc9XFobNZ+MLYYF2bZIg7+Wc5BUADtxCcJu8X2GpuK
S8JCVsio0LY0RKYHfd+JuYMSXFh08wsd6BYXblUj5SzTCGAe2RL4mh2Kr5BJMyUxro9IiodGKrS7
VJsjs4IHNtzMspduEdGd1jciJHuu/5mr7LP1AcLdlkS7KBYrkxqgMePoU2M/oLWsGqNZcigSNM/T
tslnJ0UGHE6K7NL+SA7wUNTstza8m8jbEpLnxWbjKnlOYtZ/63MMpQH2DDoMCx5pRMBcKJHpzdEI
VlAVX3wuXA7hOWQFkIO0EnWGTwIz/K3kz5r8sXjRal9x4+AYLm6b82TryVNClQbQhG8BVV0K4RVQ
hqgtkypk9iQtV5+sT479isxqNP2lXNrmLdu4e9OQkmaJDv5QgbmYnPgW4QMEB1rjN03dZayD0rao
+YQBr6OQHS7SB+ialFSduBS6RjLmGnZsbQE6BZt3nTBBI04OLtcpAiZCKIkO6G/5t/8QO/SHnajv
5DXBJvg4YxiAg3JpjRBsAO3SVsAPMebELXY+JAb9CQWUVCrBP9HjapooGum4HkIzdcOfBasdFDwg
A3DkzCUi938yQ1fkOYFEiw78YEwTUW1a/xjp68FPZ4m5vhI3bG3AuuyU6XjskK65KHHJ3Qq4Lmm0
AmyczJxkfen4Bs0ScuhyKfi/MXPhR+2mzyOMHuxcYopC9/3BBEcCWrLo7b8amomLz+Ta2ElgsKQC
U1Gvd0h1jcqGOFjX7ra1ZvworlXLzWyoxHqm09sCFkE1+wZVgYRZEDhYLTStabsDWsMiLhlWTuPT
J5lA3HTepoNxtw3yPMc8o2m+7cDnY261bAbag/959N6vH0kRoTzSliA/glRutwHH5oJF+RuP3tkU
xy/mv+LyVxfHiuUC96u9Dq4ge1Z+V1kT8bwKUaOovKrqXgXn8FXSiNknwGtmkxeRWkwFobIIWhhm
5xbXrwCxJ7/2pvaYaF+m/ki5EwERoqg9HjYQJ9G2Axwt3uSzq7lSit1bVbiCVbYiO4/jTQy+PoHB
N8ie3+Gnxg2LyfWUIm7+evAGZXte/dKWu7nSC9U3qo6phF2KrVz8u1ZV2p1HTtVWYVNd9eXCRZtZ
1LAe0zbC8DXWXCswWOAjNOHhs4apbb9JPbTKaevngZXRHUEtwT5IiL0agDwOx3fIEAVsstEJKLpO
asNxanEQm9um8kuGyA/dJeUq9sdeN76pYXgd3U15OOjmZHGFmA2WTRO/osOZbdJJtkNsldOcoYJ8
IFqSmIvXkWHM1+DEKUrUZFiOv9MTWANUG9Ei28ZSOcoL6s+Y0fNILNWyFmMx+q3g4ucGAq7QPsJ1
wDp3TcmT6M2x32Pd+mTeo/c2Iw6kJUhcQOFNrg2gKV5+6DK1IDEIZFM3A5+73DUCvx3YDz4D0hXd
nNRpw0+dCOo+mfE8d3geKaqy3b+k3cGQTTHiP21nqCm7zWLP8daIGA0Eurv9BbwE7bxn/f5p80+G
M9YOW9KCYKsJYI1mgtD1SP2gBeb5TiGUVx8Q1oRktvqAV2/bC0W/YKPxr+zg3KdKm1+UIXaT4LhK
AcmdJLUBxCTJJbgAbhTMDvez3VLLzGQAm1ia+g63cmU0IvrNrx/OJuybRxKdYm6yywwPsvF5noC/
Qoo0oIrm2YP9uFUJkphVUnB6H5F3cfJYsNEkRAiJab1F2nZ4BWDPD2XTiBc3vkE+pLy1p+iK7vFL
LJ+pCY8x2mr6418j+9fQtecpbepQ65A15ZHpEiDFOtP5zhxTJXA84fMt/gU+geyM7ADMRMwVtZFo
fp8h57t8cDQmSn0/P1SAhim3y1P9ERdqOv3+BC/lNQFjb8M4ZbnvXFb37Y2v+XvezRMX83hzPRuG
xz8tOnRIHG0pYXZCckizPM7hAUBPSgukNMx0LYnehgkGg7B2P3EoUidWgFobnpXpftJ790qRAfU8
5pazNa7MqnQuKYjHefhPIA+eBThd1ky+vfBcq0L+olTubFGGwEc4+5Q9PfbCUK67Me/Ea9twNbbJ
ssu2DmYQtK0eUlB2jENpUytTpuno3v3l+pAbYE33A2YadvPY5/h2yU9ErY2R1KYFqvWEXwLUyzcL
beUPiWqqjGJtCZbuk3k31DRscihwJ3sUyiby/puc6MyYofbqUhiUdmFAOazZJ/+kzyeOL/o++3Df
BEjVmZcb2fapVR6gFp1uWTYBfT2cXuXBQUCVbMrDtaRO4YFZ3NLs+kXOSgyjCXDMAO6nooOVJUdt
pChlep1eRYL96gJrqyOSiV246OX153fsAlLdp7Z1EGREx7zxRXFBfxrb+7tIrixmb2/+glZ3HP3K
Y3PtsUZBF56TkVHc51uq6Rhw7kQOICTr3hMEngKCysCuCIXauRyy1PfczN/hgG9xwWG48Omzzdo1
omHYLCmjrocm+5QLPnj54pJxPEhnVdtwnq4HLmuxThVFvh4N1zJWD90sM2dmn4RCaJsLbO75Pjdw
FfH0f5n5zsPsphInyMe8iaRB0qq1rg04zxTrWjDcwIHR1SIir/s9X3gYif/4R6qSEpPmk3MORLAB
tUnjJZlZYZGvGpJSkag5YuRDQY2UtqVzjRp58SdrRKmXMQksbUMy69J8kCFyxUa8SktLfN42Euuq
Podxzf69RcPLWAexxFA35FQ+JleqSJoufRwfl6cv4u5iXABRVxiDuyQFHLFdCyRUjl4AD8/3/swU
cnIpWERTjKqAgbKtoQIMo6AEiNaL74YGrRUTmJ6WlRPh9+gZsItUf8/76gqMMJbHSDV8n57raT2l
PqWjT5IIDckG1t//s9yaGONgp2bwQ5x83AV8G0pw2kohufjYuq2E5SEFzlF8TIlC7skMzi5t+jPp
krJJsfXTc09sgUpMeQeqRDTRTQ8wPjcoQL5vGOnyxXyq9f7rYZrVaEbcqDe3QoyxnJyAvAGBtj5X
d/jMJeUsxmerJnZ7WDShtm8tktYuLt6Jaa0Xysmtf85g3ZSxZjXobDRk0VeF0zvSp5mg5BqKLAMb
QFnPxw2pMf4Ikw9sp32sZXO/x4Ykc+n4HYLOuD2sxux8+FeeA7mh/5k5zNcuFfJa1MqgPK16EEEQ
goOtL4yz1KhosZLCeSRPMW9Lxm+B1H46nVnnGj1j1tJswEQ/mgzj81yEiYyIInWVJH308lCTn7Ea
rlL5L9E3LSxYaVsYtRik9c5pt2+G1TvUImRlj54jn/KKdSLPmKk1HQjjo8jHXC///S9FDesrky+P
7RoIsgdd9TtYy/c0/mj7zOqw3mmtxGt3XMCikVG8XGAsGcAtERVdeBsVhH7II7V2VUsUbO22m6qG
5qqk/SBrH8Q/Q8t3nReXXzfb5JZf+TIsAFFJ/kGxmWV1GFGz2o3kY+jS6PmX1JqOUFJ5/js7YChX
g/lE8zc13lLfHUqgJQPa6xtcL7hsuDE6kzm342KazUXzx34PQEzkymWt9erqO8zRuoQuCBMNGBjk
TKXHP8Mo6oGGR0VMkAs0bUNRBVGNfS80hdSpLChyGkrDOAFG970UXGE38suOB2p3uF1iC4tzry5S
fISD06eFRqJY7Z7ZI2pAVAZ90ozmWM2yt3hFuHUJbRk7ZC5fqAvV16KvpBfOe+GnxxQj1VWDGOt/
ziCyemi4faBj2BNAZbkaps5MnH6YWN5eAz/1fZoMZld+wY38WWRsSYPHWSg5l1OSTNcvwCtkuzT3
yhQw26tn+3/tQbri150VlQ2Sg+PmSUtyqlc081PulmJfTseFJisPbVh1pyQYlxHW4KnUADUqBCO1
YPC+Namqe0SB0IxAIE2n4+qWGbiAN3+Otsx/YeP91XBJnp039v9bsSHU4hkOq0xSo9yUf6XOPlOr
Z+bRCbobwhESKCxn6jV6qULJWw/dsCl/wqksjm+kRbQR5pHtFHNOyc77AAql8QqvI7sgkXOwNHrA
IM8ubzkYv8cvc6Iv+cq9LpZOdORQn4B+3FA52EqLnAhT6I/cR1cSafRhH9FGt/eHLfIAhFfoHiUG
jxmXDUOyRHvqs+T8DEPOW/PeLx1psWBP1lL+09aL04PpmDOjGOrGs5GGnZ55IpN+IvL5l8xivIQd
8qOYc7p0l5Tkkk6fmkSRiyvIpzRnHHEQI3YZ8Rl6zNObUhanmyO4oHTeD1TDQp6ILKi7JevWWb5r
BwhdpjydKEulhGIM78wKcAe1RPsFM2pAGWqvQIRbAqYvy7N+5ykOFXSMUr9mofcgYl+7HQGmkJoW
WY/JG0Ywa3nM4RqbegdPoDaM/GLHWlQPnvE9P8HuHCyDz4gfeEzv4mYSZG04hvqep9ynAA6vu6WF
3MSSDQeTy1305uGqwc/aPSZ2jSg81q+FHbskxSjerFRfo8z9+x1IPisBbFyk1Aiue6TNGmsd/Odx
LJaYWu0wtLzu7Pm18iRsad1A2NHfSw1IxUczVgmGfnGwD1U/OiBsbdgGravIxwUSYMiLG60CZ2lr
kzpVSgJY/jB0dW5gXlSPozplUubePyhmALMiq6CXT+KfstGtbRK86S5dI9Mahw+eHRXqciBEwhID
vbBGitMb6krBLV7ktzjGcEnk0k0FZ0my7uGmba3fZCJ1LkHPcxug9rLiqsMpF3xy2sY78tnBL6V2
3tULjRIQWaA3PGDThq8xbPu2Fr8zHSZUKCeRzkn0dEPqoklYJyiqTfmu98ySmjUFGf7qCKCJBIWx
l5XHjlWGACzwMcGrwaCuP3YINZPWeT0+9lLnn7GS8HfEFUX31rUW5EysBWHBKBdV6J4FSUMSuNOU
0uPSe3z+GwGtZYwlVvsGaOPJUBrMcl2SRxDSisexmjyLx3JeVoAIbUIqpeSQXwhcOiz4O8XzWtFC
GVJAc8RBfeh95zsclu/lKStJ0BkK1TCKgBzfZnM0Vm/s+Jz//vkV8CbRhou1PMSSX0aZ5iF2bO8X
hvBHJwl82YUmd8bJsrj+cAeE1rykeUBENkcF04Fg841tFKop9lK0MH0KSZBOOzZ2M7L+ESGTu7L0
vgtFIDiYaf+nOPyHNpbrbuc7NSoqO3PsgVrTB8lF/qUm/nbzpvbaKw1J7m8PNecwzXnqpLkWcTiV
Tg6E6aF7Hj3BCH5YVIxcMDQB+d2Tfch7oB4LI0xUVSQnc2wiYqKsMS6+yhH0fj3Er+DxA1G2o9Bs
eqetn98wkNwlbAayy+SxaRGLyTo/kbSKpI+YKfvaFWPzV/LH8yuxDq2Kj7/VktMObqNw4nVV8pdi
QakgNH/fyrM0ajodAOH/l+bT9hy/TSf7KtxBiIElfkg93A4nlg3FVM4BMneuGvfDskaiipgxmvW2
7TsZezybqQQSsSTqEclMB9mu1Y5rf5DZwYUiwGi8wGy38L/AtrrmmIX7fQDHm2zqPn/gNsabwGZU
xinUo8pujtz/WXW0VmDXhb5QmSl07GebTKGrbef4kHiXdfhkD38MBjBtA6WmFAK/eSXRzPcBRvGg
OOqa+iQ7YjiHxmUx6ljSmOyxhmwgSMIHCOulWEHWb8Ymv7tH4GhzUW9VXXSUybADV7qRVJDFulT4
WgDRpMjTXakfwu0UPHCIzw9leKIkXSNtWq7Bk+fQgYLZ5eXpxpxQ/F1pDI4hmUzxpjVuuGXM1dib
kI0uUq9H7zSw69lJVQqJ5vsqDFPo5tlB+yW2pIvui/Q7d9LRj041QU9J5Cqpt6jnThhJu4PPt0Ia
sP5/iI0/tgPmnfqErs3RvlRtO09Q3bw4fHmUxT9xDZnfF0fGAd/k/g9AnVWZxsEyreC/oMzJJXih
wzsnDX04UbAgHMhs7jjiM41KoAeX/uf0b3A2gxgj3iSMrzgz/tVVvWUyMGP58lbmv6KMg71gO985
dc1JPFiL1EH7phm1FlwWGFYv5GBm98gsrPpmyC2eq0TA2MRQzxgra4TQqAUXFricutaNvnQVSc1k
/JfssnwnwQRub768LieP5qhX6QM/euCrsG3wMH8IaGTzNPPFPHej9R4SxPRrRjEpy/2+r9ZRoKUj
+354Xx0dKlTPR5jgped9jTixE6lPAA3+ue8Pp+N58P6xnBFkf30dwqxJFJqOp0919NpjbZnCsrOW
sHv18GizeRbM8RK7R7T2csoaV3vBU6oUCKHZF9uvI+bRQ70hqutOramW7JHOFATNsdIwpyfo90HZ
lfsLLnAQHnjRq51LBrjIwU7YjcPq+x4xWw6Gu82jc4i71q85ehSAgNTI1V9OcJjXv0V8xoLnDGbX
d6gBi3DXMT0dLrGGtWJufiuIpP1MMMUe2UsQEJ41L36loHQUyynQgOJR494EU2H2zm1eVrl+DW7O
AXypgL4zDV7bI4gS8w0rVF61l46Im7UHuGBSN/ca26YbVsswbdkB7EePyUQ1mHyict2gGrA9s0f9
UD4kQJOtqhkz4otrnX3gqraX70dHxi9PB/elfOBDIyjhHHqM8qkdKgYbcTAU3fFO7k621dlaRusa
FRrKW/EMD2qTm1TdRLF8vuJcwpM8rsCFa/ckuogj9oOkvMZhIE8QYjErzDscHjXy55NqJ+r6qd33
mt7jG8voBB/UTBlfNxegNTeuv9xpoSYM3BA9S61UkkKAdCWgpehyXY+AvqkVXguSB+kWG/02rej/
xm0IZKvERhEzza5QAZH4GndZ4Po2u9X6HNmb5MIokdb2UAOT5m1En9Ghu655s8raL4RbbePl4CLg
Fw+fInSk1fVsJup/tSLtA3pzvSpgqlzTPJe+g+4TiqmlGIkJyV07AJWhyhDdJtjxKSPsnQaE/h++
LSFgqtY2lWRa40Z3j4Ean0fzVrHojkMR7jFglBfG2urcguDpz1AY1LHymETacCbQuiO9SRyHJMoq
AFaeBBhM7zoamfGfDHWaDc0S0sSk4EL75uYK6VXjlfcrYfUhw6wIrRaCP4XoG/b3pEpeyWG/VTft
vXJA5tD+fBLUO4qAvUKlOt2LJLhLjPzRdPa8NnbEt6JnJCu0M57INvutgXJN0gTR5tMtV45XjXKb
wo/FqG2Gm1oSFtnovVaVh+Ok+Lc11nkvq9/diL8oUOuIKDPV+vuZ5jotsD1z9wmgrTnA07pOjMln
CI7XQff13GEKPyYSVmv7w6fFN55zdWbNKZNZXFV06DpS7Rfqeb66snLqilSlAOdaYwoMJJDTraTW
KbDmbhGsGvd7HJwCr1x8Co3iX5rcLC3KJqyqC7PaHakdFhm3dZJ1tJ3BXzuNcjZa5L7+1/7iEqMm
KnhMs/Nde7DkiQmBNsRXCTo3TY0R+coAJtNU8m7c/QYEx/VpvIpSqEyBmNTnAxtz47OCYMN3Su8+
uorJNF2EgTP8nlVIhPwX7Ebmzumsx+8qVgf/3DzbeRiIKwcn/BWWolkVWm6zU/IDpvwsfJqPJXYN
4v5+BYj1myB/ZIgW68Wt9v8NXxK+1dipUhmlDWEm4puSzqWEBagAtRCQsHQD51125SO5Z2rrrNZH
RwN27mNmB6Y85NtkZKO0jUS7XW6DkR+AmlmVqDiZJk2yb/yNcnrhILFaqXQ1h7QNsEwQrSe8Gdcv
6bme1yQdteaU68Mdf744284efwLnBsJ4LjhriQCq+wzevwR7ZZzeRfMKlsxugZcnDNJCFIF4AdoW
81352Na7qLLxiKoShmHfdHA/U3khdCZXIYpTzBG4QtszpMGkkUGEEjBEAMWyzi1fbU3T0g1MUBRd
B1qMHAqWNgSQqtErGXGG5Qj3OZejDF5emPIfmVQknx16tVSVEPra5C/iMhfQHcus+EHum2ivHn8i
sIQBGRTA7asmYvnxFOqPMaovQwXsKlHSfoT6nJp9BUkesthr6MPTCWmuYBl+RedRcrDrWKoXo3py
8Ao7Wby82BWewdH8pTVYILVOdlajNhMbn8r8LtUcijpU7fhIZ3t+OfvFU8dvLpzo7eLGWYijY+Iz
0FK7L/stE5+mt8aYGA0kw65NUt6GlQVlT/qlD1oXzPOr9ZbtP2dflQ1/cVB1oC8trb9aev/rdbDD
XzPtu9CZiqFuk6nQIXwf5eiOc5YdN+/cvhKFJ+CgvF32DeKhywOpQdjgzRWtkrtpjypNQJ4jmxJF
vMfa8K9qTvCyhZTTYniozaXfD2JFdXPGw/QyqGiySv8+RTeMuTbrGtQKomIhkTtyxZ9kslyPpXV0
s/OWDngz9mrICdOE5DcBfvM5cneGdWyu/ZHu1XkCj6UayPSVOpzP/3G352H5Z/uBfUfjHoYUcAbP
fwuzM493PAnsvFnX5e2a04whNE1ZG1BYDVG5W9mEMpF7ioY4dzhrMwGtxafx5zuusA4t9whDvKVy
Amwhj8k1ZFM6y02l6b+wgiupxAxlrJZcYHFsc60BjhUICmXfsuhA/XzSjz1yAqIIW2Q9h0GxWB0a
QTcuF5GrzUa18TjgrWW/7Mzk0NJ32B5neK0nBz69RvCqLRbwd+pKzGMlYHDqJHF5TNdqID9xSAft
2sGBJgsaf9yG+BnyScqf7bhnlqm96jrAsd83UlmttQET83lnHWbtF+sfX+zqDRjBqdHI1mHUnLQu
sj0cuimWoj6HAOh5NKdX6nVcI169N9NBZXgYFUP1EPdzaVTv/0nGganr1GxoCPnAeRy6nI0XZ8xl
8vDe9cmwO71tMATEQdvvEqn4Nq1RvBwvWl4cei2+v0t7gHMviT8PAAFR34PZfVoTESYhwczAACKN
drer2mgQMR7hTzsv4iJANWjx4qivEhdcZUrtvK7tUKMC0ZQg5MuX7GRNWxaFpoqwS6fYXHrYSl1H
n0wmdP2QXY/68p2Kia2clnGnho8MCnvrzODwrhbKr6inDsx4CYdUCGxWvhuMLO2yiKJTOGfNRX+0
hNBRyMrh2e3YIwCH9r131IFsCUfBX/gTfLNqs+jEpH3EsDhC3x7N7o2hWt50F/SWld171HqxMm+I
shpSLC4jpg9qqziwlbOkcI0pPLrBvoIzXXSRl/mcKAhUh47y28ocpA0L12gw4d7bCvKo4kwK7+fS
tBKNqBRYm9Klwn1GDTagR5NDUmzfnGmSHUU8YI6PeFiiwAMeGHI6j43fEhNUmLPQ4PQs3xcMKrDG
RkSgjei/G3WDUnuCobm0t7uxlOaujRT/TUgopSwIhs2jsjCH+XieSAHBAA0sIXRCOhu0CxFmMi8q
CjWRxmWiuhIVfiseQNzgh8fovyiM0iUDLOw+ka6cjNyj9Kxlhc55+fbavAxS2osRkuUmmiIF3O10
V9msIKqQtSs0JpYB+Gus/iCo50jaUYEuzwb1Cp70mXJa+DbHx5jgW69ounDYXvm5MjV624IX/ja5
r9s/9vPL46aYXNo5akbt1aWRMLrlF1uGjBj4Olt+7gBUYqh5g7YX1NwmQl8YigDx2PSuwGNfnI9H
2hhb4PR2aMAjv0xL3GxX9xSpO7QaXS+AuBX9ekhPiya0xh+cozYolOyo+IbK9ppLn4DdjE+x7jeJ
TmgsVl1MlmyMv/pOft2HEM+yFZFpjMjcPv3+cHBlEhm1moTPQm1wBNRV5Y/BjL1tnC/SOcL/d/kn
oW5M0U/PqdWJBLsHmIBDr1XixFYquK9DOpSXOCZLTFB2hnDtQ4886k5r5Ks5IICmhun4kgwWXlxa
HjsAclZ00BCSqPXlUBwXbYC96DvkZYU0EWFNxyikVCdCW2vfI+OWPEkG4lCsvhDp15OAe6wuxlJi
bM0kMqpzC7qV7inXysVgvoH73nHDR9xMJyUc6c0D2e6iN/LqpGrOVGYKzwBwJwEfRqPtBKikyiCg
HfX/tA60/2kC5sBkmyvb8zHnxvG5mDnYfwDLO3vjxunr25kt+G6xRrFcqocb3z2woleF1QLJRouj
V1TLUFGjgYxcDoBBqfk0kWjGso25lLfCFZa564cTWFKPozoo3oAUHdq0UwfMV5ZgAQJqaUl3ZWhB
L8XJd4i+seoNWrFf+7jyBDlyEzoHAZtWMB5GR6gZ6uWUVcg3HbuS5zJpPYdbpSdOCpBNAocfT13H
lYQzTva23D2CehJOReSXJMVNdOUWcLAC/P1Azdt0DQ3kAOHlG3laPY2sOydWpDapdLW5565rrNav
zyDlQYhE/koGrez3QcTnECFfhy230vuZmVGL2XtuWFmg6bzshhqvcf8H/+Y5xtkj/XmGUDBA+pEk
hTgFlal6k/o3lqgn38FM1axeUJFWzcHixPdqwJCyLAnHuNg8KJlI8VeizXTMN6LAxH02MhhaeyAy
rUr/LI2fgu5cABWOA8PkzpK3Kt6aJ4KPeNKmI7dVhel4q4rG/9U98l8+nFj3obAf7urS0va9Hn+n
0R8eCoSlRvu/2Q1AyWGcNcmGkXv5/CJ1BU+MBSqzjwbDy+RPOdVg9IocIFPo8lx1eq6pPT4yjHqC
pHpn5PrJuysDw8TkUXcv7GnvrgZ1uMSTtzBqem4s4/HVU5Y59n980Bw7FKEWGKAahgmMnRRYaAOd
Q8UFh2+9sIXvcbslKnSdtbBjCgRonud8o/5WuPo6Wwltfcsrawh/JWF2LCQxUA6ViXEaV2CBzWcz
NnBHuDSTA4FkfALSRMUAhaMyFl1q198iDkjvkTDWedhwTYhZ86azzus0qepA143CbvnTxapx7hJi
uGRpyxtyuOhZL+LWhxACoHNrp8QI+4vbdy7OO6dXBYBqkDsUR1n/IYJ0Rf40zFCMyM+NFFd4GsOn
Z91lrBVJkWWnzQk8C/P4hl0rQjkUfGaUFmL8xIsuiVqWLTnbFYifysARAQTTbTSdSk38OcwZohD8
l76FQzS8BteVAV0lJy5gmAOL9GquBeH4ysdtOoNYq5psbukv4MoE2PrZFzpFoHccSrykR+HCwIGx
ICUJYa+mm+ZZLqdYx+LcHAN6Ojl0i11dQxxTPQk2zbRUwi3SYWZ42K3UP6rT7AnXceuYWvkALKfc
/9O725DDEz0d/fq8++q7ZJsi+Qu3xklgvtY4+gEiyJjWhqBe+XnoefT4dWbyZY8UPO+EHmxBYUFz
UTjDmi4jJx0gtm4nXk3Jz932BtlDFh7iBdELASvsy6cBoYXegSLB0H2mYKeJmZNpD1YWvQ3iJqpU
ZKnP9Xf7uMkpPd1qQTP3Y+MFQQORL3kWUg08cxTmYUpWb4ypaLOkadFJ13/5yzgsodplmC24ZkYa
iHI2Jw3KXgIoaWTJYBPv6yFfW8QwsyOCr27wJQ0zag8LHNddLt/vi1ezmPga/UypnE97E6hNk/sc
GLvM8w/tDs8Anp06BaNvlgxmFav4fDqBd5E6/C8/pjw7tv4H3+znl25mkMUM/4kW9TVal84WDBBj
hl403fJnwdmILLHfeIwS8KYY4WSpu4/xCb0Y3tb4VXFAMV30dXXrZhsgERkVge2QAWTxtNIRkpgf
o061WTtzge8sNPKTxJOVSxgxye2ZOr8T02T3n6Kv5TACFxpqf8ncA+mLGu6c92SndGYgm1EQdBo/
LNN3wQyZGq+sYzGSd2TpVmD/XlTACno9IE0NVnRypiE0OfFocCAwVE/VUiJQENrqkGa/5grTRHJN
F82nN3QVU4EZWmMyO82OLLEFHFI/Gt4ZtfmJWb13brIiqqqF9Nj3rmc9mHsx0fiJno34H4b4dAZY
iHTtaOPTQzf4oKQ7HUIdFszrl621LU0q9h3iyPs0qQH5zNLTFJmlo2P8ulxdygk3AoNID6nrbOUJ
pg/q2Hq1B3jSgpCFHcEnnH8NaqC7xAv71EhyXw57Ufa8y02Wne/3bglbHbDBlOLqHDbYf4FHjI6W
vxv4waJeUrLwxK9fvcsF+M0i9jwbnKuN+looQ867g8dfY7yqvC+T3W8PgNygl/CUCtZFukk2Nvrx
gGuyNezrhX6Pgv8gILA9bLI0V+BWRkGsnTKCiB1pBJAh4SZM/WLBIAwVLDyqIEb7OtJTcWGPefyH
I6kTRmuR9ZOdXVcSaPo/5OSwK/vFJn+1XBptcUkXbz4czz+aafWfN9SKAGdYxq5GJ07DSs1Oh5Ff
6rOk9VncvA5VNGkH9UtOGrVE2lRTrjYQQnVpjPdnVXdjzi43crDeO7gfqV/12f8woNpp6c+4HJEy
rtOl2q64zaXDC5dpiwG6pfy88wsTdJNW3X9FH5sgyzJfw43OrYNXEc2nms5ZWh6uSXzitmcnK3KH
vlUy1/GSuF/2nQyTL5bRWUvw4y/mwTeFO7MCEbiA2Qvb+1SPKtQAz9Iq8MGZCct/dhuTRkT4uIWD
Ne2FyYXRiMo7erWbYZCN5YCijV7Wme1xDgWr7jttHL/rjm4isyYU1sBBm7dEXZpVoZKhpPZoFdBk
2KJwmPX16+WVgRhQO7gBWV1uk1kqF7dOg0vnC7NCzxXV6F7Qc8OPU0QFPkygwFOen1S3zimGDW3Z
I/6cL+4Tu8my0p/485EGQ8NynD1tBfBok5apanx6D28C+UqxAHr4/MBla9IlFvDCC+2gJKGKLkGz
z7kxFURtEeRexwOEYujttgLFSWHxrX2irujcMFVvdIPZMGMn9t1t1/96y7cinGC/rYyLFdN7RtDP
BJaQX+2VqkfSjzYuoNSCsho3ZNjDU5OlAbhydpXeDkr8rrS0qP80efEEKTb2Ph/FjVFz16eda0cW
Smx8kEigp7ZhmV8HPc7iVd9X1oL1e3k5VFt0jWOnLb5kFsu5wYTgJoh48AwPMm6Jd9wK9KIOi6P0
cOheLp54PbZ6R1xQVgOYl17mHB5yZ2vnVKA+WpA+jLEHFxmfmWUf7vj8ryQcU0+FiZwJSh01RsY4
EdM1RPysgYJ9jA7esYaDiGpeG8u3LChQRN386yA30oJLOQlq/FRFfHy6EKZFf/P0c5bDbIc0pwxF
2eP1gNrn+EUA3TjgTymunqmnxkPs7yQA4H1//denRAcamOJJ0fg7wXAx6aI7FAvQxccSrKbSuX55
aKC/lbrU7w0YRw2HT3oQOzGk3K8c9qO4V7ehcxrKpNLUD4+5ntfh3RxkXrXAJjCMo7Mjgg1K/7C5
rOhK10cK5MxM/VFsOwmMlDdyK6ibj5XA85o2lcNAFIOigawITkQbPdZ/epgbUJ4amhGbxNYyXHUo
Hz5Q4ktvI0Kh+FYn3CB0OyEiWzykhezxJYQY4O6pcP7PmptuCHeIxCV85fg0jm1MRSVxEJ3f0AYS
03nRNW478IH1Khc4qzBCCQ97lXLpSSq3bhL9wezaH8clcq6QdQQhwS6k3TvNaryCmICcikgXzLOK
9cpr/E7MSACWHsRqG2HwNSgKoABENiOERVXHdXopHGLqVnEBmXG3Vni7YIq8xjzISa8sASeqRLAo
+jnB99/EMsQw31idhCaEw319DXte9s6t+DeZYZWOQsiqD7X9hhbOsk3V9zgA7KHm/wBropXSX2X4
4nzL86WeaWFRVPTTATpji4JOyCk7ZZN9+AnVBwS0atNyhvkOIJjma48cpXgelfM1wcfI/yuvxOlq
qXzaeq9jo2/JkWpK3eXz1OOwacQwlGhiTGvysNLxBIotMSkJGrJ8t5d3j3jomEZ4lbKOQTzHOaaG
QmELjxa62B75bwX9c5eGwcOW/dWIEtcCbxeZpn0dXBEG9HFEb+wKpa4+ZPbEnYBHZvrZK5wZpO64
xNPNUuNDQlMty8AFBKLzqA/EASpsSzJ9idQOnr3VmyQg/fBOoD9hP22VQ+jw8xdllR8HG3dz8i8C
jM2Tys7fqgNZ23n4fe61Z49WyZz5AMzgBfi7YUHEVJdwnhbLS2ega4sDhMUq5UdpCBuhqeU7+KCR
sqganQlr7ESZtGp/uguR8KgKOHqXMbjyNWtXq0KIyCnyhPcZn+ceh1JciJ4cLsn56aXZaJ4JCsGY
JYOt4znJexuzm4+/6m/iX419Hs86QFagxDXVnHymSIGWWqabRu4reVJPmp8gEwxGknay2Ew9I25o
goQCu9Dhf4dI6ToEwNqa3rC7bO1OtwSy6AOBHxpqVrUCy34AAvmn2/JqmAOFMjT718fjP5Yv81ve
CKALBTM3EpYDxP8zJQy0QbE32UvBiXVrBYlayTpI2tzff7jlndGLxFGSbKKutw72gL3Ss1XFcQEc
xmaCpCkke83y7bGhDVvehdz3ZWgYlsTvpxXdXnuWtmmGv26lbcbtAzhzJd1q6mLvPnxCVdJdZccx
pPcACvMkEJeDc7WQTA6wGYoKxDByFdEbu2e4Igz6Ke4X3qTH4Sz3NuWFg0jvz69MXvERzrNbTcqj
ThTtwarhEwsjP5AJ4GmD/zr1fP4P6M0TvszODIoo8LP0uscVaqEJrsgPC1hIAYy9VmwlTKKoZF8W
jiqsFSAwPKqGFtHqoulXfN/aM15KIY6PeBOWUN5MRMEFMMp5TeRvVJb0mXfjaqhn0Dq9pRIB8VU7
0c77bpY4UvZ9iQWXwC0wDg6HsJ36ACCUSG05dVJ9dYu0KsM/iYIL1DZUlyoWT5StcdIxkIwi88Iz
ME6hDnZmPZIMNhf+WCubhbPGqOyg9TmFH1CizwzANlyO0jKFN3xjckcbHIfJLIinJnSBwZ2et/jb
apwr4UKsHLBJOTghHUJvwILwYFHfZbgJiSmwBefmFz4Awiw0FPXkdlDNODS4mWv5YKy9MNEzHTLF
7p4sEX6MI6mGMIFV5WzflF49qwWsRSjRBWafCEjx9bSqNCPqfWzur3nSO5lXfXpp3fVqAU2UfDtP
hGbRu46VL4cXCSvwjqq5iatGhll9b+pCBLdSWAyOunBKfVoqow+1WHL0PfwFb7Jqd8ztkz8c/BSz
FdHyhETNQYkBhBGRMk8qn5XmAckL32HYsEliBznDAzYeSc9NfLcARTkUvWtuSXSaH+p+Rx4gvTjg
gh/3vp2p+DzichcogOqtwfT5rWrpJxOyY070662Af1atgAOA0WTEgrcrw9mpys1GVxJnkREjB9ug
Mp4q9ic2bckiWQuYHwglqo1ymoY2awCV/ETcsG0u9EXDIDdzJtSpBsOPXluQuVaW9VNqxFDztBIO
VsSR63HDn/w05i563KhvbCqk8pSWN3PpNnum3vpl/2C4zvkG9jlSkTaidQ+WbYx/qqzEQNPEtEe2
2k+29DubOfuM40o2hw65PD8MDUArH/kIJmqDtoehlfYIuvXE6zCRYN6hbMW4N02OMsz2Mqw/m+jW
ZD8mH0jVx0DAXpu8dKRZfHhKk304Qp028DmVIlyFh1B6QysbrIYzQRIlf5HqIpAf6OmUAiQ6Drz8
JCncz/R/HO6mmPMIx2tdTGshEzIsBnS3Ecz8w89QoXXcRUyPpiqsZ4acVT6v8BVf8xRs9wAiw/XF
WCq6zan+wLIqEsRtNNvU4h4uxhcEy2LnI51luUNAkAwDOjrdk+6QMkmG8beDJ8qnTBMISmX2YKIs
ShlyUAv/rLrDz5IyiJ4oA/12DznB4VdrBGsH2lBhL+w9vDsx/VGMBFACw6+Kpkw2jplrx6e8Sc8G
is2MJccqx0EK1RrMr1dMNT1UGXN2GVOoirs9HxhgA1Mx+N4/UfQnuGDlcD4RzxURIopa6GuGYfog
unOsh0NI2ovuGcCq1Iz6XwFJjpEZ+guy3P0Lm1cgSZdH8izrfki9aaE9sYaQARPpBifvreUY/E+R
vqjJvUxoZO5/s7/OoCsk1ztfIV+bL0vMzf8lEXGzZ6o5zH+6V6Ub0vuClD1VabkAjPXXt37vwfOa
saBcvC2fqZHpvWJULR7K6wiecaqvYLyOWEtVxmXsTOKythQWDOhTWCW7Nk+2SCvJnVGcrVMdpyT9
dMi6ZDXnGRHZ87Igp5DC5b8dGVMpNuy2PCyELco0640NOQ8jJvt3GI6a/TCPJVkwipmtfwJ2mj3l
PtAOvwbZMcQfMg+YdlgfsV9xDVfb2FMKDynHxg60HOS+yMgn8im7Wlb5Sug8j/3nx1dVxcktch6d
uYH1JObpGhPxvgwf6BOkbmjhhXB6SFt3GHSBvowFtjLVC114laNAfgmsxeIN20E+V/KwZxIJLAjo
NbsJ7uc9/WGq8p/2hbWnTBHyhMh4W7V+CW/OPKDxQOtmXQz6ihFjpnD3GY9o4ep5vMuLE7TBgnRA
S/Tl+5v72SAv0qJ5QzVcEK2QpqL88IQXe5LOmlr4QsNTv8d6SrAIkuGDtqzWkq7Ns0WNObOCtZCE
dccdljtZWYO+4zlVX+PShPNpRgJ3ZoyNCHYlDTdIXMhxF2sYAF0K4oaIt8sovfReiHJlxfg8JUv9
szZ+1T2ZfxR5I68w1lkaXTAxGd0+oH77dcUOlkSvWgo5dmMi9bH1laI5gz8BKNNjtSabiVPZtt2E
yKFZzgI6Feydk3idLN2aXAFLtRbQblcI5U2l/OFK6le9i/uY/ZGviLCIFMRm86VHqKvxuw6BenpS
Xlvm/8pnnhWJZMMxt8riy8FF2bhaBB4qTQW/Y689xY+XSsGB/KYeyn7L/ReJxinhnpBHW++rWuCv
tz9b0IKA/yKH//FPGRUxYBZMu8JhsNgerLJyVaJ7y9faI0NJz6b67XD0Q7QXnRjiRr6j7ZcbsD2q
FRXVKRuXtZmqK9govRDpUJj/A/l1CkpdNwmpVZGQYODiCG9NAp1uowdHW8JuQGZB27HuUonheWTl
TPhE0cwGeNkYN7snWX4HncK9Cyf2UEqP9JMW+RXV6u03X2u6c/enHRywLRlOHooI8b8T2YkJM8dc
vu4lbswQVh7Yk9n1QMFJgJyMDDtVyy92kYgGr2pwiMLPu22TANJc/p5kyRg+9w7QerPoRSz7/EHz
/473BgtaCzJCRDwUTQ/gKfSe8oKAUnPuGYogDUTsL395yxBxtUlLZChPU9JTlp960eSVucBPw2qC
RTfnYuFxLdML5e6BGhG20givAf5U8SV/QqlmhGgm1CenHmj/c6B/IEtS1aBiKQVZB2sv6eHfFZ1U
BDxPafOMe1hUGRc43jepbsb2H6Cowe2m+Q8khUzDrcTMDBDPH8Trxb9gME6mswnqH17dqPGyK8dL
fc9mrzZnt8OxfvfuXtTTcQCqLWZKIQs+yD7/3gR0ILTL+pbWsk3lyYc0kChoQY9PEA+d/8KrCs7h
3M5xLDSD/vaAvncO16L3ApcSbGKvLvZgPe7vB6sFvlta+38vhKWoov39CeRMm/2O4h/agKeNAI93
3en1EnbX+5w8nv+5rLTcnNRv5MTWU/V9LnHiAQfbiTD5z/hnDGQgrEfbaMZmbhEQW5Nm1T+xmNbA
wUdRy9/bEjLjImUd8EYGX9IXJTyjMAOOFLX0D0CRMCFTrTDxGd4R1XdTvOM2ztV7dpuUZuqOaQwd
rGf22EbbtOEVQlpf8m9tSnXRzZk9yS5OT8QlnGpQ6Rpn+vRXSGgUQo2072OCeoKJoxMdJi1a+olf
H/2Lolca+2de6IvRiFiIRc3hgDajRAmsPLdwK3cQFltK+5uisdHOdlXeJviHxj9128H/x5KR51+y
ftKNtTA2jJbaKRUFCMLVzvJD6mewoBGOggEy5rmyUhKQOgObppIC/mZ+i8uKJTZsLRf/dRVMjpAk
i0O/4UHBb/IJAAJqkxKIaQHM+DJwMB9IQ/Yu22NUqXiEnPr/hrq2REZC5CY+0nKRxxRlK9L63+lR
yT7kL4rja1K4KoQyGJRPsGhWFLic01jEpr4Lx+8zn9gLPT69uoxLqpebIjt80brOxdBzGhNIYkaX
96I+q7zFJF/2TgupaAL9Y9sQzCUUZdY7ShPJAUKinEnaSdKoKFuks8lVt2Er/ogDEXXQIwrO2THT
WIcztFawWpv8leWFuP865nwbmxY7HzlOAuBlJFAyZenpUs0YSyN47XaZ6LWAZse50np1Zn5SyEgN
ny6RSFXe21rejMm0WpkWGyBQwX8+8Zn4lDSqFwRvZICb2LP10K5Kb/hOVgSdtywf/DYXzutQ/ehp
JrZppW1IxQJO8eE0sRtLE8XAlFbn4kfKyD0r5tcm53p6eWikqtNMDG+jt8I90fDr+CBFH2PPh1o/
9RpL5EvOWUWvTsTSXisZAOXAW8QztoaZpV44wYGs4qQRDIc1dJ/EAnGJgBjDPjWCUrgbLyxFhl5C
+1k8dljowRuW4Kh4xNXdxJlBkcIbS/cMFVh/Wt4BF1yuDfjBdo2gCkHWAVUqMuk7LGLtvW2JANaj
1RlbRoB05fH2hbSoDXkVQuprFudTHilgFYcJfvcZIytNqfJ+0jZ0zkKX+20nwHiMBu3GNG0zLH04
ZFVbCQGdCX+hKALwje1nd00ZjysZRglGehn7HOrSlpbvuJwPmvEFAUsijNmu6IoJPQLym27E/H03
PmXk867sQozAeWe0Y8KI8GvHfDPrVTA2yYgZ6tU7iQjwIJCKjeG8nBLPVoeLWo3sNmgVIpu/Fqe1
Fmoou0LVoj6sQWTQTVb2TWkblTV22W1HGU2tv3N/LpEcD5BtytBx3teebixyGyZ0cNXRGoodfPzx
5n9VKZ1rgS03V+z1KdyPy8BWjzvLi+e7jC5y1VsduUscI9NS8vLBW9uQXRX2Y1vEhT8eODNvX3n6
g9U0+CBaW+ZcxN57cjcRs7iaU2WP6wcZ1KDtCZ/t1VB15o+7BqpMXudygW7scfwXyy2//swatYzs
sFEuLXbmuNBilxQ2XVn8egcoFDAFDxaTtoDL/+PDxcr55ybfzOXaXUDJaOmLv0cu60y7I/+KBKnj
LFZ2nhc4YImgxgBnBNINXTGZA81YV5DlHOhvOFI9Jnsr5HJ2fKFT8m9rDVYqg9oe5YfpWRKlMCmK
sXjpKaSf/8QayJ11NuWJKWv+sCp1V1+IcopTnKKzUqh+TxyoPXxqWpCkwLQEastqmgFrBu2VDxwU
TXBNn4FIWQhVv+VMD3oVkKDQJus7ePF0XOH16L6OUKILheQ8DbraOl+39vQPdRMh3oYyk0NM8PHf
ZfzFeYSlwefoEPr6U1XiFtyb9sPX2B84wFjyTv6JJnvSW2iyLjuGl/wd1iv4A5uECYCwol/dX+wc
GjKTtdfMNM1woUSHiRGHvvFg0+gM+0sZyUiBYgiIttlkGcW2XNvIJRc9lc+eX2iLRXou5KZzYxWi
To68edL+sNkPbIftZLsfSuRjfrfp+Ms7gaqTspgmlpk6KOBEzjSDX/QUvxlA9Gg9Or/HZ/2xNseK
iofXxl78OUHAFC7mJonrJZSwJi3fWghXr5Q4kJFlFVIDCYkkiJ+ecQw3cOVPTakUN1O9ZBzrKnJf
hJ0Tt6JmuqOta2QqiEyT5GxcYcj73A5YPc2f0EwplIu8OcxaJo3qCirQnMErPR5RQgipgSb41c8z
+U0Spv6TXo+O2qA0ca0XPo1k5i1ASjmT720tT8ui1Vd0bQrOGgn0TJsDkRKN6OmNKn7FDmPmWB29
5Q55O5LWJwryQ0CDVfMICx30qpQPTHKfnRQQtadyNr/t565NgIhHttYckVV7nlBcJXzsmKaT0YJq
oVAmznKp+qna5X7jWIoRkPAoBjqLNraqHFjO9pTKToLxQ8Msz0fpoq8tUctKZmlucCDmVfGECzLI
eMzs9qAfiXjUvoq5yz5dYotoz4Nj8IOSVbhi3Q8YcTAFQRZGgTGpa8r2f2vYyfXVOhVmisTcB7S4
cyO2uFuXwg30DXhbuOVNPd7419Iv6lKCsMziO5LyrcwXNSV9bRi5a2d8qmeMY3Vo4r0MNElWEf3G
kp+j1/02NOnYvIaK38jRg/Y5S4MdZWKUHgzo9kdt2nUM5p+Ee5ZiQd76rNx8MGFVLVAW8eRBdC3r
JlyBhk7dLqCNkxMeSEQHlcqaaQ2hsLxB6hMCYzQFms5X3/a2Eodg5EnlltNps9J/qrCplFG9LWb2
Dio0ohryHbjPjGpXU9Zr26AHRpxT73XYyZoPnaMpJF1xQJuDt7m0FI+Qr5YAeqiBe8PvY8eB3bsV
h4nR51lxFfV/T1nGenczRrbiMhZm5Juv1XKkc/OSXQ9q2E4uRaaY7NYg38/BOK3q+Hp+YPcXpXaS
SH0GyVB/9tLUMgt/v882kgLnFoPqKO7iOKSFmGb2R3X94C/v3McwDkhkW/4j0GNHjN1FthVf31BG
d5ZUnq8Zil+ucYK4ZQpFh7pajAvcpKbOw7uk4da5l6JgzlrlZaCRCvOz6dfo7O8CRSnlSfhn+r3f
ikQtoQpz6RlBd3Fb2+9JCaxyviV7b4LtJiFNo6lXxXOhaFTW8w9XlBY6h3w53purlxRPcwC7SHok
ahQnWUvk8cuhJvWk79n/bLjw1ubKcBpvga5j2+PGztvrX8D/5diGbX+uWKE/czjoRHnLuyWjcxA9
XD5MBOCFhpZXAo7g3sSIq+bujEXViuXn3pkxxGcoq549gRQQlBkkYYlkFi2cG41cZvc74vCEj+sd
/HjLST3KgMNrNS1Oqy+PXB/BH3A7tNedhDBq3BdzbxZPpaFhOyrtCFSWSy4L2QYbz4P1XHY7DMpI
OH7gK3x1yWhISCsz7s/4aLdPRoX9St3D504kkSQf0/MGl6b+lAHUJaYBmMrTr3nlIlIfA+pOByjp
80IWVoCqeq2bHkKsUi+cHBmOg6D4kAsx9O2jaqk4kTAPJWbc2nTf1QWDnKD3R4cGE98ptDmckeCW
iPOapTOjyKUPcExygIvPESB3q+3oNwP/ZPw4omvr1mJeSm+wHh+stfVlUvt0AoHJ/hR6MpwS/tWx
rAtkLD60elhlmWRIVB+PjfnY3LuJlFwD+xa66sdidh0nAjB9M5++BMFTv5DJYDjxvBpmnFtrUQsr
E8gJTxqTfk5/VVeXc9PvEh9ISjrvXSzT2KSTACpdpjhhcSF7iHe1Rfpr+PCbR4YI5wPKueewcHF6
TDtpQ78Bjc4iZc+vL/cVfdKwmKRejLJ1qMQjJz8xVLnLmt8Ua1ooSJWRmNYpkb60askxm0llMAwN
NQ81GJ/LMQ0WG8pE11dMreDFdC5VOMpIQE9isUGPpZoDZ2/cIX7IH6CMQURfccnt6DtWLy73ATX0
C1wMFP1fMnRPwLJFU7M5zIUbYQ4IoZwvG840StoLiIluqwSZItz+pElKkJKE4lF5EiFFghkXmA9W
foGqIxv7y532i62rsw9ntLnqVD/LEP7rpam1oWG4uAh1QsX44m0zfm+LaXMNIGAA52WekRCPx0t/
rxLLmrDJUeKPyq70X6IVru2war+8vozBR5VY7RqjPFfB2xEMDLf5LM0NobpFcB0nt8Aeeqpta58N
V9QOWp5zi1G0eCvtb75PXe2lMz+vLtZdfiGDGsLkom1zuJVkWtKu4PQZb7OIM52tqX09QMxfWtwK
SbsQTYsFieZZbk5m4TFo9JRBWzo9BmfrqdUwx7HHSVpftm6ifcNDy88KhEStcXK1AW8awYV3MY4m
DxkP/fR9El1t0p7k/OrpxJag+ttPNe1pyuMHcLKzEPa4Btgd4/XGxGWA58rh9kFoTleSpkbo/ifE
sC65rdtC9C8iLF4vRywENr2CdmwxYv4qtqQGpxwQOOeLf3qLjYGcOfmDF8sVJXJjQVyVydO40QvV
PVI8FudYq5JAS7kz+cEtfasJb5gCLViEs++1QF981hjrnUE2BjdqWkkgCzIxlhF7TWgCd5lFM5z0
Tk40Tem2jD9W2e4Eas9TiKm7NTxWGkoFYJ3d+vO54O7jqpNTUithFSRG5R+ys0FAjWOWR2894o9f
goFQndugkcwJU6pyvXcn3yS3fcDat0PzI64Xvi0oGoSFxYWGDT6YmqwTIUpIcbNkQFc5pgNXz74w
utE4Xd4VgFPU8EW2Sxo6tNFducBmDVkJX0rYLTTlUGFBTjHxd+bFF9TVdIbG4YZZU8lk+NA68K2K
32jWHSIVFrM+2yiekBmmtaIVazzH97CyOdGviuaBfn+bi3PZglWe/cT1LoEaMxf7p9AINU4XOh/r
DsCsDwv5oBTxAj4nZ7KYHO6lgSmU/8J3Afy+PaT4jq7nPFK4PGeio9Xrsx/Vx/oK+YhEj0oUv4K8
JcObD88prq2NevzmiAzqjasY2/CdLG6krX8JWW9Rnx2ogfcGLlaTFDsa3/maBnBTlhiA+NojhUMH
OKNwNknYd+tOOYGnfjE6eGDeSXYZKF5YlLlmcsDlg9yuSm6CvPlT4T3CwXayMrRmwOMC9RiRzFmr
zxXSntQUxOwMleJxM+gZ9L2ujJjmXCmueMuR0mXoaz1O3g3idiA217k2Br7+Yn2xFI893FWwrkai
1XnXcDDngp3CNHLQkFLdxFunsdCJm0+V3/KXW4fKi/AvUPx+eG5Yz+AfQlSuhTQbQcIO4xxLmStL
nQ6+qR6FsDtqQXfvk6CZI2ZtnvXG+agofjWKzXkyQAEowqSxvNt+b6PuhPOdQ3euuzdIVXiomp+z
xj9xyZF7ylr9BQKcY+cL+cYMM2KPf0gcIy5oFOIOeWklfNBMH+38olaQkKy73AtqYzYto1BbP3/N
9WZOpRtTz73eC96edSw0YZ+mI4nlN3cWVrL0xLImywlSKiV3xBgE5cwb6V9vU826lDPcERQRzrXK
yMDft5Nx/3IMNwDmOOXpadivBOLW0ZcArOzB5i78mq0jQyC0F1MtZg/jvBkDf5uk4MsGSwfNvWIb
yx7PBgnvQjjlzi7mWZeLjTsIfCROphMVGcebGZjo1lVS/auVFVRwQDYlMfn81dsezXKUm6zCnQ6H
O84MeIpPLLPRYX1P8+bm0Tz4Ox/Hz/V2TxrblVIj9wXixRGr+I9z/o1UdcMHowxulQDOjAASRY96
A+jH55B7ICzEo7w4UN7widSGnkrDTpPX7GOQoVKWE14BsbHq3F1B743G8EgvPnYwm+JdQP//abNJ
sChUqp5PIVRkRsG32sXOGCsDsv0ie9qRjoag1XmmitIwFESO4n15pLRygxdjwp2jmEEUK242H1Aw
NcoDT86e2lpzTJsfRNFBqz1VKbzz6P7zv0J0pi6i0g9H3QMTb/LyT8ZwXcKXCaNphRFMFgxMVPQo
ZZ+jsNHolKy++UCDZ1hP+MxD8EPoq+B98FTa4JCieUMQIGkNHYaYQvmioSCzN0lncWg7Eg8Fg+Vb
l++4slegMdUoO/bqb6T6Mt+Fho1W7IJGS1gnLULfL2RpU/CkKK6ar8qHlsJxNrp/EYubYcvIlt7V
F3KiWYpJb9AjPpvxXUEskknseJfuc02C78wQByjYVhwMWC5+Atezm4gJK+74E1KSmZL2zKHxtItm
q5U/jQFxS+xTd9CGk1BRTYVkTcjCWc/fT6/MPRCrkh7mKfT+KM6p1NZCqfUZ3ecMFKRSI5oJMyYO
XQkPxuFq7W3Tuo0yI1U1ZPcYVb20Y0us0WJYq6NFsB1sgRtxa+kWhPXjtUmNDXqhKO2ysz9zpuG4
r3/QKIf/R1a3xGyPTUQR/HNV3c8yTwkoGkwli+b+4RWmLIWPwF/h+PrabhXpWhosPb33h9RdXYwy
z1pdUgkiaBaJfBi7JaeYtjVqFPDdGpBOHplwDc0sH0501LQ59PMxIdd6ygDLNRWP0XuPr2cZLLHB
1a5vbphutNnTCRxCJFCwMJEthDH6kPKDQ83GV67vM6c0Xn63oc9eEoabW8yhWzUB5H3FHg+DVU+H
dXOREXXGZjSbeERu28BTkbfbFO8AW80b0oeHUeYnsegQvjPVXXuy9pWezVqQ6aMP2yyQaAHIakLg
6+HbWjAy7WlrAX5NAtKFY1v5UxNOpr5XmeXfvOCkxMKyClj8N1Rv64YkwXzW+U1IrNrMcuxH6Rmc
Y5OGn5rdf+Ny4HRad6k39zXl2uwC3/GIxNvQUqik37jLeK+iIEpBqJVoyrOZxEMYC+R53Xa1vgzA
7XvudaUetnbDbxrUl5Yy2RRQO36gIMokBR7k77aPgt6mSse/KLK5PjC0Dl1EbkIQnfyVLSQ2df/b
95Yj7jHcF1WBQ2ek8dU3DDOcenCk+5OMehxDRV8HiBWg1+znmk7YGK1fh2fSbCKc4I119YREGn+r
60H9CWpSe1E30nOb+1hNnhPq+2AEQp4h6P7Vr8IOElvcR/PVixXl26y2r1n7exGRw8e+lfNgWOPk
HZrN+ZSmEVP/TaxcbGn1UcR3YSf0OycyLvfSq5BNytMy1eIdaDHxmbhvQjJgwUmYvaXdmVFXzNVh
MYtr83ud/9267SXeEiDqsWnRQ3eBDK8WbLBoKsXsN+c4kkpiT8lOaV/IYhUjdxSKPMeTDDyPe0vX
4RWLZAPyS5iiDq2IosO/2GulSxDCJh2wyV6WVeRqHeqYJINZNxug8JGc5GSJMFa9hQmRKs9FWdMD
Z99tWrLVNdPMAioXU4aPwEHkN0D2K+BBf2dBPkp15yYJRWInqnhYcm3L4H6SasOU+hdMHrETcu8g
KqNzrSUq719K+FiFNSTNzRrv+1S31LUftePdLr4hBmk9ayteQjqLEQAPW/Bp7lnUPDrccHUP3SEr
3O75pHkMGBz9tKVUafVNJOTV2as8+afqUlIeXsv8h2c2B4G/iTIowBY7qJCzaH+6/6AMZlqMa67h
BP/y80Joi0alt3gZd7zss/2Efr3vmarPjR57WCrhzwK1GkCZ5WpLqmi5ggecCUeRGyGkePbl91tr
MTRrayDt5fnLWYLbwXfqhh6zwvSRyIzBGDCtME2b4EVOX8vFP34r6ho7jwgQ69GK8tN5TGa/F6lx
6mxsu2ShbG06lOYRGFZcPe+DsRRZc/ogn+AnBiQEzREEYuoNSldOPufEHVVx7BGvPGUGq0tM0c86
Buf9LJV1o8wMeoXS4xe0zwHAQ7CModkMHKF7bFvtGKjlIepaJoO1OSfec++r0N5zVlm8JzSY+2rv
MOhQ+1c6cXuY5eF0fHYOuS6n/6QhqK5dDewtotE+/lj+oo6f/+GnSju/17WcHHiMHbvGCjASwrr+
quFZ7MYdi7hbCQAtYtrf3liIK7sphEwtEHYSW/+PTk9HX9UU05AgY3tzgRcvza94Rd9dmHsMdFxk
waBVIS7Tj2TUhV7PyFK86hWH/y7V+SoIYFoHX0ibnaXGwhmPEJDjv01+9WeNhVXw48W3RMZN0RSn
dyJ/8vMfAndYJMa5DWfuOFwsRkWPZa64H90E4lGg8Tbhq/LXDgMPw8/Ih1WisfQKVvkOBiSct8Xd
kuqSexIPCkIWN+Ku/V/3oCBNJVYySQ7F4K7ydv0oNHGCU2tqU9V9g+NzsTnxaeW5FIwTRAhJLX2r
mfuhBDbNQGltMi41CQ+q84/H/TMhWhCn238WlWFbEhJCSV1pPEc7nsV50WiITkCkHXIwXe/5QzsY
EHNEMqsPy+0Nd/0s44/X8lDdIp9vmgJfETrZ9ykpZAI/MkGAKzNgE5Aj/KxwaEC6nYJQFo0YT1f5
L83IbeqHNG1/S8FRdEI/pwHD/qi/742LqLUKNWnB3kGB221TfXmz/8dNVWKzm3ceaz0PfHPJQEuA
z0JRzgz6dK+NPiwnNxB2WAzrmNfSwd+2wQXI5QLJOB7p+O61EJZTZ16TRhuezfJO9GCIhOFK6NYD
S5CCZO04C2OYkNl7m/k/L2APlH0uJE7LywfwIgrG8ugOycWnnkr4ucDVsiGcCqIINt1fdVx1R+Ez
2kEsho4LbZCfdXbWn3bfEqnfrXYI91xsJF3QIgd6/0tnUJgf76bcAovTezaVpmZZZ0Likok50P3p
lsRdmj8SuNFcS3XOh9ZKDZdLZxSs1aWw4ytRLFJdOa6Njwqu2k0USLsLYXx8W0krm393IpnS5Fe8
XG0jP/LghXaRntOcAZcbx53UR6A10O5/HjtWHL5SwOAcgI54lkMrq9oWNR8kirek0Q1A/BtTosUy
nxxGw4aBzlco3rXnv9bsLZP85/zqkx797LBCrlTwpW+sSoPnszs6IhYEwkKPhBUMPlsOD71gCLV1
HBNH9EonQw0xsTqgP+zgqcI/MFYXNiwuJhWhsAwtdiB2zJSQDOUYNXUsgd0eAzXcr/o1DTIeavpb
rE7gwEz92tllqmrytvqZ0edWdGcCeqbEL2SAwN5/swDZx7WLN5y+3FLiITIGFhpg8RYCpojC5Q3m
jSDS1aDBSEirFdb25tIcqqpHgoRCuRbeq4twDYZV6IaExkHOZnZuNY5WxrGNWHutNTo/aFswWtmG
hF79TpfhrsoUe3ZBll4cvBwPmW8+HR2yvm2HSo8mg3I2UEPPqCfdW9eMDQQitAw+oLBujiEVsw7i
LWPkpNxusXTqqC1RU5NymRUY/3v8fanDbyKYYhnggaCxu3I3D1ioUwF8DyI0aLlDiNywXWG+yHV0
jrPJ1Qr0ey6DAbBSxFJajwCtGA9awhxQjkSb9CyEbc5CXtwGu0/ycg0RDOA5AOKGZpEX1blA19l6
8U52sSCcDEWucFG/vm+pXARnnVK481t0WZW9Do8sDSsPdVAMCR+1NnuEdaT7aVGr/NXRzk5dqj1R
0CVgVtwYzTJvZQx1XTdXzLXNWXHi8oFQJFRN1mfQl2/wCgoDqDL9x2+PLYW/NpH+FaWoaPILHWlZ
3tHq4v9TQ9unoGGuEF4BkR2yYAQzszknWjpaYWeC7f22xklbKNMhZzcmeR12WG2LVMxJfSeWnrFl
rnH1+SXo3ds1b6rJze1xm4E7FzPIRQkxgryvais9g5SC6qQqq/dOxmmkUrsWR4KD5n5gysbsC3z2
G5RtbobZSqXi8FF9EboiEEC3uPA9qylNflePc4fxnbXdqtZh1ilr+Ej+Kx5zhIfDBoI8gLGAgJ7B
G6xeQYi7tH1L6Ovpw97dtM7fh62bIasgd7SEd8e6WcpeJoaCWVDm4ta9GfhKm85Q0Dn0lN449jnY
47fYQbtEnRExHsN1Z82Y0SGR9Tx68GkVBmBtHSupxshyCMHgKd0LknOxPa32Hx51b5F+MES08eeD
dzTP+lbUZj2UDvXsKwy6zmcMFMOZUDzQTHIutWT7MJFB/9TgMY+fTme53lxI17P/tG/VE5ImVQFz
bWp1c72gSoxqsgYT9CCMFOhlOD5PZNV9Dy6ZkVJ9LauGNJ7gLanF7vJxH1QIQuYsSMYQr/dJRusu
bYOgtVadFLbKVGSnbwZLM5PWXaAOa1ZdP0+34We9UizQ8LUtUl/9ApqzK6zbvfRwnpyuTaCOQC6e
Lk0r11Mqm5bjO//X4sofA9e+PZ1VS2hqivPS4S6r/VGZCOFqTxzPYpslHDONW23MeDvhOZTc2+I1
6Uw1WbRLrH5ujkVGKTGGEeF+z1nLMrLxLihf2AkiX21ScMxPpfBv0FBu11+NzlBzGBH8Tfq5veFx
sedJwOGG2P6bmwxFjFJTXeKbKEk9uitgWVrbs5D3aw1MCPcFEAaXIAc8U6m7J9RnlKFNnLRKD1ye
vvu6gid/20oQiXFtuW5b6xZUbj2f3VevxFjckyCEN1RiQCmJW/pVPzAzUIjH30DZ2QRJQQNIIaw9
prH9WHWXZxFC0q2MWAhT90ULQUF/aktzFeJBcJtYdoyq+uABZVknaaU0OupDgiUCRiDH7mmbWCrs
Cr9wDJn61LMIfvJ3wNYu3KL5v+mWHAyM7ZKKUqlO7YqFkYomhDoG8V1vf5H20GpxFFNuDRPZv4W/
lLwNVW6Xki6YbZBvvI59bwx1o8tLlev33RW/bLRcc6mAgePDVJt/fDoNMpnhwBmi0yATQ+hJfIKg
CyjAkmtAkcTykm+9P3c+DkcfxDhcL/bWolWVh45xEPyU/zCZ8Y+PrD9dfJmSJ2murbpguJzmyyIX
fwNn/Tu54Wr0I4m0jVIB6I9rE6ENrGg8x/K6bMmVWxkmR+UjK9Pb+nzbA/6+fKx61a90X+RsgjVv
VfCtUnvdACyADy4ocHcumo1wogahT0lPAke5H9L7yoN11j5Ol0sqXNw2V61hZL6bzfTtHDmM/qwb
2BAHUNWukPgQpp94ydFGH+Tb2Ze4gQY1gJNMq+/qKXH+QcXcZ636IlDeqdRGNpiv1FKRjSE8Vdsh
NjatAiwsav99j2WkqdQrHHvoReI1OSDaB3lnz+jnDKDxysThdZvkVY11To2MRv+1H/GfFC58pr98
OBNAnO2WpIbLzSRkjiFeSGVJPxo1YS+zJulXJx18a5lNRW4RayoPqiXcIRmp69Z4SPdOBY43S+3i
bXOWk/HaC1414bh2Nc5iYfJ4PYphVb4rn68g5Lhpa0/tjcB3kCfmy2QXl+aol3j/lqOMnRN3r+Sr
+wtbLowpNdfNPFtnEhvuYTR4Hq2+LNMnekn9NXQNMMJ/Vuk6YjNjFOOaEjCxA/1FTsjrbnZwZpHL
EkOvj4WQnwkOt4hmEZ+5P7ZMXddg+0b5n+i5E4+ZWXUYHUGOivL3ZSoBzacPU3IHDWNq9kNX2DXN
WPVyFra+fUWfHpl4BdC4xSGSFXKVS2+puaZ0ijWIFTKxU/YmWl5h58vjQYUHZNm9uBx0jO1cyqrc
dLiRJkLzj31gIdsW3t5/IGPyyFt2TmorxjXiJQx786LuYFmFNMzUwHIZAfb8oQHs23aDdefOAJWp
AojKFvy2QWRGDL97nqZmBG/8o+9elsvoZ5ZMzIYdJW+4PjLN5f5yQsnL9tqNUtJd0iXcgEff+9sj
b3/TGoJzU9VtBlJMZPswxZpWXNCFcBXoqzY8BiUXIwFoG0giuBxovGynZNcuej4rrTLrr66kGP38
yKnADHXGdY6sxVE/4XbDy9sVQyuBdznTPGBjh8RZH+/WG6kS+jP44EphLJNTOD9Si7jwKXUgAtZE
FbowWWzkzBuWG9KwFjNwh+Twd9fOwTHPeApEriaH+877F6yPGcinp1zQP8W3ZfvCOh0IJNgPTScF
lvnfF7B3zfv3Z1Stb9g6S02rTeP9Abcsu3QXDysz/9Ushq8zzTMFTqmuw6QC6p4IMR7bm5mDdLcU
0f01Kao4skARB68zuE5wu3nj7Vwn5MvQdK3pHNxh0CEHmBMQHo9AHb7IetrtUVSts3NEFrQ6GnLm
MWH0fCpDfP8L+aYqm/fW8j9DikcHODnvHW92On18LSydydPqarFL6/fxQM4G7ABlLj8lXlIHdNA6
bIrSRtSq+MofCdiA3M5+M/A/mDw0YdIy2vwHKsNZ1ZS+dewYe6lWRJ4lUN6rurdTK0qWNvrZBv1P
PgnPNLfonluc5LUgXdLKv2lu/KgmDOg0LMi4Mwetkaat5Y4Yp3BGCa5CSsSqSQeU5S11sXExAchP
f/J10WmU/0F4hExojbCznwd5C/cNVEL+hrftm2zMEnEb6t+6PlvblSKEyGmGpEmeC6sTNsnMcXMX
pZPl//QXzUUEjrJHOunDKAX4PBY29/ckpz2QyXsp+D5Gq/utg/3VMvl0521n5bcBvSnFgaqz+yIF
ElI6OVjsSwAA2ecRT2b4A+1iGxYPqsMbFjvpR7HIcZyzxMYeWEAi50FbcGLx1oIRkxqTqqhQIIrQ
VpdbZeYqcZXR0rRReUvIUdCWWxkd3VQq5GRXScCd6i0HN4WYFUYHbhXJM10HqlmUdJjtrJk1J1IA
rjpFNMFUwN5vItpzo75Z5g+xSlxvYj0SsVyI8dp/NJTMspf93Xz983RJVZfVFw1hCd9Vwue1wg//
KDj3KS8WeGDKtzTPEXfW8GkoS6aPNaYuorM5DjSe7GCrb8rpB93JL8vju4MOlNHuPe3O4KBTAduY
dNRNFpxAV+a+xhLc8RU4zEh+/pC7KHXFZymr3RM7bMYsDb2FydCjzKBrLbiO/2hVl60IKfomeNp9
fR0EbTnG07LK3rpn5Ld38mXFmygoijwlbs9NQ2qQaxVRrGvzbKhUsgABSlqJppd/S5zdH6Eubb6Y
z5kEcewls2CVTnuRZnwqWg9IzgkLYcxE5Y4+z5pHWuEL14vH9vA9Jk4EH49D+ZmDa9XIFGHFGeT3
6puh45V6m0wZlpBW7P4sBJz8bNFM/4xpSUVWc4VhLt0iRjy+rN+XOl9mIcipLPw1y5/+h85PN4V3
HjlD4bVmSBHB+aEDU15xV+avMf2dUAHpkl1IbVUp+zoJpFW0CoaHqh/2ZE//Lu7MKh7bQT7JSF2P
9Mgtw5jIarl+dqhF1THPeUKsuv1hZgPqmYD6hkESEEnEf+84CrjaoIRsWY39OHuerW3C8Xr3IyQg
NltfFie+1MklnYcHD+nbLU8H8CDIEM6SvXYz0EmwpbEu681wlq84ma0Al+YUqpkgibWSlwk2IcxU
t5AuhFFpy20rLIJkIX0/e81V6E68m5s0SOxegIahyn2mLUwX7Wt0/9yVhxt0pjFJXbGe2pa9F3b+
fwFzYwoUWZ+g+ddMRH74BPSzQarZs/FWjGX9pqg1aBuV7jjv0p/zsPQtD8zS1phjPYQoH9Kpjl+Q
Va4mnqawDPbM3tIqJUHZIYMU81uJj9n1bRgbUaqgsvu4cZPVq5ZDpwMW1kvzCVtFlucrGRMvqmy7
MWqVei4XYvqqbYH14JQW0cZ2/PmCeS0i28bEdYAXKhncMwPNDuJj3lNNG6bb3aimtjur6UA0TDbs
skwEBgZUx7bDwMxXWbXiOgI6ElxdEYdo9m2UfRv5xcTeXiE+3/46BOq4kRXF6ja5lMsSwTZWuZxn
dzfG++dEBNv2ZVHo604ItINKs/4+dA4P3uzVnhsY25+2rV+4Cu5MaETXUDw8BnwmgfiVTxZH/nZr
MRfhXQyKZ4VzkDpZifpSHJUNhbRbYx381+pTjtpLZxmGEbb8UmaDlr7jJQhh/OltGcmuT1lStcDj
E4moam4zCGxQozDJrIye4SLHFRvwz2lH9IIctXdMaYtEpcyQsX7jHYG7y45T3l2DGY2YD5q4SRYZ
kVSU5g7dMm21RjOSWgFJ6LDfHjVo2e6UW3sc1aAR8pQQJZ3Xl1Umy3jzo7oyswWVDBp4t5OJIXoV
5RN42l3rH9vKpW7Xmv8+2JK/hdwcQzgom0H2j5Du1hQYZUatDq3kC5wwthHZFrxJkZB5YZfKrUE+
0RgZRfSwH5Bwtoqcqzh8+r5dRrtqhTupU1XlCtcoFr9+6sF3xL4uPfj0Bm6II+dWCA/nUE2p1JVd
HvapW1QAmi2+F+NuBNwY3lUNgPativVwdTrYwahIzQnV4P5deN31YqCUVdp32AnCulH7/ULneLxm
mZtg4WGrtx+y7B8kZSD98nOETXcNiBVu+iI1h0aJVoPPPtQ2MiGmgmPwPBcLwdCoa3+Ee8xaEGL2
xMBNmHDC9KWcnY0tAEskPIDgmhHfP4FChDhKZpdi0YSP3HO/ekFbp7DFqLFTGntArJlkTQZLF8jM
IwihLf/TCIusDk+MBNLdC7WeqyTtu5gpzhn1zCZNsaHfBj/Xj2vowkOh/YMjd0Eeghb8ZLpOqWP2
H2qt+D9+2dnkVACHsCgIgrZrEFKEJA1LakXopC8rN9QQ0Vz/+n+RVqAcEvonKF6ka/U9B5iNR5T0
kSP3yywG0vpIEpqF8Yw8hh1x1fLmlUPd3v+d7SpKnllsm/r7+kpTcL2sHefVVKxrF6yNAhovBuH8
I6+GPIWD2E37RFtfGULuwEScgZIUaoI5oUXuoC1dEE/Wb5bEdHsoJ5geuGCXtCNi4ACSfXFIJNUb
jIdXqgeFmfAM+sNAcI/df1tufB/S0+f7/9GBy8CqN6jM8Op/SoOIgCLwGfqW2fpjOjBhQGV+tX/y
PUFgkKW4naGly+xy9SuISohk9UBpQpovrRBDJNSfMRk6A3AqdQpBp4yk5lFYu6TrfG12y2oR1RUL
T7hTPbkHuW+uKSlGdw1Rjz/76PxILSddqtg9+d+Rs4hgYp6SGMu2iNeHjE8Ho8Fzm7LG38xMbJ3T
4kaEaNY9/s9XdqgQmSymbN+iH6Mfp38xXskIX1z5S6go7ZNQ2FfA1Fj/Jigk81j1/WM6HlYssbTB
FZLU35yXKRMReH1LNzKmaUhBMDAfL3kEWUs8KU3kwJF20YPkFrTJRvHo/HwFIHes1Bmh9IG5ldqv
ac37DGKhmdjcN264CEJNmtvFNzusq14hBPq07iPgUKI2P1217tX3HZ+d4ikn2L0Y+pa0YVlUMwGw
IQviMcyyMwCdUX2/zpRS+JJeFJ8d5oG0IhOFx4W6LrCMxNWXkeioAmJPh22mkkfs1MZQd/H7OxhS
Dp/NvjsYfvU8JKtfvcxhdlCxbYizz8ece7kghPiunfOq8OjeG9RzkxxzjPaKWsL1dduErBMXfZLV
OPljKFtrAWnSHpOrgZcLgoW6FMmBOhR5LSIy4L9jN/vUONjPzF50REBlxCLDqN/GwPxbY7Y9hWBN
n3dvrsWCRhvfqDilybPkTdI1Ms6NTQhdx+Zola3apdFirz6TzvhFgE8ok7nM/JrzHOPqLDxDbv8G
SQ7QfJV0pfywJAqppC1XcMDF43gCs3pd7qozhgNxE2lvZKTzosWC2oBkLCGszM5ZEYXVQq0tL5YT
sd3vTN9BiZejWR2pXjXCb1i5ieKpXruRODxMZg0SqgV4rq60eArdmgStfFdrAgX4DuWTN4SqVsm/
gcMSuDrZcFcPygL/L5VcTVOYhxRoY2miMZReqjniqW5ALRJ2qq4lj1UrGurpI0rZS7nGif4pbQYb
zLXXrP9bNszCXjo6Wj2qLDgSUJunJpTX4+srBn94TVercit34n7xjJUiHhw+wVvkPyUn59mm9uX+
UutszODTIgzFPEjcGNmTMYY7QkAfuME4h2gqnFJrZ+xVQUpFb2xp4djjjgdMvyXXjDX2OyiOhvsB
9W+Yn56Oyofq4QXot1kqPjd9j21TD/l+M0mp96nUIOPqnrM10LlmvNpIenuLAzM7eAE61uR9Jzlf
wnTzeIN1/TbCIbyiPBXplJM7s+mkaqAH9IrFvbc6pGSR0IMg7TAekoVVbTfMIwUFhFnPwianbvka
LPBbmDK1KYcV1g8FBYVapjid82ts7T5c5ayEI4fyjdMyZs7X1Ayy7ZEB/RlkPctMTyOK+7WA+otb
kaXndRW9SQHDZgm3e0yEq2iyLiUdmDw8C7+FvGW5MJcFjGzqoWF8YGHw4Eg5e2KdxDor7kZn8QNx
qTwY1dZOUnu710YIh5I8br1c8LJ2gTcITXVUOJvthlxgDKP2A6Tp8ORNt2ngn77PLgUS1uoGO/6h
k8naC8FTNv3NJR5lco3z1jdiWWwTOEkVy0SXSnyg6zMF5I/jHJseSx3I2Plo555I8o4+uax4KYe1
4WAlTFv+tNY28t9T0flZI9oLcAxxED0qRWvCdqL+NitO4bZ2ncvnBRIQi/5xkg9Xaj+2opg++rr7
R+f371WXvzfuUoqn9bhVj9KlgGCc8uNSZVltrlUGg8aTkBx8k9J3TdBYy9/Vobo9Wb+FBoCkAR+I
OnmeASpEr5h+9Zw3qzn8vPB+fMAPJFiomqT04mbBCnjJzvJMmO7eEsgqR0H81f9ZcW5eiSKsdpME
kMvAs3wNXkHm0uts1kQNo18xijjs2fCb3h6QUYAvyX7+zKJF9B+i5UN+C1Leo8RMTEyFrWh/jNb7
QLdJ4/SSypFLJ00XWZPaipSbjFBkuQD10w3+Fdt5OOp4y2E9hSgdylkw/Zq0BHtYmGAwcHKHttSE
HAKDSsBPX2Il8C+wTnK9iakLC/HgXYlCOJyyi25z+SqzztaCbJripdWdRjkpt3H4yTS/ZLFQRVQz
rWkSN4Cl8zJ9mzKJeFuaKiUG+v2hwQDgjdvoz6DyBm8HPaSteB7H0YOtDmLpQux8xxLTetszBWBK
cGtIpmlBbhs6RGCmTaw9GcZOlaIsBotvh5vI2RKQfuHo9XbC/Hnn929RpX0CR6zz2KOC56fmt9B0
iPeSJJarxtnCCs0dVMwwyoE5hRxVRh7oStx5/P22MV2rZsFMgUkFZxmFKVVwdbXNbSN4anV8Bo/T
WTKs7SBGD5pqJrw7I78Hw8sLATaFAzQOQDjbubIIiYnzRlpCnsOYAyJAS3qGrXReZXXqenroKwu6
xVHW0QzXBV9/qqv6Ws0rYhxhDO15LCwJFw4S05JN4eh3VUVc/OxNOGgnMkhrc9N5GgFeK+5WPlwM
5TWcOYdbauE32tqlKO8b02Is9qAglL9QSwdGgcgVLETxo4jBqSEGz+neHckSg55p/V8n4yGI5oVs
P1abjkxUVQyI+BE08wUyOo5Gw6ni2JLaKbnmujbu+wzMMIXZ0lbBZhmX/qQQpVzhtNc1rPW/nhfn
Jw9cCuYNdMon8sFRZPa/3nKHNbBtr590Yh2IQ/8gHS/kQwVCPl5dgZfat4v/i6ievTRqp7hzd6AZ
PMvuwyF+jkNvYMW72LDn+zHrJMVQyH4ukLW8dQuKoNmbRhY4/sOJWWjp7T6z9JTXp6YaEsqs3TKo
WWV9auRrOaE/2wqzs7T5n+qPB3LpBJJ7t1dwKERrI4/zf9MlLwqBO2aGB0MMSOVgZUVSDmZGipfe
QFav1GV+7FGGOFsT/4AoIzgvtU/RCCKgMW3EB5V/aENZUaYUBRdlIt+mv93/OzqH3TBAM9CjTlpX
CemQGqYNbDu5lez6u2shEKc7KgiHhiVb4eMPgqiV9yY8WIe2KqnRbuT83cb7FDhLcBtEaFY3+1Tc
dgJpOEuONCoq7lXNaYvkRDUTwkOVfkPuTlw0tHLqVHkz1dzX7RsSMmZHtlNdgR4fCk3+BrAUDRa5
Wdy87CyZExIfOw7COLRys32wmA1oaePqCyGisetv7ObJyCWeaVBp2ItDbjrGn9mg/KVyGILoobf5
nJNCOGeJzSislrtoWhi8jyMfFHf0dLQyMSThOt5Zt20FXxfaNEK8BH/8AMPS7xxxyTsioDMXAf08
hvyNbdFLrmb6AACEdyhZew2NWVa1wigWLDsiDGRUKBp15mAjn5aolNpgh+pflLjJbHok4Jlbkm51
HynJ6AqJGlx4zgMKrLqbocGSvyj9ZumreUpO0uH3rVjDjrdyBGGxl32nfo8tJkRT1MgTG/c61SEz
2Zh4Zs7aZIhFLZUNlMGEkGXdRuHTQkzwm2J8rN1rLLTWD7GNvIj4Kjklp8Sxktk7d1+MCtd/Jz1o
bvpAAhQXbwv1rcgFNNxlLaGlZUw+ZjQZHRdDOqkhCtjZfh1pYrB+B5pXSwOkMHKAD+vpuSEimbSQ
3RnusZJk2cF5fW3i8fKMv6N50Kl5XmNKpF8swsHLW5qmV17bZwbEt6PboE/U/5X93ch8FSUr8XtK
7XQarJjIDmH6E74VnQbs7n/3IhAgOqj+8b6nxABxno1OElkGBdrXzdOdkGvIRHifEjBAev48pHy2
OGE/PwYdNeVX8qaAhuWNZc3nE0cFcSVwEri7jmkHhcexHB/FYbK3rYdZzQKeTzDtGRi7YAh0EP1x
dpkMXYQFTscsCgPBwq9woG4RqCnE/cl8mPSKij4jrjMrhr29SYUh4UsgAVvWcTt6ewlM2nCfVBah
sK9j0kDyhi9AAh9colGND04nDMWh0Cq6rsYItIZqR3WkYaMn4rBPw8AL/ahoVcL78OIrSRkHwIqP
I6gvmIU2RVqCJk0NQK5i3071uddsvQkSUeQOT4e3CONeoINyDtSes8yAEBLm9GrAwyzh+rbK0fZt
5BGvehwXduADaG4t97yKZ1p1MMWoyd0AaQWGZp3voegp0mr5ukc1hPmpi9QjTsgbMWTlfuNh5OKL
OE3tdbnbmsb47rinuFH80HWxYXVairM4C4oKm2qN18LM+iqLW0cMZyVUCXnNVMyItQUqawmZcMh1
ELx9cGOH+zOtsUkTA0lJO7TA877LufPkns1XAXMud9AItEhsIz0We+WgoHsY5DzBM+ftaTxvaK5r
xaTmBzB+Gx1FgwK7cylf6LiA7v0N1IZ50t2U8ma9z++xddtNfvixGg8D+1Q69YC7+ejMsTiNCvJ8
kPtnr5RCRbcAu5Fo5Xz1YAbObWFps0CbBPzhe+KFUEcSCiEtavR0Z6CsRdceASRV/hQvlzPe7Rtc
Uky47Ks0wtSFBy1hlERCjtYoLev+qptSUrlIHKU8yCr9xfSsEOMeOnPzut0ncKynpbwf84if6M4z
fJ732UdzT2Z70+EH1JOXST82vCjNgTu38xdgklFjdtmbnOQgyZfl6b/fUEztbv5ODw15Pl/aMe6m
V5eet2tY/qNnWfOBvFqugHYBAGFIKrQMHAMeGdNjYdcEMlAXbkCjn3xhpYi9evXuQWy8oBlXcK1Z
dnWZtFHfJp8i5AsSc12WnLw4j9LsraFU34oyIgOr1HhKLaajBXLJ3g3i1N7NlQD7Bo67o7gGJ45Q
YYOBLX48xzy6eFDXEHFtsG+2p9te6X98+Miks+3Ja+2/y28mrVV2MeYnFWcH71cwbohd1gb8zUNk
DNprVTDwSv1v/fS37ezMUAEIsJ5zlsZDZKkeMiDXE1XlPNEO5O+TtyFEI2S5ug79Rc0h6r0KF3d4
31D568GIZTJvawz8MkKV0+31a+Qs06uNjZdNraisuuGTBegX5Yo6vC2TDCEIQgUyptH0nbKozfow
h0E0sqmjEHCBCe34gpu67ogf/c7NkZPjtvybLw5uKvPXfCwsQc5N7h34GuOhG5bnPzMpngknNtXQ
6TtNSGQxvYp27+urC5Wy/eI71nELFZbOYhPP8BVQTTOt10Jgn0TTJJOQvZFw6UZ8ZUO+cgyZdmMd
Jw15+BqVQwTbQi9iUgpcz4Xn3EcM9pH7eSZgEA3qO3cq3mQLhRkY8Mn+YlZ1MDVmLP9DncRnvGpY
E/ik07mVby+NEj/o8u/99InjupCg6DW5+/aL1W0OOiv3GHEC9EZei9ZCtO+ZHp9l/hzsU730ZkuP
wpSzaFY8Otp/pgBzJJD8GI9/h6pldsHc7RAE68L+nF0ZYeEPq1G6J/epIfTtRoTYKiVo37WzXc+p
eRFHDKz9r6KzdFdhU69s5/A2ZGcduGmS+aHH9fawmf6p8nGV1HxjS89YiR+wzm8Af0+etmz+yRfq
gCBmj2eEQ0lkHngU94RzP4g/c2X9H4JNLtGgkdOIP6pmWiteZg5fmxy0S1naOV8C+bxtVjQHg300
gxpzEc6QZX1d3cfkhawdtS4o1Ehd1Jy8kUsrdCcnv81OmuEBlcI+siIl441m+1jUt7oCpDSOcGlw
UVVBcooB5/X/pNOQLIxrguBOjhxAAOd3KXXP0MPE+vXfHBKxv5XPRwVBnPHOxRNE/5dKuDS6fUoU
SPg849k7h+0NwAmRdM2vjjKE7FZnBLi9mI0fhhlCwHXPQqy0bltrmTAMqdMjD+N4J5vpeFQtv5ef
2urcN7GYC1F9b080A/1vJw6q5aLTMvqfexM5eZQ2mTQ/qdgOVm0zG87pZIJKaWeIqv5zehDDO+l7
ZMoyaG/yONWWK2cJUGPylefSlJrE4MBVvOCwTbz+hH+VWkXqvPFEyzOKmIHQyG24trOS6ybsaAP8
DjuSUIILx/d/xt2zjikbqJDPqwgZbsh+vc1FnvAmueCx8G/refC7/HiSfN2wS8k8q5DcvfIMIuxW
w3souAntiTK4V2T2tGd0KoDMFudCQj53Awi3WQ/iucsvlxaPe81yGo2bJezEMjACwuFBN0pVhPo7
1MY87ja4pSrj+zf+G1yz8753Pu4rAyeWr7G8cDV9W3UkFp+9gSY7OqDMKJb0A9elafs4O0MDPpRK
phUY00v0k32Eiqa+OTGpuZh0JzoYfq9Tz7NYeMNAtkbiQL4Q2JfOnZxUj9RRQc2pYHD0siAzkI71
AVwUmPxx34lPy04kjEOUlzqaMWjwRE3HqJln+DVOQJ+zwMZxtlTPGBC91YkTWyCxAq3QnvEG0LcU
WLtLYRP/pGyuqzjbQL2oXDYm+bsBeaNpyos+gFEA8uMjiSR+2Lx45QQ7W01XBwbeHCNir61jCkrX
cBaxFdFudkGRVc1vg83bAGatLfD/WkU4GbDttMCaX+KuswEzXH//58dl3dtvGdortSskY/8F87Ub
xLFq6c7lfK3NkpASnWpgKiFVSXR+YxJQkOt1TiVB/g96lMqB9NEYzropGGbAg6CFTH1Fd0yWv2qy
m/X4MOYjhR5B1yuSiDnTc3D01XfmUSBcS9+O4vR3HfPG3/sjKQNW0GYNO1lo0L0AOfj57gmpiX/m
ESvRnWmFHKArB3vCXtzNtJsMqm842rWKaF7ourQkS7rFoCuOuhpsGXAi8XVMhP2Y8tCHbBrlv/Ju
s0xJBcAOEkMiVyIeM3rTVGRtdhQm9KaE9iINvSmAcDa1k2mJsrhyYaBMHiffalb2+dXa3M1u3hU+
bXtDEr5XwRFfjZpUgvYmN4INQONx9fdix3KQp3zfSoPD0YU1GdufEI9cIEIMNep86AzwyNG2LP1E
k0kKpJtP7FM32sPoOkI/4ZSRWSIVOfYg7qpFloPi1CklwOEWe3VlCf2QeahWyV18ledkR6NsYv+q
edZQF9ShnJvvlkwaLKvLCi69/14mXp7qRf/mcZr0LlPrSOgHPGp958JzO15q0Vl9u2Lni9jecd6l
9gvevWWAoeTcvp5DGokoWF6tMVcBBn0kocsSDN7iMCG2bRbzItQgZQH0S3XUDWEKJzdEa4BRZTal
fFqGMfxFk3YJv+O9psrZ8FMbRlN4OHvcZXkVUpUCGdw2oiWTnu388nP5qMxgO3U3h5U8Mt+n9hfo
N7kupn8PcmHSp90RMH5Hby/KoacxhLU21UmTV064mEXfCmr/Pu4AhF2+kBj8yJzJXAqXTXBiURNp
T663NAgV2D/TxHDWO12kV+3IaPK0Xx5g6x4pInOaBq2YN7d+hSot2PDEx8xoX77z+SdwbgWkiNo0
3zAnz/+rVrqAiUlsSd8Gv8E3MjvIQxFtzfLaqlRATCVZrpQdPcHCS3NkjeHpGhqWIOYVGznfRfO6
tOduGA6yma6AALTay4D08df21CYIa6r8kNhD91Rgb+hqDlm5Ah+G68LyVRUqBIFdf0bQUDyGw9b8
FLHjCHlQGJ3p+4ouDj7Aag8/FCTlU+837IsAho05WKGvPot3skg4Xo303kZ3lEyCkb+iYo41r0Aq
N1YFaVdcW6DKkZE/aQIb4I3fuIVgIvuDgyDKpjKXQFGADezUpr6WyZvBciL8RA+sOntmqW0nZ+7Z
hogNSLNi66N+wmSMZoU/r4lL4v6JqAWuQoYEOJC1g457TzLzNkQDxTUhYADn22nInR1qBG+3LcIn
j006aHr/Cc8wXQ/O9bWS1htObSI0H24WUI4+RoaTYsqyJ9G5aNb+rL1Hsjp6SclW4D6feveLrRJl
aMfFhoZrJ05Y4vAgy9RFP2D1mMTtpLSLrAUUjwSFd0d6AECaZ00sYjr35WI7vebKOK/0M5nqOFu4
bXVWPlNNm4nZxEPBj6ICe0VQ5IVC/PptDsmgbz6abwVKYg+SR85GqS9gjmja3oXxbepFUdNBqrGQ
EU7yyOxQILKqdjMx6nCg2dGlIdre1ywLMP6iXxx6pAAA+J/V7cF+p9mGvZbVQqCtU7GNtWOTYLah
ZGu3QiGOSAs4S33u9ce4QsmQY+N2fHy9q9QwqdVrFQLWwAtBURJwlsMvhxJfBpfCLyX1eJE7d0Dz
8azq/zGmWvpHUudnmbbndAVgMxVQMzDiwcMJmgO2d4DiPqV2gOxLcittwZZd9LqW0yVr7fgr5IF9
5GsZDaC8JmuI2ZgSgvRNBJL53zhMJQ1HZfTjR8xcp4KrBSTMC4FTPFxRDT8SZzSGPeIi985q3KY0
+pTIXn7GEujfT6HTGKK4F1QBGRxol5Q+4e812gMbZJryWfjgOu4XAuyEfUNCCXLGCorDRFrUS5Oe
Vnqh+DrzfT3TvsoQoSMZj+zzDdEwfukmv9Tai5D+Av9e9aE9+3ZM4S9tIIvkr0pKk+4ZQEukfFKi
QugQWToQtj/Z4ZVinU0e31NV8rBg++hA8a2wHX+4JiFNoe546HoQI98ZQBKR13yf2ORMQ3R46Aww
e2tUjE9BCQfJYPyOcjR1H18JUhxCuiaw4v7NdA3uibB1SOi/FsNc6kmFw4Lhf4Ypfo4NBvGaGISd
BihHlCWuyORm/qBkszkUDjYwlQgG0Y94LUn4DJj7kvLNqOCWHHgklHC/r3WcQGdjlq31tckB4cOo
7HCCmSGLhM4CP68FpnGg9r6jVigFBPAPTLbfN589GJUek9s6by6JWEjszyl0HsaXukxkNIWIWys3
2NCs6f269g2MDcaegm2wJfm3dEUYgTwL6QzJzEEbBXvqbvNf7HTix+pYI/E0FipmjRoj5wfkONiq
9W9ryx6G+SHbt6TcqYMPEVoapGBt79YhfMgi5FYglebP+MIks7mM0DfRRBxKD7oqtRDkq0xogo0P
ugWvUzLYyliKMPMjYLInsynnqyP7PM9jNLW7U7ntLIEjqOAY4a2lzPL+mbDE79J4lp8orw0hGbsI
K4lGIWsMwYYrJoAFqhMNP/7hGddwBKgJEhg8Pl4hU6ODCo2noMxUh1lhxRQk7WuV7ucp4yf7q0/l
nI9xA6U95hHdbRJQGqX7mpWUiWDJMJwStdYWSqWNVMVvl2xTZLihElLUfxVDwVsTkVpKtrq3U3mN
yp267RveVGTcr8iWsWgtV/MMCqhPbdhxTkVC0bwdW3dvN5ipsNVSo/Yc2HSqO6sLlJD3c27dPUZP
uEVBlxnHBFXEG83MyZcAEeyCg+lhEhByW2dFSt3qDvcZyQfDy7+/6dxlCDzmZXtB/IkIUjV4r9H4
YKlYX9qqUYreFPwhacbtjYfLGUKTsVKj+KaqCNTjZJmgjT4PXo4Oa7yvxc0qs/h3xS1q2CgwBD4c
k2cev8hy0bWcaZzGwggnXA5laaENL2U6neEFeQgyd9uC8/wNvXwHGMvyrH8vL5jyoF2Luh5N9Fys
HQwaMpL1PoOEc1I7DQv+L2M7t3NId2tZ4XmzemDk5dgUDAT4QakPfZnb/uDFW9S0KqD3Ais7bVWT
J4CxQwv4wUvjr0zZtuy5VybvmgxMNI9gPT2R2qTWdw0ZjNqpzurBz/mizFuLpWuFrmTABAC3cNIZ
PY8uWsqvDXOr7hKH+nU7g6p0ZZ0lmg5VC7oyMOR4odUkArXdCpGTfi5fmCwlna3UStc9EAHPHFn6
GqIsPQNgvnqby17XmXh3bg+le6iagLR33ngFkXefnJmf0IgF7IpxXaTMy65+iF6iVfv7/5ysbia+
NVy/Eg5I+q9pHBnO5AWGlw+qeb24gPsJp9HTP9c76QijYntoI1GlTqJ/iq4x14QF4tE8hR9ncsIL
u9mIld8Eyw7R1H/MLhW4WGA9SeeH3MKMS6Z+HzSBoIFmv2tp4Suh9puyvGwzPc5KgQxo+qKBBI1i
wS+MBVCKs2x6ZK8NpE5UcqRa/3JCpnoc/kyrCjeGoOtii54uCGpAuA61wHd3Z1Uy4OlyFPi7DA3j
J+LryPEfpnZQW26JJULcP8+ouPMceVv/Iim5+EAKEjI5SAj+m9md+u2XzQeSufo+JcaOP/LT6LEJ
TLGIdSEpovYrEBmbP29SV+1G0JhHcsSzLgj8In3lZKymgnOgNh7b6fJolSt1M0tLq1PJOr0UHsL+
2JVkDsDsa0vQZvN4KTr3kkAi2bpL+4mHKTDjt7Us+UnvkHiBwk2T/7NpDTk9w53rakgGsblOljak
zur5JFm7KlU6DfNGnkphxGIHtBVXfnc07ewuxc5BVmI4lHpxHAr+yXYkBO6aRxXAD0SPr3Tp7o1c
tgk0T+Y27bUbFWboYw2RKxbLBBsw96Dex4/PvwsWpDzmhQ+h0y6qmKElJLssze+bHXvv2jLNcQ4u
x+wdphsM1YPUcNmjIwmVPsD3cKI2JLscgc6NQCObAkyC5s2BAsnkDmclAxR8R1912V4aJ+aKSuIH
2bg2zxyEzPgQ5HfPc5epdzwDLlUqqWaosO386WfQ6tdMx6lHRDjLHecNmqATQd1CKGPH7e+80hqS
1e1rtrU+qlaY01PTDc0zT595aQ5qRnjwimPSi8tqcjoxKV8LTRi3H+n3egZflfSb4yJ9ykEe2XC6
xTePBh2A5IMONS0A1ylPsxrcQH7STM730QMFsGfWcF/UsswIoHzrt3N4xMKGBe86YakkORNKHzCa
aGV7X7/WiwgVQdhd9hM3AncHto9FNXjIa5+LsoqGq+cO6tcsnaP4DR5rOweC/cSLusQ1eDvFAusx
ci1lnbRd/8OnoatP9mvoHb4XpMSpAulAzA4L16kOVrI1D8eQ7G/i6gFVlYkvlPubBQop2JkYP4Fy
5ds/wpqwJcDPMcqy60fykbb9Li9AXdSSszAEkNpE0LifCf9lh6LEh/Nlv5repjZ8XYq/yMex7uDP
gfByBzJG+EMWoxNtMnTjDQJ1o3s9Vczv3A2XW6dhw9U5D4PoJ8S2DVnkQZOSTCyy8DUUGJol+jR+
Vv2W4sY3JZfBTj+Hst2OdJzL9oj52b4OLtCcWk5TDJeX6BCXExD/gGawlM0KGyhJPTklmB3wdmtt
KzWvP8DSqkUZiak2BXeR5awTpfP06tXf2Q/MurTcY9mLsHf8PWJo7MbX2Hf0GeJfB77E7cQUdoxj
HhsYAAC8vqg3lAwzgM1QJ0uItWmVO6N0SrAhI1banZABP+98o0V3DUwkhG118YLaqGfgYdPjAjg7
P1k5FfzGj1Ml5wAXlD5dZsNmHGW9qVSMKz5djCOutt4wc2H1uFoWRdEP3+027EZbKJbqbddFwgEv
PYuAf5J6o7JWzRbAmiNyiYyAfZ73lQrmOnfarPQ3hAbnz6ib8h/sTjmdoLh/nr+G9R3OlLl/Ad5/
7M+bssZbs8epDAkBV/LWZptfkU4NTkgQiubO7AuiBOowy4IwnONX0oQ1pQfSJKZKatc52gbEQXBU
GW9PxzCF1bBddUy1nRiH99lWoUIJh5tDaN1PlEd80j9cG8bCzayPyD1PheL1MNYSd9BTf3ACUlEs
3jFfbEHQPGli30oPFIdIVkAXsSk178JGXtcyUZqVRpflZ3jnFbC22z/7LCyMVyuw9vTLquEjJR8C
FQ2ahK1QON+SOXAwkzwskYUi2rCjFMo22V/6B3KL3mU8eIGZ96MyrFxTLXkkg4mLKgcT7nXK9UCY
Hz2AJkC94Ukx1Xu3yVnVtHQvXBcYq8u4TykZlD1hxhwwD64xvH2+9CtS6NPettI27CRMJAmYCzLo
0rXfizRS1//bRu+68xzyF8LvIf1gnWhWG6k2fnL6Zb/Bo24bDDp0rwISbJepFbYq+T+UzUFzcdDN
Ck3Wx9qUHnqZgp2TPf/YQa//QliT0w8QuQldN0aKRYna4M3fjXbpmMyc9pUR6rkDdgdSs20XIVGf
KD2mYOGzTXSmKH94wKYVkXHCo0LyYIxLXB6LcsC2DUeM+mheJIP5AeFK4ZLXTLbKTAWKBnPYYXjC
k3p8SI4IGWw/WfU6PQKkZ9aTcZB+hKQJMvFcjtzBJaXoc8MIhEgBGIFzb20v5aanx6KYCHCb6PBM
MaF5oYXLv4PO/KrfRxjp/UzqLK/svz2YNHxegHiEMyfTRjFX/BqmKDH+SrevyvmRriLBlZMy+HTt
0kvKRC16EoQOjeKaClmkT9lzBDtlVBq+7LwWP6byw9ggzfuI7Qgh5iON//NlA6ySsh+VuXwhi06w
90L8587LiniScdbTeGk2ul24YMuTyjPdw9NflENBTXge1X3xnc7AfWcABL2iQhp9irkmXfPx8K7z
r5SJ+sEfR/VqGMavbmZ2vjjDOkS/hqc4rhnbfVh8ePuEga7czLrLLCxUgMgGFaOQ+h8V87gFyRA1
PYg8gyi13H6x1/Lbay1X5pCIZ+mP4R9sGlDqYaLIqu1Ep6MINpzml+oabeKydVbOujrGGV0Vdpxq
mYREMVNFC7rjQtTBOJd4iIhxInQF5rzbJSPzdzIiS5CSHY7HG92V3CE5NzYyp/WWh4oxFlK3vlWB
UwiIHnW7GgZR/VUFTHulycSOvU5JHER5ZuO8v4etkKCMZC4tx1SUsAa5tUdoemDrnbDfogE0jADZ
77o2GbGhnzefRymBazWbpDMF+yCIClq4fGOJKtYxfwmZfFDasOavJXcTDlzV66IIaJ0AeF+LVsng
OpqWP5j3jTrYqb5GPUCNFZZrZ2msxYUyn/WFuitYtDRerrkwVfpSVf4IaNQokLLyxqg3PyVYTPv+
UP285YUKKIpLI/HQeoMfT4cgbBIFdvgN99SKjBEBw9Xa9nMzHXbEcK4RJoQBLGypTrSPIle3vSSD
rD/3d/ykoVk9AuCp7yhpXz6ReszTisWfJdt36RHWM6awY4ZZBOgDc6MAusNZ1za6nS52b7O5yogo
81w6LaGEwmPlHu4ttar8xlYr+8nAwEE/U6DLfBkrDQ8W5dHzxnlwlwOeFfaiOR/5f3W5PowRGK8X
ItbQVqgT8IkylSrKj2OQmoFzeM69WVWnuKfRkWEhApWxWfg8GJ4lIozZ25qApVJO0ObGSNHFzC1a
6yZ/pPOvoiP2FuFOAqqLpgK5a1XsBkCECAdmSOpFyPIYFCwICUrPCbzOYjVL2uFeLtKSgHDIvhV4
LuglW/YbIwwXHH4fQhfMuvTK2nBTgxtWq+B1PQrKwpfVzmPi1ZibWwML/vSNlkilb3WzFCx8VjE8
pUDCZ/XL3v/ULSJ1/D5kP51NKRYDxBaDJcETCzUNqDDmGHD/+QbK2v7MdyKdScx5mQl7Q1I3j7CF
fri09N8bAWafBIR48oqemFoSrbQ73qnIvrWgDOg34Dr3bEz/nA7mgNBZnmIq3fjJLvQhMks8TMf8
L851li04GDsbB52Hvk24d7TEG1IuPaOkRpPWBqLRCtp51ckbkk3bSkbg1hL/a5Q0/6yTnr4cVi8A
Yt+NEH4ym6iVnhREOVqfJjsBAYQzu1FpoJagRkhyKIgeDN2Fl+1/7NG+LMCXkzr9uR9ay3npHTpd
BpOMzm35qQhHJ+g+Q2wIlAzoCaZU1d65R4GAY6X6vY8CkybN6S9FZ3jDFMrUzDZPUmhDTKoHZDKC
WeJaKVKbNp2GZAwHJHVeB7KOSYAsuDrqZhoRFxZTTCjtk2yiFdJRT8JUHgpUNgyeOhCwAgN48yWp
HW8hXMJu6meWkLkBDb2Uf5+QDzWBtG1vOIbri5RNaoV3N3QKixCm9XKn22s+iZCGhJLqF9jPC1e1
WS/pQna2eDoEyObDGSxpTqIY3OX2v3gFd6e4Gdo2Y2p1rvGAbefAaVqCW+Mbck7VUosAuTc5GenF
ycSWTMfrdczdxniKBjmjxqRsE4aWpGzXcc+tj7n7ToanVIrAb32o6dMwsT2eYGNOC5hpOHl4VNBJ
Ta5rK2rIURnb43hhZdEUG9DuTg/1K40kK9qpWrTxmIE4AnCBv7I3A7KaXytggoMSebvkCAEyqfwR
Tm9ff6mMIcySqqlNT6rS9ZMlIWBzBOIAkpx8TIejdcFfLFs7kWB318T08Tzckk+zFMAcqGLj/xMF
XzRMHh3vL9wCJ89allwrnsWxmLpUjiKAQ5YoAslQugvzthogAWIFaXiY7qBVijHktJEUhUW3y237
2grNGyBkD0ouAWfDFSnJLaqkrXbg+QlLD5TMI06R+ezxJkYweUWe1nf+RSfFoJ0KiHOTeK3KLGnx
Kcq1owGL/MlkShtekRhHsDiQDn63HcLRAdLOSmnuh2a8WWwixH0kjPRqkOEorVpwX8s6QvlmQzup
BN71wQdTyykBiVjgiYAF9FCVhwIvesCxwWen6RzLPlCQdCvrFRGgNBQDQK0vb7xLRDTWIZ7nVsSJ
YivAfNWYerNHWd4hDWLoe4nGAUnZC3Zn40sj+5nXl35tF9ZTpwey4IlFQJVqULPtFUXxboFOQ+v7
MVjUvheMKEmayqry37EKritfusq84u0Hrx2G/9xOHeO1FlJgsRNBazmWbw9Il37AsbSjjmXPp3+B
tmkAn66iqvca5EqP2bxcR7BDpoUxP/byPTA4TfxFFWbHka8gHTtOwG1FzLgkgh9t8geHDhH8B1Y1
A6CUmLBpuymeAVwbEIn0xTksaUryFhb19MaxDgtwbNat4Z4452AdM41CKEy3PfrmrQV+B27Uorq0
y4rNxgJwgxs7br9o+b42ml36OqkBcNdPaYhBbjUfpNoKXqEXXZsVIPAAe2rADG+/CV+1XztU5F1G
wae2stiu6HdqZbAMCmPs56QMoeUdj4tWrgMyQpkiYwBHiMdWig/TtXyHScLJTpknfGCEV4saSs4g
fr+vh8mkdSfH+73mv7kyGR7iJl1FaeuccuX/fvn4Rlt0YqTo+FUd9qv0oTKBd/Hcn2B5C1bD1tly
eYtw0zqxdaAONfgB7YfgmpJgBuKlZcuLrunrqjAp/oMcBMFL6jVfkF1rZbejDIEqmpW5PDahoJ6D
1Y8f1STYnKFpa5H4vtr2iTveXfLL/jnNuk1VYRJGMCbdbMv2fuWfnQdrsjRcwmGNOdHbRvEcduPj
6Y3YsVn7RnwX1q5hlD1kzfNg1Ka9m6dk3+0sK24RWdXNNql0OUVQDe3NUNbDQJi1xs2cKxYbYZaQ
hnvIxB6wrJImjr7JgMVjtQTjCHkRwGH6B5i58xmT+/P3PU5qksch+Xlwntz77Sw1yqImEClqhQ6o
rXV4pG9dwqKf4VGsXcUa+Qh1WciEoXpzMlAr78BKhx+vgKbzFx8ofhbo/CxXe8GyD3+fM0jPX+My
4OBMAQ3X207ieG3N0Fecmk3RqWvkxvvlJ5xD9Tzv2YSeHZAsZMLcY10s3cDodeqd+e4x4fTRpkry
FER97GD3ils5yHhEwF8uyxOd4Lv6GchxSj9o7Yp7mFQHgyTKkK7y7dOVO+L2idYhUAk67Q42qbJi
LdV59CfpsuNT6liV8Jy1nd3Xfk8g4wHkc2s31r1kADUnmd305egh3loUnkjwBlIMB8uVhuwwq3aq
KL6cZvh5zoMgVRaaHO/uL2L3QyLXZY8P/YdL1sKXyNQUsF6nI+FWoyX7KhFfQnOIXfVEGwyAAhQj
q7A1A8RKqFo0Tf2P8IZ+dZpSSGqXvO1CwuyDyHYAYizVP7cyvqeA/XpsT69RIl2N2uxuzQeM9k4F
Xs02ZgWrDqwTX1X1qZvuiavy50GsulvAv+8rM/yFi+MGiFTDMpi6Wun4ccyXNtSDwafiZXWpHkIx
X8fiO7MPGHCjJZxUJnPRRZJNEknA9cbA6P+28hJrg56dT9fGEC5K3H+mkBj6qcLfmphGXJeZr6aP
EUIdN0A49ORe1z9wO1NjIRp6rSCahIlm0U/ZIMl21Ri+RGZvGkYRxavnLR/DdlCGchnA/jUUFvq+
pLvfG5qHCHUIGWtmSbFYJ1GZciBgwfTUTQpGtkI4QVa9eL68pBjHyFve7IAVgZi0mrn0ywnoY+4A
FPRWZEG+JlRjP575BhqtefcwhXiLFNxkQYTHCa69/a+HdaQ7QbIZSlJs6KuNAEPmchbGjoiZ8e9o
kJJ2BtBkKOCdIOlu3lIKE0Kl3LNzdq1rIkZNiLUtOg+1kss5gyE9uXL/9kiRnQS5WyYU3tVFE6st
RmUaklgPTxrk8/HfVMss8KVdWzmcgKeAZNZk4+ZKxxMOCF21P79ovX5MLE54fwWXqT5bAcU/aL7c
y7fuPZoLdcIc5n2r8bZcDTPOdaQ7SWZ4rSFPbv7pJVA1/D0YJRjkvj2yrS+DCjm1R8hcagctYvnp
cQ47OFVEoDAydfuEAzSN72nfVPzZ9uPsIBoWvrzviI5Yy4BEwPSAG4NBOnLCLFbjFek3nTRk9QrD
v/T4lREUl/LdlxDHvocML4hm5qyLkygOWtsZdT5D5eTzH9xC+9T7Q8P1Z0S+3nWNNnpGeYW4enU2
r6b2cC91Q9U5t3iJfulQYnw2nY2XXsf3LColI3hhfOoNy3LL7cWleNUIkP/gHyhfvbuoZHcYB5jX
TRNQBKrPrOyvi6zKBsaR86yTouiXVGTVQIdeqQH5cZtzL5ScoSWqVALMwNCzGx8HtNUqVJGOdnTU
+q2vzS1kWD1RuNk2vNPuWAeF1CfTbkyZrGjjz+dC/6UvIRpNEqeQbJTqAut/V29gJjO+Yv+CsDO/
S26Upz8XG2+ZQOeHGKxw+bqmnX3PYLjO4vvWAtrnr69AOHLa9w4H8IizWs2Pv+v3zEeboQnDtzYl
4YptLLtEOgOHAaBWTFeYiSfk800mxU7+ht1T95i3rKPB8TDq4UE7fsxL7TtQbvW3hcoxUSwePu/t
z4UGEcJqoKTk96uhqgxi3dY0WG9vHW3Yade1WP9eeA0+wOljzbwrJpg07pe7Pjg9Q9JsNBnMtifT
3U/2IT4XVX8dkRgQbXd7cbOEKuhDxSgjMcFgqQNtbmZovsRAcQK3XUCfDb9HE7BSsAJmyVxqoBTZ
0X2VhJ8ZdXUHCITOpywOxqmBS4hZzNH9YZnGc3kqs+GYSLXxxw9OPJR/CxdiMbkr2mb8id614RzC
sY6kSrCZaWwb5h2tyysX2qZf7ZxYIjtBR+6pMomY6LN9mm84JV7k4Z9kKN6OsVoDhwyJla+nU+UY
vxzy9M0WNMcC0XcojnSkHUXSXJ/4fnkgEU2oalfPiyvxvT6HOeMOXAVBJJwrQILHyN7X664BUhJ7
uFsqdtZtf1X3p7a7j5lWNBo0phQ2pWWuhPxZh61XW0gJh+ik84+OCq8qa6bifCCLimqgKsNUZojC
Bo7Yc9G6E/98lL39wmzIJT2N0qGxDKVMcKRDntElvd6bw0Pn09/fswS+wTQZ8mPP9pLEdRN8DiAL
jCSVSxRyASW3RXGMFlm/xS+jqLtYIrRCq6vAnnqts8ASCNWQEI6rskfNxJrVEmPNAK42nDflHwcQ
VkLzBEWqTHbsLTlUdIUdvVb+6KWYtx5/SpdrRZ/Q4rk3CDyIb2N0yCKAWGAViUuTLKxF0Ov3HWcp
2C1PAVr6lTUrM0nhtJ96eIYaeDsOUAwh3iEUv04f5jiXazQmkBKkLmlTM6WouZUUUnULaQ8/AUFo
TW79qsQf590aj+ELiWTnzadixFA9lFxPUCUtXAQ9fTnRXZyMCyzbZGLOMglc/WGuMqQOT75iEpWm
ybrKyZwXiyloa1nxupAY7HLz4iHvZvsM3F2zh6nytdPHrI5aeofl6NlCfpxIBurMB5qbOF07+VcR
TuUjFmS8i19EGUWPEH8uw2+pB6WAUT8niNxH0PyTyIo+VqBOe/cqnIXRxsz0Bitw+iNbXlux0mfC
Q5WKeo5EN26GhDeMyBs9bgjm/nD3sItNj2X4kfD48MPokLqKye8GyUCIULrBkXocIGlTD639GFL8
/NLDi8tNEExJZWBXUVGMinRafqfdzEcPuQc95oFT/uMtP+8+u5AsUCFjgj/ga2HrpZyndl+6da6v
11Skg8zRWSmb4hrWDWfasE1DEVZt3bN0UMk1buAhYVmpGIMHDzcfsW1BjtNI6u6PNSr/K0H8C8Ja
fXeaXVSMd2ediBEGwx56vYpEEA0pg+UjURO+p8iBVvfYxf7d+vSPG+x/Kw+0D2lQKwhyqj+rvJfR
9W4UcEL5hnHaqpIEfR9w1vrSR7hzJHKasqitLCOiJso7Te/GZUOI8Q+U7SlPslWvr72mtuwZTmYu
kD/h68PHgImvSXcpNjzooqxZ8IkFSewns1S6nq7SeMVYSqtK3SxfV1LpgRTZQNJnoWK6v+3SnObT
X/YS3dWWHeSb9LwNH7SdfQADRBPAgaKgKYWgIFbtp2S6e+2gpyfLaYZeYiDElcmyciFwieu+r6Ka
IwoHxbqYu5OMkMqQ0by7MGCY2OihxI13vNnv63YlRWIA+Z5o/l/SVFZpZwJkSSJdxJG8X2igVKQ6
LnSB1dfLF2+YiDViXIrSa99zu2wHW/YwjY4UpSgihqufsty6F2OefNyC2xoK3c/C1Fc6rtIefoYb
KbX6CbMR2kvWJiHV0+hjGa0gK4nyd68Xe7KlTvyalyhkizaw0OEfD+i4vIWmuTWAtgmGA02fwjRc
TRUmnGnJWCiQdPL4BTeaOSNS0MbrpWc2uZV2fHKC95xMv2LEkTWVoXZzCF/eMGOoYi6f+k4mdrLS
DIivax8Z7UK06JyBPazWqUg5D469Uk02u9i4jVKY+KC/ZujC55hOzo2yqZ5DshwykBssDx6lkVya
s4Zn9HK867jui1bnCHx7iHwGcD4GNbk7VJNkaN0XAwF7hPNCRXk8wxHzfTJT9CXfWeaR3dJJI20p
nbwDE6RHdNkKKmvcwn8wpoddp5l+75q9XLdo4cKmzuXHYwYfmMOMY14e6cr0UsCb7jeAU1HUncDL
zYXAdhJ8k4ZqvoqvXClglEv7As1gFfj+L9MT5EIPO8CP2v4l5mw20hoj98+QaNJ1M40SaEWiHWOe
vx6/QQAhWvRZ+b1RRR7WUbHbWL0cEY/HFjYPb+9oR70+NcaZCggP6AbzqQTZ2exWO7BKTpOUA48/
BKn/ifJR4Cb8P+HSjbrrexlV5fdoK9d2TzW6fBEr9XMH2ejiJbn6xw4DTim1zytr958nH/WYZ0ar
c6dNXYL5Ff8rHgBzKKMJa2fW9KKGqP2ACS6Mlp4E2GfW+3WKkwNk0YzdoFXGpzFjf70COVOwVTdk
Zv4ggAf0YyG6FJrSI1KDyKIz1y4bzE/yCy3p03d/8XZBADMOHP4/0HuSGE5tTZwitsDLujgWa6Ru
enfRAWfj6jbpsBy1b/4L1ThKB2f3QklETXBzv+TohpEC39rtdeONdQIO5UF2aOVTPxYV+qkvmXne
0LC6K+vcZRBB6myyOK9VrbJRWEgIzl6INy+iqUF4/euDLd2P6K9zwGWe817Ql8DgiC+sUgvCOnaX
Xc7vfdIzddi05/QbobfE6Ef9rdZd1ujCJ9UGZ2cqvYhOL8LVRUs9ImEyzCNOFd6JP07RQbj4a065
qSZKNShJ7ImI6le7b/hVtMlyl1E/YuTio9vdS0fkXpk87Gc2zrGV2fGrhthJ4W6Ym5f8DKe4VBJp
XxYMqo5g9esIqnsZKbSlzuoSDzt1vaRwHN0DS6i1462nle8GZz/Z6Hwk+WCOFOe6ArLZYG8awW+c
D50eKfPoIGDq2MmjSCav1ur/PfuiTp8VnD0DS/r1Ehl3PgsLVCjhvgDvxYPASV9WNGbBWnMFJ/yq
aV35+DAMp0KflWPwHHQXGAgpMqq2qRqSN5Km2YzYIRwkHev3X3yfcSWgxGBb+TqMc5BfnfMm+ugH
Rtg1vEwzDL66SV4PGJP9yxxwLPQiDP7vzfW3Go6iVfRV6YdjAoZDasAHJaKNafq5Fw53eei3O78f
INaIL1rOXIJsWmrzylPnvynm9/3QWHA+Mar9GyACF3YS+FUqcfcRQ43CsDTdxdhUnl8ncuwSjgyY
IMwkicfDL4+A2s8o5PN3Ip67wlpt3QDhqv4rDdUhSFL1Mjmpcl3NTlt/TXUfE1xE6DAChHP9WJXK
1vUZxSGLYlbo8YBrlcq7d6xJSU0pwVnqWvlpYKI7LuOjdRoUrzaD85oaTvZYwSCjeSrZfFonJ6wK
VqNp2k/GbcbF3WZZ0+2JNT9jnDoWplZkRv3ebsD31/JQkmDq7p6WvH45DepXjHLhE6y1kSKDTV7S
nuRLwJ0n+QTjkA2HfqJnMOrcUcsuCj+alT7w6qTszr7I1bgqE/mZPeIZSkSd3WUfUdTxs/V5qwcp
qd9yF+nnb2mRAi6KlIrrb9mZz8Ye/JrNx1RQAGQYw/RCtOq0qQJ+dEE4I5TWK6ksYnxNRtOW155V
keUfGmDdHBNIItCvA7w2BKTR7/Jbix/7NQs145t1zJo+CTn9Uhto5x3flMIJgqNrAeDZFsg8FiNH
6frAVxxuMUC8vPdPqVnSZwfhGzXhIfPjoxhB9aIYc7npqW5BLwdIC3Ed21Q2lp6mp1MgpMBN3/UV
idvn54bNKh4kTyUJBBQo651AfRJp5FBnshIYYQPnIgK9ehwV24snnL+c5YE0WeOXo/iwhrQAV0ZE
NPogFT+88294xMxKyiMhtMdWBwSlTkAD4Afk6AC6Js5/XL8uxHNABTk5WuojarTnpiwuyKILRRU5
qOdS3d5Z4hoWDc5u+WNBIlCsKt7z+A7jBE3DU+hEqoMxq0J0EN4jgQlRLsdl+a/BJv9MvZoqLSWJ
mLlw5hiPDCW4zYLFAQ47Tmvf4095ZsCzkT0YV9uy0ekIZfCDAHRpCMEsPBve3BWYkmK79yGkoieD
0Wuh02XFTaDxw302CsQtTn+4mxqSJ2hZ+hQ13HDEI4tn0n+OruSS06FAnrMTuHpQbHXd0sS+s/jY
OiwTS8L7dZB2jbj0sWt6tnm0eENBAjvlakUNyYUDhxu11NFdjIJX/xWB3CJpkY8s9YKqlHDDVh6i
E5W+YQM6FHy8HVP033MkaAawWGVY56fhDbXyoezClSqvjeF5IsNH5cza3kdnIfmHH+/B/zaGsWPq
TEKiT13/vm9pfP4oNiMGVFAyhW5Lzl/wDqpyaO4AmSjD56ENO7wIK5Qc0qgMfQOK7txZ2hhGKibf
mr+iJVObsrC0ImgYnMVoiaeDGOzuUk5hs9hSiWx320rL24IzOZHODP1XwMPJWEL4ZsyrQeW8mbmc
49qRF53Rx7fvXLfJ2ZfPO9KSy9Erq9Ur73RI+9MhA29yL+Ff3Q9qwjTd0MGc8bKbOd5LF+h2Yhjb
legvMEjEn4XE7DgPwkeoh3OIQ8AbtOGNTc8PaP2fghyDjVPDq6/FPHgufmbKo7uS3NZAwgYuT4Ax
2jVkVg1wgpVGl8dNifchu6mp3g2/Wot1+f//QsSCVXObm6E4CKi40zEyrg8P+DDihUJnqAxpqkk4
2Tq1TzGYG6glBB7oQhbQqGKUoZBpstxQqAJdwBaDGU6lbQmhS+QhtXEhQ/i67BPz1tBqLfD99AbN
wtxVx3ZhS7/bSl3G7qeVXGnoUa5G36YtP5KyYeGjlCL5GAygGQx0t3gFoU3ienr/2aMzX/5UU6xm
XvwbxPfxhrXVWLn7a6C5Jva1R1nLtT1YgfEh9W96wKYJcPeyNAvwEbaQgXRAFGuVy0M5y+0y6n2R
RKL+nseCby73/Ms9zZaUGOAMBmV7kWG7Nzfe9gd26iY8u2zc9LlC5uPd1AKnbm5pPJ68dQTbZZP4
9dZZ5qXy53LYkXiu2kCOUmx3jtUVe8OrD9AoHSkVJpFE/d/grdNaO1R+pM5B4YLTFg9WWkMf3bIC
23s4dKgJpH6HnjdRkhM9gupvFSe0bXDotI9WExPIYmN/8RhU77Z+TXOyiUPaZEA86k7YkrSZIRxj
OLjT/gbxblcFzpJ73/BkR5qgKqo8jxyYBvKnmmwnMVDLZhtBUxE0osaTeDXW10+c5DCxYcfVf+Fz
PI2UxWXBCL10IZyt7tb5yASmzMGcB52NqmxBe5VgENvMCSFqc0fqT+0kT/uEVZbrtSC5JawpIU0d
eDxI+1pa+h/Jbz+vyg8Mo6+68VkppBNmRTCctjtNa3ggiWEFqLWZsN/qIukEzFZy2rw79GycdHmk
2tS2hlCE95PAN62eH1G4eCJwQRUOdVixmyqhB6xvN5vPOS1pu76tCbhOA/anTbeGj+Bz46jW4b5N
s6Lz/Bxy9//XTBiMAlyyRABuFY+F2fu2BQGERChk+IqEKPUZcP5ZaVbySEXRK043hXC8CbFzqxBE
hQ7uxhCqISn5Q220Dc+44CYIBom6bKsXaNhi9XeQbNYNx37+8PTPLYqqxsO7cN9oDFc0IHjkMV+H
50zg6DhFDF+g0qElOtqeva7n9F+AJkraak6hLtIviQGdiYerMMfSleB/Kc+S0/8YoW236ShprcsB
wGqtLXz5DlDmuKztGpxY3p3psgJKYJ2sPIF7xJ3qw77LoVuM0qypiVYDOk0pgp5XkNPpx7T6RYVW
EMdkKwZf7gVCq74Gf8L/DfI7kw8dICqpd4fzwXRJoaM/DKPEOSt6XdcOmOXkAKWfKccxTbxEquvo
brmVcxVD2mOXECFVkQDGw70Rq+DPws2YsQdrErwAkcbvZAbVwknhzsp41thw4riYHlbbDkDrXUFc
7xZzSAiuUZ5V+j7165ADVPrcahADcKXrqagftD9kOzTZIxYVoDLMr3TowjqoSR/4Q1XtcdqtuNzN
wXZM1DktRptiy4ZnpcPalMPmABBboJ5pnORU2nK+Ks1B51THRUAovKL/xQOOe1Wxzs1jQmsOjFHO
OhP7Hh1PoNiY3dJpGcE9V/F51OYE29Z9kO0aaFD68RPTFqYukRJymvKJ3zTbR44CGnDPP+Xo8nF3
4CznPAp/8cElljWoJNLVoNJLRnNTYIo57WkAdwfQLOsbyOPZs1fqWrqS5LUvisYRD/szIvoUmd6o
WARufLI4Q5KAbSJdT5QoRfpd04jtJdad6yAjhiZxL8lFrrsj00rlPAtxro1tCXXyJwDRmcaRcSHp
phsS73Suv50x5yeVBEADwAv1YG56hg3PKkha5mPxmDEN7NzdOz9FxzJlJVNvog65gQN46gqHdKXm
vXKnv0sGPOk9kqyURTuEwrmBSyALgWf8kMVwn15ibPOVpkGWWj73eUJcBqa0BdjuUmXSvYX8vFSl
xLEGVq4T7RmxTGrF4il5IYPZ/5IDOnZJ6BCeZ7x+ZCpzXa40GPNGJdniEnd0Paz4FNhxVbzJVWLE
0nXO+u7Rg2M6tCVBhuufMAv4jpknB0HDa2EH3GVsWC2jkbatyqI8sdaypKUf4p/qPlTLtI16hYpm
QO+MX4FMwwi0FOGpBb44JP5mK4H0Y/S80uW+IpYRFMAMW3cWQ5m9nq6dUrQfV7BeDoPdKC8F29dp
PPnnUT74kiOcjKgsCYzLt19wN7OHnAKgSJQzPOvTiXNHFBkVzWUyk6M8mwLfor5H9hRZnnLXe44r
hMinCvzqmVlRn5N7zP87NofvOXvRqr85Q9swX5QPo+g9w1ZoaqYO39XAAEfIcdK7xUnarTekcTCJ
Io9KG01JwmH98LG/RgDQbk5l/JBapEDdLxDVxn/S2o2BcQ1babrASA/m5cNlHKV0ru7yHbsq4aLc
p66EoJzsGTBCMpt5JggRzHn4bfkzAsN7O19jMRMxlHYeURxGCyAT+VV12Yd9eK1Aw66BgBC4C99s
wiku3Rt64xKVsTJzvBod3gcVhwz/k+KIXjtM1P588cLVsgiNGhKkGJddfxcUSRE8fZUSL/w655cx
0Tc0zYH2Pv39ekOBA55YLRyxFVqugIt7kDGSOljn2FielXNIamsdTil8N6BRNuX1Vr5n1hKDyibd
wp3P/KDTgrh9lpxamHOOBoU0HS7wvUL2glcNhG35B0f+yG116jSpxKiQqWAWXu5JiBZJ2GbqeV8E
Dqtys4lcyUw8rZWFSAQd3oGRZlRWQ4isYwuqEFp09QZQTEp6gDyGaE9Ajqlbo8nCrk275KAPYDSi
Q+FrM+zWp63jLP+FYXhpbvCMdEJaqgapeeTAm0g3wChjVnFOxbqXPUMZWlQmHXMDNfVcgPY+Rzen
WuJ/QHuTnmrZzbBP2qCp4BIGl41TsMeM0tWov7NsfJm8XEl7F6ouwK4ga363UoJK1ABwd86tmi45
0P01ZodI1V7ZJDc6A8N0v4n5khwFeq2rkJsknOU9Dhy63KYf7N5icAS8kk+2afnKVue0PKvTw1sZ
3xvnP9ycMvztftImQ59Sb/lcBBMs3VwoeoXZZbQNgx/FN8OgtKSOQqSJUl2e5WchCSnfQZjwZnLc
RpcMmF5g8jtvRgKjU0omnHxD6V0O3rKGGWVHK2XZ/CZOqaky2/tzs6tUiz+5gnN9LxPF4bKDniQ5
cLvZ74ijfqLvadMeKRldH47KTrEBasNrFZONstr07sDSxX8R3c8ZOPPkr37QjZKNmxkY83eAFkA0
9vOU5QpB9kw2ET6vhsofAcRGVp5PKIrex/XL0DnEnvgtcPIHHY481Xm5VdL7hhEZhOEh38pTxJcf
EeI56mHZ0MorauYaBMDh2C/m6a0nF8WYfR/qtjs2+n6mn4yH3TZasmOyzNQmU+S79iPaAEACokzx
OvcKQGLfcgKLUDP5fbWKa1A6vgfJr5eOm6b11XxDOeW70grJMFoGAILQOoW6BdvO9+Cs9gWZIElg
RMLOzt5/WiwWe7JzvYwavdhtssxjJRVEJaSnaP4fA+zNHNe9Y31VwKK62goXL6TbFhk1h6FuIzEz
8+2DfDu2fz1YJS0YDW+RUPJlGZ+v4vLiNBfcUMV5CaQ6UpZLsBeFgEJzE6DCEtdryXFvWxkLySYk
T6sclClzoFC+0O2nkPrV8tML/gZt5C5GZmHPFkuYnWStRqfy6181j0+v72D/4o+0ihMXGkRkFvUG
jB57YTaVpmsYgc39bxRKg5jWxXrRvgKjCXQAkW7c4KOWvmZNAwRVekfRRTZT8bek0j4HP/1Z3Pod
gj19lcB5GErpzFZ7+Z8Imzb0wb4JbfFpPIZ6g/YqTqK8ceonlVhxgc1dVGkzrmpLOPfKMVHt7w4h
3A188AH+yIhfi3j6F0mxpKA5qYGAMc7Z38HFWyCVm15S4qt5c+J3ErwbZioPHdoBCkVDpZ7yD0PU
+Jd8qtXQSLzF8cMxwHeAX7P/4mLSO9pm12wGHkbW3aTFn7oYMEb2SjGdm+qcBVR0Hl0Q4k2SYGgA
Dc+ydBoaI8Urf4+AW9qxXkdsiK3Kry8qyWon93Ld3UXsRmRNTLO2ve6W0hyPZZ9FTh3ppl7r6yRQ
qE6wgucFQt2URoHmYPnFsnyEGn/DBBttIz7Ua1NxVKbs2nwP2NXBCtbqF3peqt812gqyMl+cX+NR
qsoZRmfW2lgUjSrfplAAMVxXej5GOSJsD53HzQRvqpksnQAzybY6+8Tr7S1bormIpyzHtWumyefF
0KrFCsJpi+RQL2DXGreDXVRThpgElBoaJlRnfSTmbL3QWPDMZYD4sf3TkLTbE3PXTDS1AKNBmzoP
aqbtOkaouVyN0aYGV3f0urUWqDcADr4F0Lo7E8jQS3nvOuP7eExFekig+1Et39wIX3buHfWGQCmj
YRv/ctNpI9JYBUrBmMI07Srtc8yVCrgSlHJtuY2h7ttMM+32PL+pykEC0MGpkfOMlmUU4tktwBkM
RbzDRz6K3w2Ovw+UsLOUMn/4k3Xfl7tkXhg0dATFgW1WYBWNAJinV4TQA0BTWSOmQ43bRxqu8pfu
l0Kr4OB0AnOjJ4aZgIAFt/InVguZzXc2ppU0X+YgC3/jy44iMfcGG3+ZTfgXJMKp9kQISR6e28OS
+r5oL0C5QXOWQvRdTg/E5nwfWKyprn1cfX1cJbkUzmFvMCFHn1JGekesEaIOcbRDa711jf2dPoi6
RduCA1DDRVsrrHPji0FCPHVaWbxIkQtX7IGpp0upicG/VG5YJO/p7snCRNwYijAiknJVmnUbvXen
ZzgvwYuv08fvUfcmNcGznx7em/EHmuL5o9gPRL8EmFjTywRGGp0TTGObBOUqMoLzgmJAPSATveMg
ZQyDV4ZbQtwJmyENevVnw+RR/nhjgBQFzQqx6iJjGMqbaMseEzUKl20pfeZfeX7N9TD9iClivV34
01ld6ZjgjhBGIkdmTyFQ7AixsMYUmFkjgsuM/8jjtmwE6lfudE36jI2KLHJvS569yv6rKmfxbYqU
5E02PuK8lI8sS8mLXFfLm9tw1unEJnQy2XgLKIVNQGwKGsHaN/ApZyee7V5s4F47mfDbsPN529aM
j1szHzplp/5Esq+g67Yt/1d1K2Aad65Mbh/JTQw9m9syWJMQhN2Z1GohtTs41mpaUCHtKUGjjihx
o+Hu5pTLzPZrD0hhZB/dBxBFITMZBS57vsEAxjCuk+Mo1G69d5Rw6A8YE7yw45DKR6zFcdMCjKBg
g9tmk2zV1qbzWLqkGHQQBpb2IAqqUAl+zNe7BSjiSm1ZPyFVfAYEbCQ6ncB3Z304TT9uhrQECYDX
dnLdKRoQX/3MZ9abVoxXr9UPnTG218bHCB3I/deOzAoURjPc/MEOTfH+PCeHqjTdAOznk+sZhl4Q
Xc6ay5Xwj9txOrnxUjMF8PYdf8I1JIrOAvOIRZjS2fbAux32XGlOKS+J9dNhPcdCuTFyvFuh0dt4
g4BFpOoURJJIQ5nnpybl1lJQdrVL0iNEQgGWC1vAE6g0uNTz9DABK1/FOwVoeh5jghdXIKbvRdiJ
a2rTn9GkCF0CCLBfVCCULJD6mlx8y0OuIHBvBfvtA5Eb155Qw9fCybi+VWff2omkSv0DFvL4Nwb+
XmtwyteZGweKtKI9kO2LecMhTZRq7aHYSBOc8XnS+eXP+h/TrFma8kDH/mMG1Qr3zc8EwzcTi4rb
MpdoblTwiyQ96dw7olIee8ri0/e562n4qoNvLRRzcfqiGfxxuI7eIkUvpxU5dHT//lYmi/wpa/oi
8UnRrcXryoRE0uzr8pSQEXo4LdE1jI9Ta0eC3d8osCB90nyHWvQgGDpHRSyzLUnTj1jMDW493/U9
SQu9tv+Z12ffSSKu9K/AA8VAE1H28cBKLlm3zH4il5Teu61JZzKkBtxGrzuxlE7y8LkrdPPOkYu5
aRQ8QyLcxd4yptRQ1cYwMo3T29k68RewNxQMqAcXoIvXPxo9gInafgmSWbBd1Tcvs5x3hf7s5C2Y
wkikU4FkHThX/cKGnctwATbtIUTbYUv3FjCUXzQB3grqlnkV8es7Uz3KBf6BtAjMsATUJwaWDKBh
I1pvctKCZ4OHzjGtGqhacyHqHMBrANU4y6RVo8fauWyXgakqx3xpWD0CQ5Aui7KhQjD1Y7kExNAk
hpXDUrAnXjnzA13vW3NZMvIauWDu+nEw752XkJ6nRT6fxlkEX2kNXGp572RfpBCimZv2KqCj8eU4
thAQC0D2gPce0g3sV27Bk52CKAkXGstskDgn6N2sLNXdpmxuiWOo+4beKSmteSPMkXnm8UKVIcOE
pF/j4VjPMjDJ9bMqGzYkN3PylBqKTSmdyPo9/4tuDgZTAfBnbr/lS5VcCTpEGMNb6G/gabLxd4bZ
Sx74C7ZHxG3Ta0gh3e39Wj0p5ld//RhwI6CfeLG+TRK516n5GXi7LdphN6FmiMdrJDfhuVqLYz3u
aH8DXj6u8kvPMeKa20XBGQYINbLplkoivzBiPNrPhE/sth+iwE/e36WgxPvB4Id6RbPcXxgnoblz
aMEUwNTzLIDb8aiNxsjahpzVQbCYixKBBxZkq/axOypmUmzh261AXuWFthz2ChD16pCsBqViyV46
TDLuARlEDNsv8m/ZvAn2uyaEMHQOlaZDzsagfUhN5/EAtBjrgLWIug/h1TicEonYryS71V47DNnk
YkEGqqh/LFetrAo/YLwiVpwx4lq3MzxoHscIyzOk9vn2tcBi5HzeSay5wDX9YtxuB+z/KtCiQxy5
Q7PMWYLbqxhaiLk33PZ/C1hG91KDR52w6kFitS/bGgJ7EeMV63m3uybUhNOBXo45DUDBt2MQusn4
2T8HPYPCJLW1riFs8xqhjTarmR5gJ6rwVm6qRn4xhibdHVULrFs63T8E3QfO3QPn5I67GDkY9MzP
IDyOvg2nV4lUUt1cGOPQZ+ZnZapZIIzhZtGc//6O+GwkJmmlGZVZBlSxjDyEZjSBZxHRC6JJKH/S
wVfyZntcHlglT56I3qbhK0hqdzHraMRF2gGkD3CG+WGobzdAO0jh7XUvR0XUBKxCfzyXcUjebUeL
5T4xp4i7FrZRuTceQCKU+hNw7ovFu5cV00MSA4aU9rA5dyN8Ca0cMDz3hR4x1lcKj8BLcccX8Kj7
SNgdM1XcHqaFunkIZGd8+372yVqIfUDbSonJrdoHu5rYQrxWYedhYzsq93j9X9K4ox2DFVp2wsCF
WLesnON5e1m2zAZcGrjSlpyPZk1lB0tve5PaLoUqvlBO2lpexfO+fzJQsLoJPf6/TiDLMMqjETUR
Yzbym2UkkagWU11JkquWe98vdZzUEUe9TRMdxajix91cd7w5iCbfNhCatEaIe/5MuoPI0jn2XnZn
xHhI0T++bp401oDdl1S5U6legVRm1yffOAyjGUuVakmHV8wHblo4oRxSNTmvNJJwrUWw65fFz3bv
+zFOpryc0ZSgd1UjKfgCPaAl9afFkS3b/1PLmE/UF8gDbVj5gM3kafwa4B8CV/u2u3YlkeXVJa0Y
M4hLszYOOoSOuzfYZhRa5KOtFvW67MtQInJUhx4eAO+K1QfTx0EtwGQZPh6qpwpKkmk2DiAMLDaX
hjs/4H7itpGekUhqHzeHaLt6m8dGircqsaeoLiNIU3QGzh7RNBWJfUzGaChHywl8DJ0OfaDx/XXV
hejJYma0PujMdt33gvCZ1v7xHrHTTzP6Lwj+012i2ZJY/dHrB+4K6PVXtuDfuB55q9dcIOWOvcKs
gzdbhWM7Ny42jxO60xCj4ln1GmzYyR2dYTDgfcIgR6VvZP0NdSrGBa7XiKPFs1BB3/R7xduKL/LP
+kSU2syACArKDqbMEmbVfeJuN+lI5ClCZL3P6YCNlzBeqXoh2x++NGaWgwMGF4AXZ4HDTkn93qkJ
1V/zDJPEb6Uc6mn+EFCbGPuQQjqpTwgd3mB5ZanIM8vbU4A2SwrtRDuJYbc+iMFlO4msoXSDgpy8
jSa1Nr0n3p7YF8+f25bAwVMfxnN4Is+KH6XaMqq1YIwok9MtH+/wFEU4yquEgzFLIpvtGt/C7OSs
iPCxtBaK5wMOZo0ATjNeDaCz9wU1LK1Iwfaq5nPRITLHI9ZtYSLN+Wq3nGBIgUOV7rbOu2WTGNjH
KtIq1SZ+ZbgKMVLOAAQ+2O+UpqddkG7mnFo5+s/2JU+jibV0fcBXhr+SdwexYMehbnqA6j47Oj8F
WlTt9Ovz5bNnoQ/ftuWPlUoeKZRoD48186tM0mCNVYr7qWq/c68vnPbuFB76Er+NRaRhu3CYu3wu
FN9uYbk6SUpAW+0IN6HKbnAyShwnDwPyBWZ1qPipoePUao35hOgfd+99tQHWZ0zaTKVQr/NckmvQ
WMIpYlM+LyAIxSGkaMlWh6zNYFN7QV3dy6CklgVbCmEAaxsB06Z2hOTl+CAvy3PH4SFKk0x8lm58
91SwZBy7fdMhQ6u+wfYujGcaGQB/OSH/bUVxHtMxtAa3Bd80Otl8ZvZeTl4T+J8YLQs0fVZ0q08j
3ZlPGF7+WfXtQka0K7/XSpSMsC1Z3w70qe54C7Wc6j7JoYrj8Pz5Il/F2lRn7WCOLXCxc3KX54zm
IAexAegvSYS0Dj2FZxNZbLXuQMKtxoHksT2XufifgoFE6CgLqnZWtBHJslzrtoUE7eyyjSIgpWY0
WtlC5a0PvMtQdb5cCs9cJyxPTYAB78fpNgJoYCP0J6P5QXQGg0Gms4UFqF7iSg8AIu8n8e0Lwc2G
5bzcrmhG/0PYd9/fMDpqVSIdJBHdKsMkiDk9ntooJ34vNVORl6Rx5EGwhVNqe0MO1s7arr3dj5oD
BqGWtWjkzJZ8ZjqfFjvhCvf+Fc1PzfbngM75MobiUWeC2WJudBC7y/oj/2qx2bf5IiF83krbL9jc
aWFxwM2U07JKyCL+wzSyGWxHGIwT7rhunX0ECVxB5iSuTEfSgWUqI1W5p3CAXU8s6mIZdB6xmL8N
sxhxp4OlI7SmOKbxtbEufpfGb+gPI0DwQDXfoSy6MRnKEkCpEbNvK7s0BKbDKHtkhX38wl7OqYiU
tSk+XCVNz+n8yvxYyLyzdSwvaaT3VfPb3ItuUvIYDXd6C8aZRF4207EOVKjEQoI8nFGIVGtxWXOk
wkgyyRs9ZRfEQW6EcZOZPm4++VVGZBMyTmzMJUKYbhdC6H6roKZD9rwaF+uxpulGpXhstPlGQlf1
03LWl2GSpORrJfDcHr5Y4y/tPMzzesi9Md9n5nXHqHCvLcD+48EQ9iqB3uqrZEEmJSBMP3k0h3lq
2bkzE3At1HWFbA7TRJSzbKWSJyGxlSZUnnGOuXtWtperzDwbHjrXxlOMlXZ0DRainInsKVkuu+Sb
EC8dvcbGni6arq+7ofJnoTwwklIGP5oBu6C0uhs0VxduMqWVkV4Wogo+3CCD6mCHczd/vmoy+0wF
1xjUTBdz5rvlmhKTuPnDQhjkzrBKGpLe/9WR05wNerPMKB0J5IsB28+mbCgYqRlXQD52SdnFvV+U
AN1UMnWCHmhTh2nDs0Uk85cnEns4VjsTL0gJ8/IdPlB3z4SLq4s8DyUHDXFiMsdlUDiECib8RxFn
Si9dtDTRPKSRhJ5lvTeKA+U+QNDhabmVyOGtINj5zilN7nkamHPZQX8Q59CxCX1f7a/3IuUCHzos
Zn0ukKHAhbpc2JFV/rCAI/mf2rlcUU7fJIgQCFTT5nBmUh6Rww9rEba2bwIyp5rKFF1s87nb7ixq
6vftBeQLHvLnx40aotw3Vv/zQSTx27rLEUwfxEXibxJVU/KVjkABy95wCm3jHJvixvoOuM3EP9ss
0+UwPWQPjuN0gaYR04ejqPVMYB1Lp6qJeG41rpe6JhQGkhrNS0t0F0A6ys3NDHcjvD/G1zUqK0j6
qEHpooJIs/1Uz/a5p3reKF5uXee+ZlR+EQcckDP0tLrdnF8NSc/62iwTT12EfhSrT8UIAzHSJTI3
Pq56wtJLILUas4cj8PrJtw9GV6toBvnZ9I6k9HKWStn+BaIINwa0Dx/k4ivpVFZekNeR/eDaarVd
0Emq9ecG5vxQp/oAd0VceckXgQKme8e6WUpVd/gJZDrbP8s871w9Ptj+zqzmGYdiCP0UeIqu6AYr
FSXT7Rebg16UQUkvsI6pMsZ3izactrGGSK86a/fyl0CvhuqDkPt8ywOSgT0KbrhLb6XicITyPpFo
PhBtPp4/LjeieBxBEUt8ZW3JS0TauLD/R9Mg6Epv1eSpLx1SkalyeC3XgH78E+f2RmeH/EknSI2E
jJ4YEJZVrKIY6c12rtEDt+82oWKkWAccDshEQDI0BtxSMsPtaP9JxNxyFVA53kHld2Cf6WGNk+Sr
DPUEsexLTclmX73ZCiI5S/ulbSwXb+ETH7g2dl7kYA/mB9Q3tsLjfmbmnV+rjghZL3vL7BTeZvLd
ij0pinWimQcnyKXFJf1aekWXlyotNOlBtg3nuQfpErcja0kntQXQGKzx5ywH9Q+6QS8ugxIZVJ9q
GzXcsS9Ye1DXBduNkBtl07ak78CYRabsUyQaJlbRt+V+HsjtATUn/3UWQYiNId7dF+9aSzokT1Q4
sSEESBoZjYWYcEGir8682oBrWH2VuF2E72Pn2oTNcp8a/clw2xYkFFB80YAGeAXuCxnhKBcrmwLj
OEC0ZeRkLJTEYQKZy/xsYWgFq/kXn0yW29/8nU5gfPzyWviLfbwGCWB2zri8XMDn6B+vE7ieTSYe
efEQkS7OP/5IO7911dfHw7uwCYxLkE6x/ZKfO/IJTy5PdpUkv52CukQr9EYRvmuM3SG99EoAknGM
6dPf1ayrqORDcrFIY/X+POdIzuMdvrTCo5ABYPgWbTx8lMTb+xgfaNgO9495dEv9AKBnuQZJ3328
vBnl7CxM4k0nwRZsHvCpqySd/Q30iNuYjqmClI7MSv6ocbKICroyNetTlGLv0tmbQNctXbwUqOZg
Chw6sLCpbacpTfEedRovWr66pUupXN7bualn/SotyqlVb3m9sHuJF9cG6Uk77OyoAdPk4OooUjnZ
KDEh3DJ294VR7y3uElGfrUjogC9QWdEdZBb23T7AXnYTTeWxUw9dXIp6SGnXuKQsIJnMz9QZ9HIf
AxV9oIeRaleyeMqVBHaa5Ya3yyf1yOe1dnH45xPJszGqGT0t9RBr7K3e7LQMYzV194hvVRgg+IJY
dTnKRRrMMd+oXIgavUygoGP2Vp2w3s0p4VKhE8pbjaQjEoC7XhzYbxeU66QzLX/hZNuahAy5mwVD
tazYOnRiYe8yHU+VZGYgL+QdCR6zpupbOEoETAvnSU07JCPvrzvsgheZoXQwdfsIa1qtCME3e6wM
FTqyJgPdKP1v9DCU8dFjcofMDQGNgvNqpRkESFj5CLyp6wU+R3AOMujy1qFMpONBpleGnwL6Wtep
z4+hmQpZKBUs5djEohrtw5pelKS3yVqrCjG0+7dOLiQLuerOx6drLVDtWFlfPIPUMoBLz4cFHzqh
qeQsaUN+kxdR5zWkSqxtLsvSSsbdvDUCPzm4gUjsCYJrTuvjWrGlNcPyR5HKOJM31fqnik9q92wO
nsGV89IunZLYNiwpFZlkB/+uCwRgDM7beYL2YlAYcg0+6lj7+69Rr02MFTNrkKdhk6F/D9FR5+pX
m0p9gFgX0yKxEWjHVijOxkADX6TyLtR+A+yZAm0u1QIMKOiaAdTpXchvUH6JsYBuAmLTn3Fw9BWd
1R+eneoV2BQezcIWYzUVyvUIxWpsJbx6c82ZwGfFcqG2rcgpLoVJjQdobtukQMxmQTP44F9nZvlJ
z4ApBOHlbhtl0MnmWUNsoPLMKjW7rV3xAWnjoyG6y96a+KJdmLs0pURblEUPzJr9sjOSj9EQjGHV
VeZAx7oRFOu6AT8+kQHmRaXbj/S2FiTDm+SSCdwJSNZS4PxKAaF5D9ZXbUHsseGI+uEhcKFz37vZ
cvdLYjX+yvhT2ZcrCBDQosnQZ8e/csyqsnkM5YNxyYmhWV4qJqicygyfKECdxILVf5SELDwS8SbI
UXIqQcO2jqKRQT0Ich7GhDAM1qnwCYr+9Fn2bnj8jp8FTnzi2LPXJkEr8e39hXzapWWHFq9OUQPE
mDGvnp5jeIusTlRsUF2yZCQ3YaEfX7k266glff8qfSofNiRUm2AjLkWk7pa3Y9zzvtlH9uVwq1hC
nkXFWKFOLXPUtypW07XdWgXATQtRnUunG86RIDLmuW0YKDqZkg9diImDeGP5ru6St8hKSQy8g2sj
LIL7e1WEPSb/PS+WszLFvkmhwr/X/zMITD0vaMzeSykslf7KQtc+e/zw08+7s+26kNohzlK7FoRE
MtOBANhMsU/QeqB8Dw43lNTFfYyV9H0pnqb2t7/lehYnXCIHwqx+Y+pXs7u19uUm45fk2oat4dnF
U8vCe/q5oOOuttuWY5Ge3ACILxSa+2IfW5CJcXJaK/8oqoGwwAIbSQOA+LvaO/jm+hira803/IVO
BNop5ug9x3sFCIvc+jBP+3b51F8f4RfhDIVB46O8J+LpEjAwTh3lF7ddOxBuPjRk9nf7Vbpqx4HZ
+YV1utudDhBOmogdwsDbs9CLl5kUUQMBaIgWy33Vx/lN3estq9gl00FWaKZrSxwQcCNdRKJsd014
0T9UvLIPdsJzo/vXhsR7cRsldS6iNJ4kh5wtj6Rie3s9XuDS9tIYD/bI4dnkeu8mGMY5VKE49nKw
jbwuAOx6vgDw5V8aLO/5ovFwfSkE0fF189RQ+LV3tYa38pUzJrzePRk0WzZ/G/UolGwtKZ/25rmX
4ZcQKdUSgv0MlkrzW5HdxSnh47+p3AN1p4w5QrrzGRmPrGCm9gJpnMAqJfCp//f+kY80MoIxaBlM
GwTKEp9GCf1EOKWJyCAzHA7UzaPrRxyM54/GScExI86G82a+mnKwiewZZPo1GxPDSOyzjkpK2sah
qycKsfH9LbaaRuyaRFHgC+M0vlgbekui2dS5OUXrqq0dp2RNbPHV0/rXqJHt9TtB/gPkpNhBViP7
Pj4/ClKc4ESlVDqDSocnzvsWy2GF1NRz/aHsukPHhZ+s8R3cVRLbU7mk31N/tSeeUXEBgEObh9ng
/kAFNZoqJlqpAnDioYNFgwkKGjdMZr03HJ29fyWBK0E8dQR25vV3gEFsmPEfOQ+jxW1PJYaqPMe/
KAUhhnS+Qr6qlh8cuG7VGBBVeI7MM9i1dCeA07LVf877ErtKJ817GU2SyodFpfDiwLA0FMoQcijT
Y1e+NkA+B54I8NA6SmlA13JgmhkdAD18NeoSj679Qk/EZugAM/qNnRFkd+ZHeFomtIogM6esEuFT
gXXOpWjkL82u8txy7F3o4Fn1i9pjqQcFpb+VFJ/49OfLl/YmccXlRuES5xNi0mnrGuXtb93dGHMf
yLoU0UlZtwJY0CIZURWSvS1liXB+62O2jjXOMf+j/s6uHsjjzQKeRKHsxhCSuhKE69Xa1utcV3CP
E/9hKb/9dVXBNtiC5zlWHJno+0QC5AEmNzYNT0l4VCS3Nycqd+EprsfmEZq6epaxdctOQPzE+O+N
Qi1BTW5tKLl6sfCt2dm7chh/qObq53ANHH3utM40k8DshHTTDQvTZD2ZDnxCLZUjJEzKADyRymNJ
2zubT78ME5rwu+f0wK+EHTRv/i6RTMgq6hVEYOB5srk/2ZHPOY2LwPD7VQUHZ7k/J5j1umB+VLjI
QuNyIYyQjg4Bb1nBRPxiip9P/YUJNmSGpmYUJKzcPrdQ0vR8clLfNh9m79+K8rUeeo6xrU3WBKiG
NQlbfWCzzVqoiIEQDy3UwLUMVA3dT97o/q8PhGDI+uv0/aC8/Zvp2RL3jukirZUieFrjkARLNHn8
+DcGXlf/BHC5epgOQa5+baPJfm7N2yscg5zsaX64UiOpPReA3DIl745Sp1jto+7NbrTIDCTtBBBZ
k9KWsi9fkTk7qUdDqn/tp0R7Aa6COas4Im5Jvzuoc1N5Xc/7npwb68JhvkFfn/OGNh6Ps3SP7mzm
2NZ2vyv6wpdim0T92mdjB7iwBLls4LIOBs3PFJNn0kYld8bhVDlOn6xeImA94v63dLGWqO4fQXJ4
l2ORw3z1W8/HscRwM64nhrqyj1PmrNsn7QUl4K5I6PyC3rTm8Zj1w9RlEpMPe85hU2OtRQOS39Uc
as5FMsjVa8Ug8k1NLxOXEPB2Gg+sT1DZoxiT2aTJjIUpuU6VeGfxRzvpMy5Fb7l6nXfHlXEHsGmy
g2ssxERVrfDR0dj962QfDk1g5ldsGjhv00kKjbKtsAV50+PT2h4GChWrTXEkgCbvDVhcqJfWk6wC
SK72gT1T61a4kYUz7ZUVgJW9C2mJ9z6p/B3WdElGGAyCFDGVtPCt8ZanEFUUwMc4iGoeLEiWwrvB
1R8fvVEr0LzD/hqOSwToyktA3S0m+X9koxlsNwJ8MLE5v76TxqxRDoEAir5zx3DXoTdFsny3QvPK
hDaMqbtkK0LwmWUqvkntebRl0RM9KrBtQeQi/DRoZC1HDx9DDyTO8PcwY+LbMZf1Q+4OGJErGxVZ
XFl6sZVRkmilFXfsl1XVyAC4X9OdMF9Wd3+aCeWS/d+XkNfH9Vxcns/+RouSfugQuj93zN+rzPeI
4UD8otWHfJa5VrhKYyX0OnX/9NvesZQvQPAbYcj+RTrRCu17Afa6/awH/E2z7qdU3rc9GfMnNFEI
xRID/rRGPsi/QzIJ/a/dJCi7niP5UkDEekHDxrfIskx8qvXn3o8cal+wfkh3AQg3iuMFYtsFrk0V
ATfgErMKKY1Hombf+IMLWXderFQtDoTy4O9hMp+I/hB9yDV9JoUHszf2OhMID6lmFcqYiJD9sBn2
rmYyFTtnl0RsXZpCRWXq0Fr3K/W6yTOXYhshe2WWGWcvFA7HXbAI+stCas24xcYX6ouita4LIXnC
xzLYOllYZerwHLSSCGuDzh3XhEPKsYywktrobmugPgdUbuPTT2s9Pc2dw9t6wipO8MIXLSVdDh+b
GwKSTFYaSLkBpw2CuHd8Kz8QUGU1g8jz9n2H5QQUm3tBO9CXn2DNV3tvpmldE2XTxMTSTVOw6Ae0
3ciwBtMw90dYOduC9Pji2MBgWTp2j/lSZj3Eif1we/jvfD5Z2Z3NbcXiJY3EBtkYo15v2ZEc5LWp
AMGNzg9HmRrXj86GvH7NiUvkP2uvxh+TGoE+sPpbtHCCfb4dJ1VdOzcnwz9NWDNeJ6XntVVUuD/M
J4S28dXzv4YtZB2Ms+PM6HGm3sSRgQAJWEGfr4Wgl1/q73aAfsL42OCN6itMOVhOyeRdeMVmAnFw
GwwClOlHgZR2vW+Z3uCU/wwZ2BWrDdKDwrn5REqND5GkOXAztwgLbmZCyAKq3JK+rQQuQAh8XAvO
yNvRagCliUMeHzT6bLLKTds9pDHlIGLE+pssGbnNPrLil+qMWrmXuZ8ZbiegKCkwBylQUZ9E6FV1
nym12AGAnTggfB4ejUZumvZ8zAvdZYgjIr3d9/jS02faLgE3UMDkEUfuD2O/ZC+4ofJuVf1qzORY
AVt1dszZ9C6ATQvPRixllOcGbSblLEhJPHRrcx0VE0Hx/PLHop7ApnCC/Io6X2g/myMNRy9KFuGp
FGh2Vv7ZL8PQl0hjvjq1gIrVmj5ig21Hz1J0FCi7LLPIGzdKVpLDafRKbfpVzmEkHL+VtJEWe7Um
xEArBMI2RIkOWIAiM1kqdjpeoggvuuTLGlz/fUtiy41sfjeTTYh+kei+EU598gGLzZnqXvrK15SS
RQhIIzLTE2/ACb6b7d0n3h49X7fwUFT3prS5Tt/wvjKZ8MIRjU3/7c999f1V18aTze/nRe/sQoEa
0XkbK8LtzWUVS+jpBg0Xp5Mjk3VDQlO7grV6G5eRf2L6CoEEM5pS2OLq1q4LFk1zHQni7dPmV+HZ
myuFAQFNFgcZwz3tfAYlidyvsFLKhKkNawi8cLUtAlusVBsB6DQVPHVYyITxp/fkNMgYmNKjRUTL
RvFI4GNb/VeGPwm8ffb9s2aBRhom2Ym28PjtAbK4nExoJWC3K6j9HLAu1+x1DcbNWSJY02T7vHP3
Xbp6VvpRbJVmcdV9GbwuXqFnWNIUl6NeX7wuMGxBLUTjthN7fChcQpNeMTcnXVAScIReK/hl0VrX
xFs7L//rH387pM0Fa0aEdCMpzg+jx+PXqYh7/fVJxC08ftF6kHF1ZbWrTg89k3Vo+QCRfqFgElmk
L2/uDdtD57c0SlX1wF5TXjggumI+3Ceb5uSkcX5hVQWqrMof+iQH3/R6WAzjZ4TMGTSVYlOIuYWG
zFjcaUS99ZQRqA8rf6cksAvKQ5fvouLPfsHxvnskhbzc2qyrHF8YGTNyjMk1cQZUm6ClotaGzWPY
Qq73xf5Ps3bhTduMMWJulGYrx0e+zp06mxTE41kCdVsycpcwXrDoCIvhg7vyPs5gAMJsO6SwCYe7
voDaGGtmzI1btZXhEjbSRa4molJ37SYM1iaT6KRhSFrydj4sRWlTF5ZTZEYJEW4MTLpF6lJc1Bee
eoJG0fRM6Q0EUf0YZ6WrhdKvlbn3lt9Y4OfVLx6WoPwy57zP4cUi4ncEsxM9zPy62ZwLOkKIwaZn
mLFsTj+nrfcDlHbEyUikg96Vp4p+xHjvKrkd452Wd2Rso5cdVWyukyOQ3kaFmHZYUSxK2uRc1jRA
XCbK/G/F/HE5PHDLOvb7QNngrRSK7iJgR4wdGdhSt9A8RFMa7cFxk8r4v1Fg+/IxTXAb1nHKttMw
P+g1cmoE6CKqWCOMwEN7ecNtbFnpqYR5n1Q9DaPQ1YIpHldYU62yQhE94uRVz9hQOL1BjzwA6IU6
PAXdhTu9ut0IqGi/Sex1Yc1FwxUy0AfREMh9s5QbbaYnsd0etTQdXhXu6LUKrc0Csh7hg8u8ubSW
DWQVpPf5r1r1KOD+EvU9EmGDU83dCLIf7wEcS/kp3gyIjZu6e3cN57PcpOry1iyyulHH82ehspxw
Hr8Oo9xGczHa/tF5F28496PpwCEmNcdwFzCCX2fmlBoAT4buaxP+U+ysvhngevwHdpNXTcP4Y7Tv
l6mqtgALh0UsVS/i9s4cftZk2zMGxLlpIf2nBAEIjGkcAwc7mFJM307JL1A0T11kjbWQDKVjwGfr
8mGwqPPjgclKefa81WIbW0GXW65rg+Sz93vJyib5EyPqMx2cZH1Qe5fLsh/ldxrowQUdFIGPqpbV
2NYo+dqEaDh0c6voeXum2NrZaEOAspzPFn7vHe8n1G1QHKYaspYbDQPMjFamUE3t9cHb1HttjKCc
HG7/hSIUymYQnAxXEaNeTR5BtAWMYQZg0Di1vFmPQ3WqV3lmg+ejWVgNipfnHC6w8/Bef27rB6Rp
JRuiWhqQOGZXYr1jlMeXqSRm3ZF7nOWfc1dUSqR+IJXhkQsn3oYlcWTk70qmCoT+EG264yzuiXUb
eXz3mEYN0bMpmDc/TQNOYh0bN8FYvMZf/FbEnkUFee8fG9yeDQfnow+DifltCMBO9PwIFttLgDgZ
ZHMqNbcqMzcnpKHvNrB+PZZhD5XIA3k36PKa1+E25UsvOLHNtE3hSG3h7bcE3gfLCaGltkYe66g8
yBbD0qHhEvZrx7j38qwWp5UEwfxdHEtD4ExI3enpT1V7npsgTkmOMAD0+1fOQqGImFLCP+wB0Uy/
NGisUyJ4qX8vjQoI+w5tkw+LUEdh6GXqAbsgnwoQ+GhTW5m3GESZcktP6yuefLG4fo97nnLrIhCP
lmUDWaOCdpRvHoD6FEoO2jcD+Wz017gplGk+ouLZhvpy5ZvyBsIICTvlBcsK6F0M9oK9wfys4b26
jmsk+6n1ER2bS00mkFO0GxfIy3YieKc7a0dMR0EPIdOs0AjGAzipXA70CISKHBBF7ymebPX8E8y8
/2XV3U/RqT8ZGILXdAlvXfLjAxgHjyYfipnISmpdtVEC+Mt0I+pkX26cnHXPvo5p6N1xmzh40POX
iyYv27veivgudhAbhBNhEA2d0b54PQb3fgywNBxGl4zsDPeCan74055WV8o/rc/dc+dGQ2vZpvvN
CLpr6Mgf6bUSUD8ar/SmGQaTuTcFVor3SPAUHzgGN6gtMU4rRh+XuiAXxH+ykIXBybvj2yzHDfNM
9r58AWBtuESIW1A+43e6FYRjFN67Jijb1N4Q0CZUoMx7zTbJKyerfnTn0jCb+N7wbTNUVKoSNjn4
iEj7jcUNW0GOGOAPMNTPiZ21MVZcOVMl9uWP4zvV534h4A7Qf/ey+p33pFSpAsIFbLKiNxYsNh3w
Tq9P3NJ2eBHDEokWLqGHDU1owse61yQhLV2rnd4QweMpB3e0oTC2p2T1SI9bC/CnAgqF1uR8x/Li
qcYsRweu2XOkt1XwEtyd4UjH0hAoCMfbM6eGPJJnSJdCD/ctcYfUrZGhKuXEP4y/xxsxA7fonuCN
uYiMCd4tpcp7WK3beOTVjxXpiqHRPBS/vqbehOc+AX9qT3PdY0O92+F9b5QNbEe0CPbsa6NjYNT4
w48PGscUcAML0l2HTALGNFVfEMOO9ENnj8xkuD7iDlmPrYRbNlb/izlx7KA5mJsY66Uy9VUAY4EW
9MGIEFcxS0mqk8k4ixgiXhepgjiScNdr+VAySLkSZwiCD7l+CkL8WWykvv6uxv9tfvPyIiQrqlre
YiTjXEWDMaFQmLgKwG2z91/cWHWFrFiDgHDxspqZSnsHOwwitQ82BTROlzFYqQqN41Rk1/NtwipU
yNG1qlDloVz2pOGX8zNGXYedNlenjd2wlSLTVdY8nZ2TKBvsyiGd/CQY/U/3gtJhZbPnZriEMN3Y
T99nsg4dmqQqS0+HoVC3asyUht/hyfkLhdqxH3ACnUVexgr0TpwMtNiudyfKLTOIK5g7RJ/I7c0z
pnDVrqxqsNOGpJ4EZuCacqS9XVVEF6ojsFmwin6zYryIYYZAKRvei2TAL2LVGBGWDVQo9O3IkF1R
3T0FxSm/ZLvgRj3HqNqQgybukM9D5bumho24hekbVbbGqbM4hs/rYlLqZkBkTyVKzAYMw72C7A0i
c/cqh6uYn7GVAw8tOA9TAG5UPfU4z8e1or6bE6BiHrNxNC2Of2rtn9E/zKoqlbiFuIXnhy5TYzj8
5O+NG5y5IeklZfBAiiLgTTq7qWoaLvN0+OKOMNir3cXR1L/XOK74BmmGnW3fv1DCNBM5Xtlbr636
oyJ1wkXabCF7S0TtgWqSOxaL+VBZlwtOhFhzQrCOqdU4U984BwDXs4e+zHLmszYbes9ifW1S7BT+
ya2m3XImMw+OdDTwNLe6FGfLkOn3MdMHGzH9V2dIYKC+TsiV3x3T7DzFP5IZ4eiuOWqNBQg2ibrH
HfXirZlo0HcVyQ/cDIGsHKdUGeD+O/9bx+7x6Eh2y1hIb88/9oKlkf+SyTAhR/URYwzEsDsvDleJ
dp+NbzdUqNstNh+tUGcwNICy34Kf+8ZChg6gl0jNdHADFAM8cH9i/d5jzv75jfSa8D9PigCfmVr+
QRIOvd5fl+4Wdcl/zwNmktHoRe2xs2dPFdiVXNvvB9ViGqUm+nSvZeCo5iA2RSUTk5yDFzSHpAex
0cWBfG3/9+NTAM+ylmmakQ2n+jSz6Hfox1SOiPHHhQ4mgh793KNnRtvpBDVWgDzG9QdPBBe0/Ddx
u61ZH5bTr6YY4iONQZhYSskPla3AuQc9LNDpecMwquO/3ztqHVdeBH6HABj+tbLsoE+ZQZ6t7ELT
FPZrJdLXYnllzCfjeUVKdRPYhbY20Hadc+yqW0HMxY9dDNTAq2aeXMD0rkEslwRX4L6DxBlT9L8K
0VoM5hFmEeUs0nqZABdZ+36VtOj4s6rEx+e5g4cadxvtwVPiW/o3q4PYWThPq5i0BqJ/WoeRy637
IVykVEN1dmr3KK8zSS4Pe5hvECPhAEEA7RNoPekm3fg+6OIFnI+8A5p69IPu7QDUlAnvTlTrp+Oj
Bh/bP/knkeqk88GVuxIBA/HyD4JgJaH7J5CNAbu9zIgIIUf6qHYdHmdzDn9EcWHcPUa6Zx7B32N2
UFbkYWW3QUCpgXhZtSdwQ5MnPSQ23K4u1DBAoixUaU3r45dwZV8Ti5hwKPytIkUb/NlFv+GRSapz
8zI9IRdZsvVF8SJWRPRFvefjo5mvZkQQ+0yzvmgnQkqzouFdKIh3DCI5z1wdym9U8eZNPd4YUx33
uB5imSCl2TVVlvz3yc4Xj3ujtZwSY+jTCQAic9laAvejFTScapy+4NrWSArdaWVpqvtffKg7SWid
hrBKMbl0911FgV2sJXWpVxBQxAi/+KTywfp9uIkMpzlxDjNTSCH/1XMasz6ubusLBkgbYx+bkrXP
7Qlw7deEGFYg55oJQEZk13vjJ7YOyp+OcKBP0xJzxTDhfoGcIDQnSceJ9Ji7hhorxjjxMOKCUM0u
+jXr2ekRt//Tb2mzmehMrzmfX0iQcrswUz5bUZ/hveXQRxYZyvg3Q2tPpZyxv/vAQQUNROwWaDVE
B2k9nUZfMrPlcxZsxFvT/9z8aINtCVlSmXvdTaPJ2D71ajPuzu1+dKuX3pRE94RSihgexs6zheK6
9rpmbA9QpJSNq+wSJ65tFRPqCEisW1QG2olzFzkCGEryIF2um6Dlg4yBccfWYzmS6wGsKOulUdiU
sF+9flFyN4sLSNxL4TvTlxfhgNt4bOboLei2AB+/1FOWFoiVSRVSLXVYtqrKcHhptGVT1Ykz29Ir
Vli5Pcx/f+Rz4KmzjO4CC8avD16QEKWAMlX+GLPNx/bAU9SkXkNg7SZtvPXWSI1MCRh0TnydFMKw
C46kSOdPH8VKrtSdt3zh0m96g6FRaTOYAwp7dKbbyJGDnOMnmNsZGILX1KiTeb82F+GZU2idIERB
rhUueXBVmonMnI2EfxAGO8f7JZv4RuyLb88DjhrK4s2biBexnBYwcr0jrtg9yEDv0eXkw7Zh+Qot
GmfALxeOKhSPV5ga+ULna35nOup/We4mgdEq/WXeBHGgdrQ/YA5/hR3PyyQhIjtlq9sNFLKD9ZXf
YEXv/RxT4aMeSV2R+pl89tktvD0b0meqXeTn7ZJ/arTaJ0EQQAofomWapB50yR1lbrxVc50dJ+2k
m0eB4pAoeHor47j8grpavmfUgk+Trkdg+h5bINhBIAIQVtKGzRm7OQR4m32P9ehBeZDfdW3M09s/
HAdbjxnuU2ZM1pBhFK2pCIpHSoa1+JYJ+wtvA0HoAdfTiDYnkwNtmnudksmz40GYMM5bDMrW0myw
z//bvYaHWahVPELyilvbRmQ5t1PimzuGrWR6cERZCs5Up7pOlFvXrc8ONQdwOlUQ8uk1ifZCCOcG
CX/fPTCzFNlwLdfnVWM9DVXrwVU0EQRH/Kxo1/ohF6ZiTbgspgpusTmDyWW3icuoU8ZIHeDS4wga
Z3ohSgHtKA3H0Nmt7sdWKKe8K9MPN7BLei+KNkZqE4Zva3LAmCX2K8oLS0pN+K4vYJQwxYOgqbr4
Vfe0EvZzMWgmRfTdShbxe67WT5QRBMd49LDW03l5AyXjRLPvlt64Mq9orBN8+ri9QqdWODW+9+/8
rLUyV2ghkFAi0xMEANksziRN/uXt86qRHe0oeQmmDxvNKfK6oKebFB7IhHzllekYowbDyl9xoAcU
Cb3sJeP2A8BoCPDq/bM+0xTsG65+rZ7KyHQLA3HxhewexrLq4RgNn8LM3e2l/TW40c/Vnyln+7qH
FNH1DX6Px8oK2zYy+88KFuHRfdBVZmsQHiPAhvHPcofQsXTOsasffk1GRa0ach8za9zAa1wuh7rA
tBYIi8Ln6HZ3gapJ7NKJ27uGjDEf2ZNQ6ZXjPY6duJYVTfo+HDV4njh2wntVxZzp50kqt7DXZWZB
a+ZYNyHuUuSJCJAzGkxpnvU8GGPzjSkDfTpuhNMDturqrRFDiaAfyTIosMHor4v1b1xhTRbgrcuH
MMhNHR0fJx2XJumsWRqI+rVaY6uFtdd3KGyphYoBcfsiQE7GHzBmVJ8kFO45C3vVNi1WQiA0rmgZ
lNzlmdkwy2Rcp5PdvuRQWDYVUiv3KAVnY+22W7nMfl7/HNCayeKNR0FE5A/lxSPjHUGlK+VSmYxT
EvXvug7qtuXcQfvsXIy28lUzEDWP7R+WhF1o79Ud0DsrWUpWZXmnw3t0SYNov1IzX7icCU2PdTh9
2q1RzQBB4oc4AixFmFmGLlCB/P1f1wUWybPcGPg1e/LPgN2LFcw29lCq7UD9XeKPc1vLF4ME9kCW
RSvh3H7B94IYCXAKwZBtgmT4/C6FOGud5h4c9uhxuCKjxiGN+aKRAOg63Es4RhRaZj9skO5JIZmr
ZmXFciBdcPFAR+y3OSC0ReTD6iR5yCFI2SykPCa/1Zzp/gXLtuq+xI4g1bX9wtRqiHSiE4CdKsVP
+0PShA/bSahh/Sgf/CafGwgpSLb9hTVIUvAtjJCuHpCXZvxLgmReXodKx0MhvR50UD6oBP6nz3ak
CBHv2pRon5b3AueYGy/faDc2nAuMNRnrm5bsnrDH/Dk6eDGIhgkWPuwEDBFd7HbSacZtDMpBBCbA
O4HTVLf7uE7XHsQRBOt0RZtaHS7Nm3F/h3nyKKjXptcpuin1TqclTcce50O1s37XjXpoaQlSOhE2
ieHG5YAcRNSUHnfBffyyzxm5oQaAsiktQBP48SiPBNYbIM3WWdcaVzOxZjqvxVRXQmRLZh22chYI
BzglFMZj4mxUHJs4KbmCwJChA4hPTehgInb6OHtVhuDrquqHViuaL29wyVt+g2ICwPHo0efaAMt1
/m1BUcxqBjvGyXvlwGsaHQKSJEBJWFXRgE3oWrFqLtl7TWEvF3lqSeKm3fRUfwHN7LQuq6mBGh2M
aQsUHOqPeaxAycPYtLa1xb1/rijrYC/b2gQXV7CNeaCXo7WRLwv/1dH+xzUsgia8p5xGVyhsGJbq
54VkM+TkPafDytgwGjMUhIvOjc4IoZPadTuoX6Z2MduNpqKoVXwFgMi3lwIlM7ZaFOluRS5Ywl1w
wrD1M6NQOHeysComAwicvSnaHJB26+q3lopeDTda3sndGnnEaYm0Ms1xzCLrhqb57Vf/UXsfzvxa
73MesIJBCY+G+Eo/UQ+kCr75QMgu8Qrc4L0IYKL6TKfzYni5aQ5TjHDlFUIOqjDb5F4NeSu579uS
BLgxnuSG3rhcgxyI2oaLwy4enjLazMYn5RonENVAA1dxN4iq2FOCgACuCaH6yjDqFnOwPfd2VsqQ
ksONcIfstG2zujkis++5BdOojv0uP+krKPHgVzgQpCgUS/HhxfQ32oBbthfdYLBEpoo8TCklSCby
Og4yUXrZn2vB/NSKJxttZGTQNO2VuMNw9qY97T8zBxFE5nqQVj89YmleMXT9V9WtzIn261PbwoCh
+F8Pyqij7zFv4+/ZbxjNR51KhRMCho1dlmz08Fg3GKvgDTLT1aBrjmDFhWseMiFzR6nNeN3sAerm
8HUXU0spBxjuWH/DpvRQAtogz0RyI77JOU/Q7FJTFvWlkymv+aFGJ/hrqfbp0y4BOKZk3UyGOMpC
SCB/nhQmo+cWoDimmXrFNZZJ0gXtUnl5OtslTmyURTYZlFp4E9rCxvF5VTtG6fyVzEIs0JO+SKw4
6wHRzg1U/2P6VvK9no3f2SePNPB4YeuGi4li56qnuqBXjDq8ooHPmtuD17BewuCUmRCyChDMAn/T
VeSnkg/qiGnHbkY4I8JxNRpumxgS1Ft2dl6F/ja0MMowOG/nqC4T0EJCT6c2X3tXE3Ozz+DSzXWS
MsUKDg4GoozhXkqVxHF61qGx2rDFb/8a1AUjB5AqTQzkeNWhrlEjyV6i+J7oLxwK3FSaRk5Mgu3/
ilzBbqtwd85qkqSgUSozMQF6x+q82uPsQiUVL/tg3orqmt4pQil+3mq6rPEBgrOtSlSgngQXEcbd
gIPzc24yOkbyZQK4DFbRkDeL6raK0XlqE7WzsthXd22N62odceNnWzVq5PNTQerPg396GXbBCR+m
CKgZq2KMFLzVlub0xuLevZZuzXOrP6I+LG5Cx8wznmDkbXxf0QKmswms9CmIIXnmDn3uIkX9Lwm7
0votSTT5eH5xUfw4tLZaGobCR6ms4f6r8Fh12ey5L7SF1b2GXCo6tiHLrxCBotlk1/pDl5N9d5qI
2NK7LzS0bYoopsbmoTdimM4aYVISLxanCi+WJoW+eMms47yX4P7Oc1vO7SAZYEgN9dDjcrO1RcOF
1QaqI79vHf+nEO6iJP7YIXM0GAFw/eoo9RQ8pD75gqcOEvATJXEJ9DmX0la3Dx456Pd5zNiXMvOg
LVjWxVc0x8LxGIyWPifebmGvvBbW/z7erINCaV5xo47sP/SP8vhg1HaTQXnwH43RCaLlICIBLkGw
YNW5E9QwMfT39io6eM+34zW5UVHuq2+hG+XH9ylBFiNVJVjEfaAIn2llq5CHcJ1MdG+M39Q71emi
jYKMQQuygL0lQCLl5nIOtIgQoOydAqy5DjI/SSQ2TXXmOBq3zhm9TCHA+BXUMlL1MS7vUypQBTNL
+n2DzO6bP3LEd9ZJQIyFYnTRyOYTS/4Vdo8v/iheSXQCxflc6YDY7zQZsuKJWHU3O9Sz9D5B9U2s
5DzF7rHwz99EZUnr0WlvWz34Mb6szIv8Xid2GWY+eMxdyTFkZqz6wZasd0OKFnCunyzeQsP1lUKS
cNVEmVKp51WJ+psg/YJSDcvxg/2M1pbFs8c3ohT3imVitkPg3cbgo5zwOijoZg536s6kDCOvXkez
cPfGEK5gZ59yzPhwvBPc3yOfNEcRVr8R6crjDS40IjySD0o//mDXOv/+6YfsXJLXjdRtnAD2s8z5
do3DBHyJiYh6eGrC1XxPArguz5ll6dnBpCPfnQ2Rp4YmPR63J+0m3yVIH7zgM8KmJHCD57cFx6iC
bdoVfO+z6anUlMXCt4BBjMKM02xSCfTXYoLhfUWy4wy2G9sn841x3zzq0Nmyibqm/mRouuwQKEqs
lj2xZYPtQdwGhAraHWEfwhxaSlixhr3q357HT2C9g/D5VZYF8eVTVMgHSVPMU/knnqselqVsLSht
lzJgz7ZXlqDMcAyXF3gYCKcI13Uqefu0oEKzT4+XuzAAfBS/4gNCraVldzwfc+Fvp/shcyUt3Bd6
GXGHfRymx2eu1i5UXmdgyCwcCUY8+22RZDEm2VnnxaRvblu3fLYAg96DOopCfURCdSrzHcyo0I35
i6WLsc6izRsfexhISeylSnq+HA21n6z8qwPiREoPjGVi7RW4dTpvP1du21Ynw3slkftxLW3gXo2k
7nHw9GgtqrYKtuwyprPXMRTd+RdViTqd7plaN6FtKQQBW2Jh6etOVW05ncC6RbuWseGR+9AcXjYt
gLYOmFhkneksSmfTeNq5FU/gErQRMNE6T3IDhWSqlOW0DkWyYBu6fR/9mqXTZF8U9ODpxKgS0gRX
kZosRgv8zncLMSeIOVngPl7e8jc3DbEEtDjWGJuSOveiu/2l0/VyucMBodQ4HhitV+YV7jl6XMXD
u56B3T2Sfzf6/LlD8TweP3cSpeDz3nCpcpeG2G2bWeVOASZ3cOek5IY7zD0xHa+LOiF12hOJyqhf
pbkYjC7dpDVLiu7mZbXJQ2tQr0o1/USyQ3Ifg8Ig22X1OyAIIBtXAp2/0GC8QZpBDpdFEGSj4Uqx
NZlH5YKt8cQWue8514T0JJbtkh/8s08Ga56WO89wUcyOyAaxL5wn4wJMvh/08CqnPdg6xjcV7Nsv
EQ17Czf7Ty8sgi5I7F7b9ahesel7BbRaREfo6mwlZA9Qq05VKG/5Jcj0v2I4nrL7FFYLICexmiSM
SXzS9zqzv1hqOEmexYE1OZNVKZP42skS+t5rmHLtaz1EgAxlUn6HEOwV0Poq2V4SM++7CBZwtzBu
bt/dkTnQoEyiBtJDEHJja8hHihsEgLEA//NQuuGGAGPlRi2GVeIUsIvatgwNCbX6WxvoSAjH7B49
VSoTQpPztVfm2H5cbBcz7IplHAsVD97wIjiNdaDET8D6HVNRYRivdaKsEfE7JKhjMXzv6rhSYzn4
aLro0o6dTXlC9ujsChYRKfwE1JLncx04NuO+5ROhMXXSW4GXlga1JgW3Xpx83WEQGId49obHrhil
sDlEVV+dgpeS1n1avChPGrrOHUYWP6qq27QYkgv/tibH3F36R7peshx1v9zT25RrtEiQZr0S7Ryq
tU4rKakW/QcH6wqz8W63phBQLWH6z4YaDkf1spRHHC7l5ZPLHCsPjcTWkKgTvdvfzvP3uIbrWwUu
bTt8KC6EIh12fm5N5WOqnuiBOxWvDrUZ+2SuIYNnRwjKbCYfYMxWKIjafqSNi5ww/GI9oh1nqIho
lw2QGVWbwJZZBiLUIncRYT3Yy17BhoFIZH9G5AZVhAytRmtHiBElomBse9xiKQsndlNHc/vrnXco
hm4Jl1GGpYN9nmJkcsbmTIIeQ9ERs17c2VKG54EhAMckNjy+dz5PJdo+IO1XLiIby/HUChO+jMxM
5RkKETobec6NxDtmK8KgX3Sbq96qhWSlYRL4FV3SfQm8XbQmoI8r2S1Z/aZvgW/haAPwKEf2oKsv
p/VO33/yVl/eRy4WpJgZ3GnWdEb3+P445lNb6GgmHRgcD5PYqYCX61JmQGrgzKy3PDSw2REQjpN9
FeA9rDcf71sjk0U112zrdIiF6lSDA3j23Vy5D3YlZoKsC8NJDlzfzJu4UGjkygOELolcgAna+Km9
Rg7yO8xFnsuKpSovmYmHtQOy5dZ2H6fdxR4k30QkPRL+gOYkECOeUQOuZwYtPDg9fY/5h5kY/Zpl
5I7Qiiz+26/8h0PJNW3e574ouRCYOcgyJL6FACEiS7Dc6fwl53NjdA+TwXtsHXYu+zbel+K631vo
sSW3uKpbzBq2ZrXmMJA3wqO2w8QBN8A/F/DYNodmDkEZG/LtiijIo9nmhNOwtVAXNay0cmap84Ve
MQDAt8sXY6vJ5pMs7QgHb3vNHjovPqsdHhW01STKhiNmWZkVRgSjRdCGAnOrrL9H4lXb+KUn9mdQ
89Lx0rNZtflbO/uKI0Se163fGpDZfb52GpBFNd0E20t06PIcQ2bUbHDa9yb6nTlXffCytSWFrJ2e
arTgte99kLfBs1eT2Ug016fR/cBButx532wq41ONkVtXYwQN62t2pgRDiEwHmWHKcGJnbcrvYjkK
SFqi4oRlTFqiC+iQrAhaKWBMF/fmPMtyrRVDycBJWkr99ZjahAWN3/shx4k7iATY38/Y7FVdmC09
shMJHN8tCtgOMHpIkMvTjZSRaXele4yFPMa+Hsy8+ZSamzj2DuHxGLyG61QcGR6UswWVAZXWuP/t
8JJ4F+swrZQuYBM/+Wo3Q0/CmuN9Hl7dbOs0Fcz892vWkGu9zP9K1aj00rWoX26C2B8NL81C2i9F
jJTJgKEBrUn0QT4MwlZBhgJZVMgDNc1v2WVwWfA7iDivUxGlProaDg4JBwwAvPZ5FsXbdtGH9djp
6vtogix5MUEPRKwl4dtF2TIdLHQ/e6p9IQaruHErnSRXPMJ+jjCMUbSzHeNsVp/gNLPW8Iu8fJi6
ma/mClPxwjQJ4UBU5LzYk8I3pTmW1M94lgXrlJ1qceL17M3f5JQgHJPBS2DzcpYnaKc5iZ/X/LFX
kQ/7rKl4A553nMF6YD4O5DBvQoqLRuK+SPJske3lJsygWSYudKQBMx59RH+q34jA8xx69lbPhveb
zKxyS8K/0L2zSg6B4hncbO31ccHlyBp5Ln4nuM0WFKukGRsDZwnaGrqXZP2Lf4ThKtpuPhk5QQyQ
161QcFNy5mDeE9VGculUUq7SnrhDrZu2JkBzIT+8fCiUk/iR7GX5+qjpxCUuZGCG7v8HJL+yVLbf
92XFKcYtWztMwSz1svpZ3NWAQmKEHh3khelTNShwK83CbSxfK6oXdqG9AR8SEWNTfYcL2nWkTJfR
6YiDEptSZq0Ifwy00/loMFxWNVOZBDRKyWomdJhGx42mtebRtHqmwLgCeRKC5cWFkeYOTBs350NW
2tImLrBm5ulvfdsKx0e9GzuR2WaI9O/Twv6lOf9eAdHu1aTJK83GYSNqPjACo2gUHmN8mJpz0Bci
5v+h9Z3QU5BCL1AzAeDpwJasl2vH8IJocK2ZUdkVF4WIQXlMv2Ah9vZJt51H/Mw7QFvKsAuyqJ1g
KAxH40C4GiIZD2skZ50mltRYgwvvqcxRiqwKG1eNwP9emcVrb2+CuKKfF5VARP3dj7yF1vOrXU97
o1EzxBiyq7rrnjc7nF+U7PvCBhkH0CEPXViAwldFx1w3UpYzNSm4BQe/Zm1zqit0ZxeGBEDYPo8z
S1N2b7Yx194Ls2AgZteusCcqVW9HJHWFazFioikZ9zNJKn5Ce6tUSnZhPSoK7nbAu29AOc9wAPYK
4nIIQiYPOxTyvYyluSXfoZhkGeRXwsfDpDRMkeJ2+q7A1X1QCuHhmO/To7X00kNZrRF250zEFNhg
qRloxhAr9SB8QGXzc8zurabDeXs22pvasjpvsUTRneK0X8HWsk4T2w5HqD0kiuMwWTxL2GFOS/4G
do4qFNXrEdzGGqgzM4+RP44qQH1z0LKI7fvqnUqGkDeLcT04qzbAOAfivr+Qbmb9dHkzh9aseby/
I+iWU+rutPTHecmwd1uCQek0nSQ7xrjctgCHvUiDSUUCEvlmMKl8VeJdInC8/pRIMIz7bEdybbW9
c9GZGTz0qhz7IpqBZVxFQC7rOmrScQir6y0Tb/lICuLseSfgZ7TE+GzAKwe4S9kScYfFeR0/Kd9w
5cpMtIkvtWWYxeW3E6AlbrTnqDGHQtRTXjm9P+Hz0bo2vCRDvc4fTKQD0WqeKyzPABu7qUWfSyMy
KX+sSvOZ4MvFCTq1w/h4aA2SbEuFb76wBLdvkm2CmkqMexXR1Bbn5Jvxi60pQ6/uUjm+Gr02K0xU
tfvQRqPPO+NXbO7plLX6HWgQCtu0c8qgWeEGT1RkT98b9+eiMYAaxCXY3gCqgWHcp/LNMaAi1Gw3
WUDb+fQspQ/RjkLEbmNhBGDBJ8V43JbTtazO5Ef0yfASyGdjTYhd3kp9QZGkSoqbsy0PYQg5y2eh
e6KesUcnDOJZrJ0vXbc7hmXrCyBuTkG6cJBk3XoZkNd1iZFkQFjeCFu7FsMSkNifI6G4SPo8Dsoz
nHtrcuOSuJuYCzn8C/FyTlRS2IlpdRqLM/qwc8FbvPhltfVCPZlfoOyuHRzqfeaqriQmzWlbulxR
VN0RAFIVw+vST7QKrhFfdJUdkRbvO8xsrsztj35ariypKaYhaHvKkz0bxv2HeTeChB8xffYkYe7T
n5gm1MbxXG3zs3B6iuxzBVQrrTlXlufssGR3+lekGJBaDgMaDaZt7Htqq0ccIK8sFoLbpufRNYtv
R0ABKsw9DQKj7aQG9/lIjRlWQZ1MwzfShpWxlphUdaSJWW8afMG21QrLs0IFpWona6cfmTESoWzw
IKLTG+8FT/k3c/dtc+POGuWvhyabluSfuwAfCcZESgyH+DPyJ9KY0ONIaYhOe1OUN4sL3fmbBZp/
etj9YXOZBW3qrXBlt01etsa5PDY1tbXHk0LgmHVIHNmOHzNF+JxuVGQ6M82wm3lRc9MCvEcyMxEV
c84yplam2groxvoM/QaidiIoSTWP8ecAsvgatBmWbh8LpBsdwjLLF3TYz/ri0Rm94o8HI+rTjX24
nPEYUhzldLN+jQ0i1tJEE9cmH4Ga8y90aPA3ZPlecMDBjJY8zR4vQndq4+iXneSraS3fiN+0yS2L
7de7Vq9L0QJCWpGTwy9JVUg6F2WGAbbQ5cp7UyIoVGqgKo82qoQjt7MWLC/K3Amd2kj15na68k5H
r3PUI8y6uvkmhI1gc2i52OuSp6B8lKTRXZHqZ2OMf8nc78xX3gPk9oEQNv9Aq/knAk0AaTOQ7zRW
UhhTCUkPOeswFJK7cIzFViJVaF7/uUHkPh/bFSFkbGdhZKRMCZPa4roydwqaSyMS9vzgnIWsXm3i
l42pAaL0BtstNyHMrnJFDeSL2JUp+6UUsNkveHw9OIlbRMcyZ2OKGV0V4C0daOCJo3uBJ8HJBn/5
cmUdb1aV1+ikm5mqRdbOXv6sY5ASyZhbDVSJEvmFbUe44tmH0F8scle91Oy/3ktK5Vt7QYWq9O7j
55ghUBNZGaYmiSujG1q2bgQmWalMRrloDR58rZOeuU456C+1onSrNC5Iiplq9d9HPIPp3ViS1aMe
KtnuZTkZDwg/HSiFheW6QUeLDB78/nU9t1GCVeNtVTTLZ6RhRS61CHZ4SRERobf6jRuE49HCpXSq
NaHVc4Ls90cdDwe6wYc2ISfNBeEFF/6/IL603KMkZuJX6VW5ADVqY03frLVfVt7K59v3E/Ji/232
xvwLBTDXNxfkts3RiU7spu3Oguoz+u2UwduU32ANAEm321Dy4AF3Us41ME94n+Eg+mfTeEp7l1nn
XNsdEvJBmIdCHymVQmbn2H7D+7fxeJU09KWbYqXlpoWENetsIuZV+w1K2QWfjhJ1OwlZONabEfOB
vmNi46NdPf3e5pYoWb5idjDvgthCFoVCA6Kc4jMKrOo2Mwm81xmvj2qIu2I8ABMdI/PwAbxWpSWI
n9wvfp7Dp6fDw6UJOPPeeqLllLW/4etUs/8nHfsuNDCNpuz//UHlQoyp/58sHPVzN2ckuWvsPRSh
Z1CkHR2KvzrNSLZoNJd4snXfL7aIzaqfk+/p57ULV6HFbWX9N6u5EyWhYkq5LZtczd3vXqaYe8Wy
VwWjuhb/KVYcJzTb5qe03+s/SDjhWt+b0GecK3Wu2oHT9RbEoVlq/WaTC4DKyPxKVoevHka5c/OZ
9HIb3v36GgljMYqfIzZKmkj5c+iB7wFxrm6jh6lYOK2GDQmiIucS6u8GylYwuu00l2sj1r1N9qhc
sBQrnwytlO6+G5k7X3bo0GwPJA2vLf+GOnC0Kn9JyhBkLvkhe8W4WjJdJLc6wfTDZR4MN0dcGrcK
6tih8UlevwYZB13Q8you1ilE2FGgbzdRGxkieo5Fhvy3CbVrOfPvjIBM+nehZLK1j7JWtn1wWOz+
6TCQBDiifBjdvY5+agC/o4D7lsMV8gHx6v9a3q0q8Gc+RBWqWWfRghCS6VXcKMPlSSMBNpp6fq60
GW+WD2F1BGBzZ+Qy5AmPchj3Bde/mquwIxmfPZoOdCYNKoqEU7hPRNqhfwXTP8tUjMbG7NCKpv5d
uf8ZZgtYnNFZgzGNqA+3cMGvu4NHvlT6pfjNuQNW8ZG9MpJ8nBO0o2UnMUCqPtSkxuPu89JUhlao
BT+a8aV0GeFX9QCK8/Mpioib/8UWQHIxH+8iLDG6ubuYWwhl2jiPQ07r331AwHgHQdRFowPUTphN
lXyu7akwVBnokcuskrU3yEj21+BTTPLrd6dGj7OJygGvOGcH3c0ekLKFUGDG64U0xchc4jSHHx3E
ilFCL2A5xqNV7Mr5MyR5+uoSEsGB4/oGNdtXoqf72B6Gp/ZsigU5J7LGyc0kJ1YG7qVg/ckuZ3m9
fHSj0N4XlvzQ7kRqv7EdTf0skoRc47lRBiQ6cEwauNvFXlNW7UbV2x5fbx2EyiX+ZZe54z5aTNaL
NkxC4REALEBO5DSSC8sMq/C3O+t4p+vHOMrHVmjetRe3IxickQH3++Sy31TOWRrw+4veHyeyQujt
UzExhN+OOpsnk1qOJFQepIx1sGLOX2bw/0JawttlRA/NrWXGSotysbZ2v3NNrQAFqJEWSLVJ52Ee
c+TMW5leL8okVSYV6FrRbJ/TPtXnxPhWnXf1FQkQRg6dONFsiAEYAWbFAwdyuZ6WYqiczLOcVhlS
qlEdCEYb4eioMezMSjcfUqOBGwPsetpEttsaow/w1LSiw7IS6YhMRsYC4QI21SRr5T1kkqcTenio
e50MzNtXEbR+IG+YAHniIJr79EAfN+b6NCLNDDrjnct+m5QQT8oEkd5iEIzfF+tbeUGmbFu/sK1E
9kY7iQnrZuT+jNOCgTBvkuprePKxM3z7lQBQyrNsC2Az6xy0BKyo4zLWhjoaJNthQiz0OWZ6vNgY
IA83EE9soUrawGTssOYgsyFCLh7LuY3tg5FnPKMJxVi9AE8ZuazATCjx+Fs2uxwaAGOOQU5SJbzZ
VKx5MNpJDh9bEaU3+06EUHAB/yywMHkZ6DA/D5EFfyM61paAZf7dhRbfx3lJZVzGx8lzvp7DBkO6
rVo7C2LaHsPxEzewz2lhXiRmGPZSaltXjtx1oMdbWzuRZKKnQl25Ci8XK3pARnm7IPybsfTULd8e
fGV3ldHW8ljF1njCQmfJ621VHrex5D+KKu8o0/FeeDf1wIx/skXbXWAExq5HVNqXV9ScVtF1+YO3
1uFuOLeS73eKylEaQnG6gV8RD1z0gQqdtOB9daH+Ujh7UtIBU2KVvPmMRmormqRw5UEUrHrggxoE
XXxSTWq9HSxdIM2dTxUodR2qX7avsMazKaz9wSLjP1YmiXdB9XOOYBFXj0zdlEzxzN5xHP8Nzn/t
tUId//GUh5ISfXwWy3gzxkxupdSyKQw8QJu8aPPdEHOIV1ggU7tBGLYB3XGBo8ewJYvJyB+c1mFJ
WlBeagmEAJlpWp6nkAMrnGXgZFpaLhf3AWAVgZKEImz0AISUp2S3EdCsU92WQVlyd39IVrKWgh+U
AA2sNVG738kQITPApbIsAGL+zpauKNp8J3uay7VqZYBe6UrdJsv1bXQRRvywE6W0WRp2H97tM9aV
Ag59kzdUprTaAZQWGyz4aHWiohmL+FDEAjpEUbWC75Sd/AL/jsK+RXe4gT9TH1nMZyOg1KmDJ6tH
1WLtjtGLuip+alfpsbqVRAeIrFDi2/ghou13JOlUJRcUphMxvbby+n1qAQeOFCDmAQgtxNx5tBF+
4sTMh7rZmaJ6iVCODf2GHV/LIGDcglNqPDREgvZPAMDCRs5KXot8MRswQnozqWOa4Pbyst8n2Kir
pTPRzn5arr5Xndn1XN/oh4031zG7PSXVK1JaHfRLTCPueRch0o48Wy0n1E2kuzRN/XGIS2crVhyK
Vy4ZY0cwsx8wuHFCtXfsLnj/KZKE69+EPRiyxYSQPmwwnONymg49u1Zfevptmw3zR6MX6eFyzae5
9FYX42tjYfOesKbEzryfFtqdC9bMT7+nWjvAfWtbrlSAvrAe/whbIbWtlpLqu3Nb9OkWB6wztTP8
1P7f0MSXAoqwiCdHWn4oYb3a4346xtfbCtS7nzx7F3pNqusMaGkufiZy5Btp5aF5xGFmh1d3NT2A
92dg7JihcdLdQMpphNRDuq3M95nlUb+ZZ93ifsVYPYbq/f+2r2fyk8PUZBfuX/Izo0i3xwFsj46C
MjlcW4ncKQpfNO8HuELTIsHSMY2Ugr9r7IR50v7JHVG55/FnYaivFX2Bx5susXNQTUl45vcfbR0c
GRxuMOXku1D+1dz0WfzGYfO4IU4X6kX/+lQNg2uy88WAMwpsb7Zgi/KH915TxV0L3wARSLMAAw8H
WKCwYn+TACqVL7AdnG5cJ+rYgCGjq8tbpEusF3o3LV66CNgbqZhkoNBRNSK5R7JRV3m1EdBQRlrM
av365JfX4vwtqgw1ZKA1cNkUFhIVN5gnrqE6RNK3GI4t/BwjXffXNQy7p+lrA4UXKHU5wBYkRZm3
fBw60x+fZqC+vXtFd6f9arfXJ621qbs2flmQwJFW1ZJE80IKm02SRGGUQXzi/LhaVMZC/AZOg0q/
Q/VAyp94I4WhHBUx+nGjqHhw54fHHGfojXum67AEq2SS1fl3Yq00sDZMs3tkPQZQ4hM0lCJ7VS3O
cD+QKPir1LpzOveN8bD9UdCbZZTbXujxN/JB0a0trfOBP/c03YaBwZTA3EmDqiYCULaAa4AQyuQ3
9OUbP78mijH0Lf7JqgaMclpfvIbM/xC/+KgTVxq6HaLU2eVIbrBYIkevW8Hc6w7JFboWdH4/KPKu
A8Ry5Cgjxxrmh9tsZjbzhWvgEg9xUy5jWqeewK/i9G/XklC6ouR5M6iiEzqFJzux53znDdNdhHde
HFIS6MYKqjfAq1zMPiM2yFGSyo7K+z0aE1MUhUMSMe+caiiRGle32wpsrjLGeM9v1Dscyk7ZS1IM
OILyGstUXO3LI1k9t/tLGKGEh4GgYIpjMpZEeyp3/t6yA8rlkPXRdgxsWgCP/P8hvdsuXG77RIzF
6tuOeKiUTBVHV9jW0faDnrOBbGYYl9VWI+RNCSFSS/VSo+E2iBtV0BOt0YL+jpJj5T4dU3l+7Ds2
POXxIHCNWUmcb789wvFtonHUmJ3c/gxOPerog5YZHcnWtazDWbe2WDFASyK8QK0b94kocMBCAFwJ
Q19xsFCI1wIhYhBhwAHvAuMmUEkjDtxvQMp2SgfqkKKVUgM5L3u9cffY/v+F5CXjB1yF5YF1Uofy
zspsMFh8+mhTYTS7mHmqZUebYWROFPKrF8sSWjeh1Ei1CoFDnfUT3Eb3isYlmqiQqQs+xrKUCrZS
z/r+BazzF1MYO1wJDIzpHEwvLcNvpZ1G6h8Wf48/ZLr7uozkPXDkB+J8Rg+yXb33X+R9MQUiIHlJ
uKWTXR19f80bvsxMpD3kndo1mojAfnr/fFmJE8FQMJM7TV3VulG4JuduG7TySY9WHue2H/ocliAq
Lliw21q50mLjaCIaQKaW5xsNOUrZFEgnp2NrKx1vN+JCTQuprSFZsfQUl7MoaufX5bbWsiuE/bL2
6vKSqcj3GHHLsakSxDhYocl9DAu7DGffob4nDl5o8rPvt3CDFpIXvsYvbII2AVgTe2LR2o+UYRfm
vIJDPkyhdGjCrpP85H7fWVfQpb2HTFDFN6OkmGkPiiHQw8/XD4CJAXzst+2ZjIcRyOOeuDx+nfwX
gyNTVzryImdv/cPYy3gvKerhA3Ef9QWIpIAxZ1RHprHFGTEF0ccO6ht3nnRsJZN674eBayJ+1+/6
E8D0c0sKWocV539RfYN4/Z/ZAXteggQozvivXdNS+Ujo4DdVYIOkWtMGTcGy/4Y0ylzW70VjZv5Z
JCJJkE+2BZ+MPgHBXJNl71eTwX3TiosX7bv4JXd9zk9FlPtueovLRIJVBXMFtTjlz6qxgJmaxcAP
IfuFI2pzlXhgdD0zsvyRrpkuMVqTLS3oMgHqf3tBFLKj7g04uZ1fb7BfMn4iW9XrQOeWnItCNccv
HFveij/AuyFm+rcMf0H2sKUXqLYGlte43vlKLMwlxKIDxdz9MTGBx/GZdsuI87Oka8gS8TL9WGfe
Uwo26UCZq+IhqG+VdGqFfRBC471F8IovFfrsF419m81CDFwPS7fjIfZSj0nEKHes2/TArLPY7uDH
ENTQ9Dg0i8Y/GBVaaIa2ZaG1VZpoVJQMaQErcg1AUBaTiY6L4SMyX1ab9mIisQC0Btp2mv911U9Q
kNSV5BrTQgbWtrS392bb3eDBbCD6BTfs8pGdtTIZcsFukVLrLpJS0BrbDkpJ/bbVNd8XBGxGPPTt
wpk2Z0BFijZOG2tCPf6o79EJIYtljPabPOhqktBA+6qUMooaxyNYDHNEKFRzbfyber/qe7v9BBfT
tXK5Ao7KNXZgq96WOfr/K/ZLoQ3J1mlRc8wDQwAReEQ1pcVXFccC0pN0/evcOl6eedxZeOXk9qPC
xO4yZaFwIHeFIUHD08N3ngakdjF9lpe3d7pnUN/D02l7qdh9oglFsvlPY46dgxTyf0241Ese0rCA
Cy1bznMiUtQ4p2IxHS6BIAeLcRqxo3t7wkGrv3WqW7+TTmLGAMx+fvOvDZO0NN5wzkBAjvsIXnFd
kseXkKHKsRf/g+eA/IKZk49xCOWDKkXO6Vh1j6hwSKksP5BbdCo1hXxjZIXQOEvLSPXifyICFK7Z
QL3sLynNjDhpi9r7dQhku/nsOXA8APpuUkBfDiFG2vOU83IEAkLvnSvPaPpM8c/Ptr6OKNbZMsG0
xMKmc9YBk88rTGgqiefMsot3SoslnPONw2+pE32g0AyDnjF6cVhVtQ6jP0WPGK02kGpcbfKbYaHh
RFVKzbzdJk4CYMhAbJRZdV/ABgtvZ29kDTKBv3nwJEwtnqquMauAQw7JEeWS2+7LwULqpKt7Kjms
W4MUVfeBZeVmNP/NhB9S/OXSHuB+n1ggXJbnRXs1V0hwhDP8XVryV7/QzzsnZvvZ1rTQaVQ73xYM
9YkepkFHS3OC1xUhWOqfstKw5aWhyAQ6jreafis+d64yAKwPOWvRLbNbtg5LxLNy+paY3wX0gvSV
OWNcK2mpacM508sVveB/Aycpd1G3Mq1JZlhugrQK26Y/usPFMfhCipoq/DP4eJ4NyJ1AlHOZIrXA
p50AR+KSqMJeRe+utXrO7MrE7mKyj5n1ms3LGfa+17dijswRlhc7+Pp+763aIN2dJm5nmL5nMHA1
ISJ6XQS3mZFJ9VvSpGU3jVNdVkIdC4lZuZZK9cqHJBjyDdtaIsypwyoqMTIedesdyoectd75UdS1
dDRc/Ca1cI6fFjsES4B3HBN1c5s0zFnApM4kr4d8Q3lAX3lD2VrA/6Nc4+PMnmFDuFbkIPRRAPjw
7MzR6579xP1YOY5obnyMe2o45rIj50fCVJvnOKlWUtQc8l4UONBnbXU7Y6r0pbDfAS53nZ44Q125
kutxjSw/POb/vGOVEms+C3qQGaQlgCQxI4PxgLINRNvrSbix4jwd4HAT0XfqTJ/fQM5kgf13aZis
H2mMzgLGZ8NMW6uYc2fG2xrSYZqeEeM2GEfrUcxprceVpg/wDqwrNQ5fj2z5p6kQvcXBhcYPWFx2
2+HvZ0fgySAecuBZG97j8W0PeV48W5bBNYQaIxjHItdrDN4BKotQDiASM4v+Xpw71idEWbi/nOGw
WP3NCyBC+1Xlo5DDVt+1xUWvebkAmZIjP0j2XaWDYHdd0sgiX0ugxP6q/Iy6F9ErmAETXijccKcs
GMimyoV8yN64pWtUKHh4ZyCedNESwsfQeuKgeNHFtIt4vdgEuxOFOcdW67ZL6aiqCKZRrH3ylHR6
v+x65Y9fDDmPfYxFDpFbX8LNToe6e7WjcuzXX4oUnKEaG092VdmdHwWQfACEK1kyViuN/Ys+EQYN
ZceM+JcxYRKiX6U9VOesYnPUqPvBtUc0TFfi3LRdw/+w0eT8QN29zBbKy3RB5T8zRsKlLm/XbwmB
cYkfJQUQgtdPUuvnpk2QeZ17Sxi97zcAIrneg3Q4WtVQaejpivp06Ovk2XXwN/C97rdM1B0F/AV1
fWodfHVX5l/46Dm25MncItDCFDCDMCKWDkIXmpjaZ8EQnaslxVVIHrVxAJUy2OuIo7BAzttTTQee
/4Ac6ij9teVHbioWU6V4FclAJLDbFKUnmAm7xWZ9hb2E3+kZMPKFK5iNlcuinQ2iLSQFulWLxbuH
9kfW2Kd6mQG0lcYQj/tdPAYl6O9FDMFVu35pgQP4+stjCuQDovS9B6ZMY4MmWqiK3gPsLNM9Ga2Z
s5XlfKKLDpZqOgyzjbq9EZkfSv4I4bIQVshjdKB+YPu5Bin6fit4nj88hvgeuHG+5q7BSjSHqWhM
Kp6+xVlWJPeHOpq63aYM2JGpAVk3+fIfywe3UZ+wPh+Qu7Q/vJx7RkPeMHeT/PSR+GPWUR8b8dAK
anWZ6UOvHr5DMwCvJbg1w8jeBM27Uj8vU/0UENBxhHRyN4a1JJMi23HT3djq+6lQWIL0O/gubbhI
4iI7UzCSVDYkJWykKLIMv0/QehiC9lpPrhH5DXFrDY7/GF+lCZaOVPdpexVEVZr1jYwas7EpLBDH
GHsvfGgtPunp7Dy9DHaRnpucAkEUlXH0kiwzP7dJ1A/9f9FnMGntZEXQjIkCzh2OhR67/JwwfbCi
r+IIZy5tN6lGlbGGD6/FjIbru72pb9Y89htItiDNWHdmA6SIhWTxnfE1Mvxzne9UJPAS1hgcc8eB
Zqg3CiaFF4JZQEj8Wo0hfNKcixgnDkzkM9NQBH8JbXadgF+lRfVLwTjvjj7x/vqg2/EbgMu/fQ3x
pWVifNEqtgYX9yBiH2VTgHRyNrBQHKW/zqqD+rc39swd81cI3JuepHkXFohgBfABuhuAooYNHt07
rCUmWE7FjjFmiakBwmV/1oxJTaDaVEh65eh1/02QITLeIvvicUxgDiaw+IZ1Uj68me0d5Km4hTBt
sdiGZ6flUuBVxnVrRhKBhwwKuFgm2ZM1ln44GarOnjqFwQobIw4Gm+wtrs0cUJ2Mk2aXJsBxpoRC
OkZvDNXFCxwTvEjK9WkGXG+lO0ugey1MKg72yAzMnhtDCP6+DUfev9qv9zMxKur/Thp+DBvfY49l
RfeoNsPaXoQpWW2j2ZMDv1VVCVKtl2+r0kWZNSj020kgJMu2en6AFHZxiNrrs1xB919KCuwY7OKX
e8DFwmT4qdtB3TUiqUcKmSfzRlPrgAJ/CornCkz3YXj5N3VG7+WHx090PXcUnYo2E96In0JH+kr2
76VsOevfZeHb1pDRTdgSg9WW9BYx1jen5DAWphdTe2mPBBeu0wjjtkr83zCA846hfJyWdtSHixxk
eKB8SREErlxh1kxvXGaSQN55zEaDcNZ1caChfFAbnvsUj+04uOCUKzA+YXV+23CyunJGNwBZpwQ7
0dLgYt78vXSHCOFA3/VRsVqdbBULnAeOL7LDkswigMI4ulcPyJBxacdbgcsllj7c77208GfjiRnO
2qWsjv8d01tC1JXiLvrcLPPHPoRoH/xnQAsvcWVg4ZlllqB8pzo3kwA6fJMSpcB84tO5boiRmmBo
Ah2h47zNtFOtIe7Ruc67lYp/35AX4vdSIbKB8flhgnJTVkwZt5AKaRYfB69boqyIVOCTYHhTx014
WN7cF4C7x7gcv7x8j3ijJhFMjTRj2niZC9n2lMPlMXp/LFRleYs4aFkBuojqrNZ/GkSG9mN8OrTa
ElU0K+mXNkWScx698NoNhqVQ+0G7+SOXyxDUhzMz8FPKlzMRsNwI/Tn/ZFb42FF7FtaIMtO8pJXM
ML6kHsKswafXPT4XPEmcGcMZiYwiYncIiWUURF0k1uA/YxVFkg5i5FiScN6dwYhs1+wcD6R1TzTS
qX+6qfudyaBZ/IC1MvURJLo+CDHZfxZSWfka0nWbTt+WAj9lE6OQHiJI3ITzOIbSGAx84+q2/szS
WnHIoEGfaY3n/UynVgZsaT6v0j8MmL0geL8D9D+b1TZ0+MTrBdElRGkkFIo36LbgdZdd7UqgUCCf
cDCk0PI+FGd65bL4tOOaZmu4VQwN+TupUPmmla2EVw9xwmqGV4iYshfNGHOoCIW1V0Smw+qlDktm
kZohLFBFMnzgtpDLFDYhPBBQvhynPVKRVMmGb7FNy6FpAPcUErf2AKTjd9TziesgyfWSDf4AERVN
jH/2Ld0FU55CD4O3UPZntcsi3F8sM9kl0wco+8kxUh48tyPQcFp1Nvjfich/NJCsna5xk8HuLdK2
24L+i9sv5AjZu8y1xlC2XRcL7yfM2ECb3Ew0HSaVO84aFwLPphl8GWTEfg2wQ2eRA05m8ovb9A0I
UylLksXLQCWLKrquA7yceLwM1ENDcJay30F+bw4g9tuMpFvbJ3+8nNk4fhaqBL/4D4TO9/tl7vN9
KsLY+No75SBjheZUsTUJ4jDDMkI1brLtbZHuhIOSRMF1eaCYyOmxxj88DyI/4xVntwMNeJenF77S
CppN8ph9rAYJUzpHBzE/mMYfsy/RLHAg19tw9YoIS3CxWRuZyCToitUoQuSj7383+ZcTQO0z2NAa
ECqz9mvTQYRIiR4gV2W3rhEsHLKAaMOn6XI+fO2o054Ielbq0ibJF8kiJuQcHm9GQzG3LqpyLr3T
4WvKyyCzyvhJx9slxprlFHVLQopn2WWeKAg0/76u57peU2EuEaSkLNx6SWOoui0Nm6W/KGW9XLe3
Z5vf5bZbgJKhcE1kI0GXwnt3jB03skzn52/B96CtNdu/rzKR+Z3x8vrL1n5kkGMu8onUXGs9GGJY
iPfuzykQ2c2AQ2RlMv5BwZp3ziFDPM+RCFEFvtwltOQ/Arj6KtSTlAOWcyW5NC6UUnxvJec5pG92
avjdz4EwkJ4UieIrVgq/UA78IY+6DjlaaNLMyqkCoD2MaV2C0+VNL0xhaLaRIc2vxJI90oiMCbYs
wlZlp6hc2k4wH7Y/V+hRFrmgmjWPkW6clU34OBt2sU0Uo/pc2qoyEZ9+OxXGAT/brfZ4cgF92tuU
ZKoZOOvXETe23DEFh/TuUsoZLiyc59JeYIuHZNEJGQfQUXzpHPMxxEe8JmL5okhSVul6VXOs8TRA
yAVHGau0K3O6AO7q7IWe8PdpLfz5r790ITyqjccBM/o4c9h56l46ypQAuPW5pPXKOp5EPxLhUlPs
LOWGYemVw9+VXh3KZAVW7DOLhNuyLPyhSgZL1yXfoNW1n2eCj+1hOffZOoDi2vH/9eYTbMHmI9el
7jYdeBiyTCylE7Kzqu19xctT34AOjkRo8FK6C99P1jyRAjFM4y9iKA7UjqJZ6bMcfjauxOoIHGfx
BuMHFWs+h1pWPtXVUV/yh7DaWU7ooXSuo5JBJlR2ShxFeivO+hTFXT01FSHajRTVty/jEHLO65h3
R98qEaD4zKH8zEqru1LlXxNwOj2gwDxGXYGc4JuqxdGEmA9LuWUXSg7KoKvyEkYIhM3glu6UG1MA
UHBIPEMEKh/34Cr+Msjsls2HZv4cOPlhR1GFGLbOo6JJVghGZy6dyWSHlxD+yGhW4ndBLfggKfBa
EBxxOToUDVa8WFTYLIRpIh2b7s0Ape7DlyZse+Huh8fdUFhOKqD5X+p8j7BxO9wvPYpqOMBFGiRL
bj7db6eL99yV8PZspVVe93xrfr7oqFv2vw3vGon40WdDdPv43D78iHtDSYHAx8XLIiaDcErmFVu4
PLQrS/NGl/x+lC62+SRAu64oVqyvn7DRx9rl9YpLutGzhKjnZ2tp315XH4IFghntsQlzdFw1RIjP
ZSJ/UX4wjYKOtTXmEmk/bcXNJ6QhLFtG1Kv+VUSIGLjG52p+qC6AT5sbUxSnvbNbwXdzy9TpGeUB
bWQRpD7soB4nwP+lxAeRaSr8EskHpXAd0q2LDhMVLGGegQY44iaN+oXNWKy7RYaQVMigdTJFRntg
JIiUgJ5nrmraN9aqqKkt67QHJIzPsc42jMWBn0usIKCuJRFLi2042Pkp4xDCZ2rvd0xP++PGD6Fv
yXb1gC6ymZ2lQNaTQRI1OcW06plVXX7xnq9anuXZ9fZ2F3kk3d9UiiChvfW82Z2sni+xsWo84rkR
afZTpq+63knw+z1Ws8Q+FfjT9jyfjrYsjjZ9NF1AuiiTQPui7DINLde7QtmRleQ6v22HOfc/BpAJ
AH9w75ri0y9P/eRjdz4dPfR8X5/6xm2vBqRsSbIv7JKpoDds3OWbaFfS36Q5TPtwgiwQvEQQaltU
njy3Tci3X8ZNF08FdIMYIqoHFyehDBfDpagyHteMaSguC/x63ugj3dzEuPdeMaKR4fKdFH5zPKOX
QsgtgVnHpPpV1mERSeqGRwFiefy8uzvA7LUnnAWP4tm3LCs3aaNt4/ZRgHm1mxYTm2eZm5EOwCpj
TxxVBellnnKGJleaud7qOjqfoF/l6AEGQ2o62mk/JJ409Hp41gayPkGZ2uWIC5BrnaXdfphxYhqI
5Mi8TahVtw0PHzcRJr7L+sgJsZ8shFjsGJ6L9ksTmvejPLe9mL0pI0o64Mc5bLzGPzMlaxvCmZXc
DMAq/Di64tVs6Rn93dGnz/kFYUdCcHJKz0FeVNk2A9UlTrjlmV/C5dUWox2lI503E+xMY546wQ0C
XNIrvm/TKWfoQDkhobmTGe4pZul+7JtaguT4n0Quxtk9G5168wRpsVfFwI1tHkTgT5gApfPzAup9
+NpLs3GXmBTsrdqDS3fZ/aTbtnmuandFcOz71gWSqkmxNuAsH4XcuarWbHrXp70OfyeNHMNZLFTP
yIoxbuAKPm2GnkUR1xeef9dZdCpjyb2cbRkjlYv8cj2xHkTEXZUkD9eTN6zx6saDb6qXT9xXWJJ/
+18fdrx1aDbAArp8G7Z448Q68JZR0jEDTWm14SwqdjLVntVPZ2gglhpmf8DffSf18vGcojkEfUZ0
b4GWhciEviG9vMUi3uHzAHoqDWmbrM6BFVgv0zw66A/fcOKKooIFk8k6NRWuRhM4SvJSCi12i18E
PSQqyZyCQKOjfEnB7l9FzOBpUg4UMJ15nUynBmib69LB4xDURIkomP5GIWCHAhP3aadbCegBLSG/
0yOSa/msjmUNeZu4Ehv6/UCpVQAg+PNsOesb9Zdygk8HK5Wy+Gjdm2MLeTB4caW6kdHwMHISzYcm
GmYsYfsv9bGpWiANQYhfVB2cch9amQ7ZBbMz67KvWyq8UTZq9ZIfqj/sc7gApR3b+QwfAm+m26CB
9RLmCc73dx/KQe5ruppRGApdPdm++XQUZx0+sJdja3dJ3+4J6dj6d9YW/+yYHMXEKJhNjawbl77y
vACQnGCd8VuxmeBrs9uqJvXewSIU1Bf7YXelbzOGDOePj0w0uCGYYIfp8xshWF5Yv3BqogHrrFlY
DXCIcVhtnhm8RibCNg4pfEa9VDkijf8pnucRVVn4uMPUkg/CkvoDizpq3U+CgNN31D0tfhMorZdU
8zPd0pgHEJyhw98VWtcpLLJdoIRqN/F0rmDBpX0jKvcRuRsai7q83fbiJJajwxEy5tYvSm3S1Pe1
bQWpzrSDtTxTz3YBLtb8dnASOO55QZVwiHX8H/b9S0EhxQZ/dOQkHRoTKG9MzoTMQC7GOZN/kt1g
IC66tKJt/64B2Co3zAeT5VHsBIuwora/OKF0k6zLbR7DNlWcRhPr53KXNdY/FZ7/pqqxcDJ++WFX
tPSxjZTc3jsRpc/ZonEtIcbGrQOADCo1hHkllJt0G3akvwX7MOPWctcmOTTBPXLbEW5JjL1HgA8b
MCr9pUPfmLER8BewJod3r9bZllLG1hBoRsCZ1+e28YOCkOrrqYpTG+BtrKtSq7ZARB71KxgWlmyP
rEkH7MBikOaQGwpeNVetQH+Ot9qUm8IhdLYvpZVEiNR4ei7Zb8XA8LjZYY2yotCErAAcu3iu/IhP
dKJbpAf/1I/jn75y0w0+1/fYRZfxnd0bFeVHNGuCZY+xXCKIGqTHNAW49IZhb4AWbUKuqwFDipBu
FBb0c8AIQ+MD/2Pt9i9JGztsHkpgQuIiDOvtLSOPmTv+zELDfJtLItTSLtWUs1GpimuLtM4cIFMu
bTqYEbgbcprXyfXTY7gwy6iDiIIl8OVA6x2LlBLsS4tAPoUmBDNeh8N4a5/ehJLmt7cXMlEcbDO9
5buYJsAabBdhAL0l7tt7c3Kh+kUtqNEbuSgVU5h/L7+SDmJ9K+TedhGmqOvzQdAboo5WqiwtPpqW
7twK19Cy0nonT1fltiO2GiDVbcBp2YjjdqtistEM75WCC2F1PBAfzh8+Z5ytqEdHlzwzNBps4Rwx
rZAHacl4WLQI9hMbb1Xqu5hDMFMITu6RN4TpRLCyk/TVSnkSKwPbST58drh5HY9wLZ3aRolsKLMq
1zSumHbORynlhSECzqqd9EKe+h79x02AnRraHTagXpXnG1vdAstTE62BB7E3uGJlsQdDw5MtVJKi
a7NGpgQ52QgEprezX759kuSLjZgf4WWj6G94YFfmoXC5s9tSdej9n37cnOcupor+M5tUX2VWWnbh
XeEUcD11qzGg8GeRniMtgvvnBfsxlnQZLXhRn7d4UXDswf55F57eThgr6LfvdOhbI/JdvPgS2AkI
PrONBLVK88ZVdtk2ngdRvKP9z77cc+CT1Y9qax6971YvTtENpb09jgJ4TF+V3Ka6RhMoLx9wVPcX
h/nUNrjV5bL7EDIQxJvVYAn+z40OdZku8aCUUqv6gqDwWXOVb2E+5qcqljy1ACa+3nhulMKLAzV7
J9FW2af9I+6gKHKoVTXmAto7WIxkovj6qOtApIIa7S5VfBXb0kNuoLGjGWmkPtUOvyFd/7eZCbPe
s1f/4JEtQ4hDHNR4IrHsIVhhzgA5OTqnWReqKVIGhnS+2WOsuqgLIZx4RicalU8hTq0332/K7OtX
mT9UzBRU7xTQ+UYCYwQohFB3I+jqTAkzubRdP/aFZPR9hUFLFoxESAwKNU65b7b0RswCRopOF5cs
POhiiG1sP3m8a+jJTXfCfy5xpmNWxb8dNdqMBEdHq/gORUGFi90R4bO/QYV0r42/VDT+IJQrZO8i
vNpCTlgnD0nDPpP6TXM1hB4u6irk67smVHHMtEYVyce5bRNmPUg9v8NMBFXy4HIgZjGv2+T9W5j/
3CvJsPofwqrn7CkF9burABzxJuR0PpOETqqtHd2gIAKFqbk8/Q7IJgpYIfEhZYH8VbJph3+jmzH4
jfWhANO0MxGaxa41sMCizYrI1+goA3v6xoIo4HHwRsPJ5FRpXs2uz9GPIrkhNMsjMo41e5G3ToZr
YiGPYOXZyxwllUCilXwbzmBVF3T0maAlGQeRuRg291lURKjVXi5yjAybXC3g2r0Q0yFRDkA8qEgl
J3YstvpFO9xoLYDAVhQH0TfqlF56INUeGnLKw+jTGsbFbFdAGTZLP8itwMxBjWlzf1FCiQrFRwkB
yUQaU967ySj2HbIYJix9cs5DjEGHaiQRUyGPTpDZGC1HSEfxeAE9ekyLhGEmaoD0SBWukTFcOtAT
K+O1B3tdAPoqBT0cJF7wz4917D6ZQxWGrBTC1KqA3iITI9/YsBzdGiH5zSS/ssy5Nmoeus4EMQXJ
5it226Rx1mvCeWfqd+dMA1hEgStGEzTnLGWv57XKPHATsr5kjl+K85KZWyWZ/xrQQ9LpVCqtR/a8
HfJm7zLjkrGP5R8juv33Eopgpu0qDLXlC5fu/2YI+9j7BJyBXa0/fe3qAW1jZQDaH7XIAWR288Ii
BqIDiUFipnOt2ubgg3RllVDtSRCQcd1uYzc1MXLKdDkZ2JWV0wLaJLCWO+pmVmC8lzAzOYSBCBch
xfssTeqMBP8iFjsKCWxdkt64bFhGSzPnhhzJG54o6wvj2IuY2MQ8vRkFg9Y6Yi/6bF9lLKS9pXOo
1/+WGleTi6c0+sXpXXRV54vFIccoT0erKAlVKhD+uD1QA9/smxOoRyhRYjS4eQmyca7P35SDAhal
DpChXsRxBRTaWG5n0vazOlJLCZTM0AnqK74wAQeD1ri2cXrrnWIuWjqfk7rokxEwOcpnnigyjRS+
/F0QW8ftQGFl5DdHyinPAK3swxLaKFs+4LfXaN5EdLJmdaadxSCVpERf4DV3lX62v1nAmuLz6TrJ
ROM3OFoeXWfFEYZFgX5aqxikHYTO4rcSI7HiYSMo+vtpu9GHoUjBufHgXi3ZaYXJejvGpHGvrv2p
poEJLUPX/fdiMAEFrnNLirI+4R95aGj5dr1bUME8pm8KAmgd7znipqD9XqyEt8GY19Bz/C0FPGCP
HSfcM8dLKDKbx1xJ2oUa3pLwwwJ/2U+8vk9gi81bF/WWyCHv1E2JgPyl8AZq75LKtYxz71i30wPo
1AEWog9coQ6IzNp7X81xFocE+VmvxCOQnw3LSB5hvyyHFDrDhlBpzCOovtWc8dUkcRF/hX/ZLRC0
5EbV2YvxXFixw3IdxQCDogvv0p70SCbuh/Zbewo9YtQUBOifBb01o7isC7VNy4kARGkN4IOCg+KU
1EEHVmw+asc3M6644jwgXcjV+DfyWh46xac4j6b+RQ0Bw48hT1wT1nF+YxqDxuMvaIjkGA0pI2ue
MB5b5eU5Au/mNQNJ85NfZjjeO3zaRRkZWvC7KVDHgKOe6JvLzyurF5zeD2M+oy5Rjk+IZQJJTKKg
Dc46GAa75gK6c+8HRA75yBJSk14RWlRQaYffyGvHtOL83sXtL5aV+rCnRmpYqxZd5fR3IW0jB1TE
61vPC8aYU0AUTqV+ejIRFxMGgZcbWmOuKpkveNf5amyJ274yqzKneO3GOI2AV2FxLLtPAkMN5q/K
OgO9mb5wdFgvehS/RTUJq+m+41ultJoQBviOZiPYR4b5+/gue7CClKujI9JaMuiaVhfFhuJkoR0f
ss0xHN/50m/lSoUijOtG8mmFzvHIrvQlkd4nKJy7IqlRFf2Du1wwLW8ScsHdMVldHE7JSuYEFoGC
hutGs+3dxaqXBpwWeMxRTD4i4KV/DyvN4RqSy2Pdv4K+PlBHeJkjnW9L2Ll6HxbOHwB7A2Z8fb07
wYJzL06CK1lVBmxHdrf5bWpfpQZa2IlWqo4HiAudVM7NXR85E+SSjpNDMU/HFsIbunMILXqjXeES
3zYZnhqexwNgHTUJR0VCLgcNN0lAlOwVS/X7CQCy+DFAgI10Se6shaT2ikcdpN5/LCEfUVzcGhvo
jlvp+jWY6EaXYDNoN6rGLE7hHGhgqwS/9SzDSCkvDwygrQj/zOoNz4uZ/Bu6QpjpUkLya2qNWqGG
3Mor9dUgH9G6Vw2wdqQ5IGzbHxCWLgMyxfLkdv+5kZfG/sAhIDx9hm9wqIJer3rLqq/wCjFu/InJ
+GV5P1JmV4bE+L4H59NJ0KPLXrYnW+/DoFfpIFN2yjUXmI8pojX4llHSO45gI6R5w/b57pZjhdJJ
h35LX0nq6bAyRnW1en7/xBh6mrTCOnfjZ7cd9RLHniPcg+wAODLmOTl/5GQ9GG+GdGjvS9D+gW99
OuUaKN5H1acou1/RKKCRTlozrqpNHzyloqvAUqyloQfF0XSgU1dFrlevQDIsZuKUbeUbQYyXg+b7
sn83seWfOkVeBn4RMgUZagGh7nDlcxBE9k0l+8qdanB9CKQlr2NgpWSMIe0X1/oXR8UKnTn1gKlH
yOCuFow/Fo+1/LWHrF7qd3i7yepMTPHfn4gKMMW41s3Qo6/DWFnsulV+yPJaD1xsGk6tiVPM7br8
UZJap+xDClvisjGHlP1adtLaHSn+nt6wOu5CakhrtnVVXl2TLVu73z7MQJZe4snskVKsjw7yiTy4
klekIJzYrcfDWhEEu60wA82cQ9fSZfpjD65UkAVGa/LJeDyUupKcnQYDORbkEJPzGLluWnxaiZRh
OGe6USs6lEpO6vHAi2EjoTeNYrX92MeQClxo3U9SkORHc9eB6So1tywh1nmNhOK/E+mAULO6OzC3
l4MBkNkN9a7660MF2asvv38dpWHpHOWPbvBtTo7EgNey2f/2NFy8eswJhIRiO43yCsjBfaqBMy1v
IYGoJp6vsBo8bKU8g4xV2JFuGPTUQI+UYsZlV2pIl4lGl2z4awzda+ZpIJ8SfR8IAijuzAW3bYDg
EA7FQ/H1mAMBAF4CdDHcszuRckoKvhBXZAmRXc6CgY7WSmzl+Yp4LhIc/IPFrxLvU95cSXF4G/qi
ObV/PaoKM45RpN5nr2qsisCKfcVzmoOYL/CwORf4GKV339f4ZmwOS1liBGnjLHjV1sUQSnAHSUcF
Q2jNvmcbRMVSi2rgDB6Bgf2oaSHtaq/ggoYo9TUdxZ1ZNawEeuptqikcoz0nDFj4sIPECsF6nYcL
imeOFB0aVhJApTs9w4x3So2AyMq503JUC6VCqq8fV/tFPPpfSWZ6LuYHovZZ3ejEsbXTqQLD8sUp
bM5KSklJwlWZpVOhOp6H7dZQTKAR8vssi7hUKscdywMUrI0w0d0ccF3SJAxXJAASzbMAT5bBUocM
b8gsLC70epWKKcbzfuudnSCyig62gFX08CzMLTXXx8CpDt1YQzWKorvwiNKivkefcsKQhd/GuZpu
TUe+gv1QQGISTGwqJ4fGB4ZPEVfxGueG8mvTqwXZpQWYFTndAgnRmJpqAG65FoXCH1Bn1dcPQZfC
3ITsKFMLJmM6Au1WJ+rE41ikOsCasseWG5DulkU9bBt6b7HwRWmSOTKtwvkvzTL+kJ0MB3wwwdwJ
8/n4QrkfRtMPWnnJLmwEVvREbSV17FQJvJiBhyxy/hZU6D3N+2qqbzLvWVH3O5ByAwgQXlHIhtgm
LXm/6dK7cA/LauBuJjdKm7pl6bU3z4kHxbceK3D+ap3xxWOVImvrb/uFu+azko+pkav97sN74JZa
9alItQswxy2Aj9J/+zRbUflR1bYW+cIQhc/9eZg3cD6n6KzGr6x+1FzfGB0yylFBvchkV/jqMoI4
XxHQJ28yV3blPx16Imq6GIEaSCaCdq1FC2nXQYSGX2y7LbJQtl965sssKrt2WZet7qBoR5v9dy+P
gypWBUJpgAS2o139EOB0QuEwep/M6mkiyXU2x1H5AuWDRBOmh9b/25GG95fgnwCgdsnxuGXHwxE4
a37s+xAE+ZanBL+OrhoPRpwHAAXpOifvN1y4FtRVRZifU44o0P21EJsrTM98R44UOD4z6O+CmjT6
Z7RsT5Qp9DKNXjuDbX2KRjnvOZ6nRAXsHDrD/871k69E7R4XinnX+NCJbdnSpj/lx5JIfsCbkW34
VcZjawG2lzfCr9+knBpjFjkRlLsrPBqiFRNNuWlDE2+oeT9GsqFIuWxO68iUwsizrcPb2BOpGZJL
xP2+pVLDJj7F43F2W3VTFSh+CD36v91k4MZMvElM1hXmiNlRTTCgrziVA4cHrTzfCtXWXXwOh0o7
5NAPc909YMZw5lTmU2ACJ4b2zL8Ufuc+7IanJ9ndy5LWXGKkXjYlFWS+CalSeL72NDXce0LqUxyJ
wzQwZ5YS+CFX0jfKyraaSLM6IFGhTzpt8YGEnue6eBTbRI2IaG5kCq6vxE+/SvIPc1UPD6sb4JOC
tU8MRdWZNXimkaUl6ucafPQn2w+BrGbm+WFKIuNPw3QbHdbrvx3i3Tx2sHM8fPA6OhjK9w3Hyhxm
53QFwR7EUGBvKzKb4fcpbg9u8VKYRuugmMvr/PqJwMDe52IW26KmSebhzqCrHqDMkdKiaMA/yrsL
L6ryJVofWhnDCu4PLOe+Tt5Hti5FbGsTdQaxESH6m5hPotm0dT0RhIEeTo/B6mTEORjprlvYTeRt
3mm9dpxtiVC5/WnbC5jf3Mx1giRCDM9xudHwLG3BzoC61/TcKzJOFgboHpo3k1QNY7jJD/z9M/WX
PzUZMUKLpQgVCt11Cnujce01byoqoXrMLkpGqc15aEfnENtLhv7SG+nzDx6iymynhtijKLEP2uaq
SUN67kSUlFnZbuWxM3sttimby0WHS+O7DYL+yT5lwVmGVNQIkfFdhYopByvlwGTOXbKLuLdoLWiS
RLAV1kh4zh2FQ8pPZe84OhdTi8v0TYUn/1CMLKiwy64JzY5h9aZgl/0L4hXcWCZds7Ric48m/cS0
Icz4MpLIm//rPdLCES2MFOhmMnG6zMqdZsSsPdQ6X1Q7VXwgftNZNFUkpXfCtGKVd8LvEYiwBQTr
A9oKlOsX/3LcfS708gqH1H++s1JFP4zGkAKSXW6KBgJCco7QLMSsXO8LyJlNH6bFotTbvkcZEzh8
fyOcXOCzVBzrjgOgdwEGmSyTd9lF+gab7LKKDDhBZMzbF8dYV/T3RlyzQQtif0dL83hJvzdSSPRF
72jlLun2bQqdOpPdMyygIHhd4DihE6Ry87ftGwti+zkQE5FUSB5xeP3fTeY8GN+RqvcQo+9VSloq
7sENhlWOW9pntWCCIO6r2WNiWCwtzSlCeBI+ZdgeFPprtYUQMadZTcupgznM7gaiajGSFnIUE1E7
kftESi0nJKTMNpl2/E/b4Vws7SIHEeq2cbWrgcscoKpTT60bxaMNIDaFcPDNX0wt8OEAWzGoslBG
za1Pf4808rX8foC/hUabr+JFmB4x8AzrFtEMMCpwbNlbjllDH7ER5texg9h4/47kqL3r9cWNcKu7
opiJbQQU6kHc+sOF6BHkWDLXVETiDNmuv2GZkWm8bLlDJ1oO7ZJIZEw+93hCqCLm7z4ZlTDE942Q
GYn9NwSjSTnCvZEuWIg1BiVMr3U8mtcKiefnyoPZmL8Dy/nanBgfm+AizYrt6nlCb+BqIAntw2hH
M6eT2zo920V5wXBdKNgkUfTKQo5/ke/vyRTjtan0V8UfSCU+cMJLj95NfZhpO7pBe/Rwb0BrJHzw
cwLX48ni5gHZeHPTyo2U8SbWBEtJwK+UFHv3npmMdfWutsRwaxP4rD8TTkFU/5D2xEsHtiDqRRgV
jbIdS67ALRs9w/Ol5NfVtNz/sTgaB5XPIAVBDq5ljm7j1AytrGYWfQF2J+i5WKIN/c3LFRPcVOHe
YBCGbsIy/ouE8FiA0LRwZvPrl+hU5BCfqIlAMbWjl5niFKJx+E5HYJjZWo/Y5psb1St+7JpbCrFc
MO9R1YDo7kKPXBx/diuIDxrDQanNpZEpZFH5NUBQxJ/DhZUppmkv/iKRsl/AowgNaZenaJHJNAX4
cK1Zhky85YgTkqXJ9mMNdCEwTeaB4pVM/tB50NQb4hAxMHPWcag3JODbq9xk322DPggTaV2YOPxI
Ngn8a4ZHClWGhyyFsJ+91GDQc98oJG8OEZRHp1xCWjDZNbp56kqi63AWlNH73TAT7jkV3OohnYOW
0DqnjYsBT3x/THw1Wix85k/j/0+GbO4yGzSuAaiK0pGrupDvvKFbglPddR6jHTDZVbkgrD/9qqpq
UxDveRSDH9L96BOwxRoyu9W4wMTDW8wIkOq5Ga0gz6VgpQxKd/JQ7v5PKjNn13Jwth5JBQQ82/pl
itJ99qkvutp7Ajr0PMU3cFEPyIWpjw7UKslrfhgFx4KaGOrak65g3BeTcX6B42wpFiFv6EqcJD5V
dNT3OUOTgU7cpnAU5a7iL20W4gKicdAYkyUqk9yXxm3REbE/T5P8dNHZvv3Ae5v5RAMelqLC11Ih
RBb1Rt8ys8xG7RtWE5kbZaf+BaFBaLqG+GZppI5lTjKmNlzvx9guIILWUVR54Nmt47bAyGvFRdJG
5M13FRoZGuecXw66QRZ7nUUNb7BjRZ6rxhmPX45R7N0oXOJU5iPQ62JVdunitWvSdKeFZuRlguap
fXCvZw/GtX4ico+vo9a1ysQT3vrv9yPTLE/82FB//pZOLD/G/vqqi0DozMAKR0RO5X6yRIXki6qa
I0+geUAUDr64ZyHbLuz2QkfHGYtcyyp+Q8Lr2Ot85Djy0O4Lx0oRLfg9VsYf7cgMQxvJJBVP2PD1
GINdu2draaD7Yfj8cNm7e/pVXZuJx8rvm2xKOxcv4hsSMvwO3hKGZpaCW4baq5GfJ3fEgMNA+qc/
ylZQPxZ9YAIxbEWHLYpO1gX7XhnVKxwj56+sGCK9gIzFUex8vbkLr4Fef7e6uL7BVpuYplSy0TuJ
sXbY7NdS7+RqcDyYZmR9WwuBaU8xH1aOrwCFyWII0aTJ+xWnetzi7zyCCRkZrxU96JMozUKvAiSR
RRz9ZOi/4VHyM9ZwCmZDT4hOsZeY9sM5LNA6alObQ01E8WJME07WCGwFMgj5OnMUowvQnlSmXfXP
xwn272xbS876wStk05Z291XQbOTdGl2yHOed2HyOhZ6rQn6ejFVYOWlBYQTml4wGzSAPAkuuIvyO
KqKUcFm1aqFdizmj1eUzO/vOYaoQJj51EjDpM2P2RlRABEP3o6fAn6qyccOiHvRjt3cjgkXBOS5a
I3dbtQpWrE1jZarvPzO/d6vnQ9CMa/AEUlZ07ykGPSHRbp4ifAF/EgBiWsKyPM8LnKozJzmP10iO
gwfkof48MvyqBYI8MSKWydhCmd68xmbiK5soiWs90Uqe64IrfqrgMof1mK1kscGW9OC+pVvW+dyG
haylWDfOLRLgG0GjzWQJHENuxB0ISbmrJVFRDN7Fwwh1nw9njbs7tmiZ7RKk8qxHnXRCAbO9pMKz
49qAhiQUVKxNCXJ3EfCtxcrYrYT3NSq5pSf8CTAS3fNVDQ9idkRJTdKsAC0GN6T2vCa2sprabTvr
Y/Ykino65wAuuFMU0YDk0dTzr9Ecj2vkCmKdWMXwd5u3TvebMpIxLpblAgTLKOfhpE9FiHo00PRX
d9Q5vnDZ5CU/QgoLrS5rQeFlhTntInPdzN5mjIAYTgvpbNtqv/UTLqPnTKbqxzi+aSgXyRPaxJW9
psDpay+nAQVnRUJbyeI1m26uIx2DxXzNTCEmerc0FRMpux5HFKCW5YnlG3GzWa/1dDMpsaR1NMPx
9P0EWNdyF/HqeoOkFi52QH4WRCma3F0oxs9uJRR45IyGQgVVwLh+HwQ8EVZ2M1NE0fNMAopyeAoB
5ef4mls+rjfRkNUEes8TdyXgjnWnHYPrQMhNFuGTkM0KEMj6l1SWo6HELACJ+8STcYhbondcVxaw
ncMKntUGABRUSwhWUsXvGQpm/lYCTfi6VKoZ153ZxA5448Os1xZky/z8hgKqkeiY8i3lx0UdfnFi
TxmdioQ2RKf5gVooWUrw+4kVdqyg9osX5GNhhIawC0Ie492oOMtc5e3An6q7SANQfDphpUPpixjV
kRc1P0Ga0yQxiqMynZ2+KCoVEA5zqluDutqxv00fCmDA03M0k6itkuSCi4UTOpWPPwuvzMIA5sDz
bZasfISqOpnGop0qxeQ4AJjYRZ75wDAyf4VAFm+drJd8ChYKYkHY5rWnEG2A1fKLtaus6ygZu+nO
y1TSy9XII7jcs7AyIeGwmJ9GRzog1N7CMjz7o2dPViY5H0YITwK0Lu0wGsprGoZIxg0R1MyNC2TE
HHENFB4f3BRfAyVQB/T4boMf8TYW+FHQPy3iz3H8PbNfCTNGeIf/cc/VgGX8uwH33xcIn5BcPK/w
2WcwEBWnNYUeL3a4H5YWn1ZGkMlTjrbZNrMyCEJtqhVSMWTVhK4DU8+062pY5rNjDT3jxkEEMQk6
EURW4KUSfe+DSJn0aht0R9czNDRSlNEi4pQhvvhmBSjPLVJPWGd3gpgRHx56EMGbRxEoREs2Dfc5
VMheoIRim86xVEVwPyJJnB4rQf/Mr7FcBsXkEIwAKDp4VCXdV1+4A3wEf35tT860005z3JhLpkBq
sYLng7e/tNKms8RAtnZRaSqdoZE/TcCsKqG2BEUkFn+bsZft7VzlH1ZMUP89CmxvPRGGXniUzHeh
LXHXAxTm2nmUQg8ESXARHNPAPBGbvkF685D4PHp+0fjvJnPVgsDUqM13/uaJ3IZI8GMdqonP10ff
yjbYOPO5a7ziVqz6n5GJU4f0wrENOx8Q9fU1rdy9WZxhfba6ssHikK3ttulH24Gigyy+/wxbTk3C
bJy/z1F769gP6PWecJCixkgB+8LZCX8+5xTBXGM2na/pHJQdfxt/F1hHKuECaZ6u3Vk4Tyd16VqY
N155dw7PSSZ1QlfrlXYpfaTnw5y4FUrm6gr66MdpqnwnzjQxSNobTU51y/MN6FtU5rZH4jr/2tjJ
f2lyf6rjLmruJkaMXxAsTAf5bFrQ+ceLfks3pRvkxH1naHH0YcXVJwXRtqLiajtzGISVlvNi1Skf
Vu5ZNAzGjDpPANfadp5+KUEE6KV77xVrHx8oQB98BbDAeRpWSyNR28Yt5eOoxfqjkjpUDHVmVoW5
H1jW7mAD4Ni+AN4wXSfql986m3L2Kv1V2nlek0HBwBhRKHb5mJIumP9e2qdEStAEBR+2yEJaYvAU
JEw5cvfgcj+Yyt6clzpwrHnHQ8a4+7lO8ShOr5OjVuhAz9ZGXqGYMV7+P7CECb+ddteduiyaRRLN
nHPGhGLrnxW8yxrINm5HSleyK43LQmW1/TmpIFqexeL8FtTiHeikd8oYcLk8+Dv1t/ndA9xmS2zR
tDotxT1StREOlJ1MRohMXt5vT0WeonnMzMRwuTzcPql+AKX0PeFngoznj9R3YqmggH0JIDMdBCfZ
x+6ZBFCaJF7pxh88UCw/i7mZP5Vb9TPTy0KqwYJnPTUOT8Dn/tTnnGq5Gcmcn2bYtu2rF8j0QZY2
16xokMCiNji94OkaSZDSzLYIzJvXBGs6cVeB0Dqb7Mqo5O8wyj/FPTiJ2glf5LZ5Af3OKJcBdI0h
YQPzcXR1w0mtSDwT98RmXPhDARWPiGUcu3JGj7NLe6keK8DmGadOo4+9x3wP2GTlq+GTTLkvslaY
VKrqSD8fRJC36pEcen2t/jQaJMwyEfuezy+li34VqXa5RPPrimZMNH+RSri54LhXShqdME3TR4tz
XSs5WGiwD1pu+6a98jbUEvSvlwvEhW+b7DBDvb2nzAHMf5beoSzcdTDfXQ44l2Bhuf3B6wXwi9wG
uUQ/pEGRIXRaf0k6X+VbDArUXiYMF5tm5EhZs7KDZ2kXVnIoujOi2/fQj5/w1uLAw6yQCZTKeIit
XEkdd2lSNT+zLmoGdVsptF1/1SjXHSnTTA/cZKnHWnunAF4uV8Dyv/JF3J3+sEc3AnJTa7gHfj4c
3n5ywju9XHAxuRF+mpj0PJQkLTCPxOrIMC6WWGZ6mxZ3zr5i2F5Oj1QaMMHxpereLeA/pKGWEzWd
6xUiOMHytMGJZsx0W0fxPzcgQRP4XRD7xYmoqIoPioy5MnNKWdaO5BNxtXZ2Q+qXBi9su/JycAjY
6SHYtLGuMeoVLFz8DYpTORl9neTH14j8aH82NIAtwB5h8nS366PPMWAU05ul/8YGzooWqKqHl4h+
9rqzoKDaaiAnwEif8EXxTJ6jSrqPVNfG7tHLrXBxk+Exz+4no2wiqNpVAtGT+GruVI7p6yuiP6Jf
5+F//g4Baa4FGQDNZEXC/S7dMhH7K/ARcw7l6IqI5jHjsQTWVi8ZyAR90PRUI2KAIYNS8vjyhxBc
wAFXr+y5n7XizdAR1z3cqzkowYaTmQwXGNcNHnt9ywct1FxwfxDN1DB7GMeQ7g2ON/yB2FnvYSNS
PLw8Nd9eirDNgQ37uHZKjxy0Flli3Tobgw/1yDfb25OODYoyjUVVaY12PLEKcW3UkczGuVrxe+CB
vEW8AkltYlAf0EhcqsrNC3k9nsVksbmf5JayIzuL3m1Zk9nZWuXvD45dI/tn+aatb69qu//dIgJ3
QMQHUsXmzHke6TA1akhheMEQyRHlogAj5ZKEc00gNRZclgwuGUVf1TSEphSgbyleQfUFVu1dK8kZ
yACSfD4/T4Do5Z21/Xl2CFSZWc/MEyIkUhNK13w1KjZaf70om7C1cYYqQYuXV/unVIzXv23+TJR/
X2q3MAUT+SRcl0an5K10TUcwMHvfboVDmQ5JKnQm2pFW2SJM9w6aRXLnMGExujLx/piHescwpTCO
yacdF60KXG97znR23tfx+wq1jzqE6e2vFtP66GFN8U/TEfCNaIFu0TfXsGxfZnoONFdCuHQ0kaE9
JutVvzyVRsjo6IEF09n7bOtolfVu9isf0k86qQU2tZFp7levW9qObVgsHLadY7PGrQKs8I+g+fU/
gixiRKUS2aj/HL1auPz+wU7Wkt6ZoDsaqOFuCNozqDji0CKo2O8k+4ouup5SXnTOGEOF/dUQ6TpJ
2quSIGyvoaCElIRIh7Zs1Gh1n5+T5kotrY+D52r39/zMDcCataEiuOehQTy8YxYPwj3ZadYAttM2
KUhhIMuxPQaHFO7w95nV8TbLfQMvREV9SegzROKZJzcLytRAVKCYIKfO6gQsFkcAzzBFay+WviKZ
u80sRSIeWCjwEzYS7nOnZK0VZq2pFPK/njMNm5WcQBuNHuBIY3Uc1RomXNiA+QLvcDNtiSBL8xA+
vM8oo0n4x4t9GwzXWbZhQY0FpSJQGM2lVC2VrXMf5BsoELwctNFWZMDqoZx3SRe/Ty6PuLxhPv8A
3PIrtVckl8LbgW4tqUxGkK/57mbRcyBMrF+G7H1oQKH2igsgsfCHSIWpoRo52FV+xVkmEx7Oy4QP
vah/9pjd4bV+rOx3IRWtmQJRKeV7jbTgBNjY0TYt8moZzkZ1qWS94TyQAXUuncFsEYo5UWRUioaX
QTxjcMo0926PJW58ku1XMMDzcXosPEBWAZmiH/3F57ZJ+ePI/4fb/Egk1W2qTKLkQxuj8GX1e7tC
Ds86Ha32MCy7F5R0u5X+ci+tsNXCVkb9cM5s3BCIFzuRMRDrd0QZ/mA5AsnGnb8WRlZtfuj6diXn
oMtxNM9bMyiKCbIH7V+4wL8+/YTsay6HD9if78B974K/G016t7QcuD5mvayytEC28F0WRU8NLF5I
+8dA4fht+a1lDR0czXGohdBX/VvgN+OpbHSnZDmYDuyvBEKAw4V/1xDsioTwQCgCxZ2TakTbkfVz
X1T/CMklUXsZPG3gxOym1XOohgFDlNeeOYtgpoEtQu2G8sC//TfCU0gOFeyk6YUX3h7839mSl96k
SfpiIhhGnxr/i6W35Fusfk1/t3+rlLxCOj6mzBJCJEroO3L7ujC2U8aEjeaNW1Rq0IE8kMLNekCk
Oa51Ae7mfK2vnPOi6k6w6pzwlNjy2qfHBcaWw/CSD8D0cQaF668wt3yF+Jo0omSSKTPwXXd7jNxd
b27ZFK8ax/n8xyod8/wjmcqHjJtc6Km+/EB/NSLohBBvjFalDGCS9zVQNt6yL82gPhEeChZRUYz6
ndz2/V9uhcWZaWDG6AE4bf1IH6d8FJ0bTMinlHtet6xkIQVTvGyn/hBHMJEP8B58Auw8iPUUySf+
+NbbVYTHP1YEY4GKfBx2IEDbtb11l54YaP0L+moNQAcjpS7yz3kR05f8PRfeh4nKaIAz8R2YNt06
vrHIx2dht+y8SiCrPnRLtfLmhd+PB5NoLmn+Lc0UvkOTP4kAhbr3xX9KcY+Di2UqhkoMoLtPZSzZ
7jrNfDxb1vwMCLMcb3raxU47aQ6dcupc1ozoyDMeBkAyO658eOozCgIxcNdnKqPqcagFs55XT+ur
N6J8hm7wArW1aiis47bK5l/D2SNLWzPb38kUoNPLsyRm7tFOLm7+IZ9A3uOU9FxVi2FrSvJ7S5t4
Bd9hGYOE/j3CU3WlamN7/i0qOUOQ2UIAiSF8+M2SFOqZS3KDP9YNCtdDU1Oj2PMUm6orNaAlJ/sQ
Vb9a/Md8utCBF/InXRG9HfzceiVXEJavL3G3KulwjLGC53NohP9BaChIysOpzal0qWEyKyqmDag3
6HxmmEElk3OTuOCXMwSBYJnuqONoRINxzDI0q0EqKVBiZzuQx/fxRoe9OpwA9ux5cX4meftuLpVs
RJSwYVmKaZ8lkAwAOeh9O7BjY65+KKpWaDWF53cwiZ/6eJxK6+JnuY7FnANx1R/y84HP1CBs7VhE
Tia/dNy0JWFmFFTxDg+4Hb/AbrgAo9SkcpOHIPzSiQ9wrHYDUO5smd1rmlomlGOo0dUUUP/4SyFl
0ZiIAS3JmuVk+tysjuIrPxyQCylisonGo5coa/bEuNw3hJz2FflBhU0w6Wjaey1OsKV6XcYpnJ9j
WZKffRJNZxPyWltGOoiGt2zyGBw29mEUTYuIEb7plo0f7BNkckGKp0AQg9zfCnT1RbQQbUWZj2cA
SgYEHBhGXcHYy4JGYFk1ZuMnBb69jjrHtXMNq+VRluigbXdUxeX/iwqpEqihK8AukUeiDsxJD6sC
3CF2b5sL7dfV6MmAwrlS5O1wCjKKEeXBQ3p382XuRaHmgz6gYmC2/niiVmP34cmXRI7ldLprQQRK
a2f6Md9+GdtlKLnespZpqK84DLNrqmpShD4PfiI5nZEGrVBRrb+NKCHuCXMVl88E9QgJnTQhOFnB
RrtyPV00NNiQ0g+aw+uX5KlcAATUtecb7WO/lbI0qMxff1dCcJg5XtlqFUkhfwwKN8aIKOVzd8Z1
cL/iVu0atmNd/ymi/6fFO316rxBVr99mVqovoGsUxsBu2TGde2NCPCiIjwVDiOq+w8053ACtKIUM
+d4EKPqFQL0q5kLrM+SZHIojtzMi2nJgYO+KUaFeSoq6l9ATKqdtRRL1hJML5SUuP/YSIgeDVWCt
aQeiqoOWOMnEuswKmr+Cv3vDi0xq/jtvY0uvLBFZMiQKakH5/o60jDxUzSYiEb45AAw7x+i6plh7
1PHlSY9b7LFBTUA5zOqoxiHCk/YqNB1aWpMnW/FmugTAFL5/xh9QTyuWsFlFxndIhYkTEm6fIh59
awQdO1Ma+RwfyVwv7knm0iehMxSlMV8d/O8TxunxsnZPjNEYtNC24+rwOpf5TA1TKPGxBDUIl0ug
MjrPigz6hp0aoSXXBVzFd/jgsssL6XLzr1LeqvlA+90nUHojVCsXV5U3+m45WoFOo1ylLJTH4cox
/8CNS895rO3Lic2B9cUARpwMHRpS35F14rKS0cL4GdhCjPjgYvIpJHQGhHg7/P6LUyiuojNJ2Wdp
b67Y9beg8TmYlKoNGOK97wlb0WTD4OTeCl6Kq5jx7RPSi4N+I9fZhlqTe5O/6FkzcsJ/d7jRCqvV
nSc6UohyyOchDCBlXJtY+deoELKIvOTCmh/rpfn612xrLcNc6YWR//V2ePPfgR1Qt1IIDqvH3cwd
+W1S14gF7TvhG8XqMnQtRuEACZfzX0q/ZPzJ085R/6H4k4005GPRYDUiYHtOpSBxIa0mnPzm2Kgm
V68Dq1SET5l/Qxe7wjOLmEKa6tCA7oLNTW257b0b6E27pwx1LdiihC68cvmwjZMiBHdi7W+OSyCm
MX6nsj/aKbT1NjLSqK3bTjCKw48LLj6wEXq92daLiBmFXQHscgXs7/g0KU8p6X3m5aSd4PayGwTw
ZXbLjaxjtygKdcKVuFCoYfASk8ZUqjyph8u8abvoPhTGq55s2SFxNoXXqPBiX7yn1hej2RgXLWyq
YWGXvrzCH1M1YSEiztgeoNe1sleju5caH+WakYYnnrdTU5CPdZVufwn6/yRIY8a4YIx/0yTXKz8N
PyQ502G6MJHTiSho8jifB5aNBeuD+P1TOlEDLzxMx42Fk+DGtT4GAMKJU3KqSo6NbDQMewJ3aHb2
j/CdXqoXYm4TIUEpu8ySvOuH17ae5T7CDmWSyyXiMHx6gaRP4FyDrtANOHbyZ1jr0MFy4NBqM8xF
VsROEm4TI1pZsweUcv9PocXyO6s0wbwQRxCiqFtBk3XqsESuMUSYS1e3P2Th0f2qw9qxEfqCyuZZ
KeDua6KJSxKOufdgTfyI53Tb+iaibctz3bxJHYl+90fi9txAkZe/pjMkeqvAW6yRBC2CgEVyMHW7
AcUVmg7POQxqAxBdS+PacIRn9ipc9Mrp+GroVCh10iRQKvjytt0c98XbpFRjUACDK4vrdiq+h+jj
woL+Dz5nA27U2lsrTVQJe4iRQ3pTWgSqdJ56M4HNofPkyrB38H4lo72R8n9puh2YEH13OWyNZl2Q
hJgFESueHglN5/FemcXE3u4UWENsFoo6Zi9g/z6czsYXcnM7mLyjIz1rmNMTHW0/vfgE8fhUjQzW
XtdUsLY725cY3p1WQktBBlQks2yc+Y9Kc4sxKb5jqDCakQaK0Ad/oIDISiKtBMoqswy8+7+3h8+R
H4H4y5lba54Zb3bEzEAKghcAdLjhnPIr8RTJ834b0elG9+/KoGgRDmwx+f5l8zRAgNSdQJCKTQY2
zCj6Low7+zSrETEbvb2ZJIC4bFCxa8qdJjPsacGBKVIoSfnPTz0Aed74pJF2NsbrBYcln5lkvWC5
m61Sm2E9TbGw8DeKo8TALbcz9ErjL/9cxelu4t65xFayzxJHToudFT39OToTQ8ggwLxHEx4P3+4x
eGmofXrzFHFzbEQqJRZu2EIKs4gnKTNaDNd9ke+d2fM87aInbddRwtsFYQMzbQNRcoZlpf3/OKTY
N1UkBlpCvFSkasfKWo3nDHPat8mJw6ywsKH6ZStxTM9igPTrfnk4sZAESkU6fzCHnkKM3bO9MoPe
Ts+AxC9TmLYz5UeNaaqmXGH7qRqP4yRxNgdS2DmKEt7KcDyh7t0EbNX9KjiQ9jCBkMiNtOzt1gzL
dAaVcJ1+bQCbdGhRzn8eRKYU/1om/cnAv/CkvyRcQfJ+bnhMWvmuveC/vLZtCjD7VwiHLzR0tnrc
fO9Es1nkNtlWqTPaQzEDgzN6lGbnj79qdrKZdg4gk4c23/sQmpsm8uPlfOOZ52O4i0A3QNFk4ues
8e7/0Z3VRB5dzIBVo5kSnh3VvOIkVyN+lYYCTJ+RiI7ye7F2W09yzkO0UhRQDixxmdUBL8J1jbtg
WlXEviBcu+0ewObPqJ79TPZg1d40LaixZT7G+oS1ePQGTeWYShS6SX43oOPnZenl7L4L9123GW9O
m5brSP5ELQjRoicHYmmQo7AhddFW1BkNjCjLM3PiSE1ux6sfkmMRlqpeZOqyVuaIRmqRW6639pr8
sPkJLWDxnDTjsCxRbOEtvv7pwDXZZZysNo3+tjwYQX2OEXgTwTacfmg7Us0SL69fGIMdtyGHo4KF
7YrHk2lxaHzkAi+iVxK7JREDudhdzcuD2gpNY9N93jy5ny9PNRkz/SiheHi4l3mlsx00LIZhJ6fA
nYldI4/4mWGt+dh2dEN6wmHTFWPM6vvDNc/S6DK6o6dewTOR9KzAy27DxDaG0XON6On5zfv1LplL
lSne5l9LZiH+gAnfDeF/+NtMbFF5h/Ht7TM5UDhKL+gMBAsWCLxnqxYKaVqiSaXau88kkxRSVSlt
OZAUuDNe02KrP/O8V04YsNnEkHdfoLxtjsuy7/bvI5l8oxnA+3tNQvzsw/gXxiEPDQSntkO8kjWm
5jJ70pPSYv9VtEzyFvHiXLUO/cai5Ib56uP555hiIFTBo+JYleEmNyKH3lFtqCrn5I2CA36bGdk/
LoJBx9hx/PScybvv2+p2b0aRJflGE2T5v5TLMDZykCvyakDjcGK4R77WkFoRO04bJQOlR9n6ub/w
9j5m81Oul7VG3a9Xkryv0r6Q/W1ZNSauusFmcCcJxpTQfUfaadyVgnXHxVPJ1wk7TWAf2xKvecj8
/TT3oSPmcLixaiSpJU0phaMZxT1q060rgsr/s7ncG9LkcAeAOuIhswXOlBhDCyxRCIwqbXxaj8xC
HxTubp6iH6ogBsXPGktvFUIw3FFrghnlzL614s6pjk/rWiD/NLve9wQjoZ83n5gl4x40nU9tvxDX
B2f4h1tlGJ8jYfSzcrE0oZu5y8MYk+OuyW1rifiyVXHLe2X365piFbBA4K+OsyfmCb1E2bYqhulC
z1qEtP+q4R33XAinlSKWhjNWj5ymVtJWILWSvlMVOTmSpX5tuAG72A4bfA4QuzCWM+bqZrxhu242
owJRpo6pIzNFRxHzJ7hewY7Uf7tKVsabHz5lfWFiIr7yvFMp7nmA/NI23FC/eO7Vn5E5ZA9Ghn+q
bve/fC3t/p3PNygo/6srpTmehOKXgM96+a4gO9FCon1UxMeTDkduWqMUlX2P8GuDYmD/jP7DaWdi
w8EE6w9PawSxGl/jg5hApA18pyqPRy6f/ToqJB4Og/tFe0jXM8Kyndua+Za7SUcbfkJuGRSYuh8v
k+eFy5ZX2PWd2BEgGl8SRiq592qwrtJlbtYodbY2m9sTkdgHlJvAMAy3ZFQHqlTXGDvm8Q9BCA2p
ZXalPFhdsIDm01ViUyBC999ToCGiykDTaK1xZsO2AbYIQPjnbRy4oSjnVetC53cSsohU1bs6a7zk
9QKVSI3rkr2TTVWLiH6AD9omY9aRu8gLTntJEbFXAAEBT1gAKLcQ6psyNTLeXjF/Tzm7sz6bltPN
uLxj6Yq5F4pNFEKYgnbcrEsGDsf/InSb96WBBGeyXVYHetokZk08J1APZ9RTY8lZe3yuNPAX3rPY
qoi6YbrDDbjnQdjmF8MXV6b+RL1A7QOb5wN4dQUO+GFwJZmJ44Ftugex4nQoFg5y/vSganMabi0/
FYVCJywgMNe1ieCJeCmtvBf3Z/Gh/uQka1XJSwysxV+3yVmvJBr0tXsmCYceFPVGdyUtCk7Xzb8T
a/zY7vqZOM1oEUUW0ZiczDNHSuU+9Oq5w/P7ZvyYs53n/V+32kODri9uo7i/MmYlVVCaZppDpbGs
acK4T8UuhOHBS8PYly1Np7DHvg6fmlqAfV2xsfFWWkYqpIZQynJgVzKVtJMBGe1/0oPPrVF9IdYs
KRhFl4+SQxynWLZXL+MhW9iX/lGm382oNS6eE1CV4d/hPsILUy8/3M67+NIhJR0j4UpW9IHOSfaw
BMBmiBEvRN5/6gd4Ti2h++eB9R3uFrEOdKllJiJsFq2TQPv+MI2fWnf5fwer8CUYT4DDnsx/HdPN
rmJsK1OVFgeJHiL4qSGLRor4cAt2VseLTvv5WBzdlYYAnCL0nNyHEuFr49Wt+UlU/c3PI8LodoFZ
5R+4Jz+L/WZtrOM/J8RAElEHWGDvxMMF2B1dcyy0CPuf7TuAAT/hmZdPQN+ph4fcAnSkMzJ7EF+8
zoFPJ4uS/U0aZBgAN8nvLgtlwop96ZUtOQ8dmdq13zXr+VjnZsEQGdxT1K2w7Di/MYH/uB/d6btn
gr6HgU8ahhmg+W10fXtotXnSW26F6HNgLyus8kOKzUnmAF6q7ZV+u5QratMCYUIlXDo1VKVL1EGC
kixUunjfJSheXUqNQJtKPebV9mvc4W2NlcxlVfjezmpC0/R6ZG3YRipPlC6XaWvl8nAIii6d4O1C
+mS1AuvcKg4CtzTvuwk1zEhvZ5hiZ9OsGenW9uXXSA3uOKrMTRAxcbUPvzOc4C9k25QGqcODfyfc
33Ey53F50iBhnxvanzPBJray0xKBM/eMgO+kGX7RC5pTzUI9g24fCGayr2JdXwJ1XViePR/bLBeu
6dv5b4bvSmfOlb2Hdn0BVUBT9eft6K04IAT7f+WkFzRM9Mp4Ltcv3li62UbKz5eXhrQpn6quHEhf
BWSG8BEEGAxB1RKfD8u7rlwgN9TcsEhH0MQxruApF/KN6lwQzbsuBbOPg7L2ykb7QIny0ZpGrZQj
d4B+wtZyppq4fRNMWaZHD9u0dXANTrKh3TFbavEqYeuu97CbM6lzYlGqD1s6F/F/R0Rkt0ogaRIT
2XL6syWla0sNp7t/p0NQU55qdHTGx2W55T2/rcdA1divfFDnnNBceXNj02OxloaoSDVghYGnXY8g
njI8oOa+9KWBSZdGwiAwSD0OoFt8kB5C3q4FHmRx+SXAYNguSH7igInJFjBUduN5VZGnf0jj3Xxg
d4TybsQHfGuf9FeqhbB8aS27PpJz7g3S7xa7e2jH7/I6K2ZRA0ln3D/aDfXqtUbX9avYK2vqwW5K
9u+UGMXSEwmQRtnyZDDqwX4qr9KaWCFDvuVicO0mLQHMPtef0WMCmdbT2boIYIv4ffxPVp4VroRT
nU4BeVDMu64+wBBl5L9MgkqVDLXHkq9JG+avst/dttch6FKaQbxnVhFysJBv87ojBJa088LXd5Tj
+mIlgTp6yj08pah9GJNw+awUKoz3tT8lK6YF3M7WXv7rKopqK+9Pd4PT0cb5GnqQCO6zO0D6EFn9
Rn+95Aspz/dpA0+h0wMZP1HnuOiQqdhEpaUSRwuYw7KkgTtXQvllweAjq0mks5Jv+xwz2eHPcy3j
IeyCMHatk6wra/hgC0TR6OyFaR0Yo2i+9thIZ/nKG1WVRwKvRgQrnZN4UOmSUYdWZnsPlgiX/03z
vNn6RK6hdN3iydYxGbONJJX5DTkdoE7Dyu1WsU/J67f3Ohj3XCpgHr16nhq11cw/MtgqeYWmxpKR
GEBvdnX9P4zCvC+W3Z/9MN7SLiZZ6UyR2RTqISu6rsdAEucWxpPiGexVT9j4A7ai4cODulUGyV+Y
nlEnRIziLU7f/GlDfu5mdiiXb1NvJ+zG9TcPtnjlj05diEQXV/VXrLL6oikcyVZM3Yh9OEuOs3B6
zGiwLrTp+JA6GGBFnjXPyPQ79jnnK6nfiMSbQb1YPXbm3JsoRTwBZ9PG/4cM75ngBM0/wNuVPbvR
YnV7en1hVSBc/jtOhQom3P45Lf2ej/LdTxtltpPWsD7X0DyZzneIq0IByZYf/FqvFybuMPOOOU8P
uUrfy+26cg4c8nHDHxgYIY0N6CXS76m09zQaSBYpvoTfDYRXckgM2zInBD0WKIgkRhtRL5W0wUZH
CKkIUI4z1ldhPDqvslkOgdAI8qtr+vgT5yn7Qc09/FrCgxrGgQsrpbjaJbv1ilBtegoOlezA+dar
iTqa6sOOTCg5bsWBTSEpY5JPiiYRx1GaRpBgZn85SdWMMoui2mdde7PQmMLUL4UBMwxuHkS4bPJW
um9NIBobIjFezD7UTJ3+ZkmaC44PbrVaHVgnk9O8ojSes3XBWIPpAbjsnpD8iss1Zvl5H38WKI+f
mQX1r+v2nu9s/0poiOtuT0QcbfKX+g/iO6WgXNfZyTHgShlLySdl3+tOssz7ckxdFrBZLt3RlHM7
d26CAYLHi5vXYErFIN1lZFLOWnb45pYEkHfPVnZBT2xo5kRSJ05IAD0L7o3so8WqDMyA1I0eSPSm
h6O6UUdlkZbaJ+VdVsPixDgGmZ5H/CmZMKOzybn3yBycXL1kGYCztCKKGg1nzuXcFKgMHI5TNPkB
njpomFfN6fgHG7meyanQF89rkZApdSkgm1wNhTzyJhvOjTZ1/e0rk3gJU3SSHzHiO0pOH/ejFbdG
RUTGXa1hS+SdPNoj6iKfgoRM/cKqDVbaD47ca26sJFGAwQNE2lbrbfL3ICLqDDFWv5hBUVKVn9dM
PufDUciRyjVRhIk61XXeWo3DAoTx3rPjFgyXkrZ795ucvVhJc75gy46voFo1N6g2H1E2PxEUQybf
EuFN2ocBNzZsivyie+YeU7TYV2P1LVX5GdNj7+LINB/Kag4lgs1Eu6Muh1QD/MKMKsPQ0/D8hB9d
fIWJYXY32I7aCkMGGfQEIL/wE4EPODuaXjXIOeOg/sABLHPq46RwWz8B1vCexf6EamSCN8e9U6dt
+ey3aJpfb6bXlI038wsiCnrQs4Ot6h7rPUSMhIbljcbYZy9croOcdoJ+HBCb4Trm9iGbVkdbpzel
taBpHMUcTz/VxvBrdl24VE17gVJofFp7DzXwOlZGlW+dKKbK8JZuxlimymO1SO41IOshCYt9HBsx
x+fWJ7SDuoXNpEgbYHqTAlyCMfNG4CT5nsX1czYVpjMYea+hYtiWYc9PUqdPD93dlqpx+cN99VpR
DmV4syrW+X6lAH/AfACkGC6XAtz6B7vEBD++Ra0XsdsE17FDIQ1yZxTD2UF4sTAyM0odjIDRzbvz
41bJJkFYniM8W6OcHjqvdEw+emZssKIGKVIupWir8P1Tn2ogeNCnzKNjnycaIGFz57IOUUK2Xrdv
cS5g0ZrgSvxERZB0iT2GpjaRI5ug9yDJ4Kv+cjn01PEiHfiEUm0KgrGPGFkIY9L9un/NWSeBZ6FI
MAlG1LY86h1wYd/u5M/WSbbQVVke1oRQqktLsL2/uEJ8JVTvuwlq+62m/v1NVMrH9+CvXTzE4+uR
gC8RnIc9oiBe6Lb5grapxKus/BHnCtYDYJAVva3+j7W9c3hpwtmRa7pJ0ItIowW6CFRu3Iy+M6J6
7x3KMnN7V1IE1vgNJQOrB6IqhF72qAbbDvISXC9JHv7UxEd0mYLaXy/veM4lZD0jQM4Y8SeXDatj
9luaao4IHHHkggU5BWYWjj1bsGglQL7DrdkVHrF0Gk2FrYllB40REUyX1rEOsAxklkmlaQcY1sNQ
3akPn/eYynpXAUTOf77cdVxxGigGEL/Z05JI2Ggu9avLbntM3cYCx+NXh0Z8wBrEiJVb+lrj5HAG
lwBBvlMyHioyF+yVdyyZe2vobzA48Fx0CB3Ks60efoLp0dyr/nUTAjxApgZbpec7o3xW1+mgtgn9
2Xaf6Qq0QhCWWC6k2mlr7aLXzdHuqYfS16VyTLmLmKVDZQrHE9CSssVebWW68Ugbtk9g46jaX+J3
HIUC9pkk0BT8JMSx8S3cPg8Lx+9Zl85kEogK2kdTh3aUEhOYdeB3yH94aBGix8Qh7xvx29irYeTh
NyEeE4Rh6AySdPktK+lJOeW2E5qPv0BvOgAJOtIKjUlb8N88l13WjAaBHStEiWNTnETH/qVUxiov
QNGO7jjvLTm9o99hByRy5mrgIQW2INiId93CSgL0VWwUB9DlwE51tP7RFANQOB1GnI3BTU3W/bO2
XVX8ZYaZRdPZZF2lyiUL0jSMDzUrUYlz4ofKLeUGVjwp2rQjbI7mrpUhtVomSYI5gnJU48HKUBAw
6gA/IGK8gaaC/M+c8yaZHMGk2vDCtAbEc9NSoKmZ/PT79h+3a2ENAX+PhOuom6UJeRbFxtDN4SVN
0094gNsxn+kUioLwJegNHGKjflVcahwcgGOtg0xfZuiw3YdskRlw+WsP/N85gecu5h4rdlRX0dn0
JSLL1cnL4T38MwtmHuXJjVTVgUa7uU2Ll5PDsNpy+fUtX81ZAO7E6RCQKmITkyXiGLSnnFOtFqlt
aD3Jm1cba5NYJmgHdqUF4uaNjEO4iP/gGlc/r1UEea3alURnPv5PbYp5gLNs28p/IIa9+xMQ1UGw
wLoheeJJ4GSbYPNtcSy0XIBsZvJuvcURO3i3NH2n1Imll6P4/9Vc3ZNKBoVhZe5IDP9qBwQyGiaM
22iEQfSaA1ObCGN2ayGnq/4Uemz71A1tGXuKXqR4zF3+dNSDkuOo7tDWoLBrXLM006+YgQgaDStT
IWBj2hSmH5pTeHvXERaOp/31le4k68uAKsuycmfCGkLHoA+/G9Cn2DtlRNeqMoFnWk+rM8XSIMrp
dMfOLuwn3wxIHBRNC7qRVoi449EOrkEu/A9b1femXNkqtEPxXV1Zorx9xoQbnaR6Wn5QWV8Fh8nc
4r9XXnXDlmysRystQ7hHhlhWCuie9xea7RY/eGdcLtaIRBy1mupQFXYebRJ2rdPjBiScq5QgxeHA
D5gap6wDkiG0LD9HWkHVSzzozPLjzpwBnKMP3GhDPMrbfDxAgoBJ8cTz/VwnqFHCRMOvTnJ/gC1w
iNMprv7OnSe/4q6u1IVM/mihT6Pgn4DlFuOvffMSDdhkH5zxWhiFHFiKlhRVIy87SYJyako9WsWm
D6tKwH+r/hPqBw7X4b6PnKBrBA9WsGGaMO236MO7NmHsHjye8N3RtxeD4hzb55zHe4QijXjhAXL3
B/34cT/LjuNGWjKk1GQorRbAuNUtd+DGBIL+j3TwbjA+lmubEZYp9Nu2icJm3LCgpcDIk+ESFrfF
HupBCkw8NVUPtfD7JG4AhpwGx11Y953Cw2der7+pJPURwu2pby1EZOeOi395Li7nfeDDFxJ60OIT
axFID+YSG8S4dfM7eKWBhjTTHsCdVyF5s1WtHjWs9S5UtTTn1TPFpV6tmDEef5Z8qaFvCg7IlX58
++5OBGJyy8PT0CmEiVy434bTm78xetn0nAuDsUCco4U+huaC4ETeAOByKnT4hwuxtSpuzoY8rfFM
yPYge47CbittAFfsyUuxoCJnIw6ryA3E+aHDaIOwiPi/ygzHULQ2/DyZn0Y6xxOmVFPpdszM0qnZ
FheWP178HDvJRtqqKPYrmW1007R7rK3+m1u8K4YK2joKW/R8y6l/HrcdRc3YyzJ6kmcbNcTeyS7g
2IoTOPM7FkcvSAaX4ZtHyrSF9lxVJTnPOECHIZ05hPoXRcOuhZHZ2EChe0hEHWZUkCppV0stc9gT
mloaydjwwMzxArRhHd+D1mQWBRRBFltg7QM6OhizldTsS8xMHrNeFA5//z7gNVWfiwRNhoQUlO6N
dycWNQwNNET3G9uQVx4ziIfbnPlrC1HSaxlaiLYNmnIMFb5KSQUk8gqqMuf/bPIVFcx5DpDPMxRf
IZQGB4CkzHolil//pueDEsSL+iknoxLUtaTiWExfrnUJom367J99R+gZyI6dx+0XErs8lSG8r7wC
XH4P5Ffr7A0alSEgEyC74QNCKgJw4S1mF3vdg5Vl1VH2eRiFyhlxr1dF1RJ9zNyGofgUglJdyVrY
BiA9Eie7EYPXMRvgLm9D3KvNPa5dvpsCDIe83wjPO6EiLTifW/+nosoAjR1gaMaY47RIgcAxd0Lf
Vlyi6WwL4MusB80UuRAoqIifbY8TdES6qcNIFu1nV5eJJcOZuB20nbsGb0FuPWa0hJWbXcgX6IYp
7w4LakVkIAbS+FoddDd7SWlPvgDyiQb53RNhQguXLQ3cjKQa6fJqzlPqMLzd+V7caENcCn9LVwuL
sww74+Tu378ejgHfEIJbBysqAm5fIFL4/yeKVgjEiybu0xuQMqkT5y7Y6gGqvUmj+rD5EMLzfpqj
TDPiu9XD6yguhlFPMqgpWBSxqvbdSNRRrdFWYwsXhqgeRuE80qTu192BtxoENn9/3Sv6LPTF/1ox
sFwZLRD7KEVIwkGe2xaurXCJXWadCd+ehnc9uNC6zilDZotxyOU4ng23/5MyAJtSI9ZtlnCHu3RU
FA4PNwtbK+2OTGSz/3HbFv51WT8gcO3ouRsfwVQYghzH20pvJ4zzfM6aQ11Afcm9JIF9k3dIASxU
mZ+eJ21FvUwmhhaha35hkokzz39uTvKwo0PLmi2aZQ9LZ6ByOamf35cT5OO/e3q4UJU0NTL7w4S7
Zt0A461pwgXR2GuNdgPzyzoCu1aWh5YHUlgtjqggl5m6gaXgI4liO9q3euRyq1ZVjV1acwF6jt/c
V57o8MXF2Fo/++G9UC3QMaajbIZRZi3V6B2Vf4xpQ/wZJPPpcbEg8GPLUVzXIEeNPLlh9s96yohG
XurmNPLV12qcH4invaEZC9VMztgW/rvAr7K70R/D0AB9fz2Nxvtfrx6+SwSb311ZoJcDh9z1mVND
8r5btlCLhl67Bfq3wnERL1a5z92d5EfeDNEM8ThlJkycfYy/+fIROVg8LoZwfs5IE5EhaohNlPzy
k+Rlf8s3BKE7COPjs5R4vg7XqaIShAmmfBO6mnqv7nrRl2kdRB01fda0GfTNU9By0vmuMpbvBPdE
kHMwiybVIANOXCl5D43u8+xN0wocU353CfImImqjWcWjMrZQSgQrWQyKI8X3X2dVRjDQ+lfgDy6X
jXrPSLfu1bGbiUr+l6iU22zcr9iH3qOquGRuwEseVokz+jMzu48dmLqbRBVCIPghl+T0x/PaaUOR
ojWyAckT/UAJJodcTyRfBok5CO0XGbxtgGkPtD+bsu086N/pEYeTldPnccxke4y2NK9VIo6ZtRTR
P+OX7lMDw+PituLotufJkf9A8jWMWM9OsjHW6H9VYrEw5b60Uk1uHUmqe5XGUDjQMU1Rk5z77bIX
u5uW3ilIqdWN5CGEHUGTUfs/KnoS5V1AbDMTpetmkSM24ntSTgv9OXCirm1U7fPcW4pZhzqo9L+n
COSFPM9scFa5OAs5c4zAQycaPguikfi+PJJNqT06IBF8QSsTOlcrvcUt/bCNCMpgKJFZnfaZ/aOs
uHlqoy4g73oJ3jMgeFPsqNK+VWREYTP/sUwwPf0vrVyddDT5Edam1dZFck5xNLdjfvy3J1oHgEyx
qjKWOVrl6+ZmdXOKo2KhJnwMp2y8IRKCWvqCFQA/j3P+u9Rd6UQpWvK6j/+lD4q9frfLVa/EKvOF
upPazSwoF9mesry2Q6AIWhRcKYPe3lhwAvojzwOgBR6juQr4sEUcL9gxh8RGnhyD8bcD0ugL4Ya4
z27FLwHFuLv3k2j6IPBs8UU+6H+ncngrqkzNk6h2AsGLzPZNNp8/VNquNgqp7ilbNscJm1/McmpW
8fXoTusSH7+FdNuvHdFUn3qOxtOrfrVoSXIrmuWOeSK5F4tAd5ljUFUC6A1fig56CgaHDEOrSNsI
L1nFrilQyWDn0LUDbYAmTSS+C5048moSfm3iIZMnjJ7sPaXP9xlN82Azz4kvkmh3ulTC7G8sldWr
zqKIhgBk7E0+sTcRmY2b/XdaTb9nU19D+6z4CQZK2ciBCtX/uuUX9HZKIIPs7vR5Yo/TuY16WxoK
Fwff816KEh5pP+cCrPiOr9C1GzNIaoFv5ARDREyQfPr+s02o/cq0G8C480oZ1JZlmk9NylesyDvn
GpsxzzrUZjnsAiufFnUyoZ0RRO/GKnstXawUChqSzx3aj7IXSzn1LGVqo+DTWGomjvMZwEFeuhdD
TdRmVhv9egHe0SyZFG+FYzDVtg9mi/AIFcwUKSgG0yipsw5Y0O8y1C9xCCXsKD0kxyB7doYXb5J2
jyw0EKLshbXqZ1Jnxx4qcvhj3svGfOOXOyvGKThCM/AcQ87x1mxHt4HAUsl5kchlv8XrMw0huoS5
ispBU9l0c1dh2nbZHII30Py6kqMn5ZNUyoNlCNFbMjtOac5VlV2FJmM2IPuqE9Pn+4brUOvLI6q+
tu8mpWxds0sodEjUzOJQILkyEO3eQ4FYl4d79JTYbfuxxnN2JXdMiWknTwQwmZ9u88kcQ0IeyPzk
4bZtP1gHon0rsTW67Jtk6huzdLAoeWEMUBWIvzFXMoeZpIytCSNpEQQAGuK9r9yNLrhk6XLWPgbU
DAYV9Iq4dsl1K1cR48dtd7d2DHlCk5cUJc354mR5XfEtzTQNEYDlMXsmEGO1WxV9norTWRIjIIsw
oOt1L1Yi3ruceqvyMxNPK8Znf+4ierEL/xu8OvdC0O2YQmslsMCddVVsIs5GHoHAeAe5qLyDaN7O
fUtNkVhY6Hjt2eswOYhWJcAyoyXqzOhN4i5CWbg7K6tmy/bhFP4yErjhrvQXV2z7zYwkqdPq8JtO
oHcvdmFxFDnl4ysLwbDyxsZ+7ciEtdNUczabp4jacPWMewfOZOs/XnzRbU+I8loiVicf7Qoy8B99
2OE6ipNKGDIvSNf+J3Hlnz4W4RgN9/N724sCy3vBtNFvZv6vrK66TNyezwmiTCv6Bm5DUUcGgjmQ
WFitYaVhSxREO+FgRx+aHkvXi1/Cj4iVODIEzDN90+1QmHkF4LzgC7TMu3bG4yYZ4ZiosJv2rzoT
hPN5+kdKkWj8pCibjUaDV7W5fO/WtuZcAna6SYNmH/y8BDc26wVLZaSWeTIPyCskMuAid5E2xMzR
E/4wDcp5i2+2GcRnEjFMeU67mg6zXYglhIa4YddDjCCrcA3w/FAaVaUK5MCZjaHMe+73C0LEj9hK
Z5iEwOCyeAQb9czbD11y7PT2em/z+xJ/SyopeIawNiqCKMChmoZOA4+StWimmxLlneOVveHOuKXd
LZheKAVmDBrQljThfi5lu6Mki1oJVWGnKyGfF7TiUGxprVjBPf1zsSHezw5Eqar5RuykOVqy5N+K
cyGSXmYU0p5gR55zz5D3Roc59CZEM1f/9vte829Aokjb7WbxEa68y9qH1UvQirWXvSTH3GftOUcF
LG87QR2SKnYHpox4wxLwToQBM3D56AP5Rgk0IoMGo3Ij5qMDN1j6BhJbsXgSXfnDk45pJNKyJghK
r81jydeTN9tPGw7foJc6Cr40oH96parkFLlUzYGnGPTVVtzN3OPWTuEDOaZE+WRa4g5LG/GGLESe
MfkRhLZB6mQeDGWCy7VfUA9ONN4b7QtRjOBcWPfJPhqeVGgNLzTdeZ+CVyEh8ESkEnrIgWSwt1uF
CMfdH/s4S2H2PsfWuo0yaNY/2KIg6q6dOZC1oB1xMiWFhNoGtcl3JskAChnwIY/gIqg9zK6+rX2X
LSaXeZgSmD/aZgMS1S4s+/MPpRwkIAxriK8VXHMDuQjEqZ8cWddAJttaMJaEVvbk2lDRGOF80toB
tYfYCS/dujvwsKOiwZCcQV3ZQUurHSrE8Y6In6+wEV4bwlz6vd3yzmqsgNEh+8UL1Xa5j90bg4gn
sx17E0Nn1MbgFI0OiCuQi1FS5lZv+nf98VUqLF/fAy9vkaBhwnUFOHMMwfoIxC6KPnf5YPtv62pG
K5sQ76+n42T6ntUQr20B+oyZtQm/CR5SEgCHNYnVetzcaX/fzFPt+9Do24vvwqjz0Mbh9naSk83B
r5wt0d7P018W0Jx97HOQBHPCoDswZbOmdJzJL1lWdwT63WZqRXvyTRjPxISbw7ZqrNqfdPwakHI2
DPXXFlBQ3cS+Y+0BwaLSAcdJr0vWOz+K+It2RU0Y+AjmQsd4oro2b6Aw4NZYx6hJobXRnDc1Y8kg
/zG1HASYAUtDVIUt8Booh66+GCFy9RjBAHoI8wVql9UhDQGk5PIjPycO5ucDQSMLnlwxXrcknF/y
cnjb10CevTydPNpGAjZat3riLcasuhZqTSBa+ro6x7JdfvcqOZlKyt/76oYEKZrF2bBQApmAvg2e
YhTMjx3/FBnuuFXmWuAHQvTNu7CRftXYcmGoAXr4k7Nt3s85RxbDA/N1lPsSrh/rHFuI5DjySd4t
LIY3uEbPdAknsBZX27maaZRibMruX6O7kOA+I8YEsEyCQamPxkSneHw3TCufWfXb9k5KWgBOvsH2
Z8a8ovxqndniAzjGig6T9U3yMSQyKvYXdCq5gmnKr3AUnppXAghmu6BoF7GEgFsFi3d691TzWyUK
VAk1dI5ez9k18q1TGxwt4J8l2xPp8S64F5uuPRwY9Msa6f0tY+zxGpf51DDzmBsleJrfYNd/ZGyE
cOXgLJLtl7jD1WpRDMBz3HSWoKEmrh0Lzt0u9AVz7P8JQtBJMRRQr98C6m1LC1R7NzQPjQsWBwJF
GD0LKKaboCfKwo5twji9Np0bPG7FliQ4aIp/ytpOZpfGBnWta1C8Hpc5NNgQ3qEUGWRQ47kmhufl
cZMnrRZMN611mUhwqjPxoTnFw7RqT+y+uYDPpiSuAVx06pP8q5XLw5gA/jXWfgTEbYmBOyILstXN
q1ol4mQPmAWwd6IMHwkPXo5hVo/u/XybtVxf1ENi69qaEvTqY4gdmO7TS3ZmRvJfR0YhZY+cafBw
PTXIYppsOuzwknBXLPJijav8HSp59iZ6rtm3+VTAj4mwz3zFJNnBp7l2RLgoxMdqx3OUW///AXrb
y/ve5ZSnmqVjIm00KFA9+ajWWqlg/hbInw+Sl5n2D3FmmOMxKlhQhpoNzr2NJKhJ081ggJZqMKYU
8/LXiNtpp2XXBeJch6R/xjzb47dun17r5USI1MLq9o1ZxNIFUNJqyN32QcDvF7SOBC14aqdTIl7U
gF/2Y1cXsmA3lf0btRgQfLqyAvA2digfzaWKGTW9Im4NwbViIrX0kNUEtELuvPHXypkCL1H6QpFN
KYqe2HMGesW4L7MqDtH43CJ/bSZVJsdR6H8Lc9EsQyX0ZA8oJxEnpz4hIPvCIRdfNf2Gxq/NBlxM
FuH9z0rrGeBNBU5byRMo7r63ZQ1jG2myIYI9BlVtd7TiZQ+uDbPxpUdmLEyFhjF4vaKPC6XAD9fR
7EHps6rxVSM8iik85BI3kNr8BEGdDRiR/T4CFP+s6sez9qwOHEGGNELUHAxku7zU45/iMDtZ/6rO
o28UkosfhUUh9LkBgESba87atAI0k+lKVYYY8mF+fm5ZxZFCYbcE2tVj1SYLYoUWiZegLQB129dP
eaj1m/wVGiIhtVSCHC3nIPVO+f9zwYon6yhvKmvLj9/0TMpACDfqskCyeB7JcBG70tNJF8aMKHYm
CNm69JyRZsgNqoic1pCPBa9wFUf0tt7Au7yUm3dMbwSTskockJgVj6nkDras7k7BAd10TH0P4cl2
R/iSUCLIiDFUrQKiOeVGwuI4FZVw5IHxbZg2BQTkNYsj+pjsEdbqu5qyyBEj7eqaJjIVZDBh0WxS
CyEaJ0vMALP1D0BIQ/BW/E8xAUnw2l2zn4lcb7B1kqtp+GekfbPLLxeRItmWmLDlZ+v7dP6KsmW2
R8mItkocrOHn0BeBJVBsKl9FVRBjJg3WdfMjZMKbfqqvl+a7yPlK8nIMmWD2DKPrMQzbEoXurvHe
BjnIEpegy3cXQ3+uDhbZB9cukvev7u7mX2DT2r32oH4qObEPJDRHrjOcveYaPlTjid85ogr/auRE
HpPQdMlnHLPKVPxbm9FYPwxQBa1DjizcD8iknPeHzi2Cz39pO30jmOMU1++iO1Wmw04+Pdbsn+lN
kw6hjRKbi5CrMrEPYJoNbRONH8eX52E0VHvgPCOKERBfMwxf9w6bFHzV1G46NANhX4ajjXvxLMA8
q950oUwXJZg1fJYhEOVGeKoGLNi5jt9T2u8GVxCnds4ajQeb2VSIsExRwmuT88Zy/XZW+reChVcO
X3Ybi+RqZDhVu+WMssBozTXHv8nDu0+RMEFxZwAolnRi8QGN4zMBgLarEHBYU9iGi6CFF/iDc1kQ
KSZcpCq1BILoP+7muK5uoEYB2VWBW4eyGTDmR2tKdiT4s4MAz0wze2j+tbeAa9qjriIaJUP8/vkq
2ZN81a6tkvNvxklWhQMw7+23+bSWCVTKggiUT6VhqAlVRQMXxsowa8S6p4Mvhqb/BpoHX3QzaCYu
ZGfFiKskC/hH9dOpx+ryLVazULCgpzqaLWUATwI9eW6ipKXA1obWto7HMbl9JnEVSoJABWQp7wD2
5OOGZs67EkI3SC3ez7sTbtHFvZSL8pfH9skkx3FF7T/MpEF6ZuhhB5ItetdgOqDgSh29dSFXWc1y
4b5yawY0aAgquic1ky8RFnOLESO5AbiwbNwllsMrVk+fx7yJtY4k0rXPC1db3i3WUaCTVwqVm2Nn
UHSofRzppmITxFW2Jii56ir4e6QolLPS6fXAT5hhTudepC3aXrU3Mb+J+KTmKiYlnEt/p31LfuN8
I5IEmjYpwj6COozbsmbrDdbKq7UCGa2netWdI+04XfTar6qdUjnIw8Czt1Zvq7uSHLWwLyMdQ0bM
7eF2W1kpFrxncyZsA34b+vpyJ1DsMBx8Z1cc6F0J852/MwSfcDMywUbLHv/zUAVZXxI33XJ0Sa8G
+jobm/I7wk5B8kmMQMCOX6DCAY5yMWXwRKLpJ2nyaIs//6pJ99T752pjzn2ifdrQpc+DvELLcllV
bFY2bepSRcsVfIYzcO0Lt1SGISQHaLFErhhIpdF9WUSedgHBjCvEYx/MCfy7wc/1h4J/+0tyKVoh
ansRHC8s5fSj2Srhvf1jgnMYj4T1yXQ7Qfp7uUWIGvFV8tCZnKJJQPSYD54ODq2br6wk2evpqSqX
hlNCXSx4Y3H86hQ3vD2H0SatR6wOQ+zplUnZTKIhNV9yovC6h4gBCJVMH7zoofWjCHTxIjmH2xaX
J9lycRH3n+RZNJz6j/fAnX8MyuVQXqd7Y+RRMi96B+w2SNf0PbLHE/CMhQ+l4QdlR7Av8mf0VzKi
mM6H6XDjkgjbutAV2GXu95Fsek18bH+x+/CRdOhVGnb0R3vG/8EKXyxfsT3SNgrocTsTZxowUTe1
RyoPTHLqNhrGo+b4+u7j6Gs09yDyWksInrvq+7qg+UKLkJPn/iQqbgQMyNoGqILh/fVEu6sohbc8
ikYGng/W794SO0/6JQH/fOyV0tzT4Zt4Ir01MF4In8KTt7g2YvB2TSXcxXQIA50d3TZ53+WMP8xs
oYvg32qNmc8cBQCbdYezoqG5Dmqy1gInTprpixWrCyXGJ8LWq1pXNBWGS50IJHKJKlXQCRIICiY4
sIpjdK3dOQVdIs2qqPBiUjVWOQ7HsimeP7uKcXrkItZgHZREyOTZLS06E3suniPtGx7FrBLjQrQD
eEYmBo00qDnUiFJtJcpZFvMLZPuibssvTZpbVVtGHmP/19J7Z+MaRO6VwMf+oD96vCT/c4pZIg6R
UZtWPJq3TaTduyI5dZ4doxE2CXpVAsVtL0EojgPcD6DuWSZRpGUM4M5+uHk1ZovlHjaydfpJ3tVd
GJh2qF4gRJlA1/REqKmtuoG3qbawfCWZQFA84j3GjAWdA+WnvgZVNMG9skhp5HyxlkUP24Yx2Da2
AdC1UJBedQ1gtlWEtYoJEzLUdvu/OSQdy4ouZ5y4+ISoSj4eHTyIz5P2TM0ENG7RTP4mTgZ5CwuT
tNoriLtQQhxZcSVqwCXMmBA4yZjjpPOw5B7u+9et7Zhh1OehdJQEAz8wwg0PFbjJgnwEfyYPg617
yXxLpyt7CWmGieDDw2X1/FfFmxKzKr/iU6+pjIM7y7ppndXHpM9zr4tAdPWJUZmqA4f2AAp0ivO2
l6AH4EHDxCXoAgGBtgOWbsNH5q8pDt8BV07NuOAACzEgSMWnQi+JrNHnspy66NMf+8jp7izqktw2
A1saShenfoBhrhX3mgObATnksk9qxjDFJqJuj9NEgWRInkWZVaFulTDRE4R5C4woDVcPAm3hdMtf
KrvuqbAmjhVn1bzJtJZLJ4tWsXGDiR6/6T1UfynguVNrtxyYPyZXte60iLz62RQ1u8pfyoERdxBM
iUv/J0r3Zs3paGzTj12g23OYotCO/sEb5fqv/cU8sGkYTFzJLyP4nu6LjivRRoirwetqSdzokRGc
tiQ4ui961NCXZwlmxkGOkkKngPMcpQBocqmTWa2MVE0MVeuWRwf4hInX5DG+kmjqEO7botBnJg4C
AEa5YVEexhuAJ+Ubcxc1D2S9+aCVmPINKuWvTtRkeWWKjj+hnJ3iG5Oi6Yp45VKSZKwCqtSLFZ2e
1Un+UC4SvY8muLVDePkCDwme3psgC29vFfOtFXyplZdObzgo8cyKuzMfa11glQxf8a4PrzQZd4Cz
90r6JACemwmWOmGGt3oeSXylAupg5dlwVrWsTJckUhe174vJEsCQsNk96Zih5c8yyCJ1YGMLvJog
GLJBib1VKU47aBk4AaN/k49tS198gltD8MjncAt2mLHdJdY1FjXchmn9fnZKvXSr6/wbdQeojJi+
DXn/sYqMS6b+mWfG4wYdx6d3ig4zAACfuVvbHuWVxF/N9bwoprIMPvvIRKIR70Y4d0zMgf0tV+mc
uS6vW67elpG9KTlxtB1OvxM+vBPmOk62s6FCk5iBitHy8idMbqwgPux2l3B3DIRJULufQ9b0pCQ8
C7JQQbtTFvYHIGcyFpIxtrKpgXOtV3hCPNpMTcQgzLl4qP/kk2ZRpooSaDLTymKRryowm+WyZ92h
2ccZuOgty/+Fnwgwe6BKm36RiSD3+Xi/a7UYhR6sZgMEk6IGEFo/e3vGNe9Hwlo4jYEno0W47+Gw
Jd1u4NTGPnpHSJbzMItPv/qU/SV7acngVpyeVXFoGfeZCGOPanmU/4WEsvybrSIDFg4eT+1kzzph
g/BkvGV5kC1LfqIRTp4ISedc1aDV+i9KXid5C8uYVIbWxGubC85nT9bYFq2r2kgj8i5GehVeveT9
OA0iC4vWkm7n6uikZSsaD3WFEeriCRoUYrMmLoaU6AszL94D7a8spmJx8OA5nPMt84tuLHoJdtlH
ne196IiwwlXUrdPkYi/KUcBQ6kZYE4iTXrsEERfJJ+sExfHHWFGyKf0ROPK4kX0raxK+t6Wy07jf
PG1LhkqXI4qu5LDpV8JFSZqqzEXzEOuhpA1dfScDNlAkG8/zWinz4U3zGz/GoiR258kAcqgd8EOj
TkYhEt4CzvdSSawttGOggAu9w2tSzCWs+SD7pmSjMotn3WcgIAOcdoVzwovwy9y4PA0vKSnqVdF8
+94mJKtkKCHuY2CFTHY2k3X4+B0k0Xjm5A3ThcF2FeuZMBxbLeNModxBZTcwYSOilaGXjevVPU1/
HUrTSCwGu/tazKyzPVEbwiq7o2aseHXCEIl71N4PVVoPrNYoe1MRlSlw1tL8LDGd6nE9ZGtYzFv0
L31Z3uwlwOal2IiVwonplzT75Ji8RGjwgo4Vxkkujl/DXSxXhu2YlqY02oQhC+qVjg+w9mcrz05a
Uo+4jD2gdFxTfTo/Bxr5DaraS55Toj9hAFM1+/MbBA57hjrIgndOQ0b0YWBv+7zNKxh0ekx94pez
t6fjWdBA6adlpkjjRNzfS1XmmECLU+KzXGkesFUBNHamA9lJzLk5YJRm+faGJUS5XV+NGD2/LBhY
rlalrMkcPVizaiJatUqbYGsjEBcLZfqeXoi1On6u/0d41Gk0kX7CKuOWNpeIeZVA0ERDHPcfPW01
TGE6iQnmVmSm0GZPNZNaysNuTPHeG04d/FW3O4peMg9t1N1M0PI7NgHk7pq6iJF+37whoNcQ/gHY
86rf2mdA+AkoYs38Dv+AscNRQbWa45Ytvv/sMSmwlNjqVxkZs0g0aVE6SORVIuVcWwUf+0xhC3U/
qlvz0YCIqfRpv3cK+Kb4UI3dfDU9yqLsSWJZ3R014hbvf9vMgcHgM+VEuAhbj/1aMe9oHg0FvWJZ
N7AB/lZo+dXQ3UuOZy9BdrTWsFw0ZuNrhqYdyA5i+HbTdAgHeeJfSW3t6XUBdLoIuuV3LzTDCsND
dYAqGLShmfgxm9J0p+hqjE1Wes7sgbTE0C0jOTxZ6nUMzDTEgmqVHmfr/aL/NBQBYx1MSgBX7pRT
otZHX9W9we3wv3RUFOO+H0ZKD6qNSVwW5xAQDSrzBRg5k1BbA87PabJmbt+T7uBJkp+6gGsfji/E
PjFWo+CVv/Hg3wS3IHgYur+7PyoPH1wle/B6nqakLZymkp/8gZYgA7gYruQBrj3kAVDpyL7F8udm
D62Ws9DRX0OFyDg97YBLCRw5u7fm3H7tT9qC4YmD2/RQGeUhLU70FW1U5yeM8Q6v6eJ995iO2sKU
zPUpAjtEtZx3JD59q2qge2d8+6JhkDOwFgzgDUWnXXwwjiDLnlZ7UR5fzF75OZIMUbS0FmKdW8Zn
9gnA0Aypf0r4+XBbuPUKKLVjs48iXUIG22xfpmn628ycUrUsMbjKEQylOuq4Ttiyfj/NeItS/Azz
xBwO3gcdyj4L+nBKLwzfoTwKYteXKbahJ9S5McmOJKP0kZ05LxDrpPOH9UqhKA/zfbFuJlofN9Ds
O55MR07eLMuuZjBC36or+VpelFpFccHJ89BJup+iZQXdHA5vOK1vx/Oc6YoGiVpcedLvz6OsDto0
IBv3OVgOnFU5mBDDgUe3e0PhOQHDN7kQ9Ni9AABeIDMo23e9qHa93U1fpyymnzGuVL11ZuFgHvnp
4Vixrfjyp9pmtn2FAe3HBVjv/DF97N4m6aOD36N+HL2JFnVvYLd+eY+Q/8Hp58J+PxYwGNRKmn0r
AAenzZgboDM2vdmVGtgtZNXLaFhG3z3WAnjCo+t8MVOU+5nfV2YM73v2QoKe1b6wLLYaetpBDwht
PWuOKNlfqzWRqWlTJsXH90xDFi2XcHa5k7e05Gg2BmtXHkjF5QagYc88u8DIoBjW7fQberRxWfby
CXLD+eQy5SJT+m3UQpH4Znk4waUBAV8c2dlG5zRY1b64dpd7cIqL4i2wijHiMnJiiwvofwyPRjIn
3yndtLbgdmJC4ZSCnCGHqd6bkdK6fJnKEK+eMLGdCMJ8qiz3l+M8C2DToNZ1CgPACytNStJq5kuB
e7FXH6R3zeC7zpRV1LzI73CpmPZQ24xaIk+jVkyv99g2nejhxm8MOKbjW2vmBBWUDnWOZ/P3zPOG
tTwPDyAJW9NkxHpXkZQS2a4ddeVhfzNntHPhh3UuLi1g/0Hqc3gSXNQUYLsixtFrZ5f54zuQZGrv
Z2peQF0CDKM6UkMbRTirgMSX5zIsU66gawVP9pieZsa9MZS1yaXox9hMRt6JRN4P3E/Q7oH9eWf2
63om3inrSiKMjx2yW7wsYeo6UwL6AZ0iHSrxQm2/yGUYsVf4BHSMC8hfFRZQa4jH+NCoIjjWXC+u
bs9XedIMvLMdswkdcOBiqQ5FIEqsdKP8KN8rSIj0hBgaXJPrFUMZzdyhH+o6u6L5KmxAtzRaNP16
U1qhyUFhkHuJ2aiju6I0seI90xOzG3hmINon+w3O51wTrIQ1DbJ15ym3ZN04Qh+kME2Vlxd5X0SP
Z0ZV8+kwPPQKNcrhZ0diBn6VVR/4k/1EMFV+8OlatbsyhuYLs/3vW7IUQxfr8lChQ9nEiWfJCJrC
AiVeZDve7j15LStHRZRP54aRU6Iz00/VfV4SekzS5RnEJIXGHVB64ry5jXhOXeDwfiLHGjVUWLqw
kOb8uOZsNWUtRmb/km5SPtosXzOV2YHxCzM1QJd7T3BfwxhwnfeDG+vtN0VETGseT5BHN5eJyA7G
QYj+ZZ4UtU1ePpJ1eZZM+ddHWTeV+PHU6frCbYF1ZE83tIHWmup45b/9Hk+D0oV19x4+a8g+M6ln
Ya+aiZUyky8l+0Kn13/yQP4FcaZXhN1oIOPPdYSOyIA2whCfdCzMFtS+FPi8/fTB0gWYzVqSS+Ts
KSTd9IMf5D9t64QqkqflO5vsMRC2atvNTCFcgYoJcAQVDiLxmcdNe1hQAvBWIiX7ep+3DTkdoBEv
H0gABDgT14zInBGNqMoi0BnaMFOdm5NfuZkFCpyXtymaGg45gfpDYOgcybyJZkMFH1eyXPdaU/ZD
0f+/ramUa+7yPq9C9TvyPWX0TyifwWCNpN3Z09kmn3H26fWbyLyIf8261BZwE3TGaUmMkv75buAx
qFzZu2RNxSLRsSpzsGHIZZuVRWoK4veACFcQVpjYxiKLJaX7tErnhUNCYXZI5eou/YhsqC1ZZuS6
S2IoqHPDVoqktQW98SkLPlt3WNR0uSS2/qRI7/cCnWon1gNww7mRYbL/Acr75vhJwNzFt5Df3CZ6
XNKGk6Q7veVHztc9lBIyo4fYDKyT3WBfc56Ys0oBR7E9TsvTy5ltBSz/1fUAcPFQL7ARkUYjLDx8
DYinmD9mqeInfH3j1ggpsX1JF1dqw+C01Td9yfoMMln7XcYTGNeWE1SCae3MrPQ6wxWyyRhdoRrC
SHgakQwZhp4AShDJTrhquPRs5B0RiWP/uCPslVoywoJ82kGvAve92w6lFHuFL7drMpEN23V6/w+D
OpX5sQWzP1UEGYpYbRp0zW2Fn/God+IJKNCcHPngTvL8BItMPsWcPqY9QQcuI4yKSaXFYDz6I0DY
OoT6d1csaX4HvziWnjYhP76guJ4jhrz87rcFkN9pakb4rFEXMrKhR8ja/CQ6IHmujmAtvc5Xg5x0
CXOfu42HmO+bQOrrlnJ0UMqimIR/WV/udUObBsRqV2iNHX0uEWxI3kgeeuRhubSpDM4sVDytAqxR
ktAtbnRxpiJgt5J2AcyWI8Lbym9B8zLW6YwAerYCRf0/sYNjyAFQZjiDpLupepSqjAhlLZ616LUD
PcmH/5ARswDTIuXb3/vcllmMlMYrNQRcNsmGE5stN8+OHUWy0+vRs4irBTZPzUyv+g20xUtEqa0R
nxM0WqgzuAsdt/JZf4e1UKmvXhm6ix9KAduhPWHNK1YTvaNgIctYNkiTvq/85DxccMPCWhG0ceM4
RzxXfztT0Kp/awuASiNT8cFqvOLclbuYdIdzYKWs/zYOtigzc3E59jSeLxFkyji7lEP6qVVGYs3H
R0AK3Aq5+TUS9y51NXKkTrMX/nED8oAnDl8aqgNLfgnqHLXQW7Z1QGzMvkSMNuLr+Xo51IqwJo+o
ffCI+JRoDIwizlW/Cqj71VOkz/ZiJp1Ia1HjC/zTI3PXlPcG3nBGk3sv/mYLdjzhaMDBhW1QJjse
ZCmXCTA22b+sM4D3Wzjok9gvZeSk1BcmXGAUOImT/2ZROVZLE8Y2R0DwlPPd/gzcw3Ly3qjfWJYL
CjEdL+ajPed9E+TcTvuRobIVuU5mKyvwWBwCvlinovq9x+tem9/go8BVvF3X7/N0JYQSdpVvAfu4
GapXimXaMAg0HP5YBfXqDQcWFHND6gy6PnfrK+C/ro0HLCLAjZT37V7fxqpjYRDjR/DL0kAMqSph
JNQceaNgqX45UuDU0RUyvISuAymB8ePmKKpzDzkFpMzY+I7hfdSRugNEMsGmt/fAgcfAOPiFx4aH
5/6C9B1dlTZ2d5GV5bcVSXIxoKuFKhEgvlGjMDahkB5lhLlEFH1kB64L6VmwpYP+RMcMU1efqh3E
Sq3cOQChukq1p3J0AmpMJDZrAWSJkKvr+NBk2zupC5gLbktjW2iR9DJQ53/1g2xIBLvt5j/iqzGK
43mzgHamNu1X702+ZKe+3FOlc8LfF9rcQiU9135wVA49MHSzGGT+ff0zffUL8r/yerKtHxa2az0S
xxk1op7KQR4rkmJcaAd6tEovxbOqGGrbYp+lVgSSp7YWAj3qHpXQGhCoO4DzSIN7ARuka50hWOXk
Y5MKLFrMjOuwTaosMFwFf+N1O/hpTvlmXDaE5eAxIvfCGtY5ESqr9JVAQwkMGvQMLkGM8pd+fBN3
5LHGJlm3GTbcNds2Dkd8VKGA1L12biB16ssecY9LWV28v/2rhcEPEGOM6zdDa67v8U1tb9OHWJe7
AWWO5R4qF0a/41vJ+GykoVKUXo2cukg9YwtFoefvLb8C7O9d52a0iIyH/Upo5U6XzTYkRP/l3dQ4
76U+rea2dV8rvMFdqZaZ2BVQJyCCc6ZtLbZwm2VBMaCUGaaaiY7oYNnc1jvgv92uf+/6FVQIXjXe
5aGOZK26vR9QyVo0JWfTBaLXkIiV3s47PakqlroZ6UplrIvlxW1crWUbLis0skAhUIJlzf8RBPMl
hhFz8LO5qpfRWTO+AGOCVNJdLAw9L6GyasC8p5KuPVoGSb30VsYwaKJZRWd8Y1bGt751FEsGb6CP
RRABD78GFcwljXuTZiiM9avEQmmkcMVQPzH3s/qagZqvoGXWMIRN5czRtqzhw7K6Z2xZq6r58jBY
mXgbqnzTpDGc8xgEr/pjLDHLhoJFj5dXya5csfWny77nEQ1Gtnpx/Llox+t6NAUeV5o1vpfYShn+
kdT3T45Gqcc7wn9FA3xQLcaXyE40DVg2Oeh0y3aXz6PQuOE01XTdLzwxud5Hx8RVo5Jyu3kYdIZD
L4OLKioGvS1YB3zxyc5VndxxjRskoJaySw8CxtMfqnB5x1ag5pvg5SH7LWOHtOle9HkvV3YjqvU4
arKdKo5fZSQAXTtslJWoXh/NgvSY2/Lrp761DZqPVRwZIdhLNT/zMWlcxzwrJmL61gBrpKREXXuD
ZopvDpwx6WunMAX7x8+wl8K0cSc0ErFDrWVOT+GALCgmbl0s5bW+rHSnPLu7lqQHFmRcd5MUYBRX
gozWjpur+WPTFGrIS7c80GLKqI5tmILUz1owO1PHLbzXarm3BcYiYgbVy6sEz9sl3i9Nt5lQqqM3
DWLsMogj5XQSc3O127RdUNXU5D+9K2ThGlU6BS7NbuBigkBHWBHGEn3NcAOLUWQNRrKAlyQ6/oeO
2rgqzOsapeO8fEX+uTHnMC0T/e5jgZpZePIat/l1bt+y8nZyzBdL8m7a9G7Wt326zQu5RECC/Lnv
DZ1CsO8OvckJAP/uyKoFhGeKJhwe6qdpvMzpdfaYH0Q4Ms50LNgQhhdZnN6eomOsuvvA/yjFyh56
Kowts9QKZrzQv/yP+Bi76zvPNcK4cYl9O/zy+4hjCix08dEPj00ocLSULS+SnZ66AMITBHFClkDX
OS9rlGa7mO/cIAuGzfvEYH9gFU9NOvfU9gllW3dwWGPtWjKosDTT+5VXtOjSHQM6z0EbHaJ57e7Y
yOzkWj/H5i8dwboBQcElGAIRrzwh9dK0EufUVmJNa0EUGtj2Ptg6ADEvAaAAloo39r1Rv/bbBduG
6MKyI2YN8wnSK5exC0Jk+zUcR6m1CKt+TlLT5gju/VSagZRxXMIsZolJVaORd6khx80YFFeJYlB+
vo+W6ax5h4LmhrNtWg4d2ii5FB7HW3tOE17V8fzb2q5z97x3DYHiQV7/FGiIPsCfUNMhnInvo1oJ
97dOXvET33rBe2VvMOEZ3uT3aGMrGbKXDFovte/R9WDraets9Ysw7+52xcFroTAJR016meAG7cbg
hl8+lZZrZQbM2uiVgTaoX/FjN2f1SuNMjln395zxTWM0TvpeAam/VhWeYhubKIJGJ7PQQuyrbQof
cNH8m/a5H452h0e2oAaKJbn+fBE9v9Yw90E0l/5XOGpHEdZSUrA/MvvZtRSekn80tjZPz7saGIJM
wO3GkkrQmnA2OPhRWz4Cq7Xtvc0egL7XEXyQQmsCNakBvDZzXnZTecX/Loc5z0qahDIHE9z5gyXw
2mIh/bFK7hr5+SRWFCBW1Ybr5Wt8yn6cr8mu5sJf6j6AO5uPs8FCEudc6frwfCk9IUWNpE1oaDDI
F5jBwYsH+aJdafnI4qVQ0BrZtyBmach/AlDqxkdKnblejTx4HkObA2xWIyMgaPlY/TGp6m6sBtim
b5PgmD7kf+6+3b4QhJepmXEMZDmClS6GU2VUV68uwwi7KURThYjfhIbewtCLAjDUhNnviM7IpGUL
24GmXcg7uR/92qU896ZiU9KMh83pBxqKzvW4gj3/cUucRUlBSjc5dhq9wR7Jp3wCi2qZoTMD56IX
mERAANqACe13bj7M4Nq6RaA+074o1yBo9iUJZEdRtajqM63Zlt6An4rpwhMgKWvXdlDdGzFFHebi
71oMpBgnR6GHptTnRQ7CGEfadpQfChZqodQ+Bu+LtE9leoOza1miH6ci/2IrfywS01HjpYD+n19X
yYti25pf0+vt2fyjkFCy/BnTQSl8xqsBvYao6ZX+f9l365qmqFt7/0/C2D1qZiaF2xq4hwnvBYCs
pJcEmupPF75G/fWc+4V3DD0NuSNUEx8SM1fZodWslRd2fzA4RntpbyPhhrIl0VnTMz9ZY2L3dnZU
kR2QTssGvlN5IF/h42fCShtet/s2dE/apzawdZesb5pAJVZz8+tdNrZPMOBP8RM8KzgxW5sfO8Zi
+eLldoSUE8/xMb5xuW1tzE/dxtH8dX0lDh6oLIIksaEyPD74gidp4DWGuWUsYGjiuXsiZkOQvVhs
E6KY+I9SdQRLAZoOCK2ru1gyFEgWCqz7RXII2I5ZdQ17RhLiZKf63RHldEPUlCaIzP1mVMca7Vcc
p9QL8e3x6CdbtlGI09fNW41hxUT9zMSy0are+pjQ5fj3f9suNIzn+LGQgDqdn0dui0mghKmOF1xs
j17oVaAuB+hZBbKRH6VCQk0v4wGj+vhrmfRXN6hJwIvJc1yf+9kTEkEQ5PycaOo93dK0gi7IKkvD
zuAX0F2yVM6zMYZWxbMaDvnxC6KIyWM2a08XkJPMjgzYqyb4OJ+jUIH95bqiBOE92wyUnERxjYAG
9Fjre0yNaDcBwceLFtDPOkaV0l6PSju5LAJm31PAgdkVtILHgCQeeIVCDstzmkfjbGvNBSO+0sic
ug7AtXhvYO6oNVaJx+AXhG8gpRuULMxdTX/aRtxnO8qbHv2iIB2oivA/6knjp1azPQb++d8Oe9RV
fmeHbBUJ6gVb+VSma4JG5g8h/kJ9HwOQHojNhn8deKx9t9ggAdWlNVrdLNKVbwu8YKByAdQZC7IB
of6QW+nJUKxd2IBZ5kmL4HQxI0Bv/GI9Sd+NGZORGY6diKTvhEEo0en/W1rQ0hW+LRughG+1lSVm
vI9vBfO43ytxHWiuUGmbgoNnHt1I7/Qt3/ZZ39IUGyWf4Kjc2l/1qrDUiHluQQfBByT9uHgzoHpH
KVTNp4JNJ/s63+qhXsXnajTOd0qoi8hom3dfp18pwY8CpRntkmjTUo+HrSYRdHMUL0N1WYElBzn7
s4ZtEZixdmb1NuxZI68E6bwtmcnFT4kUct74w4+Nq4MGOEIyX0CAQKU3UveeEAIw6aTN2iwwyLZ/
UhICSsuyZxk1qUrcMwIYjkIagrcNZOg2oAzqbQ8RAOGGNOaXYYL07WefE3qysoXLZBUUheOMrYji
354Ox6klEDMkwVOSeY04VE4Fvb8NRq3YHAG5iIk1yTuS53F5K5zuDdNJKH+3R86LDVWKuVAuPma7
Vn/EZ5Ib/6bs2DcA40EXjoKIDDyQ5LS6JkVHR6Gyg+gIoRLfjGfC0Q89TPzfKNXlSW8EsHr2RnN1
EuJq07i9kQFKPHnep8GDteUjG9LYuYnzYLU2kPk6u3NDrCnM+hcUqZ549Vq5Su9QtS+UWwByMvA6
5IEZuQrtke8ZOnHhtpkAIqc9JG6rAvf9rftbCOZqU8sNIAojhTDTyBS8PyDCmCvWdgGHsQqyK0l2
s5D8YMf0qVLmK1KmcZClzlXAm6fRv5sz6C9B3bZGQuxOK8vLsNLVBKf+kq3DgtX6IjotJXYrZPTx
CnYbebb3mxMYKzfK7mMIixjAMH9DlUcJ7dW2F2COs5ULe2Fp8Lg9V4blXg9Hq8D+Kejd6sNcy342
AhxROTMK+xq04/RXrUbwyJ0KxeVxYitrem/skUWy0ORo6kV/6YwJ7oHmTsaUVMViWhBuy7JxEmib
N/7Q1fhA9TY2YX5L9SoiV27JWXFiZwZ8ER4PJQVGLEDeETz1H3LysQ9UPtBxfJTi0jmjWCdBabVx
jrJmLQelJYwwVglIG6Zc3iXlu8pLM4pBww7YEiLv1Nvma/WMFBnMPlz+9ydFTKpwa0TxEHuC0Hix
hsncrPFFirHl5bfWYN+qnX3np7QHbyihCuYMGloCDqusZZA9xWtBEtQIf5HRdybMd/r7Vlcf1s0M
1dfVCN/FgWjOy0HCdDNAcjzbLXBJKCbrGsGiXQ75kKPIbfpDapecDQ/8IQdS9OY8d8G7G+5qTi1b
bopMewswPQpbPzqUq2WakbBfNtYtFyu+Wrk+NvVKT/ELwCA+pArxTJsn1GPlwl9nJIUCLj6b5JK8
yQfMoLHJSU0saL+XIr5217eTNF2lawDvv5NulwLEsOjSd2csCwv4Vce6O2cLogYYF18Hx8covp5e
LwuQqBDiy6+zJFIcsQ8unrSoHuNRsw0M748V0Epq0vBWjem6VS14/5ajUTUIAt5FbH1P08mKDoMN
L5bFD0IzwhtLtnhg/rbwlgIzYERYRi2xNbWxGYujWAC0VnCpoRhCpOSBtNvmzg30T6qAS7qVZoX5
dVLXTo9Hl6I0/v2jyTMW7bzXsBu0dzEbsBjjDNUgSBJoHaGNtr8S7vX881ibjOtYRx1/937/Lpt0
7Z2zTkeoaEsSBZlDW8n0JVxMfguQVxeTIVPNcQOsOPzzC/2goFpqGNyrZ8sT2FFNHAeHpIxBP27x
P7YKX6tl9IZeOarjowcTb7yCMBvGmpWIH6XhMfkqHKA9qBlJ+mWu9hJFLyhkUx8ACUTAY8K6Li7m
hLxzeefs5XZy/5l3DYUMLU1deFfgtEuRPzqAp0XoBnd9INTrRazZHTp9YdwfawJDhM3bo8GoL15l
3aFoni5eNf1dwgyDf1XS9d9NpXfWaFBujkQhl8RV6UBS0LHXj090HOewR0RGODwKzGwIBXrrs+c4
PUw/bgjNx2BNzLJvTX/Bje5ldlK7kUVNqodLfnGbb7tMJAu6PE5hPxQPwK8KamnmP8TZWzRT7e9o
eUBc3rZdKsi5kBXT2qQlE0VvKpIwkLJJuzi8FYc0Enyg9Ud3iWH2BwFVj05kcoDZ+XuyOW7VE+yd
GTAAPrBGLYwabZ1kdEcBO+7QTYm5UjdsLcnWyEVdIQ/B7SfLrfaNWbR5VB8L0erL9WBUsLL3t6Yj
vhgx7lwFN2lnPGPdZUmbkzHk2D1GT1wiXBXJ/OhHMkXTivwXxwbb9wVxAMHIG/LJsbx2XPTupxhC
U0UWoOn+XlAPruLx67fp7+IuTmeohwZyV9wV0KP5nH6v4SrqX2er0zSGw9yx11GK7JdJp4MHI13G
qv9WkWVQHoLmyVWaIXz4wQ+o8sIsMVTCFNnNTeTeNe53E2dT3thnskJSoW8bG0+AS1TQY0Cy868B
N/0sXCvW56pgFhuTIP8DDBoqpHoEBnPVuIJ0Q3wfk1hk8CerY/7xBePSW6wBqJgFDvw7xK8xAKB9
i+5Nk7xNETkYkjrEI+e7H9hQibIww2q37/4illHRJhbAawQLvi0A8ivaAZxhbumZ6SiqY57EzIK0
eCYPSBo4xoN/LHpzulYdL121hHKtjlbpTzxaN64x+eKdoizCPT0WvuqgYLWUe3cwriC2RFrhlt5m
2xdDHmeJdgxNf0ZX0SdLzL1QfWHoVQQG6jsMs6VanwZVHd03kYSvb7iUTlVtJKreze6PaABXSPcC
RuNo0jcBQDu3I+m0k8jQVc72Wznfj+iCpnvsLsfpn/akEgHNCNtccXbqIwH2rWBzQfsMRuo8yEXs
Mqad7w7to4O6eti0ovCSPBwgChP763nK7TNq+SqsF8q5osRNXcvKmW2eKhnXzIVt4BN/MKxtRoPT
/3aiXmNjxlz8jTAvPZWH4RF53qOA3CEg/k9Qo7p+0vQBHVGlTAHjBJyU9zLj1F3sZCOw71CcNxuZ
JBuop90d+RUEoxzW0C55RynLD7bS6pCaBvEmRnj4X6Lq7nYoIODGT2grgMysbyP12/+PkpvgP81V
Sd1PomPe3UyFjRqdZBek/+a2G4ZGQgSBv5X4WzeNFizgozoDyeGq/BMUTK1Ti0ST0rl4FzC41aKT
dEiKc51Pb6CFLCm4Hl4qxtpHdpLEH8aLeGER3ix5ciWndnRV2hJoEI/riyifA3HkA3ddHHFvHNZz
gYiPoCw/zWEE2tqEI6GUDKj6hj4k60hPdzVfUh/uhhDiLuHVgr+eZbFzHIKRVU4crt3HAJ45lHRm
2AeFtuzxtrmz7WDbk+xUPrsIcAjImPXLwa45S7ksaS/xovi4dhyaZqHgdyypltAqYEqwzA6ZNuq0
yCbIHJTp0G0KIwBSCEEeAdH4Mtm7G+efIyZ+DiKnzIWWImuF03AVSNSIjF3OXCJIWilUINojP4zI
Mpc38mX1W6goPyQwqNKMMurrKGgbHgO9IcJl+YUVO1PvjAbcFsIEPRhGkNwtC8QWjyPTe8qbnanj
oOUDkY961tJaE2cCMec5T+k2OBoa9jR1GmFrbJkHEhF0jQ2eu33RCd0IWCiH1BRHkU2T6XrlHo0G
B+MNd3XrusEvCOJlAAbBUkWDWCPqgbx26eG5oCqwkT8NpcyyuU0X7VBqIJWRaSwsqQ151kmdhvMA
JPDRa+9e7/gx1XBg5+ATHZpnxACg2yLvZgUIRuPofMdKHqN2gHilsvgZIFzHWY8JtZHLd4ZQkgZJ
TWNnAiivjefcSLeU7Qz6unE6EkhvlkWva+Cdk+B1nJR89fj+kpr75kWC9rgnwQ2IsmypNhgEAK+A
3QMmoBc3fFfGfRQvGkIdI58LzZeUqYJMQFFehdueQw8WAkyq0kIUK8xywMIuKQsdxfIkBwTFuCd+
IxZqXU3AjZKzpDe5TW8yfR8TKpS4w662wkfirsEKYXfYFiwSzCb/hWyNRgLzMJAtDlO/i5OCOO3T
1KOKBEUOv2dGYtvM/LBX/3PumV15IrotJiHzKra38T7+se+1G8yKTbRkBCieE/j9YvCaxVSr4NW4
9y8J9BptgfeDxxx3Ebw7M1SFfil7EyUX0mw2J4LeyEKdgq//P5riQM8QUa7HiyfsQX6Z5j59kD26
oN+xt6LAXxKrBBbNA84M17l33quEII9LHacuJJO1OXsFDGVfDtqBf3i3aQWasQyPg2EAV6bm3FQW
x8h+hZLE506Iod/ao+CwTMH/IGB8l9iuoU2a8RqJC9WZk2i6sNV1KpYQ7c+FQQllvaMD2EKrLJoP
xDhvKIkSl3fsZqdQiNCDkRMfQJLUfVRRgNiSJdNCI65aTi+VqfAPvEMg99QfgrkYSPhXJfUrfRPO
h0nwel2NuYaMfzI7NdsxAiWZ3s2TyAqHFJHPFMdAIgjdm9ImqBvK9AiwFAHu8o+4AbMalYEpTWbe
Am5YZ0o4tXY7mt4KsrlmUe12T4CzApMDWFb5sCGRItk4+8r0MZkN59cRYOQPBI/EkuhSYFgdtuBY
hUdA2ETG0OVZr/YBkvrVgaktxaBa9Lf6nXUlRFnO9Kw9ZtlzYUDLRxIKlb62Saxan4UtVla0kBMU
iUTmXgVBt9IAtm81MSXFpKGnvYE6f6vHiPo/M6ZwerBzPOZNhXSxhPFJ4HW5ODpZ9g1bKKbBnWqG
tCTwKj8beCXyPYXBhE5n1Pc2yraH7KCWadMKdCgDdmuJJ4It9LZyNI5qVzuQZ+lvvpbfXT/++SG5
fNjNnBUhFn2bpjsQB7HdcF001LlNUQB54XNQ1lzs2jqQVTDgjZkhzU1A6Pm41JjDON4jTANSDbrE
NfQioDlaEfNl2+pQlLW91sG9lm2XFlKv06yBehLnQN9J6781LALxtLaQynpw01FL8LOh+NyDW8lS
+x6hFjgMXj40vgYzJch8YP2eZ6Mk+MkA8Yx+ibv1R40H0ErvUaQjbLI7SMg+S8idzlOoUuZebP1/
pu1oWW2ZJA+xRQsvd7an8wejYakCdeff2THfjFkTthKJiVyaI9/fej8uUP7mFVVcuufpGH28MoJA
/rG3QlvgKyVsM+hxW/boA4ajzLiOzmK7Se259x92vMD1je0YKgKODB/3wNTmk+7PDOLzVy3j3RDV
8mLwmI7BPScrDYwyOluCnYcbRQ2l+TaXcHeMKX947RHcZgXt02XOGbyV/86jiPZbVdZfRqwSRlpJ
NwdH9aghAl6ulJEwtLoy+kyCQYqYeOTE/0SqQdYPbbok8Z4Gr9FieB00eVmM/fNSEtuK3IZTwWHS
eu/gqE7lo++fB3/j7Qtar454O8VIT5OCv9Yj2fjdZ62a9e2l2PfO7tZnRswO5L3bjsBYcQ/xW/+t
ipKKNGJgLhs9PlY31JuR3mN0Z6VKnQGh2qJIyOMjvi21RwLPCV9csu58O00QyZsZlR0us4HIodCw
vtpgbnPKkSp8crH+FuRujs3/OyDOK1XF4XaFSJhAmutJMxgP+r7vvMEecFU89A7VQjHyZ6rjDXfm
Es/VB8Zzod8iWWttGSo2QY1KU7HpwctC0xL1xHTD9r/l4UtExi4ZHG18n1gyqp3Yi3GzoA3EeHTZ
DXtV7I6/B7EXS56kqrmBRqzknFAQf2G9cv+uSMzBtvZIoUI47YwncbspLFRM/v7z/DQCCgUoxnqf
XLZE9sP5ZKbsEybV2B2kyhIWAPPjRcnL0oIuLmmp8gqvyvX2vTCDu7UvSdMncmtoz9lOLzJ+3uwK
p8GZF3usNGRF7g7+xYLVpvE/t6ahgIryUaP/1Z7r0t1+zSlzL9UfY4xTMdqHjrkrGK/A7OutUR3d
QUEmqNQ5lMFQz5hqaIPKBo+qEFxk/1cdBbv2Wotu7G4fuKsxbox/qSWJ+8+EIJb+yIXXsqBzMx2D
b0WsBAQ1SZqWscDiYZbLJUUWaQ7y7IWMOmLNrVd/W1554q/s2fd1h8Kzhn4itLHlUlZ62ulsRB6+
CNVWzT2aZNl9H7+Ef5LhgCuE5iN2qpJKC9mdnmF/Nwm5OqtHszlSG+leGDWdp7qtVzEdoITIxfC6
lOQtLrMk7bzRgIi1IABmlNOQ/+DZGlrdbhr5eyCQT2Of8ewYif38XHZ/WeH7LL0mSXkZgsLoHZ6C
Zgo7nfP8/M2KaeaTi88Z4qrxm+Q1K+wQSH+8XQ8G5TjqDXMQjgwq+YY/rC7nsM2QftXBIk1qa6nq
wiF+OljZ0pxXfPVDFh7akt7kOKGSUwluggmy+OEAlRD5Q4h+MtbcbDqYiKOGEinTnExYkhRjLisk
zyvqwKKsaeKAFt+d2eaaMIwU45sFpxGGPILjknxSP7QoMz2bsriisMJEYJ1niP9xrIVWOSgAUFV4
CNW3wL0/ZnQCFOELIwi4mUVor/qapaOGqKgP/SgBDiCG7bR+WkpgiOt4kckgjpv9Cb8srOzIfRbR
g4CVO2kcZqVeLcVyAy8v5+DRQJB1R+vqmM4zfVKtMMCZ8hagPIdCEn7bFdF3auKYAkzcS91nsYOu
yU1044eW5+Fo2fruEi2LHaIQa/ITEq64gYxrmqQ1znBcEicYZLtGUwS3NL80V4q2miThPNgHO8+R
0lemytItyWeYLTWkm98N3waOifQwoWoTKKzEraWND/chPemO2goi+Zoc9yiRMSu+v6ptKjITC/j6
BohbVYoSdmcgasyBXwgCvd1YicqaMxoUyCKp+CUVy+l4vEyAfEOevtgX8d8SbwIKQ1QobsYLnihw
I0qDaTz2X4PFvgQev+Ir8gqFfYfUR2PyJOsOq9NOBds4ji+8xSAdBDA3wVqtEtRPZHohkpSxAebC
QutETHXqUW6Xo8PYtGEpuaVhGEi2AWQOfOKpvenPN4KFlEZmjKj3boKJZQts+To8jiJVNN4albN0
Y4BUT0EDx8BOEbPwCePidFAjJ0p1fKqj21WSfRi+85BQQcpoArEp28BqKhueLpHb6cZpWVgHLGkT
Kl385agmsoPMztTwhiBH77uRKy8kl4r2q66v9QqxYJuMIGxw8ekzvfHW5NOcXjXnkcqhbmEoSBw8
tiEerXY3dYlIouAkeH8eTZbqiE9WkAfJIANjJuT+o6jJhJjevKbOurONnCWsEIC/Kr8U5+CCRSQj
f+2s/vffQhJqA7USlmjDsrazloXykR5jbFLVKU5fyeyRdeh1HQNKUZab6DANFJz3Hwgy7MJRkzGX
7Mb8EMpV4iEjX/J3A/nbxLDaCfRM4BRh9D2TC90rEKdAQUn8ZY/S0Rfq4DSaZDPEelCepNO8Il5U
fVXw5qmfLh6dyrsa4M2eYlotli7OEjvYO9qrycwwLJjeGHJXuNnbw/0/C5Edl7dGZwCwPijSRtO+
/I6DvarRrpRus63F/ybGj+6Wcw+0l5Mjb49jbm7dSnHvEri/DI9FTXI0MhoPgf1cF6DbyLYPdqAx
sdEC+91xkZ7KCJIx9wjf+L5/NArProfYnOuqpZP9G8d1fum0Ek7TRk9iciTxrdMq6+PosQA+XPUK
9ESG9WjJjnmDj22iP5hBcKfFvyuzNZsKBCpeCI9hiC+HTh8wLe7Q3GeB0kkvk8tgPfEUSSdcwTXM
SRyzc9AKqHyCm3foEKUo0gr8KLjGnaKx24/X9zvmATOX48SnoHYH33pkspk9D1zHo40zEPRO+fle
h7L0WIad9s1wO6dDHF0cadJTVSK5sFMUken/1TS3+g4vgzWwB+xVKeafua1wBJIcqOzwXOYYat1y
I3USVunAsnBWHsZXp+fCXWBjbESw0DJeDUdzpr7HD3Aw93O03Bc/IGHR2SLD7+Ec6dnBte6nQcZu
RJvySGfgwU6LgL5cU+WZc0xR3EgWrNhtC3osFpTyeOsjUtX1udouQsqBN4xGmBdqb9YGpTERXS1W
RdfcBXtxSyLUuXuvvhDPzAUIYxfqm9LuhFQKTEGxcvokkQbIi+7g2LlZQNfXm3GmgGYYmPy0vJme
+z4bCke5SQyZL/mYS9RHixtpKalGhkj48KITxq7M+LMzfbUrwuEYCNmgi4vrBifWxUKCxBXGZWjT
ttiA4RnzNznC0/5guB9PyuVPl3xkcCvdHOQGfLq3oM0LrjfOEBSzPRqy2NH5lfeorjCY4Hs7qGbH
btr0zZ+Musq54AcSXEnNMbmfhnZYHrNpt05/dD44yPEWKazZ2SqyVu6/NQ5azsSrONSc5U8y1zx9
sD5Q8HsUtX9BWHUuFOov15aU8Fa0CDeCjjmM1poWS9k9xIiUCwXzsClMpal9L5bIKEiC/YW1P8Po
BNlKI1jpqD7e/xv5wzw+rOTNk+4yJ2fKkPLGl/5IDSjeiafuNCtMKCiC4wmF/CBpAu2P68+1l1QZ
nbvyGn73R9uKBbaBgsKtSU4lTk6YmqrW5BhLfGn/qSzkp/oPCiNjBzSxJWCvtmtkj9Df2r7u4O96
nhAVvsFd/wTmm4rmhLQ72SwRbzbBzUiPsg6LyUtcwx2KGKod5nax7EDOZ2A+WQ4Scu8MdNFlaT51
167ladV28QvDaeRZLlMGJNq/f/kXfVSdHhzAu78dkph1pux7OQsgQgB0EYbFcPwbdrYRhKPm2QOL
4moZ7dKTp0BPtt4x4L5YpubpcANjI9cl/G4Osp158pTtmHnQz38Lt2ZdXc0m/JrNUu54ZRVt0In2
ndFZZYgrusxVRwigU/8eoYJJ4/B8ofP71yD2n7VCHe37uNZI3sTq1i8tnARHEOkei2eGkQ1kya8y
KMB3x4NEt8DwB4g91BatM+sz/AI2rpvy7zGkfyj16dzDI1ATGMti7QE0fb/WZC35tqPcHvXh/S44
1YuMKFpoxC08H5+FwBe6VG1o+fXoivba6qF53nr6B/xNShsmHiAUEAFjHDChTJkzmFjT+M+0Y4w0
lbCoqluejardxJ90TJ7gQ0IYzmVd/P5+Xg9abqrpoZsm32mfy3QlqjXCp3ePmVK77b0rjrtOSA4G
6JAT1de4y/G1AibqujMX6vRvBLeX4I+ALOggVjN/oWTnYkVuy9ZJUDPZUhsa/KoKT2LW6Yv+0j41
AyWv7hvdT0q0OeSne5FPNZU0CIqTZfkAC7eRYEKMkoUgXw4UsxdvYIf35y73D8ST8mtaoiE/v09n
YQ5nKqgM0d2TATTB/3WeRCxZqqUm+dlkoKNewMv4FDSODppE0b9NgnOTHY9NEjiHtQ9VXGQPbZD5
6Y6oW+qszksIcMHrMXCN1Na/vjUYOjCsfHT9qT8Z4VITJ4SG8APPva6Nk3tzByZcAI3exZEKtJ1u
c88KIZMY4v4zACa/U/bMKMo0kxsgKtG3PtYzShP0lrtL53h0huGlUuarthag5P+HOsrcmS/89ou6
vCL8Hw81JJVysPs58ApiZ1F6zQc3ZuYhKZ+5XCZ7kk5ygaVk4nFM1kuMIQxzMLhcDjFVePhdTwBw
na/Vyzwk7ePCm6oj5VlJHpXvovy9PvoQ2f+3L3qCU/0+NTvdfcmYgpH4a6M+ffbEk/sD2JVy4LiV
2Oi1agmaBEmO3mbTWx2jWUnWitqY2r5vlaPfZ7QjhnUuRDfI47Cbu5yAKLNlyna2luVZ3GHdMec0
x4nTg/jMZbS72JIsOKuA0WJyCryK4DZwT+a9KJ3VOGJWnC+MHVz0880ZXb1T5CvFOTtFDsUMHYda
xKVYZbNodvW6A5b1lMWRxVjGEGj04xFp69a8/bhi9aKmscXu7QSMOoZa5JjTeuCliLPRfz9tCAdY
4AWGfClxYRCcuhcPOyOW0YdDehHZ52cRxlxUki8GdtUtzDM4xK/uhSumcRyqIORwNj2vq3rkzmmA
t5N1h3/UlleAn5OkndkSwD1ZKPv73Ck6kpQqAJUgTMiyVmJi8guDPpf89j33e/SJlncKWi5kB/4V
x6WtSWOLx79XG9r9LRDJeCT7A5BDFwUEUXDcON/k3b9bD5bH98bWcn48xV+YvIdFF29BhzPJD9Nb
y21Arc/4zUjUyuvAuY0zVlU+etm5SXzaMfe+wrTyRUFJU9TN0ss9RdzQwCljew7B0IQAHaLhu1Sw
SNEngqrHR4ISWsl7LKS6tZl27RnIJ/Kx72ySiG/9iLpvl6REpys9HinH3dHIq9bmwHRv2DcCuA9N
KDYw3e/cCpUoXywyH/7IHQBhflOCkuFL/4nyIC/ygxzgHKNCesygQ5j9cfO6GavuAfn83NOO7xYc
qhtVyMabEZIY1y1QyOWx8crjPasJICbWXMlC54IljR6EC9QEykW6U2OTL9khumNS/YrwMiJVpHsQ
BmYDgdaQfjR3L0ayU86Yrn9wMvaFLs7xUC70bnOTBUy37ojL5nOpMwSt2d4Q4PJhhuAUNjfunfWN
kA+bVaFJ1Eg93kOA7qY2KZpcpy30zrPxUOqIKaBLQ5wJ76yPGdEfYLTKxcHDuIc2WEPdtba5ZGiD
Or5FRPVVdvIDaZZGxIqfS4TPDjxFsUNMf5dqIuuDen7TlYhsLy7xGlw+4mYY/7azLaS0TptSkOiW
Jz8dMkNZX2hjNuhXROLID87jzkcdWZtIYNB//r74YTvjMYn0q+feM2WiCsntxPHmQJRmlUMZkOE0
Q+EZOs4k15q3aZSe9lot8lQmy2dTGrYamgkGvoUWfdVLmGrCpQFlZC2QNTc0qdbYjSu5rR9apgwe
zyH6edZpKvQdg5SLWyA1SF4PrEV7lCyp/LF0cebRKIzXgoTKBqI2xOlFNn0ZgpRpSv1kK0pfCzGu
yG2HxAcEZ+WarC8t7hKAVG99gdtQ+wZ568h0+fy4xvEqVRbtGASQ8nnifDP6m5f/ghR/sUfm9vDE
0tGDXlV6UE5bpQbhoCLLX3SRVnd8ESUru9Ac7rvArcTieCN8DrmFL1FK44MBSnZseW10I3UfKsrb
RX+u8Cz5+U3iDI4gpmKS9JGp5jqYKybJinqrTX3MhxIjqDJ72fd00IPPqX6j359hnIr4wRNNS48n
MdCYR3TJK3i5LIvvSMTjJBJnTFuSg6uqfSjJ3c8QHUTpPiUjx5lf8zvfOGAMpU7d5xZJOfXpjgRJ
UiPFbQJnpsYbYVxjl14k5I5VCJ1O+yr+ScnZjxEK42nXhh1+5DEodiocoxf7EIZm+5Y+fzSKQ3hy
HMpMlbpimi+KAZylbnPTeI8ksz+H6Y886d6kgShAa0uaebdAxo1CtJ/+ZAAaLfbyQj+Hp7K4Y2PI
04MbOTEs1ok49ulPwQnudDhWmIbHlEMTKgJG5zTvjzx7906FncgiMI4HtsZBMr7L6QEd0diAiRcz
OtzCU5QZCxHebL8glNUXqseKzfdUBPYk7FkQntBM/azh6ioixCUQ2CGGxlRn6mbpW6VOW5xlgnoE
ct7NpXo3cCSl8X4nJ1TqNhc+ub9IcU8IKdEiYH8sF/rDt8HFo2wDb2SRESwEMKYsbeVQtbxOH83N
tEejYW3L+eP7OmYT9ICCE3sRKJ/69M+Q/U2aLsJCgjY0bothy5/IKvfpxBweJQyx5IeMALTT13Eu
tG09ZDfYBv7r50jGluYg5gOjHfm7zdQOxRdcllvJYlRqr1oBVI3I3QHWZL1nNtWJc9ab8XGvXo52
zzWypz2MvIZQryRX90m+OidCFmuw5r6FT4WDkE3agTQuZrt1I8DClQCT/DdHREOZtmxFztm9SndS
LZLJdpGx/MFU8oB2ZFYbd+w0S654xpVmgKj9PpRHMAVvn4ongtr4o1TZTKjcFyc0bvuDPrsWN7Os
Fi5WFomuyXHe6fe/MFmqPG9NZij3w4XMiShS0aJA2BTZURE4/dYRplCpJdC6A9VRkQgumiutmoQq
/WDPh7PUuHbA/TbrXs4QYurlJDN7hFR9Qz1F1bGWuufRBQrbgvVeWO3HbVo6pyMYNQza0yWqEvFe
PZTcwzXqpc0yicWgotSr79V4fswH01PBewrNDDEbibsz37GMNRJ5s2g6wB9ap6TcihVAgkLtJv/B
Rdea8x59hWZz39nz3yHLcemAtgSo/5k1ifX7vhRT2++Mdlk7yRoqSW7WCN0XvZyqfiOFoERPc62p
gro7iUoVsgt020zD02d3HjTKqjyfOfkS3TQ1Drgc8Q5ZWSNsVh9a9KII4T5JsOqKPoa9SZUWWEej
E+Wioh8K7bl162U0/ap6PJQFAuwgziW7UFa0l1Fqu5mju3YEsiRjiKTmuHoHecyinLkMdbdxtgqq
+GNtZKfcJV19qH+6llulZh4IfnWSEfAVVf4v4CMBDVumIE0R5Nvp5AJ0ZnibM2zA58eToDLB9EKk
4WhgKBDVXHZX7OD4P8OaW7rHXaZgivZzR9ik9krZefV9u86CZpOtABH1T2y3u48UksiRfAWcCwz9
WKGG44TicHpIv5Ro7ClxDxerDImhdY4ERabREY8w+36X6m7NGoIis6SURFlG2jSUwf1AUB8hBSut
CZ6giv5e64bYjVwSixwsmbNrsNWR2yinjoveIWsm4k61fnKixdA1YySH0PGkuAfT+Onmyx4W3Fql
M9Fb3C7EUT56hRA4AMV7d/zd5UEPZBSYhL/LXVEiaun1E+sCgVwIa2SeAPihd0b1oTZNDovOCGbM
7mAgBU6AWmeakkGoG33zu+vs+nurpHvCsUCxpKi5Ns0mcC5rUDVXWjFvxeX9QpxKTZuUyCvkAdUp
04/7UARGeU4VTUzdz5g/oKKpStE1sgJHxurHvxGOvt1bMaHGp9o4HbDFCbaH2yTvQwMPYoPQDdiK
IdxCNRcP48n8VxCh9beAU/1mq5cEMlCw+zldKZhSz3uqUzJc0QbL0CC4lp09Tz3TtuSLOt4FbAA+
FdfOk094KufitY0hnp0eVzvEZ08FFN931N7HzkIngnOOmj7dQW2aKCc9dgh8G1u3SGDFm1O8JYAF
CqxiJZpITboMkrC0SNP2gvBPqj/QFgvIZhRxT6gEOSknC4OAbJPm/elRBPEulT+/eReSW2b3+fSH
WKdR3xZgdr2EO1aQKLWWQ/DkCq8pP1N5pt2TasDy0Ty47PBJFt2kBf8hZKZVV3nF9GPE3//4UwAm
Krmt0ppruJpHc4X/8CKWB+6SausWueQlyDtlhFjhSmqmi9cK84w/e0T1l0WJX7nn72wqvK8Wnj+L
GK/YXF0hhPsLjXkj7mZGJzzCTA5MnwDrhTWJzg5fr14PMz4RhNDKfGM+DwzXypqAz5PfqOhkqe+k
QCIYy42BFDXVRNpwGvtOTeYJKd6SvM+YfvTXzbXVyRsC7wMilTL/QzXt7BE+6yVd/OPRFOQWQkme
GPLksQMV+bkgwp0vsbvgvNGxMsPpYvYV3l123Lo/isxPOIZ28sLMjftYU9dpwWdfXQV3RQZgTd7A
3QDr5K/IRYLC5jaN7VclJoJkk0OAjFce2TnR2uxEQz8gazNfS3Q55yRSdIHtE9Kfw6ltdAMYqSTq
/OFRUrDWkTT8B+j1Asa3TDSuJMNDxnaWlRDdRQppAeOy4z+CxcHgylBw4kpo+7iQ8t1K3w9Uiw4M
RzoJ/ldBLYmLwhRNVVFVuW8jAFc14RUjbcqnr8N8fH02QNad7BOPoDjLcFCjipKMWUupYM+BhCOc
VmXKAz+CryS95zt1LPoy48RdxBBMmuYTAMg+CV9bslLYc4laTZZ/ms3ysORB9w4mb0fTNIBYCdDK
V/P5vE+jcFN9slzWytvVPj5vPi4vzBqDaZUS3AAMi9hV8LkusmBEYGQJUasfW4uSb6Tr4E2bKEl0
Ja1kYuVAQjEK05Hn1euqHTxy/s7z9sqMAZMde0RlZqn7BQ5tYxoTQzBNjr4bru+9mvllihKb/ZUx
EZ9pL/SWWDpcKBdsxfEmJUz8xpNeht9CL2NoluU8LvxaeoseGBykUJR/ABMhp7/aOb6+DYYqkzBg
JUMDV6hO9tYX3p7fj9m+LLwF0NpNqHJN7vsWbf4cQyHYyv7k+KTZ3DwBbBxR2lEGpWHlgl0g0LMC
RpaPwCV4EzF2YwkS21G0x/dN+KQBCtRL1WhgYV2JiJEY+zJXYWetQ2sIDztmv+v2WtIIi0zwMaoI
bkrsJWScuf+IsF1jhKm5kGoB3tPd8MzMRUAoBuspkeAy10YbXt2lLJLMfOVkCa++0NNMnfPoT1SO
4mGROYwd2c2UiX8bPMg/prPSbwpij0iuOD4PM3FMF3W9FAwVIUt/qwKKsJ3WxxDHR/Zwodzl5hE6
rHHglr8kFzqLYDT7LAxVzbCu7NBIIO4A0nTHXQ2TPXhPcY84rnXIjiCP4ZLX9jRi2u93WQM2HuTN
3qHTaWfTu5kHBiz5XZd5yUJWRgZ0lvpltq+QwAfuFXJgM55KjX1iuiiBlCDc5X4LsJHAw2e0q4/y
GSU5Y86y5EcVdextG97rSDROeEICMqxF8cer9NQSAfRXyQCbAShZBd5YCKO4C9Kw4PqQUEs9yy3Q
11Wg7JsHI5bJZHIDNlwxiD7elAlAEvki4FXW2rEMdNHq9CLRig+/cNgwpMiz3vbEsGol45nZf5ip
RTiUgfgJEOB5X5/ytlqGHQy3+2yJFMu4eyHiz6O/n7ipWusNTBNjpq41e6ruVMT8AmJKyoj1azq5
w3gUeQ4ZkQGE2xLXwUIbJydt1dAOZptxuiaSl7/XJ7faZIA5/D2zioIMIeUd4RCtxZfrtjDHyvB3
j4jsX4p0+xO1Yv6Mkhv18PM9T51WOk06Yy5spYLdxnGwUFVxtNxWeA/x508rEeU9o/FOhfCZp6oQ
RnT2BFYbXYaPrtvzFid32nD5q3RhVpyVmk2K+kafVB8aodWu09Uec/o73F/HefQq2RztqIBlEhpT
tPV6WRGos3NWPisMoaOrBqevPhYVztp7+1JAmkivuAs6TCqOlOEwXVpfGbmituyqmWB/gHyjDp7t
vOX00g7+NAVLLbqgUbUjHo1Qd7D8kNS9n+qvLDveJW3bWqbQNVxub28kZwx68bXRKQj3zsD/1cWU
IyVZKla/7XGmC3kUs7zDhp+snz6U5/JAnde6c7MOkA1q86vko6WW+qFc+4XN5JPJLAx2uvonrqVO
9vQfYqYLis9qoeobgfICdqC6xJY114qF16VlkRGYhq6CnhXM+koxAfcasIdBVsvU4L7TdDjhdvrr
fMz+sf/bHK53bey8OZ6rpmv7tEV4bLbsZmzTgVxKBsdZgLuwFx/xDx0qTgP/D7WYbuXlVqlyxZ2y
QET+Y/a56WePDgCTzqvoFH8mp2rU+zjEIspQnpDAM9TCtfrXXNAlHvtj3LqW/u+NuZAjD1DHIBdA
TlnKP8QT8s3oQ41BevadjbXsi3F6OMayqZGK9QP6pbuVVtRQEfswVXCkN+K6FG3XXUhTz7WyHB/j
UWlZShgtRU2F6BI0+vl+TxorLO/WP+E7EPIbgIv2gYqrVsy5DRleALw7rGGTPH7nEgKGVvDlabVt
BABTixHY0g9+1FhrfMJiNC9auwos2/xdtUWocmk9aLLDqp49930Z5YXEtLtwsfZaPbM+4gE5L80C
ZLcPfBFHelUcriVdjh1e6KIIZ8m5CO8U4CmtKpaej6tf06lnSBfrtbb2cJ594oKlHNJxXq7rNKt3
cQdeRNdKYvdtPKD6wpml3ZDJDCozx6D4HATVt+sRx5eyBLiVUyMnlYraw1PwQRhP5UsGViXHzGNr
ligKPiGwOBfCrvRLiUgPfqOA4MRFliMEk86Wc1+vaUvlUUplVH+kXWiH0UbDR2eJpqG1EpemneFC
Oyk8Y75HJPkAm9o9R/F65aBuEl0K23eFJrARpBHRsFEaGZsJq/qWKgR774iF0iwsAgb5g7MSnjgD
bnzPg6NMdHxWZgzIHRlKWWMonqzr9LM4yp+rkbdwFJeQKKGdKyu8r8hCsBTfNsydpNyQLfd90pDg
RHuZSCJRLSKRO2ricz30AbWjaGBmDrJv9JrZsWiGNmeD5A7Dw1+NInz0z7pH8rXsccvSaV6aKxPm
FeDir1kWX5MnmFE2iQ7pYxby4tERTEs/5K04jNa+uyYyH1N0rNCRfxJvGdqM4ozJEoowHvTWNp/m
/bZtX/yhDOF2TA5q1Wmi8zaPA0ytZShDSMQkvhdno+gBfC9wvD+jevMLBb2s5Qcmg7SU2OR92QMi
OWvZD23iSdbfr1JG54foo0S2QzNvsYfdElBV/IHVXindzu5ro2I04Qlsd4Y4M+Ks8QFdB1NmTVeB
uy6c0aaQGzav2jOqcEhoEI63OJ5OaXnleiHQgsx+1bkUT3TMjG7YLLuW6WbKFFODVgQq+xrdZ8Bz
8RrwLqH7gOy1E0jMsTn0HwZUnCFbF4YGlby3XVkq1KvtbNoRE18iBPC80cdRWT+c7ZHXLBd/KPNI
pGF4ThGzDEqXeqvqqiP4ijw2w5rG/V5rRby5N6LI8ZiHqBgfHlri8cw1ZZWRLRg4GD/NdDDXy+WI
YqSJ9GT5cVCbZAsd3ZA0Yom7zWwHD0wz6I21KNO5S+ik8ZQWcIULg67T6qkH/sb/g93pZ8fDMAjd
NumNM69qE6iTx+3ly11OKUi/Lrl/tOq5DTR3hDs1N6hu3CtuM6chGFiH1eeC+dsf8W1O07ahiZ28
ZYoSRo3m3V0UZFgSu68aXb5nfKU+VSUBsiRZ2gSIu0ttKbg0BKKF99yzSiiwDXP5iJPNRWTBXvp3
CNN/3mnoJXoG/piYzVsoZPVshDzNsF2d/VfjtHQ8F845FTkz/e/+OO7YqJ8+jvLQyP5yNFR8bJdo
CvprfMiqP8yI2j0h9UckFo0M43os+Ea1+6c1sXd7VPUxpoe0MnGO3AMQHF/dUk5x3YKAM0DCcCnA
eJOhqZ+ris+7xh/mTueYAA7WV5T5v6Tvax7DSwxnHziuJe70siWxdRJQ3Ao5uXwfq3kTzFgGR7Gf
pPCH7/n9wsKArQJA6F+7hgUBEOm3JLeMzMKOigx0Ma3n6hXrWnHOgfcbmPWlxQKEILsR+9nhLmvb
neyNTPkK1B14a/aOcZ7kUJMfQWlimdC7VbK01ZxOfCrNAyVi/2iq5F/NpevZzGbzphc0mkgHXiaB
ZW/DsXfrNCXVMPwF+cLOSY5UEz/HYYCTNxGbVUoiyJnxqYDuDV+bH4XdV1E6wmjmJEVY3wRIaduU
l2GX4U/jbKw+6zUvsPDQWJN0RXsJXbuq3Ip7LK03kHoYCKiHS8I/FtZ022+dPikFGSclX4zCYgpp
MFs9x/gts8LdKi3NrzpesDamehB+2sN+PvGfSmcjk/td4Uuj55NFCMVMYRzMOli6c6dKQYXx5dnm
B0lXY5SLbRefTZX1a5vuo5n/s0RJSwPOnsYqJBZtYVbwbG6PBV2z76Tz1ozXT+kt7tmqgehTqjLY
qum96TLfhq4qnJcwPf7FxEv7Q/0HdAffVBKogWDtCpRJclXL2SscD1t2JUspXgbcTV8SSAYfWy0g
BxWoPFiuf3jYrVc8tewfnLCLRLilih3beZDbUMhqv+NLl2JOz07WMrGuUcmv3BSdcIoBpL8AX+Tb
APCFI+w80Lc9IwpuahP54G2ool2NqNdjPTZvBoX7ARKFsZpKbNvW0Grl8kU+K4mmv/FKXX+XreVW
TBv8vwd29Bqvmn8zBJqaf4TsolHnvari1JBeALqWs/dLmL3UCyeiTCISbOdFE328o5Vb/aw/m37W
DYrTLtXiCjQEVbJnzWNi/DGhdZQRAa8ZQI7fVOAfzu4cHi9N9s9p+arP4NDQJ8WMKw7MJ2G+r+c+
bhkwGcBCJkP+A4ep+dc/0B9zB8d1yEPph9XY9NUPmnsDKOzpQqvIpY0WjJOPYsf5d08YsuChi2Ep
DTjmiWyHaTS+f6TvyLXzjgXlsC7ClNzW9dq34rZk1DpD/5uUSut0kubEaEx+cxDFjIC/sAXiie+t
0RmdX2exGHSmUuWco/5flyA/Iug8U0t85B1ZN8LM6GnrCBTWs6VWtuXj44fp7LYV7R9DiubVWwTe
nYUyX9vjDs8lfNpvWuUgbyPG/sxO4G/+2krsh8zFQFhLnL/mEwPm1EEp+vyx/Cw+sg8ciJ7OzzqW
1svt8j854js2P+oh01k6AzzvtMTkxRoNS42fo6DuJoyS76xGstF4MB6LQn3P9qEbWZScYwvThKt/
XK9mRW44MrZJAM56V7zXSfXapB1dFWOOa5exbYfwikJ1WxQjTPlnNVs+KJOsuDMUkLiGNIoaqs3X
J0QCtTfe9mPMzZhpIZeq/4YF/alNztNdWKzDGgcjIQeMVzvBPyNVpxvkulB6M6vp5MwEps2BTQJf
ao2+Da3p/NB2uTYUAhVucN+bTOo5sRQ6KQyqpAy6HbfzlXSGTtFhHRLkiguuiSIzxv7fsgYhGV38
YooMSmtu5//fLetyscoMqmhrXpv2qa/1s6xd6fEyqFCAIqZA+Wv97staKxQoIeXSh3zeuH+pdxj+
w8nfhVcNvLL4TwOrzhSu1Gc587espsw9C3KYh3rd+7iHPj+txGLtV1Z5uswwOVheIlzeSpSLtv7M
3HALP5SetlTwQW8+jn1yuyaw2tds+PE3Rr25NRJwXmC0M90AdE3Pb5vcrIXhLbvaPhG9c031Szv4
0+yTXtAztWhhkKF/w06IePBCgKFLV6HQAZLIcgTvg1X9LRzsBfJJkXdE/tnmuGVZJ34YBsUUPAdJ
LrUqafl7qctEt4oA4DzKPyr+wN3j0lXDhqClFe9WONwh8rpHEVssGPq9vUOBuMoSKZ3AohKaOgp5
TTtJ+lZutOhJ2AoMCh8OsLYT5S03iFpiEzFbXjJULow+g2I7UTu0/GnbhUM9wGtt+QtehjCPniLj
E2Y1tUHMNzf9uUUE6u5f7lU+SUAKnidQOnu9C1zP3fzB2C2Q4Tt2ef7i71q56+JwnF3dpsfLPJAa
2SSZLQIblO5NmNF2RyjoSzyRekWq65v8NzovAebJMXyA7lzIg2ejv743HDXmmwUbFNYHVU6qT2rW
u4WNlJeaha9dfqUnG3ut6U+eJLEeef+fbYytSOkO6O70W1rJHgx6RceILL6dIZl+AhsdBeep+2i/
7I+Da13ENHHLLa8CN1mgzB5wW9E69dI3T+FdjALtC2kzhf1fAxKNxZB6ADqs1cyglzdWezGkdkBn
q1eMk9kzjpos60W8GY4/PpwQ0fGkTbDx6InIuNZTF3keOxlCJLxonbHN11dgxiF4wg3ifMWUMXHs
p0SfiamLfhAWcQ1GsQLWld0Pwa3GvgeQE2IXNBdooifpnOc90d0aDm+qF6JNZOGupazXuSXMPWXR
KU5U68YHMpOj1QR+7DR7vmlORqaAEJbYpHLjXZaFGbqMPSNXKUnvg/aPgmzQMkiGJae8BjUje8xT
gt8JmZ4d1BTGd9faj0qaDhy3ppx5OO8ps4Fg84YWooEs+OVFBVU7BESLwOa5wbeVDunmUM9GDnI6
Wt4NkAFoLqFnDtsTJgX2Lx1w/9b2pE1qyUahjq8GXBKUmH9b9B9xH8AAgGETzXVoijC6UxCIYdDr
Cl56ZMWU8RqlPDTnduLuNq4QOWYMBCJXnrrKgO7lFPMGc+eKI3IATIXOJP5i4xavKIzlnmhfeYMG
YvcMuop5mPaFEA11OQHMfJSSOM5EnYf8sC/pkJqwj3fPvyzA1c4+Ffywmg3wKQN9Ijf0Oofu2euT
VxrJKdsPulmhtyeNeaZECyYQfFXHQkAOCaiXzRjE8F/qYxBn02AwpR/NKJpV84QLP+hU4Seha9gL
te8bLXWZdtd9Mu7QYz1ds1xr0vOLtuTJkwnUGL2tKGCOIhliBUltzndTQWQ0/f0xysIATB4fSVuW
VPMbAI9Y0A2oXO8poMfYxdGkEoUyAfzG7zKQz23h3wdbHWNBes7JYdyN3YN+SO/9jt4jxNGscNAg
DjjylvpZeKuzZAnOvEpNUE87L/g2kV2ihHlDRVjUlrNuO2zSKTUHTIY3DUilVyBnnkB6hUQHyyuR
eWBjraQvSY9z95qfc7/0tCzEukyDoZc1I9Q1RMqPWdWI9ZEjB9DM+4v1L7iNibKTMb6trRcETef9
8ubx1VCiZS4h3QETVWgwfyH/FzCz0UoEVS8LSKbW61/21FyIsIfe/xU70MXCGjMs3H4L59hbik0q
JrMp/hLzK6u1DwfRH2NWfquOjrKpXpkowUXI/vJMFF982JzZgSHQZXv+pW9cMjc2idFKkk39yqn2
fxuaCwz5XOsejascZeDGFKQ0MCbBSvV9FVnjTvGIRZbWGcwGP4snvYu0Jem54BxAm6eGIq+p/+9I
U/oXTWdx+qn8ApjHckYlazzRE7BJ2VTmXtoeAuF2BkXtT1/UYvJLH95CBHoIAq9yWxS7whApes/W
oKWmIJpRdbiScUZKn7XDHWi9ZvIOyb/kbwEBrH1aZFRd24DX/C/Ut0GvTEt5zr2oRtaqaG5tyBur
3xXABdWye5Q3R6Pnrc/XqJha2HgSOERWJKn9x3/nUW0FfEAT3thpPe9QfyWy82YDpAIykeZhXyoQ
dvyOxm4xxfn4HWkVc+jh/oUFhCkUBdvurlDLJ17YckfHsLbOFcvo8hq/0zkH7HJDNbW2kXIJcAwy
PP0A+6AfJ5om/l0q49dDZu9AS6o7pQU4tUR5E+Gi3Ba4u4Pa3SbIM3OFQ9L2ZxzFLle10ugl7W7x
V7xND9UIMWH1V9J8zFbbYiQBMMdvaHf4AiBs8Lq6/19M61jXbbJ/6czwC3xowR8JHipQxjodo6HP
wiX5BeTtbdp6vmx2q1PlCk9RzpPy4uIDJv1zhHypgeg4p9EKi8NSXyQVdXlj3X6qjycab8yHGlE6
+jPlFgsSwI9GuDY74F0SioyVUzMSvbff646PVuIteUf0UWVBIuJMZ7AY1FLPPoGVbdD52KAlLnvH
ZAPry+kalIK7mAdw7zNl6etH9r8o20PvObhXy0BPWWHFnbhpte6JJjuleLTQCTDNQ3ZVDzZCwQ/X
kUuF4tHqQ7Qzp4MTg8Dxzq7eZUi4FDB9fap9/Oz3VB77qQZstxEot9ti7jL+TrzN+VeAe5PYZE4v
Vbs9EPb2nitI35miSaBUO1D37O21LyM8jE/QdcPKN/QaXlMh2zOq0NTuBcriKiAUTAGJyFQjrD1Q
qWA+Yhx1gC+Yxemmmo20jKhlRuMKnzrdj7TbmjTEiRBP7LePOjTXEl6Q833W5eDQZ0bu75w53UnH
sMv+gZjNGoJV5/KFAg4uMOWMFELiXklsU2P+DHby6E9E9tGTXqm/oZYQmXVxU4UkfDQBKpuVF6Wo
kYqQhnxCr2Z97gOBGDEeHoBVhkc78gKKFxLmfMlhKjvCfHkck9Zz/FsB1q0hslm0CobtXZv1BVvU
tOn7s51DIvj1MMjfQMc+e1sZJulcJAyzJxShlUE3+ot5yBL7jJNPi73fls2KICox1Q1h+iX8H+uH
dDynPntldbp1yOuoGgsHWiI6FvPzSDTIGoQtDjcnkVfCfUO89+At4ITPIDbcf5jFK0AB8IPgS69K
5BTzWrCkpRVS8qDtR4/LSX/FRM7morih4SWWr0af+wto3JuCXP3mqRLk2aT2dtLW/jPwEG6tYXdn
mvb58mmvYhyuvlr1AaeCwqDQiiHlutgufmReN0pfAgoonDztDmA7gG7RalOLKrKY0SfcdupsUKy9
/7VDYWbrhREmdoZVXXpQnzqphOOcapeZ538g6oBDjgnY57HDs4iteJ+DFHYK0345iEo9uJTL12jd
O+WkJfl1TTy8u+CaUCJjCLwl913rzNPt1aTDJYghcBMHHEKzUqxbJR0kfMhgO/VAPRIJ+QQbeNEW
sDraQHSfMJmAXC9fzxtVhqH77zBfOILg69CPGcnBVPLnjIiMTeS9x5lBfrf8Py21hpavPhbLl4TH
YUbKhBAe1u08O56VGBLZVvI23wuaFC4BO/EKWvS12vlg9u8+x4Vfxb19YsSbcd4017D1IUImB8iV
wKHSYLhBe7smi4qmX3PcMpDR7WJq8imOsI8GRnxJo3tBmD5iU+3Oc30QnSYk6dhROvWgjzK1FsPN
PWfB9de36/gO5PrCGk809ptYzU6RfNd16jyTecopR3gl7JQrIDm5r83QJf3c734k7KW+qDiqkmSn
fToTdA30U6FcZVOGiWSNo44Kpip+wqlk4K21gBoJG4W3c7uunXQ0EIHp0GhN5RQ86wGDgW3AtE3Z
BxnrkvzTmIZN1FdhiJiEVYM0WUbxKlmiW8dAnTz82h3KPdyANAW6u5IhIYalMCJfnXfA5NQg2TKb
QyHGujTRo9QL4m+m0NmH2/FV3Y/G1/QrF81UOakm/vpNEzthP79ZsSfhC4Wpchi11+RhgvZz/Xtd
RcjPzjJdJE9fEQsffOxG+g3o00rn1LaOsEfY0NwMSRvl1B9JCGFGJtvAj6NNTbw3S6yk0p7UY87d
XVAaoh5AxxAaEZ6Ww0L26mr54PQgPNNAmjpdh53/fMXASyMLoAJ0A5crTMemhR19gs9zeNIgo4ON
ov8M9cXo72IUz+kW0acLA3Z0gN5vI0a4CjKdHNLpEVRxSVwsmV2dUTDjANTDj6pnkltcSjxMTpJ6
Hsvqt2g44xrt0XOmj7Wh6Zv82scQfkUUdRlxrxJfKcYxirQ8z6fx2CP37LwVpwH0ctEjI/5CT17/
C//+ddcDn48zcssEJor/ytP587gnOSmdZ6Xtvi+A3rOZ+U31J2bVccWNj1i2l9IbNWuIXTeKj93u
0W35MqROr7ERaA/YKqXAPnYSiFmKfrNbAZu2nISIFctainU1J/GrouQfxpfEBbzR16UdB+guJh3f
9g+k2dxWTfmCwAnKFGjzbAUnNWblneUNNV9Veip2WFaJVqwSrvFu0dBpMHQM5zFKdSLCYMH+oP65
MoQH0v1opoTRmKRmxHsp00rgEKnCMiQ3f4wCIs0LjueHu+5FT6Arpx/N59/5I2O706rvvi2BIGrh
7vL9OtIwPbe/Kir7a03lDUDsf8i/42HK+jhlFmysWN9vFG2SJ6wUwHyxeXDRxp7ZxBscea7XPgiO
Vcyy1Z7Vr5kBL/V6ddFP+sRqzexsftgXXgXjxRoNiNdKTsRGEDN4P4Cs3E1nd7EiITZm72AgPUcb
L2WayJXqOS776m+6rGuV7tkmoGJ7Rbeb0cMcIK0fTxCtdWaELqu7HEF9Svvy2LEDHm7qJpCf9MDp
BUE7VL5nRDOpTu2Pytxpfc0h4Lq1Ns3KMaF4DGfF7VRkSgYgXQIPuHxJCurNKYahQT84n1flNHgp
2rELnAToDeMTTUY+81o6zrMYPOEE55polTHWzO46xaDyCBNw8RIVM2Fpe5K81rhnYFYRcj8v4Aek
bS/BkaBT7hafGTG4uAG6B8o6zXfSPjyTr47aEAux8U6sy0F7u+msec4scD/hb0NuFojzA7wF0ImZ
MJr1s4OIFmfJklP1YhwxdxXsa9twooM7uthf/xJnxB1JO3IkpvxaA1/8g4iiAiDUqJrESkBnPwox
0X7gHeGm1kK+ReRJCAjDKn1Z/4nAVpnyaeUykmpNZmtjy70tgnYERKaGY9bj1Vqc/npEEmyVsvvI
75BbVSV0rE10LMGfN6oaUuC0JoB7jO+PV9ciOzEYi9xu36uWD6TBeEZHTVihjJkLn48C45ZrVZM+
3EY15s4XKLVo5DvNqYacXsqhJHpaNnpalZ/gKttQhy8EH6HumL9fDFOBgUbXvXctkI/5oJ4T4Pa8
WXa64f4rD3vlcPcXICORsQSY0uYrGIqPkavhjj04XYxDvOBbs0dGY/ifgPp0KYiHNbdbcuGYef//
WWoOnN2Tp/HZ/cMIjal4oSZCZST1Vq+dsivznSioMeZN5x4eUsH3N2BTH5hdVTFI0ps48bVjsmu7
KgXQYybuSXhfB5IcEcpp2UYm4IYtDkoJqFIMZl6ekah4zvQaLeEuyS/Oc4RIPcjwm/Qy2CoTT0rP
puRD3Zbm/KHXN2MbwZmAHp75RTxViWPF039bnJeH9iq4xtDThIuZ87lLahexjx6FTZP9yThB8hH4
yiwhFRQpJ7rbI57lD3YHxNiCMFQn9UAjhU/tvODOkWRQvRn2lO4U8daZ1qE223sGufFEuXXJTway
AV9DUu1AdtbDBUFPYIpDUz7jUyqtvF4YQqyoeM6cFqDImTNrFcJzWj2RXK0IkUmH5NR+IHcAb80o
GENEA/b++vlUerdONFuh0CGxXslfRPmP6BKBPsbKsnvY8TOtM4DZAnteJZ9fZB19mHeq5y4kk63V
4s3ypB74EFxYBueLowwiqnY6YbRXg4l959IBAMLvPFPcPFV56gF7lCOvq1oqIfXbr9//nAnRNNVl
iTOwS+PlVqO7MASfaZnHqBJbs84GzH/n2eYnOepYT6Egsa/SslxZSmnylQDwkaeyPdMb1fHiIaOf
PtcXq9Yq6mhy5AJBTjFn1V9gMSNM+cGJsGW5qQtmJAOehGWwy1N1kfZjY2Iantmyhds6DY+n41BS
u6Kp1mopBtAzn7GBG6y0zSIFbaRQP6Lj+7iR41TknBUvXNWXYAcMebWXmz7ZPZHArYvyhenC6tiG
bwyyZ8wUTDqGB+H2SyuUWIbw3zindlYQ2cW8+6DjGFnLQG+/RCy0v0kaexlix1CgIaCuWNhqhETU
6oYjfcxSTX4mGhFVMRx3jTFfvBz1bQb/a/uIQkBSnbj9GkcBqT2ZNRHlpIJ9giBUaz9DevFozyN0
FAqctj93n24KZLonsrvdoLV7KnbJIHXu8+tAX7d9Wi96tWd18TWB/OupuhPqW+LLRbxFyXKoXizr
rlpOOSjIkYX65WFH+Jol9Oj/9OHosBZ5cxljtkQBDZ9c5deKoak9FuOsO+M/9KF7esYJ3O04jxGP
25UjXsP5gr/Kiw94ByFoYLImrdQp4D/tElxBC8G4sVzYqndiVAqJ6/h4kRoiScMUtKAlDiexqOyG
Hv6jZ0Wme1wOtN0YVptg414UX7Lo0iJNAi6eqU+BFi8K2Qa32wCr3vp2fiFWt6HSt+5B5OK4pL0p
MzJvCzt94HcmEKPlI9uiYbm001Er+s1XA//Xf6bSbddYRJ6wFnHuUu+/oFLIzs6PScJfvgouVUGC
IgeR6yDLsp7M9qe4JAEcapy9dR10Ii0CNKC3dc//dfC9g4Ca9auc1QyMe6w6VJOpJT5d4f4Y6haq
IA3CZrD650rbo+1PhkYqjg+BiJnc9eqACm1Cf6h0//GjxuWRpVEtGONaBobmhJidBcRKfSbeXdDf
wSs2EUoDSAKYuN30Z1jnp5+8trVJhZ1+qZSnt7IqZTPh4sGZBN6HXtpkF5g2XynaVv3gDLZQXy/L
+vSvWCsSnXtQ7n4984LSrGpBFmdnD7EmVEpVgns/hs63sJtx8UkDvqa4CzU2rAsAJVQE+dkASQ0w
hOji90iWI+iU8sY07kBN6S03AwY3tG+NLU/ao7QaTiD4eoarss66iitnAct+0jJA5IdxilweqIaY
jNYbQzEWCeOYgJyfl2LXw+RhCABn12p+MeTq8E25cz/05Xa9fKphsS0LCPVC0Lc/Nv+sa/+Hbino
7d8UUcm0LhntlG1E84rLfWof3d7UzYjw+0eLfhdJLUru1n3dfnrlulOUHrtuSVfYNLesWX7lU9R/
wumwK3VA7XcKQVVlFGFjO2BmQxU+PQIGRhWyVdo+yvnWhpd9/kRAUpg9lS7ZpxriIup1FrXtvSpU
7pOYWTIQw6Ie0T56mEzyIe938Vh/6sfcJKDBzQutNRTQcIVNjXFki2WSL+UGi8H78dX+uVY8ZbP+
o5AAGG/Qyqbz/e9TvA80bb+5Bm8I8q9Ax6XEnmpU9eyOY03f8V1linpLNtW6e9Bj0eFrBg31Hs7m
6Z7eo1l60JBtLmGRbh7v9EqIc4f7szpwUDHXItjQO0k2+IUCcfkahJP3Yb0TJvXmWb7zCrWC4/Q+
LvIPT6eiRi2GWIqubliX348UcZMt6u0NYchK4M0Ayessqy5lKyz+bPUNlUnoVmAhtr6A70nHOYjn
kbJ+xn/KMtd44X60MX/w6w4tdJVe/b3r/O9ZVPkwY9DvibRDuK2SvzgxNJ/BLx08HirpIt4geDMO
8EAk+J/QZ0MpK4j5J7oK4Aft7gZ0C1QIbo6GtAwVW4X4hf70hNBKq7vN9muw6euB7EWQmVfjdDsm
tnW8CfaR3/oRVOTw3DWk25iCYlJWiR+hnGUVjKGCch0Dsjwp9sHSCY/pSkK5urdP+UmH5XzUvhiS
SbJqpdV3UNdIx1eBUCuO6JNsHNOjNP/+17xZKm69PfIJPplLjphPrJewcmnjKMDjRl2XFJz7SU7H
RHbhiVAyDgXfY7n9KBk2UuWEvBWyNhziDjB2QNa4EZYrvMl/KAh0n/plHe8lh0qBOF4Lt/mvnmdK
VoPloTGjXswfcAZwFDoRlzyh/obGzR6YKu0nlq6Jryr/xMzZO0mNTRThIOVa+mtWinS1PQqsXg8m
+sEwXtpzORrzZcJ66WJXyRyU7r8K3aaiFNJANvXbqA2v6jWV/XZPasBVD952QuY5PJyrLu+qPUC4
yCJX975zQoklGNTkmszZ37aUDzzLHMruwtei7ZGj2CeKRbD+44xN1fCCdMKF50IcdUnni0qxHuak
cNb5ueJ9YxhUsGMgNy4EW58Wlb2J2kKZOezFpacQCUkU5dnHGMbRzc9wSNUzvVAdzYq8JMZx9Rpq
0XAZ9MXtwAVDHNQjWLsa08ven3aZeqMEBFJ6OQrMc1dENc2/RZ97LRpw0Poc+oQmLM9XeIGxZ/st
l8jngFrsq01wALI/IL/KAQLQ8kN1vQApv7/Ay8IphH4oUreXh9uWPEskbSbcQHJKbFPuDB6lZZYR
V6KgLuiyDht8CxGk/oALisNZ8RjJKjwkscMui9eo9qcgV3cb3Jnh7UE2kuzvK6dusc6PhqBdBulf
iyMaJ8uOUiPI6Bh8UnqzdcY9HJ8wXaAG776KuC9N2ZE0KytWqjC/fJJv2NXdZ3fTz3AZUqv/7Epp
xauXNarxilQs4X4q3cCcFVodga3YvwTEqVCcjxSG2D9vvuiEdgKIBKbCt8qDdLzPYGsbye+ufjM7
I9QqyYECzCf4ecm+oddP56/moO9YkaPyZoei0nwzURtFYtyMX4jolfqxJOcSdtoyrpLSgYnuPHo+
lwnsXU+irVdncA3ykQdOBHxLAXmd5ldaDf1xvUMz+BYpPxMmk07ULOUdsvekV6sCbNTu7UqT96dQ
MXyfz4VXPdoXSfbMW1HPZUS3u2EwsAb/ZFJ7AKTXnK1hHK6ubYiCnHqm2ViFyAzUsMmHb0Mo3sep
9bHP2CC+Icj1hWuX4qq8u1N5ZC9Q3Qu/1nXCoCR/sk6cRY0CgkggmvqKBt9fEC9r13GZxDm/D8fi
wVD6KwcKXb0CVXdgl6++slTouvVmZN3tDFxoVFoVHEjOkKklUcylSrnZ6exhpVbTa0P9pVW1glNb
oqBusejiDrZfBW07aYowGAKLSJotz4TaA0USThGxLP0AweUJUX951NlQHRvmzHDiVcG+2kXZvyO1
Ks8Q0SUL17Rct1I0zbC6+UAX+N7Fq4fiwj2Q1FvgTH4j1r4OnAvFbVTgTLDzqM9xIHlSSyN77/lX
goQldECq6AQh78cUdO0xMJQsrd2jF3tbzTFhQTemnHzUciPMJ/sXrTEMBIO9y+83jvIucTniwjsc
skbhcOBGMtwBD2SYnCzUz1M1Xgxk0XL/7+T49hdSOvPqUVsC1Gbt0Ii+rTnl35s9ZFvKgx3vlQmc
wE5Mmys2k/it8OurUhBmXQ7ke5R3RFVcHWdBa4u4PhgvNv3Yqx+SjxI5UC6SkN7YRdtHWNRAymf5
evq/VqUA8I9KrAR8gHqxX7wyOUUOZOa2SIygS8g+hoOTkwIRXMHyzSxEM+u/b1nbsAKp4i5NlGsq
a/sMP2pk14O3EJF+8ag4wUz/nFIRywx9ZtY/Sunuylsf03nwTEFOqThQx9VFk/pmuIbPsyQvg1Oq
A/GfiBzHnpYvI0z4tT+rdi9G5CD/r5/7MiBFxf5QeivsBfly6MwDb/l3MQ5qmCd2fHh+/8bR8ndE
NMyMKVOLrVKNL3d5y59KAMCHKo0UW2nYVgaH9rMzxbJRHuS+5mYvNjpwY4b66YBp3RJlN88fm+hC
rzP51t/ealS4YmtLE9CP3LSCztWtIxJV9taalSfpMH/Le7Y1/v6HTL946yf70OvjzGBmi6B8zf7W
Sr7hx6jYsJ3LqV48MxSF9RdNYnBCsT/VxKG9y4gHkmNLkkDRjj9VBHDR03y2/sGVYZKfwVh/MGSu
5U12zCGtB8Tj21/+aCyW21+HZxhAcUdR2tS7YeWcjpgqGPc9gf0opFEjCOBLiFZnOKkZN/mFTF/5
RoRi/qEHsEFP2ND1dZ59e5XTVenR2KFoAxHvGuOIAoPAyNBj+3J3fpvnjdxhaF0kzgh7JCmVjXr5
x+H3Bz1RsoYdp+h3Dp6iLj2Oi2E8SePfZQ0xLHkLFOFLIlCnwVc21/CNevREN/xiV7uZWB5TMTaE
M3Al9hnhjBkdwwmCRBf09fNsVWdU9xBsLb2KiLVFyHzY3o3g/V2mBseq7G3gS/m75gdTEQd+z8qY
GzuIzZpLGrg07dw6fG56c1R+pFkxB7ZLH7qTYfxKhhV2CQ+Vu1FY2xAAzCwIpmcodMCxg3w9How1
s3YVSrpRiE8FIhdHEZk75mKrlZ+QZoFu1nxIEF4uhFSUES4akX4fjaZW8M0wqEj/e5F9LtgcHk0I
NvmmypBs90ZoTC/KeCF1s4M+WqIYvc/CGgnj7uZVAVm99FVuvLIi6Il8bT+y5icCw0yVcKJwz/QE
c647tPjKymtBLVeZ27+O+hlNKQY1TB2JkTlozvTt4GJF+7pwUMKDZWaUfykUmvMQnw+p84J/kbMv
2GUJR3x7yH3bNd1ZE9YkxTFVl6NB91XV/WbsHgRmoy44TiJClHQSVEnG0PNBqzr44goiA56OtD8v
X0HyarNT/AbH0XJmKzYE77oFw889d1L1G5giJCGvXPNULsIweKWlGsqTB1nm0RBc9/0r/oseV1zo
tWTGaWCVJs+uKGkDFxoLwBrD6YwfdKpNKC5fRrHqe9cG9LFcDWO49V7nqtjPmfoSEaI94JjDZHok
FsGqTQbdCFjV1c+pIHkApFwnEc6pJaF9xd4x0Lt4ZZd23beCaakIEHud2EODlkKC7w8IlBCCr6E1
RImDAN1TrqVwo59xXeQb0aU9ECLMZd2fXpsFujY5XzLwgGl7hIUiIwWhUg6hxi+RO1F8vaShwRDY
beHdNRPt3ZagHrkXKog3wcqkuDAHtvzVrBt4P2/w7yN96HrD86+kRx8D493d9tS6PojwatVCPnYr
OEVDpiodhzWxHf/54iOymSsHBs4WlkklnuGcolgeDB0p8kKwWm8JsvuNKqjQUg0RWUoNMDGFwrTR
UK3zok7cWKUIjawaTIVf4v2xaCcb05HGnCLXFX+M/Es2ci6pqvOWPImOt3UzIylGALexFWbcoazS
R9dfEecqUWS67XiFFNQL6AvWhyCbIWEPYfDuy0/tUw49WMu51zoOPqW+dUMKmWeCEQb7pyyJ7qeu
I9Pe8iXsLPa9iToqD50RMelh7bGUadINz3RZkU0QGboiEzOwdFm+OGuUhZqqNPTtp5rJOY4vqk6Z
b2Uatc3tFItMCyjAuGSKYL0VnmdMjYgcojQ8KbLG6+Dgu2lu1wZqT5/GukBVuTsWXExfPQHUw63w
eFEGMBtGvs7znAD6qRRgYIrseNwEkFBDWG0mfKoj6weW41RJvAxrd2MtLZldRmVaGXM12chS5pyX
MR3Vhbt+LofzHXqL2uiLSAWQPux8vS/cfTCUZX5i86yrNHc+jfcUz7zZMMhtetYGNhMnB5oOdV/y
4PtlwpqxryGuL59mGICkwd0yXc0Z7UHLP0LrEFCOiOvPBtyO14xP2GRiDxpJc5lA2I3KYxfmd7fs
7IY27Sc6waIo/sgvEPOO5qrqNdqRyriMF2Z8LyEf0Hj40yC2f2kEq25sw0+PMHAEx+FqNHOeAZKy
FH9Ljnt/PgzvNtFFwxBsPXpFnWk8SJcfXcF2CbxGvyNrQX9VQYi7k/ZezYe86DAlNtlr+HaSzc2x
OfPzPtXvdq5QiUoBo8h0/6u5QXC70JVIv+qXJaWA5XtGfBQK8osjEu/t7fm+syyzfHmpWgDJCzFF
8LsmC9yiHPq/AnaZ+bZsRLjqz3hCjyDL96EVVOARKlyuzXKDBwIb/8mhnMG72Hd7uHinXRhpWIS4
TnVzt21LIb5YMOCYowx9UoXsMtTAqP7QVfZ2u2Fslg3Gio0CxeUumNPFn3yEIiop1UzoTj0xwwm3
GIfkRKwg/0nul1wA2F54/NFzafOhOtQjDs8UAlDpKuQGIYhrYnSNiiELS8UgVdll2vfMgh7wwa50
nngPdpXfUYQZAr7rezEgrjqpEZh1+s1XkCbY+YaQ+J/YWciB/rcZHg0sddPHGjbNQDvWnW4KXs+b
MyALdTA5Rb+/2kjUbYctEkZ/Ys6DKDLp1UPAr37HxHz5NjdpDaFJTDWcQTLmyixdpVumEiAxCbRq
giEpKgE4LL2NLYOsuifpCnlHEMDFCRgw7tPI/KTfuxv/aI44fLiV3WdZpPM+gaAmshVxhLCMZYae
ssh57zW3IwIKZFYqVNMPfqfRtYGxtlonWboK43O79j7h1SlR3t8TwSkGnU/vt8X/gopfcar+GORf
Ecya7YMIenaTDkvh/NWKid/k38cbx0Wit5rdMdE7OrJ4HFTtnSHcHwu6NZfkCGZ+FhjeaqtNpBhZ
036o9mnTZsE8jT1TZE6bqhkvuluce2plPFChID4ai7Thol/4m8VzcWaRpqciOnyQO6cE359ErbXV
0m7+Z10qT52zVdSn/cI/JpvjilwQCh7HNyQuAVFTzRk+o4MTEOLtg/Q2mjO4iPopdx6IihanCVYm
BxnSddMGbuUsA+hw6y3YBF2EFAXE+EVy2GIVlor3JDL63bYcrsRGvtTFbIM9u4+Gai+UZsB/Zx6d
OOXJmhxVOG0xbIO4Mga0r1B3cRNyJxDVJAY0ikLNO3RGG7h22sC/5xl9x5JnRBrdmnfVh+2v9QzQ
4uAWkoPIdLUgjVnaajNChC8mZPBA9x6KCwRbv8J2K5GNS/uWexdYvWpwv9zi1H9IHhCxzF1ULqiD
xWRoW3PNrjmqioFTTObQudfcSzqXbET8VhBhDXJMxqG4gZE1SAt4cL+DQpdWs6cC8eqMidHeO1Wm
OEEvVoblfXRpd880yKrcOl8uSpsUABLxC9NjeFf7PfoOSholFO0yx1mwMQXV+6ix3Z7v2UAIXJ9C
nhEfOq4znRjudqJRpm2C7FJsOcIyrXG7NYBgGPcfDsKuDIrYZz3F7wRoOQfy0b5Q+tDI950DHrbe
E6ByJXzcqp4vcp8e021Sbg7GV2SKGH7DGXANaturjG/sUleEst2MLzrs0TlQyAzoc3G2FudjSSpu
WQxu3g5pWLhaF/TGnbkaL3fn2ggXUkLbbgnN68WGJ3NqNtUExpBt7y7STlmQfkc8dKKWvMgCFjfY
Ub19LjZ0zIf4orn5DDlS1tv+c/tbryitqueDVR7yf97/SccIYU5jfY4DCCkiI1HILTbJiOSURmqP
rpzDR3P1VcKQcU9ZtwsHMJEIcQ5NfvTRfOxWffarPeTwoTPG5dq8mYvnr37hlaQMwG9UUQ46M7VP
hZf+UgTIOlzQWmwGw80qYw8nWbOlBFN56IBmRr7aKkgapz8f6dvjpQtQ+Jg7QxLbKi2nBKQRqHdv
csvg7rk9TTe46DdJqf44QLENsMwctQgzIp9PMheG9WpUJpKW10vkp9sHt+OAL+PB7c0Jdp+/Fhae
/FX/JvGdR1hN2/Z+FSAOeIW+zmYl1twHIarmTUENSIlcGC9oA1eTvLGqb6XcEgI0sgYh/GCRNzDv
Vu/kQs10TGJIzwzqt8wtAY8tt5LwEUwd9NXZeCqcH7C2EZ3xwXSTf5f0ebHoQtprJnXoGkIJOqAO
3X54g/gVvPvayMCzGiq2BO8QBcLV1t8X4IhhViNAqGfLSXPdjvkG5PY4bbxfUN4fjxgRFeDkJs7y
/1SVhEJtyAXuSL2ijWG7RxqUc3XBuwAtaP/snEF41MtH3h4m6hYOBTJnCVS6LmxFRtNXu+teKky8
0E2rHPeGwaxrHwvGod2gAp/D0P+DrTRwb0fc0tBwhnRwwrbd2Fo/hlPTh1Npml/M6qxKE17wgACU
lIbbN2yY6RHwAooeawE/gKeMLIgLWtsgbnKnwjd2/NwOJGClu9u1cLWFUp3xTeRTG8qnjcoBV3vX
OEDHStUl6aiRYVuqA3tS4HSPB9FBAuUkxJttGA/oQoYG1SSd1ZHzYGN6BxHJnkdhACr42+4seXhl
iRpeksXV7RSpHFDvHv4cGQEzN7srH7BWpPClVoPdg0+Qmc97YTn+ksXsmOJOF0Ga1wa/uQUbw1S5
cdEftkFIkhJsEkry6YHR635jbRp28f0EopqUxRys/v/336/WAIjYenWwxGXu6rPTpSdPN2AuxwUu
SJWFkRlIm6uelmy4J6AjP6L8nPHYyThNFMAVf1AdOzCt6AH5xXP9lqpcqpLxueaHA0FetbTHgnzv
BQRda1gjpnvlz/z+gvw7s4ZMSkfGW6xuSuxZzyt+5cvY9+I/LduzsSpD35HBqLLkIWYTxa/A9mQB
FCGIeTJDRzff9ju6Vy5vpWR64Ex6J1KRiBavXWxCefBdylX9irZJCDBfUpT4uUWltUL4o67QXcCe
eGTMjSmeqr5OukPx+k3H8WzdJ3RiCMeUxlSBM1saQ8mFmXrJtOdG4NhE6J2rYpmb9etuZ3ezAeYK
AuFyPFLfQpngdjquB7cYg1zsCldrtXpfFm5nfoJYY6ilkwDCp+0edkp4sRFjk2+HbZTX4lWY9Vcv
GCinuEaOnXEHLuFldzX0IuDWQCyF3zZmif56zmoNiiIOUau5LggYE+tzXCa6D5idEOS9PlO9uEI8
LHaWctF+FdIiiVWUZbdGMUQ/hRHktkRJjhWuuaWeohv4wmNbr4SqmxKoIqxTh6VPgeznwUxRn265
Ujr2gltfp8AnzxgZgXxDuUNA/spHkPOp4iplI3wC7iyr5zp7nuOP7QgK7Xax6n6gHD12GjWTclOB
kquIFmc2WPUDL5eZfseAG7sMUKq9xeibhJqSfwCmaIU17/T+m3MHM0Hk4rdH/gLZ9I0iRvV1Z2ZC
TlcsA2LKSe+WeEDgmqmsZLMoRgaIaLXFh93/EiDkhUl6frook3nRBPIYAzRtsUcMwA8KnbpxHvjp
BdM8t/NUbUTZHYXQt1h0pSxWtk9a//HUjTUSONB+MHqS3Ns6XzObSg7sO0s4reJTPSxYBZFoWa2Q
WjhkrwL77E3eXfrUshdYZp7K4fLQhZaxkx9dlJDPxpp0kn/jijgOMTTf2L4EWoGtCjocHjuYQLXH
BoaqBoxQFSRc9YaYzEGZWI1T/TcSm2qEimu5dvuosOQ7uKid7UhFx+TF6UMBgaacVx0kXUFkejtu
hCkdPS1lyDuZb/o/s923Ql6xdb6ZU7wCw0ANZtn93d3we50UBgoDmeDhmQkGRoGVOxeXeUOYh6S+
+trjI6hXIHSe3+iotX6pHZJc93SEfwMvdatBTgJRcIi8W3qvUMRQQOiixK6c1mcB8AFhPv/gYnbg
8FxmwoI8YGkblcP3MbBdbGGWUmkSIjdP4e+Rw6AS8QhYK6HI3MDi0xuiYp8WgK9+l38q5gsw6Y6y
7GkfJZ5TrLZZecVTtMwJ6vv/7EASGaIl1rgVT6d98fmqi6lJntxaxII1a16g7khwkgbgA4T2QFyi
eEQ393OTGA9LYJxjzyjPRGph6bjidr4AYhROiVMB5iE9pranP4aLIKSJGz2GLnULV6/jvK4pK9R0
DvrsbXdnCeTF8GCG2R+3DWtSrCRL1ovYf1F3spb+3PznFqEEUX8pgM3EQMmTC4ZY/Rak3t1kQdpY
K9ntjIZV1wNoVQ6hui+BK7uZd9Rml0fL4XeML2It7O/3K0mo0bam2XXHRrtp+T1Q7T77hGA0gWk+
BRMzYPTx82IBIBmehPD7CMNhoqmcnuEMZRCxc0kCkOqbgsKY9fsOdmQxebBvE6u8B1HMoXtjHhzC
Vu5QkQvw8DJgYAc6MmpyfHa0pXwJsR4eFuf122fDi9VdZ9q98+gf2GU6BAM3aa2LhTQBo0iwN6ru
EbTkjVc5jmmv0Y2waCd2tOUapYqLrUcMPacTJL+5rhTC9hZnHKC8Z400aHiiJ5K3MbqBN89k/OBj
VCakylsQ6Vl+MbpXHCFXNdXXI00R25FrZ1lGIbpEjm3luipUCzALQxe51aaKfieMHphK0S2jQua4
C/ItI21140XEjkQmGe3GUy1Afm92WWpIlaqc9xuJ6JUTwGy/Uy5x4gvmHQaPdluRuulMPIb08nMH
YAA6LdZgrKxpHs5jYw9VmHuXhsn9zVflnuKhyASHIt8qDzraJRCesN38qe68IK80k7MatkHLuHoU
FWBCKHdzRSmilRyx5btNvs8EEXzSJAR6s8A84ZR4tBFn21t2RNd0gNYnA38PWZnduv3raOMtHt7b
D7eXwm4YGIhUnJh5nTwGwej43gjYuThU/m7ZfYwd4GR5EugtKR4D9f3Ku/6qmiA/PwLkLX/+9KON
O3DllKzIvLD1OVCDbT3CmFkb3bjIjC8XNU9BMnD7W7GC8fCg+rHxLMiAQgOKAOKTLyVME7WRGClt
fjPC3HKOUM6egVh20t1HWcu59Bs/EqS3jLOM5wulKhW8R0eSreCT8zfaKXxjSvrzfoPLZrw17D69
ZmBxIASJeIFJ0JGDPzsPIet/MHB+Xd8N0MEK/UeLbaFfIXxxd/eMqhiSbDnS5R8ws9fZYns00Aqb
QhMQ7qTvbvo0riaB3gBcVD/EPx4I9T50OjwWKoa26CMMBv+1qtVN0ytOGAjxECvsioE7SgJTRWMp
EpqE6vcjtGqiG68qWSliCL7dONCNMAoCfUReo63Jry/GZ5t6cQHlDoOIlyOKQRXjdEwUvi/7ypPH
grUp9GVA1mmP0u2I4nu5/QGTTh+NOqdNa2pO7s0Rqbe9BC/Rkti6lMl4ILNX1RBpUy3xMWadEXwX
sEWchI4fqhhXdM3LaxoHkcTk7f4W49YDeJJsVW/iKPAv8BC80aDTrqjU4QYY9aM09nN1ktgtcfDJ
c+cAiQ5qn5gQS1MBz3BMVdnX1yPu/NzCagwYZUQij0uaWI8X4mh629CAq/aFdt1sn3+3l9yOrwQO
oewTDZKs16dgCue6E2NOZC7UC2dJgB39fhhKvv2St3Z18DZyMnSepEMZGMeW0fmUGFLP2FXjo6JC
qdcrv6umG8rhli1naAOYjhmt/JnBAUmdtG+il2WMkWh4Qy6ew3Eg2wk+T4s7YJkNDGkgA+F9GtSr
IY+hBmS3+n7kUUqwwabVGEexvxth4u4Im4cYTk7Hlhg8L95AWE/s/tZXN6xXHlbOlErErQ4e9d+i
NScAFe8J0IKaZjXM/9d9G0DhzceEn9VOOLnUQ06JUykM+TSV7ji09JEi1OWq+g3fSvtAG2mTrIS/
MCZSnokJbU/OkeGFsFDNUbxsb4oCLErKWxgN8c1/O11IXVdyfhuAu4GwCwy/P+oiv5WLsTVA9U1l
NYqaotMHYLO5lIjvfdO/oNZ/jNN7JaWkxubAnpbPlgyD6Mx8CZ51Bl9PCDXmbcZ+TtwsBSc1ho16
tx7nkqg/pcC6ZVikwDe0fLxbiacMaYRdB0/HnFXbqDGOvtZNYyEL8QwvWA+XPPZAu+eReRJeG9oR
Ih5yEt9eEwNw4RdfjebQE1qMSK+pN7YQBzCJveoGvE8V7hq9Oi/cYUP9UXQouST1H/aiKCFRRiB6
O3w3VTInlbjkfkuYWY9CsYV8ZqHUzVaHVzgeQgZ0kpkFwYgJybB3nxO5qpwvfUfUBK6tA/DDdWo2
R119UbUfN3fFmusYB368P2lDaxOJAkP/LgTo3BHqH5YzrY1vHLv2E6CuTSEF04bhmdskI0rQ7z/f
n/KsaNM1rE8RsDq5u2pnfSifVGj4ARuhiJMI/Um3epHELgUirWHsS0fvtSL/xECVnW2uKguwVAMt
Jz9WYLoQief2XlxdQ+XpPeL0Z0CtRQlul/95n0rWNv5jcYx1s1aNg9g5Ps5n2tbrhDDGWMyBmIvo
1Rz60PJK1VQdEp3GAqMpZlOGqnNYhulxEzt4+Ih3WZzbtQm4mMdIugtbnZl7zeO73wQNOUOEdZ9j
56qBAwXNhkOxU6ybw/Q8g79QyvwCGWiSnPUQdS1UYx3rmejqv7/IXPLqRpD5y9PJOc8rQ87lpjMY
E8Bd/a5qWjIPr8xz/6pO/4jAY3OgdivPh+1xct3bCxGUcnVOwOa+28Cm9P42f6UD7AbJRVhYZdBR
Yx5cofv2UtRwtHKb66cRdWLGaKKmttIvRbmsTNvoQZCTbpT4TiomxtMv+pgbu1hw3zmgyFRt+hHo
NVO+AhvnPqGlO/7PvfUYVQ1tggKNT7+hOweFjLPyKfcFM3navESluZAtVonD0t3qTMG8AbuXspsS
axB0H4dGDqLj8uUL+5jrIhRN2Z2csR8tnrPSmT0iI9gsRyi95IpgfJYbP92JmSOAek38rFRdVX00
Pm713Ra8aNS8vJSaJgByI59eyaAGEvLuaK8ZSDrRTwaTr4gcs6U3nvZYcN10q9g16J0T/tL9sl0Z
MZ7RebmWnIeVtzjbw3ACM8jjp4Y6yY09s46b9xfRwp50rw7Tc4eW+I/muCx51aLQB8kU5N5XQFkN
ql/vU8k2l6T0mKLxR+rnCLum0xmQOVDB9FmyAAMPhtHDSh6U1Oz4jAl78YazsEnGmsyJzWbrqeg9
0/f+D5whQNPj9uc3xiGlAiNkWJWZkjn2+hcth4affv1jZWEwwSjdxHbS0HrTSqG2HYiCJzg4XSjb
L0rbNl9ZjLu4NyW0B/sBi2un2CE0sWmTGoP7Qyw5QWIQO2igowIDmsNNi1qCwVlzJfVh5ygrkgr1
BtoFBPlQDTBhpnru75OJSpDVNPf6yq7OsQcxRWTR46BDrLLT64nFimYdWRkENbx7xhi3BSkXIjZM
+7i1/AAm2vYisiDi0ynC9oLWroip2LUcSPeNEsg0BWq/IelFPpBcJbBswiftD6cLapRv+VRRljW7
lWvSBZZ8rfXK6f+ZstJt7LAfFydkqYAYak4SYXB4gwUa4j68mipntOjKCuK1c7caI0kfc8V3V32t
kygrcOUDPFtHmJw85mmDxHYsmYKu/yQ6+Vk4fAgYY9oXJsCXlvn/KtE9SHntBV0AmvNfJqq/CCmM
HF0MV7OurBnYO1cdgx4U3qE+UlJROihkARKL9PI3oT/XYEo2AMeX1mq0ONV1pA756DCK9o/8n4lv
I0TiLt3Q0P+4t6m646FMMFD8hs0M3oR++IL+2IKbHP0bfMayxvg2X+TxyzMonVmnmcBoKkcRo4pp
cXPiOuAGABuYBNZKZoQnZrP9Cd06zxvq9j/KQDnhnAr8qMVA3GZq1ooJcdYuDhX7nqdfsWYVECxk
tvzkcjrwK8Ucg16xsKiJbVgBRZyPxXtaAq73VDDDFHbsI4TH97j+KdP6l0e9awI8f/kEm9yRkG+0
vazE3pGWHfFFo7JBJzUDvkanrTzxgccaLnSIk80yRNouGE9ZX9xCSkQlL8SJ1XKnhx/3a/HJi8ee
00WtRuvgmseu13M3QBbsM4qrYVD4T7du3zo/WDlZLyaR0Rh5qomXGldc4EXryY1mnUT4u/M4+dMY
nGVUADGeD17Kx1JDoQJLyj/gVHOtIoFV7XQGbDK7v5HHKOsSgL22Qv1P6CTEumGtA9PM5kEp+OoT
FsGlLNRcgTn3+tjKFzvEiv5U9TsrAuX50Cyuspni8saiP3lpt1oeSasavcbLtbQjtvNNHZl4pqw4
cCmQ9B+vdxOEYq+DesrNaDG189R8zSgDeqCVyD5Ez5+nVb/hiELHxUCVq2CWa5uVtNqHeIaxbbD2
IzFEI7a4+QdkF6jWmn/BIebD9fqQiDF5K5ymLLiMuxITs2DPuzP/PlNVTHbD/E2pgFHuv6Ee9FQe
bnpwZbICZ9aRqdoz7s6SGL0uyg3Oojut1btXtoDJ83m/OPDjvNi1w7gbdbZRpXdVZjCs3PxGn/lp
3RhZ8zYcPP8hfLmF2xB53kVv8tzMB3S3Sf4UsF11ybPV3a3Nc90yDoiWP2Zh+7GwYfOayZHhxVtf
wyjk+kxnTkXEifpohUl08AGBJtpvGdP4gGGcbFb8N7iFfeEypmT9froKiI9RCrlhXfyESvhaNZhP
UBeLoJfik2i0jh1l7ib3e2HEntWEk/6DMzIEkG63CA3AZDhVNEPhvhMg9JUinZKZMUJ04eDIZRDD
cVAU2i3loCOB2TVt1QTMabniBZACKdFlV6Fe2bz7C/6fCrmoU4MaZL3Rdqrvt1wGH0sXsv+p7MZO
660ZcNnc+F+x7WXW9ZaaFO64EsEnEvalCFdYJ8TJjJanW/JAhpsY+H17UKO+hgAOANAVFomufbem
l3BhsGRpEPeclZ5YX1YVyfUUXtf4mrt8tKEO3r3PGvtF8i38lluIlPNzwSafXqwdUe6XCcEB7QZH
nn4NCH1c5Xd3xSOXJUyO4e1HlGFIzjAzy9GkUJ5Z3McZfQ90LLgHYZkE3Td+VCbrx2geANXLEDKU
s08Za/K+TMihCVd7J+fBOGpm1eV94qOShA7Mv5ZO1FNXTEFc5DZtdmw0az3woGVUEEohGE0oxsx7
u2OAQ5PmycgtwSkic6rDG9QDk7rn5adUwdSwEpDYd87IvHFbQEYGNcm9zK4DE/1K74bwwsvWhCjd
Arb3o0YZZN96YXs0Ui4e+l7VETy2n8hCzcpfx6VRThYo0mEj8C2sQ4+7qy05nwaMHb3loPKTJlh4
/a2oVeawl+eG+bhzwsGAkduAQJY/twM52S7707YVfcKSccRPULBE3/5jDivQoaBYPRY4+XGQZVEZ
a4Gdo8IXOCuqJfedtSYPTlgJcAuslGv18OsjPoOmoSpFjv1qXg9Wz3/P7Cz0eGcz9jVaoPsri0B3
y2v2QS0twclg+gT0YAHMnxtJwDV8Ty4upDCh6cKvcS/Kxx/eBPqNBKnI7yiT8db+k0EUuFzzFRo4
1ixyiQI16kFQ5743E8kSUQ3apiY4a9nvgx8thbLoMWJk1VdjUydBvfNnv6Qr2pzHsR7u+4jgpxiF
Rjqoxc+Dek3fmL17puOlB08MqgoqV6ACP/wOElnNwLmFtRRtEIk4IlI57An2NTrPLybr9tFBUamR
qjpj/9qJiPVINE11OV7r7EkoT++Bj6fT4D9ZgMSA3u00ShzsawJHpRG42P8MbzndA8EP5Op6Stu0
kyaDIIC+9K1zJdUsQZNvuHXWQlV9x0QuEyFRhP13te7QO12SYRRkisxbl73e51RCyVXbbiA45vcL
xapgqXyFG2KVGPhciAHIKX2bicO+jyojiUbMP7n9uFne67ET1mzKhZzEMQGlnUOT0hm+RR6p7UhO
GVrWRxgSX8wgr38NhWAzdmwLf+EMioc6ttvQZymfq5RHWTvz9QIJdZZ4n5hXDj1+YhCvqPZjMJ6k
cBNqJKzhmE/Qu7vclqNSyAhiGwj+nPs0p98ohNyCtwJAVlz/TiJFh8cRw6mEbxKaW3WMEy3UnzKW
eTcsYrVsN5UQzf/hWWxWDfU8+ajU7WUT0oW7pVot7qjYfYxwzEimyco8rEbYVmnpyjlH9lGDVjtN
bgzquCjbKJqY3bAY2ADouYlb5OiZCjmR1HhS9xFBjCg9nibFWH6qFBWX/4VF2NxDHjCGQBJahLs+
Bj7dgAPaFBD/h+NUKMeGF6RvNKW+IAkTvrmotOWdNFzchbCC0vNnGCV84RJ9oBTWOTf9WwGQ9ZUg
Xr/iKwJHlI72vBY8MHVYxDsMQ/lYjEVmkk1/ruZhPA3OL/Sc4zX10XgwKjLFzUu68EA0FSbKVtPk
66ZN1V6Wz0ZJIHyJ9iIBqHFijl+ukkGyE8dv3JRxf0oMge5c9BzYAsg0EUBxZXzDhTPAVbwhVvUS
6d6pu00eLW5QUGqsIJuHe1nNwYb2RMqTGbKXBJd7BT5bk9NKw0GxWCx+fg32YrQAy1FDrpYeo5Ja
MYVa+smgMzlR1gq2PgdvG+FIWx+fSaAe2//++u8wVilSemrz9nyJicQ51G14hjRFXkSfRxvySLE5
5u/KIXC2lTXMIdo3rSbzzS3yuAF3xdbqaONMk/zK3aiuWAZw94hFrEZA6P55fsyl/cw+Y/wKr/+4
8oeNotSGX8zsB5u/Lj6yqxwM8J92jvE53BTzhlvrhPr9+dW3yUQf/+Kt4bBr/Wq+224c7Yw9Tu++
AvlVTsyaJkLROnt0ag+0Si7FkO8KLn4CADSynABPgdIwYfxTJYootHwlvq5lZUN93H42a4EmxiWX
tcSIc65MXUoE4HbdfzRcHVD+yxcIQrwzYFiEtxtukSi3EVXh/L5m0AgGFhM3ipQIpvtVHcJfrRSg
bgBn+ZOlwQMATBjplyy7muI3H2GWTfzLpBKUWzTzrdi69zHgw2OKV6ctgY+6awSmNwv7dcMAmH4k
VrgGRPrYGAxKQLHoiHcF0MLisIKUSezkQRtSuZMdAHABGvPjI0EHjrtomu2TgBuZE0STDuxw0GE4
dpVfbqK6v3xffCQQ9o5ZntEDFGuSEt5VjQ8EBB/swmcxjfE8+p7OVc1kXn53MehlZwr+Sy7GgOQh
jtN0vXg2+SSjWwp6yvSUrmy6kcUXVJ2o3eQnSTnLHqSg9fcpWbgURKQfJmIxFR1amPY+tpQgphsH
HEoD1LQCOyKrEtyJJivP0ThqCrC8XLhqjCOuvCcL2F/+NEft5qP2fId6Eucvt6wdv51rbA4L8nFo
//M00SwdEvWDI7mUG9KcasyrJgCHbeCE3lGWS3gazGNAlEgjdLEBWGJFmfKj+FqQeTaR5jUuctyw
fTZ6sn0ovTeRN3mEI8PaKtAxKcIWu+8IYKIoHT5GjG7O3il1RtTlfLWEjBoZErPzs6/hzq1Ezmxa
sVEU7rMzKF8RVem5wPtZI8ghV4mMyX95dDKTAF6N9LR8ov6ql26vUjwY6i1ALW8qKhfGDHdpYoHb
xpq7LTvCBDdpCNbM70QSC1y2/w0GJVVRpGO0QSGvzsrQjZsNYTTe5Ehpp4nlBlhlZyhbsNF1pfad
oLqvaZ4ASob/Atbmlg8zZDkrW1jXTSZxWcuWiPRIv+H5zuEbXmi4lJIcljcwVtcTbheNtSP0UcuS
8deoYgmqFj7h0ay1QMpWlUv98ZWE+puDVNCeI2YtdkEgQkG7IE9t8DNF9Ls2AVWXF/g6SE3xMnNk
GT9SdQ62SgIBI/viIF6+kb9vzOELRDxAS/B5hthJa61grAeT1AZw4x5xPRP/RA9vOf/gnOeaZz9F
lsc3OdF2NFgASO1zbAOdIv9Cbyz9neifp2k5xgrw8oF73F6J/85aeioG7F4HChfgWkamke6X1ok1
csMUspkagN8RzMftP3QbihwFVZdEBk/RCmh5YZuR3cQegwlIzMjldrB04kV9GcuxmbX+FYn2ddZ5
eEmnodlSiD7ZZZvMHVOMN7Jm4HSJWQFXJxnr+LVIYZrAemPZXSIG7oiIE2BHBx/c5ywLHK/zTOwd
7YMJ2rlaVnEUnP4rGxlMUXaFCGi4VfJgWJRNmnRfbDi/GPfx1qp9eu5LMxJIdho5PpWIEArjV8K7
ccISIWMEw5NdXd4Nbqs8nUOJy1aALixme4LBVJeZi9QZ/8Wgb+XfCVqL/tmBgEN78a+f+UMpFX8R
YcAWyMmjxNaCpzb1Z13Ql4nABrGJvtDGONZ6KUWa/2713mufLL4VjWxsWGBleFC7HA46foWy00DH
1A4txfTGaG69+OWgC7X/UiRAExC8SN3GI+ODQ131XQzIJPC7kgT2pV51dEBe1rMvOizFQcAEf8ih
ptEjPPjM1odwCbl005e4M4zL5wwll+GCIDKVMh3jV08p42iLT8kITA0V3eLEElmhFYDY6ZV95+2t
6gdSbh9+rqM0YjMW0c5l4tTiC3xy8ZwoZJukfvuSeNe7hqqEQFz+n8XrvfqtkIcdTfl9Ub05Nb6T
XYyei0xYV/F+e252BgiU+KNfuk3GrUrOuegLevbC3WXXS7klQ5Lxfc+xa+Id8xyeZEvEprmW04+M
5R4ivM2us6urP+L2mK3IAaHI80pqxKvOlsZFvWKaSGBOmZeLjqnsOQhBV0rWeMjZqDJfZWoWnHYE
LSa/VXeMHcjEjeLf65UMIwK4SU7RPDdkFeBvIVMM4ZBXSP12FcCBftjWRf9SjpMMKd0EyuHeCUU9
RRKQWNpRT3avbYBeEqJcd4ZJRFb5zWEKl675BNY7wHVTa7ieI9RkPf2nuU7X45q7p0gBfHsGrKU8
oxtX6R2flXjvXg3Qjjmm1w+ffYYt9OlV6gcKJacpUeyQs+7MEH8ejAFSoEcXJ7xz9DJosTVnBHW/
IAw6KB1TSyomSPJ+g7DqNXCb35PEH7v8LailHvNZO8gGS5g/j5MzakZzTuh+uVyFrOJjx1HCQ86O
eeYLo27k/vrP5lRyVtfBeBrKlEIWxO7tnhWkoqQRy8s7wuB2Etjm7Oi8XXmGRQxDOkpPwOyCGN7/
mo8nkttS+B04w5fDNXoTzf9BIthVKHp7++LPkm0bysJY1oJ9xysAM9pMgabic3Y3MSrpZg0hX5Hd
wqiOEwbYySmqojhbQGM6YxKJSuqjYj8l/ruC6+BSVRmbQ5vSkq7eBqIX+oaLFXzWOKZg3Wd63cLA
rRhZkPZ80DzReVwXQnrBH+GLFiFHGIExfcTQV18yu+pXl0EYWjk1dbDp154nagt0aJwkC9rQuSqA
aIAp44rqSAQNF7ydw6yPxbPhr3e39T2syIAsVb5XjTm9ZxXEQu6rWouk7J7Db9Pw1wqjSydIWn/s
g1eE7Aw2YmLZS6l7xD2+7RXCnjI5py1VXcH1FD3+j5YiHQhfQtbnnkogC5/p7btLQQuWF1oQJqEx
XBchvvTg4g4lgS+fS4BOuIeBwNVAIFMrSNeismnwyiSWud1/hMIXKTyHdtzTnt0tN/CxFMBhpd7I
EtX7XIkYEezzyk+uQFfqa+kA5GonCqBYRtZLxyhXpR76IqqGxC2koZeBSMF18T20q/LFEStkwLEk
rUsSE9fKe2UWVuoWQRxtIcHP7tNbJLUDaA1yEP0W5VVAmcATcqxdeNyOGUBBcCSzCUblYuHUNeFK
kCEUJ+66jneoGP3kE9+/OpYDlriPWT8d6xr/cNt0yQvcdz4keCDyIpPW6SZhrxhPFfTh/AiUwqCF
NLbSfZ781OymDc2NomOQBysH7Yzt8ytSVvTJHxMH6RTj4ONRMKEhxggl8XNuAHBgAdLsLWBr+ofT
QG6PwXbQ8VxDhLHingnXgK3obbZritn6Gt60vDM/b7RCyQ82k4NuVXeAIuoMQqQbUIiCy91Zgua6
MV/wjgTpW6W5NsDIJGp2vZne+XEua+p8+EC+GKDlyc3lcr2NCQbPF32Sfsk/npFRWASAgx1zWy21
plijRLqicDS/oaVYjNzkZFidWzO9UmRGWLzVowLncTQfGtZ0Okr1ZRBba2SF792JcWVHMAP2MCWT
UEfLrWIIhlOHiNHrY5Ge0VsgzRqueleoD947EBHBJP8gyx3Kr1H7/Rk+jnqsWNNmZcDTc45FupTH
fnBevrNqSKWGViHaexz2EF3Qq57h3nk/H0hdZ8Z+L8cp73YLl37DJPXkIDcSjdG7qlt+WLpZNygd
8kC/O9X8UJdjKwZ7S+PaPyPfrYm4k8wrbohEOnoxEpiCWJG9mk4sVcGMo3tfGuDW8vl22BPpqxBI
PERA8ZnFTFfGyW+STPToHctIpTb30bREfoRtarUtpmToLW0qZwnsStKCKsxjQJ/qRxflldOlhBCu
KChQ6fJnH481SfeWpX9+iySN3SJWIxPSzSah6DajV0mPuKiJuANWBbjDkaoXgdL8tkOrhs2/gOTO
G19MvMgfVrQSt5WBMM2J5FljQHwf8d/ZxyCKkdczJd+rCCrRp/41yjk/znuEwKvKVmDbsCrUCL+m
Vif2+5JlbDGm+F/q5WD0Drse89eJrgKP8cSFLowQrzLiQRT89ILY9LlcM447qpIT3wGW1kT1pOmh
rNehaUGgXlyUzy1dwz2ItURy+lx/1hW+dlehRie54cy5muZXhXdvtsn0lIIX3wbVCndrRJtVIfxH
zh/Zv0OAqM9Lm5wIX3NEHreH/6qYruEo3m9PgXvJrxsqWEiGpUZgoIjiIKplFipIKtfj0qyTITOC
5TC6rvbWwXXsMJb1De+ngoUqbVA/NlPEc254gPhVK2ca2xa9fbVQQ4Wljx/m3/VDH1rP7PzosEue
0YOVvJ7cztUgb5lGF0QrmnhY3cwHC3QPk6lKFlQ/j9SaUsdy2YHzq+YIOzLspf226bDmoocxfurF
Sf55dq2/q0Lv+SdvKvPMBBhC0yiLw5easRZRXIeRoxohKNORaGvRR1AzYQta8dErqk7aZ73TQQiJ
ggS6yONGypXdiZE+S0sZngSMg5xkzGbaQK+y2tpkl5yuWQ4jSok4EKkQ/5Kj9SVGOikRdZrVf1MN
xZOf0ytwqG34bK6IrKiZrFWI0xnoR4OdAcKZMETYSorQOEmLQ/XbGI+AlEw6FAzTCJG4fMbSN4CU
5wTqTp9j9X7FmRJ+MWK2tDn01GTYJmr3x2M1ojJEVRtTV4mtLKCqT1DJuz63N4hAwaUh+s81kwM8
XRNb5SIICi6VNs1eyaZ65Qz4GmICqToHcSY1moPwbezGZl5Qz26HXSg5co3QsfmkgDV4XS3lpLws
znnOCK0n7b+2HgB/ET+dFRHP/qyCll0Fsf1xGxMYIZH0ERweCTBlx3I4tikn+zmVj3xclJGbNOeX
b4frh6pZsVmHJ36LPCspYmohz5ClmQi18IVYOibrove8vrjg5QVNSVbZbko9473CTWbQQ/Wb4gmf
L0igf365x65VNWEmxTVlajuD1u80n2mlV7Xaazyfzuc1VHfVq245Or6bwhLUP8WtXJivu7YEYacx
Vlhd10rUkEENRE0BncPK6aANNs0LSuPwd7oyXjx0v4Cq5r0BSBEtPWNIwDNAjPJRNdFqryIWehri
F29qzZR5GVO4kC8u7gJ5WdAApe5/01Mbf5EsKOkHWN0dmIbSQafuesRl3XqYGPmD4DMVZdP4Av3o
lHya3sM+9NVux0epnlZb49e8PFBsd9GNkTgPTd+moTmG8HAjcwPxrq5ltjV/vX71bTPKyhYg5i9h
g31En2aC0H4SrVNabGTLv6UUWWFVw16DMsJFcVEE0txWyWfv92Dqt6OaDurJY6OmVXHCuorp0BvQ
AK1AHY+G2WzIXXD/W8AjayA8unt8T94mg06QG05ml28z99yUVRmLNLfoLG1EvkhqBN5NyCCnDITj
NJaFEn61BTDGzVPJf3RVXhTajOF+uM8PK9as2GahOBzXARwo9Pz6oKAb4IfoRfQlJbq3/hqeLnf7
tW+5+q37Rs9Tpt4oedEC/9tDhcXvNhongx5mE+T9EgGKyvy0XndGMRONZVRsGAKtUgcbzvZyrXOV
dV0OcP/qDwdHR8wILEaRN7Aphil3s4t0qfoI46KyLlswVwVW066PQ8qXke0sjcHKpbV9zyChA/Cp
n3fXcQ8c9K9UdgcdAHZHzazE54W3x7yWfutggLyBjPPeo3QSy/XijIkArOM8Sfc5icaxGYZvBGah
ouWdCNbBtreUW2WImTMXjA+/AVAZ6sX/oCBc1AYsudwkzW6nCIeQRuusAEvVatG4KLvBdvYkZ7Fe
Ba2ujvL0APdY4XzRT9tfHQDKDlIHfeLm92T5zzE9x8ensi1IVBWTg1QNPSD6hJLT08qvmARYH3y/
MbE1jg1V30U5PdUCJHKJrnwyOM6Wp+/Fpvgd64hcne3e2i+NDIAzcUTv7/js9+z7+ECJ5nIF4KDN
o27s/l6q/nyoBgnTK7EuykmgGOBHLQuaV9XcHEnjryHCRyym47S8V4POv1AU+IG/zlF8AxvLtNya
SpvxLjQ6ZnaI0LzClSANWGys2lib3pDhrmxfglGY86ZDip2wPRLniDc5JrscZuQt5nzhKqRQU3Vh
eLyz12RWyxMVekUD5c846AtDzo083KEruBGX4+4ZCi93YTNDBhhqxku1d686kyAh1zs0ab+OK+/m
Osig/eET+9PiBwHpX/KqZy9Uegi1TshKETWweQAnbI74ZeDOCRVd//dWDgBd5tdKMmtlWyYnRWiR
hnW366f/sXwj25vo5IeSQNQMFzPQLCUW4SCy659lTjHvMGsu9ME4NkwXXF9q/Dh/9QWaifiu1joW
XtJEjfzitq2KfFwsEzpnzSbgzmhbEXBUYccsFZTiKf9n4qkVCkE/+JafKD3rujLraBi4AKfwevAp
WDt2n4hUDu35JyVK1auJB1aXy3B3KYD4015i/7loUPF9ATNktQqQ60DsdH8qztxKNUJkSBgy/sxp
QowaCOKEgtrRturZuFnEiZtpW4ywAgBm7wYoA2ICM+Qc2IG7FEohkYZRUYvLhYdPf98AHockcBR7
E/DxM+IuvzvvecpKtz1d3HtJcEzLkWeAdiQntJtlhNd/XUJCirYPuA+6g7qTyWiJHhbR60wCu4O5
FLvlHIkfonIlsxpnXC34DDvP3WrCNOwgk6LukE45vVLsjE1DHvZR+bBhQ2wnHS1FNOfm3s68I/PN
FmFjX6zS93TCgXX5yRyqSA2dyqbmqtZxuxw4u0GZqe2aNbPL0/c50AjWa2an9z+V+2leqJ6hcjjN
M89sTLUpd69SelcZHCTfXEiQ6ntv45fPrkFylfwcJaIdO2zQlCisXbktGwUc8o40UYm9dmu48h3H
FL3XLYeDwgBSF3XtUm4tdG72wryDM+26U0OPnpnPOM5us/g/gTO+mycYIZFKkIBP+Y0ciV2AmIqQ
HNYwRKrk8CVfRj8rab7zGVjSosIhEleYyPB82w2KQNk0/QKIc56v+oxrhdHWIWBVC8Kw2NC1lJW/
3nLbWoOmF8YZunZP8OL2kYwN5HQ2aR+yyoPjIxvTqKL56Mrfw3yghD+w96de3PfVrVfOTPLUzVgv
3q0v6BoURcYFokTlOi5o3ixXSqFagJymFR1hgy1nZ/zAbi5Rim3eElA1JMTHisP08HEZL0lcM5HL
bEe3cuwBaahYVz0G3kh5SY4/Gorr3IRokxSdtk/Iyr8i8JSXI2t394qR/Bt7qGTI/bcNvtq1C7Ih
iclbeqSYMnQcsUiJ3QPyZRmbxlulV9QMDfc+p5NwfGwHJkblcv6XLU0S2vTy2k+Sc0UVhFNwEWgo
c1wi8Fl0c6bskvRgx2wGFCE+sVye2uW2llrzgXbdFgThyMNUa3vk98d5vUEjUYzenQaqgjNsO56c
SH5ff6kmCTcxaK/ENUAV28q58TtPSn6pJOotEmyhn4PGUeqs3jmJAcMm5NAPcEZVyBC4p+9LSLLs
w+69MAcNJRLFSci2hBS5SvThfKUC6NQKhyjh9fvmMX+G7qo4dIV0dovNq7SW0UGYVrtzJgM/5bji
3dnJpmWvq8VTpi7CqnKbkmEq6KhUHnaBZLjlaZ7j55fvfY+kkhlkeEUmVU2vvqyfOHiYmYhApU5O
m1zopPOBmyu4DNoLvny8WCbJHKMUV64GDDiLHDUaC/SVxWQTFs7rJZpcSBms72nMIJ22RmUjN5ji
S+Dn6yqyjMBn3gVTt1qdl1Hl0p9ONHhT+CMP/7sQr+HQDp8D3HU/1dcs8X/WmQfs0/WYARjBj07E
vM6ownkOwSE2YIctQFWATo4FjbuwgGmYewx15H4GcSSoSSOk4lkvT8RUKr4s9Vwxkr+KFu9RnzGo
RXDhydl4MLB1ij/XefFa9bRyN4ZEZMUOwnTc9DssL+HK3Q3+43Dl+hY/G8up7fb5vIXbO2PAwsoQ
2UHAulmsiYRjFDmJuSxx4CZ8lcFRtDvS/axCS5lruHwHMJtTjYTz+ITUtzmQJE19Mr5dnIOyGoTP
fUvZ6khYyf5zIdcAlIyQQUJLm083cO8nFYkuoemN643XbsBkjVTKA2u6umhULhh3UTnZIyX/Q3hm
r9js4yycGzFqHf1aJCPBMVrVX3qwPN+lujA8tBE8ByozZM9/Wn5ujNOPq9PadHPOl610rkTiKFSr
GkgzwDyApulbD/uRttIdOzwh/A38HUCgEVIcMyW2xPiIWidar95V+hNre6PdyvGzMD/Kjt/+dmqu
vK/r+yELftuQVw/+S8AOGC3WcfpXBG5ThWzfOzcfPZ1/0WrfpbpLlyiWh1UQs/PEzDOwB+RXvy85
3Hy0g1GE1a8yLbEBDm8ahT2xAEx006vx2Enz4UwV73m4Tbti5proa0OXCX161dHYvyiQyi+N5R0W
dcymQmKasWK1vU0LcMMcWhfZLJfjpgABw7myT8ovF9w6/PNE+a2J2MVW47kGp4eZvA9QxW2htvFU
St8HQzd0vnFHzKf4rMpvcxb8qReTHJIXFzUzRU/LWaSq6PjoqEqDlHQTCysAxYkWnjV9CZB1fzg2
2eC9jtKZrQmaAhfHjS89E4yjGf3CaM3pkDuvknJ6EZJs/10xJBZxGTsgFWqOszqLOr1p5mXIi2us
lvsiL8JEmWsNSRVjFt3hnWsdx9HmUYVlRMUqjuDTgFZP0vceGVtrFxnwr8K3+EWM7XFJEiORRKkr
Eo3ECXxlxB0Z1c/2f1b0pQU/llIBASdhY5FbbOpb0eoxpv90YViLSc2FKRbOKVX5w1hBrcQjrwHC
OvAvVWW50GK4OJsT4Mx01IakV9Oi5z6aQ3MmflJMjMBB4glYmQmtHp6892x6ynkNuhCjKC6LqNFM
h3tRyR1ZC8TIgmTzO1UPdLjzlvdEHQd33k6uRFJB1nAZlNgnaVfLt0UBLAlmGodu1HSRJHiXz6fb
eK37KwgbKbcCwwjiYlXVIPLaq6jnXToLHIUClnzr+YRrjbLwcdHo9WQLmk4YKm6pSk2NaYTM/IWs
z7gx5n3EU0j5bLGb8Uip4xTvb7GnKDXbVtpYmH3B1DmgY+7HlugYuZE/w0hOM/MlpgvX+DVGsAAi
MxL1WMsmXtpkXm714UkxL1XfCXylHKl5Ba6Y0aN9LgS1SjtTRte6j+YTdemsoBSeKJdPvea7CKuy
Km8UCVnR2rHhJeOir316InJDb5eBV3gDzOQLUgZNSlpfJJT3xfV3M72W07/hy9061KDBsclIzh9h
shn3TFfV1tzUwoxPp21ZLWunXOGCCBibPnqw/60iDlHpdsiMIpdRlBUjfKvrUaECtP15TXhRDsaG
7paSYfn/rOBKSvTUtEW94T1PIJk/Y3EDXpR18Rac0Ir3CmZyLlFqprzPFa4WocIr1NG38sncrtLB
rJ4LZePz6e6H1BKQo9gClpOOHKDMYSH0IS2TXAwOwnRplVV25Of1wBYDr1Tl32XWQbsGSFPH7ddO
eNopsltjiIV7qWPGdSFOE/zkC4nA+wxTqLm/Pu3dYRutQEcCqr170zVxWL7sSw+VKW0zCm6TiDDd
HENTDiiTXOS+IzJihq9h8dC207wiN3C9hKIgwfSyukd2wUCJtaf7V0TmzHaqpCZUsb+mbPKQN10P
SuGC8teK8rGZJc98q5IXKf2bZNKhkJvFXXiUNJFPbg8yxOuHdd1TL3FmVv9Y0jUocJPnDMt7KoQq
VuqvWEVKnVlwE0Ge1TdErl2GxiXXUIRuTOQPuyGVFeZEz3MBCrpJCXmV903o7bYPGvinH620HEo/
DJaqGYXmD3JVokjK3oM1UuFOOWk9jq8B1FLf/MsuT/naAvHTQokToeli59CAn/Ii/tZbiiG3BtSW
/aOYwTqUg+z/veY8G4PJ/3PS/VjWXlF45eSxffgjWekKH0lF0w866sSZH0o0+d6lRCPPK5zKhmog
cDvefY5fDAHb7T5s30WluVRlytPrVtheYEGG3JTNsRyL3Y6Ur+bviqfRk5fH2aC2HC70SEfh4blV
hmRGlZynnCAeablsQ6i6PjUWzh9X7m5BGbNfAY3uO1/zx5yMjAYk9YsaDBgtg4qMcPZO6hJxkKZI
l7J2s/LH1RN2vLQO1rb3el4rXWaZkUY8eIAmnQiSFZoWchR3gtsJHecmp3sdR7laXuAOSvG4vWmN
UjiHABox6uqXWGvTbzUBDRu+F2sEnNHOXZlvEJVE1orgy6NrlqzloHgmO6bFzLrIlDiK893poBXF
1ZZd/IeAVdxor1YONiUWVaqFv0r38qsncHYRt0gzdAedfjTg20TGCb4P3KpzuUQAlxzvF6scl3zS
25Ht1Zq6o0l0WftWTDQ+pOeBIdNL6/pg7ECozrBhbQ4saODPPtVYRtF/34vmHSwXcSS2zenFYUbh
XklxEYPn94xbUWViP+hOdZQkic+htUcsOfwmD/WyO34rLmn/W1FIcQATe+iWZ78hh2lHTi+MnVqZ
+DlbLD2QPg+YyoPI4B7KinDa4CWYRhfkvuIcVJ9sJH9iup57KcbwiqXDazgNhNz7hmjQImu+7nvq
bpZg2rl9PKJDFxExaNI9RHTu9jZnbmqGmmcMhwy1IXz+GrJcaOCGrW2jDzgAcHp9Z/6pcBYl3pd4
k6J6HhYuLOboeACV46BItucewglk9Gl9N3MA2uvADSPBtborFczx03acUxS+w+QF2cNTJgh/J2Z/
tv+SoOpAw60hvvbjNgrxY3hjykfUXto8KsZ0v8DdBrpS16v43Rb3bWYRlprrhXM/YJj5RZ2fo67+
iGCScQ6qfuvfKDNKjWvevp/aTy1lD6o0vkEjiW1/11mtQa4GuE43KFO5p2tjqCdTFghCz1GLhZEu
TSZk9QdMdZ5C0mxAp5p1NNgdbqfAArA9YrzDrGKdQVj/rK52kIV8EtI9/05UtPG7CmBZstsedXUt
htUEBqVGD82ZSCsjf5pS49wRpmHGLjWPGwe3TbWFN6IKFvJzjopbfBX7i5OzXnKqGT3YAb+08WB1
Urpl7Toy1y1Emz+oItEuA2EFS95N+KpMytEp7bmJQGH3QtK1raL7oJeqi1J3ciwOTCpNbUUiFm8F
3MrzWrFNj44c6Qx0o9v3d4C0VbfMsqVIQcugRmaQKR7lnlHoHfLBR7qi/04UPd8TTPG2NBtF5OCg
IUSPQMpVsZPetyXpUWmOKviKYAWbKyCuL/SQcMq7nrnNTXVlyB9qSUNxS4Tyesuo1jf6evx9cIEO
W8Ir+oDRuJ2YQ+QMBpZuStT/8q1ptiyGnotpQXhhSgRgs2BF8uh2KsBcdVDleJaggHcp1c5EEdwl
/raEr0pSgBv4zvP4uARruVCim6mV1fmnt7R9Cuq3TbjRBYXqIhe5+C1liCTjZKy9vU12kXEe+u9v
JK+rkqtZaita4eEiHUri4gLrIHf/inT48vRYknzOkL5FOY0x1qHvP89Y/wIRAs1JoClF4T5XZtVw
9xZ9ZPgs8xcKVl4Eqk+0o5ao36qsh4gxpFsFKz51qfxTVLSIQ1WpC3iV56zR3X0cbxM9yyqPfUlC
mpGtOFOcXHMiYYG1ILIL2UYRsQbR5dMWtNt52gFg5WveccOo5PrU9Zqu10lmt6E0aCwDgxkOhF1n
IV+4t9189fckEQmyccGv0Y9o9OjH/QW06pK8ee4PqZqO/BO0XlUSinVZlNwnY4lrC56KMZrF7iTg
rtM3DAcSUlYNw6SvLCru599T9W02k6PkSEwlbFpBoFP6g2YQcAOGRAgL/0L+aWA+kFxN5O8aPT9D
+AX142Xm0qForEf+W9zs9XZRK37CCxSTvaXSWkKavuM+FX4rid/UbHg5lq8QXHGyhwAIYdOX0all
Uz+Yf8Ik+EBEpTgqi47E9Yu2KXPdpIoBuWPat2tQQadGnkGp+msrcHplgSACgE4DWVrI65nZ7d3Z
FxIUUaWnTCAncczrUPuMXBkumqixiLBIs2OeUmwtBZA42s/eCZr6/N8jNGo1SjRiUKsmfafvU6ps
N6xV6XEBDRjw1UVRztcsNAhDYEXsBpAwkwgZn0jEobFym3/Ky9NxcYgzokNz++l61TeV8KjR9wDh
C3+HI9xOi2FrJFVA85nVAoGS/bqp4y5CskFWGxqXrd8l4VmkVuRf3S84ZiYUL0su0SEUv9NbWh91
bEpXT9swJLhUwmYiQgiQPJV2bjuDP6KxWAMn7m0O5Pde3+8ReCcmWcSEjgUydjwiv/m61cgbhr3N
Vg75sdcCaIBpPniWd0C3xk0hiCFEcX+GZL1MyYUuws8VjbDSNW6SSHv4joKh1X6QD4D/1Dr+87Y2
qF3y+krFcnbhBpY+m5W1RSDIyS5tLpt2Fs8cGB8brCyuU21NOhppidLaFRkHKPl5zAYlGuxRAAgi
jOKjahK1z9Vm7yuValTMYVGhsXlrLRGeSKDQ0MpIUb2w9gJRYO/8aAEpss/r76Qk/1r5PwBoPRha
/kiWOG2A1+LS6zv9118jsdJzQUQipaAlbuThDzhRYLeWvZ6m452pjKtJJ49Q4DF2Msqe9nc0tiSF
nRS0WlcEWEQlKBftcWH6+MGTZgXlYQLW85oD7N+Oj5bRW0e6PygzP08BRQmFr5z26wvCtgm3CAFO
4OodpOdDgFJuasBjYG76ozkh6lXqVjWzcKfBdVypYomogVEXMTNi+n00RSNnRzA3Jr99kuJ7m8s9
B1POyZFYTwgS9Tl7jAdoVt6lZnVr7FFiADpLV24Gj+3hHWItgRuJnsqqetuMnthtHYvJVaB2hS0k
MM6ZAltfuK/F5Mtv4e5F8OBYXNUuIQuVM09RXz2xdtLTtfpWHcuW92D/DjLbh92qbMe4VtrKQvkQ
mVl7EOIxJSeLHIzIYNiLZoKjpyqncY9IJj1RFu5b7/frvcKs4Qw8GE5Wbjz/faeysWSQA6f/rw6l
bSSLrYD7/UN8kFq4mrtsmOebK8jCL4Oeg/RrMbewgTYZp2Gv1UAKT1bZnEMk0OypWDJBiTBOUPYu
aXxhBYxORtxdwVS10H+gzRMYf2Sy50PqE9QFndUGeeL9p1SKtc2g2sS3fQCJQfl/mXklTb9HRsL2
sgXYmghBbD9LseSu5KG3mYiKArELIKiIWfes8uXcB3D2UHPP0Hw0B47m5Zd6Ky04QwA7vA8LjGij
dr48TKBN7+1KMyA+Ddlrlk1uuSsbZm06VbiE9sVfJXsz0Kg89EQDwdQWn+e2NV/C4zrj84DSe8vh
zZGuhpJBv38qohPWC/lm8V0I6FO20OjtXHcTkI5fAKq6Si4UX2x1ChnMAw+EL40+ubwkRAXUGQZS
aMnY0u1uAPI+0YpF+OwCtwvAt/nmy4iD9hF5L61CAb8xuvZ2Wlpc+Psz5gorEa+WsDYREN3V3xmh
bFgUxWwpukBaoXTfIW//gvSaRg5kq23YUkaEupa5naVPMvUmxEK3ZAWdPaQ4Ci6c+CtY6M7mSRFC
5eh3XerIQCZhf+1Mc3Z9BHfC9AsikJUwM1KD+ueIkXF3BTolrv4wim+W8Ht+XvuO7C5TP7WMm2Cv
/w61clyDX25W79xnu5+KdPqr+GJBkXODiFToBlg6z+fA+5+tX6sjZRsM+2ygfdMOLTrHFeQ/MPmq
9+GGm65Ux4Jo7BlKUtnHdobiQLzeRIYgpeLbAeP0j03JPQz8VUhTtdBlewfUHOyEU++VxliJF1yn
YMjA0MFBz2+/1vTKFDhmmlmpvzX3ICwXZ7Q5gYvJ0EsF07+zjN9rcWva6zr9X2P58QDvfeR32tip
cPqqi7Adp/9ksQgMUQ+WhRNnkgKXoDzCAbIaRFOwG8vqak/AgzLXFuMoherNoMKVQmUHgTvTQxpC
aWaptkqohkqBpfS9f9ILpRk+DgxDl+sn5NUT0sHoxock5dnLeA/zbMUfbiSPAJ6c10BUioEkFvpM
BZh7cMB1VWJrJFkGzTDgXI3aunDtZZjqGaKZ6SSOu+2Cev8vYYiBRzHUPV64et9nIw4jhusjedhO
vQm3DFiVww+BP71QRqJNLENUBVUaxBGHpj1lCFBSCDqwfZz5dNZ8/TLuzxX2zkRFHOIpyUyxUVZi
ukRNJaJ4D0QisEXtZ1cjL+enZ0lDCsL3ZUe/m2RtxbALdvgPky6vCXWiu4nKInJ22dFy/3qMxQ71
IaEp+DijDyT7820LRk8s9jIR1Cdc20vdBKwCXT5cldTlmyO6k/iR4rRd/fTjT1QXzsT6hE0XXrjD
WOleNbt4Nb4MA6PED+JMPzTpvOdo3WkPPIfgPOyCI0tHgK20tl5eIl6wqH3bANi3tzWHoop1NYY7
e7/l4JuhcoPBqd1MgUxeZJ6Vbs0zca7JFRz0tq9iwM77Utfl52CbfhLghip0mNcjQnj/bRQCFO7h
PD0RZfy2hUTJRCQNeIojrRx4VruO19ezCDLOu9AuvGgletpTbRIr+rpzQmR7Y14ImoBB6ERQ2r4r
FGu+vkYZNJ6uRSIH+Klk6OejdR0hMCUJOQhZp9xFSkO48kKkgPazGfq0xd/3tqXHTSkhZ6HOaPYT
FPBCb9n/sfB5sW/4wzK8VFMkgSZpco5J1Tt4ndDSiWS+a9GyqDSKkLoETMDp/nCsZuI28N9vFxSL
KFw/V+d1T6xyys9wN0125dExhm6cQJcEop9KsKgDAzUSJXznD4Kt14MaaoFDDJi+bY8u83Qt/t39
DfrtkCWP7I5sFGr+MxcCRUKCdat/UwFGvXjeLSSXDYH82b6kwXUq4VKiYCBk5Kfz0opZv/uiB0X7
ia0gSCCOrtrc7zbREp9stVCMaKj/h4t58ZdA39hwasb/St6/GsFiJDh8TIb/HjGDOwc7NM6KyuCS
BGP/XjFW04e/iJ9Q5ENNFnD0DeF6EKJcR1q5qJwPlcx27+uzWb95R2g+FH5jUJcNq129QfTqQUDV
Pinv/5b8R2biOXe16XJIb3/rgjA8dEChm5iCG2GbhUjIUZuroN4B8mk2v7wggrsWtNJM+DL8qm1H
zbqtP/FHIwWsO7QXdbUuJBQ5CTCIGeJC7TMqGk7GrdXbE/3H3IDv8AIrUjQ4DHBoUiqtnFPkRZdn
KgyAANcWz1esQvwAM+DfLuZFbN8rp1IFLmy+e9ZOzhel4SXkKcNgghoAncmsoUkN3vl75XEBOkGP
o67S3Vr+sk2TyT6x6YikQg/U+pymDqrEY6rjo5jEa25KbXRns0f7Fzn/YaLewNo4icMb2vYR1cBp
EKjveCNdMXAgZKkV6l3XuxaXwVeabmbOcKG/elUKu2l6IUHjQmfOMbd1a4YMHnCFGBst0YT+v8nl
ttClyxjczv2MhTWukHdroacEC4Ur0bCr3TLsiZA4y2dNmiRaDd0Ji5hc7o9I6Opf619xMt103xEc
NzyULznVNxj/3+25rBY4WVrkNnOguPVeSXLUBLHLO2PsmIwH3CGOPmorBxyhJBIXHJw/uvZAJXLi
NMUtrdgMO2F+Qin5gFz0lJv+vRvxqvht7Tt5vocPcMkV62jqiuJ83ORBxOzh6teoJjkU8oSMwegq
fBjM983Hm7zeoK9HiUKPhMy7e3a0ECZOXVUOPcSyAFs6+G4WJfqPs4OLcpVHoi9wBPlx3wl56yl1
mWlA2IWh+/QGoGjewItgx0WVCatVobb5E4YkEFe4YhW0Yw8nW0c4mZf1DM3uOahtuiquQS9SkZXA
LzDqYeM+Uu/VrNNydOHbozz+k7eTVgheBM6hKTYmwGXkxwLAPEYlwUJDKPS8KYP2wAvtQipmR+9h
fcKLzvkKKuc1c5rG7TqYjWKKo4J1Z+s192DLlLb1GHn8PcdsA1nprHEa3+k25Ir7gr0OyrHO8RuW
D8Yz+iRvYxkv/CfuV82Nm5/Xn1n113YzjG2nuCs1wB9Ej8ps319+CSWKwtH3hiAMWwVCGF+p+z40
kZAItl5p1w4w3cKYs3dbohzZmnTDJx55Pj7KlV2Dyo+f/c8iW48RtzBJnhHMy4jNd3IVTfGYw+pc
B4hi3zEdpdLjpwGy0mQFJ3eR/HLMc2uJbuY28SsF3NBX3cv4o7wKAQGG0gXdle3gfqSqOyKa3b5L
FA1Pllv4MFICwhz0alJ9u8BVZ2bO9laZowLgRDS00o8nAIWhhQ3KOLRCkAbsjt01kxAkwkHAleza
Vbe39yPXR6OWhIC5B7DGNgLVNN8Jo7Vf4PQAuTHP+7haueM0rS2jnRSYNrswZdWoxka1JONBzcw6
/tkaTNR4FL4lLkGsb/YNoX5TwlReVek0aJAeIRtjITPdTnurWqFl1VFI5L/QoTcdk80zeGNWloG5
twIGOcocO1JnQPlhFZHeiXuqA4NuMe5BOAdTCJ+UBxF6iBQOalaymjgcEkiqIHYXau/g1KztQqwJ
wSh2sp5Wby1BqMvtPAKDMedBAk/N8gv/lU+0aIRq+XXysyG9SAOHojN6nVcT7QRW7/4SXy0xwOPi
WXJCewkQVLvJR953SHfs6d5bCpd1ahS6A8arBZsG47ROhT7B3J0ka4QZRTvTsl6sr710WxLQIaKV
69LFo7Xhe4SZnIRPx3nTECd3i5n7YXZQZRXFL21paL/udNj1O4vvPlmhCxLFk6rX4XrSxaRk+JNx
FOGBBX/v+gUtJHG0odBMjtdesbM0qLYhD16sAWk/NOOZ65Ov9z3SRRmz1nNG1UMNXcKTaSNYVH/k
QClP9x/zDmFqXU+9hFX4qrB3UB9YYVANd+WMgwKixVYDjeTNB4Ak7/RczwzjWXj6mfV6tsCfk2Xn
fAI8Ctwx9e0Qbt2XSnTSEnVLJdbhTuR73VY3qknvmgvL9ZUperL5mgbuvPLoUvs4ugnJVdMRd4Sm
tLjtoRpmZ8EC8T8UvENIYHh187FcP0w0I4JX1m6V6zVzAgURMULFnUYEuMBb5uzhfx9/EllzjPs0
vJhhCXN2977mOi3/qwJE0nOHDtpAuBqwMuGKZEHOLCIoe9i2VH8eatdBRfiM5jRa7DfegtZQWk9m
jbq/qCdv0Sg03WTtHvg82YF3yeJfmw9+ksInCmfRgzCaYERAs33xSJatByzzGzhMrodMuuGL7+0w
bMoBAz0c2VpzcssCh/0tZqIXeSUBaY/Xis2nDXJhpWcoQwScqTjP5hS4t/WSvfUlY9E9PqLBldjT
1IC0rvh84xzJGKWzFyvsVWMHqIuMVDEFpKPf1qSnLj8VsctK9IVHmunJ+8Rwwnqppty4x9N6X7NN
nmOk7/CDvNGMevv0robgrAuk2R8SgczmRU5PzjdjbgFoDvadeW7NOCPsyGRI5rnHF0W8pifyQJJB
FDa3yKkV6QdKf0rAsGkI39D1K2AgsJM11yiHuilIFlA9U9vEGePvouzmQry8/u3/dYJh1PgWo4Qk
wliROAS6zXATlJ3rpr0nDCBS0BsVxUkdTATGq3Bo/MkwCZj+4NGw0kngNds1lj7aFNpyEt7JdKko
JHToMIhEeYQwChnrZTKDVKRt23U72LRlyaqDLHwi+6sj3AiudXZ8qGUwDYI7AeFhGuA8vMzCN0jr
Ei45jmHsajzkl2n3N2ZSJ4A9COGM7h1FVm94jOTblTX3+SBVItT73qbCZ4cDPcEdEO51SmzH1/s/
sGAxE5ZXcEAi47sJlxwy1b62lJylsOHeUvxCbGZ3E7LxlDxV4hmuNHKKWt1248CplVdHWKlW93zq
Es65QcBfe2rgUJnYltnn3SwWXaFa9cGOGWAzDYg9xGsLjAdroE2w+T+HEtek35TdiSfG362KoMrA
5Y7E5CU3uFgvCIAjpUh85nppv/y6FQBJA1EvKfOJcrkQUbZ+70hSg6M8BxBUEh2vscFPuS5x63NE
PVRjkVy2LZp8v05yroD/I2wkoS57QPuFAtLXT9zHU2O4A5ieHsora34FEaC4/YTmkngKPQylyGzz
Q3m38K4ZemhFwU7tqQreoC8kirDRPl1KzPC/VlEvaGshmDObxqTntmvPUJKEy19yqF+wKXzqeCMi
vTYH/5p/3I8wf3wuAaLZVDM5KCEIskbG6Uv7XB8Gip1EugYV4ceDy7cgSGRrSdp+e/orG4UQFPjK
i/9TOqu43aA1XltiSFTkMzducDylBpLKbQPUitbtgwGVpKnWexZgoF1s57BSITxezEDYqfQCTZI4
T3KY90PR2EW2oIbdiH4NvQpU+ZwDjP6e6R2oi237NHwXs7UXBYvyprrv0kpRfzRgZ+m0quY70uUw
At0cp3w7u4H1Id1pJxnhHQlvnE8piywu1MQbq/jy45gydoSxHj888rrC6BYGFWdelJE66il6U+km
SjVTgAo3+menB88NqE5Eleu/JJgRFlDlJq7C9FCLiqtcE0mE/KWjheo0GNdccPzHfuwxSA+OtqHY
kfYn+gkjqcUSXXQO2b5Lu3QFV1OefGwDHbrWLScyjSaa/n3mUQtWT8/ApG6DyNb9rTeHfj8xx/uM
h5ZV9403SReVd4K7kYWigipJDQIteXDkFeGRqX1zU8+OrBn/2B96kST57jPle8gXlmQdBUF2fDK4
vB05ZW8Ki574dzyVuez1gKJMVsn/jLDjlOKjEmB3IHY9ytgnznkwXJbbKeOKVihfRU7bBI1oOIXS
hS45SBtGtDPburTzw7Iens1tP9hI1OgnNCmCv+Ujio5+eog3EMZYRlxPkCSujGeTex26VAhKqq6i
gLQFSoklP6Pw+442E/WuKP/Mp6uBWenxmc13G0DgsMxAyQCMDMatid1Uix2j0sf3ykaK6N690MGU
cWgeEhx/FuEnYVsFfFnDS6agmJ2hahITQQipZaUlzO4u2vbWoRxkE2eCaec2oWCk1txnas26+QT7
cRszcT6T5WqytyXI2ZFvDXIquLW+8LzzpxoauoA9PlNNNKdSz21PIj2f3kMhlK9Oaph+NdjJbp3c
521vxwNH/Vc9Cv3A8Rcpk/YM5CryYOwcxIx5xTz4ODUvknVzXdj+yxxNnrWNDSOa+1lvWwSGFuVU
ASl6I+CyT4OQNPgFI1P32zuyErIgZbzV2nP8zdPYLDmv1MavRAQms3PqgNfHy/kDbnrdouuGWbRz
46MrS6mjM8/PorjwpcJJvo7WfYSdQGOgbsHTaC2Q4yg9UL1pQtntAh/syXavlAU5v2fSfg/JxsFH
65oUBGWeIaQ1u0fy1zEtKDRIZUp5Ln8YMrqD/t9htKBHHO8767PsF2nrsnveBdxdOBPFRhGq2at9
e6cY8qrCVFvNHIkEpPb5phmccDEZnI518Q7DNBCzkwJhandKryU3kOFhxRW6HlB5Deky/TUq2Leo
4eVAjUjvQ38weOBH6EzKkA4TSlpWi7JI9hIgypKxbCRunuKUYVrvbvjFXA567mZ9UI3Ekkqs4lJQ
DZzoVRhY3frIzOmp8gmfjt/o5svK3PqU1AM6kk+AWeJFrEz9fXkuC41y3hv9GXer9gbzQRyodWKm
qzomJnPH8Z6Ghoo/ucgBeH0+MoNFZHu7BV/IUOLpiHE6J7EiQmbIe71mrHq9wHwHjD03JFfVyo8P
tzgX/y+942i/sgUlmehF53F8zDrOH1BLedcaM9HQIxveqwB8kW/8SvULX2j4QhP4nAGAo/E6Fn+M
H6ohdbY/FW/dAswJPWpl91ajH473v+vhDCZWMIBoGUxC+lhvq3LPvhodnsgaPKXcvHmJWGt5oW04
vRjcJ1ZKrqZgCzNuB90YJn9vWduCif5VjQAF7MZIXj2f8Obhg+wmNY7tpumvgCjDbyWLwndd5CSG
XHQophPyt1zX3BLXEwcIWFkBzre5kq8VIB5b/lU91zlYJ+5QV1eWCaa3yGIS3DwYRacnYtOFJoD/
wXA547EwwGdiGABlNuYj7eD6QrTB/Lhf94Z90JAJI9S1b2FuzGJypjB6Ij6dDDQVgMiWbaqOt6kY
mTPnOQ5gTPZyYhqZQLRdminT4vjpjtOHdpVpgrRtLvEbTl3XmGciOgsSmxn+7s598074Ali45Wjd
4l0o6ghmcTgBpbt8Qs7+krStcM3V72ZkL00Gu2zI4HFR5CZCNhGsnxV356n6t6e3IydBvLYH44rL
lvwm2ggRKAsevxnV2QdxHVxcZTLV7Y3gb2ynBz1k4+pda+5zYbtffLf9i/idR4+cRQRVmn5Z5CfO
GvTMicIC7+OLttKGFFGvnQR6uRSjGkskA5iPa9vlsJ8vsFIhALWrUotT6tcX01M9i98PsuZ5Iear
E1mYH9JZKKPwhtOA9BGDXRqBwkJxY7qmT+W5dIVXKsVAgJs3Ha89gahKHe10i8NV/TpyEVMiY1l5
cI2CKiDjpE/QB0kU9R5/1AUH2tJ5wWoj0JCtEwF21zZeXYvTMySAWdk6o8GIkfHU5xmnEEtF3eKl
FmvLzNWwtk50RMijN2+kM7oc4LQBVMF3ETDrnYzqoVCU1SGuK04ELY/UUjzR2c/7qjUo4zf24UJw
MM4IBsCknYsjpCNAypPBBPaYJMjtyIwNEGMN9yfJtDj3NLVD05sMcf1+3RWiaFwak51ozKmvfMcy
yLoJYNutCoZfArZrpTrdEXXXrHQuq/H7Da3g0Y7QM6PGWMghV3eNodrLjpWIJS18CZX+b7wVmCBI
UEan1Uga6/3DnmYaNqb+6/8Q1g2T+lLqxfFrf+27c0g32rcfNLxlkoyqaKyZb0Z4gf+ri1mlN+DK
shizUSDHPBG1sD5H7DR0LPqGCRYyAfGQi/LLY/UdWHGSa7e3zupuFmRYGM2gVFK1xsZQlRr4UIZn
kstlLgMHZsUVR48izdW8hWN0oZy+q99KdPj+WN8bCAOiSvd/eYe4oAfjZf+NPjr1dqR+jsnE0HK0
rog5DA3MtsjxRo1vzHCkGZ7+nIqFAWWv4pUOiy4WTL7Sl5IHgBddYsFkrRdwpIMJzAsumq9PFokR
ACpG08q8Nq3wo7wwksXH0TBWIpCSWdJkcBwBPdHU0fn2iKVGmTRu1DypVkj4z7kYleUdUufikeBu
Yoshznwe9F1xHsrhsA1FJyTa5LOKOYx4pCHwzkR4ffK0e8JccFQqW2h8KxC0XFGrrgZMHuMppyAN
E8ynJlEE8EiBZsrH9pjj5VluXymoaJ2likP5xz+wUcSFdlKFW7SO97H2LxaHXf7YFDEyNe68h60r
+QFPonvdCY1PeVPMRleDcCW+vT9f+3c06KlYhogytr+n6PdFtb9TywT0mUSQ5caQiFSoIAuhu/yQ
qVUiXbM44MrxGWzyqDXwEyc1OQJ/ErkQFCGx2SS6obq1DjdImWvnFD74iWs5g6xWiP1D/Hep7Kr/
uKbHRE0areaABf9iokEVjsSo1oJ+jPx7Of9iEPxneRCX9QHoa2CAaEq4WyjmD48cD+hCMnezO7Xt
kcHBqL2LF+2mrUs26DCdga/yurcZiJpbAU7w1BQ/apwIMbjAOL6UPRxD/bkN+DpA0PImdXiZnZmo
HT3svUIONVDkza+VOX2FQ2Uu0POxWLjwCXzsrZm6sOHI1i9ny5noMDveQtj7rgBG2FBWwZ0Ol9jG
vybRGQkaOoXCZ/ci0+ykVI4hs6ZIpjbHyCp+Sof7oT9wEzmhgyVSkJCtnqTQw1ueN/O6ArRFLNLv
K5oq2qqTuz1MN/+OaXDghnzNyn0Xp5js4jqEQC0ShFzuvgQrLM1tFOhKWgcb+dXbYZTvSKlF5Qtc
azOhoV0pXYHFi9lZBuwlKaSamzWMnQSg6fumFrzWXGu3bfV/BEo3x9U+cyHtpwilir8gmaMAURtg
viUen6umde7Yb69InkAR5p6ka0x80n3k8yAnqgDBPolZRDPnjwF+70w3Faqpu4O7KvL4skmkH0rU
PgBF9uazP23wZw6Imd5kZPOX7dLoc8+CIAP746iGX9W/MXFEfPZ8ksegFL3jr/yqC0RWu5O4pCYv
lb0cDjEUmo3n8HDKa3KpRQrgSfmlMhqy9pxAwwPqmQSbcMKd8ECtcPWZBpcGc+a7yF5dlEpbaN/6
+aYGj1kOEiKdiBH4jgV/d/PCwWOVSu63cUUt6OEN/OKcLR6G9efbMzxHkN7XTmocP4gOkRHeYbxE
G1I6geVp8dsfqtTeDD82UTQfMti1l91xZMf51VqqkM7+BgypTdYKG5XQjKAd5m1i/l2n2Mu5IP/8
Svyt/zkwXMtBc8WNay8W4E6pbCHSOjRhp/bmcOwew1zb5djH5nEAytMinz2tLg7UrTznLUzElZ+y
XdOoa45S18dGCdDUPcotBUdswPQJ11kHwPX8uxpMZM0aJ6HjmBPrFzbF05WeMZQ7X4HcH3ItvyMS
CHZxqbT2CytmkPYKpRKzeuU0LJHSn16iylI+Ff2tfqG4kBXa3nz2MnFC+5qJ3jrnlAydp6jwGNK2
KNctsQl8DJ2A1vi35KQbwqxF+aOwu61M6HKRgc5I7RUmWHj/XwNnX3jVzoL8RqSuEqbv0soaZ7lw
FbyHUL+DdNPOGMPZVLemZT1bI7LrscHhfsRCXQ0aSZhTtgqfddSS6BTqt0KxbVqJq4j+DAtEQ1jA
qerxzo5VWVRu3AQV9ai2/21bD3lDGSSd/hcLNDs1/DLMo+qdChZhPuwwvvxLXXDYR0JR4A8RiwVq
LSndlA+2zMV4NDIA68T3TAOhHzhfs8rnVSCFuNgDuyMyTyQbUiw3j+jc6dSx4F5jBuRM2hESI30K
aze2czAUGIRXyf2R/YtuYzdOwsOXOJZYZNTIsCINP9OQi11cfyokPkazT5jZsXrT0F4Gee5Tn5dy
NRTnxXjcmCq8srtMvyKX84/i98NBHdL08jNr1CVyk5rxg+Klr3JPBA0kYWOCS5OhvHyiMaYdmKRt
74lT8KracgU59fF7+3aPcQnh9ioJsFj78W6H43lNFpRaJ6AHiynXbILLfnYJdIqOIwGVhq3o0Vxr
tHZTYCPkRF5Zff5yU5taP5SmFbCFGRvq5RClqQG7w94PjSSj8rE1m87ICtht2u36j1OxJALKOqQf
YKU4k+2IZCq6jDjtc1HENFYuViXXiI1grxcHO3+3aBOk7BcBc3B6DxmY9FGviKNDxaKjIztVQi1g
4UQ0a5mbUcg1HAgd/EMUbAAMMTwDuYNSyQ4PZAQnGPKiLQQDI9SWgADqhfJSB2rK5LyYOt+I2FYK
YCL/0ebCBXKF0PaJ2O0vvapjBemBBIL9+me6zp6k/G5mXcZ9bdxepveSPeRsT/sTfzqamqCxnTOn
TB2o9Ce6zSDW0MM5q96BpANGQ9pLMhV5MjKvAzFUclTZZA+2aNgDAduA1QMAR+NdcuLlRG//6fN5
hDykjBIPaHHjfZg/ezvmucI0wd/RsYN+ddxbUN+RwQi1KXqKh6eG3GsFQcODzQw8nndvBg3df0l7
KRe+N2VVJjHl/BvlCuMO4wzWQKDPWa4MlZxNp+STMTW1ngi9/qEBPLTM3Zq0SP28y5aNQCrIrXrM
Q87xFBABxKKFMpzEleVRCZ2JE/dOJpqTNoGTYZ1TBWD0YPLXiH2YkQTYcevotVYeLzntHqpPYSsu
JTE6or+y0St+p4zk5r4081ibQuiT9PKWaiYRy426Tmvh1TqxDcVSe9MOC/QfYQSak4vwlPeK+bV+
bMq6FvCNDIiY+7YoHiE+Mw4oEfjscvpYcZsxej0MWW+nHf82poFUSmAS3mjsG/O5MabH8FvYlLck
s6DrGfospcZiyMVZfA2DV88wv5YYLVb2jUkv1jReRUTwYz0Q17usQItsSaBTapd8xLnbR1uvEECn
oH6i5aygjXiKN1rwRFJgPjFkKrdEpINulirQmkUSSD/8sf7CVQy1sUYTCu/AIbv/+WC+T7F4rFJh
ENF7fIDmsXfXQtuOT3SlklHOuzOv3I+/HFGipOSIcGHUGys9ovYsMU1vWIoiQCuwmPY0q0cG3gnS
tvZjJTQY+ejSbSqV3aZsN0OQ5N4BwEy4g+KuFqWY3i2onWzDNgD4pKDUSocYpS3dL6IXx9s2CuIS
dmFtS0V8ejiPik8u74JLZxRWAzPvM+GwV9ABsT/j34YOT/SUxEIhKH6bkvvx/faqzN/3C4RiPTtu
3hfIBJhP7X/fLXDY6izZYlRbcPn7ww3Hm8TSOQVhsRcxUSSAhoIo6lio6RDPIarVU55c6h6areZP
02Ui6feuHdfC48FGUpVvffphHFHZNmg/dWmFc3riDRIoYREOV8UwzFaiWeVyp+5T2ZID4UI8J8RP
0JZ0RmgnuCjFa9qFmuEgsLuODSCLPrd85yVcMRBHXCRFznEXoQoAI38UGqN52bHDTpP+3ar39cWn
DcJtXnqUhJRBE7snajwtQ5x5tvZQZ3Vf40RTzOM5o5eN79Sw0vBx5QkSWwvQI8ufqDrp39L3+8wQ
MjOiPT1CZW5AiW7WY8JdptvxHv99ySB37Ewh4r6q1vlMirUD4Mosbuku2bdZDYB0vBGFCJgrxH1s
6FBaunAzV2iZHasALuxkTo/1iH2kEUIiZ2KdB6SU3NwvPbW1J0qC16A2l4wH0Z29tvRTEemMVozw
taHJ8TdpQg0S2n0PjnVT8v/ZSwdEJNyghoaLdR+HfgfuxHu0JYJL/JyVUZ7VWLXisFBA9s1hyfqi
RS5p9U9kPBdgpQOjKIKV0k6FsGKAll6q8GiaQzDjDOxKNBqX5Rm8GAHLw67pjlix3MEysDA+caqK
KJ/Nj4FgeLZk0uem8PUOqGzfOEGLK2DbGTrNZA7alRqhPYDs+nT5R1Yc7No8O/FOZGYXbuO4incj
SCwB5DCdUUSjh3QUOPMW4M/ogkCCBTY2+pNapUiGbVMAec9Px5+t0SMWwOvf+wHg2w3RHIq6FhZF
WU5dtgMdHdIAMtWd01Ym8ug8hRWEZduhhOMdr/++lziK353bXsoAzU7s8qYWSNju6iOW5p4wQTk1
Y/ux3l/YCnrFD4JDShhRcV3WTFzQUFybEwcITNZuP14Ni1XNgAdJ3PI+BqXdGD9p+31yOjZ/3KVW
gBMfaaoK/HdlHWd84fOpZZgGuUHiq8X9NkdnLUKAU9Czhn1saK9Fw4wBp36YAMne7tSHSXOJNpXD
jQO+K2EBp0p9/CfxYpmsCKCcx7sWJzx6WGhJ+dkuNUr6LNyNe6Hs+FYc38DdxxRDDj8AezkIRG3s
iuMn2tVACFKqOE2lh76JY+4hvXSuH7qgfzZGsIKbHAWODJ2OXsRpPbIgwNkhcO1cxIuGBhrvUSWB
Dq8xLa5sQO2qs4cIgFcGRrCgp3Rk90OP8AQKc9yITBZwv/RAhRaoVK/HLUHcWFBb5fc8qk3WRaYs
ryOsGyB30fH/iBq/cA8JRt+yOiiqW0CY28vjrbH3wl7hUMdDKH9DE56DkDLvg6WRoiRnThFHFQMq
0afcR4BK49VxPTgzaztlbMqhW9/aWBAumq4fTcxzOtTggBVhLqldJSA+/LbPb9bCe8jfmyxIu5ce
wXpWKQVcdVEtgR/2HgViYWKTQLr/9VpECcien9GLIxdEB3bn5NlLzNbwbSOs4QrLaZ0tYSqKjAtB
Z5UJzdJGgwrmMWkEPozHkk06mVPMK3U6DP7h1ORZX4Qp4VRteUqTEkHHXqtZyxmvq+JvdZoK1HKI
svWr8zHosgOUGKW5n03WAmummZ8rYF7wfb9flYb6NnC4tvz6HnrwHpynAV2v+cTHdAMTSA/IZrPW
6RAYd8P6bF99Z271F7K/1B5EUNECI6U/y12UShX2gGtHf/18AIGAATE7b0/Nw45G9drP1TJci61K
4LiMtnuUY0dwcc+xwsPyYPiZImMHQWb17OzTYqfT6WhiP8QtREweLAjUmwIpeBfmDUKBoqQ5q1d7
Ql9aXay8u6MzWbve+PzQrV9KgONvL9l/ujEqsu7gpYJDJXzivIsicu3OoMfvHKbwIIv0Q881qqu6
Rmf5r5PBGb0aHa/Kh01ylN6cDznJl3XeKEMLhmrbuptBioBImqrQWMyxVZxox4jG4zaw7jY1DHEu
EwXCleCe2i8L/LLC8lYtzDK7CDLJ5bovtbYaLmegYA03dPyQIq15y3C3vtRYEdSc7zJb+chVoNNj
QrTB4SvFLNuqsz5mm1xL7JLtcaMSm3QjvGP/t3/W635lve3qtqGyhO+1cfeN6pxjmTlXYWKwHrTv
UWz6lvN6d3/lkbSSECzQnttw9ghd/kfTKbdbbjjKI8NQI3eNj59tZDhjsa1DX5CZ7w2jm7sIAOvI
+5jOXanJ/17/bZDMR40FjoKUetO5BIJ/Uuw9nRJRjhPWJVK9hXmdFxU26I62pl0IjRjbStpRC27t
tOUtcMv3MM/jyYuSVfZ+COHYIX5yG6n6oxo9iMaOyFxy2qPLov/d/x7fJ2mdp6X/3YZOrQ81rRK0
Q/3I4SmQBPZR+/eyJSF9N6uyMG/ZWY30HokLSauVJnEInqh4tggcMytYRFcAlMnVDBmASfirJ8uT
tQxamiPhxtX4ZsVocmRZK+3EIsHqDabeqki5leImRNqct0RRyTWH4dTfKhVitlIm/PMb4OK1Domo
YfyLOwR4+ZhQYTmbKvrtei53fwgozT3/q2adLeVU+znDjQqXrgpJHSmSftDwVIZ1oS28pLXWHT8b
CZ1khSuPfQhuOm9KXxz36TvoiOodYaGwpEtTClkjQ4cz38gFd6W05YcFY8oz4APtqUyPJgY2pMh4
L7AsYo8Q6q8lfWyBlO0rWkeSlLkOngWc1D9uwT8L5tvW3PF7c+ucjIusjpBSh1dMhgidTfroU1d+
C/o4RJLVvIDq1tHO9BVvIfxLz1rxL2QrumT68JC8yoJ/LWBPEk63sHW2hPUC2dGgNDODeExbbQ1C
wHlAgUC7xI0B+UmmctyFybbIA+/m0e6p234GJjBchk350KYF3XTSp9leEs45m0az8X84v52otGwn
cJniYmF56a3OTVnP/re1L6XeiglAEswjOKWrglwFnVY7P385wIz3dELfB6pbDyMzY0WkoD3bDqrV
Sr3g81zpNVW5Rwzxau/eiWBxh5Qq29TZYMidwI1+lTL2deTpzgCiC7naDHe6BKgZC5yZfh7D1y/5
6QmOqJBWHZk/9Yqrf2w5ZecA14UREeg6KxM9LAtn2lfqsDbidFS45YG99Fd2/5lv8o/sBCJarnRh
J+q2HmEXxvlF56NGsr39pJZJshBtNdxMxdVJgTwLeIrgsvvRa0qwtjUwYEfy/7EJiCsDtbBf3IKl
tJzUNaCO2KvC+0uJtdZdKe+W/h86fuZOjV809HAXes5tR9Cp9PZj9/yz7+UA5HnHPIEg+6Vy4x+r
KE/jq0FfnCPzU+8ww7wOPNNbrL8kJTVYXL+fz2/1R3lfnj9YBPMRUxEcEkDo2FdqfdvafU7u2Q8G
8Ze6ObjwoI9PtfeuSlDQIh2tc8E6frfmFdrM/YSMvK3q/HJf66sKixiFUx8BMqIdAiKYa3EmDmgu
b6wmkKOjtSXQ3wZNTiDHKZQPVEzKWiSxeTa4S+aZtxqqoYJPmjzcanVUicq5mlkJsjhGNTGnRdCg
/2CH5c8nfGOZ5iWO54FZuaIFFWzA7fcsVg4ATE6CsiDSJZHL4VWYT6zB4ru78UZgKmZ3Ev9OOLxD
ho4003cZcd2bylRzL42Voe7GXMl/1ImnSXTuTdgbX+tlRdhCxtDYhtVIVeAV3otGDLyBQMYSfG+y
BOHpPUoC92Q4rR7iGMFTE9WOIhzvIOagQpuVi9gunyF9ekceOWN8DFTiihKFihNt6k31/4dzQlTF
+VduXaVSB9064DQjhYsn3HNkxK0z+t1kmk5UbIv0VXrYdPbdzFQLMQfBP3rLlmwCw9thGAK9VOte
yZ8msLn9WXB7K/yYWfYVjIkAkSF7B1y3QSEqoc9rfyjkcUsFe+X/EC/zAWKorF7byfG3PqAbLFEp
8NoG3hEvWQZqOznGzaJiJ1kGS6MJJnE5mYNwWAnAqBIDVE4g36Jik4Bb5ha+zBXu7FOS6BkNBk9w
ssmeDrZI1d7Dg1XTX9az42Ex6lTjGzZ6GLZOm8virQqEFYBkDtzeHZIvQFnooPn9sIzn4r1KAcwT
cANAiQe6ofvjujWNFJDYyJJrrnmkRxYjgQzpYwR/2Bqi7v/AV1/AJd5yan84/NC8hUShNZwPezJC
0xi8q8wQ5pyuaAYsef5uz7YHditrNRwtp31933Rkj+f3nrWphP6RD+omZOcML+58lEcgV89U7o8F
h64d0bOP9Bwkq+EQZHe6DTU6lvfr7OX14J2xTrGrdJE6LEuB4zIlTxZWSoI7SEd8K442eSWXfVoK
oHQ4Ntm9u828py5ORV5AunvMcd97f7nMgROOJI22afADVK3847XHR9NlqhFyjCtra8xiZYWPj+Xa
Q16HHsQ17INrfAxIp5Er1oXwMtIDTTi08Brkcczav/cjZ4hc4oszJiSS8kr0e/RUkze/HAu+sBOO
a5EvELbg8PjLENH93RFZkCFGYjoCAUQiGTNipkE1f3zQr1wJod5Y4sEY3s8da4ltWetLex22IkM9
ZCmk6J+YDtrZOlWyHKfRsDzzwB7cW7CFHvOJxrjj33K+X3eAOScvoBrau50qEfs0ZFEF3kC21wIh
kib5MiIgVa/7+xAytI4ZFoompJ16FyG6EcjhzUWmXUCcGBZF8IUaeaFSJreR9pMQclrvKKEYmB1M
XsSPzxjv4cg1sbGlsuMwVL5sBrD1K+oBOkH97BQomd/beA3IEV9d/IA9Gw9yAXyeHDIMy+vx3/JH
qMKWFcvD8GSyabu/tRxMqeTsGimiZUpEWWoXpv/1QTu3vIwQXXyC37N3RQWRbIItA2XMWI/zqS8t
q6On5C9vUbxNC0XB3NjWk6OH/Us6O1qW4f6BQuDIe9T2v9TGZ8JjhsD1875fH3dvlxS8feKTXEiJ
eHBVu+VmhQ8usBW+7ARSqH53PpT7g1SOrj5qMM2/+BKXqvem/8oWgmzElbOpsNgckBfZyaJ0lN5i
0XH4pwTdbQ776tdv+s8UjLLnt59U9XOqXo/I73HNSpQJWsugzF+ce+P9snkrOwPA+EknfBBHvGRz
OCl6e5WU3ofu04mMieNPGFHgDCIqdLlb38vdeP1Bo7JX96gIyzd46lTtwI4IHQrvJUSpiOct3+cb
3oTVzgyQd5rQ4F2YpwC4qxQIU89kBobIYg6O7q5PjgfkFksfFwgFpQ4O6hpEwBs3oVJmU8WocVje
Uk9neWeiKypMiUrtkTuz/EE/L4CRGFTx8I7hU6do3n85KUYtZq10axqAqqj0behagIgm0dipbMg6
bqv0dMYJ8+nsBFA7ATy3xh/9rWEX/xxQKEBr3rYg1oE+1/6mbaxdaG0pKqPEc6MXrv2b0uArikGN
UjsvMzoPop0a1vtvn9q9crWzUcVoXu+d4sOpf2UEMGDsST38P1n9x0W7Jbl3VFDWtrI4B5zKO7pp
1S2Tdn+h8y8ud3oxMkZx5ID9VGe9Ei3BuXTU+2plQoEOJOT+lgqgPnCGrnaKjO1f3KrO/5BQTVqC
HltrVAU3IdnXiSzcZfv/feIP7/eaeHEk0yBGcujpCpDiYC02eZ6RCgwDjscRSmU4H5Ss/WBQtDEJ
TyxTA1dqTRXb+MWyALiD4Gap6zfDyIQB7h9+efx9690k0eNd9fwkJ/BbuJA8UNOIIqAgfRdPi5ah
wSEpNP+I3tfCzGFDF7JDw9Zrw/DzlfJ8PewIvSGtrI2Hx/e/UL+JBz8iPccXKlPaS9TTdN3DuMJR
vx16gXSsuqeiVVK7VtQbUYH32NltBziWqz2HkgGije/8ilNcVbkaBV02tFkZsGiG+DzjC3PLDb3t
4d2qXl3gEe3vE9NlfEBv0Qi/ninpVbOV9vs/uBKIvJLwmYZrghGhHEW2jKpGCdUEq9k59G0FLeTH
UjYgViknKr55gRqSWd7DGT7kztobWkCo9LCuQolSQnP5502WbDAN+UcDMkAWC68VoG15ZxvjIWjX
b0+avOCe/dyPEbWR76nySXZ+Cqzk7CNrfmVPWOngsyy+DcNM7fP0Xg6FFgcUP+r03x4AKGPKFJju
JuTpV7glBsEzwZDmawQ+S7Fk9i15c5lLfg3UPcIcnHZzrJNz1qRR83vfirh3Sr9Giu4mw3c7gmwg
JPWmyCHmnDlfWWkeVf4bEYd7wih0CgkHzW9msJW4+FQ3DonEaRPN/1s1fwYEXTSaURJ+GvxalqPv
O2MVUYiWkugFq6ElgRROpSWaqa4GPa+pzrifaZOeSN5W3DNXyh08P8luHPsf6SFzzs8i8WWBQSVC
GpsWwdZVWifsHdcGNi+dnktcy9G1gHOpMs3b71P2PvEzeSXQiInbVTWmEx88C5MOX+fMgPlVZrJc
EnZwsp/jOE2AokryLPrQVxFIoZYu9hHkVyYxUaIw9RYBIF3AqwvxbFPMiAEx9CBaFYyudKR74JpQ
OCxNDUUSg4aKzZbwzBWRI3+wwdNd6LjW2nF8lSVhIQmXfGYDDkeeC7tNTibvQgdmwbRAGyNTPRZx
VR9LtNOqaH0uPlgiFHnRYgKLaYbLWVR9tFizmDIfkUPt64m51I3g8gd6JtWSHYHD+PIYIb0YNIxG
lklONmHq59FvLkXEcw7Ii2aCI755s1RgI7hmvzSdguM/9igtynivrOTJFjkYLIe4iIF093m8cGrW
lr5E0yeIn9tLarPfZ4Rg0RMSvnod9P6jm0+hN4I4UUgJISdqwF90O0Qy4FVfr7443mFn0aw7KAyQ
xonDM7Vs+w4Pd8pYc6cpl4ca9sqc8mJW3khDYMnRTmI1GzGDfVcp5Ze+xXDJl/93VDCbyxK7EYl3
hDBLoCxC3sOq0ypgKvG/Abz82GkLITeZceK5knnRam7Y/Yv2faHNUY5MqbF+WmBBpHF1N9tzAydv
o2m8k1esD2UQsT+BBTcwPMzJAu/ySx6v/kgG3H+Cnr7aJy6y/pQoTIbLkXjpk/httwZifqmL7UYt
785e61d+cR8cNI4XLuUKCCKIKVPHVC4/IC4sTILmEHMbi6Fycbvzvc95hR/HsLuPJV25WK1pzd/z
n8AT9wY0Wm5viYCvQV+mGc1VIIUONO+7kf3nvhOu3ScXriQK5htzq5WB1j2hYOQ8AW2rx2jvzkjO
tQMPgqI7XXhHYv6+zG4ku7t0GpKj83INpD05/SIboAPX5Zubi8fLeytTgjyRSO9dvxbyZVzj+ke9
SnmaEjZFtyO+defbISh9V5EBC/xbf3ayynUxWwuzoeXW+L5xK/ThfPVciE8AZNi17uD4QTbxS/8T
v80dOiMdHqjq3+rTgebnoNLeh4m5YluO1e7x9Ao6Gd5j/BETOpUpD7r6bZZbd6B2WUPqftriNu+i
ygjqiNJ/P3+e9XgEcgHHDhvDP45hTqiseZtBkoZJ9GMtETPqbcRetw5Ig2fJwvEqmaUAkMpqzfdy
t3SyUB+xr5sj29/SQjVspiaDWm9eyQZV/DN137xFw91YkRgeAWjhIYs8luHn6dvQnm3qAR5cSrqT
eYNDp6utmEuFAIHgh5vZZBBwXN/p0z84DzQI8yjXqr7IPTttPnHNxHtM3M1h9h9yV+JXfDHtWy7Q
SabKQOAEz5TY4qUzDqrxSOeJSPZs2j9qn7KTE+eHjls568XX3zvdDVENiLp3CrjNPXzunBXr8CaL
YuvJb+7PMyi+HxwaW20LARt7R6VSspOSn9LG0Fa9h2m4fVmAEpZl7tJweNXPV6PHmQD6ef4bUtHE
jefEhBT69xbBb8frxQ3cZBkeSVmHalsHyXiwU60jsz0HSobHH7VcKhBmWuCGmF0nOvjthm2RRhka
n43LK9pZjNP3Y2PMyCAkF6QJhiVX1iTSVqrOKxaUAyJkSG236fR2unvY90kRubT3+I/sixe2RM2S
Uu1J5JAFhCfpfGGlF8xzBm+/oIvNxh5PvliA6c5T/zV2vRFPjcgFFQMXhLHPC6+rGmzqoST5xxhF
KKgW69euh7DBf+mx5LN6YDAlP7H9rnVaWRH60dSdmlxJaikuByqdi97J5VKrkNFAizXVZiJyJgby
Iph2gIJ9AXy4jynLu0Wwi5i+iTSK4AjMLMOQld3wsMgnCZhadA58d0jKrm7Mam/sjqbL6MUXdv29
aBMdsy4DSIUW6uSOstFC+/a7AlY1hW0mPSN6nuIIlgk78rYJcEN0jC1LfGyKZf9jrI7pNJeqkolh
bkeEsIBkvXzsBaRss25WmmhgmkV7vBIrzDQlX1AeaaQr9QQfisT6AP5407uAaaLKMgbIh9+B6dMe
YjbslM/GCj2AiBt0HEp+NyBOR+VYcInC9l+03mvPvlbhfWDAe+WgeTtSjGqa2NiDmmLYJQoBPxVZ
FZgTMmEP3rUyYSMj2JPim7CAaacjBl5RNGSLekvcVojq2og30gGEVCPAJorjpJM5n/ii+cehmjpU
q5k1o8S24FnJUtObi/V/6xvdxHKdtEJIVg6bEbquD0Yf+cLB/AbrIP4d/Q3CZEpKBB1UH5uX2Cta
Mj0He3FTV3MnK1JwddDmvfh81f9OzXb/E2LTqXR8+lcJiWbwF0doDGNVIuED1psvH3kBo35qg4gq
gFrA3YJ15hDuRYgQwNj/f0K2PsUT5zT+c1f0zcq5hsTTMeFtukpfSMw/VekjWjTFx6XZWDSHel9K
L/0xsdL3XtNscXJCQfohfp/hT4QHfM7dzIGzY7iL6Qb6Q1YHdmOJAS+rmQNoo6eLmxy8iWOwzwQw
tprYna/owX9Tg9FgcFgEL/QouM097Var3jBDQyZZkyHOzez2sajaSX+MG/PMqlgGzF0gqPUEoCCr
8HgmoFS+3DZ8ic/4gAQH0sRlEXUNgIHnG8koiy9bDo78mUkpWIOdbTf3PdnWmTbv4W4P7guB+1ne
FsrMbTByzh8mU9qh7Rpfrk7JL+G3WqBbFvrIQeiXfZPCLWo57LH4ATbs588BfNJiIVp/sRiW4qk9
JKwEUAlJ+aeWgf8H5Ctl2jHYuyE14IAGSlU5g++9rNjbNZTiLVlAvD7ZUph+fgz2A2JhiRIxSkma
66PliN+zDLWFa84azM+ZF2V9d4s4Ohxe5rI63wTryklkbzVunH9sxe+1i9kw4DOjDwVWkW+U5aMp
EW1AzwX5LLV2pv7RtIdzZIB/1GXJKPAdMBPs0C9cnKxy0McqeVHNQiQGpiMgG6rS5b9/5dYobRrw
TSOE+bCTvZ6XdsJjWLYdQfeYjhtW1gwpo1zKqYR2OS7cAd3fzcvQpbEv129X1yp2ix0pSCLdU4cQ
YeK5Llu4d7XGA5LhkUryDsIpk+VztTbNzf92AmvGtFInRvDKqpaEXvyp/ieJjHML0ygx6tAlCjCb
Y8vdODxur0DPY7NJ2QfvqL2MHRTx8QISN0hPHVNQAAPRh1CfXjPFWvfdlf+aBgZI+He4Qq0vbOuJ
WP8cR/urRn+0YpACKMJHhtDM5+/y19v0u6NefrilrLBkoLAaKiP3QbzB49xTPTwp8AgwFe/RV9zP
Euus5x6Uoas7mUOi6pVpA+R0znL6z6APYvBirAJGHEJ+wQ72ce1SjMuG9O2VI4cG/2X72s4k5AJ2
o1S7tlsoOWFCfmfaR6alm4cOVlhALa5B4n2TYCvU0Og1dYnJ6cA6GreL5idp6oqmMeEcrx7Xpwbm
EYbjbpTo/J59XjVZhl4UBBOh/raIFJydX1xYkKAWpZ5u9Yo1jQzc5fEgpu4zWhHaZiojn8Xqlof4
HaeoDHFNRPK667cm8c4TU1g2/XuioOE7TdJdtHeQVMU4J0rBFrsfoRLXAx0o5PiqWrDXaHL/pFoL
nQnEQooq1y+Sujo5DDEh1cdZDlUMWn31s0BjLt3IvQPSaHxV1R7p5iUl/HsEeTmh34F0Yi3O0AUG
dQLFJCqIVzDH8hBv+vwEkut9lSWTBQ4oktyvOtFsg5OabzC/UwKWVvq5Olag76AK1j64xAtmpalX
fCTAFYiMoQw1GnHhOfSZknhS9eR92J6xIHBSAk5VUwEwPv7gA3Q2F6vIsvArUSiUehwW14DNsEvt
sWfdP3eWvLOkYzNcYUYWzTmyvQgDjPwZgl4aomoA6elzsLfvqO7IGZFCyh0rWTLpXE/faRqFiCVQ
fdY1jtcITiSnFN1Kt0xxRRvnrx6rNcx7MkPDg5QIVSKfHVQLh5NNITPjpuSA/5ThKV8nWWdl8ft2
UsfvB+8y10oU5KP6alrIKn7e7cvX++kBfB5aq8MDJ90469piqFDxdA89X24y9vTJg3cYi7+mYEIF
PzFOzcOr5orT1djVH6/pwdUgX4rxSanj9SLzQZdXB8EiCE7b0GlJj1t/CL+uYtKMR+1Z1UKaR/FF
qqUXpzgNr9U9rzM1qBfWjQq38ERhJYufhPaKj6oFc+IdlSGgiiuab7D0bzmVTYav7pt+STrBOaSN
Ir7BmpDyk3ei0rreGtHbPS3FPgKnP5RLV8IfHBcQzvVFKLmMep/cenLjggkVguK8B/bWrYYfXJSu
E22QGHKNHz737avlhK6ChhARVsr4ypjKXgPpOdqsVohojmExZyzIJ/5GIi5cM452K1j1C9v3IMZy
9MB/GSSPRYw/Usve4BqicwYKryIl2K81vNEI+m2cnS3Oh0u7FmPCL6Qnh4CNnNt8EoeJhDKmeLQg
8Akkh7YRfHS23gUbu5paEiRvGo7YS3hFJxewOcS8z3FRQJ49E96UMHA9wVfQ3djmIpfDpxyZ7Agf
HDhXVHVQjLFCIm17Yov3z/WlozSAEWHwDjBCJwFOvfTcd9euDmCMpc9HY9tdA4UpHdJirsUDpflU
fOedW0A+hNh6TPojgeq61QiDk7Wqj4uMkBUHvdhmqyhSEsg5dYtl1IXQEV/NMS7q02OLeBfSnt1W
bWneUGXGgn9KD5ikVY/UoNAUs+/yb95jD+paQ3xok4pINc+aklk/guCrsdOh8oRins59TTRcYsbY
QS3w1AyTB1KBWsoNu5vzpzNw+iKahqiEWLx/hic2eRcZ7fO29TZ40P5teW83kjGRyf0ks95bFFrG
nymz01itgL+yQSHItGSm1ZbBB8Hlx7iCVPe7EbKcuMt37ULipRos4CoKjuRXGtm3Op4HFOKW4Njh
AwlpNNQAc4ZcCTyySWUTrv/eBYIy97aIIkbXVEftVgwl1xfINW3Hgegdf0HeslGqbA64oCt06N/Q
xp7Drkth3nYMZqieK1yJPs04RXkDrpG2vKN/7RBrNlS9apMEmK3K0r7075TGwvTc2/oInfruE8AC
rkS8IlXY9I8qSrDQhnu+CJOtG8l2NwuvoYDuY0Hco0GJK2Wto6WRtm80z07nwuDYXNo9pVRX1T3i
8tsm+nlGExOkimwYZvSGspzoX5AWKF+8el4KNTxeNyaY+BJIVtztobxlMcYR1hf7/9+OiZMmxkoj
tqiqw2foAnBIebckLyZLKsesEpnjB7u7RXIQihW6KSQMmADOSGUN+Y/JCz7w/3BOkj7Kc5u1SidF
UUhkFSQQt2jWr/aoDyWsm6M2rLdWNd4ZP0xeGxhjrVD5mSWMu7nPbEvTMeQBSR1WxzSskUPX7ewK
uMnywcdnEdD1iHdcsAVWgBFeARnVgZ9RoGCK6IEl2bINdyH9fXclJG2Get3zYu+io6lvsXp6tACP
iaXmxLt9AYlnLWP1QCBxCadamOEli0Lyj6pEXlF+6kSoFZZnAk4uPF6JhR/B+SBeYuAizhOtzhyM
rN2IKErqLVjKLVrSJOu0DbfSplOgX/Q9FhKZBnUzFMxOujOq+M8cFaZFnfjPdVmEri+vRlM66kWW
1N9lH1RLenp3Wt7xxB63z7xYnuMUUKmttffZQSdLzTAufifM6tjAckqybadsoNtpV7YZyHatwSc4
PQsj5UwMbCToDp2EJD/XR2XJnn2R2m8UVHI/W0gFuGS0RtXXl47xRsQtFndpQLzUEjjLckqB2a2f
UIVAKIrXa8VdTQ+GOZ7v7ZgDP3ucswNViT3en0PZZR2XgjOjesFTmDEvovRdtODux99wu5KfpMPh
NdVSj3C5TljO9d+DkpCO3wx2yz2T21USahX/X9Czvo4FI/YwvpsvACed/FOaNRv/XiyCbkVMxGP7
MRjR8IR1z7xAbx39o26Mlu6e6n1sUBTUOBKgCRWOskCG4lBAspczCRL3udxAT/ZYFLBQsM7N4dkA
pyNu4H5s3MlS/01jcKEfbiuoFp9ODyzaSm4QqVl8XLR2HgEY49vZFCYxFYG5Gm6YQ3oOTbbbgTWm
5SEgT7wvN1zP7zZr5yUReE0ik5aZ6apIYFJrHzg5qHH93A7jfJvGm1TorR/VQA6xyUwUMbBffp0J
sZynkJa7YCR2EDJ8vOXQPvAY4hchrh1BrHEUCIR7bHkCKm2BPPXGI40WSYslBcdkZbLYZUjcgXpi
U/iz8FENPv3fEcsPLWhOUUEiE8x1/KcRcVIuOZ4+W1lIYt95Uq6FN8OorhmLiAwNwqGzVX8YS3Ei
V0S2x0H5NEnYas2adfoTrrvc2dNi4b/Fnc++71VUcVkHowQWMSjN4Rn8cgmWQkzWVph+LlWIroIt
U/XPlSRBWkDJdJGqhBU87ofcwe+RsZHx301dnFFJjpZiN5dsDzNc/MnKt+uAQ5m3ifQEB669ArHx
hKc8Ml93A5LVhwRAxola52h0pTi22sXtBLStawiVTW4dJIDRHdHcrURPHvlmDDKBQjqJTlXSXU8U
nhuNYzlFufgSA6OlHKZKhTnXTIOx3DjTDsSNgqta0cbLQRPuo8J8HDVMTE6ktc4pc1kOgle1CMcO
zyp9z18/OfIyP2u8toJekm3ernBMAEW+4/TOQRtcc/UJYxi87y6kwQzhtHpzS9VYf0OHEHdKk0rh
63RZk2w4Ov1KslunYnM/lJuOkLp7mT5EMDPOtUFvea7xwcfgik5LA0dA2hd2Y9ul1fbrnEtZCOjS
V+RBxUWZZSfB0U9alVtQKMX7FLfwsvoC+ux3bpvlxGWnzgNmgkxWRjNUKAwHf03H/5Axp6+ug/hx
AwdPl8qGwdufzY0QV9c+ElBfN8XQja4E6rPM0bm12k9KDmglLCqdVyu4/hB7T9nj/5yfdcp825vQ
+9dTdyzzyB0VhgDw4ttyKh/dsDjQNbWk3QUSyrQTnNvS9cyFKw/TxbS22tFknuB5R1jG+kaaRwAk
Izfj1OpS6g+SmTsYhdDtj4fEEY7PB6Pw/mFXTeliLhq4zS5/BHPLiI9QuTpbS6Cq5ce+h57s/vvJ
BTXJCd3Xtbf0pXuEJhPEJemPRRUP4ooQE0j6hctaZCil2xucLibbLntQPHGljGKszcJgm7wliaqU
FW23X2GHJbTQRqBvDTTCtTi9s4dO4+nQPm8kErG7UODrmunM3oWjN3lfxehPkWv7SvdgktKDeyqB
QSrfOMj2ZT2kOnxey7bVyfQQpNSbh3WUPVoBJwRbblNaNXY5YmHwi6OMR0ja9VhgVAGFA5+CgW22
Zjjq5A6f+uI0c2d1YzanshFPq9uMf3UrXSm5T88Bfo7N81K2GyKe5MvUwC/MYTbymxR7fGxKoM1S
AjFXV6ZnKmMH3+RTE2rQhU/uHukXkk+NIYOoDehDGNpyeissy744VSoEPfm3adfLGKqnh2IJGEey
+MFspAYIdrzHh+ARcQNG3hqxSldLfvGGa6hLQLPPWwkOPPoxBE74HV0u3WOVct5nt/VyfLpGHyIn
xQ7Rx2JmFZ4StAZwhrWtzphKXkbAP4X6tSZQNP3tOomZeKUENOVAa3+hWstPnIlH7+3nXgBVgYUU
GB+ZrqyLycV9pjQNjDys2QJlXq95eyyTACq/bHy7ImFYgzVVPng9GVOxeX2xA2MQxl0cKomdYnPm
8WohuswwpcCh1SUQX9hrYOrOaOe2999KHL3owp1cRr1ixcQMWTlLDwt908YhNI5LolE4i8NnuEiN
aI5/ztugS83JPJ53J1tuijCz7kJjZEQDJ/0DD+tnBXFkSkNYVprfMKqp6L8/uN6BGNmhnmdqS2QP
zH5O+jXMuCzeOq2kcYDggIpVu4K1u6m+oNSL+ZmzaTP/BP/tA8e+l3/e1tB3WYKdfYuUK7kb62X9
bEXnSxtwjQZvsjYH0s/RsVqXqjbDlD9Kf6KZn5IA4kO/KM55hWRZcEpohlpcoJ1TfqpzoGm7zmp7
V+PkHnPuhLoFEAfQR04JDtWcV8NpDBVg67iyl5wQmgWeOiJpt/PxPof0GPKj38pBPXhL0A5wG7Yg
N0mvZxEd/CEgeEXt6ArppvKxGTASpAZvZaSE8oZoYKvuQC4yEjwx1bwT7ybKi9qhBqvbUG974/Ff
G41DT1pbmoZQ5C/hQHWDUjRmunHWhD6AFiE5eqjFb3ag6JOTlPpncnUElvjXIYl/dEncZN2VsGR/
MVCwd/Cq1Cnk6opLzvBLCcRB/yu2c29RZzZmlPA9P51DGA9fipAQ0ppSHx55dg6c2P8SaJu5X5Gy
1+utTmKu+rJkFtZthnIoP5XCtfZoEi+ud1oeeuOpvlJby9FE3qL/iIKqy0AfnYB/V9/fGTfVUnLm
KGo5NtCSPB8b9vyMf01uK2ueWh3YbX1BJ2wUSB0qTnXGmIPSM24AA4rt9LM4BZ3IRBuTuEO4kF5o
+HJ+YAsz8e/+GLtzIax64CHmvTcllaYTCUgZQwnFbvPJk6kXaJsv6r4AJsndKBQZWSgHTcwrSBke
/lzxc1K9EGj9zFBaaXAdG+ajtLCq/Hx2ZuG7EpATue8fJIQuSNMsNsQ6sXvqwkY3FyzKAWhU/McJ
OmGdH/WgTy+VY5Yt7pxaPIbMNmNm+kb/hzKu2wOn9231zJgzxxKnJxd9KJQEGewnMxEiLd739MkX
KbPOwjzpDbqlx4S2B7WVwczXuk8PrzbWV3H6DSViKLfrHUsEv7QydOUFBKNczqJiU1HvDSYB9twV
WFubywXv2+4/OLNceUjkvlWUnOtoX2oFduJ5McxK7B28q6yAFTQ3QfRz5M30UOO50HjCtetskPGW
mfxtje28a8wPMMikM3bpPIFAhr76L82qqYAZVHYpH5gV4lRF4Z0KjdBL8Rz/3HxOVZgkCeebe8F7
Ay0/FubuBKhq4MwoINVTEj8XVQ7kq0E0H+01pD0rHbyq/uTPQUp1Wtw2yLCl7yGUSSOn9Fm/rGj1
5fZ5b8b35TyHleALCmDnAjSHwcL954MUmd7nbQv9LeXZ334BAf0mnUWVdalLS4/cJvOm14faPwwA
UcKbJ3jiKOpmM7t1wnf/g6zGcve7X59cs8wHgKe5f4Wd13U93flaP6u7ofqAKmSpg/UUVDCzTaMt
8uhrOJAJH72IYkCQt1NbRQkBq3hUXLIk90/n/GYx1OERxgDpG+H8Wg+npulRwhl2358HGn7fSGp0
UtcDoPB2LkY86otbmpYArWART8yMJjMWmqB13yNZ+KVq72v1rSM1bmiXsYd+sUx9pwrn7Q+6v1zk
0SYMxyN36e4T8Z+ybG/qIO3FMSrMaohffdUXa36OAdtEylIHpqLiWH9MdQ8QLRq+NaqWpCSCiioa
0tXwznaEziO3LH4fs5ntBQCFuuVUA7pAa9pOupkCLricSn/yD5VQ7ega8bVkRl7BCJEQUrlze52p
cd9CJSCOa/0i8iQER/4eKeJuAJVoft3z/ZxzfUxUn+jFhQsLCbIaSyxDQl2z2xG2/kavNwMoIAnw
iCRqaQZEUzo8AJ0hvUUX2bRhJuXGLveGE2bDl9zPKyKAsv7tXmgDVrx083B/Zj8Xvbubh+nEhcvU
dQqST8qtVqCKnJ43QkKHfIfFpd+Xu307mzXkqPagTClT0NNE3+3HBeGVX7hUnvq8/+LLuW9PXm3W
67qVjUppw6kGRTxs5n0XwKlgiuG4mBJ3xK2ARwY/0tx+HbPlPL+3NGv6V+1KjZgoQ7OrNy+IRL/v
HD5eh8+YrbnOBQEH5pEvtVmw61kenoOV8I0mqpl/FKl8Gp+YjFT6QD2nraLhJFwAA+hFQnbEw6uZ
egoal/XHlds7ZEFqSbYYCvgtybklRSn0dOOzoiQ9hoz+TBnMsE7DUfjnn8ikABl50ACv1LoOpMzR
gChVzW9mx1gY1AB5FAnc74sx91xn6DQFGLInniYcCBmCBwUfVTBFwzKLG3koCR7qOzYxJ6eKz3H9
hu0laPk0NUcgVbxbYFSVuaTHL0qvnV3kXKea9XudYgvH8cMMTe9FIQfUkkKOvaD2BZw9AybI/9Kx
8E3VolYfv25Om95mJr5UMUnHRt4HRjazoYQhP3Ap9v4BFfkUvStjK8hJPaofupWxPfvXQze4BDs9
PE2UuAWEupl/UeoyXObPwdQVfQLV9fjq7axHRfzUsoKwfb68PIUOWC+U0RwcoThi+49UVCW0Z1Lm
7PKgw82oQBFoUoEPull/P+vhBOyh8UIsucCFaqSmeOX8hm8TQtvLKbxFCV/23D83Wu4ai5VsHHez
Mhqpb9DNQrZQQuhqbLhhuToOhPTOyRZL92bcBU6vBKSU78TwkdEBAdYDDbaf9t8W4deX6U110wB6
bkbW99e7q46sJlXzUQULByZxk5ucw0+pdx5QiY2K6qDeZon2BHHWqDuC4TWemsQdPjFoINuwSmVF
lSY1yWjtaWH9Xo3dG3Ex6BsNBg4x0heJcOZoWf1P2qMaApY3WN6dgOEwFYgY7Dqbd49eeNAlCvj7
Yo/JkMA8OL9vVysGroXU29pF0qbkHJjcMSAVuSyFYm5PkotlwRwGqsBDjndUqBHVSfRuZJ8vIFhE
ve2DQco4w4ygZUYNfIWKK2WFU+X0FGuMtloeIdi55b7uvbCCFyir+XgwQagQlX24q6r1Yo5/qRr9
uIGhsx38jwhlAI9hgWB0w3GRVzK2qZdc0M2EvJVv8dPB4LPeEKo0m5rcMO6Te8GMomE6A77ouMrX
7bvdOep1YxXlYHktDluiyrWCKGRLSKm9yfcUxBB1bWip/xui8neCefmA3X/+T3glJY5mB8F+CvY5
axuetr1Zx7+pPaP3JRQ22a61ILJd5UtmXZIbE2/ovT/KhPkejv1wl4aLwWc2XMiTSICRQPP6kVVZ
l65C+fFVm/kgdj3kFOlCO5kQVla+zTnGZ4ChEWTGuEvFUZYqqyzxcDd0MN78ayRqC9HkBb27ljgd
N6hoD3xrQKf7zceJC0x2Qoggk0XIqa6PW+wZBKUw12y0CJaJIe4FZYC8phFO1ExgLR4e6f+l1fSj
O7KyBWYUHe0cnORjVYdOOoAE26yqqrDAvBI8dG3QYFjr/QE04Wikmgzw0qcWbJ7ret+FLDQjZz9Z
nb02K4+m49fCK3z0/2fvC4zlYc/HcJsa0h3neM4gsNube/jlExX/uHNo/1FcUbJiRu6vA0+BM6nQ
Bf9DpGEK+q6qTYVbifoLSvEQWCrI+2wjNOpQYYKOvt153C+1NwWk44ziOE4DMc96aW92vpP5RhDe
3MLmzdvlepZDSsfKhX81vuUMJoAeLuPT93lzpMYnzuTi6XQb/J05+eqaVN03fBiEstk5Bg7MR45Z
qSczZ83QJ88tvTbMWHC0x2c/7BMxn/rsv6XOM+xhnS6TjS0na8WilW6xz0ECTFprb7xV/XxLBW//
r+jILlf11csVmLvyir+4IlchxOP60QZFkp24jxexxL1hem4mSY6BQKt5dty+2uAEO1FvSN4/twCc
rFS+U5dddxE6SnYrKi1NKefthOiWx/uF7ONPX0MmyrJXEiZvmH6DQRGhqyAuXH0nvrOLFO7ksmul
2z8Wi0mxzM2brHeeTHlJp/xhysY1qDU0I7OTQMN8dNoPA+q05EE0mb5hBGphUp18o2RwBtQgGUjd
5JRFwtseATOLRvZK0/44fVfeIfnr03hAmHxp23YeUaMDWPsq6X803hzYipci3HHR4owCmvHkzyCz
yGPV2sm6dK+kXNd0fpkBgmltQG8lbOZghzzNmEOg8kZPxwi0bK1bKGtAfImCMdmC25PxfkVPrAiX
kUe+5CHoQ3vPjalmQwZInUQZBYqZljFfs0te/LjSMnjZ+Rq8d36/8UtLyfiVMWmxHJ4AuqWipyC1
t2Xyl6gXPN3t+rgsEy99U75+N43MbwOjhmwkymMK2qdtPnpPs3jioQjQukVYUxjFnIBBp04fiOGp
WO1s6eLynvkbf8gWyvNvn7pOdomrA+Do1sm/6GTDWp8wjvLxzCQO1TdHNcNbvQmFWcpBGWiaGlFK
5uebR5p5GR+EXlQHTzTdjscOyPbnI1NBZIl09+w4q+A4+liNoId5rmfD9y9z7xIi8LXiGcfZCVkx
4MwW4bfTOM4A1HAf178e211Xwl/M5/48lIetGGg1//wqcnvDt0kIFb8MlKmBuZYHOsBDmcYFs9uY
O850IRrCqKp/xK7eMxoP+i1oLweXN1C2eC9/pVxAKXo56LOHTTIULlIENZzEVPsDxPtUD5pGZ3hq
bhaMGC0iud6AYHba7mOkftnxdw5ObXjJN7upw74yre090vZkmUJUG6vvjL8i2fj8moT11u7Md1E0
/nvIXrVyqfN46S5pbTz7BhPoncMefrjwvmUwzFWpw4DW6ZrtCJISvvrye2ydbntXOA6ChejkUpc4
BNYLLBvooOIQ+9SD3MF8vsHyLDwaRka6XcC+qeiWT8WiUwqmeieju5nVTcVZtB8FXH7fzxvN0nrr
TNsJIjRF1lk8E7S6JV6edNosTBL5KNke9AGAVuhIeTFtlf6oVPoNj4/EsGzDMHM4tbHw5EXbA7v7
mSGKSSKxGX+oW9IuQ0EtPflv/8rOWz9Iym2cU0oL2k2QZKwroqv4ad7IrEg/gs8dvKJSvmBvMHn7
N8tt8tnceyMDmgYSX5qNHVbtdo7CbXbfG8lupuUWqWaownbqbHtr4IYaGYavRYKoj78D53mhjmWV
pxRJJPIbL2drQapIYKcXnQB263mtkx7nxGyEJNJAUuOlQBg3xq8H46wJa0GA7n/fQSUQYEYP6lfl
627k70bSSO+PhqqT1x9vfCiJVGI0VV5pAAsbHPd2c0JbxJ79KqQBCliP8AtB2OQbCZcQ35r9wAvK
CsRBEkiGeJgAsu5Ie11hCPtGsBnoBT7zcD46j26R4rRMioVIQUbTauNgsYQq+cQ5fvul8ent0IXd
xSdaQnQGnrWgqk9WfGpMxJkbCkElHysuhrWF1i+Rtkj19xUdycwuAHTqESatsbVY2uvf9vjjMbPv
GuDYe8NK0NO9ZLhQg7+78+5M72ZDmwCxc/KYK3EuBy01uCujJbGllW7bY6DF5WS64Ksym4HuNzzL
HmisJz38UMcV6/Q419ePdEjivuHtzuE5u/ucqjOWm+UYkZFLJBsX2qFf7lroDefnimGNPiG4rYKL
9E0F/6Y7x6S458b0iro/mlFBEFDNSWHaMW10VocyTHNBbV33YglulIPuaacU0MoMc7Bit372cAxy
e3JpCseg/i83re61etOuJwjAJ/vzNzvdqXs9g+ibn2pe4CR5fOp1x2iOG9ksjclXN0Pfqd0644oX
tB3vW7g3M+XtGu++zePl+T8OwaA+U3jIUQR0aSsoAynzbDc0M6N77Ps9W+u1SIGRMWUW4be09LCj
hPZmUQgu4K0JiY/5kQWIYIeRl6h4TKtNis2N7uN8M+f7vepEUulxobhAeifS638y+WfNVfeUsSE5
IsDAlm5cu/qmAylOAzZubuOcc0BN8nRgkcfqVXGvRPfJKvHZMnkZqG3voeG3X6VEU6l20W3Hc+F/
vVtmM51kr53kR/VA3TTy0qtobcVvb4ZaPV/FksWqvCVMGW1Vpj6+Q+fTGbjc7RXcpe/fO5QHrnog
pBb/O8vtG9SKFyufgNdhKzpy3icM2ZiL/v6cK7GBNTx23x8mEnYwvSeR2TAcVfJHOEAookUFUAdb
c//9TvUeiv/MULF2JAD6oel+CvCtQvVoo5bvKyRW86IO0pmS4JwMSkGN5wPQmeg+xQnewCps9FHG
JW7AvsnF30ZEx802ez5OtLozTAzUNToDa7dnZU5AhX+1xpDRabKKUmSDXvTm2v8DsJNLJR7GJzya
8eIDK7ELryHatYOi+R0DQf4nhMbyRfMWK3ZvxsETA+uEJdMIZ4ngfCEAjNef+pijMtkEZe8EDRQW
C26sVkq4NQ1ethZNrrF/dEpy8WhLYKS1kcCA5H0sXE/dGwwHPtzcHDVtxgR7q+gS+3YoaBaNw8zj
D0d98PfyldtTXB4rtBBoKcpSYxWQnMwkSsEfzZ8X/efGJ10cZmyJ12RePBtJfBjdqfAnTCrYR8gV
mKPL6A8TaUgvYo7u6Czko+/LFf3x/7I2h3wchu8HtpziyhP00C0I+4sZJiI275d86OUQfgejDb4C
nX68iHYm1RbMmL7vFungktW6QyKXDp3usaxSTwNSK7eAo/hrIxbXmODXJxOr49pVE7bRFS0joRI5
ozLMCN1y/XzJLD4M1CRRr0ck7p9QPctwa5/OSolenwpyzXBDccM6FnNFKejQwb7AvJC7JrQXU9eb
pdRhkreG/ZOvFNbdI40L7E8iVwZrVn1ACPx47VVgyRYs1nGuKzYBrjiFT/wr99yRishZ5L75bt4y
+L9OVj/5Zyf+eSltMhnzNStsAyMVNUzd7cVaFhvPyFMf694R7szgIJRRuZB3ei8+Nv1QAgNb0htM
u3YsgO/KlJnB7Czgj9KCzU3Qjx2q0Vy4+IOk3W3fyubKtwLLj00rbqcEok2ZOik2bOQymXlG2yCH
g+ORq3Dta3LjTW54acVUlKWSwhJyYXJx70WxJVpPs2wsHVUhw0KJN89oY+akW1JIX8RX1QQEpUW0
L79nu0vCKv+LPy6Cf/Sf7ah/QjWnKwldBW0tW7GDyeJbQ1hey9KvZbOpsR6WWi3a3JNkaaVy+6S1
b/B6XT+55xRY66/yW2eJpf/ds+x4cUi/jX1SYuU2tMY7NW34lbP0QJxjQDN8NkaBCFszuBorxCpM
6n9DhurgQrrtm3Uf0U0Jpj2GS3VFJnYAZ/prBO1kACInvXbbc69Cm+pJLVEnX7IEphu6LKc9fnoA
jHJaeTfO5uatxRhUkEWdyLztnqckwyVrsUqXhoixwNTf1dX6OWDElnfCm/1/c0sb56EjygoQ05XL
Zet6ZhSb9GK7jt8Z68CF6hZgFQuZQgfZHtGbiyiztGRHsZjbQI8RO/45FXL8RlwnKig8z43ejFcd
b7xGfGDIA1zs+P3CcIW5HnY8mktflGFS5VyMxGhBnnGaf9pcEpT4LVq3nT9bZVUKzZ6zHayoKH65
foACALvo12OB7igYqrD8rzTXDzhezlAYzMqMxPqsG49N7vRUMdFwJQuRrqQDZo6VfQg3v7jfaRkr
hoxM662Vq8ipZPiQvg2ozrLDuwczLRppHphDs8vaqlDJmROpchVWpsFFVZYeGGA9ZXsnluKKVip6
HhLAEYmhBPzcaH8zPH/wozX6FvGPVO7TIBEbw5UqdouxFIZByU21z1lqve/x0GawqoX4aDXg0THh
e5iNUgC6yyMtlcV7iK1XzTPEIkSfCNv8lxCSfabicwzButC/Yc1niHQT8VhHsrDRpu/0NnKV8JhU
zPAC0xp0cBmurp4ntqEXZnnDzybW4WgPdokeHuSI9JBiIHARa+Q8Wp5tQWCCMDJ8gw/Uj3oDhvaT
78P6GrnkK4123rtYmAOSFXkRxqW0WPl5hkR40Wtglfd1InjU1d1ymLAIR0Q+H17QKu/OfS6WrubF
759HcwOC95h2fsQcYHgwwwrSksd1a9n3ldaWn+m2hAva29WaLyl0vnfQMGM7IoguybQacFafK5Mi
/FKQaNIu6cpgnQUnxiXqXOuA4RYFDErB6+G884PTzaPnnpBhXmmXf9k9oCNRYv3Pfo5oRYXytLFy
SajgtOz6fvDL0yx9cFHv7vxqZLHcODpq/TL2bUHe9wbUPxjS40w0Me/7VoVR7Ubn1v947q3azYvQ
jOIppgiD3AmbKad04GEuM+hts4qoJY4PJNZSkdDykEohSwZl+SfeTiWSqAX3P2bxeIfh2+gro1kS
6VLW7ggfVqRQJpo7AO+JbMx0E/YSd0NGx8iQy5N2AeSFKPOB/v4XAuO55wU0hNQeTA0JsgERnE7x
PuN2EurwZpUQcUTO6eiH3A5DW7SBylSnkZHFIw5f2r/oBooHQCeBJmZetwbec8UFs7TbzzGJMKgQ
JsMFF6Ak+RWzMKUVQWWgAA+cFdbisOurdej84M9kdJWq+H+OYd0wYmOMZuMHJc0vaV55vsNIfbf2
Ow6NPeHT+mvGkB8ckKmYNu1not+sdiz4EBMSQIrEAajPhVb2vP20xloHMGbiGYUxsq+9cSAqhaNn
zhF2kuKYr12FyBI8/s9dncgUZaI1FkTULBuE6Pk2Ngm7hZnDlEUFY6fkbKMyztgp5SY5GxbrKnlk
XnHWlGlh4auNj4qU2Rm6H7CixmyZM7OxN8dWy9TGN1thiUsEVbJ6bhUcjor23F2h1DflR1cyBVS6
NSbIg9KKUHkQx+sdoRHb7Vud95MNWqaJznw/5HQY42vg5eTeFV2zSbwZ+zslYlX47BC/NLNP2UQh
j6i87aR5y7hFZuSzj9bgPVIRq7pkkjzsL+XV0ogDnVbEeVRF5b5CK4uF7kS78my5yV8+3ryFwmzZ
rLRA7BzTS3Cpt2m6kVeX6gbFS/o61olvidpOUM2rFEiaUt/jVfBHkO3LtjEPuOblY/vVBZ9LUGPf
xVvbcn/j+uxdV33VqhJUSxsgMSgxt5GO1f5htORcoHRRfDvV2dX3PdiX+m9KiQO9nS6Cl3eSSoD4
2Nc2O4LdVqpyTVWVQyP+4EWqPk1JGp1b+hRylQTPj/jK3F9tl/Z27akPiEefk7BKaC1pqgRCCKKJ
4AUOUiEn2+6PEyBi5LLo81eOAHeLZVTK9uAxI4rQeTSnOFEBhbWLDs/D/JzzXan/N44sP9oHGNiP
O1R41lL9B8qllnVLXTUlmekwmhA2dHwW+zGghqa5SMtZ1kelAyH+UXzDWkPQnrmDYCwtzXs8zsdO
Q6lOaCmvPE4Vi+h/7PXEt70Pc1FEj5scEsPhXEMuA9ZKPRkJN1/x4XKLZU/KVRqlu4hyEYuVisiz
xUJ/VR3Ktgq6cwWXp17+v7/vHPANeI6obv+c3syhZaAO4jAzcfNv158zwNCiTWYMOzXaeZOS7/2/
Of9dRm/LE+1t45idSxi1swum2XiBxflaJH7WFsGnTWEMDmhGc8ZrDg8w6ZxlaxCHt2gJg7DIkVRM
TN+7c7dB0yITZkgybyZaDMzCZ+K0aSnZFzREnRu8CRW0VazsfJm2MO76YoUx45nvbggQ4M2+Q1LI
FDdQZecZk8Awn5XLO3EgzDGrsYF11iu2T0njbJJyAM3wzvaRSh7PTYQdDoIDfdEMCue2iMePF1zj
PEg5pMOgBUlPpybhp0w9kYVoLGeiS7U1MJBDctOVBnq0IRkaW40aXm5P8b8XqvskOs7nksw4kQGk
ppXaFYMHEfI58FspaRA//HJ/0qYazC3LGPckOIxid0j8i7XznkQ1gurMEYF287uO8k0/bJjnKmTK
0PIIHBytH8MuNMVyIgIC/M3BytAnIobMcoY8uqe8okfArrF2pZcSzuQOJHEiJfY4pYGfhH4DFYxL
94sg2FrYeJK4DAaQhra5o3ivWKPIoytN6Z1shcoO4Xm5jgb7SRqOxVDRnn6mBgiBHjjpb4W889LU
kXlayjIhiNBX/RluviTP+EQsBHEqpBKpfUBhiouBtWaDjHtkp1PQw/sXmxeMQzJtEr30VBSxhRjr
EhDmWvqXSgwazbriLuuIOeQKdCECxL0FxTkQ8IUL9vhwOs+OQv5PUM4MD+IzQCspMdvknJRuSmGa
hFxEePqEpkY/RutO1vvUIF9plB2UVMPMWw5AVjP2ji9FkQ8FsymjZvwEZ54TD5Pgtv4jovR0dL0F
NUoNgm+W6nVHUP0EUufoNhRM+n6ScJa/9WU9lC4ef/2bxMAskPPvAHQdhEthetj0qzzinMyzihmO
x6kDVn/CV+M7Uead8v3AfpiENEqJAXjED8xTtunSs5+wmcMdfLbGL2FIEG+gjPXl9LwAF3qYgGjE
lWYRtOC+2BlgP7CtsP+P1yr1OyYAElr74gyQOAbSRfOZIKkvEZoGFS+lWDWd/eBxgqo9IMiuUopM
LZqiL8Myhr8tiX7AhQ1ArZE6n5PURYpq0/3lb48MVwf+Cs8KELOTnMAvxYcSBJh+zrr4RkczuUsn
HODKNdBpV/k3ZlSVxFx0gE5/XeACFbSS04Hjm/+cNqzKEWTkl8/X7/ITwe5+w8EwONFfqJE9NRgz
RPT5OsCitSm/rH/pb2tyrDSYGVqNmhPxPUvGDznuVJV6DpFbqzrDSVy2h6cF3nrBbqu3WwdW2H5U
r8KBLwnoycDGcB15/qGAqMeOTF3MvPZlxum6uotdWPQk/BvehfKs8voIAnrs5gBZCxYt7eNNiIHk
OwzHqoxySSs55KyFP7xfDlimEjjUVgOKdGwV3dfe9FPXHzFI0oD/J53K0Xn0g1wCeNIw4hoW11Ru
7J2kpkGnzX3UruE2jKAy+mdeFfNMROoKjbNSVXp9ex8xcXDB4H2rEVV517BoJY+SqtnAcog+KU85
8Tcs3D8eZhiQtfV3zMwxvMEcWKsg8QDqtvrr06lUSdY9yvEjbitCNaAJaw3gZdlj9om81hJg51El
vz/zrVyYVLzxT3UIFGJ8pusMD1iMJ8quKM8CK4SWM5ihIwQB7ThmrvF1aXCAJLvDeBDooEQ36C8s
J1bgPdxkCYoTmw31zM6lcMm1q9jtSidhKKv4bBLBQVpOEUm58hdZDGjENUMRJyw4RgSS4JguIyd3
Tq9XyPq2oO1Or8zd97Rpgsv95wUFT059lj6DuEMuZ6KUy2wSfZbYOrAZvDB/c1A1vEF0dtTf9iT3
smXdcOu6QVWK8YJgqKQZtM1actmj6dyo6ZIO8gy7JY10bxr3eXeQwmDsG2mCNlcx9+Eq2NI+xLni
iPNdABkvestpSTxYZtMUCc11KsClEXbJamMs9S/+xgY7Zj193Jv8KITAByd4nMHHJRd5Zd97KO3+
h3QjDUu36Nz02ZABfKyxFXcML/UiyGJnOdnNePSGLgzxLdOdJqpL8OcahKu8WKNnKghP7Jngeve1
xXP8oetZ1g5RCmQyA4NruR1JNHhl2g59ZhSnzFGvSSDe7N6m6lkvvlVSZvC6PZiRxKhwRhTC+jy0
gZ98DhElxwZERSXDVUW+CtiuFnukjKMkm1ctO16EhAiBrpH4hEooqd5QKcucXbYOLzL1La4G5QZP
E1q9i41Kgve5LziNZu18zuqu8ny1sJ8Z+vnHJtWCElYImRVtKG8xZO86BdLhnOyGXkvNk1GIJTp0
S3TN9nqmhvxc17wttm6NbfLIX2XlJ4+AuK2pxfN4V/gLZ+xjoOO97QmwZsRvWWeCwb7/qiGFc9lw
qjPOvK7q+WVvO4IyMCB7M6GgyXCmiTWgT2FpY4n6/WX2UDI2sUEZHZqT5UXHe1/gzOnpMZymEobe
vF+7wxpDu2i/okJ47zVkFGLj/8J4ZA3j7j2ipwKWpg5Z01rv6eNPcUFuEM4ru0NWzFGfYFIM+Fey
ecmYVt4BFttWH5j4edJK3uMFAcuCKzXKZXsbSUKxB2MqHeYUwwEiUGeILtuTiTzCRtnnieYWdaZq
St1twOl6/HRWnHFsILT0f5zvKPq58HAi8MITMcocxPoBXQaH6fouhWI+NkvP+MZG7B4YjhdMLwfp
fSWZOx/uOJ1EdnfVPBCHqRjvBJwXwyXn9PMBQi6SravnIURF6ut0yOjWtqqDzUKFv8hvnL0Oy4qD
26ls3FIHbAOtk3QeDieycJspuGzczvuNkWX7OamwGqFo6XSHJOYxKkDOWCpQWG+RTEHPSxlaLNP4
1N+nKX6mNgJLTk/4X1lwJIPvDp89tEwXn3nQK87wAKY+TE7XoLmclTIukDUR5IEGG3v2QXi/r++n
ugv/Rb8CPnaCNgJ+VphY+X7E+Zj4F0rPFTo/2gdxXQzSUdSEO8oXDatKcbxUO6myWK2/bBta0BfE
f4nz6OO2IWrIvo7XnB7CU7QRWjsMIKV2FGA+yznb2aWQbcWnorXavQP9TQIryA8Jr8wqyzUDHGFp
VtLnLhJ2rl1pekYA6dQu0wRpNQZPEpqcC/37a4r6e2D9uQIInuvow+u2hw1HsBbDyUeAjd4fzE2i
b+9NlVcEAI6SiSPvobtnzFw8JWCcdmuzSlo7ETaJ7a6+PJxSjS1HL6ZiSGLeszvVaCdC6+kCEBEE
su9lzFk0imMoZx4Pp30/HFjhekAsxkqUZOiOkIja0+JMvIOGNOnl4ulduNZQNSBsi0UHH3qmLc3c
lKXHVacFKM83w7Nwg/nsHF8aG685aG2TrOQ+5pb+9FxHID6RJmp0IoFbtXuS1P3ShzXyuIn80i/d
KI9Aeenork6DBJsw/t4S8FefcapO7aj69LY19bNkEfH08hTRCcT7Nrpbi0xbarJZbIfvGrVT9kxs
RiskProhFtCDQCsdxKGHEnm9dzIfEOifRZkblLc1/5+Qgphya1t8i8p8u2n/zpPRrUUAfMFrINwm
FKIa5sG4KWXEi6qD/PLdFyEcsZcPbUnUt2I9Jw3yR/w2wGkKLu/g/jZj4aalGuzhdVCFCa0IDTfe
DBii+yTW4CBf6kCs+y6bW8bzX114AQVlJMSR8Nw/sasWfxHDTf7z+rbkUr+mFF9tI1iYcA+k2F4l
idDVBUd4NyAYDGz5s2L6cx+nh/YugkES8ZzfimSJwU60UlKv9PMiIQ7JkRKKuTy2W8SRK2JGBy7j
KiiXw/UEkWcQJLWO0bylDIAJ487auEDeacHX5TXjVDIScWp58DLUkXD/YKceDW8Y90NxQtPlAed4
1Dvvtnq7uI57bBvaZbOnwgsAguAVKhuj5zr0DqLGdlOsapmJybbGWBT0nZQ2CludSBKH8T2k59he
0BNlF4iF+E5nHQRdHdgJzQ/j+Mdeef3rUjwETk+ygYmuJZX+6TZf4gy4GV5PDmn1io3whWDTMHOG
+AuTzQsbxmpmmw72vgumcRSeS3au6mj62bAgyj4qrW8qd/q9EwOj7vv60qqX8qczxAFPiKoDQHgb
jsHQQFoGRiVgD0ysoAljs+xpPNPr+HVACbHw2IQJbiT34Zzh10wFoxkoxlk4HYv+xj7y+tBUn1JZ
2soejfin0j1wkDJIF61sBR6zfzVtx29mvkHfR4lSShO0eqkjDaL3VpGjo91AGFJqndvwJeEfnnjY
kVO2pufEHy9+x5wdAwAmOC3lOn79SvMreUOca5B5hW9PwZLQt+6lil2PA6QCP2iKkBqDAFGvJD06
UzwZ3zG9ctJ9RhB86ETcuV7ADFjKlIRGg66vx41LYQYCTwXls6yaVMqzlrWqE4aEqS8rihey5Puq
4ZOukiwH03qNNba6PKuk8aflsqJK/FJeLByioNxfAy3qzghuc9kvvaUFK0Q0aH5nX6ylwERsT83w
nLL8uRy0lqu3u1N1XMCLL44jYY8jOnxfqgg0txPpoHSCfTnz2ctXIMIlmhopKscdSH0xSi++Yadc
Ye2WtsOloJgsKGmnM9jSadgW3729cX4IRsLfD2mopqkl3Fi1uEbjahkXU0KiONzphkX1cUlcK+rk
39d0KBX1tonPCB3BovZq61Iz8svDXn716ZccWnSL/wgnYqat/JJLZ0VRWK7f7rHZMoogOe9tFyNJ
csZvPG6zrsPz7z1EvjB4LmqTV+7z55MVC18YVvTNwDT8AyyryrI4NvOBQtzKv1YQaZ1SmJmym//S
tPpLupy3UAA/iyJFEPZdSQFCB0WCfkqgJazpCkleI0ldlxy9pwubnnAMZqVpbY5K1NiAfyBfllam
tYLLK/7Rp5PyCU/OzZ9Oxr27ZbbDEUFcTHSBc0WmUPng58rcCVD5iYO1n0ltZn215eLOUZpNlGSc
C/7lBvE8H23yYSS8doxJI8sgYxKn+xwwwtHbTA3xata4gLKnirZsaeK0zOaUoE1gbkVschGEy04g
STyD9QH/9ywgdJ7vcCiRV3z55CigSkQ5NB/a9lWPxRs75CGWjJ8QL8L6fnreVnw21pOU2+sQkJDs
FEU3xg6rehm58S/JwB7Z4EZiP+OtAQSq5R5X2y/drpk7MdkdbSkOxtCGB5VHkGMtGG0O7gDyEfQl
nsGLrfuHpMnlvzL0OV8ZCrsIf8bIrf4IDf1ZduQNhCtFCGP14d5t6hceCPmuNh+rVL9LVEJKvvaf
LtqSSODG5bvYc966f70AbI4jrify/QI9QsuGdxK6EZz6Xe0Ae56wLpdT99YKvmNcCnfgqKnZvLqN
I2yrJFpc33y9EF8tu0Tvm+5izBq3DKZOZTNZ976NFzvO1PHb4MiE5JTg+QTxNxUVE65+qP8owwxV
uTpkiAqh41R3kjVuI6ePJyi7T4XT0jg25f3TB6Vv3I5g2+Y/oy2KKLC116oDnlhHHXtHwatHkN5n
7QuVinKrNiVXXKo3be1VFu7so+PLzaPeJd2EnkLO6kSWOtdCV5vQm0T1QhLzP5Upy3Buz5hoK/mu
CBFlnokHkQfg3yY3QrQmC0mcv62qRGPiqZaKbd8lg/2ZS7T9rpJxQfX4acayXVjMWBE35eIemEAo
hWaB6Ztae+ZH4RltLcVM0+B3P7jgWSsYLJ/1XJ2etHM9lLyZ4Ss8DE2cApmDj9DgpnmwMgUMlnHK
ZB4+D6GDNXsA3SefR2ponATPmtfeZ5Y1+sdP6WYDRM8z8k9h4B1DvHRRkH8Rq4CJZ7Gz70CHb+ct
8/Z0La0UYRgnibSe6/8DXIZlmIGvW6EAhapruCoNdg+bJd4a+ufs6GysdXGAe0WWvtHSlQzk5XGe
cuQuNYafF5GTewbJj+FxdQhZAhEBJXtaYzNGMNF5az5cpCN7mJKh/QcILnGjS55C8megJTbQDsST
ZROOrpyY45fRyRmyvIHH13merScXhhKEJ42IX0AQjcOkZifUXoyZ5SP+v4v6wqMT8wCynIhz312H
WKLFeWd0JiP1oaqeETPuAqDLZRzcPwhaiQSRjxpMB4boML+V/BBZsxJeTPvr/p6Bs5istkAbXp0i
qdNwSHBLxtWJ88FQQRNLm4dCObZPHRkRVuuM2D8zVCW+5fWEZk3edBIU1mlUl5le+IpT7FCnb/pO
sx/N0wdUGvvJ5WtDgavt3JBK8p4ix0DUz+hT6rAQM8BqCcP21gqtkdHp/kLVC4WUBlSEnxnfSoE0
1YH9FSAvgiDIkYuOnO+JzCRvEYvx8qps6XhgqLcstDj7NQQypNlClrmVpHUzfxo0CqnC9hTcMC2K
PUyV6OtdtLairprpcOu4VXDxdMEKg53LiyGm/Gfr7XHgbJ2cpyu/Aw0wRtRGeDZivI134Kiv0s2z
bf1RYWW6YiaPfgwE9uy3RLAIAMlLkDuTdXoLjmfWF7SoFxag6CIh6aI5xtgw8LG3dBxTjQdvlYg4
uap95DQs0O3yJZUIIAl1A87zJyAlBucQoS0K7/nNn7zcsIgkYy4kfjU3ynenhN05m+09OSZt91eP
eDuH64NiXGlB9IV/LXVN6RNRq8g0m1IaQVUhzOl0vIkfzl45WiQZOxDnm1dWKnqtXns8EHa3jRK5
TgDU+btXH7gl2X/6QbnpDh8Ud1snA1ibZ4EFEaQFgsRH8JqHrCxks0znOZlb20AvPY8ev0sc//Rx
viXpXZA9E2GZt8JjXYiTesyEOF7fQoHBwderx3Jw8HWvP2uU13WoIBr8SDoqMBq2W/sp3uYdDt+q
eWO2QL7UM+yq1WLXWdUXsZ9r3fvuE1tLyrrvURdzDfQhy/vgO+MAhmquIlkggeRm2EXsqlLFuIzS
pTmxXxwDWvOgaAaM1EwI5qwSl2CXg5ZC+VCS04+DGV01gpBLDunYbdcCc6DCYklb6mis1V+zHW8k
if/5yMU3jQxw5OSrGDkSc3GLhHd8Yboxc96e1SDJxd2bRGzP4BYkSLEfs/L7Ii/Z4wttZg15wbV2
2Cfe/GCnSrBdFhhFZ1k7hjGFpDzYNWbhaZUjeZpCSztSniXc5KyHZYWvWHzlFekSJMudm5FCtnl0
E5ztwikQPWSsnHXT3sCoJd+2yzFKLUQKXFrjmZOW905FLWAtAa+KmXeku2K6l3IxFFdNX25MJ07P
/7EPzPFPduowUrDSuQ7FLolP8YjPOSjS+xuwrQH6W2bd4cTJJ8gdXJlTN7r9XHV0PKajrSfC7U52
WJIkzsk8Ei5QaDt6OyTA7kNaImj7pfgWW9ThJ5gNz9jj/rH3KprLLPQk+lJtfGU9pglgZKDeWWSl
9kBjH4P/0HLxc/avYkCgxj80wjVgT6ZsNh5LunD8Mk4WBORbkT8f46vlCtNsEqvIxC+KStEwHK3v
XMk4ErNPNRU37lthQb7aX1klYFPO0MzJPhyOGQ3KyRpJbwG54un38WFuZmF0hOVfjTsDO/Swacjz
dhLAEybsctLRikhWP8C2Xwm1HfPoWxBdgugCOpub6Od7mhx81HnV+ln1+EtsOupeaGaIjFeJJmmv
Jrh2rMQhf0aIKqsMatutv9v8sVf7RInWc694z2f9xv1QNxbjrPw1JVr9QDdBEKBGrlGSmAd1Bqw4
f9dTiK/9RFSVHYDBqrNwW1AC/RwgNguAwPH672nTWMcJJGqXxw5wyC8zt74sIrczIRINi5olTPRG
7CkVBuUxyXAG0uQxLvSzUbLGvak+ua8iZ1bJlljQv13pISyqzsFwtqq6l7BQ0lvZR4ILYYBPaPfC
uJJwVkgbtJmhQb6kBVWmxwDpAvzfYzP8nGV7xiuxBuLtV+qDNAX1hcNimSzH0vmee7FAbi32fFTC
3cPsH1Nekgr1dnHJ/eVDmtYT/Tg9xDw86k4uUCALZtmxyYodHPXYVocWyU2hjOdYtr8udpekRq95
znTAHeErMR9Iea7grQZBH0PWhiNpkJWcx2MtgwE5GsMb7z7f+/VnTS8N9SAJZS6fnM7VAqfIjzGI
nNSUP9IobJuhe3vAjVkiEyOp8cr3CRa4/APIe1eB90R7JYNJrSrwDQ2GtoAEka2f1VQXt1nzgSnK
oxjj/+w2J+UFN5yNEhiGcfP7bE9VBnXpDumYdmFVbmRV2zcX5rOm5rTtVT2XmZ9kSD+qJlrMjlG8
+9O4ZEegneoPIMQQZg7XiVtP43U42lyGtsLFMM8DdohYnjLXSC9N5yUNQElmnpBUUMsqq27xC6n5
nsHlqDINYQLZOq1D9O4vCaWQtkSl/yfM1RGIoNO7VtDGAusQoDwoc6fCIbTuZzs1QyulCkzHL6xL
VreUVWAYlSeLmJWf8xT0ASrjDIC4frC4DaMcPq1KIiY0TM4RIAPXJKTP/7uDjJLPo61aZn7+70ZR
Zg/EXq6k1y34hCzcyCA3+U28e1aSvjDjsPXjMOdYBCktoAVFTkqcjonq6Ko41k5KkVQLqXGT8QXh
FqmEMHtv9lSt529FldO+U8Cva20+EE56DorTvSUe+XhLmeVbSOlriYerR+0IAQqIcO3iIK0K+eIg
zE5M5LcAon+2DudHPn+dEZ3h59s+b2hGm+3ctOeU8yVpRXY5dievNAb/Lj+aEa93MF3KYvtmFYW9
iR7katuU+Oen2VZ/JqBDKt1n/a654duo+UIJZSNXuOyju7fEKxNqQcef7WJNwPnYDPynI20ZKtYm
+Xa1T7PbCXzfReq7Z8VlLOxiXGw/eJCOuotL1joIHYP0fsJg1cmPRzPGMTTgUByIAKstCBBy0QtP
L4eT3aibVNMdttCvcEGXSCqrq6POG2whPAaBLZ7+lUPAQ97f3y9cQ+y2VQ7jz/tMXMsQmK1X4RZt
suHMholGTBECc3nNOiNw/qWv4DLM9dgXxeNNQUBe9MdiP/qJn73AlGsj1tjpLHxCTQvrECHgbghO
edtgOtZhKwVUiciiGkjUn7keirpPsiNAi/bLDLWcyn+M36nFjPppS+5X/hSpdjrmtkjKheHZAyTa
whwjzQocPI6tma+hASbpaawS33hfc/vmg+aq/9fpsqbtKV+VZ0RC7YrRHw3oJ9YpGBvAzApZ5T5C
19r9WEt4oeAztEBsXl/89JcQgj2WuUwYB6KZYi8YSwBlhSS3pfybqCn2cKeXJINAfpANo/rVFXoN
gn0fUEfnLkieFAnvdKHRD92emGXcp/ZBTB7HsMCGr9Ohzs+g6LHl83fFYffb5l9Kbn1WCyLDUKW1
SBTPyE+T3FvQoXfTaiqXr5ZLlwHNLmHiGTJwSDZxssMdlyBaBbSAt87dDj+/nN0LMnwzTAqMH3zx
9Id6BBSyTw3v6np9NO8KcF+xF2jOTE4DiJSgZ7xq3jOJTzgk2xcChNiYIHC/mEMjaYnTvqMrqljz
moUs7gdMhhmQJnvZSbS4eoZDfc6U/R7yQgbt/xdaOxtG8fB+Btks75l9jEbqz4MJyVrINJkh7PYr
ONykI4Od0IlMvvuG1EniqACyt8RnUrip477TUctirYBT+yX/1ridUo7xYxQ8bHh37VrYUbKkANF6
YBq2kYiCDCE2F0KaWWyAqr6sPxRF1xY6gqQXLsaNCeM+Ye4wQMpBtFBDm9jKpkfEUdOazemHoEbZ
tbZ87JA5Vxa4UuP3jFYVM8jfNl7K42OxWbe7jaYmZ62s/JC2bmEu5/KaN7jgvA8rLmokpQzeWCw0
4HbI3dVppInDSo7/9lggQuRJl3+k0GSvnNM4RgO9hh9GUmjI7asVxxqvghDha4U7BW8Hf6ReiDPB
W+sHsRuAor2K2l/yPS52ZVzshgpcz9oEKdqn/BMsVjooBe51Ka1hwMGy+fkWyDvW1bK+mNaDZTyC
xoUtYf39qyVmFKXQ3HbcvG9UAdAxX0/EfIBYYffGIQUlMf8J1zY+l1qmf7QVgbRDpaDYcMMdQ3yF
F254YI3e3wBlSNCBHV/9EEvpNAQ2KiwSfPtrLzZFcMCekNHyCO2OVTgoXMrmuxHTyuMr7lFBzcx2
fHIMWfQb88UpfzVW6Pw43T9dKIOFKFnF1Atu95/mxHwnpdNNLwJ32B1I4OZxxb4tqXyLmy6/Zog/
8Wf1oqbl230/Y9aKO5LKg94jH3oW5JcxBQo2EgILwAFvaDPQjGo1uloiOkPpDt7Z4JXPu0aziJuU
he6dSB4QY66oBwmCuz7lcvZOmzdHdyxLxm/wbBrmiQvysLa77Gs9kMTOT7KnzLE6p3ICgS0U4VlY
kLSRriFznL8J7/SPJu4T1Nbel+lfi1MlhI40Kl3DvkXZEvqb3kRtaqPFYPB4sSCWh3ZKRgBw0js1
BSkF1LqoyjAtEaK3wySxOG55INHihQBfwjvZg2A8is0BUt9OKe0n/WDWTGuo5DKqfZ4RRtRP4YAb
qVQdRJcvoPyBl0pAj3Fn8kByKJgyCi/0FaXLptyZGnqq5pZ3hHzGw8anGR4R5aHTnYBoUgCtTvIw
6ZYxi/4iIQW/iboySvk+ZXTw9BKNtFVDhS2JSfivkPCRaoIBSUreGtoQjCkgg57pHlwlGRT2cdxa
nVub7ahCiHbXWmuzo8m9HSBVG7bE7cEI5npvrckylVMahp+12eGIyZyLGge0WNQMoVqcMx3vfL0K
crmT17T3cN61/Koz25nWrpgd11KOXeIJCzCwbnsq8kQdVEtk77koB6kLwVXoiqN0CbqgHQ3mEklb
tOFsOoofdC/i7+Y5kwfDecIy0txDl2X6CUfuprYIc2P9Vp875ehT4djEd8BPBFEp60SMl6i+l4+d
h5scSNoLBUI4+AnjzTpxeq6bE3gs0M8uUDi4vTKLw9MQ/YcJ81tppy7dxvJUjRsIgRczAOdKiq00
QYpVcn982RIqZMUmW71zsipInF3aGGgf3mqO2m6voPve7gLOTa/pMyfedIr2EU5lgDj6P1D3Vaf1
eXmoPjPAumaI2+y8OnEajPWe+mazhUz19TT681cdZQZNrByfVQzqepPWFm9FJJxPkRxosTRzWkfa
L3MFTnABK2j4qFaFpcjv3IZfWmaZgHKVF1Y40phXUSzJ+bISo3RScz8dgxRI9eH1+WDR9o1FkARz
pcL+kwXwyo5IekmmRqF5x1tVXYmeFmpVoUR+DOfu5fBwdA0hdOXNj0fxx+BkOzP59WtXFYWtsVmX
Iq9qGs9SBYYKMj+Gd9nhC8ohCrLoVKcmgIveM4aepvaUp2SS8qq77AuicAJSjOU2Nn+qOHVcRdw2
19URb81W8qwB6giIN07MkP5H/YrMBnJ59YFOdVI22vo80eoQrD+gZu9BA55w4F/lfLGI+K/LfoCF
cAFVoNBVF2onaHRF7esUD4+qO7gvaev+yKXuhRyOOH13NrInR/Ty95rdoLzdtFp83vwzHAOkaXKT
IOiUqLRtcGFqWm0Xl3jPQNhbgWbo6ht7H4ZurtfMF05IJiodeTtqWyo+upuIcyfMfX5cnuhU4KMX
Xl2dVRXi+K0DqYWuOpIoI69H+GzhhJjU/sUIR1VJZXuzj4J/k7+gqHTUuQABGxdxQyBnK3TMVRMF
t+xaeaggd5obNdS9vGJAAfeKmuIBGv8i8b90fwiGQecBAXla11KepyMmAIL10iTw3Nuh6jmwhvsq
EGXG6OctJp/uwcplstgX8dpcWisR7O8XuUohP3lnQOEOWphCGAHcnz+eY0JJDuopOfIzAcvqlkxW
vzLfYAORRyuBRIXiLg4GQzvE6Jh1rPtxUoTb7FVSX13oZFNIRRKBBD6dqUFvUAn2bHymRm51Q+EL
MRkV7rF5hVzm6A1UaZuascAketUK0m6MUvx7bjFPMnGBts+9MdC3hRPeezt0kRMKZV/x+1jKZt4j
GQA/YeH1OwaxuNrQFZGPQ+hQB7F7eROBcW1fGoSvCvNvWwXCo2poLOQjqov1cP27y4O40Uc55W/L
MQXyXFLMcmpu8rZlIfhCA5BMl6vJY9SgtpOoAgGztzb2kHUnrmamLKArNxt4bw9KksWhKCTzoFT5
TGqvwXiYI1zSavkUjS49KGJ3cmgcLynHvFi3WmJzkziNTBh+zxN8kHoqQlTISrk5RbOdO9/QPQwh
tQx4d19hcaMvSU8MBH9kN70TktzzSUFOEOGZA5JT8Ye6T93xOwpbIx+8DFC/MluSuZvFfcywzsko
LgqV4uySK7M0wjD2g7EcWORgKKOzOXEIOGN1KqoH1X3TXwAKcpzeAfUnR5ifdzQ6q1wzPOIiU6HW
WBchzh3rlgAO3/LokpMryjesiW1fsO5j3wvd7utF5OT+cOEqCt/4Vfb7HGiq5LM6qTUah+YeXR0d
K91NUjR7hBFEc1T+sdVhV/C+b5JZx2XKdbp4YaDDbN6Bg70Hkl6ayNSRJzOY0LJ/ho6dWWzrV82F
YxDGc8rt1m1MFjpHTUO2cmzZo4tU4l4ydEOYkkVehEN0MorO62KbpWOBV5PqLKtB+TlDoxDH/5ot
/yDt7hLZ7TBj6c0LfsyVMTLfJW1VHuDCKjah/IkuFlEK8MFpZxHX6Lxyy5p1T3GvBTLgoMG6inqx
uzkt3KxiDF7aF/uQsAgydq0pO/CwtS53p9Pn7RvwkXZd7xilBtbBilYHo3T8cTzoUQlDB7U655FW
/6+eeLALz+YVv0lsKv5WHfxRXYVayQRjIidcLVbnZS0WRryP0+Agvp4kIPifLeOoq1ha6PAbVENi
TxMTy4E5iDXWPCBGhl1F/T+MasaGsi+UfRA+ezZ+VPvb+9a+FaTU0zN2s4DTkGUVedVJ33Fcp8mA
OE8AsFmxvkeIXrkubaVtISH3RHqBw0JpJ1nY7MPjIBmMB375tP+mTHDjb7fn+ncrj4gNW+Akstod
kIeRO99zMLQnHI4X5tKeWlv57Z/iWLspA76ODnQhlCXo6NSBUjHPgLj64E2dmUZUcKpPcb6o2bSV
iSxQhpSlktLZY3+gR4kJe2aFbVoRh32PvHfdrTsVoZK35F4m4IJ73cWdyyS2ABHLTWdC2s4k/dLT
25zrvplYBts/UoMjRSG5noM8wrK5vSurq0HPoVxueIjHz9Luch5F464PwBvmvP2OOIAwOX/T4PfX
SSRD3JGnNQD2KFHpNIzfc/xOzUC17E5XZOMgzDpNTo4D3KA9dpKWjuq3BiAT+bjt6ip7wh0cpQvy
3ZqpaazsaZabkoPbypUsd1vegsrOobJtBeeU7tHSHf6WFLGb3cPoyFZUEg99rIRl/4h6FLqGUW58
RcQfK/Oej041TpgsSTSDw5JIlsuOegJ6l6HwZ5+WPECvxb9XGcw5CMpTR1PxMVCysw3QA5e+pjJg
XlkEWRjhZSJON+25pAUHbUCWkSyMqNPQmGHQywlbEa8Dw/umeMSESsXOo2/M1Hz9ou9NuU1J3am7
8zD3vh6aa3DwUmXwZOdKfvp18UNXHypBxPNaUEmxsEOz0ea5XEEhy++ishIM+2hA0zwEKwOyD8M7
1av3Bb2rVv2bxlkA9OwQMD+b9YXHbfct6YkXinSB3y/4bGcokr5iB6WLqbV5IhsSQWAMXDrJm6qQ
Xg6a5GsCiUnP0SUmwM2s1rdg8fgPatM441ha9LetgswQMnceCtAmdBee4ButIrWUU3/FTqJBSoFA
mfbtvVNRPwzo33FLT4TLxiTmboLFiyoGVfHEQPbii3IWiAaNIaXMpPGftUnGxLnypHFJWtnO6Lnv
eC94K4jWYPKSlPL49e92YgEBZ4yhSGf32wTlObbr150yT+B2VfaKUW5xMF7YLVwb5ObgEiE7eWqD
mZ/jUih6MDim48bY4Sl/ghAM148LKb0dMhX5gtdU/OD/FtPZLfdNy1q35yXDLdY1Lirvd2NfhXdu
hvO8RQ8DZ0WtXzg6UvkqWsRFjBN4HqMlq6FYYLY5+XeoNKx6+VcHPhey1qVcR5IqRInV0BtqdF/q
SdWYRK3QARZ9pqRkTMT1pSDW0bmExXT+Xxm1Xr+z8mIjMfZD8rffXFUeV5MVo0C6Qt4DnYvbO3mA
qKO7BhHDxV3uHy6LyB8LzRPMm9GvE0T1EkQo0baG0+tMplCpZUcQtt+Xd1hlPzEqYDSmfZ1eBiaH
rq+GprKJm8Vcx5jOuUDRItqNAmgZpZL5tqYIeqwHN/43E5cBQA2FKwL0DjsaI7uOX9fR6ZXYv1cn
U/ltDHWbrOS9xwrCe7uSp57VNy656Kwm/GLCbB8iuuNGnSDvqs6EWmESMKJ24AJig2kGnDquOPGV
0CxExjDrCjhxuZyBbE4ZLXUEMkacdAchbCrXb9sn8u1SibZyJfuafkmCLLHXICPLPXltavIujLLV
TFwSCNAb8jHDKPvyPF4lsoeKk5qCY77THSZK+vbevZ/FGEd2j/e7VEx/Ad8tu5ypsMYGX9ePCuZY
o7p9haXK/BKOfwaPH17Nhwkz65GwWPP+vn8jlyaNMDXqWes+glmNj9us0wOVcoTMQYvvViks/gLm
+VJrYYusX88CLzlZSeaCcL4H9LMVCN8E/YPZfqdTSmneCovpJebw5YwCcF1mi5aGoFaszQe/5mLv
VdGUKVC1JkZS6bfnhnZXvFthnOEGY5dQznUFETUvR4uJertaELAdqbruf46HAvudJMxVF8BPb6WZ
LBHop+Asl4WP5iZtv891/J2TsPUQCt6/2AGRRaZAjVL1IM04OXPRwz3YTtQlyA7FxuR482AZbvTs
sFczpXOUSvIMlm/vuTtAwoS6/ducszKspcD5esTEVRA6BMCcaswNfECz3r7W8do9JehcFsiI5C97
iX45EdjxwmE0WY7mQKygrqnJUHySg3+rOg6Oi7JK+HsOPu1NC5ZcfGrhDkrD80AtkJf8zj/90Q/7
GRiu6KKuyAcmRA52YxX5EAyNgH4plSHM8ERsf0ZWrdSW9nudTeZjwc2+WMSdMcWCnUG4m9OrYRXa
wMBm2qRixlwMcpzQVkA1TeyC/b9e9FdbW96k83IE1XjLufn54cTnz1riCBZ3tIIhsyrrGBhkg4u1
+1/q/Z3QoWiW+RIGAxz59K0ouprE2qLTTYE+cyzs784na7H5/uswbRhptXN0dteOR91k7TDVKDYw
w/03mm/VigcnxQbzq9zwZJNaCumRxSOSF/xWSWdQNotV/VWocH0291+5GuZg6GK9Hq1qS5e78Wxd
kXE6kzVGJIzX9v4UwUm8JzYy2MtGi7R7ujww+zYkfC4JHkZd1cxWGmGOSH0EDBUB1LkOByU4Mbm9
uirZehwQSyT2fhWkp/wj2KcxNchhi075Us9+wSKQVv2GJPTje7yviQGilLeuI5xZ6F6qVXNFSjpp
6bM2IWz3966bjt37fdgcUSfk1atuaKaO41OW71lMcLHyuzhMoitiCwahmPMSsLcO/c9gRDzzOvs5
Tf6QAPGVQwHM3GN4wA7F3dDIBQFcKQDrrPkEpjWEnvfSO77sut17negj+GWTKHdLDC5ryvp4g8KO
lHAa/6JPJFk/5zIPo29kkwnRFmdXMaECCSDWTsmeFSSJ51EY4Z3roqC/7rUhucmvOUwiZoC9W3M8
d0bJrhD7nFTI5tlElyt9DB/mhyar4VyFNXymkft4hRLzBrJVIMD7j3Wp5xwODI0jP5KIym5LB6l6
nt8q0vBkSm/zU+Rxg4TVfyJ9zVjKFyRjukpdy0f/0pSgmYQU7qg6JxjjR2TODa2LLZk4qJNxutcI
UtLCIYQPkf3hQPdInnqwo2Piu5BDPLniIufUKaPBrx7oYzDRYp078R4vLNpqjJBo1lB0ntQ8FYg0
3eEhGuzedmI9ioa51KnE+xYWbxRjHKArzxGxKtJxOUGrnHav/xfbffRK1+V2h9v2ROqwClNzBS0H
IiQnUavVY3J8ORxNH+WfVQKzKKoBQL9u9rjpl2ENqeTUCPv5S5x1j09+i4reDS+aYdmvvMeHSco/
6PJqn0Pin7Q9oB42U5KZcd2zxmoCigXrHDWlUvQoRXMObWvDtodNT65LNPJYDO1jtzYM3txlP8TT
u9GlJikXgESdgX5OaKkfXztXSqRJI4YC7g4a27184YsVE6Yf/RyGTcNiupeJpbhUZ4dolBHJwcGF
bSnAY4wRhaQI6GSTXoqGQflWl7Rfyw/WTOPlDL74lSxTmfClE9uA1g2jxk5AaVn0wZIs7LwUdYci
OS1NCeb8CrWrZg/2PhqCKkZ6AkXHVcNqig2ljahXMuVlac9JlTxAitVBupnUVVXRSXqfgmnkSxet
Wf3oPq9hecUnlweoHlRNSaOOubZbcHtclymlRMBITGGlfH3mxgpOAy/r71C8kcoN7oBry/1mPOd3
oz+pyoE5XnIHBPW7nf8JY2I8L8gL62pOh1DNMGDUKo/EPnf+Nt6oPnaUt4/mAQ2oUux4+u0jPZot
J9gN3WgX3lbjBasM6old5MRf6x0ewDLOFmQUB/9MFBj1gtthRkHEr0+LYP7TsyCQuZOpppkhLbSV
AXw9dbLnPpJODJ0Syblo/fMVHV5LVlYI6alVb0HdrMyWB73K/qEAXlycuoDYwiN9Lgs1/pRut1/E
ilSTY4JG+ZoEUVSOk9mJ+eU7L8eQGJrLzn4w7NtBKAdoWLCmowuyBIZQeW3IX/7eY0VYt1rLrnN1
7aglPuO9AjSeCxi/tSpkxIKEfYL2nOwfZkvPUnucNoNEo/2LanQ8aH9a3edjJvnqrHpMxGmILksW
jrF+SL954SCSsl5eN8AqscCFeEKa7id3PUDs0oLVrclQvHyQWgMOc295HTxbZdhtXeY0UgSR+2Vf
TS0CmxOB1e03Xfh8IPjoCcxyLZ8DmEK4enlo24s5gkEtGb81phDqONwZIZt9AAcyPJmZ8tSZgFwS
ILuIzYtS91OJGyxuzgTO9mzpdp1GMDxKPLPasqoR2RbKO5vpoSSoaQpmjDLO69nOK5vy/0kdy9EA
P0XyMwTtzkue5NrZ3e85Nc7+Ixu2OLRt/9vzbPV6p516tTodJAru9FbhsEE8RyCfJY4ALzV6xiWR
REGrhOoRtxORjUUjqPSLZze/M82EVeEkn+zcGgGjc2dvetpSTT79zCu1RY/t6vCJ01LDqpezYbA7
1ab5jnfJAXtnMRyfivchoAJ2YXwGLMmNHkcrHqdD8gJowle6AQLzyal8z+r3iKpcJgeWnOGSAPK7
KqcQQfxH0jW9rh2jSZiHA/w7jwlGxu/v2hujszFH6FH4FPH4ZYNfvGC+cDtIvlzMvM3r3TxvBEdc
ZmbftE5UuKuHJTV5zg8YsFaXm9QPKdIyFAM3Egg4iq6+IJmZiSTGFbYmhGrKqwTEFhhFKCxRsr3c
7sKz/8QjOvdDUdYPYJDW36sQtVB95rSrlkhaWaSmntIUM8is0wFOQ6uWjZZpR4MO7k5NZdo40927
eMH8/qjjSIi4EVv9gkDOveeHX1Q9v+cO4SZp+IP/o7KW5oawAfnE/i6zD/icGthaZ8nEQGdPMWdB
ZhZWBhKpbYfqRBv9Udf71HNIPeqGbmNzApTJLQ2gB6/kIww9XzDez5OxNYCXC7lqMljYUEA74hFM
sbwMtwtwWVCN/0k1XwigZ+VJOrKkAkwlW6Hm3l6tDSgfh/DoZhiXdxNuMOBD55kJRC+kg+C1bVIF
Y/zlGNo38z42ztJLCZlRLnoS94QIgzFlpwtRs/1KjLiUAzxPiFYAjB32e0X6IgbS+jTmwWpZ8QQv
AX0agv1A1uKWlOMXoom25VKi7J2zNa3wQfNCA1vbIGYTjmT4mI4dstTuFapggU4/w9RwGaMGgAFu
G3UHydVnGIjcFa0/+yiHXTbKt8VjrejurynZMs33ijMGEMpDAfrHXslRrzeWbJoVsoIJzYXjOLu6
QTVAFHdra4HIVfIMBWT2D7rYc7r+Ds05B4URAbV6bLh8XoZvtRKs1SsuOiORokbEWPcGt4jZE874
CD4KR6q/KgDGvmkZeXpbk60xs/AaiVwdJrDIdLtm7Hzl6SK08AJhstkUFPs3SrHjuVQxjWaCNmgp
ogoMYeFTdcgkBZNCZScI7GSqhGBu5jUvb3BwPSWJvRPGKaJdJ8lzBnz0tF5hjvvsGrP/Jx45c3ES
LWbvnnK2zG9Dh0ngxSDfFLvO6igoZRXAqaHcuFDrmhWj1pKrZiTEFfLRo71heihEX9zmJ/WImM1f
v+/PYIg41K6SabVUFCq000R7yrKJTCEe8t+J/KuKrcY9XLVxkRmD7y/VC5c7Ku5Ji6a+cLBgYDE/
WtQCMCBep5ECZvPqb4lRMw/N5Ri8QyQqsrUoksC/Wd8nbNnhCP4Cd/7OKZliwwTSI3A+6+2LyaLZ
m6+nqDibmsaeq93jsE452ymP1TxXc5mwIr6BXl7J0dgwYYQuR11lvZHhdsQuvbGA//JvAQIjndbb
z1sAiAuE+6THKps4iodSRbKuK2jgCG25sR0SAhxCqHcSbQBzHrO1aokmbS15Ugde/zdAsLdvEOxR
dmv5HwggAv8/TzxcaBDyT5kQsodz9Z8anAe54EJeWjxhM2xfHlIlCcCpAcj8ds3sGoXLXDDdgw3X
NFtldnXpg02XYcJaVt2ne8yIfO9+ugqW7qBIndleSSqjdOwVbiyAdhy4xEYU3fbLcUE1YiIJTDxa
bbk+LCEJbI8aCiL9KoJpCO+rTYoYS9HaTY77QLSDsQoy+hLwFi/5XRRXU/f4I3Mdjuo6cf+3vFxC
cSwV1vz7nxUK3nKsb6PWqE+r4BqLXmLJw9HE9GP7M9IvVYkCjeWVT/XpVo2Bq11eIw8+RjZbnt+C
lif1ggLvipyhPN2qNMIqGuqfEfSaO7GpkGNgcpOVqA/cfbTtMmZlnwz2Y7iXC8lc7/8vWG8qOxBD
DPPKFWKlZK9pg21s3ns2hbx3RhRHB+OTVc4BOALaKswMmrZUe/EBzrPBL0M4FLlbEn/t2gaUlR3i
zuMg7OdiGPV93xaocQbyxN5ehepMs2J/h3BxuyXbe1YlAHmP5XDMKrA1W9rrYBdlypp8Y9AyqR53
KcYg8M17RMHxBrCqP3EFssgQ9L5neE7AkWT+4wNZA4tnJzyxofxxLPfWIRi0U3w2gOtUvrUMVvft
/xWDN0KskyexFLMxqkGrFSmansDoWXOymJWEPt/e3eObVKlUjjX1VLD5/TDObYgH5DiM/6XP7LW+
KFm3Hn/WTHAUp3Df5OjoGsd1eOK209OnQXIQ7DnsD+NsCYKit3V9zBlXMjliNeRg0wC7CHP/N3VV
0ssk7Qd5ffTHdZ4iGTDLws/4O6PnU4WRjNws39jvrzwWJtEmZWJd3zn6YhdMsp9i55syXCvwIrb3
YjC9SAvpJPB2cGByVzT5Q7rBald13AX87PyhNm8QUR0UovHtyXEWCgMmjLBAm3DtOF8/2/gIL5VF
RECVj+jWNyOMoMyNSFdd+vXbbSd7WNu+RmpgSNIb4EZMxXOHZVSStDSbrd5wYcNjE5I8ucWqQ8h9
HbIpV4oEtbiEFZ7WjmGEDym8bv2d+PiJYEB7VLEZSAhQMyp6NThIhHkwTqN/FaaO28TLq2Gr52sG
htV/fqOwtXSC9C5ATKfdJDIJ9BQimJpw72Luyk4blnlX7fdSfczrfGU7FvCkyi7Nss4wrn98Fi6P
HC7etSFe4TJzX5ZjC0qSFLG5i4/fAs73L6AS4qf5sKNMB+JVnT7zCCvtk6BeyB8yEyVMZOKdsF4f
sypv9F6oyzuRFUzvw5lUl34ZuOeDyAHAN7SjSsVX3PHzLZA5a1YMdPpgP+Ex+Omdu5KW08rkHNLh
4DrzHj8VlvOtjffo7BCcV3ygAj6Ot8B2A+7XK1AQR7hZNuih6NqUxVjV92cXTjyLr0C5EimRocJc
3JQW2wT0dHFvrYs3CDvkZ4d1mkCtvjncuA3apyWpS6bWlGuNTgckmKehCWNSBAymST3RUEzSsydU
uCz3RwSMysQYL/1lnRjr1wdd3f0AhfqUuKUb8hG1ADGk5IjdVASt4HeMtIdZr6TmjH3GP98pNvA9
DBdEjgZSkXuqzSGR7N9PQN+ObL1Rm17oLQEX2SP3FJh8mLZ1A1Ly7Vob0tbfmWvhogrzpAomymmd
zF7OYJ49pknx7w1t9XOktlxIRdLJOjcTJRxjw46iRuIWs5mODPOhKfABE4IgegqYMzOjpJXWngyx
k6r81mKNu0ikE8vWs/ue+ImKG6z+xELopkrnMzIiw0/xKZmXdpSp9PxAT/CAptsrPZpd+j3pCY74
yNPCkuiFbJSkGiSWYQ4/oj22Tr7z8FFLn6cUH4zdyXntgtT5TW93hcZFIfIxD1GFs/8SW+0nzTYK
7kuObFj6iHytdrz3nIBETV0dGofbcqL8flCrt/aufXj3PVD4O+8xS0OshnDl+yGTTvM33m3HBf6z
GQLXwTQTQk1vxZa5JsPMv0NoCsFPQ4oWdhT4aRmNxxPCOYp16/phKYwZdf7YqdcDgkb745ZEiCI6
wvnN45cgnLgQS8/J9fueIZxhabtjd6/QK6C1aZMEUf07upc8tkGO48yQ2IjOFOlAEbIaV6dfwpqc
jqtdy1DAb4aUZQ1bdXGo5dkJJGBCFLEtQ8BVAQAu5GbSk+5vdncqT+6PG6880aqMaG5dozT7qZdC
8Fs7GKueK51bb29GdQyateBD7/wU7rvA+YYZ2qy11TQZzfOrC9bI4hY+6Cz48DpoPfRS5qsnGBG2
dD8X0OLrct3RoI4rthkCvM8zfbJUuu/BOhEInqcg0hiAfmlNjkdHefwoPzzTYYH6LJhvemx2J3XB
/P6OL2alUOrE3vqB/seBP3Yow92L2f+mZGHgLzP8MtsuSXAMi+yV+qi5zsEf+KzsbkKEOCL7Rvxz
Fmw/h4cp/7+oooptimCz0mUTtMlMeZXtX8sl51hWr9a4Kq3EYqGxQtcEfNymsAL6p2nXe6rr5tjm
l7LKiNtqJuxwP17fu0M1SeQ2+/F/1+XNo3gKjVTOMsVg1JXGRv7hGCdYEPQOWKY9BXSeAsmKz51c
7O9JqymAty/8VxHRhNdV60X5FvluvDmrkiqOWx5WMfv5iiHEiTTw6jWWZmyqGE9/tkQfzUG4iqiP
nksXRgbugqkYdo/bt0D905QqfzsNktjjzsx2M1DjkNDTlcGCoxJvc5Bagi5o23LXeX73BjWelxo9
8YLYKPckt2Kmtcd94wYnK+E3tgPu2jpQuzMfCepAk78hXovP7W2iezgXpkJGbRdNC9ALNYoIX07O
BxYdArVxlE5Q4Ztmis3lJOChQV/hcqTLr6e4RvxmendmhcUE0S1mjVYMhRS+D3AkGbk0IRfY4rt3
hAI4a6GLqRz08CAMUB0KAelaiaLX3kdUDrg5rSYPW+8IV2fd5lhoKFeFYOILXcxhW5P/xbhe2yBi
mxOHelwk4GWwj5xDidy11ATDDBB/hJyTm880Gh9VdhXGTo/svfYRPE7VotdYckjfXtHUu/mHCJLs
Oscrm3PhOZOjxEjn9VvB/7n0O0ZOo1C4i2cvyqt/78BRm1HabE7yoaxDQ+oCY70SdUQ9la5y9Jxb
a91n1+h3bGu9XB8kmtAWGMO7qAWsXwgCpd/heoy+CtacP7wR/EiPxd6HtfbrKR99QZOSBuSrNI1M
VnPOv/HZ0Y9K1HQphIUWQCXKWK9zsejcFhSIgi9l+xGnOVCp2oBmPGrcbBBYOxT7JcUkXKJnL1tY
ti0ZM5MuBBP9hkUjIPHncV5keAgtTkv3aAJx2nbsJsPefDxrcpNn9b7zh1kEx2GIwDcQF+w02mj4
rfi342Cv4qgboexRy6VOtV6QiffXy8q6LyZrojJ8a1pNOO7A4DO9RhWoPj6UKsyV6XKePwdWpeWL
inKsZDoNmcKjs1Jj4gUotpXLQfKCABsTEL+WM3F5RAyQT2nsOWXJWsvywvhxagSpTwmtbDKO5uXr
4jN+kit3qXIZCRQChr5x6e4UXQhzfO/r4LW6DttVFlX1E7SfMsqbx3kchjlqkf2UiXPv9aJ5Dh7X
4fbGpmFsEaj2VXUQ4EfRNDPELhpnxUn7XCTqOtFSpBqdQ0Ht7Zgwb2InV7TuegkZr03ISr2+SeZ9
C4Movqi5cGeGZ3L37sDk5LCh9cAnsrp7vzXbdsCYmJZABLjThbKjxn23md5ry2Wg4Fdaz3B8I6jX
908Ib+/GWnxrTI8sLFeW7NPoxgoUe6XWoD3U9UjIHWQnKs7fky4w/l1Cn8Px87vRTfA6cY60/rBq
nwnj6/HumYRFWZ/R6vBQKjKAk8gt+r/l65ImCYWaHZ92/IJvEL4AMhoMK6fZhFLKD1PMU+deo0Ki
Fd/ujI67/1/0xOFTEO9CDJL+NRXcqmRRQnD+HtDk4yPaOmHO4sd1N2vrlIrd7RiOKegKW8sdKml/
kLpM0ogRoh2Jwa40S6RPu9oqAzwz6uOy+2Aen7ATAxbbWzTd0ElNJrzMAediyNxAwbis/99fFuJK
aGOmocljIRuwfKE2MqFocJSfa35YvvYE5KKdXUkZLebSfBab19JG316f+OufrhEfug699S7+giKd
oF5V5PLVKmqvEMRDvYhEGcez9NoOPondVbOPkcud08zGgbtH9c4l08XzeqXYidySmrtz1TmhErhB
BpVSwEaCkXwz7ZkAbun4KhbUDqLaO/inmp5aXznotXFR1CYeeIIIIkP4mob0jQN2D0IGFdixJ68m
dSfl6On1B9m0vYXPam4vFSU7/mR7l1M9gpkWrv5/1gh2Eyhs9OI/Ie9fCAwpWyYPZu1q8SVpWGFR
enGerk/Lc2LSWmkRESDMAfNSSnwmkwBKEezqcYEJfSGxw/sKdNVz8sgu9iAEYE376B4Bl2zIcuOQ
cdm4oqrzjC+wBeHNTs5C3roICCs4dheJyNs0uRihHvdia9eT9v3VtxiPNG5P3GIAvnR7Ns4ewI4i
tYD3X3nwdA31KKp3b+ad6weJ9Hnh/NqbRLfElpfcH4TuXmEcxUJjjlJfvFZ6alHYAfOPckDbhvw6
9zS3gq06tcrErt7dwv9mGmtSxPhSNBzi2EXxfgwEVX2l9BgS+OZNivhKyE8e7EFBKFMYQm87zwdX
UfsQ6qrWN80KS2iqdeOZSFq3kdr9MHQ76W9pGem4NYXB+EzzaSNS2CQ1J131oRiA+Womo28OAzkh
Z1AY6oV1V5ABYDFYk2g560JRyV+Ws20+DDJErPHLR3abx+zubhS6BpcbxhY8ihAMgFZ6qONS57SW
0ObpFZfj9kbTkD6m9HJ+C2+EMiQF6xvyNkMBlke8rbVY+7ngHYIO9LvhO7PYAF3gyMntOyy7c2Mb
HodinVMafvVuFKQIb9EtvNefgQf3xoNxV9//F7OA5tfhvl81ilErkXQ7dllRbsXODwxz4HCIHba7
ZBSi0Xwhy/YfqFc9cjC9oQpnbmTmYyOYPXIrk7GcMeBXL0mIjs6BeN/czxSRjNqF9TcQkDst9ZNA
zM7Ohi+OjNCCvd5nmwQDgVmbkaIefDUOz7wnTQIuN1jQ/F3mgJk6/kzdABww3izKHMgfZXgfDkJe
ucpvu733k7bYKVvxdtwIcaTrZIxQ1GXBODbONZwXbIuAVqgFY/AbYic2tZmh0hGiB8yXCeUUuWTp
z9rBGH2oDuNjdM9Hi443oQ5KAnfHlUJmEvnGx0ek4VcIINuKQ8AqPtIzp3xZkoeKCF4A4DJmVgwF
JmknPrsYebzx7HKYAAWoHwEXr/5essbEJhMLkJF4d5Mw/udwZyTWlnYAFJKBx+SuorKHTgXELX0m
MXht7ZwXqmTIe/dHGXKGYDkHwMYYupcKsrk0mkjo2v7pZH5EWZihfx1L1pOKf8mvZxG+FaszZ7vb
CsXFaP6v5wtacYXv9wIu3A/eUniW2w189XmSGBgkj24gDff/VbIP8SmmWR5hK9SjngHLr2Rq3tBa
9bIKb0T3ldSHiZwdCxq+7PrQa1RnYKKXlkynltJO8Z/GGqLQC+F3UlU8f/LxKCzQfUEwp8kgrggk
34iW2yVCIGz1L7MbUAQAtBJeZCjOMmrMPCnKUIVeeWNFukEISfileW1mftORMgX5KM9wBzdNdHbB
BiMC7/2SCf3C2ksTEf1skkqlk2bt+1+swET6yML/C9qnJfWTRT7uQquqENtss3jjj4+p9et27Tef
YZ3DcYOXgEKltNdVRLKbi/1iU8H9LC2vFm7EmtRKe5kxq26K4FrZ95Xal/rHg/dwpG3ZoqKqBSZt
S2Q8B74ldI46rFEBwosr+82i0Iz2MTXo1fR/AHrxBHFl4RI0kaz1PWHEEFhVYTsj3UfP5HVNlhnv
5E5+LHqQgfSm6KO6hj4pOtX0aqagD9U9q8ksuE0D+5p0b0m7/jv8JKbiy53wXyZAEs5fCXZakAGs
7xnnm5zhNepE55zXauHjcPQ4VYDACR0OsPdhJNmjoaK/k6rTkejc6sO1Db2tHH2DJ6VcAGzibaF/
9PSOfnhinSnl2q2yAB3Yh4k2LTFzynXuJVjTsvWjk6DNu3qhs3CFxQc6swPB+6Q6XnClK00MFcxI
uaHTUidjNsAa6FNHMbxGmUmVmyuwUTJ7+HTeByTTACHw7SRO1DoRKplebl5fBF6lrUT+4QNevUa4
Va3ruY9arqSx/ycMf1sN9Nh96xhJGwlzYFqUypS3YOjThmLGsXJ868y8sLbU/8Z/lz3aH7KPTn5w
iZaxRkI2YDU6V7L2lUjbb/0+VmiRhJzlw4jq4L/tBOkDhSMVsqLekHu283zPYQwyymBzFZby5ZfD
c+5jf8iOTz3q6eEik9k/Be9D6iiVHPRgss+f3+I6e8wj9775qF3SOHFleKHInJq4HXsl1rZV0EuG
6cHlWJTcFasQpeu65be5+WZC3DyO7Akiv9IFYgFyjpW+3iW6Ssnv5zKXVbUADljCpQrKCJEPBmaQ
FUlrweGlL6ZNC1EQtC+6p10Y97qAI8yZyKfOGsZ1/kCSGmc+kLiKsUyArwygZp6VIc7PftqYqv0Z
oFvlrDko9AcayONPhQEhoC/yvSjckPoKDCCnItV2n0BUEbs0eZwQZTwmRoUN4D+wQ4Z5z29asYPt
h6BUhNvJkpOKeA5T715ELRqlgUpKjTB9i291PTvWn4xBRdzPIws/4Q/GlyVwk2nhwhDq1zOmNQdo
g6+0KMdzBT3na7+P/dITQO3Se8+QnnlCI4f7CHZGK8b5pIkT20KkFHnU2tdx1Juzbw2snnPnKDxM
PHDDaIzY8qhGYB1LyPDscfDB51cV0SBPG6zzJ7ALvGzhzl8+2DBN6YbDiGlQ5b3pPDQNs4WGRhnB
iZ4a79qyuwMoZAXWGhYsTAR70ffmnqhfnM9VDuqY5BYSmVRnD5g9HqY3hqLt1lXPAqG6Wp5a/2lF
YhDgO1cXLI0vUGqBsBp4Qi4g8dosOKxQCSsRMWAdzBacxrWKSauE/1cgbgGTPNHI1LNqh7zA3v3R
wuAJpYf/XkS1PcgtvHL9lLIUNU3D4yKWTagvdnBPci9zbi6hgemWzz6jvmdcKJ8mW2HzF9tci11h
ktXK7kHTFygqfHfMRRlogTkVYQxETSZiIWtdsPrNIp64hkVlbrnLL/FFtx3SQxHHTSmqEtm3SI3Q
+3TrBiqgAk7oNaDQR64AdH2Fv0tCvs9VEKlN/AnKj+QuYpiSRxxgYZUpkb8aZ5Hi0oWUIPddue5Q
MoEKB9D/SHaOk+f+sth74OQ7sWkwtOBoOqskj4zjq8qH+N5zc69VsdFaPW31tsHDSyJT7mkVJNiJ
CeeHQfwi7DNOqPMcKMh23Hg5pWWhd4+JYavqTyA/z6WE3IggmxK3X9wW1AXKjh/nEj5EcvgiM8sN
RXRzs/XsyAtEBUqYnXwzegJAgjBdvbkNanORHTTrhx64P6MNxu4ehDRoOvXtm5ssYzvClUuEcqhH
t2wQGOgGXFJB3yCn8joVSkh6bf5gkzHeAmWhJkuGj/qI9FAfP2S6kaVHy1B1DPsTIZ3UEKzSV1xJ
FL9yzCEiBbZlB+WYnFswNGMK+2JFhwhYZPjIZ9q2+dMzCrgky6KX7i2xzlQasEHG3LlQSH3uPvOE
IOzJcyq4mSfxlJWYCpO/j8OtyEB2a+Rf1uG08Yru6GZTMdJlJQmqWNQxdsGb2mZx9r7KaLDCtBJJ
jMaUqS9JCZalVG8iWwLDS1rynOrVAFTA8xheJX7L2zyb/jK4fp7BXGoVhnqeBcLAOSjA0HIA4G0W
w08a5VqRh5g3901dSy/R7mpjmkaeQTLsI035WVMPIrCotl3/HpbUn8sDDsQZKaX0gCenVAbotaMC
pBu1g31jODYW7lfC89Ovno4Qj1nnUlp8Q7dcj3PfzQF5oKpplH2I/1y7Euf7e/M1W5Mzk/iMNNRM
Ia4YKAbT5S3EB3zXz/QfwCO3q1g4W11TOYd0Ri/6JMMqR4JRe8JO/ApWglFT8vjxkI5mubu3Q0lz
2tjvnlilbvZAGgsdJDbRn8XJ5Oq22MU+ccSWM4y702UL3g8lZIpIHEI68NfqBKF4YXh2uDxVLE3C
Z3dRQztPdsj1bgP0errfoQzuSJX5NtIE52Rr6OmKAkfJ64qV8JZh5sL75iNRi8d8C79OmPY6CKOq
7gHxVP0A4Zw5vQl40Tx+q1zx1vUWENFsaRz6Qx/9ZROaltmBRR2qNqJ6xbuft8drmOYxbR4kIPtj
QM6vnbRtKZVX+m0cS7EnOCRMOWsyaBnV2I7N91I5CBex7JNXWKUM63ODXNtJUbd9ym9REgeCdSQk
hQTz/UgKmswdu7Y6J/JPYVnrrw05uTvEHAYJxJxQa5xMNIlI4EDMbau14Ic6vcKlJW778WHYb06F
AYBKCtAOcQAeIWceavvx5bbTiYqfDCRsowTLHtAc42XrL2dQTJTVa/D6eLoQ92UaoL7wW+xOzwgo
EvcWWxD0LoNPuV1c5JRKpjID9KagQcKKGzKd5oCUMKVme7N32z4PmHAwWhJwCcMqcb/XQ8CsdMIa
oZOseEka1MshVOvXghnV/es9tofgtBzkIxqUYPc/FaKdZA2fSW6cNRyJTwpPLPiJnoNOCfJIrHHt
hTDO865QNTORNpcJqEAboSCDBK9EJ6vv68sZSQX3F1mShGTzOL3GcUFORDnCDvVNMUg8oi6WlJJv
nV55yIn3OurFyURWQds7loiVEMxIV3fPS696K1GFeB4gYZlhMslxiXJOoMED91jkYWvVeH+jkezT
AhyyD2JbCxFQWbUit30jTGxBZD/zu3SmCFk6T298SEYgTFah4WQbS6K7egtFjCiJRssFxdPP628P
rzuhGwmnKAtfAlNWkEph912ZaMBACkTKfJQyh7nkiJ4zolGJ2jAij9+1lZcR1M9m6YOAOmelI7Xf
ud+Czs7XxY/1b8wdmxZLDUQ5EiV62WBFYsdA0jSDxMdOiXd+XFd9HLM5DlCbxgA9/AvsAnAJcMxy
eotN40Reb0089za1tePv8tA9KnKjgOcq99zGFYju9Hf7CLuKTYkA+eyTdw/Ixlw6XaXEvxGMCZ/G
OPh7jYVHqVgusug7+gWXVP5M9a+HMjcfU2TI/v9O1pBvMne2/5UsQzrl6MF/WzPs5CfgNnrmlaDR
syZVzZZQBRo1zIey6zkd6WFrS4IGvC06gKT4Ei/LvWMMpmy80Y0smpAVTPSouJa6w0evQEs3EkCH
6xMbvD6Qt9yWVQ6MH30alnq5pHD2NwbWV8M/9vWjtpQXBEjwcITNHXbHhvyNeH1bpX6czv22fu0R
lNo3YsrIeu8TgK0hQBsQMm8+sRwKAI3vjBgQX3h6dohLnBKXy9ZN2cVe4GBObgJgSLUI64VRExz8
uU0LU38tjZ3ZnOFAgUC033FmH/nFTvti9DVm1sHa8Ip+05Tf949F5KBOY9aipJhg0qFMdu8ROhqN
IZ8+CTxvaRVpU52ZMOvaCIWP9I4AwVyqV4TC9sfirmBPRkhRk9vCvSpL5gmjAsogeQqUXdxQ2q8S
qclXfG9hbVwJhdmySuxrbKmoIazM3oEfXpGQnQq/C6GXFej7RakQNznaL7IMiCH5f3tofYuvdlOp
eTPKfjvhHUZtUsjlQ7gx7c4vaACUJ1L3xgCcUiQCdCtKmP8Vj6jA2C0vn82DN2vF538bceYkbpsE
ak2jR654kXQUrCMjG1CnTy3Gxr4MgtEUVh6qhj0cokpjfWJyoXr79IZCo4FW+xsEOca0d1XAny2n
0Nv2HeOuHf+9Sg6TXRVytPJ2D7lCtly2gCfahDD3RhatYrXSNrQus6bYcUC9rFrM3uSZU09dFql4
Z+4OTGivWoRkut12VSPO/Uel0Xd2DY0u8IiUZTXqDOODPH8Co/0InvIzWMQri+3tKX+YofPcnIrW
SCdILAtmA98vlLeY3lAKXaamQhAMQ/9IQxOY+O5wCgcGYok3xpe4L9WKVBHUzeGvEjUp3jNm+r2Z
DtWlQfTJt/jR0feKc2vEyciToIstsd4cSnDbUXKWJzvpX79t+GKOkbjzt5oelita29JiNf8CCQPj
Ad3FE/8COCXuhLT5gqfTJajzv6oStuVwgelNjOStk1ijKBhnSNU/GlnB0mnh+QBtHRjpVZws6V2d
fsU/pEkd5olJRAoDQEuf8JRdmCUafVpFuj/xDEfcpEwJIEOXibkpPjw8UPWn++8bk2T4o/gXUlgP
YdVTrbCbETgg5FWWR0vrtxsI0Pp88EtJLFNXqVXMNDmQrlj7/Y5UXG4y00UezRi18M2g6drgq4xG
U6hYUQ8j/lc+tcfSnx6j08KD0ZVXVep6YXhpm2G3bIEtyhv4ZiUHtVK7sB1FJ6uQrp8d8rd8hvry
fayA1l5KVqvq4c4pcYi3RUd9GnAJwIqVzqiqrpOBnGCpN1JGBQ3sMq0E0DLhowb1XNkOtzXoBN+1
UMMMvQWQwIIQD1B4McZZKsBlwWunG2uxSlG+MyzZpezCGmt5kCOf3maCdOEgIUWWTBBTRVPpWL89
GZgzQejir5h0+DmnE7LufeKRYUU29CWALlDdwDWSyFWhJC6d5j1P7160mHQE44FH2sf0d+BFzJKE
MhU5Df1dcY1aRH+spwcmoy1EPBVn4EItSqlIP+rtoUz5V961SYsfZTYmGoyLhoFvlIMTqaneCVdg
6fEB6drXjY2TDfZ0df+YQCSwGD/G042/4qTyRGF/q3aStX2gGhKLM9NR4IkAwXeSmOxUSM7kb1cb
Jsz3tMlxizdwnEK8UjwIyQDeG2IlnjCnTsSr8IhB0A85PgX/3YXd/oqvFhaASD4qOYSfy7nRfohh
mi4LMV4g/cPQurnrnDJkrSgj59duXniGd/PNiqu37XXdumrvwRLh7MgSQNvubUgmDfICMORtPVP6
nqvLjnL3IbPCaUonJ3G6EuRrNgQJMuZuHOFWRisiMj6yYnhq7HVKAVT8762+6HSnZ5olTASsH+bA
dWSEelZQSMvYBR7eOdEwq2tKrxAhqb3C/7TTqNdnSNdTHRk0hHoag3NOnaQs08N1SM9TmrDfqtvc
qCExnlK3dCAASS4sATT2pXeE3dQbFO5zk22zfznks32t2318tLVg3CoxERyIOzkcxNvwIsxGr6YX
r2TBAMgviJHCQuSKFh1g8LsOedQIpTlJtbJCNV1OrRNGjQ/hj2ZXZePMugbPAdDqvK2OEP/4Dp2T
NZsZUVnvuhqDFDLxVcqZgamxgySVzqUXo6CskFwm9flFAWtIm1pF/4PQZjAzaV+DqHZdFabxPlzP
XbpatoI9bwwmOfRs77RtNPS6s50LAUXcmYkfahe/r1kGA5X2pi4Yc8hJLaHftlWpWYFlY2A5f5ES
1AGBGkE/wTRPXNwJ2t9KlWL12bdgQRzHOIdQ8dNhnGXMJmY9nY+eRkai7fTGj9Sm+9KKdGbTGri5
OQRRVjQtojGlIkqlHe09Fl13Bi12zZpZRVSMPuhdJfy6UKlYA835A08Tw+6uw12+C3r1TWBM9yDe
HMTP+FVGNp6f2lbEexy8LUYUmttmxQ7JBA8kZDTZE49hHr5pog0vpsR7fJXILzMH+y0ZNAFeG378
C2IqH6a7XFt2qh3uBr75L8qq7k/kPDV8wU3/bRX+ZLve17UWj1f8OZUZiuY5xqEw4wH1FjWBVMHg
7r5TZUNYXrv0rglTWHhCqjX4LU6tCs/emxqeJ8hkNPnLGn6t7dlLgJfy7OrolSSIpuv/sy5HclWq
c5TJ1angVg/xNraXg4he+GPkHk8NGr5irdZuyZmTwq4AJBQDB7p+1SaY/3xJwGAjzIe2kmUCpXeQ
uAAd+9yvInExnEt39bWDPAwWspkRESOia7ISNHAdozAu2Bt9iV64KeRQLUwqi+UW+NZo8uLZdmE1
wOGZgSyk2ARQXvgmLuB68Mymfywi5LwOPCkpN/2iA176FMM5/qsAB+VSHolG6Il+f01lJpPLXdeZ
GlUsJRpc53TEEf+YLrC1baXr0JTKFJsItUkuFVXXjQ0T/ruq3P4ocUGB+seVCSPyNbw0t9bLD5+m
tm9yCcR7aMrHchL6wwymXwwIs1aYxQpj3UMl1y8lfMaiLZ3G5AJCohH6UzFZm9IHMiuxOnNqJekr
tNHbaR8Eav1vSzhqG0lAT/1lFCdTJ7/bl0WZ+C+rn/BQ2QBRUxVTVc93gnfzr3Iz6//wLnBpqEXv
pMsWQqxjqv9DBH9phdiYc1strLj7RberhpIcnDJcIb2CIIrLGt19KLbmCS7Ej/Errfo8BL4sC1uv
kYf9gJdLk1s0uAgPS/B4vkcuAhYzupt0PxcSAmIh9d13b0b/MzZVieLcD6VZfCJmalDAgqnqZ3xC
MZHH6nNNJl1Ec7Sl5gO9dKQod5tDxAUtJKDaLp4UPobp5d3kHdCCLiXfKPF3ccio5CdKMDhIWvWi
M0FAIhXYU87ql+OP7b6Tobc6vv/0j0xLfsR+ras8R3/653dvyCFUux8TVg8aVDMQNyCF+12LCAsX
gksWcT5du5k+zPqMWjTID8oyYCNa4xgARs4eCLCvQGKocyUaJctkjEL682f9ham0t0pgAwPKsEE+
ALMtqMkcTZzGIkPRBW5Yr5QDCeY0ymJK6/CNWnb9rLywpoCkKVWySHwb1rgH815QSqsV/RVN3UVN
aUkH2g9j62Qazne5my/RiKnCS+YBEmUUK1NU8WfSb27qGwshXZHJUnowsM/t41cSk+i909In1KAM
stWCIebXO49urmBHVAlMGPfpo85o49BWQbQSzNyNvEmLqoycl1t+NlkLwZWwaGsGudh7bZxmalQk
IuxirvJSrBBn6mbNZIM5vRpcCkgByeOdDNnuPRebL88ReBOrtOYFI4JRaAcOZ/u1bzbemgOeIJdH
Xnq4KKgOR4kZeH2dY4jyE288VuBus5Ou95xUHqbF7wYfEF14w6XJXgZXMjA+H2zFCXy7LbEvCuF2
mIiLrjZiZwyEfD5sYxzPdwjIR8f/gen6LnXyNdzHSH+AgPNqzo1xRWRw35ivmMtVi0JSzwzwZOOd
k0nnc71BabSe8z3OE7yFyYl7L+dvM6miAgS3D3cGfRVP0RN45uhERF6pkmR1UM2gI1gOmczE3ZsC
76z7o7iag/LhhlBlG5Mq993j3MWVNbvI+s1TWhWEfUtzR/GSt6Hwvyf8xfGPyH/hPaqNstlRG8x3
9RA3yfMF0BTLW6HrdM1x4Qq9WYmPvCjkg4TI4b8/lUvghGfpPE8vCEv4c2CccoMbb1rt8TaXQPHV
2/f/QmQWKsYpczZlqBKQ+vyhlkN+DSLswAIoLexvZ9ABlLFmyrEiiRs+zTfWZ9cEuK/B3cwbref9
uWwE9DuSosxS+SBLLqNl2aDvuzRRx4JdHF4Z7NevHrTl/EJgxUUXrLYWKRSuMwD1S2LYwcZh77cp
CFUuaUHT9CMJCZzSe51qghuj+MM+S9fh+ttyxFiBpaWulKvPAEObdHa7nHgh3Qnr78m38Iuxebsu
yF1f87uoNdFpDZJ9U3YAyuakq9zR+22NnKG0zfFIG4lXje2zOlupUaToWjDR/WHng+IoUXaYRHyu
1jfcjpLM4MZLdHhMuInwtpm68NQCZx5ve7LQ86kzp0qBSqwn6Dn+jyFTWTX3TXv3O5EOcYFhy9Ib
JhgP0mqXE+eND2MkRqQ0H2w+mA2iZNwuVjZHPUsC5aost6vD2siWQRe6x4GE6PeVTSQvA8KDjBKg
mEBaoKDV8AjKT/LDY/RS3auActT2LC+u1We1Ab0TuAaOplRI8tdfMmtEDvzN2mV6PFFm1uDfjRfV
qQDW89MjsHrvDpNp0S4OFand9D0A2tYuxdglm+ALV6xSA/gLmO/n2XddnB/BqUBddLVQ9tIpcs3f
Cmoq9XGjwJsWzbI5uD0/Jw3XvLSGniJyGgNFw2PCVJnniOKjeusq8PTyEuynk0Ptb6it+uctoo0a
WHOJsgPtt1cIApHQ1PtHUcD9HD/arc7TMSnLXTHddg0ue29opJmpl5Sn5oDoK6AnUyCf6u1r2oTa
wkQyF5OErct8F143JUgudpj9OU8GxsPgHogtAU67wWjK2YaCor6C1EJWn4TIa7fSX9zhGb2Hy+i7
7ZPWoRYqq9Cy7Ndu5P8UOiP/x3LDHS0+yjVtIlFKocM18sS5Dg8/wJw5qk7S6w1TVwu9A9b7hKmX
DijgWkst0R5xCW9bUVI//j1vDJJHkrjRmr66hhHJCETEoNQB73kA5+VFLOnakOJQV3H5GGPhbeCf
F870+XrWNGb/wBf6mh/Gop6fkzl2fTPkO5wdo+UI3dHxJ3lvGScL+DKlwgmVJtUfxQn4Qa1ug/UK
47EK011xk12+wtH8WxEWxN2CAGxDIsGBEuErZBTSYtjKL444pZonkmOYABkoigGSXfd2inj/PKrA
XnVvoYzvqct4jsoMabuTlxKn1Yd41TV1tNSL0W6lohzEAdKaGTXLrHWGRGYc6VJOHLgnRcnwJBHe
MkId1syR5MtFMyRWQqthxdrDQMxhqBTnXQfnk1hg0doanvoJ4d77xCvJ/UY6nfaQ3BEfAbKppfel
o0oUF7B72JDP3yZzj4FUO0BRGrFezeG5wyO02lXMMIcNtejPEHOEPaHnW4+4oKmSLnOes3ABbqZe
tUKS3JV9cozBBDrya6r51hFS0IhVHpkhUcp+zMA49OvPh0Ti4GKolYfGU+3amc4dHurmRe0ddAsd
Wtqu6iRhUigynU3SLwQ03/raDIhHfgmp6gyHb3fJVzsBnLrpbzsfRHZ4m8MKGyw25GUcaP8plFVc
/6DKcvtwwXi8/PWyqkYnvtot5xmT28x5KdA+u0NboIAOF/8CcqT37UycgC2jE6QgVo6/3ray8yx9
hgpBsVtMhPdWzN+xVBMbQTL0QLgDJmYTbMLJxI/r0XeBgQQazvhwAdiflhig+3fBxr7mvhhlG5wQ
TyDAjHpvgnjD5NTDDz+5ORvJpq3ImTx6ENQdRFO6qK+emsRzrgCREJ1IJZF51gbFHk0mVELXQfVB
MN/iweEQ75kCI1gzrAMaBpZCq03aEt6iFQka+hcsO4UAeEj+R29R+WxRW6a5MfBeDlry50K5E6dZ
BwXP0KJgwMUxNx6RM4uO6jaYqnAl6Uul9myi50JcDgTi7rpIFcOExrv9qH+MeDdsftLsE8ixCKCo
aMz3TK6XvePNs1OLXBuhiE9+NQHxpSZGSh6ihHrAUVnudThSaxHEpCccujOcjH74F2Zz4939+LzQ
9Cji2oI0F/SEm5UxVfDknyS7brYCS1P4Ohu5cudwku+oAaUmdwi7x8MSKGzzTJRNrE8zqbl8xX9m
ilBHfhirqttA+91bMh3l+owR2qmQgWelUkL/pdhgTFVvv9Fs3CdryJSGv78bnQAJDuuIJ7o2bcxr
9pIVj3HgUvSt0VEkqtAd7TsOw2I+hr1Jo7EyKDyfuP1Po2Ck4ik2VvW7jmHHqbWqm2PCync2e4Me
TIg50WnDsgGlfjR6fyygkvtgEWp4M5XGhLLNiv0UkLMkEUF7hp3glxk+y9jO2NHaYclWS0w7zWYJ
JT620dsPCUuMVur4Ys+h+GFa1Ev+njWYwNNWXHZz33/htY1lXp78mHqipKddW+8N+siHYxh5zWHx
RY/uglkDRpC5R4EP2fiEI9+4cXDnxqCaua8oG30tobENA3TymFm80QpVQELphTx5sYQZjKywu0YM
yg42w0Y8OOW6Ds6OFnBY/nzikfmB2QkHxCT8nFOY2iS7SSYsVrMeAEr4z/e1KODW5nNPWZ4pYkEl
umMmjG8TgQDD2zAr3fAyT5kA1jDiB0wgTo8ijQY1p7ahubucwrFfwM7TYcDKtHv4bMomB0OuByKk
JWynSipfAaFoyHMepovz3mj2c/9oeYPzIaprxqd8EPJl5ycTBxM2cwt1CMI60SSZTlo7xL5wRVVO
7ot9G/WhQqdOeyxzAGP9NXnTQY+ixhh5W5tkNO0pX5WFm/7+Hb/sX1cidEPmyyFYclZOZsnnlQhp
zadMXb9gDb23iosndXKPkl50tlEZ27yU3jwmKsfVlfVHQl9m2tv0lIDvSkHDpozfbPZzojW5KlsS
bLpVsttN5k/aBEUbZnvg7jci7m01WVYI96sDadXEh9HeY3Z1z3zTwi9N1T2U+TVB/erPPVJmYz//
kIyU0xIJRdwhgQZxJVL1ARIzd6yfOytRyu+yNoAmGy2O/QA0gDHcSbVDvrnezF9E4z6RKg0DX82D
6U0tPt9VL29YXJYh0E2yHipYhW0s6+M5bc3hRL2hwp73djSiU/NxHl/Ppz/2XlHIus/aAYE4fkse
CGzLiGbU+PMEHIAQTtzCu6goeYNGBi5TXqF/zFVjVW58viOr6oj8dluAQnZiXLv0rN/2b5ZkeD8B
NaHNdDJ8LRvUCzsSzd/YTFERXD4PX1Z7xWeWdKc6ZBBagiNcOrqDe3IrlO1vo6P2fEQdNjCW4LkG
5oUiwlGu8XHCEu2kMzf97njguiEveeIIQ/Eg6/p+fGZ+etNYLhJbU7Gpw+3zLuCtyGBhKp2G5FKM
FdmeTh/kco1HQoOSw0A28ZJ1L/ASwAEkcSMke5/VHlxvTMQKlS38tBSp8J4cAgC0AwfDAiF+HR3y
Y9P787jm64rn3UnXt2QRDwtpXh/gTjkm9u2Thg1H5rwC9KCuVaRyMSqqKlY2k/1/W9uK/q89fdeb
vZtvfnVC+QdV6c6tts7NbjamKQKWiuGLtLY2zF21r13oMII3lYUc2aib7POCr8S9ujuxkaUNO53r
RHNqT10k2sXzci4icA/KV7zthJZGtn63oQzd/TctFM0fjSVyp8h3Cl96dnBXfTkBGYmcdwlxAEIg
JhT1grvMogmLFR5dZb2sM02bxNxxYdOJWym3OnccMvzfN1nvYH7xOh4AYCC1bk0R3rJiJwWz1Eid
Ll0s9Z1B8hDi/mIAIYHd9kkRz9hJbmibvEFWLjn1GADW2NXEDNtJn44BaZntQ/Sve0I1k0qsAkoT
3YeOPVYkjAZym5ZXL4NyBG9RaJISZMeRAtjVGMkLM9kOkevI5Wg+TFCE1PhZE28ekjmBf9jIxi0/
TOLXaLOf/mI+zP2zH4sWuHEWkyVnrwqYAcz2vdJUx8OaRvyVYHyQCrmTaTBgns7Lrgs+UiEJkRoP
7Hbk/kgD5IQM7vAn5pvY4kgnjz3t4ZXp05fbBdPMCtywKXTazJCJpaaol2oKJQCUK4JE74njrG+z
iC4c1vG5JPobLcjoNmQwG6XsihHrnxrkrCEq3ThOEo0HgpAUM8gA1UBf7R3M6nFw04GXL9qNmTEh
6Zamh1/B6oBV2TFALBUAlczAyZs/WDCT38HvR0210RO7sM5KtEF4az8BkFghNVN8CzFLyeJdKggr
9rO7GZEpmuVLrqpAoWXNP08UMmrqH7qM+ZbLl197F3f9UW2VPqgUpQWVxL5oG1DvSS/M5ybdhfaD
0hn/+X9V2kG6/tRn06PsJMIjWWBu1Rj7A4NTEhkSbzOwYa4BXlykxKaCoIyIyzd9jPOkN2xT4KTz
bcMHf4uk2BdJ1CPWCtGWtvSLjb48tcFFNQvBefAzAFiYyLaTMjEZfJx4HA7OZNDY60tM9NTFFuWF
An3M4Jf//vCUZQZLa3m0PNdJgy/cKQrrFBJ3zsRjwgK0QMNT7krAl2D7OuwllSlw1v9tn8/NOXPN
++GtDiWRQzPCcWbuO086uT3r3vqiT9xJ3nPj00bp3gcz6Y3+LKmtwGU0UDluEdbRrXwYnyysgwal
IgsBEibnASMRwgdhguW+3jdASAwsbkdQJOAYn1Z0TcmvhPeAS/fvo4NI7+B6rkxefghbb4X7EkLa
8vvu9Hf1ZUKVnZ8Ja4LpIlKkfY1heKNCeg/jCPX+rl3zNST9O1sSNu2qQk9cPSuDE8KbV6W40qJA
d365ImR9MQXVyrsaaxJMJ2asbfrwQbgRj6t+NurwpK5y1SLI65nkxZlHCTVTAG9PXCn8EUDCpYo+
IKs5ZWZuN3da3mpEoSau7JI9rPs5XH6OQpE0OS7Bvx9Ja/fezoU8FfxUQT6uFz7va9Q0K187oVY1
W9MFlfGSnn15IXe1S4NailA6A07PNzxRhnGBhvT8/0s0DGGPHJ0zkMDx7DNDRNcZuNTynt57IOLw
htL/AptH7RQujk/q0DjGp+/hbu1SE29VEc8vBnAorazIuLxOFsjcnbqMUinKQj/aTI9fnT4SOMl7
3vjypMiam436EWmKBiy44CXoeIFUnuAG1KwoP87N9LOdmfiJq5cbcCG2vul5mKEl4A935APoh2gH
5v6F4DpLiZAYXDZvC/7YGXmAvR1atjT5sa9tIIbN9OdQtbjcEvhghja3NifTEEj3CjBsi3G4d5Bx
onAMG6u3Gxs/18OGRcUSHLjCz3zf1fWXq/8RlxiItXPeptsp6Pdh4+tQtUiddzBV/p2n8sERufpr
Yo8t0gH/KPPgXN+n29WJ+MfpYLClsZoFbCRpa6ij0T+frKkwCSf5YhuhWOeg/4C4F6ZCJqqlVoOP
ShIffExgEtkqLUnYCkQG8DtpoJTNNMNkvfGzKUkmkck3kIMx+ba4koL+y+giry6FBKPNjRu1Audy
MtpqDbVv0gQmbq3S2aGJXwPws1FuOtu3NGDOK7GFKB9FTtO/zpG1Yo+elkhB48vJtff23EdSJt5H
bsqe4Ar7xWmbYxsuhSxur93jDzhhjSeTBzLDWXWpd2VmHnXOq1iZ4wDAI+jFvqAsTGt6vpdNsJln
wn7m8a2pP4jnPvX/CeuboEiUR+m5gkf51mwwLE3SgOyxCOAJG3UDgTmAM3TsEnRKuY1n/WRSkkbg
rZ9lCxKfR0GkOUskkgk3ynHNGlUgw0tOpvfnVgWclgC5cxwkWY4WSlYq24JyBAnHrQrMPBgtk5F8
wxvGePGjyMxOEbi5MLuu+VU/xai0pMTIGO9IfeqMUFpC7P5gm9VN+O1SRRsZ4XJVKjaLYojoQvig
TPF39dycb1TOT2Uc7s44pcLIIaMYB6PRnImSLXQXUO7sUIMK9m4KVECRNRVL3ZjAn/yYhu6/d09j
oXdgQfxmYGXCkdyWyUkxbW5OTm1S13KwL0/aZtzZtJdL9LIvoLiTDXZF0d7A6H5bCpKVxMzRGzsb
bpArOBuYtGZh2bAUBo7TabzeDG3dgPMAP3W42U/V8KD976r2BTpbRkp/dFz8d+PETsZo5qYfZDkF
UZ7iOFIevDHrQC3NOuO6OYOZgfiUqKlNls6LooChxbFGQ5xKf17nwUzhoYJNm9CE9bC7+CzpvpiJ
8/Qerge6UsHXoODsKhLzmQ7EAZ/TUcvvuXqhMU5nNkmlZIcditnjKC0X+JFAdojOwfhGfHtA8vXD
6Gqw0NeAagLyzPt/wE/EKH+TD+H7rk/xDuR88K8P5wjQdNhXXlNZ8OXKC0JVjcv7sqSSxi6j7E6r
nNBnOISkb9E8UubxQj+5YQSO7F262SpYXdm8DmwbH+Mk5+XGUFhNXQ6PyOp8fH8KyPjwiXXZKaTa
Z6e7st9qavJ++dL6pu7+HeR+3VQjKRZcXpW1XB6t38K1cXsgg/Idp1mFfQ22nHgKeZVajaisfK/t
xXX3MGa2x/fbbr7sZcXY5uoH06qX7Bo95hBkN5O2dEZI+mQSlIlPvkQQRJuynNDjDCzfI1sLnYI5
Lhu50nJqSsSIlHD0FKNxx8xESbjSMZzQuBPCyUEgvf5QduCn6i5XumB9z8TAiZE2/RPezYTkQYpi
Cxx2z0Tp44DOmJuCFAZLhgZGqnF+SSOy/0JGBmrlLrROcSq+Un/M/zCfsmwvS1H5UCFeGaydAHXW
pW3xNklUYjCXFwkeo+j6piGHxQwhHYSU29lIqdWkgvGE9twiOuGvvvbFlpu+ln2ZYhWGeKbWFFtG
wAdptnF8lQcXpILZ50W8RnDK3L1z+8JCxrgUP5UdaTN+UmFbp9fJ5+IfZqcSayyAKN+tNyT6Vi20
aKLeFiBU54KTA37T4bXfUwFzuxJIPL4jpIip3KaJI8ZE6rkMMMN51GbDaVMkRgVELid7gKQfX7m6
Jmjn1R9a3oExBeqll403BGy+KD4jU/SMKp7zyOO+q/aQCyrIMX4yha8rjkIJsoD83iuSbWd5AHa8
3URD7U0958e05jAnYuqwfoYAS4lAu595UjjwNWSmG9caa6nhDaXLb5MDynV+OeN9TIVWWHBRqoBf
Egjy2J5tzJ7DTe3VTjxx7VBhilyVZx1G8esfTTQ0Brxdzd7Sysq0R6kLqnWpACE9I/wiGOeCyXOk
mfwKp9YzbjG/CKG9g8jRAKlZ7edNV4VvSXGhwN3S1UkpZOdtI3jmJEVTeZjszUaeYozwdnvKGsgv
eNEM5VLKKWZcF9aLMYun2Ex96Uvd3HTDAdZp8hXm4QGwytrWh9Nw5o0W3dgt1AbttH395rTVyo8R
M4mM0lwZ9C5DhLlLnlGXeE6l2x9zDdhVZFgNafkTB0KapW+U/vnjfuVNqzy4qtrLhbj90z6vrCM6
oWDKpXOAu4sZ7NArjYCCdQUFxo6utP5+3ZIvSj4XZoMN+yOfQk1nH3X0mSyed1+/L+cRt6fchJs9
hM7W8u+4pjcP6jlj8y4xUF+JUmvTw4MBs1yyMRqyHz9FYryINoKtrUyxhwaR4HTKafg02K8d3BvD
KdvpUMRKwdrCrqZgAYf2LgbMmGowmOtS+Sa8sNXPnVNlUaGmHtEzD9Cc1QwE48Xqv9Bz+Ue9cqCM
Pzv/pD89eaL6BtfzNplOFgdR+tXt2N3qnjWuvvZ/pTNYHad4PqQPyRz/27jkjDSa9AWlBx7HLWv9
FUyfz65sbg8lIRQKLuFAStrTgr64mr7rrKLfIh1raymdcncQ1tz5ohvvth0kY7wePyWSDIJP5iRw
mk06vqqfJQKKm03iDq8bDy01BbutRATz2R6ZhPVlVWpy08uoTalvv2j+E4QLmX3sXNx0HjXjqDlk
wsJNmQ2FCZ5Kxdoy0k4Wqy/G7juTIMA2Y4A8fNrMo8ioQlJ/38/hB4IaaCAa16+NbZsbMdwiNQsv
F0THTMsrVodsvUTjoJzINSpp/plMXz6jPsjlbbziUW3ZDhJmPR3qsXkx3Gf9188mqJwQS4E1qtZS
+zubIbnwhoq8SM6bkAVS9gPTRUduHUQFOPPmCz68xC0AowqyR1ZV48Rp0QDT5o5H1lvP7Ub7M/Qb
x8UCV3sd7P+mA4MM24zucEMkHt6zl3hkBOq2HugJR1z54jolIlzIoA2W6w4mqoiQgu9ZhAe9k7kb
1g+sxl62KAl0jHEyvBKzsWhnjdlpgthj5f93IdQi3z2l+6rBC2iKlhV02RzcaBlF00o0f4GHFzqh
Fxk5lFB9GecI4ud/RTCM/HNpjaWG4BSqbSesOrueltVWU1ZvDaYVjFCcGq1sIoUVWuC3tjVmFq0/
rUnlhtS+u2gjEi0KkNeMWvVLGtnNrq7O4fhxrz1qGL2q1XDAbbmLi781gtZP/l55Ac7tV3ZAvZ4g
RKoSPymoeLRNsllg7Tr3Mukqzmst4yG25akib27VJ0qpQzMVdBd9Elc00Lel211KXAIzmJuKY5B6
dueptUfug6r+HnObt8dMUOQhf4SifRm+qyqS4VAluV+N52XtyvQK7rNNXCL2cfuZIjEyfop5BnJ4
tkyhcwLwHeQWH0/aqdauJAsQiWgkmsJbcrrpu65Mj4Kq5W4AMoYKsqMCnXAlyJjjEAezVE6jcMud
pTLP9TttHayS2cf4d2aAjvgpyZBodvOp+HpR/uro4BLpcZEwXT8tcipPUuV7qcGq1vAwisLhoH13
zEVHknLH/7m7CkFrWDzir1rvKPDX/WsxmZQX3P1Le7CB8EpWY9D3qfGc42Qs4Q6gbXelji3P7Lnh
xtTz6hWY/IrSwZ0WZzo1osTGjYotudcTIeEGn+alosY7s6dKjG7jkzQUcSKhSnWXLAbtjzRTKyFO
jvxVD76qz6uyLPO3ZlNGZrwmSPMN5ZVxiyukp7OAG6CCepZI33KZBQubYOagHGCdXYqVTwoSKCfJ
HXBH3grlndJGAYAU6yxwVGICfjX7jr63CXzICVCvCfxEeMiwe7BQevephPkXPYSsF1hku3r1moaB
M6AxRQoibMwRimRVDUzwMVuVe3S/RdZAMzFUGktu+xHITavr4HoL/pvs+Au8Sg7GPL+EP1haLiVH
4+j22j8kUm8rE2eKSspei1VH31L7QH8kHpIXTr1j7x4FteWJqd01m/xyQ4/tDK+gkOfpEQprrlGX
YXsaG/+7cpIIwly010fbedskseqY7x0zubdwyz1gf8vKrFcw/M9dw2iUVlwAFGdE/SrnvYCMwU8m
fXPui9LW4YmFZcRkSmvwKdm1fB3wNVlR05qRAtysRuB1Nfc4E/Ec62VExWZjM+r2Zxf6+mhJ1MLw
U1gMcrwuIGyqMpjUBX3ANw6+wkpzlvBd9Vd5Z09oELsliYg96x3wiHW+678FWa3vSLZFUda7to16
hKdqtK5xUHlsIoeKdvUjPltcVJ/FGlv4vZHa0M5ejNCnWY0Y3zD68Xd4qOcNH97/V5Wpb94E0UIK
Ro/09OorPEX4MumKIlzET1QWh45p3CCoLq4WIIX7+uSmLBoviDfRZH8UYejjyk1FLT46Vkji+Y6t
MiUiIU+xNpKjHfFh4hO63N3h6Gc6F4Q+MaR7hYz77Kvz5CooXdTAlIMTJTNc7XnpWgUUP2IOzqYp
/jbjQQuJUHcZwPKMocJ9S6siLnIhedop0HGpV9KzNXC9OBYYo9w/g8e6qPv+1kjoun5ET/bZwbMa
dkAW6hrIgzKWDx9RBbAiyC04xGo/0RatUXQXr5cY2EtYaTo3VPXjzk3M2VN2Jf4SNI/vHA/pTi+m
++WfunJnz3bhCNjueJbGqIJtBgYtHy1M0A6Ty+J9bYctjqQAcMGPvLn3HwqV1eD7nvXUvSd/sxJD
SMojzYgbBKNo/I5Yn6Jspjh77rXqE79/5VLsq9OEpSDdOhYxRLpfHFi5dBxS6fPxl94fMtN1g3rp
pXMl8qUqRb4Y3YfyCs3gJW56qxdUwviGovgyQZt/1aG5m6O3r0g841pPkh4k/PJW8huCjEVuLj+x
DroMYk/Ph1mZYT/8giy0SCz0onOBIgEnqDPxA26E8r/MzhwpvJPBckhL+6Id5To2qX9s4VMwG0Ga
UnCKE2C7MwukSswxiW+O9URGdFTpdzNn2gArCn2LkYjdNv4RYsfw1PWHyRacTnBpZSW30OF4ehBZ
z34HYKxCu4hzP8ybZynl4JhJuJOC3sO6wJ/MTwZXUEu+ItNKfiOxu4AgCVa18Q+cSO7iY1i1I4pp
3f8RfBTYl8KHl+Gb4mFzdHo6Lt2QVI2Vq28Wh0MRXSI9xnqqDnB96I3gQrmX1xdnIIL0llpg+I7j
j+lrTWs+Cd+FrA/Rqn+QXV4adLimFwHa2MrpuQjcZkLHkqbUu+ETG49WNEdJ3VkHti2dog93AfbS
nDQriYKyEwYClSquc5o8coush5ooYuHS59TgQ8LUL2a++GZmDVZjdj9mYBUQpj+wr1KKas7F7c01
mxtSqcgh7xVaory9/ycMSoO8pROrfeLagUDDhhWfBeQ/4aJN0CkxCPU4oTII0Q6HKExLP9N3thzW
C//mGTch5JChoGfhiBLAjcDQcryMvEakFmEBlQrDkF82mskKdfM6TFzEeaxt02vI/d2bVLKU0E5T
tG8DJQGVI6sv+QvpBXv0Ee3mwD3KfAg3KVpRaCxApKvktNRMPHehjT+TqROTIYSWU77THYr+L88G
xNwEN8fK/Qx10sMGACrVwknOKq+hVXenl1ObZ+BGtMWcVTHSVG5Ju6FlBUzl8+fvo2HJdoc8a8Na
iFs1XWuP4YeBDCZvYTkEyI132rDtt9XWEa2L2Qn9m1nmdIJHiyI1334QdurkbCpUGyNFd8gFssul
OCgmTSB4nuWwnUI64Upabu21YJCFuWjo9D3lmGMhYs0WToQuacmYwwdc9vgCYXNh82sCCyxym7Xu
CHV5Qz17h2lBMSVIgeAo0mljf/GezvSYGh/l7EF5nfd084YjxgZr6CkB5lb0k9fgH6M5xWalyZtZ
Wbk7/kx/b2+cGNjdZ/27Vn9eykP9GnvHgk0XbvC/2Iz+eJ5hmaPfruEPqSZSbAeJGXxN/d26jzsO
RnWR9J15CQyhPOLlRDdIaJmLHyDnHo4uLYb1LZsBSNQPUJRvLQBf0ZRIVXNqoLWTPr6lzSJYb1kM
wxqbWUR29S4raQpDe/tkEgUVYarRrh+ztq05KdqAtv8Z+ABDN4gIWMiCoadAcFonJNU/WcYlfY7w
YclJP8hoF49SZWF8tQdPSiS3Or8VfPYsjRGWl7KJb+/YL7LmIIpvB2ehcfDLO8H1whnzarbWrki3
enfsXQowLGHRIc9FjQc65BrtWwnXiWslbG3lDrRiGGP161YC/lRPhxcpZlAfgb/7y0EYjpPBcTyP
TEMkY3IkjRsRaShest0tMKrm3ynsJXOjMPMQvjVNvLFiq7STOVnYI4KfX//pxWuJ/2l59TqsFTCU
2sf/b3u9DsgVDY2jeGAh1C/+mCnFy0GJgWesL9wJP/qo6ij3DbKyxVB2oc17z4hoSvwaj0zNHOUz
OInu1gECo6xl+uVTuSzXJ9f+Ac8bTqeZFdZIPVOxTcdhfjTlAwXadrkkEBbFN5maqZaqoUtWVZOA
A2AEe7dkbwjDcalmA10z0jlpUY4IH3a3uF2GtJxFjgUu2NXHw4mIlsO7pfr/gbUSgQrhkDkN0dFy
Ry53PdS3MFNVLX4wA3baC5GCTEy2uJnRQmsmxbci9i2Q9L4O5Cq2qic0EaSCZuHTjWG+q+0YxR+l
o0GjTMOu/Exzmo8VT83mKwxNgr/Ny3AyQCpdL8Sujs4b1q5vvPdN+JMIhRKTblSImmFQgti0kvzc
ErKU36efSFQK96FN7fnbOlLvhn1e/qGsCuuq3CMIGAYAnrQosvwKxCUbMcBShhvrix5ajlkaT8J3
ULq5EaesDt/gR1hBn8s8wyHpToNUyMt7aqv47sGZRXYzkVEIk9+GW3NMxNvZ4Fy221LW5BrMNeK/
Y207ACXuh7RP44doyTfUD81m9LgjYFcuTM59yPNc0ykuRmHr36zGuDXBTK9nBkywmRMtusH8GnL3
E+MFcVOJ+V50pI2uvFxkMDrNUV6RHsKvhVBBz5D75XazmamPdxAoFrjFQ+/Bb1Qm/x5FolKjjEqm
KcChS3UF6J251QJB/86FpK71F0SIetDSc5H5hW5+pUeeNxhf39Xl1p4JbGLlJ+Sz/1ARsLzlirtI
pjuzaxKNwaHh/UC3PYrqcfDnR0Bwe4w5Zr5dchOzkSf/81AQSp8XffXkQFladRisdDOMYXdDrTv8
QlB1aMrAp+0SWGpSCkSo51zfIn/APA1oIlDHu9bycEjAggZNoLt/6L5p9fG1acxhhOpCMl+UDrXw
TbXriUIR8Ay5xJQY0Cab4JNlzMGS0WES1IzjcsdOi7D5bc8Rj771N0kk02X0A+76p68b4vRrIilA
xEnl4S1wLitQPJgg97P6nhiu90pPSO3K8ep8Cdz1ukn+aVJwSZ/fvobEfudN8xXS0g0Lw+nEcgNq
F+kY1gAB4H7SsMptg9Fhm5Sy6Ff9LxlosZmO7PbO0vCUQntNRHIopHVB+qw8Bmv06PJS2ANhiWzK
IlJujhTLXAVC5BNX/oXqCLNmGkkycDZ/xR4RHMhOdZFXNEZU5+PB8/uJm0VNgmqxXR2RtA1rKkpi
hT8xCuFo6V8CPHxlgQnqgdG9lxYd0k3bmdJYCtIxwF2fm6t8yaSoK+SYGIbncXi+UZyPHY76yDnC
8g+nOCJMJxPx9lX+4uwJgWkj0u9c/4t7vKWgpeq06gcFkPFu+a3kzU3QN/W9lfGUsyZVfssXz/SY
L3B22EWjh5j+QaBesQTq2mqupPlgD4yk6RL7WM3ufkuuVEq3wIwTzZ5xFwLZp8ckxmNGb1G9ze6D
7f5axUL2u1BW0x9Blne5gHq7h0E7UyF9Ocb7JMPY1YECb9JDPXx+sGbU876KBamLbP82uuRhmTN1
z0YBFjkSi5KUMl7KNjQUfBlgZ74Elmec97NEawUeQKV1W++E5xEZFJqtOE+W4nZNd4i7wPjljhLz
LFElvGQmaBlZ9ku4ecXvnTsucJdfnW0X/UrBrRUn7MWHIfzeSmrP/ad3CYALOlK8LyrQlbOQW+jM
PlQsNU2EVtIb2lNxUg2Q+GQ3MgpaCKV/nkKdYJpdxA2QyZHkjHMXfX1YuTYQmE0xDS/8yORO7MAz
JnDE+E0w8wOA5CGOc/dRbK8a+MoGiVANC4Rqz63NR5Z28A1qhx1mLdtLMGKWo2FKEyCpyrvPYhhH
zO6bhbMWTNwfLJ9gRxtqtoNO+GeW2M31+MxnMt+xOGW6JWPp/YeX/2S45rowubkV6D1rjx/x2wgX
U/JOPx+27lYdxAZ5N4+1i1ZDE2HQacIhnYf/qFT4wEQGXWzUfqgCPnh5O6sUZeViM+nu89xNex/Z
bhwJovERF6QV17ZGIKoxhZxqr36jVbiiAMpsdR42t0fXJ4OhSKCsHn2ZSzPaKJru1rJTOKzCHZ3/
FadBw4eDiZ4Ify5tC9ygE39hVGVWBIAMroK+B9huNVQCtFMqTE05X9DGNHsiIZU04C8rAMMpyfgw
+NT4W+5ssCZcKahobIYnUjemP4RVVUXnS8aTIr30DvTbdnhxPvFMTudA/CQvn2zTnPNqBOtQXVKJ
FXLo1Dkh7R+0r+bIVcxxFf5GxnxWM8DId/twACpCwyZmFxiICBckzt58674kE+PS53Yu8XNW0MHN
b1rWZ68sQvCJHEANKNcHIMuPMKe/6h0n8r5PBgALSarhLZC7P5THXRdWkdiHOaYlBLatcu/5k7wS
5ufIXGgmkBTWEl1u6C4SAFJp/iNkembUlQrvgyBi+3Q0y7w3xCVrUX7ldFeMXNRPAtogyFTjpRwM
dlu7tGAtxXyYY7cY0SzMz/LLNkPQaQKbAbJP/Ok+RBqENAZH+p50PCa/GSQBQSE/Ey4pwtxgw0rR
cH1taUbw1QEGKPz+Sn7PFiK1iOwMItp09TcBMe7vsMJM1GwYfZq3uGPy/8G6hZrYyppdN/D8b9c1
OxdBb6QCGp7QNtfLJpKH6adKCEV5Nr2ff862pmtC59sR3dJFG/q1IiaC2OS73mLukmzmV1aS6lAx
Z8t1suK3StkouTqO0R30yeroz8mBBh+Na8rfv2WR1Egqnj5iym2DnltW/wUH5XhfWmS65gxqK7Tv
KwPyzynyMfvHcqkpiiLA27sAhpSCpQSlsY3GwNQO72yDlyo0sfK8pqlTna5B4s9y2rsFvH6c5tvY
Sb6Qr6Hh+0+5pkc/Kdke5D7W9Yhlmfp2KBf4CcZVAqlHB0kicLTutNzz1y5GXYCcYZjDkXSjCbEs
ikyD7StpctK325UxWGsm+60dVwrQXrKwOOQ2oTFpMQPUcJjGgkC8ih+uI/sydDrwhmS9bOZkZKZw
zUeBar2BT+nBZ4Z7wNQmHW4Wa3OLsnArXZ+FVh1RrqWTO60c0IX+gem0yM0Mdz5T75DYHYRVWkoM
H4f+KBsdewYqjmoZ8LAw25YLZHDuidHNcNqm48poV6vsDalPjkphhEgit4SXn2Nlr062Uq+X71qy
YbwOJ9dGsl0xIvX206ABARAZr/ukwN2kiqBI2PZ/BYFgoe7XHeHyEGpV0OPdMDjIEfa+XIbISCPq
ebtnSMjaC2lvwKxHkLSsiv24YocYPGCffwIUwcp7lE/BDeYVflrCeiU+AAmTaYVfLbK1SXQrsJEm
6FeQQ+L74RnyMg9+lHzCYHto9ecF3BfFL8MeCMsKCWluIChwP2B7A3JMMjy+oYRNBS31Cvv/EKSv
KJTjiDsMnW2OFiQQJnufOLLp0yKXGEDdxgasI3lcG5i9PqELSzwyWJGd2znOK21U1wLXR8OQ8e+y
ZaPYt6z81ejh9Qd1EQX7mJYatnXPyTMKnRkFsYqGunPeLYbu79qOWIC2CLJfOvwe/52YQ3Kd/8Lu
LmwuLA4GNTbypZG9wsSGPfDR91/VQjCzyqK9uyJgawdEYLxDnE4QsUDnILDeZIVHGJUUP5nkj/EW
tGH15bb3KcnUNG0ww+Nn7nYdfoAS2gZFlMEbkUOztOPccSQB3CRgosNvpKMtcLTXKOHb7KvHzZuF
/HWjtrCGqmW2icKj1N2tedIrPT0J8801jkrIXAcFx1kQ7hihezdo3Uz5Mhgc4kgouvI7UolvMmxn
Ia1qhfTuqjTXLhvh7oe69gJX14Hysv+VqScikmUFzbXYRWr+Wnhcwhvfmcda/aHkW8f+wjKAFsmx
cb4LUunJCg2piQ/ZD7emhzSqwfmO5mkD36IpiSiTFuMrksWh1M++e922YxmxhbdYIjZYJhsNvshc
CULfZCkyXiShaTxhm8STbBxLVbF8IKKL8Ep3MXtVqowdH1pQn/Q5WK9dNRYHuqYghDFtJZeQHeNt
IXPIZGt8FTBKPM+D8D/UQ8+Qj/yW9poQACBs414HM6wy+uFbxXLpHbYZH8tzP8mjtE6f50mkx1Wk
TLKl+cq2t8djFf5tRlv3A8nphU9oi5xEK60UQqKinybwqjG9KU6Xxxq8euzSOpQbf4EjdnZDEx/d
I/AucthSMytIGBBaMft9L4K5oSpHEcucaoL/YekqqafLZquKKWY36WUgE/wyzs0hW1gTTJ5jISZh
Y+zfQuMUrKz1HKODZN+cqmZmgDqbnYmogINS0FyrtaU4+k9XpNV/boTMPqWu4ephb/E9hZw2+juI
KLk5nK+WbBZLHEXlYDlC6WA2qJgP33qZkwaWbLbaocp/FQE7bJqiQNB4MtB7dKXrqBPUPwrOi+fJ
+FJfq1unOh+Nd0QISsytIBgb7qJIOzWsZE7qSdtqbSstrfkHjngH+MqjzajaQv9qG7u6200Gy8aD
esY5WKOiZgFa+ny1sSdnm84jBFzhwxV+bEoqhG1/+JsHaMLky600K8yRImkFcOC3blHlGPn7ODOg
PImSSmshDZSwgSz0WTFE1x2PaHD+iDWSD0oFcOzdF/hpqnOr/i0nBZ1BwoXASB9mZcCl23riNqNi
MobPPiSn3Fv3dWe8AKU2cXwwx9ZV6FSnLHeDSfZYh2Ciow5sLFwcMirQ8RvnPP0aY9py6EYnvJqf
/4fjjdrlwNJ2J0XAF7r7+urO8X0zxPqJf+YbDFkAxyv0ocyLox+/wUGUyWHtCJBROkYLqGG5AqgM
xumI7si97Yrvtc+IudtMTMMenZUSMzyF4shN+yPhtjG7WdEwbhX/y4wEfk5MWlpQicU+iNV/orFI
DLR3C3dHlucd2V49cCj+nSTtSfPbHjD1wQUW8CoB4XM1XOrycf/9s50wQ+xqeJkAm8oLMDtToYks
mgr56f7BHhS6AecPsFoY4OufthSTamOgfB/aAEzqJJulqMRPQzpw2EB2HHJvIVZljLPklrRrU/mZ
l/5TIPufjDQFMU4pHNGgw8ODSu9DbPfHDkY0xB+NqeQtvW5Pw1UHnKPgJVVUpVYkg4JGZQd1lCzc
XO0mbN0ej2OOiS1qHaoc2m8CooZz6lW3E/6AIQMKh4zyQZI3d3k36sbsSkrGZfelYMvtnokXGlPm
31Y79eC1bb+fh/dms59mU1RoHEUyXOWTK4ownhs9uqro2Lf3wDhctlrmNknoD0PB2KDUBATwf0wi
m8blaqnrXkdji//Yn9io/MsoNo/QtZGCa2wcPSzhhIYLdkbMY7OC6tfnxsHMA37sl2SG2VloXLWY
AbP5CAR9SGcttRhozX+l5zpg09JPFfo3mv56aZL6SaC6kTP2dSzZayHxmpuIfYKSnU3VLtKd9KC6
0E+V6PaH6btbhNVMRqiYesLd0Bpz+nRsiCGoiIhk2wnAzl5nElFl5sNZPGUEFrHfnvMf+asvYPud
Dze900tSbSvZKL3BmPXJZo9i8Bo9dMFaluf0xPTaf9beefXaRcIufI5FIeNMnWrc1f0qtiQlcAiq
tehErDsOkzkwyis/liUk99C+47jJMhCkOm9QthkReQAjOI/EkHLEGVuy1M4Lgk8QrMV7jWS7+9cs
WrubVo9tmnP+PFKnCJpAzRv3GVZ5hnqsufmzL/XLDd1BO+/tS/jO/QThZevZPatXNo/Qvg9AxUhj
7Xc29LchrU6zX8tz7zd+mPEX/RY33JIAeD/vK3yNMYsEh2BUHPTXcOrdIUmVE9Yc8wFzTHLL+o+z
JHWBcWN9z9VZGT9+zSPI00rIY497BSm0WCumf7uiNN225ImsSPBFO99R0HpafO26O9AV5oJyEoBa
EaGAfWFPSrX7ggOIj5FkqtvXQLbjrVmpMNWN9Jxtd81PHjiMlm5RFudbpgV0Rz7m04YM5E4MxB+5
gYfmvVhcKusqjVH4F7UJperAhW1ixbJcHmDqM3D6/v0IVdTv3Vtvyy/RugThns2TcijoruedLtWh
k0vVnb8yIUOAHQWOz3XXdG3yTc42BDT4a6VsaF/a4DL5p1l34Cs9GT29KOnLeJDf1cRTJSnhyHjm
YjIIdfpVqvRFxkWEVu0FFjLkU5kxtPmw0SerrjX6vBKhtjd/D8WK2N7/pCnR0Vh2rETGaidwdSok
3Y0mLfW2e+JBaVZpq+Glwf1t4GLTadpCd3Dt55IO5QlW8aq6duOlUjeC/qwxo5DVcwgOeBl4OuBs
yHg99rik2xifX4M42fYAANAPXfnpyHKJxjD1hLExPh+FA9xA5eO8lX4IUC2wdDQy0LiDXl1yNSyi
bCtwQCeVgzgsiVBfc+gwNxp2e+LnLcv7rWYLqkY1mvQ7Tnw3i9ytpArKYN5aTSDq/3I/D+qsyWCO
nTYNfsORr9XjoN6Fb0gyOCAabgHwcir648HaxQ2l8F560PwDmEMFQlbslAXwFB47FS0zSs6ytVqQ
WFXkfkrYAI73aqx1YsdfTIKOb6Psb/OaA8x+jYCWbeZqKIqPojJF9ivHEvibDMYUHVNZLBXDbV+s
j0uCZIaIkymA4AMBOiuFks6J7sSF4A5OFJp1U3GyysZZ5cN61IIWsjNIyjfGJCjAS95lb1MjPr0w
Ahdm8089OFiXfC/78UwzIPQ4oRXPMB1ZHvb6gzPTzt6DHgbAsKjx7OD7bT3PFj6UikOvN7bhXw5N
2XMk7PiS/JksnBOOp2wM6FJpYAGtuBTYHLxUvwF5CUYdUOHoPVJefonLn68RMDJPSMGG3I/BBjmp
lHFNehfNe0exR8q3F6daRn5BYx15V3q3HgsJPZ5rVon7Dcmm9G4ES0rE4OGsqclK0r/nT3FaHPc2
Eza2W3+mZvzIKnF4jCp1xvootBW4cMBF93x7vQ0lJwuGIIV75eK88nY+Ghc3mZdqtq8kkWddfc9W
JHuwnJZbaqt+LryBWnyUVofUamPu8NkZGhv6UwegJM8i4uiuH2nV9WP4ApVPDjscfkcdBxoTXBZt
n31dBMgrd4u14mdJhQm4djo8n8NCEqUfy+4bs02n/kr/2oRLu8ZnC9vwi3dnn6AS5ikJGDfKOr2/
GrQC9oN+C/JsxfoW3PGSG7+umlAOxSIpeuM/hlchIxIO79dxtjtCYcYJl6YZnHu5kSJsH48UNE1e
2cEmLkYOQ0TFl4TyZJeeb0hgq+VumLIGNZnQvM4fuT+hq2knwi01ZqK/OZD7xKagvg00j/D9eI3E
Zo6X2RvbTDW3Sefu4XHOz2RhHLzNNMjsO7aBPMWnUEN11WpuhngJPavAYCR1dp/smg7uXuYxWbGB
fXBAfYYFByJ7vsg29Y1/SSwZcBtuqiPtdj07Zd469p3w41AEaOPmpM9KUjOJbnz5wmBM+QCxZwBm
xADH8NZTESU5u6NG1QxlenNZyKM0QGCSY8WUFn9ennnXWvfVU443kJlhakDqcNb9C1KKoQ1k/o4T
1TvtLXf400lnXnV0hpzjtV27dT/L+JN7xfrJjqezqQkP5Bae9pQFFTO5jREIN9/h0rAx7xKdhN8+
Sy0Je6l8IMXN6aP8HdlndG619/iYCbuAtSx+TMxw5QYDBmuLZzL021VB/stOwVJrlnJh0FL6igud
sUuEzEniPk5ZbBlWXBTENcozQiPxPXyKZuiDVIasztiQwIL3OjW4t5/Sugqv7u9zEBvMlBHJbP/h
ItGslkgFseI/E4GqS0hO7ztzw6D6HnolxiiPynyH+kIX8tRl8LA4o6k3R+XdBfTx597mBLOewDMS
wUgEE1eFtcRtLs839T0+kBOrjjhS/HC3U3pLN22nLNqP9S2uKWD+uu1u298p/AqsAhZASva7vtbq
BZcCPiPkCXD12t3mJt/5uv1y3N1w//VGUtEFFcD0OTDRpqcVWtVEcTFVFGL3dShNxXuUV1lGfGXj
MKW4YyO2zwTZ9m8rSzUkiVQeIPCW2BFkYFQAMiPYM9qBGcqE1Cbb+aZqmE4y7mrcCubdZ+pf5BVO
Y6gXyOSCCWja5KqchONh4RR/XGbqFXAoAyFg0yNdukCUrhidl9C7BXB2ryElvM/Q2QEVczE9eKCp
cBzdMW+IxRDPEBKTFGO665qIDgKjKJ6OMV55djjWwOkpbOUmeVSPS+b9T5hD5yhjSYTIxDPUuE1b
M/QHJjb3bwmU7RGqA/hDivgJRdKqWzMSviY6TTlBxnn2OadNeZtzdTLBFtsw7yRN+O0F5ljB1GJG
R1V+YdZycQkSUaoOFJcS+Tb3akQEfHgxGdESKcFWnzEYcKh652/d+dfDnfu4cCmciojU86VkKRVD
nZOjIM7J2efR4NFTPwGVzpjU+y3a54fTCvG9xnZy/ZWkwZlXFz3G6cU1fqhy901fusIms9Fyk0XJ
QP5hoNkMI42oAdHL/dF9bwQ8B3zJ3zoW29az2vebOROBdylWzwI1q3qdtGdiaGXzIWZLiW/7qdzy
chZJqQpClsU9jDUDA32NTx0xbT0N5747RttbhXlyBi0vdeLTk8KUr2dX6DMygLF6IksrSbHnGkXG
kOOHuRPLe02cu5IcEkM9o9r0SFfHnHbHII3CfepJOI2hRbhWe2s6n2Q9CHA4152pE5Pu0A7XuPmx
+t5c3t6ZGD3khCUd0j6lswKDj2Cq821OY1myK9GUbDCC2E49UskZgRq8s6w9cJmk6xGZWcwPWsrs
I44RQWlAzTJLRInz/3zIvwgDlwKwI6NQUtvznp6ITrlGhZwDZ68DGjMKUtKD5SKQBhLjp5n+nuxi
l3NIcJAhkSvQZwm1fPGERdolOQpY38enToDRF5j6RH+K1Y/CZi/0KTCArPIADvdDs3X/Jf9dBI3V
r3vasVbe0pK0ukYWVBjJXHiZxqqPy1tPSBzz0HMqpJJFXZrqle03+bEYqVat1/dqIpL+q1btY7yw
8nQh99yBn1cJlHRaCS6hcc212fGsgtJtKwTGQy5eZuTKEt/72Qxvh4EbXO7WGjuodDTUa+Oaay0q
FubW0xymZ1lI3Uq0BIvIQZyTGFU9FuBe5jPik4UWLUs72aAsd2K6//B5IF4LC8k+jScfuib/Prtm
LyWc2+OZaV74fC1KmlEa4U0/OV+3tCQd+PGZFyHHJZsTGCNZ6wX92I30W4Bt/GXKvQWSoj2I/y50
zAZjyGMf9V0itnDcshpl5OxwnjqX2jGUvAVPiaG8AdgoLYmfwG3GrFNLqn8fO2e0Ih6wDYOPJehK
XOEdLSi3KNe5QD9e54bHF0SaQhwpxSdz53ncEXEoma+XSCJp0SLHq+5HrRFBAlNEmv4NwkgKdFNR
mOCy71XRTXWlFqh6zDrEsYjK/nZddwU2pLUu4E/SmgFJHR8rZIp5BKGta5NiWLTIOOYnm7sgoSvn
iQiyAw5yxjq2r0XgzRFdY4W2AedzsSyLw8jGcPWOj7VqgZGc9sYQ0Py1eEx24j9RF6p4iFmWOr8l
F/sESrfADDX9pwzLTeGVVnHcmmfDTlfwGyissZJCZ31Agk8uxEhhcLZ5JiAtHtn+p4NCeFIj4ETH
1CR8is3J1GMGsy0JqIY1qdCgkTu2K9Ncw07wGw2Phg9zTIsU5l9PdtP2eqZP+pBp16Q/zGoXUxsh
zVuZVoYw6tTswvLGsvwIYayoC/wSxQnHYDZs4mGsUYbggHVY1LVkfp/pl6y4A61FgKq+PIYh443A
Cg2LEpj8Y1CxcampGyUzyGpzFECECLoyTeDQL4ndcLOdgav4xMkVkh9saXNfZvZQ20e3K7VBd6iX
V8CYVqvXU+7wSNyZV4S9ZwTxN0u0nKFNNIGmqGPBq5f5OkGQbYkZJbuMAzkHJxi9dATP4ATDLV0F
9CE+A1FtmLy1K+noYn4sMTKfzywpEFFhM+DBIQtjmskh0X5ZdsnGCRSW3KiN0NDZ4el/RdTaZBfM
YCv8hg3ImbEUY1kgx2xEsoD8qjGqyyilEjvMtmDdrym+UKA6PdfIVo1otud1P5hj9reQqsK/qCAv
Eu2UzSTTWBKLCdwaOyLM+0cwP11Unn9krzz/bZwRmoL7H8Yq9J8z47aKDx2qNMZLuV1i9XScWf28
qGPWcujGN0IHHWbCZUcxFtQxVnrwmCLb5clnIaIWCzCI1hD/FdlUBIgpt/5efbxl3cl8lMNit9X7
ufxpDMh4gpjOfHXHs7trixCK6YJF5yfGr76kw5BVGXBydpXvoWIFs0hic51cGAYphWhq5oZwUD6c
meTV+7LPo2bCk01Z5rZvheRFv3npJR5mKh6UWd780JsUFiTFWF0WsijtCfIIHCXbtIzoWSNYNEB4
Vg5agDoDlMwJRXb4SMdn4zKiiPtL8hhhWa025YYfKjXRmozohkWqmpSN3HNuLeqhQ8tQ6HcEI1s+
7EHi5fAMCnBJuOlNLZ82yId5uVc+EW39PXy0P29IXT5i+ge8mk/V0eZbv/khWX2fFTv45uc/9adi
L4T+1wIdp08Xlgbo036LvLR0NhmAtwcK3xaU1DkLowHOFYLTGw0up9QBYeoZ4fLHmdiO8rLCXlhe
1s5bUbfnku9gKd9Y0jc5OYCrjOJjMwyMc/1k2qxPvtbU43CohKsQT8efZXut+U1o7Hb6lTdpeXQm
7U+cukRPvE/36uexN1D9DqdiG+LBefFOLccf8cua2RcEWJzGayaSM/MlrlEI4YZXkuazs4/PqIMZ
uU5e5RecJxBcH/u4tgUk8YnLKL2drFhzbiSQrAJU5xwtAMk6qh8AETo7ThbDQq5zyG6UV1oNp8e/
jI9hn+anMvXn2DFsawmoXyhdS6YzLbXoQKp3XUdGPSGkHMTHumiqzH+Ochr0eTONzvfYbSgTMNx/
y74Hiq/GRKSvpas8HMquXR2JCY9PAlSq8sfGe4HxtToWU8g2pfoazLBp3zuQvV+4oaGxIUyGaFTI
9I828lJvaF6GGxbZFc07bE4YRz/VKjSdcqWH2kw0N9aCO+MCs5ZJ6P3u5xJ07Kt21QNupJxvtXpP
i7GNuUI+GwqdRUmQAkPQOZtHWHx46NSvaIFCPdtcFi9NmUA4WFg1s2YnraKDJdpEuFFEr8zyFo8v
55FxDBM6Q2UfKyalGwjDMW3aX0dBR7/bJl3sHMr7ENRnIQVphJYzib0MJCndLFNUce/jX7Ybp6mY
y+5DG8VJz6z99Sc7zfeI6hAPrK8ouy2MkM84zccrGm7M3wXRLEDWaE43ngN7qKzLE3XNeFzJTZnJ
7CrQIaqBzLzw+jTx7n5e+Jm5e73g9M9TgTWl5kH794puFX22ujz2PRjvDRnHgM0w2OFM+1OzYxjm
GNvUsPlZHRReZKrmGKD6JCMHSrkFUGCSs7xrJ8yu+glFNenItz2vXBP5G/NfdkjCaL1KYLts+xqY
u+oSAaDnHEIo0j5SMrOxJ4cNFopDhUdki8tCaHkzZrBJ1pXMyDJ1mWr/kHpjmb9Fbcpsnt53i6C2
XgLFdePEikrATIFmepXq4hJN1qGVbSA166zv5nokKHbt6byOJUHC2SsI4L6H79owfYpSoO6DUSaj
oLz/W0tu4bSRX9AJrmzbHyGEiFsjTxDAOtdJaphhmgSUwlh/xiTaVWCVM8anTuZ1c7i4x4XW8ICt
tes42rmNT8Z4biiIsAP8+ksuq4nDeoxUtmVzvJPdcI5aNyXdXwDMp9QouVt9ZnB+WaGfn7QqGYKd
neXbFjebTp11ptxi5UDGeE67H1a4ohRbq3myKYFSlFXMTqvg2dNT9VKUy580VaSmX95ZH84zkrr8
L+35uiXcUvgwRk27nv8HBW9kN/PKw+6Fqsp/+XgE4As8jeoiomC/Ey4+iLS8i4P6O12k05+MwnWf
WgboeHQeXKcBxBX3jlP7kv6MX6LCgfBtOB0DzWJWW6TmCYkfnbZTz015FAs4EOw7KfTMFhhM1tWq
Z4GikfveEkHwTHfzJEuxmwe76zJ3YGXhkNvASoMU2jR4JFMs1v1ho+R1Skl7mp4KexjQTg9JMRlM
g/F8DLhiyekpGf5LGnyPbrZvgyhg4mm1ZzWvEQbtcWg9M5kPTITi4pXrO99T2TsRK2+x3E1aFJzS
qqo58eX0LM2U0hoeuvjuXFXeq8Y0MywPcZUv/OyFsf8pFJdPlRtAcfrx2VWUDguSBp5rnuaVQWER
4mDnOVnje6fEFAzmgqovYJT8LbdN0gvPcKTAZdigvOMdoq4uVyHh7l/1x6JDvf32nmyp1RSFftzz
3PzAblVGMqBpeXhM4hG0UURBE5vX6T1a/044buUl9Co8w4Fche6pq8NoDE22u9/P/AL6M/BY5Cyi
MfD34P4Z7apwIsNIGGj86phIt3gimqfjFIvbBs/+Iz60P4rPwOOhYliHZbBfakJR5x6x6ccaVchL
ZrIhx+qquLv81ayXQgaUS7B0GbXwptGTxY6hKb7K0lpgChLoSbQw704xPQdJ13NDSLvJVlczIqiS
sUALC/TowFF1++CtCXKfEQjxuTD7k9NiuQo1RqateU7m/pB2FaaHtpCEQ7vMlmYevrJQb+1K2UhL
TqA/qoLfK1xNlDISHcZei+nGZdLLllCXw2zlzgwLKaZn4h1yGSpV20P3vJ0arQ10HPMm4lTCtrIz
BAyf4oKacCondDDMLHfp1O6nAQNGQ2H+gC3iburgjzQwuRsj+ZA2lfyApbm3A513/jw57oUbU4FV
0tAWR2Vb0vLMap+CURWiTuPEjbxatJvB883LSxUM1ktQjd2ecqt+vWGZXkRWQE1sOhZ6ydDt4Xl/
4IYwNVpqH8Y7wWB+MW1VL0wDk8TbqV9J1ooIUiFnNj2kymXLqgkMYMXo/Ij8SOAPFWQFNXskRf+e
e1wtsf8oK6dQkekhTQqopNHkZKNTmd3REqSRelfrl03ysvu5XG7nRtFSbsOweSBnx0zJ2Cd55TOz
7XOOnjVycjz/Tnr7OmQVmdaaaEn9Qq5uJDxpQw5AmXZOxmM+X8bn/WW3a/4xjpMz9uqbh/WSw03n
2U8x9AtpAsWBn3FqLEViBMonQbRh0ur7vECRVEAPV/MmcBVQeVBxduuQtA0XkbEDsH6qu22nCUGK
5WoWdxruZcoVKe98WhuayueVrFzHWDLd7SAHHuHByN+awDGyPZrRIx3T2tjT23d63jzMBmgcWATi
Im/SJukdE2pfqu8b827doDEtEfDLWdts1gdx10RWkWi81qC+w387M/qalVI9ypIWSmTSh0y4k+X0
FcNftL5m211M1Rgf81i6hcLLlOqwBP80T0NQrkXKEmkEMTk5A3gXABKDLV/Anc5rKQIezHsuu8KT
QFIiy2YeZjhHgSGYOS1JUuR1ReO/vIbSSqsy+AvWyuXC7ZKAv1d11A8rPq4+CeSpENHoRUFHkxrs
fhlkzbQ1MpPPbkyCm3dIKlUZASPjfmZjfQVw9Ve+FcI6fT0Ct2GvxxuIx3WLJ4+Tx/cyhFFzU8qu
C8ZhiAuQqjOfw3DfA63/1ys1rAg4XHEISjarlK3VNp1cotdavAugzreucHLUi8p01ustej96Ovr/
THaIOsrTMpgqE9E/dB4G2yegWFgWwAGODOyfVrIGUEAi1kqxJJIiUwqfcjPXKNskZ0IhkxbMstBJ
uKf3s1A9pYThyujJYdzzRyS7Yp2qkK74Q7vlA7vdPZtoUCZGGvdwVn9+3d/P4VwWpayy9AffEcNE
Ajdm8g5mCIOJPKTowxvHIA3tPFmqCakEqlvr2laMOFXo32Ik8FG5o9TKLvOrocfB4GT9xjq+gSoS
Ug7IwhdUv6ZzhzY8a5T1vnKxpDnIStp6G9tZfECZLqQ/slRlZ0ZcP0ejFR77Z4iz4F7q7mAV71EJ
KHf0DebALEqwSgl40jRPuhxQ2E4Eoox1OEM5wx0g8AlnpFYe1HCjUkEJPozX1S1HEz6VT6RUJp06
491Wpdj6yUMQbiQIqz/7oYrffoNNJn0OsR7c1Lc5JO1RZ5RQf5PXD0DJkqX+Y++89k37f3EhAyWp
NgwfuHKQT/15+0/j3Kl6YJVnQpgIfLnLzImGZHIDfD2Ez5eI5CWsIXwxz2vh86TJ1PgNJNOiy8ZX
CmVfKXKTxiHy3j947AN6rRIc6kRmtsJWRhMIRKfc7v8z3c7fY3UeVZBvv9C8922a9y1lY/f+p69E
rr37rJp1KriTxturhS7g1ZQpWQ1ZU3BnbbDS3kXEb4OY8ZnlMbjyPde+735m14YBV94F4airGdr0
2boVlVEX3sD00LnMabQ7dEtnByndpLfQlKvih1ChCPtMuIaC8RXl9auP05CxYif/w35BYTAVB+sH
N9S10vnPz9seNl2+lBqNGu6oVwE5dn4lzAU7AMOM7pdIaoySLp1Qy0hk0NNWdLsegoTo8Bm8QJi7
Z6A2iITTGKTZ+4cQXEzGM2vGJnuoRrE30QVY0/4OWHUmh7sQBRKteqj5bDsmcnuTfbWk341J26m/
GhUR4ACZS+JgKyOT8kcGsEWhxWfF5NdoZbLOw6hAnr7R57jPEvpnxsuHhnbWIuMgcxHXijEtG67l
PUWEykSq25UMOOJrVEKoAXotrFbGbJpas3gtQUGH1Q2Ysmo8/1Llkv25DE2UZTbVnh+jHx9YOSke
wqxGKjTcMBip0esxEvXICBZqsitA5HmwSybwLf4w7gCu7xXvSyq5UPhN3ZOORYWsXelW+wSnZAvn
atZwwPAdEGHrA6CjvHjRWPR42tBsJl00aIQzbEQ73lEwAin2p5PbbSdJp3/3Vm0fTotTfpVEapGY
5ALG30UjIBOTg98MTHKeSDhQxj0EM8KEyoAgaa2BsSx3zT1RZMrIJQDz58euXYC6vwm21gAHZAso
5QjDgzzJguSblHxloPn1+L7L7WtY9ENa6PV7iJuzY8rUbnuQw2iC1SvoDgU8vg5x74+Cu1KUQCtx
vidfosz6g0eSQECAhWd0JCtqsv7TVwhT5rIAkW62pyVHqPHQfXmmT69bNfX4Leiy2Ra06y+V4A2K
Gsnvrg8hqHTCPaHHbKlDUR277iLQlsQUjNcXbywDU8jYK9kb++Y8eq7a0Sjf28/cnNqypdK6aHRD
03NrZu5OqvqenZCI3+rIgaWa87SK7C6+Qsurf2KRJUHGJGYhuvc+05T+umsd8zqPjdzAdg4cCN8Z
+FiwW9TLD75yn846ffRbpU22l+c2zRp3vdB3M2WHpj2M+jwvW8gGGJOuuFinEfMPW8awHm+e1AMZ
DNHYD4CBhuuSKcI47MdLQ6GSsHob42sIW6ZuodR+aD7bQnmM7vZU/6Tf9Em7ZE4xIVYR+0+ztou2
2T55sJgjmbEANMRp4Oxsc5z+b7elMxpmD58fVULvYW+LGgVqQhR0A/xxLcanAFzpKJx5uQHq+UcF
UbJBKvzL054+GVOQwl7D+4WW/C9oO61Q/v/YK2hRStJ2moGt64i1jn8F/JGakX4SjsBbJno3gzcO
AR4ecxD4BberaUj1vnNmJ0gDcOkQopHZAtolSRw1l22EWn+gk6FYW4TED4YT9I9EnpgSI27wcnj3
HKzNoPcHJZDVKcO0lw57w308pKlFttR/HXU1Ob3LnRXQQKzOD8bC+GBkkmwvqnU8a3j3j6w7MI2H
1uFQlVHrewnbKpLa6OPIhnslhWKTYkWEvWFfK3B4R9uSnGTjuV/AeN39iQxAuejX8VlPwHySuvNi
rDJ9OhPZkArFSzUdV8xUTqBDPIpScgD9vnS8CheYinOOVd8p28Kimh1Wb3ANqbp7eFYiz2ngnND0
oxAXkhbKu22RkcsJ29er7s6YfNlflH0NGRicYIbU3TZ31hsPwXUNJdUKIttDXV2TSE6X9VpH5pmW
ituNwvDU/7Ub/UJfj/dXrgccsTEn/v1XGtQNFHnxjynMgJ99olnLcV5Pbi4msKA3zx6PnTKwjzLC
mfZJwqF2p3RCMeX5Hv91fi0npJTTrBVoLmhLTwKEt4Cfwg4EnVgSMD9NnikjZMlc8yRw0HKPhFIV
j1R9uxIUEiFPvYeSiUjxidUzWm28z9ODU8PaJ3p7zimqTHEDqVcrL5xyJw9vjfcDZWEHjIYVtVoq
qlC3P6d1l0OGuvJD6cdph04mXPgQtbzOdm0XxU4/+PrVwwbzJZScGmOvmVzbDoxAMBOVcmbL2iSF
sfDyLU0n4lRh7XB4hUAK+ml3qboDmXXKJGAoXflFKN9MZocorQTLCeEiWlMgoUemwHAJo6TRxG+e
IMhOiHROU+LUqN+L17MrUAWFPkbjkymCQIYfwIHCvnvZRdpxjnMk+XzuwTyv6NL69bontNdaaEPg
JOid9hriAHWur5gcWJVAqejb2wCBOQiHdcCo1fozNovNjmai5gtERzcm5XQ8jVfD4DFjYq4JaomV
fPHdh/PNAoj/gV166C5YTMlu8OSbJAM2hzWIWjMzS3aC5kuhQ6ooeihk64QOkLXXTizHO7CSaJvw
ayLq92Na9bTTR/eokkeGf82vCBxAypSbRa0y6EFs6CtgreCswKQin9UWXzXu7eCJtdszcabH41ar
psCJYtsCaz7izBcnX04CXrSUQjGifDk1GrCCWf7pS+VEgNBelJqXcgKBDDcwaFJuSsz4zkyw1eI3
xUiVcBf9IDUFuGvTIeY9wXUu0TQ35ER70wkpK3vSTY1GfyIcqlMhlf2xIS+qA5hLE+o14UPbs/g2
QYipZyuwGcOmsUp6M10OaYe0qSxs4Qhg6wscuFBEAgtiDcZwt0/jH7iOhTqBltZ7e1KAczMHAC01
Vo/18arZYVog+M7LsMsNLhfb4mNwFmPAO1GscaMjU3TxKRDVItJBBPMi06s4B5oWoC7Y5uAV5Bx4
QYh+LVTjfyw4gPNZaQHzfKL4wStz/eQS/p99JF0xfP0Kdt3EXFxjpVa2vbGs9LqKEueV8Vc/ciYW
k3GcFMGeuBX1J2mIdsCjbMcbNKExs3jVWCA6MkwBT/jDtCCX0k8gJpwHtk7RVyWwwS8Zm6RCbDp/
RapoBp54vsehQIJfgFDjFJG79tzc3t7iwwS5+nR8MtaiK/CXpbKdaByH1AA7yJcwfJ5+YwnwDaRK
xs2msimh/fgTcrxSR8ooehbUDUXud6m6YdqQLYaQ2pRJ9EtVuViH3RVfU+wI57aI669Ym0ROkKQY
YH89DpKiFBYF3Xu6cjvvM9lxFvO5FiT3bHc8YIO+Jg7QeOsK6DDxtEDL40bcH/EUIuAAt8CYXCOL
p0Ig2aIcO5XTVYwZ+1ElZPSMvTOmVJGJzIIb+PXNJfzqZIy7IB5Tr7QSDEq1y2r2yIkoEzMpfde1
A9a2vq1Q7EUNhl4/5lVrk+Q/3joQMiJPBUrukgddDPSQc9aFjYWrVzPy/ZcRr9G0z519mtWfG5YT
dmmwHurL8no1dAOQSfQ8eYqI60ZATqv7JKJzEX4uvmnTWvWaQyMhrpOD3A8oCSH/UgsMhSoilI1v
Eq1gcQo5HW7K0JmFKnKsdF1JkmNiuTLFZRIWWmsPKwjAi8bulbExCQfNAx/j7OX7kw/0eho25N5y
ZdM/NQuvS4YYPEIOHD6FdhOGeNNv95jOn/HObgh7OV/JRl2bbZv9mDJr/eJ7zw+ttgA81GSSgzEV
PrWRBTZSfn2V3ReLXeJ83EZWYEjtt/QzWpik97Hk+wAi7w5ZA1ZkTE8GQV1V64jX2x4g60ZsFEK2
cY7yZkCexRcBL+tqEXhHn5KtqrObRdmWsA2NXkkTTAJ+tDxiMpvcfWTp89XVHwzCQpzJ2LEuvAGK
LusBI9SbGxxPeVSIGDZMJWttCUGXnOrWrEDUp7PZxDGR1VXXC9SarmzfchXn2zwwzGCCsvcIPejd
ToWc5qTtyNN0D+6XGYxATSukBWNf9rXM1fLbGkb7l0nauyuFThHZJ3i+UIGAkziDuxhVJZV+ryj6
k9Av1pPdA4XgCOaN2oUaK9EqMABc4cvClFJK6cfhorPa9IoqihzUFpau97zKpOabL55abHJhN15h
LuGdiT8HIuf26LE4fD1bM9QYm/ufKJFkIAO/iJuvdlhAPIRWBJG5EJWDf0j0GnEsa6ZqXqQaDICf
+neRdXt5DKaatxMGABxPwG3LmCBeKCjLnDAEi+HmNqj6tPKkhHfWqmiY/jRjvaQT2z/KQu1V/XyX
NwAIoV+9ZOsGLZ5r+XYqpSao+wsGLm4wsNaZdSmat39YhWlEaUVXJY0uX93xF3cQhKyG49RYgGCZ
z33pj9B7xLiweEVbGucU5N5l2q7cw5osBg4hdEcRmPpJSZ8sQMTlHnypzwB92DOZCyvFMmL1+Vwb
Ub/na2KxhjxXiCPRVsl2VUC58pMZS2hjGBRowYi8uClhDaRwmfJr7wNOEk+ogaA/MLSrkJp4Ckem
xcelWt7J5zfeT0nf0EUZQNsZi1l4w7u3yxOVl2ODecxWybG3XT0OKXHsPV3u8DVo1CAxzpvUUsyI
GurRw45/W8TPopIwjmZxQ/QCmm4nvvE+ycmAryqpk0hiOV/T3bzkZJXMZDeWaFgfQrnQqxEr4HX5
vVOwkYRwh+hcn4KRta+B9R7cYcuHjjsqzVMoXBlOlTuUR78vYZdmSgz7Ax6nKAMmTuLEhHdWbk8F
mD3hjGgk1mhIWal8VLDhVBJ653I/80sHEvSS7XGWGWRK+u9iv7TI0u0fC5WDEuvO2uealtDgl6N8
CiJvWcr8g+BDaJvwoNQ2malRimAXEMZA7ABO+fEqmCiuFyX1JPX27m1AqMM/jcJZLuAacs9pARaY
T+AM+8Yirm+K2JBoVx9yW2WpJ6G7elpGcHPqtAV7aeKWxiVdYandkzsrP4ll2NEcsdNM8pFQtYbD
CS+WABclP+1b/KI9tj7hzDcdvK52HfqZ3PwH9TwxG9zcTFhcN9vXzwJVIX6IWg4E0ADNqA5IGzhO
X0gBGiT7KKsn8Xy+fz5/s0wDWIDroGj3bWGpZdtjwqKOr8eNVYxu4flz4LbJp21HapHft3uhAchp
IiOnhGQCpOnRYFNbuxr6zLoA93FhniLgMtlLQvzl417dWnHkWHMEQRhQFzb2BO8bOQ5TFI+s3i6S
72LaF8dX8MNVpC/gvJp5edhWapjAVUrxoVXhlulGjJirT2dQB5Jco5GpEQS1xDRrwoEBP6hLk6M4
h6ToXf6I5hipZk5gWb2wClHpNRib7AxKS9mwcq/GtV6bvPxemUphrdLDGo+LpVd0ZjVrnDNiFgln
XL7E/xG2pWBiP6p0XZ5rUEeYe1/1LvRmUlmAn6a/PP0WWOwsPno5Yh/5VTljOlh+x3nHiWe1Qkhm
/3zc06jdZDK5wU1k3z7fDtftqFirMSQfjQKbSyT4Xkz2siOpyPyR8HKgn6eSfsO5SGTSYcPYVzEf
VQAnomPamnNo5c3ViV+QZuTT1WjOM5ZBHO/XNAxfXQ3iRzPRh+PEu4e5wV2RFdsYVZ66sedFQGEW
w3ybmQegZGYZpykQR/blw9ftyKrlG01GWG8/95ieFRF8DlF1RTA3/HHVrRAhOGWt54lYUodgTXJS
Cd0+bwTfNfP1RBC13UfdtInVFlsMV4zVWxqgHR/vn81s+gWIECJtjMngSb6ew7F4M3LSjGrftstp
aam7lKkGa0Eq1oZM54hTI1eCg9lLIOzyAPgDLc725VKGdwsS42rMhgjZL3c3rU8dg+LUTSq9Jexr
+QPkCT42rZIiRPfaztdCaTWbnYe3T8OEiiXVZD793yzeSf23tp5uDvQ7kzCQE45h3w9oFC1SGYRA
A1wH/aHWX8/faickpylBbRhcoR2Uo9u+LQrHtWyLflKBLc0FoSi1HSRJ9HJMmaZ/sXajwsWLbWkE
EHWDpA8Vj6zm3QF4xmcOleJ6n0htz/KDvdSIJ7mAiJRK/LW3nn5dua1JhYNWxd3DcouhDdjX3+By
EHMqFjZa5YwlSHFld91zBVUFWquA3Nuu0Is1lm3a4gnSU3RP1qiCdDFP0KT6FaKO78Bx6PpWEYxD
L/9ulem5yoilv8iGbAN8SPbWq3B64Qg0WbSyQVAN4HEB3GhPxERhtJC+At+eMuuefcW70F10V/f9
E5iO1S80WcyWM9du9X7gI3maaoPYXg1jUzorqCSBqmfYhL0sO3m1bQ2iYPdDeZVcKtVNitQ7Unz0
QCQuuTED1gLZkjHWMdWofE39jWayG9JePzLkcFu30Vb4rO/T7cl68tF2HTHGgAy2OdJ77O08c7+W
iduStk6dFCS2OhGNqZf5K7F+98PGR0yHGXH05rc0sAGd0cn1jEzxqJ5zP/qIQeCzmLT5gtKOYpFF
l7Hb4I/L7PEKzalEtVuNEur1v8xMdgiFqYHV0vbABa3FeiRPAFTXNJG1uSE1iFpi7nUoiYkCO62N
wQg0I+nyYCHWr5KcADS/2DBw4yfGzxkr8NCA/Urqdm/18QJJLpS4UGYv9ZkXSsaCJC9EOAWDkUQc
9oE398iQe8zdHV5f7yuEcA7hHFOE6Iby+/6RU04Iu05H487NKuzMutDTZKSAUxYJYW0ZB5KzYvjC
RHiLLgNzJMkkHLa/OAIibDZbMlACgAzgEKsS8M2gF+WZVB32SsXOxfNciz3LdTNaiSaGnN6Err/v
Iwv3UaC73TFdD9r879vtXyz0L48hEvUVZbf/xqNUN0vjxMBlK5bZMGkk4wx/LwTNezV/RwUsiTUC
e5eXtbVJ139kEMEPQ3douKhYvmL+s8uBbzz9G+wCIZN0Zj4usjWieoZ7gvZNBWHA16kGs6ZKeMh/
IJ2mzjfeLhElxMOJeawZf69ZQQJCsQiSxx47E2Ky0LQ3ZlGbvvXE6hFeCo7MQNF/X+mV7maCcE2M
16Hcs+EIUTelFwimzXBrQjh3+9XpPWa1hBkOKJy3YONF95LoA8dlvHyT+PrK11KA+dR6c19Cxh4H
yGC9Bl3YkZAV6pWfh2yrvpvaSZaMVnI117D39SMw/eTUn62R59IzNflSGpxzbxolZ6suvOjkfFGS
bSR6idITvHHZOb65O7c2f1MFArd7hkkgWI9FHjg5EYQhNLiVU72vwWE9F2vFBIkhkhmWXhMkVfID
qQu2d0udyeAhL8drMAPuVQwSzDpJU49hb6IixW5ChRmfqShANhAWD0/EFCh0XTiIoKYt8YNJMIPw
b3Gpmh/7GSr9vbeox+frDGaK6OG2OFF/N7x4pDLIcnnGp5BP5dkKzuCcjk2jJiDHLqvhS8M9Z/BZ
TeubGCwMvz+uxA7o1Lbix3VLT3zG/P/Hs9ki2flpSB2EcP4ez9e0EXIR0Jfr6RUFVms4oyL66QIZ
EDUPEq86CAlVkuvTSeeslknfDvIDpn/6qgkIANSwQdiFmaQLODa028NLpzwlyaRgemQa5CsFr8iO
fBRoDzx7OF82/2QnxaWuD0uCx8IokD0cqMJZ6Mfp/NqRHpXGabdWqBsCGHqErFNS/PPJx5JdgYvv
wGPEd1gDKbR0ior2gK0YvHfrxLjemAU0QRqEUT/RmJfhCzzo9c8+roa6eghPYTUnqbU8zog8ciCE
VDR/GQn6xYzuSUq8sHd48x3x+xVBD+yUU/ptL8wvoIBWffiz2GWw+PWTrqh1rt2V6n8Mt4TeDKB4
ZhzufEiVKUSEbbnWobY2cy/5Y7Czi1bpuGcAeATooH3APMIeMX4kInk/MQ+qzDqGR9VbsS1BN2iP
qQbbSFt2vr9tPNi7eN/rlZ88XZavQGynHtkBlOblP2ke09rhrF2ymdnR5mRYd9KjuNDLdACuTbTa
3KP0DaSftGuNrap3KfVSaNTQV2RoLkQQuc2gJMSw3v+iJCl6BzR1xlcrif/Gnk1+v9xmQDbHhmxC
w3h7Ag9CURCAGo0sZiLBBbqURWtobERK+AIsE8SF6G3R0sneojCZZtD5FWjXJDF0tYO/ca9bdKNr
SXC1U96zojRSV8caWRAxO/zXZkFJGjM9jWYVdnzzG0Gx144cV/F/Jw/78KJu2wHJpKvIcu+poJbx
cy3NTqPe5jKuhqdrf4xEhcoMdR1+QSebVriROrVtkb+xg42VIH2QfJHXdMkPcap3kElNuPEZE+sD
DdOQID4/BMCZoHYvbYoj5UmwGadjSr6nrTy8Cge7aY35oKbkj7Qd84j/SoHEjaQ+8y1JjZoApjKz
XVoR1RpJ7CTig6ezkOBxFi4WU8UYrhwwx2mWj1RFxzxLl7hZ/zRU0etSNq6aUdbkwjyqqu3qtmhT
3yZEbatgtih8oW9gDlaa8wdtmkeoIIEurkusrv6miB9MVr3qVkAju2CfjlBExjesczCsny7f68k/
qu/LTL4aLDEENOhZkIBZZCt5t68DcY3v35Cks1AruUB341tsCYQe3Gf+2U3A3FC89/nwSkmWgJ4Y
+tI5niV5yWChB61p46snh4qBYD9Ya/dhjNWYiHHwGfA4BwC68gpu/5Y+kVa11p/cYMAlSG9q6NRj
Imq+TaKqjz9cfdvM/CUGlISQROart1ozsaiNk7YBYRw0NMvuzGiFGRf0uggnGShh2qVs7AKuFHok
JiGrFMci4UeThRLecoIg56tJXvouSzrEIWFh1FedVgn4lamxAjF5TYEWvAAbmpkFlk4OEr2r//R0
Lcq5N76g6+DslJoV4oveD7fiTlU5RjwkF/EPvtDT16ElqQ0VyZ8r1PGQOFD+YeGXEYX4NHj8aGm+
qzOR/tlBUuqC7U9hWYtJF7XtlwPP/GuKtIropFi5zvh1f7OfAZlaeYtf1pGySEVslc9n7moXODH6
NVClgTP4uTlBd8wxZxyibFhK7bcPQSiBrGd8xr3x0JSu0UeIa/fpEPBpxkL7n4eKNBmcm8uo2yQc
ZULAkUS2aCiuNzMXAl0+GB7FomMx11gUCF2rmYick8LxkHnfaBplAzG/23og0Aai/iK46rhbPZuO
HPr3MSKRVVFAXcVr7yKdXflAeXsBZbsLopazFTyjThFiP6vlzguzvaOwjXrqcNgq4X0ZK28VGmFt
M0J1LrPWWMQIsFfI8FGrhrk4czSRB5bKk1Nth1UeesrT6oHvFUjTr++zhSc8sE/5iKRcildMBiHb
PFb+MzYhsB0dGeGUJ7LxX8VasjHw3dClLlEwGBO/WxUf2Vwi2+eYxl1H/xyWw/QWBbLr+kfVXnU9
sJwQVq/CDST0fqfo7XEDsqMOs1EMkjT6fO1Lp2CjlvaxH1uo5zErdWXTD41gIiWinu9F48f+6ZXZ
xLledR5ajdp2ae+DwIBSXSnWN93Du5oRJwOWuMl2nU1WpDb7ZZIRD9VwTe9qi9xk5b0d93PIJGVY
LQuO1Ah3/DXivuhZ9IkexIcEe8eoSwfgECLAUXW1E20t06qqhMfHCoo/rG0PxycYENf9sC7aiS55
nbelqK25H41ZFeCF4OR8QodOUeUwtfynu1D7DFaSSgT8FwKhnGLDeUjdN/G9f2ZkKxSpfLUVrghm
BgNFHKesyvvUldPfph4uijELoxqCafn3julxK8LRyVIR4Vm5lVj4FOIvf/KoFrbgVQoBEo+rN2hE
YfBm8eVry3TnPgbfs1A2KthKBFTy/clEzdmrH/JufO2DepYBtceSoammxpUNDaeuN371z/DWs++X
c00H+hDYpeaVjitden+jagB9+cVbMwqOFh+E/HO9UNHfHKD00R9kq0t6NZtcTlkwLVaKzWKsVh2l
my7TBf64RL9kBY44E1yf76tOSDfhFVCAd3DS/FZVJj0WOp+pxz5/fJtSSLFI2AtspP0iTjzrwdcU
VxYJtDhxZgflLZKvfPFoispznPKObi5MMrDMAU8hFI9Xo7uQ6rkrCyP4Jy6GQ226bzPFfC+uUKeT
Fw1mvI0YDYyb1Fr4dwCqeTkrlGFqjejE7gvURoLfwDUQPuaLKiRGG7oHHPU7DvDGObKbNfDLkQP4
i462J3oA7x3R3/Fp7oGExgGFZatmUq5E9XlVYx6CCQCPnJovEiHlvmbPTtRn1xJ3QTbpu/+Q3vP/
bwzqQPHrsr9Tj6sjl+CzpmGjQdTXWQPCyuM8RS5TmNeSqo9f1Q9gIDY3M3CyQAu2dE0ayanWvmSy
FxeymrQYit1kuI8wkCFiZlh8rtoh8AcwRDFtPiWnuk06fjOptnHrRvu7G3Bf8l+Idmyi+k1x9Dpc
+iQEHvQ1qkdM6HI8Gw2DhmcPmRokFkqPZiTomGlvJitYUxZvly5RbAI8liD/d4jl6D+D3qTec7wX
pbcSvJJBZPJYH8yC0ud7KML9okc2zKKkOcDbaksv3qYV40kUlvApxXFrvraJFVL9qj0eWAAN+P1Y
5J01ee2DYEi4XQIFa4IPEMJZLgV12KP8QmMokBewr9BtWUSAm34Wsga2jpArWumXpIjv//oEtlv1
9rYq1RGvVFNWFH7jU0KIQUPKLRERPq/X+gyzmwQJDRL2jTle9gfWorrTPuDVdMNtRafMgusxhCPd
pFZy+1CfZp+YqMJ1Z+LdNHfCiyzr36uZy8/3GQbpwTJ08xtKWSmCRLJBxFIllCfu4dxBje6GLbrM
xZ8+uD53zW6iN6fq7Rw5JZTKWfsbyODNAdhZAr1H9nY2RIC1Ob1URnFnACtMWptOye7msYs4RIYF
gb7brkptY0ethYQe53+3Ibi+Bi5dD+B/5h3y3eJ6r9ExaW8fVnPT/DJQIxtMh7riGG0tl81vOzki
0J3NdnH3mZxH8fq5N5jmBWq5uPcCsn979llrNA/uEy7U8N6ydoQZJJ4WaB96viYoSKbkb4Gt6YQG
q6KYSjHJE3RLHf17ZjQHl42IUjgXgZIA6yfIqI2SBIn2+xAlmI3OIfqrkCHdhYG2pGqezwtsVwc3
+0FK2nco+HbPLC7KNQlzqG3d8kXFkFfly/jM8NDhD3JDWasKFE4XOvN/fK4mjY+b8lzY9AClpYIp
htStzC+fHkUemNMbhuMUNbn/GjFctTMhp+j37C8qZV5B0JE3TdtfAe2/hE2YXZ2aIAVT5DSqyKgT
dtUOBg0srhEnqEUKMp7qSnx/AraOmb9uIrY52baNYVSLOH5O44s7u/j9g729jpP5f44y1i8MCZNl
8hp7YB68rxIk3sdJOu7Nic4zUMmW6N9ugqEKXomhCht6KBqT694+hjJptk7IjRd0BffnRwf44JcO
bymmSVFbm0M8UmAJCcgKHRZsnBzVmtShUJYEls5xNy6fR0efohIOsQ7X2Jr4UpD1V8HxNOxlwvkA
/T9Oejfmujd3MbjH0tS2yeingF7CSDFiiGtWPNGShL5aBC/iEsHnKxSgh3W0FW/TdzKBk7HVWSvp
sQVZ/iCbMrVue5bgrybWTJT+dwoBPCqVM156Uca6uDZuPcohsoPpXCdj6HSeA0Bq2cReC3aJiSM6
ljv2RIwlIE4X4iFPBNiSe8abKUFU4VIIMgQtGVBY1+zgl9EC8rY8anhR8dnK+FqfSMNlBghOLTnt
QarmHHKw5AD46cOrtWob9xrpfHpWEHEA0uF4TPTrMLBwiYypHPfJ2GuM0Wi44a+F5MbWb6e7dq2M
q7fUpZaLSaQTEEtG4r1lCjn5QLRLoj+aZn+FQiGsgVr+nOgan2mDHB2zKqkNsTymVG9arT2wLPc9
XKNXAWqSX7YRev08Fj/i4Q6hbP5DO2ltuiIKbzuGmgVjRHp3N9SWjYtV3PRf/1ezrYseLznwnNRI
906tg+jW8b0SyRNMcXBP0aKAyw5u4sLNHcf+VuHO9UiBncKZ8aO9VBXRQC+uz3YEVAGk0VTLbLKe
zj2Z0O/otn/w6MWgWRQ8UjC02FImCJkmYoTSPKpn1qGnHY13FPpxr9bckknZLNCn6Qn7G5Ei1/35
oQspCbKJNorbZo8LzQVPKcoWokru+ZPlqljRgTddxeElKdfCJxFGLiTzHp0WhNSAXrY4T4Jxu4Qx
PVYKXW9HVP/JLIj867O+r9L3H9ZFi8O2VMKJ4KR47itvpYyqRDj2cRSHeihq21wP/t3UhtL/kLzM
PtIpmZhSgektvPxI/wyj3cEn9Ih+YAo3Nll/e+KVu3L3L/ANvD29QbWn80ZKdL9QHouDnf2AX3JU
mKAMbmkhzKVabGd6ldeCVaGKGVkAsCTECrf0SYXQD+1AbpdaJW+3p2Fz6R4a/XBoJwuOi3ZQkXts
jklFV9RptL0PNNWrkcum/n5Gi5KujdbZb3RUs+Inb+MyivBPkXW6z3RZ+5rTHPwqDSl7Ejj2gV7H
NU9sJ6Hlr6BO3aMZaN2RzC2RVPRZfLdXM/60UxJBrTnNJicS/JHJYtTOC4X1iHrSn6QUSLV8Jjw6
oipwphc4K6uLo4cpRTgWtzmr+Xw5yD1QouEFQEAzntwisB1wQjmLMaQiDPCZajAjrPoEaizMHjDJ
XP2Gm38jqNKc9wyXVcS+wI/7osed0oLA6+l3Ke+UZSOTiYITcNPBvHDAKSNA6iViXa2QgGtMdBor
3D7FY2RwrCvo2FMg2pq0XMmUyjR8gDWPW9hP8NeezTf8VrfntqTJufLbTM88lGuL1a6lWnBp7qOF
RJwKf77q3dORTAHfjP/4tfb49LXMTOUk4nbDJ/tp7FeBvfPo219fTcNN4Uv9GUrufp1S5wMRJrxJ
H9iNLEn2NgdftUBC2cx75TDydKrAR4dnQ9orJ5CwqAzjUkdwxiNsVIf2QUBjQDhQlTlx8H6tu3la
FiQWjqWuQY/GwOihBPaCaa2XoNA2sd5ATHNR1CWjM6Osb2PBKQdEvmrfLwIB5E9lWaQWe04NMGEZ
uSY0yR4UReS+0LTvTlLXQ0OVxV4XWEjMdvR41j4LbeD6zj2FptFl+RQ0arrlykCnUcayvjcF2iJO
dKopgkl5YzzJotvplwonuBukkB2jvpar4VJzS/TZJo+Z5klZXSJXEpSCmzhw2Couatazo3PRQsWH
c8MpQIi/mylejuFU5BNni3T76Eta4Oiix5Ocr5pgrFUp2mVhP3IUpWyxhzLaTnldxf7MrQVcSnID
AIO5wk4wA8esqN0CFnw+yShIr9t/1NdYdLf7WbCeggR+kgmeSJm8vR5wvAqwe579+/lxhQTCuQNh
Tu2wogRVSFHzHLw2VpB7S3s1A4lXTrjcOq406HbpGxzusdcddZdp3TA0CJ+t3RkTNSFx1kE4Td4P
Nl/uqbrj66Uz4F/GMLQ/FxgwTfWXSiMqzf7o4HVHbY2jmXoqw2QwuLzgA8ACYcb1hsPY4029Ivtl
IzTRbmn2CKVaPkTZpIWxre0zLXVPGONO/7/8B9PZr5Ry/U4imglqAehOIjlAy2ayCIs42mOhzPKF
2h4m8UOOfYOQ3JssqDxjJmnzPr6kRb2+EoZh+MjAKbOhJuaBTWP9M3r3pexHGRejnpvN4VVMYVpQ
69YheIymdafyt2W9K1EgpRTUZR1H+t10v4egqRnGGpfSWomRd8orJmqs2jSVIzi5joiGRicvQeuH
vQddKOQDVYyGqa9WR0qQmQ/fv7kgvcXfOZznBfOJuNJ2XGME/6jO43qR/D5bs/B2CrPoWtGnPmGc
Xl5KF55G96a11W4yH5l3eykWHTP2wj3cBCJUZARQvspdN9pDs3fc6yCBcXY+uPd7cPkpvBqrhNwE
2Dg0kvVceCww8MSG3xwRHMnPEA7uNy+Md1NQaCQy3LzozJ20gQyoCqwgZN3ikLvCGs4KGG8F5u4U
ptjRg2Nyt/6sz6H3cpt8atNP7TzRhu48OqsVQxDuEoPP1QbfGZbHMH2/PdMueAT3fsJNjWuguKsH
JrHSeXsf8ozmVw2K3rOojN70vCn2YjHS4Wh95OYZrGtsRKq2GmRV3zd+TRNGauoz0rgkNDJ773y+
R8LWLsX74iijSNxH8Kh3NgZAnrNACaPDAAZ+IWsRyoJZ9r1hyzsbCK0eLGHrHCbHcxE5BveNtWcW
7qUswJfyeCCwzETDiUmG/Qb45ePj88bf/mw5+9jTSIiNUozgGAHBe0Fz9NY7UcM+lTQcuo6y2fTj
m66yPhNPAebHP3JERNyrJUX/rh1M4smRPIf+WrPgdKq1rwKlOAFXgvkwNju9moVv6oyHcHoe8LcP
97UPtudx0xp6I1CL0nHy953p9NDOT7Kq/SPG8I8V2mVLWBIDE2wzb/K4476faGEVQtlZzpi6bKkz
s/tJOhfaxhXt86gEUWFLgE8h8I/SXwUqkxB9QXLM5siIvgv70ikGb/Z0AJA03zUXm71ves4NyLqz
WmdrQU4TgfeV4LZdF0lETgE7b7qTdmNUqiDKdacRdA2X2sQjG+u/IbOqjJWFgt37lxPJfTL92RBU
Ofc1gkJs6c8vj1Up8MpGoEL/wlYJAB9+ESMe13nh+w5TOlXidGr78AAYEikpGkiRZvIAHU82+e63
CORw0glJRAxmYj7M4rc3ZdYi+vOBDb73BKulYBAqy9RXgEOfUplAYyZE893x3paLmBhZDiQmfEsd
ny4tvSHvQIrdvoczNjRmk/3SrANMobsObpXcNtDHhQTg5h1WpbXGHHz4scqIfOn9x/iYvQoML2sl
3a7QBgCc76aeqRuKGVatEnn9gI4DtNPXtE84RLmhLffhsUyITRE1+9k+kHIGaMeBuZQx3eJ3QnaQ
c7Vb4oIV3W1iChO2G1Gypycsp/rkdZeCjZnMRuytn6NK9lbUtr2f1mfmhg0xQ48EWckrFdeLmVz5
CZqBJ+pGCiGM5ecFgVAVco1vMTMBLJ0NK44MA1OOjQGgxXJkitMAeBQUcvgyDvNOGFXl3XgVpvrH
GJt0PQFQxUsofJDePH8oNTajHw1/dNdGkBQmnZe75g/EpPCm4b3HYKTjXlVk8D4A2r/mVIw01s0r
Eh3LXlp4MNnXGKw/3tajEv6r+ms5wufk7T80jy7kN7HvdBMkXtiJ81JZ7rVfSvusmgs8W8t+ue43
KGiD1NnLdBbtR0vOsmPeHs3jPEb0m1+Lyre6mM67Dkt02c/ilQNGse6h9IrhG86AOGs4VfvD0T01
+OpCc6pHwYKud2EXHIWkVp/bwWk1ANApS4yIimSn1C5HZhTUkIL77l9aYsx6ZiopsWnDNSnlvfkL
30vRSJW+LOPF++i3tpl9shjWFf4MY1GEmxQI6haPQaKLgeC61kNNdVCWDzcMCbXUSSEey/jW3ujq
C7PGgMyTJAgRye71Ys1WGxypvMNFEaPO4hBJlbQ8NrMyjuhtOwoVVoN4gO/eNSP3VIidRqDt4rVV
DGuyj3m3Z+DuvutkXw9nQrZwB/9xuaccr2U64NYScFu/NeAIF0JnF7AnSQljWc0edwZSXxg849sQ
WXverlgyvvoFLQC6Lijva8cC31tRul2AeroGINvd+lyVUeKsfduH7kt3+nz8buFaet7p8pcbFqOt
kkXkln0SbXsMcwGpuy8oTqoFkRrLWXeyDGjBdQAW0UFyGrEDEXR3v7jzKGV7g0vg1z/CwKXWrQPn
hAFniuS11u5OdNGsVCjEt1KGCDzojWOALM+mRJ72rTG5+DQeFPqx+Qn1Zs4wpYiE8xe1ZWBtPgq7
pt723sj7hViThj5RBvnTOgnhxB5vPAcuTuqthT68PizGe6NL0uA22qTIGqkSXCTcocUWGJKHOcrS
WzOnoMyLpwpLhRt+64bEG8j7gDJSYHHFhZ0UYfYR5JGjDdo/y4WafWxxMzDVhoJ7qaSPAzcn789y
R/gyQQ6+BPcIeswUvvGfMjsZ3oIRpNbD+BOIao/OC11xmXWUxsDVMI0EeKcp7YWC9YZ7v1tH6O2l
O87rI6oVLu+M+Di0gmEGKKrNGvxJOlU5b95BgcgikT/t2TtT/S24FAl/2lT5m3GsrNkwTWO4+fO3
D+pz3bNhF/eXRTp7vg+25DY8+E9RYJo96qODpecPjNGkk9ToHZ2UzxZedf4LPT+1cboyIyJ47v35
7Ur4mw87r5/bDQ/EH77P8kluBmb4jz1qTWMYxoyodlzzFNzBEEhytsP1AMEWyiWYTuWQ24/AOHr+
JzV7WivpMZM/GFL3/s2QnGHIF7xj6Vw6uHP1sYqBR0y7cxQoxWjsVUsRe5VIICYK4cmCs4Ptmriv
ZDAflluaVe5PT0NxlYdXCEBgpLj7++DqGZPrcGwQfqEVd8YcH2juLZJhY5T3JPfLFsr8V0TkG+t3
ZlR9QVV4hsF0ljet7n/ueoStPjIoanQJMPs6oKvFB6oS+zVKSHZPEsd8M9uzvIdKOWTW611T9BxT
c+ykC4ZOXaJTFzdL5IuWFNOAc6J03vtTOgNQX3pm0LY1hW6GpmC2qPWN11+imOPzOmeXl6n/v92A
QJMH/jxkeiCbYsFFKhibnNVjkEY9y+rbMvOaIM8VoSTXfKOHmE6W2JGDG/osR1dTJSs2xn7V2TGs
Ico1bwG4V0cehztWTCM+tpcKSswnbJdXuNqaCS/Wl2kMTjw8lKIR9lBjGKzRAXzOOmmcZnKWhyf8
vUeh1yovGz4jnJfdmnKU0LjmdMBjbma6pk+JHr0ie92LNogrIPgLl0iFZIudH77RvI68y4QuFZhz
bMQBCqfW9PppGFI2Fv/52p4nr3nWpKZY8CmqWXo+1lFJNUL1Hrv+sXg9scsKTk+H2/KbQG/qeyQo
lko7wABqK26q5uiEsp9JAcTb3SlEkw/cqN3sUV83822t/nv/ELmmq9CqvIp1hrPQINlqsf0hSdgu
zXSLQWMbUe7z6tJJmi1RC/K4U2eH/95pIbUhsDwoGNhxikhE29eg2qpV2nS46XVo9l7Fs7VZ6zYF
BDAuwYiYnspax09L6Xn7WUOH4EOOMHXWpM8jXx+jEzHCGCj/8cO+x8Zbpn1fRxeam44PFA4Lcttn
ZamDdH6O01dGMJZfuel5uAV7HY56o2ef9pMzIVv/ZwbC/RKOxbfMa/JBxhiIi5YRu6II2zMwG9hP
ETXi1zMK4PRG2xeX6UVRcvYJC9gVeOFgNf5RHJ5FR70DOu7NpLb4/HaVy/bVgqygkQBIqdH1zshh
C7HpEkSHvpboxb8XJdtR6Y5tQI9u24zDQ81simdBwbZyhR2+/mTZRxVyScXdYU42I+Y2nOAI8KIC
pO8rWIwneGKUdycza/KUSh7uul4xvRRsi3qMgR10VlA1ZWICVNePOTN6cDOIVMJsxy3R2B5BiHhU
slmgxS3MbwdVq1pYmL1LWbrisw4OvO82q6gW09DaxqwQ4kR0F7ntxv9+GYtO4VaMCJayYC+723im
E4KEM9b6uuHLvLtNr6lsnhFZnodYc4H2OwxEowYkC5I/WrJARnxQYJiMMboo1JvywIw0/Gq87TGO
hwG7/MBpNeR4bSyvA0Ogy5wb+p5bPaoDKXBvhRMqwEnZRJCgj5LNMd6hBPkjkh+AgenOHsUM1/sj
NsavKE8Pd9tNAw/3/n1DK1+VqDwT6esDmmxkTO+fSwUoAmxy0QCnAZ03lKXkBfxLvCaIQvRk8Hh8
axwSnQBBJh7JumlFp+RgZOcj8oGUSufvkvj0wDBhtmXRocSaLiSJTVqcOKtmTK/x7fCXCcg8FkOn
y0CL//JECzm13ZUGXqJt31xzG6xiwm+3jwQX1IQXe3j7bkFvFGj6KPaBzNcnLC57bI+01CDqEBvo
PTFpIVceN1C0U3BO1YE7PAibKL/peALCoHQIGNS4blo33lim8tyZfY7MNQtsMg8cdgTrWni6tMEQ
sR+qW2FK253xBfcdg9kBTj4nLnPtqH3y6CFRGvzITI+GG32H6YRZPHQtfsH7y5d0GWfRpYAL25zD
fymC2usDT90j8Puvn1CNn5dhnQ8NYQT+qrYobycEjkKZI+5LUtT/MgNgyfOdwl/Q0VlK3X0aveQf
a2BiY5pBK4E2BlKNu/eKxmynS4sIfDcduVoooxjtcM1MV6dmhUejvPPl4h06zfy/m2vMUy1JGh3S
7Wl33T5XwLpRxewlfAqE0bzcesmHQlnPP34G8m2Dt1nYj8GeP5YyXUrq7xEpcoAryvVXGkHu4i2W
b7f3O+Go/g7zGlUBeEg8Ncd++NQWhIy6eikSV/Akelv5IkQJxpRnPph7kbemPQRqd3mSW/KgQi2s
rGtOSUfyttsGHkVkJichDxOXMAw1GNNkJwG9Mzr5CohIrz98cD4FkNWQenCn3vR5pwiu8sdpccw6
OKmlSS5ka7lTl6Th53q8sybwBXRb0T6dleiCVIYp5vtC4LZxal0gfBT1mBUFbsR1Vkf5WBU64wRp
geSXdgiAgTRoYx18qwG5WMt6lk54FtqxhR8HBbfUolZ6tHXri5OCbxILJ0X6ngYdtoHinAiH7m+9
Ku0m4Y5B7Mwog/xFNzkFjEKMmCAQd23MJyQi6YCih/gDTVarIRBXvX+ct8xEMq90u5LQTsxCGEUp
Euu6zoT2xO9CDu2iEPgdQO0evVxBpKkMvpvhc5DxV4VA1r2ESjRfK1mjoVidqqwhPScJgSi6UVCn
8OfBvVMj0MDcErMlmcRdLZhfruI4LcU/M2bajNJz6d1elm02O4SONOdG+fYucgg9+0reYvXwgBIa
1mqLbTMzGQx9ORckcgmBfwNauTW/AKNxwa0CBOD6C/qlIJNL/gxn+lIDI4S5VaQox9ni/a2akAO0
IkE8up3GtQLvzq8KMRmWEN90RApECB2EzjrxFrkc2rMP/h2z/LqpdbOg5UsulY7VUYAOD8NmEZG5
eiuKwXdfz+Eqc94AwJ9lb8rNDi/MtCZ7qM8+g+Za+amcTquHwCINxUFj22j7C0OWLGUQObd9C6iT
9d9brl69gul4iM/HiIrLntdfmqYhBR52VkjQTjQEnTzS3qOiPJkLG1WC6F0Qpec5vu4alXywieEo
66ddgbIvgZzFLaSK3DWR5QFz3fOXBwsv7kCgUuko8hEmhBmS3yX7uWq8KjoWhBHfkLItIBOJr5Nc
SVcIIq4oCvxm2Kp241LX6KGIeFA5v1PLx4f2RzepC3YmmKi0dpVKlWuN6rH8D3pqsTO5o95MRu2h
4MzMbVCJJsk8bawDQaDeZjHK9jNrlPA6Zz5XEMVcXERvDLFzxjIGUBVtZgKbxK4oYZJo6hyp6Isy
Wdg4oE/7oftXTh3D1K064How50tlpv6x0k4p5G4T7cVzoBvQ5uCwSfUi/OTKEwldd4kv+L1I/JCv
cKl6dAHkEttCzMLr4U3IMOCMzZO+YspATLRpo9/bCVKBTls/ZedwVYUQsXWyhZFwkyLJdKs/5Iv3
R0c3PSqnagHWKsQQX34tGIB2qENKxAr/Sr8i+TMNTd83Mgz/iULzsn62ogZIiWpmVmAg9sWeCMZP
2CsiRwlja9eIlowAAL5mltjvBnqxa/q0l/u3atVSTQyEIuZ5MO/QqI/dm5YFNijrJh7wsUJwuPYu
zOUgw/quqS0/u8kbU7sebNoXk+YkgSYzgOTcpAn0In5xVRnltC3Lt+l0jAkyvbiIMlhwmD4lrnx3
vst8R2788pfQ0tJ9t7RVnxECm4nk7nqAokwjexO0M2t+qBYLdsDudgmfdKJngBPXx7heiVRCQxeU
RtIanhjDbiopT+mKdcielEwvVs0l3TIk10u8xeCHOqxXiZteivSWjTh0gPXuU8YuSweQ+zqXu9Fa
6dFDywdyi4HTx7D9XKOiHOwVaJFgISotNCUoWc4dwWyacbPKbuOrLkLyWZsmGfqhI5OFg8v85HEx
DDUphBo1C7ZsCZmxYggb7RZHDt4Cd+yAACya6p4LwrgyZ+HEGGYj42zmmtrDJVb4TIMkF3h94o1l
aNf3RBn4KHRhwnTq3eltU7AsvMKWvnC6iUizHdckM2ij+8mfcMAOUaEn6ygRhq4Hc44o9a8uCFel
QeqTjUo9T9xp+tHs9na9fPVe+le4+0UbrYScvZLezENVfLqGeEIxbWpSsocazUuxbyp/FBuLpbC3
cv4ZiYOiLqRZ+3lbE1YQVp5Lz90kWOVklXIPfrT8wYwynyE8E4vdqEyGZKnkCuvRtLTy87t96vlI
aUzXkxQdoAO2owOMrL/CnjtvOYp+EQVno7DCjeeTdwSa5buJM6gxWcahDDkrPidkzumqX7cks6K4
FDV1lQXGJ603xPjC5bJeoDpA1PYtwrh4GsSIJ/lT+NoMSaN7b8HR4iQSQ8Lr552awhH12JOCmiyl
9IaKHKDuuZgiIbExmG1fo0y+QQe0jDPrPrlui77cCBvlPKTU7AWaotDcttdxCzG+yx+QOe15u8SD
Xu/6rakAfboN3kp5dE0qhrSZhA0pUV74oVv3RZUniV/TbVFdca/SMVy/cDy86mH+sYlVt/P3ZUj3
zg5Z+XTR5uesXYhntBDsXD1d2jMqsyckJJtEAgzeuacfbctQh18PHItSYPKYRLeXoAuYvi3/DDWs
qSYK7ynoW3AJ0TwdNdLZcVRN/C4nvcSqnfZODsmd8qkJx0+r6Jn6QHP6K+UpxPl92Tn44BVXNG/y
KUtB6KXr59VnBBMksifCLlpHxHiDky9xDKXRmyCStI6uk9+7nBTx9TUH2tg2U53L0pHJB7xmxt3c
RlBtmwDsCTguBQ0FJdoVgAsuTcf9L1K/9PES9pejRHzZWyGZ71nOFiHdYh8lpHvJIxwfjhXScqxJ
F8ZDhC+tkjtcxY16r2XxWill3H/ybbaEn/05xkgm6eRWWcUm2IDHPJDKhpDC8ypBX2fSaLda5jBY
lcZBWSzNXms8EBIPb9x+auUzDWE80yKx/wxg4GSm1NAaOE3O3hCCfGCXTIgP6xDB9gnopXKCv/Zl
aqoio7h+44KM43yq6+s72usrHn6L5sySqOK+9GzWITtBUycAB04QobjmfxeKdmGQeJMQWR9OwxQ5
QBcTMM+3WeRDkEW5Y5C5GRFZ/ohJONvp5vnacscmAHO1DKHvaqT9o4x3zc4tz6x5Z1nTWhjJPyTL
Igsl7OAdHOS4WJAKQwiUNQxNoxZ8R/EdzzR7PK0fv1zFqpRPV9pyIBhcwDLCT0jJ9sEaXnbJqN+4
6cgo4Jw9PMovV+j43omO5LGl1gJfw9jlCi3vkh00hskT3DOZ/jn2ZBjwjaO/DoVykqEZDXeVFtSl
cLpjdHs1bMb+3OFrvu/XUK+UqMEQ5Ywej6pgBdFZFouM+GhTBEgnikMt2Xlkmwanegcu08ugg1St
CNThc7PqP9dv2g1ChnZGJo24rmAmoMbgE5XX1iwNqWtgz19Ja8qlX1ZVAQCsW/CTmbOi2jlEBxPP
mDs/DVfhBkfErrzNct1QomHNUrIggXchYCtyMWcKUgqKET7u2qOuv1Xw4yZIkuAcMhrNh3F7SHHY
3j+4p/n7oezN+BJOzagWxyuu2PPMkQFKjO2fPqFZdFPwvfc1Mv0OyxDP2uClkNMxiXsDwoccUHmd
uqpOtixnec5c6gJAbyjfYTljuyNmPbWDHJaGmdj8AjofwPb60LaWymaFvcsRmVDExdeRYdhwX/H8
VMD3wAa4lCElu+V5r4lAsjaLJCh41ysDVoB0xt8sfk1EhFMj2r5NzS2G/YOdXoNQwLyrkUlh7cde
8zSOHbDoMxLmAi+BTz81UH+jHTohswmZ/Rpi599AlvCJdiN6ucab/avIimxNbfTYGfIXslsS6Vv3
J3vsGHYGDFalMd8tdwH7GnLQR03AVJH4NP9QdRsvEKgZEx9oKcMxRN2c0ohMzWDboY1DL6XbGSW3
VVSD/LFeK7ozKoGcDIUL9Pf6nPLu8VEu3/16kNrHoPBpJdK9gpI+7D85GMUtCW/uhaYcf9xmWoB3
vUkKDYRg3N/K0fIuvPKtfykfLD/CN61GqsZTcCqe1ElygMd7C2BNjnH7RO3ntd1VsT88dzLIljBN
E1xdX4N7YtXDuxmliLsQII3efe1he8S+y50qXt3ntHyQjnUwdtHNsr/UZsYh7eduOpkYNGBcbvVk
plnRutm3ZD4AEm2VtJq/BmIDoNC7G7vVfkhArGzHpBuPy4cdA8ZVZCt2E/YPBjsPyZsRB4R+NWy/
IWhY1W1UPBUFCi9bjwNMr5PLQjfVSFCeOOiFhbWw8dwofqbDT0KjFf4drNB4saNKGFo+V0B0yyRG
rHZGL8JbLIBx6SBaOyw+95Uo/HPkPztoroJxE3fi6SyvD4z09K2wILxYJuE8JX/VrFjPcBPDi07V
ttH53aalM7FnSLmma6ARGh+7XTAbInaCgyiBOewB4fbLyOEQmPmUDkS6uKSDfg2fRgk6jMDQ+LtI
Rbgbo3QtLuJSxKoTqSeC8/74IXdyHayRujzc5x3Fa4NVj9xX5rqCZbcOBD//nxAsFrUZGgnN/hgU
d1TF+VpCDEj+X7WQPHjVtKzxB1LU64hGhgPtxhFTZHLbB5q+WyYDhVtrgClJdsipWi4HQJM/e/4n
uDi/S55tyKV7qYnkN3fna8GeAfilkNPoQ60yBXnozUHILFOflCla447Qxn5f2uXNstPpZ+NayqSK
kUUgP9bE7y1xrM1Y4IGt4aVBSlrgncHqW/BsV5OELuN/4e7QYjFVa5VsUJJQu7ezXeENgziTd/Ye
93zbsxc05XgA6bmaFclQ1cpMUuAeAuzgmxSWhEb9b40KEBfutpHKfqcoFJhCtaqjlZUBB/8SAiKZ
nTW5/BPSGWWmtKY4lZ/z25e6AQhRDALb4norA5XXd3oAU8zg/kRc/Clrb8ypBpDdNN9p29cxjADN
e54hiCf6mM5FX34uUDhCLhFKem6bLB1qolAKfSHhiBk47aCPlLOjjIfe2sUdBkbBLGLmCY/V3qQX
RvGNe53/NSxE2fJ9f4C5lzYaCkdBFXOeLmUJLF77qY6y72VV61NxZk5UAC2/R0n84lwmQix8P00U
vf2zMfJStgAcmoyBCOV0OpRd0IuXubQp+qxjYi1cGESW39p5C+58wGHM02DuTKJrBmVaFGAcGS47
iwpkbdupWe95W6LbGtBIjOVqhMQvxj3OtErG/FP3Dm7e+9rpV+e2mrBXE1U4VIPFqOIq4j92UZNE
QcqI/2YtwN/xYLFGFfu0vuLY7nQgtoCdzyZEHs4l2TRIxKLMQJcGNSEIeCEV94W2g6OAVdSU+dF5
jbTldIn0Iv6qHQmG437dwiNUGmNRepQ2ockZHfh8liOiuq39+oo6kc15YTlh36DRQBFETREgLA49
uzi4HofMJ3Ii/09KWa8whnVGmUfC3xYt/Q88jeNcgrKvVpkQH8v1CszljAiyIqo7NlFu2G0JPyTa
6RyxTVYKbiuPboDRoztXn+L2sClizhH17cpPFO0WMz0TfOeYIFZLlur2ZiPJfnq921ne6yqAFrnI
yTqGqn6GyugMQvdeBZapbdepe69pEhXuEHHkU9lpIJX01XKf3AmU8VIUiyavaJdw7Vwm4ayBNHwB
ImIoeh6pakFR+pZ21EQJmT919WY8E/qwYZrITTzfkTn1srp98zOyLp/304RccAXElpdy9/rYez7+
K39ztFF59zVCMe6MTxi9967wfEK6BXxMqzmWR9lklzNV2wNa1j1dbDPg4jAbAju2bfSjx/iQwYUY
WU/1TceGqS5t4rVh33M3mBAIAjjHcZE67mvK6vr1dpB/p2mH/DrQq7a/0aifyxm0k6Q7EfudmMlM
jTsw80w2X+Y2QRLphAcfEZ4wS7259gziSQLwTEGC/VDm5bZ/yL+qnpwulHJgNBO5eO9PofCt/G81
QNSc193IOZ1XSctZpNg2bRzhy/eQsqm0x+2lfEWao1C4c2dnbpQpBomc1PbbOOiCVxqToGnOi+P8
VH/L380imNbY4wcLmIfNq4FiZNXvYADmrXqHQtD4FYXYVFVjGc/8gOkc5j9hd0379AX5kPImrXjB
sQkhQpLVNeqiSZHHfyT16t5CyJm/0nDVHPSCcQLiJHue4CZ7GttCyuxP51ez1/XTB25Mg+fW/EM5
kPaIUnCPxBBZK+tkG7f07BKa7Wv8s8HoGg2Tb5hE6QBzAbtqV5SXREoLYAhsyoQGEJZY9JdV2t0a
G18XgHXSWq4YMUZffJuEJgnB7WBa809NGzWBX6cm8iwKlr9tuD5Vrepk8w01KgX0tZ5n4DE7TDFN
nHzCUmLk9V5bm9PeYtpF8jjAECE/bjFayxIliDJ1r1Mpc39sd49UtNs0qkD2ME0UgGrBNXeo+l0p
PUnjYmpxGaN7LoCe9xV6LSsOY1TvPNB/pKcgYrpE2moYY6xzhy2dsC90xTVM/sD7s1ppZS3gPyVW
wxTgib/KK1b7Oi5InHGuhwHi61X3NLosdDLfqx+J1+GADzh3QgS42KbVVOnS5AwvOHmdlKst6y/c
rE+b88c/7RxL50/k7pIAWZyi8XumeZ89dFdT6xazenQu6ZHEdkOLsWytTxvFnMJid7ULnKpr6x5Z
gchtYWAshM2QUudtnqH+GuXEOuU1788AWBZXKRnqlcHdX6jME8nfbHVx0zA0h9jJQwFHnxprJ8kf
3cZTacKyiE9Xsj1DymQDALrdf7LoFeMvCl++5+2dU6D383P0L33VgbGpGbzrVy5obifPgn+glhF/
PnMo97PLZYgOF5u6/lcWhBTVWSsJ7rY4ESh2eAvBO4z6xa/W+ck8+jmmLuYIh08UltjMT56TxMwy
Yjc5cOpVkPRFP5YzhmCmhTQUxrfoCVTIoyHDZCOYwb2sPuNC88EolqIlVbIb7Itkr7gk6CM6QVL6
vMmtraiD0ovK1vWCPaNW0dcaMta4wB5B9ZKCL+MEYr+I1scUMpL6+9jm8Gsee0zhw3jQGj4UvUL1
QyzO7zAK5sMTVu8E91QaYFZJIrBIJZxansTVadIObEaj3tAMe6giFygC5l/ZQt73iPtMIX/Oiv3A
pQCV+dA9vDq5691m5hedv24gH3I1Soq7e5HJawVc9CGadk2GN/BcMh2ZADS2gr3y6rD7QxpT6nfk
u1l3Dw67IrOJhwlSFtRG9OoVRUaBDLPmvYe6I37tEKWpEIn6bI1Vc+FetlfNBYATWfg8XSQuROga
LuBtzUJ0hfbxv6maeQKZs+yKO77GIDEpI1GmuvPmQUiHWKsynDHcGbXDL3iDsSa679ZHtcF3E2Vz
1Ig8LqOWKg0yTrTGBUKynREKnC9HHx2qVZeJVEb0+baRluFFKlCULJE6NOIjiQNJe/AL2Xgv3Nyf
50powMafCPFZTmldnYpqbsaZySiOedfAtiN34e6Cp/MnXBMZc9DqENx4564XEDLv1x9II66YB+da
5rG9UmzEVdmSLeEkIGbK+TcI+8usCbljLwLZWfrW38P9GwjEZYmm0M4US2AZZDciL3xUSFSKW1nv
qUtRN3ZiiMpl8FPH3QLEpRI4cS3RFP9LRZAwZkrzsq6YCxTktZ4hNsAlBIwDiGJPM1523curBNNg
qjCcm2uN9qssP6EuUjC4eLFVn0yVJIcpUKrkewHosGGQyJkpyWqloZ9o8cmvQW0eKkn+S5ZaFa9x
I8pBp3VPVJPp1icC71WH65Z3jmGZtsS02yXR2S9TwzpWoZnIu+d9VrrbNDP7CpbmVDlKTcREYWT5
OTwl/JckITnpJ1GBMttS+7TzqAQbTi6VAKd4KPnNUE34lmRQx8U9xU9UVK9j+gTfiSQ3E/yadsBs
l6sR8ycub4kI6x+G3mqd+kxK0EXo/EqYRJeZB6aJ0YzEvss/GZtlzh11qupC7ayxIFyGz0S4K0WE
5pyRYRQkEO7tCbphNZhPpkbpeHfbBc/oCPfGH3E6cj4yJQRvDF6vh4UHqDsK+QfWt3p9429wDfSm
drE7Pzy36rfmlJeXiz5b7qrWX9jlQUZx9RKmQ7w1vnD0djpxusXmaLjwf1x/w+NrTPfx9DkQim1z
sH/RqZKGCUYEDLyr4EGwSdLCQ56Y7QDwxGlvFdUaSgIDIazqXLwRK8OBfIbPs9YmWfInXp/sQVVS
V/tT5CX6YeiBmw8PruIh3SfPrAUHl9fRwqrJnciPPENlNTMdYjlK/9uKxxAeZ1ij8giW/fSYmwnE
YfxIaIz4SNAu5dxAh4YSOTbduokRCCn88erDBcGWG2U+u0zIty1+LOFX/wlEwD1Ueiqx1yq6ldzj
Qs425qbXlVokCGFh5KSiZl75X9YK6RahlMmSp0CWEr+kIFOIspvbEEyEdHz5Y+Rn///lEDO0IfYq
yxiP5C4Oec6Jk1+Mar0ZzFhgEi2ZCH2gG+qZK+cBdWlLiJGFOrBhhKApAW8w1JPt9qRBQ3kyjXSg
9TmXII8l6W6QPxCBieGdGTJaLSXVHsKYSFGwa6oD8CcSEkhTvALh+yywlGEL5QcCYtUbbcp41Ng0
frhza6Xr9+pN8P3jzcN8CLHtOOUYB0/ll3cZg5/vKUxKqhF0szrazuTbEZYio2jw3SYsVuJt6djA
jiJh5RUIxQ9IAGcbbE+cMiraOlSQv20Vugr1X6Wh0RTI6KdID8XUwY8xpkQ4wNntWpV29NPAzgah
SywBFFMgxV/ZxEKM+DWxMKLlyZZ8N4HOD46E86uJ0i6dGxHF29p1SYbo56R23NDjDGJuw+LrLmxo
EkjV5FnxsFDa/yANh20do/XgjlTMG/F57fv2N+ETd5qseoCxH7ug7glAhxnPFfnS9VBzZmoSIFPw
SotTc9rig1LBOYNaeDG0TAyHoXqYkANzZf179N36VRK20G2ajt+w67uOxuQMFT3krG9YuhHhq7ht
ma4WjzpDHaxv/LSRA3RYq91SAd5WgJasOqT6s4FvjTRiexG2z63JOSXDyCqHnyQp8zP2NOh+Y44M
jeAP0mn2e6VR6EO+8z6p4f2CvXXuklG91VX7zOYb1Nqi1b9+wUDw3o5JJRGCROjI6IHmkXDqaFmc
LkVObFQjgmbXbuu+hSiAKS9rq017SbAo4VZyru+p3XqFTQ+hJyEm9D0WFvs7iWoOVCVSVj11k2E+
g0fFgujOkaTBLTfbpgrNu5aNizH7MVWT/q2HA4cGf7EoxUkDJrvTQN636kmJWgpAvxJreLpA2wJw
KPYU7f1pWtdTatMaahw/lpR3KajykYV4OK3uelqGOnHrHxa7rpE5EFxWvQSQls9Jf7dMXOmqORfD
nPPjdUxspGyJUH/3PnfxCFLZ7t9/zavmhENMHVUUy4NdDx6qeNG4NH3xMSm/ahGDETohwGXf2y83
SnSuJ+r0Q6whqvGJrwm4p5cefs9wl5z+gFEPbfXN/syvTiLFDlkQTpEnH/sKHr4mP/S4aoQah4gf
4NM6Ix0QJWxLEKwbJHU8xP7kCVN3hKLmmDtWCM2HGfdM0Tt7aZURefrUAFY+/XX2YnrvD7KHc/52
T8FXK7tSMzlOhDumKNzbR3PT636ye3SdhTTz6Xb1Ueh88gCDq0C76Rs3vvtc+EARWr9DGPNdRYR6
Jw1L+TfO1OLTKGkNJx5U7l4mtvE8+dV7z9KiqBPRj6WEkonyVghXErckvXUB+rf8x1soY7RcU0iZ
mf0Ufk/mm6o+BlG4+V7J3kEeXSSrBnJ/o5ZDASvmK1bge1lm+qpmYqt46Nv5zOpgNDPyiz+fffMG
gWFj9jlP5geQ+7tJTBUgeSRSsEzX3fiNXPbvW9P53dqfBrxIIjfz5XQGRtctF2LMakUME/mhAuKv
VU2nRz374uIjEa4fUvelkXhJuR/Hu3y+p3EWpHck7oyL8MwdhVKRdW6EnnAGU9Oy+QA1ik3FrW3E
Q/L2huxyfwHQa5qhUqfGOUiogJ2sMIyeYaJu21YrA1mVbZHYsGiw1GPTNs4RODFCN8TjVj6vRd/F
4Oy04hvBxMhNhQbq9V8bWdQ4KZpQ37F4nNGq4prGu5XrTFGQ5MN59Koti0yNK6srdm8BxP8GF6dr
88uxVaWdda40iACBPKtWfvZrKTlxiy7LfTy0hovzhdpFv12g+iLqbiQgXfkY4Be98jfl5y4FrK9x
0b/AtUNvPXBNYsjIHKPVUbr71jKkkOPSzIFzaiVUFQWEMb0RrUyyAETU6DTtv8u8p5UULMxVmSe9
I6nXzCWm3MVf6/YaRKG1mMC+Gp+62wK3a6nlh/MC3mtzP2aa2mv6kr4EdmLt/kHIjjb9CrpnUsFg
P0Tvv9kLII+UNJhYtMZ0AHIov6Sm5ErQNanTW1czI77W7qMpLL0Mea6VqO0mto5Q9/D+JfOypKb4
QabU4TqginXyfZvBhoitldqpfSvzIWv9l3hEl9EuhJ+zmhQGpV7DPNjE16EHi5d5r4QjCWm4GZxe
1DvqjRFahXFGkYxwnmufIt2zbuqS4/tiu+8JyGjJCvDb3+OCIzAbr2jURRWxl6ynBpmiLgc185Fk
HE/BDxS+BbQkwZRyGwHQZ4nKsHoCzLus11pspwksfPQ4Bly/vM+WwNIhrpxzWZpScRKqpDZxjI46
db6Dl0W7yFk5IK11L0Uy3bHJYJU2oakgZKqtqDMBwCD0lDTS7yQWQSvZpLzUEkSixC6CDs547v6L
RjKBaKsCBnzHfwb863aQtNiT+sokz1GLLfc8mXxIMJLZI3SeTeEzpZKTAUdiC7e8fE1Wis/3pZZq
XfdY0Y/WGimKQbjUhBiBR2P4KKYS0dkSCT23yaPHVbV0a64Oj76+/dVhZXZsqiIw6QpXs9ajhkaq
g8m8Oscf7cVSFEThtggFfiCBr/gVFnpK1kQx6lu3+c0+N9JSwFSq6Gp2Op8dtjLa+KVIyGAWvrZi
05Y4GUVtP4iNb0Ci9ZZU2UcdaWwe1iV5BnWnvsyRgnAJdGTMuw5bb0XLcnFTyktiG22wQ1Ub25in
Y06B4ThbO6hMd5jHVZ8CuH8+uRKd2J/f5Q158BECI9BdT1CsSd242Zb7KSxqkuZKD7VPbAw8QJBQ
JEUCIfPZUiKC9VEsOaQkguZPk2amvI6gT9TNp3VoSyMdO4+E478hDe/Hgjgi6YzOMfQbT9Lhs3cD
Ma7SlOC1qHhZGquHKNZ3GvGPN3qpqZLN7x/T5h1kfV+vGq2SZhDuk83eClW+CMq5wLcAQAxOXj9z
bfLwUohLZH/BZe/yXwUKCIpRSxiLm5G5S0SQrc+dbZfZZn2R2ssXpy4/YAYu1a041wvstK4CyCW1
dv8WWU8u3hK96+pu+QCNKLcdD0YoIZFSxvxUE2kd3VbD2sHtuu4N3nUeOaAjTrT26pCT0B5BJhZ2
kxm5yXmBbMDWQg5Mk9ycpqGeY8kRhw2I9ffQeGYKh1+UfFB87KFrZBSdk7K/31aYlLjY/u7Z4L+M
gfaksj7qC+U7ucSxzyVEyKaQyS2YN4sfZXEYL+rvvxbfoZB2DfGz3hUBZbzJpV8ABOLG5yG5xeLL
Fb4yBnfmNRCXi4bi5pSfSRjRNqlnbEqvGa54LDhrsSstvMfiRajThsmVjoaH6Md/1xCQjnEQqpZD
f1Aj6y+k8FA/s7mDPnV156p80+Tc7Mdcf2hPeVxcuz4hWcDUL4HEscscoKu/kWM+MRHyWreP8Hs8
ZWOvwjYMU/rPluJWWYrl2/gkU1DisA1SZlbCmxj6RCpfTKdSei7RDEvK+nq+kUcg9qi+0iyRmDVx
+GarfpuLMHwnB65gh+oBUDxXNbtPtWJyhNxq1ZcjQRHmhjpS0PELrWn/sCQwhpiKHlCIjOKZzqes
h+NZtPO4C6CbNRhUmgzwXA1hq7ObH7tbIS+d9JLmYfizADZuSiX2/GoBXZI9jDZ5Gzb66E+EOuBx
/fvK5OusbxGDuKbaFXiJXQM44cK06cKzfUkCUpj9CBQu//ybVf18C5xuGnIQ/pSJzsw2vtHZoGeO
VaNY5WFdOCUPbDCeuOA/2I8dV1mmvqipPdaNmiEIEgK+HLJVrqe50q0Q6ItkDwnvimcU6FTM8si3
0VEeyTU2axd5XnDZ3f6M8HoroVBa3ujOmLrymKE3q1Ll8MvPnFVBuOd/rr8KoDteOdZiiZxddChW
KEoWEcr4oYDQtsWJTLg267Xo/ADdrjRUGWLPucl6f2I08HaVTPlSF26rdh917HriXaddAXzrZoRA
EtDKHW59Qlx7t3Xf+T6xUXkporvgeoeUpQyK4l/nFaKmFHWckRh8oQQ9wCnuH8ykQh12ZwzDw7BF
yPicsE2ra2hdEOGfT62kYu0lm8lo1D16erORZW8f9d9OZTjCLrgBLiPt82C8gnaFWTjFGvIxpT93
CUiG1/rnTQ6RxiomF8pRV207XMDHg8cMWyhv2HixypGUEd2X63jJz9uW3qxHcHwCnLj5C0kL+Svf
8uzJ86H/cdZmF9/+w75a9E2U5e1v5M9hnrs++9O5LAOdNkKe73vynq4jdCs6wuZdfLdNAzX7q5JU
sJJ8/Y5+RTCN2+VrY8VnrrTRZJwLUDYne3R9/p2UMO4u0J4f51yMSrHNGIRGO5jf/epga9Z0VJiT
La6mb5OpFZ1nlsqKRSlQoVzsEdEfrnV/4flUGEGLiXRwJPrvgkYujzPzMh1NayN9I+ikRkcUZf3H
CqTvqK87/BWWbfEr2rEwD71pJB8OR1xzEy1DdP/HDtFc4gSYtJt1oHc/DPKQ477AxnnEx07UthOT
1lpU9kDJ2mJYizWqWb0wNwovs61548OglOEtClH24Y+NbfHQRd8YwVYATYLF8NDY/BRq6wZWx4H6
Z/teUEHRZ5f8Wr1v6cZqWxYby+h3daOm/WZC+EMLiaIyWf0a78G5I3/HI8ELO6AEF6QRppCr16wo
UCBJQXnNHnyTYMUXXjTPqpeCgs7vjnhHg187ZkCGBW/Fsc8bh2yISzHir1QWkKtkIdEnDtSVnF+R
+NxFgG/NARvEStFo5E91gk5GKm32kXTa56XUX5crktlL9sVK+2ejXpOoItb52kJW62vL2osI7MU0
Yn55IDKesy7f/gLqL0A6BOVwLzwR9tQOhXsgmXEVsLXf/k3jkC4MBrD6dWXb1ODdeX60O45y87OW
u/jKaCKA7ekkArkPf7O3mLV7p73F6NFudP+BNEokULgyBRqkQGV2fYV+oa1D1E4dwoey9LDNR+1Z
qkw2S0c3dRLake/9FRmLIDEg8lw8oo2Ul1CbGfBHDAfjdKrAy7+GGniE6V29vg7nMtghDp3kUfn3
XmhNGtlOsWFV3gaKYnMoNFtP0tXilLIrX1oe0+yAsQ/lyl86ZJF52tPxd5v9tJFEF7Dh6xwrrnVe
vJWFK4+/qv+WUh+IcLrHP+DcYjwwODloUdHg7RPDgvHiPPoZvJ0tA700AJNFNzBzY5hy1E3R4SYw
SR7ja5qdGMeat6KeJa1taai4ELRKv77MD/01hIt8WcAFmf0jSgUtH4MJGJhGAJgp06lnutqQ2aqM
zpxF0BRUzsTAnL3dhH5YJ4tWgDajBSGxziDFMAO9jqLS7JjFgiITd/OC32L9u9ZC2BqDtZ0ZatzQ
JKzJf76BOjmiXOaD3ThQd40SqS7VrPaz8i2zUmX8KkP/F3+wPSajhMSdL7C1hdU106b3Kh1cOp1X
RpWhbRCs1mRTDulP+PsRkZB0W0lcPcpFPkTw9B4ow4m9SdSZQAV5n9qqQ+zPZTn3DAqdQu00aOSt
rOOv8A36wcGyQq7fCukudFpPgiM5w0YTWzF7PW5nNKeolcNK8uxxl1CEKPSJZ25c/WCIMQoNn/23
yqC1sWQvUUT//P4EQJ9aeexfAU7fkPsdFSB6gdmlqxHYVIVmSblL2T6cSv/6X0uSyC+LVeHOzxiK
GIznNcfBO99Nwk3sAnCDS0ouxO3gEoxoRrfE3vPg0O6vH9AeQ/8aVAUmzeG90Z53FdawmyiDFN1C
13DGYG1UhOLXFAeENaPEC6xfokxL4DLF0YXRcsI38W4JhdTb6JfASWcaQObPnnn0Zh//z2NMyaKf
7KactPlawbj5tuZSqbEQjqceD02E3tCkhWG8aEG1t9cxua/oUK4/Mraa/dxc8KPNmKHZK+J+45v1
rsrAMGakUgYe0J3T0hBQ4GGgxqbtZ9iUuKqReW3hKWxk1BZOaJ2gM2U4CkNrK2MEWfpp9YowL3K4
wWxBUgxqSBVjedC3aXI/izlvaaHyt4vGcih8gApcXSbBc45Z4aYH3bYTvQoXnGrB+1k7Ygc05M24
kba/6x0L/QPHEQg92mn6TdAzQBDjR29lE179jjSFpiQPtvNPiaVceoGvqLHSbldEhrfRw/GuT7To
l4PAYENxjNCBCLSHXMV/7aTLvqe53Rm9PseeMJ/LZK/n8D/ekwDHC2QilqfI7iS11NJFweIMkANF
gpgz3OpcJTFcnblmYqZQhr12sgzHgPN+kfePWqo/DKvxQ5AMSbh0Nw/ilkvXuYXQ/pBFNYvACs3W
nVwF9MvFILO4daz28EuKUMnZLLKY8uDdcUFguL0ZPZg2KqOEtrLjW9PFvpJKX2EVZfF3WYxjSWR1
n23P/gMyRdoa/5SE35s8H5s5EG0F2bsctKvekgw6eIN0JFErUv5Gtta+TkrJxFTeGK4/VhB+e2Q8
TPjbSCjozaasY7rclUa51ufia5DccO7dRe4NQDdYit+meTry0RtAlIERAA9IXvNkZXAUzXnyOTFs
XWjN5fmHeOhQBm9S3iC9sPpS1DNCy3cGCNsJ/qRnoVBVacZ+XHmqwv2KwXSWte93WrahESHfgw2s
kHYwcfWsh5DDJkGS+TkxVLsEWgdRLjpQrwUZ2/LaEyxotNxAcWrvDDRETiz0vqYR4vXQdxvyItVL
J9cdL9c6uqQYW5Cb9S44RC7ZnWIqCQLe+ax1rVbgNWhFIkN2PEyp1W8CIw9CrOJdCpCg83AkYMSd
afkdJ/fdqYvaeA0TaPb1/ZQDyXT/WnT9EmALtDLwSj5T1RSKjbU5HM+d/Z35BpAvVJlWW9eLkYoa
Fqzii3CzfQnncZ/6Zsff0jpCrAH5CO/kYcfZKlhp6MujhFzIcQsRF7tQno8cg+ovBGBeMXuJyig/
ygwfMNvceEMoX6+vVYvF7lXeWH3HvzJgQ5G8hgtAzf+h1hOBOepGVqVmTqTBw6/5HqmwFIJg80t5
uRt1fmKzd4Jc97+M9XwJath6pGYVDi+uXi0p2CpFsVDZqDuOUwnrWxU8ZWN+JelRawvitnHzFtdv
wNAOJCdAvWdhwtf7Eiiajw+C6K4hYUArdEIimTzAlW8fWP33xHnKlpePhkipim+AAQAd0MIvT0rM
yTemECTuwmVwaWr3EeqPqHl2Whlom3B+N1KMxHLMJB2QljevdVqzS8dxszgbD8pG4zc5mERLe4F/
v0AHVZBsQVb2jfMdmH7YKMFMHHgcku4gLZ9E8M8y4WhJTcGhU9SoIBCq+WAQnGU45roaxZ0WyAqC
e1K1IYDsIMvCHPks2tdCDlTKVFLJmkMlACE9+sD+/K5cV/EpY/3fGjH1GE3BU0ZGpeCmLdy6lNrP
NX7dhzV7KxMz3J0NtEhKLAFZzKUj8ebMVtW0CJtr6uanLMVWY0Ki/W6QYQMJ2aYY4To5E/N+5oFg
lEDDu/aC3jKPWes3Y3SSPRp+aQ2eqU/65qM2qLDJYiV1YTMIINIqh+l0sKxIoUED9z088vhQKOhy
f7FNykw7Iv1VjdNJOoD1hXVC6zVY2xkM/sR4WdRFyF3udV1Ct6CCiwQWNs646fHRkj7xDf+PYOnN
UUe2KQ0bv9PRxyYFV1xdwhmbAhgpGXp4qn/OgEdCPEtCD3UIJ2OlrECSl6yenaO7FUg/YQfrt64J
ymZyLBlRMed4Zdv2yrm5yidfsE2tNVqFLYwVMP/gu5JOd6/Zhck9A6bb+pJUXTqSA5eMS5pS4tVa
JSsSNmWulaUrSWyveRtFkDnQBHW1QBP9CC2DauXi1kjiDsshjXVaUl6HXsJcyMfYQZQeqIuUegTw
C0rt2mAS4ToD3rDL4wsUQcsYUeyfjJ5FYexj/1LF20UFgFuTQviMpJ7USwk80KMxmepvcGBvJAuY
OFp4/4Xk4G7bkyO5A6BAF50C7L+hzrgLt+z+qxTPAi9ylq5+PC9IFpJBOHnHScCtksP5ezWk9+vz
5tsbru0I0j3eaEHtrVxdIkATE3iWIvgLr7/kQemOB/MeTGL7HhV5OXJRI+8+nb8nhYb+Cu3r7vCn
QoS9/50sgrHPAxpWImlTEgz+d/YdkVKLG2byS1k+cCbQygCIyBNOKAGdCrl9fD1dCKpgP8Li/Mec
nYma+F2Of4j/XDeSHg88N4wxBlbKPO3v2MXvHbG5wH31LuU49l+irNd+/8UL4gmWlWAzO8tAry0E
O3ZecN6WaoJgqwMYKV+akE1944Tzv9bVIYfH3z0cOohUClXJEEA2yPjubnFykONxgr247engINnN
/zja/pEUQ3RHT9dT1RBOGfam5FIlrddmjFCeqLBa6ASOttClZa9lW2boySxfXlJkUqeOErI0wu+U
dRlaa7HFWesoYu+qzuCfafMAs+PFsqUHalCuDRimMxe8EGPPbvhK+f/mUjOATuh4pFKvbAGia9Dp
HVvrPH4iwdsHzq5xgGFmCMrALw998gt/O3sfG4P4fhwgpNGaV1QrUpeSA22ybrbLBGHgzNw836Yh
P2DpjAuzcUyYu+hH4JN0UVZETDl2Q1FOH5QG/UA8nWocSABWyZhD80np8+f6VKQ36ZmDLK+pu3NV
aLLDbMBIxkvjmvAiNj1fPU42dhLtdNrCwTMzMuahw3cZlOK7MCLeFEf8UgNYIvEfZkzHMeiCmObq
At+phM6XJPxx5mw1HUhiRh/Fii6t/pITIAO8spz7uIJQdEa/u2G0aXmAR13zJ+XH/kW3AJUr2DjU
ewKyBSh0+1x3OfOcFRvfu84aQr32SPCqUAeQ4atLq1NoYJoIVpZM3sE/wUb8bS99xaoj5vc0E9+X
JuhSfnMRU9OrBrZGIleAe3F1tN1Y+P5H8CrPe/hVLWBRX1l28kLnAIzDN62lY1oeCLO9LsMtllSr
SM6rswGwtRhXtjwWSJ7m1ZTErbNFyrVZ3RbCKfLnOyuBJ+n7SAgB56d1iNFQmMbruzPSA6ryiRDR
MV6iTirLDd6XoVWRqt5OCbs2jMxc9proiacdki4whfAD41o3WUKBGUPIDgeaOuCj5f5QcrgPZL8S
ygUpqs5AvcJJ4a+KDchI1gu/457wwOBDPbbbGbHjA5RWuS/OogwpkP9wPNjIaZjr3gTzqlx1Fv/0
MGCrQd5YvD2HYDaD5UzHQza9D7biuFvqYRu7+DcVIBHkXszUrlqpmig8Yc8Xr6hNpBcteOIVMA0+
F2tFfrx8YRishWYBLC6/ullPM36nvbliGmpCeiHYr0gwJscOhEKJZiTIOOkKf7pGAdAgndEthkYd
rJjO56AOUpyXj4OlZZMLOKB7dAZ0KM3RszcaLDl0gAKGsxVeOuZVWB0wewdr9rB5VxSbX8CA8LOE
mFw6bhRWiCGfHyijLhc4ZP7M8iZ3JKpK7hCwqalWNG8m9UM2RD2p4fT9Df4eODDD+Cna6uUbsbMX
Ugzzrv+4ge2GkAzn0zXWSDUCTV7JCmnSRSfr9jknXF+zjTJSzSwqUFP945rCTm4TFoJ773U0jeUf
PYM/hRcV3Z/wByhQa75IgVepRFYGwSpHmdN8LrEGzeaPapCqCCnuynP2M/ZTlF+QhM5kWaTsUpzw
zHmpIl0Brpl4N7gjU8UUfyCttixQErBMZnJHMYzAfNV7AUNEEPgw0Qm3ahKQ92bUrSZWtdpoLeS3
0Bb77tbrQceslL90GkjwjlyA4s7XMzT4KoulnnWILOCbAV7ySsGedcnlR+tb/tbvwzCF/VmKhHQ9
dnBs+N+tMnNF5dWbgW2NlJ09CCT/VFfGiH/GI0KYimarLyKyq5Nl/Fm9Eo054gKwnsk7VnGt9/qk
FYGZ16XpPizeiNk5CHMKOjRCT5kdLA6miiX+kAx5WLFi4WlOSZABPVx57cPbmek/herypuCfiDCb
rZSq6mCt+CYS++IETFn32AfizAfRMPBbqg/70FL+nJsCQxS+qR0ajcfEj601/2mFGoKnK2Q7vwn6
nxgvrQ1+XN2IAwq0xQpa7iXIIgMuKbNhBgzIBZkMuW946E5S/a1v1tVKResU7azOs9uK5LThebcM
/Q/vgSgbWPFQWWc8EqLuvw0dFcHbuMDoklYH9CPyiwxBH7V8sqPuFCuugAdxAih6exKds1IU5E1Y
j/H3C0PrLPu6NnvYyJGOTpAZ6VJqnqpRdf7tbztHYFW8HKstNLejG/HMk8wjVGSLihjTvTQX9rsz
WkLqJuUSEz2Km/jDr0z7bOBKuCIITi3HvZtmKO5KlyulLqar9jkA+EfVJg8hBoX4glxUalnW+3He
C+C/6hMgw0aLt0FrRrlcphgGtFWJSZnDCpkYxe0C021BnqRDWCbrDpDne1fGFunXsScPwBOg46H6
Q7+nU8fZjkZaDoljN6LkmSV/ir70Yo0WtVY3Ajc9Je8wxL9+Egi0LvxCGd/EIJu42qBQJjMPIdpf
xWoEeLKIFKba6d2sab4bEgXbtiOi+nlTUaDVuU5DHL8gI0IhVjAXXiIInS8JK6DBlxo5YkAzm5Y8
darceoiAUzTGKdiuJpQKbQhs1hc/AwnxOElieLVu+5QmO44ezKisdZMvyrGD4F8fimwnAPoLzDQQ
UvK1Idp49D+UTqfdhNLXRAiINvfpcjYy6Xw8sxxiFOW5aI7ASI2I6jMtv96a90HbnY03KUUWuMfD
cP6Jt/yVM/JtVJKYWZjZbwYQoMyc+4kO+XvEnU1lOcdnyyz6Jz62aOp9IsqWxdCvo/WShSseoAYv
7/MGPRWQyS2IYpMyikYU0R7xxz9dXvH/Jtulzcc7KEI5FvRmqjP1mnXnYFKS8/0DVJpMJH/1RA+J
8tleHgy3TkJkJkxah0ybJzYIDKoGJ41fa3DUSJ3zczcWspS4XGhi0IcINcfc8Mc3PuOhjMqDJMTL
JM1zg03p7Di80qXIYky+LX2jGNEt3KTqUUHQjSTCp+vsI9NTA+wQ2iZ2UBWPtNR93MkgOHKKRLkR
OSTMvSsmVObtvhV4DF9zCbps9CXFYBiYuA6rhHqaTMddolP27YafgFct1N+m6GF/1UB0uTn2Xmex
6K1onL41Rk+YKN45FnB25cp4yh2GcElGy5SqUsH+X1cflnLu9I4Y7Zf5CtY9FUKPt3lPnxqFlrjS
4N55wXJhki0avZ66I/D2wv0Qs/djzoSj4WfYs4sIQclrsydZXrB4+iR6lPxWWrPtcFEOZI6x1xfK
TbnycBBcjglspbh5YKb7SH894N+/U618+8m3VoJG0/TBgjpbiS6u+T7VAESbXT0zIjtn0yuoH526
885Ly60Iask5sDhyZl3f7rPkQD82nk2b5xnKWQzW6NNHvzDVmdHJOjRoimu9rwE2xghwK2YDSBN9
dXFFSthmxaGdZ8qHDxGWDlAMKXnLqD5IanJhQAHcg//JJIZXzKdI7eS//fOTiX/wg2aKerleXolA
qbXtMChVXsg6QHYtViiqBaBfpLQkjiJQ3yYmzMmXH/ipfvayOvTNdzons/58eOEfrVDGxIarxSsq
xN9vYr/+LkdWp1a06JOxK+wBVj3tvlsGnJf2vi9HyiexciCuP/1dkhrpeptUHukdI0Yt2sw+dGFz
kyqB3DdIDdE035/r5tENxW1dOA0WxP76QYGyEO7yRoAoUMcfaxUuZXTrjqowFQl/25iWyOK0cv7o
xSHSQTPnOp0HAhwMatPf6uyEfd9zKQTOIAxsrkIGIDuNTlIOXH1/q2b7G5sAIukf8KwIdzhDp4JC
fWY5PrcYj8PhdMgPUNnU8fB+ogtAXYA91pJeJ0JaESEwv3Lzr/5merbQl6zmg0S6/AqFf2GifeNy
8lIH0SOpsN3HrvwQ9kO+RDineeAZHP911J+4As8cVahjyvBOwUX6e8LKfhcKINU98GYSfrxznDu1
LEofBXwgOYJqduKRFP9fL0bYgl3YANtQljRr/2cgdLW2msbnGpfMJpxIy6XIYM2darGbdbR3OKGm
b3YoZR+yeusBXM1QQM/uAy/KxwOarXUdppVo3Y4C7asL8N8uFo9sSl8Kr1M+KYKt/AqGOEDkjLZR
3bykJjl0K6XAy1qmVsX4cqb4e7vdgskrofY1h1bSSg1eMlIcJ5GnVw9OM2x1W+agJWl6nXTHk8Hy
qSk4w1Qe5FZbgfgVKPDWpD44EKNAZ569nbVI/m5kY6idNCNlxlZofMzbnxq/V19ayWhbqW+DCbyS
Jq/R9hnIsN09I9KEi51m0uNkhKD2LAdS6BIOfV/lU7VFUzJxriS2nfmftbsYgq47irrBmgT5zwxk
IyDHPi9BnNLg7O/2/6sEd+iXo1Q+w8EkoK6xyKHjmmkO4l1PfIzlpRsq0rGpQusgnaKVZDjJem5p
NB1d8LBBIz3scS/bxZTNWkCVDLt+1ujI81zM9rtCJU5Yq1NEs4IKur3thbQdEBTaJ0kHEEQBvkbx
oqsQld8UNZxi/gGXCyE9IdRlk44B5rR4QO1WaSandfU4Fk6aTORtcMgrEbsgn+SrLcDapKnK/3ee
B9zw4SZkgIc5QtuXJ95KY7mOjnEQ8P5XmSiOgdEWRi+yeyf0KH8yfxW74c/hWTYLnUbI+e7jFcvV
9lDivWbCJIApn5UNaPig+hIptcg7wnNckPpU1T2uVG7ORa2pLmF56S6FA1LqFkPatc0Ez8IXrUhP
ND5uqLCA8Y25i9h5mDbV23kZkA7x0n0Hzgf22ndlNIUKCctETV9oCBdzbApF1o9ET+HftateXh/e
E+6yHpecPPIaQl1cAIrYqLeaFWPt0CIX3Jlw/v8hNKBul8gYeOqq+JAERvLfyxsIdWsuJGcQcsqn
W9ftThnt7BKzHkU2rLK8wTbOjObsJINZpUw8eXk6InnmCaXlepJT82BLOP6w3FWwACzzedR/pPA3
kHQg7W2y/BSV6KeAifEAakOlL9KqG5oeyoB/VgMLliVtBzsMMJcixZE2GgPhbBYNMrd+2/h6hDy3
YKMt8ioJxy/iovzEXBs49+HEz3rJ7MPciH4vRaaSh6xRC214GVWsfOvoNPvS0gdmqqhIK9dn+YCl
df06XQRXFrgz4+3gl57wXdzpeCwWzQXYn7UN2Z1wPmS83MpvZTDDBKk7SKcjeEsNdzYvstZNx/pl
ISkfCuwGifBpbphyaqJTmSxeu8oWmv9MbHVSpnfdyz/tISaN6md8yiyCKC2gbOAlqoAppic26q7m
htfI4OgSrjSStLbj7kZ7Cpca2pFq9D4RgYwcBEKYxXOX41xsIigMJbF5CtmjiYeQgJ8rZKHGOU07
dui1m0Xez4JQc587ZxC+0Y1x0PUg2A1suOwYLlZnGcL91kM42uMonY55sZGdKaijOcyDCJvOeCrK
d8eCEF3sNEA5DxqjGv5SOt2+U3brPWAY1LUP5/r6VyF73SqFLl1H6B+G7SgHmsuzx7S8OV/Ish8f
b3wa6GnTMrAaxtjn5eBy7cM5IQKhW9CZdIJEz+XhzT2IBicQIE6736x/1VdhZwC3VmEZwQACWcIL
2W2gOCiANRzoa/EGsEHkX+eGEvLZG7ot34+J8z1HIZvUklfeZUsjnoUkBABEUUAf/hYdGSw52OXn
JcTA6zVU9+pVDgUNwWovz3y/ByMazHrAiu8X0Q2F50Yq/8YZTRgxKRFNwINE6Q35FrHetaCwT+11
kovG2ATPMgp/XSJDKLK/7HI+XaQgftC9/zkJle+r8sdJ3brEhRU8NWD8aA2AHWgy21lJVXslZwrO
+Lh2VeMsA8GzcINQcC+SJttzDJBhK0rwMhcPP3uleZ+06XTYjTBCbhJRmdi5MYW2lfaUG+05dq6b
fCe/PmG9Z/WxaTg7IJSPafFuJnnbEp4+fmNmRxF0WHCRg+VKGDTjKByYXRCliAfpTz90uwdjOX8G
nMSD7W5V3bEQysASqg+SRt5CUCyq7BZzIjBhZQTYPQM2Kv7zyIBbwESqCkmEL9idxNrMvekmMjdy
aR8P5nTGhUwN1XfAMNfYlnxHmgeF7b0zQC4OROYMNV0aYSZ7BZPuGu6B4qyUextSJ+9YUFC1OwE8
RXDreajUqfDJNie77IUCQf0USZMbZcMS8pHRd6vwKqUy7N4I8shQQlWXoJxH7UPHnOhkyD2T/RMb
rFPzv5Cti98QS7D8MMKHK1D+oIR11csevYnIcSPkkQ8BwMs1Wb28FY5RjWEi5L65kHCxf1FPS9p3
MgTCtFW6AFYKvUVwBqll0lzZrQoRBlfGMZi/uY/ktZPBKdPTTw0JfMYOAz/JDnfP/gG3XWwCzrgB
o+baGxiskBGtOvgKIVbbwT9IXxmZDhBIvuo5cEabnxwVClwXvmkXv8QZAUOEZEEFm6+knijb0Zkw
LqTUnHR6eNdGkE8py3INcCPFpdJPmDDJ6PbfUk99oSpKjlR6DYNVc0hM9ivUhRyFkviULXTJuXvH
LHy2h5mTYGzpw4V+8hzVI+WgdXl06cnZmGIWp/4V3Ik6Iu63Brz0INAtdDNo2bK3mi1NsawhH39D
NFY9crBJu/ESLYHagh6E/zpgWTEeS8u0Ph5nkBDbTYAoUibSUb6UdbUisT5rxku48dFop0h+D3aJ
mnu3uZfaRlRw6cY5wp/v+381v0F9QGUU2Pju97KmhdevNBbwAMKd7KUM5462nUZYgZNxsWVeQBJP
JhjUmDjL6OfOKmZqb6lYkQjcrWIDaO3/hqs8mitNcH7qkdYEDI4MJb3QQ2e2YyvYxX4giPgeZEHB
QOYUbul4qX2qHJ6ByKrVr5EI7nkH2eYAe33gU7LxEpEuZ6LdbhI+wY/uUabgvjGADsTkPysh3TLd
v4tg5f1CpgiD8R4Atwxm67hMbsEX0Osx7GtNgw40vmq1+McslyrqrYSpZVF/VaAbyyl9El8PR+74
t5qeyAK8U3bzYjX4CeghJ/Cp9WFjljeB5UDY5r7ZntQFomPcLs+eRxWLwU3WxnbRqCaS78Aykea9
6nPoSJ+WtdYiuFHULaIoeWGdEr4uQgfO53h3APhquqL3pjv8ev1gtUgAAwHk7Dq2i8XwkgwRz5DO
hUNoNVTxKkrpj3i20vtNp0sUOGl6hvdnt3tCfzsXoHMmgw9AcfPao/ehO83+eP0E0ztsASCFins8
bA8o/FUsZWDcW8M1KsEFoYzmGgaAjLlO/ApkuxRil0I/IzcmIA7UGl2FXeFSV0mZ/1D/6O+YcR4d
fE1FHELr+Kke7cV9+5rAcz82d4C+A+EvGWCxkhORRF0bsUwNKZE90Cqcn9VOJVGG6j1+zeRK9rFC
HZmgRTFDPsLgfVmjB688nJXIMIoLeblXASJiI5Thc04mEST3ylq9E3qHeFJ6PedkBXlvFAYcDYq6
wXpwKE2+1xlQS+6JB1mmryeUzH1cseLeboyUsGIXvqagmXQvEhIfm3zVkn8OTbn1+Ls+gYtTxS/M
Ad++16DryWCmT5zyCkWFXKdt47fmy+Y6QQ+zAvG98BAL+249/lIBLvWudcKNJPJtpYreu+Lg3Jc2
fVMSs18uieZ3MmNhQJCHZZxfhjISBzKsvCB+nx0iTWdSC7bC9goNtdgbKHguVH7lU49K3WtoCOcT
pP0FerVP0DJslh4SSDtHMsNd17MmtN/peZBjyG5UhF8y1VAzBZmAYbe8BgXY6bZdH5uvb4oqN+6E
759DBP3pITxLSFEEE8bPRvVtCGBgyPppo5YMIA5dXZ6vOQxeCZXksZhh4ozfDcy21NuRBW3qPr8g
JKvAGhdGaS1tgMcWwB/hny3nsvAOV1kMqZIrxAYDDYhkyplYGogjzj3qkrDeIMsj9qPepSqk8fC9
2VkbGVM5yk6wzvK4tqJ+A/XZDVJvjS6aHQpxFj6B4H2QsJEjEKXZ3hSScJ/dH8AuUDrBt75b3qKH
li8p26dUoWFAm+ZFshn93cnDdwPC56fFyNugmA6q36MRc3nfAuYjtTbOwUeXoEHr+yNx9lSQpM2S
Ly+ZPHlyZfsUPYfgvZPSac34QPfIuT6Z5SUqOu/4RwjWJVrecDMitKNnE3ar+h942LX9vR31BzGJ
6gtUCVIzUH5YAz3ATux71HLwJS2Rg4772i7pGkWCPGZzRou8/9NYUjfGDooSrYisORYTi6CN04Oz
FRtyF/gy2rTNLCMqGJFdxwIIhXAhZP8T8I2GxhqQ1ZNWDrkSAXNKRRSGWEofVuNjx3nzAngAxa0G
FcYk/dxIzRXrSi7xYCMsMvLJ2a030mu9HzK0GO4m++RsT160J5LW6P17+0KaOFf2VCEAjG7i0X/Y
i6lgfd/XOSvBRltpY3yCt8ctwzOpwBPZPR9VamNSY3Y0HVukFNSmr1xZ1+uiAktQv5GLMivKGl/H
P7ooN9yg+TXT0SLfBb5cmqeD/eKp0xViNjfXiVjONpfOOOr+X+vGjvTJ1GkjWjlhqip5HVq1Leol
7GCahqAy3VSVhrc1sE/SB+aK2i2Fmi47oAN9SDFVGcpgAYGGWO3dQe6UMI/k8BUUXz7pa/RjbwJV
Td0LqepBoxPf0ZconpMcnSSwjX2RNem4x4CQNqZxIuj8AyYjdqaNmrKEUM7vWXxKXTsm12QnJ1wk
bPIkBYuLh1DafQAmCk7jabDraU/4oJCloEplRxGYANMGcX2Trj7A/5piM9KeVptmjDrJh5wElX/O
g7HZsDTIDjLOimcCVBHHoOgE4h0rGUX3H9ul4QV+nBGarBbYuNPMcVy9Rv7NlHfss4Sj2zVOrs8v
/0dJrftX4iWncPbEX89vSFoHudBfSsyPUXVY8qtAYo5Cuyq/LZQeFM0YIb/oDpcw+qzot2nwMDlN
pCIANds6PUm+kk7t5wZY7DCbrXrid8+C6Qb8HTy481kxx0MK39cYaWAXFOlGdcLG2Nl1sbNK3srR
28FJW36ycAXmZwVxL3t9yKFxJJoEJ+af73sUuPMu9KUowR2kxTiHWEeaD154lZxstbeHmUrC6E/n
/9r/M59LA325zkLAhFTF3MbWoIMinly595fzV/pxOqgRjqnMXR3OGwAHbWMdNu7nT0gcLQWqCz7I
qjcrnfHyp8uRAGVthbYhW1KHCNZ29OLDM6CUKtDXudwYyk9+msZgdy6TwUXJQYla5lDqHepkrqq2
zqdlB5S/Ojslm1BEwJKEZkMUX/HmGjRHmlivwCH02nqzTI5dYhPLeTm1lMDUeSvJKwdyVR0cqLPx
lQoMBjU0nHasj12LQkcei6GBKKzG6juSitY7YptGcQA5WacagQt8SSp1XGXM3m0vYfhlvBL4RYaU
+Xp/Enp5sEhx86jDRxWqNtZs0ZQOVvQwl2CRuAye1tG/F5iqtpD1/dq1XYj7Tn4TU38RxwauXbAu
BYTWV7apcrdrCXdG/CbIyQQNALvY8F0QFfTlYesBdSu0NBVu3qNqkti43Qo4v2oqpL0rAfx1AsPQ
4bUl+eqvuqH1KDWq2zCFewZmIffXQXI4FdkuKZkX7SLJPiHqPQl6TyPphH/bNQK+o24wtPViNlFI
y/yf6GZ82ImypjKree41IRbOsZVgKLupKEnByLtZk8/KJ1G8MDXMoTX9OgLX8e12ywrig7C0RBMP
7l4tXP0K/egQMIsNy8L1wzgPmNjWZCjYfNwzECTGmmM7xAway+Bb2+NNVCmOt9Ga/8318dXkFuif
Qeo41w0DSs5bIwMCzpOtNUuq/kF8JaRBz34es/KtAC92j9DqO+rZwuSsk3A2mGeBkA7lH+j1j6ay
svr4Wjmv4nz+Ikzta5MPGZn06e4SRYu5xlocL0MpZtcEaopl+G+QWwe98eiL4gTgaPtckKmJBI9I
XT+nAHM7LE6PvC8V0uDHoC8mNqJVNqKt1wZJ2VPBWE4YgYljcAQi7HzwkFtJYl1DKdRCUSDYz6EJ
oPxP2YLt0AuOWyPj+dUJZgx5cdtVBlC61GSMyHj6QoB5Q1DyNBmJ6+yz2rTwEwMxR7GRbjEWtWDo
WbO4CTQ3ZZEkgI0bpGkBu/gchtUt1+5cNOEmtFZudZPEwekgLgq4W4VQzgexXfjOITIO+18Tyxt3
mEE0uRiq8JRnn5PwKekuFaLARxx4QP14K1Oz/hjnETPf0/Fd/DaS+KkO7Pv65euaIY+vH4b2dFBo
eFeEr4dU5Ot09brE3g8AN9sgtsfTeygQl5DVhGw4ZpQ8pHAkP6YFauO3BASe3qwf8ITPdN4gxtbh
BBUixWk1ZYOAgUr/7sRhFNhtEJkArN9yOmzbfFl+3wMg+cgXfwHaR7rumpJxGayRTvYa7gOLgKna
Zw7OBP3Yun4yitEMccN/SgWDPjWP/rbNUyFlumj59L5IEFlMnYLm+94KufBblgNOkpCtfDM5Z2YE
sS2wiga/7M+3Z62DW5IGpZaOD1V/mxMSgDSsUg49ClxZsWQRpOZ33m0fC9SvIhsKz3PzP1m32uPk
w8BiGvJzZS2J1STSc6hpi5+3hEH7gHBC3Sbe7ix5KeyeqfU9976tqkCjfWxPgUvhPpn/vz33wVj+
KDnGbGxHyqhD3Ak23MZhHWalGtY8HqpXt/rf8UhA5tKyOQZN4oXAUujOOMIuhpGP/kdqLR24q+c2
ir7VOhAdeQl+IK6yss0nAyGLG74wz/+OKk+iDUhEQcSJFawC7Dm0MGmgE5uontaecQn2cPvYtbI8
6DvyAfU/h7sYd0AxJDXkOM/o1+1bVq16X4ji1XQA9vq3PgWaLkx9DzNmfVFy6g2i0IPWynZWhA7R
kGcZPeZNvjgPDP2E8O6a2OZuzwcpVC26N0ygWc5T8e6tu4I78nzEXUVNHFV3Q2/gR5AJLJzofooR
hOYks5uEiUjlNFUjNydFuacVmF3deaMJUPmTxiDLOzSLjHqQmCMet9Wsiw66ZBcXfskyPRpiRl0x
pNpWgaGz/8YiNXUAgJ5rJISgluAFiOOH+Vdg9kcaG+pXdqqE3WGb81PUufg8KKdR2YrbCnlnl2Cb
d9d5ZX0tCJVx9k0o2xqMDNUvOanV1wz5aOc/d6wBPYkYd7Ejq8100Jwhkej8hf33ozRfwVoL1YrB
yclcTCFtI7Yu8Lvdua1LI9KHkcWS2woqGuXwJCDz6vN6OmZg1sX36jtASFvSgVlW6D1g4kZ6IsqQ
vk8Z9V+ba0yByxCfosEL3HsQI98FLGali27+BPfkv3aFk7GaxIIa+lww+5apptYEUkiy/HweGVAB
z0+PZRIyVQaiuHmGKyql9OiN69+Af+b/zQLudlA0QFnzPT6t8Y3usLPOQk6+4fiZN6WeUcb63x32
Vxug2/UDV6DtWGtdRmiMiJUe6G+b1o/Dib0UiI7HZF+lJLI2bTsKt09c0uE2rvAaPvYygzRLgSo+
/r6L6eXqwgrHow78jDk4Ngca1aILaPogilqQLvjDMJ5V6kTxdsfHcTNhCSiaBBwNw2heWx4Gdgyh
HwNFGEsGo1xpEn2mRixacP3RgUMyzvvTdUgSGnPoJVms2L6A0J5DsBuSkL9WMC4jKQUHjW8Qs9gI
blHmaUu0hnAHC8HAu7a+9p9BVa+9usjm5tcA9pQJ/YNF5RMkUqsZMQ35McmFN1B2dubCb7/+MEAK
s5klkQaQxEN6v6GNxNwAgiqBc+oa54XqdcyTuMFB53KIaqUTMoaLTf2X78wNxvsnoTwAfFMbGOs7
8zWKzZqaW+WUl6HAFPAgdXb5eyfSMFu48WKTWcNO+FYTEU0qSACBAAIrXGKDiMUlM+rjV8ZomNZG
8Y57a0aKjiNTHkdjk3k0wDJRGrS+qw9m3eRpSUtBQHJYwmUWSDNBe+zrytIfq6Xde3SjfPm6fWkJ
0udmpPyU1fV8wJXUgxjT7z8a9PNHCGdgM+07k8VIic6znxFvL+PuNBI/OE3a6Bw4P6Kpo/qZeFI8
7Sz18t2bAmUZJChKsMi3nJ7d4md2fj4T07aNQ0iVzYvaWBsITjew8Eg2A6qrvwtqfHAnDZq45yeK
ELkyV/AHRhHt9WSMM328574aUDaEUPWh4bl5YQTSP6cs6idOq6Yqv53xEmpFUq9iuNQCHgJjZoOC
pQJFFU0prC/qGdkaSL1QnxOK3tKz+whPDFKck6z8cYxWGuRvrBDEF8hpXN/gGq738yuesMDa8AnD
Ry9M04IuHjqpUBw/SeO1OAbN87hNq0iMhaQrv8jyQbGYe/noS3NP+KpO5eRiEv4rUnTwbHs18I0/
93F0LsBvfsqhHqHLXFXtlEn7w9JoBkVD/8sgcJnYkXSx9byVoE4Jb1sYtEb92KxQqoyyMyvD1Y59
TUDbFri7g9yrs6N5VVufpL7h1/crB3+o/H5ZebHJTVf2n/DZjcuibxuLg29uN9C/ebv7kNkF8H8p
qge5WR4VLpaT/Q7lgEAb6osKRALcH6jwoBlctMwQXEgz4FiG1XthoxqSHAuf1EYJ8TgtMYNEz9nu
q8BewHdo+2iBXEDR3BpXcodzalBsbBN7mz8V+HiIgf2syFbV8lrb+fl3UjPqa+ilVkBh4l4TctWZ
EHWthfQUQYc4AFhXr86W5lx8lrGVjEI/sKzdnPWrFWYjSG5P/jk/wKEAx3Zd0XoufRIC4InzSd+b
QuNkV1ScWWkvCOCVx3xmAF0fKPVxFkYaS6dUZn486A6S+PUc85s9AZrtUcHh9zKe4y/GFz2SUwmm
6WL3caCCz8FnNY9Xyn2CaUNL1aL2f4q6M8aSfuQt3ao2jM/sZP5ekjo8/EhG3e9ZbK/ksvVIGpnQ
B3veAdDllfG3/Gw9/mvMMGFv71sktk3lWGCQphPgsX5wdQFhRbvZH8FyyWTxo1FiKi8bl/35NYfc
3j+7i1Wu3mAbrJbmJi+4WZ0ZCbxxrTkQErrmYb6f3JBbVD3By85p+IevxQNWQCYDug6VnbPg9gg5
GOFv0Aye8MFmloxQMIZHjiIuZWLLH8ytBb84PzFjN9DV1m02eYEbAl72RK/1kpUrot9EbRZ0Bqs/
GBBA+CwJGzvbjYbBAu1w3LRN2uLDtPuVU/zi7RA4Hq3qZ2v9lJXHwok2Vn1hrPhpfp2lR7Iskz9U
aIFTYm/eC85WSP76upg8UOLhAExm2SVpN8pngzh7UxVy0kEpoDsyIfJpwClk8zEkFu+W2Ae5l/kM
jXQhKzIebinocb3JYGVTTd/zwyuTBm/PD/3omw+uES9u0b0bTnjKM9feIWrGnwwcALCKHb0QrrHT
jwX89nR91utKkuPRHT0NpIdHz8v10ejcFxIO5gPZfmAvzOqDTr2ErlN3SpOouZUZ7ZoBF59k+Z+7
J2UYcQH7EobYYOc+/s4RkLpNUj18zKk0vowny50qu31Xz3XqSjuwAcRVYXpqmgC1DQnB62luEzZZ
+DuXhNeiJzZ/NOSH5SK9/CEGJd/0VeOm7yJYOYBb9Zvk0GpnGQKz/5afFhi1MUDE5f12e+2WWuYY
VH930LrSYT6Vkkj2r14vF3sOzCZRDvw5gyIz1tZshoaWD0vuJ7Iz8sHIZREN9qEWsBTv2xlAvk5Z
1YgUwqqnpCCsgrz42eB7mIkKP1AuMlPa1NuZisUZT3U0Z5zrqzy2nR2Z+jx+rHCmCdKFXJiHB0JN
ulSP3iwghlRnR1/cluHyvay0AYPQYVTmVkzzHfe0FGWEsMZoZphKQyBOEfCaBLaOF9nw2sCsjzg3
xDoQ9kkiQW29FUMhiuS4k12/IYTL0MECcYAxhIFCUfSr/eyDycYGx8YrtZOZuMB7qM+ZI3F5p4t2
3pwZbnCYGdmRT2ng3zLxYzPtFxpgA5FtzlsYRBWQ7ZIvJiA2trGkkuJQ68cyAnmBdAd37wUsD6qn
80gr3dUKUKzYnRaQVOZ5PNljXz7AX2PG5Vy7CpcTli4ZdRetBCNZtVNxKqfsFyBL7rivXq7wcVhu
llFxiCGDYmurQcvpFgsYGgXI+ssebZAesnb2rqPXUNb36HYeJxI0zs8PEN7gxa+Q3eEmyu2YBlxi
UPw/X2820ZEniziZAuSfF4wFLZY2sAjNqBJV/+2ysyfifu+zV7zWLupy7hDaJWuS8QG4tTZG/92P
RjzeXbX5P6vFxnzOLlKSO1lqwaFrt1WONQwuSrFsfkUQlk2zq9I9YJwkFpHKoSVb2AAQ0SNNgKJ4
KqL2wW/Rlfym85RdIj304523B4QagAaLVgBt4n1uUgr7JJwuv4QhrpNeUkAsdhnWqC9vlL+yfqZS
p4G2Ksgtrzr84dArZZUrJ+fG9NS+KklQMPsAqib58qWCbk/t6ElOG6J75He94xwUrjoa+ISmVxyt
nN/CApJ61xh74aLX92cM9SrKhNRvPJa7f9e9pp6erif/R4Vuw/cX6xJOvJyYl7epYwNKMQoCBv9E
s6UmcPShVzGi666y90xrnuPc8/rmFdGaq3HIvn8oyJF4T03JrF2CNJe407xO/1xA/N3MZ+pMmze/
oEIutPZjvGwENR2gFFGAUVfrzC+OT5I98g2wyRLyJZkngG4Ck/RoHmAOhBAJqgx7hICIMiYJ9sde
cVcTOE+uHSpzM9N/j1vEqtZKtfWpB+JO0WgYMM9PmGkEtOz3h0IPxvJZC+KjLJFWcEncXOczxxb8
aHWiWJtVAfBJmggoY2MvtRHTtQV5E6rQYA6IN4h2Qa1E/qsGdoGhIFreSddSv7CfrZrZzyPNE5Os
qIRauMMrU1iO1a6yO6+Jqj51vCuGLMH5J4/IgB/slB+oDmmgTzvV7y7LKgiq8Ibgc76OrmyW5uY+
yO6K5L10ieb/fGDG8Q/u7K4SDGLTCajLTIox27di/9Dc9Y+vJQEz2C++U8NWKrIgk5jHBXrWgK3t
f61FgbImmKo12scYq0luiB1hu58ehPUKtd109en1Hwqz7uytpdfWxzKFIHO0H2o6DjOtE3SEeCtg
Y0bjGqclNdztttK4c1lUiMB0KGog7UORPcZaJDpdXQmMy9XsEzRQm8me/ieNAWoJbBUEeO/7ssZV
R0SKZpxi0JcFxtOavssKYUBhJBAxXp8eNybaARcdqQoBYOoJSgi0yg9YAda0c3/iaCr4xkOT5RL7
XS9n30YfbAJmOjwpPIQdSQpHz/IzsuE9pD4RcYZ8KNBBRLQ/gQ9/nf6S6XRPTmziandUoRVruPPw
XajtCBn6p500xLi5Go7W0iy1NJIYuYcyjPPQK0h/ZIsah+fmNtyebl2Gd4fUMKto6cupjEmVUSP4
/DuyN/JQPuA+eZ9SEc28wul2dcqydi4qUtMimgVTkdS+MytmZkValkIe/SfbQ63g4oQ7wAAIJRdl
yBzO/Sli2jjmmiPsrD/f9fFloCj1Rd9nhqJfJnvSkyGUtqpFQwNPsokI+EymQMBEWqeu44H+HKY6
kaK6IzfCznM9541CuqkTAMk59KUJeFWAyEOlztlcJw5Ch7WXIBea9rZQJCC/71Qqoj2SGDCEei7K
LvJM1V4gjMZrjUk2AYlSIBDrDE3FNEfpDEZGRzj9fg9u2zCMXDSieGnGAT1fIWtR0LkCGKhRpeyR
r8eA9DEE6w3i2m7vyifbKFPID/xZupoEYc8VGTvsF7rsC7RR6SnX9ispH1uRMUWnejMw0eQlLiqv
sKIA7y8kh0DJRmzYqFrKyTlx65++hhgEwUYRyFbDsbnADVIQ8rAjiROE9X8XkLKOnix55vX30HF9
30QV5E8g9Xu5YT+x+NmDUei7d6UtaQG8nYw1DpGc0fPNXwMn9C3URBm5cgeqzq5z+QLElM/VK2R5
/0wSesnrXkJ5ub3gj5SmRf7g2bw0nl+xjBdFyV5PW+hDRMg/oohGg5pgwfkoG/qOV/F1D8qOMbuz
47R+1QE9VmR8Q/J1NlzOUmSaSfTqHz6HMnwPHhu8wrIvvppJDb8oNlxH8BB/l3Jh5d+bG9hXLGcm
H3Z5nGvGS1yIctD2cE5kJjIhaksb/iR/dLtuDn+sjaD/jrL0vCUfi5h0IadvCYBKT4Ne40UGbkRg
mQ4iC3v9WMOI9+EG6TkruSufqCul5IXfcB5/ySxSC2QaNOZN9cZqdqihIrP0q4XbIHFJlSzPtopm
o6jH++uhiQxsmxpYK2XH9B2EAcHHm5EYsqwSmaHSFrxO0ZS2uBb5xPsN9CVKcYIfCWyJmebVk2Lr
MeqCaOjGFaqa9GvYpFURPYmwgo3FE1gr+/92fK8kZAOnyTLT2nrxt3478ihGl/YsuKaSLwckvUd4
oqkvWy7Q0zeyRgjduwp9gxyVAWDL6/J5JKP0hnUaBwZkrBkynT6lMg9D7cf7xZ4yEfOqkxSaMd5c
mXGHRDAGDdwGAZbzVhYyk39zYfdQsHUCcXug61j5JtuOjTb8aH8chyYL0+obxKO205VHMtyIMNYb
elDc6JdEB4suop4KLtuY5fsuY0MUujyU7dLeZNLbRiFgi/qDZ8FlOcsOEkmb7zsE6VjCCe2uTmi3
WA38s8HnEQMtz3UTYpfPDGTudnjRe/KLs9ZOiwn2ymlV/JJsaXq4Lejj7B7YUQgF2w6F38cKbwsD
mEDBXju2pT6jr9zVpf98P/t/uSOBT0n2z3F+d1WhOC/PEN88/AJNtSKmCCIDvsADPuw6YvDlKB6L
ezSvJzW079xeeFTz1j2MJh5m/xsODzcSbsMZ7Rucr6W1BjbLowB5s23kZevPeOojtyOIzx+7Rl4J
Ya+ghWDWBLjEB0YW93atZKPAlNlbBm1ayC8ta5HOJklOO0xTrdYP8rcA/Vh8lN4y/nspeumdp26+
F5tV4kDwugazwhzjwoQlwPGslfj4QWASgjCLLkSebSNboC8i27JHWLIEeUq13cVrpKvHz/1Vwy3X
dYf63q4BgtCaahxMQtzIM9a0YOmDZK0PBdm6uk1Bm9mhMA7ufq30OaVXHawgyvemgGo2q5aDIF/H
iJ6p/HRfFD89LeuXDNvm3Kv3782rca4XPRmUlbDZOQKZkAMhvKP9pu0uDK9IhjJKGJ7Gk8DwkSLU
4VT/Qg6SdcQ8hSxgqOqwuz0ltql0pOJ+HW6C1qRaa8pCyJzXoSLpRd5gZOjJsAjS/zZ00JYRlzrf
u65bV1RWShYVTWKDJloh/O1xu+zBMTJ+7XpyNcqZTLHrDmN3pq+PIxUk1bFPGX8Akr5It4LTsCur
nCoEg4mNdT39liGJF0yi3xbYNltfL8dL0yG6PF+WrDR/t617mbSJIqG20Y5XIKD0iWGIMCs46CKP
Q//pUJs0hGoKHLyaHBEZFp+HHW3ao0dxtpDBY87McBomGMtW0OELzpBS06qOUmqKHH0RlI4iT5J9
4GDrBL0jUDt6ZR1WzRqLcX0XvPlYF4VMJTdDihBxkTLF/PiWie23R46L6FAUxFysABDBcrGr58gx
MOcqiblsjWtPQWYlWxsKoTG0tDwD99DH+UGXFxi4K9v6QTB6ApLZvPlyuJzXujRCrg8ET3zC0xCH
P3ZFqXnO2kRqP8VwmymDY4jxQZnoP3yw/HHY2XntGqZyqd9yWjsMExODgbkDTE9Ztt/NbIBI5YqD
z7KdJKQ6lsYexUvckEzRYrS3lnX1Fpr7R1HiJMUFN2fBOUEQr9vdaKLJUZixcWnlkQU+pSAQx2Sa
EjIoo23AIf+kw1XUq/ICjBackjxIsTzWXP1VnpgXUh0jgiR+SaRLKZ2PVSFKyJ/OfCVkmPdiWbYC
tjJBn8izrNrr59xIw9a1RdiEjz/LvlsfCQ6NrM0BMNf5FFwBakQ1eohSwz9YZVItWk9uA1svU3Le
km8Ktfp3NtIGKmz1qVyNsbDJL6TSHjMwio2Vhrds9fYqBUX0fhpEv8F9Rp7ZcmF5OaWvXHc/FbKa
Un99sZxB9dvL+TwpLR5+zmsNr3/m46XPybHi2BG0kU6kP0HOZ1YeP1+bd8Zk3U9ayHprYs5JBdjj
3OhUEI8ScVC4t0awLmx2Hd1bGMmOR1cAwMPilfU4xAohiD2bHjOTWkHT8ocJFa5Eq57BeN4wydAe
AsCXpc8R7q5XWC4+331y/vAou4ZVIGfD8kXxcKTJZ7RYiJEamKBVfrr1J812oZYUeeNqIS8Jr1iW
a1To3FqVEuCQdM0Ew8yl0qB5t8xbCw3Wh27kKIUk0OT2Wi9GmoXzVgqJeVqA3SjL1NhHpjZYWub/
b78jks8YyadxjenWQcr5DmiDVitKpyQwoMLAG+AUZI1I+71ZXOha+6KmaksnoPkxYtx/9PaQ4crr
cOCo3w5svnCyvGPlykBTDwe89ItDJBHo+FqZ46HO69a0QVkesJ4BbcS/y1aj/mdqjzHBHA8QE6z8
sazy6MgKUDwQpzpzp7tR0bK4j9z9d7V5oZ1FzfRvCAY/LXNyhOkirFH9b4hNevx1OHYMoFHnDbsH
p9AhT924TwM+B9K9OKdKqjUQ8u2rzsGFx8Nn5gEcyc1NoT3uMyBetpF2+iwNNWByjDCFY0uRqfCf
wv+rcwdlzaPPeI9Ie+p6peevuk9tyMuQ86f5uPkTCcCdIKagX3t5E7tBAdLAnHftzFHSFq/hljg4
o5ZVFD9k8sAiWn3C345JmbF5rQZcBGRaU572hhimqvoufOe7sOJJ7qxkRQMp8ArgbfT/oKoPRYM6
pF73GLb2eg/JgwksvJDQBGVj+nhQpK/ejtOsdG7OZzrbJTZbGsLSYkCePmeF5oaOksEf/Ep8TJ/K
twOrc3KtGqcSOp4ttgO829e2i6cFnAGv9sbcxkRyAjyiAqGz0IFY1eLQcFpMSAhk+L3gvHzNcrJJ
vJcuLaQ8Ws2mb/evVLHL5Twb6eCYo5OJp7UTzYjPS33TL7wWKiidUSAqo0v/lkbPu3BvBwdYiya0
uamhDUgtOVO+nHhEnYj132B4rW/gDc1e3WirOq4odhnAoHHEAZo8P46+bl4f5v9xQ7S2Il9VzJsf
WUeKSMSYFOI+CR6eifrI333RBntFiBHIRYOx9c0GoYVnYckIpxpnmI8xShcKvbb1vmnz01TdrP6S
vkT0SgRo9Hb6Gt5a6lBa91445Wh6Y49pCXsUBWhTdiaq3dHnO0z+srZtKi+bCcZb9jIPstYBdIh2
XZEd9M9AGiw+ZBMHq2cYUxSTI4HDnyq7MSMSzsofaglHjTnSC1ikcGh4sa+jYfD4DgcQX+Tn5ttK
hDIcCVb7NnNdgT6pU625bGmOxdI8Z1hsp788OLrkWrvFPh9y3bvx3em+vjwjiNmiKDbJv/Mdc7CP
EN3TyKNxKNJd1/g8PlEAKRDvIJNeZPFVWQk8jlIIX/CZcc46GQlXUFofjyyfUOVSQdYwyv+ShMj5
LE0kAkdbYgJWIJR8xGyDqJKQz7WKvUXYLZw36Da8ajzxyOVYOdtYU3GFha0DOtu2EuzZbcBVp0Gf
oKf9vYMwhGCuzkChXyYbK7P2zh7H9zw9YlDGUVn/eX6s79qkHMMgIDe6p+BSaaCzeFCuaISl32UW
TcI+wjs+CPZPY9Oi4jEKkmAyRKtxxdzZ3POdUM1+XL0N5ikgsoFLhbLQMb7bhzwG8YL3/XHD9LAO
ooVlcVkTyhFrpaA2SinonpyskzUgQR64jx3WY4QHudzHkQvNLyJ4khV86y+PuRB6Y/XW5lX5P328
PIJnvfDX+OST9QLfreHhCb0NF9KJ4JiGc4XgceJWTbfJbDACZ3CD+4TwD57KSc/u03C+zIfkvPaw
LhnJ1EhX3KF1id9+vpXa+n7CIMF0kYk381fSarPTZXuikZtZnm3DPaALageYRXvkQPzSWQl428cl
aW+wSiiAKIq0hcA8tz+yhKcmIjaGVQ87ADcrBN6ZuRdRnzxdlwdRRmxvxfJ2NNTDQWrH+9UbOFkC
igoy70m8VMCOlKjRbPztKWBMe1CeR7bKZ0r89WgEkQwLFnIaR4QruqpFM7dxxc97h7u6FUxA38Rc
ZExi1CKv5U9EGgshuOpZYP2PB80mNZTggO4644P1ZOJ6sEwWXxi+hD9zGSAOJStRB2rvpVuN9Ley
vOVd7MHf1ynHroan0BVu4rGKyPlKo27VwqMmr8nrPxhCHxQuzcbCAFBb0bsuTBcpBok7bdQMBxpP
2feq1jajCSRX5YdJlk5rQnHC94rKJ76qSX1sYrhn8n4H8LaPBXQ/cpm3vcKW/eUiTsHRU2BZw5zR
AToq3SX1RFlK+QeCjBRVI74ijVzm6txRKyxiRLb5b4l777ULpw6SjLZmOwmA2nO3p3uo3S/xhZuz
KcNXxWVLpBjUmWGb1fjn48pryVkHb9RCJSoV8gZw6NBWIy+QJXr5pTOLyS2S3q5723nicstJPR3I
Puv46lUHl9FZ9v0aWCaw9IKw2zCxUWM0LbdXy9GzFSfdXFUGe8gY8GNeo0hAI0Zg34wFK4VrYb6q
u8N174ldPSoO6YPf2uEFcX6gNpcQD1vOkY5z2aUFhWtG9hduU+ANXWh8O9zsvEUllkGwIzeatW/G
o1UKB8MqL2vErEzToE0tzq6IYUF78KUo22G7j6f9xSpIiSx5PP8G4BsC05gX7HLekTvJOi1DM9yD
uofPJgCxQ9ijwTkT1OUs9s7iqFOowOLByNL9onIv+fEp8MHg/AxtLIE9G8QJ+ISUU4Nv0GM1JY3u
LftcJYZrMEwbx2myI+Av5v9uINvv2UHfHSMH0QPBJzLSjYaE7/6V+I8i2biIPajDNPl6T8PWSWTG
bMsxxQaXc3PL5E1hpWWuAGGNe/zbajWPmYlJ3qNMJ+I8eLczBk28N8I205Zm9LTN39m6yZs8Szpg
oQbn7z6Hi9SQjaNshC2sKwP1N6XkDe3/8PIg3YXp8zlhxfCVHei+kT4Q6Gi2ntrPnwbW8+73Pqk9
9YFeT0FCDyF8dRhVh5hVl8lhPeGZNRlCRx0hUmsT+lXQthWLqoTJl+MXcCQv7ae94poxgrl92l4m
7+rEG0RryzpWPM6l5z1vLwwOTrbwbCg40b3JPUENZZrAgbQs+cnKVZhwNWJCneSnOh2hsWOdppBM
SqiOcGdYHJ+y7QRvJuYAFkbP8f34t/jVDkyVLFvJjgrsxUOaE84+GFk5sGpBGtNKq9l5R22n1ocX
KE8u7lBFJ9DPpHMPzCLbEp7LQ+bfRh0CDdhRBKE90B6/JGJyg3Wnwor9lXqh9zeyAuciLYwvGUEW
dsrIYUwPFd+MLHIvr6U9cgNSD95Xtf4a7YcDIFcBdkk0B8cshpgEuc2oqm7hAg4Whx9gBP4sm7Qt
VfnDJRu7O0wRi8wDb/U5kaUXxc6WSqTzUl31SpnUlMuwdJ5UnqGe4QrEMjDRxxuI8ZJnuIDJ4Y78
hM58EY9eEovadsHWuIjGhLCmY9QB6w8/sTBnpD6HA8EAp7wrO+7cgsWpVmK7zK0HTrFmFLqBV16T
bifAkH8gSH2PWR6KdUghlGs2KIhLbdmhS4dE5We2j9GPQXR+Xa0UNKKAY5xzXKxpB9qV4Uu//HeS
9gXjT0Be7rJjNLNC7jfLra46GJDFpvQotSrphgA1M8NoXONP3nO2vNp9MH6hNo+YltMboETTAerC
S1HW1Af94Dl0dBoVm2Aw3zFwS3j40OkFIt932K7BoXo/ijFOfPPbQSMHz0pLv59QQNFUq2vXTPTi
zFA/FRUBla3WDAJAjCFLuuBOegKW1WW9PpY9LcqdcPoGeQZkUXBfe01X26bcHgsLb67tAKuAEZiR
hXimroaEggEHDsqaLNPmn+MUpL4bDrFzSd1xBfaLxWc51MuyNyDeLpNwuq++DM4vg/7rVtRPZvHX
akaHHTIx1vKSDk7Pajjaa36Z5otZem1ZVFeQCh+TAEfJeLva5GBK2On+sRofl1rXOuDIFfVmPcrg
JhmPofYci8Kxv6fWaf2Pns4Z4j1jBVXqXVubBycNpQTjuXRt23ZLxdgWI8xRMxWRzS8v/JKCPZti
kef0niMecmv/RdycL1bP5BhPZIArBmx/qbSwQDPQrjJ18ruhDlt5bzYaga3oHPSct8IX02euOtz+
Ev1RLoNkhvN/Onxv3E3UCEJ5dRHp9gDGoDzousooLxTrHoZb+BcXJRhfuxg8JU25sqVMLvGqBUTx
EFU5KeGagN/09ZE8CF1zHHRY+b1tpAEOR1aKfxB9aNWrJhHjwyiAil9GNgWU/+g8cCuDbjKRCkDE
0BP8dF1YRs3iBuc+SbKy2j18N5J3/H2/fHnGPcYxv3w9XqT5jOTHMGCoiypw2TYzW1i9q8j8KDyA
Q5tcD9ylzu3MRmmZvcAo3tEULpRHyo9FKUPtvXOC7wgCghVy8bmhy8+6lAbhLH5ovREmCzcXmy1R
fmSzfsfDxsjBjIKfcsDYMejUCdiJxm5hF7kgLCwO5asdVEyFQUDCv5exeVgBNxJohIa8R8tCz94H
XtRTADaH65kH7cGJUwSg1l89C/tkZittwHWTGhT/e7eSqm3YpbYwEanre8LeCNvryiNtMrZHaePu
EV9zZ076R68EpQaaCL+xGXCZfbRLCnpL0bNIoMYpL6PCUFGi9+e0Kg3m7uA5RM/Z1iSLKxjd2rGi
bNKucy8nYC9V68f4WS7CVNLgHS0ULRvq3bsfrxgImo+VNHt5cJbrQ8NhLfBToZFcz7B+sSEs/3Pg
URjNtIJurTax/EnbZJ4sqPSjpo8bPbPKDIhHuxv9EvBqmuKhGtuf3PLBIPe/qnj78UnzISfdPO2j
z1Uy7uUN2omaF0vrXtaVxgU1vYTkSLRn1aIAIDu5Od2LLQbWxUNh3smeT/fhOWb50504O22jk8es
CPEwg73gkup0aUd/fSyDuk0y1cST/r3kD8vtyT/q/nIl8ybH8/yec8VTHv6b7fdK8Q3ifwPh/gDs
l4+UT70s+vmP2OANHhyEE8NOR2rX0ki5Jrq0QsIMjowq8cJBBM2VRix1jfrEuz0CbqT26fFWc2wf
2KdP3fwJuRcqVEVq/RTaQUyP23jgCpD/d+LRSZS7dLbvEohp7bP13vriNnC63keO083HuHZvvul+
fZbrARvnL2U6HVB0iQnu7glrkROzSn9HX/YQUk6agiqPqFDj7cDlrfQ3yxEwt+XzTWRR9TogekkQ
wcriBms3Cz++3+o2AWzei9WWwQYmqfKwiOdSx0tg7iRec3AYsYiVEGmSpRaXZm7XA9WrqMxRmLl9
5lpNJY0zLGQHGJOKeKf8AYCMg+HmMewgnmon2nRxpRdeNjD7gAfcmDqiaA6rKXCQHyGc7bBmVKV0
d5n20Z64v3H4mpQ3mCwmeFk0wxl/cdkqgUshbpnXQ8CwNZAEhrVJZeq7ifEFz0ZJ/od2cV6cuhF8
dGuGJ7mzkWQzLUwqTe6l8non1wBxq33a3scKsZqhuAnoLQGUXITFp5IJuV+Xg2CajpiYd4YT40fO
E7NvdF2BCSgqmMEB/9EPI/xp4VJZZZs8Hul6pcPtPT+FR4F0GjSeGn8DXK3UrG9ibkmnhIO+8Oil
egFr/2GCxNTYFFtaP1bWBwsT4izfQT3E3NwJFTVz1osIlGzMZ0e9KPPGURP1Ttufme5Fes7d2aP5
Tk/pZJ7XPjx0atbx4iA1WJRWlTnha2ZvkFX4qTA0cfEOaXhAYI8WtA2n+obMhZioMWgyDvapoYeJ
US8D7gOy60RdtotmgsltRPCPB8XszPLXXNidZhWbwii8k2v+26XZHWAVlI8zfCOBnaeHMuPHoQsr
T5Y4jALiLAZxiRdXATeLHo6mzMFemJ922XMWo/5MJx+jpjUIuEBgMNXh/BuY4jbsw7liLc/cbXAq
QUU4vNZlqE/Zw0StvABltIEOX7hsKGe23rAJrKxO37/1MimZ/l0uPr3rwltWrHivbwo6Rbs/EAaq
CP2UY3UUgWt+/l6T4DbXLiOSEGmGWfzekUbJy6pHR2U3lWGWQRQZktg/Nxq6jdUeyPxPcm6KGhAk
ZHlBvkrq5Oa6CtRxMoAANUozTCjtiO7WUhbZT8qQ9XBAs4v941EP/RLEzHKX263BLAqrAtTpDcOo
rjrI5+J1w9JQvc11tPjTESzSEu3eXNeSKH6fu4iIA+j7wYCoEZ6ZRfleyGpYTZiq6qUfglDqSkrr
73Jt+2+YdORzdLz5KU/LI9TomaMl74tv8xd09nFXCkMrfLIZTuDQWmOAvVh7zDxeJMlyzP/vEW7q
pzh73m17xD2LlRxeqSbfbBEaDuPHaSwztljyHLU7PCf8GdvN30XL1rz7x9dPOWiDexMA6I8JbZsu
pqVhB7dDJt3Uwe1IbQ72WUJ8MZlxbiWgxZFbI220PSjcKUrrfCyP/610AlbsiTHtlINmJ14MomKJ
Protj9amGDVtb3jqnkC6xFdROeOk9yWrinu5yFrXguwPOUpfX0/8dxN3qbaK3osz1L1fKL9dDpqI
1JMdtV3yidUBEyMXsSi8HGdaRkufOaL2+xRlVoWsOhXrCdULsD5DUYd3ayGjqq11iZgp1KXxvZvG
9Kt+EiRwus2CGMwkcPN6VbJ5eEtyAGf5m8QR1NBOOSb5wu8H4rfSFZ7fyLMIQLgV3u+QPCsmuGoX
UaOCoAjqV6wWAG0N07x90RjytjV33AVhAew+8KbqOQZKlnjmSvg5/d4GmKkKZrKRT81ZpFpNfIt5
RgfMQUVflXmMu9uwMRNJC1dtLZ27IwI6PqtuUGXq4vPEccW661zUs/4/VhOwEXwpnV1ilK3fHaMU
kMBfNXjR3ARQfYKjAjlJkNCxVGkwdZHTHuCf2TgLS2DCrUaVEn7VqoiTMPWG0z5U87RbHHm12EK5
M0y1X96F2+q/uRFW60KgNj4nVI6HndAa7YtaPGL/RHIWOmzy01sCkb4tUtulNkvRlyodmzI8bs5h
xRAalaTcTEMKoAiP44l4YA9YrkTq0+yu1VbZ9MPVfWfNF+MqfsB8KjgsrCpzmCwLtDUL7jS6zNCr
lAFL7/Qxo2CH+ISElod3H0EibfTZeuSJPQ341ygjIYBmb3hia9+JFcxYa2FccFhXxG8k1/vENG/w
mZYGbKNDEsiLal7uyuUpguh0z9kGlUdhlD7UVjo/oNIKPn+TaESAf0kOA1Rznunj6hFkxr/GBXVD
9ARnRTk+Rc6R3NmvDiv4MJPZ7anG3/ek9Vf6oOIgtaNGnExJ4DBTl7L2KQgMOPZiItonc27Ac4Yx
2q9PoU28FyZsgkm7IRwaWzi3QCjGw2TeZ4bfI0xhSvxhZaaeKeLOCBbACfCHKyuQjjETy3deMDKO
UGS0zZVoh3aqabqfuXwUXl4frPNn1tllp7s1yRl7f2sFcRiINdsQU4dO9lhIdUkANyP0QHXALd7L
bYxGVVGsDYUzLoCLKNw9HrEZAbPj+6Rdp7ZVSVwoshSR56dlbhoJTJ+dkVbMRcLpO8iMmTfpPtY6
CbduFTSt0ERMAZMzo0JlntQaMIU7NMfE+Xsb1ExzS2Dqdy30n5ETgFZP1/cKhSdPEbXwbFcg4Eh9
9g8E4V7p2PXlozOIW1oVhXmUaVjzI+wLWjR0xmc6PTXqUqPJ8u61/uFxtC71ouB3MdqXRwf2mksv
t6HN2ef753oIimobyhgLbcPFlXsYxljV2/59kJHTh+LVOc+sCElsCrGkR1RAzHWIqZA+gCKrW35v
bDGhvLTZ1G3Iy1up+WA0B9ODa377enSXvb4zS1dI+TA67EGl6rfep4zXA3888u4+0KbLCW+MJ1Tx
q+di3214YF6J6kFZYD+UQJzgeJeoAM8rwSKfkU6PNC/lFeoMriebkNMQ5/HJV1GJLrlnElj0M0LS
RyKCSu6Vc0sgws1mU4gjDw4fB5emixa5B2tVkr7TaN7Tyf+0BvVoWngm03SohVISOHDIoPyvfAZd
tffJH2wh8952wiysI4ULYbu5vbvZ6MJggkXhiSqGK4RZXnRUZi9oRoel82W/tt3lzKcIEzdbv0fD
rEavvAZ4vw/mE8sq2fnv9orL8nTYbu7VQM+dz7X34uh9AyjE9X0WYV+iE+yXpnS8JGUwpNTCTFiP
w8/2yJdzpJ2MjB81wXxQVJdQZbyaTmPyETXkgAZTfju814zhDhmk4wSQPd3mvD2GW1Wv3CB4ZxNH
+DeV0gCzSBPzRQ+Z1ApC8o3Vzj+zmlbkq3HUmoqPsy0OnVnQXLrp9K24KQ3CZ6NZFTpnxkwF5Yyj
aTHAb8yXUagDokCgjobeneClP0w/Rdebo+vaI1bUq0afRDzVeJW5IcrAMCGYAHRmp1lcQ4rmH+eX
qXJYOxnGm6ydJjBmVf0Bsv68FwbG/VvcXZvrT2wbD60Ch/1VnEoEvKHYkB1FFH35noPqivPZFXP1
NJmIn/M8DRTue68p/dh8ie+bsawirR9FEhrNk4YYNEJwEIF1hRQp6nJ+q1Row390O0MpcOdUxoYL
4UK13ymRI/TeeDdV+srq77dEH9E1lAH0mhj53h1r6xlbSt+0T48tIasJ58/m393lDIT5dV+ReAgM
SNV3MKELhaV3yBJ5hY3HrIx1/PtlvZ7Vc7OT2Qqe1JleHbL/DiH5MeU9H1MHgOMkm0fy+ImO2I8R
kb2nU6BsTvS5qpL2ZgqrdB6pKdR2RqNbKiOHWnLR76bL/VwsmGAbgPKoaCAElyJ7UsqSCB2DY/aa
Cneo3CzBa4wss2y81A2mp5/ZZpbNO8YokrdqWeEST9HQfAlm6v0BtvmuLDnx2WL0mnOtNV3PmyKs
DacRwCSf/UEAkbw+vQ3YcySavLpO2trBHdOfTXXpdC8VqIGLiRE7FOxrZpUXNfFksBmV43R2CT+y
HGK2itG4v+GAzB97JvdRczKvtvqa+QTSfJ03DwfyccntbWRGxb+jJS5mMD+dHP4mdk/jgsapQDkE
Hsp+XY6wlecL2XYlaTm4/q7LTmFSDe+eMiQbqip2ZnXwa06ZHHhvOyYNF3+SjiNBayYIsuoujS7T
BDCtvFu7TgulX+1V1PH3WlEnHgd7aaoHTARSA45iy1QTA0X1pj5b97jcFZ0OxRbt6ElJECLGHlKP
q6TJ1sfHiyWquWN3O+6ss01OoN7CJJwMnctf9qxwcUrq+E9uievAzVtfga6AVlPeahTiifQn6aPG
qNYQ+6Qv9yvQfgr5cQETV36P0bSR5g4bhMKQbI8rtEVZ/zCJ6aQdYYglANNYzV3X6Z0Nd70Qjlco
QkkaaA7eNGzkVfBPn5sun7qYYAPLZD+5Cs7Pj3L0DroBrhwC/oqLu7y5OrnXnt2996C5/cr8Nr7f
ofg/vV93N4JmBj5PU5TfpQbn/Je8YgTYe1AtdiZm4rMmGFBLH1DwcGm7MXkDL7RAd57NpzDrJYFS
hcI4TofOLb5wqbRDHj3+w0M0T3FXSEXmnWU9fIATTnFolf1s90bjn1+75y+CAB6yaN2tLz4LsXH0
cGR7V2HApCvf8K4q57ne7/HJvfIBHSvNeVXrmX+KpkE2kY4ymN+UEy+6jNZBOBj4Vkck5EGbHEqY
HemlmwpN0XslQatG18IV0pOC7+dekWbxtbJEXNwUGhC4LrOVACVJNU2rjv0/eWFojqB+xaiH6R/h
kpKB1XiV9weRwRNbQRPXP6UCbqs/a3OClWmzNNEUI4qaXSEyDU0ZSsNtWTOeFjp4H7pOEU+vUBKj
pFbOKQUTJFabCDXvlJfQKIVBEBj8NM1lmGFQOHJTL33phBd/+y1lhIcQpPXGuZJnN/ouYeaf9j5M
6491BVX9Sfjl4UAN4jN7pU2zLixOgadVbhnKyxAfGJnPwrCWNzEH24qTolfmEHWJzYkOtE1W9AU7
+EpLGJ74YbzRXSbAaTK0go2eXIT+EEfUqTz95VfBFqRWNUqEAmlz2u2T8FBJxteu7iCRD5B2DPSL
wqCiYKIJbNv6t0MUiuLyFs2yDUFmvVxLUU10QNI9txcJvAGXQSKp2TYwLM/ij4j8GLxyhYinHtSx
YV+1QDCPSGPazuld/h5u3v/2FONazHKKW1ZyFpjta7cIMViLsje2UnvD5JfE/ERfasKBpAi1ErTs
OmVD+VDwFGmc7kUYe3FSbEGDzrMxADVpDsCcloRBXxXdOkx2UdMXjZ1u/lmV6NZJz2gy4s8D25MO
qiFLVFJ8qRL+vvketDthtorRvxr2YqtSccZqB/hrhffLnZ9EOCWswN9fot275W2jYKe3SHd+QKlk
r1w/sbecRk1pgaUEy9FCNgyFhh4nDpyrSuWGJaupnDrWGwv/jsne0AO0OmXDhUt5nBSGM3hFnNRB
gTJVH/v4v1JsN7JitYBbb8LIidy6z4XOIHpDnL7ci7jBohlnNqQQRs4TYgx0osEO5y0eC0yzr0zY
/bC7SVR8rEb3SNblHLz6GyzMmSrYQ84xSEjAqmkPq+256tpIPMXIR519cAeoguLR8ymJHxJt3UIP
+iQggDxB7zd6Ga6MUsHh9hUSNYNRqU/mN3045+qu0OP/E1L2yFCbM0dDJpQnNQJKophKMfp/ajHQ
C9eecWzpDWycx3ZXC38Xm7ws0/l36kA/FCNdZeBcOp6H9RqAbMfbHOuPJ3qReF6yDK6lwNkjc7g1
oho9HMBRdwnZ/2lGWckK14j5sQTtLES1R+z9sgDWV8QRfNNde0HA8a94CoHAtsFesG3lUfaorym9
fpG+pMspM5splmaCi6FfmPubtKKGG3XROUGjzPIelxG9g8IfpSWoszEUla7Hc3eGSyQoct3+TsPd
w+HZRgf6ztAUMD3hN1XSJgJ5/oBdYc/FeuDGPy5mzkmG3jAPdSS3ArPFFIvD1NBcKK13PpA6wYOU
HZIDRfK8f+9A7W18jtnl1mpP+0Wnf9LMyz7xExKAcePmjDfdluQUsLDDDQEanTCly8xNeSInUy/i
PTXOO2q6mcx01LTp1XNncSQNKzz17+/SRmF3wHmCteBZIk6zeHMhT7CxHcaCfZQoLW/DKkqihWML
2ahSMW3FwY+7V0yF5FSJHGsZgiam+8pIV47holu+bDgjGNpbuL/V5TVnDbFSBEvhG/tKOvaYUI2K
jeEP1/I0sz9QlKqJd5or2oAwSEbkfZOmEP7aTxvgrLFBx83L3GwXm0Nl+sOe0j0ajadpROYllieK
0JxCYXIYGqrDhWdWr11EOzmoL2a8ypUCnAPtf7TE94rh+99t1WsqXKc9HuXufJOXNOmsYzAKs54/
86bI6hVNKscUHiQdLRpqVjzJlcri93UYYGFA1yoSD9VVJaitBAj7xPqmFfMViBmoiCcrARNBIvjx
lV+mH+fZLCQWruJnnCSl43i2j/xoKvq+1hB5yQGOiFyNSej+NvvVBrPI5RqmGx0Z2Hq2WhIuUgeJ
HjIu/4Kl/6P160lUCsWuagAz3NvTCMhjFa9QVaIHdbd7aqn11lS0MLb1tN+85k9kSi2SUM8BowUJ
0fEVFGz9o+TVC6cyqT8D8yQZtt/ZgG3aetMxDTEJnZ2WayWjwcmdA/3Ls3NhS15yXBw/V0RIHKRp
IsohURtLVqcVsLXc5/Yd0IhOZMl843vTxxvHk3QBKDXFY5X6fGj9gaoK5Z/nAQ4ZCCDVK72wv0O5
K/WFM4itZkUhaA1Su24yyNrxQ+fousfxMyWlmTNlCNcd6WWW+C91GP1VgUW5Ye2BiUZzSBy6kWsO
ND9MYL8yZsQHoXWWyGdENCNhEbLEh/idVTWX/pprerEI3nIZkjMOUvj5ZmARe0AA1Mev7JkKrXv5
3qvkAj800sk/Nn9ZqD2ljVnNrvLs7OuAle2Bjzl9Lmcd4S9GaXvUYVjYcsUx6OQI6pyTCFEspTFQ
KVhFuTtvuAdatphIDdO5ULesSDyYFe7kEFWZUvVnfNg9XS010JleYdHzbTU0ltZJrC89F2uS7FWG
lI2puGJNclFNFKtdw/sI7F327XTuD0LVVDYdp+wglhEDXvjvnzMJ0Y1UaEjoHJ/nI8hgnHHHX6v7
HZnDh5WNyDHE9S0kcJ0ma/rMO51wto40ivsolfMGS7LU3Ua49mcWBdZgtf1tfwQyyZiCbXmoA/8c
TZtOhL/VAgPRwTr0mIcy70tMoEFVv+qWkBamZM9JVP0Q9xmFccSsOr8rGlDZ8Gs++XHz/3HVrnrs
n+KXrfRwVGpx6UE4BQ4uEBODvQG0LZq/edo8btsVID/BbTWC2aqiqA7HMrGxQnVc+OKLnpaZG+/H
KQERHUEzIzBPLggesk+PdQ7o/wPNS/4razYR42eAOFM29bT5E+j/nJ1Glj81fg6zc1lWkMngJ/ZM
cAP8KWYYJvym4bFqL7Nyzu88u58RYsWHv9mkumJy7RM+c9oex3CdVQrbBFF4yA4YqlIBwE1BLvjh
pnaHMdNEnZgIs+Y6u56+AjEr25ensv8xRITjwkTPP/T5kXgxERunn6G6K2+qSTZip6G44ZLyY0Xu
IPcYm996hF3eJ384jbCa8Ps/GE12af/lmHEQmi3PwpkPawkOEK9WbpQ2vPYHDwBprW0W3p9VksxT
uUDo9V9ANEcMomMNNQSn3mK9d1QFfkVp1Byi3eUjk46jpU6x6ENAv1B4tmPTpN9O6Xi7z60iVZk2
k2Cpm30nhYO/E3flY3yBuMwjCbqVZiTKOvsSJDFpPEvGfdoF/haiO8RT3ymyiDGcGpwX5o+82tMD
+wwSuoDhj6dBq1Kp+SwGqAPpWhnJw6TBK+/BRhEMTI1P/xY8BbYpDI9ZX5kVrMYvcFM4JVjCB38G
4PnNpPDfPg+6hFRphIFfx+qwjn2uYxQsTokJsv6iQk6ZdKrTthdxKJDunjUVOP41CBPjmQvcRLnW
TaLeFHLFW8HPjrPT4p/u8yFnwB1bjYnIABIck74e0suTghuOfWDDSACgPIiaS9H+FnrcZTIKR24u
DjYc9Hhrbj9z70v+/11oX44wLVpxZIHdoQAxq9BVepyy2o7/1oVLuGymA6U5V7XFcm5YfKQM/vf0
6onzk4y0ojrA9LqiJnkaSjAKEpn8o8Fa7y6Pw+uaG2DZsCseMGpHmrCMZAPIEFT7z54vdoIT4WEp
58wPeUxF7zdE0Hwla0+NWPE41ewm5rklIgma/8TTNly/xn82qg4kDJG2CO2jqDWkK1WFdyGTjzfm
HFxrrHlyeO0rVGvnRaUlb4zmruTbyQrM4CE6aZDk8PTuCk4j27Rqo/bCeVaZ0bWQn1UFwj5Mhg9Q
oddIv+SN5lrJPdc/gO526hq4urO+N87/1ixsUwpuUmTXUVJTlnTUMFeQ1BlIHh1wx5M+vBpfmTzW
mfCgZesiyCz+TzTIMnEzNCgy0hNQz9H1utT2R37Khy7iAwSy+lfwfl3QHRv7iSgVsma0ulGj41a6
UIazBd/IP2tlG3ZQVmhr2OaYgx60LyqqHCZl759NMV/SBWwf/w2v7sYNcS9uke0CB3XqxkZeR3ze
7hx6uhN+ZQAVKHuUxiV38CUZGunBMKnJlnMyMsfrk3WvXkZVCfM3KDF0v2CW+3TZulJsFMrOYjza
JzPnCamQSJABqZ8ZaZLev9IJUogFC3DjrtHCVbXMVu0NL0Xr5aC5ov0yqFulhFsgM08DpxdnYSue
wEAxCI/ruvzP/Cc+9Z102KG6Y3I8ZV/hPYcWqkiyyvitObW/FjC5T1zZ/q2Y4m91noGey8Yp/Ub6
Nzl3qSisJsT/St7/QJZWT8n7OdIMoH3r5WCnlnSupS6rccuvu19e9iY95GxSKLfE8xLjJgNrC4Wf
0Ec/OXzdkceSRqnFy/HV70nOaSVZcAG/h51/l9mQ38nPJtAKnsAM8XAyqLMtJslcFSYttSs98jvS
sZKNKKqbrm+XJRfYEXSDAXKSPAVgIvNxstIuT1pgaJ3wcLqEg77xslEg50QcVv95gSoloVsxQLVz
BiANG+Wu5T9Q3IL/G6rCwmyiPL+sJspbpn7HaE5urCWmtwVRw0oJ9f3zcbPMPZjpyowUD8pqUBz4
7778Rimqwq44I9X1hgsuH2AI1MJ1gujhiaX7N0pKy3caTQLoBCUlq1qIEthxtzDrbnlW8gv9H6Jk
4IEEbINYILCaNxQbPC2hxGRuJDHeeBAqpwdM/wU/2JI6MxfCH6T2sdJGgyJKJ0q3N+FtGWRR3ZdM
sSMqLpUdVLERLhVvyVgMZkTy7TZxmsplddZnqabvmPBj5pGvEN4rZNg+H5RiiC417JiDb7DvQf4r
sYFFou8qj9aUYvs4jsTuNoMo+kTe8Gf9J3oI6in5ABqxMx6I7mG3uqOSCgSKJOAUBd5hrv+VG+01
jFtQY3jwdQFoj/8FfCPdooBdMfphTOmKtP6cXjaNhwG6B2FoWwFuRoCJ87vJOUtXRnox2rEABx1k
awdbtZgQfzoBRdg8Bz7kQFdLwHFgJY/h+rVT8gHnfReRTj9AEq9OQ8HESj9/BSPST73/ttt6iIbB
fAHMg1MVbxPHnyLN/v7TTMumh5jAI+SMzEUOPiuWgOas8f8KJMs/ry/zjF5EStSE06dt9WS/BPwD
uJQTc2zRQtIw2p3iW12+wUCl8Al6FkC31MtYS38b5/ILJufj0ZWGdWBmBlNmGUvVXbaCnZCsom3y
lniIiHlZ2cnwt6KvDNSlEC6OM0J5gDxN3rMgEDMUq2PqmPYrUEbUeADXxBykuWuKcqRMUCS3jcVV
hCmv9VNuGgqO3xJarXCRY7KVe7fVci29SXK/9ogNoXQR8KHAo3OPbPGqfmGjOnQ6zIs0gSj0jo7D
yZRnEIhXdU/qy6/4RNdQy24wYkhuZwtzV6454q/qktYOfc/Onjp3sUZloqvNDI4lhUJNn7Yq3Nes
+w8GZWzHWo+GgMhjk7VSuPswGhc4SDE7mlTwae4oNwN1nrSTTLbTBzw/oRXWb2Zf8b9iaagVA4Uo
0O3N+ZPIbxBmDoiu0eJiv1fXdo4FCaa9bprZFEU9gP72D1zpq3ML8J7uK8lDkn93wF7n30QKIhJQ
4vfjEulEs9FTZEg185XCqACrlIKPac4qpCbJFSDKKZlsSkQKkzrzI4bS4xqPLh9DBKxUr16xS8qc
rwZnIcsstAQ/OuPnmsEqc9ypVXrrLTWht0glmCN+kMqX38TdNz79Cp4OOjkjgKXjyDSz6Gl1LYzU
lRoEgjXr15RD7FDsAvmQrMw86w+dtjmq2gD9tMYoP4POvlgjI1BS2G2jdN8wv/u0LSJ++juyNzQ9
4aMYMKvYvZ1TMBDRiJobxaT66RgmUww+34Pc8Qx3DcVTfh2/dG8lGxBZPq7gM7TYUOiGVs55S4DX
qyD1abMpayzkABkWKGukA/whEMLJV9fFdgHkeS+bGJ/p5bfDVdBY75VtGPR/KAEklxZAHEPuxtIL
bEOkq2SDBhmiiFg4Vo3OpMoMOjsR3j1B8s0uMatRq+aK9g+RkLjWGGPOHwe26O75InCrDXhsmpGh
mYHEg8Lo8EI2TRC38/Xez8vsnC4mIfo604Hb+4b85Vaf5P04aFh2yq5obKPlDnA7w4hBJXlMRV3g
mqtgZ7ng9/DJwyhZJ9Eal3kWJyvCA1U3iMBjV9Duay7zVnjwidQmbWLuxsz/ltBuScFi+v3YIoAG
zzeec6bTBwZL8B8njWubIuDfIg7j3e81kpxdaDpRQNyqHBKQQEchJO4FZaj1O16rXOUwDbOGAUJc
mJQkKzxe7at2jNUXnVYoWEKrL04oeGXljg7+VjfG5YRNbJ2qelEm6leJ5RUxnMWKy+XqFSc2J/v3
W5hz/tY7Ult7CzLLbSTWYaouQYSqfk6qzyip/LssA/2OwZ2WxEk+g6GRoEo/ZO6vmP3d9GXP1NuQ
4WCcj0EqoipVv3/HVtFGDeukEzrmDtL4XZDlg1FkmoeB2qv72nqdO7qxIdMQhJZElPmU3iGk5Ewo
VPfIjUs49cLLGeTBp+7EMJLDAvwFcofl5STK3zR67uit8gvDSHMV/1IsJgU4EkOZH1O1kLhmVCaz
TIprswiHM01Rxev7xrMRDNK40FXWfQM1QJ7eg7n9imi3fCtIL4YNSnFHG/M7Tx+bafKB9SbeWNi+
JHUQ2gL3LAeOXrGiQTeIdOK9uNrilbR1T3GSJiuDbqDjbH2y0jHBIeYRR31Bh+Cbf4XgFTS6lX1O
fXKSRzj0AYnd0gI8nx0PH0/uHz/9uj6QNg5mK86JFTVhx/cnAevA3InCVbVj9YDIqYUqnqJRBptH
gz6e0zTu3k1cHSbWip2iteKen96HIaUMI8/4hdnRxNRDDgyIPBpR0SUjcL3Iy00qSAJVHZHAn08o
PvYFdmfhkNn5W4dLOQZ5Srk1BSdRdMHfrdxoY7n2/ESZmHFGZHLpm0kDJXa/jWfyTRfRcPNT0cKS
pmRe77JiKtGz8mO3SrLTAb7GqQpXyFZuZ/Q/Eo5gwrBf8Yh3MiUCz5rV4g1eAk7uzzewC8j9oYWV
v+TcbcUKJkjL58PwEB+Z2ZmefFEYlZgMmfeQ/bSx1KB3TITnGmTa2Ly77Yi7/kPGNwnbyONj1H/6
VOaUl9TpWSQCSjBrLX558JGIG1SMiTFuTb6Q7szXKuv9wMWzRGJJ/EgUw782Ue2oKIQHRipG+0yn
OjBBoTWhPoK//iRnP95MjCjWD63anZtJ64qLO4XdFI8xLPDWRhTbkxOj42ze7e3DBEeJZ+KfVYx1
vjaIJzBzCnavlMIXTUD9HmNN4tWiiDjx3mVV0De5NcfOpJVRFDTG1W/SYzfV/QI61L6ejINKbBTL
vbMD9+6Kg451XX6BzDqHJroagnyJUulOkK/em6iEovP3zxyfjODiiQTCf7yLhYPHzv0Piw3izFMj
XYEkBXUs0DI9MpbMjHC8QKM9y6k1FG7hTLHzc3S6lKsF+5wr1zbm0gyBq2zZs308VBTGxVUrVMLH
IBu/DyrnrXxXSfhn/cSID3aF5VniO0iF48I6doSPYbtKh/bD7IqoYAv8Ztr41CXbR1aWQsEdHHIT
FgntLmnN3jRXZ0y3r88MW/QqfHDsT2g5K3VJ9OzAYf5waZpYaZsoXGuh4zZgzdy3Xau6dgmvcid3
TPYUTJXmfvz0YGyPJujV44FOSJ3x1Y14dHJhTNf4MBTttVejO0Bfr9ggqiI+pKwZFXshAFe5gALk
TuEjSWOWg1NF7Z/4P0j2eZBnLbmTvCkMnH/wmKns8Tv06MfK7Wik/3wPcrbnsmzs5klyfjKskcGy
J5T2VZoblAAhvzIZAwzNSmcJtqOxb47Cys2qH3w2aC5lercIQE3jvgfESHR6Mgps297CZoPIGaZB
7IkRf5WVMjLIonNqz43L7jGMfMd9oBMSOLpPujtc7NuIBE+QYBaDBrWL03zsO+0yBeQLHOed6261
h+QIQEL1bYu/xJiMxNfJg3oPDw5k1ZgP1DcoFvz1G4qEJRVh9Rtrb+RWf391RoSA5yIdOLi33lgs
AF4dr2hqNe7Mvop2vTmrneIikJNgB3OHTPjjvKH87hm/0I9z25xm/h4mo+sBtopydYWfzpkWQ9qq
wWHcJ6fRMLVJWCf6hXh6TOROTEerocWC+k77OXWNGARWdldmL8h0CqiF88HqB9DqPiDPN7FWzx+Y
u1CttCskNTJKGgEO5WAZkRF6++ZGrcDfE5pbvwi1FfQRBGikPbLew9Wwc2wsIeElqmyTkS/ypgiw
Oq4k479rsgnzp7DvL74l7ixi7n3AyGniqam877PWnCfiy3zxfkRg6hc/NwOSt6wfPV5+vrDfurWy
0utzk7eaRtDvh/JirmCcEHQUNJbguP2T7IxBSbtWA++uZpvD7tYce92i8yx+AdtFk7ulRPOxTzcg
8HGnygJFFOPM+Du16SVNOp/6b9WJ5/IgWhTGDc4ThsM6yDw/LC/pYro9GlKI77GO84u7qOaq3Bca
kdbZ96pWzJObvIT6Gmnp5SGN39asA2iEFjtakK576rkMz3clNFcqTTUwv3l5A1DWrN6ESSpmPbt7
mN0piaL3OBO/etBQbX5piijsfTjhjJUzyTWVPplBkltsDawrQ469MoFX6MVeGM3rneSmcI5ZgELO
6LkBdng3/WpBb4EaTjczMkYtAHbJBiW+elgLdRSfL+QvBJQeWoVoiv7TiUUXSqw+8hfjifcnRQbr
sCspalhCMstiATKyC2I6LaLAk+RtAIVyGJwrB3uEaCm0Ht0MaiR0psB+KwY4HLmu36LKm3JImoZh
dWjxwNxr7PszsLHaYUEbZUhKS683whsdXQUuX+mkjZ9+pw3T6KfcCM0JIQwmhjpyKLXLAXwGBKry
2ZA4LHYzDDlXbLeo4Q5C8jxCLaVQZpsZqKK/VPGA71Y+LmZpgd2156MVTfHgb68eByy6PYP2dWg6
D0z7Ns4l50kVRrL5hNe76mLAv6x/DV44B8GE9Am6gTAQBhvHFf+7ST5nBf7Uq2PUYwqEGGwuWuj2
5t2SjQsCcl2GNo5qY4beZIw/UXy0F6cGHcFak3SG71mHn4w+JW8aAPuvowKijVRAfzAzE8JOwmzW
x7tTI0qPu4K7hUA0gSHVCYFiNLlwQlMYOqcwqM9VN1vqf1hM2F3K/9dxqwVkhVOK0qt3qfC6zlgI
H/dOFy1f3xPwQR4sWkiwf91vI56znF5YXbBgmAoktIx7+v5GO6u5he+n8/aVGYYyPOzSJhYlFb+j
HjD3qpfanctZCWHljJVGkMh/3Us9iXZ+QyVCZD9/AktCf/T+C0zXR9jy12Y/+RH+zPNFjVDjpYoA
KE5NfTs3TtiCqDn5YBHr807YRvsAYz/jZNVS7+9IuLzs4lWjZHBel7hu/F7NAsD09kxJ03qgUN97
LNcbe29vCR+FwnkdGGG8gW7bnnYi+IX0daX4VjaywjUsSTnLxHWvZXcRD5NQv+TDYnk6WYzo/B0T
i8O1fwbJpCSlJfYKEtcl90nHqly9m8SNSJmF3yqE01QQjgZbc64dDbf/TCsG8436lPrbUtV5fIPT
x6F4cAHKDxNhpfcXHv0izF7Gv+UaYr73dG7vVAp0ZzUxedbL7kliY8soqCQpYvqNpdtbaYMv2jL7
HazfvJjXydxUSSqxjvPcoiIboKXBtRfL4oOjNeFKpV3Fo1UBKq3/iUfCzznTtwyUQ48bpAj0ZNR1
bLePn6UfAN+rbkotdzOaDOSOyZKo7p4cJnQklhDuIdArnYaeZBwXJyvLyTbRCR+tO9vedm16FMOO
iDioreyY9ahUW822fAY3uM/c8oySf1iikDQVd+fsseiu1CGp84124wEaloHDAKqfgq3I2cPGcmPL
a8K5BNoglsX6N7ezj6j0JlkMsUMP8cBsfEwvO8QNurFPmzbB0M+Z0ni/AYqaYx8CbJOtaRIOkahM
o78cUgl7bQrxfFHiN5Qbundb3LILk4f5H5FM0rdLHoa7AnROL1HIyduyiqTJ4KbeEGFPosU8ht2e
trGuCYbwugKmw5d5ErbfXRVbwH8hKy7Rou/sW1x0mbZZsVKJL5pLTnIq/LzNWBXiWXS0IczfvayE
xvvTa5tHFQlguVW2hWCDkbNsnVoAagrs0DdZDwi3ttV69ThuPtyow4IgECxelQYRnOXGRHfUJ+NI
4gP8Nid6evQQy8hD1+RYWsMSOx+pm3Qmfbtoj/KzpS2+LpXjhRgMYNkk4P8S0plJtH0RcTdCELVg
+f38uybgBUja8bMsfVGBU56Sxb3uYs3k8YXdtz2lbZOaoSv0Ww7DcxGIZBxTf48S+IUF5G3d4Xu0
1BF/uQsXuZn52kGf8Ng8x29E3dp/UbZQXZmkZioN/VAAqvzJupNp2FNRqDDj4rbxLCbBxCZBzVJ3
GJexHuPjIbSDzKBRXAjYZnEH3V/rqHJUHde95Bpo4CIzEJkBKEqBs6sV+DPg0002/+f5KPB+7QhK
S6P+BY7y9fxOnmKbmd+uIqLINZfbkSc+JOD3eJ4sB5t3BB7dImohz77mzhxTGdQGZOXThNWKW829
oeNcjnuZWR4yQPJT6Wc5HHw7rCkUFhj6Rp5R1mJtiBGwwJOxtv8ga5SnTUKcxy7GbqeOQqEJJGbc
QG3QqziAQ0pC6KvF9R5kFrDSazoR3AaOS9Hd9518/WTDLKaqAJufeswzInbX47q1eOOto+JUcpBS
ixJnaE8Q+4wDY1L1hF/o1vL0nHL+taPz3OHEpeS2cgG6cU7OaWYa6PFA2JlOp2McTZZ/2AkJSiqU
qkDKD9hgbF/j6fBg3fwgEEjetvVt2oM23f1RViJgeD8JJ1QUajGYL1r1tYpO9hKqKwbuVw5+5OK7
nTSUYLzOkcQhQdhzK58HG6GotsF4yGwPUTm127TOmz6Ppa3jLDENg7pGniIQ7r/MDUhig/L7sKlm
DiG5xNbX2ll68hUX5CgFyMMHKkJVwhw/6xcc6Sajb44i10PUfmuYS/ZF/95zBlEYA8CJVSJQroX7
PGvAPA39fAWaB9KsfsDeUXqbAQdc+gflbFD4r+uQTHQQPtPkrrn62FaQvGD50OElo2//5/zTg94d
2+3coeGulkk+A/FxV9GZmz/yKmGrrWh+HJYaC6Mf+xS4DtHir8GsoxFwWxDmPcAyNlK978foeZMJ
93IecFczpomt0c6TnYqgS3Btxr45g1VdBO8ybb5g2QcozUFZQWBQBdGBTiBznq9a54XYUDN4QprW
2pB296E4g1byaxcQ1Nlg8g0ZbaQ4mmHmWeiojNZql67n9VLjGL+/5doPusYn93juzoTNeIxJs/1+
yTDTk6seoEH5lTHNvlOQiMQOcEFl5gQPGgbhxTT4LEOn0ndDh71N/EzXwHDRK95aMmB32eIYj7rz
kSbVaaMDXLRo7o5AG86vanuzEeVSO/+b6ufzmxwNV8O2URektrKUFI219TAa1J/zUTHJ4upKElr8
9NzHiWq5lN8cYV8w3eCgB8uq/aP1jB7nVY1liYvn71FfIu026aceFoLY0dljpDBJCSulOSfgxemD
yjw6td5hfvYmGsoI4BL65oJJtEILVoHmVtIODlo80+puPIOSCbCtIqj/aG7Bqim9FlGK/5fjcrQj
ca9J8qzLYU7/QJRNV1euFG1QLlJP1uscjBWM3mA7Mk3H2QJaKplcDqOwWqldoG5XwyPF7E9M0Dg3
OY45y7d2tbF4t79mYFzoVZYoKMhdXPdK7736S7qgyc6PgmMtHq79BtMQYezJNiOzZKxEEQcKAL+M
MGV+0QGhJxMWRUgfVqTvPzpoZ+DwNserfs5sxJOzoeiSE72MEBjVJ4FVL5uFsum9RyQSa2DmKTnK
RMfF6cF1XMpYyGSjw5FWgAS4MCKnlxQsqM2TyETUPaWb8nH2ALvxS8eeXIRaXJ/QlaFr0+5HWm4+
JqZULmSZL6UEEgBexnbQ4X/Ytuf176h/jIunN9921UYzocfQslJ9jjrs9PXS7n7lkQK2SMnD76Qw
Sse6uKE8udDXX4QGleAqei27JRcbQKEZJif177rqIJU+4iwNmSdrWSMcadxej+d8YNoODAxEGCeR
55RZBZA1tM0AfVmZHyh7S0Wu7kHGZFd+c8hNYw18dqLolTzoXo0+wtD+8DTXwc3+cpc5wlnbkxEd
gvrygjar+FdimLfT6qIkZ6IMJ+mqNgX2ZE2nv5qLVX26F4KoHsq8y19WO07WFkS9gYbG5pxki/+r
06IUj1jbU+8eYWT4UZtUIPI+r8EJ4AlADlv6JPezPvl9RjTI5DcRtJ5IROZzwDOkJ2nCCVZR9Rc+
rCv5gFNvW9thn5ICE/p1C/5rWcR6WwrJcKMcCfBSGxDDAOyvpShboznFu4sIXAM8Z/+2o1rDqek0
tHvhFUyPvYmiHx6bZPZ/j2TVTwrFPUbI/1GT3Gstf4YzwhRn7LOcU12TpLWdDQQWtu/pPmdl+oay
/WGzs27MG16frSl9zQVgmGyEggkkGKMYBqa/CU10jPyfCO6WB0BNvJutdpyyb7ulxgXKPj+eG+nb
MRz6nbHJ2HhCl3L7dqzEzxMzlIGs5nUGVOE72xV5W6d46OHi+yKvtjwyFi5QSXFVyY/+vN8Vwaaw
pPBWijPjT6aAOx1gDTDCKHH+JK0eP2E9Ab8Qgd19VjZyDTVxXMUFSG9wJHuguNPvsw/mWFTCQ7jl
BeDvDIOe8uMmC/emkFBlz6VrWikJUnoy7BhDKB9s3zNzJ//gDHvUkbgxc1QLWpcnTOP4hvUoIKx4
eUuAnoIe8aTA8ChmVD0DpuUWFOVRu8alDqXzZswWgOt57NKt+H7GHyRYkHqzN8F5axRi98+RuwT4
h2vQE8SeykkL6Ij3Dc1r/dt4eH9Pl0xplYTB4Bu0cam9YbUFNBxaNwojvf7IbsJcjSUqovBRr0aO
l0wMtojrPxXSFM8OxrIL+C4GkDP0JrVMYorhXpY4EuZU5T/2lHt6aU52rZTKDSIboVeLnV4UhRRN
mH3z9i+B2QUQTxur329oOfJfN7PVb3gYKBbDZZ/64ki5G1DTEiMJ1wHLMAuXi3TNXgE7gZeaMa7d
OpYcLVn6Hfw7Dr7+AWu04HKMlvSVQrho4RLm2eCBAXiqkcffqEMSgdT4tVfkSahk8WIHsMsycRMy
AJmFe3EfN0jPqW43hFjWpH80jvfIwPMvIsXPKRqRmJChwJr2glMomN9f1E9phel7hH55IWjj1Wlf
CVSdXOMpxGSIa77o8xRFqETLPG0gq11C9SeZ9tDiPula2QFF/1FFCoIQ1mSzjunmdKNxTh4vrX4D
N6eu3t6LGVp5+4Rz2Ul2nIuuIYKW5/TE1YzBAHSPSVZGC8u1IU5foApUsRtf3854cFZqZl69o77J
ylVqnLaAitFstQ2Rg4NiMHz9ugL2y1DMwDNqh1OBNhQXpDsaExYlg6fbACXu42fTccz2teXI9BgI
ZszBVfHq0Xjz8K37Wi6R7kxH61BCuSZl/FCcjlbOQkt3PShjEVadp3hrTAYCCqHB7pnJi6qDpnRp
gt1pM9SFWuemj9jYo+BCDK2atIYBBWj3yDdipzdAg6XE5vFYy4IrKFfRPdkGwFSCRf1EkVfNnFOX
rZzy1QwAvlHU4fFBEfFcvjyzpHT1xuFAApoSu7KBFZhQashcLZNAXAcHKownZSBjpMp5LS2tHwER
geVK+kubeUN3BOZqk+KNNfq1csKnIMU0F+5WB8WQ7tfpgHirVtT9AjdYxay+fuTFOvvJVtsqxHtw
DItIkZNrSrzZZFlx37uV/E+2EsXJDkTVgbXZqi1IQyURFBgLxXspdFjRyUX1x4bD/70sZB1IVDQm
6Agabyi1rjQEpa4IZZ/y/MW8mA/zr10vMAyMdv/OQS0D83FyTQNCmBauHEmjZYVg/Zf9HGyGKn2m
JfTDGguzwpXTS5i06MVcDQtovJJy9hXbQ0qBjwxb1axW/itFzmkDbQQfnbrRwcAPUaGWJZyMVPub
sWxi6iSE98smub35ZDGrPJCce7If411gckTMb6VCVbI61TD94hX/o+s4SdGwykrTcMNeMgHSNoyC
dE47inWMLvu/upjY5A8RvWZg1lmpc/zAFujAkSll2MSB378ftSlb2ew48ejazSDCe7oE5zUevQO2
5NwEJiss634NlsnV0Ms+/rLMbcwPbx/IydeoyhQD0yzuq1t5Qf6OaWc6GO/xSG+BAdgizNS5/T4C
9EtcdvptBzVBX7qiRJBvGnAB9Xa5D/D01rxcU5QA9sO2M24sxvjlkWEzc1eZsD7oPGSRVwdQAbzG
40BInBu29nXCd0CjYZSdHT9GhBKsTkUzR3DX1Zsx0w30KWQLiRvnRAIw+wb0qrqxk2E2DH66yd6S
2n7sDt8rKSJoUse7W7BBq9VAxPlA6a/BRtqrVjqrShWW0uNrd8KubaYR+lnsWQOC/JoKo8eNBcgC
Gvd8FdXonTDq3qcJFDHfi9x9Eo/sZ2tt2sdutOkrZAqTPWiOOgH/XevhFrcAVEmtTjcOBJ1f/RC3
tgmQRYVlPe0PcweZPLeEd/BqyZ35Gq48XMWHIjaCsGGWyK+BSp+dRWc0GC8LayBgYdIGz5G+5Zvn
xLe05oDxghow11GAuaAf50KMxzOEcBYyg3PWZpK0zc25Lm1eYxypdDJgtDcq9yi+bm92b9ZEbNM5
4gm5bdyhyeEKqZloDfmg+01BACJbzhpNz0Isl2S42Ne8zkkXw57dzCKiJMt+6oZkbMyh0ei18sKg
k9G6vs9VpHe6WZD59wI0eE8bFG6Wt/0eoWC1vsliTKQ7RvzzaJA63w3rzMdiGCHtNiiit+7yd5RF
bdwunsXeNopzPbiUw/rgD2lsRUBz8vsUlntEjpShzXsTnAvl28ppWgCYyP50AweK8QaKSrPCnXhk
uDovjmdYMPENjiVhKcbTWh/GUmBIJ35HUF/unIOqasvMk4UFchaBYFdTDL+sWpDnn7x8u2hDqJ7g
B046IISkwmoQckvd3lfDlwiceXbNJjnSXGLQQ2VRsnUvzKJcXdaKRx71fqJYWCBkcAZgBpVeA7x8
9klg5YjEXKkqfQOIpXqx5ZAeXF9HMYRe/9O6i7t5HyHSPrQaYY5bNIUhQ/3b5BPMnZoNl3UzR6su
V2PQ5/0Zbc7keEQryH4PebDovHmEwt0HCW011le2GhkyPRKtnE6XbpaMXFFvJy5sFlzvmkz4gWVQ
7wAdNVS0RQLZl35WrpNocpzOZmH1PDACOi4xAktAwlFYnssvjedKhNuxZJHZLdrw7X1TcFMPhR14
8WVb/RlgkI545hp5TU3pUfJW7QEHzmMDeGCpwyhS8UXQfsMs0WagrkU/umKq9a8xoOtfJ+CVkjqr
3GY4lRWf38QBOzkiBPTuwBdZ8dxFker6grP0tXhAyccbQD4k1p0mh3oK+qZjM/4Hy7bp/DM9ntsE
mHJ1MBwrPScAEiLazONnSywaD5+4mWqyH3TID/szsy9xmnTYyKnOagA0bbhjGUr7LSHNl98t1H76
2iQYB1klz/i8x5JsLAiv3e18PW94XWtZkRha29ZOFRUgOQb6/h76LgIjQlQBkt7PLWeBG3/p/907
cvbR74GauZ2pwO1rSnUrmeGTvSn4lhXEsf8AKXn9NF07erDXP5ES+1EEDb8EYK1GDIPXQ/VNNnvd
pcX5SAow+X//Fp58CH1RDfNIStGqrFwY2AYVFe//GkVvDmEXh3r4YzsHk2N+EqPzSIN/emU1rAJ5
bl8wH9BxrwPvq8m6hT9vq6qQIdMIrIye98AJLrfDq5ZXCdCF0rtMB11dIm5Du5fGqRyUmLvtQfeO
DwfyvbW0h0KAaFxuCwDLIjMU750cf8DI496VWNGgcFsiXmDpGeWfZ0Sc/7rm0YHZncScYubTnNXr
hamVwLy+YI0VQ2S0QmI9YzY3sEOc20hIkkYF0LxJqtcA9Kfcp/e+EKp8QAYzaKULzy9MQhi5r90+
DKkwz+XjRfKkKR4T/Ac2akxYeJHY2LcsgNM7H6bGu+yta2DkfquerxYIS+VkDfblJdyHdwN5B98X
9Rk2uy1LQiyy4WwJAtfZF8oOGNklBQXYSFlgJacnRxxF3o89kJ9iR7ovETwFe6UAvx4FjZ90G4K9
aJKvVt7hnl0CpNTHmiI5RYcTOFplUGyM6I63KNWVU+9d+baxyfRhOxjc+1Hjnr4kC6JVHNxk+xHZ
AzTyUCfbvNH1S0xbMT532p4RbrlH3GY8wGAJAY3+2RuCc14C493mIdcGBSsCivGNZO2//SnPMVs4
/A2tv1J98kCfaZT7OFBJ5Znv+Ds9MoVhSGoqlWtyiU4dKrwySvjGZVTrZgdrWk1cCnMr+EA4EnNm
NzpHPm/jBVH9sHeKp18PVgYEHKEVToXVE5jMvEwgCWjuZSsIoKI4PzL4r40NwRbn5wdojX//RL8M
qVs7Vu6xCvVzW9tVbQ863bYCdHJBfgW93Dds+Zj/1I9moVj3GD8LLPvR/sFcf8HFxhziMNBtJIpj
PuOmaiUaZd9G0wRoTgNsEoTfYClujgJlnhm2u7AH3p59rV0LFjcVhawGFvqpL98Vj5mKDW6PIbe3
mVmwPIlTuPWsivPsvwTWVo5PyfGMlJk5v+o+sszUM3zValT/X7MZ8EABe+5iZudFaHdo0Xnpm0Mq
pS6b2fEmVkrfu3BQsn71XmdvOl3WuHksSq8YCcwfag8NIdCQi2cu04Mn3e1imQjNYW6p2896dyyz
JOSSBEs9CYXuZak+oobfag0+tczbsKPKt5YkVdZqfEtW9rw+sEq1eDzdrF6L1pwx5mJBaTP7WAfJ
+PqEM9dxRNG28JnNXVSWrgToa/AzN2HjEYlGjKl36AlrHuQB0LYIh6QIHvZxwg6iPqOcQVpCmUQ3
KlevleP7/74D0i/GCSyf873JG7j8RZL+tZQ4qqCtLOvo7Dytr7x6AVwV/bBryUknz9w0Lo/C3wcf
QtN/Bq+p5xxdSKzk3/gK9m/XySOR3nP/jjjOT/SOXnUuE3iwCzlCb8He29gkn69/uKLs+cfaUQ0O
YXPsXDmvUDs8uVCnMGlw2YbjrlYv+/SncIsRdnUnNPD4iOGVwVnPHB2bk65a+udvpKG744tdN495
ArcpFHekGJUWoP/dImEDxmld/ldwrWVCKL/xjhiYnn6NLT7C1sgEqtEkz2yz1PhrpTITW1yIpXx4
i0iufNrypZPy2NU1Bc2BLunLmXOZpU1ll1UgL01RzBTEvrdwJQMI5/XlXqAR7i3RKpbyrO34mnc8
paO+hrHdXROICuBzZKJa9MCEqhsUcDlaYpQTm5Bfz9yPbtRRpZJRgv2naBeuJ3C4NbmYroTTUIM5
N0BgHVmn9GQ6NPu4afzuTmQuZhMhGEiFUHx/gGQgwHDGUiGdzpHwPfmJyXdTYlJ7iUnnQ4+3MFw+
f84Q3FslahRPhxhtTaPRUL0OgISvi0tbwt+ZDlHzLfgpoUAYDnu+3dSlNyK+/kU6Swj4FGLih5IS
E3sdNea1xVT3NOJx19OpnOCh4JoiFW51GVEZqFh+Nf7ucKFTiWhWcHkcIjml/im2RHs73FWJEiPd
rYHEoj7Y47MehL6PBjDPGdJlc1dV5l+6Zl2T205wpPchc4x9fxteW6tv0jwtE1v7wkicYvi11GNE
6Uqj+aKdO7xQo+fl7RRQ6o3OnJwzfP+wtU1g/tMpQ7x11WSdovFSgYUUnFTNA7cYdlT2kvduCCgt
GWDKgm1PbIF8OHXKbzlKqEybrB8BRu7rUCNhp1RXHY3QXacBgGrPI3PAgEJky1POMaFnpox9BvJp
UzBcbU9IEAWR0FjfpAOZPEdlMUD4m4TDROJarlrGQtgJFTiP4REQSRXiO2fLGFkKxo810MXUFTxu
jzjwzLaKKfWi3wgEVIvn/1sQ1MQpUmlSfLrFkZtauJxbVaNi8Mb28EAIhHDOAyq+LwuVOPEzhAb6
6t/qfjB78Yn6nMhf8vzzj42ArLmZLr/N8vidBG6EkTwfNHoiIID0djfxraB6CJb75ChmMDdzATYJ
1ac+ROZH0bRYLO9Eo066PFFuO7pC4va6/Od9WdzUgJXGCoWeIIKcUl8ivZnJaxIaQWWdRqTrvdTa
z2qR8cAyczctcmONGPmzq9BpZ+UKETkd7jDd+NTfNLugrOMqZ3LV2oJQS4FnL1ck7STdqvZdRbaK
TB22AAsJwX2JlXmSf1cQdZMHYITONBSolMzKF5gJMe6dMWlJemryH9j/U5zx7RLsuelV4xVTpykp
Qc+Wb7Wvtr7H2etV2fE2segtC1IQAJUO+qTGfqbn94PN1buL8Lgp0XmLOAlhlQWHeMtd7X6nz3FQ
vXlRBSs5UmHUQmIWLxh9++uvSggf83WCgAxmv8yAaHJE7DCguvIxsvYnaeY4AeTSFl9An398cIsA
78PUuozkejkoTq4bYn4IIiLz2Om7qezmM8xTg/CAf1/HmMaFMUAiw4K/N+vhcGE+2f2DLfSYiNzr
3ID3wX1UH+s/5YbNCaX4eVTkbL5DzButvgr1Wab9lsuIENc2kk0RufZo8KxdOLoI7WobrnE+TkFs
QOvzhhQY9R23Onf4PwsKt+xNovKkUeHLarvI7ljbGM1rfuoLaK0j1VwzPQA3fara+h0gYZcpZbC9
A0tChXOv/EueI71wNyzYjczjSyFFdIta/I3/kd9LUed6fULzQf0UXcwI2bKI3Z5ESsH9mMKmXfyF
9j2vm1KU0GuE6ZMcNyR3AA5xrs9zQ42D8dth/KggEgBxBVO9QkNFqVV6Q8UP6lPgk6fyc6U+OWGi
DKVmfUJuE/cK0aZkwrzSxICBT73jIRnDy9PgvqcocqqJwur9vkN0jFlBVA0bk4NywhQoYWv7wkLc
yDio9DftFHehGHFscP5wI3A1LFKoQXh3aiQBjAtC+SAjmWwZUWnCzsLHVEdlBHLBag6zZ4c9jvQQ
v6/gR1rhkwj2vOgl5k/U6PlfDI/xuqgD7lA+a+kexrTEj2B/OUkiYYAZE6SjyLC4nKhs/LdsZICs
RG0TnqNwmdEI/g2oo6mMC5kth/OcIccoHPNymprKqCqo9YesZq/O4Wmt1J12JFu2JinnzC+dvzmh
eELOpoRKnX+ZnEiKnR+DopLKdwfI1OEMZPJ9Fs/5nAhQuDwJiT1NMvyJ82EeDzNAYrcq+I1HioA9
P14q+TRcdHDx7jggsNrnCzF/e2EwMW44It+AbwL59dOQiDpvkEPVwMDmZF6BBBiPFJiIh5HsZrWN
69YNNPkYWWxFI1CxOFcjhZlECDu7Q6fbJ9SRKQQhG1GV1qWgv0S3MVbf23bQoC2zunOZSLqxUg0i
ilxcp8voODC98j74B0+QAEtMCHysDy+r8oOZTN8UquhFzybfQDlAqOVXBB6bpZM44QF9PTs/JEPW
TQ4ufRUjPgPdkayaJU2GENYGKI+AWXpi3E5h1SphOeWR74YBQqv4+BZEoJeh8l5ULDQgiqr/WADR
CldfnqkaMu51JNUdmAzsI5NSHZptuYKnIld0kWnJrDGXShs3a4X92vAbsJ2M8n0fIromE5lDzH3s
/hbQyDTzzms1OTrvjmjvW8IESAu3CVBTWr9XJiS1srV6z/YdOVIxzrL3tOw8z9JjWVVMGIFS66jV
z2vF7nxC8HTyehCXxnEGmDTMbnW0aUqoVGr3dGHgknB+yXbnK+l1MmtZTnbLHplO7nGEI8CWM2f2
5y/84HHTimFJ1QBk9IhjgZDrNFtDhRNVNPVM6Nc1scCOIGHXOmMSDwanYyH2DCJXtX1is/zYsYxd
Dk5p6fdvZyOfTorAcPD8hSbK2Lhv44AS7jxkQC7AO5NA3xcYAKQJgvcpaFY8LGkU5hbKj+GXh/Np
BF7BDylJYsix4MaXmmosWh7OhCvAfsWMH9vXjlKwB/MtzlmUMRma0C8NjCO3BBHZvXF3ijRsAWZs
oypf4jn9DejZGexx8E334KsOAr+pHCogakAYC9d34lpYadYcqs5XYxnDU7taLxcUIlGJVQ7KzBXl
wZuf/pSWjENUEkFnqqND3gaeD7qxaPxTrUrOPGba4hqoqzi2PogeYj1pr+P2qczQCVXK9LdHnHEz
0omyFGIYXhxEZRE5ucZlOGfNHZcE0L4//UJ6zI5gYkMyjdQNv8a3wZ0Jw8p3jnQ5/9SdzSi2JTA0
JWDBVhWXmwwrNZXzMxomgMAc0hrk8+5EkG/zx6RWCgck+02WVlUhInUbUMIUYkN8VtoWneziksr9
VPwvz19S/J16wPx40BYUKwWglS87pqNJ7DGXEWXe9oGejdJzzCEy3JSa+oaw1eMESaUJzjmq9C8u
St0c0b/Z3idOGXC4Xpms9yvmJPcljqE3ZvXN6sEiWSkrkauGaIIb9w3BsIOzLckaru08QDALkcte
PnLSX/LMOwInJKscja/81TpkF1OLoC3J/OEUBYZ6kgGG1aNSWT1NfuksE3S9jIQQCEhlaX3wM769
PXkAkeleEJ1OeIKExxAWr9IX7HL6W5C9/R8zNbzc3MzYzK93sRVVAdNVzHwao/CJDSHlsK9EPlzK
uZ00MKyjFWJge+rhizZ4cojVNUtKJtyu4A/uZ5ATu1vhxhMRzdldwQ2Y0d6YWgcU8bAg4TuXw6cK
SeUVjyp2NdDAkjWngpMZZyuilRDn7VmSMZ22PbHsK6ZV+gT1NJ40d2vR3UAGwP4AWQX91gQKFgOu
GbKg/ORATcWWXjCggS/a9ZEvXKziQRgvcGSiVl4XONF5J351Y6mKtyIKtryxJjh0eGHCU7kvjcBv
DxEagPm0cPF/kFtyGtmBF/47UxA7/oZTzA7UIZTiQ6+cxNUtQxQUKK3Kcbj0vInwvMsEAhunAAxM
fjHc/tnxJhl1ov+OcOi48vwbU/uMNBzma1flXTTb2+EKyi3Ftnqqm6zl1EbQN4cBtRHZ1fUOWXxu
lzhLofgXa6tj6CZxrlCRMDBz1W4GObg/tOhi+RyX9z5hJO9zQ4w4X0QDi6a4bJWqViUEBSKF8LDs
E7Qx+aPaUv9EIIOi8D+Ipcq6/kn1oECXRWWogwKwYF/jidnTLF2Bx8gDTbiimHqXaZdIamR8+Vwn
3XV4tc+CQbWSuvJ/c3q5PDk0GlwCqyRaU5dI8OZJNDMB0qngnx9EA5vE/gxxJCu2+sdoKClg67Xs
5L5e6eZvaRlJEXZE1cCcGaLMT0emNteaQM7MkNyADSLzizk6FA5IEVex3CYrrTweGECz8/krW8tQ
Rt4U+bU85nUDZNCEhhIaujG6zYqz2w38WPFQlyrnp5ljTzzg1fQbjb27SZf+mzblCLuA0Mg5WdHB
+CjfPWl2vsejduUfD7Jor4/4sbKXo386vXEQKhU5lOcoz6ujf25j4DYCGkape1QqlGaO3WhvUJWN
FOjimx3oYbbkGHtzhgrrMN72aYIR90M+IPM5QEhv38BR/BTyp9iV/4gsJN1ZGrnOLlB1K6wDrLY3
w4RIT9xQN8/NiV5/hnh8fvsLH9euVWshcyGCc4dqT69wBfQb9xTSMtfu9GsFpuGbJV41iJjm1OD5
m79hku1zWibDuNGaPYofRBcRNUZwa8K6Imn18O6EfcuBwvt/1Q0qYDs9T+bHM8vjVyakqzZwMOia
fFcSl14kQyWmvu/80x5uU88i1JK8AvENTxItZFYPOZEWvWufpTMxnkwro3YAF9AcfvzT8+M7aKN0
qXZIOpN4cZlZ3Q61X9N03JwxWEN6EnCVBf67/XrSgnHT/KXc1cHgATHSZsgyqX2e0S7FZBSjXm6x
tHPirGnpCQfNkp8av8YI/VEqeWEOGH1l5klcr8WGTczu16u6M63AjxoMGhVWz34mJ7mP35XncbsE
MNQ0ZgqryGmnTuH0Q+0xLEacfm5wBHXpmj2JTZPSWon2QNwGWenOe+n3NihKaW+LIPUbuKBRCUeF
LSmwUo1nmR13MRnXybko56hhvwLa6g2UWvwuvZPmLlT3ysGIfigoAoo56vJiqHjePD7rZ0ikir7p
mVtadKHoMGvT36JGNODgyfvzEpwWDQQSAdjn8RKONwK5xa6EPRL5yuQD83mkPuT5KO+SwFyGrIvO
BbtM7zLZlM58x8BCV5T9AhMtxr+zcMeXggj4syNg3qeKqDpuerQHE7LYZO0NnH6qB54tbIS0gX6O
/nw75ArtzjZWx0+GUzq1adRAJOmOwRdWOn0+hLuniED91eVdVm2DoVzhyozmcB9Qnh3B97BUFUkq
IJaOwbnkMz16Kbl4jcnGiKnwlbOtXlF/Vd0OoTxsYUBaCUZGglj2uGnwogpwSp8PfjWganj+lJU/
82qK8KJ0WRpJLshIMrGkMGJmOuKKmr4Rrcgz/5da63lo5DCm/qyNCOe68sEb6o91+cHKectAm0D2
A9BRxGc069Z0Wiq1T/J7ett1fFuxk47fT1nugUPn2P51On1qHwZu4xTHbdJN2X+Z83M0smaUQaGs
YaD449GBhjgwbnpgrge4w9A7r9u//s1BT+UEIjBNcHpaqK7L1JFRegzmwWgGX1thSAP1TqHcVet5
rSuz7rZI8jBk3FyZdvvcnX9VjEm6Etj6RSWnpAW9jOrgiGhTQhA6BYjB759dFTogcnW02ehnuDud
HXb5ucIVqNd5IraUCSpSaG5qAKOAEHnkS7275LsLA28qAQIH3moJSgt4Q/J7diyJbRG+uB3pank3
c7a5p3sWRkPYhLckMO4a3XHPGmtJ96mD12So1VZ35bEouHCtMxhAohyBZN+iN/X6ze64pn5oB1MM
Uc+60JHU+w7xHTbTcCQfOspu6nvcyFf4xnZsbYrwjyVjMkVcDqwB+LRngWbnTZNZyIIRGq0Bq0jo
5Krzv/fnh703l/PuTwXPq8Ytqhs2leSkan3mEXN8WaRinBESCC8t02tN6ewlbvWcCgKL0qJAmUic
9eiRxtI2foGgb/FrvwFcxZAddscqPN7W36dGzZzTBeu+G4JCWBs5PW6TAM+lh42TyYek0XOZYTfd
bflUA4H6twI+NxcOElAS/6sboFTVJdaclIGbguB+xaTtzYQCOOWFOmSkQwxNBb/aVCZkmmY5y4MM
zaexTbHjDHfXfgcrpbrA1baoGLsyo1Nc+B+0nDTe3rIuX91mABIlhdwDqYzC+CaJ/QTVLbZP3IDf
2wQDPJJgFGz0VpkKMyjb2heaCMGzJ3TOUwCgZ/9PyHosHX5jrqGCBtLFoBOp5WXVOg8GXgitOwFi
6qvDAbw7BKNc9DxwT7RilYEIVh3lbScRB6AH4QE4TMVnr6nubdoejA19FlvQFqlljS5NcAEpx+ja
31VQSOFt0Id7t5n58kxiSkpwJy+G0470IR6cf09o82a6BSdYPg6LtO5Pnt4j6bi7Dv5+bQpefpG4
AaoqBjQ2v+exZhR9XE1Xm5vlS9GkMN3zuZWVaokYo5rTy1759no8lmYgHcsAuauurCVULpZwbwwa
Tyo5G8umRrCKCFEBQieLJjoIw+cynidqRnrsXbOhW54oCNBcKSJMy5Q7/VXoBIaNKhW396AIcZV2
uOyMD6j55eIlki4iiypsVyCftAaylLOxDqXz7CRB/dQbFWUpzzJv6OstzUwGkA7yASZBnMZD4Qp2
rSCtqUeH7QslbxwYC7SVvwnMqOn4gzbF5IILjb9bY1ldlCJTyV93rT17j56qM2RVUTm/rb8mfNnM
mL7Qu3BkggrSrkytdobw7tAtfveLYmPr1tE8D1qul6m2Ey1YT3wzTZc78bpd9hz+Q/gtP5BDNMQN
4epFU89zLNpqlX3kXgxEf6YgyVOgPGuy4uip0mrzqIKIUbXwUxDYjLZrIYOXlx/aymjMBm6drUqz
0ykdxT8tifGnoUV9CQ5fYrMIyU5uQK4ALrC9DdlwhTRbB6xpHyTwIJN9Om4gx79pzruPLqWNIPQ8
qOhqbagfKl0hwQu4iATh3szED9/v2X1C9CPkKa1rDf/PREXBlM3Nh3TvEzPUaXSme3XT64YFSZNx
ZOuQdqowMEVZXw6jO1DcQeRmANVhRQazR/KkPb3Y/jJ53KxtpZXdEtnwIv+4dzc0hjcMpZY0Q9Ru
cbh5FhlCpyszX7At055G/E8vviG3h1P6A6Yht/SGXWVQmlxajGuFTDedsKa0iqzk7up3fwHrWpVW
fFuiYoAtoFEAFntxsJRFaD/8FQYelVzvC8uaAa+g7pIya+IkTabGGpD/eWt1docrPd80IpniZHXy
/3w0n0lAzHvkOGUtVogZxlWI1wzudpMRVMIIQXl4BqyJrR++6UZoKLnH5niyhmQgzeErKv4qpEQm
XpHUlpAm9VDgTTd14i5aPp1V9k2IJx3eylJqugzriXFvdrzfmGx0ItR+ltdQ8qvJPPVvlONpehLy
USEiu1xnEDe5qf3Xt5ANiFVsudunildE9DDWy9wh+bT4DRjPuqTg9EwMVRzr3LS513jOSLyUBCVm
7hvqhqknXPYMR4SKAG3+ULvMSv3FvxXdoLSa/OFYg5Udp9oO9Pf45opBxGOX1l3pWu3M40ONKWXk
I/qSRzHZv/S+LSwTeiK6VTYYQdMV+X9NfRiXaYU9MtivcIJSbZfoD9FAlcSgvDBFrLgDy4kAgUin
llsewfsCHDG3B17ipuQ7g4jE7wn/DaJIjvHr+PAf0e2POkWntOHzoEpY4dm6aTPGiij+JwI7bAhS
Qn3g3zvO3p3g8pvGKOZv5sUO0kzlXXe09KJ/doCVHH+G2kz91FlH5gB9MBOFKhclDyq+H8KJ5s9U
d+3yfCipld5Gra2As7wPmtvBuKgf1AWFKQnKzng9552Ylpx5Rd77zWyeZDK6a6J+0nm05WQiUG80
qNmPHP5ZjQCZSkM5OI8cVs71WTC+RhbEzUPsdKIhLJjfOQ2pfnfEs/41wP1fp+aV/kDSb5tEDQLB
gwoBthEdBa3W8TjfMQ/LsQVJxqRwtKdwo1CUiN3AzDowvlpTQqtnQLFMOedw+pZV4jWt3ryY0K0/
j+SsdknV6r1ffXTGTdBKhMjkUXPP9xO/8H/QdQGyfAg96zl4jWVEQ93WrO/+14vsYIZLwIC7jhF4
bGY2dMeuJ8Qycve0DzcyFen/JsWBRlRS0eHy9oqXWEuqAKj2wGVuUB/TZhRjqjWbkYV5/Nbmfu1m
Oad3WrtMYa+XQYuDuWClG/G+tUWVlcGg0jWLEK+9YewYNJo2FsTtsQCIfuylQaTktaTOdw1Lfnq+
9ynW6stEtR1KxKd+tmyu1uafRI30XhfcBiy2mQnTyh6/HP5AmqnDnW77tuSxjOBhxp/AcVevsnnx
dyt0+1cBZ9MQ4UKfisEPYWIAsJXEY65c6Lh+g23qJ0Q5c4lqRcRFtoK7IEQtmqdRblt5NR62W6wb
rweHtEiU16oERWW4xdrGqqqAM4+5vt90gSzK2IXBeFLhvD+G3FzuCp6riv+w4KbbhuyFZwWASQT/
wMtb0dAwOvXdZaGbo0DQRN4Q1XgLRU9ZiZ+S3NlH/y4lnojAvsiruhVlfN0tBQcgYC5DcOo5BJgc
G+2WsSL2MtaBUGQH4M9FRIHSJvevMMudx8b9WHjjds2iDCEhW04pOmvwWHpZ/7YUSklJuuK3zC7B
51wnCKqFhs62dKzycx9yri4FbRHqyMa3mrh0iDEsgOJzvAzAjSYAfzxm7iOUzuX0A3xywqp122Po
lbRrKd/fIPTFL97bumKTr/eBoaiU8bxy/Ra0DYV4c5KQutCwEAIy+TfxH/qW6q2QZZSZdAgYw3pI
jyw+Y3iC/itNXMS5Q6ZapyVFdxqaUnoE2Gwo+0G/lM0hH56v+QOmg2mul3nWiy4iAlccsIVEQLP+
4Y+Yy+ZLYVW1gXKWaM/QB+224zdPsAv4+NJNDuRN9NnohKZMpBaY4qnaZxbmpTIBvB+sT5YUHazR
GYA5z45JR3RNnuC/5duUBUkWLrwNaeZs8gYvp4HFpxQtLweFdnDMq4lr1SRsAzfp1PWFjkP3L8E+
fXOl+C6L2Ne2Nm48HJ+81QLnYHzwWCQ9URUF2qctBPGXO+oG+7PzAtXSQ0MeknO/QaVlePuTXYKq
b7hRj7S5cGrvbMb9neZIV6EIXoeqo0u1uHZzkI2jqdM7P1JSV8PRyEaHwN0tNR0h67jCLMQ+N5By
ZJ7BXrWRy1Pxw5leA+SSZLnsk/OQBcxBJ/aqRdhg45GH7Xrm0YBVqglVj+GmS/AX8dwZY1TbaH+b
RQz7RxBFbK78p0eS6448RO6AeCSRDjH4h+o3T/dkVmTGtEG4OQcEcBaVRnnXsv0hjLkHM0B38SOs
5z1lf9UOxU3QNplctF0tOnOFECkO6rZyelHEtBvOyqLhwWMOV4ilE/OZZz6txcjWxNkOak5mPO14
p6wE4Z1/g/rE+Js2W5V4Cae+gWNSF9LnPHMKjq/HlxFWGbsQ/UhNN/+JaAEbx43RhVNIOW1VicRE
aW1lVj39f/FPi8bv+tkMvSCNOSmxthx8KeX3/Kv1coMgkQgnls4YjAKRL4QfT/EEVSte7PglyNbB
+ivvcB21PZ2uSMk5BoMvAtNNUXkbKu/B1sldjgBKKRP8oLAaZPW+pvZZ01qUTBOE7OZit6mjaSxG
JjbIFSNq7uqBHcUKv6JDW6onTbtgUi+kLpuOrWEJe58/FBQvxgCSjZcoAZiq70WKPm9G3TrfHrws
aWKmo2E4JMrtgy60ezrEuS42WscaiG8XqEaobeKioyW8Jv2RyuaIOXBMAq6zQJi6QN2PNIf4JNKr
8nYTFEcY/oRNv7Au/eZzDQtcjg2kyCRoTs61JP0Q5X47BCZpHbqQJt7GC7ihCiEyYyp7kNbbXGFC
l+dItpriIPnZu9N251y4ERkkTm2r61VfQgIpkHNjIpKw/Wj0N6wvTFYIW8uXZEnqL799wZ3Djjpr
0xs2+AWDwagsfrt2fbRoDCnQT7CZb4+17+3QDqwBulaxu95f56im80B0XMkG9wjFnOEIME8znL/1
Y9Yy/pCpcZeAJt0eb+OIHf2P2tKWTebFO3nh9jtXWRn/3QPAYkeyB0Ci1/dHVA1bRDTwqBXXRz8o
JhgMh74bXd4k8HyPZ8+b5mka8aw6eHZljE8LioWkuVwYVTO4K9xA9lC+du2LXzi0WxV+63zBejc6
w56HMdwZ/B3vtw4boR0ckOEDBgPjipMUIKCmO4Rz6hPVArU9RbL9s1x/9+ZFZI973tjCHjMJkVr4
cKCITkjzyfPq2Iw9uBIu12wOUJWKx61WbGtR5LJtqIC5iYDYWP2J2X/PUzPfEmkt1FbLtcGKz0X5
NJ8rQ+ER3IMC6nwGS2R/DGLufsyEjOVe9y3AvPlI28crFOksXRTCMXK7r3TvxzsDIdry/XYFEJ6m
6U9sBRpPVrWdh01/r1UQKovkAASiFlU6/xhs1lBhfDaa58hi2Sk0NH6paURurcmTCdtX/KF33ann
m+ibDS1L6rJTQ2q6tqeIgrfTy96rgADtT2ehmYb3XrAfGEBqG+D5gc+JL3hLQwPI4pb9FqgInN7W
kjHv4YPbbmvVi8pCJ1W/xOvHa83uP57HWYk7SpZijDV3lgIQETXVlg/qUMP1eg+DbGB66OyYfKTy
1t/C6U1GYWdc5fuLURQeV+FK3vNSGZ+TRPBSVK+qHcTNmZ2SKPO3oosz9pStrz1MdA/UGjySw/4g
ZWDwm4somBB1AyY2GWZzbKwgeR6NV2gSuSwh7NemRKRSDPA058G/0TvoLwyvOZM/BaE+ryOl0+la
5FNmLzISGMoPqCfzhbYxNQS2U50uwVEyG99qKVFnd5KBw9gDCAv6NGbKE9oM3fRGvYPBaDwo+Cg7
81R5/83YNsW/Z5owbJ7vXEC2hD3sHu0vIsaVg7ZUzxWv3mHfhiQq6Z2ij4mwgVqoAqRrWXnfXXF0
Z2CwZIf0U7uc2C+A0M4Gt1uiEX9rSRXf1eQSgj0a+ovJIIi/m22I1ArEA3lYSMzPVY6mSK4PjSaS
QtxPZvWI4m4h/9teE7srFfURWVygK7HTNAkoqkaiNPQDMAs0lDxkrJSr3yYkKapJ893XYYwE4y8D
dSLMJoAgcf9YXolGXZLYrzn/m4/eAFL+UxR2jHYDTbL/o9yxKEjrT2cBvjREuMaCnOLQoThzy/W2
nuyeT4nqUtA+zafinQ3eyHO7wm4zu7NLdatC1l2wOcXk1AAZsAZAsIlUg2yqXQmzzBSQc2vQ/2oI
rR4OFFAJNp18ro0TJvVN1c92mW+oRwyRfJw7kfpwEStWdDo0br6UmG697zXQSk/QertBIfXpJNvd
bAg9FEg2nNfyxVtwE5RqS55HlOVZWwO/NyCp6HdhDQOjVzUh8yhXaKMntCrSDaMACtUoyeruoEpj
WxueDZ/+gVfKA7b+oO758CObJFwuF0yjObd68FTwx9e9v8tZ0fdkHgJsVbFxD/vvRxA72VCs5Wvh
y5mjUG1m0bM5Oc395fYFM0dNxS6nmwJ3DurkZ6AUHe4R5+AMCnGDvM8YWCbhLt/KK6293lOOhGJw
BPmF0UKinO4rkxyiQYre4+ZHMIpsjAxeM8zTE0Et8Sm/IjcV1MSTyRSANTliD7jpDkJ2KXaOMcG7
UXesxMv7sOcQEDwFN0w26mMA4TEhMLU9ejvGW2lSCckNq+SAWdJcPH5B+1xJ+xAfl8RmoNfDrHpu
nfhXufopagJLr6n/xtsMY4bZaiYxOSL+5dt+rpMd3T38y35HBHgJpUSCDtlvNfc6CNI2vghqVLhB
P/MdU+jQbODPTXwWD2F4fxuhCHnH8M3K4J7vyKCU3lajxY66IsJL/JE3+g3iiDNxarSH/BJcdoYs
jfWt+Caps2ugkf9rCpLiWnxz08bNs6k+oqW+dlbFPKLGdUpws2Yw75f/u/VTWumoTmpOtDG94d+J
vB1gbVwrsNKiScXQ2fiGAafL4EikmfBEa50jkx5+EMoueU1jSsmewCOwfIDONqlz/TqR6b5KalGP
UkJr1bNLeCwnkYOHxnrnbZFZVNQXOm0WkF1T1OJMIdqR6ft+tOqDb3xr/cseOJ5BTqCEytukHhMf
dXc7vRSsJNVVRMvDwDTUY2BSdabjZIqY/2WeSaF4BUFuighQnt1NJ+Ax0sxxjqqvOuwVJzwxn74D
mc12Hp0VzAkK4bQ8Vu1HDDlJH342lFE9r91b+OIQiO4wDCBzNxy1aMlk01qDbtoXSEx7CLUN77J8
9dfMERiSdFUgMRUaL19PEaerQ8+M5jCjMQ9md9P/KqBSyd0pOJHy2M3sDF4MAdd+HBas8bJ47JyG
KKuvdGU5Ls4/jaOkpsy3nhcra15LXOICRo4DyA+Yqo+1XYVwEZSKUbIj0tmE97bE7JenvtWp1ClC
74RWQL3KYYdwqiJ8Q1FJgT9JBr6tByUfxivJ0vunAjYgfvbd0UIViomMGx9RIdFDhU/gH5om/jl9
7rq8+vrbmbl8y5Vf2Bc8xOLila5mCae5D8uvRiRfk1ypCSSDEukNqRF/w4lTxuTgtRyqStQAt3pT
OMxmrpKAmMKWmmL0rx1Co4DN6gJEVyFLB/pNU/Cw7RYCBxFejlkrl54SJhhJvp5JoVdOwJjoeNsi
GGJ4cIWdQLQkjW7DkUSFeBQWetebEFXdlxdBx92E0LUaLORDi3vhjDvJrhWjLFJz9BiJhnG3me7c
+dI/Jy/3/Myo3dS6Op5EXcSdnuuuFCx14WRiPB4TQc2tCblOMgVoRhFjK3LOA1TyTWzJfhaS/LEE
cOjQWm1oLyYW4Zt2bgxqL1sMIO1eZTV45GldhreCrxQ4meMEuScv6+IbGQvOUI4zB1nKZ4lqfKUo
Ggrn0pbXCX7UJB7PfuuMEdh1YyB7LxnhMUFsZfqp/RSMu+CSaLsqi+CShQT879HfUwWfdU7uTtPG
nHgdXJYxz/PBfBqf1wa9uSCuGgB+Pn5tGgttIMvMt55NpE86hsjnH1CrNEGfI2WGpwc2vT+W38re
ys6G+KYV8PyUKOgrNGJ22ArXChTBBsewQ8dO2QGbQz5aJoHfkJmH7B212lDsnj+9S2xADC19+upv
kVxIJvhuWpYYuWEzY1myinNI9er6CuS7g5je0R9lA3Bt5+IK8DV7QG02ArRTvfWRXa49eHQu3gLE
o/ewvMr/sKAAiSb7WqLrePmOm8Yq2EMClDTGr2K0q0nWEJfKTnvyNaKdfWKRAuxi1sDgVUv5q00f
kLi30KpFyXeXi/nuPuhjR4wGwiBf/NZzqOVlp/lLeo/yj7HLEhgYMURFRgLkwBOA1jHZS9w17FFe
e2ySsYXb1rRoXrxOlBYg+KA3Q+bsKEYbn6jwTmzHUAv3Xz6jflq7kAOXxfWhlhEDf3pNXRkey6CB
Zv9TPfEEG9NoYzIW10g03JAVBbjanPwR9qCXonldV66TgBOaPFOHfj9elsSejRuwfLy2OjfJBRtv
OEkozYDZe/2yd/dDU6yCEkFIS4JX5W3l8Hkw5ccghSB0xXT72eYVpQcpap5XVvrEeFiBxtBFiR8r
nKH4rrs0vikoxm16R9vBJZKP1HzMxlk0g9or4+DRKBXLPvtorI2zQKdIQJMXHQ/Gq84vZJSlY7QM
fGoIu86lhdFzV/PWN/yhGmoYUrl0Wzcop34UF5BLMsyDW/EiKfUZyZz5K0eYOqARzI6zNPo3a33T
5gxPbzuUwftJ0PsNktLN0WpqjxPl9usNKXLzbjcPrWz5MPVa/TiACPXqDFlFN/6pzci4oP3swh/T
3HT2UpXW684rPTVgCxTRYzqgBFRB5JSCb3/wFHkvEp5b9JWNQS1zLizBqHSAZrS8DhFfMn+xNu53
W1lWctzwtId+eSoNVEw/UXZdFWDXtoIfQHR/ip0LtADOh9bHfuS+icBT56Dynwd2BbdiQqWLupc4
L/2pV3DyOteuEhcGUZ8y0EzJ3vYu44OArpMRgNbwJtam33ur82c1fj5+DOh8NuYpykwD3RO2rMOf
GEc7RKrNE1l40nNl9mHhrIgP6EroUhS23hWcEvkdSxejV0sftIA4trFkIRMDPmqrE0wjpZIR9zVT
b/P+nyxVpMXAx+qmzqtA9Jk4y9mfLqqOBb5zKudCpxprJDVsivPrsAqGwwtzBBpJCEo+l6mAk7G9
Stugi7JY/8iAr/KWqa/XQFXeFRtnhxFKLOOMcoX02VFOrjNs2mbhRFXr8vSWRtrF9Kv0Hgy+a5To
vcsvzAlupz+oQ3QEGwko17avPn2ZBe+DCR+q5N4MDBLMdxU5Vs9qcq7XXGMt15Ilvsk7pylAvAO5
tmPdew3NapyeHZhFopWI3TYupglzeuKNyNmCQmz/jPPeQJ1jpEHpEYeElb5PfBSvHHf2UM1h7NLC
AD8r60RJl2NzK8z4JktpIVVev8jy6tIN9xpJ12fMbBZVAsjS49Q/G2/rl7A/TrN0nI6G4hcFjPce
MFlOWq+PnZmg+0xRO7dd9/nVa2ZACMHqsMAO/9512xNxY4Ltt+yVu2QCtzTyA3/ogsxVM8ukvBzh
Hz5TfR5Gfi1Q9Vz4zgtyHS8GVK/4lk0MT/djaRgNdb1YHWmKPLY87cIBEq89Wzha5L8c2lIHt5Sz
DjaO59Z6Rj5SL7FeyPOgmzDUwl+eWwSPnXGYHgYpf2+32Whzzg1NsDktPYJQ3Ocpmi33FpkaqJD+
0M3NJk+YWe7CSx5k4yfUj+EaVpbRENiRDNC0yrer3grC220gb84CiVPS2m0P0XzJfE7kuDwMYOxx
bhVhgDiJ/eSuAi43E1J80YOuWK5t+F4k4tt/gNimFs55WAMlWuibUxejTuc+R4+7k1HrcEtFt5y+
PV9kXgGtBwVeJzj20opBY0LgT15oUcLJRQazJW6gnXYMbGk6pIaNRrQaSJ3PWe807+O6+UTG1QBu
fj17hc0IIjNLtZZftWS8DRRlc0EeGz3nTbqNbkjpS/O+3WUv4zaBIhhQkW6H32A8lzBAG3lP+pyb
0D0AtDlLwfiCwsStF+aiR2dC/0Jl4F8mvk8YbPAmEL/7sGsbgimVkqP7WBftsp0wrwAAdgG5d5CX
yDf58xiSRxDKzc19zjRWh+zb5JP4AuHA1fgYJgUBuiWqa5R20UMD5pW/sK7GLJFnhiL1NbU5tvRh
ICcnltpNZ3VgUoCznlfX4P0ASPmE5iGTV0BgE1fKdlVAk/+KaP1Toy4cKrnmYZDxlW98ynistCtG
3HyHJ6lEnNzs3GTQOEIubd95YE702wt3EShJYhGxa7+rGCyjbysDUlV22BgfxrAmwIs3XonYSV1s
GIOHt49VUoisYMVNLmTM0Qm/fFw33RcxaCMrhTP6viD3+oAJWM2MjSCJN8WhGYmyOMnk+/atONiC
k9jikMKng/trhOraJ6swMpJppY+NHu9q6cb8k4S4JoDmf89bNONEZsGOeF/+i8cEluE4l6qm8cjJ
v0/Kwch+juLMyYPWd3BSgCbZnyqur4aTl3MmYibhbz0aHXOFLPxUR9gLcdHcrS9hShCNACW22O3g
WqmgfW5KVgBfavbNZykfXXyj6CjHCJwHThi4Y9wMP2KuptpUkdkU4ip9Eq7/5S3v2xyNUJ8xQuhc
V1VvHaOujaUfa5jtZuIAlrkIdMShHLtZpOM7Pn2WVRh+CuHYf3bXpRxvZzsMtbHpeiMyxXZMmbZQ
7LAWpmAV+Pw5djWO6vwXv5Qs7D/Yglt3MYqSXTbKsTqJQWXGRk6Bz6xICdoIitnZ/oec8uOptcvu
Ni5uaMxV/1jIfJcZl5EWpDuBYOfFDht2GGBd1EKR0IzjEmsweoWAa9VSqgpN9NGQfZgJqGe2wEvj
+ELPDcHWgd42ONNFogMXR/NsmLxCVOU5aVw0/cw0fwgE/X/98YpmFY93obXasr7OfEYuNH5WguJm
v70s38j3tJdKsUa12ujBpyDcERluTfJK3ny0ykNYhYYFOr0UJdPmjneDP3XrL8nDcVhdVd/2aOHd
AvNzqpIb8dcn7LnWXQMKHpFRWKbkeU1THbEWlLtrZKZJDGFg/ILeUqofr8RP9ab66Q315sWD6dfp
W9k5fb+UpNxq65Jo8P6EYgmJpIcN9msIZCzcXJa4EkkphCY9Q8zakOC6n4xxwtLpWq1LmkxNhN9h
+nhI7fxgZgh/EWR66YoPNdm9WuCuL4cN6s6uVDLwAj1OoIoH5V6EkmIKcO4kC55yuxHsSLPAVYJJ
AppI7KEG6BoHJhL3LW2Qx00+gHw/WC5XUlIDJ7jdM1URR+Ov/rRvHQIwA69DwLqV3VlHXPCvIU+J
iLhtmTpi8upMILkH7CMl7SA7QmbV3Awc42tl9E9Had/uN5uf+h0wj6V0dX/RYuXMMqZwAhVik7rS
b4LvfTothBdBEBXB7stZKvbH31NRNQBFxlUWj9NFmuMdsHUx6D0ndTbDcDKOanFngnqqdOx8L+X4
JDVc7U+SE1NlioS6PZLf0FKa65+10qEIQzHfCsMBDFoOZS5sBUxmxsJSHg0jStsgKIQkTxU0b0WV
blTSJi7KGXDAOW2sQHE9zG8Gqhag7KW3M4PMMCqRxhxHKpxvHDw4NCPW7b2e7jLGq8MTqCWvt/iN
WC24Hf+05QxWlMkTz6wK8Q4gSbjVySeTyiSX9vluD0Wla7sU2wIz3WbTw1cthURXEHgQImxlLdMw
U5qxWqc4W1PB5oCCJzciz9huv968ipHFes2rrWRfDAneQLplqJMifnRT8jOodJ/KLDaAdXBmPhFJ
AZpSz0O/EiP77UsdYeUT1RHFYGKciTfR2NJypZIlr+JDQuqCX8ddwuDSpM3jVZFF2N3y/jXHF0jE
QE2H15+8dL4YXFph8w+GzQbbOixjVS0DjtE2qmE9muhwHsNgdq4JmQIHz5e3O649gehszmgp3FpO
AbqqK7qClIvrhEAYnqe14ClSDN6QzQDmZJ5u8yyfMRYdaZTaIjNvuV8N+51TbTchKRe32wu99RF5
Bpd7qlmxwmvvPeTO8CwczWTFQ4ZHa4oB8OaQXk6VEUHacUZ0c1cxw6AOdvLShmI5s3x5XHmI+Cpw
cts9Ssg6zXtAUySOAutguqWlwkmJ6m8Zx0rlKZA5nFBI6XvxzKTzYUI70Kn9qkOCQb/v2c0Xfo1/
NHL4CZIGKYD4yFbiF3gRiFxW3Q6lvfuxFfOgXSug3+TZJjJPfTpgJ1yrg5yKdzi6gvMmg8lNGHTI
DMKQozfSHqkK4s1Nhsg9+O3Caj2B+qDz8BQWKk1RPyiR1EyY8wDr6rFT5/ZHIpuiFSowvb51DDhA
KSEj/ibNxNdPU32eKV9pMbUQEFdY0Rk8tyZReqguByB/3kiSdztKSGtIELBz5mEu8s4QF+M4GyUe
HdDvTDO+1zUh6FNPxMIyBcB6APlCG/pvvl9rCfwkDwB1+7hQn9ZQc34Z0HClnUaEQmpXjJZHJHMg
FG7ub6j+7/a3EJyTQIc3oSmm/vXuYVCWqLC4phYx+hrvOwd2jG0wkFO3e/xFdogfdnIadeRndMD4
LSSxk9ECcRTGLvIMkTqsBoQd10eeNp356cRDPZGrWjZa2P9d8bEjWld3FYVOVUa8FDNDsHtB+n0x
be/a52fwIYPq7KUYi2lnFTLpJbS5BgKjijPK5ggAKnxXZlATIDhEohEU0ESb8Q4ju59oRGtL0rRT
l9dBjSu1xVd58edbN9aiNowr1jNpCSZIn/UKcXuc9tcQ5pW6qfmnpqh3iwi8A797fX1fkNpMf5oc
ZQmF62w0hvy9hr0P3nkHbblUn635+BNbc2ZifApoy8Ytd0wKNZmJxqVBDX5Had63JSCNkHPbu4HC
qKnFVpT4zE3IMNawauyK95O+0Qcm9BAhwjaK7g4m250QdPu0LjgMBcFfI/CakmROfnoma7cNNq8s
v4fe4RZDKRKwRsOk7lo/v+H/kQROmwPKtEdqGtXNmpUiZZa/Wp2LsCdRinYO3iR5EKXmk866QBrG
yA3bTbTaZlRQoy7QHj1kkYSma9p09/c6ZS4BqbyRY8qXdx/4xNFmaxuJJvZ5DzP9GAQgGuL251s4
KcOpyUCQ9v26Kz+do9PG43SkJpObXqCeMN9DmUeM3ZOZd9FqG/CWSgjHDC8EYS/tyJJqZ04gNPHy
fZk80ElvD5115rj0JqrH++Y4YXZ8x7zzynXO/TP0tpQpsqWTWx9lwA9FbzAY7//kBoHVMHqkgTwJ
WoMcdw6IiBEUvvrouoTc1FhSWU6nhP49zpzY4IzcewKZwp8M0h5NTVqOHkSb+YaMs2QpBOoaAHgL
xuwMCENLg8VbZatY6HM4J9vIoW9FcW6O83xvzG641m3LgmaBRB4lJdMTTbnW6dA3j+sQedbWdy2O
ePU8+UNpSgajh0lEbtkX97w5YdNA3TKULTkeFR/+PynyL6GvVYJlQctx1fGNnUkG0i52grdg82AX
VrFoiQM3oFm5DBe4xJiz+q1ALsHI9iMAvAXCJGReoTUi8XDeaznFB15vuSUHRMO5lgzvxdu5wb5a
h4ds/V6PLppSaEg9MmD/0Tu0J+vsxsBPGFGRjAuaIsdLev1lRJt/kYe0+zW6WW1NYVUTYbJVqDAQ
VpTov3cm8n+jPAQBxyNiYX3QPINyA6+aSfcax0cnyO/Vw0Xw62IpqR+jUV+XkxTKHm7EAMUNcO1s
hAyz4tkd6dDNZu93/sYDNmEwJbK7xbAzJ3bC08ANYI6oWVt9s6W/0JQdB74yClSzNpfT4KaZMGVS
PHEUeJXIwNo5+YzyjF/b+BuQSg2uiTBQCySUFLZo1BQOb09t17VIE75cN5b7hIlTj13f6XpIBkoe
pQKuEwRdInAz3TH8eypbAC/Z7Od3Vbq9DeQzR2ux2k4C1Eq/E8yCu809qze/rIsXdllLzw9HWD06
2GtUxxvZeDlvRLHPdlKUmV/h7p/KCzGn0HS/h37jVwfLJqSCS/6LcGUemaFEJMbu8bXUrgLf1a06
LcWxO5w9g8YrNgx9QwDi2YyLXwWQARVtO5DwDGWCFqRqNIdKe2uRZ00DJYIhDVwgVxZgjvFjSJKZ
rKgUbrTtfsrXTba1KG16QOuJAWpni7q266AMJini4kEZm0K7JS/63vLZnt7n2/hgjlCz/pBJ49cq
0k7lOgdqE6UWqhgOnzzWSM9LpTVJD+paXEAGbOdCyikFExqn/lTPWSEQkiNpMRTv/rjiHK04hliL
0AAXi3Gphuekiipa3BX7TR08G9lM/+Ptr0vL4yF7qJn68I3ULK2SQsND6PJexFtXlWNbcSon39Ru
5R+pgMQATBHxn0XmqJrQVSfaJHS4480e52DifoxV5K0o/DOgzRXirZHDVFNuiIGhBsxQR2g/Vb99
HJLkh5R4RTctqg224wo32yuHgoLngZ5wNIKcB3KxLXwI+tFimIIQiFZNv3tjtV8cKK6HeUlgLxeO
81Bw8A51v9w449ZXdO9ObjuWljAo8e/esdpoLy6KHenlXrYRSF3oXlO8p1cLhek74NBOXbE8rBJZ
PEZqM3kQaJrTTDuwEhV/s3s5nSsNz0cNuyaqhOc1UwztFbmZPVXGRN7ijqZMvPGeNnA2zvCfRGBy
9lPRHraK/9tjr9QsAL+S4iqjR1M93/T0L6TML4KRPX3S5bT6+/YvyQyr+LySVQJnyi2JQzxXMBn2
7MCHrrTavnkjOt0rwGuIh57Ht3/4Ako8MKesJ+PngpOCx9o3KRvV6dAiuziuf91q9lO5b+Hzm9Gl
a9KEHn35YMS+/PtvCUsltyI1CiAX3pMp5uhU4YH/CKB357Jc+9OrGigq89I9bV5KMbQS4aU6V3Br
20djzRdRUrJVOwmrWpz0Naex8tyZTYbnvl7oJKtgNJ3e4aQlLtJzSYn3D9+yQQF/pG/5IXqEzSJo
bbB+r03goIH0CLrYvVpRDt/CvCF2CdLKUgNamteTv86hbm5K8MfQq+paFOlU5+77NPWgP9/iXwqV
DdNyc845+a1RgXvOCGQliwERVb7y5nIT2AoMIrDKvq4h1wLX2UOPu/BFNsTKxcCLT3khJU1rbfxr
mAj2zWpX/6XDwQPQjESLapLWFgIcaWzADyiYCcEVNw8NtH49te2Wydnz1trdE92Pj5h9sKrRvkVl
07cWPh/e6DR8C6sgkz7WKaVLOaeiGYH3gHDit2ESSnMnOY4VRFkfryj8Bnp9B64sc1qzbeEXiz5D
MuBJ8lppd9FFxZ+P+vCfE6mtkxY/msjVif9hKNO5pYg/VaGNHDEOmKW1z8nn+oCi8go1lpE+x4W1
X3DS2JlRLgHamuHpDf4RIthPkuvU/IpovAI5Al5hxX8M628dgKWwu8Gegel+WuSHyIFv+bIPYaQk
+A/eRtzUaN8JeQ5oR5eH82hSESwfeWhzJSEPOKIxK54qzkRgbhy4neVsUtCmw4CifT5z7L7PwIiw
1eGP5Kr7iBTmY66YY1YVAPUnk9V7S4urANXjOqmXsJKbG5aDCDP15dy3rowu1tmrxyjYqACYYvMN
44VEX9VL3aeYtFlkXGJMKJaxXgGbCC4H/q4ykhyuwQaITcN1WT7L1JQoAv7sFjJ8vNUelEiNQBx2
+V8DWph8boZx/Wz4/YePWKVaf2w1XausE0zwXN8KNrdgMArzZsmkJ26M1CUEPSn7uqH8nejRaMas
NsMmdBTh4YgrBXow4duFPsRKaxVQb4cP5buXSVxt8Yg2Rb+NDWCizT9UicISpNTxl3NkZiacr6OG
8jNN7+fEE1EuxdU9y/W71e96FP78sjpxXTbcN72BBGsuZFl9zBD3ueJuv1VMkGghsQjc32drdIul
aJ/DyDCiW/O9N6D1xdw8IfqxkT1Zep/3Zfke9KDNHMzKmB3X/4XIExZ1GvVnKWNIR6rMPu7avOHm
DiKtFHkyyMPWXRNPBdHnpd26yA/2s0/9QNDvY4r3tw+N3ds14a94h7B+ooZ005ftJ3D79Cyj1S0g
uPeRRfVXNu2zhHDcrKRXrNIc6UR8dLUwiQJXYgeti5t5IDuh5pEwaKIbQBA+1m5mI61xSmthB9XU
OjaIpLWysnWZ/7bUKzfYigu7SMsSw22Ynbx75V1DOHC9vJgsv7vyN1fkP6R4Hs2ftb+VlrJqzofl
z5BFVmx8eAtJ/UIJ1V085yxU54peHKdn+vKcCwnmaiIyiaBlMHOrqZRffKptN0Rz+SKHA2NhtYZy
8j8fh800kX1GE/e/+Vm2dVrt+b06tYQjg2sUzUiitsPzp5UKVdqUdaa+E/rtjmm+bC1dg5p+9WO1
HGgVDB+OhGKua2Z8aLjpQRx7jIrMJ84ihq45q3zeKOlQ/75fXv69k88CqAytTas18e12iyRskWGA
xin7IOudtKIKMO7r3IVkiSkcPWhdhBBn6BA4S38Ao5TIjEFUF1O13y6mO2ZXVo6eUQuv74oTSwnJ
sCGFpxHpt8Lhdx9lIhl5ylfRPlq/2WG6sSIU17s+ngqIApwp9OJMMQtczYtw0TKQbno+jujJcFMQ
w/f/uCcq9CIYrThymbF2P+5rcTYuGUG/pNdt/F9ltJYjEZuaDvbBTyWPZDoH8jwenyRJnb9/X4Y6
WoYnDsYW8Hvf5/0ApfBelEk4hQzHIF/fBTpGwzuItcjtqnY7rpwyGYB/hL9PZME8fC54zp6Ty5s1
2smK4plUHprNQMjsk3/KcC7pynqYexCjpFGxT3kke2ZGhR5DQNtCGsgXSQmLPb7le0utIfJFwdld
d2mn3es5ybvOXeT2WP8v4quuMRn0roGLkXC0VgQhDr6hO+Hl7T/v1QOqfqHUx3HYulvCZL8NXFDA
ISgVTAyghlGcEhdVTi4qMeBPpz9rf22FOUBepDNAgTVw0g7kx2kIia7j4blbeuVqZtcSMJpaf3vU
f1jfkRFpYSxU6r//Jk+R30UMEPrz0SWSjq4n3yQ7KtdI7U4PD6sHJTNsFxj6X830E0qX2Vg6isG9
dk6f0PRDJh7tCkC7adObGkIvOIZlH78znMrrRlNBuA6kln8+ag+fJXq0Zpkpao9aybcKqcjb6ZGz
RONkD35Kwn2m9vArX+qJhRGLmDa/pvqJof/5mnI2qvK1ZMauSHjkGlCeLBOHZH3U6D575hXYnkrq
WhAzn7p3iA5+DGw3b4SV9S3LCXfnNSZ4Hi+iOUoAU5qJhkM0duF66sb4ba2/tzWCu2cZS7pluIDT
24p1VnEg9TrbKXOQ1mzPVpg04dZLQ2K+shhUejLgSfy9iNvXXS/SSmXFazm2DPF6JNgVX+V6fecN
5DFLPkI/VpKtvFvY3iL+/bUsmwoz0BQ3DYAOeQ6KJm6tCWjC7tbbxZjYUII8h68xcTr3uy/GtaF/
UxlDD+xgmogwsbDKnlFaL2tqctwv1ZKanxjyf/lvoEYf8O9BdJR3zSwdO8mTBl4IB/IDVJk0Wh66
soKrlF9AXxta+ut3512OiU3gEbg9cdb16RVUY+mCLX0CPPdaXtQ3VeRGO+AItpBpJB+zf4VD7l0D
xIO7AE3J/TCQ3U7Vrl26euS2nbvQE2HMjwLy9ARM+MM0fWZkHqTZg/N8lWVoGxdxvvGtb22sdt9s
lSSlzF/keAxxa0Vz13QEyzKUCv0rwM7skrU6cknw2KWwqbC3Luwsa1eKCwwo3/g7wTQoIGw2uJec
Q5QFCWo/0fvf7GUa//mrQY1MobWHfpP8KkXcOCNJeUnYVrh2cPnJW7tixB0aM86GesPUGDuxIKR+
aJ29/z+W90xODLxpYb8o+t5O2CZe0zyT4tSTL1AlMrrxNLo/ZjWVR1V0zCRcEFekboSpiKIUw4Mz
Ss4gBE4Wyxg72nDpVxn0gBRCjRxI5E/vAuNyrUz+CopKbO8+VaXRgGSUh28WnStQ5eLECwcUobMQ
5nnhoZa256rxQPUg8F7k03D6jSeCb39DBixVanW0ooF4ugousaWRw9HzR+BeQ3bJLRO3J7J5d6N9
MsaKeonFNeZ+xQqBH/Pwls9QW51R+8J8nKi3/fp/BPwQ+NH6xudQ+UTxb0Bm2EFzvm6BBOyxTPVr
K90MtZ+wm1PWxjdHa0iInc3+pkv2mNkjxI5pABBXMLm1R9q3FMFkGa+xNepRgRc6+Y9cbqQpEGx0
i0ZHUag3RdtgPNwYkMhMENgpOe2mzx8db+PWV0Yq7GrCDB0+6RZ9+QwHKG5u858xIK8GQDYQkZ25
wlinz6No80U9cNwTP9Id6p3CqynOlXGlrvs38GKL9Kwqt6vF9E3g6u9Tdp9g50jr4lIIS7LN/jJ8
5eo4sL15mGS6h12n3g8QOor1qrXMIWjmp8RKDH9Cv9/9pnrsJA7SmRBKllPEPbROOsqK4NPkP7On
Vg+yvxYipN5qBH0Ppbf7m0kTnz1GUWC2jmeqDuiv83G8FwFQ1r9S6bUU7zSr02hNATRcKX5GKpDo
pEB6HWDl9QGT8ub3ShP9u9ePzrfxI4nZJc9gByl+V5xRGDTcVvLoL3yYC+9yQK9+R0vOMU7oF7Lx
om+ze54rscCiWLw6CV9Noqt1of5ShIbSrCBzLjk0vheEvZnWKRIt0sv5Md+oZrhWzXkrlg9BJtrP
aYsfLfJpGEO4sZckpYqosv/Eo6nthzKvOk3QGToAvb64qD15JcW292pp29Fr6d5nhuEZ8aHoUQek
ruTOqezZoiNp4IyqxnITPQ7wPxTeKdG29kWqFBFpkHIRdY2q3R3dHN3AB2qGwV25K8mnc2yYJ0Ne
NDBx8WaSn8/Xm9yjWPfVbKAG17tF1zUM5X1WFqfcTYG64gOts19lxpolkNpusCe4WOwtKtNkqSlM
yYxXo+QiAyv7xe+zuk/S2DxxetlIM8Bjx1oKvaRNFy1rb6k8LM466q36QTD9nF5ns9Lhzaqcx8eb
4YfhEW68QdXVpgnl24WegDdJWbAgGSEvIINwHc1Nhkhu0k0J6iJrNjf8mc6CG2yLkxXUzr7ML9oL
p0FCiwKt8CEKUVu9/RgXB/4PNTZrdvLIuA5FgdkgcNudQ2dtGsh8cU6t9bGT9SlzgkZde84fU5NC
HJ8qHEAfo7mREy8d73zGETdV6vdM08RbAHvtDyR7ZLO/dI3ct5/LkM0qmgiQop8G3Nff0j/GdPMD
u7hXSSWknzv1koyPIikZCCkRe29+fWsfaKz6HQ7lauATkRnYKyw3k7famP4oTMvkXvSHHd4OT8k/
5FGrREeLEAV0bEZOStXjImjDHfdICzEUmUvqOi0fZ4tP9ViXOFNFj5OTGKL178qFWb1xWYHQfqA+
jDKQ2v3YZmPoFnrmccRrJN/zIcK8tmmw6tu2WPrbNox5+pVd99bHFiNoDQuBE/sGL8kER1lXYQfc
lBSy9fXeaOH1XIcXQrx0/CnGVgk8UjdikuLnC/Urg77bT9AzP51BXmRM+nX5dqihISTrsUtSV5Ao
kSdRe8Qf/TxQOyXgrSUirrbq7xgiHlej2Kw8bIl1is+6Jci6BPUDBF0xNLHU7EvSvzNsyRn9KaTn
u/D5qyJ5eciZB1Dby2ZP2MgCiJn9eMW+khkleFwb1O4Xgxmqe3WEvnTI6p+RP9U3Qfc8tu5GOTQB
eI2UIwNSU+dtHtgSdyUAhxEDUpE6nNPrLO0Yp0WRvKLmIPCJWx4yNa0iZp5yGJrfkQpqrZy15II8
qG3hdR7GFj0hObk8VEd2Fky5FLIfXx6STUFxtIxAGW+IBLai4pqPixOZ8VNI6Df2tYtq4tVPABcp
TP8bXNBuaV4KWuaCcXjf9Qwt1/pluGD2I+wT2SgQ2nEVXq49qVXmGVUa3PPfpWChtuA2ohvliEiM
JrbWk1UqSflYTWcWk6gQZFfzQvuPoLlzEs7kbQiObIyzBOfu9IJZS8inIpOL1eNAAhzEHgp18Rag
2P72/ftlhoOFTYRta8L43t4Mk4UZwCQEAlDnyX2iRv/64GqDefyZZGWzfjazZHGMZAikXzI8B8qt
j3g8DsgvHyvVt2GaaDznE0IiNx+4LHLcv0uA3VT/ap/7f58KuyEY+yGsuJ9dtqeGzZzRmiXGTsEg
CeX6g8y2YbVCHmJuINYSVMroFGmg7cRWyYwS8U1+6RtboYxHHnTBSVejmvswrq+b2zmHntKmn/8m
Jba/0l7aDj+cIzhhKtX7bCCcBsgUA1R9qCL57c38xowHENmVVXshLHUBzQZjz6mdvwgXOG7vt2nH
MOaoqR0aK+a1vqHBj3cOdyL4cd6kjzE55gc5wWvDZhR0E5jKvPf+4JcOYQfF8hZS016EzRELoGod
kizoC+HG6B70lUzyQ26KicxxGXNJRg6tMGQ7uHfE+xMq9ZJDmdJ396BubtKInQcegEetkH7ziPES
kZwnXLG0t49yzJ6X3O6PWdwbBodeHsv/Qo6lbW3zPsQ6UDgCAWyJgLy2fI48d7hynayYhye1b9Vy
iOr1rVPPS8xTnr/MfkZmU4e1rqewO7lBnwk5yBDWlJSH74cKDeYqf8B95A2r6sw0/2k6ZTY0mjJA
xBoQLtr5k4mJxIok2RSUlLOvRyfN78ZILdLANLVhNgGb6Y6IVGigXn0Wr4T5tM/h43nVrTz7qkYe
rwtAiVJcfMrOIkB9CTYbvK4PXoJdG1XEn5MU0rOW5M1ImSR+k/JZWTPD+vbLqHj2Q05ciYIfDQL3
fZk5AGpjnMrDS8bFowj2l0r0y0ZslqqbOQdy7L1Xn9hwQbn6jGVK8Jgb6qoxYdj/CRpsVfaYRakO
werjNp8Hr8Tv6nynPUA1/rHlsIDEVaXNE94ObbBjuWUJEihE7Re1Pxn2nVJG0U3EWY5E4te+aL0j
vkaU78TnZhI5t2HeaOwGS5ucq13MiYkBjH1P2eAqhA0x9gHEMt6rk2RQKRwFf/J3byTGKO+g/Eg8
oAxOuKso+ZS5UiR8nQMcvZhia/zgkuT9277dOO3zlt5Z3GLmqKb+iZ8feJpQvRNgmhEN4KlQQQ0f
tMeM6Mt3vsP6YYRmUCETIZRXKHo1k0a2RkXGzHoSvOPYVH79OWvBFSEXNq1CV96L9mlUVfgEqbUo
ts5Ib7Y7rzeSXQdNtE21EvHrgidJAUQDwiR0j4rFwOELfqOYGrd9gmC5fZOAbusASAAgZvdUl/w2
avmp4zymj0GYR0IUnup//Nj41z7UeOi5DDyG93fqQQavuzIjEMez26QwW4OANAHKRHcLqQ+2OiMn
Z1so3qkzBJP4AwsjkJBDoKwhnbPlySwxaLPVI/Zl7b0VPCVxfCgvm5AdCyzq0kI9Oswxo392avf2
G8EZIY18zRhEbEYV2Tzjtm0FbIQGqTnnvfKRHQ7W+nHDRx/ALACgpYirhcoJh8Z6Ub1+u/YG9j0w
kLnbAHZIAi1V5At8vxNCEY2xRAGVDhIKApKWAEOM0RvH3reF6f7jxYmydPB2RSi4BXCdQr8+osqh
rKa7ItF7ao2zBhkblgTXe29Un/btMD0/+eEBnc75XMtamNQ5HKxBr/OVh+Qe0JY2vF9xKIKapZZZ
xkki9QrnRBgVjhTRCci6k5qQ5dFxk00K/S2VBO7eWXCda2xuaNBc23BbCmQ2NUfjneK8WfuPtg2J
kjrk9NzgqjC5uCzxaPF3IwPccC1smS0E6z9f2km+tWjs7lQtKXh4IMF8t1nmoOZfA2zmsi5x5Vf4
ac5GJ2d2Z1AZ0H0cSmJPzhekpSE6WdUJlOFqpMJrtIXdeR0wiSnbfbjb4ACInDvrcpfuvvn2qy2s
qELaZybYI4OO76GA29sbdwca8epduW+TbZcBg2kzQdLOaA8MdpY3rippSa3bcvE4/Kk6KF8bE+Ii
TxS4D7uufgJMIO2tcBFnOEKk/r4eTQh/9AraLNnWJuID4YbLJwfCOG7SdOrf6iU/6ma1pI9+8mCj
+5vBND8cq68PSbdjkSsMFd2FOTwE16NgMROHaZGkLgNThX94FW52Tnd+tfbFw9ZD5LMnYuv6ECBe
H9QzTfhao6Rhh+N0c56uJm51YYLams9LE4UMgu7fTfgx32yC5J3582G3lB1YYEoj58YaVJfu87vV
g/v8P2lUEnFCsnYuf12nX1a+BvqBSauq9/lVGxsS01NgLAWcnLpG9GxENTuIbzxisRCfFkkeo51Z
JF+XVlPQ9oX2U9lDfkfzP93SIzOOX3DXlRsESV2vux5217L+j/0LgGmFlsuBd7WKOLTzR5tbEwaN
reHLAxg3U4E83TLXGFMjbtwXInF4WSg+hUqyV6sX0VPS2jh3SMMSexG4tXZSxEbC68vZhGfGD6/V
evH9i2KTxZlZecrh9yyG1oCqySQfun+7e+5qpM6eFeqkfpVlistiJ6ZpMBP8eCu8KojaolM9Gfdr
KKVz4vzcwIQMg+j495mysX7/7K9l5hUWuO87SOR8CPLUPeEQ2v6123ZDFfqgXYDw+v0Cz7hAF91Z
vn0KMY+AhIyKXFNpb5AyEyFkB5Zc4aYh6+HRn9fhajLMCoL5Buba9sy5nBN+49ZPmk/vOYnf8r6P
8KLD0mMVLUzAdT2PYy/OUrvyrPoBOXi6VvqUW6N2UphNlM4jhO3/IK4Hy1PxUtdxa4Q4ORSVyRbi
ztq1HiAaJXhakSR/+qzs5oQyOIuo20PZr1iP6kdXnJhokx+lqLIiLLHeH+xqRRsmOMARIu1OZzuN
3WDQ03Vtkd6p2xL2zkvP3Vxke3enLWc4fVSNdR4h+NKBlYF+Tgz3U4mcVND3FzFcjmFN81eoT7uc
Oox0S+Q61VQ62RK8Wxy2KdxBmTqSk3Wm/NGvxVLHjhjAfDO4WQomxAM0ooZdbyw20dW6YU0ZcV3h
ZOsFYUfbuI5n1zpoCyl3iTYHZY+frOtih6AKVOBddyq3ggmZCAsC0PITk9vpPvOoqPlTwT9PtAto
raP8nGH4Jy5BWKUVxTHZf8RtNqtrk8rBJaAaWE0uRDHnOxr6ykIw9sAsFYHXh4dzdTb2V63P9GXH
xpixOdK5PKI0r9pYCMnEPCXc3yfty3NoCgENGWv5R9kGA4g7SRCUzEipjyC7itKdU9dTFuUxdthE
rFmE3yrQthbB7iP5JI2ji4H2fsCojwhOQKlI48l5vJu1GRuJRp4Xj7DjKVTUD0CH0schnR0htyJV
ObMvJnafwig+kaW9UAAH3GGHWCs889YjFQ652a23E3c+atNOQ/fnqvZ1xtCysV1lXdINplRLc5li
iQHYCrFBxcpRJSZAAUL0dIjD5eE6S9FfQXPDBhN917oGPZCTIBLZnBrfcCiaHQwmwvKu6SSlBtQF
CUznlpEGQEXwOkH7IgA0Ivu6yDw7Tpbe+WODTb+TLQ4t3LM8sfEpwYdeSYSrWQW5ETn+I2F91Ttl
QIJ3msXW26Uzc5DWAaw1NB29MerNCYLGoGaIDiL29z3B/cKaKGl5gBfyfeZD4KYLRgVhA+NUjxC/
oG2ldwF8Sg00ivmf+jHX/paqzKnb/EEXZwvSWpVyGAWUo7LLfomBsZDNv0zAg2AuFgqIerKSVCaD
1mueDmFrp4HzkAEuiiO07dDkMD4xeU1zS9R8JTcmxNf46xrd3AlDejBc+0PG7cuGUVEGeMlwIYnz
V9odaCL0MJAfzan2TPEsd0duPav6FWIZEwY7DEl1vjEnqUPyi9MHkZMfHECoUv42THNGnOpS8R9o
NHQ6E1qB65d+Z8P1yyqatMKWh2rdmiBOyNLT89OfDiaRIwR7M1yrlxP2D6j2RjYDwLZ7mjue899H
4L9z24PU3GVR9thjFnfDRFTmqo2g2Ryfb8azMFxvEg/7SX8eqoPH5qb9fsImNE1fmrQknELtjia9
ZcOx9tDpAuSvhPM1dK5qiF0xEOyrtR2KEQ6JhbetReYpQQltbtLeZwzGux2dPz0shv/8+bLDGqWy
6nRXDQ32AGpfmaHAndjyxCT+bAvBCYR/0S3mk1TekBmNEyU1RTAZgVIJPsTKa2zcT1AF+9f3ce+I
na4nnaPfpFhXtq8NkJAiO8Qu8ExbX2fq9Uh/l88Ov3pKJUhcZn9nnTDwWegh9ZjqkM4W1wkxxg5t
1pcegwnFaQl1Kz3pcEQwWaMu8QqCEnOtWNB1hYPaCdMeeDg5ObPY9jFF25nrh0sQ98a8rYEi0JGk
TonCGKZr5h0hj1sdwwOKjkMNUE7j2tVGI3P72IfGKQgW6SdA3mSCF7Q3iF7tv4nOc0FNqdIuKBU+
rlNXSMicpuM+FT/Jxo5mI5W4iX39RXq81NXTF+Rec7qyQmxqRy+LBtJ8B5ZjXlxWfRKTT6WDkHyj
MZfe1AJttU0zN0rl/RNGCHr/2revtDfXNg4tMvShRwN8VVYy5N2J4Ld72Q2ziwNPsOkGieYFBLbJ
M2/JC0wvDhqX1YNXCBuHJfaRKM3j38jAqJFlI55tIv4PoYY/XIYf1sPtdDY+qGxsEoZFOWvr0Etl
m9L8NJjvNYC78eGJSWPIXG2zDw7WSy1/eu5kXFGRlMWvdyT212ORC9HBlKQxKbCKqGk7tq8LYUVT
9I+dWPTKLkiHXCPCudzYbj8lrJht9AU+FUI+GD/FYJqV24Fr+4YtrAG6gUrZcMffWPlB+B03iyZg
jaZKbscVFinbI/3BqN/8wTsOmc5iTKYqknqrAyBBIjQhIWmStOcJDruzkfPn7qD4fB/f0BVA8hWT
bqVKTtVpL63PTPoMmTh/5K6Wfz3KWFs/32ihvlmxg4TQ9+bO+UrlXog8dRxva1TZ+CG3zgyCyojI
JFoipw8ndsemsO5o5LvZfXx4gBHppB5rmhnTWP8ZStDf+R4qskvfYzgmSK3FdLFTi39Cou5So52l
vaClG0MS058bCaOt8HRHdxkL/1XJjm1jdMGxE7Cbzt6u2du7Q/axmVOX/n0XW0S9y/Sv1goxlBfg
4J04WqhSkCis5dznWjr4prY+I9IpzmjEogFg/wbilO1dlcV9QM7m2xvtCkZsjBMw/Nic5/F4S4Iz
L4GDyBPd1lPQJKrbEdKfx3F0Vo/yuDH/ZAWTLAbTNGSg2Buh9yPJ7gedo1o6ikNKfZKlZWxaT+26
ORoMF2CbUwn8wb1ReVg+m7fGpuXaBLR08pbht3aNYXgblsUZkHJ3OB+G4KeUzji+OOdvlF7729UP
DsE9fwow/U7ecuCyUvHFuxiJ8itEs4IIscO+OcCBqOQMozbax14+f8XJFXx88W5YKRl5biJeWM06
l/+GvHZp7IWnDqUSSpAkzS9tOOw9esSGYeKQhI9ujVibvmwaVp7s375gz1mCXdUQTwic+Ia8hY3X
HWTuZg4ktzOMbTCjIHx6f3T41VyoWSE7lY5fwEEvT5q+bvuW/+JWLWvJrkm3xB3z988naeCPYoLs
5yW4HydIlMkNDus/Io6ewKlYKkmdHyozW9BroIKnwwSpMjeL9LRJu0n4dAGET0AFMVaOtcLl5fH4
xU6CGelyCI1C+bR8b965FwH+B+qBrak2VwUSf12wRDjgTfUx72YlY6QY6qnL80LuNkx3lkA8+bGX
wt61Bu2NtsxJTcjscZSf4ALXMbOnMcyAaTjxoS5EQ9fpAUDrzBP5orDwSG4lcxx4vHVXPjkdq/4K
zVFq3PxgBx23FfFBbwhaYXXdJzmTcO1t9sqc5iJxhweDe3oIk3eeWjZkqMSBNu4n6HMcZekB+qRg
STXjj1z994R/i7lPh2iLzsoEo19wjy5+EtO2VFwF3tiXOeieK07wHAQG8yl71+c+L7XzfvYn/6Zu
zaQt5C4z6oq26XWSqBkRuYTFuC/0G/099vrQoaYgY+1VpVv9vn+/i+VZ5BgXyHDapElmpphhNWw3
Ctpf8f4qdUs4bp5uc9cOP5QCq+xDeGkDQbZ3kDrimKMmYe1nRWM1FNhR9p+YzMW4NVVEuZFbwFLR
wOi52NJ5qCuSUJTDbxuEJl4guDg3953xKG67cmMKuUlPs7x2STMGwaP4RxTHqsBcAfA5ZUO4R3z9
buxesH2d+hzGdEGfMk5eI6DGkZi3WTuGa1qt7K3UwyezQJyPbPZW8aja2fRt1MDUMNEZ6AA6adLv
PQQ+ZY+32aI4oUK/ImDfHbOu/gNwVniwK9xnxUe8iqQcmxOaScsiodiSgKmHKc+6EW8J6w/miTBT
6F9+6qt+Aw0jcFqTbBF4ET8TfMW3dDful3TTTLGxZsnBMbUW19KwC3+mhBlsCOK/dggjfmcXLXP4
Uv6Hek8GgUqk8N/AAVBYtklKJsC8IMj8L3SWZk5D2lCej0gnGPCCPTyrkqTl5y0KXjXQzNWeGdvI
6pPFFD2yMqonqNWW+FqIlqy+k9JhDbnnjh4F6iLhODJzLtjQPmXxV62/oBd80DmjzfwgS2b4ZP6y
+mvve+gRJ9n//pmmIyHwVGJIvB999LeKmfqIUtgUkowO2m3vLLa1mpPzXSBNZ7tT52qGKwSiTaKi
jVgpAj0rY0FPkDiiRiq2259OpaE9/MweyvlTE2BJxTbxcz3Q7jeppzDDZqU4HX/CXreFc521HHsu
79VinYTJcBxQi8lzFhuXJVBI+PfsQUhqNk1HdY5vHxmfn0tnJNa+3N97bTXKvvtyySQS8nYPEztN
O/gG2pbRO72pRuYg5l6hqkG+O6qhdyoKulYfsX4C9Lm1gkxPVQTNdvjpmG+3A9U5OsPf85kT4ClZ
7aniaKMprmUr+N6G8gQRphWEiosQBfML+hCy0HjHhI5sfRxmhfQfuUrimt5r5EcktoTv5fsDHqMG
fcI/Qeni7SpK/8Gt12vZEYDtYNkiIXs+FjPd/9vbUgmowx94mfOG6Nb9Mo8MGgr/7fYa8cuJTto3
SeDIuj6mPnoFw/98D52tFdFCBXmHgGcNGSFRxLvVad95/1LvxYLPf3mpNNZlGIdgB9SRhqJ69E60
D64BSjlsQyxUEy5nUawBRUN+vmpV/1wOdtmk4GG1o58VnZ1reH++pvRIMGa9Ph+Fvt74rL4/9TYO
rz+iAHJJMP5Jf3mrrPYMs40ljy50tD9Sqz0Us9jtAaNDg7K3mLKw+gL7s04o1jDKT6kBhDybB2QE
g81LqlPv+f6VeT2uECbf4I03GGEOaRbUgWQf4qM5W8VDCN81KMU9ETbx3eGCXZojnjzSaNPNjJg+
Bvn+8c2WCTHSpeZcGEFyU1HDdkYc5JQGYzqJdh4kRSqXnL2KF63MeUzOhKW0FFm0MJrgQvhFVYHi
PxvTx4lNJCKKP53qa1BTDLEPT3ERRrFDvVQaAAtW44IkB3/cnsksoxB8iIB5sXEIST1h3yeU7Ug1
mN7fQ0wmcy2S7yU7zPHbLvu99nSxP/0263xcsdAcb9I+GHmlBzUQ79KsseY3kAAwjW8iQgCrWD0R
+pOU43TbBOBjKoobUb+XTsCgmeZ12GO7u45n1zUPOtKBBiKkyitMyLF6/ge564K8tZ/Vm7ChNzQ/
42dU0+FSl2qDsH4dhNfTUd4/lE0V8DZ/3YCXa9A1iajQAqyHVZv2EOwLhnm0xVR59Cxh5qu6wiHM
M2uYPjfckar3tlKyvMHlxDjhvgpJtOHvSG8ONKNBb1aUUFIIuxKPGsj9D+xG2BJ3druo9JaKRqbh
6wK7mv2v9GeVFNPAyL1ZkZopw8OLmrybAN/ooXV9bcY3iiJ/DXrTvPmZ07UwgNkQXiuxWGWpTd6Q
1m5fuWNJ9czlFB0ZHEkKzSGaCKlfMl4DpKg9mVZZ0SMFtI7XlmH+KFqOGvsA4cq57avi28U7Bfze
25QXeKs3SH6B0dOAZf+aZwFVdcuQLceGU2g7w1tSZIGb8aWUEupVTc6WOVjnzfLb0/4ddFRA9tKF
m707EFwVeR39u09c5EpYg5vEsdhp8nXqXetF2TnNYG70CAVoR2JyXdeljsLhxgFdVRubAv3Jokqe
W28bDZuMCQ/o5dN6/iXDNie0T7eh0YRROZ+W0swdfsMhv2YCTXUxH7uGtynRdESUQbVcIYpPbDVI
ymsHxomxPsvz1qtijX4x8r6bD6VFxfVpUYN3w/6CAEXKmt25slftdBFTBX77NRn5qxpN8WwrxRuU
7VtQX/nQWe5Br7FqbkTjtuFQx4XJYRuaSqlpiGOjOI/OgG+Ho/KbZ0eEHLWAlR3IL/5QDLKJwRBh
idbPw627SJFabCg6pZciWTk6IQ/HhhosED59xGrCkifg7sQx7GplTx9aZwzJX+7nuNWaDBttS2oG
CL0k2n3b/sT0RjDgAD+b+zn4Fc6WQVJ1YlehJn8LFVoG4ltIdtPOqtSidC5sLMKFHdTGk8Ik5Z3I
ZOLkZODx7R75JgQ+Jg8vqfBIBmhom/xRPcQMZOi4WRyjJ082J/BYUB70w/F7yRsOBm+Cu9xMz8uj
phWU2SoYhhXTLjWQomdmrhFIGiDYmiWhyiO+fXw81TTVfw42tEa0VCO78pwH6MzbZVpxK/B3dEIz
bQvsnTvUBy8O1sRRwhcbosE9TRU5v3KCTvl5aI2NDL5+eJAOYSi6mCpHYvrKyDDr0K1JH92LtTJV
Az1U1usqKfaTiFquMZOjvre0A+1Qnap6cBnvKeXGzrkavDDGFEInpoy4+lt0A9lvfSkmfVno2Ojm
1fQz6ab1Vhl9WLt38MJlH/pJxsNJcVC4oN4XoetmL/xFF4iUTylzpXFCOq13Wp+ZafT+9BFss2ks
6+M5bMOdmD0apbG36/kvBIcCHnMWq5eG1JdWjCFEk+O3pwHDjnPefEmlakMs7aGAqKLtHk5f5NCD
mysyN5LR2iSYb6Ci9uzaIRIc2+o5aeWkanOv9fJi8ElV0gEyjHRWp7y8LQvC4sg670RUBSi+8/we
a+QWO9llL9SgWO5O7X3vgRg1fiVeL5R/tBUNICuJBs8jav1YS3WXs+emZeILhDY2SLDdRw2Y18/f
RF7qaiM0NMid37jZ9SiHzT/SJUUbNLvdtGnLY+s2tmSXK4Cl2OcWaQKeXaJ+phSRgMbegNeGaKx/
KP4k1VJbNh2W/qRC4VEbd1DHfrppkv9xBRDZZzhb3gbseygo9isPBgwV8MyEH0CoyPyWv9YXt5Ie
etwYNQ6OtC/wjI+EV6H490RzN65eq7djvYMd4jIM0tJJhPQDexYiCBZzcu6X5jwndqnt2JrNdN+6
5WY7CxfJDvrWw15Vwd/1UEhTp9V2acIpt8bMCpTR1AL71J+jwifJ3AiHwFXNdtB8x7yOnNNY71aG
LjNTlhH3cX/ebwdd7yL0G9zlMmjt20dxJkmwPTPRMU6GtBc8FPBwfIVok6+vWkmNh2vw8jucq3XR
l08ngkPMUBiaH3L1DVZjRKCpHcAyTx9kwXdm9qStzy6dqv1fwOSdutYF8HHiYulb07Dd8KQHuAUI
r/5YvTonLrvc9oc0icSb/r1ke0x8ZuRf6VdxlpaV4YJCXCYTFr0T9mTNWlSB3EyqGGWfW6VMMX2p
h+lSc+Kk6uMZkyBTuUvVR8HFbsPysu1QsdLb1mC8/adou+nCyKT30+iALnFE5sxcgI8URp/92H/Z
ctcJsUd3cODScmpI9EFrkxp5GF5nZGOo3kyPpHB8M2mn2q8vhyXIqF2gjoxzBJEYYdRS8QFGZApM
8xUBl7IgqgRbNzr3EAlDQCzA0zdsswuGqeC+Cv3v/VfveEMUO/Iv1RhTMSW03xMCOWhceX6IJD8y
g6IuPNXnC9B9MCENIl70CkQEsqY37xMsUOY+erjEYfsijmohYM6w+lbgFQOwG3XFXs+6g89Bpbx5
lsc1n+FCIvly3BOkVFhZDNBQTSsLn9oXn+6CgjkPGREP6C1Cy+vT3EEG8E/dVTi4gMISUd5WNW8D
4baYUda+kRdfrNZtgBu6OB4uQSLqQST0KSMmWTWLRAbt2xURA62CTJnOPTY/JxM4HbXpAI0tIemU
ciyJdJuCzMro8/t7hBjKyOVFr075IgE70D+EnY5aiED62d+NdYiqoxAi/3Cx8QVbw/strCnIDH4d
MohzcvJyYtr5XdgHYGpNNba44pG+u7cbGvBkdgjo+CSQvtbn+dNIqjHbfzvdwIak3lUkF4DTdCXm
95Tr0/UjATxrwVVn6rq0B36JKM4bBtzguOfXDBJouOcJng1bSUqHVw9osigP9KPtiiFdP0FUWgEM
TjEg8T2FovE91DU2T8wI+Rr3CNPiXpq9UB0qntinwrXWewoSXRQUnt9EMArgjCe+LR8SKVgD2/yE
BSfXt3Cu18EkGDrH1qQLwjkWG+zybJHHBfT13b3dwmqxK1CP/33ijXdGhlG4hZPvqBYrQkuLJdWj
kpegfYLbraqBCizXedwwLkHFMS9Y1w1B0qh398WB60oURpsK7+KHjQrQpuTzL8TNZ69mTrmjMtX2
AJSpMwk5+F/gP9i0L5YQJy3zCgy5BpQJsszYLF8R+i0zfRtIVG1MqOYz9VXhoViNOkh5QpR2Ty8y
Gl+Ile8t90MOPFlfiTD/iS+hmFLp6K5Ab5Fa1s095E5wif0zGfmY93o6Kg1/mxPEyUg8p76+jCkI
mpQ6R6snGTyHIV7RqEyljXUM48PMvK6uLhwuBkgo6bgEX5I3wr8Z21BKpFpDGHJfv9E48C7vPOaU
OAuMG6TR9Pe/PJZECF2Usr5kQo5b3z2RuVOtKAVWEYtyR0QMPE/K6p85htI/L6AmN1i+PaaIf4j0
bcOJNlj/op24yunJFRKD4iQTf4aMKZ8ecglgLcmb5RaperQje9pyB/EfzZAP+ePkbIfJBqqXH9hn
mH8hqVpbVdqv4+qOk374i3SNE1HnamE5frDJY05ew6whLcD0gIK1S0BvuV5k3QiS9KDorMtDOEJH
jUhpMLX0wIlh60zPNr3jiE0Xu+RyRY2jsqhflyAfBfGNFucqwXyvMyHh5q98n5ypRCkQUOovnLkB
s9ae5pwhgt6CYahYP2ybwrpLkSUSh5PkU20FMqYhyF2o/I+WSeBItStoW9FCqwXIj42w0+HBpco1
JnjndNfjsKx8jBrpHEejmkNfCOE0J0N1f+TB9jTXpQ+V8ReJkujyke+E3puGylzoH/U93skoGvb9
X/W6AP2JBqDWq1E3fM1NTAQSEfPPXf/1NA07PznFILFPhi1ulYG6LpAf1OWqtYa4XjKdOk+3ovk5
e7lXltgQfYpDXJ6M/JysX5SMszmyCb5cHqx9h9njCs/mvQWS+DdD+o2AfVOiLpzs7Lkm7FLOoipC
63/ZyGo/HpfaI3AW951S76lV59fcRmOjX0HDsh2HJg9YEUeF+RjMEatmKTOQ/zHZ0vW1tYpgZ3+W
VO9W+XRS3jaDsQxKJzSBnBMKgAT5pX0XYPntwSsjV9cIlHdXDxLBXgcfWTjtrKllCVQOQsB1rpkh
g8nwQguBC5iz8j7+T3NSFw1elugLW13eFufg+LyNresl/gjv03rzRvPrNn8TRRBOHTQLPM9zR+Kb
oNcmqfStFLsdGqwd/HH9TOdNI8j3nc3Oolds9tc7TLsgeMFXxPVqQLcnSq2V3b9D2kBsbyX1SGN1
SeJxsG5jbKumbvXE0YCFdTkPiSasDlq2vU/0Cb325Kh8NLCyZ1UJNr29wTOWvNx/GhxwX5IjinmA
lvP5me4CkqdUmdBCWlKAAXvqewQznDAnbiJcEUbAArTfQw7QMjh/yMnNZcmo7smwFex0RjVyUBQP
T2fCIC7kAD0IfO4S6PchgUmEJHB60+WT8qJad18y7wWzTt63cniz5YWgoXSejRJhjyD72NAloeQH
f5ahY3+jl0IdyE+8/O/Zjl1Yjc85+qRiOeHSUwG+kU86i/xs5NjxheFlP6U+R8XL4qPVHZ/nnWni
2I1erpblOZN7d82BcM8sVHPF2bUy48vPrkpB6HkBFgx+6G+qYEskSJ1qj9PQjEn0NJ4YnYpWLRKo
wa4IFzSyPz7vujwytPVaGnubhR8wccAaIdpRpztyBujGvrq5w5Rb2iTfEL3rpFzhRuTfjRp8GB35
7E8hu8IJRgpN6Yv7ZBmXrHrI4sZ4J3WsH/N+yhrvEhhCNionDNm6dJVt3iuwshJQtcBUWFZUTDY4
hBU2cpXaCGZ/Yk/aq4sloar8ZntsILJ7uRkv1+20ygiGHjXgGDCIMmjX95GrAnm+ZtNt296xVBOr
jiS/Cr0lzWYDjtmUT8OaI/sdYdB92DOWIJGiH2lwtn00eoNcLKwE/R4U5DkxMBQYp3OsFVnF0VuQ
xN1NJcS9wF613BfMGzJhXVTFcXkA7qspzOF2iwYN81nl05z5P9h+BepuJ3OKoUJLCGJMCnB9s3it
PuRGN5crAyjwj623o7IWEnMPXKEAWw36wausyrxZnJ+5Puz4jFRrxOgeuLPN/jaziZHWaEezQzBD
Rlq4kdKIQyqq5KMDb7czI6EmFYj10gBzA7dLAcUljyWXCoPqyt0WCsl5lYcDtOU3f+oDtypiqvfv
knb47VUoagezuBzDedMYhpc3+Ow8EnPKUokC92guJDlx1PVhu9KvLLZFQs6zseMTrg31s6gc1mV7
fBd9v8koD18XpbZpPKoa9CirpY64qt7+UPNgHbP3k+xPAnetn4giES/S+oUTwzglRnFxif23spHM
5G98lAECd23fGp/zmLlhikdkr0P6Zzi0u0T7HylPx2PkInaapmQblzwhPK2C8cVDVjHY2wc+1vn1
Az/TgIHRrbVdELDFw63oDkLNpmb3aqT4ye/oFDf2SJFvsiORWVJjoXraFhywvyX8Eze4tHtmMGn0
IXiPunFldLuIOAYWil3jDHRABe0QqBrWeRWToZucIrYR7rklpawg1ALl4Tz2FJ2+L3b861B/eWZ5
Xhtq5SG1yxpN5UGjWGVnCr6Uf4mC/HZEZLOgs3BMSobHrizR41KGc3nyl6fpuKZLUVKTGR494DjX
JSc3ByIOx06RO/Ux/i8Jk4JD05BpnEP/yC6yNNnied6ojBGmwOmcsIfzjw0UTKEXrnKjNq3dCJYm
F5JJu7BVhNB04Jm6THwj7DG76G3qhOevQjyRTskRew5BGN03eGwm9upFPasuSRdasSWZwHjAIBhu
mqMbr7Fj4pYeVICQ50Yl0e3cuoe/0EqmrJz9CUwFKlbdV2AM1Xlk0o8mJHQPPe0KwO4arBTekyyB
5+UV1FTzN3thdh4cgvtK28SgExjLGO2Iny6mD+dCrW2BCTrpaOUqw7jxE7nEM26MyTbWyVEjMLTD
bCLrA5iZV+s8l80xtneHIU/05DlYTEA7Tgpv1pZ80EXJzLtdiPK1fu6euuu//hU1uNY2S9buGdPo
ErZwt98tewkDqNc+UsilyOdOC3FAOTLlBj9zB5E1zpf9HdS2XMuzWRu7N4OubkfZZw+8naH/x6TC
6snNr6U8lH5xGsPe2AnihE9OElsCwfrBxgrTIJtzW/Cj1O4P3zWw5rrqOoeAjorzRjeHRmOOvDmb
Zt7lT2BCXUF0Q98xNPrGJrG2ErcLFEQaCd4oLMauuVvllOAeoGWgjyLJomLKP/OP3cDVZ2D0AfTK
vH5kUmtmCHX3OPu+WTG4v57iuHpzBRX4NvPqAZFfgpL/+D0XGL0LIykiZ/+EYKYMiwpqro+xvofQ
T3nj/l5MAERz89YVRmxGeV3flqStsA/kdnG7Cbp9lEfaDScZINrY8K/ADafeKeYO5MAlVJumMOKE
N6fuEV9t3Cc4t5/QquUMqd4q6JLkMmrgyWBvxmi4kDcnyLFbSDo765CX1YaWLconvZq3kH9NVH4H
CeqOa3NTG0tdsgGanu9l+SZ95WzEzubINcScylhwtWFl3f9qoxinj/A5+vY7qTxhCBh517YYajD+
yoxEdw9Be0yvyTkOQ8fxdg/bTH1CGmFkeGyO/aVi0KsK6R7hkCvgDGIn9sDZAy5CFvsEeCm2aVT0
PO3/d0mnlAS6s8QKO/U8bcsQSDucIPu/sz7iBQavSEK1hdaaHCEXXVtP1TdE8TzU+Hcs8jMqWgLP
7Vwc4WElOCbjON05cGYknvaB52ujJoqFstWAKpzSgrh9wGlFVa0cOAWC5DBnMhpOizohvVIzhkFy
FmZhCSdZdaBPzylQW95gdmDJYdOOnr5oLeqRCk+DBWZdrLB2hqAllIbWY9hIDBK4fuUd8R5SwdU+
PeCW66wNz4aFQkOHTeHIUiCdj1nOuL+A/htNLwZs/zBVAGXETilnVEA071rNu0CNIh8xILvOBTL5
hXnuyYhgcv1KhyCeYtrIsXvP9/Zh4LhMGKcXcE2U0rbAbSlGLxQIYuXZ2ENhZGbW7CtId7TOSbfk
K4+rKUCHvEW9ETk5xzYUknNRqTrVGprvztaqyyBVyahgsSYHZEGXUq8CjxO87vvSpyBO77PQ609O
e/KO5siDU2r8rfcBBwwCLbP/A4iapxPS6kxonQePHksZYOUfOn2AMHsaot2ra23JKCvNpM6/ZGJy
9olsrAImcTLz/Rewwhvx36LjFCbPXMVQWJcHVkk9IGl/lsJpw6eQ2aoyfxR8LQyuhBGf9bT8dXkw
Gn74QSXMpQfAPNeiLvSKAfnVj3GsBRokOCYQnETAQYr0q0CZcK9XjggJvWGcJ+xagHc79hEWqFaY
cLpqzz9Nn02+xN0X4gaDTOye3C/fPX/PbFeBrbT9R4GOvU9HJ5xuoE9r531riqIU97QGpXSY+5xX
L737yqhGY64QT8WBGaw7juLsnRyB21yRRBTjeuGyIvrsDMZJfYkA1HV7Nb9YWzaN8ByZPqyN+iRS
z8DWEbVvN9hGYoLX3C6CWMp4twimsSGDruI07haJox/uZ/NAwOAH7Au1usR7osdVkkJkYmP1/Tdb
76cLQdgcgoaCt70jtTHgOhfzZ6ZGv8iZp/4ACZhtaVeFpWIGei1Iy0VZ2X+DnKu2d+pua75Ac+wG
t2eKKwtl8a/4QHPx9BnvO0Jl5hW+7eszqsfHgpA2P8dl3ic7tiES0JHJ/EYf6tENjxMNwhTP0spR
CDVDjdHrLVaANr0f4o14NhhJwmU5i8naPcyr0ZBV9bt8+YaqK01zos4zSHgPPLjNnJuMFrrZgaTc
KboA2vH4FJ9epoVFlFXSLwHE+CNbCYbyXjOnKppst1Mn49L36ZoqKMgK8qzfrNokkkohMN6hcQVA
RkNaY2Y0C+uRIsSk64JujPHQ/TKAntyuL4f51NRnl5MpT6/SUhQJeG9DUeW9RG2A7hI4P9USHHwk
2gnmCrz/q4ZLOaoepyZn2cubNSM8DWj13qbN5/auR7Y3urSfpCfKPfUTWLwyNk5yDe/7bNsdJ4x5
+w0WUEbVrtQxF9mzHP6Tj55IQDtolcwLcUcW3wf8IaS5kWOS2vsWJfCNQedPQoKDmTRXZAR8oY0j
dN0VhuPimxWMVbJFSO1zaCJzRWdhYBDldsH0IAk5nXr0t66o2o8Di0I9GFCutah3XILRC+2qsqOZ
iCq9zRse4J7AwZbbj+q8YmMQ4Cg0oh+s7EjAvmZKmHwy89MatdkDsUTxoF7fV3qGLc7+BoxN32W/
4IrK98cs8FF3FMkO0BDWkHTycG9CPvKZCVM2ILEgyLd1tWm/7lykuu0em1hLBbGYm53htjYFcOtR
Mu7SQL/YVJfL7zVE56kQ7xZRGA4KYxHq8ZsYQ+f7qJmeykBcQ9s9Yif1Qd+LK70vT65mN3apDbrj
T4M/JcwUq3RiHnKSemnku8oEegkzTXCP30MaO09sBqig2+y1kdfs+aMdPF3gy43B/ZdeIJGO2Cmb
09Xf8WmstDM8mLc7P+97DQhlJMBpDIXauJfopOPAgU3qzDHptFCYJxsl+dAtc8zfWbAUyNk8SB8D
AQdm9qsgtBfwn3avpBNnY9Z94aXs+GUqsh+k2VTE5qq9chRVODwhCG08nIINtjiEgLYLdjcZyGjY
8Gj8u1rIyKVOaJr607+CkhaiRULNZr+qIZyosAm24dD1NAfHdMSij7tCeR0I/F3WttcVhp7j+sW/
EuHXulalyJ/KDxTBwX69uzEDDn3CQTkGG1S0T4rh5G0uzaJIs7ln2iKOv2s3SScBlyI8S/O5wDpX
JBnO9v10HuYEXg05cGOcMH9KcrzFYNirLzSqb9cQlh5RxS+wFIETX2PHizcb5ckknayTp2N8Xtfe
3KORpEXixy0tlB9ePPvcwKqHgFx7mCajAeAeLbdw1zKrlw1+2nrcyXE+e1d2Q/McUP4JjlxMLK6I
cT6L0m8R2Q3SWp6Ip2W2zRQ+09Nt4WHD+Po+b77+y1zxcY2lqCZQB6I4s6NIaSb0BeChnOquivRM
eV84xHWW8Y8+ukX9V8a47p0cHCQcgPn3ZTXrzfOWptCi8aNI9077WOgDAza4k/ThSias5O3SHJZB
j5jJOJfQ+dNRLPzolc1Vdz39wWZBHbMFyXBV9RiQgYMOxbwG+Yrf56MY35uU9M4ElZ1YjgIdpJkZ
vgDdkuEhR2udq4dnMneWHENgt4UabUoL5PVJ9ZDkUwjmKawGp1orcYT3JRBL/sqU4j4PnU/43gv9
urINInbLv3Wm4P+J2G8JOFkj3eyhK5xX/lpwKd569SfEVwuCRVoScwg8a8lUkkPE3dzV27CBjthy
C/sSP71fCViyhTH1xG4mrOrroxSX/H1gDV2fF5qj/zHwWmMNmBdZSuOZzmEeDO1cfymOz7MJJATc
bYQtJwXmPZUe/ZuT5Wf67CUcCVDPut3qlj5JMV1iNV8GbAQggMSqUTE1eQoELxR3Gt9Z5mYrWo9R
q7jyOojYoJqwayXjwg4f94dmDQfH45wk4q3yQ6RWEIxq99bpLuZ8EVvXZ7+RiJD6yirk/6YDH5vs
2nEE8z1L2k3uesRdEMypkT9Im7rEcHtSUGDQsezrAxJ3p1qKkzZsrGsSypxMgZhHpP8SraFV6D2g
8oWJpyJkulVYKtMcQrXgfPmU/W32eM9FXQ5/sgL80zSiaaoDik+S9MRw6KDK1fL2IpbmFJOhuS6n
xfIqh7BNtb8fP6QTBS4m/SymTZTgMw0tgxOd/jNGsbyffRJjFI4+vVjQG6DCLl57xvBYD/NkWhIg
c4EACSM9fVpOcb6c02DwprDMP2lLJZZLihWhtIoFvQUSJXmwmv6IwAoYEJLpzjQc6C2QZTqr3lp8
OWewD5CDk6UaS7tw4FBQBwqkUdJsl+pQTDhUUXYNCqxZH/p8HghPqrty0E+ZIGoE6E5lQPCxRuou
DHxVKrVpVTE0DofkSnyrgwf/f+WOdpP6GPt4MAu+MuLo12HB7cLTNve/RaHsxbWSKi0RugjQQklv
mMDaOCsc1bwAK1CXSjzUiSkOWH995aMYepeTSYH1qnU+AeXLClmtvkkcfcr6PGMZRbiibKn5stLk
JzbZaBAkeFicFLusDMzcLDKpkVjAcCGJECCUuH3kWwxpqAM5Gnjl49gxmN+ggR/D7fE3pKurFk/D
0zxuOzXhHfS6H0VUPjoo/l8PB8P0iQYzmy12aV2cnedZR5rHKBp9vLbl9j+ccSEz2oqadwynqi4w
lBe9klf5iKF7qfaihlo2h8Hc1X6HFxtUFpEIKQD7t9OzocztRPzjeVpyClWL9+gIoPpE+llhNtQB
5ad55xQqManwgHsuMTkVf+uXZmM3cOfAXMjfI2cqlo9f0a5zDVelZLG6qD7RtvQn0dsLiIwun7VW
Gn5mxe2V24QfLpNKJ5WUFvSilx1xvWUu7KwUvQxZ+zLpGn8itXBJLukyweFQhw3AueeEpIm4t//8
ymkpPHDN2pSc9vhTVgMfHoVw9vN1obeIJEcgNfwwLUWZKnIIXYRwCj8vhaxln0opmMtJFMjtZ/4F
X6rh7B5pEtnmDXvbdRuqf+f1dNU0SqqIyW48IuWnKzJvCGEnqJl7xSLP0nxafR2hMMXy8NGSsnr8
sXHQ8U5ISQfS5eFEVPhXDTQMt5RzHsmX3w2Lq4ustDUV6uKNZ+QIgdDjOd88VGznrToctYwBrv+Q
RnqKLrnb4+rAz1H6QHbxBAqpv1nPrEtsFkaScWdUz7q/gk9CyF6JddQzSLzrznhnWOBZjh6y+TLB
yIwcu2hs25EgNVQgjq2UnO9JRGr0OEIK11tkF46G+icGOnVU8SG7Miw+a+fkG+U2vVSkHYRrLqco
ujknjUHhhX8TjUNY9PnneVxW0e8IvFLsLgF9LHFzdR83BmS0X/ZEl+VDAc/mr4Flg7u2OFyg2jLb
XqfeHVwfzjBzkuOQShQAwWjMi7jXtlNidqCGpnLunAdKTTQ2lLW5PabxE7QhCr73TQrVg2jm/3U3
8zfQHreE87s5IP2WqWXqfkPIqamEGy6noiNrFtAQajThMbyOIRspaZr2RuW/rJi99T1YW3lCtApo
43SKGyPqaAuL/ZCTaKIFyypXumlXUD/kDO9ELDzbBx1ZsEdYNP8C0GHRYhmMYq0b8v2OJGkPJ2Ti
SKN3SZL+MWRIKdyi0iYzqWCE0damOJKs90QJxuYKYIkLHFKnpvRHMypEj7gKoJ8rJ6TR+/4b+OGA
k0n3ZF++bmyoXI6A9daPVyj2eE2AVSFZea6+Zqpus68omd8XTJZ2+NTnf0IqXVQn1JcLs+0hbXF2
IQtB+JqqL9NXFRGm/plsznUSSXAB2icCrMF0AThrq99fR11SVkHl001OphEu9TXvSZIUpzbtqjdO
YH3Ytb/pFBGrK4FA10LtJT6UNSN5OYjHLfIWwy86eHlp8wk+z34oBYuKYSRDxZiumPxsYjj0OIqq
Mp795jfIOHrh0qYThQSA/2Tidpi8VRILX4lLoNqVRvjLC1PaY29Q6AjJ31L1pZy/m0diWb30xLcp
cmVWlt7GIaIf59rQ+vpD8CayGnowfapu1ujVd9O7ltLvWbpBDHl31NngrcYAPkjhbtkN5e2vXJC0
n1U+AS9MsdJg3wEUwjApBh/5qfKyROgruTQwKbEtxILEDFBC7tJbaa2CafYDv2ZAotitlAFG6Gxz
iwNGr97rQfea2/pieM7wBcmgChb87WAkiyUrnAFMiW4sC5R4qvtEw9y8qlqEzHFW7AQnU9AcVNLE
cTW4bVbOxHFTqU+AovtyMKumic2WQe5vX5B5eVMECG/bUyAvmtLXP5ufpb7ebcBj70jO8xZ4TEO4
GrDRJPD2HIYhevP9hkbv5D+VXPEAJXj24P3Gjlziu3dWmDx04cvlYae+pZS7FS6YGNkZEGGNYsN8
88nokY/QnhQOCCwugJJ3E3IR7HLi/Fzgs7znBgNtXmm1E9bKm9tVKx7B1kG8fvLTMKbrF/uB1wje
vMZ0DYm80nlagcHdTZa/L9/eN0KH6x477108IdA9WPDN+L3LF/rDKjeelGRhsEWIG9YRqm4eHooS
V1vRvpp/MLtBkU5CywMuSqWW+9EvAhsJzpwuCj7rbZV4JIS+bLA4X2Sdr8p+ZmWyL4U3yI0nCeX7
cW8gKmC0Zx+xcYZDwilBKQJMap9GXH2aSxyGL7D4/l0C8r1DJkhfBESiNOBxkE6lTqWZcJdcbSvU
MGOTFZV5lilnxd4dMBEEM6AYEzcyEAOSeF0lLr9otumS44Od2L5j/EH3gfPUQoag3WumYHZEF9Kt
AEVhL1VqeAkFLnsx3ns38uXcJLxqp2UN2LoB+zDVATPvrt6f0GhCZKN3THi9A/Ax3kyUh7y6xCUi
iNIypTvvYAO0RNy3Csk1My7Zx5S/EvF6y8PlSBgkTkyXI5gXaZD6+02FVIBxQftFGqioF8aNFD47
8Q7yibZtC9HmPVT9NxnkaPesU3KVe6VwoGCIJiDJl+JR+8M5Asx0FEdwINv35hlISbimCs3sEKBk
iNaihNhHEP1IE5td6t1YUfwWbgpKb5FmkZ6zzqFfIyQwjWJgvXBhaGnsd3fTJkVVf35L4tNkAkUs
DEVFMbNEszcu/JQeOQ3b/4lJ1XJQ0LOv0EhwxlvKdHOpN7v8vyNQ7K1JVug6X7Mpx5TjCvZCOM5C
nOcENBClkI4f5uhkZYlmxIf8gcj/taBIXQwcd5GWkVGIb9bURkh+ofkUeQQrqzp0FERwGqwyBUrb
UuXC+k4XS8jfEf3hMPk9JM26I3ocsrkciIhCRVDt+j3vUh1Gx887VxdR0cbuy0ThlpxSSiIrNL5E
ZBpxbtuDd5medoU6ak/TlsZceqPFnMHj8VaTdEJxcJ4jfmlA7LG5NH+OboHfYp5JDiJcttZrdbqR
HdFSVkIzqDAe1Msf/Iyba1HARCs/vFFzHJOwmYshQyJ5tynHzzYQPtziFBbzaZ5cbLHfT4S4IYt7
eBzGMk/+psjsg7/zwYpMNxdBAfF3Pi9WoLWW8VB0aXAZHJ6QnpssPP+FE0r9z/MxPxZ6rOxbDrcy
3kFlaHjq5Aapvkkx4fidUcNjrZt5lTYgWBIsI5jG5BvnLcSFzKszMdMDrZx+Fp1WZR+Qur68zdZ8
Dxc658YjSwpLw1dp8toZ8SdlDqwcEAvsmKbIv97cFuTqK1Ux59OqOv6FE5+8MVOtezhCE/rcu449
GC5lk7RjHSqiv/Op/AK4LLUfhq2tbpDad6xYmes5FYN/m3vQwZDaOqEPaGF9ciNMPgpC/1V79LZW
j3ZaS5bE5eJ6kjoaQc5U1n/isRP8rNNb0RQ78HI4IHDzkx3cBN6sI5V+z1l1we+xYQ5Cw/2OWdsG
FNlkFcE0kvK/SR0DCVwwgmO8Ux0n1BS64I2tVZpPEqQ/zXPzkS4nvrc9GMnRqJi9lS4ec0WuyVTA
/kGcLFYjk1MOOX39+W5ajPf1IoM7RqG+rkEYU6eX7OuIP+aVVryZQaafMjW2DPTZS2T7zN2kMEBt
CiyTnqirwkZLP/lIZ0I88iSTmUz1jgoaWQ0vXzeQrcBQiHpa+Hj8Mkg0/NonUVK129h3yGsMxIGn
QXRLdSqN3d4POVMwUgm3tgJBl+sR0AgJlWPfs7uLUgxa0KSJI8dMSmyMOrx0uHRAowAziaZePKT2
D7ID7BjTo+mWe8TGtD7fhpCuOY5x15IVvGSz7ukzF1XwthzqZprzzM0DdnOYbG1i2HKsoML+VuB3
wfXikspscg3DN7BTFgOimCmUarq4OXGMCUy7fqL+67T5COrGOgDDtU6nfci8EAwwThRs/QF2knIh
epTmW6JnDgBJS1lHpRXfbhL7sxd33XHR//Y9F6hzxSk8+cC2zm1LKFy/m+ivhMqQjykCv27wGb2W
z2RFGongdWcnGrfgLfNRK1i0S9zRW+Q4AcaaGZ6pTcHLnwgz2EBQ/fDaO/sCIf0rDaL83NViGgYn
k7hLkwPLXs6jQtOECflZxnHerNQQPm+MNqfJ68nA7F0zCkiocFTo0/J8SqroydPrZ4eUgKgjVmch
cSt3tFvDcl1OucwW7DoXl/48cBLnxtz132JupTdkl+AI2OXbB4+EC+3MalULqvwrh5jGfP3U+oBs
641xWKw+KqZVOogHky7/705JjU1kzuHuvEHqFkTKNQgFbymJ/+a+1Ugp+3U5SmJ5WNI+TjlBE+mN
Zrf/JQgfXngqniUcbi+VkJtZMLo10NvfCAMI78iqnzO1QgiTarENhyV86o2NdQ0cdeG5FRhPrav2
QblofBWvPsxj4S5msmi6C9h4YfnZZq//sgj0qVWQlimi8VAAfq+QqPbeIR1K2t8SCdXytrPwEDb8
vpmeC9E6SbBsYugqihhZ0rxJCRt5HFK8U8PXL4JE5WKDXkkvtBrCADMnoyvOb0jBMesRsyWWwzTC
DbZJLwV27U0jbWJvwxIrwKQZnkj12v79I0Pf2ensEWtf5wQd+0i4dolIwpll52srZ1LPBzuEawc/
VktLTpNLHc2o7p3/sYQXjwypKGxWmMxabuCYS/h7kTUIOt3BLVAjYVQlrz4nY1HmHnPax/yXDsyP
WEiWJWC1yzEteARB8i7t3icZaInsN/A5Ol4Kf289yGchkksiiPDEXKpN5kAnLhP+yhUeJJgoVp19
dq1Xiv9GSM8hVmiPHOf8pdB7dQmsfZhxQ9x//LwKQrbbHAVBzXUYXMa61BeRedjuJLf/abQRzPcu
rgW2HEEAhWhR9KvIZ5m63+w9gjgJPDVlUX+aVGgyVJOnqRfDp1MNo2qxfp2s2GsBy5ArPgoYp9zy
OFyDIpRGD+/C6Kk/WEy4Le74pZmRKYWGn2yfJnZyQdZc9KXjGspLsWWzdV7BOzYL+8ewl3TvfO+f
XHv8BaJ3TR3TkTIy/1sCjcU5NT8CIVrNXWo1NEsDFHquhzd9uMe028CTZ++GlBYIPH4u+M1EW0eg
6nVl5tkpLFw1gXKLeG3dT0IOT7KqwcV5EiwYlRc0sy62aNTl95zXfAVmm4jQ9Vv08iya78k/HxFI
AoxrmehRhhhQ3HKz9PxMV2G1jRdfEvuvlsXAZIOEP94uEiGsUs300C8t034Z/GFnAC2wATI8CTB0
QHdtUe3oa2PS+iiwdA8c7h4pL75rLONbV6qQcDEJ94NxB3J6MYZeCoU9NVwdGDD6gvONbMR/oF3/
8NnJG+C6qE0WHcYVXp78W0uQphKNRyCsIdqCCO7J4jEY+4UPqR1NE0MuCZQyxGlboeMia+BRTZkp
UJTxaBcczV3vhqsAnfBkE/44ABbUjsKQknDhesNgYWqw5a7csJU9IDYYVLm0TgMZP0BC69FmPc77
nfi6F8SU/4deA7ChIrbSwvKghHW9w6XTRSJv7Zdb6x50K4R9il3idKpqwL517C5WeVJU1kF2v2iZ
OEyaxLK+W4JPdlLsMfnixM80yeO8GPSaR1KIEMZGKGO+HoVBn+JGhltlBKUpj+zhp8FCbnIkrlqM
AJbM7CeAsCWEDNQwPEZqHSX3Q9EVXPbFUqKrb/9N4MRVYysjsQiFu4aj9bmkobnObG3XcjCjxcAH
2kk2i0Q23jds7CM5uaYdNvEynnhrPbLUONVoOnBpWXuaSdDqiV9XmqoLDJAnOKpDgFAxkUSIZhg5
rfl0LeOhyGk5qYsSvXkI+Q6Xn/S21QVcBffOKq7NRbzTbEqkALHk+uS8gHezf+/pJhkVp2PPy/ew
MeRvpgVdo0dPnqkVe46ZferfYtP6IsNABHpqhbOdMpoAOw6SGb23Ft/8NWcyZtJmGNuhkJQWpKr6
5ZvCsf/VYgLE+l+saicgSQy29mz7bO3CuwXIQcGhUeYfYwMbUgHT0ziFyO/tUPFQ2Tfq7JH85rP5
t8kfJGwOPA6Z8xZqEwri85/RTTVsd2u1BGI0RSgWPDpi8pET/pDpXYpXlf6BFKs6+m/EjMPbmPfe
Fq0qPdxA1LlO37/NZNpgGjVll1tnvXvpCbiClju87cK0+xRZmctuCroI4az8FLeX6NZhbHPOQvb+
71r5XljLgsA/LtbilH/Cw8kNNpU4hruJGhyZK3htBxeBYYk5UTiUKqj4vu0lxGvguI21WkqWzAk8
Nh4eI2wmAF0tcwO7H7cjPI7EO0cwH48+AapXfDLSxUUdy+A+tlr0n2hOXiLxVVmxFed/LvfUJXeQ
uwFfKoVG30QvYGjyrBy79s/Y6H1QrvUM+GSoY7B/FAEJrywdljRcRK1Y4Hly18odMs225MumZoWH
SGwPD6oBjWjz0uSA5NlfouUT0Pl//hbZ3Tck0PY7yAmfsTFKzqdGxcnrHD41Z26aqeApEJs0dPd2
JTjhzjusDBZYTvBOJRWPQT3bJa/CIO/asN4Im1ri8jueMW4QkrEQqW2AEmRXGvhDITHhMdg+g5H3
x1dFwKGLGRNsc3rMQdepMKrtrrJz3tdsG6FRX2gAQEmNH/0Oix+OeqzFIxLSuFI+8glKpgs51IZA
rqEF8J8kDx7+FnPobKj41OHv3nJGt8K8Y/4VgGHy2cZiZcFnOStHbGP47r9w9ZVLu2WQiC8F87bx
bIlY0PRYEbS9qk7URRcelHWKz5xaLWL5D/0byA7S75aRnw9gKQcxZtwf72/05C+VPc+zj4Z555Mr
eqlSHRHGq6CfBibxxarLZzm/35GYCv+epFUmW28VNmP2ALBqEN9FK13yHuUaM3m5HWSHMHjsgBKc
PEXvwVWfTG/DIO9/Hpp9eSkEjFRr+/Aq8lpcCE7e+0/hamZHrqv6QYY9htL1niwikrM1QrRXhaFk
GFimlSkmwmghHYDiutAWs1T8Q/SRooBqIBQj8EGuVYwXgkIIKf62P9nVBfRC+Tn0erFqCfy8a21v
ramVMIDjtwg47orC2UZgxOjCBMJ+7MGIFQDx7kWzWsFhfP9jrXb5lbwYWapVF/aruaPl1LVjna8T
YmaiCpLEqg5VfWc6aGconOYBbHiVDYcOk8zF7jrYFjOmcCtcK4O/iMfSP/YOUD97yyZrNx4OBOHx
I1G1UlF5sD9FIFSSmPXF5ey/hxorZICYgTSiNi8991d9M2G5P1QHua+qO7xOiTIUYB1KoxsKobuZ
gnvVu40hSU1iwTM0wqKO2/GoIsEt9oK6XDR7QI0CdMqUu0I/BmKTm9rHAhdi6IHxUzadMfnMjYMF
QJMKeRRvKLGgaH5e6SR0c4XPFkXC6MGnfk/BcPZPtU/oiZcG2FeBc8PqVVgQqQJJneZAd1YAjief
LfCqYGV0YPxLwMu10y754iinywjnnd2th6eHQvOxCHuFo5PWszY+bMaleeyvP4vANPwDC9ptZESZ
kY6pPF3RlrQalzfgbN3zqIPFArvGe9LNoZzv4Iv9cl1Al4/25cGwACvfoNyGqvBHald5B4kVkrJh
BCfs0jelq1w6HvaWy/OACf3SmlOpkazjbnfMtOz6tudtDaWOyXqBhvqedMWWNMgmLNyCLyueFVtM
TYOE7Ubxi+Py/9gZuY/ZS/JvUnr/OvCDDkvuvCMNmsyVEV16+hr8iwfuQE+seXU8PS6MGafIVm/w
NAy86USLR97vE1fRlhWNcAioY0Qn7Bj83VjN8wbtKDV0nT+F5kGoEri0ShpMncf4bVuvqYgsTozq
PRa751+eev9MqZiHIcx3XOt+SCkW11PBhg/MC63zBIXbKB6beaoCSVue8HWsap9emhC8wBG0wNMt
RbkmAJBKDn81x1eO/lDF5Q5VKdiynUD2V9PxnG0/JV0apiAV7JZumX+S2NwUhKcl/u2eWzza0XDA
hnlTtQggaTpsSHsTehpmL2kRUd0IKAZ5NMizTr3B4rXT1sT7DqmcFQr2kcoxS58HKSKbs/GYAV9G
fMN5vJcD8/wwLHEnu5yGYz0OT6F2nHp+Q28p/U2/OOK1czbBzOYy1Fde0tfq47Ia8W/+ZFnQrlfn
hi1Hb7ETsSNWYwtSKu3ekAagoc5GTAFxb04syWG2OpMttY7tPc985qwSExfwTsLQ1/C6xm16ELCC
4q/UwpvePz+zkzDQXr+ha4LFKgvgtqKlhbl3/VP1BKhx+qRb0ecZ6/vHh0ssD8ZYRyIrl/0GLYl7
Up66Jdz5aASOY1IXRG1XNYD+EJw5RxmwxwGTb0Cnd3n2fj4c2fUKq4lmxy6VbqHiHqzvFGCaypdT
eQy1Le0BMhys/VuIpbQbYbHnxqm41NjaCyUkFyLB21LZP5y8nvBmQd/gnLUnRJnC7KdQc9+ZvVIj
FmMBjtIswFcp+zELfFfJ3Io3UbctX+yZBomT8mIyk5sT9xBR2V62Zhbi8HWOM43obEoaOOEd8u9e
4UI0NddmCCtrLZ5RmqVPTk0Nh+9ePFGMD+PccnvfUo1wCpNmqxX8N4qF40GBjuTYux9SHQyMpCHf
d61w28Gr/ofPnRGi1AZGqswH/r0EqxtEiUmQ27eUHTXmH/KkEq7McRp3BA/mxw8xlwtNZO9PHEqk
EOp8uS5TSBwAVTNOhg+R3Ez72oMO8elde6ZKoeV3K3aikuBOC39rfkmH0PT3iXqbwvtHNpVXt4qp
Vh9yAAKA5ycMdmIqvUVhyky/uQbp47vF1G7aWly3ZoVi9QjrrRHvL01f5fU9T/+AkKg/TQ9gCsfp
snKZRW9jRiYXiLjRxADOL0Jey1NwUtj0ug0DAdmZCOfUyZYWc8tUDxZAjNQ+hRVmThz1NkMFqCiK
fWMbwHSiDh8ySZBma5VJRafB5kz+Fm8FNY7KX/ZYDshl/0UmUdHFkVqQomz4Ub4DULbbUbpwjOiU
ymoXqtH727eN4xUcCmdAPalDNZehO/7n3KvsQehPSGRMoFrB4iD9DKSCS1aZD7QmxicN746gl2MN
8iWcDLb9pMoRa0531mjT45LtUV2WAFaKgTJPzshOM+1xF6KOCUHOsKrw+tBCUH6GNApFeMjjQtui
kiJrqv5QMFP2CSbQeUCiZ+OpRxt9cQ3SvZO5XwCOU6NxT7b1X8UeKKc5d4wxrFYNWgySUuzqx6Ob
yvaR0Lyv/mazlbfh1MsZxcIX8y2HmeGNtr6BUDLPyqNxiLxzh2niaKt/s8eF2Drj3fU9Xupa89aG
73S0fIxWfquayLxNK4qDaP8oFiHMSLKiBlESMxECsWo704JUhzrcQ0Elh/0dM2A4+YDUC0Jzab00
afjgsVTafdy2s7BctokkdBzf411mZPpiQq6F9RH+dHHke+nCtY1F8AhjzRm1xIPciuZQcN/ZRo9z
7sYM5PbwDV1WHu9yLE2+GfqHkxzhRFweBTS514anKAWmEZWN35ANCC9QEBvjL7XiWAkRB+Gj+pgb
8H1GT6iiJzZvJEUZobbuhnH2ao3JLmwoYddUmbDeHOWuB0xYBSuTKnQmc8a6lohKPWjjT1QuQnjl
zAbeM3ew10ku3GdKMJ19fmnQILTCUvEwGZ8LeILjoXyswhlS22sQf24uy9P6YLpfUIChw4Sh+xs5
yyFBeqDfNknIm+E+JMxvb1v9bRFjMo3Xk6GVwZjhlqrnVJey6PrtOQ4B7Z0YeIPcCrpZXF8vDWBr
JOfrvMJf/t2vyBguSf+fpdfC3FEBW0GovD6jakSYYgh035ZZHujhW7A1r34yfuT8vx22JREUardh
PbtSoxch6+ksZ1VxNvkoJA+5aa9b03jmblIeubclBq73pWjwiCESXS+gyHHyi1NdYi9HE8KPIBSH
A9re/3SKp0R+BT5FUHOTOST+lYY2xi5BFvW9P90ivCzFwYMu9qsi7PUTfDgcT+1ozORtvksJoMRa
qc+xQaZnPPFBLxeRiX/0LHxanARcbQ/FZW2ql8jb9BPahaSLnxVvK+tv42Z0S4lIDoZ9jyLHAa9g
rJd4tM7x9zz/XcVoLE6Is+wqP12NUiPg/K3+HfMzm/uqJtAKNgUgyRNu9uoVMTufJNxf+ibgQQTE
4QkERr7tiGxeQDTyF2cQZOGWBxV9kqmh0U9pMbs4qRblfH4rRL45uWoSoxtHPZEyS7t7pLlyx5kU
ZzzCM7R5YnQwcLOFODA+DsDq4VRd6WmldYjxPIjaQxtr2HAOloS1o0xoD2Bx6XasCoTqwbtExGXS
NpYsVNFHjbVHCdB0auFMEcSqDjgVTq8/OQ4bw83L66QhxmWLppfDX0Q4HS1gxDhCw6516nsq212R
1+KqqL8kVaMNJeqiwYkXOksBQ9sMySiMYd63I6hDPx8fQw9M4DIvBYvVvDzd/S/HYL7V2m6tCPHk
nusqSDvFmsNBQ9vFKl2DjLIsh3Cf0XYivVQxy6e3Rp+Prne8zAczyQVkoHT3QJveVDtUjPrOn8zs
SLHCeZ9ZqLfXz/4iYla4iCh567DkViDfYtT6xvIj8Y002VNHkaKNE92h5XN+anornuOkidRp/OAE
rsyp4fohoxqG9Hy0YD9hw+LPL2XXnLcJlFH53Qz+kX0pIMvfY+XdR3oVDIPFBr8e4GvNuGvNuAhI
MNQd0todYJ/C/qGWck0gBKPhBkhJVXLXRZAE8hD8qxQHgsyOlrj+7rz9mIb56o39dsU4hD542jnp
O5Bz0INqBbQZd2cttWd3X8cfSqpXBwxQUL2UDL+ofTPx6dxqSfpIMNGikQcsgUmOtFad6S/kulAF
a7s6uBM6TqGTx0GoVjU11ThdHKD2up/nrcKXO36oo/cjdVrClVzKvOspNng4Xes1/9yqociJsI4d
AJjxd4HrL5tmePlOc/6TtDRJuvor7xbYowzfQ7x1h1DESMy+4jAuqrVEQ35ZuzmsIYYH4+98Tjso
CdlYcPq4rXP599PVMHC4uiOJEc1O/px7o/OIaKMEBZaVXBxP9hRwW2br2Fd0/Gt1jhlN3z5DM7IH
8Ud1Gr5dNjnHm7rbFbea8mUaKbsS6JQ0Bi/UD8oieKlbdc32AI8rkhg33pvU8UuNsqJu+McyRFwm
yiQq2ryg3+bKPRcrun05w2GlOcaYmegynzkO/XjpOQPFCxTkdGb4kFd0PRz+odYK0qhBIapb/8tz
pEpXwb7at7MPG33XeVky+4iliNq++ElEkdrCM9CVuKfLOGF4RB+AYfWU0Gp83btcRRHuAU+1iqDq
EtYNosYRFPgzRHfpXLV+lRY32Un646Je2jjXRf6B0hQ75B3COpGoHMl4noWZTqU9vyVDFP3H226f
8jaPAm5l20meJm+Jyj3gpxGfk+1Aty77pe6gYdvpvPVcQgMxPlL8Lna5/xSho7j3UZabZgxo4wSC
YUqvh4pxQWknx19xdLeWH88zo/JkTd1h/Lw9UWtNv7skEtR5nKheqLmpJulZ82eTS8hUXcdd9DXI
nr73suiQTcd2dLeXFdgBjhMYRuNinrr00XVSUxvTgwdOKDo3iNS1F7gL6Z0mhI8NxVZkkFPFZvj0
xroUG9iQrratRSzjFiJSIwpPMHX5GfpxgEbqVkwKtO/abq5/KyV5iocoMZQvL3ejQgisCgSemYNj
R/1VycJSExaPVL8vUYaToxmDCEumkj2oxNZZjEa53ZWEtBlJByBsD2hpGs7EwxBfH/LUQlUA7C/5
tLrx4AKtpZR7DNfEqLgY61csy0YSefYD1NxTwFPU6ONWWzAGIM+npzPNPmOzeUug5BpUXHviojhZ
l/hekmT/SxVrgFbDe7TMOqIU3LWiE61yE16C3l1jnROhN/Sscx/7QFkVJHhjNztGW6EzlVo9Ixa3
jFxLIcF+0Pg/moza9drkFIyAP2XRlAfQa7cDuFqpCAxV2/Y/+tfcnfHcwqmK3cszUoRBlUCQIWlb
LSZ6uO4T/MN1+5cqZr8oU0ZuVkf0bUvmeXMYYDA+OsPXXIIONsC9u5POF2OfiA4WBVvB++c46z3R
wiM0u3H5ZfBnNEU+0kmYBu7SazpXfjdP+LpIu4k6WC3cZ6afy1vZiVXrqdGdHxHRJILDVzShbFnx
oe3YNTOwOLz3fjASIKOSpLCT11wPAshBliBwrprrxPwlVw1y82xyAymnZwUb9gtdjYuOhlsX8Oq4
XOjL0rjhJRVbg7Oc9udStW5ni0LOxQAQ13jyFRvrpLlsrl4e8Dh+0e0eCsyPAJQlQYIl1+xBP0D+
bLdUwcOGs5SXPImePHAnl2IU8bk5IxsJ7a9CyjwxjWVGyKlW7788kiyCgp/PIYc2Yr6x9LAtxt63
c9s5GU3h2uIbJ9uwOyGL9mH1n1XdawcRZlS5WfcqGbl+bk/uE1zX7D8XILn6TyrxQ6b6XJZji3fF
3UgVdKGAnqLVzkKpsZBL1OftaOckePRccR36DA/NzOe8l+qqcpxfTIRd+Yk3XGyN+NlzUPOPSQfv
aXV423Vyo31SnpXlrbEGEbct5qVChC71fvtrxQ6CPbVf8hd8kQm0g+PJ2pjpqPqEIoJgyFOMvgXy
pKXVMdR4IXWxtOJxX3w/qV2GvcyRkfB2vQBDBUCznhbzdhwjCO/FuxDQoHTSVyeSvUyfd8MAfaBC
1uTpIYrTSrf0Hh1Q7ZfiAWqK16yqZZiHIspCqqlDxNTdnoWmmmSGARrQzs7zXCxIvcGeHFoJxIg5
qGTBmCLyUKQLVmiITokEIwFBhZoQxD4T5cJlE0Oi1PT7zisHgN7WzDjq4codggMU4aIMzsQufPCB
EnrS75edgvbg0W0Ojrhc594ofHtusqr8eQPFFjTHFRyJZ9YyG3MjvC+ARqbo1ps7KOc3Vag3KObj
Po8gvLB+r2mmle7ed2JNpAPvv1UgMZkIINMP/04OpIdAfGSrJ1y0YC0sUuV8Eb7NgbC0jeYcTgkg
GMja3f+WDJ/OyuK/rhZuO8dNYlucOLFM3pPy50ca+IoRBI8/V7ZhJhY+OAAW5MMnlizxrzwHLPik
/vuAYaVLrhZXJ1oXubJFnp+sHqh306DY8n6hVd/3FFGJN8NYjxS3GB7ZzdHzbZuQjPZF4b3mXeCC
kRA4doZBnIMM4h5mrl9EYm4cEnIAPjoC6S0r/J49ORt9a9VG+Uokh1OVdmfR9TEq+5Rf/irlyGCu
b5C67wSfuPrFGva2g1ODZJwjDGuTQc1dck5grm4aGglzd3XCEME/tyxj7bD2rkKOTfalWpG4iVMV
VUalPAcGtC83JfvUOBMe8D/tbEAULKL2oS0+ZuVKo9jIEzye5tTCmgkMP3CeiGovPBJRoD+Jqb22
VxXFaOZlMO8bOu+lqPiLCtzVnHxDFt0UOmr5r0LPLfAPH5VC2oU/qCdGzeFJmbeBuoBTUGqyQcvo
ry7q+fHiIcjGUcBCaY1H6qTqL0X+7TihDru6nTSC1Z8PnpKnccvQNyBJMoqy0Av8aucIaPsdX7Xt
67KSyktY8vZa/fjyP7xvCMcMsW8YhKP097N+8Jb8uAd1dNFK0TUb6DA/yt8OZeIU5s2jiTpRRAcK
P0dkHETFfJQBl0qadO+1vHmvRjnosKNu1Y3wehsFVfVPl1Dgi1Mgz89GjuKHYj3WDokL7Xemdwek
PiwSuRL8BtkSJOCsZWW4r3gGJieYLOFSUnrAmfK1voix1WwY9+sA9o9bNhlAjWnmVgnoAiKImdjp
USWSATTrckm1CJSwVSPEU2s51IDwhjmHoTr+RwXkRrdRtB5vjp/nBbGrGEHpt1tIomlo8vTwABGw
e9k0H/wXEz0NFSgR6vWEAOxncRjOCD5+lFuErwAiEQ+WGbPxuFa5rC8/Cf8GzoPUgGIt9UrvraNi
cPIkv+iqs+yUJMEvwd2cmqY0n6SJOYqGI9Z82uyvgzEucaPJhbqAg0Ygbmf5NR0fs/U7c7P16wqj
fa7Lojcayh25x447AZH+AMqDJkxl8PMQ2E4KiXJ0CSGgwyJxYiBmBcycTkKT6gpnMAKM7uJFFTMv
GW9L4aL2v54jh1eU1A+JBLni1OVwabXHpVosKIaOZ9G4jJCyMgWiwoArXVs61cKmZp5l8Emc2jTq
lMF/WzrWymzY+xBFlKfZBNdB+d+JIbW2D3FstxMPdoIscpCwKl3vApRvPtHRTKIwtMCh3rv+Hs+c
xfFM1Cis259HfHTk7c3PnzDOoidm2E+nVmPUlxgsx6t1Q28UJz1r+/rc/ktqtkZmoPWzdBUOnxu/
PGuyb2yXtQlDac9OBHVnw1saYMyxdrLO+driZL+7WEsU+dyOCqMbeWKBzqj2k7upuxayY4M2G5W3
Z8pjmWT9aP9hq2YC+nZGPxKSkPAkIhc6zLIxVYLDm0QQGoHdxzt+2oi4OIqertzZYneh+THQnAw0
yYqezFsCJStZk3zIvppuRPOoaBfJ612bLWumskSepv+G1rykXpSdU52VI+VC9yoAq0Smx1Gkmdpt
e8Pf59oMMSYXcw/nvS3LzgpOaPBtY8/GBremdEm6uG7d6h+7/HD/g26duzrB1OmtyMr7F4zTX03v
fVXezJurRXfQhUc59Z5hTXbDk7inEtmBu3Gxf+3oDhcJSAzk61ib7c77HAzb0kQ+RTa8YvUdkC/s
I0KVpsquRMNARUlWob9LxNAgdh9f9mZtkYp5or0G2u3Spy474PuWBH0Djxfs4i0FVF5ZeslNUStH
3KtllkMjYE3OgEF47FFiOUoDmN09+mgvY6XiMel46Vho2PFDOxGcAjBLTlrHXzjJirfbmQl1bpyc
DJwW1mOdKcr0t4TWucX3YAMozOwcsftBcz5ADyashBOXZOgwu8sVJBCIUoVwE8aYfXu7o7HVIMJh
2svWyVYb44WKcYEM1mAPLhXN2zffz8xXilp/Bo75tBabm+WX8GRXf1AyR7TrXrfQuF2ezA+eU++I
010zmORwnK04OVfczfa14Q5PgGfhycXS0djOkk45L5GuQ3tsAH+IeVFMpqPIJSwZTq4uYsRi6LmM
ZLhG4SbALNlL3Oi7Yo2DXnAUKldCMNT23k5fGhCcpyURkat3TOY4UktEAIW42rIKfpJ+g2eT9KNn
QB8eVE0sz/wwuWohGXhnofF307iFCmj3JgZesXEUdxg85jqiQm4HTqUbawd6kZulrYcSKJDwbski
0mrmWaPF2551KJgKiuxbVbe4pRMV+rNk/1Y+mVwkgXTYkzaequDW9Jf8qH14vff3pJLaST3xco7u
AWpXV5oZXYFAA8xgj4TWJ5ceVIQTWWnWcUhb5BijhIqFaBfskeefogezKm8HpAPKfb1RPus5tzGM
2aG+HQNeJaEbkOs/NWwDBdEHmEvJx/LCCctbqJJpinWYWx0vPMiZmBk7Y8SoVA+yZQQRSyd7yVd1
qXFFoPTNKbtLya5A7HTWx1RorwpGe5/RFkLdw51RThdtRhVkmWfBAi4I43ELl0edGCp5grF2MSuN
fC0S8FarnYe4g8Ylsix16ydSf0lDw98SaMEa5VNxohJ6wRI4C1iBY8uqnUxNtt/fQgWGHMgfvztB
5Qy23yJJ27s2HUl4XAOTWzBEL0uTDkhg56hzm5Ru3a/Nq8TQ2PPcoQ6NheZ7TOAx5vHv5ilUUDmk
L8Krfb8JPr9N14Ws2qFCLzJ8KzHcM27BHS3yBFFQz/gXNT1YFqyhlsFAgulOGRdIbKx6ldwD6RaB
IXXjclVcqzZ3rTqjcFe3TyZRBeRHhunFe4vfH5wY4fmCkpVOgkvBu4iBoXM+/EsMc2S8LzrjmpgI
ZJ8Q6pipCQpZAX2zagF1Eq1NwDHbkEbPwQ9lkIPISAGd11BSxOhgyUzPMfF9LwJOpt/IAaaBnvfg
zWnP9EwrrS1I3OmZFqD0jfU3CBTCjzkVz+Cd3AUFASWuM2pmJabq0DUpOEXcoUg+YAHinQ8Tmejy
DVNxULTGbGvYKJBHwb1/IMr6W+gbRrkcFqqp4FUX57rZLt/rzDjILMKb6KIQRuePa/ITlxfKEOSy
lZTd+2/0Tu73JIYrQsPPY2VX05UGDVheQTOXDkUp219+diSXylEuBNNyNIjUFiI20h/xmugZat63
DtjfRYmkQs7RXf11p2o+iAKNnj5v6C+6tMUXQ3HvWXHkekQyeFwwp1MReJVirCdQaw6fiFXqBsVX
WZ5fJs+1H6CPnmT6eFgTmV6FaVqiFngoKWTtR8ZRnP970qlxpXflDD7Z3yqDbUfe2OyyVqe4EwBX
fr3zbxSI25ZLFCyfj38njvb4FreJEW5gOFsFywrFAdRSs1Eel3+BNGrLlLILeCwWvslsyD8WQF+Y
V1p1dMyMHXZalHpP/GmXi9IbWL/X5pbCMqJtPBfTBCy8VMHo2kGbrJ+x8g/m9suHcSevI2R/pvPH
PXRCkEhMeNg6VgfdrTUgs2zq8lZKdis4ILsqVxutKK0gMcCzfIwXSjqxADhoiah73gpr6SL/iiWT
VwPKJI/mUgNoj65g0sCzaJwDovfFCKP+nn0FQ/dcTCFlMdv0AcRwTI3eNYJNImPWzYh9yqbQ9Rmy
VRVHIdfv89zOtBOBViCEim56t1W6UqDbgOOzrmD6miWIUYr0CPifG0ZMz+yDTW5XMCY0jnfN6XqX
nxwqF34AHgt5E07HHra9z0t2WvGpZgZ2KNVnM9EFnr09cWOUxkZfb7umKJEGDTX9kAj+tDl+YI2Q
+1ugAMFSbaetQvSDPSXmeeXdvE0VkEdKekpWO68XmLyVSmDGhvDOV8vKVlqYS6zpUspnvPqxJd+H
aLieodFkwo608bL1dUqNVNuTbRrAEqFmI+RVNeW1HreZ0tTVORTtDEp37DTkaoMG+F+xRPUw1iaR
uE9xmny4TeucTlIO1EJ0pkSbZ3XxsFf/QHSQzufoyFOZ+A+iioDfQze0V5LbNFKLuC1y6Mj4pbH8
rIhzgFeo4dXE0Dzi6kNnIhbTsymtiubYnLF64CYzJFMeG+uYOXCEd2Kc+0UzQuvR0ONhETAUgz/o
0sFj10MhZ8jKl+vawGO7BpWN6c/vpNiPT1i3B7DGYyVkHNuPOamvUMmUUX3bXb5S9P6fsNiuxGKd
0FyJ5bRBt0rBAobpFKwU92K+opZxNPAyk6MckvwCjtYmiik4cL4q4QFKcjkcv+9jz/Dnlw/TVfNW
wn10OvhXJJIUAGR6EzVg6L7QzPKNWmeAWqfMmrr8Flg8rWgb2UR4ieIvDifv9k3cKYZ/UMOjTVEe
nFIl2cU7y6yB30S2T5sjv5f4FqzWtvd6eH1FsA2SvtGRXfej0I0Zp1zPNqsyHtPBrErlTB4B039w
h57Yz4y9UKNVFlDRB9aaWoRnvi5xClZZ5DtZswtr8ApAikypMv1y2vwEOeTBWYS1v/BDhLkb61Fb
1utFWbd+6pWugkDAPBFK3jka/ZGZOoK6RiQOYuvHfLO/uRZySf6mVg7SxSiL5TDw8mSAJ40fJJmt
zZ22SpG4FTKHS2gFKL9nlHTDdkL5WEq3VbQvlDfnfOGqjjMu+93bJ4hoP8uOKT/bnlK1/Q1vu/5B
TxcWdVeGfCTrjrXRSBMqPCLsm8BLu/fvkcVoBfyoug+NyxM996wuDFCrmxDHI8Kixhzz1SSp1lue
SBPMgOHnuJoWaqOWyARws7EplLKj4Bsv9b8MHuJ3AZT5lxffyB0o+tQJ9jsgY7L3IdOsN6dk4HjZ
WeCkSdJUGIFaDKrAJhEgAaUfI/dbgzZxrB81BIAi7TNqIzVbDPR8Hr3MUQz9ftAAk2uYKsxgnuEi
jaQNnaV1fN91apqObgAKsUFzl3wqPcoVOUnC5wsNVqfryZhtB03O3epdA+VxMpOAZK7dxX73k0Hl
SwXRlVUmBn2mzzhzS8wNCmb9TFjeMNiNRuQKzp1deentdpopljo8GLXJHAgZnbeDeMAi/4wl0SMU
nxgVrhgxWEVdrnIFhqBPRv+3gTaaJMQZqQOeWgW0Du1GAi7KBg30QQ0xnKi61EHzuqngo5TklKM6
0L8skgTfyXjE5NJ+a5FIgbYbWmgw5p+RJkxOyYvOZkHcU6e2JDUzpq+EJV/wvbwSTEW+iMmgbXcO
Nnts3x4eZyo9g2DXRCm/qXdPCqeHBtwL6WGEY1WLLA++Y6Bs0efpn9Jj2hjc3TxpuRysgObvwnKd
UaOWqq7klKX+wuEaS2jDzf8cirEMOE0U17Lcdccjuskwv778R7Wq07r8qm++7S+CBXc6byExgR/c
UdmAj26I71yRALwrzJvKVeWkAVxNL2Ho8c9Rsq3tulLypJLMQ2NmlymRo+vM3uuZRI37TkOLVWxp
9bOJE9lkRtAjWei4AcrEPepC821Dh78XX81vPu1QdboRm8eU4FqZDNeIdjRr/44LBkQN+dhd74g2
5bOOceLZ6BM494R3FxLpSvqz2Pzw9p5ReJtx61BxdBZzPp55HBrA8uAkf5XYxwNMwIe3Hl0L3Y2L
lJXYscvSNecvpGLEzpmzXi5n5I0xQlB3cmB6/e817qv5w+g7k1X3nlGgQom/7JelD/nURz96UJRO
cuRk+GTXglRh7Z8CQdgEO+MnT62z0EMl6vrGsVzDQspSnuV1KqwI2wFL20CdZQRtjSb5pDvHZNXd
DMYwFlZKH+yr21ApbFa+tvm3lGaj81tdPafJ29zmU8Hyc5n8AW1j00B9KfCvMFjVoeNO3/RmQ1k0
0oWMrZvyCp2xuX3u/6TgcXQNUlUnm4gjQ4bSGKC7SGKRlrC8tkjUsXs5m3uwalxcscTTLRg0UR+Z
+xVlXhX46zg2PkbeZsWgf445GTEDkiX9HM5t9Ce1DTFfL1LXtPxJptaD2aTAUTpWyFNroC/gZcDH
ijZKr2+Ss47qvraQoP0RWuAWtEQUX/tihygs2UXfx0YZBNe7mlW8BWGmpxMhiQMPjuZXdCksPQBP
5jf3pQy7aC+yl9nQfk9pXiSAvvRf76y6hKduB0vrO5yKlZKMbhZaZUO0XOS9kJtrSWer+aD2dUU7
RJxFgIzfaWOHDxZxbwmy2VGAMgaBDXibrhCSLlnX/NOR1a+IuZLw0EllJRuGLDn4B8r8Bh9T9r1X
ArxK7ozYmBgk2oHD1/BTczyEUfxMpqcK/ms/bKH4kGXr2Aa+JSlSd4eyEQdp7wXyJn6xIVShoqzJ
zocgWmeOARJI65iY8QN4eRX47o06CgN4Yy/S9lzOODCZbDHUqvJgqDKZO+2rM14ihEx8mQukHX1t
e+9DORGFHJXGGnub6bWGSlW4YELgEYa1mv858+3thmQNYjCO01WTP/YuClvJkIXfX5dS0XQkuqUH
1uDN7OujpgXS+p18jcZihrDiplAQouCHHb7A70BaZxIIpw6WnnPdUbILCJud9rCONs0EHq9IlpFB
DcguLRCMjlYWIIiRSt1lKqnXNUeOw6B9vnkrZxMwb5rqWv5TKu0z5KB3Ec6/v8sDZjFPFR6vtuQ7
vmi0SQRTkRwUXSrz4kBPy5xGYIZzN60OBaZ06GUS2rHvMM/Dps+d+S7xUZcnzEfPJDufBtAtug9d
FKc3npstg45+0l/Efb5+I2SD6ULDixr+8WZyPWXPiiSHr5DRQIzpyNHVljFWGS3gY0kqQEXiFB84
O7SfRexTa9KOzRJhJexeZuECsimkdvEVDbvllMkIaatjCEXNdu5NqkEtvyNv+Rc18gqBBHsFLCHp
++ybbY5F65h6yYi33w1SlszjnBH4xkEGMiEt0TteiI0nnoa6uIepb03bKIae/B7heky2G6rYfmuX
3jG3xguwJ5RZt7/Ag20dcg+WVzj008N7speeOzqzvrduz0npsX+Vq8wQGcTNzapvZmgCgQ/5gR/r
rgh0NXZmH/OGIXuoBIqFmyKIReJxvcQpfxJbe5thCDpi0o1IMgJ8mfey1oahXQfUZBGToF3PVX+t
Et1PIWfZgskL1igvex7AUD4SFdllHQVDm6UBmZC80T5fRm/53MhP+QPS2X/AALHrkScJnIRvZhVb
6kfuGXOZBAqwTmOfx4XgTWyLY00e8gNPckM8Gv8YN3xGkuV29a3KSjitbvANBEEltA19mSi1Wqw6
PZwFkdJaOxO4s48Ym90kPZBkPzLSv5Uz7hSyjwBthGmbXFLHH5T5xKo0bPcXGxvNOlNfRxYnlznc
vwCtAVinHNxme1vny0Q3MvG0MFPQnXFoNm1K3dte4wYu+ItZSiznR3Je6qAxPXPPlPWgyZOxUIv0
1/d2NqJr5xC7pWZ3dTf/d3i0d1l0+w9ON36V1hJvGfrTdmWA2zd8QUGPlnsmNva/VmcfbOog5SjQ
ZxrEeaGoPzcDDC1Z8xqft4col7sMjaYB5gNXshwy1M5YA+tTBWE/z1dmywj2Bmm7KYPHLFDgKHuu
hvySgEbcHUXGkon8z8e5bBGEjoHmRb+9tjQ7dPnzkdVE0IZb8U1BGJ/0yoiYSQ9L1HBAjwjwNGH/
u4wM2AjfR5JoTg09TKhXg5do7CDs7lnnqP1yT5BScz/QXwcfHjKhb6X4IUBYYjP7dOORlcdg2CKr
gT2oWYmBMcfapQqVtGR9eqzE1gUfIvFcxJRqU3Z7zzEJ4chJh1zq2L4NchONjHi7aArnioJ07miH
RQnz3kMr77k8i4p8S7nGhTQ8CK/aqMoSHhOs353s/H+0SqkKkAav/corFIYNfKAQKIucBKrDPXvD
dHhHmTDmJFQctSclg25JsO8MjTJph2JesB1+VHPvzRzdTVpCnJOWk6J0ptIggZWmDozSv+T0I4oB
UBz6tMPpnEf1DAMlPsJug282FKpQdHXA4j/zOYCbyGArRq7JI1lsEP3MlUI7W7sHM9DQwLSmMkKy
VOccCHD9XQVXZxIVQqjMSPO15V7Eh65E1AwZxtk8FWOAqBwaXzLhejYJsVB+6HKQotEPKZenNH6C
dFjcS/bKzhaoOM5bBPf+ysMi7/cmu/LVJFIeJ10Yu0iMb2sZz3QaKSHSfnGyspFrObK0tihmsY34
hJp/2zNy5rC+q+7Jzf7mDqF+rfWZISbdXSAX3Bz/1h0X7r047wbsHnznbiLMUf89rbSr0HxbjgnV
wHYLsxnl8srwxKT9+DLbXjcfMPmglLR849seVQNNn66qTcYa//0yybbiJj8yaJQ2m3b62pSoVL7y
DkW/semJT3sXGs0Hg1+GLf3MbwEkEU3pyR1O2wBHXSQSSq/tszzhytAWlITRXy2tmKLkfBNBXFsH
iBKexJVJgQl2J1ljJDTrhbadcg8YzqAwf/4pv5fkekyfOsfuh05c1oFusgiREFDvu1dbKScCbQII
YZYE1AaiT3LbhVyQMtLv8kID0L6RUkKJKcwA8GxqGzCyB6XfZV/lRtnGDr9emWBVxgFqResMS7GY
vgybylSKN2QJZWh+OFbc+Oh2s62W8Gix2rTlfSfRMnkDidiGvuL4AomUNcg4JH5rd+O0dZkj+zgx
a5Ik0+KrOddL4puCUF3W3QVlQDCm2t7Yzti0Ld0dWzFPoN9S9kxJz8JRuTpp8jLhNX4p+qSoSWQQ
g/VHCFD9ReypuGfSaZvJ0+LGTKEqVb0pvvpk4Ya+UIC2k3oT5Jl7MMFnTztkDW8olqd95vFtX6v3
BG/qO3XlJTYpgom9SJKEhn5h08uguqQnCeik1lAvQgTjmETwhgLxS3lY/weNrQEeSTqi6bYDthEv
BHA/ALYOcl2oELosFVnCemiqCBl+rVypIoJ7YtNII4Xks0UMisrKYd+KPU84zSO8DU5cpTyvXKt7
75LNSciKdMptdSs6gtWDSkTil4Fu1wc3oo8CU48uL+9kcEAvpg55cAfo+cYMSsaRdFmM5vJ7+Ubd
Fm4+o9bxduBQMnDDAfmzBFV3KBPZ8PJK7NyeXeHOz782ijpYF8dPzYpxWKVFFBPTSMHOT0feyJrH
M0favTBLrof+o2EEV1f4mCVPLV+ZnrsIQiACFi0uHMz/zp53cT63Rh0jNoLAIRIGOqUUDS8SwJ+l
5GVyn65Y2fQrH38XxVUTBGJhI5am1hDalFY0wFrn8Q9uy8wfXCk5nAKJy4OZXSyW7fhwNnv8tbBp
xAkcrokirqzTdr6BZSHL33PpgwhJGIKN6Te4wbmYwObam8lkXAc3XkBisvMTlMbLxzt8q6uUxrMz
ElLcDHL6FK+X6NrZWFxlcXjIfF7xLSttU3qKWj36Q7MKKABWc/Ox0J2aWfWgY5QCpLuguKibjUXG
+GSgZeVLzb4Gz91hW1bQB5O/9VfRU2MZpzl7Ae5OMipj0WRfU4Pa7gKBctlv3rhPhLq+mFz+bKtb
SpN2mhJdew5s+bnkWjKWnnJLfYznmNymUPZYvGftHPqOy/+PdeRm49un2wPEkwdwKWTYfAKRkOH+
xmgZApLBdgM1fuH547n0lAIsraCKoLTYKxHiKuYDvxwP4ZjDmr4NZ2Ibt7E+RKBwZ4GycE9+UPzQ
8YnRXj7o6+/AmtMfY7eLomc8GYa/HKDqD7N0wY+bng7KBV3rrcZh5ixye9UaoBHQ470JSlrjrcTB
lvPVpOmLuWzgG0MA3Lu41T6d6OO6543N8//A2knYMJBmoxTJejJQravyrFY3Dw5CvPX7nU+ldWV/
8BGQzunueLwm1cZYIQQTno7NDl57xN/AJKsrBPiBoJCoZDb6XjkM+Z0uJoHuJicTOe+CfAZhJTIv
qA/J8NWWw+in9PqxgDJyvmVicKaRqfMBMSfff0hlbBk+Xe3hxEts3+1crhL29dtLHri9u9mbjrsp
DYTmnV1c729122wOmC+5d0o7kfChP86U+ioPCQS8dUiJbdKBCeoELYJPFPBhGLdb9QLU4hijJqX6
LCyYIxS0yURJkDRTki1N3m4bz741RG5Hv398CUEX/gDEaEM4czUkuelFqMMm3zKvOWzxgRSotSE1
ZAVGxZGdlPysveF+KidDU+F9WWd/muX/FCxiRmOoievhgxf7RAQwqwvzBExZBlP17gWiwNjcODDb
YS5RYFgEF+EhKH5nc8HDLKsEgwazmR7adX+bZEMfbzDSVXSQQbUEbCwHHhJBB/wlI2XanCTJpk+p
K5XrBO9dmF4O/BKZgTTHyrQ3dulmmatk4B8le9tgD15DAqsqo/47YHPO+sA7/6/OvaoxVJvGRDS5
FIIJH8kqTxGLOFGrMyTT/W55Ni6DV66UQfH52vZ5OSvGNV+GpPqnxLIJsvZuX1qwsvm/ORI5nCna
DBQT+RPhbsfKP+cesM1lZBJcUK5HnDUWNDMjD+2R+OkH8xk5n3LuqYazClDWE5xBPebT9AG7VNJ5
dSTyqH/1txzjPKLV4ObRTVQAIzkYpSal3zYaCe7F/zwsGWHlMT/p218VQTnkHul5RUElNGScG2rh
kqGz+73h/DpqFoLVf3scDWakMcuTbUHxlhi8VPGUvuvX+4c3AvG9WyDl2n/iDJuCoOudjGc29hdX
bFXqKPHXJ6LU7IpMtnmjnZPIEtbwfNHtlk3ZjIom1NY4P+kUhTNyVPWWuKuIHDq21wS1JiysPmI5
IPGG0lFoAcyWlaVkSaPPtrfkuJnlGb6+7yZJu8kfZDoEDEh4kLSLNqXl4D5Yy1y/llFxtZdUOvlz
tpket7bfsRaUPxBZuiOHUao4WWWjL2ehYdmLUFEoedfpXA00oC5mGLYj0mkt+/AxWlhufFxmuG3c
FB5JkcxQd4cljVDHXLnf81+oyrKPGL/hzWxVaoBkRl30e42zG4jWiVRPTNuNKtnTBP4maeJUg7Pe
b8komqU2FOz06xb+xZ2XOP9NkoYwzu9tkedMjSrb5Khx+qyCP/3EBi0EC6UmmOiVvSy/CfLdHmc6
lm9TofZ4+2qq6WFbJbShd5jNMS+qrf924yreBDxUer5cNCsR508qHTDF73iTsbbvic8xd8eyNABv
rhcjW/4QjNqTZELuQchdxkd5pYtaAT+4CY0pcoU5yEF1JTwOP4MPpETmXhqvZ1Hxw+yzDK6Twpvo
RzroQTZuzmuNeYQT7G2fdEz6ZoXdaJ5qq1VGUTtBhr/AxZgeGxKHRRbEUIVk7JXOkyIeYI4UvXLi
mZB+DufpEaYaG+tQAh3RgfwMSz2o5GUNMcSwpieFLRYy7su4dD7yD4cf3m1HRXnf8C0kRaqq0yPQ
hxqip4x8GAIxVbAFokElPRVwahL8sFDlQ1CrLn04CBkeg8jDm+3z6A3sgajDIchc18viwxqLy0t7
zvlQ26epreVT9mxu+RnLNMuwNZr+bYijlfUZ+VoIiIRCqJZttBnLOadJUa8287cGpT0/yfbZw5dp
/3rcb2RzXerbFzVrvG9GPhl3CmwJZAwrIDVKMd5U2PtHoBO8UlZfVktxbcLG+c5b/ivs8THNHizX
rE2HpauJUf9sgyXU/9IPLu0oM1B8Zvc5mHRWQ/VxZCYEBp7GhuSvRllEyzu6kq3/mq37KR4x/Qg7
KtlZCd31CFxuMuhGpwSpxhtrJt0rvdWG/IBKN3b3btAz/oilOdTEp7kj/ADLdf3KD6IpN8YfFHva
nrghoPuKaKsABGhytBETeqI7/hu/NAf7++/mNTVjPy22U1/Yq6YOKqGq4z56vd7/+x5EQaz94hhV
kjszkDDWoO3rxsAiNtqlG5p1JGofNIgFWjBMPLNBvRSyNg5FcLd6UV/Mtl0i3SXQAVtWZmV2YdV2
ghthi0z06Ns9nftov6ClhwQAByiuwzMmTEU+o6JSrSqbU2rZC46NAGigdy4s15NhiTaNKCueT1zH
M9jpnMlpNza3TShBhICABT1RCZNljf/1bT9wsdywaPGU7kzmSEoeT+fzfwzSVx1DGMRrWEP1yGy2
Byr894iwO5iftX+CLc6RQiPEhgJZzR7gK7nP/GXK4InWwRociGe87EdOVZbkxTjd+OD+DOf6xgC+
X+3jc+bgU0M1FV+/ZibtGk92Fc6+HcZRP31M7xcHjUuuMXpuhvCJI7sIrLE8z8vWIJRo8H8nqmGt
XIJtxXg/oVDuMejfHCmKxUj+MJ6zCFqQ3+sponrvCEGNX6onp5plxa/LhqITHyhbGGjXERYnKUrx
sBzvalbApKazd9xpkxnjTXkMrbi/inDVjHlkXk5KOStLZ2qHYC9wE5BcNglDF85X+OEWpaRfOagI
H0HpPZtTIbX+h+/LFzLyGYu0HqBfcVwLuXHS85uTYsiiwaotY1KlJ7IUOp3N1qwU8v3pN8FMuhGk
lz5Z2YSYsh68rNwnsAQVVdxHnL9pkQHOfOJ7ym4s2l/9TmacLAimlc558EkdKODuWYMVAIU4G2ui
um2/dKp3rr+oTJLpTfLl35oIoLU5JuDdCplZ4wIX6wn53uysFWknejT0j8oS7l41qkM0PtiESmV1
FDWHNkaYldKsG1tIQYiQUoCyK2QcVYd1MN2zthwvrY1DG0so7cl9YTy1Beva2go4OapPVEkbT6mE
QWqzVIzvEJo/gJenWM2ujhR+stVTdwhbrodlgNBFniWBpItZwu4I49hukTe55cBsm39M/ySXuOG4
exFHnzUWY4MAdD94r4eB+BMvT7FqnH83tnimq9z3x/KOwOFMOtdRBxJNzHi/c5cy08rkc7jFi4Fp
ACPZCQbMc54Tn3TLcEp8CpstoLdserQSdXy/ijwXZQ3z4UQae2yfsyFkR7ieCGlWA9QDTXlebIpQ
1JmmruKXyLD95wbZUGIb3XlKPoQPTEtm/inX5JMEjZLEWIqd5WkG++MRwXAefCUfUchALm3PB9DI
IalLtsVGaOXf9Gy+tN5wYnMn04Tf7e6ccjex0lu1Uvie0pSjwtEkxoxva5Xu1XgYCkrlCSEJst0j
/r1a460p70CcGt0dR1/hVkKJyEdjXGp1BQv9DsRRpUNCiymoSHbTrbhCaCJowQZpyu4GGeXgOcBY
pN5EVI3XrTNcBUhRq8dq6lxAzMmoHe1RFPu0w9gCxF1yx0UiiKqk29sZx9Yc5Zm+VK6RXR9gYpK2
k/xbHhktSMWPUVdokHCaoBMTB8CfbmUQCNo4x/psjOi8GprBgHuaMW1MBxem2HCRYdpAvZ5OpBkw
Ic86RK4UR/Z9rmSVaOqdFVhRWowisWLRzj1100gC9I0WLaZ5xlXrE6QYTmGnc5TDicKuh2QwBa8U
U4qFETZU3rpP3UeDdddyOMb4BLAs9/DoSjM1V89KgSaFr+aqhz9bqlBILwMbqF6CAIxYkcWIP8NR
OBaPl6cL9zGPdyFHacXwjazmO/IZIoN8vVTfLnIKhe+yXQDW0xx+JHmqSousG4vjS4S/UBxXIvKT
o5KgJLwXaumuYCz2rsk1ObofuxWJ62zVQIe2DLgi5RFIn2riYOBgM5qtmdQvJiIIN/Unj26X5Jl6
eTVI2+6M2cBoKrU7bQrRsi5VdLh0PYZe/JQb6R5OW5SgQ30CYPRB/Qxp9jrTR0anHeMVRJBwQcdG
SMBfNtTRTDTbEP00+6BC3akcnwCfDkYJ6gh9CvPhcae2+pwXp+kF7uD1WsZK3cop7NrO1fy3Ad0s
Uxo4+Y511bBXeX4VX4U4sYr0nkUr+aSArNhVaQZlmcL6sWyEu/ceYOJUaxV5vjyeNojgptBtG1DN
ivucAcHcQZ4OzORz7cKypkxl75QsOmRsHmHBddnItGRK7vu27kPGk/fZ0V1Ze8hlCFyqW8D5WCuq
bY2X0rIyXiqM9IEi9ne7YdmQhI9FrRgDxVhsf8JAcozZoVtxA/f8QCADAmgGdAbM/WYGggjdc/lf
1Vqc9b24DJ4Aydyld2Zo/C1rX6yV3kPPYCkFF83g+lu/O7qHN8++imKuNKZL1Q6zC3GaarZmFzX4
U2WkJMmmTEtGMj9NspzyHFpiYXJFnirX5CKqx1ajdDQ6oi+SSz6n1TNEMZnrcQR2oNc7GT5ilqJl
cBWU9cRnK30W/yOwmB1A+2TtXobbOCTomL+nPo3b7yLpXCCXPmQznxwg/VDQLxvJ/giawLUUCqku
20UiX23hdn6B8lMxHPe0Y9740uKazJ8KCXhoDWhoXY/wFos5F0IqpDHHSzTGrhlQcSlYEnZ8fFr6
oSs+HSBIy+LyeVK1VmUz7LWwuDCJnbuWaxMFwgGH8bhwBidjNQuS1KEw0V/hRJGz+drMUiMnw+4N
XiDjvUOJHjMLSSN3fpx2cP/82v5RUYdI9NGdEAvhLWjkaSvM+/UJYOSEkAzvNrxWiiW8Pu+QB5EZ
X65ZfaKFt7/NUMKVi5n8q3NyLt/mfaBpljIVyaaezwMLnSfxqg95EP3kq8sRj43SGGcxzKE6JV3P
shj2LYalDb8sSbCzWEE2ap+uvX4rEMzBV6JMIeXxZWZXjBE7OdoV3NOvxJ6q9IlHvo0VzcHDIYLC
XGNo3zQWZIiFnKqNYUBzJtgNH7fMu01p/RkIw9juopbFfZbTuKQLIGZ9JNXscdC/DHYQnC6Xxv67
J+smznJL/EyF1wx/XL7IZSvcCYXzCSIWmppMkzLAfd1stNZX1JcHi2t33Z+rJhBfbyNEB1eY+6Th
pwWO+fR5Jkc++PlO3bHxcupc+rnuE33AiOpPAB2KlfHBTyU7rIhRBsZZSefMl51dWLYQNdOnqJa/
uEWzzxiONNgO9KnhTMBB03/TUC2oPSXYmAy2kNxpj0o8QkWlcm7mCqvES/9NwxrMTwx8Bkb5Q/5s
iGcpgdtPPwp1d3l8ElgWjIuqRapqvjo3Op/1TJb2KiIAq8qVIrt/8u97vBFNejha4qmXQvOLo8u1
IdH1BDbBz60xIhBek5NtmrYFvEBfcG91M6fwO5kaKXAl5XLntN1DRIiFTA2x0xBpg8FdqjB/eoP3
HS5Wx9c5LgMdsZqOps475PLFr1OIrak3Uc991u6sGCV+qq9x0ItXW/3GB4RyNTfapdYkawvNJi+e
30c7Ux4cTOuYeqiFBSrojEgHNNyxatez0IqvORtHGUez6fdMbaFTFiGqRFP+p4JVuFvAPc3oNtgu
S8JJ/PBepbdWEv8Jd3Rz5/ZMiCSmfFZgVMvzEZStbBwAlf6KTqofQNS2UaY9cMav7oR6MCHZ+jiy
8g537NVm23Yrc7gVcOcTDJtJgk4R4uR2FtUyPYiXaN63WKdibKJJ3uV0o3GjMzaH12YlDKEI2So9
tPuHd8lCkM7+wPzm37tanCxbI2ewrytuVi+mrz67FJ1jS+0LcAwdYWU7800aytjM0yA+w3juwecI
903ZQODDwrWNxVRm0rZacEI2YMWIwlJv7Uv3gRY59fNf/H5N2c2Wfo3mFC16x6R3s8jniLiKZRPY
v7NrMtVGfMZWTf2tqzi21aFdi8fbaZ2Ettg9vax/iONWtazI1G1QUcLuPvV6kO9GDf34UQpJaEQG
uVZZrS58YcA/sIRU12yUNA52lJvdhPDAXpscoTFXlhA3jcZSGptvfasekT6OIuFbMZsa4bTElFjK
8IF03UqHa8/r7pTI/ITQrzU+8oXiddCYwDc3SkRQwLFqGybXzVXtewRXCezfKRFYQpl9louX0gJc
uWYeojGV8BnDKzD2ycnnR9Z9kor6js9AX4/9QmPgoNES2wXMkSnUrfGj4Pqo7uI9tfNTNqyZZXf6
L01UxJx6tdsPVtaGAY630BOsXjZcrtbWZCbxz9xJ2epNzn+Tr2lxNd8hsyzmbks6mEav0ejlxAoV
X2F+ih6DZfjt8LEXpK9xloIaGQlodv3+VHszrq/80rCHuTRjqvok7cXWsC7mj+vjO51oSKaIipn4
MGvXohuZIqmZpEKf1tC+hPFF2MSnMMiVyUpWOqFVx85ackQIGZ855jeJKnhM9Lp6H94YBhJVzAQl
RqWgn57i6/lq1SsiULUfSLX5oulUKs4qXVHrz22RMp44adsIE4UEVAfv7E7CTCItYJee4irbuUuF
lzv8VaWVCEFCwmd6Oo79AZ8MYwAMmroMpb+YyKzm5zc7nMOF2PgRPL6HzinMnueaDcwODIi4gklj
7PbO7hFGIJtI83zNsUuMJO1m++ZglFyhyLAeGMshZmh9tLLGYxURTybKEanWVMs6/IiLDjwHQ1P6
ZQlOtYyhc0g+mOFi0vtGBpHOwcYqb2TyagFhJpPPR6IvUBLhmGk8cj2DCKkhjs3QKtQHfAjgYNjB
AsiaZC6ngMTm0o61M40Nacwf4ePkzgTc5uCLK4fkeqa7P2hWfSxp5Ovbnl0fJmpbA9osL0uU0QNz
gstWhJVuPc9HXK5o+LmEfWztuh6mtt21Qddwe8gtFq1J/tK6WGsKd24f/hCWLbBrTnkHy7Hps/TF
X/Ta+en7WG92XB4gizWpR2t2LPZqbLtoULOjoRQaY6qB2Qj7Ajba+uMNB3Uqqdy75ySXa2XTVmNs
uiCDP3sjApniAiVr0ZtNpmEEZ+DLEP9i8PctfRItSB1MfEo2vDY+MdvUqpHKxjI3DeHEwr5XIsDd
H2g0gX+u7FUpDwCsAkycBAyVCYZxuLb0JbADok2anqT2w6pmaSjdYELovd4oOKJ+qi67iQJdEuJf
PYRIfH2ziGBethLl5aGgoyZbFruzKdkVEnYDzH7gzsh5dPhYoDkxNUrshtwyubZYs/5rbH619beh
QzM1v5UFdj0ZQF8jE8dKiQliyfpHgrzGEqXVdkLYoC5vyWlhQjuRU/P1nDXSQWMOssLoTUgI+TKg
IFJNJRyuLbXRwYTVglxuH8al65UH6E1yZADxyuYhxr8A+z2PcqdhnsxireG6I1Oq4FZ/M6sAiFgg
Bs/VgiO9StaTMGMcUFx0VhaHp97LA0h2lrjlTR3YaBXg2eRsgOS5B3dpo4w7jW0UR1pZ2099GJiC
qXdD6kes4b8jufMBqXZlUXT1ZurIXk62TWPz7RVPssl5US9XKT0s4IlPHzjWi4OPU+JaV2iwCXWZ
rt8LVksZjX9oJaykz7fAbMoBLR61WwWfcDUIXJorLvrw5p35tQaWeF17QMoId47zeHIzud/zjYF4
f/Z9ApTz7OjImAoPDDS2zTvFQYsnO1laxf3S4OVPGPFgvDg0z7DY22LB7bm3en9ciqHEUm3yCw9e
DjpujEfqXXW2Wqpq6UEuPHaqjmpSUMfduH2S6KTa5bC2EnWny+yYGY06u3LBSWI7wuSXlPEE+VRq
KkHXu/jhi24v4JMEDgR2nWyLrIiJ0xL9dEVzvrPPHfDr/t3ec4E3jnw+UKcnd9SkCXHhev2PdeAg
L38fs1KqqfM9We5GfOOx7a/EhWKeGz+7yyt6GgCeIt9tlTpiqKzaYNpU4nUt2LIbIVIPRAsrfnHM
JONNFb+ZFrqu59RRI9e2cSk9IGZ54FM+3aGuCymCez5LD3wH+0TmSfs9mr95gy7burcIpDeYawGB
oFkE4cbdCbAXc1YPfwZe6Sd1q2vfsg8ukZsDF7xmA/OP53JztYtldVcQd8+m+z1qJR/m+9zpvnIo
o1olyS075Zn/nXzT0RmVO6xc7COgnjNacahTpJBSovV2bF9EbxxGzdeHXEkuinIk37SlzfEHeWOX
Rm4FwpsGMEVUWYlUBLm5PP/rINpd3J68z0p653kagbvIzT58zhc8eZ+qrbYG04TfkxldMAsdg65T
3Q+k0pnWF1kRLSZYc9zpi2WXaECW6jXdMra/B5w9tEekUmFyoLuuux/Zd7rGQE9fuidU205sFP3D
o+42KTkyYlkANnyC493lv061xw0+n2kqImIT+DnPexucPJ7TezcAwvhOeuAH10NZs+KVYzXjIRqC
N+n8VPFunggHSCASap1b+zZr4Xosl4bMjLA8zndD96oAIU7UEv5v4vnewRuRdcjYzGT12wvMhQps
5uir8EHLIsDuNqJzoB1L+QGOanosgWWHHsK2GblmqyBUxVeOP1eefehngdXZCKHTvXChNDqvfiW5
k6n2DWUI2ZNU+w3pQftEESMRzPwtqDG3lQopQ37aDQwrDfYnZNwTif3GLctQsWX9i0trdy4QRF2s
zB5iqJ2HSQ5de7EH27qVzKf7Mlbf75ybneV3HwrGyPl38/z4UEtQF5fAiAv3FbRx+zGp8q8b61eq
LFzmnfo4jcAtjbVMFSSXteF/19Hroj+26W+LW9d8+t52N3QNx4xkEj9n9YFSxkfmxrlMILiKFw5E
7OQ9KRw0CB0dbDhoGq5mCmNlqsEy/d7/rYqYeaRZ62xmcakRCzxEaHjnSOu0MLZwYIpDg5mPZ2sc
5ZUDvf7U9t7QfDHa9riLGbbGJajF2twDrNGK8Et3Z1LHkc8UWQsNmRkLzDvQWDPsIDOjkuMBcFBq
DI+BDLo6/PCJX8IIzIwm3m8L5hjTRa8j1JLxlp8gjG84jOVuyadkkA/PidueIcDNgDZp+Xm5XuRO
xtwRKgf1af5bNghYE4aLzvzq4/aMOs4i8J6igC7HWWR9jn6cVVeIuTtU5wVZZ+aXSl8NPNWufbP3
6ZkLYjj6F81sowr7K9mk6Do+lrrPygrwAu5S9WYbOr+GsEyf3ezbOuYnDwmEU9HlXl+UmWt4Btut
Htrwig8lHPlQ9/1WsqcCtrgDIjEnGq8chnsxJSIOBg/BDlJ7OnZVaPwEilJ3//XOI1HL9n/tBo3M
/AB+dtkM1h18yw45BZkGgGTGsNCYQ9RFEj+fpHsDnj5ewVlcuQ4ambQ29Hx9AXAICUGltqkFYlPt
ikfA8h9S0SDUAnKPzOR+7kXGpflJ/yLjDrD9mZbPjr59YhFF0daNEZ3fqs3wAdcVBOoSWP8Imnls
U4vdOjD7nl5vFZkVDFEMvM2De6hkYK4OqBsRwlHvVnHtyEBlvoGu2+jc/GXx1xq9iTTu1zymdC/D
YFu1lK3+NivbfkkywhjNltfNmq01YBy0EXPyATxpSvfjrj4AMxFXqXqxW/4NQRCisT+1NBPjKZZJ
/7mLtloT/qhb97iQYdFFLBeIDNd9Bk7BfszErIUhu6bOSBvNh4ingjVJ4IP3kjGAf7og8l+61KVo
RnHixLheUUDY35mfDJh3LKc6T33bmHMVlyYIhs8CJNl/DKNYfJggtEIAaSMBTQCtLVHk5r0Hdxq0
pkU7v2r+5v1+1HM/hEx1YnJXBHmESFuHsUNfvOiJDAd0AR+9/Rc7mBTk6OhrVvlNyx+v2BGRAcDB
b6dDxy2NFjuK5asBKksKmU2h+L8/Tc2iJGYB52ng+HqI3cP+o3HuWjJz9xCb9Wn9mufaj7Qp2xRC
U/sdRq/kzfqU6VtBoOXEsm/Kt3vGyWZmys2VvZVH+hfMqejO4SJ0A9ie31B1VtPVc0aB0QGRduQd
H9j6bwqm77DgcNP7LElEIJfPq4g8noVMdj9JAAzh24DstQjK3+o8ZsDxr+mE5/i6eOKNKjGmsf/G
oIiRKveDI5LPFby0l91gb3pwQ0SmgRmu51R98qHHIxyzX+ZJ506K60Pe3pxHvC/2e6ORqJmmhlJj
0xTHMaKV6N0IxlP7OmVkzmIjKlIlIfyKtMk6Trf8hmMxsEyrc0HYRVcom0hZXYkhhsWeJsUNFLPS
fQ8eFWa1YF4E8gEOvhrMhDL3hi+qAQyHzoLuE88nJIzDsX4du0KntRXDNJOTzYPYNr/TGkuVjQj7
7BuUGxSHTNOHub3TtA4QKDRedK8qpiNaughsems1B+RZfEBLzwLQHQk/VVJ5IcWHqoH2HIBqjPrC
5F+YdvcdC8CnwW2MFjtYNjpLT8xEbF+7F8hkbFCmQi4gc/2Vv7txia9dYDMQaMoXlT+aKsQD0RNX
ivti0G3v4dgPWy4SoHAgdbQlHHuqNaaOsOfYp9lUh3HzSVPfa5myMcG5DlEANMO/B3Hr3p/eUaCm
IcgNLvGg/Cj0u0UXQzOg4Jd90v07pPX/7J9z70mx9Gc3zqoV4f3e+8LQBB80pO19jWohveyEcNGD
w/35/SWHCBi0ZugHhc2VePj/XZi++VKZkWtNBhTf5fpDaF+cOqsVIzLIV3pCU30caRXfvI3u05K1
nho6pnsrqJyYbrdbsW4FrhCccQL77xW4xJUAHvHQkTZS1HFcLuhxJevniF6QAg9Y8acOq5mZyX0z
Lq87qN2rmwmjKgkbv6kaJKEV/ej0lgDarUzclOIZKvnlV9KHGCieu0RxlFqG0TWkFZCa/jNLFL6w
Lr2J/K2mR46dXWjcNIUmDQ5y7UfBffpVF+Ahs50VBDnTOlPRMraReoM/J46tIfn3CRwb8ukB4/AK
EM0+1xQQsaOF6EK7QMaDtzh7z627TBgJj5DsLeOw3bLvte0qaqQWljPUxyqNSHolig4fXw45UYMZ
aHr4Y2+S5U4uplVsCfH5C/MpXZpB6FHFEqo0+thD0Qs3fkR98xUIaZ0ULxVfV0Hi+ArT/ejh5M8h
wFPDVLMerlgkhIlHq9rsAvbRxatKBxNud6T5K63V58jUlV/XxJfSvTJq5PTIKbLkBqxjUkYASaA8
HQ2+3MmbhTecJLX+cVpauAT67svGSpM2J/MUW7MocSPaFZft5q91o6Zur3wRb6V8WrWxSKo7T7Of
n7/f3wORsMx1WfSjtqmu+xI636zSOikYkSBrpuHj4CF7ZgNB/EEKhSZZcWimWgJNvyM9ZmrPanAK
SZoWBO6i3RDuT1CJeTAdXokO4BxtEi7/8gqfw6VtFwHCsZREkkDW22KUp7mH1SZ8uT6yL8XM6y+R
HEOks9LaBKSL4gPMjAAIwIUpLx6z3BzQkeUP6EvmLgPikb1vCvh0TtMUhrt8l88te7oQEY9GFuid
OBvY1RVmz5C0KiM0VX/DAU4Ozb6QXpFZprq3SHz5QN+itmhiYqFEGCt75RehzMmP4dRKGlakRWnn
8+5G2wAlFLBBGdM5xUY7fAlAc5Y9liHqlNcRu2zOXD87TmE/kED73pgLafxvhHSDadBO1Use8mLi
kHiCvUthI4fV8uCBhEA6R+28PaF45UBQtEAYa+nRbx6VysJymkwNI+R1CM9JSl9JOrZiYlSDUvae
tyLnj4ZhqWmAewX3T5n3ADJCjONqEMTyrOLlgPm1Czwj3WjRPae7AR3AsLlhnhmkd+bFlQpfu/vV
Ai589q2qOEL3ro22Ki3s8p+ltR2zNbTCBZoF3hf7Y/leFLEZCOV8wW+D4angBv3D0zpCBWzeK+xq
aQr9m439zFWi2YOop3I+MAHVMqTj75pZ4sLJ1P2eAhNWYFfgs+4FGTygwkYo1auPflUZfgen9mG3
/5j65Kj81H+Y2dDSen6hC1cIDBGRg87rEumZ5SXQHZSOXjgLH12UL/yGXSTYXwtEXuJXs+CsG5Z2
dXcF+LR9PTjKplJkUvkGkHKAydCGPr4ehz0YuntfQQYtRLSwvWi8h2zLybTNMJd6md5fgndn+jo9
ouXCQqurijuaqu83oWaYKc4W25qpy2OhYu8kMupofI8FPrphqe09ceotBV5JwWzD0BToNmjMutki
SZWu1o8ZqBhamQg8jVuLr/CgSYZ7kWoYKh+kbY0lWJhBQ4QOPjiC1EAY3JHRKEmxqsMjteqio7m9
kG/28p7e5mtGyGZQjNYnY+R1kV9TpnJadeSVdImIMrZm3nj1NWRqwHw7jWjq6y6pDJLOhzFSvOwH
PHaJR+xM4q3GkOhC0AqysyIch/f0U3yhI9lidUJBDxB4AmtnAL0cUtgeqXWseBNW/LDqGt62kj0/
biArixYfDMYS2AhB6qKnlOl7kfxTl1CnQ6frFMc+T5os2VqbEe+ZJUc3A6jZsiCmfpI4fSxcrgHt
lhLpp7woVmBI6alUrBHSm0W+mJsPneaMpgkwpiHUHDeff2x+KG/iMUtaTU7M/D8f6G9pv+VFGoB7
ym3Nuj9xFvdOcoOpsuKhYHZEXQOwM7M+X8yH8P5f89L9pFQK3YQmZ8LmEYYCU8wh1PwP61kiHvHT
76OYtzb+gPoVxZ35a0hc+DeOZqTTMx9y+z29d8+hXU7rvdZdpggTErM25ufIFUrM1rhy3mn7jitr
fgM4zmNxXzsuHchZMNrRW+s+g/uRx1k7LYUIg+N7TWSc3MrLfU64t5UC2vKtmRF49PWm6ONpvJtV
46M0gjExkDsAhRu6F7AmOrPqkkHR5OuGZmokJRu3Vd23C2F+j4QSQlKF4ou+7QzkMWl58SlfTfRN
ST7AevO837kqebCGeSWOt+2aXSYb2Khw+XkM25foJjEMNXsJ3rHBEwj3HQjXQHEKLAR81zAx/k+g
5qm/U7chKndrV21E9agcfDfzdSRPqDo0YL5wNpTFGLNYO+tLZuWzjl5nHTjBzmCqFPihbM7NeT2h
ZkUm6kEYyR4VkqXmKoC/qy2fo5g7uv+q4x+YvZ1b62Iz5YPNmjvhv5UprL1XxmC709Yz5++iNXOP
v4Cca6bvOCiwyb76XMjBfejEvxg1wLNNeIhFKf/T+LRNb/CkUKE2b8APHImIsvoTUD9mOS1kGva5
TA3xPwhl29FBS3eEEQ+B68Rkt5o8nRf+WCQvI5KcyBNwKsKyjaK8erWBbiqqsiRHee5/16NZRMbN
asFNjW68R3JPODJIm4Yw8Hcwuokvqm/xSygHt7UrVsMG084CGeKz6lrFnFB5NnYYyDUX9+FLWnYu
8xXv7THJgxu6z+vt3nWJwPCk72eOGqSmjRs0kQ8ulwzLnkE78LcYvHWmw3c6sxxaWopt3poHf6nT
/QGZv33Y6VTYRH/4XMzJpxCbmM54GvyyPLNYO+TDB96mHCvSOT8z+X7dKl9kram+i4mSEbWADGB5
N0kodsQ8UYz1eOPCiGJl/Kj7bjYpQyqokd5iYrB4mV4a9g54Qq6jUOy81qL9F/en+tpMznnekwAl
99kBMC9u0QDcDjSpTcKZr6JaVzNzW5EDiX1dSSIRyKcBzqOPKHCwdz0h8BiY233RSQhdOKTSPXph
2nGRMok+x2etRqVA4JuEV8B5weHdNmtAliXYKEuS57S2X9rYaSyzcch0g5K5kb27qz6NAakdtrSx
LXa1nD7Uzxe1PNmGNljnOpXRKFarHDZNkuhypxVG8SihA1IphGhzO6IQ4gGzgXNiyr4wWR8LIRNi
WiaWlqYpdMJ5Eykj1n0HPIlY9Ma0lgwnYrKsEQk0VrFu4QoHnLgUwNWrZbNw4bMkJXSRuBWl2Avq
znIs0U0F7hEZ+wzmhuS9uSCt5mAzxtUQlv+sASggMRIt5kHGJr8Pe35p5qnD6ppvrMO04PiWkiMm
bWqg0F6pIGDrKM0ZUr4+8HsvHO//Bynyf8meAr0lDjxDMUpuuCBA7R0lIsS1EWdNc6s88VjRs97Q
m46h/MH3wDhGwrX5yZIwRxI/vbD0kNlZdOLWszEk26645KRqnfQND+lX201t6EQ43IqI0CIBdK8Q
3JSxW9wBkmcjGHEOyamQ/tfCgV6A8RLfT0xMX6a8kSPVeixhCvsG8GwvQCg3ViDlJ16beDhwT0W5
zn7oP5ePP023rhTXUXSVkxvgcvSmnr0cPfJJZhdGsD/fqfdu+ylGtlNBiN5BIlbsfOubtw2qBF6g
smcbzW+yUXL7ReR6ElwxmUC3kKey+J2GWvAbPpgv6vgd5XFFbABmXZmvotTARgjQwCxtAQXjMoEs
KEPireok8QaJZ9q2RdgQ1kK42CwWAeW4+ZjvuUB0koR4ODswd8VUG7jGqqD8DPIP/gK2zKwOqbhU
MI3BpV+o++TNXnnhS4kK6YP5CBu8ErbcBOJFVT/Xi6qsZVl/bRqOPMqIumFALPqnACu1nyPYGgwp
ayEJnqOGVHJqJ2hux5SXx4mLO5ifu16t1MVIALnQ9GHRrI3j23NaT9UFP+MMGRzatfFTgt/nY77T
IGkkZqyPKMZCX7AJTvutMa4oXhKw2vAX3qM1s0gFZS8N5hCUnCFDfxHH/3plaGhBP6PE5CHRFosI
hr+IGIhQMrwsaOIFf3E1nVEOTIfVZrTFnSZVcs6QKUIDkabQ5gYwzwQcYoS1iz2XttDFl4BfbS5b
TqYceAJ0jDMKNTkBT9iCPifunHbwxD8JIS636bB2ddw6UshX9lUIh9Tr58TrVvA/442MPgRQeq0j
ymXIFcATY8SZ/TIILdHElq1YIr9xDV9YcatoMtWv6MjbHWMi3MUJ1fTBDqzLjH4ivytll//H9jvK
aXF6jJOuJri/AUKWNQHhCTGjndPzRbOw3/Hr/Xee0NFlwCoH98SzgiFIYEIRlPMgsj+1egA4f9PJ
N+X05ppx4+rHzfkPdxIohTKCZ1WmAvWi86pYs72Ukc7gI6/7oWUNPQ7iUma0NiZccap3dX/oQ0M9
ByMVdJAk4SaoRAs/tMOTO6gM0ESV0IqQBUeg6Yv9FaPEOeKBZync1U1QSxNXsS8YSWyp71LoVH2i
4K3NT//EMi1pYhst1yAMsOWWjdgxTG+OcsWkmR0q5Rygj0hVEbn4gPErNetPaF+5M7pYO0kDnytr
L4kfNQjsACShVrbc5gWW71P3DEj95Aa0KEHL4rV6PgkF9jSr3qpsI90EOc0kKHj0xZkAu0ljhHlf
xfn0U7gzev3y84UnPfyWgbk5+z9M9ruwcSLx7onad65aUmeZsNEUG9knwGDwZljwdDPc8Tkf9Y4H
2MMlY+CaT9iV6CdkaQ8Y5gVzwWlH2XPhDarvvPuNzAI+DUlRbVtXfPKEYVuYGMZ3RIv36c15LO0M
FeeHcHYgMyJzDcdR+wtMxVB4FIJV7gHbHTuV76/yrQ4vZcPABKzjY775n47+fYmJ8MJfkui45KjF
EcsgvqRPAkNKUcvF9n3MrTMwIs8bdnarETdM2+gQdwpOL6Vwus2wEca9r58+vKVRn5iU5I2o8gAt
hV24UkCBt0C4YufUkwSywSmk29vlOghQLFjmFuR2X9DN+laHy7taw+SV9Bcp/PEnRJAgh2fIpXFV
pbFnkXFG43sfiRTcLFma09l+LQU4ncw3a+PwH/qbRIZSFyNB5V3v1ucflHYX6ISVH5/FbkeHKerT
eTpCTpvaf/VfuAbweQu0SZMWGhnldZQy5+7Ag82Uc/OuiZXGpp/0bL89mwIKkp5W10vrOsyYbJsO
QwKFGEp5a1N6hncp5XLlcolvUTMruCJRr9GYlJI08XV1OSR9IERgL/g4S/8sIquFADu6Ag8PlZjE
HtGhljMRnvhmZEir02WiQMX6JA9HZPqMgKupceEnC7V2oBOsZ9XJVcdR0LzMYSJurBbdP8Ykrz7g
w/s8vdVsK7m/nfPKEEwZ8iYsChhs73DUI+VdaFp+W5AKKMpzyXJR8Hhf8BdsMtq5nnYiZfLoWPkH
PU0Tiwstu0s1VousqgecZyVha1l4lX2q+kTR2VwX2663dj9aEX+hro25fO0D0jkQRndjiDSQN8DU
etljrZMmekCA4m0xxZQ8SGR3/zl1UCIojJUrnMVU4p64zUYArCZmM8PKZjqj5NUpvPLMlts+Yujl
Y9zthmNp5tL9Nr3EVZuLNGULHMarwgx8utLrS3ycZQUIW0ceBSizp5jiVbyuOKlytjFWFLn2Wc+C
s0ZhqOAR61j2wTJ9IX1mUVbfPqTxdMJEQzv3/l+qa9dTIedReItBkENIkkElTev8FbnRryu6Yk53
+0Fgb0csTLw+/HqXdzxVtpOw60a1AIKDTxCjZoGA8ddcz8YE9El2cTrx0iLGEFfrkIyq7sx+MYgc
Qiuq7/5zhj0QMnGU72/4Ow2/6n5SPI/C+7v0oR6xNYjWGTE75L/Q6CN0hfJZKYx2h6bZk1jym2b0
qEVqBBvefT7zO3NlABIUN4gaYPKu57UfCA9h1g41/HgWwNbubYnQrXLpnA2v6twINd9cNY4J9/ny
OC49+4OdHKVCSQBBQt/9Hv/01HhEFOmyV49dR0DSe89wTJuA3SQseykKhFZ8MbEUd1dNQvHQ0jMN
wbCTqm/cTR95p4RDeWlOxZKs6vc9sP4Vg1UmuiOuRi7jq8cu6QiKJrvfCe852hLXM1uZeQ39Q84U
kH0Blvh4g1v73VlIGIfipZVkk2ZH2zEAnH2dgfPNMYmr6/pB/FVJEZwZCI8qC95IRW3HTWq+6Qim
hFDGE79zlGmMl1lN+hwISr92zMuJqXVftpaQ6cxsKXUFPLIOaFfrMHi0dbqJfTkRHA/UV/lZ18VY
cSK1BYr+0L61JrDTTDW1kjKegSrLaWrg3nF0kUkI76PfcnMZ8IsTQ9/avU2cmKkdvjz9mKZ1V/KU
HnWBVVQiZDe/6hkFqf4Yw/qcAJwsFgzd8AB70Sxy7aDuBCtn/U046HdHYVkrKqI0PraQjmpGTez9
M/nh2fSk/CZ8/mNvqp/NC+ZcdesdWUqSbBqkTyBP9y7He1vlYF2idSEc1cGiwIb3BhXivkXQSk2y
FShJKGGtN+VV560hfAN9CZK6k0414DCuTX9as2ujplpb7WWdfK6dOse9fw/J/RKsQVn2UBy0bYzy
ad8MUrxqCKRjmZtFMWcdu2O7e62tQhfhkP9INswsJOCPY5T2cVUxg88gcDcLJw6qGNikiO/vtqKX
NPbsAgmWZxXMVENFhzLILrTkJL2iY0oDsra0NWGLcjiLlkuDYQDAP81dNu1tO5NUjLcJZidpKhMc
GyWt3N7FZ6PA/tvBxFa8kX5mZGXUbWPu7fxtHzQhrWI/apGG43PfnVfJAmak8vuk3e3jpRLt0BIN
v0oQaWpe8Kuq6+A2gYwZBvqTwcd5UN9Wk7IIkzz9RwPgH9yAtYi/uuT1j31iodYhXXph8RdcM3uX
ecgbXvLAbTipu2MUwu2bHHTHo/AT3xR4J1ebra3vGyCav5yK+n2C4fOBuDr62pIDzqd+2bBJk8Kz
dZ6TobhKkemvr7I/1sl3HHTSa4Cs2PXz1tLSK/2iASd77Zt9cM90gpTvTx3fU6PenSc+QYqiZzUE
/MEf7KMmYstE1jo36caCC6jifuEqQSMLH0/vMcjAmib2EFWwV00NE7gQr5it5LOFUdXBnESwklR8
oS7HXscAhaudx01f4XtePK4U7GWp52hl9NOTcTbp77qDySTsHSTOEZPV7elZIJKd3L14NZuUnjoz
qF7rGu5N9unMUMaMyW4c4JfPeCr+8LGiX3qztx6WeQBKToESkhkGPXzkzTnL6OTMqxVmLp7PwS+x
wE/9AKrTFmxyip+N5B1DeJ7d9vrP7YqxDhbiMTM2kizcBSBv8rPAjVIVnWNgoqBFMDZxpgmwoqVd
SOEQRL0QqAzPjyywVm/DV0aEHngioHluU6nqRBABAJIYTQYhZxTu2TVO08x7azOxXB04YqXou+d0
NqB90dyRxVsq+Lazc+ulf6TEnug3XLKvbF1f87ZGNcNNYjYhAVx58HFZTZ2gPWl/FAZcUViPfFVd
OLcqnBlDuxgieOiuwbJMNAlvaJ0ExMS5WUYbsaVVR2sWTl4GZBBNFZ7zzIbIS6A4gMHcSsGMOzhn
BU4ECD2W3JaKGEZ7Gh9ofH/Y0XCTBXqQZlpArw4L7Bst4PtDGkLm+3VSd/n52LtSiT/74Cdnj7JZ
BWFgrXHk0CfI+uvq9Wc9RRQrfvq+GdZNJTrnGjMP4RZmLthLLmR7S2gENRJEF1XUcX8dviN11gEg
aqVAr8BA0gEp68Qvxvf9mhC3BrM7VI/8n2+XgiP2N+Yk8GejiMj0hqzLZLErB2Smcl41W1RYcoix
bOIFxZMNth5x4EMA1f8bMwBpITFRz0vcBCmwuHSYrTyv5Umk2yelCqz7QyQPbuMey3OrvE/tTk3u
uhTgo2cr8o83swd2PiSm9Wc0jTPZpyvQwhgbFfQ7HMkTGM1ZDpi5zZFXO0aGiosTMpBGkPBSktPz
MO7Znnh5wqba9+4nXqqtvlAsc7qpHvYa0JpuYGmQ2uEMt4VMKFGlvwt2xw44VYlWZTMHObIuOmko
P7Yym0RjhFXh/CiZ1/kexQAhMQv+X2o0UNOQXzNrA/++fHZN/BqJIP0KiDaMyVQfP4LdyeT5PKZD
6UTAW2ohdmk+zFvaqw5l0swCXS9ONnSegCxk3RGo3JzrpGSwgtTLdmPeTawMsh1r0bBQEOMSZKHp
k1O5ERUi//ABik/lYNTuLGUoDLhDkXkDxaaYSYpjeDZXsJJ6R4RSmMksQhUjG+2ZDterAB19lKja
KykA5wd5pxh3j9mTsGBZQXbOZWupe3nrZEHo5ohMbb2X6noCTlqG+W+4OcSBTbWKkVX//vEyZaVY
IRTGsdgKyqdSW9jAPrDM9qDxKf2upDc2ZKQYWi11VUzOZjatzqBAgNVdWzlV5FLSZ0vVlChFhs7I
S2hIEhl7Ez3kz42EOiTImq9LvKaWZzMTzX98sUlkjmxzj9Kk+fuZEMcOjj3ci1wg+dA7ntiJ32Vo
Cmo4d5DLt3LWC05ps0YxmG2vcN9o88ZQhhmpwQQyY21foPNar43S2gzFNfqnP6UqMmP5PhiyA8s1
eAtKTewTvvfmbbOVaKKo+aoHbF87hJHKOQ72jVUKt99hpnAZkGruLQRZp16clyscWOfY+ZpPY96P
RKa8DGoXR33Y+pH94Kh8pP19YLo1ALjgFyrKcHrS+4jhoesTI45Chd+EC8OFoY5fBC2jZ5SR9Hn8
fkhLZNsbYgQsPNbL6tl4MmzR7bryST707rFADWfeKUL8BXVKCbGwewDRo1Oo/6AYpMstRnRT7Uo+
Iv4NUgZN3IoK94oqIRLbSUFhiGL+KzhhgxyEIQCX8qySf028y4+S+IAWgvAMMmgNtR84iUVsVP6O
tU/mKzLt/gum5jb8RfN6hT2j5cC5v+SIiN2xQfOaDxmpowbTuc4FLMfynyv12BtYKzjPbWE6RSYm
84KPst+LDJVwJ39Ny8iB4TFCtaAMn4g/ZPgpj/e7Zl6g21mWJnCN9uYcWOr4ka2yHEUzFI0tqL2i
vuFfQHCxEvYKKxF4FMQJ+qrkCkF3uHh4+MNq+fFAzA7EsuPD8qt34wgXs+wD4OgKQ/+1aWmkn/Zi
cRH8/RjBWfM+YS/Is66qiZQ8cw+ocmnafBWJ2GKlMW2OCsrvyEh7FvZmLYKrcPgznJoeOPG9fVJ/
XvawwFs+LcDtSucQgacj5dLKEhVG2bBWIgf4WALSiM1OGksFPp/mjseJuag+cw5OBjQiocdfWwd2
xxWFVCdi29A8MODxkZfiziHT5FI8OwqXYeS6BQzkod4D+pKX4EIs13wY5olXHVVwlU/dAsbHcMV1
FT9AKRIk29rdHtgogAxWTMgkAPGcvQAcXN55a5LLCJ3QIaZ6PWrvLajy7ZCRtHb5HgPN6wOWHOV+
/svDxKs3g/Zko/eYc70ohhpXzFjWzTlibOT6I8364G27us7L2S5F7a4PlbU2ZUusoZX54qeUvkTe
9uX8DBB4rH4CQYz2cMncxiDkvlvzD3PFZBka0N3Ib3FaLz5qy2VQcpXB6K8Hf4EWA9W2GUFlawSB
1uqzsbxh3/Bp9Jequbfx0Wq/3L9d0XmtI80PHr39wTni+7ameSHspTZC7loqX5bgyfuiVt5MhGTE
89nQvMUxQWgsspj9Cq7r9szHfSgAjeUiLXh7cnoOwev7zjEGrIwuXSsJ18mND0IL+w6ws6qnib6V
O3Lz/GucGF3flcdp9FSkFKW75EpdpUmzNa6FtQz4vyDhNS5x+24NvLFc3Zs+J2zswHSPtHNBNL4L
l3JAYKp49rg0YEn5/0mD4uYVVJywD+a2XxFlXFi/JCXIaAmC93MkH7E9fV881RyiZYDIiJu4iB86
tUzsdZvDuQ4Gb8r1R2AfVQsv4KNguU1rTivNSuBkuWeVHV9zMA6L+W7jC2zBWkEkXhajCDv/bEr/
GQKVgKgftEcKFFE1KQ8fUN0yj5WZc3MI4g+vwfN+FQ+39faHqfik6kngoWZUEXkDr45VgWdYtgJ+
7sHyQ505O5Zi/2Y+W2xrh8CfSZB78RzHzza0FUnXe4PJjsIduoNpsVYKVPWIKxiWnNZp6SP948kj
+VR3jxVuSE075VaJaksMNnpzpc6JnnFQ/2T0SjwL7mCg5B7V1EtrB4LRy4KMumRW6tUFFgALp/8/
T4P2s8DOFck9315Q5N4vyzf+z28xgMyWUAuCcdKkx3z82pj7j3TymmLR5/IRqEga8HSVEKeqtPDa
zzh2V+1I749OkbFMIZfXluZsOQsuXHm4Y9g/movBGTPkHjzcGvSoiVXM2SHLF6j06DgkkiGXaJRL
aVxJJE7XOi7SQ1sN6UOtEw3UMWTE/ly2oFfGnQDXHD8d8N2CEeIfHLQgjWR4v8KjijxIdHENB0Vt
5bE5yiqwJL/dTKtK3wtgOiTi2yw+DZ2rmk+t9kUFdhbB1JUHJDt7dDYi5sphEOryo6j+7X/3Q2bK
hrENagOfiRciomkSmx8wdC4sMJcz4C3WInOWXXTS9SuAYji7H5gqURf/ifmwCxmyjw8JZ1H3bdOv
AfNUA0V4tgjAwF7NSBsujSn2Dv0TSSmHOGwWacO7thoNZfvdDK/SAlDrFYtHLGDe40CwcTAO4wGQ
GubKNRsDaha5SH8XCKc6mORTU7wt9Qx+3HgNRD/2NaXJaI6gnsXjtyRvU7/fwLQumkSOrgXO29fX
SFZN9gtjdE6OlP2W6Afwz/UezVvoNS5sPn+GzjOa+w9/gi8YQ88/XmT9j1HbehJ76paNq9pQfHCD
4dYUg9Hy75BPBeOUY9dk9/S5dzzh4bwzWx8nn1MeHxGbxNAFuuj9DqXBVEZdfrf0RYGefKOLkGjT
XgqR2sITUczpA9m9n0J1ln8oSh/T9Ix7CqHn7KXjpdPioXK8fVweOFLt27pzZcUgmnfIQkuMlkJl
6JuIakvtkXV/Bhsz17JajDJEsXHz3NXYVv6IiOOiEXW7iQy1TIo4Z/152b/mVEeiLPMljT4CCmxV
F8DN5B2BbSZYKPtWfTMs2cx0xMRKoXe7G3bNoiNY6W+bL6rSsQVdUQexP5veTvfRbbmPc3mHdYbH
GIeS7eIX9JtCQwwHhwA5LbhV+3guganvkrdnSXwcGfkH/KqXvuDHKKb1b806SnWW2ViHcJF2yvKz
MQz+4f15XWRC0rwlmeRgNNAfGDQaw8IOsu1uDLxQGF5SYY5RTMV85jqqa+QygwqMAo6QXFHyDK4Y
idl8xSiD9ja+fv0EfUqdAGiKuzy3FOrmT8+IQ7X8ILwjFvSuiQwyaiP8cZzAx982Hr7BVxZHNWh8
5dCb4U5UWmU5jtGfH2orhXD2OL7ttjx5yXPs4HWCxTKEWn7DmE30pjBJdfIkXB345F2stizeTl4F
ucZvsbNRETU3AQLqGLHSYXfoeW5LTcfOY7slfOdvSEquXs2/gZF5jem0sFEBPvpEzqPu/yiuwQj5
NnVBLe3pHqX5KkFQcPrTNySokefyXcdXlE/yaZ79kMVAEM7/V2dBJgxPDU7O0gIvu2QOBgju6Wit
g7ffHPZrezQZU46iVhWMnAGECRl3VfqJRmfwU8ZgtGjux9PaCAFyg4aNT6mBFA3FEwG9IdJuapuN
PQdnmE+VYok/nGZkNvCGF6G4m8ehQ/UzfJSpN5cltpEYfzRWJzK1aG/x7fdj7Hu9tNc6jqiPAn22
sjozj0NUAUd7bLBT8TvQibSakDGnJbQ9RYUZeC0qCjvvc2/HkTsvX9PThkZHwzqG5RZcG3T/QBIb
XFdUWY2GneiZEfgpl8Y0R/pX/9+df+Sd2Pfa7FDpD9JP/AL7CT6foMe5j0lZ5tCbIKyWot3PIfpj
2zx4Lz4kX/3NmZvMFA/eqoR+65YX5yflbKX/LLox4d3R+9APYQW79kWR9/eKu6n1AjGgCfJJ+q82
MAVLnrNCx+Ukb5O94LJ1TAWQAzCbLwlM0k/TmtTOSxAJEFmS13kdoy+rSY0IEcyHwGgr92N3RR9R
vnuYMQNWIZEB0TZJguEmYuuhnPqPNuI0rdL2HAqxEDxARol1syhP9Lq6cFlA4p1MsTlWH4T0BZXi
L8+s+K18kTSG45GY4f9eD93IPTfqmE22RzANLFTfOSXBlkNCr9CqhEcS8Ots1fCF4xlLcQz+UmmH
iNFKOgx93ALEpjFa0HmBhjMoMpoorozXil5YBUdpy0ybuqC+E2F9YRG0j27urTACB6hJyn48GJi5
i7FEQfqEfRUrkFj8DqH6jUNSqxXrrDkDVZrdh6Mm1UZGD8EAQKNznJGVS5/O8EwVDU6f1RgIb76o
8Y/G5kCBTb9PY/58WqOR1+sS5QLJg/MyTCbac0YZv+brWklFyxtAcPDiHapahOnAUJDBvXekvVYH
IUnfy/aVwMudRbwgAK4jouq9WhJ6Sk05pSO8aCbQOB5meaEPtEG6P0j5rHcZhg6vuyKHcbg1wgFZ
1Dgdr9U/c336k8RdsRXvk+RhAHTWbbK88pYrd8GO8qgk+FauNETk1lVM3tiHU3t9NmaqnjQoXsll
+QP8qHYMZnwXlmAfyIUttwvZNV+D7yqJJpM0nC4smpL1UY60vKaX8uYfArNDgRq58uhL+QOpesSk
kdzayNxZ9c+mjITW5MJipb6UjzhI4ighaCNBJ6GCnD53NkE+LZZWUDq/NOjkaK7Hhw63oyahZMhy
QI9xL4Dms1MyvzxToqFvxYsztvSCAR4ITughLjeYcPf9lWXYPTVtIiY60nFR1h7UnFreDQIHRF+X
f/2Qd0FFEKhZCI4yGC2wX1ygeRtz3+ZCGDAue43GnRU1/p4XPRZvcrhvbylN5rIrBubYEljFr8Xj
nZJqYxDMdIiCbpPSdB2MVusEM3rm9p1ep3u7ftBNW3lp+ZLkhgKSFMiVUQLsjeIASGgq9wqIRARI
auWsOm81QC3OnNOKKD5CvlMNCr02HAzHySEff1hBW8Vzj3YAmKYO/KlR7rhWYJSiZN6JEeCXf/Ck
ussEaGVx0MVF9QxYroLAfdo9UupBdvUMDqiEqa/bz15h157KjVzUB4y5G450q8Sy3BwIjaqhSrB3
A/7HACJo5KSXcp5chpmF0ZnZhQZIr0pAFVyV38cw2ykVb73zXDY3NPkG3yKzVhzwQSj2iwBYaRbm
PMa6Hk2cVB/kGZdKob5jRubStUtSx+LEzc8nvlZU2VJ98h+BsnOckEIAO2B4rEBIchJ5SFMvl4Ze
P62TVmvtIiSO2iqhODixQdEu65LH/IL9FMlyya/qHrPN3TvA3ipE/DiPgO7Z2n/cVOkzGB3c7pLB
B+Vu0OOES5zjHLMQaSd3UUG+2qm5AarfeCH8dZ9nBzl7EP7KVtG/4hZ+SOwFYAV6SGs/zt7ggCwp
ks34sec7fDzHV0QzhFiBFWIibkadPVqwKxbPdliOXP7uREwSCr3RGk7e93Xit8UZxYKGFhzhqHYr
FkNOstij/ht8eOBOSgabPJ91jVxzIffpDooRyQqMWJPPONi8Lbx1YLPDhR7z8HTQhPS6j6PA8GBR
EL35qfXoHw4sDQs/4HbJQ1IH3SIeEFQlIGAPLZJ0XhqJfKoSl0HRNBFUI6W6n47yavawqGq098l2
p9cWIFZCGRpyXXIeCLRiFi52v45cccrrdul1xJPS7wygfN1+HqU9snXkh/B7C9egAvjRbQpEBQzm
KB9HiGlE9V/KlA3/lVO1H5ggqxNK0rjDhDjkLGkKVCiKQZCxYMzc0L6dHkyQcpaEVo0ptRDT5ON3
7rt+EJ5V1Z3OR1mdihrL0wG/RGDSIzyYnS/PJ5qNY0c/pzZ8e4mg8S3+ud0gbmaRA9EQ94knO6Ub
aWhWn9KS1QO/C/Hp/VEAOwmif28zXJyM7hTUZmOwbO4nfw4SNxjwOZcLLMyaSsfseRapn/U+nnqu
C3YPbILvQ8QAMW7eBVeHGWj5Qu6NTZQVvTiMjYmOaqdlq7b5WuYlZ2trzfBMFPolf2g/wLGsw1Dp
Kb3gPXZT9Ng6oZtMb+7SHX4pDeYKbMc+rpjq6xFmjuO1hmMkrrUmSznAeid5WLaIxbxbv+Mn6fFS
7gbECNMdaARcf/Jtpgx1bQ0J1OPMJwb+8ig5gXXuln3kEcbCfxwNGsRJBfEr03+tCmQfDDgAG0vx
wrk3tKdtT/NTbwq8VGNIcJ//J94KOawIxGctWtcQEn6EV6MedkCLZB9dq9kRk3SRZ68YILtJN8+D
MS4z4Ts3mdp5YexsM89wOFJ1C+3d5FgnEL6wVJQPxnn1ons0vyaUkGRwKv60B/wmQaC6n9gcVH1K
Gceqw4UgX9EeaedCKITigj7tu+UkzzzK8kacnAoQOPm7N0igHVQvylAKk5egYPyfEqhdEDyPLgxo
RlsywtxdFBHVEWFPeDBY5RHjs6gs+prftt4U7BL9FsQOuLB+DjgTq68AvcGwWoTmdfTeHzMEXBpS
2WvkQ1i/uqptO8vrCvIJ+uTDGcv4fnq9Y4JMcjGbFhzqojwT3Uz0NIL4Q9q5QiN5NHIizBM0Cpql
nZswmWm9zUpgH6KqFxKbd5gDpW5sXZQvZi6jZlouNBBwsoZzHYoGngfpiwWJFreVeop3UGbt47lP
E0poWANtdTCx/OXYu1G2BERAEGfRInbd6mpqlR0dAm+ND8SUoSDs83UcRrpxU+T8tz/tHsqKb6Ie
CnRuDGPCivkZuJgAnth1hjPOBucQtMKyD+orvVncNJw6NarL11YzTwhD2ZxZ+mdq58zi264jbMtf
a1lQ1NE/uXko/4EUmdNXRl5lpc+9NHWKjmgvLHqUyWlgkIfsXZLmpUB4eVbhEiHy2xERw+bRJDfh
1xf8mc7E5xKDLrUXb1/s7UhxgEaR+f6VYWQsSyu25q7dljFumVutb1BqyGJ6MSfNKdAw7Sp7Taz9
jp9UzMheIkZh9HOZBDQRNwWTW+WY3Se3EW0l7Qaj8ggQq46MMTJOTmUuNqKuKhZL8Gfp8cGyE33O
xfS0XyJCUVZNOTveQM74jcwdj6mEgj0vMm9A+eBgr+/q9988yIPVyp18txtKPhbeqrKhXSN5EMjC
lZ5DBvp6DPRZrFW/Xb+AqvC8HPVAqHhEERfQk5wb3osw9ATKz3ZUiRlYo/jeFbkW9KWAy8w57+MM
L3nO1tjubLpiSq1/GQeyP/MXhMlqyXQFcDHxWw1zZkx4HJm/BCuIk8bTJ2S2l48vbaXzmw+3ZETg
kiKU3wo+AWYrjYnMuRKchHgNGkKQDM3QW8TipDTKL7mtYNKBCRAjhhgOSbmIwTxmRoUp3ITExQzF
OaCc7L3euS5e3T+fAAtPaEeEsHexfNCkEhWL8UhnBp/Mi3Vvs4lhb9uQC/4q/wQvPwCzD3uwZhRs
LCuA3wAWyIk3U0ZCdlksb42FofXM33raBzeLtHVUGVGwFoDb5OTdkvBKP+TCAi/xSOPerY1tOU2/
+7cRASWowaww7htnfijWmS6/UMllHKSd98c9mzOy+QpF9GB+TlDufNFR/YHPfTbAV1DuVPHKWtI5
SS3wz3/iLHfyNI7QNV8vdCLrnRqnUIkUTFoxEH3hBkB3JIzWXMRzElPZaTFPGlPAzzAVdzRKn3+P
udIuBJzAh2VYIit1ZvchkNgY0nJOgsMYGs23A3GaNL/uEYZ0KL4fc7RcuXzAUJcCc/5Bd0FH9W9b
XlH1GoK6lhveKBc6JDVIwQzx62/USkMswTSWIBYzRvk+mLIku1yZfIi7gfKafcxO6WqBkCtJ/Pve
i0uHJQdP0jHTiG5kPdqpO10+ghlg4hz3asxIaCGg/GqJCkAuD0PsuoHSzwhXEOC56Ebadkhqf63H
2c26Iv1t5ZYRKilqH/bQcQnnvxnLBWAWNlyPGnkkJWmFk+3kZHNKbaSxuFIlhKYWSjQ4BkbSX4yW
IMImXyT9+Lp6v7ThXMZlm+KVr5pN9YuS1Gu6yKEwIFurzaq7QVeITs+nXi19vOZ6auKVKz6ymam/
3YmeFyqEqfPRtzr8KBIpsS+ntxyYW0pqrH2KEPPcfUMo0wUKvlsWoa/lA6r4BsLS5OHeehSz/zsK
0yAk4qwFint8k0zZFJ7OFev84gYlmX8BMZQuFYAl8tzXeQHFJfAOL2YSEHq59U3YDomWfmdIaJvu
cXBo2BMaHs2m1WpqbgLvDztkRhGkedfVrl42FWrEKO1tAyKgXA1X/79avCkpLn7GDCtwvhd9hpGR
zm8hx0o5hw1SpltvF2qBc92qqk27/FgMsJlyu7ZbfLfx64SL/I7xGKA0jhRdaZ5TrqnZEu1IR5bP
KtBbPbOW4iRnmL0PfCBl5cDntBEOMR6xZEPWbmx3OcT522sAYzjj3d5JKDlvct5nsNhZ5bAsDgIE
NaZqZ8av8gZf2PgLaTdOxdNDvyop2gdYh0ijFVZ00NfatRG3TkD6FtT6TbLtdJSkOehKP+xU3Twv
glDfY3JedIDZynI6FWBFKOuns266kkYE9m1/NREbUAXnvAhjc8Q05CTCD8TtDOD4/i1jdFohGl46
6/mnkuqczg7IPejNLYxJWjYT+rAZawIxruspxASXVm8MkCOPyKpQCNxUQ40rVhO0/8F1QWe/b0hz
gKNpWm8CRZY2EX1vAHmevmvaAZYwQXBkW4BIgdtkD57N3fGCym9wnIlbFKZTT9u15oelT2iGVgN7
sP5kHjJockHUgkQylqzwB9XZdy4qW26TyBbFOp8VM3xICV6cM4xTDd5w4B5qyGuAqUQuOHO5VkZk
Y8lZATApHPssiJwRv1An6mYufpEsnowBPt/cIcaykxckOPCJYZ9rOqKAow9cNpvHkYjKaPpunMZ+
Iw8saKVWRZlS8IMwinc0MXLppDbXD6TIVi6hBkHS0sIXUflwvvw4m07g5WLRCn3+Y6s6RsZt0rNS
q0kqjvprgSJr8K4eUBbp7O8jgboMZ8vSt4NHP3pR60szOIV3znYDrn44NppaQCBVxltlJaAEfUxN
O9tkUbpV6+KkhrGJxVYcvAltzA9D4RIphsLK/kH0gr010Lt8IqFR1vF0+De4gkOhlAcJfB0njv1P
9DRsbkBOUkcdQZZVUva7OspZ1kT7OjWJg1Q9mgHBNnw3QE6RkB7i2/XMUAVrQI7D7s6m/gcGfgJ6
ai/Rt0PxK6ULdkhyJj6PJvJMeuiXltcBAo8kE28UgYMLQSZh67DYpfXG404/8+4YTqrkz57uKBOZ
rUIQptRHhmr6yIEG3TSXX/jCVcDOVlKdy5BqGHofaIgDrL8DLjM0RY8ZbhhM8xaQ/eMStPY5wtiy
A+JxDd6F8NQnrvlG9AEzlM0pXL0B6JZlI5BL3HTEZ5E6STJfAhmr3h6ptTMjAYWJLPMyW1Q2gWB7
1hxoOmIMtsqIBkFyz9fDXpJP2VvRKPeG4rYDi6ff2epj7lTGSIjovF695xOWyNYgq+otQqH+9Mi8
gMZ1cEsZKVwtNew1ENrSveg24bVmy5IatqaPB3+fWgu4R9rwCFdsxSVRcTAIiAoaBCvzKMvB3Zbw
RGoZS2Za6DBuUm1ejIADgTf4HG2HPgRdbnY4TVXejyNHL+M5q2yoEhMBBDJf+t9wMFJ2HZsH3KId
w2sL4FtYzZ40MCGSC6MTMNHCUeA5cweboD5PWgGiDz5vADByAULTEsAlKYzwB9URLxnl30ACQQVX
6JUstQAxwMd8GLuw3F0L1NNXK0GoWWmotqG3gS9VmxN8OMEgrp5CH8sQRSAmDL2VXSfdxFRYSkU6
xJOAbhNOxL2l+9/wazfJDdLL0RjvRrBHSzQ/CF17GJM3gKwYIWPf7wtMO5vOn3dm1beLK1gcfK3C
sJJmCTr5LCvX8+krmQvHEihOzJRmSG+BQS9gWq9p3SRio0mshluvIj4JKcMHd2rLvx7utIQCFhkY
SZDQTZpa01TJ3XD2d4nJX3AIxk2JA+e0SlEtxOp2nvx90vsLwvkj2j/q54AplKTSJzRqD0ayPLX2
5PMexWdn3lYa4VMtnVtceUTn09UqEU7leA6nln0+FUCyL5JLnLsXGhqydyzSQ3Iiz3uGshhHwwDo
U1lHn+CpIGoa8WbNh9VbHmp4bI5jiX29UJeIZ+LztG5CfSPOPKhb9m2Perdih3yfD48jHJl3FgK7
ZW84Op4hpHEjqB/GxNArNpVx1Dzsy1bJqpABb2AQzspybTv/LEyvmirGRFwqJePVkYfHgDTNgb6p
F+tIZrdNN5tcvihizq8ety6oZvJuRjztg471oY9gaU7moFSi0IK31UJ9rs/C05OBGmkYecA2/Igx
b6/ORkPscH35RmHkW2YrK5MvS8FByfbV9yp94PQqruqVRRJemkcp6QGkI03XL97qoYIB6xKIlB8A
RtPeS8kLbBQ+/VAPaERcqSrx2rhqXl2KaxU+LvESL2Lvoex+i5z1l76xC7KPW68JXQp43FA8fgYQ
VqISmPJgdV7aSoytsXcm45dsHExMqJdU4RPxsRMZTW/d3i/KAK4CsC7hDY5XpsTbHgQSCyYUszt2
r6vvGF/OSwM+2AfitM0ph+VFw1XaMG2yZC9lV43cfOkEmkNrFTbhnicYGvSKMwER+OkBIOl31ShD
m6a80ac5h2GyLmh4fCkcrB1pbgySyWcOgBSf10THQtTGt8LyU1H1imWN1JgTkBpDkagPO24lTKKg
B+juMs9XHzw0K7CfobP35UUdSQOs2WReT4JyMMYzo6ZGlQ+D1LGyoB8zcdRVN+pPdcaNOhb7JTXQ
a+HriWbcUKeVfuuJl+mndr6u+3eR8FiPu0QkU9+bJJ1aLUWsO4bXGkZ7DBznrDUQXzqoRdENpKep
lamA9jpVklbhcVu5r+RmoD0xxcDOzUaT2hgnz17w0Shh1jPy29f4u2XGdaoVhuon1HFpP6+p72tz
53mvnQIwhQlfJLlnkPtdRtot8EmMM6dRdcR5fQVoDOvSJeD4WG+Bz7Xe1G3Sc1uP7sAxb5GyYTmV
8pT8aOM2htVv6+yFEF9xVkDPaB2j1UhA6AVKVVYkWo/5o11mIiF32Uho3EppCNForR5CSklbfVK6
2Sj7msz+Y2La0/csUXXVxRV61W54Yq8ecm8aLP5Ac8CjcEc8J7iIoXbJ0FpjIJqvZrLOymilIK4j
gCl3OqHDBfAQxQBzDqwKMWLYub/Im4tuZ0ilH7kmxOViybgjnx4u/qyEKIbrr8xickZ1aVaE9vpZ
FyixEdCS4pT3e6AqEL5OAtwPwsyOzfZJQLO75vDPle8kzA6pIXWI2rds6qE/zw5J+AG4n5r/pJ96
weCfE+i273iLKdi1tn8yRksuhkqDhFp2P2/Hm9tFVi2jgf+ZHbNryxwNSSiYTxXuGzIQdR2Wrnnb
QwxvzwL+7MrsvrGSIuc+m4ir/eu2axqFoCMKeFY+Jvh239RKQibYdtRrGRWMgBYL7NcPA1ioFfK6
PysN/rVmvvOXcgBiobx1X774sKq+ZZ3IlB7kuhh1OdjQc+f/9hLBM3cY5Z2Dbw4U1i02aoV673MC
9o87uq92IeIUYOevpzg12KmDpwt8RR3lFL+UNBO5H2iuq225DccC+P55h6tDkW+2jVdeH9/6EaTy
EF7jRdrzdydXIR6/46bduBN6lTNva1pmrZ0Nf+xoWeJ7RXpC4DEF76NT3HKGaD/EZYvbytpyYcmE
RRDDYeTfyybtwmBJyJpIRRg+fTlInl7ez7qozoJZoCofDauyG8PEQCMSiR22IKJmCsYDwe3xk/YU
HmAtHLIVTiFWVQpktuUUAmnb58rtvm2Mz+D5TrpdSqJ6WR6oHKxxm3kPcs3uCrHqMAQSkuUlPlCq
rDqUwlynAtqoJe+SlD2BnGr7RrMGAdtg03bdFad5rjtBBPqk960rFCFvhN1ojCmevy0Z1f8bawl5
kF3UPDBgupeusc3cbPUEDIjfynSXW+pC8WUro2mpGpnf/xhE7qb4hIH3BBgDj1WuQwpFMk1wJZYe
YwVddcBB5wMsEObDjpbdOpKq0VzegPX7QYOXktUh3IT9rO4Bv0BaIhbf6mZLLotmID3Og08aZaOe
AKWu9PrOV2vh9+ZFsvn88y7u02hklZXugtGoLQcVD4PNaOxDo5JIqApGGKyiKmQ68I0rSsw5d3lK
1wdkX7//3mz/5Ct8vug+FqyV1hXrMJcvOvduXmRoGlQ5HA8V2JZf22ScB24ddnHeZJxlg4i33Oj6
H8wIyOItEXLeMnv3riiJ8c8p0dHNUdsQ3+XXmOYsUcxA9nQYYdoPP6sVQUU5osFmnqVBPX8t3FPp
t+5SHbSetsqfFxfVG+vmKFn8+uyUx3P5CO0YL2lJTvjqFAaGm4DRYFaLeJ0YwdlTIEUYH+BAVdZs
3Hv3wAfWQSLm7MmKYWXkp2o3OnK6p6sfLVm4px4ipC57/tJFWCMiq3r+Br9cHFxaprl1LeTkos5n
YdC0tcoM6AZ991bOA5zlveIoEC5zwoV6LbByBpTg4NnznTPLvfJyl7H5lgRQF+kyK7bgu/LhYx/k
lHLyjvlHIuKh9BTNEvP6w/cMS/BINMY/8r3OD3FaULjWU+fHTjzXb+Tv44MHn149yspEIYGz2/ZV
/VsFsqBoc3OnVdjEuxJ/s9u5qs7sRwZEnSBkB1m6zcz0hqeUubog2Fp5Og5v2c/Sy51c7ePDXDKI
Q47YzOiFx0kjk9w3ytdZtkjB2zYNuu+kiNlUyuOYXxrD7CbhTkWFxkmf7Dtt+k1WYupIXOXdvfzs
bVUVk19Dhz7n2rzhEIsFYgzGLClU/z3qt3DU2hspaM9QvZcX7YrwQ6CtbJtwR3+YdMN3LGV2pz5K
yS9t6YJqLrbOb6/bE9ZyNQHQNf2hy6jtKiPV5+qIOR9wFwwWVQtJcN6rwt8C7kvYZRbESt9s7JwR
YTHUq1gCK3Sgcr4lSbAR6S5p0JXmlWgRYH9uQfWL8+grNBx4jXR6KlQtQeKO3JA1xvcU0l8LVWeS
9FtSpz40JHsjGziNz9yWOBd+OO8BwjG2gm65AZOmfDJIAepZajQU38DVJoWV+3ottxPmsCBRtfYc
y6P3+a4V3FSaDgbBTklmU/gQvAzKYRnQXWLnWvmHWBUAieHTmZ7fqhrszEtHf4kkCef5j2JAwcgp
SaVO73wYVNziJju4PDLVZyWwdVMiGCZWlVo/N9Fv6nkdi+bjTd9J4Q/g5ih412DADxSo4hou0yHn
hYKgQ+qC8BaMEMi/j90dRkYZSBF1Ck92mNy6jLLQhILMAhL3jn7wcbvQwzqGNwmPXrogBvgc7MIq
zHYrBaD7V9M7A+Q4PgLIKDkoGBgRTmaW0N4uA2GvjNQMiFSSxVneC6OAtJnmVUgvn/SmgROkf15/
RSbZMhVd+1PMQEx5rEx3CoQCAtO5NbHTO4w9w5PqECX+sfMD/HMYkzImqNqfZshciJvsUyRWclbk
icyiIujvQRV4JSVmNW4xryYsQZwIzUwCu78MYl3DGucXU3Hm0RqOixw8s+HUOcYeN0h+iLjUXdns
S9JlcleqTiqHewEQcaN9m7FV0CIAct92VtXamtXxIiNkcd58pEoGMsmKKtsTEnjba37qDoX6ofwS
EGmcjZ9McUO7WVUHt9vCg0pIqC7G4cNGehsZEGf5+ZCTOkxq2K7mpPmrUp4AkJzcwh0Q23gTTVeA
b/PAY+y2slbY2un9ywVFeIvuQ3z5atpCQVl0zMad2vJIQXA4wVSFdQoKnuTZDZbc6QQzs/2nEO9V
tC2R6Rq8A068selz421W3qOgNCem5+vLP+lzNvDV8SRzzzCZENbemmL85Ez7SOq4wi+rNiwH1sog
Yvo5cAaXRiYOrAm9gc53K//z5jtJpLEc/4SeIdqZkPid8PpdDj0dkVYFmnHsMaQE/Bj8UoGV4Uu5
42SfXmGwmKCQypO1fYPYLdvWHS6bQLriSGlSPAGvnWtGdTPAo/o17XF68J0M6aPJc8h/w7gs18Ob
lOnhSEUnuCDHox4+mU7+prMEYZ8OpxAKCo2l/QqSBfrTI51+Umo42WYCyShWpAOzSfu9fvO3E4R6
/EsObKeVgApzDp7SGTE81YfHgowZ60BfymLEAC9UI3VKk6cKFDp6UFHTJOW89EFkMHISdsdw6cae
h8Ja7oozcvc6w7WgLQANBof+zWO9IFZSRN67OwmNzfuGdYV72qalJNe9xbiCp+ce+1DScVrCkTkH
IqyNh+8aisZapoyHbISfOQzfV/TpU2W45rFyLJK6aHUbEAchFxIqrL/FdF8aCbr5Z1fLjA2/9sQ6
aApcvhBGD1OLnITGZ/UzSihZ84ASUl1A0d7KN006bwB0NU+WMokLLzRoZZERJhJS4bQE5EF6EJBg
LNxR7EjfPnhiBqeOklra3K1FmEHx+/6kuxT7ncINITx7ujdTEb1kzaIF9bl+5/k+U9fWdnoz8CXP
2ooTeHWLB5Yui+ARL/Eql/Tg97fQsVwPNOoCoDWn8+PY3RcmK4zStW+5FZfuCQjv/qJhBHEn5nMA
hYrWHpYvg3jZOSfjeDJTbtRc0zdIojz2p3ACg6jTUbSVcX73VUejp31FEztsEGAEZCqICyiBeaWS
DIsizrl6qjvPfcb8v0FaKRRtC0wITDriD/BnHeGZ7tDaEs49Z9JQTWR4TUjKGkSRGCgtnkYwOz8N
8Ksvqptlick2y2Y/OJHVrTvvk2k3b978H0ZM02xdXZMxvrJA2jzv78X20UOJnrxOnpl+g7fWNEhR
olxLsPqf8/OKdmpybeGl7yv8rsBEaYpmxtR0mpjcL/JMR4iox+62yZC+o6koU378l0HeQgfD2ujG
JxlBd09uLU8/AJNxRrPp/bPgPPro2BayrdD0riBgHSEdvt7qA68ZSIXMmReRvuUdM9l1TBBrP4Kq
UUBwc7ctYXdcYA/yLAfArdHS2gc1r5drvOQ9UpL0b9WLqR9m7pt4uP2zWenY+YSYfm8/POX03eDd
04L8IgrBqgO34voFNCm/dE+MqsCAbPl4d6i30/rTzxZSjlVjPjgWtXzoC5Pb89opzrTDuCy11lRk
w5QG2gHoSCo67pnBc4RUBKog6vy0ooKj3ukXgoUbsTamrqy45j49SV0ZOl2IMj7T2Gk6bQTlTvM8
X1awzeH4jmc9QQEFr3yobX5nutQXtVsmw/oJWH2L7SSDwYvBhrUGMwswyaJ5sfLRLYLnUvCYY8hb
nnf/EbtfsyNJZ3MZ35EFGiZ/mNyROIv6tc8TQyPgmSzCnXGcKpHJ5+nuCZURbiAVjXMcoOQONLqt
hfk+8jEl2uR9clCQ5bPxvTku1WtZuCYQvLrHF4RPvSdFsNueFQnKmYaNKtvpeBzAuV1DWTtFjWJ/
IJpNkK+FfrEg12hZ5+4FIBez/EGhgVW3wftaoYAXdswMp0KSLcEyWgZemqP7MLUHukD9E5Xn9Tqt
TEDSoTfyXTHeuagfrXnfcCS1iip3+IErAxKXKXYeeJi7i4ZJC+b/qX1s/BDe0uo9zQpQ0DxdI/F/
JUjdaMCZRZIwp/SJm7K8oPGVDR0HttyWeHBzVWPLLPzN11MSzv4UkwGklACSlGCuIfgIh97J3DOQ
gZO1uPVaWNKttvqwY8ojSHmKlvEuzWwvTmgZkChf9Px7Q95pBIeovSa6Fk+eDJoswY0KvJ5gnjzA
+kIoS4YtBc41y9JTatmetppSjeGvuK/XuvgJUJZSYKr124axSp0U2XBzE8sZItRirOgQ0EiKWElx
f2103qqi3jdasm8EktDH4GV7uVTIPFj8fE5rsVUrGOZlRmpyKEXQrQyhhFKm4jLSaIF4XdJD+sie
VZvTw2g+YjMEfw9MHtVKnvfl3kqDOibU0BWu4tS/DWDL1iqqWDBu5UbmrMmIZHL+R2ZJOa6oeE+V
KsO5BwV6BR6F8mTqndnGWTK9d5UalRQJihqENWkw7iyZLpi57bX3a3usrrAvKwUYNQ/CTXlg6mGa
mOILfFhnITOyfWzEcaYPSKJ3HSh6xhL3BGmJOhfSKrfstaAMnvoicnVaw4fmLmx9NVRpW4aJnVOB
JZlVLWHTmPDbDxE5wohYakEuAkw+s5vuD7p4uDd31yV0x/90idoxgZoG1vEfDu6723B0P1oMrHft
CnqAOTRcdZKKUIP/IMfhEwXQWadi9s8zgfd/Yy2mSNoVnX4WTIYxdZ6BqWAc6wwhYctcszYCTKFP
ApArBvCiRQTyAICyFJSAmbBNKJv+xT8nxhoK0v8dX5dvpld/KNxlh+qQdAMUqyZV4ovHyGSCtnSq
n2gBAhtuf5KSIKAeyAxdT6ZFMP9Xa5I6nQTsXuEpxIZpf5QWtbNQKkawhM2GtDav5fyhAW3COC8b
aOWnd2DH1J21ojC5eVaCW1pQdS/6UIDJqvpR+5t0DKwM6ZA+gbx9up2ne9er1lmc2uyXr9haoNFd
BQlTqA8dZ6b0sGF36FaCEB99jazPezZkDJZ0DI2pH+Lkm3qRlz0ou/dl1Pk7UceExOifzjEZEPIR
rBOLHeIiv26Rh7QRSzZzbZhQBnibl+lhzm3tiqhjJFuE1dnV5oGAbogU2+ybQjsqfFIFTKUh9rRj
wuI6/2P+Bg8g7bSOxq+uPdDi4FNzw9idgRZMinziua7nTJVwlrZWQ7MqVuh+PrJD44DDh4lTHj5A
Ogu1NlKVoTel8oYP2B78eAcSfqljDYCz/0IMT+NnEAodYuGrXR/Tg8nvQKk1zevT/FBIUWZD0/GH
I2T4Ya4pkEAgbyhjt//MrJOcdtpfJVIBBeh+YH3sh1HcahuAHrS3q9SqpCvnlOrrpnAcb2B82uR1
ieX6QX2t4BSX3v/VKBgpxB+gDC61VkzctmG5UvxQpWh6b4/p0NbytQfoYBIwJXrDa/kwb4uGA5cP
l9/KpwADMyWOAd+0eGJotHpKvhvv2Z0BiUrVUH6fcPoT00g2ksK6D8iI63dqakYJfxrAH0r8desf
mpoVLIItnqYdx7Lk40/UfMz2QpGpq9vngYsEbI3SSZCpO+eUuDoz/1JmBTJQiyuJQChU9CWcyb/M
sgwQkr12tjrZvtwMO2Q271REUbVFCGxUAw3sZVRmYo3DsExzqzkhqShpQTmUsEqQxn1NqYDzE3cc
KTfcBWgmshx69IlGHuviooWhP+pWGYrsy/ekohUrY9Q3uDvCqB48+tocdFt8/FwtYtHP7GdPU1Qn
FsvRZrd+OigyWFZxxuh1xSOQ1lvp5I/Vj9PED7r7CrF9xaGzVZnJLCajj7NCD7os9PTJKfUyy3/i
4ehep9v1goRtTvvVp1tfebA6F0ybVSK8xZt7yCoA4Si6m1yft6JOpQKmvR4aGYm9enoYOaBX6yhP
TJKKi6u0tlY6BAKMnEQRouAx3Mv8mY8gPa/1kkgmbgdO8MEYBAI1fgdpqd0uPMNDH1GN7EgN675B
E4fL5O+/NSTStSOn3SKy837behGMU4zkmdVtVZZ1mt9Jjrk9GGFMJTQwHzF4z/xmSU9hhmQ18iJ0
lINu4E8by7I9pjQi0VF3+xb9EPcwJH+nRjLTxv7A+YgIdCaYnWfy+qPCzPihl9Bzu/3blHwyt3oY
u0EwkXVBBTgb4sE7pBwqXds+ODXu+xJUgDdjKXABNBfZPk4udJN0SsqBkJje80AcaAVHaVQTaz7a
0Izt4yMig8XtQ+Nkgu4+fpVwG1UTdWLhhHFtwRdrdjS79Iif9ZmutJh29vtQ37WEI8OO0xQnV3aa
L5C8jelXgOAESzmwlqvrLyJD6jYHFdCD5Oo3WDfVMf6rnzHHHSzV075PYQcE1YD25vSnjcOtifzl
HhhV7BJ64IE01Jc5d0r5TZsliuE23mK0QP+5cP9kQPdrB7foxqvDIgdYv9RYjjCEkhXKny1wQWpz
tP/zSnCczZovzaVeaoWe8+WDxPAIaQMHBCi9cVZ41bBEdr968N0OpWUnZDNRjpho3qh72Oqejqvx
q8MoIe3agoDi71+IJ0u0ATjAdGjM4z+IjEUWf2CtbbaE0HIx2JCu8s2GFxMK0JnPIDj8QmqRj8Fk
Ojsqy3AKORqYH0tNz5aoAMtNyPd5u0VjD3jmAcUfM51tPY+X5D4d5Be+8w6ei37kPbGYVRtBPQtD
Uz3BcXLKHL0mlOU8xnuQXG1KiJjFv97inHJAXG8xE9pc1Dvyb7+TXEQQav0lHikSyK1U8ROU3csa
03mC55AdMseKtGjGaQDlNPVxSqDi7v/7w7GjWEwdLdFZ+i2xvR2sbr8uWyhwPGdGDPQteLirLbl7
S/u/HdDUwR/DSb26p1BpBbEmDtG55QVN2NWqvnTbc+TUZcwg45cYULjqjdOsx7p+csNMsDvBaxRN
7AS8trWq4sHf3XD/ey7YFUUQAb8dRNUVRdH1m0Olcv52qgiz/QgKGuame7AtIyPq588W/Znea9UB
WQdGxAORtLrHocroazYCDlGRj9VebaGF5b5h1JGh5pwy+hLSrivESg7zH3oikoGd1bfrw8K3Kl59
islwHYQ8nCGhZKbeIRj6P0i3SH0Qbv20U5wtHbY9sgP/V6WxbnLk7KFGSqXzbtLnE92JAKB8ane7
qPyaM0p8f6AurkevqmDja3heIo9cGP6hKBTAHoJT5gMm9+HCt2ZvaFIAg4rkfllTv+DsbXEiEgTE
RE9YUgT8cc0VryqnMEhpFHZ9zCjZHK2jabijccyfs6oBtCIEwzrCjX3CNFQYfnk22uilGNUSCmZU
3/8RmVGLD3Ma5UNDUG3T89+JOjmINycFyBmj605MILsYwWokBaElccWi728PYxMfCC7ISGJPnKLI
ob8Ev2VBGUIjOWG7WPe7YUqrsdlb9+RoAqDXKFxO+Fgs+3tXRmol3q2+kEGQJ/ovU3S9Kd0knFET
emRiuKft9etHmZJ3lx/JVDtGm4iGodQ4NeJfwDZQ00pke29lX7IUapJc3oWDXMRggjeVzb041jh6
6Uu6tHbvFj75oJWqxwklARnwczaj2ZIlbmMGeB9PK9s/yl9uf4cV6dEClxjRWbQTNucgG0bi9FfJ
ZKJGSPkT8GYReifu6HRfFB+KSCiLnS028DD2fNaE6cverP69ku9rY56uuLSgrTAz3Ue2J88gnr3p
o1V2NNagl3sf2ex6DIz6qTM1t8ZfaNzVfVUqpY4QjzMiihKGe1/pDxkzsEYTfNzDXo65fW4ZgtFM
QDV+oXOsNcg/QlKRSjKsohbjj1H0rxFk1elfjXaYAam1zo41LBDpvcaUKrVBDWsCpqq5fc3yVH2w
HfFVtJby3JSj4FCCRLNEzWVEiMue1IQkjWnvgtDjs7Duw5NGfsErXY3MI19bC6V6tqr/LyMcrKS6
yRhyjohKugqp+74uQ4k4ubazY594yGzZzRJxQEjy83dGx5uUY3wQSr8QGYqQivap4EedsdBls2/o
y3k/O4916LLUwLcMmPjyPfugW1waTmxa7MBw+KSF/Y/c5g/btTAGPAjDo/xV36ojGhjh3wHQqQha
qOg0uslj40j7b4xu5Q5HXkguAkM1cf6A/vNyL8Jc2mORqgCnffk5np5iGW2nXPlMkokbu6BJ/DOw
BlOw9uCUXZMa0Db9T6AUZCPzKaKm7hiQfX1oZzu1DsGzxFVdu1tgw4xJdXkFK1qL/S27mBkBvs17
TkZbT4rY1XiJxsqQFMmHf1YRBhS7TZWR37wuGQe0DCe8/yXFOfp9+kZ/MKQMEEZgpCH86HqU6fS5
cZgjypsYnPABRxLG92RMkVZMXOwqJHpOMHoYk3iHVj38tC155tdOUKvWFWIs5bnbRz1lrx/PAJcC
yd/ur8YL2+aBL4jkQjic2RrYnShcGgRiJZvkTU5bW5EYEpaHG9AQCByO5I9aNS53PQhky4okuQ/1
vb+cQlBK7VrUoDyoc0E6LYM36t/d396TDy98pO8P1ib8QkY3XiUar5a/NTe0EbJI97M3CVJv9Qxi
AUsap/A7w/EtRZSSPD4KyMuSBJBlRy8XEonBk6Ij4EVvSN4S+9b8upW0LYvRl7z27u6ybcckfMIK
uMA1qeBsT7srI5/BHlUAtYaj+yoqSpWyAgPFodCuZbVOulVkRDyiFqkUO9/MQ+nGAeY8MXuttBsM
wtRi4ReWMsB45kZqE/bkbo/AkVBSwmSiSD/pIr+BfC2uzA4Iz/4ELj22V2nkF3CH2/vpztMMsHMc
jvwq+E6U3JaSr6g1fbnk5SQSZ43t/GSRlc6UYcmTq8OYZMzKQLOxzZPeqIXyZszhpiQJdfJzxH4u
tFMKaF8+MB79MWrrEloveVprzR2VDs306y5uk9iMViceL9BCrdGflxnu5I390dpcD57D+/7TEKRg
BuFitRl4mKT7dg6ojUEFYnh4/UgIeigJZ6N78FBHVIWg0HjoJSUtZ7RCppYl2NzkGqiRNS8c07rd
DidtGzLSSK2eCnrcS8WSJ7AMqD8Ot8Fj6wgvExtoUgvb/g1zItTn92h2xTxzc7Zi6lTpcc4VD4cI
sROGlFSlWA6TM0GhI0Ub5f3TpVTPUW5Vccwaaaby3dELbLig/exihaCbh4wihJlPc+T6sZAbyAGs
Qhe09DJwrWz4levdfUQkMBRieHYxzMaTDX9DwsppXOLXDPLBRzugi2yHZUfFCeSxNY8CYzmy7Q6D
MlUYgZFo4oJ+IW/6UY3+vCzK8iLAlH48nBidXox5zpKj+X72DFseK8IRrdGksBMcigpZ+hHFagLS
UxTTDdtyQbCvP8d2TMot770XcEthOJJCt8BGeA24BSZ+CsaHQMzRMpTx1Kd2YHq/cR/EaXz9gSNu
dL4GQs+RcllfXeTmSNkTBtbcnz89FukTNljSzX93rpIhixwyoUVmmaatYbsEp0QWYySYzAm5cji1
jIc3/Vp+hzgC8UnAXGmA4s4zRYIe0tlHuBhTe8kR/jP+tqE4ymonWwjyuZIjBGxkvGN22gXKm/YE
28QYWtCpARESpW26YTbJtoeEsqbt3FBQ7sCF9evYFtar3KjJD6iSzY0S5DFbNmbtw7QhRq33ViC5
RNUhTv60Cwj4tPn7yqgyvLD6GnLKPuV5WSwNXoTqB1E8y9+GsgfYdOIo2l2pGSiU3s5oRepEbdb2
cq1XGgFZxeN0v81SYS0cRq2e+o/32mdoqTuzmHj2JVLltAgyCQwn9YEIHFGdWqlojFe50lZ1janz
lO/hBT4PWzOR2OdiKV+u4WHttgc7JhckHcJzfngG5vY/HnEpMxp8E29KY8kGkcs997O3vosQK90w
UWPx6POVMtvFb6AOPbYYZ+0RDFy10w6EP/rPw55LArdQG7aShzJ6CNpn+lQ2s/vSaKCMGqr5KCRB
T3p0RqLAemPc70t6yauawqE9oGTH/fb5v/R2auKqK0NFXJzBT+/JkcA1MxFg/eh+B55GFL8l+O//
sZarHGgy4ggLLfy/MJegCo0EjeAz0Q9A6Opb71zJzSTRli90ycDhjv/xppCCMFT69iimPN2nLhUV
Uarvi3J3Y/uhz/1RN+8cfiDU/eX8UP/Ml99r9OYvqXrnc4upUl55kJhTepyKr1QJYb40PtDwkr8u
IerIBPtVh5f7TUCBoJN6LIvVMOUXgVMc48m1X0bdlLZNmXM69Q212pq9VRqFbemXSkRPjrbLgwWo
PvYOHFXtWiY6DytImglYyrTpVny0q5iD/RUsUMaU09VUo9Pkd4WgNFat9S6jTy7/1rc7VtefRiiy
fJ+Fc7YYfARYo1xgUfSTzBHDvEm7fNZXvQG46Xm7AWgUIOtBDrT3jhhczWzRtKygSDIcV1Sx9Fl2
s8rJbIK10SEI030TMM60WIxmsV1Wm8hkW9Gcl6WZeK2eUqFDptBWkvvN6HrNHfjkTFvGOfeEE+ib
uq4zG15NPgZrsHszjv3Olu9RwIRKwXx9AMETtieeJiCYFnn7nUqQRuzz0fD83H9zibk4Spa5OZ01
BY5q8almZWlwRSqWpYLf1nlS2x8kvLUk9ojUvdsdqappD9txpeOpFF8041GniGosAqa7IAWLalMM
cwuerh1nKiZVRgpb7NWsoXimro6bCyE7JM/OlVopT0uqCTpFgN+VIitFl0RyxcHHaOhyzzjdE/KR
amm2XNrLD4Gdo7eZnUgV+97ePoXr5gpg3lwLoagUlKnqEZxHEIzZC9FKeEK9aIwY7ROtr6z/R7EN
ZAyJtmo8naXwq8oJK0Fau/VVQpqe4c5f+SQOIdspjclWjodh0Xq/RXlEM4Rweg9tOMhZ6wnDMoe8
FB9CJfHSNidXRveO0dD1OegnwX+llSWz7a54tZdTSjo94Ku4ue17AlPtKdeSpiS8Dqf0TkYVJJCK
WCDdZhVQnxPqk7cfuQtfDWFZT8tbvjjsICwZ1eLGEK2WSbJ0gV6XKjEH1dopqPhfd1LJktx2a+iv
s/RJN9iAJk4o5eHxA2sEYuxX4oSYh4Ul9MHuPFN7Vix44MzepeEStDDUYupn3Ggupq9dmDOa5n4P
ZgmMuJ5cYOzDEAwE9yuB/iczY74sOp9ax73Pq50YsemWuGbyKUszRUCjpEKYZ1YP9+l1e9ozLUH2
hKqBxGDiwSKd5JZdlVMq42P+iQaBL1cmmFz5vw+1DhzRmNrs+dfxRMp+7gt/OZDKYtFMTCEUDYWS
QCjn5wjNbSUdr7V6ld/csg9OwTEHYo4d+tj+TpL0xKYm8KFfXtH7fvK/b+dFTf8bfhhbDqEk0Z2+
Tr73RPsE4xHvKQrJvdMyzMgE5vKU50FOHImOrtQnYSv7nWxuKZl1T/28uChEk5Fejpw6LJRtJ1I5
Wp9rq8wBvrKnWv4sZjrPW8GJUjwN/2RkzhiAknq59Z8atG3OfwYOqmef5UhYe306ks65aFgUdwgk
qD3z8vwUHDXUtpXI/vXh8i7QGjy7Vu7zXdsBzPz77cpuQy+WZmiXKl7YMCjR0bfRX5LEU8E6KPhm
vHkTFoX3n8R6cyMpLS/58zjZKda5GLYtd/aX0opOM9j6Q6l+8jhcHyRWSm3gjHmLSfwFxs3xTv4D
xwN3eUPaikbNaJjgWIHaar3FKBwC/Edu6fqubJiOUyVcCQxfFc3Ekuwb8G7t8DV6t8m8WDEsmT/a
rMZ4Lfwr+oP0yAEsZDuxg9oUdweiYixvPivwZXlBt78DeLQkgcmq2i9b/rl45Hjh4xwsyT/CITzh
x9riy4wu9nKn0VCoatWF98fu/qBDxAe713oIYyBoPeVRq9bTEuHOnjn1FaJhoCvsEXMnlCP7IQuz
Onxqk8Z3FqL4noKWZ6ah6tU2Tc1dWnf03mocsFR3TPH71g6KBhaEqkptqonvENBq2KXV8g9LBxRt
waylaWeEJlmL7uLIUb7VjYqX+8h8CnI4eKJVnGcUdBrsWCRRZhiUAAQkhbxLQIDOVrVZ10Kiv2VU
TAm6ZQeMXElGDRbtyvZCqZG50p47xmD6NW1V8F3NEXZcSHfVFxk9c3nI/8nvlp/ti+n1vlaIkGzk
YbQr6ReNxOScUE+hXf64nUEP5mZP5F8UyyfguT8/4rk/gNWKlN09obr/lsX2GFPS2bAjUs7hfVrW
LLvUvvxcmw0Oorg9GHyn6QErgCU7ytHlaL7Lfy/EGaQ9l7+lv7RDzYI/G8GQGM5BylwVRjHXP0aG
0DiQhuN34uX8AVq8NQ3zxy5sMCYZjC0iuY+/A7bPeahU7VENnopB278MIx1/BvaQR7u7v0j8kqeY
NbBUwf6MWW1TtAWFeIvDkr7aC9A/vpOCvbufq1thc35zNolXd6A9kbdS02MUh0Gq3VRvK3O7CKV1
QkX7ajCW+Y9oUPrqLHo3vV2Y9zsNcRqh5tnqfinoa+mw9/5+UhKk0dPzUgDNVoYD/g1FUPr0fC55
FceyHHaZ/5RryssV5J4wViA/0OhMoTcp3+c/Z22wvzCUorYyQTyT6R0pw5Qoct3I+/lcDLTmVGny
6XDMy65uDmhp4XLeOgnm84sHTAjsFeHxztwGLTDXjO38Jeayin/1IQTGhT3ztPjqccgvDOy9SQ/L
UopEvCR4dV2H00v/KVBSgO+ererc5osUVBmRvnYb+fAImKiOO5dJt4gul4W0m5B704UHJA5rViBy
KKpPRFKzUo5cZNRm1SOfNrI+sN8fKJhY+N5DP0zCniG/D2tutnpjaoQP7ysJwdIJy23hRiF4J/12
5njUMo4vQK39DV57X9yd9piLcNpMweiXoiC6K1aRkKXGApzddD8hRkjXGHoHVmSCJZuri8hZhlqG
4Q0sqg4C2t0RUpIkTpgxPIkWYQYi43H1qDbloqAM5eIhHU/m1viiiak+tdH+c4Njaa3RsQnAUQQ3
7uocwcKTH7ehvJMENIooYSIjWK6CGXtfol9XI9BWJu2giZDHmoJl0mLhQ+fnlk4H2InPcr28BToA
PNzjVNmAVPCAshlheWAZaJ1/dzXlU0/aqPiGjKolaa96a+P1hkdATVyRBRjbj40feEHT4lSP4ghS
qd6b/f+TT7/F10gE+l7i3k0NH1hFAnFqTW4BaoY+YCDG/5/xkuYdHq5kA3rwyZFlv7z+OnAPYsbD
xQLG+dknf3GmOnf2ZVetXbrZ/r9eyl2QiGsxTHGbWdFOp5kdMszbF/oa3bAo4OcvvByy2eHVxO1C
KwF/UdUPge91dSCe5mSfogGm3u+kL/OVvylQ5h31yU1cZ8zPDQQBVlzLRhAsrIgNafue/xWXfZbM
wZtuXfCziugeVToShIHssrn+nghl0/8w8dRGjYYtdjEMW8F90qjScVUUQOovIE/s/3lFfhGGyn7H
KZ9h9XY6+n5d4JukFzVwZ304S+yGkYjn+4IzHNdFl2Qn8xFcjxd4zuQ/zSwqnFNU0p0b9I6MsvVK
D0hGwlgSIvAKkzd6ZJEzHMjsAS04/jEEq9aC8tmcxCns4DEX2RlDhIPgBLUmsSxQ+jYLDkX2c5g9
36vA9+FQysi2rEWTKCtBis9Fl1ENKhRzn1ApfqtwTZxNdsqZTciMp0S1PHkmMAi6ipiX1KkAVHX/
jM269Z7oYeUQTu199DNVYHtLfELZPZS6ksRoxh8Mj8PCAcxyAQE80E96r3MwZFviQeyWpSlsJu60
dFMbJY/3rAi/1eMMGpco8vc1WiTZp6kDeknSlS5+wMdS0xy2hUb7soXE5CfcH4JfAQrYO23JWZac
mkszCAlTlLWaqD8XJQ+BpZaoJGUT47kvDPUkNKs9WMa7ImgGTI6+KRsuCTLK1qHyMgrb+/iEUNRL
qTKeZgYPL6kM8DUDNsS7Cyljm4qvJFwoqiIt4oVNTG+0W7tD7TsqU2JUZObu1zkGvJX27/uLl8uK
TFkvY2p+ykxG1Sz4NPyLeUu0h6vzNO13P3Hx3jrQ915m5TC7U+IwzDRVAIQwyvq9gQr2BvOfw/NP
JF44VvA5ri8hLREsye9o8jw2AHYHXMYPFBNqvXBI1N5h3pUsdebAjm/h4z6FAb0LkZtlMauAqHMs
+NZspMErWQYqGfhP/t9R9lMCPHBt2zd7m1GSfqiHGFbisFwKgH/FIl1YzLOzZa69HJ7GpWgEOkL+
yBIzFB221bpAo+er7juudiBgODs6V4eeKsiHkbxStfVbm9uIGnhfxetAQHk7mcQV8rSbgwyBjibI
SVW5cCwXFiguvUVvxzklmIxMIgwi5zhKoI0engkfUhxnRTXNPca1v+GlwYztp9kUhKLJurRRYDNt
1eEl5j+sadxCGCpktQdTMq3VMRazzo1wZEVv8lXDoJyYwBqKY9WQU0UUOXP6eKWuZIzZ0yNE4tSF
kQEHCc1BBg51VZZ20V1H+XDgS+gSdRwTbvZjqwXvwue/iiX/p8m/WHiRV/8gygjVgnHvYkXQQICl
KOsnJU9nxicUD1Ot+lg0uWBSZRLzfI+dzdRC+V/Z7VR+AINCgQzMG8uWRdjycHBdDwxxp7gQkd8U
4kEUwHqxYbIeetURjAbZXx1CwHeFdCgCTtB4GPqT9Xnvq69U+MyhUapgzX9IZpmbIIt6t9c4Bc3V
mL5YZnreaE5ksOJvwJJ/ENHs6HT0ZUX3o7InM/rOg10oh+C3I/RrIc8/PseUiGV8akkgB37mWf8O
pEYQilawHKCAZNBlaCdF7KrQ7sYSUWvduS0X3bnQwVE5Vgv/MvbTUM8jUAlRuLcefGVMmeiwAQbu
W0WJb+6cbEpeQmrtNogor2DZADtibJS8Nf5e3SAdubhjfuapfprWbguPMiszuTeBqHQrXV1D4ZPe
lDWOmNxoB8veJJhaKRm+Xp/zvcVK6IsyhBFPsMr6beL5ZE902KdO6I0zHRcdIWAphbWsbijPYqfT
qUQZ2woSJNzjKLBxsTriacVV6uAeNs9h/DB2Xsj/OKc/pomi1OFD7P+WGykgmZ4EHkRQn0LEKtJk
TALTZkJMUcO+dRM/cffwlrIqBSUC/O5Bl9qK6fClgZf584Cfk5Uc23p093NQ0pAZPciclgC3YSm+
Pl2oQjAOJPpE27BYTrDhpgo6bCxScMuiAJrKW3t3QEyeOfSjiyJ7FuklyxuZmKO2vOwQEvgnnCmf
OTVpD6m6oXRQ4+WLJ8ZQ2ZStlEcQwHvBj1MP62eD7/z1zvjUySeJ9btVBLNB2Ylvy1F2VBwFYfBC
jATLhbWctrdlEWeydWTUXz2cJCZXxWFMDVAmUnD4j78uEZQgAi5Sk6HbWdtkrDJC8etxPN4qOtVn
QYfzdqfvnZu9DWJPUD/ebRrWsOGMRLB3XUzFF6GXCKHVLCQYY6Y9Em2aX9PnoMpfV8sj4tSc5piB
vy4gEUEyepJNzdIjXpa1L7wXxWlHRVezFAAlyHmpyGHpQWz+6pNw7Y1whE13wazK5tgPIKQFMFuc
MDFVRxDqG/5L+NNWtfpIGUs5S15KRmdJmo2Ck6PtPKl9dKBM8mCcfjJfePE4Yzl/JmjpRD5CHg1s
o7O561w//S00qu9wxx5jm6RmXdzxpD33lvKcPh2Sf6Y+Cq7yrRMjf6SGXdzbbaTUkzZ7KGFLuzNT
nMaY72x/GlgWuFxNWlrBQz6IWRuity/sSBTtMo0MZmc/XOAuUnK6bSns0iFzFw7dFxCq8PzPk6hX
BsJV+Ze/qbkahPeMw5AINhmOPV5xR7+QGmHijwEow1vz7YYnXOwedky0YcLG1EcZllx/YJj4FIQL
MY6p274OjUUERsVpdUwLgCzJTFRpeNlKDcdGb/LqoKRViEhSQU9YmuGv3SIBi7TCrPLTxlgjaY+u
GvHccXK9lDkKvLfGNwOE0LcWDCooTm5BWQ72vrPf1nSF2c+gyZ9d7621/80ThuLCDSMUl/RW67yv
smNh+veFsANrzOhEc6JbP/tnWfA+ntL6DRKW4PBPmzeWG0dOi3i3lBdxVVv0E7GzVxFVTqxmuEjp
mQK17LIuz4MJTYUBbqNFmrlVjqXcJke8TcF5a54TbaOzmijXpOj1/i8A2KWIwUHg9loTefhX8My9
P/XGeXyIlijSaccPT91VgE5KT1g6uRwvNwOx0dwG4J3qh5rpbSdtCovzvVbfUUBD6N2pUa/lu3RL
j6HH28WK78WiNtV8LiBmi4nUn+iWJXEMNkgqSLyXydjMXXzfwawrI0Y8oFknMMUp7CFFo5tNa6V0
NffT6rQ28Z6M4mCHZiR4FAkXU9HNuN3laNemEYRuTKGaKBgjfvkj5FEa46P4KxennoI5eB0vhsmh
qnUK6prwOHjWyrSpUkiO6OyUalc6noEkHmMVxGlTZtiauDxH0/21xgUZRA8qJo6WWsTKsoBISnWg
EVHbIpkKjwf+ONoOiS410Du3EMFc3ncXsv9mbjd7YKZ9+mm77M1pHa/hp5okfCyNdoGaEQgVcIaP
xgB5WbJhCsY4igKTqXGcKzHQTUVGox5IIpdTKqMe2GtWyDh29FVa4Rb+jQCeQi0Fi/F2XMwVPf2t
bP5WsNR58FMSzfo5Fy7X738TXlO6amlorTCxIQffWvD7fmLxfo7yFumhmAgh7L+lgJUXgUKQVQZZ
nlrPX80BYUhabHQOf0jQCp+V7OaeTcDXXA6R0l4egruOzJeGd6qMa78cTE7AKMp6/9Q7Fd4SoZoI
CUIeYM/pAJiMstuzORsoHpNka2YkgWzRzeine+AzXSrXdrTAYIq3RfstKqaS149fULCbL8awD+DE
m8YGlJ6Jb6kw2nOkaz6AXyDgDfskEVJBEiDqMcB6YCo6UNZmbVJZPKyLLfW/mu/RhBxM2hET8wB9
6sqLI71ks0zbIXxnKKTQKMF9UgR4o71A/b2PuPP0T/pw2uBkGby/uD0lUTxD6VNPXnPs2BnO6i0d
AAQttH9eSGn22H11fe0JxfiZPMDIrwqMg69pRVwHmhG14QeLFlLOxME53KoElSoAhLA7zehnQtvY
vtZ/0yL7s68+IS0OaRhKLxWZYVAYe6iqov7B9xPcu8CNtjrgGb8XdoSe/TPFAlLUW3RDbdZjhbm5
OAwoosk1XLvv16jCDPmkUjPEv0nOQfIvfs1Ymg3neoMdDwyg9sYkHrADh8QKB7iinbduuYTOUzQd
6NsWqAFnuufmeZBuJZDe+CSwiT0o+pxBly1z5mtYlnybb4oclhQv79QajBlluIPZB6EpFj5tUAVh
Zsl9nk8/fBRZnuU0UI33LkRPmgEZz28x8Yfr9CAxz1LS7nUKZGxHxWlPOEempbIqG0O78wKGdqDz
ziJUv2LyQ58tAmhowQfF0/RubfOXeflXeVnJrHEJAtQAEvVjTPc3ik3j6AiRKghzLD77+kWEEW8K
Ll73ueh3mevRuXGoA/DCantWI2+yTzrlNP2KUEZm1g1TUudtJ27Z1Ul1mb/jynAPaC3GscgleEg3
D0JFP12HPt7LXZTlZKZ4SgVIgwGXGd82M29jEdNGYeerKpZmdLZbxxWvzZTK6WR7HE9faLnAynvn
S6GSi1y+No+yqe6H8FtFAnAUagdn6y24EzZZK2xeYbDrhbs/PzaBjhOw086pDj+f4LvN96QkDiiS
U3JAnsEnzrC6aRl9MgeAQU1IVvpZ7GQKhOZJgBTPr9mQLyYvlYhZrjPT+ER+lCw+57qUtaeSvMjO
sGiocjZvggmsT54PibeZp/oJeAx5DJiPqq5IOmLNK61wM0UFnICR25BtVwgx90rvTUw83UpW4HwH
1S3x2Fv8eIMCZ/VZp2fsIGTo8olE768AjSdVdpuU+x9JZ38OM2vGdN+dqmHUrpG1J6RQnljypckd
v840MBC1xGA/0/VJaiY+0J5CO0t/MDfObMelP9aTUaH/Y8gFCEE77AxU66GQ1l7ryss4cKEn3Q7v
rgxmLqu7zJS1TyfYUS41Yx3qAmOANs9F4H+PQkav0XkmEQAhTFVM5kLjXxVkLicnfz6EBGCvgPqJ
k7B00pqeGy//4MbNN7mP6Q4sOeafQHe4m4fIGSodZ2KC58xqJ88XSmJSadCA73SKMQ8JeZwiiign
fMXHh4AJAXleT+DjJ0GdeCK/zkBzJUakjDJ4i1CxmlKcgemYzuUoTNADwgMzhxMVU9xnbeK0FxFq
AJ36JmwIKCCqIE/SFT3dXq41cz1olU8l+hGET+1OVnIZIZLds+xO2vXcwkdq62BFHPO+7OQi5m7A
JiiY3Kj6d9HAB1BOEPSmPMTap/4mcmIG/R4jPJ/eo9KUvmWdr8bdFtrrYdzeMdgPeErCDnAR9hXK
Qla3B51VsfEGDaCvF1YD2pO6ykVZUoKWdakMWjbKCY5LBNu1tPQT342DIUc3avY77R9wizQ1UwUC
P1dxTB2macS2YtyjznsBx5lVpW+I+h4dRFWeSYFUTSqKp+/jxU1TOGi67SyrWvCjyjo0F5Ef0HmL
IgboCDcfz6Tr0hiiZ249TGQmuUkkL5JYRWAhPm3UYBG7DMypDKAWH9/jDrd0MHLYHTzStC8Bk8ND
uVnhA6q5B4zVQDYdDSHreB6Rcr8De2xeFa3bYAvWUq/uuP7s8CScPRdmZGj6b6Pe5ltgu3jJT/LM
gV5kJ3gYK6Z3zoo1JWG3jVpcVSv66da1+CBc3Zu8uo1jtgdWyZCE0Urx9FiKPI82ipFJmbbbbAQ0
q6ZysgJ5qAaWdFCaVO1L8QfW4P44JIIrt2grFZ8EE0++rKAaT9kYyZOLADKLdJOqWJgApHRC7MTe
iex7JfreF07nWW886ECTiV5ieTkmZyDZSsWB4UO817hRlkGM5FZ6TbR4UQiL7ngmRjxhTaiKFlIq
2naIMn8nQV6Ajky/W6Pi/IoJIYAKVmKNu2NK4DSrxKNlbG25zh4vBusErMiobQESxC6vPtlkzaai
iDaxoA0Km/q82XMyJg/FJwlbYvXanRuRdzxvck4yxhue6rXSU8OqUHzCQ94der1/bakyyF3XCM+w
JlE4CCd09QEvYIMC05BUgtvixPSWnn+wKru0Dzk1dGwWf6Zv+UEfF9LBzkU4SRBabKGPY0wrGB0/
xVzmtz9xsikKIVad97eOg6rYI6f/tdJRrAwHaKNck/sCOc6oWu/zRZX1AuF59YL3X4z2t3tkRwtZ
qjo09LhAjmHembXWCwhJLE7n6hfy66X2tD51CiAzpYqWpjcaCtJRZnlysiuSMUYjzQLCUHUqKxKi
mYa1Ln3gXZ8CvLR0eKSdzGyZMZOkhr51HGK2PBSi6qiTEDGXgOpsbOCw0/4Gqg2ApQRPUdgsDeLh
W1HplJPhCCbf3REBCFOkpGWMr9bc9ejlkugjcrV5Adt8GX2vVFudz4J4v/gpb1MapkXhpQJb0pHo
LgNrj/oDr1Oz2FmuoSfiXYmM846ZTpUZ5EoR0B5l/32FdN3V4WhSEoAKTne1IVC+FIEDsAtyvo9F
VCmIaP3yPFmU3HLSjnaBHtnIzeIipgFO6c3qdrgJdxspOBUWaDmZtfpXQYTj6yseTxWJdQmvuNUn
hP+0Ki0HtJAa9HPKd/XumBymAsLiJ7lIn1p8+qKQJGX35PwhpZdupptiCB4FTG2uVU8lEGZaGEl/
bdRjGFdPaB9PR8F9rvz0De66t+SIgjoGUCxtWrSCppbAytCWnX1NuftwSfG+SZNnFc58adJ4Hxr4
1/vJ2rQu9uera3lUB9bRT1PRb/digRez3ehgbeFLyc2Od4iHRNQP7b4vyiM473dp1sT480sqgWcE
shFvW6chBXSv0DlFEETpMewh/k30/lIBCROQ7YvRGTZ30OuzLXuCgOvqoICU/EoHhSEDUDPhq8JE
NNMWQf3zHB7Hm1HXLxhvkGbSPgjebcXCAf6sIrIWd9fLNKdNX6BTJNWZIbUKZdnTtbw1T4JUq8i4
FAOWh8Pz2l9mQnPD/pBPpzAQDoZI1Y0IMQeQU+XMiBFw349kt4Ttya5w6Y2w2o+QkTBX+4Q5IWaI
QXbFa3yg2L943ju4gS2NLfz7b0QLFBkIL31wBetAO65xKTvRnIP+1tvGftHL02DR1jpGND66WGAT
GtlCfp/vbFXQNB1bt5JsFfVVNRQ23hbU3EJdd/4LapSimggrIXsKh8EvdoupJQCh8CaBu9h6wpTm
1fZmyC1WMynDfeErxjEQfNr20iamrMOrmh9E6jjOF9ekWblU3TMaC+NCXHGFHSnowOWhJ/8S4Gqj
RvhS0KCwEU3j1GMj1Q9dBkxIRha/vi2GpnrqU0xGkrtEmjPJmZNdCfBTNHQ4hgYkUg4e1cVsIpVE
W0Pl04fafaQ7qwmUahFtF+B68gtz6vn4G9rQJuA5cR8G20cC77TIu06qSPKys/LL2Ra1F4miQmaq
OPaELnbPHVP7IjwCYl4Tgm4M/fdKVOzq25yDw7B9UUUTNQKhJ6B+GnPUx0kaeCG3r/Eu1pKn2WxM
Ip2g+fEvHpO12HSLJgrGoUIoSYPm/CGBDbsjzvY5ch2EGfq9rKdm4Gd3qLyuBg8UjqAq+ilNuCon
f1dq2r6Vasct69sO6hsbuE8IzQg+dpVtcBjzdM4j5giTpU6k2FKFbsz7o1DmpM0i3OuhHGY1n49i
pY7b5BGDCO+4X6CTzsBGn8MkPZmtL52kOYjT9LPnNl9+JDrEECsCDrmlQSbAAoZ/SDqvr+OPIrMq
EpXo+jbCIEsRQqYiZuyTZL0eIGH/aP5/wdCmSq7uiSp1aAx9MBJ/PNb06JlM3LwQIjnbNV0pM3lT
A18LOFdiwMh0/1sHfF8CUUKwNYIRlg4RMgbUKpMhR+RIp7C7+ci33dRc/jaiiQO/u2P2enbS9/0x
2PTBuxmcS5ivYTqeQV3S95sL6WzHOu/fVHCN8LqLV2wugYatWkCxOtyXv+QErC4M7KnSN3ccfj/W
VoXQWazzmSfci5kAARtt2gLIRMTGJN5bNwjrFHv1ls6v5Q37JKazZLmmxSWKlbZGpIbMru4t0xkE
ukEoEZ1mGKm566yE3sNq5TkYMfbbZcyYLRPCCKtoU7hN6n0nbEujTsS2cICgWO/r07WmMJZSGp6T
2PsB/xxS1z029T+UGQC3bvIfge7tLoU8CRLpcIKJGNTtJ86+87zYGac4JUNF+utksDZsxq1Mpn1b
Dj/9AFqyurga20ZnwOd2E6vVBVGD+wVELlEhmYpSVLAnHKNpnFgkZwVSWWkW+zc71vrEksFd0a6x
jq9P7tRhJyy4X5EqERDNYoH/LlpJAZuSqHiJ3+VuZK5pfhluojrIu4jz64OehzXc9orFTu4APfDm
+eLyWKakLfz+WxGt06iFlW2VcqEGbjByFlGYGdkxE1aiX7kUdKv0Tp9RuifsPUxk16dDV/JfB4cn
3j38Gem6jF18aKUteQLQmmils4mNgzMvVTeLlmNK+qqnTnPdfDX35LBJuS2qBTcFYVYDdagTvtrV
QMArEN5pzfZF4L/1CuH4CUNB+C7tASS3EcK2OOQ03dh3ua8mFgBMND04uUBgpSwt/OqJzUfguzZ8
NNQhyFJXCIMWWRRepJ7/E8340++Ov14Z786Pw+5pN0tgKW+OmWOig/bIFfc1s51hJgUKF0guDiNq
MIbXlOqtLTa/hzkpSlshvp9kuZ4O27Wqp16rhvIRvVxqqSPjlDR+39ZhkgskSBpJn466NHzMlbiA
TQ6J4VBQ/Q0Jod/51Cw0sogh0NLWs7XPQa02sAGKJI4YU3YdyVG+GEBUKlINCzNbeo4oysBGF+tz
zK9Ex5eg74yFJgrIx65LiX1tD5Q1krszplHID2ChpbKsYdjXBIFet+hkiOpfKBZC5S4/rzXeFytP
76F4mhr3FAY8G2NvRXbtzerkBSnQX0DqwnWcWH2Wcq0eW8q4hDUOAZ+an/DCNy/SoIG5NiV6V76T
U6JBh+eu1mEglGMvp117XWAM86FzNzUzqPy6ibvVK6K3nJjxa009yA8RqOseI5F/Cq+9tPMiSs7a
UlmJSbNNvMSpagXGqwK8Y04y2cc8+gSu3EPi4duqwa6O6i4JlR1AmggBHJ08zNDE/3SnGvfyHTkR
aSoY82fdCs2795gQwhR4Hvz9rWzwArVKBFeRVVmCBft1jRMCj8JpeymkxHvaRehNGiZm4AhA9sFE
UDW2cxbzNIKtcah7lOrZkV3wOlw1Ufwygmlx568P3Sw9PFXa2RRrLGW2TTpBRL3M2N990HlQROt0
/5fEl/zYYz1elNgkkHBGlixlr71aq0LZ44SZ6LqgTvgCidOBDbTNGti1vjuL2RsruM8iyy+lH0j4
rSYbOyjUjbqDKogn7tyJuxGqe0ZLvZMPEvjeA28VOHWUcRmsVNSkATnZ8jVxQ6NigNmNHztxYu9s
vW4B38yAcUU0I7d50fEH1ZSMQ0I1WhkKZ9M/95x4BaryJsDxC/P2+lvoRCmNT2I8/XYPM3If6KuP
yZGKwd4CNzREpBxjIWHSdmtEFK+x65BOy/Bhex9xCIP7LvTc8QZ20oCkmM+44Ymxy3oOXP/0nurS
GmqjwNWEftO7I1patOBr8ZbTCYbMSXX8hG5bvufVrf1c/Fpeqzw2RH5ASryW9V9ADMiUXHZE+v68
/fRz3fZpsiUzTwXqMCw6Fj9ur0a1soX31KFSR2izAOD/RQsM+UBlb/DOHrQFHB8mH6EDaHBJHrz+
XWGQXNDtrHS2E6ETujPzHmdZD7A0xkiKq1USBHWtffM8iNKGXORhh4KrNLQVkmrx5i3wfS7E0kDV
DZeLHzI+7/0sWxFSDjISswUpCbxlNFvZMMCqNtYzWwBnsMJsDSmwRoX8aswVtJVJcO32ynuD160r
QcMXjpCKK4YoIMEM1GDqcobxYSivRydxljUo+YsT9xqOmftnBjqDpunQF3DCOgWhwyZGu0pETc3V
TBUH10Ox4P7Ouk7lrMTmtfO6DYGj9bfNxYLBJbKrweLX8Wk6ixhLE6WB0KelaFU7mx4NM8Xrn6ng
3WhXD2ANeQlxIU4W74y6QQX5xV+ZlZS3wcwrJ/wWUzo/usqJta4a8JDLQvHZEgqLHlzp6BBUlX41
8AnO/o8VgZSvQk0tOe/CnyoeCpUgERCobYOuhTam2D7QjIPyNOzT+a1cxPITSQFkFPwKPpgvNVYU
GoQ/ot56oZ5rsxVBjGSoDKNF9Ui5ZvQ8yB9uxJxYOfyolW4m826SLIIt7Mq0QkfwpF9haCUkFP2i
XzSoemwERqol4IKkKQ0/otqepggG64Ne+4Kc8FOyVffAYXgUa4zw4RPmRSotWTRqmdrpQo49yEVc
pCYF+qQfFVNEJH8pQL/4k9i3irEJGNvQSeomFKFEr/IZjLRh6RXInpLRmX5hN4T50YvfrfROOE8I
eIkS+7o7Fs9lxOr9nIE0f8mhUUJxO9AQBdLqlsTJ0weLE7ke8PaVrubzcTkVZorqLsqNEqg3wToY
Mw4FF377ble/JgsE+9MiQ11gMrC5MXNxVa+ydNYft1j2PQzZA/GaH0+umfVOxcoCCJ3XlZNRdBFu
aKmrojNb7DplRtOtS6zHJ+NffGo1py9vz1WorOTFh+nl2YdcHp8qN9Cx8TdZyTlwm+tcHgO4OivP
UVkXg3DmbLeO8J6elRQEp9OjmM8e1grlU44eUP67NL7cRfksLK+sfUIoR63qPx2yEQuRFpjvvmA0
C1Hby5jvF4nO6Cc4GHGd3y6Kqpab3OT53JL89ssR2h6CDT9tT5T6JfyBtJXMojBYtDDQNXDluLQH
5hH9WydXTQenJpEbe224wY8xojXFvriuSiMM5LSR+RzypJEAGwXdtkFA3lLghU6S7dWX4B99ijaO
AumEwul0dxiF9uvcXPZgcMumvWVWL8H3Ik6fBMNRM5d9v2+Okd2+fNYA/WzRWwC+AlmWfwJqBdoB
ydQsTbgNJo3yeCTUv8208nhVCKPP5PBOkIJwGwBI2yvhMPqfIoeHZvOWJbMUDaSWTivt2eTWEXzW
DtsdL3BS1wNjm85JhEB5VeaMAgA0SYVkIVfsK0YhQN6LyCbU+cewHrXUae5dNH4FP0eldLCkB4Mi
YV+Ldu8EP0m0yDMJMr9hvfOSthZN7JEeOX22n1QEdpK42G4TdLFEcAjJ38qPJahNIcSRLDK7hgTq
PcoxUC60xt9JB1ZiGJed+lka7mWtJx/mbuamZhKDZgilJCHUPV4E2Kv6EGT+EaCG+GbBre4yP/Rz
U4fiLjkynRRCKwp8QVsYY5uLDz7j/mmnAaDKIyTIR7tD5SeBboy0Du1ivAInPpeRG4W9MFRleFa5
JvGTJtGQK8kufIZi96DnL2IF0XGjZ1UFjQgI0bBm/9uObMihtKa8WJVK4NnHeSkQN7Ua/yhyOiYC
M/PWeoPXTRbJH7TDQ/gk7TGZZkXF8DsWIX1QW33OWvQCIlF5E/Hr/faeg9bmuPjfQdPYMnZGYF82
R0xRUkl0rNoozxF+yuS+s45Nz9C2omQ9S7wBSqUnymwpdYyF55NHChwX6+aQ/rh+VGyiXKZVlNtB
AyfzZAsjd7obKyHc6ySgyHcdJ1Xv2Sx0x3HdZgr/t8XSiZKgQxUnNU+/pQ5lmmdQzzcZDcYbD0k6
QzAdED+wFnFw3qrQj5/hE09kXnh8+JSvqVG3o8EJx7kMGA0yEFvPmUMwNCKrOSRuct1kyySQXvj0
X4wNcixjd4NtJ6r4J9U+mc0uvI/h6HpXdkXWMgxjGixMjLSqnT72RQQTdcDQX1BVxhEI/QTQ+Be0
9SoyH6+H8GZAfvtanvtD53FA1iPYzCiU1lnd2VgQeRu2++LvE4CfiyD+INg9PnQYWTfvt0yb69EO
G+Z6ShTX3FtzwW6KBSALZCrmratDlstEFPKYWrfbeB1vWMmAjloILAgAf3rZh3ERfby7L4Xt5gR6
LH59NKDHwxwDkIS+osYgLnNVWRiDVSvTRi5GMUaLPBGKJj+ko2atqmVhLJ7FSoQK5oSrLnjLDOol
U2USCcQbtnhB/NQP05f8S1CAp5t3AqoQMGqqEpFBS/7uu+OoIFOo1s5dDqx1y8j6GT88RrqmL7KG
JyWHGOHdfmy69FrJw7n5i0JuSnI7qbe3d06HRQFCHK9UpQ7MOnoRZ5FK99oahAwnlw1dki03ulaO
qybdvC4VyVX++zcpLJziMH9KJzAXnrbw3UF5jvD/iSASrZDYyNcBNeQfu4X3QN4GiWEOn/GZxJAg
DCZhbS3Kq/pYDVky+AzN1dYyE1sx3OMtj4INVymvZIWNSYHp//hDweARZytWy63NavWV5WtUV3hg
iegzJvFDVNkse8bHhb9WCYZjXzYQYa04hD/SXysEu6ZIcFBxRrp69hH3wDgYrfqWSf2vujOYqo2N
XRMjJyqtJPZ3AdTExESk46tNHIjJfHjCMFecqQwbJh6mZ4Nm+FMuukncsyIcAEYadAbVZd1AHeAI
qrBC8QHQ9F/OO+QoisdFhWi81/9Nx2Ju7X5iSmH8HsERS9KCgJeyjApB94HAOZh/+iC6F3AJf3CP
US5kQSMDBh66oyOBGrlIazfsTBa2B17vbpAK1zgMy17WwnlTpKSw+Rn6hAL0ZsosTBFKeCXvJ3tS
2flw2VExLHgVNrRXzb8bBRotQghvknPNWHxaG31g4EwwJ9FFQ9YqZkuX0gEzNbVKGxoRZZjY41Ds
gvpQesEHQmM0Ts9v7ZZYwbExmqcUaJ2fR46vL3E0i/2N0rmPe9yf86KPqGvgnkaqsycIA50bYeGR
OVMTbYGyf31pvXs8uVTEpKcupu95s2oivbBt2qyGfI/nwhkgsUk+VNTj4A+A5VAp0dMba34FLCWZ
81v/87VYq3MAt+JogdpyNUVFa70iyYC/RVKbYM+eLFs8hZdEZCmodWDvLLY8kX8DCark2Z+6Q/WN
7cqRrx8QjapCHW9Nga2sthHitO99Wvx8AZHRcOjb1Ac1bUqDN2qFj3O1VjFLQuLwCV/NSfuw9rUH
ZNzgStbGmwNWaHdwiflvtTXWhibi3ZUwmYFvKccnr2xUfhNosZ53nLi8ma3uN1lFed0d4wStbu0r
agMmWq2rJfz3ub35a5WqW77UuVcPaN9ng1bHwEQX9X+9vuUuhhu22jpeMcBbdv14rg59Ysjt9eds
MDeE/mlEvXan4j27S3Thv7ejMuSHIgLAJTqvQY9Rj1Cj6MAlWpkV2N0Vqia+e4XFAhtSSGu6IPaQ
Ru6UZRkw5HrMjpDetjW9CGHtZwshJSPTYeq4vqN4LNiJai09yQoqVh5uIQvObBB4zoBW65en92qM
ayD5aY6S5GOd3VXsgpTkzuqVmSLTnoKDaI5vJJxie6PT4r/u+smGnIzvX2ZFYHz5A/z7nC57XwwW
Tt+L13Gjb4a/akpRwuoIjHVj4gQOSBZWhWyNbBBL8makrPUJowkVpQdQI33ogV5l0FauaKnqyaOc
czgcNA8O5bR/fCt/FipqbSSZr5BeoLwqHiTAmdtUsVYZcdU/RyIKcBSIZbGR8yC+AWuO9s2AU6GF
xtdJWi14y8jQizffE6WNWJOsFXEoQcf8j7gxaVr9//MzMiQcF0hDvhDGPqJQMjXuHQjW3Cc5kh6N
l4W3EBuM5un5fwsWb7oB0OQhbApwGrHlNY5aHsw09TlJBOWk96GD6Q7DgAPyk+J44sv62FUQHzCs
8tZ3t+KIJ1wEjRhmetn0YQ20bXnsJGT8FRJOZNRIVZqwpQgdqnmPubXbPSn6PAHvw8UVKXid49+m
pu0KO+YSG43OvGqfN6omb45vo0XCDu+1ljt06sJ2loj/+H5CKZLu6xFi4eWu28gRVA20uZo5NuOj
bCHGmyMulMUuEJmthbW1wKmlIwLutO5v6Tfw6AOwAh13rl11YWh/qJXYtUD7lu3BmAReOuy+o95T
Y3YgG3kJDtOp5G3tS68UfGp5Z8Sql6P6eZdNL0rkkI9UbukGvYya3/dhZkB34ovawtZm44NY65GX
4gIOaewgSvxMuz+XAp84v+sH97RVaL6+JB0vYFT+ufIuVkIRYi914VZY9ZdZFZuyH4AGleyXL30b
IIU1QbabFn97d3IrFt7fLn/2mqrAuxcis/zeX9DbVdT3nbEISrqMaEqzIIMVXoxVjoYVN5L969gN
hBJK4dzfdY6xaaQzkmCYxf4Gn95qg5OzChwnQXz1AvcVIVaigdWW+emXSpxDDt4z6LTOQAzzfX0j
f0p0/69iTFTpayw+yJWPo89aBiVxxDZT0IbWgm6kOVtOvAWmxhII0T/VHBd1br5SBywWPpTAF3OC
mOa0FZd0T9IbpHPC2HeSTllS6HOTmlz76qwfD4I+/gJyNSfM00cth0mjoq75fuPnFMncdt+yfZWW
munURaj18EDiziZF01Gr+P3gudaIUySKAp7UtfpUwU+XgvpD6snqlDWPWDPagbtFHZczMGfykSqq
dkg/XLyzcRo2dvZMbAsZnc29PptTWBUHvisDln/GLDhviMbvjEB8xor0l4gb4VEE+q9EI8znbjPK
yrq0RAheEziY63EiiS6ANFihAe8TLSUHoize5IQybZjF1lxZxWl3Egxe0dhkpMtXfmNxcJ8YpzNs
iLju4UilkB5W+oP4+v47W4TYxAVnD4/y1LBNvjzt4KDE7BAqhbir0ffte3RRtrot+QIJvvea5+07
dtP8gEe9SM1eByoqvzi8eu6F29wDMW0v10Qg1/om+hwDVqrzh4NUZM1H/qKYWZJ2aIkBTzoqCdzT
xLsPUPhvwoftJ4Bet7aCH2qJZV+grVpI5pCjuM+x5hwABOPcplG+dGg0jfJDeDeGujPlBsgj1c+T
295oS//5hpDDPzZB6dP64tawD50SFaczK5fZt2EDLp+CYyr7Go20JP0zmpRzrMNqkWRP7mLSRawN
nUnefyOuZYx90jMWNKDW4UleW3jEE7Fvq4mcGNcMx850WNEBW9zLelvmkdyeQsmIGefcaQoPyhH5
nprKEXeKqPLnVYKqN2VbN25tPzybdISDox6FcNxac2hnpVMs57nOFAdOcLu8a+AOgMtsCHMO2VTw
zbsK94kxvnLflagw7jq4/p1Vi0ohfKm4KyrSMfL5D3EZLqH5Cuk6/u9Zq3iMazlxBrXLGzT7ezG+
cW+hQx/8PtBIImCj5nIQa66Lx+WQ+PPPdBBE7BAXT5CD4V5hb2jELnYCWenYPhzv6LtHynjNJXMU
qW37A+yeIjY4Mm4eFiAMPYxqgLH/WH25CRAK4NAuYX9UMVXaWhn6+DcQj6oMVwMQ4GXh2CIQZ5B4
guyZPDkRmEiWN3mWe5sJOUaK+a6kLrBzbH7ksKsxuZesa3EOvuzeek+HIhR+64776aFXHUD87pEA
0Iz/UmoSQcXFJP915VaMIRTMFFetaCjo3evB9tkSa3eNrsyaG5z119JZirZ8Ywg7WRehLvYxpG8l
BoKtzZuI3KkLeJPG5dmfQu1lZekD+jyaeB9rJfaf214LmOlvT+W1akfM2cKEg2Wcz0p9YWOm/MXD
L7jSuaCF81jErkPl9fxco0DAlEh8919um88siDMc5f+AUPV/b0ZeY6x+ohHqbCmSiWSbZObLS6Pb
JWmDu71/0Q3NMXH6zOv3v3L7nxxRZFfusFs7kIS68nn4UxF61tRu7FQenFcxuz53B9sGrkLm8mNz
0JY+pSTipgRHm+gTtYOtO6QVcNoN1MZxGKXUqilEXGdCUhVwZbDPciXr19W10jH/ZqjNzoxAA4PM
yOZwm+YlgzyWpAevNAHxSd5/vOstl1vEiZE+pTuP7DcVOEMXk3hqts4/NOo8TGTywH3aZnjW8d/h
HkzvCZEFMIy4Lmf7yFGENwp9dMkcx7u+SRe05dwtP3OBcSIvCtcjyIvZSoDa/ecO4kKwKIf++NWd
+fdPmYoSm1x7e8wP1fG0hXmVvrks/I4Bgr5tamco3KQ/JZoxlo6tlBgwZnADgT6KwYgZNRxA/fHt
Jt1k3MliSPbSUQIHJGH+WvRJ6gnYiVG+reHGowkAgxHhZ0IWzyTbWM9PrXofMEUnVYHRz3MGYXyB
lsSuU8fl+htpQN4KRM2V4vWIQHRn/FM8ykX9qwEvd2ISV8GQDM4mVFrlE0UKYyZxMnmPQsVx8i3A
0DVwYrYp2XdMk53NMSF5+nrKsrM2ZDtPySXjx7N/cOVaU09fYSPDhglIhDC/4QfkR7DHzoaKqRtM
VTdxnQoXubYfYb2YaBLhxqlROhJ8iYjynDFNmRUwK1VHmGL+o4hNL+GFrePIO51IOawPYC7Dk1ah
aBWsF3UExlxl/Im5hvIy0kGlEOrwiDu91wZ1FRe3i0lxHOQrzl4/ehAsIliSTHygrFnY44ZTdEZj
vPO5N5J8z/i3DwGfAs/yRHS5Yn1DB9YPQuUH/IEwxeI/+DFKMJ9pKo23OKeJcqQTvzQNnKjA/aVy
QcjYTAbzxgqo/HMjW0POWRymcS8/g7SjoBX+Lb+jiBfvrF578cZy1Yx+p9CptD+I2qLrIA03F/dP
kFFVXtarfUpF/dheFTZZsyFUNrilt3ioy+ODiCeavED30Yk2P+QQsqVIqQgj8dG/gWMcRe8RtwXn
relPi8E4j6TaKoshgNyjdv+GCy9aGkBimhThNra3F3N4OL6+Zh3Zaq8i935iuh1sClK5BGJ74Jgo
293MgHWe7Dzt7e8aQzC4YNjppAFm6gcUQ/RkTSmQmfAw/mvJmln5vF1aUfoHvEPhQURUmGoQerF5
Z4nD5CujC7eb9a7SRESwC3HhboKo1qNYN2c9oGdHL1+OgHOj9vY3GaxJRbW4yrg57QBi+WetysQ1
UURH1OzZ02zRUlTDyxmWIRTlbtzM+Hv4OWfWZOS2VazPgFRQIThBO2Oqa0o+59lVwuODj8O1t/1w
r4fmdNbXTAc+d84kCYPBBbqvJrZHIdaLJRzZxMnNmpDLJiBn1GVA7wkKXc7Wy6nsvrRo1+f36P8H
l7WKEIw/4KclBqkfio6wYZUuy+PxGcFl2/JWZiJgPfgkIMFmYFX0yzOYUYCimKoNUFmmsDFkQ5kQ
mWT57xH0osJU3x6yGFS552YvxBNfUDu73a+qmCAxOWdJCjkzPoDGL5imqXUvMLEviZr1s4PcP1WA
yeGhMmh1wgU0zR7iKhYaFXMavEuH1t+jQQcDPYsb3odEzWROzVTe0NVFJismaU3hosiimnYF+3Fj
4XQxrlqPyYa2aaEhBns137Uxp7mgNdKTdpjPxI7UcxHOA/nu8t5f9J8Vry23qH6PS/WtlefIoiyz
Heh7QhbC9t0EJYT4nnX6BWIUd7BicyUcgYI80ywIW3Fdv8IhzP8qYYrJF8heTuD8gWMC8duNtzSf
cHjjM8Cc2AGBoVRkorkQwR7y2z2i4FCzKxpx6Gc5wibjxS0oOs1LlTVW8wza0LH/Zhip/8u9fFph
fozZjbZO5V+Dk/rGM0/0MFmNCtT0DOAJHvd9/eZc2X2jSdtKoqatCYg/GqmBO+9Unn8JRLtClidp
qwK029z0q7hxc0QapLp94HIl8PA+YGX7VNHk1h6jH8sNIzFFiuyPKuJyXznO3hTy5r1LK+u1CWYe
3dIbmYBnSib23EsElLo7o4i2N7CzQ0JT94RroZrTFoRCqd9UMhqKsUgRUwQ/6xj4u6Gbsk/6OM26
Gkbh8z4T6xvC6P+60GGdaBzLn5JpbSwvvO3Ok+B6VbPHyA8xXI5mMguqiNHrbgXIPNnYLAQ3ZyP5
Yb9l9PEICj82Asw3VVJNfCFK1jyZa4Q49ovoRcfHMW7ENPsnSXfi5OOI85eiBDqOJL5IqbbXdYhz
qMZRTE8Ir/9KCrYQBg4JfS0fwnQdBliV72KAkEg7XzcjCvNXWFZVNaMn5wM81hlcO9d1CjPPfjcf
+sSNF+YNiYbSA3j7+BIspHYadabseomL0x84d83Vboolzxn+sVM1KmMsbKoNdIPX6mCy23CcYVH6
+3CgKuUZUl0UuqJaaQl6FOLDJ9ID+fqlZZQueu+cLrZHgpb+aqHKdMGpV5tDhwZH2wjc8ocwiwjM
Xi9hW1iVQhG6ak8gHUo6gkSRC8ZWPIrIgjBf78AoGKCFI0zWyt87vMQIk6j3NPYfYHXBg/yPdB8J
bWtgmO8onzqQyC7uEW3GsMR1Qs01WTvY+s7HczgEqVIV8tCVM4nNkQI3fUd+qsUlU6czHrMXIvtT
oAVn7MzgeFS3xZ7qRyHdkBEUH2XBbk2PwBHLixOHYgQQOvwI5B3Qo0Exbf2h00yrNgqLROQPHVOl
JC1bAymVi6pYF5Dhb7pFA2AVa7ejlTkuSZyExhKq6Foo1NHQYy2Z8H3m28LHvvt5XT0tOal8hYFy
hnf9lzffx3xePA0X9E5j5UVBHY6k3UhRqlBHvPvqodCB+AUQRzRCtcm9DMj32njnPo19ueXAdBk5
ILVYZ9bRTG4Cwf39fhzuP/AzMQH1NFr90KCI8PYtqz8BbJ4Y1k514el6yhD6AM4+nemjF60uvBcK
mmU0BgVx142gMaUDxfMwOYNInEgh626wVkM1ou1gleG9wNPhDbu5ezJgrNtFzhdyqeKWuYxxlUG8
fpFwwQfLM+Sd3Wm0nE5O/yq5ibi4haNELY1c7RXwrxDZwO9TDLQJk/ELfomJL3FzjUaCI1jGwbAN
n96mLoJQORPD3Shvjh27BGZJm7sCIwATT0y4u9Nzv4/JUTOqWLqbfx8R3By5tbQhqGFXtwUAQj7I
L5981nInA2IsoFfJB3FOeSP8oC0KkgZ2SZ4gKKgm0nrRmLYElRCcdhezL/tx/WJXdiGwhlA1Oytu
fJVfzqObjH2wjc25zBWlLJiNm8hDQwYKde2rbJVzAyk2UJSRBwPIZ2bt+iAjDH6RWQVQITOx2iyO
E5yYQ6Lm63x3cYsN7vwa9JKd0vdIS4kR0PUccAhpMw/mU3UXjoe5LSg2CQJzYNNMUaqvYd/ivHIK
3sDv1+LnAMLinZ+Zkd1oHqXXYGXTX4l7owBTDjgmJDNGvilRkk/Sr7zYP2Mj+LXiRTDILE4t0cfy
TKjI0KogIxhlj7OTvgRbxme7GR8Gc1C3BxKFtbzfw/uM+P8q54S0DuadENJcoucnp1meN3buy0xs
Qg0sV2qu5i1OBws8I4HXapK3AWKOvqAJJh9+4Dk0rGw7jBS2ql5/4YWfL8exNzNFkOrLV9jzlnc8
5CDgsUA0o6j0vROvLTrfStnTvzhpkfUuL15tDgxnXd/H7nyqlIslM+CBD6uBbZp4HuIQ4VgKlMMA
uuzPxnYhDGRGyngWD2ZGYRIYrH2NanV0d8dCTdkQOccKtxb8D+giFO+9sycvYL8d7v/X1M53An0L
hjYjAbiIWdTM7rJr5TesBEP2qwPUk8zP+Fk/rT3Y58tPT2LG5C4TLgkzfc9FqJe0qrl2mM9WHFu1
osxCSItbcdvsGbWcFSB9pV0heJ0QMHLqycq0vne35ssGn1egkNm1Oo/yo1YqL5+8aKCIt8q2dzv7
zYlgPpFQ+sKoY1tBK0bXOM0iUZL5QGlbAsPKC1IpJowxgSqaKM91LKZR0rpgky1oO704YFutU7pB
Gz6/1fQbTvuGBPgTfOJKpEejK+9yC3L1gqDbAlqt5YIQ63FqjjNJYKIuzsUkuNG1aTTzCgyKsRLN
+jJM8nk6NTES6KOMHQO1FOFOj073Pmg518zstsG2MCXUnqLWlHgTr6rtdU3YTlLXwG+BlbJ2M8eV
Yd65DhJhP5ROo2//4RB6OLSDWkc+xmSOUEI/ZStjXuMNR2KClUlnqcp1hNTgoT3dLApoL8tQ2x01
mf4kWrYWaaq7XoeJCY99ZHovYyUWBZEZ7mpQ+4uIxktK5fwXdydl3ecnXhof0pd+LDh+42opjtwW
5iK6SnddGSJfGRCkifwHFq61n0fx5T5KDNbIcrvTPmK0rTJXj5ttSgZAxOEaBGvLd8p+BJsH5LBF
+0tX6ARmGfO8ymLfe13BQ5uMVu8gtelIP/HQ9AkYiAxQgXBrcPe8nVqz4mIk+h5q99TPuPaodhW2
cT8xka2rVUsEerDatVLGNFy6uo+vy2uTAC8bmISUBdI9DExzjcG5pC0vZJ64XseVKmmtdQ9j280s
75uy9jE2QHVjRFdYQ6up4cx/ypcjtye7dVt2ENb8wF3QcVFqNS7TyGMa73hYbwNt371cLn6nFjDU
NH+8q/QF/TLzHeesb2aNMMxDlJuLEh+dhHDWc9ZV/f4r05VTdy+TpX7tQkN0xXk6G3hmCBDh31ZR
NMD9djxl/OOiPtnjIJ+c51Epz/5EY5GsYFM3vQU7M66b0j+YEAAqQrixFZisyfT+aSNGwFiZiDYu
Lt6czfs7ae5g7KrM5QTQpJh+AP7dB8/VjtUs9aIw2pIxQ5y63LPaUmZaCg4swlboAD8pFFhb79cA
PyOKDdmj4lOMrCpOLlxCUJiAe98VSp3ry3xUflxKBQzf/hCDpGTKn46C8lMFxZOAA5Zz8NSkGpMm
61ks5VfbnXNpcF3X7/Y3vJG/zYqh4OREqJwWPIFl1OkQw0IqafflE39hlU0Be8iIyZKAGSVS0Di6
YZBntymTiVGyvH3YqBelAnS+H34gTt0lpprhvRbt1okj4HxfclLRSjGCshoYqDQVjvqTvpzi6wq9
3+0+TksElCQMkaA9H/gJnXHcwVbCK0JwmOp8Q9znc+ZQEhAENs3RcTm3VANVMZf/RyQFKUvkLsEy
nTNU2ajNfzAMwVQOY8dxYUlgGVta6noIKEybdQdaxHQib8xFVbS8raOh6ELdSVigY34jolBFrT7N
Pb5wx69UE9AzfruGQgBcTrRCBNPZAO9o6KA37yd4dPPS8sLQJm6q9tOkRAra9wXflAX6oYHd7L6N
nGIV9dDCpnvvokg3ouUqQeqEAi2QYPRn9hqLlC3v4a2G6eWgNZVKwBDKZhvOeSkdMwDtIvhIK/yF
X+E25qvklWWUrveZYFgaAeHi8RIBc+gkYZEbGGFY/+JM/2OEjYMi1IYXIs0SsB6+hje43/5shA1q
fCBdUNmOcIXjQaTxCZd++jGg/9Tsr02WSU0QrhvoZZv8iVJaLO1r7Mf99Bmp+fltJ+7YZRPi1LEz
+y6dSvLwn9eOmwi/UtYntqIza9iob4BNskaRlxVEZsLGk5D0oqEkE25yKZswyf3ohfe8ml6Ebcsp
z2YPb32bwK9UFPQETOQf1vmBBFW018HEpxzMjFAccTXZavYNuZFUCC6i/j+7/LMiJasnTEGNELnk
C/ahIIPSLixt2dVHgcCPg2Hikhl0sh723fPEOSOEFunpH6880uwND/GBSoQutIVUi4mr1NHL8ywv
BybdhcGWyh4guQYt+AxFTDegCd1BIuMzwnm2dzhabGON8fOL33xVUgWnbgg90mYu16+dWJ4gLRYz
OV58K9nwPwvPlV7xSmMoqWbdDzC8ID8bPyG/PdofTnswcLWnQwT0bAyJAKHuG8aUGJfI7cLOgQE/
IynGcdOjK9ITJua1xucS/v7kDsTUCHrnxQAQx/d3D8vyOwpMCz0rVKyCtG9zrGc347sWEqGPhWvu
hoExFLyPcwP481elM/Avg1YksGk79kBwgpR5OtwI3f5ZNVjpaYrYZRJCU+clXWfuGKIpCDPGcWnj
AL6bZ5mxgThbr9u/snGT9j1IsBLSV8OYISKDX6ZrzEtOhgDgPyLgwVAPuLinkkxaSiuqACQw3YQj
XtmCDwXpyDirPZYxK2mcyLjuj1VQo6apm/yUxMUnvRVOmrl+sWwR6ViZTLxz1iPUgy7oDueASzlg
5+iFqkutF1trrDHw905a55ZwOzqSIBG+p0dmTbunAx+tK2HTjLajmX7Na0aKdBT+7ftUirgzy0Hp
i6m/SXrRTUM1hG9ojL9xqovITHKut8Z0kmfd7gSXoj2eLNp7t/aEbxgkdivMFdkSbDf/y73Ngo90
9rD+uaju7zaZYJ0IcW5vd6bKJ5T07ILM2Zt5OPq5mBrGSSUIiBZDhzRi2Ywrdzujgq2dwUigLfGv
TBogh2l8P4p7qHEBBnAezL2T7CUaFMQ48ZQXnoxQSDo/eSdsCe0brjSjh3c6FLcR2cmzkEXe4bdj
iyXUquv9sMGaxeDviEbnkDVMa+GgvsEnENQDuG5ZdMGfzmn+jZ+66c1fF0jNC3vfZji7ugxkX7d7
Ydb9hfyC9jAnY+Xx9mKRhmCUXMjuZ4NsEHYQdPNSUV4YWfhI3KqwiaacOVbY9ZixPb6hZXvTWwUW
MKMnfjRFsdBk0H9NDVz50DijN4wu+3PXqhagiyPm+8JRHR9zaGS11lYz7/aMhL4ztjg/c9vt99/z
2Md2Wy6Y7zSL4vCm3w2ozti4kQebqU7F/uchO/G2403GW6LVilT8I1m5YtmXFX6mQK9mavwxZcQ2
Dy5LFXsp1eko3KRN8p8+7ekFBsXJLxOHVOTTreHap/yxXSm1CrC0ghMzuAuJtzXFVYnm/W4g4JNz
kTyob8VZdK2rdc/wr59hi4Pf8GoA2G4HGrbA+p0Re7TBT21tjyfTD0ZYRw+44kq2pyXbEmpcy+iK
E3mZEmMKmyBF/IRhi0cke67JcmG0K5yenR6orvq1Ha5DIibjQJ8tm9l7w1I8LLR4IoTlhMKvE+2O
4vuPA/APwDn1spCkq+7lAASLR97O5XaIOi8INqUX7yXOrM3612e/3fkdA6XHUDNXQEdP5qZtfpS7
1gVI6Jv0tXBo9fTGyK/4HXQHFmMD0h5RRRhIRUXVpC0glChxzQM3OVsAYCpqTFJ0nygLpAZ5g3x7
RcV6I5qz3yjVV2pmTcE0CdY1cJ/PLIpzpiPnJv1INi6+3BAeIWgUd2y/UPKUS5Aobc2uFDZ1Jq6G
RetxuEL/byEa6/DMCYraQrhjBojzHK6YmpCOKezY6jgNTinafHZHX9jXNuFXGWxNj7U/l+mT/RKY
6Cw1Nrap4WBtpv7jPLyZyxN73tdtsn+lAEnNYwkbL7U/iLNnSS3NFAQt3yxg0YlvS5ufmBp8O4lv
YfqJ0r8gXpsmW1X6d8h+ub5rJ6mtsOEjcAwcm7QZA3qIE+wGkmSUxscVOIAxwOURUENJggVdJT0b
3Y6rLF42DWYilNYkDJ8Qwz0LwN8k1WkTy0sMgk2VjhdXnlu+4MCLcyE8rWIeEDEDc23jJEjVExzc
+5XYLIMk5uAF9VNDuCjiaqwfyWXD39twsYxv2kzbKQXmN3sDElsKshw5tTPokcibUq+/nvwNxmGd
ULwcOCRXIXMzsy+5KgWN8GqkmLDVCeylv9ohHL3CvsHALhjuMJ2XlaMsuhoqbGDu1Ivkhsu6ICHx
qwEWVOcQ7ASCHL+cY4goloWIzkKNWk2dLc/ny9PqfLIcbke5Lr2sVJGwiJVTULZ72pt+Npy1Q/qR
8dka0l++zPpL+tG3THEUjCz8X0uzquyHMtGAXSAtqWBTKDX7GwFWTcalrijqa/IGBS7U26bX2Tgb
jqK4OM1GsSJ1bZDxwWI03CBKhQ/s+7tSXLPZ+hq8x/Kes8LoB69CHSO+xbxfqYUHED0XsUsG587i
elzTKXpbwHNHaOTSNKS2wyfDtH2n87k0wIB0Du7Wus2aWKhh5MKxWUzH41iBUhCWNiY6tKJLR02l
nQXeW27L8c/sqwHFpFDQHyUBiNtjcXzQD7IHhxx/icephD58o1Vdui4mtIA5hq/TbadHzU6t5AlA
2M+s6CFLQOsK1pC+Hc0anYUvPE9yS0cfV5T3fCpiRxeLFjTY7MpzW6wIgzEFibG5Rf2KEzU1dyHC
FYUMCJy3XUrePEAT7Dqt4tDNKN7CD+15THfAquUbzHA4MaNpRH+D6DfuM1BQvcB5XQxa2FoEdTFK
LCutqUqnUd3/dY/qTmtPX9t07URHy5Ipsie+iRux526N8jfnndnSjm5rjDBWPL3mdSlk8q0yOahG
q36QsZp4FaRranGEdlpoSzRls/o5jrLFTh9lrEqMqJxTFjIrjOvsZvMQ8DDLsMQxEPW7IJCGU4ru
zIvWYT9mqJGlzDYC4W9g43G4pn5Jd+yLEFxsdQmIPeMWJZnqHnl4CrmGyu8WPFMBw5jV4o8CKbHM
MV8qhVE1o6KZMd5PsuOrVu0Ae89UNPw3drU6UmiHvpUA6ub6Me8S3Ubavb/l0D22magwyO4jNpT/
IA0ZYlxL4dzOdqGvCGVvUDChD/jxS7Ez8ruUmiIz+RkgXKalhB2vMeq4w7U3SJVpDdJ2TMcFBzTh
GPiWx2OsK7w7W8oVpmqad2wO5EboNdtDSQ8fq5s5+vnT3vxmToMWTSuK1zW97y8+3zPFwJfGURr1
1mLSn2kxxapd8CF2J3ZjpMIHdhz/A73KNfI2dq/zCZKwf4GmTZT9h1keBuM5Ji4fveFaQzlZxhq3
wHRorYwOaCUnHNvi7oplCqWCuFvfbGRljRAelwSojxpLAhE3QQKiwY+XEoRuAFb7pCLjVDL6ydi3
O8e8KsUwtZVszHvGbkttZ8LqJl8z6U5+Rdd/NdTVp2N6sd94kv06FdvVncAV6QKwOomKw+0Z7Nu0
HhU7wYCRnkokq27KmOBMvcBZvvIImObuOINe7lAaPz3rEi9Di0+t6MfRG5z13/XpfuCLujVJxAUY
VW0Fk352WGyadhP7ZUgdyjFIXuJWeqqHi+5/xFTcggmKMSNDLCD/HkEb+zdGyAdRS2nI2+cDwYGf
RLRQrxepcc5xgyZDnxLJHm60/6HNrvRtXkqG5lOhnvfRJZKzqXaUQk2zqakzoXWzzeRAFVmBuhf6
Z4qLrhUEuo5e38QLq8LrmEm5rmKeRJTjwhLymnbPmPi5Ba7N0uFu9KNce6bgWs7i/xpzTX+YgwHx
UDuaNRaQ6DgbaT9fO2mfmpgw13FeL0y0YY1fqp8z6JhPJDDuDr/WK0Qtw3VjEns64FeC6o4XuSjD
6gSQIceDJDcwZlMr7ZQM5I2iwW9+PeVsERcVqHerv4z56Bp3XWBjvDMmLIlD6MyzuKyizd2OMO/B
4xXeGQ1iPYajORNc4Ioxpd5msKX3EId/i+Un72Qgx79mRLNu7a8Vca0kZ/gJVLqowkhOEQnYrblb
BZZXAMM0M5fObfl/AemhNe64C2z/CdNB+uL2A4FY83EhCF9eehqSVqTYdC7xK4JDni5EE3fbUmLw
CvY39jF7c+EpIg7AS98g2RG3m9kwdYjbTRAK2IJwBBmX/PtEToGQYQkgv828fR0PUAYaB+Z1ifzU
9ur5kP+Om86ygjxC2zBCsz3yM1NgTXT985wo7Gv2lFTu05CHjhV+sVsAUNGVBdvfZKHWMmkkRLfI
EQsg7RB+jjowuawVn96Uo0LkZC6hcBgOsYAMytmbiNZGwdnaglbYcnRq1cGpKOALf5YXp2NhmMhq
B3kSDsNN6IcWvEOVisKW2mBbqY0Ob76TdNcgbsmJMZ1KWSMAfHxYbV/vv5+bio6eF0x3oUUK/xrY
8r6vycLK1HooL5u5MkJcOB2p5ORZofCH3HJao86MMx9EFEqrw3HrGhDlxNaaXuHHa7LDmduTY/jR
bGAJyMcfe4agbvbT3nMIJ3cB9WOmgjvE4wX+8PVO4eQh3wOk4pPKJVjg/D8Rmwcpux8EpuJpww1w
7UWz9NPJn8+GbDY3M1m76S6tz9sy0vTopBIFpShTHsLSgc0UuraWM0yHmSLBZrtT4u53LlUa6LEF
Rl/8eIu+ZRt3NeRGcSslyKXyQsww91pV12Pv67W7jK97qX3b+OGljV4oHt6xVh1nLxhpraz7RtGE
6iCGaMqZiS4dfLGFsxQvOFfNAPLiJFOtHd3FeLYvxvJmeXEYgXSkrmjyq1d611jFSgBdlOeE0zfa
TzfsaTSfhkbM8zf4i2LBLtPO3XHSX2l2rf8vAS7WdyXPFeJAU89oQI1CUad2fd1SvfgHYV8KPNm7
xLA1rF/HjccR3ZZTmFk4d8RMrME4Uux/t3281icR4sZPd39v72Ba1LnpE+gicUc4YUwJJyTTL7nt
3JodEYxFuExCdzlnUoaFm038oPt0iC2tiqW8Ouy62DNpcGEUW+ISseY8J80r6Vc8LW7tw1gpjUAC
WYKXxtoXHllN9uU7g4y/1eO2+DKBs34YTDA6umZ5pzEfxAJXjzDr6J40KumqCwlr2sxL/Eh4c7M7
OERdizBTxM8i9pQsTr5dw0Pmq6kqpaALWnTbA+htonyZIoD0Z7sfV8W8rhRyYvfwhe5Cfgnu2oab
oqGM1TsCJdWdNufc7rakErDODD+dK2TZYka/F8dC2uhYZnlnaOpBp2+XFT6WXHtFiB0oUnwWukcK
byfsJJl9tcxIElT9eYq4lqCjoZ/COshNdetM8/wFWaPelXpfHYk6X5BqO+q7sSlexZ1R+Tm+X/9q
KvTb9pZewxxH/ebNApMITzHnBz7ZXo8tAi7ZtqXV6A2vGLYDwWX/N+5Qp2OHfJ0S6JQ+0+rQrVZf
LTe4yxCniBSHPI4fzBZ93zr7MVJqxBJVoos0rcwX6KMYVMGrl8mifuya811ih7e43EbdZVJEw2Tm
Z607pWJkKIK8wuNqDNWDijs7mK1rJUSa9Ib1R0F4dn0q7Nf2m6YawpKbn5hGZIQyahxlpRPzfVNZ
D/DFPsjR1zrAwib+W1Hhqvwk+53yStfxu/8jx2Y8toK/cbxie0ZghLxCN1HJbXQU/X+lKtIhjH3Z
4rY+3OXPlsG2Wwgczc7/g5RWNLF84rrJZK/o8tjfehDerrUEUfN5DsVJDowlNX/mdYAtIOsOHObW
VDXD+6UFz7MC6f6wLwVQJD5k2l0U2lhRVuu5Ie/iEI2iGVUqnqdpugzb6drB9/mBEhu9oabzihhu
sXiy2RqkFeaKeOm7VpEg9eJNhuPvuJ+S3qGxE+A+Sfbw2hWT3NKrPGUowdaeTbojOwUc7vdLObD0
SNswR7IT5SqOoJb/Zo1AKdhXzCIIrJSJUMeRmRZ4KGlS76G3iPm6oTqPBoeh/liWje+EeKU1Ipib
1G3x7IqC+qPbvqgCxHuuUEWrolgczl0AQSPbE7BTNsQ18V8kccFeyguTL1k0MNcYLMwOTL9Zuab3
6k2LSEuwvBmxWVRudI9B1n0BheUXuJ4II1mpm8neIQrMlvzr4tzBsfSgnliAWwUXuRinjOnoaWhE
yTGcZMGxuzkZciwaiIyCAbYg1qPwz1FGd+6bU/MHWGTiimpCV8e6+yzfiqpLutzk9hYbx7i3mgxo
P5hLzOWZI+OikCpLdgYPJP6J7ztn67vWH4cEnUcxirsJ3JG58PKgw2+KPz7HBaC9yfbaCPlJjrPh
5BnxNV+RJ+/fECi/LlBHBwGdL9wj/aYsYot/yjLPB4/nLozE7HxLGfcHYW0/rdFGkU1SwxAglAbd
MWn4shLire4+xiNVGUjJsQwzbnJ09xf3t47NyY2YwntzKXY2m9uypE1mA0Y3PebL4tLiqRsJ+MOK
kPff3qdJOEkQDkFhTMOffcYb6p3ulaWC9rcQ/J40SYcK/dCGiC5GmiBmI1pfK0gKbKw2e4ba4dCH
pjPJ5mce2wY6b1NcI1mwqQYGG2xiqZTas3syUU9ns1YCNNlU0fZTdCc37Pg/sav78S0BkEU07k3/
HJBa1fRBnzjhLsuxD+yK+75mJrdH0sUN18yZ3Rsi8/qXtAGLRZUzHSF1StfxaO02B8rUOKyXPuus
eXBFSbiuRPHldQnTEUQuTetw2xbIvtr09TuZoXmtgh4enTmdyvGctrbvAY0s0N8QRbRZieCJX8hd
lZ05oYSpbyY4egogDIIoM6t5PG4gHyi9j8kJyLB1WEDQPUEBvaj9rYszXL23vV3aHwbZYeRcrNwN
Tke7WsAh6QFZ4wddaWoqxUvdYtzokEIZPL5VltGw7gjcOt9sLEkeVZ0PahSwWfGkt9+oqhRrezUm
Cy7TUDV3qgCMxn79DFAuJYtmkRmcHyGRlyU06BLSo8QXcgJ5mNpPJpRKGvViBKqY22u5Hl3nMFxq
T8xUIGqgliPV6OrAL4lK4IBjzMaokk/9KSyTsK8z0WuvrOtQn9tHmPNL56M2gDcF2W868Qc351Je
wihEZ1NWGuTZi1ZNlazpbP66BhoKHMraQgiktlbS8rbnSumamjH4a8y2PWeXMcIAae/8s9kOK2UG
VNZ+4qtsK66Z1Btg+LfaZ3f4jHxGK0D35Vc2fNDDLAxno/+cb4zB7Nr2/67kLR4Md1sCEpVzS3R0
AncYgR2lzgvy0mnByb3r81DOQzUgrPuDp8/zLFbvnwGml4MhGi8OlEttULNapkPTmYTuD+auuDzr
2/MOZLayNCmeeWxbmERgxRzscfBrVmXUzWrpQsN4/4nB16z7qnM+XpTO2nPLSRV+fC9YVt1uoxVs
0jhvNIvttJ0/LX9UTTHdVH+7ThvFZDV9UEe8TpJZUomN5ouWkX9CW+HR3OkNFrYTw+R7v1fDLw8k
WMapjSO58VvVI6IXz7OkbVK6zYYV0QOg7hBxokNfBzJIHFOMXXdfv+6WDEZH/OeyxO8QItPW/O4v
xZ4kYBIzijUXW1c9y05jTAeDB9hkGNrEh8tPKrlZQAhRHEexigfOzj1d5cACv86f61Fi68zMA+dg
snCR/0FSFSqd5YDbhquYTkybMxNt4O7HnNmVLJMrJKz9t2t+zRbV6rqQEoSzwQifhWdhjUK6wPJQ
uaOGtp6tViQ0UbJQ5W+KQlkZRiEKK3n+3HZbpUEt2uIKH4L/guXZ0wQ0GLE9LjuDFxDv/m/vK0wN
B+4KAvIsylHZAKN5ChF3Igjje5jSqRryBEetOZgFSIfsdORKtcQB+FcAW7TRaD8M4VO5Ufa9kEYF
mlLVTwAiKye41wXSnobCcbEGTFj/7+jiQqInlI4QGn7+TQf9CTiiYOvW/+clPt9xXXOm+TC1j4/k
9O4jUQKuPnBAqw9oelkHCxrTR8Cjts9GOe4RdNfEly5CnkBUMh+5AAwUijsSZ9SqNpiwrQnsAWig
e8lOelUtXLtzTFuTyeN6Tf0aI8IXCw5WPUAIOhz22+kGoWVg/buUdxs83UDc56A2civoiq1xh67b
ZZmj4iC1GtZdwysKGDVClsVaFIIA2ehwU+Bz/HZeu5rHFiA8YvJyVhyFUE5EnURIYCSmYmYIKqoT
rt0Mo4bQ6N020IqktGOMSxJnUkbVEXhE8GyN8JLq3z49AYxy1WPi4UtVgyxvP9/f7zhTiG59lT9H
XI6+DAPQxhs3dtZt4jF7lNMQqy5+WWCparAV7bqeXAi5DdLoOR/dWMaVfkiDX6CjaYSFvAlPwsIR
acKO5q+D4AMn+x/zYpIv9isc+D/824MaA8IviQ/Kfm0EC6f8RpFnmJriXnMKpnzk+yetN+MJouzH
FwQBVf3zX8ASa2wqN4Y3TcS2zTGZ3Taqpm72cnAx/G8pV1kHE/azFCrO+ubx5hAzCEn1CjsuORX3
vE4rIEUMU5snsO/SYcpxdAIoutDTDxjFOg4po/BJXUa2JjewOQeQ4UHGok1Nuhh2kzE5/7zu5UgK
JA8zaig85czqVCVl+2sGUNfygWXYtivLFxT+RfiDh1Nd+iVrIWtWAVuP/L23lrbGtofYo1f9neDg
bes/eKK73zRsz/aJsIiVE7SKKhWfgrPXnk5cAM3Es/fc92fNE2qm86dORV3DAGU2Zz3xu53DgLBL
BmbCfjt1A0vZXWEthVXq+DGiX5IS8YPCM73ksiUdJSRmy95pcWAuCfLHoUu9Wt2VqYv6/gqPewR/
3Cf+IPJMcYS2uJnpYamTOmHiB7ERHx+xaDSMoWQ4hwq6qacxRY0ca5meTQ1fC0QA5YTjUPBSLuzi
OPFYvmM75yk3mKBoe4UOQ6hraVm8bbES5W8JUv2wKV/qVI2HTQHUB1KXuUfzsc9JLfEkr1nMy8ZM
E5vaEQ7TxwFxFOWJ5THh4xk9r8yMU9AbeA/0VG1ASVqjfEaNNFV42dDt3F7x7zU8ZQtEIyCCVF6w
oxB+Axr0pJy5jus2s1oJUgyvv5f6Kr2sO/aL0MZgDQPqlYq4LQ9r4Rzh0JMog5FP2zSRqIEUmoAw
HS7TnYUn2wGAnTu7Hdx41EuAG8mME6IbqcB37bxBNnABD0D2zjLXidmltiQykwZQxLIOUEkmnZxf
uvb/NiAAoivFKsNUEb0CeL+FIClSNxC+xk099G9h7uqlXnU4EHabkZENlJIBSaDkkWJYqYpeBTND
wNCg87VWx+FV9yv7MGTBzho+OEz6B32Nbt4lR5GLBdi5KfKj94I9mN2II23cKfhCEg7kjEp7vC5+
T6UGt2wdOHlbXnLaxgLbMDiWpgqd+xNLiyMVJh4SD1YDjDT0JzVQ63Ap361lfX8yQAm4XsVUg+Nr
mLOu1JoRM3x2T9QFGXqkQ74P9H0M+kiRrgbaWgKe6KA878cjZsnFOfozqhHD8K7kh9pxCVmCi0dj
8Il4rCp5Ep5MF623vq5O4cUeLyejqcfjK0hlZWWjBEYzcqbkH86V8kDO3+MvEsgRfpU22dhHm9mK
Wn5zxarkI4pfAwO3B/gTiiGm5rqXnGijqrutJnduCKaaWiW0pycO5mnuRKUnhCVbZzL0E7+UcG7z
qIjOhd5s51mu4h0TOI+TxBX0vLTA5afvDj09Ln3cZcy+TVIwjhadVpVG+nZSCDMHEZdUNgokVpIN
20nIfKvRJghHfiG7IaFS2YB5sPXzHnmHSLnBto0SN7TrgQRRXVxYktCQvbkYxa8VaHRWPJ5Qt4n+
SvQY3LWopQPL0cA2joL4ikyC+XM3u9by4t85uGstAGNaE7rNmhKs6Y6iz1UEPyTNZRvC/vjlfGOF
CAnL63wggZt9o8wAvJ2vs50nbTcmp/KYnWijvCAP9wRtw0l6SzPTX+BwedkqPp2hLjt8ng6Asrk1
OBoRXlowzuL1EY5zM6x+JiSANvPJJjx/QvVoHSf3QsGkEUdCXR2hsYdG6gsA8uT+CZtmSOkJ98wy
vY9uILpzY4ayd1Uq6tw4v0YFDcjSOq/+tJMY7vR8u1v7x8lxgneNWv1e9xcECNzz1+UWKINsxk3D
W3JjHR1/3EFjn1VNdAQ6yszJaJdfQOTTdzjq4tBskH9n+XPXhYGyrQxJJnMH8a63+2TNwEAYaneM
gkTFiPOfx8P9FwJ5ehLg+seWipHeWdEgQtezSFscQUrgA/s1czze91Z/zxgGYjXkQSA1xUnC1oFz
Ms5f06Zq1gVu4nHf44bqhpibtJM2hlmUOcwYSEdqKcibj0/11ZSRqjoZuGJQSXeDw0oV7vb81Bhp
gvC4V2MS7Y7Ka3TRLLx4wXOLrn/qrAwvdw55XzBqX1bgfSr0nSVGAuVJPA66hZlfmoXbvJ8uYiSa
FJ9luJS8vxdqoU/EVoFHydp7/vOwYmnWLNcypOvcCiytrmbDNhwH8W7dvX5s6hW2E/ZI44WJb4TS
Gl62Q1cV3ExZINhE3p3Sakq88HnwSEjYP3mrJXJ/dp2hm67f1AzuovhE5sVmXeOaoJThMdGTQfqy
USo6IkT4uuGbfHmloTRUqQyFcmfXhFJTNGyt3KJK5TJomjsfpURD4P49rAhpjq0RJSP5rxgivS+j
jxEwgg4BewTE++wcQnSYt6Zw15iu0s7bwLYMD9xHwuNaHc6ya2yCdhhdkQM7Fxy5x2GVVRS82ZvG
XYJZBW3P8mA9xOS22wOpdCM8qPsN5a79sjLbGNu+QdOwLMIdc+mOjdcnJbjG5hBoouazRJSoPNnt
YRZrZaT4V3KA1uCulXx9BVtimHNvMcWzP4A1rucWPVKXb9SBeUMo1iCXV114KOOxKn+b1guMrZs5
BkH7MgRVEvH9FSgYgxO1wGxpf3M8f2kakqnRopCdY01CNQj+68lxPVarHu+D9lvSrStlhgrYfYh9
FerNuXS5iq3wxuF9h3XbSaOQMp89gY2ol6s0PvuS6Sb5HmI0EWZP/421tnPOUZRNlhTgjxd91ORC
aF8uBo/SH7MEGiQ4aOSneOctyXAUWLioIhL8QZjgk9v8FvsUxgoaBxPmJ+X9mOSxyQ+M4ee+HrTu
lkjPE0j6Djkqw3sUs7tUd9hMMoow1lSepiivz2JEG3pB/wirysrWru2JHh7tdAPHbt7OqyM32QQt
uREkb7ii3U6J6UlTCG21Fsq7Rl88I6mUoBVbS3OIxC3kPAtEA7BP/2V22v8ewXZnODPxihq+ke8D
F4is2TOXXcEYSBKRFn3gug0L2qb+8UKMUb4oOPRwIwXqTOkH7vXjRt5sYFvom5PrgdFHcS1QugmD
9S/Cd2e8M9olbGF8b/dIHEafAya+12XrBxAQcY4R8Gk1zQNwetSegIYejjKHYyjScHS9SkB6D1Hy
NFa3+AP6CVIeSX1Fsa5aGscx40bNZ2h1KD8BtIAiSx4tl2vQzujRX+N/G/sprIjmPF9qwJ3HGA2W
RDZnfukMqYKA9KhJWbHVn1VF2OPA8I+j4U2BASdIWeUuTws+AXTNVlnyt680mwrT1Fjs43BxQpTq
jEFk7ixJWAC/FQz7RLuT2yBAlnzIGDPaJ3AC3tckZFxl9H536gAiXKFdg+PEtKPUa8n6IQcvuknd
kD067OLSQUEQHZUUZf/mPZbi6lPg3bkLECJ8JO9H875YSbREDVOAdhnBKoZBV1Tb2rQpmAmQwg28
Zp87J9xjt7A7C8RNbfBOp3uw9GmMXPsgOqnqMWH94YqHWA9h5/Il+X4zwmBCruz7wvBC55kyCL0W
dOw63hVLClJMkzupRDUlu1xdRn3VbcGyHy4vAGUht6X+YUVQUf0fPVNpIbGMEF3JJcO291YqAda0
rx+5oqQQ7M2XQtxfTWdO5SHFj9TVRhZcUHUqT8+ZgkGF3Hwg1BMgnWRmlIw+R1JG8bGDwsD0uVOZ
+KpJXvrvLmDZm4ZnH4MwoA+XVyj+4wmxpWvagxlWbCkL3/erwRwINfxI3Bjj/fhucTgFHUL6z3GC
qqJ/DhfhFh4zLz4UnIJgFtXUxiipkLwlcNobyURByVgbcziTp3IQulRg+fdGDexSPamgaA/Z8/RZ
T4iCgqpI1/fA635MAwpwW0L+d14V7CK4+iQ2nh2x8k8VlPMI/IsaVS7Va5pLNeZdKB+FwiNQESWV
Z6oXICsL/pexY4NhknWv3aZFBXd6KH7fcOv0ubsOW0fObxJRkNcKknA5J/Rh4KYmGgAu4TwKRZGH
9n9j2oJoBECs1BjlEo99ezqvFuij1tz024cROTEEYwD7wFLtLceK9dpVpbaOGRSLIy8WIIkIf3lS
WfJ9QEOdI9sDvcwT8u7aY2x1C+Cz1XFBwd8+MON2HonfVTmF292ltLpblYD3RfWtg566qNpIqEva
N357o8Eg8o7uT3uSRwHosuh6nhttD4tWNLFbVymDPJm9ktFwcxqWp9QInOGRohcArmN9Rt/wMQbe
cAQlLKhaY1VeD4DTJjlxp8WjXAnczMTVDaFgQJEnHUG7OEkcj4ihrJxBLMd3tCMiDbxUNYjY6fH3
cZOduMW3KkmmCVh41Eg5xwlpDoo9myrJlptSiTC2lJVXOHd7AwXBxI/4hTcSSwiFJgRH7r8nhaUQ
RREdHnQC/Gj/0vhSuN3d89/y/YIlQS1YzQzO5EXV4Q95hgil0iAqXc46rCrySU2wuep/Gvq85By+
IzLuGre9Jr/vruIixrkhHSsJPDL7A5L45924oiZhzk7ZJgnANZ6DruQwkyu+VzJtCqlC4laO7uyY
EmWuxVcKMe99zPxq0q1M5Yn+uNMXtwwgGGM7BFov6TritEPvz+F3vVaKbChKn5fnEmeUlewdMUIO
UYAdINzpksOm73wOifKZgGpLYL+0z206XikpTH0KqFg60BXgrPag3iMw6gdFlwr/zV5ixUfHAjJr
ivFes88W1KZS/KaD37cHdgX1LAbj/t79dToy0PaRDGpALVrPoA14VCD9VJIs+zcF3n687vdvyCfc
ahoqgxXA0UOmMdRz/UFq7faMAJCZXwLt5o46YSHuNEdCnGdicOUPbH45ZWqp/1YtIfIcebThqTat
QqfRDE36caKSxqWcn4UL1MtZZDgeM7nbY0rGiacxnxHqK6F6QHdt/8NLq17oB/8Lxuvoide7e/B/
NzMjnoy6QJVJch98OJnrKApUemtseIohumKx5+H1uSNUsyrpj5IcHNDdiYqCHeq2uhY96hOmKdgG
i2HhsAA4jXJMjqL7lqaM9bw3DkFUdK/klGhEUTsN4rRIiKV2EopSL/yhU99/4XhWdyPczg9xXoY6
e1/lM7BxxqKbTCS8B7lPZwLoRJySvK33PkGFKZS+iIy2mV/bDcpgB3Wp4hOnxwENffxywZfiQtui
hS02b5DObdPjryOJJz0JWAQfto7CjzWVKn4y7p37l5v76av5fdqIhqEawGWgkdSmB1/LRPYHLeY2
wautZIF7VsU5AbdxHR0+b0GE+3sdpNeTMc5xCndaQqIvLltEKvAtZom0zzOBEe4UPbZp+Fwe1cLG
cestmJx0zoaVzkPIUt9k/ruZbrkaQoVbMqw4p+lk0S7/CCW/7sCKNgm7sn+Vz8ABB7giSKOyp1Q4
aFU1k6PKnRR9h3Ht6tIxzfsiu10wEykZqmvxi53FgGF7M0VdZ0VLAfCv9ldyBb6jCWb52vFebjnJ
yMFsghpJ1FptWWrkwwIugOLDFxBK1u5CPy+B7/Zvg5XDUehlu99sdzRc2azLikBDpxWwdOLtTSHp
5dvXCugz3DimmNo4PL74SAqEXkfX/FETCs4Yz2yvY3kyvA6HCaSzgO8re/VNQ8W5kWdcJdy4h7UY
vwd8rV3cB9oD1rCS85wQbyL9x8N27xxeYj2D09JWBlZ9yZjcUA1FxvtwLIY9eqGR08rM+QbiP0P2
iT9FdC+nmoIw5A240blQQacoZj5GOxV5b217KIy5whQOOD9wHMjnJJWpR6q7Bopu1+rb8CHPowt1
XUQ0I5mqeOoO5+jMJdrKcL7ozE31+KjzDPs+sovgrknCDO3/gjKz6Mw4N60oUrRIa/iEb9ZHcX3b
PwdrFYkHFTS60/suQuVmBcUhFIv4cAM6JP12CLikHYA6XaIs4/Hd/EvctD5WKwyO6C8BE9qJv6tL
AUBwrTvgFt+/ACPBcHgKdaVL+D03YQztuLPZI66xyZ6Hr3EoQoFCaITvq1zIHMSxDrakziPM4jaG
WYExyoZ3JcurqsfDySkw/NtlPEXfnkLaN6cmESDT4WA0CPlAD2vqeJYKVsKjtZKcN0MbKGlY4vnc
BIP1NTjb36pimTBVk5LvWZG7wZzkul6GW+Nu/aAs2Za4H9YYzxzB9+2kX/cGT2hRqEz97J3aVbUs
eBmJ0tcUy+sJMKbm1azFh6oA3i1jXB31N9dzVT8Icb9Qwzh9bg3FtKgd+bLAsRMX6DG51Cwfjz+f
96lkrBya/YuAmuhEz/CUbSbvWemHd0f7LKQglwwFzgf9VWESwFUIMovN+2VN57M0AY4wgB+Jm1vv
iyNsWL98tplZTRgbXG5GBGF+7ciVkhWxbhq8yB97SqYm1YIEsx6AHtue16uqmzbXquWXw8RmGQy6
o2yIqdHuf772pUTkd4y+RBAl5XfXpVq9DaqmH+OkyqkwpA7JKVccG3wn5mctO1b8S22q1Teh8+Uj
rqsQNyJdECcyxtl8B91B/qlZ2aLNOT7q8iZZcEz0gLwCgvjaydrpc79gi5lhpr//9RVA0OL3GzDs
pXmB0ngR7fg5PsF3+xE3+XWZUxkwrw+3fRt1J/avHQ4KXY1u9BsH7K68dKvHUwrzbpBDlw2dz6P2
cTX0Hv89SP6gwKd3ZGKR5DxtuegpEpcBMduy1I+hJfKTnBF8f9qtslUu7ZIlxfaSRNnQf1kZwOZI
pPKlSs+ozed6Efc/2rf9oKgPV7d/RrQaTX/0xzKM7RvHxvL80jlrMuAKv56Jk09Wb7j5yZ6zYrlm
j+FDDkaQxBgFbpiWu4TB19NQtFxM1EGuWXrAeT86kcnBrkL4OhsIMox5cBhdAIyacaHXY343QZfa
UUkyFescx7VqxOb62ADJttDgMpppkc8GCvgFSGVdl0B8dXevBS2HYz8/YnEpWMIcIWnmLBTBtegd
LL6lF4ydozfx6+q1hRodjgxAXPg5MhQ6xfIN9BWpPTbGCWqzrVhkgZo+f/pUAcDgfyrkSmmnsQ9D
vdGB8fjPhQQneKEXP1ZRqHqxu7nUuzqRkq3JUz23Enoxx38NlO97hvwPooMaV9VdWMNLO+eQ8FnM
ojGOHQ8k3DED1jNCedoyrV0pUzgcZ/heMOOuTmCE1GkjXvWWO/8NF4zwIE50fMHukEnzjy9BKTS/
03VvPnhMtrfUgx2MHYTfPwz0gzLweCvfmRFx5KlnvuUfb2HlNVL290sb2sTa9Ong7fCnq8tHdot7
Yy8Xv9soG4t3gOY3JvgBiKGFWDDijgMZZSxeeGiZXuip74RpANgFZu/+ICAZ7NTE0R7YEthztcmW
5WsZrH5jJeMw9Dp40oUumWJPmEjDOXbPWWkJ0CKQwNnpi0YYBHeS+nHxB2Chu7kIIGyc5P73XZ1/
j15v3AoLvXCi22I6tcPNuEvPpjhgdhGFfsTPoTPiqgWpuU90ZfwkB4Xalu+oFX9eap2RBSRGqUna
E6qsdg9fjiLP9BpfkLOf4fPQuAjP5J+jUURHKMobXRNOYNVOxXpcvOqRu2oKzXe6cDkx73UZRiGN
gqzyQ++ZR5E1YCc1/GTuB/H/MArse9CBb3/zVSoMEYoKiFIi5tKNSPMj5MiSLivPxw72rqPayR19
rD2ogt7/QPzDAMsYuGL3rj1tplNWym9NNPdTSDsNrzdOB+7RcM7e45Er4ASSN7PYIiV3uiTSUpPm
4273jLNWYIRhVqXw74X3XwTDd2M2mKAbHXhyKB7rcWzLjMFXBHu1GHdhGdgv3AGzlSXVgMArpUn9
WfvZ3CfDOY8AthKLAixzSziclavjzP9vHkk1dlyY1xTHG2KGt1lzPRUp4sIlam40RPL5qXrgLkfg
UpXdbOUJqvK+Y5VO5b2J+oHxbgNXRV/KkatkNK6VIipGJvAiWJmLLk+o9+ixNU/72OtmclC5MlgE
FRPWckdMwV5KIwLZpQ6yFs+qxYs5jOQfovSCR5Vr80CGnwpzuN9FpxvBWr/2KuED3CujkJVMyyWR
+nRSWy3ayq/BHhIy+KmvoI2QsRngSTio3sPIJyAquhIhpUaTWNwTweBj0+L3ef/F9d4fSYMs/atw
LMGzLidkOexe1cKi/bvhbWpcE4h5OEt7WZBXL3wROBmPC+BJyobN7WweVb9IE3G3AmpoHJwxEJ9C
HQ0jW7StqByEg7Ud9ZoSJY5LEtDTuZfx8Jt+SNRAc2pDVlhByvyDlgGs3d6ngOt9wGyqswNvbjt/
DhGLr/JiLb3/+PqFiZYc+NjqJZcefm1b5er3yUKmQgGJ5L/sGLwgX2vIigw1n2btXA3fKPmDwF2f
S3nF418v73caXxCzRTJRBVYvZtHcVWw9sHG6e3NfxkP6lJ8pe333yBSswwYRgcpDharFIKYKwoXR
jK6NoDh0I/9+FtQnAmTQk7PSNov/YgP0cujqzURlf12zS655YHqdBEV+hPYglcUkLSpvHzhx5HKa
yja9w3lcFcn9vLCKGUCtOWQpSbO4oFxZU6oN5qFQ5rNqocnOBt5qNucsl089DrSmkBwH7x84fYP3
v1hDd4I3EX+IXgll04kFpC5WkZ+7DSc2dKOYU/TL6CK6JlVEn0PSKqPD46wXF3NswgR0q35SdHfU
MBynQKXDwYijzm5lDDa/JIOBbQDEJv9xqTblZIlhWjFeiGYaKBXUKhqkCozaKEPXM58BzP3i6gmJ
nppKAl9kK7PhZlogTTvqaXi16RovdZYri8kVwosPT1PptiS0wL1hKlEEpqkWqRaejSMLYfivtmrT
A5QDZ03gf5ke8+iayKAUxTFHldNO7KMR1BICrfSlCAtKJiuS4xUumPnLxu/IBfjiegLaRxz70h/Q
MtbAh9pu6qyB9Oi97RZgW3Zh25XNjafYtuczfATABrI8pIC6cCJ+HWMA5LDDL9gSijbt0ZGB1Hs7
Jgxs8jhSHWimN9i5/vOOAhMTPB8yh1nA0qsmvrEhXLBcRT7rgictOTjhvXEiOvcSFXlu3f6ihl55
eXJsGiqA3OUTVErXmM7FSYVIVFfRC2iy6SO5KDZRrhRRed6SOfVs1qaP9WKXWLhwraLLAdsOwA2b
oOaGFwSojRiKNeJdk9xUaBtzEAjqnPQ+gufC/KlYFV+MMRi6X63oOSVtyAdLuBNqBI6L+GIau+3o
pHAZJQpDcoVKB5RKlfv4HibnNTvMQ+UZJL1gXgiWza6EnG0thvvYTnD5tvRRy9QORH1QTQ3vmJnX
4FALXC451z07odzyGdFVn/Zb7NyF+RUvCpyGBxbQLXx6f82mj3H1d4q6IZp2i9YetEpqfHwDsWPl
XKGyaXXiPm3g5BzvzkXEo8xvzS2jhIbZf6RepkZIVcJK3ZxAWaabs+vmdu5UHnI/fTKVq+5u30sJ
mQybgye0vwkZF1xLyhMvgZ/zi4E4XLbH/KaCYe535SHrnmuqQLVs+4i6fZ0OlukdHd/dDiyR8EW5
MIf2/sKhFt/4v0EWyLFd22uJf3hwXZt5u/JsdYBP5teknE0km6GWepk/ZDIjAVBupnkcaJdEh/bj
HFGeo5WhnC2M36vlGXGWWaWccJKqCmuGtWGFS8PdnfMjk2eWWfodo2V9C1WXjM+DYifjPKFUTTaj
1wKSWGzOFwZmHj+az+6EA2hOVX12F0aTnKMMoY5od9K/FGDvdVRcZLg0b8eK+CfoLjdHqegZYLhX
zKbLpGp1TEMdw2oqRzWwATCyO+v86qLLAPvXpWCEU5kBJ3kI3OQAJqRzYt+T7Y3SlGaVud2AYlHB
wfPIdAYEBcCI7oX9DcG914J1ErXI6EJG4UM8c3JBtZdTFvod0RrZ8lNFK/81qiYmDwMJk2+l/vpn
luTHUSNu004Y0UtzxHS8qZJx0Vj2GmowlLIOL1kp8914P6cQQNVCuW2Pz9RfGijqpAXf/NtQL6Qa
DuyZL5wQDNdPEN1/su7UiC1n8ruqZHRVVAEvXYXMamLmAvloqUwQpVUyTqZMUeuBN4yiiqaTGzX2
iHyBQg4yTgci9FmKkcNsNd46VZyjdY6Nyp06HWLLFgGM6GqVGAmXaKN7qH+VTxsqEBZD4fB3n9Gm
o6HA8e/y69q0wDNfI3a6rp2JwR2OOLfG6vKIpxs+6SCGcpkUTbsRpGEPocIFexgdBB/Tnb3QZNah
RhCAzGKszs5r6HfiVi/UoJBId38quf7jPf7HQoh5868vGHmPx0uvRzzhsNpubPs1CjgWBEu5Xx1Q
VX6Wbd8+RNuCan4FY7k7hpFnuWp7VfT7BcYf4EW+ne63S1GAdSb2lFkFTUyjb7fZNRaFtJCOhHvp
nybAhH89q0WwlYMCOWiUeoodl03EIl7fPKa14uqO+1FHr+f6AXQ6lRbJ2kmHl2hy11UvNSVJBiDJ
+SDIYJR9HRbriiNzpSQj+XQ404tHnRzbfwDS/+VWiF+ZnoESGEsQsYqEiNFk3N63AEo8xHpBI/ZH
whqtbuftQTF/r4yeWf7tU3jumyqfiPKYkcO4Jm8aYlJEzTPgOCmCryqN8OQzluAkWJX8zRRLUqm/
cb06CSqlLzHIbUz2M58JS+6h0Nd2uEdTNGPiDxe1XqLuCJ4uRI2IumGuTOHoYWpUlv5IpdgyztfS
px/l3vEQIX3T0yVAx2U7lJWBVgOA6oGUdu0AlMgE/Ov7hCJH7js4KBHLyzKI60VxKk+OGAZS4ttY
uCMqMQUVYg4RVbOC5dBNKQwfuhQd18FKYyFiPae5ZrNFJZy/ZBs9KEd1c3LIvyk1CTXn8YEKgRWS
y6Jlw1UoJ0kmhOT4+8tnAJSrC57j5zXQR4K3cLKIuccdYYCY8zSgG2sSTdAqk6qF1DvVmpIbMLSC
IIgM1nF/0xP8pFLH7DAxBCG0v3MOTLX+NC3aOuUE3qBhMVtQTBn7a5gR2CVQYYIffxA0O53vt6uN
Gxt/XMVGx++boI2KqzCugclM5zSvazMTjaLVVKfCGyWzCG0JFVeJKDVbji6uFBHe+ln6KMzeZSHo
w91afMrmsz4GA/HOqeRzwy8dO7WuPxtW7mP7LLOKSr1X2d7y9kvxORt2/YWSgZixpS4zrQdglzBn
+K4Ge18tUoegwUqRJYqrcbV1mbVoh0QCNXOVnl5YAY8PTiODQoCQx2preIuwnWF3bKK1M2xNkPyM
bM4ZS6uWzp2LD6SNZHy0GTcdR5SxMlKtiKOm7jPOVVx1xhcZ3ooiaorTuCck42VbOnNv/HED/M9m
j3mVEruutYD6pLAXeB7sUpDXye3m/4s1X52PEcZ6ZdDRdBzLusKrxvS2vlHXN5vDtGQ8XBnrgOVK
9LSTza7KopGBbscUHzMPJd66PnZKr4wo/ak2jePMvepSBMfT6GlE6ZQWEYyEUwr4dOlI4aca1KYc
jcFhYQxVI7Dx2SuwJq9cOUB7vaYrnXKjOytX2Lhym3logW2QE6k2yZWVqb5fRW55hCJhxHkOMf9h
/E3NsTUbJUxYyxn+hMdAagLiiozrpxbBhKPE6l9pvrVkMWpr4D64sMPvyXTnZpWTN5mCc8Yd55L4
fJ2EomPkp2vYSAplkJaXsu/5j3kzUhO0IRP1zJ6QF3FHy9oYblwUsUq8SmLSd7ZgBU0KwEciS9yX
LKwDYCzpVYaMznXPqMpXr7C+KZw2DxetAH8IJh+nxpgreeFl9UyGSbbCGyLWIH4JA/RvtcPIO/Mb
Tw4hw8oGuBrUmnUFLOVzS/WLAeUkKS6OVFNNe/+5pFQusShjDDDNR4TFAGVzGiH+p/wY1yOvpvEK
K0pLLNHrwuOyds/NROlt0/w9O6sY6quG7XUPlFFUUqdYvZ3s0rkSzbU63AXQq99ooXyqBnjnbyq4
33DE9Edk2Kn6zYPDGkSMn/wp6Zk1VZt+MbVtxd2jUOfV+EMOcjZhGAWQxP423HLBLGhjYen++LKf
vdDQ63DQJNvAogCua1XOogC+FZZXzv7E/3VfGUunFulODaD6c8m+cbAA4qRIkYlDnf9YjvCqW856
9haOTNkgg7w1gLhNZUY42tQnJvNXEqiDO60HXm5c+a8EHgtOpPdj2RtpXj2tpC7+n2GE46eyYAqS
1Zr2D5gL6uNt/PHPldk/lXz/KE55sCGTI/3NMs/+9l3IdbfdLXQ/WW0vXnVZhV1OR9GBugzECIxm
eGc37ar5+j0x8Am8JE/8qwvyHO1yd3Hll+OCZLcXOSImFFiWJyFYScTa46lRWXpT1p8n9XqmkBWO
Thte+AWsCvXztj28zIGMNfKtOJqMkgf5ENqN05M1wgjyvsT/qFFnlCLKZPEtRffv9QJCgWbabYEz
lH1zBnHK4kUfY8ROovK2DBb2aFLkAaWxar53PhidTB3/MHSCF8w2iGvcNCfERnNEjtaJKGP+TVMg
S3efQNyCohQmIR/2PWsEkpagDuzNoGIZ51cMsLkD+T908bUXonDTVI+uIMPfoY/ACJu47dyWhDHx
zRyUFARXoa74TAeIYrByJYzWLGW3UDsZ5458lrJuy8/UBkMAV2bIbn6M4Zd0FUe61HxsqgLomUxd
+AqINQHxqzrfhNdQaG09cObW/Pl1nQUqA2pS2V7Bxfozt4uWidxeFYHhpgrO1QtmNx8E884kP3oY
9oVkmR3D8rQ4f2edpVHTGf9CVL55Cye0MgpME4AfM5cxJ+6q6T5sKHWoKlaQRNDXoTE+x6qe9slI
vUIb0FCGOimFdwgr3PVVUKA+S0dOqor2lcubLQx5OVvZ1ZUFXy9sPI0RHftKjq4gKH+4lj6TCqWK
yHTk8RpIbJjLrsfCPH0kDb1FPTuPln5jdZQOO2vXGKpSKF+Xy7+PN5bWUoJudNT0j0lRr7pUkB6M
2lsvIsMjyTW7eFuBROtYFBdYnmjxC/o0ZNAw7j6EDsgRyw4PG1KohdmL/ntsAp3JWyTcNxz/2Qog
rRack5pjzkqG2sYKYS/kM28laP3+6KNABCE4j4cHvLIMNBOez52Y3OcYfo4Ajs7TQvczQNj627oV
JaPNq1NK0ASl6zyqDGuCQgZOJkAmu1aSHhHKyYkElPZB7aRRZKsXz1NGXXNe7Tn3H5i3/myJ94X/
p/vrI1hmpELNSdpdAYVDZHsDjV/WSoRJTHLrVr+2m/KLGTnj0OJHaXkE0SaFAaxnUyTQtT+U0nBW
c2IivMm4BJFSBQZMJaMstc7eqpmBDisVnj3SUgg4V21kORE+Qg1pH4IBDw84f/QmR9PqrXW1/sQX
bVMF3dLDJ0DytrlYoSQCXUtDTNYz2Rb3D+eDnKRg7im9G7sW7UYAnuCjJk05sKz/spHn+86yhT3E
2fOOzhh+hqtNb6JoluN8Ystt81w4gpvqqDyfMINNQvYlFSFrgFsGIB3K4xIw/KEZidTzpN7y1oV3
XVJh+h4KNPcbIcwFJ8qaSNGLP0RK0sZyYorgYT1VEPBk6JDd1mE0g0zmQTBN7MwWEaOEvp+iNtkK
5ltFyCWQFAX7DUN2yJMiYwrUqfOuEHN96G4V7qObL/YuVIkEoxkT7ei1JOokxt9LRvj/6ofUbLHo
4AzxzU+peGgz86lG8MWduzMkb4GBaX7P2lbdTY5sTjReFQybe0SHNXGxV776B/1+r8Y/quAc5if4
96GF+ARLVfOOi6QSOvMDQvbAW6RCtyjGNda2An7tmYOcgRdSZ0DznEVj4dGoWUkobUEfhzATeiqg
3SbylFG1Hjy4kjh3xDkNDFmRklF/FHHuKuM8AiILpSNrXkkcDhb/fJmxbzcocMWV8JwGYiuK8NTX
cnv9BdydkK3elPTfniWB5DGeI8erynurm0bixu1Fp/S05QkL7k27SYOlB1JcxifHdrw1y0aoD85o
rfTZqVwMim4Se2CDs7H3PdjR0DILzkJOkusTP3xvKoMhWDCLlfMTl9O5W1X0lEd1+puDVZOvTkA6
k1FVVRjYV0mYrZd8nY1VrMiHOA9GtiBrGp5aZopbXYVpGpjezI/EoGviSEHzKl+hnwQjUPbTb4i1
C5EYNpMSEjHNzVgBvkzzLswtapdCvFkWrXDaR+S36iTSJw7G3PCJVYJNBQ3bM09U+b87iU6YN42R
QpkJZe28dv8oymlKNh65nLEj5pE+fPpvvaQX4z6SyGTly8MXh8gD6BirLiSFGvzb6XfOSxYrcleT
8r9+l6/U9nIfWERRW+rWHXYFaySuJFTZI9NvyKdBDGhU3FtRXqNsZXbw/xxzPMZVXV/QmIyaQ8sd
HVoH3v4GcYLRh0Wxg91vAgu+SdgtHGYC04JHTvqscYGo18PFIGAC9QpSvgWEJtSYHTcNXr7D7n5u
dozHxf97Sa+4WYH2dPJDRbcXZgNwg0k4H5r1T2QV5g7a3kfWdanQNtZUpftNGCRjZqBNmh9Gq0TL
FzzDJCwr24Mb+tQP9pqe8VKKS8hU0OLgyAy/voiU6hzjHJISGZW8N8p3Fefl+BVrsZgzoHNZ+1oJ
SA8h0vBqt8ThnO6vg4zMEkQNHlobZUNCgU8eqIlRMbICKODBdA418lQJgLDNLY14Fz0dBqGDRNj8
t8vFQgQUA8o0VBHkqdnfx6LrgzOrG/3b44kMSd6Ur/5F89sqgCXwwfXC9kJuBhOuN3g5gb4rmp22
4SUmmLfl1nptKJr5FQxZAtNe8+LGV/g8XD31YwTA0dxgyp/BgtqfuOrTCA+QQYbof9TUVk68A+mZ
zetuF1O6f5SARdHnIcXKNP8F0vzs9Ik6/HmEqIQL9kDUngmyR8LfQHy23NWowh4bR88eh3UNRxH1
w6PsnPOejUBJ9gFOQ2Qm7MZAtCVt/GUrYpZW11rDdBuYjCyEUOUaXgzbL5H7fsnpHpWQX4x6oCcE
XwVE6SlTO/dHACzgjIxoLuIMF1q49Q2yMRB51pWXslhkPQ5gQeNA5N+w39DYgNAGo7v6KdgbLuQo
RdIG1vszpcCSPf9n3Vipa8FeCrM7tAw3DlKgeAemN0PqQ+BC9B9jW2kdjESkf3+zndavDhDXpI2w
lkoZ4QIy1dWXT0wgDC1EdwNMf9HXtC4pqApNVgcwxXEncPw/XhU073EkH1N67cYoeraFii8O2O5p
Bp0ISWjqXAV6gvOzBXLbc+AC/BqaOSH1XMvU1ETG1o0Z+rQ4IAoAUyl2lNqQqTFeHRIaBZlNTUyJ
T7pOV3t56eSk5mz3Sej7yib1SPcAcQ1MJwzBaVN0UDGknMJsf6SvfhDRAXzdXvntLNO7lsvEwN63
YlhXtNzCI/zVkBGvxLYdPngsWo+4GbLnwvJY/vVqneOPkQYtzBzl+uQMvEe3uU2+mAsh28DXzEzE
yEIM8adJ00xPd2YNnaJT/0MbQhBssEsbD4dIDXv1vwZBpmBWTFOPpEJ7GLcN5HJmqR0eUATsDvLt
B+fLknzWAhiyXo4hk64CqjY2riDeFrwgvZz6KsAlFrTWyPJeyNVDGk9/sCf3B6k6nm+c9E5fPyyH
zcWXRKmiSFP/xQbFd8BJuFUc7fk64x6EnE+O/8L7EIXuhmPsFZ5aFBcK7s7INgbCg69oG80PGMwV
TR5W+ZxmbBcw3I9lEFXvWEfnXG0z5L+zMCfoHIXkbvm9Dmogj2vdbkl/Jb5dI+cKL+S//LDvJ/Cc
uJSFJeLaQ5BsFQIB6w+/QKrH65ewYPCnwvA8CRLfmswsHs1RJkr7hfz5Wr7LKYImL3UWt75ip+MT
d2h4Y8//Y21rj8rwgMzixMwPOFzKzaG5J2ZF6ZgGWH/4pcMjhihHJ3GzmNqtE9/dVGrV8A6LLFR7
zWWM5tV+dloUWDUghrv3fTmX4+3c7nfIZX502xI69P+cyR74y19b/Ie2gH8EAboGRgYlBARRvj24
tbUEkhyYttGtLWSqRlOK/TdAK3g3KSSBDSzTNWFn849O6K2Ol4Jsfjov/KxpECQuvVqOVZuDQBZ0
10ci11ckRZQPuOhMxahs3XowOLvLfx6Ib1QcOI5qMMFC8U/dEX6l2I1MZAMlCbyS/D6WkzpOAhbF
8lKEvbfb8aTYA7oGDe5eEplK+tYjaeD5E7IxrdzCdnPyP0lEIsdUVwM+RzMVm1PN44Ey7EZRJe/U
s8hDGS5ZszU9wxFCLLmADAyhsPz69oDxAaTCT6lLj+syLZIZagdLNWkZJYmElCqxTZATNnhI9y/G
bAkhFbynWsnVZKvAxwTSX0vgLsRALLENZTcX9Ma7j6sO6qW6vjpl/sUk5WeSV3nS2ATGVwqauhAI
HS62Sz3wd81VPsP4sqlmyMOhB8lVLFVSv9JYW0Y6y3zUWwfjwpy6LgembLuv53cKRU1InNyG8Lor
vviocolJAkOO+shI4bw+reHYOUD/4wjBwIWdXfMBfCYRmHZ4giyxEjmCJcY41WSYuhxegCDnHrEQ
PFdu1AthU7p5Rc15DO7uX5MoyQgjfTUuC56v061XoGug4tDG3UevniQ9cem4PO5bi7JspPNu+13T
dzq/kY1/cLNYBoi9WA1dkqJFydJRBYrxKgxT9QqH9rA1NxWimU9OrDDPjINBVhHJ8457HNo7KRLj
LM+3BU7dvqAO9bgLiI3Dd+6ZWgXjuHxOgUYVGIFsdX0a+3WoX/fRLpWQH0HFBckutZFFC4KmaYkO
lA9wD7LLRSxepmdZmhtOQVYkMM7BLZEDkW7YTP1xL/qMLLjSkP89V3AWGgbOxR8t7KMcG2Db9srP
pFL8gPm88S/GGpc1Wrtob3+MlFNcw6AhRCovTd7AN2gdoAWyuyNymfvkW47BHco+uLXQYjpYLIjT
CgWAWkHpsc8Jl0xVTO08QTlvqszLxvtuhimDwgvEIL7pOHknmpwSQ3KC1owiw/Zhatw9e7J3Urnm
6KQQnK4hhzbBPf6NArz7AuNjom+c0LPKUZifd0/2RuXfcVytVVFgbbhYqUZvAiF+T7b1mki8wtrE
a2TeK7GtbJJB1cdZPMHbBeWRAsCG3q+X4Sen3Df8UIu3b/lGHHhH2GSU9uyh9IjMabxl0ZJUcHQk
Qo/MpyAE/vUYGlZgcCF7fDsPfjxqbcWs6SsruT8/zl2GHJ4u7SDbIAlVeErXKtot7tSRxcbmt+q8
eX6dUqxHPn/oW4/4FNwKOOmdRVIxI3nNUu4h8LUyebydcpsKdw1V7VjaWA/OVH9PWJsvk7SD9nVR
+jdH1gj0Emlf2AXROHbs6nUh6KsHPuoWriCVai2/e/2Ai+/GrZx63g5WhG43PmLxHHsidgw6zphT
jdLoys+CtMbiUTiyCh56vd3ZtDKFKhIOP0SkFRetIa+q0wAszCykeH7XiZ0PRyhidUo3t6qNvuaS
Xc8i5sIdlrJpXvDQHCB1l9lygtFM5aJFK7kv7FPt+oyYSAllrCnHX40G2QteIcXZAewLTJzUuSjE
zv28mKBVVwjsk/kTBTiAqqM/xFKOwa2AD4SaMnnH2KjR22QMTqDutTnGgZYsrznV9N79e6vDa0XZ
lNjfnwi5abMLHJL4TMwzYC+hOUzphWnvuEVCe3e1fEtVcLXqbrNUlLlo8U2SR0t8zJqfV19MBK02
FIQZpr4fKcBG6u6EWu7DEWJdXM8Fz3B76jCQxkAr9RSxribQpvXPtAcQKM15NeytXPFB7VJnPGtp
19AwHYT3ENfZhYcbwMrtPyYFU8g7zvnCNBVo07UXDgtPok3gYooA4SGdrNdXllL2x2UzoioUnsPj
lRFBsIIDRkZ9A5Ae+bCuWGxDbxSw4pXixbbf46IdKCGZNu1hiC1C++ocasWIuW31Y5TltephdDNn
OW1h1tfopTBC5rKw62WIt5CVR9qazDGCravxxdgFzIQVzpv3XNNTXWy8h/DwOZyCykolJohLSQ3B
vf/wq0tZ0nD1mn0MShSAomn2fo3uyycv8yfxOurmO4cbY+I/oduDzdUJbBjRpgLeB43RBE2bzSO/
sF75ixxy/yFVo6h/BbJ7vaYTiCOadXU14fZDTA7wqw0hbyQ1vOzCsZxu4VaDHoc5lyRrBgMJg4Kl
oyTWl/kSrbYuGciB+XzRK/wiqaEO+s+MCsYkS6wKsiPk3B6zR2FTrgIFwDtRUIyX2YbfyOk3u/a2
J3gCsnR40xMr6EzFH3VDVmhu2CTR57oP8YE6k1FqGHigJ8xOSSiSk9d+QGi3mBvMJQpvTMZGn68x
SOqaBBoYwm9ZFvVdpJvDBfGAn9F0v8JT9jOID6amSB6gP61WjmYUymG6JZlnhuTf8sJiHgdYI7Nw
SjgRo7MnmeO1thTgzeGQAv/bgqsr+tVecNqJ6nE96uTXySJG/BGB2PQ+XeJboD8IMaD4bcgXS0Ta
9ny10N+j5w9c0pFcXVihLXR5BUR0fkBK3rSqMKd/mAdZx5nsnDJf/2gEGvnhkS5h6urilJTzXDXF
DrQIJNi8TZHSfDENuNCvg5UgzrJgKdtpg0dkjKmQd8mfwlkPca94m/9FGq+fMIl5ynhXDAIhOyqy
sZn0U+PabgyOIO/7KdFFGVHZCreFGXx6AGtrAWnpahlYSGRGwXq1EvhvopBVy8BoZ0UEDUXaqhwV
U1o4U+mrtMhGpSZ0COROXGnNe85d+T80ceM8v/BsyC/lwV9gT0mJrDkAlbeIwLnz7/t7hiH1mIHR
K3ojW95/KNL+U36X3PeXaoiy8BMkbnamHFUqOIkHMHmcIsVehPbCmWkeoVgQstAv/4rnN1n/0hNL
jHofzBj9GQ7hJqlcoYNr3ygxyQ3zOVZJD1P7K966Ra1DyPLinaDNdPqF3Fzh7qm8D3aQhlfqrEjB
/oz7jZNRO8+mxGGyCYCegf1DMCYVvxhwBQG5en2hL4KuNMR4hCppqnC26JKohuQGrQJmUuVlphaZ
j2HKroKjoYYWyfBox4H7ANB/kZC8h/PhVapFfWf+wunC0dKDVd5IlMnWPMKd0mIdhpfjpyT4tEgQ
1iDombAxsZDNGqrqcdVugCfu4fRGRySLVA/Ef4492YzmLiAxaCdeZnK1gKQM+k4Gr2jw4fu8r5zL
4n/7JBZPDlCMBieTHCMrf6O5oDyHen1ePlKjaM8Rm/dSIoxg7Fh2zdSLXLdJxzZEkztjUSgvEL4g
iW37EQOsGYZmtom7nEknYilWjEB+jXOXr4oAXpr4NDQg2sGb7a4ZgH9H2WrWi/8wfRYxRQm87zG4
l6XG13PlRObokZfOwfTT/pcns7C8GKsGjl/Xq0NohEXqpSxSPlsIs0rmOWjyRaRNN1wcjdFjRJO3
CqCgF3d0Hi056mN/2MjlGVxpsBfLnmDG+442UETIyg8MzT6H+xnBfWLLkX3PvvyUgc0TG/HvLkkR
q/wiZpDEEoNQoMXGRS+kXKUtFE5BVXko/IH8VSi1f4c04dYZk0QNh6FCc1YJdG6WBsXz2vIGJfak
a8DUu+cUVwwlPgSRwJ9wK9gBurRaVg8ebUha1YVuMsy6H21odQ33cQKGIAv0IC3xihaP5BMWCKZZ
jh/in0ggmaS1v5UM9/jKIUPhtKmcLW16CWCouXcIklzuLZf2VhX9OvVWz4YbHwUA4L7IvWeOoQbf
AqXwMw6G2PfU8yXBNM1ZHMyB0QyC2bFo2gtg21a+9jHFMAQn/1zfCCWf9zy5j64609QIK4cKbTem
2RH9TOtBCK5/mbduwTrDSUMdn0WMR2X47FYAs1O2Oiq8YYqA7sJ4VwVObt/8ccLjXUqYPu1VybpS
vCps6wcn4T74D8sW2rJrzIDc0aHY/+1IoKu0RKom3kBQp/Q31Eji5oM+wV9J/wiCF6jOEjVoZXYG
4JJ/t22tHEO3R2v+fpDB2bPgVZ4B8U+nO960P+D/5C0yA9ZlogBQN9fIeuJNNvTCwJkfq/A3yyCX
Xd3z6OF734fnu1c+ixuz2tLGndoKHMOIQaYtEf6YTLYgUHcVCgDtn7o8FiOKZ/Cf0OF8g5OvK095
nXyzz46YFi6xaFyH/nT45kSg2k4LR9c2Ilbwa4zFUNgqB2Ad0mShhRqXT8qbMzjHrUJxZVyOF6Qq
G4XHtsEUPt3LEap3Je/CpDsnCm8PM+HjvD+cfHtFmvckYzubGj8ijeM/vPXHZmSas+zxFJEeT/Xv
Wh0qnjLDwUxxaqwFJA3we37GA5EP1dkffNM+BIlDnQGB7btFAtbjth7dMLaJcRM8FktZOl2re2w7
hz8PcisNNqpLTcKPXKPrC3bKEYwe6IjcDheNanI0qgWADpm84GNQCr2thp29xluh/Ji0yAeL6wu4
4meKoZb4OTIdyp6l7CcGKfBe6Dc6yzKnf3OavvZR12K/1j9jWqkVi/SxCzfjJ/erfWsX2ZhenIQD
OYpyS0ubndPcqvZ/M9/WG7/f3CrADNvJ9TB68R3Vu/A7KUaIrQBlElpngFHv/0UmReolSp2WsGOa
FUy/NY4m4bhXP/v3ZGfd7ztxP+AdODoTaJklQGj08/msJ6hffOSr2JaNkJlSmqik4QvvrOw6QyBf
BduLnN7NSYm/VSI6/hElD5SQ4gLefc5fEEjh5rdg78QjKnKRIQSNMaT89Ikl2o+w2fGZFsARMfdo
XJCR5kYHeBgfSEAI1sfqUiLBRF5+St9zN0tsQTx3gpSEqsF7duxEVn+wbIeGzhIoxKDcuzLA8lls
6M/Z2kS5mj7o0lBEjUw6a/2EiDs8O2j/yFD9bxzgoUftj+XcSDJAojJPdnRbVQjUqWYPae0UC0fc
PPqUYcGJ26XIRiz3ga36S+VrmteC9o9fIyVZDtkrPUxNGhw77OohGR7Z0mIRFkCL+Lb9eR6KFYOZ
otfPB6iOT7r6LGSVn2ETdkLNCVX1yWLRf3tFeGlQleLpHrlAEtE3wqymdRTAAOwcs7QCpR+CucSa
DBiaXCztq3CapfCLQTe99h6Jy38oCSR/lHsQRwygdgtpTYfv0H+P73AEF7MljCF+IbUFNqQXzucR
LWawngTP7RsmatEbkl4FvMCNlbmxZMO+4QuBuMyHBswimtJRRE9Yjt3CP9viF6KsA2i3gYNbkPUa
RShvAtbMqwKrzi7zDr2GRb2g4FSN7XOnt13jRbMlx+8kKfviGshl2PwAxfsPQfkwbbQOy/KopZwF
Uc5HRLXNl+/7myoBI+g19YyioF9Fqd3156NK5OlsGcLXRJseLhbqfXJ8aIkBzO2BGNb94OP+/7WU
RPi/F8ovSRPw01VNDEAkISipLsUJ2KipRHp6zCJmZKi+N4Ug2n9LziZJ1q/5iBWeLRyzMrrVceod
a/OYCNldsNuKkZwZyvM609D9I1/G1EKOutumKAbmq/mcmMvPkwXT8UYtIMYkq6h0UTr4so3AYnuz
bFGpEllWa7lZMBnQZfBxxjgesoigo6wGLdoWvprGzV1e693MWKXfmOjAmH6uURz7oRzBWhg8vS5E
ILEdM9itFgtAyAWQ6M2+JjVCU2QlQXQYmqAACfSu2PdvWVtu0TeDWbqCGMYbuuS99sVTZ66sBEWL
FeUeb45j+kMiUBTqS571fskAPEu8GAkqZpZL+2Krv1X7UCxiKgYB7gVpMGvv9vv2Wxl4PdDbXgN1
i0sd7liCXUJnIxWpgUzihocfX+Fm8a9yjDxtNUSApL3szKajFOWoLwfm5hn8UXnEXpKma5LDV5dV
tdPke/nItJTX6k25JaBmDk7kqzsjLuJPJ1Cg4UquyB6pymvIQ+YzzQzUFp6hVS7KWeKvR4PuMm+b
4spKvrzD+k+UPLB6REYpIeAqrYXqtBbMSkgOcHPZ506LSoRSflp0TSuK7ClDFvkgSZWlEzDkDG0g
rKpq8jW1VeHryZ4EKRHaGuOPNvk9c90az4yQ5mJL7tI+uzbY7LCvN/0UDSf2GCoSZVbODfC8P5Bm
tB/7DRzod/mv5i5UzMStg7XkTPWfTR0a1YDHmZMMsKB2fhe/xT57yG791LPPlSFewJNGnOrfsh2e
+OyyM3Xj/GUxaT4hEmGXUfSB2dSDBKF5RDVriP0X6qXAd/KlZgaF5Jx65tnSlslunWxoXmhaiRKp
dsy+sC/fzzdhhU1pPC/3w5OkJ2I4Xydw8k7gnjW71R12tEk4POv8dG1SKQyAHn1Gb9GHEC5xDBoG
FE4CkebQFVBu90OeAurCQvuTfEoeiSQr0EwrJjk+gtCpTVSQ+1kMj0mX3Am0jjsHvbZfsRdlil4D
rvgMa0Dban3GizAF6gPs8LWvylDLn9u/2NfA2Ani0lJL4paqPoT2hmnAraRKJ46NOk8Im1Cpp2VT
VsGwS0M/TxmrYmpt3m82g0RnYokpZmFnKveT2qxZj4Ig1WVqxKlH/4Pbj3bHQrJ7yn7y3qf3pFyG
YlOy55VUmau7pGR/UXH4R5cv+iV9JWzwOSPKaECgiQx87K6z6GlKQdWNMpD3oWJAX4QSXMyGC+gc
UiR+Urspkz1dovB+OpN8OmorC5Sq8y7BtRAXOC7SVmv+bjLDy5h8Y2Rj+5RPgbU+Fb3k2fdhXT4q
AoKAq5GBTFmPSQKyboH1HdepLcDQmRwVcxsTSi6HTytfDagpydV7zcbRY6M5EeDSvpGAGkGWuz0d
jksRv7dHTAGwjixJjrjN0BpzP7qTqMlGh4W7o1JTiCPQozHpkqjGcVy1YTZ0y7o+6OT1Gp8miD1d
nnuUhCGhYnJRWbp+7ePr0hcZDjt6o09ODKovIYwPzHJH8PHJpGiVLDc8TTZAnOmm1EKe9t6pOAZV
u41MdBNVCpK183/TXaWpSAD8Td36lok6wBU74mK2MhB/sEC1QVwhHdOWT9WpJa0PzryZEvrT6x8L
S1ZZy4MFeJz59vt0nXmhkQ3ElJMUI9gyHAstZ0all68RSHxxKQtEwJbzi1imCE6IwfQjXz4fwRKE
FJtloijDScSk0BeL4uPYpO/96Koj6x2exrwDQT9JbS2Ocdo8gOtjJIKqVo+HMeZrNtHxmiYflaD2
7JNxO4Av3r1tGIu/VmKsINgNU8u6HFKsGDHgWsPRc10KONhzlkcW9dnwXcSc69ZB84hUTVnuCJb0
bAg+oYY++K5Uuvk/hO2LimNhlrUMSy4cRgvx8TTjxiFXTQBFRrsPXncudlN5Oi6oSrz3yjbNcRZs
71kG1qRwU+ypiqc05UkRIFhpEiwDUPAHM8oOrEEJ2q7Ba0F+tgNercZSMb9AybsVdmUDrZR8oSec
dHGjFGBTQRBADpK2pL2gZx3YtjLEcXPcKGpUpU71MIArpPXpyb88wbSk+0aDS7644tMfOojsjzYc
N/zBsLsJPoZ9bu2TOOgsRTwEiunRZOAPhmAS1IYWoMa/6Un5YQ3agqr49qGTBLSImWXSAB7RUMzN
6x5o8/TDhxNNjVn7EdAdLtWSUDABwiDJ19/yosChjSLAL9/sVqnpX2CsIkz4wu7n4d/opJ3xR3h7
VlPdO/tMySbzMW+AoQkeDw+fyWov9Q9E9Bo9amzaAiO8cecuvJPUBtqkNt5iejrRoGhBO0vJHi7f
rf8QscjIL8k70sc8WlL8hyXqoYfelmQpcj62hjMK3jPMsQ0Z3VXcQsGMRrCPBbSlqDfaTCfwi0mO
JOgtJx8AeZB3QbdOzuyJMQNPIwwD4zw0Ipxsyx4JJj5rwBUyX8S7tfGi8n9TxgSJyCvZ9rcdQ8Z4
dibevaYwo3EEEwcWRjCUnxGAzZe7WG6t7kHMR62bVzlVhC3Dh+ectakomnt6b4/sbGwmXJUOK6wj
VFl5sZ/4dRS7tdw34Jb5E47RFmTvNHP4/YzKxJ//DGjC9r4g4Gr153/QLjnXq23K88c+HqUH+exY
Bs1dh0aF8L4q/49gsH8I2Eg+9mu0K0C/TwM7eMEdgLTQtz22b+ajrxPd+z7msiaPGstNBM0H9XVA
pOm5KMnbEPs4jLXddg87ycmcvPRjpwsOXa+WryP4eeUGXrwT3+C9QV+zGIBZDnI7/XHDqxbupsdR
OKTKPYhoi8Y2jeY+we5MLASCegZTzYHI2Yi/odqR35k+dNODDx/VuW8yRsbShfmm+0skAkoB9suN
IK2ND5S5BJM4Yy9Bn/F+yBg2cu6zqkEe7qsFLLN8bZVBVlAVyjo0wBelgdZcC2DDCIGt2G3X6xBP
4x14jIMJx2GDDcBg7TzzcEQabaRZh5XmFfuKvj0q/oYgGAZILNTr8iqFgXlIYHOdEzYVjig5XCvt
nl/IIoSxCEHVad3+VrmdpSLFIUsypSQ9XuUZht71a7oUz0mfZ3Ddjwct6j77ATJXIl5grYsqBGWY
XsrEjRe2+JIkIUdNpLVMQNMqmFF9D83lDKVl9Zf+bBQg4/71XnhmeK72HRJ9ufy09Lh5exGEKIgS
qUimlC7GmMXmauuvIx3m6m2+tu+QrX9mmH1XOGFlHh9AjNjgkJvPcqhdWKuHp0Jt1RkIsOvgHfmM
q5YdIJPBE2wlKu+NtwYo29g86z7VHCK9gFIB+S1Ooq0XpnuW17YRe1RMNm+nTo5jLZXC0ax2+54G
BnzKiK60PLzZSZHJpQUVWxFi1oEVYMMyITdSN9SeVR1YnR5Gor8ut3i03+992I0lQrY0wurG8Q8i
fyKU12hRsEI2eZUyY4FfYgC4mFgrJYKFN91fiT7+iblj4dtXx09lf/Jn5/gmHlv0v0Rpf4WKCDZw
eyjRTJTync1nM73Hn8huoh+ydwsdxWC/+Mn5Qo6MB0FwKcxl8Gp4iM4EQE3IS2xTVRy4pUvxQiPP
up3Mfp9LPpqifqxxXhwi2C8Ez6RN6WYGzJ8yVnwR95UGN2lzGKYI8yLx+Yv8AgNBnEwQ1rhjfmaV
snpsltxLUIw5DgXQIJm+RgUcO0oDk12XY6mDvQrhKaN2Rm61vD7dE/RaubggA/uOUD8wwn0dVvgv
/VSRjIiK9UZTMhjqORH5YSQDTb5RVUH1Fj2RLZacwHWlfnWtqpkcel5nwjBI18gcpbBzcmKndv1x
naAxBq5HttQUILMfVkvunYGe5W4EYPh2EGLiwFKdx6A0RkopHt3acpWwWae9+9AQkjqGmGpwyNaF
wfxDzR4V1XaIwzLTWiVoWLahytNPWCQuVFQO9C6Tt+oZcYriAcOJ1U2o4nk3Ny771LoK1j7rPJsF
a5rIFbby2osQemml6y/fjv/PGCP1QywSiAKlfkLysMYdzfytakVRryaBcTCIFcaCZf4/7h50ZT6n
+pj6cQQaQ9EgOgJ3mNMxDdCEPEp6/7cnBsoTNj4q4B4+KZrG4lrufiB3CzNTxG+WwdTvCRBynr5Z
faIwjtcLbRe9BTHPGWHUyAkHciO3GvbYtlPrqR90sasFVasQwWppOPEMB64NwKY2N3UZMhMmJ1yz
mZDRksbcGrQNiTIqnesvkCt1RD9kb5XbwJ0bf6da40WG7bsntLuSpCajZXUGLAt9s4oOFikwPb22
YflTfM5r8V3cHshfA1GOocnYvwgv8gORYNe+hUlPSbsyptoaW+yTOZA6g3Vof0DE+oI67mKWAj/u
z6QgvXZxXrgVSYazkx09Oabb4rZ0yhmTE3vn4j/uGHIzZSzvYYbeoMcG6OFnCSg7ZMEetP8CLoDY
z+z5mSLaRExkCJ+BDkyYj8ooaRx1qD5Usum+6KLYYPRYsyUQL23x44WX1FOIvxNWQsvXgz/732nZ
tV+bt32VU9KkxyM65uRLsjKWZ3k9+zO3w+u+2y7CGYO7/c27fTmQc6YOIDdRUfb63NvyigQ5b2hp
MM/i1mN6vtBBRChQ00EpLkh4gZruYNtrLWnXbuz489G6vCeboUCPD+ZYz6pIlHcZz3JnJHZCC6An
28nyLtZcbO3ImwhISWdFKaFX0nroLeueBufzE7rj7I0nKTaTz1iIMPqJKj2AjtruYgWTGAs/N/A/
VluirQQ0jhH7JgGm83d0spY4X4i+K8elB10ChOgx4DKrZlF2kWeEVbeood04HkLTREggdYDZg6Q1
UrdMIR8fUad55e4kQ9bzNYpYv/+Kp1LwQxTSphsD//EBCRNt5I+pzX719v2bS5Q5hHA9IZBuNxk6
MDqHPawa+o4AtVyVf8ihy7HdYXrue9bBcZhon7iyJ8AwafgyRMXsy+H+6VzFS1jUafn0aMAghW8W
3wT2thnWDOMsPfqeILdxcQGKX28rNU2LLarcR4JYBXqq4VcEk9Xc1FM594VGVhYEZ4U5vEGr/bR2
0WcFrB2zDbgomhpLis95JvkQ07a3zT3XFTutl4wIAPUmZUij3rdh4w7mDT6Xo0cmEtScGz7KwOXS
icGbdunnGsdWffcPzy/ufhtId85o91x48rsx3SUIBZFg81Khom6G8F/r5Qp4gbImVor7QH+DFEFD
M5cq2O7zX8j66bC9Z8tVdxgFbiK4CuRmEZ9dlqDIgkUlCs2iV1mva03EseWYp6mm6gUzvVqstcMc
CD1C6Yiih99oFZtolMiQ+YW2JUxITg11wNLeNy0zvOA+D+Lcs5XiVZnTtuSFwdRfmN/X4GMjIU/o
IT8DHgViIb0dkBocA0rEB2nFQlwOdg1HAHpjAEfOuOPyfBk+pbaAoM74AbxddYxGzRTl27Auxior
yvqqYjgwo+a0O0pt6IqdLLsZMJ4lrIYlkfHUhczYKUhbXubNULHzGpGOqRdbMqXMvh479OgcPBPq
G39/L8USK2QMQH4Wxp0fG+OCQBjYzq5GgfApJv+NEmTGKhbPXU3mx20wIBOQ4V/SBr1tL/4grhEP
vC0qLV6eh9LMH5JDtXN8pZ69j2rwysHugngZIG7wMzfzBGf1EHp8ObU6HMD4rkILLL7LhiZpvbQV
JUm27k6STTR5PNBJbFUarMDOUT5IRVpmNVmFsbFox41nTiz+C8DZajX+OyZERIStmH4Ozile0tG9
g++hMQAynW4rIFlvZbeUiU74uDNTbibyLurzue79VRP+Ad7mGxIBPXlBHpnBghSKAwknCZBo5RuR
uLwhpirI+oKH0XtfWWM5S+cH8paAONm7LY7BOLICKzNCbdtSrHNsruxRDN3Du6lXF+uqZuV7V086
CpzOLiYf7mZ/icfA3zKqzX3TMP5Z6POtxJxTKGLV5VbcNk75HwahSZBaTjAAyBnKUe8WXTL9vwmH
649G07QDbeEWzndNeO8P1vx4Rwa29xr31FcwMUVXavh6u6iooPIof++OKlBm7HNifCJjKKPFTmtU
mCYOxXKMY4ff6CuXnLH0IOrDUPgpi6U9BDGUh4CpODGQ/uFOAPkHn2p7Jw1r8+7V/6coYw0hjBZL
QemaQ6joo4eFOhidYWe3vckbHzyg76R62AJ+tZ7kmWWztKBNVXF8ICYcNL9Abl5zHuiwgFi4/pBF
2nmIr18MIrsGHsxgEuovoJRSKQuukvRufy0SSCGDwvQ2o5BmN1zhCTcWvL53VOzdoPkw48p462nr
rMgpxk8QcxgGjbH79L3zWvmOcjXoYygXTJyQg/UdsN5c4T72XUAns+KceLiBYAoQ4jB8Rq3Mf1MG
cDn/RgX/4TzKyha7dzcRQU1lAg0MFRgnCiXQCtzJYWwsDYo70LLrPrq730PZG9zv7m+3uQzkRsEH
6QD6jTg7UGRYM9Z5wvadoH2WXf94nYQzOoJ0xTQQaawOZdgCfkHSdgT8ti0TyImMVSX6/40oeVP6
uvdry0CBv2x6GkXflwL3KGiBbXmd0i6g2CAAumXoA9BVG7LWSk0AsaNlSwPOtHlKnqQuKYDSjxSZ
cdkG9Jhlpue95K4gJcpeJ9PBZy6hr/DxUIdrBH0MxK5SfYQl4nlmHmZ166GOlEN7ejaWeovrKNJQ
6PbY0TfO1dI+8tJySxSMuC8sv/iWc8+MomkYgj8/98e60jKeUuSqV113uhMvgIpG7IP2cUsRugeT
MQnDAx4yyoGFAumkVlxsiDBhIkacCqT6DkZDatQbYB7c3qbZngES2swCqrXkCfph01HYFKpTA9QR
1rObH2AuQFzszCi2dAZZkcsUj8Us7dI7mRowc12jR1RC3sIK+C2ZTwsEwVSsSaAOCbt4uDZFoso1
g6Af37bcQwqkOlF7oiZuhq1i7Nq1OOucVJp+hakRJBHu7VvMUYmbIn/LlqwYmx9ebf4kQfLch2fZ
WVv4BLqeJjB28cuAH4d/D0MGSYMYm3He/YVlEtbnbCmNuzoUBb7XYvcyw6gyQ+hDnvIBWPpDXI1f
DmDTEs06bb3qiwGfK6uK/DGRXyIdFd+Uq4U9xyV9W97sgX0mB9asmBdsrYYbswVyGCB1I0K8N4tp
UrQl4cpb92mcGAKT9bi5uY0SouZrU7ipM6e+zBpDXycoVBvMrvTKZFHonpUJNFgYwOml6n9+4e9C
hZ6tQvHt8WmirJZO0DXFTqcNAjU7HWBlpy9sMHlV+9pwfZIoIH1Gs4sIYkpN0rzcLGrDoTBiqWBi
X82e/v6llMDmuUjktKF2Y5BbzwAFHuJbJo4EaN3a6fJG2qz5EPyvK3eAmDCuy9G26BbSbtTjTzQB
LqcLld4I2Y+hfOfgb2VSSWx7nv5xRN8BA+4of2CcbubXhLjSCdJ5MiJd8StfvJ1/JXsA24OMCPGw
xCo5VLcWFNzlwR0F4e67mmf++VYvaD5iHw4pe1WjY7VrhSda2VGzy3mHdrb6EIFDExt8euIi05su
kt9Xia38/k48O0xvMtcERebUp9xGOrZCMTwfd89Gmj5Uu3swQJWrK59SLHPySNiXwrsNbtqEoNri
sdN0Jh6z9d2WlEqlyVTPq5kS9Po3mV1bcSHdLdUPGSQSv4UCf3kTqcRiz2ETqEImlnznyhfXHyRm
gcwTE1RZ6J6CkqvtPP5uFLpEC9CbkFguKxW/ku7InzXvxeD0JVGb/4pjnVF+EEwK2CVz1KODPq7S
KHMDAmhoecdM7dO7BhaxVJwcUSgAe1jpxLXiBtUhae/l5+kjK6xXWQngG2iK2HDbyTFXROLjxIvA
11jCmarkbyOfPgTniFlA+ERdogHj22BgLougVz5nQ1mmMFyMh749k+MtaDxUBoo+fQLuUcROG0X5
tbUPeEV2QaXNkb+oVzDkpxs5sNy6g4ix32xW9nUCL/Uxtg8VvmfOn/BGVg/5eW/jhkHYt7dcIHAr
P54tJX3kTG0nvbW2gUnTzxwriPeaU2xDI2xlt4/G5oswXfKMve6PXcHBsZcPvryyuTi3chVSUFKN
mFKVwCnCzUvj0pnHkmIWOfDZYDzh3uake2f2mZ0AyMu3uQYfpqJ/yRgkX7ziteYPsV9eR+lfYV0C
elTrPVa04jhiBjBcFVtweGnsd7Nq+Ng72zNeUb9811w8U5kVTzGmSnq4yigfdBjuwm0p5y40N1R4
2KOva9bve23X/PGt4lKZINlpPG7Kio8Wu9Kmo2FENvocvIfR7XdRtIOEZhzAPQInij0B1THK3X7i
4sdqI5UnAAMDJ+QgWF7wgPoaXjIYoRnpvbuzzWN+xpZHcDnOw5rTZAuFepuzgLZuSINbF64iCe0j
TgS5XJddqFZH/hEENKx8rv2iJwH/7spQe6PsgMLS0jy7q4h6ZRxSH+5WbFn+6ll/nZeazMOBlE28
YZm79kZQkagEifjDJEBuQDpf/Ekb1CE67gY1uwTxDlCqkSzEU3zr7qVc5C0YKLheRmGf/U5A/Xgp
s1z0JTMA6cNpFzp/ugNfRkgdUtLGDz22e9565PZUC6BuvelXhuahX4KlhJiKM0IcbtggmxTOio4H
GeuVAFOrq+JrbCkkARC9fglTOpJsxZ6mvjRZUFGhxKcuCOgLDS1c4VFDv0+s9kCGuSkn+fPd2OFB
nCKIAr+/Sz7F2ka2ifp/DT2bp0C82AZuiL4ntSN1klSM0lIZp3tl1U+Yy8JNJea1+8zrQwAKY/po
9nvjX/rEGAyCzJIARB2dOjOGkGjQs01hyMA1RURY5Er4G5WPcFsy25NvR+SeGW7IjiDVWLnhfKk9
lHA18kcrHxBE93oJolcAOyaDHe8gsCE4fiAX4NfUSXHUNshUte9HB+3FjKKrn44NhddvyvtG6g+c
rZ94JJGPLCcze/aKwu+dFRlV8okN34yGBU3W5264DgbAs0cuO4PwSkaFvJcgxYmN0ezb1hvhltrX
rqi+xerD9CT9W3nQyJx6Xz56wDvloJMmGANuAPN286KvS9v4LTM5faLcyFiVZ9fo4kYDTA5ZnMkq
7X97MK8+HQZ3xEUTjGbplK7ECpY7Ca0gprhEMIcxG6sum5kw9q49YxTJvycUDeyOxWS55EKWwhZZ
wEOaBjjWEhacYnoXP2ZsRsc8dw8PuVXZqYnNuDthqjoShMQ2QA3dyoWUBXvN5gcJylrp3kEGIlh8
5HEA7RZtO7mqGbl1r4R0Y5qChk9CTWENnfJu3A33VqEMykdGtrKwyneH1PeL4umcmIXeA2LeOHV7
nHSZNSoinaeVJxPUKbH5GCF3aC1CXXq5vlIZQRmFGu4WEBlEkC3u8LaVmZ1ZGb/BjsqxJE+FXYpU
xj7/DjPyWtaH/1Hsz89bBGvXPsiVmcxOe46Cw52KKI0zNwfSkEL/EpVwvXySsGLUi8HWp6lCCoEq
W1mJuJbIeuiGvc2Oicz6AIQdW81/psafOY8IM7W2ER9VjHzRGhkez8vVPuzRwzkNf6WmD0A5LCZV
S7INHv1QVG7LiO8XVedV3IPQAFHPpnRptdNStyrqNGxAOKV/WvLBj1F8ujdt0zjWGmOzA5m11pqz
hiJijpxt2mLKfw3zV8SHGP0oHXB0YvQO9yebQlWH4oxwY+BNb2TD4MLL40gTrieT9TtK2Mg9eqWy
NfueXk/7xVvdxrVjq7nAQCiDyul9i6tZ0eq69k7SA2aGX/kjNkNQoqf+iHlt1AVc1Gd9PTpBwLYg
UVPH64NO3o87+GYOeBbmYh++4zZ2X7CeHCN21H24ctkYK+uqCGvKeGhlMBM8IO8AnZ+jOBfUzDXw
xkFN/7uQWsSAFSdSiC0ziwjs+UhnXi7/NEvzbHYbUKfYJYcP735z93OWICftHlYc46GyU8UTK7gw
U/UVNPalyzalmW+tvLkWZRDp4jp4eiwGDeZPMrZtvnS66fsQ0mskS6Foy3zddFEU+wzTW+JBHnZp
jyFdvXNfy3Vb/RmHxPOsDB58H1bwE52yjaN4OIK0le36u/XkpPQqf7LezySpphbNa9x/cnGEZhTO
69Bfmm4zoABCOu6nAhIG5XHNrvsuYM18NL917WiFwrs3MtAWJD93t4uXsXdel4zN+cWXkgWVAgGH
00Ar/QiGmbBVy+3qXcpCE+VuMvg6Evd03IwzBCkhlwj8L/Do76/2rLV1tOaQmHlmNCQHDnlZJD3A
DF4qaE9hSwH2xBdCfHbi9IbmlnBD+Lye/eoqvTc3qXqm8M+WHxlZGx8WrBuPEslN7mGx/cK8xJMj
C6xIIPkEMfy48hMQI4KdMqO+vGc9LgF4HlwJ18Q0SNIrlQMyT0zmilp1MAeC8Qhy8YATkMVwpCpD
ANjmv2Pv4i5+c7F5+Qi00CxUl6vqP+YRleC3RlI9R8B3+JxrQZK5Yea1Y4g69OocOd7sI1/jpzEm
YvISjYGo0WavUPrPl1QL13CacmUyta6qttUnQb/OeZ2Nw2MmUqdIlT01VILZLlFH69DwTs2sAogg
aPj0UDMb95JXmPNz62tT+As7/Ykf+tO+z44KX/xb9N+ndPn/KSegr8Uj2VtQlTmowUh7MttYXEGP
dLjFAXt9c9Moz9RLmykOPUTnPsL4ACvJyU4mgahtwDTCCRIJ5SgJ6h8jslgX1RjoblEDOI1UwloU
Ov2wAkH/sTTmtDO6b8SP+VqaF3mZdVYuenWCxN2qaEDHaRm3gcm37spIxRcw65A2HQLX2Ze5qizx
FGwHyM38Xd+kZDLbOikXpAA/uvhGViRhjPXCwn21uQhYLKX3s90FZiv3h7Z5KzLYZkrW3UUElwYa
k87dfwOE9RNQCcG3Jk77b3IktFEztJmXGhm9P9HptrU6rQ5tLZwcLYe11v76XelR3ZFvC0pBZUn6
ReFVthj/Y43WpEqKNJAs0IVcInrlLRwVpfMuaIpNl7qZve6EC8KIAqlp1ekr4AJ9dwWcvFYRcnHu
tbe1EvnH0U8diTffsIq3RRPlCcS5ROyoZJqsDhEVMz366zkMQzL30PTNu/OR+jLR/9lYmjBVTkfr
NdmkRShnD2giPAQsooFtQw19+Pck2pWZq3Vfw8zXvwImWk2H/rgbVnQCr5gtHLw3qGMATFvfH+re
sYGNLQISDhBamC798ngNgSQR2pyiZfL04ewMtRBRXwKENGTAO+jR1yjzssrGTi3JPfqq/w7yb/kh
v2wqRwyiAAbT3wfEGy8FeUcF4hkuYeW377glAOOUsn+TOXWunryG11ZSlyh98QjkT6fUSRXVXSZR
KTDQ1t08Ur7bM/VTqFQ7FEKTsgMBi2H5K4i2YS+A4PKwowVvjEvQUjkyCdlTKFrsp2kKS1I6plCM
c94HuHzu/hg+tOVgKKByFoCxpZtHp7vXPITuU6XYsOP+dUZKrQyJK3UzgF2D9UpKf9tw1DIcpNB4
35STlTOe+83L232VTObOJ5oLUfI61BjnHZwYNmhRhG/QyjggWsgZmP6bERgPhWGtiDbJgPwAmMbS
GatbiXIZC7aEW5I5bEjQrcOMHRQWtekFyFsgvuuFLFRiqfADv2qoujYvRvHBQAvjxU+Z5nevlUMd
dbVEkwGJ3c8smXaXhgzNLp0iDiZ6fvkKjWoXH22C9LKRO54jgIpzCb760n7tL6CrleSckdOeoLPe
JuijzVye47RHDsbZnJJq4DE8Kk5ey64431PYjf94JczGWD6QVPvoyAdE5X2sXdVXmjRSgf3NYdtk
N2ClgmJEtjZI1tZeZtqFtGZKbzRry8JqDYkI3fD2LDaEy7XiXbhxEBcMwy02AlL6bdh+iyghurTc
nUGMVHEzomJ/4f3bOJAJ/TQH88ATfpODnRw7K3Xc+Bg1DYAH9ril8f1oJGdYPHmEqnbZZxnE5RId
dTxirjnvylByVugb3VUyiyjzrcrTISzO31GQzYXjnh9O0cYnRJNkDb9maHqzKfHki6iGXCIP3/2X
/gTgJIhfQk2yVY9Kvj0wSinXR3PEvauLPeJklRgJkbx9vwCdhltvGVWBrLxEUhEmBCo9uDGP51av
Bn9kveezrbvDnR0eqFT3RRn/SmFkSngRGxaLqdyeXCBIZywx/rjFhypEUcT5QXLAWaAgpYvTSe6G
n9wWJhGIyBbj2xLgDz3Ut4fXQ2X3Hrj0VCzI0K00vG9ihi5V40b5YAnSyfFnpPqc8Q3QTYYzxnzn
iFrnPg0LLbfFuslkphpxslQAs5mSaNdjiG55xuxDvuM/VHucB0v5LM2/mOMSVbq3F8Xcr8uDm/bb
ZQWgo5rVmPFCsnrQ4HVHr4FWdwwwnVwrz5f88aYvgQwlD9AmTq9VUl+WLkK7N82z+EHH/QxbW76N
EPsM+W049yD82oInNXcO/2KVdLGYBcmTWWTIAll9SDRwRy31lJriKiIjYlLciUwDyOKDqvsxqGuI
Qd2CEbA2rB8Bw0r7TSVAcJHoaNdnvosyAh/kM9dBHLUOILuk3vxWRBjM8gXRutDEpcGY5ys6Mb+u
5zmzQSX3GoQ2O0AdJG3FBAjvRtqIP03nSuQlManddhtJgxMzTDGrnr+m5CnM0F91hqKk2nH54onu
zTrSMb3NyHO7Ox9vTvXEPm9YIYmhrSvjIlO21fdwBTsPPncJePIPtoiEJ90v5KRYzS7ATGf/Z2aQ
1uzfJMgHQplEafytwAW0yXsyl6KujjdFqk1fHE7fKFAGCJmQ0zzz5NYSo+6rbEIaHBvABsaGJ1oM
C8IyhpTodl1TVYM00r6uNUpfHftDSS4z0CZcye3K8HS/sbcB1e208gtXTFaT/Z1WuG5uvgYVRuMo
DoOrTg3XypA2gXNzuDdKjwRqMSbkmqgAbLM88hkWvUHwHYLh6a7uoOPOJTnEHcjLdbLbLS6v7ams
bFHgC7r62bGrWGwL5jVJFP1UsdRJ5fGHctBfNpLLiKM5Q9LcIHNzf+bGPLdUhPG+HWTc7tzieYUi
gZnCq0mt+W0jXHzxRYo6PVnTf8Lt9sdAgZ/kn7XO6lb9eJdq8qvUO5ZUpiuZh8AKk8JZABRAvZbs
pmYMMAikMpTAsS94I4aUd167IAEPR91eRIKTeolYNI0/T2ZN0qMa1dP8OaJsi2xntNVr4zE3DjMR
j9eQBgJpzx0VdlOMPbUNJxIbNaghn71rn4y/c8/c1tTubmqvG5d07562BWBsLOdKBVG0c8qerdtU
gfl0JDOci4isTiCwcMPESghyZgsEsf8sWbmz9EVu6WlHfssiuGgy+xmJTFhcKM1+hsMKufGXnmOD
l1jd5c2RQF1keJCuwe2PmU2Wx/bOV7x0PxFJbhYcOCAz+Nr0BlL7DAzJ5/6TJcS8e+KFj67Nz4db
HDs0HrClpvd9roBr/MmvpSpy0Y1aRvy5dYcDHctKIqFvJ3KFaHfEMRxJm44tdmNGoHnlLc0c+pX6
1Pnh1gaRznQPHkbtv7Nv105bblKqy0NXUbTPSs4maNlcN4w/Fabv1rLny4IblA4pe+WorGcuN0ry
Q4SX0OwfGHXIAXmUx7ar7jNz8OQmM02RXKtA0U2k1j2mKzyizjz3pCKwsLOWL3WBilHeEj1IBOjC
HtlEpl6oL7CP0hdrMzq2tb6TVnT+w+5eMt+FDqc1gk/8LU7HF7ITRGIuhbaIOGc4idrUQbXdJfS2
OEtU98IM9hIU2fzGNwbwQ0GQVPPGC941FPW4NQlgNoVm+Mq455twGABioXTg7P96R23RAZZNjXYK
VZJnBHz5OcUYIAmIfvKq9LJG/1S9vrsCfn50hckCNL7ckLQHUOF7TnFQuGaFGGIqf4pfA6JN935w
2007drcnR7l1C3hwyKB7V0gAbMR9Js/2fH0joNqkBBEAJLXM1yCb0DhG0KB7lEkMJda66W/Bv+LY
lfGCCc7tOCopN+fBoW4bmxcu0qTjwbOHBqjLflrN/OyCCV2L1wyrOpZaGKyN5KVfJzZznapgv5Es
kbwqesYe87S3RK2q8eR1Vyj0kAEk2zy0Tb3E6di2EdcTju18w/QsN8X8ynkBcMbjqaN3Dcw4sHcv
AEn7/4WI5TNJnnT3hjk8N2Dt4LN4Nq6Bsat9D2rl4Cf2AlPxZCUvPno709vShF81uQQCObLute5A
bZl5QwbpoNRH3gbXC2PeRqlb5WHWfICImNtaNbWrEzksNa5pwPN7G+f9seAzYDH9w6F4xTb+BKcL
ofxSq/JprR1cDa3+KNSSghlokfAFl8QbPtnFbbE2QCnSDI+nb2oSI8R3PTkGdHOw1NM94LjkUQwe
wS39AjdQU/iyd9BMo9a78KtAZnOYfw+i1Av3rTPChRgtQT43bG5f3vvE8GONDhkS7+JhsO5X3K4h
RSXzfPNZbbAy9c4fceDYoKrVhpkc64fIiPoA+oavPMcp7dNYQoR34qPBiCP+EPLn0gpIJWQ0XBnW
UlspJloSTBk6c1uHzfJN/i8E0oPEb6Re8uTS5r+yBif1pClZL5jjw+nYFMsNQ2Tt6pFrZpi5mjJM
pNq2JJSiriD/NJEHmwieWGmPvp5NBYDqegnJCbQDWMOoBfZa6aha6Pqk8KcnjB2DDgJXsow9qRao
RIOFFYQ3Z9FLNvjG5g+MYvh6c3FcXya12RRGVMxBrFoqaqFZ8+YdoBh/4srtEV0SX0z0oTHKT6Vg
2NPoXAmMy7DnNHDuaj9kA70aeFOls2I3qLrqxZoslRG/k6g6hlF6ivuGdzHwp0cMqF3Q2BN91YS5
8HGNnQ9h9rdvg9jVFHU2R73rmsbd0WKFb/Ld0Tbmk3mnjeMCqHOdI2D6uIof/H+JAolGwWJDsTP8
gcMtOnEoJC+k5TFNBgfLGiTdeFkC0scTsjWWEJbmO12SuUP1pdaMSd7kCJ40rroj0RoGb9WnPwGC
c8TnuOCTyfOBydal4B242O5M/rN60TWpwYBlrra3S3ZInf2T4cdy+60HoGvmROmRqn7adNLcdSEQ
AnqQQrKOw09oBDLo6YzTHXeavtFrEgXOd5mPZPURAaIAkC9cXwY6wWXLzkLVIl0/MzrJs/Ljdbts
bo16SPDoxpbCjXVf28e1esa3I93iPzjmA8gHG42MtqzXYQXGPF8nMq189qurO/vqLBPs1FfdKljx
NcUeLyQbCe3k3I/Oy3QUiBY82GXvbOVaQY+ihtKcKhFds+jkUWwhACC46NzxPAntTwBlbfolCIQT
ZXgMJDxll8g61A2DTqEJvkoCbhdS368+myGp6WHFGhjiqlaIB4w9xMlVgUSkIJ4BO1b5uj9/40eA
rtI777tV8cty56uF4CZEzL5p27SQxIUTVzshsRqgm2Z6UscX0lj9ALWKnGjyvzW6JiJt3sXAhIKp
lGlyqVs78CxCXCXEX3TjxjOQ++NDV9kyRiYKBKoFzQzRgtj5LfkZBVP3RTctmnQt6eDnVrmJ690B
8iRKXruEk4f+P+unL6c1pkfdGQBZiAK3sq2cpVvqi0ZY7moDu+JfMh39yHCafJr5HwPwoaZb2Ypw
m3RIfHA0M4vHuW6DTCfBdSRVLw25ZJ9/7wxUgZTFVPGI5L/Hu7DbUioToS8luy9fgxzr9mn7WKKf
bhWFq3jZi/gvqBCW6xxpewMphbJKqI2xti3XfTW/X1qBdG1nyJwQdxUPhGsAg3Kn/aNYLn9nyldO
jvh/9xRIG2l59D2sUbQiuUBzzft4y7ztI07yjh4RSurQ/GC5kjfGB2CNGqDf/ItG2RRBgWxnc40V
DkEidFMflAwBUkPD8T/Iqijgl/i3lItw47xlz/eg4R1MRv8NPO+FsGec93fgnKJU3n8Mv3Ysm++F
PpcsZ2VJkENXb0UfaT3h+vrplJMQsHxGa15JXKH1ZQAu0QWYRouWmJ4CreYZK22L26gv72D+FZAy
cDUBF5a1WEroQzZu8EqzJBIsiJ51ExQr6HP0bmtKUvbOdqQ5OrctMlZdi5G9NyU/bNjb8deF80e/
Yqke4sPT1Oyy3rIcuslqHmUHnFXayUnrQFkeoOTPrlk/rh4tPUWW43H6hBSvNLZdR9WxvzrS9n3B
XryllE8gV88dDu9tuef8ZVjWzu7ttT+ppzn4JJTJ3It/rG3/x2+t4Auv/tM0/Km3hFzQe55HO3ih
VllIXf6avV5w8QMDLQfV3k1D+FKOV9G+qoshnpQVFxBVF62XYgGNcALYBX9IcbbMCp88XXWwYRNi
S71vqT3zrxIWo8hAOm8wRGTu9Gns/SoT7sBFnAsPyHQ5J/l1DltBi8w1Y2sap0WeC69j9rxtgHvt
vfyFDgkMFPt/YqQFpczDNj3oe5ZnkVdLcvUfhiB1+iq6ijmaPx70V4WMCt8vk+sR+Nv2JGhXQLL+
Mne3W2hyTtfLeGRpXcJgT4vGQRGMjWv30qcIQSxwJ2vbb76P4Y9Tbi9T6qv8akoovI50+mg4Mf5i
HBZcLEW94Tn6X4cQHnP8SKyt4uxL6Q1FhmSzwegXcIBn8uTBBPFK1mvwu6sAPsENtvrtmu/6G7ge
XqY6D5anwkVl7jMRN9gOUWuYK7uo1ujBf4hP/nK8IeMAKmt0SuCLB+bAzy5ta2OujZf6pYkM5OJz
lWlXaWTc+Qlf9UD5OqXOgNmRgW5IceNpBATKf/EQb69ONFoPljZA89BuM0xSWVasJbIFyV7hWuPM
GVoKF2FMPWVmYADngjzLaJNbE0vCTWEdiJrdx1Wj4XWZ9gLKW0b1ugUMGPaSeUYYtIn6y3J01dXp
pHCpGd5O2Ro4XqWhNH5gqLTdLvpiH/eDADZcb8syO/wtx+1MZhXQdxbs1yxSeIcFEOuqWInrE5s3
Arr6EM34AZIVEB16cKK4FbEqUcA2871P7+F8Ew0o0P93+fjGuQ4Oc2X6KZEz8pPk/tEstgr7wP4b
qVSfDH3aCpTK+GAu1rQLcbuu+N3KjdcBh+M627j5lZwxRs3vqBneOt5naFJ9lYurVpRz5nVIGo5l
5t2/gWHtJAFuYjcnXs3cfzAZrCL5jDnSbintnhqBURsUFrm5n5z2YTPIdcEzBl1Es6eWdka8iDTY
l7k0ywt2nlLPCf8kHMPTqJW0aH9CQjIAxW3yMIdSGSm5lIs/RLhlq7M6BJPwy3fJxHc0F33k37VN
4NMUXbhKDt3VTu+/XnFYhpiUcHQ8V+mLrFBYCgIC4+FWL6f0CGAR2NYmmsCooukSEPZhCpIGpELS
+TNoVyia7KW6HjD7W5VfmBxJfDUHD1/YOK4zRO/R8KbfuSX3L4jIcrQ16paCoesCxAWr4lbjs+el
G2zRwYZld3ELxneu97uQdOCvC+BHsAaykLqPQJbBAr+bgJefrLYinHcf/NwGSsC+qy92kUyiO4PS
9lgWRuFq56y6iSrJCtW/xIKxuZpImxihGyawITlhBSG0zsed2+P+S/IFCGXLa/u6p6C46DByW2qQ
8YR/vE3BlYDI3RE3y4K0OtJoujOUa9m6aU3rfc2xMwPrXWZ4JDo+RAvfAk4S8b9rEA1kkbfkohqT
n15br6DNuYiLtvpLtfYMLZezFcMbI/QYDyDDnQR2i/HuqKpqmeVgXBMlEqhOsvtAsiXK64MqUfIn
4pzPDJhQfr6ZdJXGQ2qOAujkmO1GJiOxUAFu7a1u2pD8nH2MtP24twhIttaqKnsHOGDzcRisP9z0
bW3B/RoEbrIOzKjk1No9xHnUkIZM/niHeVk1H+PCRERHl3nj4fWfiN8zsTXrxM24Xe30qs4/7Mf4
RgMs+kBk+XMFlajdE0M1EsgQj0h/OtSqZAysWgKbODPMRRuPBMP/Ov0PrsHIF3hmM82NC69RX+aO
FZb0KJ1X3SG+Pm36xakPQvA2RhQk34P/p/BProxrp4g91R0AcNvD6IV2YOA70dOWSMGfDZogKkJw
tkG36NiVvTtZKY1DH3kw4exZ+zFftM3D4BAFuaE/PB5Pd7vRBSUw9SAag5BQc5zGbOrZBRUrWZRz
2uVaWHsniTNw3BQLxi7Jq3W6EL8XqUHTY5bixYNntDovUvmbLfLjQ4oa0LRpBDqgmhFiA691g+Rh
LAk9kncoD9xGxcxovnzmwkmHOqctiPtLlhDm+ZbCu+rstDiO7pDZkzymicygx5hqhK4IzizbCqmD
9wer7OTVYBm0F80VxCT2IFHNi9lo2U3JV7o0OJMcJjPIfUv/f8DBDgY8FWJAwf26rYK48L/PS1ob
p38Tzk8Rp0Sja7DGXz8ljc0eUdiyErHuu1P4DXUG259FwGHDmBozVtZ/imEkNNIuE9K/TR4BgJ2o
PvilJnnTEk+j3AmFzbRBqr6GhkU9tZyUU6DAonkv3nhifviZlBIBUu4xSQVy0hD9uWsUa3ZoSyjR
EkIhDuMXmR5z9FJThy8uclbf+oVR8mL+GcDnH1uXcK7vx0ofui2u/u/WqIA8NVzC5mud3XcfkhHB
tiGjry3uz54Kcx6zh3DgktdRoJcAAAFR6+aMzBMCzbQ+pVFOeIpx5F6FTuhlhQpPyPCchyH1gQD/
qUbxekLQFU+dYIwLswhQNGCHxi5E6TqPZsrMJtxnxylc8vgYNKxdcmX8EgJRYDF41O84cg2I7DHM
OMBKeIK6aRv4OEwFxdCQYLuCn/avMUobr2E2OW6uTuRbF/FLIcy5VUNs+yCpjqy+cMl59JIwCFJw
JPL4pYsrqTnFum1IVslYRHLzLPv+/tyknkY8pQ6CaZvUc05FN1Vtocj8mv3INavUyN+bGVW9iK6l
H5vxqkXDWpDIcKi+8Yviu3+sYpafHYX6gqFYtpLM8n3plux9FHG14qBkqTk7jR1iUOFCKGfZoZsg
BZnh45UOK4j62VhWopWxXNnZckoB3u8Pe4bG/AocWYBbBDHpJDAuOT2m6WP2KoIRcpEvj7k9tAj/
8YlJiKTOU20K7tV+q9ngKLz7ShkQy9EmIdZGIfECtaOHLf0QtZtO1yTuPmAxjXwAxBIYT0p/XNe5
d01Ji9p7qvlRePOtEBi+xu57LonQgbjlRsuu/2BSzxB66p6qzDNIAaHTTaEu0p8B5sRjZPXcDHdQ
gix7vmjzLxHVkuMmKV2KfFLNXpjfRq0k6heN/E0P7vBAH8MWvmtuLwoygrRGKtYWjkHvPMmzo0bA
CC2x+nPZW53j1cGgcHtcsUt2wvN4mCLfpVemo442dFKe6oJ8Up0l9NwJWxmtDl6JHgXK8JBUYnB5
QQCwbYWbUgUYfVf01N8xIiQ1znkCXy97R2air7R1SUG1i7me9ohaVwfvcW7wMk2UfK3XnAIPaRR8
/EX5CzywAwVYsEzh5HvqZ/e+75eUL19sAihBGRZyKvGpLeGEQ60szkBKCKjoruaZ5JOsRmJAfkL9
SCuncXfVr5HWGJ8/lukLm1FlIaSS10wjG0jj5yBYNP5U7G8BOdYDozb3Y4WDaI9bIN5HSLFxGass
ms6pu8MRb4vOWzfQCSjpIMFwYMxQohKvhuz4gtgVjWqA+a99Y0zrfUsylMy1fz2SiIVWR3OCkwNv
wPIrJuAise5fIa2FSOjuWkRqQk9lk42Pa728x2D+m1XX+xiVREKc1QRcdJ5MiZefhl1XR0SbmkIg
0Ct0YrV8oQ4Gh1lWoozZ2r/Ae16nChviRpD1Hpj0Bt9jiZz4fdmXlcc0SemGZNIH+jk3by72UOAy
KfsagjY35dt61Qdcn0Ys4Qvgo8T00wcZXHagRTaTQsUEF17uxfVQEkc5Zdp7UCvahpIGMzgkpC0T
oiMUJTAi0ovGvXtdBPqLrPoK6rfhIgl7s6pYQctFACa7qWDno+rNE8+d093wdXnzCvBHIWLiF0b9
IzNz1JNwqZuCZjgncBSrJUa3S6IF+o6GMevNGD90evVv8L2XqQNSbIHmYOBnDOJl47qF6EZmox29
QXnOuL2gxjzU+Ksd+x45Wq68P7L/a4zK7VDnt1EDy1bgl3pTFXqPois8Br8zT1UKz1psZsvUKCZK
1S6i0qVykdWLm3gmYU1JuAdR3Bhg6vWdy67tnUAvYSElZDaqwMTU4b5i0DsBIacW8wtLscnOSeIm
NcZ73B9xPkj5vfRi8K4mHcN5NgxFEMXIwJHC1R3OZZtYBz0pcbMT9HVzs38z0AjrsIxNtOxhY2nE
OI9HooP3V82xMzfLPAn5nMEL4Y2sykzZ8wpBuVU1IC0BoPz/Ojl2n4pA+vtSKBY79htUHxaQUchC
en/C3BPClsMFXbMwc32r9t3qYRaG+JNap9nA70oZn3dwUSy88WL2OF+WcR11z/Aq3kiWEyAEuKeW
N2xy52pO8r/MVWJtYUdonE6WlXneSUKqzT+ypKXZRu+00vAHMn4+Gb6c4dYGkQ1+NJEKhXMMBP9P
V7UkowpnhXNYv1ZIbHPZPNCdTt1/TOUM5+SCf9Fkec2QcXcVduva3wMuHopNpCA664jzya2r8CWI
6meS6JFd94OiA5E73sPCkw7l2cLjBPQH4Q47q6BaClvQsVqAI3Hhn/EYVMJhdHXQqVEawWNf8Bwg
dh2AjpZWIJFOWUufcHUHrZviAL2a8QPLmEkLY6k+y6HnvTV4jL24wTnKGHd41/1M7Phz+Vq4DhhL
7UrdS2J1k2agFNcLyP7QoxAIHjEdN9hA8cUnBhWhMyfCO6ecJPj4VwKSurC9XFsAJmdNq4A2krEm
h/JZojcxRPrWIdhNw0SZ5bBhxV2U9Vhr1Isn8ILJdgdH69LUuGd2hPIXrze2ga406586xThviROZ
YqJbX8cSt6MR+WKzreYT/XlnueBj9v+fQKObFmXlzk7LB8DeVyvFTjJ1CjJQUSXXMpffQkPp81bD
O5IVsVTnjjL8mR4yy5Qq0MI1NKy0ClxnuJ9li+5JOpROm8hUOEeu6ZMj60vF1qsZPHhvB1TZ+3h+
D7mZmNCm4lMiXnyu9BjKEDGnmGMiFqHiAhhjccWXLiQs+BUt2s/XGKVTnfwnNbQ5ZQYjnROah9YO
g8U7siOj2kF8kKSvHwrY3TYudSHfVVWdub9AxoMrdwBQvx8JMiv5TlvnoqYfY/oJSkU/e7SRq6GS
fQbQqGvhgZZpBFt0ltN9VJKuUW4JwRfpweqBPIKXo48ip00z3aEUvZjqas49ZguvM2F3yJTtMvb7
od/7DC0mB+Ar8U0IvARi0oXU6VVe/y6g1U4CYCUihCqvJlAu2k8SC2SUHG4KmjZYCPb6ZoD2Xdn3
RbMe/bC5VUb0+O1tzQfxAck8+TfBsB/bVljgJgl2rlAULgFIOKQM7q1UaxrtWZigcdX/OHmLUWqZ
9J+ZXWnP3hILwxoc+TIYeAh+z/Q0sj8RaEauyjJrAwcC9dUB6fIVqrI4tHp+zvRdXD0FLS4ymt2+
TzQoFt8x00DIKhTXhZRpx6f7Zm+Ezgw6ElmX6pPB8oFtKnpeXV1p5cH4sDqu1/u0MMhlV2yUDg38
iCjuzTUhCfSN3olWbgiw5kQ1Xn+xbAs5FcndgifaTx1D/14XgHxWY3HJtLl0p3NXsMQxFvaZypuh
RZYd+iBIy5abi5P838aWpqlF8+YZdRqsnVU7hkBRgwcFfYQHZSyJp6XjN0mFNizTeZV8sB/xFqAv
1RDoCB8iAesUbuGxEL3iWVRyD9VTbH1W+1G7Y83hW3FfLYoZmKdKu4S43XdNaqvygh8WhgoO8gfF
e4bS9uBSIhVRy2nJo/jAMdtt0qCbfJQMX+JIhnZGvm3Y5kFUKi9BTQ5CO0jsqcz/QFkFvt6U6OT1
H9JBnA8gMbu5kiwCKROl8kCBNYFw6c+wPnVdLnAvDyqNPc68MK8iSXFXoPA8yLVh9E1ydP8sLOw1
250bOz8WMAAUfC4yzb9MQml21q3BkuzQWvw6W4naVmpg7oXTBdwUEqTFqxzvuYUiXbEQXuPa/l/K
2MAMtPjwcw36W4Z/FGBRD1ODjdtKZVyTfuCWQNTrMKbTaSj6mrOQzaPesUQyBlZhcKJoCn3jXcv0
ZYlFR+GFbPaDxHCApnbPj1D5M78Hx6JmPBHpeJPB8w0OZZrvTdHN4pvLo4E7NzfXslf7RvATo5AO
0ZYvD/yu/0C7CUwcNBDsgJ0BNNVTxipzqrQQymalfunwKI1ELR3+MtWqbqXx1C3WvmaLFNtaU4/u
cO4sIwY9f0vaduRBxw1p8QWsDNiTPZ1RNyj+gTGpfWFHTlZvqd92rrvTa6alhh114ixiE0tXP8vl
CCaY0/wJMp+m+4yv7KlmCBFUQH0bGNze4Qn/QUfhBjbDxQiU0RCAnvoQlI0q3bCdMX/KXGJAV4IB
oxEKWckkL1QwtYU+2SemH/1vq89kjWbWx95RuckNklocWJPbg2uFI4bqjrkPhFVUs1dR/48CVv+S
r+0HC9c2y1d2ldJfQHMLJ8Scp+ZWOKUspYfeUNkW1b/YrqIr35H/2+5E10YCCsT/idb8Dk/1H42f
os7SLDn3Ii/cm4X3cqRrxNtaY4TtT6kUOIGNbsivJxi88I+Kw22es4FV1NbpOhmK8y0ORkGOB7Wc
7A2yE/lMReiczdVqg76TtTJqxhiIMR22jUt2NkNh38x0+oX9YoxEaTJ55qTNPxlHjM8xQeNmB5n/
zEJyPdxS5VGoXGOJuxrY6cLoR2B7/IreeVsLRsAGM6rkUKRjvO1LveqTKHzeC9m5a7HBJVGwTbOs
RzPmi4e5W5ox3PjLDn4n4kUiKzVT6xwipiuozvBPD1XuVLIuWnE4HQv56ZelDuDi5SLUIbXV0mxn
oMGVopm45yweeFzviHbydwJut6OakHioJLHijxvqJQ9zqYPer9YP9x0t7fNo3F2auS6XljuCbzCX
BHrxiSuj6RdViTsSwEk1zn3DhgCkTA3xibxRCj1KxNDXOiHN/JZ+Hvy71eg54H2ABB0DFUJm12Un
YiWFSKzkkshA7mFw9OAo8JATrJKN9FP97rK+fDdarFf5ojUi2Q/Pyp1dA4Q0AlqSHieVg+ZysYbi
JXoQSwuC0lRF1sT359XCf5cphY4z9YPIFAd2enbLw0Z+jNa4MDONHtMiIV9pwLzn3EzYf8Ts4E9j
SbllMbgvz2ub8tcn+qzAi5tZ1KianAdgTPPko1/68/Dmg0i6r9dUWr4Ub1kr1FkhdUH9co3z75q8
0YqlqvRZ6cAo4OFmdTf6XmfQgPTcflKJXco7HO0ZivQR3JW1IJMFVnbCAXw9CrvJY9iaUuUEFyTY
AihUKU2UNwoEMVbdj5UJZqfV1FxU7KudrzIONf3fEnsZIIWlVprhqJysEwsgIenf6BfG7pUqzrXZ
fldyX37obBN4gtq5XFIa4EPtzi5uC2AG04O3sCvnVctzxT8xgVp8QUyoeoBMHU7Kl6ainP3h85jJ
O1Xg6JOsdW9aPL2/BSPzchEeSqCrDf2c4Ln28BISHTn2RFvLFLUP9hMHGRQj2yfoh9T1dZD8ITrs
skF87Z3/xmzf3SSrKFN9rnlFrTacSiTyfkUtEaVtUygr8aGoWC2uTZfdS6Fk0t91c2QxG3Sv5SWB
Ae/R7nHQpkhCd1YePltKOojwLOIbxUUq8bPpepxeJH4tkzgslk5a7C3l3ilSgFtQq1XuNduftOS9
5UwAvJtCaHxf8bg+iVBZ0NXb0pji3LKW6qKw7/C2MBW7vLN05aMuM//C+QtxUDQ2LEgw3BvyhGnp
+VbJYTzgGVS25HS9oMhHyu10rgbVQPFqVx4QjDNARxABsuMkvnjTpBpR0jI+DSLbTeksk6QKZT7W
5jLQICX9lzzdJzJkF1Yh2kCkveQXE6thnqV3TwVVfTO3oegQiEelJFP1ltPxITzJQOyPk6Pa0+L7
sKlNaokCDNZHMf10DOiPJdhFPgjAc+I9pxlmZlQE+elW6LzYlk8nHU4pBhC4XnAeywqnmhtF54lX
+5w/cDKkLFVdWxJcM63P2Z01yizt7kiy+x4IOjDj9rooiTe/o9XRYnbYH0SH39kCMaiBe1jeYQYP
7MVhkcn95IQyG5OpcLOzPB46EOEOsW3sZ8LuBEovkQDt3W1mH4lyWwlnV0cdaNOCPHo94mZWpI5H
8pkzxFeH2whq074CO1x6Dw/sY7hmI6/r6k3xYFAF/IbGoomp9OkQv2WfOBPnSbz723rLDCXXeJpC
z5bJsaevxtAfj2WfAx8ErmHcyXo0pOa9ysz6ApZF9oRrE4o4MokBwBluP/0sj1SaDRJp1H7nTvRx
ElVe5TkdxYaUWXO7/EHJDj4WOYlEKx+lbxbwxvx1NDoPkdSLm0alXxdaHC+GjZHmxW8/UTN5W+xK
93TWZiFlptf3GnDMrpsYPA5ASva/4CW4UWGxVg+rAvvDtvAO5HA3fQ52iGPJ6NjWdiasvJQirAil
5dAKdDn/FVk/VBQwvT8JSO0qmTKnAXlX8WmEQX8mHe2eOJbKPJe89gcEkYOMzNrXygHdYb/voq/g
TkGuzVTul2e6yEwprDor+YzQh7lZVu3hFkEr4EdpLxPd3gh3aS/VYzyI7vp/ZPe9QF9ioQ803thq
MupMfvp90EiGu4ByaumLP3X6iEHMoq7IFUf8PU78fQrcx+rzNA2MV93Iev+/9NXV4JOHyFkMWonS
tDEn/blB7V//Vz/8XfXdZ0Qr7P1/Fldsert3jDvbzbkhcKy0WMYMYwdwjYx06zrmgodmDLzitGEH
NzVoaynxh6laTaZVRhRbMGNGdEqs7c8CJTjZWoMcKMAvuH5OCK3DKKjW8P5XXSEWcAJJmxuQsurD
hog1nv/rj7xf3eakffPP8yRmBnKc5Se6RdHSTWfTFafG7DGkwKZzLCA0eqC+/us9tefjV95xgjof
ifLJv6hJflWFReE5nff1srberL2csRtOoZi87CMhqwj+/aEVdrPJkJHtC+s43O1FRctqIVSBq/Fc
oGPrlOfZTaRYAZXd74jQ4K4dSLRbAKHFWuUZB8m/yvw7yYKFO/9G+2hHzQ9HeFOCZWmvkf6CG4Wc
lZYqA79UC9wRTHvM7XAYcq1bVGzj+D4mtxHtV8j8KzvoOoI1tb1B32sl/WyUynyUt1MGcI7ZrOxK
MQ+5grC0/xqf7m5DYYBzvSdV+ZRqpd/13kJ2r2NklPPNNG60YTYdubbv4j2CQWUhtz+7Pgw0PUya
XblEK+VkIRKwpxj4QNdXELcNem55nHgSeKEIIfA0/rbAjq7lWYg9i3lBOiLT3zvXBhfjsaG3s/6E
Iyyl+AK/CwoF5Tlg23VCnUMh84ejDYtgASzqW2L/fKB4T9L+MT4ym7aEMorIMvuNtus3HMT+S0iT
3zWYGV3LyjIlAa8TbcToelmq9P8aYuQ9tEQrtjwoRktF+AYhel2iuh7GOWlFRM8i/UBq9Ainz1f7
5GPN2Q2hjbnTkoBVT4Yv0hFfWwkZHsZ79omN0TH+fi/52IilPGVf4UBaakUfInCNzkmc2HJ18sSo
sDIreYeqN/6c36Fcjl8VXCTilCUK/wYlNFHEvEaboKWi4vUSX3QMhQrBkzcxZgs4Mmbjeu91OLKa
2lV8o1nt9PsQggl5maYtDRaPbCvu5cDWeNzlEepgolDvY0PdWiAZaIX4I5EKlvfu3m8MBavLdy+t
PZmfPN5oc1OvirK1ehQkC1D4ZinTy5BuBq3iz+bLpl8nIlT5zJR+BZfEzvzU+paHn8YXwOC6l8YA
RGk6TN8piq1KfVlpBYbru+AnZYfgOdmnOkCaH5/MVlnnryip0XsiOSajgpsXewkx+LdfC+gDXc9J
F+f4QPOU9xq0E1W1/b5zSBERRpnd1wP2VYnEMRM4AFO0jeMmPIYw3IypnPAJRy3TFxgOVtCNkdPo
oB2Gh9KNTwn06m7/lgxqiCuI77gxoGSxJ82RnXwzK7FzMNX0PWetr6Y5Z/hd7A18Ij0IEJn8Qa+D
pJjXJHqgCUS7YwIBNlxBiCMTnWg7y7lHnLiYh32k78dy1SS3gtJjBmENO5cUZY29AeKWw6RYwUq3
hhLYkdvlt6Lk8In5zdRWfNqk79Ddu4vxhc5kEK3x3LYPaceAyg1z8ehV2+gfUWka77CwDATcvN53
wRSojhuRxUUrVns7KnZ9evAKvAYr519WPHv5zR+3Fj+fTgyQct1V3hmihXiMjhGxCVk6KHM3TTHt
xmEaADovx2LQp5LLOvM41bxFLXUGdkbOvQz0O8FmVsbLtA5d9RkNUbI5UQ54GagC1PLoPHzTiwXW
/CRAG+fV5mRopxVupmH30WeVUp5Rtad4fi3wd1HAaxavw7dLF8mRjee+kVM93L2gaK+MNobW7KwD
3MlhMgQ9rgDmqHLNKe9tv2UyGeXdq790WvX+4vyzjKpxe3iRFFMp/I2AawFFLsO8HKspZe+B/H7E
pu862Whgyhd9IkCldp95nRVtkkr8wdwQwEU2j0mNjvu+cZOPnc1USILCWQOulv9u7sU/7NyDdVlG
JJkWCN7OsjMq4KntvAW5liZZqc8eNxBzZGtN+TLWu8zkzghOWjqM4BBegN1foVvLum8bM+Q1VsJn
Og4gt6cfwIXoFxGK2qZyy7CjbmbdHwQhitCG82qXUoZK7Z+wDzHCOBZaL/gWio1FyylrstQw5YGj
+guVKZwL/s5sl3I2U21PmreA2EyFvTQhr4cN1s654Wxn8GI5pkwtsWzZMS/Sx0VKkHnnkH9jKdgl
paFTiNMS9twGxXIJbp99/BVBnqFy54XGsxb5shJCarSUWsCohnBdraXn1q4QfffG1xgdK7IJ76+3
mROLmf1oimHJsqF6FYJvACWQ1u0S5q8NSU2ncTLYru4u9VJ2N+TdjnWfBy6XcNAr2zbyRctOGgbg
uCRisp/IBR6l/ZlaSGoPjOFqKz7sHN117Rh33c8TzIYP1SY5OzSxetsmeJyT3k1XGuhCposXsVeG
Es889aiL/FHDk0MDFyHc+wkSjxrGyPJjIL28jPSGgHuepOeaGT0TTaA6y0VdWcDmPdh+RXMZx9cR
XIC5GynRRQ3PFOitK6EnqPzmez9UDVi+g4q3bdd1XSyt8irPNhdASY3JPdNblHxRCp2WZHkyDsDz
XFLiULT9MPnZycqH4kGEvT4TXUg2w9ACXRbafVu5sDlnYcHxP95AzrEjZRDt6xI0uWsxSG09T4Zn
VHLW7b1oHFWvMTQ6yxl6jpSOvXZgK9iB1RM91aHfZmVSqbH/UyOZ3qKBduSdhofk5asg3WV1uoVD
I0haDUTv2GCsp7ruv2Ib5SPd28vNMko9IyRqyhrzj93Zmt0TvlBWAyx9gE4YtiIjJOgtTjIvoBH0
ICRDrm3ORynOlH30YTiZQB5vAGjizcVm7f5WTjeReg4NrCgCVVQ0z75PxuDy1+wIhQ+/De00ikQA
+Jg+nBAZnu9tH/8vU+Zd1Xb5Q7YHBoBEaf+diN8eDnLfCIQAAHTdVpiaisyW+/9n9Y5NeGkkIFyd
Cq3Ry2LE/CUM/+O8QVXHRYdZN4L7NuBruWCZX1GCrEsoC5Or2eFjoOyZevvmsKw8/nDDGrZnR39E
U4bSdLSDAr+7owNxMAaQwY1iSDzjMvuMIczBbUs3jjlLl3YmKwotrX5Pwl2FI8WU/Z/8xjWjE2RK
xlgGLyPlBDN5MbRscKyq8ZV02gSsl1WASt0aN5pKZgB/B2Nef98LrD52m3/i31o+rcfhPc51a8jb
b0i8whSd22rwvts6FPlcm7Aey4k4CXyNlVY8GnCpGemCmg04K+18v45yspJW5ibTqh+87jWfbDN7
bxv2CMr7MGOrLRD1xwkOMGW98jvYXiP2wzk6971dmn3aOeHlMc+M4BzQ/tksl60NiTvix+zzNul5
s5hmcI+YtK18S5Kmu7GsCD9U2qa5PySGNurMUuoclHXqatVF83ZEkoM3NLNTDGGTgnFowOGHcBEv
ic1i8Zsi7DxqXzGRpHG1+li+r5L4C/K19uX9bp24bft2HBo6b0jWCCzuNKsRH7ZCvy7siWTTMJjO
Y9s+niAfyuxPKFzEh6oEpqBcIFZYxN6IjJEXCCvGYhUggVdWUqLW7AtTN64knvIYuQa3SZ7umrgC
VqAEKR/rkjytjhLQsDbwLKSCxzS0HmZeyOOPlFKNK8fFAWCk/7xIWCs3cls04d+IZYP8fqOBG0L0
8DZiwGNqvbHEYCMbbZQ4uUK7eIJYorodhqkfrlz/RO1a9hr/8+xGC8RPru4Qwo6l2NVJ1qOVSxQ7
TFP3h8+XKdqGGugTucqS7SaHMKjvD/IJcZ2+w+mRjZ3p+hcr8DbaAdv48mu9Hi9tFTUp+AhuhYqF
g5yYjdUUR+WbP0+Jl6xF8ydUa77QaoV+U3Kczfhil+qxcVlY//9Ac3nWmO2b8uE7Xn9dkHROd++X
a1qW0BmZGCr6eq4Q0IZqutJ2P7jqyZ+/BfmiXCOxQ4MhnZ3RXrCTUADCScH4r9ZNiNVldQdiUftI
ibMg8Ea/cKhUBcRzZ07It+H7Q3vDFC+dPqxF5TxrFbz1E0Gdc8+SnYZ7/q47T1M2jxYhfO8y2Cjb
suUxPQX9a9dUY8HHaiWcYefsRhDhFseU/Ei94cHLdecqD5qTBnXvYiVSXyUuRvVdMV8zHwqpk3EF
bUHJCoyRlaIGsotM7oXmbpgfb6ODHe4nN8UffXL2pGCRzEbTiijkQCUZHE3Eabzx3G0/jXWV2Kfl
vO0XaLP+KYFmFIlS5NwOWxkB8e136FSUZ5ypwMJnrjZbc1qsl1qAFsUSU+E6haJa8fUP9j4qvHLe
+5LARb6E1O4igT0eLPZK1NJlKkxjLBc9RSGiy7loJx+M6L6Yjl+5PXK/+6hWYFkhSHWUoNBbxLmD
lVCOaEjUtlNATolAfdVOiQkw44ZpN7lWUsHXJCXgd0kcFKvVjacp/cBUr61ZGc3lnp/jJtJtpq/Y
kQJDeifXlrARYpN5/ehTNRY1YklR08Q7pEfuGZlXTRKM0ej6bm3QUtnmf97g5oxNZxJDXItPdbYL
LmpZbiFYt5rjBgFFy25QhE820ORVydBYRO5pTky5Of06xMD0P3xkPkl+g5DDcoc0l4hF043TglHM
RTCJ+QPWckBRYYSCUnLcWHpDrTR49PWGyQt158oHnGYXJV/DTdeL+/8l+qZ7zqKx7DP2R7WJNJeV
qV/0SxxottbP0Li+cvbeYm/nGRrRPGPtftHY0V8kH5y/n1JMvwLR4LQ0IjTnXgxGuy6CJjKLLCbZ
dElKP3ymG98TnrMOBPpllDXKSeR9O5sHycdqavNLHrLc6H81gLo5z+z/Wngl40Kv4LljZRyaFfrO
gtVAccw6WGkaupcv/8ZKxF2kPZq3/J5kioNwV7Afqfd+NqHxlj0qbLOPtItEw9D2xtC8EECOFlfx
1gmitvECDTqnQa3dSaR4poD66DoQuNrlpifEfhzzFjXNmh6w23R6KKP9q6oCUsj1QfRTY9jeOEO/
50DutLnUVSbYlDurxteHEN0YGx6Nn2qG05VCNPxSUC0BEDcxU1WRtRp43F4Df8cee5xNKqftntlx
0l+7WrvbIc784/ovI5uyWToMjhQTIu/pNoRwPP/8f/gnuY/wkugCLTD9Ea9K3fwO/zkmu6Y4Lith
drx12wyjv6po0zmAZwWSw2cpF4KHlLunTQxA9+qO3m6FScT4yTTmFJ98ZwjPgr+pO25awdoX0de3
MUK4eSgj6/hADseCFZeHULCnYO25z6K7SQVK7+v2bZ5gDJdZ0acbRAXuj2H9B+ARpHrTdCgalrrQ
osU45IoBNKx0qLkrpCrZOTtm3vCXZiIEJTPLhJGxNyOySndIIvfnUH3oMxXM3Q0BR5S9MSJYmjw0
+H4JCi06vcAxkczy1WZXmWmKeS1M9dL7klb/HSbhDDAw2H3lwjCJz3LHdSNtP1wbRoyqZXVnUzZA
UEIj3/fH2zvpdjil/k5f9XXpL2xuOioob5CMNbeFRsyEhkvPJh0zITnleVNKbW1K7reFbrgMYeye
5vULlOmnP5a7rqYQgH81/r8tjIuyN+wC+cTxH1ezTpyO+GbvwdZ6zXCYxBcbuTT2Wn3uYhMlmPZy
oVovsaku+nVLSWsFhLvnYBU6ko7pk4pSy+/Ov8EO0yYeWfL9GqHeIfd+hwEgtZlLvKZQQvUG1jYy
rRTg8VM/tza6afN74UNsQjn2YqmRfvg20odBYNQFNzI2L/LcKD/ldJ798p3Va7GZl6xxKljjPVDm
6+iewntYsB08eR2P00KRCygnLJ9BYLYLw/j/mc9WLq2b4zAY3Po9SKZReL8fraz3esb2Yr/LoUZn
7GJHtie8TaBkI9rMl2HMF9GnT5aeRDRyONp55iIAssHd/JR4nuZ5HuIiaOyrg8xtmtTWG2FlurIc
jWSljJxaz1t+9JB+uGipwQVfYbVavG+ONGsf4+aWm04tWhNuIvGCEBVPglzQ820YcuIFVcZ0KT1b
Ud2WomFoJxN1AfGFqo/Wq9r3fzwz1OLMrPA3vLQt+/gO813RvxJMhfTedOTJLVfRk0HFLlRWX+eC
xsK22kN226GX//CSxvPlN29MHOhzRwxjKXkQ+NmQpygaJXwSFUUtcokM5q08s6Bi5mH6AR4tTl2A
fv8s1+KKAmpAm4t9AyoukNMjRoaLJjivanUqTFwHkrrQz/H6wp7/x83QTBUVvUQIems/EBAD565i
wIDHM/7ZIZDXqqju6B9uGdMphUv+12mGYvBZ6KWNQHlE+tuekkiSa3cypopUeK92/ifzaz/B15h6
po78NzmKR2Er/nWrqNUaJ0ctRvgN8plMT5d2stBweekIaf6jBGEl9ePbwCrV7UlBEPzhexJNdWBC
09Cxnpyq+rtQPazMKwsrMwaB8LUjMEwEGzbKBRTN3bZaeRn79+/adTanH9XcJoBJr4VjRsxuTEaT
HWyr5As2QhwE142R7FOkZphmUJG1BJE7GaKiOYsgKIcWWYZzPNr8rpzYqUSK1J0KmXC1yDvUFD1l
ukfqBQBWOQWOOU6rx+ouA7CyH7vejSBENYi92nKYriMWT8uWJHoQgf22FIDUNugS8XIFHjVMOrps
yVBqc27uov3P9MwGJx3kP03CBdDxfSTwZBEDtJ1rUcBTornbpd+OkGe0ADT1x3cqZFFWVufh8Vuf
tQHtvShxK43k3YEsFLF2ZTNQjrxt+8XmD3wssNbPk9zLK/h1GDkzZd29b8Mt2AeyWl5yByNJGZD7
5lKBzXfh68+bsexDwAz7IrC+l4eams2ypBfkhOzAKrL5JISAzy13u97j2koeay+hHFtYVmC0ftzC
L3u0NYqH8b3nPvnSeIxaBBADRvBqdMgtbs1ybnSdedTt8tSEvfTbceHtZXwC1Ge7umnxbY+GcCIK
ezVULxoDLsHKHmF8Srt1FFer4P0YuZsEVB+QevmUNniQsUQdMIGa5Cj7BwU9UIsWWgb2dOGMl50N
5LfFllJb/ZVuHUeUfgvfGH5Tm8Ep50ysF1qvD458McxmouRaNjVf36Ldm5DUQQAuVaXJn0xZi6Aq
D656ZLihBkLx8qWmQaYDdqXK+fExpu0dbPOO2LZCobFyPBMe1LHrRVBYwZ9jpG3NVEXAtSA5FyK3
v0G+mK3MqCVcx+1ONizLXy0lkcXJBsZkBSYfSPaMkyeD9YCaygMlGbIUgxcWwHAPj4L3hCASO3Fn
NaQxQVx6FG82KA0cbZoETjOOk5xt5501QnfhUowEEcVIc/S7iOevIM669Rn0pagi5CWsG0jYA+tr
XHzissNXs5DBs0EB7tHDRLC36cuCUiAPMNCTVr1KVROpXsPkL2y1zIi3mnHIJnuDwqpd8MnJPhQz
eBViWQcuhsKyyN+aGGaz7pnBsrCLFbbgJdo8MuAqFogH0VU0Jgn5LimLWOmvTZOgknxZY16eWDFG
ZvdQ+4y/HYnvWfIIfPvzdHn6mXRqk0k4aPYNqok5QfVsUSzVG3NXpLXNXN10KKQpQBabVriyKwD9
JyEf/FF4lQZ5QqaYsurHDTVItqdN4XiLdRgE0LIEPRbtS5DfzH6HWGNgYm7qPnTY1MJmLbNfGtib
y47nHVombzVAlAmaSKT4UBeYuLdn+b8b8hIGWodZLEuMm1/1WeZkE73Yuodya26iPOmgvW23T7M7
u2P/A6czBNcLuYKWyWOKyh3JiLLOZMNj96OTpyDiPKYVgwFVW+WOjL3yjTJEc0sjo1WMAkFkz06B
Wj5celH7iNixQYad+e0ehSxdFXr2l7rqhePwhK+gIcRjF+8qKA4nHbiELK0KVoGMFP4S7gv+sa5A
gZKmkTWN6KikU1dy+x+ULAw5T1ypx3CM94C9ZRFyjCUlmTE7ght3w8aE+Em+Takp6/5VgomkMAYt
+/2QpKSIZQA/moq1PY24+S0oKFtg1mz0iN44yLj1l6wlU/AsUSiw32aPBOaOrQ7g9/Pbov1iHhk8
lvSnacf45bk+B3s54NTU89D9kyGg/Ba3P91O+JPeEYQtGutK33UtogHoAbRc42l1cTPvtAeb4JuG
HTsq3nq+kgnKjg8b13+wdiIZKIbor6YBQnvMFt1Cge355uRhueB+XTi6xLLPUWgdIhfLh21xwmNv
UMaWqjFrQuhsCb8xrnP7T753BfhmAUC6agAfP8cb2OlVNO+lO2+b4jnYA/IEoUgbQx1kw+47924K
Ve/MLlQYNZcwipRS0q7Eq202xwjd7tP/37CzFDuUCtFf4wsevDVWxvoAkhPHXMhC+n39XG+THzdc
Rcm5AL3kYy4NaKXBvmF6Eis1mzaNHAmzn53osqEldkH54QJmwwm8U+m8MDy64tHAyyWRKI14RAxF
VBRNw9MY1DM6uuMWU0D1fiIioMKZfFhM7uxeDEqpT9i3xyijMUIki0f1qtBiYQE15g4MYc6l0Y+1
U8Oc4UQ9n6FARq25ZZ/2PfaSiq2PTcGMUP2ESqJ5cziZFzKpgbHlOGcu9GyKuxSh6DX/6QchEHF8
bzPDGQpWSssqmsBI9kgmrzXc0AfiILSY6c70SJB5lzILhxA5A3d/2L/xESNxAY+PoWx/wi64cr3j
4Z/wq40Xj7h6fP1haudofVNcFcT/i5HBE5N3oeyEWZkATP1ovMSonIWhMG83PFPeNjROVlmStIng
8xNqW6t5Ri0TGHf5bVUJEZPXcWGIlXjXvNEYaRrwRotSCX/fpujK0b7InnTXPK1kCDx1ngiuXijC
p4Hx3PsiP+kh04H6xmeSMj0vuQW0IxjBtxZYD5MH/9pr/aPIg2Av3sBFQ66PVCgqy3X15bRtv/uf
qUiBXo+yW0tZCYzH+V70IF180MbrbLfA+RYnL/ft5XvFdTZlK5R4FHpKQdrZFKDNJ9ilFVcjo46v
EfrNq8k3nPo208xpJMRDoEWImTLFhfUhhsFpgDmzy7g1Mxkb40Uq/PdeEwbK7GaLX4zsOCtMg3l5
sEA6c2dPr2EsIvQxQdLWp9zenT7/tC0xc9G+BkiHzYmWLwgwbNclxB1R6tm28qa1n8fF0hdPDlC3
uMsPx+a2P4ZuWSBRuR7OJYUF70PAICNQaP5Tge9PGc/1LsTH0ntTKzQ1gJOipL8fdYn0bl6H1SSR
pQy3fDM5TwLRVP/ZvDvVXR3IMqQYTMZUeVl6M2Wdp1tFQ8JXi7utAAsvvN+qGb+gUC1dIZM3bdHl
dEd8HOpBDMkQejh7lLtJWVf61BIbKQxFNHBQnZXGwHIY5qzixdOno2eMJEKd+ACfoiDeU+bT4DLk
0tTO8mc+2+eUGBJdTTfQAhQxCzDw4a7c2yjSC4iB+23FXmP7TdDpGyolyDObYlJycH/92sVB7yi1
fxjRNgyHrcYI8WgfS5soXGtMCAX5fi4EL5WOCHyIequ2KLnYwj80I9srFWAxz0rthSQg9Qnw7o/H
/A5WCVvbOpJzpzWAtVOSXG9aSjK8a/LcbDTmVvK4GuKn50SSsqlTh0LEyoexR0om/EwnW4jzWt9X
kRU0ZiYPYbhzZOwrLIRF9wW3sPxcrI9w7LLn8VbBuin0pi/e6X1LHDaAEW/vszVzSBt2nG1eCOos
MIUQtbSU/L1jM/MJCk7DdANeURlW/rF7c/af9IDXThGQJN5veFgS+wsSJMrbHWt8jTM4yEHZAccj
gKaLgxUE3xdc5Bm2+6er/qr43m46Fsy9r/LkjVcK4+ak0eOb1cOAlWb5NraOuQjsY9wx2/dFHNWq
fzFW0rTJaA2PtWb+MLlABoLROzU3EX1mqkxVycMRzeSDBFuV8QrTVbGbivrmiBo4uMK7k+dSDcAn
tV9zV21MuwbaZHtWs0YQwQDRBcswgl+VtVBoqKmtHfV/2YBCCMtxkisqeFNrZ6Wy3h+PEVS06EHr
Tscwor6wfkuVGxfgIPlvuplUf9kAxQFq6SgZCF82tWBrNhveDO+W0y8Wpir5FYVsTqjLj3k6d1kE
yauN2daVkS3wgfAdAkiIxE6yC39WlU/Lilia8UwuGssGR2Y9pA1dOc7kEV3PdSnvBtg5OiGPtPjh
5gqtWAmCXOICi59qHD52YAdksYstfQXHZV+poR7/k0jM/Q5+3t8ceJafjPWhE6CV3V5DzqYJ5wSo
720wyLS+F6Ilc1EkdHA5t99sqMYjVwf24OWNcggELASQ4d14Mc1FuKdKQe2C9xiHlzLKYgQrcT6J
bcBcFD4vbwUuEpZmVXBsiYxtvEluwVE2k4hHfZ7KzJu3vZKxur9An0LhCR4aOrm2BDigSSedmDFo
uwbcuiWcSJRg49A7IiYBBhHLG80uzKtHTTsaQzAoEe/CQz3TFacc0siyB8/Wh+I8qOm6iBipW1OP
Y9lB8DD/WCuOUz2YAABVZvaybLIxvLLSDyOPKDo68ScQdYFXBIwGlwgFJ1mpO9hkU/yfVE0DO1ha
CEgnhl9jBofNlZMB/jtqPRGHUuK2Lh+Bjx0vy1cE5dAsfigPQzsHydDYzF1srfxxOJ32FBikR3/l
L2OQtAm6B2AZU2eOJJDjuN0VdOFhKcgLergnnyg2xtTynMJMAT93dQtfPemsxwl9ksQLDXbY1etc
0rumKrLpA1rKGLA6X0WgnmMuyuBXleyuBp2O73vpam03hUb/iBzulUXI3WG3ObbwWb+fwnuHDeLK
UWYq4jJrU2M0Ea4ZwpxxahAT8AOvYSb8eBePW86RzwLNO0GBqJvazQ6LMULjVtK3m33ndvE5IR2y
iRhmFcCqIC8Iv3RHkWIJ4xvtgQwMv7135VuXcfYzGXBvzgK1pgcLqLlu6UxTDgXiBFypO5riXUC9
Jwu/t+9DkxRSAQHSHge8yjt2brCeu2iN5aNxdtBnGYmj8nIbTnD/eXezxGoqg3NAk9QE5+X/mGV/
6m9q/hn6XTXw38B+0V9BOywldsyeTpW3RCr6vP/eFIdvacZ+vr3lS4JL0/1WDwkKEnqX/xJnVPCy
RkSn9nfv/VDP1QWdkleyfm/lu3muM4F8Le5EPunou2MBC2mmDyP7RGarN87+kRXP0PgdG4paDk49
DxPZUzFTD4w+2u5J4I9kezpsnjmM0X6FaDw7PQaGyaQyrTF4FROG8HbejJXJ4sLMVePx1MPIGVyh
/W2FqY5lUZoJQAx0Jyq9ip9+st1vLyg/BeNl9jcl9H0nJBvA+8EGleUyHxZzwsQOHShYVmSv99/v
thLf2dUDWML3plY0zG0V52O0RvQWioX2TTeUsckFnWniYW3pRXAv/vyxyZgEE21JvFZqqm1vubFX
zrztQT8uYFkPe6dkrTrx+cEWNC+bKvgsoYX93lLV+6CiZ8IK4z9b/jpNk6F7sTb56GYG9rhkVqUA
LjSzb8LwvoO/ce7l0L4spo/xi9mg00/UaGxNOQlhMFeXy5h3FOlLvZ5OupdvrS8UXtrfowOtxx/2
s+okM9cjfEMknXr90oUST02wbEYuwn9OTW6qamAJpYbU8D6JmP7utZXc40fS7URVmJOIzsYlu4ge
9Uo+1A1GQHsaKNOBOxFbLYvmZYDuMmHEuixIdV+2ECKwpfanBDgYSK3D2ovaXPoSUJmz3a78nhGm
xCwIL2uI3q0O626NZnNsRLuGlb2HV7t8/qnopPm7Ohs8g2UVNx4pBjE+rEABNivtLSjm+V8hA2Ms
9NsPZWgsJ7FlIJXu0I4iAlpr7ovKBI5yG5VyryCiC9cXhnZAB/fy0jZH5LyTVqaCDsdrsAj+d+19
M0CKFSX3wY3BnY6gSB3Vvmn+WNEd6C8tR77hAFOe1P4IKZ8E7k9tZ2NA57K0Ev0R4MPVXff/N/+Q
MVnBHzqbJN88d5Y0gVe8MMsAb9+5kuRybjLpPtAgswGe0MHKGs6FDCocWharJ3IS2QRKA4jcb8KL
XbUqcdxTUTBif1lKaBkZB4Ld62kjHjiVgsZHG8WOO9o21Db3vGZIfQk2H6KaFYlkPJA4dRZYUYU8
3/bRAU9jHvLSaL4jZSBSR6qQuffNQTDT6G8LqokIfLQMsbDuN5aUpYJuZXkSNY2w1vBN2Ueenbwa
B0jbEvmolCLcI6/zau/MzrJ6c8ykS9S9GZ35Jf48cr2vY5CEBZA3/wRCsKeWWDnLW2ss7sY72zbr
VS6HXdPXf7tohP/xiv5dK1KEFERByjIkNSuiYM7snerswJVlTMYF7ISxzdTcDWHXiF+DXWcxEw6Y
R610lTZn9Ff1/PcuN+lGTW49wo0dWHI0oKI6m+oCmDuUJMDfXQ3faIZSsMI+/9Gx5UnoAipVLrbM
Nkn4TFE7R6360l9jW8hLD6TiimUnQI8gY3TA6N4xfU8jd5KFWBtOXJvFx4NLs9+UBuVNAyitXNXn
H7n1qbTqJtPU2MjZS8Fre4uBEM7YXsDfjQMNed1uASXncMBzmFVgcC2Tx/Q76ZaRQ8ZNNw3Ged7T
RHRcZx0eBxSqu8Vdme9tuPjuSzfPhMRogtu6S5QMYvc1smCxjMAYzQgqPECtBShFZmtIObTpPqVu
GhXJkJoemKnkXEYZmEbdkV1soNsCwFw8s3NLJG3LS83qaAVWy3smEjRXQJLfpie6mV4Lhasi8s7m
th3ohJcVJiQl9FPIYiTbPwnADZZKbjuPgTlf954mJzVK9GnxMuYPLlqmdfUQrIlj/3PzTvqRu+es
qqbUX0qXpT3FpoKkds0F10O3uR1DGpbkVkma3IQF7XqW1qN4kN4qii9WsXIi6XJnX+UUEGWcDAUe
ieGO+QCDr2tHuLuRddQLCSnbbKMbqcsgSZNgxKfqfjxd4/U0DWXFHviQwEsJYljenx7Us4tHAXFs
58n7ZmVyLbn9VS3NRMW1ar3jRz6kiGnSJYK8Q8x/+go1D+XKZPYwuibXF27tocuhXESjROYK2Bds
6CUDGOgLQDVS16b7myikLE165WZKPCoVMMmaqxF8PavobzYruR14+s9eQ4S0Y9LtzJSULtUMdno7
iA4WgAWk+kjwCUKKjQGygRdPumekW3R9dqtDlJTWH/3OJeyBK5HyPvOrvIOLWOcGElNq4ZyW4OCF
YuK71vYnswIXA2ZcmA3+J//n7Nz51etHG/OVfV9sdgh9FBieVNfoNAD6EUDWmJuq1gj+ZECNflQ7
fK4lsxb3qMUXTXYr3bxwdFLZcw7pK064nKk6RecD6SDFy4P8TlMPl+KrjlvT5BAVEDSLWJoAVktV
eCoGDgqwIqcUHQDTltpBlLrvO7RAo2mRNukw0nbA535glcT86RSZkhJVjiKGGqalINXGP9cJbmPD
QH7irZoOsbviRgpR71HGK5KwaqUaSs4LNYO11QyhWiM5HR1nET32FJezl0SnAV+9tKvcFU1va9O2
Xf9LP2opDyPSKuNsuPW2KnfceF8DrCwWJpj9HI1wNV20iFDhxysckLA4kWXMCIaIzYN6m1bv5vbA
CGhKELVgZlX/20endDKqb7jXWPjKN5Az5GRalcI73990RI2i4yLo0bS18Uyn/bU+FTcESHkjqim3
mspdIn+k2vDypPRm7KW771Ig2QKGdi9afFEKyeUVDLtIzz3a/iza73+KFFvKMFD58/SiEyKuH9NC
mOZZO4qdHtRNYHjkYlBEJydWvQt+NXbNebrrdou9oO/qDoIzWhR57pQBgxb7+TW8Hy1e9Cq79kic
TJCYYnQCDeZhoTUQVQ0x0FBy4NiQ7YCIp+9Pk8lnT3Zx8iQF6DOlpzv6MtWRlj3DAxCpOKdeZWit
5ju0namenZJ3KC6FfSMLuTHbUn3JKXvT2eS59ZJUdKs0ae7TaIyL529+cOwDAp/QkZtbA+FwZhy7
7b+ndyuJpTZLn1yLMAgsTNStkBibUaTzrWDJdtXYaRdXwxcxGtubj0WdJzGdpebL0ZBJKCCLrtE0
WmuwldN+PBDy2cVeM7uwG32J0HHGbUhDFnEVXEHtgPCVH+NcsK3Ha8DBDsbLQAU7LF25ujaokZDr
1EAJZ2BEBKziZL2UdZV0LJQX81+/RfeSvfFdfRdAJ2/a/71yq8WqFEgESDgVleOVI4UH3JWWVyu4
1nfLoekKQbqGTzM2//EiP7v75Ts4+j97xxmVX/Fc/Jc4ESYaoaJ8X1gJXnFWyTFucrOUk+cNsVdX
BXoDA+Ks7Mc4J7Rs/llyctVV9mZ/5gph+T4mE28S/VrCTJ+fsZNdOv2dBhPVClEZYPtQfGP/fm/8
1LxWBPdE72T1FLrJhzfLthdppxhlexS2+eFCnPv46R1tZMktCktG9g14UGsERM96Dtr3B/j/o+6p
4GULZphKFq0vDLfnqhRKoiUkRQEI+pnaWou5QpnGpZPE0YQ3Jm/cIgG+UjaTt0Ffq388Kqoiqnvs
FspZMu4Ex43lMlsFKsali5WZIJH3Z2OzNRsb0TpUbXW+dlWSBRJ4hdTreHQcWSJ8b1r4cR92+P7y
8IucJOkcUsTYcVWTbhf6E/4unUHYJqPbVldWnEo+MoHtyP16wPySXAeSwhnD+gaUBerK/jnnL2+C
Tv/NG23bGmGqbARrhNBuUwIbk8immr0PebQM5aPLM913a6ls1ArSFcYKwpyvF7bLyFRl9uDRmaf+
sEUScx/y9mqiigmMC/JH8M/a3pjeJD7y3g5Zr/WYa25OuSYOi3CBEU/o3ioOuDWRTjUArZoV4Q3k
Q9iMkqnyiyjsA61o7DKD2pze3KKcTfRYxNIk+wNiO88wrc43UYj+mdu2Zu8SO+MrkE2HSfg7RTTU
l5osbOz3o9U/KmGDj3kkvhr4HM+BRZqzU1Xoqsng4bztNgGSEOaynVk6M/1Gg3ZemZwy9m0RUL81
OWHGXTSqrTWVrkud+hpSfL0xXcqMESPuBYGwDxaQuoZ8+AAKiRQQutTJFcH4cjp8l9S+XgK9a7hq
3AcB5KDZQVtVErWjm5UXhO4qx5uy9Cl/kex83LFAL3xHAqNJ/yQasQHi/0OeBC1PonaeA/hsrmu9
jEae0o19qYatQ8EpDiNbmoU69eOqz+NXQu2KWFTIW3eKN6I+6J+ZHwbm2mqNRt6L4oem655uh405
k4JKNhHYMrKZ8LgqxoSRwdPxZ+dFL5lfUHgvxPo6RAK84jWIwtJxOAuzCOfYmIY7Rv8M+LmJxzRF
NsHxvhadQwtbRRNxaU66jePyjSr+RYMJYyoON8H5jsTGnao+eAbYv7bRZP+5Iv3bhhmBFprXXShe
Ywet5MFodYBvOXkR3sVz9HSWWjatW1+MLzj9hf1e8HzlTxuoecfjAVl3R4u4jfdkxPtj7EWLOD7O
WnCrXKG0yKjK3f4TlZjirdyk/8Sa5wR4rurqTP40inMcNSD08FtqXNmYMyDCZCE5PbYXL73OxuM9
CEeiffY5KF/LqMV6hmKKbUmIbTMW9geR1eZzYmi3KV3XkCParqy0ISmdKvcc0Hsv3aEqEQYnS6ge
WyidLBBv4aF67Pb3wlU20XJmoqbrASFhZS8GMlIRaiAsyIV5H04ekHZ3bE1y2drRBYOnHGH6XAjw
ROYofh73mZf+roSVLrQ8trzMXQ8/1k4uXX98M7Qt9+/6wAbVZFmi4eAtmFmujGxesEXeHzTHOBfL
ueG8Z81YuqTu8qRsJZSLkcsfwP6USMNCHZS77hfkQxzVADaHBJWdrp2Np6JZAyUjR4vLdeXdmka2
Q4Jcr+ePwJREtmiDIwDcSf//5wirBMP6Wpnh+Jirbz3nV/XHUHD50HyRi8bJ+VZ0FTfYE07PeLZf
D2zBDDwLCX+S0+QUg3TyTFYLjeYH0vmWdGq95qKkxHscLtqCyreSOW53aabaULiY+ljgir2LJaR7
ts9oSxYO2v4zUFu49tGBCmXT7pzVwxpgZM/C5eWLWhODUo1bi+puEdECMb7SSmoDY6YMzh2mgMDH
TFJI9wpejGki3BzAED/xhLi7XMRveF/VzbctJHylbIj/8CtD0tqFXSEmC3utE/7zU9H79rc1MpOn
7ksaC5iFOJPyJbAYP6WDeMLrAHeZbuYZ+GfJ79P+eBvQcSY+NzVv8gDlQM17UZm93MVSX9FgLW3g
Vn8uR+gRCBpow0oOnaE94RdOPEu8XtGCyP3N8mB6j1XCFiox0yJ+dQ0dGsTyBJnP5I5DTZIAYEoQ
6P9G4mbGjVWhUYQfnj2j4MKjnFQhdD7yyn0H9DTbcUDplp3Fyqc4iq5epMM45wKWhD2x902PuZkj
reZJ55gqNPsOOwBx+zDDn0FOhN9JHdQ7QbGDOQGSbznuIa1677XOA4AxaKVl0qDpZQITux60aG/6
Q8P7rgQ/HV5Xqh0Re43nsYK18ORIZk6BDSL2oeywmj/cz0dn18hcu37xWd2/81/HwKRHFq2VjeQk
EdTrcIlyO1+5WBIZCygX38O9nODuhJtEBBOBT0jf+4AWU5v3SeUOJbrujVJT07vViawuR+yNBUSF
z8D2/mfGOMELDcXuwbY6z9uVnJcFhRxeqVKIkYBe7X+hUbfGJB5rKkntWKbNaaIGNshyIvmKhUf9
BeJueHOKvzQTro1nWUGRb1Z2dTs32TrQVlQYhUycbeWVcrcyqcvH1noj3TPu7pMFrUvNzOU4M/s1
F9uadk4a3jtYwxFwf7v0mEF12oUryFSd9iemw10s/92kVCbO5bOqo8YL+f3gTAGpdB80k+s/jbty
vVUTVmA/UVfzr5WDlegnXp4/Nlb0IuXomsv3aisoCmljsbCVAIDi5nIliMSOID+iq5tKUHivAhpm
gEAdXRzMu3NLOW/oJc5l0KAZDlCCsBKUVIFAngNzfZJnsMjF/MYMn5LpUh+VsyiAdy5QyuB+ozuL
NQaVx8Miu9ZratLGyrznxro0FFOTfzqorwWFIz/x6GvEdhOoK02iT30LxbGqVcCe64v1Rtzsitn8
UKx+EiV7vUn81BsiKKde6gjFFORdsFuoD1bceZjHt36gMgVaIn3ghZP0DCx9yrA+VUqacZ8r+qE4
AFIeZZcVbKZDzoRJ+LtcGMKJoMqqwKm1FAQekCtwvM05SGa2ecCV7GmRDhsHAjDSx787m8ydQm3f
aLnF1dBFRoOlQWDb/TiMjzWt4dn/WSxs8Vi1IYk4c/RwOI2RVp2iVAXqAWCuC4ArVW27mikAn/IT
IzHDPc+Kc9SXyuBgggl7cDrAYlzCffjdQIllnwYei4V78tZQ6i4IVOmS7IPYl27NCNZh4OcDRqgK
HFw+vdSQcm2CMSTwgOuKv6RUSvnjh8eoxLby2Ky76IMKKLpVC/q4KbRnkcT+0gCBqL6G34eA0D8f
TUTuYlEDT6gBBFhEzU2rXIlavGmKRTwlHkzzoxNnLos5l4Gpg6Qb2ducne/3Q7ZIVVYpnAQDewLo
54snCfGXidKmf7HAWjhlkWeXDue2kLy+Q5z8M+ePbHKyVykAHTxVkz/c9BHmemjSFUgUWTjOrlJP
vRA2l9Dq/jO+lLb9uuKKIHBpld41WGJsewF+6nGO4OwFxX7zOeZSC6UDrwPtflkcbFXAbZ22RrS4
b4D5mhLZ1+9zfBmBgt+iX02skd4/Y+x3f5MIMCCJcbtMYo9VeyNdOFSP8Q3BMrLDGAc+d5jWBHta
wbDX+N4edUGoiNDN8AIoLDO1mJpZeHAR1qX9PJ8qQUBSuuZ0TS+2EtCC5VxxAd+MYTJbBpYvk0wc
CAhpfWFhNQyKYF4NFQnJZuLpvcIR/vPRGanw5HJDgnb4b2bd7KVgrNEd5kE2EU3za2C7xQ8j471h
uuciENPL7iD1OWAZr+c9ZOf//6LSbV1Q6aRVf09u+MmsxYkGJh1Jqcyfa5qXqAG1t0DrH9bTO6ll
n3bFZs3YD7Yqx5lGAe66bfMZYFszEl/u3vama68hf9rRnz94TJzYT8dSznFv1PNBwtxMI8/zL7Ei
b1dwfx0DLYBQ0tdCXRvAbEUZ0GBnuDCRzWI/Ox3VNP0X+cF2ifZO7wYEMzb5gRSUUOapVy38bHU7
SVIhzKkzqPbdfA/2nWDsvD6Llx7FfTiorRnoPqQdaT9lOtAjg4sFZb01RpBVy1Lx+e8KkEYVNnGB
DVHqKyU3eaMnMyU6PnglFmRWaqXnrdVyyD6d7Mzk9SqHJdcFAOmz6hizxshLNDzRRthLTmrUeBMw
JJLM33v3DmCns7z93AKkGw3rsX+dCRQYS6iU9jCseHSkA9MlwgXuh8DK0KTU10jt9JzyS1xnDjN4
7eAzaVsRS1XPcIgF3wj+SXs3qfPec2IzTZtWfxZ0YaMA5lyfO+qcdBWQtLabEd2Eq5rKwbpLDib9
0UgSe3n5yXJkp2yVs15n2EuAFA8iB5c2IHsVK8Q5tG3PyXVFrgo3IMQubodv2VX9SpZb9OjxnJEQ
io0zTWVi4rwtGFdklKdgd9JJ8O/8hcIa/qvdE81LdMxU1QOM0fJMC3ZPLW7Abxh5VWkVFvEvdeKe
nq8PWZrI5b1ZbFarGXYuK23kgtdJZVNGV5tuMbosotzTEsqYdQ/D5d/Imr5puqUK1xtQzHFcG5aN
HNgCn1ATWdctgHaGx/1ivEME5IHVbRDqe4ETM7fjiazBNp3Ci0glETbL9I1mnKqN+pl8bjDt+jLt
9xGdoJ+7fcFVb4P1eZj5lAOHJ7n5rXCp2xPMT63JE7yooPKouRi/abl4UV4LiL4e8Cfih4Sa9+XS
1jI03Gk1nnGj7bcGoHhUeTqYg+U4natI0pXsS1zJpaarhhp/tdR58CWGjPLLZDNJyPXcTR0+9KOG
3Wyij7+iYx2wrvMVsp138FrSJd5zWtUV9L8KyAWjIDOIA8zgq+kBgOpko0PBqd8DhPX1e4GLIZzs
3+byIivM92Vdqy+locW+h3Ux3otEHGqpXK+HZZrjdeejvzMS16qmWJfJOuOu+BD9mMWxBiewvmcj
a/Hn5mf3PrYykMT5ihFeY42hB6wtL5EVf9VW5cykR2jOMmYsWFcU4eUoAhX2zGMCQL6YMYuAhbzF
qLRMgQ4acIM9qb+b6A5b5XbqNxizDjMbUYSJE+9pVFO/K+pWAo7oArp0x6Caj3Qe6gQnAQLYT/9r
Wyg9ohlweSODG+KVw8j9yswMaF4Trtm0vPFnLFOoiOAa9FQDyDCqINkdWzCrY1MihjWn6cL9O8h2
xb5qlcnH/BVq0ubaUdO37P3yVwH9zUQzstF+iCamOhuhFdt9jDrrTXqzZ6rm17sVMG+2pi4OK6Et
vXt2jfDw41CS56CHiKK0lQn/9qHG9eLXsrFf17iJpkeWDKV4c/JqN2st8JFDrj5TefKVyjXqtItx
5wSK9YYYRahRF+ewRvsl5beQGjBMLOR3VNI95ZnVhl6e9wtoimSV6HsJEyzQlfBBvMdK9I+DFioA
y7iJYef/xiqZLUB32mt6MSh4IPMpoBHKArJozg2DXBorJLXcYZT+dhfbmLC66o4VbpHCMPzquewe
nUlnmsSKoQ86SfFZLXmT4rQkuVSeZE3w5Qj0uIei8aJM+WBuPdPlVzCrik7TGlb4cZQcx3UK7zZa
0prdEGCyQwTdpXNBHLmZ437hB8l4lnvYogyumZ5fKvKbnnCZU6zj3kq4//LCmjK8EF6VA/xZ3vA0
7P0k0xd/OS8FFHPJ40QKGnaBt0Goelut19zV3GOcKNLBesfQ0Fr0TRF0I+EmfvYSvITtu7CPFtPJ
aR++Ewwc7S5IqC/l1UfmLK14DMe1E2TCHQr1nZMHFO+PJ6tKgs0Psakot5fvP0mD+tvinZfpUn/2
b/e1QWRBmtTkzOBzxGLFlt6ZBRkTg7M+norJ72kohxhHy9Vs4xDCICB/xLne9Np1iC41IvTcw8ix
gE7hQ7YEA7fULAnOeYW949xNqjHXzQUGRY//IU3dw+paKm3KdIzvAbaCKNhjM4384kpfzIYDqpzW
kt9C+wdIw1a0KfrIRTqtH7vid4rBomhlE8YF4k5X3cWDp0P5hwnTptq4sc6EUhpOfdEmQ0rFwQ5n
inNL4aNqkB6TpJd8B5sl25MTei7bBZolzkvtLsLawcadGSHS0ddNYilmAwM/EgTWFBlx7squ07i7
nz8bEMTn0bU+5wkOXAqCiHIA6d/Ha0vHpSoBISEFWtVucANivzE1Nyfp69fciBVMAnv5kNAmMUSF
iInb2WXCi9jDnWrigs4A8trST50sW9Yir+RAQAAVvfjsp1JsPdUYOWeIjxfPeoJ43rIm12l9pY/x
Bif1kmwctNt8YBZHuNmQtYVhvmNo6ClYvOmqan2HMQROX3wNXd8D5HPz049vp5NHUYJmHZjbufkc
oTm3LyLSgW9psx4N5iPO+zGGqbIw/d4312X/Qhhm4x7FfzmOz4k5kEk7QDqI/jSkXsfNU+vAstLY
jTwjGy+Cyaoox/Aelc2b8LAP9ALqYI9m9e1iY7bmZpXMJ2Al+XMApD0X8+/2MQbsbjSGSyOTtMj2
h6PMv685uHbyPV1nGjCLE63U4H4ZnOAfOEwcE1Jj9eM/mQxlcypzm7MHhak2D+qXqyVsRcEJUW7g
iigdSTAt4O+tE+wugrdgf60ujXa3G4L7sUnMF4t6kfrY/mtAd9OgGKbbfkdb4bcBeBZu6s9PsQy9
nGd/XH2lA+MoXza9IX8dxDw02OiOhcPwGjIj6xPPcWzI9hu491u4CwQD8H8sl0gtIpXHJnPGB5+l
eATCiRZ6HrXignHV4V1YKbx4K511e8q44h0t2Y4OQ7tzR9xDXchihHVE2m+whZq+GFlRIg3G8O7Y
3NQuksOOSzu4xlEe46GIo+j6HGYXnrrSdDaC2d0fakLFWp5HsZaCN+c8iOkTpnSwehEFIQYi1JDM
BgqrwWViwPd6imDMVpTAknzojgUIOodxxrzwBUbbMpBZO9PA2HI0poBavODtcNjcDJEqa8YGrIXp
3B0MCRDALYe/3ONLVUFOTCgbJzvhQOida2eXrUHkJ4zP1AWUPoqRj71L3EjeZX3sM9o3vVwfGDGz
e90AUik3Yb0RJNNkZbIUyRl4pl+GWodcNHX9mnvFVu8uhLH3O1EAl+Olp3QxbeRuzcwd5VDOHeJt
33Tz4oDv2XgLIWpZTxNcQPAw+vsd7kJ4qzuNdBuKoWvW0GViVUTWiMJdazWfXsOXg5uV5yXPjAgX
YHGrpPoAFRxB5+pHitkWnq3yFPMrqvqxz0JwIcHc19oxZY6FsaxPM6yq7unuIDWvM/eUngfBD6XN
nJBN1sHk5R1/kxXpr935ukdJdUtvE3Yyj1/12vvvLkJl4gJQF7mtFB9HjuDz+h9rbzQ+UNQhbhxV
UDtmAmtxMACYDE2WrEVyUAmb8xJYFKq2Ezu3hkvX0MpnS7IAe7+e3iN2BAFhVowF0DF4KBc0IofL
NIYCRDkzl/hVEjcFCprB3oZND6EGXwLRThE8PCvTEzGoS+tNg0szYnUE0dnhFe51AEb1pEsCfpVL
QYdQ2M6VNduS98nVtvaON3mxJStLlGmgsw5C35WDmY1pPpmfZeeIt9CNS8LD29IVr6eavDK6mcfS
kFBP6I+EQrld974ShfbVhD9YfrlWEzKt2Rolqzy8rrR/nOw1UuDFk6b4E48cbeeF55AmFWAH9Xy5
S4s/s6NOsg7ivTxKSkxdC27YgJRRe+jd5Lp7KJ5zEKUhnYWhsqd07IKT/A833PwzHCpLJTTa5gT8
hX+/950I9kD4l3Ee/BzNsX8OE51ps0Vr5NuyIRJDYKv3Spq6USW/nAlzNKFodQxGwzS6QXG6wIE1
ZygcA3TIkXwH8Aoz4te1+kU0MsJMSoBAr2AWwgZUuTgPaqEHqzUgX9EMcCYR73aOYQALJijvM2bH
yDYTDBmRaFpWDSKPYN/Yl/sK5kgtkAwCTXRbMi1Ixb0PR0fssuoE5uMsV/m5ibRJnkE7EakArOi1
R0qMzMXl6wodFVpG4CF3Mvqy9Rape6ni2PU4ftq4tftsL3AQ7f9uVdgP2FmApLOahnPWz5hBCJgg
EtmIRA8AKWDlgqeHJN+hVyXod1MKzILa5VijNM+pzidj88g7g7Opui7k7os6yHlvaps5I/fiqIIq
k8MSyEj1oUe9BXVriWLaiz6WRUQQ/mSvB8hVjmTmvSNCpYvmKR+3VEPnW+oZWKE8+2Y+LknrlRL4
kCPMnmKHVRchFr1qfpO4KyMS6EmhGcxJ2wJmgGodjSyUewXucSCLO0rOhz/y8tnOwJFLpPOP0adD
/mS0t20JYJEqLI9rPD/KWoirX0QD1qkIA7iAiSI9QKqBqpN4UTxo+VHZ6YSSW2yOuXRHYpWDnC6U
m7utZ8nsuKifLcng/VTR+5QYnjdscO9IPm9vcx5/lvbfri0vzDN+3Cz15Cbbit9TnEc8wgOyENVf
zen450pAvr4/4hGnDo1XELxdSXNgao49tXCTg7MhGatLMXsh3TBm7R53k+u47bchN2a4Dxt5PocF
1gj0zbEIuS+3+/Cw8rxgejrzPtJnPFip1BKjbE+oRHFuEv7BGmw4TWsedJwwigKF8cPQmU2eho3q
uEfcne9qI1CWBtzb/kwFdZHWWDzg0b36TTmf9db9jETW7DN/sdvpOpEzqeezjSGmGsSSSdpGJi+N
Hm3xWFbhjtL1mLWz35YYBe5nNycTO5elARAtEE4wt8EphiEZRB9td6O0G8JMSafouoVpyb6mSEIf
V1BuZ/UvOj8ptGo49ocVFkT1uP+ScVn2NsLSjzLlGdDhkAd6iTf1WqazCierXlSrDc3u4yQOOi/I
sc1OeoyOz1AKWoNxEZ+WuaXVVMETvo3lvEvAp5P/f4mS3pGNW/Z3hMLeeZJgXsMtR/h5hJbPzhdd
DFYmpzMJMPp2OArKq0iQ3+eINCFRVy2RsjdM8O7GXWo2+yDuGrUzZuK7QS3R0WYtYCsTeBmRuI3K
cIpqx7E2iE7DcDGvzpEhXFrpy/z9vnIB79P7Ikdrp39R+mABUR3hN0EmxWitJPKfNgXr2YbA7o74
RsMykBk6n5ShtUWGS+ESRlhmoPbf+wbBhgHcSP4obBLp5DPpR1eRDfHjOY48b94CKtfXnvZHnzoE
lqs9OghCfqssUw5DPyC6AeN3Z0DvLz3ztXXzxCt1dXnqVrKiLKCeA2zSbUn0Rj7sOAJaR5kGPZPK
S3DEmCcSSReTMAx22wY2H3Uhjz647kNmVgld9OnRgxSw/toIcOKn8Y5ivBhpzj80zJviGeUCRbSd
5UvZacLhUFjO747NKTTrIvlb8Smhnomn9bqQAD9sdDU9GK6pD8SxDGwT9TOeCq/FpR2bbSaXtiNX
MrTboCG3g7qLm4MaSgaIJnZpWV4o63G8YBK52D1WHtVJxgg5kHXQLelAxvwzjJseiw3xxoQJkjLB
dOlWCC+z9bMa/CdLagWZKJstnB4ndhJBLL8XS6bg80+FUlRIEC6FFObLZjFdYBM3QIR82c3d6xah
ps3Wxy/xRQdHyMJjdYodBkpvvcFWJSSq5wrJlb0pL2Cj3tQY8SVQcNSWkK3373aaPhkeZq7KGvmd
iwraQhLzxvIfcz5FjWnPwRIe+DoKC5Vzvu6S/Iqmnbv19lUnUJevqnGvxXGUOeZ0Zac0pCIvW4Jg
1/OhZGJiJJnwmFu8RlvUIKKsbN7LW46dqqq2B+uYwH/5zYfsq4wLT37s94yJtV4uM1n8jaXRBdVt
ysbWXuK0Djt0GLJ8XC3y6mXyU/EUKcXOaLuUY523sLgCmuHPB94K8sVCnjUV7+lfWsLFappda+i2
nWzNqkS9agWI6zpbtFKcguZYPyFgkny5fGuyRl3QsmgGPtFjp5HJYvn0l7pQa3Bb40gOBs79S9K1
U/wfS7C9QOAzuxPooaVESpQaWdQHvUyV4yV1rf79+FLFQPTdBbqG86MMsByacgml+Wik9lfZWlWD
k9ols2feicGhYI2LKPBOGwj3quK7GWuqgu+NuD1y0cbRVj2tV/Kyal+xOIFL6ILOoD74152qZLWk
X5oPZJPTM3Me8UOIccZKyKN+fmnDkEvsihGCTqPjICX+AfXyBBwxbaXaWi+YHbvwLsvfAQJl6o0m
wsIt+tNwC6K0H3OZSM8rHReI4qPyuBpLc+kTQXJjP2TW64DSRh79/tLZ853p9YqRP2RgZOLUmZkO
1BbsZz2M/8l77JuBtFFnwATIrmWcZqjbrQ93EhVzpYjjkpEG/q160YQOqU8fVHMCMpyWnY76P4Kg
vnuD6wdyEr/Qm9H2ZQL4odJ8g+ewMx/ADZhOP/lHpeDbBQSEMhla1+97N/fdW+IA4VueNMhXn7Ey
wZqKgK1Dmxj/+Ax30heNlsKNnZNnS9QMnjWURAvhhjcvyso+I7hf2yNh5EbtU0fsUtEjvprTp72m
dJk7MGetkMEwLnJ+j9/2GmDOTCvBGte1nVtpVUEr5GrkrzSxhcUkKhVJkEnKpBJhgsFp3lh2Xfgq
XnDijbwXeqnAE0PKhKsaY+cJbllR8zxSy80VXwRltqz7157cm1reTbK0Y1aHaeaOytLR6N8NvHG5
lB09mAP98g/owcLuPQw+I2Dqzs5V5llW5wCveCT11fqsDTrMu/qVfznhvRwEH94vR3Nd1yyRYWcW
l9XffQWTqOs+ymBlCrmpsmLphYCq5ZYveRb3So2YJROq+gxgLcUnl2RkHoaH+pBvmYc0G7s26wCq
oKrZ696iPEEaMVekuf62FfAK0M32VO/7Vrj6vgOs3yL2FZqM1Qt1mSm7ADU1tt1Ox/0JUTiUc2k5
/EQNNa1fVgfPnx5xy+gOcRJr9HiZlg534zYsOTAThQJWpC1fj51gU+wnQWo6rdVLWfxDglndtgmg
V+7Gr7POgcM77xZgzpr0hqiLIC8AJkmyVvnSm5a5RN+E7apAamtrSYkT3LM2Gm03n8Mc+g5Iwejd
QdZaGolHxQsUpSnvwieMASk1vp3vpDPhF791iDPSeajVroGEmQ90PbaT4gecgz2err2Tr3RYEIGC
W9S2U3WNg3j6JeUARagu/TMF/mOCGwCnzaKk17FYKq6hz8OuD6Xq5VRbvRJyDuKLLTLyo4KQcEay
PRrhaav76WRkGACs49SQdFoF1v1EGDWn/GG0xl4GDq3gX6FHjbvCcZX7komOpiyI//jA9JZUY1Qz
BzMlcUj+XwMQ3MZ5MdQH974HaAFx/Cp1ZYNfG70cr3VJzuDZi0EQoiWuMSwrVWaCtS8X4bDkXNmh
+X8E2I0OnaH0FMjJ5xAHQVanX9eaRkNLxiQGprhnqtECta7qDCWbVywkn0xkPKvCTyFPBUppbbtm
UkG977sq4dFE27qgvVFoOT3E5DoCqqN3xXsX66+1dBSwPnzAhquvLAeAeOpp7Yx0sUc0CNgQBJ1v
cMZdopByCg4ZjWVo8BejUgqezZzUMRCSan0tIuYRWKDEHfropl8n5T0u4DPwtNeUs5RO3aMEh3Gw
NJupD2mA3phD5JeDL3zEDMMY5IFtck5Fgzt3/d+JPFMaSj6D9lKtJLbei3LPvG9R7ze24cYa1xYj
b9BKCSVydIPixfys2e055mntl2V0KnCnaklUidmST93R6CGUy6X12ZkVZfIyQlHlemYigH4h3Boe
tCkX8ced+UVaSy1RbJkN72spGvtaQuEbC9cknkQIosFpu+tV3PfmcORwJ8AhNL2werNOWdRwHTDT
7H0H2fS/Q+seH8n6ZGsAF2kdpBAHL0ubH3uL7wTuYplP9ffYZzNifj7DTerbKP/mIABQ2Wa5b2ce
lLydhL+Ld0qYvhkdZFi/RGfMPk/I8LgqjXvRL/1qytl67d3ee4V2KLV78EXib/XSdpVGlNLn+a5c
N2dAnNfg8WCnBrM1qsp+UyJYXzrCmH4o3bLbCdl0gbm4xfw/VRlwD1GzSzrLnvZUJEdkvDHgViyq
gbFGoDCcrUpcn6d6WHDxiQAdBWa2+45K5xpeKc177zriycuC2UBCLMdc3Y+SWX+j58xqBX2vBwcN
gxvr2FnzqOPj0AVTxNm0etjiGs0uSEqPxYbL+3v23QjYzJXmyjW/WMMtORQtO706LebrfDga0XUh
mpJx904LmGhTBLOE/i0XXU8NgZ2kxC0MRpIF7w8xHWVas6TEixnE9WaRbv38kkJvlEaGnvT2q6fY
JHVdTUfQW/3BgfvmTJI55DJUTDsJXl+uc4SPL7/QZJMc8Pud04Bk/C4sBMK+X3UYU3HhLCPPbZe3
O1Ba7intDok+HAiB+Ep3pE6sbVcniLHdwOOK8hlMbqJwNQhoUGiyYSbMmQ02SB9DwYwjJ/VvRp4m
zudOHY4xq+NRsGfortrhwJedy8vJNCG13QqkasEFsZafbmikTSWW1IsQve3UUtcsqfnOht9xEzW8
XOAsIIUf6Dj1Jr785NxzLrc29257xZOkA6kWVTfrDbLIcL/qNxz3BesI+8nTifBUa6V83wY7tusJ
+pvwQHy/ADPq/ZEOJV/Rw4KVIdaoar5572PdyQifTuKfIdCxu9BI6O2JiAUVc5h45n6CxGd3bryj
dSI4Ny4veNev8gn0rx0nRIOTWsoA403VCi4CB9wQMVlndA93QlqfSgpQobqjmpcu6R10xlU8eGj5
07gQzorsa4pFJ20urxXdjEGL1QOJXyDSMXELQMfw7q1yvvwIDoXBM8fcoQinPikZLcN4bk0ymZNV
L7WnQABB/cFn7FVtclnyHV6ikkBOdoMrzrvZ3gORrAKrz6vpdChX5vidD/eTkqVWWAZiaBkyjjuq
M+KEna2CWCxMIEIGKF+fuZCA966jW/iUUaMz+Wsl8tWiULuqRGWfFLsvYeio7hYL371aA4XawY2h
b8Toj7rqbh2q8v8wRt7sjcbXTlg7sofis9n4X8wVDgw0RIGZHv3VGb4RQCNBBvmaFdfKR+ZEqObQ
N33d86z9HXnpuIuycZFKwFzb+9gMVQIy4VvTAbt+3B2K6kybM99BKr9Ue7N/qZmnu5dagRG1O7OC
EEfAlxVkeS11uvmSUH3b0cxBhmwRDxTJJGait4g7+Qit5EEAdMjCqsxXemap+VqthP1k81/CNLST
4mR+BcOjB6C6f2CNbQJFhKimzHzKt82UeN1Zsj+IfGxZWX7eEipGYLR/greDVoWB2ysb9PdY4ty6
mxyjgCGApcfjgfER8gTzdDR7w5UgcS+T+vnzZGhVkXmkZztsaF63wS4X3T+1iXelHNaq0iTgUOcY
/0jfu7uoNhkD96S+monmlrSenXxLugGrzsokeQQaHtIr245vbWoXdve7H9WQimxzvrlC6uo6VN3i
md7Y0SvEvLqeNTr0z0uLEA/qUAnLFjnTLExrzKaWKWWZmH1/FbPSTj+Gm1X0Vkpk0/5+iLxCt8Am
pMJnzo5UTSGxfghzUU9ZO7x7pAK9NeJjMwU9AGNy7e08atMz2BGkZmd1aGn2xbSuYw29JoV7Qc9C
kp+Nv7Ip8xDKaD1JTK2nH6ozbDYkh2Wns0k5wmgU//YrYoe7MDVCC7Ifo/8vqMPwUvbhDfukulQl
u0FuQoELAxkobRy/fKFYOsG7b4WZQonYJqvuElX8BCHVDt6d2HHehloedZ7Sz2cVeRhEiv7yvIkn
Nv3drVQfHe7ayt3Sn8cXJM1oq/aNbxu9PcQWfk4OAyCHrLE0GU4xlt3oXGlBWDEeyRnmPe8q+ouk
ruZaOlq+B314fhmTpCZ4ctYckhwxkepzJK1teNPCdwvRZlRbtko4pXdAzgFfxV36AZl2nLBTXVyf
HbbhrQWnn7uoYmeUtsjKnc9ZY7JShkb4Xqtcehe4SEv5r0ADCmiKMx923kE9E82rfniCoKQO9xL7
hz02LcVzbXqXj7trH4/4vFNPP/qonn6rU+g/9XPQFSyBw6W5F/zTWyJs8dCc/kSMsWmBS7qtJlGD
33u2Y08s0t7eJH6kDHElvAX+RjjDF+LGEI7NFTdfZ5i98FRgKvTHDJjeKJrrPGemWe0KCcLWtunZ
ipJfIJ+W4VP+IS2fNDEiwTVgYaQ+ZuMvBZpCvP5K0+bStPXwvvEPKzUqcR292l/J3qO1FNTfAhB3
rZIg1h9lfrahZv0PaaRcZsrsN29v39qWkksSSRc13o7EIdZD17+yVdbmb4qsMRNhY6iUz7HyEZ8Z
MakgQ/ONdhVVlQf6aA/MUgzORqo8HqwnFI0LhY72e6vI60JaPmuTLsNXLDdTt18CIJg1vdcWxFzw
6xcUHzmri6cLkyaU10wRXt0pQvHhHW/FnCrtotRk53L9xju/PDSRIHS1GOhNQfMtfGj/OsF+EjdR
XmG1gXg/TrwcCjaRNdQy9/QGasCS8DU4GTb04pzk8dkz1Pw58nq+z/4m3VKl+QadeJHbb/2LI48G
ZSaGrRdAp20LDAgMh99YHI6qjda1KAPPoN7nor0LGPfSAAE0qcDRKEtprg8p4+Ua1A44MH/GNBId
+GkhYvFOujgeDD2NBG+GfNEyA86DtvzOae4zd16Y1nNKRo0Ot3Bv/3bxgbNpujUBp5z0bY71knb+
fIv/kK6qWruCKRxYe5pCbw0x9CEzTeW3G2x/FLGG2oaxzvXuEZxyYoo18zXNfhUYGwZZo95he9wo
ho/ZYOgR7G8yHkhw5rALzP4TrIasGglkBXb4XI1/ZZ0cix7keDkKo3tPjd/bcHsFPcmGRIz8/f2p
SgSlMJgcrnedSUrwzUaaOrPxpsHWQa9nJS4PAOuHFooXbt32x5zAjktn8Dlw2xnffjemlbOZlqXY
2BNxfavjLTrxwZmPLHzZPhoRr5wIjiqzYfDpSSxxHDc5S4lHJ+KL03VdB7DeKusJGWmDCbzlC3kj
4uaAX/KwqizqA50G83Ku/p8W8DYaWkJysxXvWpJVLDjFyG6u+wpHnRn3BeJwm8PDudiNoy9/p45Z
2ncl60GhsRMo3vcMgACxRGVO8YcHHVWVYCMQQ4BIQE9SrLBtMvEG8w03H1k1Qa3JCX474yRQ1wiG
8oKM4o1F/gZOwwU7F0CjUykm5eRIxnYi3VmCgasBml+91ILz739UEEUm4watq3WjxiRdoFn4v71L
aH/tMBRY84VWZYZPeXzU2+6MZjHDRVVFQgD7Jwzn52bvRRDkL8DJK+ldmrdGk7mmuw49uuNdSCp1
B9hTF1KIodr/cTVASlLGBb+W8RDw3mh79OdZ0kKuMyaf+0M2UJjWGQyjEsk2s//7T5qwvxlpStYW
QuN3f7iiZiVHGRU/3/NVL3NSw+gCsYBiVTIIZbOxUGoYh0L8BO1zAOTsbZF+KEfYzDBrQurmb+a6
KoQyt5HVYVvJCytV67fE3IQL6iN9KxpKHSpaNA/n9SsgsD4khrkQSGWvdwZiKvzMNqxRNpmuy/Xa
cK0sbirl1q9bbW16WKUgx9afOFItb810J+uvdUhisVqmBQiwOL3EyfOmMpMyzE2F+fpACV1qq4MR
qctHWhyLaDL1GznTFtY/lG2Yxovue9d1xrkxUM1nhYEBm9zCKi9Dw9SyW6jLJqg7tqHgpV1KTmGU
iqQpk6PPhXYiG1Kp7rl8F9RCQVNLtGoxHxMQxnnY1RhAGP8JENGL0STROQWOKL09nwwajJgwwr1A
NUKTfezcoLTbxQ3sRRoeyVBmNd7tND+h5HuQr6ooXN5pkQvjcuyAoaqONOtgXzW0k5WeaNcIiVSJ
mOGMNDRMkluUoRPK4L4nvypus9SDKI6BzxZSYoIxPZrT19X2NqAkxOmt0LnIDqd2BG4/2rwi+OmT
D/0etwm1DDwDrZ6eBNyeFQVNkneETA/iYxIT+lcxSQCCJiK0aELXc5N5e33HTAfGL8MbEkZ6V8JX
anXzC+Eq5oqOwNwd31+FhRBay0rjp5c9ds9qEsGzf10+EhSG/UFoLqnle1Sb+1NOOxwJMnS3UFZP
iGysyiU1TOf5tZ8gsNJMeWpc4HwjeNMvsOo2VHNcXlfUgAZZJ12nNbvgaLPzyjZC+rmFlgIeXNit
yeX12/vWAQVDuBOSghHCu0pdahAc65+gS2P42UjXOEuW4Tc/P62NkCSCcprNNjNsB5D38iX5KY1G
ufM/Ju5YMmwdc0Zf7Nb78Izddh2hrvFZrLqoumHb0aggpYa+J1jJs49UxYNR0W/MiIl4Rok7SyUZ
uDI/6od4h+DFFb6hofKA8qNOhzQ5BpGjM2k7rAo4o5AuTenI4MCgWok3hvE0Ncw61rXtR74G3R8x
RaqHD6734tH28PKl3/LhDcA1hbLE4TrLOWznQBk1yuKovEaUvbb+dAXc1kZ9uXyluwQfZ5R7NJDV
YH+WXhDgHR03mUpMBxJVlKp4u2ml2fxk0xSjw4WjVDT0A/AxfnC+gar6XjMoPj5m9fsqbmun7MBf
y/HSFsZLsnSbFfsLKbheREQ/mHIIpWqMLVTQsVkXZJIdpi25qrzozVJ48rOkfHCQ/XcJK5j0caeo
6Y64MLvx6PrIw5m+oR0k7q4qoMaOxQ828jx6uIn2J2fFL+3i93EBEoeRMFHpcZPzTH8niDgMN1B3
ofP5y5h8wwlkA2IXsum/wysWK5hLvztSxZ5FMNCRpRBHgR7/gDZS3NKU10VKtOWGCJSy4D7BhIZm
eYbhGaXgpQg451vqHaLYUwbzkJ5bDKZFgOSFFo1JNov7Yt9YuPa0zxHxHhGNZiRY7WyEXfK0vg/v
DBw1I7SZD2elxuoasOxhFBCUpMLePO0ui1P1hzudMdqW+BOqnO9v2H4yXUaUIcqLzBpQrIJ76HLf
LFQ5wwsn2ljLgpA6r7jq39rRFRY1VI6YhA0vGaVhJ6XyKXLNMdkBPBHuXcbAguikeZo6qqjLOXZG
wjzCc5MnNSiElr/E+pcEXyAvvbRRySu5GnPNVKLlwIXgYZl/fjkzydNqGye91zSGQFg8L+OTIgab
xs5Bh/X8NtaP+1oCCyerzMAjGTa+KoBU27hNbkdtx4E6wCebIjpH1mYOLyh+97RsngNPJC+2jpBV
o/wkV7wDBEOq7Vm9RLxJ69a2lZdIq4uyixYgceciEj9Mhs1lRi6N6TCcD2EFfnZxEX5EhRf4O6Os
vdrGMVVR7i2yguLn/UFoWEObxWSW95oCXz9SD+MVCJQDn3J7T8909mtCcMmxmmU1kxZAZv8yJ+JX
hUiseB+idmILwFVl1CBkZJf+ZPkBr+ns7pmsRfYxiyTq0969HKTF5/kg5Lv949oTKYR1LcKdWriI
PklHIgoUuQhBWtfHb4v8jinzO+ryyPsclT0/sgG0wadVAwOAqxDKd6V7LI6tr/D25vWqdWOjzri8
l5iq6NNyAHh7MiEYyxjATGsgkcjrJNtni+QGntuAkGcu39c/V6fjC2duCIKNZKyyPlGtiu/WE1qa
qdYkl3zalSTOjBuwR7ip3Ihu08wy/PBiARnt73O1nnrCSwW7Y5LpxAPQBR0fbHv0pqOZC4ECIrF9
fnifT0VBfrg/0nRgSL1JhtNhaE2TDwbYNiNTgbzoy+VX/99vtGm2GV/K8p8GfGSopeZTE4TAtnCz
dBLHykmGKPjb2tKPKdMPK7eZqswruem18rh4DBY5tSAvqF2PO26iPZCLUs+r5A8d7HInxaAeRCOD
n95GdgPfMf69rNX1f6PtgCWsT/EvEWF/c7parswhFn9ZvXsDIvTOJobrJvFf6Wie9pzgOYsJgH5c
/Tm8cMFDnKp0iSdVy7CjnRD7GlOeCtCHqUMmOB6kqx1a0t6aAliiPLxidXi5bHOFKvkRYOF38uEw
DPeXvep3IJhhCRrMWQifMbfsf0RF02nfjiPuNkr80Ko0XvHwAST1KHDvOty04h2tK06nrl5mlPqK
aM58Y27K4iVzSrR3P8YVAwVzdwF80jl98AJXTn+p6eFrDB29tsJHCSqsu8CJ45trAW5kSZwpqpoE
iRT/cKaSINnJcdi25aVdW7/rWOq0o7t9wbRLGsAyRyMIB1QTZV872Kj1CNEnYJLnkZ/7G9BJxlZA
8R7PfuhojSKPT387JrjakLPCRR+35jvoUGDbmJ79c8NnyI2Zs36PTaY2jDWbcJgcFXFoyqCOWv56
WWVvJoOwBFWjZZ4Xyq9AkHke1gGbaJKcB9IG7dfDo86j9g5XhxU/ooTPiz+6+Srvp28sW/d5MpSM
hvWUmpu3KpBN7F0LldI3u8itKX/Qz8fe3R/b9thR93y3/8F77n5HDf7gWvJ6FExd5V/1eLH4GnDL
3n9JykecZk/x2qY3HFOVCA/GqHN8d7kalCoB+1TIg0CY1V0ddA7cR2ileVIJcbu3IViacByetXGb
T3ZuqGpYvuKOLtMRgtJd22JW5ClRUZPTspWhVtUmkQJ9K/QVCWtc9OBt6Ymi8Xl1oghBCoHkPBbl
0yChCV4X8Vle+Dm6xp7LBSjotX21sA82xKAhuPZI6K+Ni01QnpyzaRLlpIoyHHM1CjX4R3tWT43X
hmv+OKTWR/ZEHuIVE21lWD748ug0mPxk///wg+Ll+UpR60pOWUaP2rG4IIpb7QNYsrwtQPcAuZaq
YFVTVSzBqhg3ZL6I+gsSpvHe6mlufOgeIHfiUPVgD9zmL1KMZS62AOpP4pWIMM9/W3ispayRaQ1o
KLce496DQOk11YuTip36bDRGVu3stYv+PyfrNo5wlYmz1hYd2paUyyLbSHA6YepoD8ur1Gu0bpeJ
ObK9rLXfWihBIshKP4/7zkuGbkz3WDyX505UpuPkd3sWInkU7SeNH3klxrYS3OwdVbxX1IUd3iYK
+JjIfHJvoDTiu1TE9MV1vXzPsq/j1jHJADxvEdv5ljx5e2ziTyIcvC0pEoEqFuadORhZidstBfwU
1WwT/dj3zDwAgwshh2KHVkAmnSTLX07MXOc36L5+k8D+6Teq+iTdoxvt4gLLhahXN6YMYnNt1TEh
gF1ABrYzr+eRK5yINNt+VFPmVwF1THQGlAVDm/mzF6g2XO2HGNkt8pgbVX9RNp8uqE0cs8IM+0iX
+IfefyaLZXZILIfJ89bK50iNtbn/S5l5TiEENiovLW6xBdphZnC07SUJp3qi15Qmf9DGxoX3cOT+
Ysoy4hn7n749Zu3Cl2ktQDHKq1iHjEEpo/wNIxVo9d3CMzxqwW7asyIsp9wFK8lgSlrU0rwovv3c
L/OkhcGXWMpaFwj5ecaxVup77eIkewVVTgrcOQucYMsnxfQQ/OMKLOzNqkKKRfZNs/8McJ4eDuSM
8oqsx405NKxQYpWqHrVA6M8kxYt3VeJHKRce0eaj44e3RQTUCRPYqlY4WhaLkEOGSN1WYRO0rS8P
uQw4Ggdl5riKhUkygtIopN8AdhB0ORqTXIkCXqBXrCjSPCv4uPNVqtYITV2kh3AS4GjVY0ETDW3D
cPeRt7fOoySqk+jTCraCTW1LOVWgIC0axhr1IfzJomrPlzH8A/tESPZEZLkrQ/XrbI5aaQIq6Dfu
dH8zPOqwyHTWhmBbAT0++xqHJ0aETTIc/6nZx0xJOHb/BrweFOjx2QFC74I5S+Lmb4Wo0yfNHtZ5
Ft3ihsYCW/EWpNiZgvlzkX4oh/OjY9Knnoj8YGqoleljGNLbtW8dJLR0ZWHkb4FEMMlgx6zFXI4Z
gqfZoGWJMjOBmUIpmkYHBhhYr1ia9v6emL+UPOvS12/02bXnWHxtgoaFjBgWMDtbTyGoP/1BHDYb
djk7PvY9OPhzbCyVEy/gYPQdKJgFaztj26E6apfelfHdaXNiQzfn+rYUNQCZEeJKAjg/6Ebt1RXi
zHLv7/KpJoif/ur29NDmWEKXYbgyAu6HRCViF24MUTM8rZl0j2TNpCUYXgtEVk2gxHa4E0Xi89G0
xjYZDmrqlfcR8WrsSn3aLgggx51Q9F6g33LPl/ro+U+XDNWfEtFxgwsmYb4w58utXq8ZURKUCUYQ
yxfhXbBmPUYwM98uky7cw49H3gdE2Yj6cMW/NsNmMT34TlDYo21eU92EfPijiygQgD0GZUiskyks
09I4A+9re+yn4QkBdPLNB1Yj+UoSOCeGpM2kgd46s7+ahZCFES+L8Nfb5u6hFdloWmfPxybdZb2H
667qereHzvxR8yAStE0WBKN/18hnu6HGjpwmtQIvXDxLxHEctWtghrZTPCAz0wYHer3IxKn8a8PS
u1O4w62f/1ocp3jicQN+EVpVcstfp8GHe45UNhvCoJ2jA6sgSNMOrEXrUFHBty2fjucJyiCDSnNl
v6umArLDg95rLZjwakMfYei4RMDg7OtihjHEhAqz2jnff/Pdm7s2EFimM+jGpEWE8L+MRjb7nc9S
Cwht5QPj9O8N04X2sVu1BLR5cVPV+DEY7n8O4n3K2bF9goQle3elbXLdGauFMbD3uH96GrMyEzoF
hJ4qM+lxtJec9pNlZDJ7tsgtYT7ek/2xriusFxROs7UQE1/h55XiN+pHak2GcgZ2uOUBQ5ItOZww
0Orbt+Oz8iEsZzw6h2k0u04XENALICtqhh/oialYi+XHP9YEZbocXoqyIVVzkcnGnd5l0RjZr2TN
fhLSzT+zwM8OqRju4cc8fGOV4EP+Totj4ThjDPyywG7HYTFVLMzm9UYZGbfxvgzwfKx9g9bGxaCq
rP4FbECrw3HEyZ8Ol3c1nxeW0WndrOl/k0Qi5uXbo08j547ZiDttH5oasotcEI0VPn6zNwefAIPd
GL/Nv0qePeF8ncDfUM81gg6hSGUV53A5+cpihcua5mGAC36gejWoAZiXHJe2OxtkhARJ7QSw09w6
OREhNaxgF13rB/UNyWdAP66iY6eo0LwBmMGt5XxIpox2Bk2ZiGCEUYYyLHqee8JXP538iXzRN0RH
pv+iK4AD6zONxzhp1ecFnpI1UKRKcTh5fuyO7EjiNqXD6KGWiO1x4eK1hnpjXBnpC3pLI329yNK5
1GADCl1ENpjUHCxiEalLqyChUhKhltyDAmZbv/IiLrNt4r3DENkzSy8Jd7UTQxKza3AyrzU9srrU
Y8MvwJ3u5Kov4BY4j8rVJ3w+mFAQsE5toJBpSNQ/f2YePRaNg4YGhrVp7NTF6qFQ2fgprKcL5KTN
wjLOrSfH2nBR/tuO8ytgk05GeiCeM90FDhrEqJZ5M5ThkfZrChDh3EK7b1r4xXSR6O0x+Oviw/65
UcqfkNBRQVmxBa/Z/GfX11FLAB0YWMhhoJ44ZBJI4KvvWBfB4klU6MJpY1uzW4Qec02EsZijACqd
VB8HNs5fWseQtqhmWcGaBNeekiDLcxz5CsRf9/N6fGJkb1BnVMfQOWhEpENWkwvHnyuC8mRam6yN
vTh/MqFKiTthywC+WlZoRhX5Tc19bG94b2B0DRqv36VqAv1rupnYSn7wdGXrQW9HlZKrGyCmxw1e
i5hlG8f73ucqBbRhTa5OlA+mrfYaFswUOPYT82TStCSL45fVAMfXqt+qe1pgwUxUB/W8W8Ycxmpp
4B6n1NVcHPLrpZbezyg3inPcVQ/bq2yWPM5u0eNkGeyoW6ck105yXZ3i4gTze4TBHkxthlj8247p
MrIrO848Fm7cTkslTbVSPUgkVTrQc/KBs7MQzRLue/PhofhxndmodPkPfz43EuIWjWCPpx63Z9jk
LmdZ90Sld2Ly0d+AnJucld2CxgZuz6pXMOaG0PkmOmBzEx2P6y7Tg32ZwDeXD6Cyoddbx11rUG4O
2eyT4lyDNjbxNxxj2iSKEqDXrjcLaOalGdhZTxmudIVhR5XukbbE7Tr2wC7kddk1UHdFrJklYZRW
ROL68nZfRf1IOhVox90HrPzKTr1+u33hnegf31Ng4lPqikWc/s6+N0lgEbBTCGItkRd4mbKF7M9C
+JQIdTSGOuhUYzn98WlsovEi9dVZ80u31G6bMROdqT0VRTotTDoNW+DQP+KhOfWP/WE1PZDT/+dh
wkU/egwzIC49UCpyFtO8ytpdgtUl1ZUevOM3Ja/OjhRrF7cJdh7ZVJdNmypzW9XMIhb3gUXt0yYL
kP+0srCtr4gehrvk70LTKnzWLxCwQk+9jA08olMJ50RwZCx5BDa8h/GZ9I9XqmuYTSwN/shQVbfi
C+B31CeSK3t/h0jd3QKgVGvf35VEtxs5WUqz/YbpjKIfJaxH8RyRTYmnI4ZsxCITNfJELvpZufiN
kr2m2/V+QGFnMYRNXmmtvSsGX/qvOtrbJAsOtQMbtOZoLDOIzMITHq6KcaJHWFWn6jfEDeDY4gFG
h5XI9K7drWbvSVlATBXhY8dzqh/zmIMFl6M+3+VLpsDvcguHnDQPCA9VmDRWS1jp5CuODd5pE06y
DUUERFmFraI56II+KgSnBo0gvyjPZ5bN7R0jxjgVeLjmYxy8lq87ZVkhYewFHKvrTUW2F7KxT8As
uOk+5alMVNNOtQ2RUivswDDDqGeDzbHoaogZ7eajRTRNW8Q3I/UKt4CP2ruHD7y9W6ToOuRLg/di
21YcW4TC2xeQSQl8DwzFVqgmyDeRavSDza3iMo5FQfANOp1KCz0uNS49ZNXGM2An0cjT/Oz/M7xV
4oM8q20ZBVMuEsfzYEipiXm5xBlCKnAyWljWqvd40apyU9KVhbf2sDOEnU6thUXC9hY63hWdnivJ
0oCREG3/hN1eEgreJqliRsWvM6c3m/YXTuHNWY03QkKBM6zFB9gjWdDcUGGk7Ir0MOh4LIawEg5C
GYgwXeFteOTtyFArICH910L0ln2PSHZA1RiFFSaJSt9KksxBtXTd7ExjMV06yjSywgFu6wHUVWpr
g5oyaGmZHvYQwliw2uSRsGstMIoQhO+kfkzXg6bsZBMTSZ9x6bpjM9Ue9B0Q8YUq6pB5PkUGFcnl
TjByegmBssFKotcyEI1um522zkPRqXJrMJ6XYP8CIOPfE6g9pFcy41WgWpXejU6udYcKOgaPNx6j
+Na4wYL/MVUQQXR6J5AQjNMlDbIdwTN8ljJRUO/ZEQRC86w8hYmlQsxHj0KR55rADyaspjOrRyQl
QAFACMvG/M42jIJPe4NtdRX/BvWAO8ymwP52EdEYIM4fOFZJMU5vMwUhM5fF3LwSK/+xhv9KFekz
l1Yh4wwLHSEq7hDgX+ZOZr7jhIUEN6zuCEqCqDAiPFzHz2+wdY1pakVT9Re+toq/srccQRvaJ47k
2F6Hg5MdEfDicJPXyJWHGXKFrzZwYcv0/OfSS9QNTjxtZzgZ+7AXMcjPZf0ok6p2QW25LmOW106E
ISPSIw2zOg5UxE2kSVieSmzIUGPRtMj98ibUOUSdu2bMW5xwnq2tELFXvvCrxhY/RvmIMeglbusF
PFWUo51TQP8a6nDa7K2aaG6yVyW9o7a6tpJ52wIwGmRjDEjh8jA2L44PYzg3u11kNpvKSku2wSM6
1Inrj19p3h6RjNzqcgzbQS0qGZiLmuW5OdCZUERCRDtnw3EM7MdDuBUgoR5+7OknRVa0nF6ztOcg
HGWPX9R0QH7VqSwXwVkqPGCsb63/uCn77F/el9+BK0qlPlDxgsm2AbsANX/VUzDqryJ/7WakxOjN
tIz5eAm4Va8ClNrgcWiQQrbh9mtGi4sNaL30rPT4AK41+HRy9Au45kuCKHxanwiDzO5LBlUCXRJz
C8GhBO5HV3f/8OENoibmSfAVzWImTUqJDWws5p3xXWb1rLscLyHHyecoko1y4gUO4oQ7IQzTiGj9
lg22oQdt+y63xloNHrqB774nKliuiTma0r4FZPft/0SpPn7JqMvqEWT2Ov6fGeBCSoLma3kwKMQK
dsR5H3w35aY1Nbqk6fuYdEiYw1PVaMLlss6neTnI7jxiedHl8dipYN8efuiTaOzIx2f8K0iXAd3h
716U4IRRC5n2++9VPcbnTAhMxDtBHPxrVCxvBRRdTXd6WQonOdJ6/UTKCBzpFePVY6/INo+D3x1Q
4HXmZiQLTCx6Or3rhP98gXWDDWtk9RpYD9nn1BHs2Io3Nte67sXsunFf+rJvokRHbRRA7+nKqubv
CPy5NbFXoM8KoJB80wesaKO2fLbVHOE9ERPaVvb/8kQJ4EWp0Yvy06GqEZdcK7cnsXoa0EQc8aZn
V87SfdtKP21exUanMC29lZWY+2BKmceD8ylWmEgz8DsnzlWU+hJL0lFa9tciwoX4UYpZ7DC4bos4
K+1D/Cbv+vae9RmjbFm9z4ACa4NAiXvdePD0tM77Ut7+CEx9lLejUReMCaScmuXzxTb+QtaUtZjC
n6hCGBqeeRFftRPKy/dWY7zil+tJKyHC5y7VBlwy66RiT2JEFUVkqfG1ImlbF2mP2Y+qDBhTdMs8
MisG9UpNuOe11OFcOeCL/cVsNAwv5ygc+sogtFh/8nzYdh9WFLTFUMgmKB5XZNjMIO7wV8qQdcgc
zUb2uKL1tpdG4MOVeemQb7sIF4dHjp4Vl5LCXF+lThIqVdcGdJ7v67jiUIb+gJALkzMZdutabQLW
1utvGeNMB/w/LNO4FqNDEfbphh80pjY8VGPt8k8cDQxKx6k+FXxX2fp51IHzod6SPBTpCvSCQfad
H0Abt5Gx/MDrGwsmbebDWue7ppTL8Shv34IhNDKLVcnGXKMhCY1FQd/LzE3SXcRpqNkSdR9W6KMe
EF2qCzLfKJLx60Dy+Ko2ND18tAz7RU/B24wbyWhXRuPG71CKkClJ3g24e5vvKwF+NVhlCYYPl0o9
jQo8xZj2wyedVrtfRGyHI/NCvtFGi8/AVkXDjoOIMfe3NpppVZBOZpvYd5I9hVbaM4UxWaqiLB8i
G4gasHxfA4AU/mVPwFxMBJeaNycRg/WDdd5Xh7G4omSrl7mafeshaiyicXqttoW7Z9o9rr6nW4t4
HQDJz310/YTgu2P+p93r7cT9XCqwY94WAsy1dy1Vgp4ZiJ7nmCf7qtdGjPywbRm6r6+fsqRA+l3g
ejgZQ9EiH7JxV1jC3zq1BQO0bWSGy5FGlgPaFnInQoGgbMv1imYTsGcUNI9dqKF86XEpjpcvIwHb
onDmtt3ZpWU2ChOKvJ1/JUKlqlD0V95WPHBmMqevsrw6eG1wKKh6jx8WP+S1Z3ddkvyajCgnXnVX
B4r4nLwpZRtX3j2iDSfPdytVz76FUr4ZJongmw0iYtl/t5Qk2iy1KmbqyXXIkkrcpyzFEw7Y3GVC
kJOhkSNeABdjflwci0Qv7WtWcTSOqJIHN6C/o+wNLOWb6rjCleNRlaxAwNLWIjZZ7TDWCblD+g8e
/y0AsHQc4qxQrKu2FiAZfOrf3w46MZHmh1ocVMTiubI2w6oWvx2cTXq2oYCgWkm8BaksNhiWRuhh
8ySZ3BsWGCnK7Msh38ekazWWZ+c4QW96wbJP5Cdap7CiC8+AVLvlnjEBnentmo0v12SP7CPpKgVx
k8PXqMrjWr5//3soL8FKZrC1dKMfsJXoV7Zf6QvUrS0DAlpukElWXnyxPJHXQdurQph/AmiDanra
0SL51VrcF11kR4RAXyMtxdh+TJML/20SKQkd+XZp813C6yR9yYdpkZI43XbLuiHR5IR3/ZdAS4A2
VeGZ/lDPfqQxoI63AgT/RIqOJkqi3NM257Op4GbRhEmw5pX7KOhCjExTh4GZCKJYzLExCDji34u3
GOEL1VMYFAzozgbDHGSYTe/HmgjL35lOdiB72+d9h8/MYOvKPZElSvO7fzdFPK0cTGPacgxhMagH
0JUPyajOuRzh4OV4HFb7QIycmxbbqfG1c6if/aSuAT6eq06vTU5FYBt28bbz2uKhwGV/aTMgHxS2
wqoY9k/6aDxhJIInjwzd7K1g+rlkKBYv2vFEhFonxsf5mOFpYwPu2uMtPkvSJEUFFvR5IqRX2kmT
OF6opCiKy4EoBkAqjfQMe80oBEE72Y6IlxnDPkvdjg1NxRnbvKRhZ92BKdgbZCHxM1sHYwfayEq2
pm5+DOydu9jHaYY5ImOKPVi6lLXx5ZhRNIRzKnVGAqhwUND3i6cUFgZKh8rKN45b6lcDvyWBk9ri
xH3JCQ+ySRzgOjO8Yp5+mwN1FgiIOunnhjRPXEluP9Cnb7hc9ML6j9dQ9p3DUwgLTbEkGznln0KC
gqAXtl020q/WgxoB9xvve4Wssy7/1VHAFAYsqqtPAtQ2GKPf44vxcKO+FQJqJnPIQ+mvPAB2Togz
Un/xyueQwcH6+8gso34XeW62SxE1K99PkQg3KhdxpZrtWvcqKptvIkbitTtqQlQWfYuVTb82fO9s
C9FR/rakw0FOK1d69CS7eaXtoY19fu19BGNefYH1GWraEghCSbK7f1QPiUzmoGJGqgUo/x0auxID
Lf/kfEBW1kv3j7ebPdVDlIw/kY6nJRctBkqyRwazkifvf62BjKgt7wR8sGQaOru+uAsO7A2jD7w3
4oStrfx0LpMNF1XfMCGzgA2GU4xE1kLuIq+uaUoXFJVVFpRcjn2pseReldJpEYieRXTMW/C9WwL0
yhqLyANLjrE3K5ERUNY3o603ccxIso4W1FTb1UOiOlY5ipCHlNHmLSrqWKrCqset+UIHBlClznA/
RGJ0Th3q2m9aKzcPAovIebRPTDJywRY3+/Q8FgK6BF/dELVS9vQbDjIb0Z6t21ZelzBXuiKxKiXq
e0MniZiabBJ3/wGwkcDjGA6SSM4WQ69BgMr7Rt+NO1VUqzqUUBpnjcQrhJkco1eyFaxFqz8dpgia
aJPH+CNcpmFuROXlnznIK+D2g7Td+c8gcEp3FBUChf2C+dtTMrVbiCT+shVotVMRKWW0rdZl9k1f
zc3VO7jnFxUHkS66BPCM4BK4t2215xevhaLy7QVUVcbzXAlVGjjjOtJMzy3l3x2sMZ6GghPdWp/u
5fy+85e9ORJM1C0M6/+wkqpNz3WdKkmf4+4cepJ6+Z+nk7QfpWAzkZQZ1JD7yAhJWVdX5YC72SVl
YpQmAa7RBHIiDom6P2ZH4traCJR/r0NHphIjS07OljuGSkLiCYuHHmFvA3qTUeRF8xnEup7Bsxoz
f7EBj1RSOuGDPeUGfbIzVj5FsC8weqKtWKCU+aNQMihmCUQwYGW0VDoy6xrn84KH8nfDz+lZqgrw
3lkJF6CS8bqYvaZEAHxoYO5SDJp+Y6lOAjVruHqiBdW4pC0cLbocR7CIwQEFdRf+BM8PIq96gS8/
xMOmwbHhYU7qTh/0bEB/Rjrtc4aNoxSPSV5W96Ge6B4MvZfZ5Gfp/nV0GgAL98nTqPXDwe+brghw
KxwnSYrcnv3g8Hd0g6Qsu7lv4HWNVdBz5qSVL1rXer+kpe989LXQigw48wy+/IFH+FgOs0we+1JA
NweZet5BqTtiNw+coI6bIpGVYkAlGclJU4O5CCQZiDHTwozsPtmB1v3/BnGo2yi0ZB0APfQqHheA
AHOZAdPrsso28eQ2NcHDpEao9wnljuCDQokCw8RXMj6RtZlx5+SvKXXO1PeH4gHUkT9itHuGekhG
dcTJWjqTzSpFwf4ih11tDIGxi4qzZKda2qHY7TzR6Jk/yaIIcw6X42dY/g8oGT9chFaZ2SxvrRnF
FoKa/QZQ44rGRd+tmxd2AH765JpPuty3za8hHHbdQx9BjmRTqSMxe0AIy5euxFRmxaJNhFsCe4Hr
t9oIfF+bWiaoF6Hgt4KnkNgnqRXwSG6ksNDcLBFewmUyFYuqdW+OkDOfswhhCf490mTf6TaXEYgH
pJt+rDlsBpYL/ZP0webER/77zKM2RSukNDWlNYdJdfiEwGgQUDy+irPkYJzzXEUwkoRMOzMZ+Tx1
/hMuRDIlVV2h2IeVqB3x5U45i+EPqhdEvNOgW0sPayezRh4Q7/7FTKU1bK+K85QAz7a9fcvbcc5F
xIMLezr/BpMaWSo4kSJuqfzl9n127l4RzboT1Pg4H6b+UsOkvk22CXoCBPCR925vkyqD4KJT7dsP
Nh5f4Z1vtt+Dyn3KvrYkJOSWgYZGFrWqs71r1vObe2vJGhZkSJVR+C05j7spp62couMhwzj6eYqC
8GD0Ubk4P0+sNFXuAGPVcgNlwCZ4BnYWrdB3aYaK7NIUz0Iqcs7bhnfcm7+j7O7BMdCzfJL+auoX
PIrMzLPVLiEBewzrN/sD0L0s7ujC/J8nBSIUIgzC4Xb1rJcNnERXncL52iZFT/y1iy+4ph/IhmTI
ueyrMvyrPsRQUlQ+P1tnS2TAQ8sMoSn2qrUjAkY/5tXelOS4/17U4AC/cV50B7oVugH1/P4qvIpX
Lz1mYaVYO6lJ5XmaFl01/LzHMDRtVPsbgpIg/t/rLFTaFdnSzixgVxfen/s9voLiwLGcUN1ISU1i
VuvxULHhjPVDONyXEB+1I8K1DXNPgYi7qSvQomQjvAZY5Il79AAOpdQZy5vlTTupHVL4RWtDo2VF
0tM3d6nBZrPGM4f4l9yaxFIsZluhjLyMuA+YLt6xTXNQYmD/wwDWyh5vERI93PoEMisrWU9nLSXj
boWK+p1EiBYSUXVOfTY63KmMyak9MYbuSag1wVkASqkEsa05i51FMCNEgdsQ4Bg8ytdC66XyqWFt
pv6QgMR+02Hcu4VYo0+3Y0JBXedQAp5M2uq+CfjQ+zBow73kzrazmug7AfiKMUhxqG1B4kG4Sp13
ZRhn6w/DNy5B5kv8ME0aDr4fKOnvpSZPgHZYFDTla1wzhJUZPoH1m32E4e0b5rTq5KxqHdqvJY6m
t6pF0P5zIwTUa32aC/nMPjm1yaQ91+QKWFTm5S9WXz8GJP+FFXTDpR6kgFE+cMgxWxaNv1HAtaKb
BNgBjLI0mUGnsGRYCjQdgWwNWvpJ75FJTTrB7Dql76l2H3/ypAY61S13Nuihk+ErheWS48mosuiy
N84HKtGFZWjxp/+TWINQntwL3wIhZx0c+1TquNWtoyMZrs5/J2fhOD6tW/6bkS6Ew7058yxUTy4p
RrKbjZBSZ5fXlSmR1clP+5tyaGf7jHLPJV2ntPxE4TdLWpDP5CK9bU0ewI4iiYtvghRNhorDOzDA
ovsCbCjxxVu4otuBE1n92+OB8X7KDRkFasHBM8kbq7ps9vufWx7fgsFtWjEusQb8VDhh9kVAwBjE
yGCOIHMxzqGwkzkizm92uTRaSLcPmcsHe8iyvdctGVraxjAI9gat9mDrMvpLDvOO/gOyZyryysTJ
+rowDg6M94wobypgvDDdjcbnMSqcDxsduy08Sw0HkIh+dNvrPByCZchDuVxcAtVhrH7uah25Ah0y
a4GIQRrXAssoCd4754eH8BEVlDzJi50ui+rthcfAMY5ZbG+HM4jHcLmcCW5xB46T2Q9wov6UKLtT
+btPQ2kgKcisSJZAPR9Mn9NDUyEOfdTJUn8BKq2JvAg1PNhmOoWVT7+yjGN1ZLgBq/XSKfh+qJoV
2/+OVHyl5VZjeIn4HljvcneU2+pWw6ZZ0YmTw1wXUk0RPR89yoK+3YWzWvJ2wmbSMyH6Nd1dTO8w
lBKJrICH2ZkSxo2LGzM3GTMOJFUJrwr686ONg92PmoIRE6yeRyG/M+prSiCfm2lyU3/8G0JEDgWA
YRSMLn/H9ajiNg1AzdO+5NKxIdZ/IXAoTm2FnKrmnOhVAu5wA5N7eL3lZcS83bIDmBQoOF4JykAu
bL8wWL63g0eT6JgghtHfb/16YDZDT4Qh2VeWTnRfgNxdhTF3IcETJ4K7oTHNvIL9CmLUz8Ki30JI
vjiSPsfnwhGAERKRNAL51jUy9k0djKdWj7MrAWRZ6l/cAPnk1gz1hQMmDOlI3d0H5a8bgd1xn96h
OrI6DjAEp6dsOAG+obXBCxcMpRVx+vuH07mr4vMpSeuQ5CXNDMPqDYoQfkMRQaz/DTSSMT0P7iTp
25FjlR0+bg2gKVoIm36kmqtdIeVshE5XN/NoaqQkoxVMvRz4HaDEm2gF4STK1xEZE60wAGnHcVeY
YcGfyVgQErKMzBlPP6ip4c5t3AkSBgaS7PrG7hnFAU6I9S9Y8QnXSaY7FBDMN/gqTCgC4spe94XE
lDnYBF12Be5sjlYhjPlAGxgoMHZki+sFfSx9uqADYja+5WV3zLqLwQoSyciIwCPEWsmdF6T3oHrh
1qpLCrcOvc272NCMnPnGNLVSkDBJs1/CJW4brFq8zWhqCZ9u6G0vh/a4qXFEtEpTqTZHY7oSv6th
UxRt8rZNYtiqVpWFsTVmBiBUGWdeoSX8B+J8bSoDZO2VeBzYadX2hxp3ciBFGAcR0Ig2Slozxrpi
/jMgrMYZSpbSyAUpkOVJMuD54vZ9TNj/u7ObSv/0/OiRHOgAsVsQAkwAqWtdVKl2rDflZ9klGZXl
ajkhNNywRg7sSxcUT5txCvk9wxBoVV5C5kbgIZ42WMluihrvkK/ORVz+hwEce+TEXD1xfXbmW4AX
ure0vAaBjvrD3yuydI6Ko0Pp2w8sSvZwl0Uljze5AA6OE5M2XFUY7r6B20tMPlw0XbNpH0v06/ba
cZP91TCKuqzXSUj1BSL5tGwI1WiFbR4qZUDFye0+6Ch++2aLm8LJoXOL14lkazaE6XHF3VEnBKVP
fcwHm0d4RoHUqlqM9763bTkkg+24d2vnq7O2ZTW2opWuPI9t4acf3yz/VMGWtyL83/3r6X/04ymT
v1q7My7pw0EACGgqSbAeqSGX3es/7AMtLJZFd+1CBGrhXob/qB1Hpa5HVnN4eM7uXs2kUOcIfjxx
hGpOjrKVf9LEAd8huuqdTirsK/HIvsE0geZVHBlWFJG65+iknIJm4yqhELrLhaB7HfeSlzRoBpYo
dpkBQC2fvSHzeWwneWmXIMmH6gZyxwTlgutiu3PuA91ZkvGuXJE9uIDcKMi+len79ltzYlm3n8+3
exyP25Q8B4diCn3LtfoSMBqN8XxW8h2T6FOGzWa+rrX3XpBV763jjuljO7iXM25xZdeVFkzt4X+r
nkv8oVOaFd1UIC3rtJaPDoHREhU8tMU1YMYeavn6Yy1hkFsZE78Pnbx2nnQdt/NB1XEZQh3K15Q0
pqMq7JQeb8nCAvdQzvWuy7eRtSM5jIKydW6OvdSJm0Psr2ex266SKkz9zHbsk25TSCM+uLcNc3mH
knDb9uxd6udZfM2Q/Pv7jL6INdEgJ4AD1fJeC1pBabH5wSOId/NrTqGk2iyrbIcRQKDrzF+w+np1
VZb3mrMKueLto/nKNaxVmK1Tw3L0nhsoYOKTXnl117XMMtBOWCJWX1vKyPWvtbk1A8yT73tV6R/S
4pvxsDacEpliuxwaICoHWcFLAE5jGfWRGAyuD4ZQYuOI7YKCUCDeE1CnpA6CqkTDuzgWdMzKrjJp
mpXNFobEe2AFiOMwUsbF66yWofdRaVVjStH7eRArHTo2reUWbqXsWrPUola3iwStlaGpoXiIef05
D7MN7VrsXrXQ0EwlmrBfUYH94ra2x4tVpuGDDBLIiyj+M3IxAHllCHhEdgPqwaHn2CnPRHlrbLSv
QKHYbbVLUA4wrTd3WdK7nWmvWIr/4dE2MAn1CuNbgCQTLNS5cS1+4XtXMaSMfcfKYaI5/lZaLyB2
bTyDXXd7xjc+FMtqormf9QlRcXSJ7xRUz7cRrJOy52spMX6a/ccnxOebLUGQsurmZCO+LdavxoDJ
Hg6ZLRG+NO0a0/u6YkMQMoJ/kfbXnyyusx+sYLM0sDR+cuJv0nP08KQoLmMlURCgJqPbhD4D3tdV
4XjzxpuxXrkxbcsyarRnN7KnMgk4YaRQVJobW3ZR6SY0a/ipj3dwKP+VZrLj7EekvCvVtq8O3Xi5
ygfGUvRFA+p1JvMfXVr+VwTu5vj4ReIahesOX9xVgbJbrmFSsj2Dw0/4iF+1oHTCWF3axtWXSm+k
4hhYGdQRcYuAwQiWmO6xsfJ2hmqQ21knEVN0mmKB0zS0IU+Q9rEwUZCPkf3HEvwMbHT35cUorHn9
tFjT0276kW4PHJmVGmsVhnbVPz0QFLACGWgcQ0DotvMzaw0B/pR1a/1fQ0vrTOeTXYKIkomRbVJP
vgeKyl+dJpU3op1sH6WTZtjGQEp6rIiOgiy8ute7vIpaze76m+kbH5AK4K5Mu04m6cOMIQ1QSSL4
F5/LSDuQjJ0VedAzMPKlrqY1tXtp2wx9wUZlDlk4ccMFCYhtVTce5hVV/JXXr/x9CyZEQRCjeV1Y
XxDtsdifsceHhf+UAGdhLbfBVSGeMw7Xa4bukDv4vkxdMN6rOOeRyPelbS1u91Vvgr1wuZEphTs/
qFKVXOJ5XaLs+ThcmZ65/EYGxQJDZhAct15cHLzyL1erMjeynp1zqo+b8zHXfhXYVFs5tXTlLwvD
Mm2ZNk7TUdergcu0cM/e7K3njg1r7zFoot6RAbs0jttN2JnysPfWOY4aeAhNMBJTqGZER+RY42Yx
GfixD2J5HLzRlVq3zwwbXVZ79KergO/DsDSbZwpphRxjo/zwYRAJhihM4kCnoQq6tyGlFv+1Gjm2
ttTVMdBAEtCQhdN3V1QD/ooyczUVG4+3k2e0J+8jBZMANa0aycgzYkBxWUz7r1RjN7+WniqfOWDt
llnbxnWxBxmu9yAM9wm0F2WRhDCGsR2oR696zuTbhadnwTPFDYwLYOcF+9nT5crfEVt12Z+rnJ33
QZ+GVAw1PFHLiiqVDF7erhVTVNNQV1M8jkfhD8zlpF9Kqh0suan2mvrqrvNqCML+13K50+V+qGRh
wS8NjqTbp4pCr1XMos3hEQOFDhSGBl6wy7ghjOPLHg3yQT+EVajWrYrIDINRh8VCsZ3HZklpTDYH
26VGZzdeGdeK7aPmtN5NLEfnB/W+9UVe44uZls+ae/C9RZ/jNfxtdR2ahJTDUpm4+5rgrWhMdN9h
mAq+UvL5BLeypo3jx25HKqVCWMN6497Ki90PwSBwu4c9G62hhzpya/nUf+g85h2q6q1LqFxhfxws
HB50a6qM6fBLHqG3cYWAlXm0YFqHXmJiC1dolcRMJ0S61E/mqhuigZbsb8KlE9FyM/eIqaXh2l+A
Aw2VP+TGeR4yYsimTxliifjFZTQxpvAhdO3TxEuUPzOr0FLyNh/pREdOkA1QeAgdlE8i1QtH67J+
V/vKgT5oRZ4u2zQaIA4gr2I/lw3aLGcIze2RddoYlA3mXy04D9PSfq/vDHXlh9QTG+AQjzqwKkVu
poT1iJgs24oRyxaSag1zshDD2dmnTZ8ixCRjZXKV5TkjssLOAJPpTXA0SbuZInkwwmdAzP+pcMM+
E0pdZ2aD5rkjqnphH8jM2XG0QGy71vbv170agC3jeN6Dso2L3gjOd8eUt8nJSOx09mbckIH9P1Vf
kX3vK2wwItUhCuWQgC8F2xjgnMscPGY0/uiMoHxUp/95rfdci/bOyCUY83jl5RH8BesT9qY3CZ9+
7cd6a/S3WTz8UdDsn1lYapiUipVrMRXp6xGo6QD/G2bd1tw2EHuWZoVCooJtxsHLs5tSJkBsfDzq
sjKm0vzm+6n1MvDL0U68HXfGho8PqZD6sWSOuBzNX88pWjPwiocZe6ElNL5T22VRO6kf7H8ElPYc
thrVtTKGUpQ7PopR/or8ZUlmnMD6jjmVS4Z4+SepLOHUchl5DYVIMaqxtjJbnEHVU15WpmMpHJjF
FsEd0NQCtDgtFJkONhQerdUugf3eqXJTmaYl//hc4ZqVlGp2J0EdkO2WWauYAPlZhBBrxoPwpHVg
qOSt+KjCtorO3rDXzMfN+TDNeSuS1Mur2of194Ok0TYbuL4373vNn2sHkDkUxSVHv++4TSSluz0J
sw1uNQfk2nCrkQoRq99AuxKP/9xCnCWcIwSTgoSY4Mx+Ok7rRE4W4SpRcudYJLFrfXqparleVP9B
P53RswFiWnZUuMyKmhqxgGj/6iz1kAsn6n+m3T1l/HDbS2y27Yp8vynK+g21fAX2UJLKBx/d5+DF
cnEvY+zNjIjU+EwWYycQfVg/d105x4kFcwoJg65N5X9fgVgZyKPgpM+9TdmWiaH5y6UlaO30n3Sc
SsFXeaZLmooiPsS9xIjWzWT6N+gWZvWtsZQFDmaFCpCc/SNz2oNYQoFfwaIfQNoGlZ3KFgUUbahr
+58zs9pcb+lV4X4WJPgVgF/GqEWQgs5dlEFRKKgVd+ixoXlYzeODju4hVtI4A+RiI7ONAmiAn6dI
G5RDfbZE48H4AUsmel0DCbjtsEcU9vZAKaH0fBnj23JPCO2Xuji/9yrsmVSmdAZxUOlHaVnEaAE9
7sYRpEMUcAAiegjaToHI+Wl/PG0jBfTbEc+HUQCpXd8eJH54YvWE4RJRkd/8d+WNN/yXw7K2EO/P
J3p5IABFyX+rhmfQKDFxNlazUQbv8hcJVHyP3DHQgLecntKskuEpNXyv4eHnbgBaUnLl4ckZFbx2
Uxdvu0weYa4UuSGoi2bEROhEvaSgkxIFvITwhz+PBFlqGUg5B1zh2aV8sRLSaOi9P+tIXMk33dBW
DdpNOkP4tHkrd+h/th1/0ueNAfgMupO7lQ4Qb8jLrTRyNWgRwCbVSdDqveLvWfO3/rU7nUQuG/Td
+DdBelai1tGz1re4YjLzid3JKwfzsoa6npX8pCUEgRsNm6IwpVQnOuxsigq1z3HSluGbSrKbXUvx
KheyUqAST7i2Cv1vkF3B6ZugazxsHaHYP3aIObiOrE5o9xb3EfZdliBO4PGNnUTmtrWdCb9fwtML
Yp0cJ62pUZY4CGrYSXKVpqaWoHmzWtEo70E8OVxGDxYYqGLREd2wwD8ZbpHWUZnkKPfFxcl0j6A4
liwDEFxKXOylg9UDQDeeSvHcymKWk3Es9sTCIzPUWkc2Kfa+PcyM17SQQ/JV12b/cuqv9/XUrAnF
TFb6jZQ0RB3DvjZcM3435JnmmX3ap9/0CacV5a6ta7pEegBPXj08jZRZwXqS1uQvh2P36Olc/cNE
Z+inDUWt9Qj6PXA3rNuscKhqpw4y1ey1IZtz6bkdnFwEomAdZ0F9NBV/8XmPOGgdMDd29rQsfQ4f
+gqUuE+tFTZ7mXtdB6VrbfyOAGMHM1pvPUbdK3cr/mVKLUjrtuQ86jWWx6y4e93hIr4jl9oUb5MU
9d6DV9VrcuGuxhgpXs/dVTgzRUG2eplrtVQ8E0RMNWhZtUDL5msqnW/8rfJI3D3JDuhwuLzYAPYI
YZagsDYa9nUTow4yctLMz4tNIDHnnWMOaFT7sorKHmUyTeWnIeTMZTZC8RArBjHqusH2FB6zNIwe
haG92CZWMDgFCWdVsYIjH0YlxhlQVDfpzbwhQKkCyR1dGFBP1IV8P7aJAKIusyRPbxJIQgllVyLK
AG25BrRX1rJC4zRpTFq5lDOwDPtw9xG/QtLMUoY91r78hsiBMxppqglEDSEQo3yfvugO9O0sBsGL
AD/nJiRyY+nsUNZJFP9CNf0zsazNZPEBbKZDTgpTuzzDq79o8J4Qswlftm7yW9+z7TG8i2pVfyWw
qIX9nLefRPdWLjnxWWElzdsgHtGI2uJ0WQb09nfmY74sZmarN5I74TqwXgarPKxwsvuiezvw+emC
M90wmWvGEh8AaauoOJejNvbki2LI/LsZC8T3YS7dIQltl/1N1ud6qYmHRMG3Mt6DYZMkqJ6TGLxp
BIb+cL+T+amJnGOVT+8tlmo2ulp5+upmZFbxogHeKwBJHq15j0sLOhbEgPB0C3Y4ip0gfBK529R9
15P8ki+LZEZU+5x4zBbJNvCznd7aGIJJeL4erDHHSoCgVYSwjoG8K6hE6ghwbzK/qrxvNagjRNZt
CIMMcgu4LAslPUpQnxkIpsdh4vpwaAVF+9ozGbDlidPYyLDi4bhUbpMQsrCxwmdTqhQ8e99j0hG6
oW/a+OF1qHQhit9ExkrnI2Lr8G0v6sJfvERUm6YXX5aNFGaVqRrxN0ccxr2uN+qHElhEsMA3SuWR
MjC/TZrSDiyuS3EGEDBwaSTncTNCUc+CsApr0sAthNAL+WS8s0yhMRH3xWENoPjbqm9jg05tvTj8
hjo7z+zZuMtbzc3KIL5e4pvQm1eaU1LdmzVfpLmZ5gIsqnKgWTzmigkMDLPzfiEBUOA/qHrFtbQ4
Eys0ETCW3x7ZiHojR08s9jaqHlUGhX3/Ho2qGvbqfwFiCQ1Wzd/Ry8wMnTLmYBug9huyCnNtgNh9
1OkPAbEfgbnlnBa6PHlRHHBh9Im5tlRtUfPKeXd/7Yc4znq5HXUzFNNNUa+rziJ59+T1Eo6XcJrv
naMumUOOG7I9RPuDAAEGhrNWLWEkD9zqqmfAY7+bcD7HLo0YrC5qRFZXeAqlhDCR9Lyt0QniGf3d
gPO22yxuAT5qrA/09iFdVg4BRCxnXwm4t2sHGH7UdU8QF4cfj8j793TkhjhTJODd09T7LVWdNwGU
f6blSj/zYrSbWJkJtDKsprq0jJXndHHXjPY9OglM9lT8Qvg9By/2HACkw3nrLOe42j2cK9lfRr5k
fBC+SuVqFrMM20iSiqHdz39O8VpAgXowZwfyDJ6WqWS8lg+D4bt3spKXdueP5ZUrcrrpCRkOZd1a
VCn9QL3oyS2KGKMmT3Rp+h4jTx++hUWa9fmvJqgyDkdwnluB0a4cyPA4bBqP40/KiDyCSXqI6rrB
tE3BgSGrmvYID8cny7/DgFzLlOyL4dvCES9kG0nqXXBrTUmyc7a5XJdPCcEgumgRrdA9DNaOD7nY
u7j2HRdGY14dIQonQ/FEB3Tq/65RyeeLgBZF6iySRecM1Y8xqzlhFtmArepDrJiMJH0pm0etNd6Z
NiSqFUfib//kwbGjB0Cud0KEfi15ChhL5Rxx3vsSjxAumoZs4yCYYBwkVwN166V7j6z+bl0kgidX
nQXu6xLbJ4nmI00Q0fiB1DE/O+aeR9o1Jif/zubriBNbaNNJNA4IiymMbyDI7b6SAkCMuCkipNKN
gji1YQyuQ2aC2tqebAbNUolP/yM9CCYA1Z4gZWmAptkV8g9wH2v8+39FPzeYTD8XZ9WmkuluKG8S
s9taKlBhryGtey50XPkeRVzowTRqj3hlboLu8uXEqbHMQelht9gvq3UNfmpGQGArcCdjV4mVTTEW
sS1Rv1lzBT2f98mNtCjPTxIGAaAzT0aG4KPxEiRVXwkuLBohYnyfR8LratH0ZhW3XtZ/KK1+VOvS
3bw1dIyqSk4rO5y/ZtyqbuRSFVKp9RN8gkOYim6sxrWnW07RTauYnZHkDACfHKJ7pKMfvyV5NtZ7
60L1MRcBzTrwE3yto/YSb4LfXxSzvFama237EYaMJNc9491LATjv+qRiuJQH1ueglE/ebyPx0MN1
e7ZEkbi3coOZ1hNNONpS4s6jzi+i+L8/W9V6+Hg6G5rhZ2XIjbjahpsGcEkqc4MRMFU1mzudK7+E
c954vcnFGdGTVuY2uCLOg1Akd2ywJzF6mvhKNjISqQdkqIDKbjRG4eL3qWc3sJuovq39Q0RQ5/Jw
XKb5rbnlIJSheO04Icov59gityDioYjYalYEVe9KTCYGBvwjIgwXWhkk3y8smwk0LCRuf4sPxkXO
PFVgLujFHAKOzhNBm9b4ltWRvZRz5yqigQhxXLn2WS5wS2Sqf7S/g+nDdaHVWaq2hUO9ZNZjDMEv
/L0gwzYi8vFBkyLlecpcPIYayfyXdAvYu52ovcvvHwOO5a7q+aaoo5Q+Cxo7NFX7UB9802WFEKUS
E1L+q9O5mO1PsZhkTzEZqsndmshN2vFHSqSOZT1pOMSo8xSaDeSJHRkiFvOEKakXWtA+1qJq29mO
ubL13fDjapJr9cLsmmeOUB2MWr4RCoB9N0kxt8t1K17YKNRPlvgJk6DrEHUf8TpUbFQV1mkxJIf/
bGTP5MNPPM+w8HHI0Q3hVx8t2/QoFYVCijslk5sALBfxuaqO+yuVSZ7W7dAvBh8resb1ooMHenW8
oaQfCF8KKTk5ORfKxt62qFuMrvXA66zlJM4GeyslSZZYvqNvkhizvquhJ/O50s/0guDZQC79XcQ/
dD9JAgTGHUOum0Yd6EspQWQNO0WGHQnlh7iR69XGq9ucCxAIjeEdPJ/h9xDk+ao0WngWcibaSnxc
6y7/UtFCsRADKID8kctSYgMENrh+MVs9x5Ru+UQoemj2ThpmUAc83NzT+HYM9ZMmTq5IcXCDEPhT
zuSlM2tjl8rJPp6bO/+/P9F3rWQ36pLSi5kKbiNmMw3B9971YcNAi4y2d9PUjtlsrvzt0CEMMnV2
jCR0FsjbBST62vQb5akw3VsmNqPBKkLdzQcFmpa/eFZHTqHwiI7RHVFNutZXHhsDowd10oiEg66Y
O0VAt8jnYBCDOMKCSxRuJJX3gXDcrAaG56y12nA8RJ1ssLz9E91syx+iv+LKMC4WNPydvLdc9el8
K6JVSuHRrJIm6BB9DmzrDbatQWIC0APT0OoMsAVUXzNDWXUm5ZBvnATxGXJgJFC68UN3/B773o+i
6fiPuyWGOAVcoHo9NDQD2kBG/FkV+olodoXu3xzPIjCGo8DU9jHjfMVGGRBGxt6ekS+Di30Scn6c
KE2klkkHxydBtdjp3RVAr74csTpsLnfN//afPmcVPInRpJJ02S6xfWLleTujcOC1oIg91RierKYY
bcQCCPWuoEd3TYWI6j0FdV8LPsA1Md/ZCvKwtJ2XYJN29ua/gqYcH0ke+5doncNI5NXtzKf10CUg
tFjMU7M90YVS+3fyxpr6VDu0+b+zjHUdkjSTwMVyU/fg3aQqXnNI3OvrW9gbcHdPZXpq5ran8u3D
8Gi6jldYmXAOkU5pHOxveqUlX7YMiwC33+To6Pw1me1qiuoFIYygW+kjxSdCJXQ+a25PLTHrmuXI
FC1ZpsII1s0IhyqFfT9yRinK70weAy53SajDnQdbf2tIXfokjou9C53skhDaMgx0KGz5e4i3P0zd
aQwoPph4+Ou+JTjCflpVfzLeJ+QYbuAokhcJO0nJeyWW+L1D1fFBLSWhE8sTkjglM0bcS8YT8CbA
oU5fFMv6kVX7rUC2b/B9ORPP4H94WN/kidUUG7B49NYQJofuGnpxWP3IuWTcCNJq3XPMG/fSm2Dt
jqaCZoK6F4QMUWrlvVuznMs3G29SZ9rPy3B2henar2BG1WnGjx4fvAtlSPylfquOjSjFBfE92M2Y
D9yrt/GZoWx8UNrq2zFGAXi+qxVz3LHggecP/V01aoZ8moVP776MdOaezCeDtPCTRP2/Ou3f2Mt4
LUFSPkD+cI8Z/QtlyYS45CMe8bEymWZtdeUYbbWUpDx5YF9qJXj3r4GLgaPR6qdV4Dtiyp4/9Z3e
vBEQtAkPWsDzeSeOrUyVv2+DdkSSqWw+5QBbx0takeqBRIMLP+tFLiHNEkaiYb/XbZsbpy4IqPXU
foe+flwoinUggLYWj5GKf5x2Gu+s+/EgMi9rkLalnNjH56AmizhFT7DkclXXsYr+MgVJhVPYMVf0
dy0EkEyVVGKCLbSYx/yWwRn6rG330hQ/DLlfYcR3pJKHAnjCEWaNIrObTrgnYS+evy4xgQAECxKw
ecmF5o43AVU1L6HHIiMaTSvWH1D0JEQLl9ARf2yVV4sRxk6qr1sle301Z6f48huKzn3nROyT+I1G
8H4EYCDZzVB0PItmxbzdhDpxPNjIV3z3xS3LNZrpZom4oRCP4JmJBts1t3fqnfwM56wTJ4jgQ7If
tMItpgI0Jzv3V5DplDIYbbcSv/9ruKkhTwH3t5rAAiQXfFY3nhhZv2oAp3tLW/ry+lvIPcIt3eyL
BhTioTcvwasoPPmOnS/QBggjaTzpMNFFt87yHXpNNjvstYppZDEkbKx95wFwKjmqqyi0qzAvXf7U
SQsHyOkzH5C5U635z1ILrX5hZzdddyA6qizOPXl6xZbkSswg7/mOsPXp01pCg+2CrgokUB422oey
qXOGhkdt76aEHRdpU84ZMLA4GRVNby9hswrxYuPyOJIW7RWJ+Ywh4HLmi/OXuzptYytp0bE13t3A
ZiZWPK+MwgjTgBs3TXbvJu8vJFLsDi68qtD112UTlJAEeNICHVqv4MIq/0CYA6/kJCipbFA9ryDP
3lKtEyvJFBWMpOa4rRaVuZ7LraSs19xJ/doOeQn+8031nIHDJn5YXiLpZ2/Ist/+rVWRIS7iO7kM
j9KAkmLuR2b2zeJ3UEIOZdV5lnkrjJLaOSNVvjiNFCY6BSShJGrmLUyN6fKRwoFyqYWsjG+inK4r
8nJRZKCmUu0gC+uUDbot/GGFKJ3J+XnJeEcxr782POYmuRGJATJpwiQAgeggb8jRZNWH/kMFdwhE
kyVSEJPw+yUJNuDEmdPu7yQvRIU7ky6NM1jWeeOUaEZwIzoUvQ+6keBmvzffFRNgrwCU3iq9rKJk
wp9HVeUBsWdE6P5zwkyPpFqXeb8WTzeSH4SJBZLaOpRxmfqI3m0U1+ifRmG2jAr/014AQ/GqDzAe
iy5gxhkIA7Gl0Dgi/qOQT6ksLwOsSAzsjxhqorV2/dHnHWl8812ccU3NCzcFuzQ2JsxFJAEJII60
ISrJblpu78sMpJMrA1IbTaHWU+Jbdt5GkY1gfl9RUPUbMa2efrM95h1E/V5KCnvBFPN3+E+BI4aX
16B9FlA2W/Paw/Ax4qx933dwVrCSXUDStmAaules7eF6exk17gaCDltCjrxJxvLgjmXBHoQlQ72e
0X7uiPOcAOB5E/nPGZcCB4LXWzNhoIpvcU98Va/3S/EgMgeFqmwr2TcpI0Zjx9vssvMlA9bkery5
ADrlIOhaf0FJLsn1+3xmaMgXDO1j1d2BoxLrwzS8A65269aiRSqMDnz4107Mqqdns5rxpU9S4iW7
Re+1J3rKBFlaEWf3mOPQyiLVV0I/jmI6Wq6E/655kmNM/78iwpN7foL+3WuZElMg+TP9wUoPqUIw
kaD9RBC0DUzck5e3R7kktWCxNiiglTJJdS8NEXlRFt7g+oSkS5BfH/0qpT9BJFbk3NQtExOWgFiM
jpqo3bGVS2ebkB2/Z2LpkdBN8/h1wDBJQuSYCJYXRuuyrqlElHw/HuDnthm2hRPYHyQJuHWRxo3J
B5nVcaJaJBGnfEYHXp9+m0f9P0cTP/upEwn3ZXPWAtGWQYPERqRJ8Y/iJpB4OQTIIH+ExkPzWECq
llkTTAQVFt/Q++QkUllaYxUbLl388BoMKCvX8ESNI/I0WMxhBne/mTXK2OB7VrkEbRutFnRYuCsQ
BFLgZx0tqC+QJGrDlM3p+gfauzUIek3lVRlPfzxopSmDyhLmxXFgldjDayFZ2bokarWkQmm1OgZF
qZmf6yu/dGpcquvBySPK9NJVc5WVdxNfnQddrezkWtcw+468uYD5rQndGW7Dz9WHxVwnGYSvWpvJ
0Dp46uzgQ847bwRs3vfOsDafcOK9fGzcINXvsj0js/dVWfsKAZ3YYZcXjVuvR+7LNcSDpSWM8NXy
/9FoaXC/iw3e+0ULc/F9H5MEiohzer9ejWlHftGFnuF+KgSqaHlE7bV3XoSljT7aOVqi8HqyOcZP
Vt2THwahXCDWk1If/DHM8zf6uW2uPkN1VIJyF5rZrdzkfLGaYRpp2dsUMEtHjDTk8yxf9SdSdFOM
6TR8sRO8tcT8XAsT0KmoXbu1PLB/rOLEv+W676R6CeAwj4iD0MJ2s3HJYmgj2vnIi6p88OSOhyE8
f0g81nAlKWLIhutyVAAWd765hJugCwPuKBN6K85EESc+JECBNW0sCOOruZW3ukakVzNWler8itnh
IfqjYHrsIRW6QR900VTKO26dGS3nYQgr30AfpNL/x7UJ1P3aNG0SL7/sZL9vZByExCRa98T8lG9Z
Z8VfiQ5jmCehJKVtul9AhYrzBX4h9RvlGiUPARLyxgT6smkSx1rTXHUR65NeK5npjRVQGUGhTSIn
Emx8Cb5Od274j59LC0Q2qtgsFo5lT683iahTSASuiFuRsvDSxtsNoiugE4ygBBnPnD2YrysyvpRM
kDtaRlEbAS3rhQMJZLbKJGebFYmnXKHHIKGFT6SW/ZMKQ22Xy5i8JcM6Z2cVLXG74JxT+0lkaZXV
9hkAfyFBq53BIMaVEjsnVVS/NWh5RTQwioxNw1ykeRoNB/BqtaPye25KRU7RrmT/IuwsEMjdCdl5
MYNP6D8S4GW27/FtlMQt5iQ02NugI2oVQSOPfHVFFTKwgaUcNjGW7vY3HncjmCkL6B8hdI/kZPai
88b/r/zPNxog/+rlrzuj1f1f7Hf3KFLumGkB2GPR455IRLqHvtjdSAsYjwZ5frEiP6fa5raVGxuL
uZmx0Q/fw7s7CB/dbmVvFi+SaBLtwxXnPhfIvwAe0SBS2+rau0jnQ2rBUGciHBChtzKkPIFOJRVn
bSipMWJH8dvrlG15/YkGRQgLqKehBewjDGw0sZgR3kcM7TbverrVE62yPNgstnpzaoRM3CARc2Rc
qGZdSMB1iGV1eRPEXZVKZ2xM+qB+bNMXoYws0ZoFZSWJpCkHioA9AdXjW0J8JUl17eIOvmMiT7Y7
gkjrOu4zYTQrZMasM54gEKa6OAJnZZgrXLkF5tt15aAPZKO6R74stzRxeC6yJyu72KUxQP1NdlrQ
22tE+5pktL/nREFEY/yjSxmEz3+A+o278ZS7OrbuwKizGYdlashIvF31F8dJZV8OHY+S6hZZPxNJ
6wRn/e3GfVHGxlhVLVreK/+4yVFX46TYH4WZNERzWxxGjC/8B/1VpP9GdPpkkP3tjQGPlVsc3I9g
dCWZbt5HlwpazbxPqg4Qcqbq7yRVXwl44VTbIrYYa0F/7eBix6ZMyjSacOaL1xFldd0/9bIlw0SK
3pjJHDR8avLG4B8PUvnfpM1S4ONh1pnSx12urBYe64326CtXhFbgWm3WKYI58YYSzekogzSu9LK7
gPWuSkjsWKHuZ3bYEZPABCD0C/vHEjHmPy16PuaUwhsTmDz4Kih+qtSkqzB3suNRDWoher/2XW5+
QhJ+yC9YZN8HcSd8nlhTsVrvMLyMUqWLrl29iSysg6y4S3hjaKyBwsJEaEJyFtnYZdgwKGuliIn9
M9zwtghBFqZqib/LMex55UAnAsHlPT/zVYU0p3y5kGa2s53IJW6VMvloznd4roeLl0xEEt6iXtFm
Rxy/UU4y8Y1fW4f07TZQGSHoHTx5vNQJde6HaRShCO8XhcpFOUWZHz6iPsl9aWSqv3k39J381JeC
kSQE+hbxewXu9jne8XNB7rHBd2pX7q2D1b/FJPF/MDRlwFGThSMfIWElMBavksYlXpK1xSkHCh9R
Vk+O0yTRLkPCi+EFVuEIJCR+/9vyIwuv9Rtxo6x0cc3gVymn+MSBWyvWBGDiDvJ9mQ/G9CqndIYa
Wj15vGHvMxGcbpSdaW9kd9IhyFLSItfuui2kAQqHflVadPkjEP3xkByLTzApPvlJcZmUqM2vC+lv
NHKgl+fizEcLouon2WTwj26B0Q45Q1SH+imRj42NYtGJzpyXLbZnl4Pcf1KiTvR5n1rTt6ZifhUp
NRBbOMpXlwZisARSvMmp9mp8EmX2kAPeftsrbbc7yxZj4Gns1GZ2LS8ajFpMHlXGc3TVZYJDWE0B
Sel+3pBCF/trdeikAejSxdh5LPkoyAfbVn1k3efAPqqrpzyOPcgJveaRHwf4eEAWrLdjHaSLd9BX
GbYhPAgy8Poc5KD5AGdwQoEXXHpakwCUmjA5TPFVT1mYHbKEb09YAckexQvprkF7keOiaJnyqQw+
A8QanV1O3x8GzcTyFxMqLARf1LelQeQTOKHELSxVW8LzfsVcR1zse2CNFX4AOlEhhIzLdwCHo/Jj
Foxh9CT+J3VYeoSXDHnJ2X6bUgN3vate5nlO2stnwpXhduQ9Zf1m0B35taGSX2K28oaLSXVUDUdh
Br3h274GOn86A+oHcQjS2NRENOoeOgpNBUCeNtG7nYNSBN8OWlpo2VabQwCirS5f4bxaxO6JIFjt
LGjHGXfwJVw0a+gKDnYgoM11MhODF2CtTR6c2og/JlQG5r22aMts2rsGrLP+0y2sxsW6ARNBi3BU
t36i6l4rffD1jITCzc3PC07guS1JavFZR/kwc0RHVJKZRsisLCn76/S2i954gVriOC2FdgzNsBLb
h1/49lGadZkMFAkPmhEMzncJtZCL3jqJiRBeUB0sXuAPccymiR2jkU83Hmz5nWX+FJkGZcsNd2lT
PBPQfIw9cheQ4LoxKbdzMSnSk7ZHgjQexOc8AEm8Dwi/yapm8PDkHW/yXwG3OISsfpynCgXWcc7A
kriaDcs06n5Dl41EFzG08lm10CzuEeT7rvArrbRPIk+tiqH31m1EJ7CG2QeJov97rlxsjOY+eGlH
/sII6I2Q8Z/xp9ESWMGDDx4N2Mj1sJr5+KmXXQCJQqRRJLZfPIxOQi2C+92/UrDSV/Hbup+KijLh
MlR+7bH02zodQeziW7Bh1bcJnq551erlaMvWSI+BIohQvuKZd5yFoAaLRbGNTkPr3LeYwJQWEOCG
dYaR1B0bbUZZN3wY14gqCKsqFO9Vns/a/G6BxMpM3/WNZgqwdvfb/hzJU/O8/QeYFqvP3wY46Al/
MD1BlXzkr7y8DqQ+c5aKIIr7wBWAO4XsmNQrdwuh6AbCI9Gc9M8lbcS65l37QDnj83IdYGJmlp6K
zeXKB6kcha09z5gjyYey6IWufc+qG43VgWjxSNjynrfuioBaxowkLHkCBu4awfWgwJqQPNzCh086
ca+Ec5Asjhqnw0oAQlIrfHhxUu1FsNgHu2FSQWpLoJSk2KpkRLirTLu9Yul19E7jnnw1yp4HSGV+
OCKQvWx7tHb0M41DG0vePjNtsRb+Hl5OheVBgpqIX22NBS2LbJB3COsukAr6MeNPYUfcZBrHXC1o
DvD7B4R1210X3ZNelXyktvuOkjt78mg3INrlb8nicOqtF4zXcPyglRI9KcKzB+Kb4dM4rmLw+EkO
XPOd4rwGhonVMmGfv/OjfNcilI2wERGxf2krVg+oLMgCxjs1qioZ4Pjp6l04/+5zo7KFZsxqlfJ8
7k4qhFw51vt/OcbtdexzfsD/WUJfgkzWFfBvxKtF/409SB/toz6cV+UK9YUIVrdkAAdCK3gkxfQC
W4UQtWGsPM6xQUJatvB3ZgddyLHoic9UhIt03BqWIyXKkLM30QESweoaLDmcEHIyhxlm3A2qwJKn
Ao/utEuvp0qcTaFs8H2uOOyis/JPXpCs51hkds9cbPD8G5/xeF7x+eQI80MNssWFoUmTlpQsZd3/
X3siAcywMuzCY4i03Ly0db1UZHkfx7eNrwBGw6eROCRwUzjmw+PgD+Cr2/YRgJoViHGaGs8Tg6wI
m0bOdIJXenyCYO27jHgvLJ/Wb7UvnaDQ1KFJ9nEVr9Ge7ornvdLba3sj95uMc3ieRiDrxDzJ681U
SJcmyVfhpX2E/tJM9pKJvDNdemoBvrHnmmKasiupUBU+4gfqeOSuhCqynCPnVhbOUKJF3Qa+RU1H
52Uh2KhW3UwNG0CQ8x2D7+paYKmv8ZvUPulFPw1gqxS2TgobEGT8bsB43QRoyYX9A384SSAzEwGx
5xXVs2gY8fuo1MrilRTD2KQqYXVyCv1Z+QcQQNNdwFku0mvmssIFvkuRTN5M/h/rBQ0YviKQse4C
+uVYyYW5vOXBi4SpVjKgoYKj3Lg5BiJkACoA4CPiIW+JE/VUa5fdrzIRAPBOW3WGpIbvFSVSzB4k
iX69m6RSFq7zqJPHAs2IPXDhjTAkRNhqR3ZXRwhCFWKvylm4NOm/j3TaOcZXsrN2LgzCZHk6bPZV
745zHvujf9ASWEOK/o2U6EoY4C680m9Dq7+9ZD89p8fEmVikgJAkYnEPA/FGUqyDde7y6OPZ2eDs
a0vCelWktqvza9OuKNTgaJljycu3rO7UlYz32fq6snaUo8rHsuTUMzPd/FPk3qBwimoRaf9ZKzKg
9HQurLC6i0qnG3J92oofRlfZVwGuRIqwsq52z1kvDoaSo83KpPnL14XKrfn+Ij8b1Hutt43mO+UE
07fc1OU4rheZvPZRC5YRKYz+F09wTPUwmbqe5vyKlacXFHUWk8auJfLU6o0TbGqZzzpVBVIL9afF
/c/rK8KhGFBUfgTSKPRuWBK4PYwWfYgSijTcksWI+MjKTgkMBLikRo8V4IszR9DAYWKFJrdriIZb
qigikETLNjAGpQ8lBtKJFVixb4eJJuyaFoLIA3NqAfjvY+jD9YSWVF//E5WXV8kmJGTyPUrHXLbs
YR7BNoHkE+QbdHQMoLmz0aZKehcQ4yhFzg6/zv78o8Rhx778P/iug2Txf/Rc2fgiUnfF56SeuP5Q
GzJ6XghNRjIeqMSpkE2IGAoJ8t1okZckyROoVAod+aPBG3CPkbdHod8/n92QLfOsnQQ6q1/1eTmd
K2idoBEOwXbMzeuJP695JErsBdi4/R8bls5vgKJOtfT30tvR2RUhxdNNaJjqCU0PMOOMNKjgejSd
L00szhhBZzCtBlYmlDo35RjFfUwlObZrLnaJxGBaJSfre3q9E/FlsJN2t870SymJF8CVnGPHXdm2
WL7286wixvbnPg2NiBP9eaMu33LzIsCxbaJ7YA6hqjpOljK9pEh7EXC5WNPQdYknz/873aTU31Tr
AkGiZ3gefHGbDdRGUkf7SBsqADqMimH7D3jkeqQOzJzYpkNCHWQ7zZ7//Fi5IE/Lwz4tlsbv9Zxa
YsC2CW4J4CxKtZNpz+GaZ4UgBadZEvqUT8CS1r90nZla/tgu9p4jGpyWg4tDBswBlDPjmXAO3W+0
/p1xlyo+ziCzb2+d1KY3RvYmyp0uj95gKbJ7Sv0tzpYOGyXz3/bBWCxdDOR5g7MYW6uroQpWZiJd
ICOzMGsel8XJDp5KYa65k1sgf0uoXtZymKKmTsRaYM3lwZRFXTCv3P4VbOCezokeqUdhjzd9zNxh
kJrcDdmoHVqARPxSrFjMXVBY7tLV6AnQGJ4jkiQi+Y3/OtSl/t75/4rVzN9J2xEGK7iS3YIeTmIz
Df/EbOdh8iqyhfhV1jE1g0iHHnlCmDLrqUBpOHCoZtCZ/FlQQOGnt6+u/me8KquoRywgFS7QHtmU
u1c9ubkYJmsbsRzre1ZBDeV7d1BiSwWUSYQFNgePT5wf2rIDK/mdCsnoVcHN3N4ElKHy0VIdBUxY
DJ154ZdoipYtFd/hSEdsfEGYwuW5lCB06hOFO9iZHKiIMGqKHhTOs1FAjvz1NCN93OxU2fzD0J+b
TLuhLUDm8yY6lVif0u11TR+iDsyNYtyV2fTygqcxioCQe8TEzlUvqHRZ85pJPXD2+/+plkGGXkrW
53yBkBvwKS9G/7k/I3a0LV5X4WzLKQ7P5p3JfWnsh8Oa6aeems586jti9EIusEEDWrdTt6rQwKQ2
P2U+Ux3HoRiVP/XaKS52VD0pROmPRVi8GZ4ZHL34KD4dVaDkqebwq+jA8x+L4wEQ/fOP8CNsq3tR
rSCUqyhTD9uU0vTlkn+eY0NN+rqg/Ts3lRUjP7ZvTlMDdaR5JiVAmRjj7a5EgkZpKfKaymFgTfYQ
HVvzj3CkZFS+a53CaL8SM3zUDJG8LQzf9DdDH8mfrG0aP6NRr51OayJ+KBA5kCGOBwlSQmSiIuI3
UMXo492xNHzlw5koKvPCalAoDr250l2NTHBaL/dAALqc1yssRX9+Ya9kBtnQZ8HgR2DK6w7e86KW
DKKazLuZqYOlila4+KzNvayOZ/L3P/bRwhHehMKvzH8TQnjW86B/7o46X+1yY44+YF9PX8wiuQVv
fyo8LnTa4OdGNYyYiTzvmBuq/zToU115vN9UCEWZzGCIPyzuPI67BPEkaLGFXZ8GNwjUQO8Bas0F
fMPoT0wpCCmXpZq95iNc6985LHPIU1XVEfJm5lt0GpZM9YC0e3rVVUbxP2vWs9AyDnzr0FeexWNI
hFImgjGFr8lKdKE4MaB3uUSxyOTGW7nEfzUz0iTykcZHZ9DjTzYd4+lCGg8AWbtsyjBhPKkveEit
67btmhN9ArG2IqDbL7UuzUiIe/sD/fOZ+kR/A+DcfOkETGQNq9Hh+v4VhguDJNFuinlzCxySyNTT
v9vUPna0BbI4NGZ75+NMPAzLT1u69EZZzx9FJrJNGFhkpWgM61D3j0rEdZY3sFXFqiLq+DeZ0r3Z
zkewmMYumJndIM4TL7r5PuVi/MxJYB5Xilm0OmXDXC36RHQCIpr6klw8s+zQaTaALcyRwBO3bzFx
QX2DLgt3MprQkpp/Y+VY1DYxcRLmXjBu7TdE1MPLV+cf0aYb2siN81fHX3GLEHs2o1oTneIYzXHx
S1YYCIw/WjtVNQWzF43FkEjX7oRn0YUFdMUNfgIzRo4Ldf+c2R5WNx2THcs0WnRg+lGOarm56oyl
61dzhcXRF+YdqzyL4C1cMiZclt/3iT4Oh6dTsv6XN05rViek3qy4lJJNasXPVHI2kr1RwEL+U8iT
B5ED/DeP+bJBng1Jcet3nHKGbs/vnBO/0+YJYDF/jJqz2NSadBH/7GIPRWBKjvAUdwbbBCdIVn30
oDqe6iAMZdoeYSTMGj32DOHEXqYYc59KZEc9SO4sO3uMpoeVQwwvzGiJavDydVred/dUcTPRYZZF
JVVwhYN1hGPMLIXWuaMvDgFu4aeSGaqM/jDEoTHnbIW/hNM4sud+0xSkuAvNPebXSOfqmaVcQjFW
wfBGxTEmHOhG/36veDEJOd+XQlzo5P+l6ilzwh8Eu+/xE+VjXb82iw2+FUh7n8iKNAL05E7gQVD0
EW8vbHoJ/8xRyRkO+6TItaJzw6Iep9KgUu3hpWHS++lRl7AOw4fbGQy/j6Bpo/1HSVBzLvj7ghXH
CrO4s60mTZiQKqpyB/OUnVQYPtCt6ajuin+MeY9lrpqqfG+p5WySj+u2HIMMq0LOvHY5RTi/llRT
nP+010r87+bQk2a1QFvtQkNa/ZpWKfOwFpYBR92cMfIJZwRBF6VViGlbkom1F9v8oc0h/N+clKxb
KpG2vFyOoh5n0vgfU/MbOzBjlkRze8oZkkFKHWP/P1CUhjWUcvkRWqIq+RHWaeoDqlIMmMtr5KIB
zYmqqd2tXoRfRGjIzFYQ+7AlU0HP+5Q1FopHqBbyD182AxmscKvt+o5rYVC+uRIXY6wnOQ4NJRDK
aQ5f27pxYSet4bws8y4k1C35Qo9T1VsMua7aynhKca6ZMeXa91FziuiLnQ25hoiaQpo75i9954Vg
H5sYmM91Ra5wku4iuWCc8yWqpP/SUqKEscH826gVq7XhbfS77n/n5fN6kq+gD3jtpKJUKwjyhlru
Dox6wFJ59SpT/zWS+f6F/s36r21JvtIvGjilkXphrfaeNcxAvC68ey4HjpD1Y5UjxpqhC8qZEePu
kFheGl+3SIzGR0Yt3kKI2NgG3zLcTaJCEGI9Txnr6EEUkXDVDSBmUCO0zdecXfv6onrCoub7MJm4
PK0k0FG2O1ntigb6JMHoNnhy71wZQSuXrJ26jR/0allPbC02GQm2LEp8AH0huh+Qsnc4k3OY8eSf
ZIranxKw1UZfchx/WZaAx+raWdXl1Eqy7seRMQPaGuHgglV+Eu5NfLziJCMo9NfpsjvTcp2QsMeO
c8ps+qYEe1pLDg1lSKRPu3z0mZGFvDR7RPc66uZAdG4T+zdsQ5elhvrk8eyIldBZUr4DCEfOdAzF
cmFvXRXsqb+Az9ioXEAEf+XzCeJ9P8Gzxu0sCkGX5YVdBy0BQONbZScnGFjdL2xx6whAVBfBRd/y
pJ/PnjBpJjC6ItiwtDYKSUXkeyVGxf+hHaDSWcpyOx87dbuemd2tIwtqGBBa3/RHciARSerSvSrv
FeexIpuLBjfYOTR1A9wZqQ4v2YAT116PrrxQquf1ISUNjIkfsQQKkxWeMwA70J48UKG/+tyhJFai
KLu71oDRAQZPqJqli364J35iQSwHqYe07wkW2zn65rsigfgeRsnA29dIUahjgUKg+5uVlH6zq7Ha
iLq4gaQdfGjCmTX/d8VnBcnZQKBLWkML4wntC1E3UhKnIKmfuMoEYDtAm9zwKN1cNVc0XG/YMnE9
BCAbEDOshmHrjRYgayvGoDhUa0ZsozldMZxqfWBzxkX0l3PUqYQYEE8JLVfMNN2VMFblyReoTcfm
SMoGnlrKR/IfLL9rurIdj7NHJ30rUoBJ2qMRucRVJoMPQuwvwOll/dzklbmaIoePHeLnCuiFdi7d
4juLiFkHSFNO07ys+gMy8rKsbT8oeLd9BN/FWmpBLlDoa7hdd/Oajk0KyjUy9SWG0V+VN3ltfdXz
MD04JqS0CGuTL6Bho4kItukP0fenPf7C1bgQfJ2uCgxsgZPdoyeyT/jQX5QF+TXo8CNxyScX1OzR
uwjcWfAD09NIwhx1CJaBKf5fXAy3sV3sC8rz48fXtfgX9tJTVyTlQWywCznSYHztJAvL3+9ZAzqc
RmHMONhOgQfJW9VwUTsqMpPsCWeqWlPLXMWXKDfndwscBets86BwmdOecXmFoDJzU7W4eJXUR29u
PNs4huBpKfYIUsmVS5X7J96aQgx6aelJTUMVmynA1tvCU3gq5sHKOrtwyLnhv6G7tBdaDz3xjipF
VCzy7GOgddBsJ9uPAsQBmQKzLfBagDLT2Wg0MqczJaVCmKCZyWTSOfWFc2scN1vJOVEmikLPKnQG
vsaDxOb+CBAzR5tOoNB0lIuq35G0SqBlfb0PI6U94VWGQT9Wg4NpJtECItsuWAfBEQDS2s0+9EwJ
6DJObkCHwdWJQqGdSNKHhPdjreeI2EkYciGWFAvNwImkzGUHXjD+rqc0iY3Bc1gffTYwQhe1mH+7
y28bvCN2Qe0UEb4hqU5Xo4LcBQR9nNVLfe9/i7SMo+vPWe+jc+kLi4DhWVoxGr923yRA8ZU0KxDJ
hCSVt8/VJ/9qO6wV36TOEAe22OXhXvRfgkh1MK9I3g2kfnTz/wvxryv39eQ2+Xjm6mP9nuP1/jFo
bjTKPodK1vFtly7aAzPMUgXKng1wRKAqpO98MF2kmKIuRtbim5pJ7T6IEh2eX2p3aAUPGKPP0f6k
hUx8lRPSeS7HENSzRh+H2C4ds5uBwvJUkbvI0jK05AAqPB4mvmtlBBRwH9s4ipAU392QNBWm9y6a
Q1DOQ+SoPR42RTTdyMSj+6Q5aERtn/pG9G38HCY5Ak8wDW3marHpeAHMV3J0tqGsxwYVKtvyPSnG
RAYDPXxmfg6rdNl4c96OePLX0RWOzFMmPC67QCCrqtqLSgO8hAkF4Aj+lQq9pVi7N8XW0ghkE1PC
gURgdyPUlSYSLGABoTpl6UNzlm5aO5Yz/VrQFuLF0nWTBDOSgHSfmKIZ5xdtOIsbrGCl89U5/rBq
3qPcTTgOS/8WL2e7ie6NmdIv9HQRI6Lb02BFU4XchR2e8Zqn/GnH/pP3Wlaas5sLY6IHKotyFVr4
K/myF8pyFGiVZsO9o4p4dr1Je4z1BnPfkoyPaB3fagjHWavCgAE8r0MjQSX+lL6v4DZQt1H6uQJS
Ag5ebfr6pXl9vg1TfZtiI3YzfImQyy+K7JGO65cVxH3e+erfozQec+nxlVm0E//mciju5Zm0h+7M
elXWD64djJrzF5oquAzp0amQ03/9EzCpaBB0f20R5KGw9i/1nGCL3ZhiM0yjAjK/bF+RPwaNLtPz
SBw2nRhGC9VpFj1+ui9b+yLK2578Osnyjo+CMzo/Gn8Xgva8xIAnworBDW7pNdD9xd6cCI/gcK2b
OiswF/QXjJTtFpNSZxyxGcgVVOgXc3Z0nAyDPHmOzfePkOlr/QYywLzJhze/zDbKULlOiqr+prwj
UiybORmcxZQqzOYshvXGbSqcdmuuIQdxPmIO8uQKbt2o2f/Q7ZmpiRiXC6k8SNIOPBU+uV0AfWfy
EuzAOix+hxEsnkkiABM4BIVZ691XzqgjYiw/loqJ63VXBJXm+dx0HW509A6EM88n9UjCaskMAW/1
rUM4HgC5NsPnWZTUAMaOsaR9/idyJYi2NOOZN38cKFCfhMUY2x2PpBF7k9CLGkyKDxo9BkD2bmMo
cFLl2LFrUCayZo5rLkOCrSNHbbd9l/sG+xvWpE7HBNXSatDDggkwErF6jpcM3ePqniyKaw0PBbFJ
JTAwL94q8slzlv5JdgasS6W5MdavjJgGdhwyEZP4G1WMS4ODLX1Yvn+kz00eDRAixErYMPjMf7gh
5dQ1fD8ThN8Vxs+MwBNP0yrsY9psvE2L5iWlBhxNfQ7q/Fo0I+4rexv30zJ9z7/e5EyNJmcRd+aK
L8TMmFKRZd/7kO6rWKseyXWH6OKcK864UwLBkYjsSk7lZ1B+K4yOAAYNGbiIjdK/zMv6hzvofvwU
nzMRMwFEIjm9WnUAHxBsF1kna8B8rAp/nU9dg4oxWeQDWVaIXhe4GSf62SIHgwGxtnORcJiupd2z
YxJXN7gbjRs4KV86SWzWHieHuE2QRNN2D/c2mcL+ckcklk8T222a8iGTV1GkIyRs0OkWV2wJhS9e
/Vmrzvcitg2So2QYbu66e5m14SWfMBn/c7xt07R0HzbyHmemK5HxUy35P2nIikU6XDfZHVqsOjM1
skpj1yZHjog5Tt3BqgFg4aIThMEoIolK4Zx/TtJsjKyq9IheqtsqYNXxsBiOL9/2qgS+8GXKeyGU
eNxsDMhaT9Dkft9F2X21NuXPY7fnE2dLZziPzuANWNbU2kOTS2Gnn4FVfO2h8whKqQDk9i1Ga7F9
Tf86KYI/fHe7GKjpS1zAujiO9SEvY4mHlTzVCVvp/TvlDcAVMsJAZ6lf5ifVKI+Uf8WfsRD/A7wF
Wd8nljLM1+O+dZmt5a2cFqlU2tEZDgMCWDwWuq61qoB3JL9YLDHnDQSe3S2TT0gma5MTpe8gcJLo
t5NV6k4cFRiz2LzWxrzDaLmzLQlpYpKNZEH6exki7r2X0X+FrrEIHAzVd6vcVm3MBMOwkg3+OwKG
BnHeoNQbQYwRyFVTSitzjjobLqTHod9MWo/X9W73Gfl2zm1SHgV+IJ8BvoHt9WAI7OL7/9MgSNKH
cYg+ETjjp6NT6ENW/mqssD+WBeN9Mb0duWSxQmwix56jjsay3igLgMqCNPstpbMNSoIfjRiBp7QM
9iv9s3AjKEC1uDCxJQN54KIoQjbG+39xbe+/+4XqZzguWHuYdmmVh0/NchS/anNA3APlywDlZt75
KpGpGpe1fCPvtIRfnDGsc4A5lfPVJG3DIlL511y6bi2a1/TeteqcrCSdEV1oP1EAhXqjx413MuOw
qQv3JsM7SifJDsIDvbeP8z1uwIHbcHUAM7Hg6PcRCVBwcHCNQ1LIt68LgbNecBsW26uc5TJIDJRa
qCa0HfLiIRA1kBpXeNUxeHiXHnGqD/LXVLkAQl35xtK1p690Xh4UR+tfIx3SPsaWq4zAZ+7wMSIh
+k4RrSDx+fzVN0zk48LlLe8yGXKaCftNcKfKF+8QDfpCcgIFxXDpWPvDau9OIzJ6mp09BEz5YN3K
s/kzwPHC8czglPYZHb4Djj8UiGcwDhDxBVCY4TyX5FutUHPDePqHbuu3nwovKbJxA8H1RIMyEQee
1TDWN0KWUQpuVK2/rdt2rsK4fu7tv+6yzQT0RM2zIshLoglRYSs/1n67PaNFuyz0+RHDP6/UWA5A
GBsj8WOf+2nnxiO+1HrBZ5WsaurjJX4nhLUVCI+dl89tv3xGlbIL+0uNcR0m+JbU/IYjq6ufCi59
DkD25Nh4yBm3Phg99TNkplfJ0LSayzkLPuY3WkOPXNEPuv4tqCR9nhK22LAtmAhh8kxFGn9xKbEw
C0WalXviwR4K3nMXqReCGR8Uktzai0r2J/sF/qioAVrFM4XwffCk/p15FS17KasJ0WXctCKURXed
Wn1PeKSIAJytBSgwSdEuLGkKoKLSo6Xk82Ts4PP4uF7UdHvDVT8XUN7BmYVPzEpqUBDuYqcbD21D
wlB8xQy3FnmqsvYPcHUhrYWl1qpFIGQyslvQpUBfw2THtCxGM5X9GIyNY0fDXiRI8NImtExPrSJj
i3f2KzDzAGfbK8R12NldxNdBdlnzfyf0Wgc45yd32eYe83o+mbmq3Y3ez/5EDk3oHZChpkgIkssp
5zR+o28gItYSQebFHkqWKcU631oeAmeAJImzbjAWdDGNxR3R6A+pRuugq7UPb7buG/G9/6bTvG8f
BWTtsewxxudCvJ4nCk6nGyglU/scf6265v+Yi7EzI4tWVvzLx1hCwhWyIUladx0Twp10oSoYtQec
h3Kt1kV20bg5mOxqGQVShqYAoLYWjUZHovTGe4Yng6TWUDW0Dv6plW2wP226iKtQHoGe/czp/L0E
rZ/V9mYh3t5dL/YphPUFaNIJOzW91CD1JSmpt9sCap+C+cDoGqTx6UTyYaj/N3NdsqllPukML9oU
xZr1gXMzg0feWdWUFbEe6BGQUksykqlumZgZbVpFwI+9C35JmnHvbcwQgVcFoBO1FquvPinQMKtt
CxUOQPD5b/vjD6pn7YbT02er2s0F1pOM1sfCzX7xTGmD0QYozw4c7rnmsQEiH7yKkK4lLNb9PWh1
3OiXM83Xp1Vqgf0ywWszt1XYwTH4pi7XhqdIo7hETG8r/t8Hu4OOPT9DS5NCQ4U2IcoVzx2joY4Y
rMfLvLKY4R9CK2UxEHPYkdAwb4FMAPkUWFG3Z7YUcD/aFBdTaB+epft2ZQ4gC8xaE4yT8rVFFooe
L1WT2spZDoodIaIylK5mW8M9dOHafrUNKfl/PqBgQF4imdHioQCVWHzmF8mdeGP4aK/gbvYZsnyq
7/hPQdqGLYLzkihcBRmV6v3PHqf4vVYWGEg28L8RczQQfRDM5PSnGdzLvQPNtfAEiU8hSPj2/WUg
vKymJ1higGY6El3fmQw99y51gCp4b++UvORM7FR2T3FbRRk5Yrtm99U9R8eeD6QWECN62uDnzBed
MwvNzJDY1W7NbShvzGUd/DG6p/f6lx5E+9551ZHn1k+yxeut1vjor1+ULdznfT6LRdPJw63ck5rL
tNUtDJSO50cVVTzQC+lsJM5PkVr4WNZPSy4hm+tqdKNVw4YBd78vqc0jBiZSS1dBhl7P3TstpUi0
pDWFM2d36JA6OI9Ha5Z7Yu+11vlYbKmWRWTVxmwhZWZDHB4q8cH3mFzUa7LMWmS8wghEC5oo2Bvs
5KfbbNuRf6ECBr5ghi/KrlJ+Cm+91pLVyotNEo/2kr0qH44Al7QxWHQNVT8UuocdEvs0vO+4pWEx
6I6uX41+t6WAxHfWZAQhyhAZwSbY49sVNwMP8XPsmf9la+6Hhbha69/lz4MFeGmjJA9Ay11G/P+Q
JMJ/xFEzjZgb+M4Y6Z4IZGzuQR+4GSiy4/C6rO1ZzAKF1CZhUKzJT1Hyhcc3G6OIlqdhootQAiJg
GM9G8jYF4876ndPnI3CTUaynQQ7SKmjsGbA6S0xid81DIk7RMv1pPuAb3H8onJ7EZrSWFyM0v2MN
arZjm44UH0TIjCoR3T+7XaODJnoDANvB2Xzh6NVPrlmP9WhZNtiSPWjdfSim93JoILBiB00n4Mn8
PxuK3pHcSxlx7VVw3msERn50eBASGwlQTpeJY5EGgy0WN/LgjR8Hgsmc974bnR1K8sc4VsnQhG40
91K/NGFvMX3GGiDFANruk7UHYOzwrRLB5/8TBPt3K3u2spr4hXC9x7HNFxk2jSACMhrYeZn3H+wp
Q8xbPaxFAL913lx9hazE9MLkqFeL/5mjd4OBzxVsiIeID8LtJbpJgV8XID268nrD2V7ecGhQzQpa
godeulc2GWZyXhoRs4q/63PLavi3y7QRG/Kd2tvYH0WST8FmHn4wFn1eTHlp9sZh3IEDMbdznqG9
yAMv9tyucIajvIEuTvP8rC+p8WWqbT65+CCq1Zl8ly8rd5TeOpTmotf73Zf9reh9VbJe6ZuswDoq
RCcIuMY+XKrWMDkLX8s0yxkwnyroXPsqe/vGenvI5gkUbkKSw6i/Ennb0CSuP7JfdbgUtg369HMz
bjEHoNQz/ZkCMCeACO8O1GuO1WW7KRJvfjIa1tazufEPsopXZvVXns1D74LYRfkG1ENyEojyeaDu
7atTyjNjnHzLWlSONmtSMRYSxz7rP/+BxyQ21mcHOw+sIN0kWwf5LM/uBUF/AcJrd38DlLns0G7+
rrII39W2PxiN+OyMxfcGxXF+WvGG926N9foi/qRDt+pqx1D2kPlEMWpvKAE8iD8ofZ8rmsZVoEc9
wcOB5xlsEeiqUqg8Yy4gyO+Uq27RmU2FDCCql+i8u53hDOi+CKNp1WI+H7y2rjcJtu5tpavBQFsF
uM1fVKiIGUCiXPUzLzr3iqFvdrS9fvnEGiRy7vB+kOqEGFJUyvDQxdkV+guswaIPdiIJf/P5x0xL
FeXmgbw9u2e8+5thSwCDKGGbtyw+vwxYVP3H67Uh7tXPUpJmv9Afkw3K6tY2ebRkTQkZCofzF1ll
aSD5iWDfHMLg0a85VwovKlSzeg7m10MgrHOawGPzNMquS5X8WEk6cARUZyokHxcgbu8scYggfS6o
K2kCI2xBlk66EDb3Xa6GjxkdHehB/fQ3q0E9R5P3tQ/yLwEsZjG5PWB7MBP4H/FESYa7ymSQJkEr
EAB/Hu17U/T4aTuY1N8couoZlPfdKbvyWJiYyC4PiRgP0csC+2Pgstg3X47QtR5UbZEJegVDtJ3v
CqnANaQEf0osvK/5v+Y16oplF/MwIAW/QiYhQzE47f2hYPzDn+7R6YNQ0/iqzp4laUmlSEsGesQ3
rLC6O9PH6GWykP0ZZ7s8VlFyzts7qDiSNPWSftmBkQRVOZ6IBQnGCwvGTR84YzQB/ANHsrV+EZIl
jETaM7ZLOl/CHIy6KZnXy6lCRoaFMsTQIYR5yH+uMQXIem9ZZTC5LsSlaw9FeDXGD6G6Y9A6zSnE
CtbsR0ryrLiYTAA6sfPCYrWdCFCeyonDTDUsf0CRFwmqAgr3bl8Qh9vydmob5dOuKZhNQLRDPKOj
aWKM+TGm4XpELw4ccc+M5/5eo8T09asB5juQlVjxk/laJLyQMRf0G4d7BfjokGeNfGD94F5vRRqi
+8xmNp/DYVLf7P+LBvV89+pzhkDqyPYgMDMvRAetHZkUZF6i2ZBzxVuSCtE7YEQkmdjHszUacWv1
8R13mCvH1wx1KEbBduofcW2dQU7DuRpMct2bbU5KBF1bkpyVTgHh4r9y9NSE9NjX8POgV2uMHz5K
yUBk5zK/NZ95LQzsADtcoBBU1/VNwVXCPAXIjPSOLEl538J0aGIlGWalPJax87MxjHUXClRdp6Ej
QCV6pRn9pvF6raNT0d87hfUwc1lyFeEKVwxTMjzaj6F6egHegPScpDrLnCtFcgFrgedPm9vGpZG9
o6ZVmGwrPqABtNDXdjtjlfejBgKJfcp9TY6x587cAQvbpQ1Q2Zg/39kfizqnFSrwRA6/k9SpAfDJ
seiX46Y0+4xHRyE2oHkqN4duXIgoVhIQgXkHtjpgTOD9acrxwan/FlLJ7V7IDgFyaXrSRR20Lr2T
cscziO5p6xjK8Fk5Z3Ull8I6Fi5S5LOSNhOOKXX/pfkBx4Q5NuWVFP53ZJIaRgvPOz6tKvtcPlfh
UKKvRXqsIXyPrTuknNkdokaP+NqfTZeLgkdDcPztuc3LAfZXeE36Q8vb4x8z7dVrw/FsP4Z290t5
/tJVs88YG6Sa5Fl+JJLtFc5mzENGjcqEtSg6tpP5f4PKu/tJtSlUvJnbZ9OGi5poz6er1uhibMwm
8sgWHvGK3uIodhrVxHYTNOPWp7WoxkoLDZd/laR1TJWRtMsgLGgL/suC/zuacCX8Tmol8fAUR42Q
IhOfJ5mtXaiICotoZyuIxb6mqkA73tsthM4xrC1y41ZYxXgGT7iMaukCr1m7IpfMlDC5Cqfqmjj6
BTNPXh9N0LBAJOaAK8R+hnCjP/aVoHvJ8A2OMVHb1Y0+lRKcj0wCsBTLoSE3HIIzQDawC8SRTvp1
8+UM4aHXywIdB4lq1iew55QdRXIoJrMckY9fLIqsu5GR6cYUyqzqRa7PJh+xd6SzJqmU3VkN8i7v
Y/VhNbNOPY6du6gE+2sX1Xo0WbAGPdG/6+sl5VSQEM37iahuDai7q0xJU5OLYJikqt9TzP6b0qzW
e1z3Yhl1wKbI6ADpb7PNIW8XlXZr4ZPDYObRwb/jYsfw34Q5BuvQT0JWj74VWS0ktoeMAim3PEFd
2g0WayLAEiCdmdw9EQBw5iECccnTrxRHsr2I2tHQU7crAD57rvtVZ4eNBtdUFkOVDczFk8gd7yx2
8jypCS+DDxe7e6dYP8lJFBrd/J5cThZCd4N9IgtQ0gQji+7N2J1IczZkuJzKkhgepZrirO/YaMK6
3S/SIXDcL3MolAZWEULKFs+uEqp0hX6h5uSjEA7HCiRaBTZK0q1LCYpvF0ICXYR/HafXTOYJj747
vGurFuxADuNQ0MHBdcS830+aGKrofcASWmyYsU92Ot+KMlo2b7bDOUOCbwNYFbnquL66EpbHVhHo
hVD6R752bVjsrQKcIp4a5iZqspeiVQXFAuwwuW9uKuGom1bwcwoJQYVT21qJ3kM7dd5R4ilyKsnf
modsN40V1JX4WvxOmTW3GXpMKA+c0hd/OMkMAZSPlAtrTvx/mltZ9BxChJEIdo9CjJMFmBrOqaxg
oaAUNp1n9sBcUH7E4ir2q+yOdCgAyJgRtzH7x5Ul7Dtvfsh0wDW0IHoQzhFIVZE7w+Moj53byilx
qenTsXjUZMEKypRll6wiTuy/zcz36hYxWI8uuGccyljwqCcs/bYrgjaGQ8mzi4A16A5hZ1uPiv9c
AkYplHnwUh68fLzr+Nf+X1/cLyfisE7uPBlKz35OtC0ZJmZLjDKm4AHZwsWdPdvknU6cjYZhsryN
VpAa09oSNTEp3wSKvGe8ssZ0Eo98cfftNKWQU15ujNkH5oiNA1v4QhGprL+0HnbD2+Cn1IVRQlOB
agBVa97c6KLf+4KmdZFG2/l49eq4q3JYWSsQVpJCzpMOwjBAPihM2sMGEstjWFLDnwRUKEtrZ8+y
0Kiq1ZtDukYJ3wKM4ycy9l8DoxtweeT89gvvuVzqQLLS1Lxk3RXORTFYW/af0CUYCTjbiKwtn/5p
dQME+VxTDXnjXFgfrKpaHrhWN9p+GbhZxln7iXCFnB6WqiSYqYmRbgtgN0FzYDtVUS4fjJNuon8M
xMkeJffaqiFRl0F1sFDh2SQ29eU7brHOhL0GzrAFPIotPjzzjKt8/R9gqTH6EtNqp89u2MbY3b4N
rIrvGjSVqWb+3OS1E8IJEuxCKv3pGz0y6jbU28f400c3wktO/jlhjCTDTLPknWCGuMQb2TozWFVe
UajfMXYypY4knCV8QBiB4EB45p5ZFRZpQVKskM70u4Zjdx6ar1QX8hb2sONCXqTlMWp9BOh3FWmd
MzWIOZV9sWHFakcZyj3ICpbu8vPzph2dpFnPVVxO+eLEM5keb+SLVuw0NWkrTLiJJ+S8N6AcCc5Z
Dw9Nns/OZdkjsrm/IX5e0uAxwbbWMHcsy2eI1X/GZ/mwlovWlSyBDSEv6kRolxbgEOcBKRPWoBSl
SNzWN5QXDaNQX/TvqBFQi6RjodU7HaB3J8Jr9hXcolhc5yznKaPfTmlFEQbG/pOQaqF5R+yO4lWy
v6BE+9XHp/pcQfUg1lB/0B7+Lwj/3In/QVw0/oM+AY9H2Tuu7r96Mfyak+BYsHPxmi7EkZkBe+qO
EE2KqF1kJQWmDC7pzSvNKOwiNq8LFhauCXUfx1M78sCdkU+x3iVqIr1v8XQHTeBuWOH8P4JcY/F2
uYuEFV9HmHUlb8Lt1DZa0cxrO0tGgLMw1fJaXuny0LgYHiuqvbhsEeIkeJSslDjnVYrJJacLzEU5
SSZyuat0l7eAueTwpGURxMofUueC9V5K6qekM7y/9fiud31EtJTx82XeJTH8arxg2z8S+b5y/tMj
6omWGLGR83Hf1hmZY3Xr3QSPa83cSperV0KxN/wO1kFYqkkGhDcTDz1HjgXI1RwodFZ7fD/WEaHF
EWbckBu++DyzcsRC5/5Az9kRaZHpATvS0Wkq5lPa01dp1Riz9ya25+p28M6RoIIsLqLFzKZk5QDF
ZSPzTyZWxlzkMolt6i4nWKGk2DnAx+jVIn8w6ddlJj9cJECC2nG0gC5vquYaIAse9cYx5L7OMQr/
efxj+WbLl3O15uGZx25YF2uPqHlcPS+xPmnjckw9f9SkGXv+NmbjwDyhn7wNQhbJ0sirryP4WGcK
XapLV5YSYgMExHAGfn1041LxPf8zPRHbhQDnE3P+bCBx5GIPHuSrVjtlaZLUe2URzj+tKB9apF51
4CFNaGMQpPI69Pm2gDxbN1L7K0WLBPTKqbNZkmeAtZzXIl64MlGfKrF4fIPC6R4vI+r2xTUeEITf
CNQBxHJIXFuV5ejbhSygqGeigjGNxMgc4kpjSavv3yaZq8gM+zaoxxilk97PougYC3k0zYTGckld
TpnKCzuezpdXzHOWI4hcJ3zlQM4kzW8lQ/7a+NT8gkKvM6fgu26c9lP1aubLyjQG4td+hxFhINMN
xslxQFlPolTmT7edDwDgNanSvYThEiIkbhZRYqWvLEaB1rhEgnHiZECDFCQtMef1FCHQ7YXFEiE3
DCk7oa+04QMDxsihRN4pcWrCinQfEtaqHBYW7x1E8G5XdnfjoYeQcYTMOJRb3wwtedmvidUY8BJp
pQJR3mxng5XcIkDYpdCKc9up1jSt5kcLiHc4oNl2eP7qDDuZHFecP3tkZCVaawmwA1kjg6zZSVVz
S965NL4vIMucODArOCPEjhpdCkX2u2fmx2n9/7Fy/IHWagzgGPzlrOy5jfslkKoB4yqF/NsxsRik
/8c8ep/rFJ6cl3bNbarGNJ259A5uJCqbD7VNdpF0hhwUqk7tIfAGRJLDM/DvKnSqAsYLHwT/tXw+
nuwUzOAzYOUNijIm4cp47am4kjJH2OsHyyejh5zWh1uRvv7aQtB43l7T2vCJB5hqMg9te4nmURMq
Y8mwZDyvSzy+d4pOGxL6V3Cj26LF6OopAp9MCERL7M7YaVbWej/DJvBee3F5yJAWjbnhhUJwZFP0
yL6aRFE6t5lLs0+s9bDr8VO2CYbx89lXkQ8YpYrMoAqPMGHPmv8haW2EWEC0hali44bPigxm1qrE
Upa5Ij3+r0OXziUya/KEH2aZctMLJMAFb+AHA2DnOWZ1kAEcpFl9scMqQPRygjF8UzEInHDnFGXX
WSGMajE9BEr1IHOu5SdRyAEus0DizTV3qLJZluLFAy3aGVknqt3Sxsad5O/iWy+/YG+8+sxVFOiX
aTykPTs3038fjB0m9/an/l0xsUFTcbxJPlG/TZi8m4AaB7ymlDXwnOx57BwysTMLO/rXsWQ+B+2R
5/RqWnOP0j7bGqXqIHkZXF4ouRxaKVneDPCIPKcNjBIaq457f9eMeECa46vyQmPpJ+8ZQk/Pg2hw
PfkV1bDyCAjvso2tZt9YzUnX83HT5veOqqqs7ZstEJOyAoXpFJBcIiQvEEisdwXfd2C7B6yhdOEf
lFcPAFyvTlKU1gW3WRpOKqyKtp0EQXzXswYICj3Xl0I2VlbM5UbblKRUSdrfnNaRNvNISaMi181v
F2ya6pgwTw7IiPfPkYamuEKxuNS5j8VF29YmBdlHkiILKdvy/2DHvUCks2H+XJd3Ilei0EY4bkWq
x823Lp85G3oza2liyEqXlUHwXbp0uwTLwyRc1VuRQVbdJ5ci6e5BjUtpKSLJKrEFMz5+oNE8EiI1
nPjngUcafx1Wm8N7wP9l8sGNixyO4d8dzsjjSPonKxgVjg4LGOFIr/Zmwo8o0gLX4HgXYEqLeo4N
ZYT2zY7c30+bWOcCHy6wEHyDIlBrAkNKg9gvoF0lOyGevjc3+W9gceOLqxNjlBBtV6lLmh/bWt47
uiEjYy+n+WV96+ZJSswj9VbLmuLXuAa2WqZC42btj5Cdu4mzkvpBByp6zUMnplFoMEh/OISOZfDS
aEIGwr9bfvr+CE16JYMK2SWVpfP4mQxCuQkeerHh6Ze76oikmqEZmXVxtfTHDCdteBIsApwx4ApI
bhUAKolVMNM7rskq9jitv4SlD1U/76Z3yRotk8twi3oy/Nk3DeHMuZ/trmYutOtxx01qxsTU1yzH
10sZ8v/qm2NCGGb6a1+4ofi2NbMwJEWo9QQekr7hb5RglJ9k3BALFJ28OABrgNzT+l+eNMi66pHF
OQXEbFIks7EqcaJgsC2fpw7rFObRs78Iwu/+z3XXo+32WRks4ljJNSW3zigVwy+dBboGsVARTymj
S5yRFitmIT8E8RLFD9tX4YYiFr+Aq8Puh1ZUigVnAYwzZwKuF+ibbPcfZw73hHDrFevfHRNYPCN4
4UF0ZO9Xq3R1C5CUshdFRFgJN+c1sjLjAA492SuIqTcnGngQ447DtlqEODnYKt8V+QuSIny5eo7s
aSNVHSAq6prOVtKYArXFD9r9LcpZlgYrNG4NKVz12LNGVts132wrVMT9QAHdHMS7XpstK/IDbodi
iBkR6HaaBKtNzs4KZ5ZvGLT4VRYIUW9+sNYFY2bg9Jji1bE2h60sU/PCfsOZucWscP/Ey8jWCBye
7vK6gssL0HZQ2ekEksv92nPVTJIEaIUayO9jibI+6rRcsMe6JB7TmNkbO/AS7E7o1Hfbk0+QZocv
v8yNkAhRyRE+d6zDHAZPHJ9HyNUPqyLjVCztlXpMZx9n1GR/EzRX+21sYfF8o77AmE9AkiWKEKYJ
TBGyCswI8xEDp7ED3bZkCogJzvL0sO3qg29HzIOiMJRFJ+1VYI8EZCszXtR9Mai6irAWJYdC1yU/
Px4dtcbKem9D0y1/iOUtoaH0ZFTqvjvhHrhUWEB9N+0lX9erSF/ioaqoo36SWyqmTMfvbQ4/f3Ph
MmQMQm8/c+Kn1a4Xz1HTXI5x02iUwd6i0jgxiUBJ/pxTtbjhmV0oxb0Ohyf72crLmD+0VbGqyY+E
IyWIKOddJGvPRmE9r4APEeKH3+YxSZLZaJM+KtkkB1cIFpnI9VImStxHXNKDygEO0UBCXkc/eBRg
v6C71HUOlLL9JLpfUwMXFFDPe0sT/Xsh37pMIaLpSfCMk0C7GLZoN1GCiBrMRV9/NGszxq5pu9Ff
L/snH4tM1UZx4FmE5ziaM1bgtX8nPh6j+S9qDHcpUy2Va+VjgvHq2l2jLZ9XeuAW6WjFEq9RN/7A
tPE7iY4T+ZRNdo78IQZ8iVBbk+sNCWV4V60SwZpJJHKrS0kqs7ME9ZZxIz7n8AMvFb1Czm57xMPw
zDYRK+1/uDIey6gKQjNQu2WKT0EwbsA0Ds7G+92y75612r+pdKdTBLajjw+n9eDe9xlbdWCFCHQl
PwAvAzmwpSMjn+lA2OSPlq2rdp7mFL8v9sOLycHGU0j5syN6uuFDFoSLQeeNuphwGvQ/IplZiYH2
KJu6iknMKY8EjUYt+7zu8EwlVLWxDU+d/nB5/u08tS9WccH36BxbcG94HxXMd3WpxXuNPZMjpEJ9
F61eqw/cojmatFLD57KoTkSeXGLuhP0GvKH+gorhYgpy/6gSXiz/6GPdV+HoechTUbMwe9QRL+ZY
zeIxlXxK+4gPjBFtluBc3SZGJ4qIvPAoTwTHqyPQdNeXXcxLo8Bvx52klm4UbwtLix8CE5afFCTH
4rUp/7YPWJCBkpAaio0S+q5WJy/TT487AlYvR3DjDqXMvlViXoCD3OtaiTC4/U75yGWkqFd07meg
0N7Devh91Lg8w2EKIIztsfmUjmBqXYDMl3x52UM5WRTspyj/UpMwZ2vmU1rWlpRRY3Jx5ZCmIYA6
XHYyvfeD6n5EtbnR2aTEEsjmwMJpLPBLqawY4+75bixt5VseBmTbGJWHTSJJWK+oWV/MsZVesvLE
XBv4sRP6P+RcYymbnve9srgsxArgWUW0QQGmmIZHNe0pW9d6ORg+6lvGyCJtNQUIaz5b4gXvkBr9
UwDC5aSX60PmavIBKFodFLsBHpfRKg5lIWcyCste7pQ7ofkMqv6ZaPlX+3d6M/b0V4FxdIhP6dzi
BJAmIM3m644cLpTeyiDinI269IdjEdNGxcQTLszITryZng/DPiouKOYHs2fA7jb4H1UiSlpfkKaF
s/QUt1iB1ZgyhCH9SugV1AfVPBwOTzXj96paHUzMVltcdwX4dCMlP8cLRqbxchoLNHTZ/Bjg3cU/
TCYwmcVFJT49S4cFda6g54/lN4kEk5isdXe0tdRdh6TRLznp03tZjbs15R86XJq+nUldiur+Mnrq
lBw3OW0PYe2xB8jJ1X+W0t8stlxIxBjRJCPAFdbX8OVRMT7zn9ANQ08/p8GGUt6zz2sqT5Bx96Ja
MmKqM2O0//RjeDzQif9oH2HzNMWDSn0vZJw7nwRwBcpoGKC94BxtYEP+lvKKzpUIQHtIel6P2UPE
/sYCqipx8Y5fzfvVXXSRyzLG8RPtz/oQUe+RiaSE2uTO5Fv9Zk7C9vTkVqqb1dhsD51zmvTP8+l3
N65jstvwcoa4MgC2iQzxZIJI7NJOnhKuB4cZi+8DQxHbrnhCZs2ksdOPneNOn9hECacDmnQXP2bf
ETWSUCf/NfZkvuAdsaplx9jD4j87P5DyePERZZxlU2QFdiZIxSYHZhe53lwmyRQr7r+P24RVaZdV
uG9tSSTMwazdYL8YXa6uH2nm4cNAukLfZLzikO5lPl2a9J2bko22uPObAh4QKy/ub1DlOEdgbB6N
kLvOwdnxwuCvsntUE9coAbDoTgDCnF3C67Q/OO0etT7hlyXY5/9qL4gWZOVufijb3iKpB3guDLAn
jq1JF3NEnm8996fTNE//OKS1V7CYZ+6qkbldiVjoHwcCe3V2mYkMBXUrYnHz+VELoNWTIMrB3ndb
YhJaDB7tWSCHIAvvKUc6XnokqgG+A2FcUXs2toWc4SNofVPGeZ2Qy2hPCderkj+FPWkc7nYYon4T
81clrGhD5CPydtNHP/af1neuIHSncvKi5F+oMlscu2+RQ3bZ5U2kD/kynfLxCoZknW8gCxMmiGdT
ZAdvC0a0iAP3g55FjMYZejyYZib75Mvpg2GncvpVWy6rHNZjJraBiiKj08VCBZ/j4LpzRpZjqn1z
isZwigl3+WvzvnUUbtS/NhfVUc6ALMzVya3sPQEIV7eiaLU8ezVxWD2oCNC9LWBLzb7plAbZgfxJ
TPDBbUnLwqijNcq4uVrDl9XZ4e1yAiOlfKxjD7Qmi8GwkwwpHHxyTHHYGQo5dSa87bhY3K5Ny0Pk
y1wBEY9e1xsfaZpoVn7hiRJCLBrVAI2fDCtma60UfBiq3l2Bh54Tpa8xlSui26ViBtQgjKi+ORko
6ekPM5ayC11z3k+j4wTsvlq5NllGVRehp7u/5sR6hDIMdI5UOC+Z/oP4TWQtAThtIXf1dKvwVO1m
eI3bWfhFyK2jLNUbvZiPwtJgC/Ag0hlak42D4J7omwi+SD2xkCyrEAAmq1VQsAadHG4ZIJ1RJw0K
ID7t49zw5QaSvClqU+8DqORrUEE1WCfNg1Qs1+wZOtLCOWIS0GlozYK1uOFPJcozbuJcEjprBYHz
xQZPaWO3RbM018NCFQwEKkgl5Rk+k0OKqT1iX1aGx+ZRkpF7qOw9eTYcFZfjUpU5z5q3fYDM/BZk
KBhKW0njx1PgLj5Jpd8UiqAfqvLZoBbM04W0scDwmU+3Bmfkay9dp0nWFi4jRXGdRBod1wZplIuv
t1xFQWpIt5w8KMtVo5QjVRtlr5hJ6zeePKMiCkzV50wCmWwVuWJH19u3LmEkca7CjMSwOlN16QPK
g9zzs+6oZvao/oGYYCocE4FYFH4fXibDYGUJB6FbnoyNwvU2t7F3mI/Y9+dhkTuo6E6LyJa1iOOi
CyWQ5+AdSMRqjXoJiS16K8tknnyn74aZeqWWO6uzj3i62WJFiCDK/+hS5vIeBezNQSFhjSXjRrdR
BsXAJW1JU3GoMM1WSiZdYGCzJ4OMcVCY4aaBJ/G2uofiaqBrQtRpm6pw7l8L7ma9ruJf2oBOMwek
LoOsHu9Z1kAKJBVZd3JpoyZQuXRGPxkNz/HWuuj4IzVzhf08ZrKHIDL07IB4moQryXuOI6Jekne7
FFjSZzVzHHBPYUYE8U3BC+CEFvXz0k13uLtJvlPzexyXE3W7XA85fxgcjtyCL003ap6ilrYYvjlD
Wsl8ub3y3HlupCVowfijqgE4a2iiG1QxE5LDOaODR0NmVPVpuFYcfH96ykzFPlCOAYBmwiemcyEl
IyMyaFCcQNuXM6r4ffaiUcvnHLGF22VvEmMHNHrC/bLS4Nd8T15zs47qBB2tk33Ck9aaDsHPAvVi
adQNiRf0dFEOpIs7VsqlCbGTfUfn2Oqjgx29Q/oNBbeRObL5rRAP4Cw2iOVR8XlXrCCh65VdPuH7
FkXPGnQuTVBzBhM3Syc9fOLBOZPPE0L0nm0LY7fG3p9np3AOlSRMAxCB47jkipiXBKkpu3/pUEsc
6PJPSNc4ghXmW/dEIcpaN3s1cMzv+H/1C8RJAtmed3qMjJqUAUgU7nr7E8rRWq5BXElxjyRvcw+r
Ori/ba3GSqAifBTuofGZBIZ6vg2Py65wVvttuHfpqe8bXoTos/yxT+1iTmTNYv+FUSdQXlOV+RSq
CuN0no9oYC90gjEYYcnWNnNEyC78X6LyPPkOK6tuhCOrLdi8ost22xNqQWtweilsLQXj228PtuWP
mjG7o56rayUvV4mpBdqDG25AfOZAJaEhcTZXGH4CFXx8xPWe2iFfxHM3G94SZQLem3mpaDYIBOKH
mnTjZlfDpkYpKxA1PRE/ZQ2XLsRD/XhYh8dvkgzkOgy/0u+o3pcc6KVOHtOoECq/IPbbF2fvhLzF
s5GBz6cG0gTP61lwO1dP2Dji9D5MzRWg3kul38wjufbrnEf5zpG1vu8pfECyooozhyJ6vNk6IlGZ
zPwfr6yqP3cgapTaQKc4Zh++FCE8rdcQR/E7LqsXw4acF+CL11gIeU0g3GnxQET85w4b7JnydWPk
CUmwDt8SZrfM93JRueCZvR08jXLh3ZHJXj2TeXEN+rOpjFyBaZJclvoaICJQE5mU4+/juawVuXeV
S2pFRnC0zjLBbasvF+UvPBvIVJ6UuiKGc0Nrm8/p9jYNQXKrxdjsBjM5J9gcpV+kQgSESuWg4CI1
oj+9cGEao9YFJLcyCGpq+6zD4cCzzgaB3tWrJdPTTMwMKsk9Hkzkgbxt5HgrM/rRVLPgaZJsm2+T
2kvhc9b0GpFNQbb7/est6wxRWh8KZl0BDN41YAy3v3s5jDmIRy++DE30P92RRQKwvWQG7Q/EAv/u
5rsZfkQWUSpF6/fqmX7yjJbFzTRFzWBdUIh65ug0McPp6vBuJmYcP1v5j8vCZ9BJxSXDYU4sMuyS
xXrHjA82MDF8ryiRZrn3x0ZNX86+QBv8bvs2uWByvJumwCuUoMvRgnadbKZjeCjZ8/RZXhY5ss8F
9oTqARpky5Z+y4r7YxHA1Rh4jFCV1K8RNFmvLoNAcs835Oc+/d5Uuj7L/Em4NVFwNDUzr4+Ojlo5
+OgrUHkshxVoRNXsKe3ldHiozgRGFy8HNeNsiSJCKI8w6Okir7TpqM26rRoPW4Hc96gEIUNijgi2
8WzqtDs6Km6c5UtMtgLKVEz7B0ADnS5FltmpesKoHgG3wD7k6NFYkxJW4FLiv4f2NOwtCXS7TLIv
lMySIMQJfBpBSYtN4QCpU7ogsTXPreKnVMpKma/EOCcc4a3N1HuCElvmS2FXdABC00ikS14wcKB/
bZqJPOGejZWWN1dYOnMf/xDG4nLIcoj1yDr7poY5Zox2hhCaiAP51oNRUfWp5CT8rs55Nx7OCS8x
0sJvVUv3HOuV9c8Ato7eCByY/DhD+9m9px7QxL7pdgEc4eoM/Pcr8S9gsXQGZhVIJdUeH7fCBazv
dB1Jcn9Eps2d9hRndm4gmRLsdVG55fgJLeXot06j7uh+K/hsHsVLVRxmD48bxByGrLQ0OUJof/O8
HWvY62iRwmhRP5YHLRhEwsVEwDzNjx7xujyqZ6VAZ1DgAB4uL5u0NDo1gmRZRmC42muANOSBf24S
t1u5yysdfmj+ieyGUoHnSSU/2xPpnVpy9WLrizWNrW98EIOVB+6rKSQuix0sWG6DdvdxRGfBlqk8
O3fEdcFoGoaEoL0Iq/0L4VR3Tl3qTzhwgND30GjyPECFVzNu/epdoNHsRfUa5zckTsQcjc+fRd6S
JlGragAY//1FvfVLwG0g/OFa5ELxlEG2JXX6Hih/jCE9+tMYeh34TBMs4OcEdtCHzill5odggCzx
GjPrORMV+9CIP37lqwk61/2eSQfFaw4ZtUG+L+PKBZ35I4oi7uj5+PB4fYzbJZUWRTyMpSeljQZ0
BDC2OGjI3wPu6Z4hXeVRy+bELHP9F+JA5oXSstnhPZVrC+hz9hW9wh/Irjr5JB6JXYPDyXiMJNOT
CXUyxssXb8XAax8Ti1rkLfa6QUEtRKO0yjCu36R9AwR9c4pps14kLHqx9o6+Tv7XHHQuLAowRZBn
dMSvzzKRalLfvY2w3irpo2IwpBVu+Lsop7eXP05Q5cscwe3uWoNU0pKEvWlGEg90aTg3MKHxlE/K
5E8BTOapTv2zMwytMGT31HonSQO52sjsdq5p1buk7rv8gGEFlGUuf44KVMJ50wENqn35CMaBaM+X
JHlko8lDDeHPIsW4NZeY6aJ/ZKNqfvzRe1g4CKRChFOOUytx071TvHdZeiAzwhDGxsPsWXh4rAXm
X0AbWJXs+7F4904harXgY9/m84ug4XODtOuRb5sWy58PwvFlweXyvgI6OJ2s0VwYhg2TZZOMvDDK
NE4BFYDIpiv0nUI9NkRe0eKLJ9z5vT/ThsxxxDOzZ4T7wNXI5X4SJkjMlfSqCEzR7XIMHz2vigON
B08tNgfSLB0nW1Q81G5cBlyC9fhwywCYMeoADdq49M4kNFM/cP/cL3T/24nRpyf/L0HdIYFQs97C
Yp4C0utbuerC0WOlNgmjtBaL1AqnyTfEiwJJzBAmXH0KhdgAcBVfaokq1K+RrhxBk2CaLpszqlp1
Wm2rc7+LqtXxJwcvTvYYEwCFpr3zbGnPDve+acQ3RrHHb2wzdcc8FOH8fFY57+Cz/rZmz9aZIwPe
HtVVGztpknhTyDEl8zEZbpJ9id3bv7v1tRQeyKfzZA8P1ZqbwxxE2y2+HOoo3ou6KqdB1Z7R/2DG
1Jd6MmsGZGvO9Kva8STCT+CS9rcHqL4y5KdGGObD1lJ4EBDClx8ECwQkXhEFinU86mQKVVCJnAM3
Qr8wKz2Ecsf2v766Mhs1T2PYcM6B994/Wc9AAA/sjM5mFQlJ5n/KvkX3Vz/qCjOBjNo5BUktSR8s
QiW0wb80UPyOloRUh7X0FN2QWWMMsjQD41Frhuf8t9di62NaQNO1XigUc87+giRqNlIUsfyk2SOe
ka7u5plDoAhf/F9qG66KFMg1UOG5xnATPgLQiOMkHoKu5kO3ZOjQy0+QfReF/j6DZPaZhF9V1UnW
c/qjq/RIVu2y30I3bDi+PbtNL35R7mJtVgNMRQxOK22cyDOfV4HeKF5QJrJCvSn9gSjfVP795gz1
VTG5Z13YP+w+GOZ91mAb13B+cqkZPq4w8plxRCDZbOaiEvLDAGiVSaSWAlm+I81Z9kLxFEybFdDn
RwACYA0O0GD1ypykfiPBYwuA4jXwkaFNUGtRudK9VfGQ6vWTrzIZnfgtpEzL7CfwAgfqNyqNLxnp
CsyFVeq0yuIHJlif3ItLQxDdveY3RwfrnSddgegTT75MKkEUSWIgyqHlFKAelI9JNY5sn1okKtoc
hmcjUmfevKtRCwyA50dC73vBfDsTKNZ3XWTbSfBNj2gHr2lNF5MpR9W6QwcEUkC0SpLn5I4SjBnf
2xfno456cEaO7Kw3Ox8qy/MVd7grKq12vbAsB/w2aey9HgLJvFLrzljKHg0blE4RhI4PhBdXNoWq
/WSkH13SQwknhxuekkAwEgHDxSNbbskxAFPytioW6EpvPSsfR4+l2uw8Wqr9QnrdvOmmHQRQcJ+h
fGFbXSwjdGutoz42BIrySVjhCP43ZA1fymmWgTlfNEcXSv9qM8tEjj5qs7/zzCywoy0B9rXt1PcQ
zzpOelTXQY56BNnuZe6jy/ATMhxX7xocPW7lNOUekpD8EdkzV3hFJ+qXZDzaSdNa75INaes3FJiC
sE0+4xtbXAwhv3iqHLxt67ph07yHDB4r7wox0ofDxR1Jf9qiao8XBjYVbmge7kkh5m/0m5m4Cqz6
eI30kVh0JqR39sOILZYTO31gHWn5w8Y2thsocZGWNPujycuqhu/w1aJL1uzIufNGA+8zLqJ0COWG
/DDbOPCQugr57BlZdaQXScdwPV0wx15akLyk21yaRmekSeunE7S8vXt0Js6/61TXj43D8+s/GMK8
DHNuJMLywaTnqxjFprR7E2JXCS06oe/rBVJpXL+5o6jSDCZax8DbPUdl5BMczM53ry9HiqAueG5s
yjLrK+vryeUzyCWH1EmuHKn8SCKcqUKkN6FTF+AehLUg8bJkEdHKxFL1kZfh5CpMNIEqg9vW5ERk
yZKskFS2BHH1H6Q5I/N1ju7P86palXpWw2duYscrKWRxCONaU1XBfH4kNeEAJak+mbr4b+eHuBkI
RWwCrkxmPd03+zyRHvwrYmYmst54rNX8ih6oru8CR3UuN4IW0n4gmbqWszTkTjCoB18ep/e9S/ii
om9NhBgmOPuwaQ/tpoT0pukMyMW9tU1AhmTp+YrHHuoO3MghWAPtVyMuTyvE3zysDH6pWRU0ts0n
2p8SodfOPYr7PWlwYzVRNPKcq86ikwwTcejniGfUNL3CsmmYbhac8OsHrdUw8gn6KXYAeczcS+hx
lkp/1RPjzlLcmz2B9XcLPSmM0pe2MRodOFXWC0+Dhx2g3vCRx+9YiRi68XzBGAFhYdLrEn69v0gH
TPOrVNMEjer/q0VYoKhOpusYmJ7xey4lx3K8b4AG4uwWQPvTSbLZjeWR0f0E3sslxyCK+uEPUH9t
RPxuF8VbJIEPtmKss3hZ435P4Sc4meDPbzl/rHbu7mjPlrBb5kkD1+Xp0EXQrQSnMgcDTNcYxuP+
k+UVB3hqWZ2nQgs4eFjxtsamegTB5qXcdFBbdFerFY6sQnBOHrvjzx9eZYrm6mNUy0CZQ/rK7VNI
0AXqyh3d6/ofAoL9R4BNvdLser/sLMUP5VJYitnMRJdvHTy9ULHZfGScFrRSAaGv+//sKz9vN85I
24atAO93tzAksog8XZr6eiyBnEWHmDVi0HAY8LyF/NHU9J1CS9vWemkBNyYqDblSEpmlUm9oEZpG
JzfjXHJIkVnwqxYO7GDwnRLltNHjO1FlsHJRMHUjCOcVeI9VY40yZCqE9DfMh8SzggbSS9gOfGXh
k0wQnMFJnlsPPhGds8pL0q6vMiPpOFTIedfwP9qimeLr2UPIRD98kXW7cpt/3vl+sbtOwTn4q5xD
ZcYGNFfogOTsqUazP/lsPrBcvwfP5RSSA3YJLI5iol/+/i8gEohQcKloFdqcdx9918235N+Yq7Qp
H9W9zbKCY7lTB4QkvSuMbS2r0Vzcal4lJNHcOz5Wkdgr2rTg+hLWIGeosmY3/2lYZWDw3Jp3WnWP
kIT+X9AWIu11TjF9aEKHM6q32XOgrh2YwiibhL8WgMKZKJgYF7dpJtQ7NiWUjeXEz9kk7RtIHk+K
NkmYX1QwnkNjQOQXvGHC1yftBQdRZY4zjLQUVmGLwi9nhH2ULto5JJ8y65S6yunLxBfMbby++InE
LIBIw/36qkCnNeHMxRW7QCf7FmOCkOL5Wtu/8UsanxeLXMOuxq2ADTFEVgAO2ZMGJfNvrXKtIJq+
QODP0y6oF9rkObp38Ndrpzvql0pgrHpY8F14/PLC4841pgJCaKJ3sOgGTjprX7jJ947tQfBg0hy2
HmQhNUuEAIT2GhYaC4YVC2dCpRAiKwBN8zJmUffNW+/StyezFKqmapcSCdAdNIiIPKghTFvsrXl/
jaDmv5M9PJ6p4H15zYpNjc4aS9r9LrVe+mw7mX/t10Sdg+cXlw8USijrzfEcnpby14cCjkoKZhfo
T3dwL6IRYvDGG8jA22iWP7d6ENJB1k+1ntPk93pjJPg35f6Ec2g367u21Ha3ydKf23ugHoQ6kp5A
QaJu/RVdFFtCxDhN+WiFcRNZRYxc/xUQphsDRC62W6NBgJpEvNW7lSQwCi4aM0ny96jPmyvgGYlD
B0bWiOgs2PXrl+sDrdESIBfcNBdt6SL84CmaEKoXSFNHEQUJXhAlaZs7kPcC1TEEHkDn4c4zppug
RSThsIvFprcoNOX1IY0SJpvd+H999XCsNFdc+h6nlBiE/eb9gl1K6xIbx00cUBGIvAVfiHbIYw+f
AWNgaVYW1F+rR2yCvfYRkPSgB2thlCEzLC0EPFlbGKLF2pKKgfaHWCurxM3U8WGTZFNBInptV7K5
8Ies8EeOPS1k9LePCUBW8MXrLV/iYBf6i+p5gxTuNPB/kpV7nFGseo3eJ0bazBi78/urtRyK8Gi1
vs6CIuEfD0wB1vzZOZJ/VWqoEn3T7MpFKoApiT/wUiumDrWOM9JlufAyV21laOeaFrYrmJ4PCS/f
PnAUpbNDHRzf08UltsyAgxlJJWDnrvpUEgpDPWrZZjxzlKPg2XcDyDae0KEVV3WxtodyTIZy4lGo
NdyKhseN100S34XcQu+czXYAAW/O3E1oviqgfCoj93/1cL+MBYXZO51QI7+bbclXGEzraIv3vcP2
Zq2BGTu0Z6n+JTOLNnaZPyFwV1+xJbE7vpOlxXzDJmVvCTRT63oucanW8M7mgy2U0QUjeWv4dy2W
HNthFz3kCpAhSBXt2LD7RZMgfktXt2TLZS8CxQDjhfkT8bnKWeAHx+lMUYRtxztl/VlwXg0dt+ov
WKGfbRUZSbHBTmKNYc0nwSB9eVi8sNQy9YFuEZgz4zo+ik1YVsJBlfwE+A5GjaP7cswLOpDyIK/+
qJaVBlPuJVd75em+OKca/xqshtwvbTVkFw9K+5q/AbNZv84psStpWYvl+PkjTtbE3hipOGfPPC9y
B4ALn003bLSnhdUVIA0Kn+gayINId/00IlQ/7P9iCFicbiLA53SyFhrsp9LoW1zHu+WeYepLilMk
Teh0jDoagJlvgzKFibLceTmBgcEVFjcwhh0/vHMMASkeFZPTeYVxVSu0XkuPpjOFDyRo2+qnwWSL
GEEy6xmE6tBA7jGo/cj4BaZ2Mwz7GUALkqVymkJsefH5i+Z9W7P3R5ipilatrz6xCJ8Urpp3O9Et
wdKDyGMTvSgEVUAB7tokronp/lb8RY91EBE4pI4oMZ/schznbZqYiPnAR0sWQzWkkllKC3Gg/Olz
+tTLjE5bjBYPNGUIpgwrs3wVwCD0iu+kt+0f4fE+1zh0wAGW8XrRumVoup0HQqxilR3tbakASmay
NaSI5lN2c7XMIkc8gpWaCl6xSoh1OpCe9zioRxwgb8yyg2NZk1tZhTM4Sj086SivOR5fDDQDkAWV
MKCRd95pC0I22+yPR3jxxeJ0n8HsEXQpdP20y5z+/wI2CxDFGYBkS0MqDrfGZXXsmRUeD/fMNP2i
VF3k2C14qixOEmAX6XtgDovJvqzW66aRO99LdnAhD5+CQer2e/rKjWX1iKLvj/61GK2PSCy5dYqL
vOJVPP4psMC7T7ayySpft5jVzvARoDyYWYvzXDXs2VHQCEmYq8UEdpNMBzWojuSnWwRd4b3jVF58
W8XmNnK/kcRcc0u5OeBWHAJB3prC616z9UL0ebzfW1KcswDhAu5s2tf+StlwiEVukF1mBehjghBW
E14rzYx0VJerEr3gbZbhWooMarlWqrVSr8CSTMv3ao3AEWhq8Xc69t2q1f2DAG3m6etPjGCttCsQ
lXagGZ/Krgw5Q8PsR/MYl8T5glKGcr5Le1sCxoTTHaz/nGOLgh1AJjMBX3PGIBZfnfPhu+mvme3d
Oth39kcz18eKOp/gmHsXCUNBxzH1EvKy8mTvuT//kpORo6Kc242QZxqmvWXNmz+JyAmozUzbUHaD
2wdw8EXRp7nxw7A0LJ3Ut+mp47ViLxoSvKmpI0xnX2ut0UfS6I91XSmCBURWJdmNONW+bhxOxGSa
cllcxqD93fsNw939dEUnRWWpii53z8scw/81z+OhWt3/aH/F01aK8SPgdDcLbuw3Th/lkuE4ouzh
tRk0HTNcJT1lH3MuKsTdFLcqo3LhmMv7+fdubb6fOhtnoZJJyHaLI9y9CvhH5pPhMpn1leXcEKVv
8yIT5KF4aAJBx3ntbVivKPM9dJUjpfG72n1epe6+DzbVHyTDtS6St2p/PMaZYI69vcefLa5q1qrT
0mH20Q/jTNQKoSlxOrEJ6cxnZby5uVzFivq5iKrZjl3uS6SyXtD2slQlnN4kQuGkbq/gxSyVVrxq
kfUVMGkfeAa8YyTZIZ3eiCTC4KNMPR0P5oEaxgI0iVvWJPj2IrKJpMrgu8wlNQ297Vo8lfEt11Oe
S4ICBUMmrfXfM5Y4bLTDqhHewvW6mXLzbucw7Vtfz/ZC7KLfODr/pSElfDHf/dWn/6mTyitcU/x3
JKl9Xhv4bKdDBJ43yefWtpb/cqdeLemmhnQG9es3S89/ENOvtp3NiGOcVkqdrlAGow3s/qkZU5yY
VHWWTORsOlmMhRvnQemdeNba+cYZw/U9LnJhuvtWp6gvIvJntAvYtHCQNDTwpxf++OB87sedxkBn
wIOHHiSVBwEUU26xDUruBIxGWSfLvtSn9/YFCsJgZb7d/0EY6BeBscHjh2RZIz97oU9UiXJnPBTR
ALd2kd4CpENt+JN0CRxHRwWhUrH50mcf4lEeVvXwDYtBeCcFGr9XfmCcShlUklMOYysaVli0Rasa
Dm2ZzUtlZK5iK+WImfRiiZodCxn4SwWhbdeHXYL+vDDEXLqeLJQkszOHONjd7pKnxTbdGqmTarHQ
WNCJLSFl5KYbvYV94qSpMioUceHhKu8Q+lYWgckL98jMMjX/4dAS3EcF2x4YbhzR4VCpZ3r/KYOz
fK0zwIRV91+VdEEr+T/gbHCKm5lWp7Qqb9fhDVp2Y6E4NiP8mmxNRQy+SwwDeWlFIyLxFcVCo0EB
v6KbXQLjgKfvk3SZIjBWKf8cD7QyzCc9X2989oQnPpGqQz5Q/bvot3mtkZTxGxyhciB6Ut2U2FQU
aCvhKyVlAEPxEneFWt9gsbBu+Mu+8XdIRjUvwSZxqdzrg4kiKIOKm4XAuyxI3mBZcsdsJ51hQX2U
lxBNiz7KHhYQqWX3mazYAFbUgWQa8N/YjYLVdQqAPe9LNQz9C/5oDrBkm6wPvz/G85HRqu5oLiro
uf1vRyTthR5I4/C8EXJWTmsgpQf0DEwyiJPgXYT2U4lnfmo5hpZISDfu+NATEzqLUUJJJEmWS1qH
LJkDpJtNvpoKxX+F15xHZ3qTMNDAGcPHTuUgLfpUY1LVZ/sq2DKhIrroea04TQZDFf65otlCAZSh
0x0PTmpC4lQqNFOkWcW7CS2SFXWA0qQsWRkNefCuAPh+Jof2LSbLO3jNDBephcICBoKtAPtP66D+
iqqrfGbFn2/iURnsNtCtBElAAmNkfTTDSlf3HFPXv0EgTZxKC3GvaTn8y/oixfEuojJCG5F33iWQ
J/Phl+xk2RixWLd/OpxCTmHJUHGZpb0MsSRmwoMCeTqloDcV0qOwgZC/5JGHATnb73J4ua5XTepY
0x8+HMxpsY73qe7fkrzFNt1AeMOuJau2dXB1YJkzRn35C07FYhUtGU9ZD0Vd2m9uXeXGIyC81yMZ
EqMlfIUNaBZyFNei1UKypKcf4oo4KDMcLKCeJaLUemY6fkPD/b0o6kAwCUlXs9gFdYUMwLOkH/Eb
g/EHrPAtQSaKOjFpU4+/LUQn8s+NpCpxJuQEzzDLMD5vkW2WND9HACTn08z+NTffTWwC5+icrTpu
RoUaNvJaRhF4zo7N5yoPLfFlntAEqnjxW81uzd1ZrCMebDtvk28KexEWP6y2LS1Ay2XDAJVNaHTW
RPhIHmw0M3sZ2OeilKBrzgfFhZ2zfinfhI+mXdt5k6y8ufUNeQFR9Wgg2grnLpIZxmp6sN8w6ktz
vGqImZ0qz0vZI84KXQIq9prU2wlSOzPcakE3ROGbO3cIrQus9a86WmHH2BnsIHDKxN66052q3uso
FGmQwIZ1riMug9kWjtFWRIDjZdA5s+SsyFGH/NddywoQO1QE9NCvmtU10LHa9xHZ629aFaHC0nRk
56AKlY2e7xtVIRUMh1/IIRYisYlgTI7diPXQ07PGFRmVFqcuux5cnX2xbkt9O4Fhq54AdyVaMVQ7
wdpSstRXGcsQdBhpo6Dt65jGqvYAcVq2cSr9/ZL+8sTcJu2JBat5TwpmuOKwS8PTDtGRMbBwC808
a4X/GV695lJTaBotXyxmFA9kd4Ei8xRPmtrOmrqm1Ksccxq8bBp8DcrQmVXVMNZB+qXhgW4X0V/7
RhcxbwhexuagJFESrBJhJ8NB4sX0DGKzoW4gfGuzrk08gSe3p+hUz/G8NdFIO4CFQu3OJ2l5b2Ox
osVJlkpoMdnLkMskuyJhOQoF+rNm8zLh7jiqn3f7ejcBMZ9DzBXDyicdEMf2RLHU4qSlKhSo+I1N
8JOOvyfVTZuKz6WDh3ca9fZF9e6HNmJuf1GYIex2Fzacer4J2pX96AUtZcR9TVLlfKXv+rSY9FAr
VBQ0hhAchUxp9GVC/PfJMbmv2Uv3t+YecJdP/acBLfbs7s2dbGFdJqjZkWBjsM74DFji6GIQprBQ
0CT9dM23sUSrC1TpaAFNv0t3Y+BpFMOVlSWjorx6j0pnLralfi+UuWmLT3XkKSnjuXzmEkiLFMCY
J+gHxtICl30DJahJlNXUiMRybkcBks9LgxvNEhAW3LTaGKlvRelm/99zQam/JkQgujZevj0XQCSk
LYv3YKp55h737ve6bSyu9GwiacNVFEdoIVOafRYIo9+toI2bj9hggnRvCttLH09WvxA7YKM//4Mb
HCTQ6dcnf0T27Up0mMUch0yEjNiED9ivmE2JEx3yYv3c0EAZ+l0tPWU/aoyFCroocQ8Dy9lyWjCS
IkGjNRl35a18ojiLcHLPAr1u147sOn3NeMEwslErvCIxoM40bELwiTxBsozt4mQTgMUlz9mhPSi2
j4aY33L9jGf83uVbRsSpFzbc+p2S1It0U5bUMAaWMntRdxnLUtLdvMqZ4bTvXsuUMzoc3tWPD0FL
kY5BSVUCEOpwU+CT+x/rMaYjnOLvdFSrlxs7rkvO4Z577RHYFmlU9+hOctPAiY+1D6eONRznL1FF
n07XEKZn7+3zMoNi/Z7Wa2DjKqHpQrV7L1/Nzl7DbzoWgaug9cjzmOEkjhpWufjT8fh7TuqgCcRu
ckc5V9UAsOuWlqTOtZD5BSPE+zOy6mCI9g5wNPNORSBY7Gx+bMK9nYUN+raIY4avHZVHD2u/AmKv
OUS3oYLb/eeztGbWNR0NTM0gwvZFCMTHU+DxeymJ7likCKDs4xr+2YJozzF4xGXlAD0+dAcvA5r5
BSldHuVu1667TeN7VgMoGYZ4u1CgzOgZLNkH1H2rSsFEtmb8aHUdSPbXja2RiKQK4xWHGFotMLRy
ah057V6qe+CCZ9a0nf8Z56fb7EOOATauDodpND+Oz3b7ppk9XsKy/5n/EVEcwoW8bK5oIl4vXnRe
HUV7rCxsA6VCvLEnsunwBmlbrp5lX3dl5jpdmAU48wiHEUCtLr1wOPFDMf2kz67YpWRkAZi9phWx
vdFX/u+RJJ6A8YeKg0T8C+b5u6elHCsjF+lzPsbORuJ1ka7WNhyz3213YG2sDiW9dK2az0CNmFMD
62X4aQP+7vim3z3zqyteRz/K4sXI3hPy9ekrxa8ZhsIGjksD8g8SefpYLHiViVimQ30AQRGLem7+
sUe9LpjsBHIRn+DosC8Wv7aGRqqJPVZogLMNLD6po90PoDeoaHgxkl4c6liQ4Fxv+ILH5McJJdUG
7c2KErPbiUilixWjSehegP1Bg4icOER8XnvolVGYvlbgreUY4y+DBKz2isnlAtpwcrISgUxVxfT+
0bkE7ONt7l5UcpZuXrM/v+RI87VEkefOqTmxziE3yS4J9ExEGhSiIcEpmtNMvvF2dFGEm8fPzk/g
LAScCfXB9IR25oTXsMAszcdJ/rboEJiw6haWQRYUkAhyr2kSLOqln8guMFJj5bFe6MBQ7NrDjnTC
q1/hYDP3Z4i02423xRnYhAouL7rNqDh2vri3zg8XnbvEHnWkds11+Aqx4Vwt4ftitEjj29xM0Pr5
SKQPW6Vu1EcWZr4km9oZlrTzduDdakfo3W5bpvLtDyndnSlT90xmjBT9LBi/AcGX8WEOe2aznar7
Cp1R+Dehqb+H3JxnctPYYK34bJseczhLE5Ehm0/+DGRKQKAcHw4xWVKyfuCE2Vqgmg8q9k5EKGFh
zFG9w/yxHh5oA0mWWoz3hCvFkQZDaUHOZBgtFe/zkpsp457UOcGbsj0RVFJ9pYGkwG0Qlf0pRmLa
QZsou202Bwuq7zMS7MJKeUKkZeGoozQa2VCPdOel222qmEh3RTk1Vqo+lvBk5DckQpav82ht6B63
K1Rk7PoO+oTKf3PmAGZMBWr1m8r66RQTpm8GMjKrcYDQ7iqBq57EwWCHhubfyjWBSZABid5c/eT6
wbOVduhmrhWGReYnfPi6CXO9EdAhUZQPAJXgAvsc3cIvcA9tJkWJhnPMw6tr7v1sK2gc42VCba3L
kzM8Q1uKTZSIoPSyv9xHekN83TE6+5wo0gmsjT09YQrJUfsCJUv4n4tdTFfOW6JofryVZ2DB3sAc
f4H3j1OyPoqBLcQQC2mvK74FtRzcHZ4qMW2HWCDRTUZeh1mWOa8j67A4240FFAPVUhBz/OgkZdJk
s//MAB+M/sh3iN1PWfUhjzY971WJfqnAo4MpysBoZV6RXs0KQ7jR8BuCY9WSY1JuomSL3AjFyzL7
X3MeROWJIkfegwdpolK/O8q3FN3P7JPHKC7mEiytDX8QZHk4n0HApjGctl1AYqPc6LVryqWkCGdf
ul5JAC8kc0UQaZxN+1JKhtJgFUfVs+yWRHbwhDruPtPmH7y5VQNtpvrA5M6YF1e0FvDJ/gCWzeyG
Ze1wHW1jOxmxdE3ed+NM82WTAd8u5WIZPiTm+SoDuGZeCk504dh3tLiVOLRoBf2I0rxWNahSWSQ1
4DBGjhmu9vXNtmU6dTRbXiwMxOC7LxvkTfb/lF/B/Ng5Cxo+haVn97zJNmMNvNHjMbbvSQ4kkzFk
w5V54OIofTLVKb6lG2TZbDvluVQ98eEKudEt3WXJK8s54x72dzrHCoPOQVyPZvikom/a9WHL5Y7C
7oh5tdCI0c1b87hMg1VASMyPOHmfmbTpCeY3VcuWYklfiWeUiepgfjqzN1qHn9j3NYOKlMH/tkLp
7GepW+l7fir3XUV1KrPdOFFJ+rljBAhQHSylI7MILAlgywYUHZdZiMcXxi889bLhD83OTP9Q7z3t
m9og+Im7YJdHCw65NFyC2iIJi+MZ0xIafaXCcmpcV4saGs6GCKryDzG/B4iKGxICgOOGE5nxanVx
EQDLceLJim4sPpMfOXwZjNaDRKBUKv7Sp7SyaYGuOzeEjPzeR19yAaW5yAjM20cYOOme2ZIRsOrZ
fkT+UN+sPd75qrmmdNwh6172vOqsrMHKQy1dvG2QmxBLE5VbbF8MX9cyQ8SollSYbRZwAqM9VPRK
gUtpvTIcv94yVeQDxp8WqXxlQ/s71EC5t0RDeefeJRcHvWJ42U5NxL/eg2pZt3qaj+COAYSe+FiV
Nyz7bJsA3dF6gMuu+AyVbtAg63n601vyIrT8TSnFMHmeO4sR5YLASePhti8mv/K1WSZ0PPSc8RyV
zbNoiEmgvh6mBcjiTnjmVLqJFMUMASm3sWLaQgErIIDq7Yc8YKUV7DU8cWsdDTqgn2xNEWbvWPh/
9W4+bw48iDnaeMU3wDxrmxtE5QSWeQ1u/wGDkTZ1fcGPLVXKPWzXzyPfYocq0WVKWvEHKJhKGAJv
fHrWmmGVHYmK8eLg4jPYEzoHYqH9vkILgeNwxPsidMLFnx4h8EW7hiZfmIORyIgk87u2nbDZaepK
bgcfropO9FGvMo329KLfDcU4g43A2Erm7zBGgGROdcjlfAqvKGDyBDGdNQqVXrxEsI3zRhMWTlfk
GKtwA5kLnHIzHWDipLbML+/seBmIJ+PoQDw/lym0CLH1G/gq/ptrExW35bjnEyQqWoOAv9y5ZZm8
4DntMVNKtjPoFpoYkqZzeC3bN7Ai8gWLc7wT18naJRcKeNUdd++e8iDAwdwtTa2ZaepgTHofWsa9
Jh8/GAApEi6Xj5pX1fOz4NFBO8rcDIcvsAeddg7nZ4H5X1LUSIxun2Ojkw5PJuAGmkJgn6uNPS4T
kFvPsPZsDk3Km8q8AdYYWnIfEJ/kOMxXcQYi3ORSaXaGsQ9OTtRKPZkix5mGkGUUrjXH+hSAwNFD
kLthHmqUYEYTkVT5UxVHSXu5A9wMD7hxjM7kAM4lSi+qZC83b4qjkp5xas2SqJL3YVhCy9nn0R2W
4tJ+j/djwC5AvlRPZU4OsV0sq9Hf9skg0AfsVAVqLrKD5NxXaCb5sRQADa8fzThAcyzIwWITKO5B
j8XLLxLdngCECJzvw/MwNTszwa2vzWZlR+IS4HVJ/ktr1O73h/iv1Pl3KGVKGnl9sCBY8lWLqQuT
4NyoaH11rr6UxHR8UCnKjwRqp2IaPPBIVMuwN1SZnUeu6fWTtPym5jp+KYVc2+s5/rbuCzq7avtv
56uppUBo+aDa6Yi5Or1Yt/4mjKgys5iG5D5H3qJnpc5EdZOVV6swd7SWbSXQakpFR4KrbWdQXtaJ
YIOt24Ix5ztcDHPnfamoLkQMB4LQpkwIm/BccsAXeI6uJIuQ8RaHkMbVhMCwZNWyuFR+t5Idws+Y
oyunBguM2T7KBlE4Jdbp4oI9ucEKiaiuvmlvp95QuGO5afzDzCsNJR91hNWCDRPjKGi9U9utcj72
snsBUYN9Ryl+73GnJPVJ5mHXA/auCBNL2nWpXeL2JOx1uIdOqwqHuOY3HEox7edwXm1Zuk3daZPS
7i9nvCmKXpFNBc4+nUA1bkRcubX9gqgxXeL4DZV3efPKH6kK10Pv5ZBItM5LiKkflUgZq/mr69un
gTnudHC2IlhxU0zUoNX1ZYs+JyzSK9CHB8PODBRzDz0beewD7eiyrRA2Uwyo49kY+a7qgBNOPe/M
vsbk/VYcMhk08igqxLjfCqT29+vnN0dlniM52ImQ1Vs/3IGdrPrWKyAKysl0aT7GB1JaqVxGswp6
UnvRVta/pje/dDMpnphK/SCDlXK043nj06N5NT6UW58NHJPRYBVwJR2yeNT5qVxZ4mxlXLUD73m1
dgPnR+tD/iQ257ol6yZd39MXCzzPr9P75/Meog0/v5MWF8mpKX6SHOAy5C4ZVSNRUEUt1Q0DTBv7
ChakfG96AKxas2V6qt17iIeGhc3VfdfrgQrsAprpF9MqqT++EfiAage0XoS7l2il5TcPerAKU1HY
XxmA4xqj6aWFnPz3nus/NZooMHs+ntyNhz8zOCGvqgGggpksQOS1M0bx2l3B6WL8lM0P5qQqwOy6
UPRPXOsP5KLHtpGpMdmu7ZHBB9z/WpF223HlPtX2YADO5aXPqvvSth8nHU4zyTjA93YC5KWDpYS9
KqpDm2eGOe4q3hGFFAbiNbNfSoGTOouBqg0WR1zYf1UVGVsp92hyhhd2aBifH3wdjTi6FrQyXjXj
vrxOZpgW5rtn57xG6itlc3KutBw8wS3MCSI7iIkJI8dd3g4D3nbmKDOa2yK6P71iEZx6rwZjH0yM
ZZKfCm6+cc3oYyNbix0tGjISfAUUX3xu3BWekDD7ZtZzAdgyg0OHyaM/eIFxLMf/VsYM3QnkOHxO
iPWHg2mVRmrAZe4cFmSsCv/fRS6L9WemeyELn6JFLXE81DG2tIzBMRAxDoSIuqOdcm0qf0v9TTG1
Lg0pDXkSFfbX+g9wYqYufr2dyYBPWDpoRcwYhrWdtNshCR+RFNr8bAelrxu4j3eoi9QAveKwMdW8
2FHBisO41q+ZWCsbh5Hpn7jGlQ91x3mO+TzOkLUQZF6D9zeg1bG9SfoyBNHGV3MpW9Q3ZFl+j5hl
wu46EeqAO1I9Sd9xj25V/w5iKigwcMVM8S/DCx1eM9Am8Am7uyRUbJ/0LNQC0pLjkDSqZcBCxz9B
yhFL2kXsrxU0q0pSJX8lewigBFo24lh6ZVnJYtuCVRj9oOShU4Csr8MAItLsFVMCsEuivWq94a3q
Kl1YjLcKk3WBBVoucnpoIdo1DPED4mX6T2VK+KVMlc40S8SaPaUSh1ZCwCxwBDOemv+YmUpQpL67
auFrr/GOEqByIni6p6Zy79jlBNf0RhBWgeDy4c5qpxSlQdAskBOteD0V/9wLWQI2ln4YBub6B0Cp
GIUCJR8iqmAY5AazCC6+0QGWIf4KX/lRzYFgvXaLVElwjACzduZzpFDKYW1XzQT4HnrOh1z9zCHs
5qNp7+//05nP03ETYbbr68mFPdOXgLOACDieHoKfemDhDzwid1Cnxe4z6QcrVtN0AD+0eSktMHtk
hB0YVlQQs/UMXtzpDxqH7y9a7K/KSJO6WEHwp3m4EHaHPPKnMMxPHNSj2xNQ/dPKWg25cX4frdWB
QHf21RAGowtQuZljkkf4hAU4cg6TEZjeoG7N8odYkyi6pBCC49ZhuT59AChDlen3GbF2zYrwASgi
PZzS9i2ERfe92uQ/YOF5cf1dWd0gpQ2GRsiyyNotWXDzzi7t81dpEBRqtCrJu6pmvGXiUi16JQ1J
iF74WLU/pwC+u2dW5qui8pWzI9GwS/NU1WcM25jfOV+R7C9HuLYX73l731B+knUMZ7LBXutOdhKj
vghPUcBMJMch9VTlxTv0VwVkKZup2juSX66ANJ5Jer28Bxo4Nvtw3Ls3Q4ZYei4iBWfXZ5QIarWR
2mekPn/y2Azx6+dM8ZaVkSM7Kl+rkV6mWFWnlMt5Z5ADVGqeJJ4itsfZbNQUd9f3TJDjS36+2lCJ
Edrg+4HGypFs8TaBeOL1GCVi6LDbP8l9BJk34aa+yxHX0TVjyyJv1Jgx1iRvYoe9+xGJvl26MSGF
KDMGXkqbKukYi1TW97bfNIUGIaEMo6LCJemImc8L9gwj8qGeL8oslYwt9JhYCOJ/uINRLbx/ueF9
JpOklgHZ4thUZGK5N4l+f24oDxkOgA3clYwlC6+j8VIXTzTFrW/JO1xlFsIEw822cq4Pp8PXeXOE
wjj/YY8J0aVKsjboo/pjNaWorcr62S5t1pe22c7OhImqUMEHE/FBcJKAnWjGJtx0qloisjUInv8g
+nW24P4Zad68ib1SgTRMihqbQhEEqzU3XaIihHg8TzRxulzLx0HITrsAgJQ/W1gxnjyeA6xQMRA+
6K6emb5q6vxeaCngNp7n9+uDOJrzNcacg0co+3muJZ91EznmZkrolLUr5fGEKTNr4auuVBx/dE3X
nO0d5WMkNQHnxL57QCX6BzXupk4+5SKcAgAWUaMnEp2nHNjAucSmbMEmoDpoidyFw7vUkQ/kHEdp
LsF1kuyI0vGsxbTK0yexWjh6go9lGOzcq0BxmSPDq9OIBgZbWf1CptSniVJzMeJaapugpx9on53W
lVhLXnjMDdfNM5em04gOC6H3lT8niX/oTioYaa4r/ilHfZDeq07Mhtv8ZHX+fO0QHc/ZxqyfhwWe
DuwdSzH2aUoSg92EeDWYi31RgnGMoVhK31uWt5fTiXd9V7ieX4ySD+msPHgRtq5dzJ/CMMXpBHX/
EeicUDMqBnK9T7o5veyZwUntiGpgJbno79SRH6g5K9SbxirLgeztG8QtI4zv21pmR810WBJvpoD3
cFRJLp7nINv4u96GlQK+/KpwzirvUTNl8LX847COou89FGkaqhahnN2fYPPt9hPsmV8OriaJo16m
JMCiHjNBkxmXswfYLvAAs9w+mu31WtzoxTpCXk9FmzrHaU1OAHmkVDd7mGYGqIp6c2zVO/1FsFvV
HVSHCyd9A4oUqX15Gk9xAizlmG9s5GT/8QJNa+0WLWKFeBScFNx4SirXHkP/VG80wtl4UZy0W48t
Ou36YjtXClFIQkOJL50FB6l4qSdME/1Qc41/BKnCmF28UfGHFbsvYtLTAEtUAuWCFc830kTYiuJV
zDygE0k+/EF3jnej6YsjJaCX8cncx7chNNcdPV3JnLiMcJR//UuVvnu93gqFpSd7Z04D3FlpDz40
ds3M3B47cYIHKxp7zv+abYafYPX/Uf7kRBbxzdkMfu3uywNiU+Gy9ELPmlbEYIRWR02nmqVGLRt/
AY/qhw725keM+n8VzQil3LFuRObrTWqz6346ZxdgVnptnQ4mrmTUbPRPtTKBdEKZ0RPQta9nGU7N
ZbxgM/OznQlG1gbzXFbLHJtKcLq/2uhizDdVgpa/B2oCu7e3b0cwSQCighnswZ6UcuTBz+2mK1qC
xt1eDWGGadMyXMbi4ka7IpdchZPWKCR7lDLkLthzQN0QYYbC4YunUkt27MBxMLjhyqTneBbuOHi/
kTXVeWA7xJZMy6BDyNNP0pIumEjO4vYOS60hLKAdTI1LM1pAm9ntY0sjM0zJYWdY3VbpIE+zY91e
x0+ZJ0DVXNtHVy9vxMJbQ1NJlROnr84lgIMImK+PNBzcPsbrrmyCyPzC9vpU4Yh4IL+dhGfaBv3e
UZEVVlVYUkCeAKMNz4DKk/fxx2lQJF9chlUs+jm902Ua9Ny3OxWatF1gkOdXwyDbSKj/kKKGt2Wj
AdntoK3z9/RNPKukglRvCC3q/DUQydwPfKRh6zjln1OboQtT6AsgwZtpdmO/RSLe2NY9zJhBzSGQ
RyauoNgUk3M45xZnpuy2Xu6QY2uTpeUROJ5IEsyCAqMfIljcc9y8DrQYk4PaAjFtmLQjMF1m0t6k
2nXuHYcdt7x7eRdKoeIQgd40u0QzJWIXrFvQb4hY5mWw+7QnzjG1yyAT0AIVdJL4tW8wn2n9CDjg
gJtiaZWjzuFd5ZdyZWDwxxnIDEyIXcOxOBK+vL4SCqst9cqPJd1W9+xmz1PRLos4dhivuPIz1tG0
Vg6mT5bM8hoXUOGR5Nl9V64JoIVd4HL3Xwk4DFZs7gwyH4jGUTniqgO0uAi5eJU2gEwkJFzJD5NI
ms2tfGlauOZKy0CTtWyhWhry1dTRYzR+JlPAfPr5rMWKK66mIkdA7vsZt7nDmUBtQ/tj1PgNoBrG
A3aL9U1PUKcCu42wigifJDdqOYW1Udf926gH608xAz07uon09mf39QkO1WxHS8XXBpG/1PtdQAqy
GSXs7XjYJcSizSaREYeAcbLKcJVdnDvlP93NtBiu8fhJnahUnlwXLuBifHFy6t2CsqbTWX/5hqbh
lVoAHJLZ+hueCsT8UVDDR+XD7vi1f8wgVgSNZLFdppnSABll64dlsNUXfthX44DZ1F70CQD9qCgq
QDdkpVUpqXNG2OgH9kdtRT4rlbuBLy/MTMoRia1PxRme2u45L/+e2p+/ypU0RokFAAb+5+giIXUQ
HP+c3T3qD4eP45EuM2MgufcIRZYLO5I8exNkjHDTdPDP9H2PI3/7P79T3kOHmMBrnYDuVbAEGC/i
f1LJBbMUjRq8tpDJNZdo3VkJsyYxtmwXYTgBkeYAdyNxJGtyiEN+aWMKgXkgqOdWFY4ao6fJT1/Z
CtIreb7NJ4SrdiAvs8Mf/0k4MGrwQVconFEm1Z9KhEPDbJ5FSyzt/gq6teaA8UQgLQNoIsmduz13
EJk9TFso9NzbQdvWMNi5iVWd+FnCPonheGCw0rsEV7HjYcFGFQ2OoR6Wm/Yz2mr5Cizb0MN4lAZl
+o26zH/dNxYLrRnnyn16AvRvBY/pnORPAGV82Mf7K6XAQB/ClEkSh0Q2bI3fJ32XhZlkmR43TmLa
SoPW5nve46htf1mf6oKs09T6StEAdbIs5NZ8h59wGYWly4wBFkXQsCsiZhwArh+TywIDSyxZvTIU
t7Qsh5I1pCZ7CphIKiIx4G8prfFfAHeWApaUJZ4R4J/Wmi6vij2c2i/qY6gDhBUfkWPXUwABbtyN
J/QknZmvzc7205MoxuepedHTY8FO8eVlN9qPZVpugOs9fFmZ98i6oTsg/gg5OoycP3efxgnt8sKN
O4eJG27oR/1fcMBNJz3ltwzFrI/pdNBiGz50mAnSREbeVXxky2UVvclYiHCC+dtMyNvcuqYDZ4xA
4e7FWOKBQ/RoM3ahPvkKYdggR37y8d//ZMAKNf1iKGsddehmg7nUVlkY3PODOqi2c3V4WqJLnOnl
36OlmgQR3NreznBnoohIzX4e2pEJw2mZ7rPZ+2iV01CBf4rk9wlA4m1hPU/srAT/R5ctYHhWyt0E
NjtHfUIMabrxSF5qpef0nBAWZxR0h/MV9xVh9SrGJw5u0LUbCX0S6K6iihh+ObOzhOOn7CD1x0ZL
TIBxtJHQSRgtGiTFIGmQAwDAgkZw+KisCNF2MvnVc9Cbnj1QS/OPBvLzj7GY1aoarqaOzarNl2Wd
GGg40/sGiq+lU1P/PzbFc1Sj1RvZxRgPPMsIj16Jj82iFot/Hlon3lmwX9XE4hIOASAthpyvead9
joy0+lSOEr9K6YBOZI+ODA2d4v3Gf8urHm9HrHmgWUhobWkjFs5gXs8WzAyNYs2xuubdwd1idOip
m8QRVfGepMt6y85MB4JVmWvGcBiNjBQyNDGdaFVybme37NRLzBesvByR6oT85Wx7TzbCRqmDydYD
4Kp7yCeS8GIiD8DtVi3xjxdYdKx5qO5Jn+Lzq+MiCNUc5CTPBfYed2h9nG0ydsDN0i5G/SDAwOy3
+XeXV3Roqd2v9RcIoZVNoRwVT5wQlV3K6wz9rFFi5KCDfEBbiu3CtsKJDesxoaq67/tN5n3jQv9U
j0jdVTfdeLn1piZdTiTPu9nmiqzHZ33sYn58kKrzM9QXPzknwPloNrX8QoJLCCFu+CIATZc2oxo3
3UvuABqRXgaRvhv89EFLCY4Hptm/7PjAwQt/HswAVR+lqSJo1ws0u4AOXCywYECexJMhJVw7mkPw
iFwa8UehFUF3jx+a0elzqgd6lufb2hGjB5wMbeAQnR5VSHiy4PNQGaRgs1Jh1YKN4Yh8IlQ4QZ9N
Lw0oZ+DmINsrDqrydVRkltrPpCOVyy4FGS+e1R/f1VqeSBNJ4VaAQ3cMuGEXnIxwApQMWD4GtBCx
pIOUM8XVcEVjBT4tz/fCI2pVTLshY3XFz6If72X3SIgIr8Q96ROFE8vT9Q3zhYiciaN/Xa0uU479
qHBdGC4bV6JE7P8xvpBOKtc1b3CTgYL5NJOrEY2BHLS6TmEy9h0XASf3BPJFQMjiTW+DY3+9Yn9O
oWQiXMG0dIKeBGWDqh61v9jB3Z2JGgEEw2LDk8/BfuKMlqoBUlk6priszQanLnvAM+U54HeaAW3x
IegU31WBbgL9zUI46DhQBqlAFRfUc+/ZJDMi8gpOUZ3EvPiRPWNsW56K0M1fQK8DXiVNSUA39Bk6
ou78VeAqPVlsuFGgV07tMXbwd9rsBmd2XYtOsjlLk4WtDKWyCupgtlA0/cxCAph7Gx7Gljd5Mt8N
DBJGUCR93p4hSJXTiDNCfdIKv/D2cXm27ejLB/JYozar8IT6R+Wfp4fS/dnQ+ojeKSHjVAH89fYp
jhl2GyK5q5JEhEIeK7gOQmA2qdpUQJBa0ZUqKkP67pKTyLYUZWzdMPWgBYVJXvvsMeskj+wa3gOe
Ykvq6ZAqQjbVjoMb0///IIFnVbrlw/6d3mXaFKvYMVqhq/VVXnFUfEbpd1iIeWojznbUzp8d3Clp
mPPBM59vPI2UpF99l4eUTntkM9DpgNtT+a5BJbhZ1eWswXHOCnYy/BbxROxkEE0QaP27yo70XY9h
JLP4XPJY310axvuZtVSGqOEPjLDu2xeJzuqO0/s/NRKdhJ7IMu05ZTLF2HLXhNr3cWLVh/Lr8744
LP89j3VFnalc5VEyFS82NxyrpQxSr8ftsqRAz1Jd21QRh5yVUMvvljbezXdKIzn2TxeWsgOZlMnp
VOTLuwXlaMxnyoqBq4WQ4xx4NbBuaZLFXt1PT1bI341cp/78E+vmwaHupTpMNLPFLHYSfCUSsFe5
nDL9aVVbLB/Diz3Dw1ko9pSeF1O0/fnTN9xXDmuAfqjrg5NUlO6uh93y1dJhh4omHk7Qg1MXyqci
VgH/tyW21rPWPpuC1gW/OBfaTvx+v06Uupz7XYGIwq4cF8uHhzSSgksbCcfF2JSbvgJsEIu4Nczt
4NhW6CoSgfgqk+yVreuapJ3I7fqy5S1jmGAscp2MkiW7LarDoytHktXlUZk7NoHTM47mtx78MOjn
65tCg4+vZc5AgWe99/2Uve/CqqS+e134pTQh7sc2X7Sw+SAI6PbW/pXDo5UMzNj3PlCW0AcuwZHX
eLlYdTeMTOIwEzxC35c1J4nbSXhlk6PfAsTP/iWPyVYV3NQDN/36orwG3CZf0ntVjpwiFO+Ojw+9
1vCnRLg3R/5syS3M0fBN/5O/3JIlkuT2C7ES+qTM5/vAS7A2mYulMRpuOVxcYDWP8++Zpjk9Rya7
tHWoYG9BCbyAx1IcaEl2gdFWwAjkkJQvrKRniATq03SHz8ABN+7+Ct9jCpsekradf1wOOL06lWX5
Me8tsqSTZUWKxnuR/gJpJJonU2fN/Y7Jcdj6S+vAnjGWThKUjdhmzto7yQwSnExpBJz4cfL4Ak/q
oZ6PI8fgT/h7WlSGD+bt1weSYFjbujwhkJblf9cVZxDd0vCPaoUOiMnbNw48Gq8zA2rDQ93uCOs/
vYPEY7knl2Lc0kkTUgThxZDRANBcBKnxZw/cuScypRYSVoaMeBL7VQkiyO0aS8+SCiDUs9oaP9MI
d/Je3DMd9IQ8zi2I3B0mnLYVl1DTPEfeWUqVcEB4FawTrvi3xGcGqAtpEVUw6mCf6nSsI/8i3Nif
+MpM1TMMYQ/0sH+I6Kf9jZeQwAJfJWOHq4Jn9hJfy53F8S6Aq6Q4u5hS1DuNE3L+wRNnmN/zhxoM
dE0ia0s3eRSWJOtr/kns+g7D5UhcAIN44uV3d5OpiJ1HIk3J6nb4+CmOEQz1QoPdW54+OHvSnLz7
x/gij3OEe/uRih9UkKsVvvNvc/FFHVL/al4/z0LslGVRWHXAtTx4LNTcPQyg6d0V55yngCGvYOpv
ik60Gy9FJd/a8ueyTI89Pw5dxgoZAY6ecWvOZugdu5uupPkshtX72oI6/ANqeXjkdW3lhEbv0t6S
uy+bmalhOSWE026IF528FLurU94/WIqJK9vJNyKI6sw9i9xrCWC2aS1w39usM5EE3wDtFuTvFGuI
CO8IiZ4kqDGknT71chK84kJyRAH410PttGIY818LvKCe8ayVHlVZiFahnAxxDup1xOgi4Lpy4QD7
apl0lVG22nSnHZHbwtXncQnvt7ARrBgoZFUjUqmyFxY8efar1N+2GJRNai1UIQgJAlP4TPyqgl9l
5QAutiSJZ4F1D082/AaycXDKlfb9FOfBaCYfnWKMgdEesMRO13ghCCOoWbT8YTXiI2zzUPrIogb7
OaHUjk6njyLjq2b+9Cvh1N48nFL5IQagj+zdnFFiQbcs/2bGN1FXIczzM/xe9V/jdeetUNR+daQu
GOe5LVbaBSoW19XaFRCCBZZlnUFr87m4yMcJFBwW+OoAzCfC6FX3SHQ5tCCyTr0jmrGPdSed3aRz
5XxGwxfM/T22TdhXBnxSf1IXGlC5sJFG4mvgg7SWwkniHgKCBl63CrqhQ73ehJcnVN29kW2CoHSg
DW5qBk1hj1gfv8ZjwKfu/Bhe2/d0fIhXN1pjL1PSSKqj5IRwIYMkRFfPIlNPyABiOtVl3+9Z/hD+
9dp0ovZVy278oMFxuxelh9or9vjYBWnvH4PcvasW7nUGmmQsAJLe6crvWqaCHqrnE6O6ZepDLZAt
9+pr7IvThTTTSczf99JAXrRrJg6h/lTTOnhK5/sq/rCkJYvkeJ+nwxH7xtFKFL9DS7TmV0+kClE7
MGUeCJMLnjjUkqxIQff3xSPiJE2cYr30qwSDbutPusjZ0BRoDPcEj0OJoGzDFa3atXSb5wTF4jZm
YDinB+C35PHH0zI9v1yHM76I9BsRnWrbLyZqp52iRuO3mEUwDIbEh4Oo67g41pz6BdTEYTaxqFvK
hek9FOqYhajMu7jtdbh0qdITs1uss4Q731YyWdW3TBOqYJ3C5a4SmP6BIOrzBZl/FPSY8xFL4/6P
Tu6TwuhhowdZBnD9xthMml5M/Kbbh54+cdExQ0ElIURD7LUrzq0mPuh8xvF/oVsPAY17pQoSrd3c
FB7+GOQwLBsUGuv6K8GODasBAfl1wvlKNH21Mbkmq0F5+Lc8eLDj38z88KbdJ5V5rz6JYRxPToUz
Cf1ndD+k38g79uWFYfj9FYZBZq6xGi2T3Oq/XXxMcOf/X0JLHIiAuKnTXnKBfw6rP2kxbrT1oWyt
bz1Sn8CodYwj9SQBgrfcAYrCBFLoscN9+oU/VXiS4sTJUW81XJuFKTgmlhu4vKP6Bq5hHFmmK7VP
3WdQ62B9wBfZWjw1U9UacE2PQLZrGHEOqOrPMwGM3xCOwxFd+chlljF3kBQjC8bMDe9qCLe9ZcTB
mpER6wmr/8p5PwclgB4ibw6+tLqwdTTTeV47EihdGu9gK0HQLo0W9tJ3ufMI/SRRtJYFghwZbrOm
FbeeGX7+noB3ZAL5UxpjAY5CQC/8UnC7KABy39ClNqHLCuSnevWVP7bPWrj+TY+l6LS7bMFfptEs
NlQeoUqK3ueuH/mUGX53jKKQM5YfxTjtjFSfPHHwcJPyg2vEBGdVLHW3kW+beQW+MgCbYbv4JzfF
sUiUt7Q4zQsvYTlsun7HS040ModHOqAN7fyijbKia1ztOX4I63skDgKusV6+ASnOeOSFLbO2XJ4Z
CvxLThbItWGXMLUmt7c8vKtyqxGCpVC/3JqrCBlevvvCdoxHI852z06SoCmrxK19JG4WEqqufR7N
0E6I9e1h3uKNTdHqG4goaMcelPmik7YRxiqCATViXHqkRBdduv6FS2eXjYmzOAJJcdLxzLGCf8NZ
IfqKaJpLjU8/f5IeUf8utezJWR4Vec4ZkrlZX1aA/zBb6ejsJdqo5Fkr/QU1u8nTUyT0v0MCePov
OdE3i/NXxNrcqMmdFIkJilv65a5rH7casoRKBhogr03duwH4qThVEjCQXNdtMKD4Do/71HFxlBMH
pQXLGkbuTgUF6JYRg4i7OzpLsEFudy7aqM/M4rOIAZ/Mp0RvBcwhOh5TCfbxLk+8NF/hKjjL72eM
4xA+eiBSnz54c+Ypk3qGz+3i5X4l54aIdfl/+gyGyeLjq+okar/YA7IEmcnoE3OkpQTWBru3StsU
ZThrDahgu02gAg/f3KIrZ9MUbeKAYY5UHJUy9z3PtlHsbrUhEdBvGjHEnVbafhRBdUdYEeHPOONc
3A7X2ho8QBeLx295A/Bads7FOPj6Unn+T9BKklZUuQj7Bfov5VDd40sQSFZ0C8p/QdDZ6/fpJOlL
0wHsl5RB2BeeEocuJL6uBOhLvrxUNxZBFreVY7Z5l/Ym9On22bzy5nUrBJ7ktqt3wRM2Sulg/VHB
ioI5lUobf1Yvxl3v9fFuJ2SHt8TnDJyjPX59zmTjTahl8FVxaV64l+5PGWj1yrjabxdgNX7KjcSL
DpYpYEWM4wNLQ+k6PYxI4WAgmpHygRXvacJa56B509ABDIXzMNmV0Pbq0q6IuRySPI4pwt9B2JgY
eGxADXLObvxNr7g3SW2M5bgP6TPCpFPrwth7kRIlhbsLkaguxIQMllW7Lb/SWR79Yv51V/xqvC/0
Q4tDtD0UB9YGJpts+EG+6b/VjrHCe6flX2xiZd0mW7+TPIf4Ow8J5tUHOv4QB1l6HozNcozyhmJ/
yUQZQMMbX8QivLdDIPp6UtQhLAxGCUNM1q8EIieVxOySiINassg+vv4vkdY+narsOj8S8JfAzNz5
ShQ68OsJXpOVHcMKZ5UbWodnHRP+pNRztCgkpyQ598KzsN3w71OaY/oA367I0Ym9JlRKh+jcVgDA
pA06um+TAEVnhZMITZZ7Ly60uSpKZmLiaiL3e/2cSZDnHCIr6MDgJDuh3gPz0wRaw5A6Ifu3q/JL
s+kyCfXN/nzpe28vGOnSm64JnXljDg+SMZB8vEdMcAsNsk220R4zV+iauXpBXkW0C2cccZ+EkDuU
RyA5sKGjkZNezEh+A1P08CmL3vplT4m7BPBRzJTcS0WlV2jvVdSLUF3QanKmonCgHIIQEGACjuLv
icnkgMy2ZZOvZyRrEAb8X4IXioNeGsqxZV9QX5Op40qaig/foISItuKMJaWPCys5byJGGxezrYDB
AbKQppldZ5NZvKgjaPhwyxyYkte9JsqisEVYZfio2+Q5jAupZVSYR61cyVS3/rKGkBjCp0+Zef6S
F2c5ZDAcHWqfktb3ao7XBzXGUzbNrlWNNz9g9BSt9escp5QBMlgWMdh1Bsz05uWnRwJtZDxtJSiW
yQ9xsLL6b+r3xXdUfAXtsLC7PmxDIbrlOJ6ODsY2pFy/qfF9R332RmCyjPLjqxIJwPcfb7P/69sr
TrjDiBP/SmURu3hvnX0u0cSx8uVWbnfZtrkdk4uPZ1w4Ho1Ofx1OvbIzeIp9++aqc59a555idnha
Y/sTgJZHt+QtDKSzykl5kvpnUsbUhp1GHEvjYsTToboWTAQeZh0z9wK2pPRBjae6oaJuJ7yakAO2
l5H4mphC+rWsmYH/8zg233bf+91x05qZcJiH43y1zJqDqcxFVyh3FHqVf+nrMs1HZYl7Okq5myK2
B2d8QspzEAl/HNC4yHqFuRIZunAyY978nagmxOiYvs3nhLQXfmndooKhd7cncdAfS/oR1sihgmzZ
tn5P9emFxd6DRLvMQZCMC4bGniMzq2AYYKJV1IbrSota3f3jOcCijLn8MNOzFfbTjQIoyuITzux4
JwtZFAb46ah6YyYUh5nfQL8c7hNLIj/zHksUEcz9M9ElGd00XbaaGFD54ALwo1qchUjzVtqhi7Iu
hsQUn1FzQgrlVUPMwPxFmcADnNWtQNi6Xny5BnMHJpOz19JUcb9ijiOyci7TbEHqVHcFrMfqqJv7
fhXJnltHM0KpX3SuwGxpwL71l/3qAmwJ/9LCM7dmpKNe3dnT9+9U0uVWlOdZboIkPkAFWC3cH+ED
1Jii/Ct2ZELgzoJ5URDe+0swtSy7uOIA4IX303zjxeggqhUzjj6u2VE/2Qoc0AAmoAtaYLWwhP6z
VlXTxdCh333861i+8+k4B8k8O+uOZrcU5eWFtEwWkXdD9BNEy5WbELRQrCWu1y5ZiYpux9Sa8yCY
SrP5ZA0EL7VZSJrdqFxfC5x7AR9aiZFDfbvjuXj+CI8U3zG5BvL8jSN5TLpSn35HtOQCVLe0tYz7
rDv6r7+WXbFx2AWwLxOniCPcRE2IiNLfTI9XKyf7e0X5jDsSh+Wwb8xYxn78NQwbJsAnZ3jpRXBk
8VME1wtl5nJOz29FUwL/bMZ8scTHnL+t3e8kh4Kj65mpOvhWu5OShxTi1SAmz/xjVSe/bKtkXrGw
2uG7bM+sM/jafFz5x8Gc3KzSQLo1CnUG9BhLNGuooGBu81MjNT7inOC7spfzVgTAdRiCRxS72++I
PrcwaJVywFGOCmvTQlHUk8SP6lQrOuQPerRvJMv3ewvaWKehwyxrTo+3533I5zJJc4sE2qZkEjCF
UljWOBXpb0tjnewMZznE8p/U21tBbs6jacmbIEKlGNmVLV5w0Lt8rP0Pdnh5LzZwtMElJilS//lJ
MZ5L+uVDuXlHLTZ1Or9oXvrKfP+wWWcQxScXBjgvEBUdHxgu6Yam9pHIxYfErlEP5lMLw+5O92RU
swWzHVsHrBbPF/ZTbsYrF42O403t7a4mT2TykfAtGTaUT8CjQjfpLjpA1sjX3++pbxjsqKy1a0NK
Ttkwm/JlLnJZtR1EDpBQLpJHMUHTUdXQh8Smh3QFJkxfID1XF0rXpBvtFJ9nRBPtaZ2ZLmJVZhGk
1CXqJ+XqybAjC0IOITxc9AUNVU98VQqqWpa0N7uC0X7ELyXPT96zeJI9R+8Rp//AWSWNT6NNbIM5
P0EPA1B6gNtR2ZM4AC56NEl2fKUJDFliUJRA+rqQ63cJlwdOoqUivZtpflbF902KzaV3TuNY1LT0
8z23lPk6CH3k94Ai3v/3uY76mLS1JEBQEAx20ksbDFsoReHfvBRoc62L53DkanwU99j7GxpuE3NB
pGr9GbIQZn2ogP91mX7qjeablrVw7l6vzMlvszNQgsgIvxKJFIbYlvwYI7nM6iPpoibBvEX15God
rodYDVB9Kygkay1wkLkc0PaSRPsx6rFuB84C9fvxcMfkLzGNORzq7Gd8s86w0oU67bLNfLM1Cprg
Mgogb5qUYuYupxHJ8e7ceEkd3ztjsYi95Xb+VEaiLBd1g06C9aAhQ1LWXvonnz3c5twSfdVDcrdL
uZDQzIJNuuJUqZD4qq8WopjkEgDEa6JyM84r28Qd4RkJMGgY1JLGVdSmBj1IMB7yeS4Fue5MNUIx
zTAWIqN6qVBL3qeXhpBV6OQGzCDWPk0iMgXZpJvw1nPPc4yJe+1LTNVweNXkp+oXRUmWyN2p6mRV
jONIrxLE3F6hFrqZBb3ju+AzJwORKW78y/OSXcAhXnSkkm/90kQ71WWxSN5qy7WLalfGuGg4LZMH
WTsiXRJ7pArMHxEUELmjPgdehnfZgn4yvpTloz5CTW0DqpfN7oD7nREIt6ISyT7VpzvgJ0O5rU6r
HAV38W6i9HhbSPNVAucHmIe26RL3VZyz6DLEIM2hMJWyPVovcP3FrbuilUeRIen8yE5FgN10AGdI
0+dbeZH7suOTJ+RvFeLzZME5875cMgr9ufOpWQpKhDMAD9zpFv5/Cx/nWJmgC6mJDMqhVKPWLvzO
GJsahtootXTJmZ9UZflAP2o16NNQHwgFVdQ4WO0w1IIksCKMy65UXOI0yVHOXlAdvRMyvicVoRPe
M7wnjz+fwW4ajoGmOV/ziJZFBLW4k5wefjm02Np0l8+bS10hHxEPn2D3YsWrxy5Qh6mlp7804Q+z
u7xknLOVquBg3mnBhbs3RMigLa/ZLwgJKLNYmwtm4TM5697p6842hNDoGKcpzD2tMSa7KIqAntgZ
dXjvFGx0Y/k21gVr0bW1lv927KYA9aH8KIm/B3oDy6n4Ajx5MSZJsGRL97PCJQpv2H0FvHrE+cU5
Iha7jUjmmQJCcZKBbep4Ol0eNpZ84Y6qMn6DxR9Jdy7EZgPCwRvY3t0JSQOqq7HtB5UUmz7J15Vf
nwcco1Xci3BKUIjvYkXotijDqrxYHlUg71YZ0GACQZobh+MKWlpRgyb0TGN6jBRVijxaoek6sxD1
LXU4aAp1g/HgoR23qtp3TvKvZRJqv7LMLRote6qf6xuygFWoAXhPGiuzoj7W0lv+NrekLuS6PL5Y
KugC2O6f1A4KxgQ8drV2gic58kpzlxLFd01RkUi3t+L+524fzBnyA/Qkgwaff2+rsqe2vQ29mAzn
ad/QQbudec/1R4Rv6MDMQFSTyFB+cHtVfVBolXRTU+Shj8YPt0lFo3TCQUwIyO7e4oIwrW0JgErq
xy25JpvoJqeWFHgmBQXwk5svX1C2y9gXa2lzIMzJUu8jrTWRcI+j5DE4iEHFI2/0Qrsc8qon4I3H
7cR0EeHrivUyke8Dq2Hn+0iRDWXa+C0HUQvpUOYKaOZxVip0dWKxbvfkFLuPF67QHXCD+zQYBw8N
xIuA0XFq1QFWC3EX+cP17v1H6XJl5l04cXS0STQV7XCxCvQ/+FMiMtX2gwJOKc9ulIRJFf5O5Rqm
8Ub2L7yEfO0fNjjIejItlY3nDS8uQdZyFWqfqRbesQ9Q9A1lxkzsAORCB+qK7JcVPwZLfeNbSBJE
HOhRAb8Z9YnN4kyXCNDvj1ApxWhc3qDVw7kurFhr4uqrvf4JsTD+oT6t76CKPMFWiHpHB8halVQ1
Z1QsYybEbhbpOYNxyh9rUdyG6gxnKW7flPwwos6/e1Il0Ie5pFcK7kVmWQ1tESaUKnDSJjQa9zYA
5GrtdnZWNorDIujFIUEr/KosAjKN1jmfPAYVG9ZGX25nVbXE7ORIQuOUnk1XIoRvFy1iUh25Tptw
aZ4S0Mg6yb8j4knGsMhckTWz5QMyhlREgtkeDlkDuJHA5Co9vX17BqTMQ4l4kA48c6Z8pSmDYiWG
FYoM4Q5cwSThipF+5Ma6KnZmauSQTwkoGEqk+NoQO8gKl/11Y/140cn8LP7M4iQKglR0pnCL2G8J
3tDLFjD4MT2HgbUiFjYAJBXPufLZT0tJLLIhoriT10PF1Z8rFgAa0POn19fT5sFfS5UF9N452Kaw
qCgBAuUUQwVPpeI14HFmUgJiAwfyVPVAon4J3TIiD7Lf0jEKvcI0nva7UraUOltcYD8C0UJXHGgI
X79Mds5DuAiejol+4u49oGvIfPaY8TSpgvln2KWOnufM7D4Kpvl5Od1L2HJV3k3ImvxcYwXbgE/i
mIf6gG/+MdZmzyiYkTDq4rfWNh5VqTdqmqn4GxY6ok7/A4XtOJnx3k1EyJ1A2EWw8MzfrYDorta1
kS7pbNFGPZokT4fHkCOtGmTnSsydj/yq+E0Wj4rTeNSAsGe/uah/8iCH7J0FyXFhQKzjGelOsgLD
aOzcjxzKWiR3eZtSUs+MzN1Fc4gszbjqAbFhGq7qqV5D7Fktrt8aX2EBjWtDiPm+R8eG8FySj8rc
1b9zirXt8Cg32NgnmoezzkQEIWGQ16aAxaMhvjDH4nYP5r+NCrXQzNa3VrDEMTYsaoWSjVQfkjdu
SfIHillF8mzARdWvkxuLN8u/D1zxBJQsK7O/RtVPBWjpjoZsl/xITTTj3t4UMI/LhjnfZFq4VOA/
dpsHogCCUbtanyRni83sXE/xqQj2CVzuu1sNosFgBzuD808ajKcheLksJZ1h1jkIK9t6vmBHmKno
Rz2DEpK17OK9ZqbKZxvGLBsCyIu5yJQ7GzkFjledHi0uNQVDoXRT1+lmohXa5/KbJhF4EUiwT3T7
cfvYyPjXWAm09GWQN+afIlVIou1BhCNp0y25gpqpGswDvHJpSBwP0Pcy+eNFtnhO+5Y2nvEfIEch
e8eRTx3dWdfj+PJgbBIFrtV9Ynb7V/MjwE8Yxby463zFaCH3v3GpdhuYzjjNerP0aGh4GOhuye4C
k3ls77bM/1lqYkNzibK0exfRjnlEJ217iHUFuTopekXyw0RAj+jM0SneNew6ZNrxNt0pDtGEe9e7
SMA5vG9jc3lOps3DiteiRRzNI2hA9R1uOntcmtYQdFTSJSihUKeRq+GfWoC9D3yB1vvQmL2Tuisf
1wno8G7B1lFYtYJPC5YppTg+YcqL1P6MMRAYLguNS0wqMIshMYO8NO9539QRjqmhRSdbsFvFbx+n
CNjDPAl029zbg8fLiLoeZ3bP9cbBeK5IIJlUroAmgnInVDQ+zp4cBBcUpoCLSsFWUSFrX2h8yw8H
0oiAsqGboR/7SHBQeGs+E1gNivteY3FhFLxLd/WTuIZI97Z0rVV2p3xnVj772xr8fOnEeOtlbE5F
gGVlq4KFSEpEu52Rso6jUUga0fAME7/ExGwsh1BsK/TBzW0/zh431oQvW/IMKCV5R7ezs+oIxmd/
3KKxqSQvQQqKKdQzYH+Xm2WNr19145csOSXlhjSBj5q5HOLbsN1HKrvA4x9xlXHrz+S5CG8W9SQ/
2tNHEEw9C84Z2td6h/SCo+W3xH6WIzRinyyRntJa+f7jqlHLY83gJeYbDFt8PANzIZKRGcGF3Y8e
Lj31OflxFe+9sCIHhMm8X0k7ddDxIwvHQUfOTk1nSB/0hi/xz3hua2Oh9xFNwHOqmcvNtCs6SHpN
2xcNs8Z0y2tUpyrn203rc2/PtYAbD7hiYOJjWJXdp+faPEO2gddzfLf2XYm3euz7tbWqdB+802YX
P83TrCDq5jXh/s7tPGVEVKq9EC0CUkgunYz+UnoE85xJ5jL2eoqYWe+SiNlgVHdScxYuSSAmQMlF
TZ5YdYinqf2p12DV3f1NEEc1/dcs7/TiUi2OKDtweW1XYuAiqGn34WHfkSSoW7IDN1REhDHQpW2C
JWATunIibrGlEsEvIhXuvrgAWgfv+xSujXounelPVEjtjeLDTriC6I6XED1yGN93AoKlMGeVwXgQ
UjHpFnD9fO7bvzjZjC4BM6D9kDIXRdSqrGtZ/DUdnHAWAS59s9M95z64RzLCqmKc4AaupQKmvKIf
sB2Gl8MkAe7T2Eb6Qq25/i8mwfr9Gqg2Ddzi94Ettb0vvchP4jr4KYvv6ZbV+LSaM/8Dj534eAd6
H+9bFbNlsGWI9rUXk9mnSTCVESX0QnlZJH9wh0ql/PNgfNZmkInKUJSc3h4/644HNbnLi2iUs9XR
HHkwMLP4DKc9dowBv9kl37+ylc1sccTadH+ZCo6SF4uB1eCtlOKyCuop9W6HsXcx98bsL4CeAOs1
kErb1/GbGDxOOeyPRBvrK/HTecdYfIBlsZWNrc7FCH4WJr7JbeTWI5Ms/6a0vyE00+HdzjEmimea
74mYdXmEzL7aeZo1goCigTS+lxaUUQxpr1J0lyqzCIzpAQkpr8bR/sCLQAVliwBdOrKVysIUw/bj
lMqmtK707YsRKzOt1mfyew+MWnpw4VLwgEWkTc+6iA6ePaRXb4LSKncG4PuTickPNPRhcy6EdylK
VE0EwfxVh0ScSrP+E76W5RyhuqTQH0ffwWwP0EhW58KGmhKGYDn0ZMTh2sKlBYowBLq5cSa0V5YW
OE1Y17pa6duGCOzRCiqs/r9D+61c1z8mMr7Km4K2KleER1a5kLODTQ750TTEXWDH2IjL5x3nkD/M
Z0Re9dlyyi2qO2ksRVHXJgHIXrYU+z3euiuX9LJ+snjDiYQh20xbKD3nGiU4YznlgabKwVtYWZoy
WAkaZoIL3qo4elTsl9vkecImiAH10lrMeC0Q86kkSa47FxC16ZefimXoJSJyz7GG8tBuWK67llOE
934Hpb0St59BVUKR4hxJi/TZfVEb+WXlt4qoefdAFlnpilT/XOFIZq4938mjhcs8hxtiIhiqgZyf
IElu2TxTaIAxJUHOxt9NcGI10/FWkBTAkWLy1aPp7gUd6FS2kRjqrjjwo8JzRr/y2kasylSTjBsN
tZTIrHNOgeI1HUp+y9V003ytjCme9hycLbYcUkzJHe+CSGdEyERWVNdbKnakKEpvPWCLq3dkRn61
81WD73sK2TMptVf7jT0e3Ne0PWad7USqNbUebXlHu4OsmNeGJ4OxJXlcC1TEIndjNJ/bJYXyZ1rN
Xy8PqDwVpiBoj47AXtQLTLk/a4QWAJSlKmyND57E8xFR4KOSYyJ+eQdOJbUECyV1dfg8vw3zzreI
W0S9Yd6F7DqRTpedEOlNNsBDKgflgQfFY9NruiGgc1HZhhREzKAnVOfE+UJ6VjTixhFy8YiosIhm
aFFaXy5rFHsMnxHcfHt1dS/74pIAAFv0SlA7/QtioSJxLDPQorEik1dfPDgXyDe0hsMQzN82gJfw
fEr8PZyrUYuDp00rBi1Hri6StwPYYZkUbRIYW8CGjDNZNRYdPdgRZ0VV+VEQ8q/SuSbsgJyJz66T
AUCDH8+HU1c7GaU8glUb5gHgnGmhrczJbSRbVzjOTQdcrgWCO3p/ncI2klSURyylzmG2EqGtcW5/
25pJQUiUNaXzbW+APNE8N5ARjOrkY010G9lpWaHajtFzd+47dKs4SrgCj0jhodehL3yBehT8rca2
svMXEGmDi+qf7MuMHrGidSNTJ09jXdy2vMvfU6VwJP/yAYTWNGft6+snRsOVqURc29fvKGOUEIwW
/FUCoakm5GZwe91h08beLjAF5uTbU9ud5AyXtBj9P1wyXwQlKXu4gOYRIFQuR9QJcD/QKOm64IzN
WDUjbNvMRKF10z5SlrkTz0GkglsPZFHBV3+6Aw59nfWrjbDupLvCay6q7AvuBn6pKFPpzH3OpZtk
mUI4+hsRIxxLTw06ZAqmv14m9m5EkSVMbNEQGbicXR2VUn9GHMbcNvooLJ45filEnheVTWVUpFQr
W9CqP1mCLpSHMPgtTG3GqobC4APj2R9BiXNm08rUGdkWG6kisGwuzyGlWZEMc/cKeEvu+t41E+7H
OY4L/SFGT6EVSRxs1dwDdwhupdKRZFywjpX+O519nVC43OGj0m+bjp/BwHqX5Z4kljxj8S/VWMwC
cA32kCL1dVrOxV1r9Za9Rx0ppG8yEq27oU1YUFnjI0asz8o0yzc0EQCg0ujZvO98gkEMPHhfOblG
xshMkTsxPKAyGniuUwRozb4+IzskjaIIl2QQ0j86g0GKyHbbndpScHPu45N8OLrPv5aqIrpTNQe9
cVLEmn+f/1TUZJNBsb9GKhcagWqG2hLh9TLtHWzmXfFx5TJEHUyaisTTNw6Shwv90QHuXTqoLcb3
03q+TPkqomK78tsvxywlKsK0OFwAThbpN2wx1bMBViXbOpc24cpud/t8bM+4JLCeuKm9cia81zeK
/qoMOj8Z3/J4kxPdOqQZv9ZOuDHYFwAqTJvIIjGpuivOLpBVPy8T8s7M0BO4ADsHmONIJAnilvjI
AUqafZkhNjdmFKw2ONpsRHsUSFBpkBBXNNqAc0m0KtWCAiL48xSMfqwXIWHnJPkDTRvtHASvDjNs
/Qf9flyAobwjCwVunULdS3QTTpAG2HDj7GMRQXv7WpHNLtL1DrzIrABsSwkIXq1j1BcAm6/bCQWy
4uo8WrfybA7Lp1Oo2n3JmbrHd8r0TpqaMAoDxwjJY/+NPOeMGUg2ngauGydtIc2WGbR7oP1o2Ind
kTElj0ZTpQ3vInQHmDA1EAidb57HgvmOOaB9yIJn4w9EUYGSzmNk1xdVChwZ/QCAdbq31t82vnvk
aeYfQeEEcUY566n4YhXVtS845Ry/NUghUhFbz1GPUvJAGChtfKHhPs3g4dagh/6UYsjPH0anLo7A
BQpAKfB7EFHsWTgyMKo0SqOaWuhCaxg+8B3mmRMEiFuXK1v2SHy/iTWgk7ZKOVctQwS/dX7fuy+g
Wz50Z5gzeGc6B3dMwusQnWwdXRu04TkzYM2n0yiLwRTCJS2W7Lk8Kz0EgT3yNYNXlVWNpdh0THWe
6KDbMaENFevoMnvTaOW+Mk2okki6jW6oNVvf8VE+H2njnw+ZCKC7EsDK1T/Pvdsph7EWmT2erAs8
MXeIg+26eDYYL+gorbSd4qXtkJ9KRu1z8ATjFRg8nHhQdGrIPQTUKZRwxcy5Ob58ZijKfQ+bLUC/
KJ8xLnZeyD//MfUYZFu0z/0QXRlV/k3Q2nwbVWnSSo9ibrv17v0FTVRAOUjZVmtEhG6V+/HQtkdR
Vnz3cvd1O8Z5HuM4UbdykjUp+UwkKDmTYHubwVfQS46u2UcUD22D0VL5fMfzpWoC96qHhsaD6LyM
+crGsIsKs8negOg3DvpZ5kFqE+c/OQiOK2wSajoW9RnY/Og2t+OLIUtCUujIZ+1Vzbyzxxu3XyFp
nah/OvukmnG5VMRErLKEpGYqrKDHW+o6ZR9JHtzAzb7eTv/cpGQoIi5AorwafuIrloTCdYebgZPQ
EsXbf0UhOS5rwMQHtJ5Xa72xi5ORzhD7ftTmsqehpN75pnhIsVc6fs1XYZjnbhLglGKgzyC8PEh3
BeCqV+VReLqCGr2EEBB/4dTzryf4DAYTlZ5UoYfGnAuCFkCKAjbScmtqdzFdFOyteZojmpgVXLo/
U3xWB2kuXXzrJQULCtZoR7lQw24xHuOHkOta4bzb8EToDr5yl294AF3MG2VA+p9tDLXiZ3HemH0q
QAMVKmQ6UrMRizOiv6xX/lbad/0mxbrJMOFNk/1//ZMtbQ9o24Db/UNjN4rnAxgAKPMdEhIE46nG
PGn74QafiPelK9F7MlMKzyTSLpDVWOqKkLo+L3TOefEjk/sYNQKLRNfJ6v7k0KBZPpxQ4MDCLDD8
m+c0vYZIgla8RRFRFs7UBw0gBjOeZN6Y6ZFHKzsRR5HEMX1mHsq70X2gq3BzPuACtHZS7iTKlSBt
MB9w03bguFix75Gew6zxqaMZL+896+v3BCeAwN5VKeS21muzWZf8ClX4FrNmv0/HCmCUBQGXWidn
8/kPP3vHvck9gkRjwS+CHcv+lVLfu/0JlsKMoKdD/YTnSEx/FB7nT8Q2bRGVw8sseOGUqZnwebr+
impyxHgtewtaiD6Ngcq0V1QGe7HlU/Z1v5tF93aE9Ofh9IBVLXi8b671MJLHlf+ml7jsEtAQuUqg
zQNmLHqLN70XCjiQoIXaFX8YZbWYTwzi/NeMF95UwfJ+GSGOtugUa+12vFJuLwQlSeEelJRZlL2s
ihWGA+KOp4nejWn/YEsF1XmAWrUi5nxTkuKIfqse/0ankg9iLtmVTpsiTNA5bkmlOb+41LJYoFXX
Jj2bq6WcWwGqkoloZ728qMareC3g1OboviqoI63jbm3JNcHMRiwHcJFFustu0bepS9j2k8zJZpKM
k03nzBP26eThSnxRpKxXkZ4TZyV6w92qivMCoDxSwhInQAluLSb5HpFy9WtfxDJjxPrgXND1jAln
9W+aNqEdkjZdBcV0KvkHWWe7/SHbRgTh1vlELSE//PfhtxB9McmBH/Fk5xofkUBhwwNBMXVtP12x
GPq5JZm8eDGCKSx6k5XSKqnJhOwefqFq/kfNGPxXb+aMmE0wMrgyTNDPo2CBDIszjxBK4/6Yfiaa
gJHpgEZdJJLS8TPIMDZqnkElHw2udis0hn3iJOefN9F+FP9qpJ96miVNqy+3XnDPHVciarrDEGSQ
cs+QstZm5Si6024XsJZsM65/LGnih7+ekS/b8nz/Nm3qyEEbpHYBUWgsierk3N8lPUvjHgXaJ8au
ePh+m/WLEtYpg+jWgmkYE0v10CHb1YuHesgy6W/shDTtFLGQCBK7dUIugT4YlgyNsHB6ySj5tJ3F
irxgcOrtw4WUiPUYh8UXClk326nxWc8dXIbo8vqpA7VAWC4nsYeoPj3nNPcOlEBoxsbV4eQiCCgg
8gqjAUmqwFNPb51uOSVrr41fdIejRO4sxciXpv/RqWbGZaB5cfGQf6j9V2c/dr86OCJ1rZ6CEj8n
H6QG7Nh+HkP/h1frl9xSGr3nRoQbj85Ip1HOeywaAr1ylTaG24xBf64yl9u8Ewl1Mvxixz90UgUE
3r9goV6nUh5T8xSxxYTYp7fo1YL23hB3iGz6tQoIkN2SdA9uEZfe19xVd6VEW8+BevMd8OJi4xt0
4FNE5pCzpvtt97DtXq45J18Ke3QqYHQe/s6nRYwMM9wneoMAshdABiV3cclD9RFcJ6njdMtsZmey
vgQon2jSl9AAx4GWGmUvo9znYoUENoPyryzlimBIX+/kfZOn/2ASAupdw2WRuroGDIuFa+SJAeBH
0CXsa2COBcMNfcQ9wqHaHoPq2jiE5jyvDB0uNENz9yR/Gv+KMkoT6hA3ot7U3v+6xQJdfLogMLvx
05GgDZJBrsMd1YICypBVjX6lt+q+g3kLcJ1lq3GG3QmMlpZsY3PUFo8rogeOg0yYbRLXgG6SN4P1
SheHkYxmmepaFuiJrfKQtl2Q2nCNsGzXU8wu+5qbrxzBsyWokr6HldTyLZdlWfUUaa7BQ7szjAHn
AP6DFtAuUCOGKQzzgBOmXalRUDy/QaP6AEfwTeYcAE20x6lfAPnslEheBlGqm+daW3Xqw4ufNovQ
YqCWnhKvzv8rUotB5dWnQemmzO9D1hvubEguBbshOxpe508vwV4li2A/mHOaxhFWPsLNTFmrC5ph
yokDTRdtOwUqxteiVBOLufLnCu3/u79Z6WsDx/Kjif/Zs5PiiU2zGldNvIbB8pEdYDD5PbOM6mSA
e1Z5q/9IjeoPRyLmUjxfLwCOdakbjVlm+bgi15v6DLQRWKdBawqUYZy4wREFOZxazwVjHcXF/BPj
8I0cqNl3/ImFSIst9pt7m+XE6BBurlO4gZJamqD90urqr+kOyZH04Aj20w/wFodZNkuoDokHzUaq
whCEDmjt+y+kw/CpXz6BjYOb7bvsl1AIyUgBD8CcxuK+jgn400jDh+aYEWf/VzrtGZ1ioDyIPRB8
LibyI+W0KC3jAi0XKvxGmAuOQLK5BTtVJkNi3iIDQPR2b+oEr4SaU+DeLBo6aEU1eN16dxirhAJH
RTuIo4WanrnHY5ZB2bvB6mydXmAZJL+KaRNpPFhgVCN5POOwxmy4x5KDVm/clMo/0QtNdKZiA5bA
GGgyawf2s5Ly9J1jpwKY8ApCfI9waEsFioObpUNiSwZyJxc4A3rXgq93G2SMe6EQRxtzzTIqoUcd
McgKrGClEwNMnLNkkQxgAnsG5dzFa/usi7SkyEiJF+DSraXYZFK1wRSifZhArlvtjYkgBEnNRSvw
IBE/wtmWSWiGIh/HCgDu4/aNTdiaqp/u1lSXQ84jo9yJnnUZa+1fwjGe4LISmgMI/PVg03eCsIbi
nTOXL6I92nlGd+ZCFrXkan2oH177J+sWhr5dMSkB/Zy69zf/Swtufvvwecwxyh6XjIAoYSX5kdyl
oNeCVzeYhv761rVwtlj3d7B6zy6Om7yiurqDx0YXp8g6h1nilOqEtva9FRMFSs2QLrIXTQ/NAiGz
0u/PN1qNh5mW9tQ5oZKuOS0/53eUFXgpgGg7Vkxwa1DmXCigF3XKz9VJTi8sGfhCgQzut+kWlgKU
EBOek1/c5dQ0gx3MUMrYT5nm6/W2kQvQJeNc/bFSZS3OyiBbADkzTWKAIH12lhCAKmWu3mjSmKES
fcS7ywnvZUo0u2EJvWVVhKp07Io82NFjJYJwH/d9EUzqu1sbmSdgrkb6MW+5i8n+Mn+u0UMjURO6
Om+8mwWYVVgtwS4c+OUfmaOHHPH4SajtxgNrwrEv70OwJLQDY3GgvNC++IrDKDSmhgkmmzhlMXti
wtKLI8Kpo+5BTj6XuRVmNbMXstUwAwuW4Vh3tuhDmMF6lUJ2kTFtQ+Ni/H3WzWCJ1pY9nAWNW0dL
wfJf+g9BGvaqsNAanIY9QAkRroVEqKPxDlQQ+bqiMpdIRxZi/d7sy9GE0gqaUieK1VNRezobsq/a
/GsQFgfPlTTOrzkBMOEpg0vNCwaENFZc75EOdeff5yKS2LZMqZ6lQUBcYolqFguZJ6Y9VQ4ZY9C1
nNBTng8MCldLlVJC1i96LFWcSS0zCyfUGKdGNS2W6Y+9QRuk8lneHH9f4980xiXQzmdRxmcaqpY2
ngfTdfTeZ+SA4pTsYW91x14PRAr6Our+bwgWSfYZC1ytcrPeL1hzbKcj4Fu/NpjUReeQAYFAzC5e
+T/cuD3AH1k0xfJcB3DxFdLc9z8lkj9lniuy8/lQA1cEZvfcVSDca9cCBCH8bUeLXfEm3qRLuAoc
+lDvRbACgpawBOKoc2J30M12DZ9GgiUFiV3AqwwoedGLzhqpm0hKgaVtGKDGt2q++uBtdc9utbjs
u2UQdM3fcggQpDT/3q21nzPAMtj3KX1DPM3/qU7k6QK7sh9sA+A6rgdbmR0jhwe8v4pW3e5EcXVN
CUdjA8HExHA8R2wU6VaOVb0po9GusPxilr/ZiCDJ3FAcbyVPW+q8LF5ZGX7NVpOuc9O0wqFmFHyg
VGmQsvi5oasHYbTTpU58vCd9teg9bLLeMGBpubmfkexRCfiXJnylT4y7Oj7o5PHxoBW3CE78B0GC
rjq31M/gsFb3G+T/BZBjnxCxsc6P0SKGtdfMBOqDfjh6ABSUjmrHdyEf+XaQ7G0dBjmhiMUzBOBb
KJFNhD3rnloUqTNGaBwdtwHHRfA36gD/ERrgmiDzzFUItknmQm/WcjWLzAsFq7Ep0nWyfB+I4Iuw
LCR5dc/Ox+HnDw0SAyZQUqhfcpyiqtveqZWEOSpTq4/5IlaEJBQdVT16vWnpAjAmETHp12uz3WaG
PTV+IciFWnJlSfNZt4gd++ZjooUibSDPvU0Kg/wuDMniv4v0qC33L/KdNpGOdLYIffQdQWYK40ID
6tjmMD7CKkt1qzXIVMiDdbgRFBH9fX4wBNKpFpTaA9osXfvv4/uicvMMzPzE9la6gfXKFO7tCKVN
ukeCA1c6fKYISOHFmI6MNvydpFlnLnhtlIHnKXlozFpQ2dPZcPCGX8h3OF2Sa3V+D7FloTUG/SFa
kCD3Tf8dNsOeRlsuQcM5HjyiU6GVsUhTTLpZnurzQh/BJKANiP5aUWvI+tmrQLHF/fyHSj5e2IwN
OCvxa7ispp44iM46Suj1TcQsdiR3ErT0JEKo9QM7OOsQPqRKgyk5zn9Iu4e+a4PTcr8PBci5IaUG
z56EMyyZNRAoQKg8g2sfkYqbfjq8+BfoTNzdsv/oeTN3rwwKx2mAJL7JeExuoo689+q4mXHWF2X7
aEUSDyDJfrUcozHR7TG0iGiSi7tHXxlxPGFgE5gGzUUVSVXJxIVzwmwDxR5khE/i+fr5autoq7X2
MJZuSkjzt+pS0G3KsFA0aar8/tgUXTRCet2qp9RBYEQh7FgMvQ1t5vPHxF9tRvYw7cSF3Zm1nMYW
F5Hqx7kRU1AXRVPj7QWkJpk+GNNoL8jhY5WG67594ArFT/jUOrrHSI/DCXN7P/gxbrbUrz7P59Cw
UcWPs+j1Y0UtlSUlVbSJTWvILfg6bSyoTqqEA5dXz+bNFIeWqZiAOAH8+mBeyjehQYqGaO05zuPC
8+A1MXYQrf68AC8Ua/IY2Lj7SlgHSacUoGFSTJZvu0/LnNMFbl8IAy0vg6ZmvQawTSoZk1F5gPV0
cXA44cAtwhG4iVlXDh8czcscufuU4W8vIzstKjAuNixzXOn+Qw8DOSKtzkh1KSJ9Ze+JKzt31Wb6
jM7PsUe6yjbBC5TPDd6MEDykIsqzbLD6QumP/Db4cvAh63L/Xy1+0+lMZHVS6E/vTwfxY2D2lTfd
jddaGFZx4zzxhGRswdK0hID68DYj/LRraW/AeUrdNg0TvdUQz85sdiQh2L6PHCPqw73StFHIicrd
FQ3gLKjI5ze5iSnGZ5aZX1QNMP8PlH3drYKuxRb7c1Q2OY6XAZ0/mT7Y6BSA3E9TnzCSMT/hxOFZ
/csi5U/sqHGLcMTyayXCNsD/qx/wBF1qEobzrFrJ8VfKHWhuf4xipEdxNu4Of7N0HpRgeAq3OrE6
Q3BmMITKeWhjpH9Pcwnrc6ScVM2IozgasYF2vzFqy6RUzeML+KCx8YcVbhJcr6ccpsVFaWzgnQ3/
8nihcK+sQKLkSTJ7A5vXh/1OFqXBjKy+6ESymc8sKC2ZppICNoBGdK0VxxVq+DXq9BWcsR3hmAmZ
rVnnWGf9nc1wqJ7nA3hQ+allSAwsYxk2lhUjdWwBf3wkOsUDRd6Bs+o445lOIgtSokB0OKtwOBCh
1FpP3lS1pXz5Nu1BpmpPKhuKnpz1aNR2dyMo0+VTkr8rAg/O54iIFg1y6Qzd0RJH78BhQ/nX9e65
Uhe/FNxdB83EkqR32ItbG0LhOt+MJ7lOfMvd47cwHzaqBqKcT5oSfknUmpvzLbIRm0+vSYfzWyvq
cDb5Cbbrl/+xGoYgKE3Nw6VMLNppQbZCApJDnkMxkTN3s3yU8b+bmuLE+4WJRZG8qYjGpzsNV9ST
+WdMjnLG+jZLwhjgxE5X+ig/q4ElhEJNH9i4FbU9FoyDhcyk6+y/Xn5SryYj+9GYRcg62eN36QPE
aRuovFiNEKtnYqYgJNrmwDGcQAPUjFM3Zve9IH4ySd7qa/XKbj9MElTvxBluT2rx1kwQDIq/68CO
0smmU5hxoAayYxy4yI1064EpAsafGIwcOfbEUjnfAXhC4MbJP+z1CIAPRxuO6WlwB5U03Rkgha30
N1/j835jY09rayLXbgOYmXoGTFD9ccRqx9sGs/aaRDLQyLEM/XZdOHRIf045i9RtFaz1lbqG7JDy
v/QSLSFk9wdUl700+z0Qe1de7h6HmgwfuJL14ThFKapZ3cY/+CMCU8+4UZxVVnviRO9PgF6lIIdr
Awjlv8gyvmFIk9ZjGrw5xJCEc2GGC7l/QpDtCv6uPMhAwplwflb1ISMFF2rCsjBwvVfP4dXeHEgv
XWNGsaI/vmvFIJj2UIkHNSUHbq8C4UTqZ+u5Pz0yzL93CegUIn6UfD11/fTzDjPW1FkR7sU3OQKV
Ralt13wsN5Y9ugEzdwZTMP3sU8q06szN+ZtSFcmvwbCOpgamAxtpNSd91cRXWKVFj6pp5PY5YuJO
if9+Kd4pFNGab4CSV2WdgJrysDAdYml40sKU/dndBW34I2/5XLl5uxFTaYtQ8dYsYEDT7Vq9ZirQ
iZ51dzjuGBRyTfnkLAA+D+VuxojMDcuE02JRAkNIRRgjIJF71MDY9N2Bb7fiwHaakpuQ20OFER4Y
tJGpS8LNjDijLzCslzuIw+fJoazyRwlyAPOoCuy32olj4O0viZ6+Oa0dffa8TSqYsFRJK9HlaAqI
5MrSnAtaPq7sT2ROT3R6PL35CQJWqRgh29C7Jn4iE02mWO3R8nkxKc55L/qYF2vqyvgTk8CinZpa
E7VrcCn59Avxoq9KbJ7vqX7c+BdIx8sWOxmVkOkCKPsWgFQ/E9DrLsKDEKD5P3u3kpO/3Iq0/HSY
iKQ7WIMFLVsmYPAl+dlypSr7FTnDVRaF4GvrMyrH/hzheNcMceFhlthaNUwZgWpcvbOxrXHrNqtF
GW0JUNEbO2Qm5BiyCvfKaHfXEuj8JsgBcCsq9NUtSaVc24061iqIsE77kUoZD7KDlNHhEpje+pha
0PFqvAOq2AvQngY/I80QEHG7JUpVQ3Ovek1DQHkOawiL024N3OecqiBU1jjyrx5Yr731X/7H3ZpW
IZQ4rknanJf2U5SZp9zirTrrIJ7H+eRiEzJBBJNspvctf2F1r/luwdNqkCojxH4hn//1qQmF9jGV
qH4MAfRnaT0KQKS4+iSK23WJnzTHLxoxtHCE+JzOHJdkHwRgIz0nMPFGYSsnXSQCae8pcb/vBmYL
GQqBxs206B3osoPokqVeTshiBu+3jSISAht0fQgxjvvXxUqa4Rxxlk3qGZM4u/KxCxJUuOWYhQHK
LN/NBTf9xQcACkmYTC8Cf6P0NjP6Eh3GVzwrlLXu4CnxTTBZmXzYbT9SL7cul1V0Z/JCRzqTxGqK
XP8fKWqkJ4tR7CjCVN8DzAy7vu14aNeK/AsxmJSz+aleiQu+UBQxgviDZKZLQPrH7cjCRLPptQh9
ULCxPwKmx94XERNI2NL4z4mCWEEK62lhj/Q2J6bfW5spJUPAfIJBjoLBpwxZKN/0V4lEa/Bb3VCY
UEmiqp+MLfgCg2tL+w23oXg79t1nefkV7vPJuTS3vDyXFM70Dk3r4h0n13mvxhNzvaKTB8j2b5oC
dh3aTFJPhPXNvjXa54b+iGObjqha0sgKzV96KCnQXTT8xJrcgKzLWz/9ca5BomxINLvojHDbsjTD
K6oPEOSthRRupDpUcpMDUT8x3UomgZ8obb3w4Ob94v4R+Vfq3iLJLKdHUzU7nq0eDUMpruu8TkNF
QPTJlshHkyfz9ODUnI1J7/LBjblQNYOwr/DRGJ8x7aoZzG5sbyeq5Ow4g5s0uIn+gCKn4RDztnzM
zCIky79UoWZAEUk5bMavtckjMgErIfWvGe0fev84UgcHcvxSLxlMS2AYzYitHDeXV+gz903HPOYy
g2Ywsaxta9ztemAxG0OhEB/XlJx2mdR9FugZtrhOytQX2agAPhSmve+zza2uvLpeKiNaYAnQtPvY
YP4opvvImKh8/I7jjEFRRaGh1FINm8xWpZqnGcmkhOGh80YYKpBpI0JQ9IyYHXgS/RXN9XaAlibQ
En8qNty00rdY/x1YPlIJApr1VzlChapzJIch4a2aHa+9X6IlOHaLiqMFqgEwWgvyjydVku09RLXr
fqHYBa2mMgh2/yY+NFuGT42ZjutYqTSejb0dkp7HBasJakpE3UEQII8GJth3T2hP3NfSFhsVHgND
MTWpWRmcCrPTlCczF/DFi7e6FLX3k5/MzlTI0VQc1dK5ewS4jRXKu9dyfFJUAzNELM4UOkYOPqbs
opFHCi/+wDBEwsC7i1D99EFxUkZ3DxxD7BrxXD1zL9vk+NBPmJX1cd+/NJ/xBsNdo6jw3sKqlWr5
jN1uomtDCa61cEyHlEgaDB+tmWN7Mtm9rTvjwIYaCb+0aULclgoMMYHhV3th02gwJPfnJs5NkWUb
C1aN2JQvdxoMQFXNGhccn5rx2YGZIPwMNaDLQwoCPosUQDVDr+zgfgCzo1vmkOiWf3OJsGaYZvb4
OX4O09PTDP1kXQPacPq4K/h6NRsGn1oWJOu+gNRzzhPOpnrxp4ika2Fi1JV8NeoE1Z9tnDtjHofF
p1dHfeSBModsQfcl1YfXfYUMwbhZABY1hgDm98mx4MZ2JOg1T+iPqdeHEUuwU2htpAoL2rn01CU/
b4F1a3vHIZmqc8ILX2T+9xUJdDJXyL+MAq32PppvkDU4grBGAP3savYVaRerzz15cYpo2HlkuXVl
ynoMFj84KQWzzhphLsxsuBJB4CMWKsY6omnn49fR8yQVouAVPrkZti0Z7phjUK+D5hKaUfBsIKvO
r1oTXOSGzeGFcx+Sk2yV6mNgSszWpKXKVOtPRLKZze/bM6lwbgvHNoKb7ynD+LWOSD19HLp8gMPo
HwFgqEoQUE4ecV/yG3PrEa+1ngXZMUYi5VEPbSJFulhy2A8vPTaN50GRkCdV/c8Wc8UoEnbEgw2M
jwkg72Q2tTPJ7fIxqeDsHc8mnxHsde4ik8xkeFYKpG6/3M/pjZLQxWW5YEJqZHCJeVC0ituiphKd
M5KinK/Pzhwhjo8oI4npaX8Ms76PSGa+bUInbGojE/i6176HHe6jA5LjGwQ+TVr5IaoxfLaeVgDN
c5Nz36wNYNjsO+7JwLDQ/93vF8zvVhEXPmbbtmLdIvfpHCVRL/VmBmd8ESx1j7JCWWc+PPDT2fnT
kbceOdzxAq4/xQrNtDybgY8eO76hlnBKQaRAqkmHUfjeREXsWG+R5dpttxXG0/nn1bCQ9AEj2b47
bmxRms77GOmFckCeDaZXi9Oo5+JALcvpEJYgZF+gGJd3CvruLxa+zD52OBqOlBOM4ARGh9LUlsDO
KCG4WmDU1oEV7MTGcz0BchMAgJHT1fQTlq3ampprMFRe1dEDQEsgU0PLUoRZycY9asqgmvjTlAq8
Bjk7XKzpDN9M6PTyLxM4tHKHCGE3O0JoKu9EI6mLq4fKdqzZ5z6Dz2RCeXeX9bMhsJT9xIOH1O3x
tUQ30Y8R7Q5k6WjmNIDhjeKjhAcPIGcGtAntVOAmNItk44OtnRLRYStfYDgtsPB7govfPCbEB/+R
DCjgjw4uZrsAYKddZXSf805aHgESdaLkSRc6eupud3Ho8CbBDuZ1sLopSK26GerjE4bUo+N2K8Zm
/LRbGABsH78AXn7MqUu2op0EG8HXSkfgKUjzWJQiRVZ7q6K1Vpn/8TcIbRqR9JDfsFcZZNfBg1tJ
9yZgmfI3DUCCLWVatrEIkswOGQB2BOhvRT2naGVExakFUK7iVL/FSq3J3rzr3fWROAbbOKdWOqi6
nZZyLxjglvPmeZeYtOd1Hv48eSKfav9tbu9WhLw008neXe2kOxEMVTVLkno7J0sPvXsg3dsQ0Fsn
wRenMKVQIqOfNA1yL7pDnxCLiIiqFhxEazE0QIbSt4G2dq2YSN7DvEj42hLp2USclwW/rlJv+TA2
jPmNHsfIsUIYJN2ztjlQx4vzqD2VUtNBxSVayf5nuHVfRyqiO2GwRVHLoUkm9w/1SHuDK7tCHgbd
0eMhtw/jXTvg3YDbbtVTS9eSDxGjxSfpJ5QuWhadhPTJ1Hm5gpK+5iwQ7ydrFeVTCh5nVBAJhsNf
EaXBDCXzG68nULcZmM0GFUlXTaXt2Bljn+wCS80Yisrq4QtAwM4kv0JgG5kVhgWErn18YfL6nm9b
iq/Vbrn4+9seaX3jwZjqM/yyOq8DaaRxdtyCK02N1Aet5YLk0RJQBJl7MPFQcoh2fVFVXyREP5Tw
rqLOz/0nTfs4yETm7j1Jyulc67SvFjDlMsVQ9tp95Z/WtxnqhHobXGXaAJe/nGdpaEkRhtBv1OU1
Cir8IqL1MpMyIXUk/IeorcwTqRxxtSKRUoQbxADgS3MfZo1UW0tI8RQwTditnCPb8Hr9N7ivYLix
ISh/+DIvItWrC1EAZ8sj04OnnBPiteV2QR2TflGkLg8EadQWgoaeffABhzOkYFHn1UhygaQPjvTT
qzEx6eqlk+4NtMnnyVnURRY1QYZ9VEw4El6m5lwYnuKo1PcEs9dP3WOj0n07+kB2e13rVEgF21b6
rv0wSoLZW2LInHqpFl+ms0LhgXV+AxSntE52arrG+h7B1A3sXu+1Bbse8+6BauVvacB5oKxgIzM+
FmM03X0arCU50XgmJd9Ay1beWZh5j5/th8ALqRejQD4VEpQrLELxhJlyqrRZVkeZGu5TZa00gXlB
jkyKCQIyDud+6lWka36GevgbfmrlJ7z6+SotMEZbO7vSti1vYpTOQ4JDCS9cXMmkOUtaTy7lzK/Q
nghoAJ/rEkq5fI2bEViN97Aj+dtuPSXwfP8uAFK8UqzWfElph20Kri9wzT0+02/62t5IwoRPCwPn
cN5e8xtw3XQhoYLDNC/HUlZ/NcsIDWcaGtMY9Z7ZZ4xJhWluXold6syfHWIE4H/mn/8Kv1aqVs2L
emYh0LovqrcuBR2Sly+UTNuSmtcQKB8fX8gnIbcLHvdD8XMUoCiF4zPiiqMECvWTDtGfP/NFVIen
lUK32pz8VI0RLMB3Zt/IJDb9PlaSKSrIhtgaFpLVC+8UwEuJ+Nc+bg/n6vRB5cDRyUJ2aEVz3poz
qwQimQDmqdNg6fQ+nlZaY+EVsekauL6EAT9Xo0mNIK9AZY7aeBIUQsj5llTr8zh0DS825a2VlsYu
AvO77PkLpxaGiO4NlsRMLQIRQIkgIs2OKwAQSF/QOnyWITgAG3Ob8f+2hJzjM6u1IM6WyKE4aGID
bRbpvY53PLeENNNaVpx4jsTIrB4l5no8H+qQeMXj/hAmXw3bsunjqJHx1BI34/6bi0914BZe8a1k
Kee4S44ZOzF7HVUnIMYpzmdAhDyQt9RdxLFWXq0M+SF8G8oePSzODwLt5abGOjtBLocpYZ4IX0Ql
w4RiIpSw/cfCF7+7gc2h3eyQqfRgKacx8lZu5eceQBgpgtlDMWBghNeQe5naI+BwrVhCxtI4YQ6N
SgqCOz+VgV6oCSv9j2tlXRoDLwbrwrQyxFZpoFWK/ucblDA9KWuQpP0+KY/tDLxoHDc2sNFbJA2k
raqIUmTwtDXal56CNrcSQ8ToKKonB3PESayIm8ONv2nG393OfIak6xMzmGzn2l2swseiD2idKcRR
lfsi3rAYoj4p/DL8/mZ6JsLMF7JEBm/0gcy6qI9h+1PWWlAPjhwwEfz453szBdcigNyO/kjKO9td
KNTd/vOieSxLsEVIDjwak7fYxoK2zrHAXXe8f2WyU0FajRvpKV5PFAJynTWGImWHGlivDsmc2tli
6JfAupIAMKpfNE+YhT+3aS+MZL94YjCKggCZYOoEUCoVS8BFpzRsiJ1JblX74HLusHnqqvpsal6b
sUB3JAk9HphWRgJ6t/fjmKcbfIcr4/EHtB675zgzDxiPSXOmRIr2R6syHmzQw4/tHpmZwze6Berx
kvxV+65kvR99jmfh+iKxRV/Br6HZIm2fnXxed4ZWn/uDQG4UhSVWXTC2iwkSilkE6lq+LMJXc4Z+
WAuLTg5ru8kevIClPsvKKtdzgnafncE8smZ6DB88CmGpxaGxTb26ZqQLgdXbTVl1fuzLsNXqUSF+
61kKhLscgUOwHJOg9qBc/nA/nQInxghY3R1SY4Xe5v8sCa0n1459ynSv+KPFnrBlofS1tWxxkjL2
xGuezQHF0ECihOPIwQorkFfT/KonMSWQuvIc3zKI9ZFlJfoSBM8KwZU73R24j19YYNvYrUbxfa04
LOaQV/MWxwxWQzUm3E89GsPwAoyst28aOA1NZUtDJSFWaxJsGdN+XqLQ30XgqJ8CDS4EYtbmFvRH
3i3hcEd+UrbMocPmiADU1QWiNL4CjflTjlPjYSh0hObNOcN942feIyuDMLEOyzGSccsbcu62uNY3
/p4kt3ly66DmXzkBHL+jOgH89zG1ATH4jsml7Ok48Rj6n8BSBOIhQkkfEh9Y8HuLQ6U9FMO1oKJr
0vkmyuICHJ/vyzQWgicg3LA2Fu1Szlguk0idQXKgLP0kVIteWqx/FaEjLySoAhx1cyw6Yuur2snI
tPW5sCZ+d+YBscqmOtH0OZL8ISci3VRm8jjtCPZ5jh8lfQMigo01jAV6u5VdIkevuoroiQEQ1kSv
9JvVZgCuuUGszIT0Z0nyxzkuui9SK3dvaOtp3kJT3fo9f7QUzogxlf+txMRif2YABAO6pvIxm5M0
BR8X0tPpSYfCMa1QQomDVQIDOWG1jO7GwE7V0Y1S6QEv/0aW/8uHEiT3Qqad7jrpqXOb+Gi/L286
5uwtK/pBFxx6rB5ULaxg1Ecij6f1q0gH51lYELDPWL2Vte3m+jUHDkJnVD4X0V2T6diw36ZRDZo5
YdxIGJbtU5W/GD4UWud7wel1ZvLhOhmkMLeZDTG4/WUyKZ7/Racm83iXs1xnpMq8uvN1njdGVkJ7
ae4tWb/qVM7qXKhuK7L4Ye2D2YkzjiEjXWqBlfOmdE/RxNoonGxUBthWh1iLiDiMGC6U9ZUYI9Ew
ENxNiSGWwcpUMESg70A80xn5qMb/TAxcuT1Qj8nzss1MWGJ/GQTxSCIxDGpNkUF77mbRdp8Qqrok
t31FUBKsIL5HKD8C71pg3xrYhOnOaRwd6zLBE/XVo3VUT/LCAP6//owZetThMYUm60RuwXGNa3mk
yF5T7P8SvzlYn7HIulidvrJp++BWbL+eEsrKh7vhbBTQWr3oT/mNvA5LxVYQom90ZjGQleYj+YnQ
ZOmlT0JG2zQ84iwMarHiUCjFBcepAWGI3vYtqnNOqbv+X23iLdpo0fEH6J1QNqbhgqg8NEpVTJkb
Ezr0QDPoRkUDm8nFtZK7OxngQ2ha1ujc31P8jWanh8cxY2gelNI/AbnKlsZCgvZG4FpSq/j8cbGK
n8Z3Ca9NAtfwoK35NCHOoEbntYUzflVNDiZorhuzcSITqhC3VzeBh/bxKY//rNd9FGGXrsmrmOFN
hI2YcyorygUbQPodDb7z/zi+92nj3MROP0PDRN4SlSjAgFnsUJ8OCFWjc+C0hu48s2vkRHit19gd
YjSHe3rvJATa7H4fnmAz5wsKfrkhRv1FssgwIAe4u71HwDRCRwq6MAf+xPBfEEkg6nZkHbF3N0cx
tsTJpGoFlrHQc+xC1FjK4NWnXoNuMFJ8DDJhSaPfMGn+p17S0kRTiOKepiCXTjtH9YTlAKYVFWtY
8yenMBxLgfXuxCfF2q1ZXIzcnWwYW7t/UAYB4SE4tl40c4ISjskixLM+X7J9Nolk8O1Oed6zT89y
LY7vbFoN/1/Qq3Xn2g1XO2HKNJIwceYAPZbhBVLSWwiiIUDvEB7IU307EwC7mhyQKOQu0bACdxBe
wiTDBL4z31NLEv4/aCXNe26r8frqfwuL3orqKYsvWTRXXR+oiIgqQp0Q4UjaA/mGdzpCZGXuejKK
3RxVNFA8zlhwZEnFwWZwjl4RUySg8AwPE8IZbug1Ctq38mOz+t7CrxdLNNUAEJ0yEwn0qLNXuUsD
fAmM0shMMdEdoeC01cbtn7RLKdvP/RC04T2M4ooVlhb8FgyH4ERH43AEtHNsAMwQL8lTkq4GpvKY
8Kps8maKWu/NY3MTFolEzOHvwesNcbhTZXpJCqDIDCSy9VWDvMc2pssXuT3JVJr21H/HiLrOYxmV
y6aDnR2eyDR3NvcB2bwX4Ebm+q1iivSCJ5QLIugFXnV2aqPgUYL7BZEfwkKstXDZUFW4LXcWFO0p
W1QcN6uufPQQ36HN4gD+HcPamziBxMQ+eVIWk92F8DMrtwLz1z3f7IWwb1fN5c/qeeuDKCWRoey0
0hrGEbxvghALtlXs9Klho0RkoR95nEJkXGha+OnVFRkLuPSxBhcWgLyZUhftQmCtwN5etKweTeDe
wRy0T5C9YsrlGqQud/QRpdVKmjNWN4ViLWVaibwrzr+ALmr3bdEKVr7lGOHhi+YlMPb1ECxNUFJT
BgLCEA6bO5Ynd/Bx55Z0AzERjCKUZ/cw7lQUHVGnnvh6ODJ3sFAEgXQf9fnVeuWYnAn8vsAK3nDw
LwDs5oMknuY04RsI8FRSXtyQtncLmdH4I+Sj+BfgjyXO2r0jMCgEjHDuOb/oKVRAoAvRb9QHVFyZ
/lLAc7fZ9F77NSEYOG9SpXwpVl051BAfT56x/+FQtV4iMrGH/ubfIhoHkvZEWkMkQsck+aGznqhT
hJPzbtlMXetj7C+pwj2hY1J7DoDwu2LHy58XU7tQN7F+2Qtk3N4anEFNyv9ZHfKCM0/ZuzGJe7vC
WbJFLWt0+ABNWiyzxAV9YR+Zl7oiZycLY7Lf97zR3CTcuM4BFUUc99OgnuPsNQ0iYS28iOV6952D
DMF0tKQWZdXXOwKQp/iYC+XLBguiv/PD5s7x18dMuALFE+V5rrXZ5Flvuhtk0ib5Gh0W1VdOezw5
RgY3a+2vxTL4nfyI45PjGjOhKVn1IA6yowTLBugKtLL66toFKUQIgPjuodL1Y+jIpo7g03BxYtFO
zqqIu5WcfRYuGoa/EJUs+p1ngDd87buOcOUX5hy9XTD8pANgYRe8nJliMFpLxVPB/lddrw/4nwG4
hp1U5+n3eM/5Te4O2OqTYmbjhqRy3+iM7hof7NukS6+iQNN6Qf+LW3diFkj4x4vV1QNwAjJqw0wd
wKU4M0tHEmaJGG7ORgya9pCyhbeNRVw/5WWTNXXggBDTCC2jwf8uXRTQYZ7MKM8P5NxgXcs0/XS7
Jy2eUGNbljf02aF00DokkttrRRhHphUyFLxngbT8LYemcfakP2l5uN/N/oTQXDPbGj0JqfUf94QT
ajo076MK/eP13vVPjUsDwIBqdtMTRyc3v3vhgh4OBzV/3URROeFHngm9/cGy0YRGXoqVK3LG6X+q
4J7DtLmhMdVr7ZBmavWX9fF0hFms9kOqzfKOqjA+HoVyUfKYDVtWV1GYzqSFxPJkLYnXKo7gehpq
dUzQdLsn+Ul9mBJFl8B+q8jXQx3QnKF7Erb6+JvTyrIH1hwWRFdi3ntelT+4vjilwKn1aqZesfit
tmElGIi6fe2hgia5o079CaqntoaTm2d2pOnELQXNQc5Kq73YVIbZWutCYeuxxb/TgXqekFJ4Wr8F
sKY+Vb7o6+YHz+YsXREZ0dXGv2B0t+fAuqeAcrVZp8KKk5U8G6XNB3Whj9x/U3ooS2m6CQTjKd6j
1ScGtfS0CIuZEry4dVY90FyPsL2m/vW+/XoalGnEDRAqXlZAqLly/+Ln8kOMolvdc3COwvtaKTvU
5snybbeQXStFF954m4H//NisDo/Uo3+Kj+Ov5/evmkT0AvvmCa0JUai1wK21EjQktetlIdN76Cno
XevKrVwNo4eHCU65BQd/kClPqVzeXfdGmAqWdJwH4l4vNCVEEQjy2SoNgAaoEd7EWu5q450hM11A
yfEAgP2iJM631B9ecRn7LnIj6vG529g/Btctz2W4dyMtFlWrGeDFXT1f9dZD+l75EZUPkMpz6Xra
CQ+i0UQlhgpXXMl4PLxy1wjf3TqB36uNEcplmaVY7MqjPWQ6zjPu205qFIzH7dio2kPrNAKq8yrw
9+EKZfE6eMnAcIGQEjwU4hYewRJsRgVPTdmAQ+zuq+itLhltKuV2D1wEbWCcgBj+tUBIlOU6YmWs
suqdF6vPyN3Q1RDsZaOZIOSbEaztaaSfCkezLce+zuWHY44Syxjr/ZyTAmoa44VtrknqMQLee/IF
bel/wnASzfO9H5tyTKUSjL0r236n2VFn7ZI5iNuJZrTjs+U1yUnRXcqvorbRDYYz14WUuvhJL/2B
mjHBfVE0DHqzIowHlWZZgd1Ct4E71vTv744JtYAREnmEtA0taQpkmn97lGCnkxT8c+XBSegBVxZR
dUHZm9LVtjeTaAyvqVEjSTZVHKORtScMxOBM7ttxTfTnwINNVSFICPOsMlDgqJGTgeePksSDHMc0
jyvzzjEFgBLF/ZcGM2iBlBhNJOchgajf440cjitIKE7aTgv6ZZv9EUw8q3rXPogo/hsDytLYBjrC
Jm+bWVdcRKRytRMOYlwMk77j4xPeUFFy1dJBxhmwpsEE6Flx9GdzwTJz9dclT9Pt4jAMhw4grZuc
09vB5ZZC+1AvDMhY2DdRE0JOd/mOlP/VhYAYcgc9ikQq9Faygcxhypay4BeuVo62ewSWCeBhXeTJ
hkt5Rwm2Sk7M3K8BR9AIc7qpYG2s743XL0M8WU6lCTLJ7KE6IkbaUdrS5AoPpUCRs69bGm7X3kVh
Yp7WtLJLh2SryaJ35axez6D9xQ/mP50L64oAtzOsC4zMSHRbuPrnbUc4sHJTR3Msy8SDi/rwp/Jp
+JBwhd7JprgicHQXxmHnutbSc9CHOiDqSrERYy5HmFY7/xl0m31pul6QVpxLrcgeuvL0ZJJPQj0T
TRXlgz7SlR5Fy19bsJUCP0JP5/9KE7Wi7qeGYmMgf+RKeW58hsWSgMJLSOR0cKVnMmx9HjO3vsC3
NqKR/dV09Zy2PnF+5rHG/ln2Gsol1HYCdeLfeZYl1j6GS8ZVOOM8oS8gMfiGp2mIpEBJH5GLz03R
u0iiIi4dp25Mduuj4YboxAzAJmQU3fnKm/dpXLTFOr0STzbuRiN43WAAHtvHlolM3c249HU+mKJn
sN+jAFen19sXYbIW01oKz2XjGzbvOalznwWwmgqrujg5gRRV0OvoF+f93iwxlIjbLHm4eeOo8H4w
My6MAe8NvySMbBWWSjfJacq+uwggG16a1GWTm+XzK4I+enAmrwcB0N4G6uFwR5h6vELOaIkuUIgj
6Dk/PYGxhJAqf20SAwmPunVAASHkPzXjUffgT5iUDEZjJX06nmBaIYD5AcgPzF+acxYeLcWZxlDp
yuE3LsW2EG7sFIxgqCWa9kiJEvN0FiP6I80+8ysY9OFpZ0iX+GWR9XEQORDXuVkySPefvC30HKDU
PyyCFcXQNL43JdxoOtFhGgpJfYhnVz4Wed5+5xI36XxfDuYg8FpNs3D2O5y+jmdK3xhdZrpz0NSc
/SYh86Qdw39bc7ozgfpU0PCKcWbQt/RhLU3otGF96cPXp4HqwF0MPnj6kgbCPtV8AE90DgpC26eY
Xy4shZB5UDMalYhLKaSUoGDjAXu6gHFNE4tMfEcGi0OBMDOeO3ZTHFGCwOm7A5VNTLHdnq5tQ11t
JECx3Mycek8EFoL5uogaEmGlHLmhdKDI2MyfOt9SdpTJyHARQhyq9NlIzbdgGYO8qVEEeCwg8PKZ
dqEYcwaZevtf9YXm03PFrEF4zIxQMkEfBre5Cz9/n3nm7ZhqtK9z247H8PzPku9GizFO5XuqiwBk
8p0k02ezBARJx7tTYqC+uMtz8xjocLXseF6MGSvO+WWcoLjGyY90yQF3iSRxCpslLLte9eR7qQxR
GXn/dQpgJJwgeTLJQn3KtuiVZOynNju1Juvj5qjEa1aroZPNfqW7VdQZsVc4iDi41hz29QPDhDdz
K7LiEhBTKk8Sbb+Z5G7hsSe34W5+V/hDIrGdubs/lsO/08xCZmGAhEjsET943Ime5j2zAOwLYBIQ
l4GNaF1pGq1Dwhi93tHono69j9LYLyMhun1WFV9Key4yxaoStbRvKdjQkaIQHk1S5bu5ZNT6D8dk
VWEIoWPhwAlZWk/1Bs0PlE9gdz3bmJ9/l03OpmoZAbt0DyTsI4ByuLUNF+NR146bHHePSpKL/p5Y
DPKzMhRqWnFeyOAdFQhhzSrnxdlmFdsBYm9g5PBd4sX9/MrrfM5oNedsQFhnq36KzpIlpN5uz4qz
Qto3CWYcYjdSR1id9lfAKdtrg/XNdUffSLVxOw2noL5ziWw5ojyJCh6SyGeri2elluoT4z0kaf2a
tXExFAflKk9SAG5THJppcZsmO6XLt1diFp5qJKhzTi6byxaX45/Lpmdh3yB1r8aTWoU4zUDr0U0E
vBxBfZMxQxRfdALF5kJVq3i9kJXwwtVjwQckn6FLWxOyfAScqPtediW5hXHZurQvUorcqlb5+1Dy
BI+tfwtsFlRvIAyiZuOwgWY0OtOeYkMFZjorJpkKLJ/Tq1KvFKcOV1IFmPRJ6tESY7bvId1mO9p0
JUFYefjTqRVdQWvAdAhS7useGvjiYA+1gXHgCnhNAtEJJ31kh4FTJlVNkdx17HdDbfgf3UkKc3XV
Pzw0VHXe0kH7RlgQ69AV+W4vX0AysH8jksrA1s6oW1NV5iToBPpfULUdlD363my2fEz57nUY7VXG
nSBfqpkakg6qzkT8fyTVZDoyvEY/9ZDWCHVdMT844YL/u8D6BaWQAL7KvtnkLMR6ZwDuXXJeZ5MY
gRdR2ITkJbzXFesuyadsKYp2rvD+FRbBPyyQUlIhTF9CNWlUUxI3B6iXwU0dlQC0LNdxEfADpm4h
QZpoimYvSqQU2gXQEVXetqXAfu78LPmnvAyocvgPoQDX+FXfoU7t5q4kIcSgfpIHLIBlu0WRT/0u
yzmdma5R1vKQzueFfe7GRJNZjPTCJhu3Ou2C8BrhQ8WBzvPqj7lZwugKrBUJOPdWaDgO+o0a4fly
1l7UoFHAdiFV/Y250H6CNEZQcYeye7vFil479F74euax/DCJ+19HmvTQdNAFhyj6z3iWQs31Pdvw
uX0HuSDvMoQ4Sh5F1Hp65YRIuqnu0qihuL9KGQjRaVPFMWaMIH5kiepJvHLZm8AdmvvzPsNaRov1
gm1bQRX9Nba2sexoiaQGlnwaFCGCzVzHPs6aK7suqaRYpzg0MxqWIF7errlRq1yNJhEf9bngTQi6
AqXcRxic8Rxglnyhgp3XVGHOT/DLEw1f6RyYvHxRyfMLkLvm4alEaB3Zl4ZCmJ7HpK0llXB/7ItG
lvoLVex3GFRP2MWuZtkHaONK/Xj6fS+pLLy25eKrFh8aNHQtJP21K2ojUFjzm952zY7vTW9eDFax
pdbakjzWneGJcvTGBf1o6yeKVYAbR9/ZlLi3MTzryb69wtglSdJqeto3X4VvrgevdjJnpPf52eWa
IlTK8a81oQNDNfddmhU6Mxh3dcumn5y7s8Z2uY1zNaWOA6iM/tmZ3SDvqz3LHKs6u/tXVWkq1D0a
dKlxvdwgA5+m9QiAW8hPT/Duql3Z9PbhmCeKwMlPIj4O2jDQreWgH+WyMUtKH9X1jnkJYhD3CMNw
5RGywN6fgpciwN3sV1clpIESU57+9XDbdW3AlakGp+lpLB+XUGN3/IvzhYHtMcafXK3+cPSSwg2D
2JQymrRJe10qZmc3ixAbWPqG1p6sYOzbyU4OGHDyeLcfdSfkWe9rzaLXHlRRhGRL8YN5nRqfaLWG
q+EVZdJZ8bGu/dU0OP/92E1DLFMmwhP+HTDdHW3p8fR3PebaDqVkOCggD+eVERVYpU8g9BIPDC1P
XAtGB5q/IwrGk5ynfGTcKRS/HTMq5vP2wryqp03ryT4H+XgY+EXxSrElNHyKOOS8UYMMVOyXpFK5
E81+CtVtW2nAwdSy5bInNT84irLaag9eXNVFQzGYfOM4OqaooUKtEd16g7Lf6jyb5qXo34e/fDEY
R3O0MN/PpXsYajRHDM9YaTpgCTPLxsIzhmlIGq1Y55tgQxjdqluDSr0cUjqNDrPh4tlRsWp9PO4Q
vs2W3GnEHChc5/yvDcINoMVCYwd0xgoHBh7xS0f1UBaJHnezbfUbS9eUN4rKgpEv1gdMFz9egzdl
PytFazW0Wefa0vQTwRELmROmQBLbsnl7mtDPwXd////PPJGBsjp5IKG2/x30HpOFK6e9JlBuMqpG
53c8/37HIilF7AAD782ac/i95owubQSSnJjuHlsu/jDKVa1j2MpvdYerFMq9qfPJbhLvVNQc0koR
MV7eXkV6KcU9dVZGjcAgmuR5B8TZKwE9FcCgAlgqiMzyCmSctgAPOdMLlPUmYutJ0491tvJNL/5V
IEFs/u59mt0nWIWvkni7frOZrotZMjmbvBBOfZydigmz1Qg60lU1mTxJp2xZZ+W9DFxdS29ul3hC
8heinr548UhC8HDjCuY8ziVObxS5XgAEHR4//OKNu2MVFWBksjxMmFobXz37THHw4IdhnD5n3S08
YgWMS8Vuf8XNRKEiWOuf9JL9En7MNMFH1S5q0ZJBpp6xhykuDpvvaktNkyva05Uur5tA9muMA97n
XIlJ/seaMn7ZXuEmOfYraiHH5njUriEDujmu5xwI6YLGEuP0CUbKgfQ9gwac5GPncOyvVVY2S7mr
zSjCKLoAVRHD4T0njnTGdmZJkH0949aGpgUevQDq2Ta7uFM8CC0Vsr+Yj2USwXRvWAUZF6qNRpTz
JhPWTgXRSmANjzYdfjMIMsmZtI9pnisstK4oGBGWB7gtOPzf/oqI93lZD6zPHcQYmB0CX28AvLTu
Q0aIPpeTC+AfhsbySKxpcIGegAqrDSnNYi4PhMts2la93w1vmkl7GbQ60y3S3XG7Tp5NgM7LSwpa
sP+ihL7J8dqBcdHMTF0+PEETOLwIZwUdy1t/0RyqDLznJlKrKvJDDgx6r2qtov6p/3voXdzEQI1n
JtDFi5xiFzvj319rPlNZkoS8aNYM/v/ewD3qsaoG8Df7hyYGkX7Ndc1W3i6QZ803rMlVQESexxKl
ayFd74PmImoctDYNL4hkdmFblqd6AyFnd9A2/1vphUrm6DOOBfjX6Eq6K4m5YGMKEWC8AamuQ0te
7PkqPODProRs+Ma3yeQu/16ju84DOzit3pq2wFPCWpW7qLyaCHW1vhqdmfcx3rnTThh4xEmK4Ipy
6d0ju89+aAPnEj+DNs/b62aAp868h6wgNQcPp9c+mSMoemhHj/4yxhQii5S3onqzIzlzE4beB31n
SEN847Kg/GgN+n3GQszuSf/earC6fnMR7ASnjDvkjIKZx1VqpzOpmaDDRB7Jgq3u7cIyOq+l1iKa
s+4yo7EAZldUoXH1uTBag17Gu3FmGQuCfvpLmXrwQfXO9XRK6nTZ46nBwM0TdAMLkWUEkC5DQmke
Md+O2h+/bu9nBMMbUSMNKDH3KV0gLcLSswj4ZlM6FZUgfN+/aFjuKES2YsK2ztosceNxKCN8SbHz
8Sfj3E8jfh87rWoyF6oHWt7BPqBAIGwhrcoTBfVM6l1cRxkiYyI2u7pkzZ/Je3t/DIBtQ1xr+P11
TFSxb3I3l9Adtqq3dKwREn2Lp8AH9MEKKuwOnhK0Oi3UUEjF6trv6XODaWit2/7EvYGwQ4JYJ3zI
xZ5Hw5ssGXpCjTx+ClBrwPdltixdDAYfsyyxMY6EbmFwIsO913/LUilBrzSc/U9D07IkNzFxJw7k
4zl3s/oZuoKTheeiFqCV2XfaHgGAGcK/4rG5g0ZhgP+07VDrSZBRunwaAhHRlHwWNIpxlLzWEGlp
xisxHg8H6StqoZ9EwbLqYpZE2tXC5JmCWPvWcv4scy/HNyfS+2np1G5WPUAJFzaPHBXGpDv+/hN6
2oIPXBcRcI2RmevOwfH8TTpNUNpFxzBUj+g0V5q60FlENe1c/PEoKhOrbemp5NChJ3WpFc7yp0XF
LeA4xgSP8p6WQBqvgFRs97JvpCkO3Ai2OaIphXnHKtAH2bL5J6qKPIckiwfWWwdND20uBWtM8pF/
GTCwuL8JJiLDQW325JDMb8LnxsINXbQNQPw9V7CtYoJrIlXVf+Hc9NlMj5/e7gFGxp861lPVKDxS
eJdxEzcNO9CsVi/NaACjCQZhxM8aUGbPnMikw3zNP+W06V4qqkAaaTgpN0hr9eV2vubIL6mXEobj
A1vkzofyDwo6rR9yaExUNzbgJJK0guTDWRY+oCEXFd6+aNIbvDtaniOdalof0Q8CsZAI72Awo+PG
m6K+eR5vwloa+bPOXjY/8G7ynXJnKx5sFo670DlUEpRTHnnsgW3II/G9j9SJGbuKEO5up1mpr0aB
5mwsRLo0sBgWZi5U2ze4Yito6Rezd05XVAar+DB8gl9HEtq9jkJbKQlDMSTWgzi0PIgSYj9qzCWb
6w4/yi1+7CVmCUUxZwTpoFgPvPeynBgtiH7LksD7eS/Givt312BuJ1fKuZhEtSlQrbYffKaelDXy
t8X8BkPkWKjHH93qvkIwRSoWf1Ge1XQMFKDfChUS+Vzex62EXSxFCAzzf1K2YUICHxtpt8tbny8w
orksDE6b4zCr2cMe6RvRyLkTgRvs/P3DSALv4bbOCicK8cYQ/j2/rXYQrnpdflzcZPCH9Jc50b0K
V6BQlPg6r8j5JdtkThdvF47AMEDsdy5ur3q7RSg2u6OL/sH8yHHr3d926vRiTHYH8AoddHzTcI/9
gyQmju0nenSU56ExClyjFlavY9wYLFN7TKcv1ozTWm182Utewv3daFtthUmoE8YxDBy6lyhyUeWJ
pGZ83sXjttEHkYJNraoxTp8MV8AKCu7Vem0vYsK0/WarPzZb4vzjGcR4evVe1+RSZsFf/P8Q+2vy
1u9MPxb6FJRQzndXLygcnFCODlsaNiNarzo8T3CZFx6gEAqU+8mwdrwJ8Iu62vWiLeqB2+EUrtIb
6EDI4dZqqgw5YwgXZN22cIRsG10MxzpGAa4NfQg9Md1lqHrFfi9cxbC0YelzqGoFgN8CTobYiXyv
2qVoc+Q9IhGKSSlSgLgecl7Iawx3TkHir2r/n/zFoYgOCAss1YkH5lpVSz6zB87PFv4sh+DQ7hj3
z1cDUau1salYVef3XewYKWDQ4ms+C5zJZOuEQhtVAf9HzIrunf8s6IR8ZdBcJnAOKb1NJNgvX/j9
G102dfx6pjvJhSCNGaf4S41UKzjD5CFpr3zFhrz3jDmCU7rwg6X34lUKCUHGowHQBk//ck/5hF9Q
z4Rr5ct4LiTF8ULr+u5dyv2nT8Tryscsa2iB6JCmO+NW6vVqihWqme2chRwOu2ce33X/ZOUrb9v/
rio+EuqN0qKLC5zFL8NgZRa2/1a0uwDPYnF3fflSCcXhBn8sgZuZIPRxkaZRo6qJ/FLJnYwcyEew
gQUlWR5i5G0K09XKIn99ZpJ0SzL+8HcT98zEhS++VanGPUcJDBxJtRDnXY/aXZ9oz2iCC1/RtrnP
dbT8mKL9rxkFZjkFMjWqysVo2bkn/3ARpOHXm+JyGYJr6fAoXCG63Vl9K4VXE51JN3GN27gLjlsM
oBjEO701hV/1ejycqFxA8f0FVwE0A8vvZSxeDytgmhUo1/fOvmhPesJZIKjtWjJZpgFAm3fatybP
OOS0wODa4XNrOEzWUjn79BZU1RMTW2JyaLNdzSOrrNKnomZzdZZE8cjDshhQAUZAoIbRGXIpG6XC
jGLM7J8QO6rmORCwZqIAthSzEzfKJIDOtB/7jeA8w4Bc/KjNW/abOMHZ3/rE7FyZOq41Xr4tH5ag
Hr45b+1mZLGuRNXzmTlIkiMtLhQvOdbgip9gs53tskDTNe4Nu1AcwFE0HqVABxsx8ycqyhwWkh5H
xIG+4D2xa/j+akxgM9qbCh84P6tOONCl8vI2LuVPZ+v6L24QVqs2J+YLREucXWPmYZ+wy495Kcei
YuE+YulVT/12/38m5vcmyNaAC8Aw29M28FXewEGqCJ+eNvJWI86qE1gsaik3GKuh2tVL968MDE70
dPWObLKc5IDSDCQ5k8EEdmUPeY8wiIRt+wKZGc54ZeVyPjChsDAPcYT/00CY/ptT7BLob6Ya7Bcg
2xuyVc2xJdAzKtzLK3hTNWDHqaP+iCSsRqZIkPN+dYJ0LL9VgAKd+Sl9P6VJA2eVSP+QlFYK61jR
QpQxNUsds2P2xcD75dXuRePMmA2Pf8fC5DtnqrtiRZyB7OIHT20iiq8f7S/+JfIJpUKKg3nkx34t
ZccS0wziCUOq8ACLui9EakpEbearTj5eEdpMlszwiqTbNFvJ2wI93Lv4Za2bYEcR2ojrgw2UcHI9
AYv6S540nEAdsFwHCAIwLguzryQFLjXg4qw0sFj9nj5PGnxaV/wYZ0ITlo01b/M8rDzhu10l4Ewv
O7LWZqkld/w8JH0HAtXvx7IVgURXAE6faEuNi+Hbrlof7Nnzt1F/K/FJQY3dllxQn7PwiGOLHWBl
fOK9FowPe4fpvEPJb1aKffupSXkR8hZvsHWba/IjT7r9cH/gitBhStrL8w8PA9EQvz/QaRpPbQN/
zuktrHfGCU4tUirmMuJM8/XLx/OP0BzfzQ45qXfyJxk7jUD1j9pjB7PK+Q6Jx5QppFDgwPYJLzQf
F3meeZRcmdKZZG6409ojUovABvQNhzdDsdBdRBwJy+BtyQIEQDlXEKmKm6uLGwb4evijyBEArnY9
DDbq4JtLRqTmY4K+FWcFGFJprvoFsP0GI4gA8rYNERq2TdYAviW1+TPdroHjgS5u8bZBTNGqhwfO
pOWTqxfmRlDy1O8I5FLN+WsbPcMDiS8epxCQE7lq+yWCQbz8F6GpTaJVJbthb88YNn5DNkXIE+Wg
hKxUQUy6CA4/vH21LZc3uF7PS6CDzdFzu9qe1nA5csCrEWtKndU8JzoicSKBjLH+aFDa7cy7Z4Yd
rDGX7FQONPbL42M2KRezsNLp2FbCvp3OdAhf/drLDw7LPrE+WrqhnXLLhUsfVCijiqewxZKKT32Y
To5IsA+HfYbIZZXabCnCVGbvFkK1v6UHOxO1SMvuNH4Gf5dYlB5IUQ6ZYOG94aYPqGkUDry0779V
ql+RoTp/4QDOZPi9gJd9+4+kxpiQY73VEB+fgVwyABcrW8P4KVS9s3TRgSSuDjIJLwGp7Yvqw6T0
9nBA02/jVXtpzMkFzz69b+qDPhRJcERy8ZNjqOTann7nA/JFmJLn6kPzZs8M3YzuxXwJ62wcesdM
x6c0JmcNiNrH7X4/pAaJgG9LneX7isKeGxLgdtcY5xEyEgPWPDiVYqYvcVv6Jg+0zwOAXDt5Yg1G
Vj5BLkJTGBxteOZbPiPzKZR3JuY0+ogm16a3WM/4W5DojzgRfK9+YzzcxbYkaPeFXskxvWaiYSeG
NL3JuSeIUvXDKGKsPqp+WVZc/zWkibCMJGX9GJEfT67yXvQtu8aryHyf5hfOkxJHJEDfc6+ML35e
WnJLHcLtiB6s5ldS8CHAgDAZbLQ4o6BrMkaFQChHt7lq+/HwXdkewW9+PKscynyhorYPVNiSnD5+
pejdUrsBjL04E/pHrSOgP1q+pinLtTcRLKfqRxgCiZErfNepZN3OEHJFDJJEfQZQmpJJSUO0Gdo4
F9vqOOVqsY5xmbw2MaURfa9vIM54+80V4VSPfXIrtE7fPiQ8Iqdg/SOIJO6YKMvIed43OWA/fN4p
P0YKyZxMaeyEaXYwkv3gqx9Y3FKh4IT/ZCuCoOD7/lbSqqqnmA64v1VaomGQtJ7QLIg+kJLAl+6X
vb4ddjvoH4Q/M+oaeSbNYzPwclCSaZDAMxvEWvxXQSftlGQoXMUx6XQp9Z3ElVPpNVCfx07S1gyP
XR9jgNn9B/JZLtuXsKNqfomLzj0nqL28IiykIZ7mWmDUQ8GXbtbz49+Z8C46666Obmu2JtdHAe4Q
gznWXSbL2AiBx3Kw7wXRxEJD8gxD8jtB8mQ566PQvLVEEBwO36h589IS/Ky38y1zGib3bewp1MbH
tHS32ixewNkhvGX56igtN8dKdqGx9n2sesGWiMMs69Hhi0xQXFH0cUvGxDJXLkD7wdYD+uFTsiiU
jBVPzfCvr/zH8XmBFZHxUcqwllwpUiT1TG1NePvbVd4grnAChKPZmtUZj/UMemS28O6WkYwQ1Vfi
jDBPqbDEwsfKuh0AM0QAqdfy89mS032rZQSHSPTRfyztlN0F//6yULx7VhckZA5gzb0EkiRFCvFs
H1XCC1KJpn5Bkwp7zBMXnPR0wfKb/4alqYEadpRYyyYBYa5daTJp9Hc5jprxc/HkFsvyOj11ZiOV
ETBH87iG5pAWMrKEjFuCcBNDoQwiFpcDO5qeyT5y3E/f0G2pW9UibDboI02B8eQ2SEtlxlYD0Zdr
6UkMhslSVWhhyDCed8EpmyM9KB3GOHO10zEcJugY6032t8Tp2+ud10zMDKeeTNY6caDgCV8Czxb6
X0Snrm/cFZuknf0FiV5i36YhVTjLwjH9v+hiWvQcXDF9QhgGfhyXe8qvV/ORCBo+b6dcjXFeImAU
n/6u5Fczu0GIbQKQlw8PNxrahAbQjhm3gli49bCIYqPp0hRby8Xm2TfUc4TMa/3cg8V/mUxk0R6z
qfYpV2eyfvUi7Khz4DbcPjw8S/SkLu2MM6CoLmHZTuIEKAzQUnLGKcoXJiC4IBkEbQ/WICF4anHd
2ZExCs8X4d1/jVlUANqgXqzhJWhDbvUSZaxZOIFjMHpEZ5831Olw5rdcEk4pyY/LOOaQPjizMYpA
aUi6wkiFOwDeqQHTSZCsRn2eUuWs0jIfbaAjxHf222crkPUA3WNbTVJo6XqHLmZkorwwwhMbbeU6
T+RxHElOSn1gjfQgs200e0JZI6TskEdej+MeoffeT8I+X8MoyIgzdDEq+Z5Nri3WhEp9KHAjWmyg
i4prpEJ6GryYA4rJ+Z8hPXa3Ge2fzOzXG6XEo82TVTu7PjbUMxZWK/waFlncv9BO8V/qmchPnAt3
sauMy0QKRV/kSYd+r98syMiRkx3vLrfIjt3nb4GeeG+HxKg7Yk9+uIr8ZhDmCAo//PScZ4lDZC0Y
VdUwvyB/J1rLdtCZZN/QVqhmNT6KHnznvS9wAJCBGsebYAeLhuVTTHlxzHKBJOwklsPTn+1m3YXM
axwk60+SRtWnXg4/pawc+DDmtHvY5VgNpgo+A0jfrZPKo8TBIDa7cYsQXzX+sy3TFyRaYIoPyTKA
4nS41f7LmO0lyo6HWxcVFvmA+zN5klGVXmX6qJ2lF+egig3f1MgzqAxmT6sdb1UB2vPvG4xBMbpk
FNc653jKJ28duIp0bABwtzQgc7xwoPSHUJPj7KNUoyD6pQ9fJxoclbjBYLW7bQJ/qBT06ewgpeK/
IJm9aNOzQUMu2E6XCGmRlwOZFNVoNUm827fzji5lcDJUhE5BedVJKlbLAi5OgZBgyjNTQKCNFk0v
g2a3/ibBftz/ViO1SboNOZ2QZmqhrlcD83iOwb1JxxpKKc6bBwyzvhw1k6XSqkltFYhIyVQEbv1v
CQ6TnVRlMOySO8/hQXGUNgKNeAzwqZQVYujFPq61x8uVCDKrWKpI8wfQ+k8MQVn/5BmQsWG9fwZY
bGS+1AP0JRxKYy7pV7yH90Ni5rK/AyicN3celnz1Ryt1WplUo/C/w+vFU/xLw9L8NmQL9moC5O13
jII2oEGCJEfL8nodxRVp0bEwiCLU9p5BhW7v0obfilqLWww6P6IJzTvm43lc0AVGI8oImxiHBV6r
ReDTWACg+DtUotjfm1tcF5mAgdF71h0XVRgtZZz9+jqmnVCK2STsQh9wsGS440dJnNFZUkl6NLmz
SrMBEtdD/RowKVAIfK++VBdRlhm4Q/nw4RD/j95m0GXqYPDbyRxm/zXfd+aPIaWociNJgAyhz1bk
WSoXgURzzvJGipAzyBJjKNgCP8hUtAxeXVNOQyKjHexQMlCHpFZmcA2owH82YZOv7DRp7Fwvz6sn
SGdjnG2FTC2pjM38yzlu6/xBsh4aInEr5zPKkLKUq9HK8Sf42oIho6A7iWyf88I9vClYcxK56Q6I
g+sypA64wTW7/Jpxor6PeqNlO13cLCMYrO3ag4I1YVkXxYZZRmK3NskGNnJ6WmYeo6CnhEL9MflV
7jrZoC1VYiZlwd9CXk7vk+piaQLm2BdY6T3Z/bjmoSrblbQRORd/a5Ks0/0P0C8jEbxkAsR0CE/I
6FnOnEXHN5qAg6AXI6bNu9+4KSzs+GoIO3OLQuot4LLfYuSujNjNd/BPDY0U1q42W25jvHXw0pAA
TkbHDuDCtMZjR54J0DZsYIUGDDIn1mbQlhg+zhfRXLqvqyhO+XKdLK+oxPfl4WCBdnJ7DTQt2kr0
YSfNOIjkFpggU4X8ABn8LHpYoRdat3/BmckvgdRJge6lGTGSABFoGrxYxgtWW7PcGKXqNas17u7D
yoZPVKAzyZF8vH/IG/LUkTIR0ICiW3VA0OPo/FuaZOip1idQ5D3hyKtxvQgY+WasgmuYyJZJDol+
KxRlElPl4oOiOlBhqSZzDp6p0Vt6+nKYikxhtfGDJ4N5hiNqoWaANBnLQdcdq8QWPnVcC9FBYemU
PjGWFEkFZ+hfkhOK+c9hdSSsHwA2ugqCObLTf5z4UsB/Fl7tPXFdAyhu9QZJ4pVGA+AQO25gSoe3
+uNBija9tNdND0KXYGBDDvcHehH4q7/l739mQTN8pPrMG+ZgnnjcSw4feT43hUr/iijej0sVzWuN
oy3B7OR47IpIFP8nTwkWmzi2S9CgKzfcPzRVlvyEjWy0dg9bpQ2J6hkjZiRlwEu4NmajsfLxDk/j
KjrON8n3xtJtgr77NkOv3fu9iz0d9sMx4NgCvdIijlGiI90ShEZfV+teERn1Q8VM/Hp9ZpsqW1v9
w6hhbnkXnXa77xqXweDLjjIIfugIB9aRSxbeCrF9aRUXQ9OETOMQ7qeH3uIUOW74jL/YjZC76aVz
dAljp8unKIrvcP73sm5v2CXhERbUYgCAyUkl+wH6UQ9GY3y59S81Z4UOOTUeNY9X44jP49nZ51pR
dt7AzIAvs5Q5t0mvK4Re1YXF9yPxrGomZhnfFDtgDzjvU0AvQXPDt7CkYkCiKcPbwm+O2aN3Q31y
NcDxcYBuO2q2LSLVL3ixgWzMV7A6Sz4C8lhkIhLgk1NKaLLuxZVG9uUHFUzytp1PMFr1rgN+2eHn
jJJ98vjjPUAeI8D0QdN4dD5k1FEN4/Cj7oofQpZ0Q/84k2RebLRLIfXEQQ79r3Z/ESsIbBUzhGFq
jqsHfhVCDJdqGdtu8PeVlydT1iiNrjI1nXFqR/rabFPb4BxfugqMzeK25SHbG1j8mYWC1ELM/J09
nl3svWtma3xThJd1SQYvbVxo8yNayKmP8JCQcg64RKQZVLXiciCP+YNz0mxMYqJK5VzGLrSJQNEg
sYT/IVhGCRi4kvQZ69lTOxTMXTFS3/pJFFU377p/mDsX95BFTON3kanuVGMhxX1/mCD/MnJNwUGj
mWqAK/M/J+AVN9T/eej10UQWDD+9BnaIl80Mp+egwUWB7EJX6uyO52dR3MRecxmfxlRD/02HCQDw
L7E9joEHMtLAWmYjZarUheCik5Z6qiSyh/hwOu9tbRTLNnc3j+4gjXvkSTIE/oa7Do3YB4tmFEdp
gUafporXYDhAc9JIEnqBIwANZX/rHwrUwffZQp3hxuKWJqoB/GBBVe7y0yi8zgk+TKoJN48S7t8x
ShC8i+bfDBwdEeSWcuwujmKn5LCT8T9iwcG/vhpyHtN5lw3i3eefyJ81x2VcPIhFFhxYQOukMLbs
DrKkBSLPr+4m+vyPl3jc9aAnGUqhgpCZ8PMxPmNn1aLb9U/eRUQW/tYijDKxHOBGEC2VrXR26bUa
mNu8geZ+ltKXJjRAumx74alWBJU4KjRNQpEsFg6Qv1gbKy1wbM9ac/iCaIE2sFC67w8aF+axETLA
Mmu9U7JpZ49ul+UbkfXUwKpKDLiBIO/JV6nsdZfdH9BPOmA3NIS8cbAhucdAdWm0uUCvoRP7KCVT
iNbAJ9I6T6svhFj95sCd3kUKqdqMybDWqFwwMMSX5PopjiKzDv7ULC9cXE5xtOtUFkYOWMc7xFxj
R9/fzW6J5ZX1FCA1Ii1KzLeAf6OyQrjqYxvB059Fcph+m7TZ8PzWrfPk2B3rL5iIyiEEFrKgl5ZN
OAoeQN0hOH3d45J5wloZds7Z2FqPrU8y4z/TXVZ++BJ7e967mayc2TCNfsPJ36T91qGlVuQilrNh
nX+uB+UPKfengat3W2EGY4h4NiEBNz/EDh31Y2hzwXQG/KmaraeosuEkU5e8EwO4guJ6gUu0exuK
lsGh/+4LagtCv3gMF00ZVG3e/oi4Y4bGeiGWFE10la7UQq8nncF3t21NR9SYdxJKgdodk1SGN8ec
eHJIDCGWmZhBbbIa6RpjbrOaE8sKTXz+8lnaLUJNpEBEYzY3loHM/HQvLbdR8xk8FrQvAh7JSQa6
ID2p2cHSbzSbCSCy6kuUT99hNr8bOEtSoujcStYZ/akxb78B+bEOaGBIUjpZymf2niDdY59ipW7e
tSS7cWjZmBFpgbUEjZD0afi7wrU3n5yN++olblOgthkGa9ng8XSZDO85e/wtpd/6BgkUNoNg9/i2
0j31h/PJ/qDS7HhksO+UzyurqVdDRLOwWT1vnV41cZEA06KHG6pxK4ETHZDVUzNVri9CXJnuewT2
tk9TSS5QmWoVvlQ7zd9rSljnZ4UfoqiUMqNupuf5arwKfb3Jj8XAOjKukmn/CaxjgvMx3hZTfPcw
euc6FkY/68Zu1/utGe9TDRDwz32oJZzMzZkrRGJrS+m33YrX9UjxtDhNhaxJqfdzna7m6egO8EmW
zr+X/7qGGgxlLUAtpKj7Qyyq5v0w/eHeh465V1v62FfKvb/zN5hMLnQ6twFl0ddP1LXFKbZELtMe
f+u/xS4p4OvxYMJJorhAHl3wbttJV0F5P8mL4N2aa1tyuYiWPuzAxzpXxiYYXF2MLLhWC0/oGOjs
2mEkUC6XaXiTmOXOjsQQ3xTpxQBuYf0nhllwenEW/lyKkT2jc6Ui4HAoIyrDtV8rKDJZbrR0a0X9
JC7LuPlPNpiK+5fyWGbDWKrtJwpXE9srHqxrd5FNxPcMmJn5UGSaUEWQePXc32KbvC5+HdphnI5r
YIw7RYkxulwNdS//VDnqNWpvik76ZJTlc5mONZuzjYKNM+c0ZCE7z7XyN/tXmxtuKDV0m4uLtf0S
sVFvo9J+RzfXGRnMTSkLTAE0VoeEVgZwtVKD8gaf7mklWx601XILEfcDZAPPq1pMVAodjqSkl2TZ
EaftF2TtK7GOAN0hPT7jGQ7zqlX7yEHrjJq55USQty5NMJ578t6GXTGGH7NbyRi81F8qPniEp5oi
BACqLi5rT87Oj/DmYkYyr3bwf42z9ivXr5xP8he+a/AdlT4YD4l21kXswMrRHv4IcYohttFOTfn7
JLXOLzbVC+lMgBAa0JptmRDXEmy/Er0+DEzPTtfdvsTFZ4Enkyn0rh5MQH8RsSgImCVwi5RDLOk8
GRhfBo9ZCpqBkljBtclvY9kJaWVLbBRB12wbevbVp0jydIg8GYZKzSn86mnayg8Wx+cZ4EujhFPr
dSyXAAFzDQMGwsNN+AFlXJ06GyOTqGDuWt0NlAx/+L8JBm/sXeRkWckisM0bYPpookxbQauMU2u5
cpFor9D1vLs83TmmnPbesHpl6z6n9o2qB12NlW7gtm3exvg/Ft7uamEwvNk5pYIxL41ZML0nJkZ3
27eKg8wX/guKeojMQfm1xNx7OfqsknNFO38kkGE9EqQyYKq86gxeGPJreUb6LgijJFF4Ec4MLPjr
xsjbDM+/0r/wEeO3UiftDiMXAQTlCQtCrg1cg7E+NyzutF9+INOnSGayam8sDjRO2HRMibT/hQaM
9UauVbd3BL/PAKUM70AbM/HiAN3GovsGozFCCBfMj7vJ6+3y3L17Gd7n0DfmW8JKYuCn7nPiI9cw
9ZS344ToWzhD6hXTXUY1eFe2a51RTooTV593L1TbqrAHypnHyDXqCdHAHrpUmAFfsb2bKoSDZiQu
P1pxtff79FE3SgEo0+YfUes3jiyZUQ0k2tMP2Ip7zA8iuag5FZktVyZewg9Z8Oqa8SR/WCqtAdlt
+wDLvF9ps5ioj19jzaPSs8/EOJ7G6cz2vGyJ1fcpWSZqR6H76zetx1Cash4uw91TUo3/2zBP7uMQ
Hu+w0cld6CUv0PrS9a2lJK+9FtKLcjPTP4fIlUgSBM7hT9yxBHBAf33nAy/GftwqFNKJn32s0AgC
hCSOTXX9b8BlEzVff1bqtPLUbI7fLDFxhYnWt2gniIxjVroplKZdWnACFbJ9OoLaqiGJs2FyBph+
xAT+NfE7BgY1VIzhGUG+sEvO9U4rOOLgYDxw2kNXXhwoKbxhlBGd3h9L5ANyQV7Y1ZZuuxh9ycQf
pCGodzxq+cmzIzfWO5sOAZGJXlSjrDcCJnxo7KGr74Pz0UhLfd7+u2lcCoKxEL7IkAP0d3KFPTma
ewDDz3pW5hK5F3c3m2NYI5oWDMyRgJ2eKEn2AJOTWtsET6tXI3f2oY2UBLR5jOE1D7+HoIjc2XXN
AmCrX18QXeeDllFltMr2jhb1Rez3Eqtjw9O0nP9l031cj4tJHXX5mM9yyGXtYUKaheXA0a+Rm9UX
V017pBS1eY/OU+/WC61RUX/Oo8s/iGF8SWC5e491rbjQWchZ5eg3ja03yjoUmWtgt4CasgB8VCLR
bapeNXhQ8kch2GBDAeR+jIdm2lVwWM5YlFYOEhVDq5YQz3zfQYp7fDdVOfhvZ2W9n3zZmyczSWn1
+UOBxDzY72z7ewcDX4cWY4IybBkVnENB6zf+iF68OvmlbgD5yQfi/av6FJLIp3nmcG2D+PnBfCq4
J3RX2F4sDOjfAQtqdxi71pUmK4tjIynFcQ9nrVBTstfztg0FNEQDkqtgCk+U1zd3RPtIYyzRyVr7
T+paqysaS3TApCUcSRAcAcWWKhkEn2hu6C+iyqj8ubzNP5zLWYm8aOvKRhoqq8viBwd5+gvfRXjG
cBrlqZknoofJKz76SOkuMdEOTRkdw77mHdtICcLXgNnH37oWsHJXp8Z8uLvhHnDY+iIR7nZZ9JSO
4itIBd3LMlqbEeFIZfjdDJITvpqFLyO27nEBY6o6um48zuK+IjSMT7Bx3MNSescPM5OwIVMBR7pS
+ScZNLujIYuLEwTX3q6f8oIcJlGAkS1OQsfCxvP3VsQDoM7R7Fz1Ldd61NIRZWI1mXCzDXYJg4yV
2bre9pHgj9x+AyYOnjfooifPeXKQeOYPIEEGOq+woZDCNtJ5I1mHCGjI6736Jp32QzW6NPTyniQP
MsWPGlcqnwuU+1LLNIoUojOQMj+SCzsU0b8/sIow7azYRGihJb43NKRUT0NPdZGqvp3svx2F85s5
9uBrqGigMqCuelgSy5CFiIbLQJvRgjSm1tRd7q8wkaA63J01etXqcJawN5JTnnRLBHO9n4l/hA3x
JgT+2CRCOca8UCbptG7f9w0vvL+5NUJP0QWAa8dyqHKEhNFUq+ntgo5Qh6xrrPsB6mjBdSz8/0jM
TmQHO9idhYNhnkOr8dnKAuTnNPQYZljdEJMcz8948hvGoXUXwhpMAwpt+6vXPtFDAXrflcjo8ZU3
atJ9uEOxNKN07XBWuAenw5s9SPMH2heqq5oZjMBYH1QqEzGlrP3wBL7CJdjVjvJIXbJ4jPLR1Vs+
pKsp7N/iZJJc0xBEFewMXoOJpd2EVMmiWvIr9UkgcE+mqUA2fXAhKQWhIBlIo3Q/ppSJ8sEUdr82
m+/XdpbE7x8IFXqup2I4GSTw9qfemvKB6Bhy346pbb+EP1+9phjhFZSSb/MWEj6CzKE32totz8AU
E1h52cfpSV/ibKv7iUmtjjjNSYlePkwCF2euVkrytY4L6cIR9yzc4mX9esOl1eFMcGI/TBRcnte9
bPagdi0ksY6eHgYRjljiGl/5a8NPcxlwlalh65lkFJYHUVvayCbYGO6AvUo2+BqRJkYa+OCVlXuk
odlmSmuZ0IJDJPLXp89o9CTGZNjXBAxrUQoizGUewsPPmAcgFcLK00i7cw+hm5oRCXFR4IEeVcwj
dmEE9Ay6QFhJiPcA9zY5SzF+HZaZvnuNAJtzFU7Vxq129CZDPaaRw+ABNlVHC0k+j+dRUS8tPj5I
yrJp+WWJTQJNLRzmy502GwLEFo06qxzPYnUga7MDPRLOoEdTD697dnTAtHW8pXFyr+45pWJoYBRJ
1AubAjPVETy+SXmvicT3SegNOM02wBo9VRAm4M/HtPAly+1wrje8ETWfM5Ks9/99FGBo0xM1Yiv8
bN81D7wgFQvVSML6srnC69LrjsBQqOmDdSis4vuqY2gPraAzjbgvzzggsC8sTBZ/vyL8NkDxVwia
6twFPjum53+FbL/u1iis++dfd3ostekL0f0JUO6HljFEs/bduihCgaOumO5ZFvMtV7ts3qfr8Cuz
Z9gEtNnf5m9bCVGgdKjp3klCvSi+Eukwc5J6JuOl1E/D5YzWyQRalYtGTcDe1pkpZbwWuk3IpLOb
yOp1OdH0p8Ydg2YmvbDbyJZUUag86b2pitDoqWMmoBbbZA/o/+djIUW64gHMYeQ6Y1/Fqwp9NKBf
tzv6p8Jyk7kKe9XadLFhwlkIgZ/BO6fj0XR1Jw4qBGsUM/+FishCpU1/FnXUQw815z4LhyzXVz05
w9Y9ahxtWOzyt85TFVa+xU66Y4Eay10pMb8XsqANPFjGFy9jCPWsF1+NcNAKIzqNR0Sa66dzS19e
V3PXOFet4XmKq8+BDMvn+/p+1cFxA+xBQZbO3LkOUnQDF1XqSnj57iLwYB8nXv336bxjIoVRWq4Y
b3BvxWlmQWxF42pWOPHvGRETsm7zENKqVS6YAAQjuIdL2OrUpfMgR472LWux8wgQjp6JX2bj8+OY
pBokvfYGzUyDj8lq9gQsTkH1+UMWaJXGCTwxu/ZClvXg+8co6BZMFqhlKwuj98kmqN4tQctYeP9Y
4qaZwvgcD5OjmFSbsjvZBq/JGRjg8TLtHLsYymoVMpeGpphAtdm917O/JEdQtV0UZlOOEJi0A4ce
yQjK0jbphuGunE8cEAH2opUjNKR/I8OdOBMaWrI73xERTyMrSYVkhnJjJ6p8ilfBRBHxBBWRBnSM
vAH4HiOWDr3lE6aCy6pa7G7WvHKvfSj+V89IO/tjj/4L01gDRrh/ZlcS3z/aeIO699c2K4xz9WOs
e3m3sHkThCnM0o+o7hYZhOWRfhaLU2IqH2GR8GRtWAcVm2IoWvTbv5F/NIlaS3EdZn2xs1f3c6fX
eBX/9n0oVrzQDH99dzzTVxZcZ/e8D1my0ZRIIKq1rUed5vM5Ovx/T7kEwz36r5JhcE5HRekdWrKE
eRmA5GtLLIhdAAnLmAwr7kjtln4racE7Vyj+YVeGLor49PMONoO8mCDU5ZgNlr2mcsJF94ArANbR
D0Mfma+DHAtje8ANo5twvgOih0LS0g9F/tIzJSePSnLj3Q1IJRGMLTBSt+FvV2gyGyMyNexUzRHN
TlI+fe8JofQirrWSwAWqh0+egqT01OWaMpGnf6vdxdc8F5J5bu8cG18Jna56vibstnv9SzqOoLMW
eDuGbHaDGDmKvPw080D4W4fFwawrB/P13YLlhs9r30K9OqC0Oy4Tr8LyOtdi36rLtCzQGJbR8tMr
yZWgrR0aarJftJFlKN6O2IdCJxzOUieHfrzibfsFS/V7IClPL9wp9bNI/N40CS3TXtpC/C9M8wBc
Bo/0IN0v3TwhSc/Wf8Yinx+cWnH9nS+I+Vp2hq0469JtoAiV5g0AhueVdKm2kmMPDRUpfRWVi+EN
reuyzJmJ6yCRAkMigP4vecTXCsHuDqsKdih7zmdhGZ65x6i4eu4IwpauvQCgKd4csKymBRtV3JBi
OmKYM1PY8jcdL0eEJsKpjRKUaXmRIia0a720W31yy7LxGKsGauBQxv28PjuvgWRAl2uuFvOTzZ5S
U7/x/EAks+690YsGcynEWT2TaDlzck19ivE509Vn+UD3UqL7qtqlsGjLvx7iXfhiIZ2inTQBLQLi
TjPVDERrUyNyEgCP7uV1qdMsZ7q3ej86Gk3muMxDAqSqDBwKMVCZTOeN3643O9IWCdqT/eaTIsN4
Q9R+OgLB9ygmEepB7zTUr7aUjnJfMqTsxVDC6Ro1/JOpCiCHThPz/edRPVlFJ0hk0+yt0IT8INrM
nFoZp4U3QCALoN5LogbEbBBhFmRw06yaIEVMt1uZMq1p/TIvOJRWAHm3p0L1AeTAgW1tSt+TVvJS
r8OB7RAvFeaZVcpeCS7zxAX9bz0Vfid8rTBS5G/AGHoX6mzfldNZJFQB8cfwlfEoiux1Pw1zEvG4
9EKUZyo3/WnXPFAx2gKHe57fePRSVFeZU0GfYXWsVMdj98hfqBfGcMyFy47G4e1bnXXs3QZeq/pa
ON2S96vQ7Q5Sd0aw/47w88z6vwFeZba8FuWmjqgFBcGLtGuS9G9zUkWqswsI1RxN1mAsTz8vHvcR
QR5S+l4hgihQj35VXPr7zvJgqaxRgDpU02LcNFoBz2wRbOO37z4JBShplsPDlEiAEhUDxtnqKgFl
VdL4kCZmQfAKTdDUTjg5eqBrtvDYSxpyT07iyhSfvLN36Wf0fBMe19R+4qE58p7OKPze2PERE4dU
4X0f6fFiqs7S0TAbL6eF2W9tsRpjrlENj2vZ8aJbGmayosAgZGroZVSOxBaYJq9qujPxeSrrQ3Fv
YHdVle81RQErmzfdMUgGzAtIF9B4oiNcgkE3XyAx8YC8UWlj5diKjxd+BMD7+cjA53h9vhenBM0c
yJhZJlTVohREthwQIMVCGrKN/mQbKJBN+kg1/c/VMXDs93KNs0/7louAQFqVMYlaLgoLohsMpKaw
TlpprcZCukorR0dDmU1EbF5EtepY3r5cblUBw6IutvzOK5i09p46W7CXswaNptvK5sTB+buG1PTU
Jbz4IpjJjnqIjmEBY3XnQ/+Ki0XuPnD9W3lCttw1t5gtbQsHebxqk9uMfWdqGnnOefd+Z5LgbAHe
/UNy6KtpN2A60zPKUtXlVpaGoTiWksFLEhe6GbfBd44z2TOUzcnLQs3D1ZWZADJ7o0WprVnSRfpM
i0k+lTUXAKFaiaccgRP7aIOM2GlhQtC/DNyiJMtp1KIctjeIsaaNMXgFX4DoazS+XgggzJ3nLgGd
lW3ppdueuEIFdqXGYH2oxDhMfiUPVXAoKBhOSqi7FrUrPxfuQ9ocqxfmo68p7vTdxBsxT1sPvjQ5
+iX9wOf4CbFV2qW7cnvcRjLC4uQaXQOilL98WpouOiFXTWhdxw7wsHpy/w59Lo3wsm9wFOH0mhbi
XgmhSE60/WItVoMU4zaek/Ox1pvZe1uwnpouP43cvGsbQ/JkzBuXgqxFGiTb9eEzeNq/vW0WIg34
XhY/yDskTbMcu8XeFbuB067qp7RlWY63HtJwlbZ19p/QydUz+kzqlRH1NM97kEDfY/F9+TWvGNT2
Cs1CnenyCPzI/yPTB65dz8hC+XxjTgB26u4uAm3onQ06MjFATIzSAE/WNKj6EXj0Olewdjr/3e0n
YUz+H9lrGAvjxEnkUfIVLq+Xmvgb1nB1zzkand4WNsl+5B3QuFalKKgXoeNeRDE5zxpOe4+edwqG
bBImkurBpXAyVz3pi4iaIhPG5nw/W0iCCQ+J900qWrBytyTYmAhplH21TL1Pp4SdN6ZoLHT/kNQv
jkhfJZnQ5yrFBG6/SmN7D1usvZB4xk4vQJRdO9w6TQQOMhDdxy0tbPsD+N1jMdWeNyN8igTty5L3
WacWlVS/tHUDDgrBLDlckA6YzHukbBF3VRihNCVCD3AjWKwUyir2qBYPz9EPmHp8Zux+6rZfchg+
ZieZEGlCi6sIWBhkWdM2cSec+2c6rCIcb2/Vf46Bk4Q4EF4JXSemotiEZsHh2uQIj7TzhYDsXnfO
zYxuddLF6G88vd1hBPeqInF1A3PYBP0vq6n3PMa7N4K0Fo75y1EZxN6jL++cMBpf3rJThqF8m8Dq
QRKIdfcegMZEF2FQoGJgaePeTIz6vGR393wXuAPkS3AtTVv0Wxeom4v+ge8Ggn+h13KBi2f4ot4+
0IVfXuXBrmxf6xW5LrYw5+NoVtEFyvYpyLaaq2l7fKQYR0Z5fhD0nWQ45TBEJ4FEB9pYuX0z1uOz
RxlT3f36IV08K+cC+ZNqFDElNRR2jfoGRbSRfNN5dlew1rlz59b2GB+2EH9YhfoiTCt7ZRvEPubK
OEpnT6uJd3j11ycIRcq6qAX6pF1lghNl+nc2iFXu8vr1ABgod1hqO4GduFW5KNj/qEizQPFSCdjj
Ey1JtMBsjlbDYsQxRCabq+C22H0Zh0HIcsTlEyRdc8Z/5mRypaZn/d8u6eiGKgG+peU/QIov8PCH
Mz1nVuLzqUkSnYK3Zm9BZp3vyzmzJKFZ5cz53AYbwAfIkF3TRW7LudC9lDAxeZfdXfoODuisFTYk
ZuMBWjWriFp96s6kSqqQZUifcH0J+qLnnhkBC4XWgb3gkpDSYgi6jHPhn2X4dGfBxh72kk7VoJqB
wYET8Pr87iKYDgaznIj33EjH5OmnMqxDIgQAAqUD65LIA/HNRSNIxr+ZIKEyRYVL1YwzhRp4LYJt
vPNHNL1XQbO0j10f+R2yDWrEaIDpRYYk+HuRtRWRt3VvG35si3tXvDzdJ/y0Djdc2DHIVNh2Xvhs
ZtTRjLrz/OFEns6BeXmLmQq5tI11sT6wHx0f6n8bPSwAI7GqqOM/PPrSHcf6kXCj9GaOo4CgMbOb
OBtx8xCurl9zN9RGe2ZExq0MtmKeRb5nO556PiSNJkIV6rGmIQe76yK6pRmWQq7SFZiWa3WQA58o
L0CH7KAMIBUuT0PFSiAvZ0miHGpv6m5wrUgUWO3JTeEa/8H/SKGffZFz7onE5dD5O9E/xmCc0KXG
GY562fb1Al5+IPU6g71ytNpDGZcI6hknTlbyJCM0VAmBYQbkdjvAbKetRsv9GDuJCr+ROVsjC/hT
sQHWO7aZSWrlzAPgcrGn+W/UrHUFZPEZ/bYxrky/z3bqvPaY6n76fGnG20eADBlvipsDGew9d7It
VPmnXZ3CgSowL2Ms5WkLPq8+C7Hkch5BUEky0fi3/spxbgqMW7AIfIXo2/3ph+2OMHcmu4QGT6Uq
9drAkqkfQoyCYK7W8GVBQf3mD9WMYYk2JpXf1IKbqAehRC6e14HIavhWmpzyOp2NzGTL60G6JFTb
/HlPnDoXutT1eeA0BzU+o+Y4m1qJef3eEPnp0MPbL2vt1dVFW7OzydAKuhw64Fp7GqjluaRZjWFy
1jscY9VLw1JcnuHw+7AzbRCDnV2L3uwkgcclAcBwkXfQqz/L+VPd5naFssU0ei8+Y7nMveYQ+CiC
+BzWrYLAS13rXo5+aCd/KrdDFHeQGkvApykZaJOV9X6UWYNIJ0b5nbi+bqd91J7PLYcTNPKOJa+1
g+ojBr/FwlvXF+yB2YupCoF2FgO+ZQ8AKBBjnX3DLX13wY50T7LIt0FHikX87wakdFtHAzRzZEjB
k1apX+0o74WxLCoQ5mHVuB2XV1XMeB9RR/Ygj/nlvbaAttHJccxnaOqiLN2i5Yx93DNeIuwSgS3/
7Y1jzx6Tjrlbz3mkoOyiztBEDDA9XhLSKDsduDdRJAtBU+RLizr3LFzMVdWinOHNKYPOdPt5f9zJ
FKwUmPvApG7dB98vNX+v9APAQeUalIBeltuvHHRHfnSZkb3E1fzYlqVzXTU45QIywn4Z35DDJbsi
r3zT7qyKESaZNuHvJGdrKmxzPUaHgbMDaMcm3OvyOAP1ZGf/A0/4CTl9YCM0gJEgKqlxy70c46YI
ibfGBGE6uz97ABnEFeZcc2JxgqN39qD6wg59BxrxOLMABnKsrQ/jx506rnlfd3NKfVbfitksJO2o
qhdwk3QrKMXA/8IdO/94uWwAByRdmVZ9t8stJn/VIyvXjkMq0U5IJdgz3nbG2/2088sEFFS0TxjR
3Z4AJ7kAoKItIvj3Y6VqcM3HAc4y5y0v+EyoduUQeazB57Jf54IXkMYH6Wn2SP71xtBNpJzNAeGw
0sS95D5DeQP1fXDl19RVFENWvmVhLY3MGQTmvs7opJbEcdOAfkihwAk5kGNPWS8KHTOuuVeZNW/0
fA1lt5MbnYTQmc03+1ihwy59/PFxNivz+opA5KcFd6SL5TfFv15/VXa3X4mWn+Ho0IpJ2n8wVp45
q+PDpuyczBgH6YcKcSjihOK5/+yKH4aBmIul28ZtVYeSYckZra8BFyKoq06ONYOdJLtqPk6Xi7QQ
TfQs4HKxYt2FETrNkQLQ3dyo+MktTV54JRc+QfHQV7YGAy/tRjKhqyljxMj/Mt1dRX1G5J+qaffm
58rzzkM7lvwV2w+szNdP4pB07+O8Xs6mamcaIfd40qNNTGJDZdoSc0rVx5hJX49lpPMePStaYwKJ
ORgiStJ4M7epi7cNOYg4maurOGFPmvYbqGNqPGPfiVqDdn81yIIR1y2HGVTJNDMVDkxHd/JgCx8D
W/XJELuB87gqBQQ3j56d3xrbFSVMPPxR+sOCN6cbOSWZwqPOdIOXQqBlpGRboahQ8LH99X2VY070
5smRF32vGPBjBhvZr1FHsDQF0Sh7W0vyAPZT5BQbGUOx/PP0gl4G6Eu/fmsspq75L3fhUgtB7LrV
xghUq/fdswbyaQMMlOZpKeF6XZr29+Ncb21tlxSNLi6HBY+P7TkeyZ8e20+l9bphOkSnRV98yQHK
16sYMekcrsetkXDhe8rBwI7QtQ7iPFj+YCBTH749A0FTycpPOBF84mLeG9l+Io2rkFLLRy/HCDpm
9y4gSnut5+9PGopHX6IHtJA+Aa1sWFNJ+6UktK6lvRoJeyVMymJ9nBvxpj9o6qlZ1Chx9lphXI0Q
+K9YbCGcjcFfVcBGJLPn6XzjJ0tYMoQgDgrIjmo50M+fdbIazS/kXz3AaOc+ZLWXVJloPDiaO1bo
sRc1Pe0Bo3a71p8yrToZr7MASPRghR8+WrYjLmSfrpfRfTiz3E0OJudijXLvHDyc7+gf3laOTlxu
CEqG6xJHFt1v/xvFQbbxB6u/sSP3aDYJ+PwXcVjZ2LuIu3H7wvUtHUF2qxtQJcu+BH5fCifEOyN/
Rlchw0S+pUmh5E+EauAZx1bEUp6Zj7LC0gRsUR9ahNTTGC2L9tcNofIH7SkgbNRM7zicJGSG50V/
e+Pr8JuMfyvAjp4tnOegezcwVw37HK5G5Gr0CLyV5nhv1lmseUg2VjivzJl5q/DEyelAx3Wzbivd
IUn+jQg5HwD+eeWfQqI66FmpWVlYN1jZnCVZsUnoWS0s0wmnN0kvtgwjbwarbEzVRGmwTeEJNoTR
6s2FTVP4WxAOpDzvs4LugU/9UX8LYRvLEpn+Xeio36mQ8LL8UuPja/8WL9LnRveNAjMgzEXScPh2
GR47/Y1/IoUPF/D3gIIiugCdfZbs6cEveLaIGWbP6t6JqhhPs8XRhCmfVDMB0yK2GQMS5fHhfS4i
RilaCkdiENgdMAyebzmV3qD1B1l0wNrjl98soYQ8w2cd/B286zEEY+/F95gHj3OJDV2kxcMseKfX
e4YMeLnNf2HGbMWabu5Juu+R7T8d3bkTp0Zmo+w1JO7E8HKd/5Batu6NOdlFIvMXSRptAEa0HmJs
455mHBLXKjmYA3gInctMzRfrXWROcQ6YykQuQ+tvLMMum7nfUcd29o+3D0Dk8CfZQP2r3qP/1Bxl
z0UC8r7rMiiReByKAJ5HYPRywoci+aHKuQqI+Yh1po9czXUAgfSkFM8onyBn5Bw8bYlUNO6IQ20/
ztTLT77k7NnXM5+P+OlKAmoaXHWPelinH6GWqEH7OftHnI4lCF+JyxilJE8o59YJNZy5d/Togns/
TTGRqF2+/oiDHDTPRtptoOt+5fjXzoi1WMR5zQ0eRjVM4ksvxyRP8oVPrrI0xRzUnUlACItJej+X
z6lQ/HBkG3/KhEm9qizOadsJiAqftPSpw8CafRNQKgLYuIIBOSK6eh86sG5oz5k+2n+oJRXyq1k+
ossE1Rt8fzcsXJP1sYFFBJwACz0HaTYmSzgOkHJYJIlrT5lqPohnv5+zSKryNfB6eiRV/853xxzB
DmIneeI7U266Iwe7a5PhjoTB4yNSd7ECbJFuJIFR2GpROnJPkGPM7Lulmw0i2WRmJbfwI6aJENN/
VPZzY/GhLIFN2DZ0lSf5j5lG4mBpqfzsJn2rkFsuN5uFSE0j+LPzDDIkcDKIMFWGS/hjzdBFZlzb
l10WMgb7ALDkyj3jwXZ54X1ujVuOJf6NcRb4rZglLvtCV79gqVQayUp4MWTegKDDNseNyYDHsFim
Usbt9+BkZCQtfk8OzOww/vYzsG7Z4u0NC6OVU5ECJ5UBdo2EruaLNE6VzCgZya39VAFqRgQMLMyW
6cXAXqt5AR/ZeRlS+2LgWtVV7F2PvS3eyHBJCu6n9vHyZVJXJH8lQSFfsoaQUm1IIxiq7IZVOC/I
pxla6+oFos1QjjGcDhLypiL0bn4hwLXIMklFzL0ZjZApAFOvRSJ3jv+Pw3IXEUYPGZ8rfbrE0zxy
djelhaOjhe/xiCF1MG+eeVLjNNtWVSfqoa940zmfva1pXS3R+bEe+9y5UWcPJclzTvg/AD9z4ck5
Af9vHiL1+oNRSTH7P29manf2r9H1FgjowmhZ9lOoJj/PW/s/woEhqx63YAE1L37a90xR/uKb55lq
zaakto+NuIx9DrcGyPDTOGaYYAu/fOKIktsiItiYklTzcM2suc1IEIKOKKnUHTuJMKbUD/GAW54a
Ab4no8ybhFdPbOSM9PoGJhxDggPhMkZvJWxzVQOombiT2EUg4jgKYyBWUp0fEhmqZvhI7KkcCPMh
t1/W8Xi9dQaAGzYA0W5kfHQdgK3cZMEo4KR5AmnzIvy8U59KSQjt3wuJ587UdpDgV3GS7ukxN/KI
PfCZVUR6kApcWjBDqdCgKpVTR7nhCQg3EyS4VRAMs9ek8kcTn/Qz2Vy4T4/Kc/mo5roHSiJzY17h
YPAsGTrXmcCpAebymPCChEjvgxDWN1k57Q8e4KUJMPKhyIXmx7MbCzaA6tH4WqtnikbBnTKU29SS
DIvXINZiyQXXR7Kg2zTJJuBCHu5phak4wcbowIVqlKDJHdpJ2nfE4WfTrxzqNrXX3jOt1/xQ8CdK
wfzXz913rVBrSbLAzz2dmBk1OR/v3lEfvrb5nMcLRkYu62z3AtX/gYjbOQiwN3cEHm5+/niUXqCF
1SYcl6rtYsEPL6et50BwRJxuD7IgZmSkIobkjwGJ7g6nwSq4ZICCgWT+VMGjlTW4MgmPWy1bleBw
8Mkzr9Vdf9rk7/0WftjpnbliUZ4PeLbKH/dorkkL3i1jNWwvor/1flGkP8QARTUukMZLfiqyUE6D
X72/Gbna9zdbmJI1vv95x/iVXzAh0vqjQ209tHFRbeKF0sYHYPeNQaLGCgODwgyTU3AluzU5swDi
yexLlOHZSZQ+ru8/rBRWuZv+MXAiPgi59mFDTfwMHW6Fg2KR9GnUJOkeD0WheMnZHJAbqjoUXmGj
qIu7DKxBOirwpXs2nULEXX/wUodP4hbRT34LVDMPym+x+8QEz2AGuadJLpxxiUBl1hoemUqReehL
VH4KhEUFqSrVWbIGyP1bw3bcSmdjRP+Ssy3bRg3skuzIEm4+9Ec3F2n4mkD37we30vn6X/toK+6x
przesMCHzXjMhZrpE7sjl9uwOxYqlioDO1QYUhIIQ5rgGuTACe2hyrc68xvQB/WO4YbXzF7n82yd
+vjuOhLiTZqNjZyztXGRMuKUUINW5fZgpX5Dl87K+6Zu3NIjxc2j5ENuL/euZUwIQI0Dj7zi9gvN
nq2uiERu+FM3l3ipyFF0REHYVXjfAPr5rq3cPHXQx8y0K+njCtyMQW++GDnHOuEh+cXvsOdiKs0C
r5Xss2MH4R2zOY2HQPIervCrdqHUWqGaYqPpjrRoGcYK+4sbtyMIIQ9FAEpxzwnv36BsGScUiKTZ
BdIy3BFUtSA18DG+5Y9g1IqXIMqrMh72YT26Dk0RngxyD8aPt9ZvTeydS67hFToi8ePm3mRp7QNv
RxEB0Hvq5x8qV5QsVmBGCoQmGUTa1TWcE+EVe6/KokHyM30vCtor+TfAtV7a+mwXV+zN3WJxSvpP
cpUS0cDW/DYammGwdAu+DBrAh+ohsAZ41vbdXg060QyxqZoW6enmcD5JQ0ioAEAMZfwZ1RnuNXRG
OAiOi/1O19DZembQL8P4+K3JNyp8IdLmUmw44ZX56xyaVHP/dFVtVaAKezRo9qlSALf6EAYDXuhS
Vk7hBJoAqlOKkw2uxH3pZwROea1hxCubGDA296+kVFJIPH4xqT5Z6RsP569X6SBhw5LVtTHBiabB
h3rZgHFR7U3NL3GdpoQJ4fb6ZQMFlUd47KomXsImoaUz4cH3OoTyAyXH0FYPSoYlioCC0yrWBjow
2DIkMPfCHRyQwzqvcoHrS/mQy0h4KVEhOTiRC08eFKUDyTvgyUVGgnvJpFBcEjuSZCV9T8/6bqTI
G6JzPfvmjTdO5cJkHVLTX2vHzS9FBN3tIDgdbCLDoEdmtoCpZNYPXr5i+Ps9HlrDZjWJcExh2Afp
r5yCxcUa+zrUDVPE5MotoJ4ViNn/9uKy+eDARxY7ikSrBdh7d8/Zmq5Gfyn80olFWthqw1YsvG0+
C+O0lX/iqSr8gzj5neLh/gZixg16g50sMF3Y5ZWoL5xCq2uURHkTJKTgfcSR7xZcXFFo5PGxVIs6
GM/vSbyvffz4szvUS/xUBgk3o/N9tCFwoysGOQXStHIJRo+lDH7jW12K9cmMFgpll6abbZe7Dy2R
pviCOdaGvTdal1P4Gy3x8+lVe6TDwi/KWHOrsTv4B6DRYDVBWgXnvdTI9JqnW+MNgZZG86QT90fm
jHyIIa7QJRMnJrHbN3TVecTPGto8ln12/c44ly7sxKWUsCyN15FFyvbwDxGFHfQk04ZZoz1rKMxG
FInBb60U8TwPZKKYbX983HtWd+hr4zvJFhRaCJniqhYULjtKmXfCCr6Q833FlJuxax9OJlbgaMYw
gOuITs7QMr++SA0jJdb9+vnPxJXWY0nsixCmTRpLZyDSPM6xck63QO3+CWEIK8m4GKtwZoePrCdZ
ngYE2J02s/2Nb1NyyuDxKLq/1wC76Xn45cG9mwaCG2b7kiNfjOEO6Q3w3LRpSfGsPb54I212LrM8
tQc6SNkBJn/VGszwd3FoGJ4PhP/aWq6m6ZS8nSk2ZIeWlqMIYv98qew/3q8m1/xnrIjZdYZZUcQS
qmEsmLSqEEIPL+kAbqLleOhXQnSnnY6aKqfzvREFXjqrJ1d+ezT2imkuy+tVGVHVjW/dEMiQQnV1
BnvGw/uruM7jRFvz6V0OoWqbtus0Ehm6vApiIrAm5jx6h6+xcZ0BOzfNDVgJkvqW112BYefMeyCy
b/FH/3G9mUdKD8HmMOwiBC2L4Boplkbw63aqD0xgXM/C5AQOEGpPtfvFogKhsw2h6MCGELPxNEGH
m/3Rz597Zv1WNL7edDHuF7GvQJeb8zYck6opR/DgmiZngoU6cNIgSzCa5AoAItkMob7aLct+obqk
PEXPqa7DpKh3e55fMQ1KU4bZUrVOJazGrPXspbEFDiCYaXdBJWeYSyFGH0sRME3W3006iSGY/29p
0f404OrbisvUrwUjcMFwxmPfn38jTUrRw6Iz6pchYHhrRYdw+usymV1F+XkMfTfccR9PSVGk89M6
Kq4uIyclnHulSBSsnhuLkOwt9xyTYq24hwBaZw1KZDi+tPoJ4yGJXTp49sR8MG362pWfrK9oO4C0
rCR9Z0213RC4qd0PAcx7x8w2Cwprr6gVS5mKWT4zKB3vPTlq33mv7nQLmS9M0GFsVQNID8FSwtxb
0tTMZ4RcTsPEXE9u5vH+HOCs7jh6P1CiXd5ZHPH0APYwJrP31ModaDXfHOBrtFa52E5ZzRFuP9cg
tidpHJ2EfrylgTIWtjjhmAnILVkLIoS2qMvvTaFJJI7pdZpmlNv9htAwb761nDch6z5cH6N1Sic4
YNGirjW+H1hI7pjRmbEmeUkcpp+2xVYC1cDlmN/EnRosvSIQ+tNdwtXXZe5aMikBQK+Tl7/YjspT
TLR5F6LS3Rxg4TY4EBXiuwS+bbxcuMUMYgBRGDI0J3ugkpbXKuHPthWMjD/Q5dxcV6bSvv1lsnDA
9ewaTa4ZdIO0sY/dF61ALK22C6BhgxHeUKN3o8OHLu5JpGxImpPeYljYnxQ0mvAH7L011H6RryN/
Z6h7lKMHGcBlnL2H5lSyEmmVIVvR57bRMUZhU9HU1UWKRpbiR2HcXu8tdHG6Vmx9T4ZnJXisCLyB
xxe7EENSBi7KPkubiEqX+Cv9C3oSPrlRM/M11eGZY505rT7RdAcuqpRtvwgGmIu9Bqv1jRJeDpXP
c9S8bhHBoIawWr4ufvJIWlKjN4WdxGrQ97PvCk70LEmDv3OyDLYJruNQyuHj7iTRU5RZTZ1Dyz9t
TrIhP19nUuxeBqk/WKaPaE2BNxu+Npefzc6GEByBSOFBueLoYjlcoHRRR2Oxw3z5hQwLPliG7qxB
9iOW77VCuj+MRDYsJkVijlRlJPDUpbLK/zKNpKh3PscuUtpDA67Aj6EYKVoy8SMI97+OZ84dQDRT
MeLuzldGtTakaihJ1zPsc70NgU88QJr/NyKnlQRQDyWcnEq1saAfAd0IBqbB+8SAJUvsMW+oDNu5
D/n6UG+moy8/VAu7EqxyO5nW9RIl7z09Ez7qU+dJqXuV+b3dZQwjIj0UJWgvrtkA0sZCXmUgxj3j
mu3BAVSsI89FEs0OSx7zw6ERJkH/Eb2isoVo9hheXAv3YW0K6p97XT9Eu/2TI6q90VcHgisCmFaA
qJzT2CGPIBibj1eHkk06QJvbSfjalLY2I1soK5n/uAi9FsBjLvEI2lwhQIJJsyRtl8MWfIJZJM38
EoU7yTE+URZosjAN6QbGe2q0eRmzoXe2lk8vkbT3OpSZeAkl1agjQ9AO3uwOGAr028vyokUBePCP
6sc6/n7Tvaqot56Yd4jtdKBJ/aMWZUY6RVjC+2N0dA09jH8nBUjYMuPa4uB2I6yhzgGXxowr+ZYi
pU0PGQcbUz3OBONOGFAmHGy1F/yc5Vv3E9kmQBetEs5EZzqWVfoUcbzpS/Xb+x8fllrhHTin1yR0
jxF5sL1nwDYrPprt0PyUMpv7rJZVpfHzNGuqyS/6stxQjuLU2n2/iELU4zfgrQneY3AjaKl7DM1K
UfhOnTKCev/U5w9LgwWY/Rr7wA/XExqOj4tXfTsixbtarWPocYMRJP0nNJT2JR8jc0QNULyswmH4
VuRY6+GopCWCY2SpXa04yptK3hVnSHwOOf1QKkI5/SkFadzG6N+9VbzDTu0IBg+IOsIE1bjBVB4H
Y1X7GZyJwwJlhKUxpY6Pe7HZRqZBq0tNaQJD0kOaX0DF7pBCZ5xAzHnbXVRO+slqmyjzUKN85l0L
kqJCIcTlSr6HwMTU3Pd0wgr1YZodaH8gDX2C8ZrXwetjBOPgUvDx7DQ9VhY2IoRw8spCOASD0HQj
3qAQwRL58kNLcenYoMEAgj00MhKKpSa4z771RqtS+42V0gFCOUmE/V9OvUoQ/ASLLFOOrxnJFU0k
pWOKOiHo4utytAijzOGtFh1TBl1TNH7uxfPs4faGB9v0/wb4DyTc/8+G/xyRfHAKkoW9PLJl/h5d
gsimZ++LLeTV+ce4ZqeScs6tzDk9CIBWQhcAfaX3PwBQmHUj87KMEHdOE8RKgN8Rtr+J/tuBgdGm
/UZZRiORcI6rznSk9Bt6GEPfTf8sbvltCP3jR47D4rolICw15pg+qnvIvxXlep8veXXdAX1Q+rot
ukt7X0xpr3kNCTnfjvg7yKrrLVzTbkkb3QaIQ6aszUmEFDVvhlGg0RZoC/D2GdMHHwyh0h2eYTUj
QhGZ+dRN1wG15BsuUAaHJBwYYm91+RbsuoxiSCIeqt5evv9W7BxDiEzf0Z2OOiv5Yj1SQzypws8h
/H2x+I1pj284+Niv+woexxlRoTnhOTFenZmQIJnx8fux8RI10BnwTCBmydSUJklti2vS5I/fRhld
+MoJWHHCin2WEECJ7jQzbR7SokQ+9zsQBaQ25xy7/XUN1kWxt8NPmupYnuT1HyObfZ8pXToKRsA4
Dvs39nk8RriuEBM5io0yYO/EDyDAN8lrGj4VHUOWo4U52SA4fqlMADfKFONAduG80LM9m5jQRbUN
LmXM4gg4xVVg6lc4uMmb2OGzpbx4YuVPjdR7Ojq7mzoFAyTaM2jAohxsiPGXzIhEaXYxLHIZeG7l
aGXzkVk/1h0X5hRDnGpZtnbKJkvOgupzh568FHjQ3lkSk1NQtQLMdr5/YWTlepJSl8nTAGDG/Lgg
f/CmX23X1FHiC1EJjxFrJGpzAZdguacX6gcW5V4UTqPbfpmM3DYBSRB3VGov9sixhCnbTiJ3Qhna
qC0kSL9Dc32Pa2ee3YAOBAmx5iXSEI4auku2c/UlkFTHg2l9VDbiQQwUsiqE/5mVkQqKijSBBvBw
dJtMyyBByvdt0jeayxQz1Ayn7LmS/sNn5jJv5M/3zd5OEyQJOB7VuQNk81xjZDSkx0cqrPHuCbd7
J068jdIDzgkg+hOS8iIyZjWKMS2pLfCSfS+CdlmuZt2RxZ9ARUl9cciLBdof03s24FP+nPUXSXfu
doRk7HuZv/9uAg03uT50ViPLyM8iMkWfdxe+UBPEIxEu6YxCRTdER0siMw80uYppjXuGBbsKFp1q
FAvupkJ8urArLwLm4V8RWSlRcJvtJcx0D4AKr15nH79X55DbuV6NI4uluJ9sLMJAK4k/aJIuFruo
hJZDiKvvxFgFaGEX8S50ftZZq6kYmJK05Bfql9hNo8trlrt7276UT7HqeryZTNzgIiCaXh3s4ZnO
pQY0vZnikisXbfuZ0gsvishU0q/+cBjECwZCuZ92wJhE+CCDhExoe1+XmTYqXARfn6w8mBmJmugs
eUgzeBRZ54W4l4plangqUrVnPww5cZoHw5PTADYP0Ekp6CrpoQP1K0tLMoyrVAhSy1T7gYMxtXby
3fJFMLCy+tGgrOC7AkrA4CfrsOIUGA4vN6sReqvrwABWtSQb3WcIb04pA6mOAgDuImO8E/fabpSo
laXgIGUrFKx/phgo1HMx4jyJQ6rmtjkKUQWXBbHkwrYpuzNpE3s/7WjsqmLJfcqE2Sgn4l4nZ471
gTXu2sEAo6v3kV5GSIVMqI9rqy3XFzry9bvhAUca2PHpeNB3DjV+2GKBjDDmIkfonrBtr0UyOVdH
LZbinQz0TB8sHOXYcIwLFHM5XYn6EBss5xz7xV/G4IYBjCJcK5QyuhB5KUdEI5kr4rQVdx3QYGVg
+OHNfFtIMnaK9T7aR+idS+xFKl/cr3fOf6LPDvcdjKIaFQJqoFyCxXgmt0sbMbegYkA2uRtBra25
SZvdy1wAatCgSEN20tRPGSCJ1Znj/M7M2pVgkBdJyOtOeKAqe4uU4NPLEQO8nAvOaxc0A6h3++iL
AkHArY6+8iGnLD+uN1gjhoKftMoHRL+O9QgqAYJewy9TgO+xYjaXwv+E7O4UYBZ4SVVd1rva7I68
yZBfSXdWXYr4k/wi1fB/zydZT/BUGaUvZ7uExKbBLMRyceQ3XG959G6vbjcJr/sgfkLaftpnRRGw
Wy6r2jhJnMow9JMiTtqW7SxX1Gm8zZS3XZLMNXY3IcVObaa2Pb5ZkQX3XsynH6HLIVjBJrhH5ueR
+wkoL1uV3gqvJ3vzLqtYO4Uu6AXvPeg8nI90qyfPPB711r9YGbPVpT1Swog6Ay7Txj161Qw0KXQE
xXJMWIsJwGPj7NVmOUvkKhYzBarTqnxQ5Za2OpcWbRWC8KlW7n92JqnhxiV4AFtXgtbaHshCiiip
7sTLsxtsnDlaK7f5qzo4X1PQVSv0WB7pHr1Dt/YB9jYq0sOLdfHTkh9d2Iaq2Kgs7CX2XR13Ng2W
5MIbwJzhrbB8ogBvm+E8xJpvCXrBBNTkPdq4/mB3hcm2/XR9eayTUyNLx3gm4fMnU+S+BJv+aAki
etW5auiI8S0TcTdwWldZz1BuBPDVRCyOSfFOVg54eTwC8rX7G8GL3VZqblwN8FGGF7+kfh7RNeNJ
40ZA5XNWavK1uFDHvEzQDlXHl0N2mBLKxJ2aU50Pf2/eSghshbJ12btVR/DxfXdRz0QqEYjyHkYD
jF7sBn1mHH7BFzytjRt14akYqDvH0zbOj14unjINaZDejw0l1w2Y+chqzLuoFpnBEF+gsBWYaUy4
fJvocGWCkCfvXArTjNCgk31Gnmx0xfJ4OQddjSI9NNYIKFUf2+AmyGKwpHhIuF8y8TFC8E92stL4
kKLhLoLnqJugu5uPLUzbTHKzKTC03ogpt4NwSsMveZWdkViCmuf/jdfdm35UZB7U5HNYl6MUnlu/
4UvraeFlMaAhVE4VtKvqV3Te09QDs+ER+aK8iExGd1MsmnGINXez4zxqs9sCYuqNTx9vbqQHUC92
Fyj0JfFYgu5oflEJg41T9+kQCrMnRWZbxoQkFYQPcZTPEyYvkV+6kuPlbuM5QLVpKskYBJ4caqXm
yfPdONX18bwwUaELQChwRU4ioptYLYd9+JnxxLGY4RapKypsWmTyPxglwo7F2t05BzmHIMTXUwgb
fA4BleGNKmP8/K886pbJUvu9UtFlRYdG7Z8S8/3H3G8CPzwlbRt89LTxMhWuhFh9im9c0xZpNSP3
72QL/BKbxzh64bmQknweQ3NaeGlqh2G0NiH/ZaLhp8QTcYRIcUkbPay1E/3QC81da5DByU+slDAW
kMpAgvdJCib0whwoikBXk02gtJqmukwsswNA5b7QHgF1vTdEN6j0YufMIjqhDNteRfWvKOam4UjF
mvVzNm3WlD2ldYukSN6R4p9XCj2LRf98fe2+eP3iC2DQIiGieJIuJbE0nl4fZ3AVA9YN+zY1KR6m
yszTIuAx/Flz36ojF2LheuuW37C1Es/TpVqKXMcYc/h6V+qc/CiU6/bBoLe5GIBFE9mZ1SQLKPqx
N64HaLG2fbnOuqd+oApVNBcXVj6DuTjglFd9QXtD+GFRAcxQTMX+qTsqcAHRYIh8ub4dYej0KY6c
bFizDeP3ngus9zxaZnrqJuGhS3D9d7IHUH3bru91zXB798n3McGWBrLLWaBqkZdgcWXFHJ5C6hH4
4Sz23FlLO709NQo5iYGetqzhkMzStz0xPaLQQgWKwNzHIhJgG6lvYbet/QwHqs/waOUlnyDpObpQ
1fth/yDBdA5eBEerAL5jDvrDUBWCjg0VaeDWoHNr4lBFGrCg5bjAnjOG6b2Br31EbiOLlyMvp2VR
8kkSkf1Xiiy1sS3gk+71gJ7lingeIX/KyPDx/psj9NnkmTcP/R1oHUJddqIvOCRLzJJDX6eMUIt1
vxAhHzdi6hjJ8GUlYP1Zj0SejimFKdXGWANSFIVjorx/JZTfZpltNj/OGpsNCWIqmFOcwmuNldif
AJ+8nkBF3wRsWXJH5qMaGYc7+57YiQZyOdEzL3JLrSXDNTAVL26IpQqPtUGim6PqwbyE4ZZreWsx
0pgyAlKj/OBqHUZqBLKSSFGHggsNv38mCfPKsiGpmRJV49ROAkvnKrUGkO5fB2Qfn6en2RhhHV2s
Uo06XdnOcwc5vZ3uiDLEdJ9A2S+h7jCUvLJRtWjmv9vySxLaTZozCJOLPWOPIQYps9FiRRKAgDt3
WmLpbkn6fcOHbXcJINuk9x8jjr6bmzTahFLvGfokBBhvzcc2wIWOFBQsu5JkmjLsPk/B87/jrA1R
ZBK4YYMCW6v5m3b/62I/93z2+p4XddCVgxoffRGFuwsLroC4hSqLy0rad2ELot1djAUKl4EnMzyX
3IZ5W998xc0mkbhuMJ9gz9J+rd1JS04UCMVho+08pWaw9gm1FUoXPugR2fC9tcX8Bim91v4z5Sgx
0fTHFvfIZq55EL8JaK9DzJA8DOv50pT8esUIN5E4dFa+Vp1IC03mRL+4X+y+ybQjvQIyoXEOzvcQ
VIgcug9V9dI0EqE+nr8c2zrkipQJm0BNO/CJj6sg/jnZHxIqOwYxaHvPj53GdZuC8Et3DItpi/JH
tjycFgi3xHjmyImuYRI5xbuC2P9HPLuLcdQTWLGVYzxpHP1nQfKTGXA+dqT9on7RHLBR8/Htv0DB
bzqZK+yqhsQsi4dVjpzLgY1rdzLEeDh+eor1H+ZDaympGzD7A84qHxWKG+N8HYX/AGFP/zUUi6+9
CUzjQtgNPgwvoiEl4Kc4RwFJSdZ4WbNqK9egbg82YRFW4s5f6VSinRE4jmwZRorNpkaqxdtSsgQ2
n2eWKnyb+9wH9JUXr7G1xPWyGBRu6WzHwj34WK5PQ64QPnAn94viY1Oim/To/gUPu6zD62ns8pxZ
Ys8HeHZ562K4kw+oDRstKgMlsv3VmJKQI8BTMegbxOV9PE7FytdmY7PVFSgx6pVzOZXKEyKsCDx4
7c1C0iAh6EgNZx5ULqzFAVczqSFUAsjHxoM35kQL306pYavIOK0+IQZKtC5ABuWsYakUXdVFfCIv
IG7g7TXD1kjupGGzYCYe0RrjCgDrXB2YjgW61bxvRHXXNxK1HvTzCqbqG2nzgeEomtOXKhzi/uUl
J9LY2TBQ1QAO963u7Jv+07Cha+82waGhLBe7PheHF7XI1QRwvX5kQArikW+alDz3jY2Ik4s4NjfJ
Svta8DgXicaDQNnoeEQ8Q8KWz2PlAgIA6alsx6vm5XXIr4p39B4/OxwqLoXGejdEA1aqcDxcNNZy
mltC0YxydcIPTFye1wMu+laLuW/Ama8D+poJK8uB7uXSgLBYxWOcvKN7Eio0mo6Khp5d0yuDmcat
LDEV+RdApxQA+S/xOwjLrDbOI7Mm+sTyokrghYoDBWVSrqA5gAuMrrxIg3Uut8GN1/d/LI+Uiz1o
ubhAOJw0BrMbG26Lwzb8rKbu+zI30ba7kRXBIEGFK3zKYh7dywe+warctHP2dE7X44O3lO+Xos9k
NjYzRe0iAcSvzSTK1NxCUL+bcQNWS5wlUzboKVyCg5o93hzj5Ewuool3/aEjDcPDo9beRyBcOi2D
b3EH9xPou/Pt/bEdQOp9IAAoQaDB0xEZnOgGm7WZtHqk+XiGTjQYeK0yTuD6KoxNV8Tukbv8SOQe
Ys3YzygwbZbl0xi6FutQ2eTYM2K77nJXKTsl+esyjZLHLT42R6i5cHGAeViHOD8KJ18phc8MMHEz
BZyDWiaIFqf7M8Yai0Pn/LfXBuDYOJ9V3tltCi32Z8B9N5k6McFq40xm3GCo+qarTJXcVPkvom40
pElqb4Qo5hA12WoENOn6T5qSnACIeZQ28zZ4KzsjmGyDIyRLmFvxsjVItJDE1DIkRvMe7YBCyGkp
ssBvJTlItdhqqfMu9AugtU5rxOjBPq3SJmHkeVjdz014AF9iJSoPc7V6kaEWJXhTmwEngApO92Rc
FTOlkgiOmR5phqErHgSIYmQ3hqEqVy9doh0dmq+Ow5iRRJXATbtxx8m5ZDIEvoCyDMmgKobPWVnN
w+z3+bcWTvAnRdEglM6XIttXyg60WnDs4B6jEb7/VdP7QizNdj/hgbAUMfkS30aCNL7MqaMFWYzA
eOGxzk6k2kF+DvCKxGWDz96YciR3u9wGcLTFPqRpWliM2A0qCcBKxd1GCS2UV6iTxZba1+7FP8TC
NZayKMdPzEIuuQMnG7uZMSNrwnQu50ssAOUeU9zLuLz290XXP1VEhVp6+2JJkG/XdynNWjf6yGmf
XD5vALl6XvD8EdbVFOWN3BC/TyuYobx7jn1eDx6SC9pd0CFGqr0yFU3lk3K5Ul3bdPA90Nvasvie
ImNtubkY5EAZpe10fFKY5ojKvQ113mJXlw7Nm8nfT01XsW/MXdUuMrNwWvJPdW1/7WOQpSr+DQgl
ZKc/KqKdnT+mWeu2yywxWFScuoL9cdimidm8+rrv60QR0bnEpw8wyuimP9IiDZYrzdL6HNVCq6YX
h7pg1lBjPd1QDaYk7DvbsU/kqhGHS6oKSPSNXMX/sIkEnVvJ2hCIDYQKAPWyVmK5r8PrrdVcF5Fr
no4wqCphd1Yr+eMPhY9BqocdW6VgBRoTh+QN5A0ep68UTkpc3fEdWZD50d7Plk2CJwdSVQ7QZ/20
oo/f2ufOkAQQ1HM37AeWHJwNcdaOpK2gFWVPTarOrXN8k5bDUrjOoBrblWEPDeisDlJ52wRbW+vy
sNpZNalUnepN2AjbzGpYWgfKJFiKTxlpgas7tVnhM59+AMuRv0ayweYY1+KztE7HAXD3KAQB1fsl
VurkX4F933s93rnJXA3O2+5PgZchaY+osfUa7yX33XWrUoREBeyq5HBh+e+SGCWgnyVJ/nkGD8LM
oFe8mUuuIYUfLVpJXKTG7NWM4eiDMjrGlZ/QEEylTyKT8Ml39rlJji7gsmz6mAC1drrogkRX2ihh
38syb03hsVjU863xNXZef55G/xI3z1C+Q4HHrRKvZCrZum9lLtOQJS+7oLHAbNKI/elN7ibdRRR4
LZ38sWU6vE5EyKw3BgsqpcP8wP1We5a8mbM0XUY+xGS/n+F4XkwGd6bAE7JUFNS3X5P+4jhPM06E
cO8NTMs4rpcLH+Tu7QibLXwFrcfI3Dpby5K+lvaWMuZCjLJp+izJ19ELT08Tcca1d/+aC2g9PDrf
qehmqvhBq4W7eFiCcp/MyOQy4K0B12lXBx5ag6A6FOS6vyUNXhmlrtWRIWtjYKYCP7M6bJVowcAT
Wxdacjx9GZ8l+7a/AVPG0PkqfyXPDFptmVy6FfLARRXzgVulqvpSOnUysNBSQaRhtO6j0oToTwx/
fJFdVkyfi8/fY929xmEZ8k+S/2GBTpaPYskFqn1MLxCYmchyf4P2fVDxbWhI6+JP95MOJ9FSE5bx
omDiBUI93zEhUCLdchKeJQoRUrUwuIlDCkRruvtTXM2elOV0X2KVU+g7g9+SdKhPFTFR4tdp4SMT
FjDn8CVwI08uKfSH8oIAs6GOr8fh8zA/mhdlu18Sluu2K/c3bTPmgKB2GbaZKa4dO/P5sGx0tgj7
iZUlybjMAwu4hi4DOge4M38NvkXMBe+/1nP4qwO541wjc0dSHICPqE8pCtrx0Fs1oiw4jIu8oDy1
phUvku3/85sn1GQFrCnEtGNEbuu14al/fMwpL70EMVWvmohCgA8BNL8IAC+w6XkHdSw2+Qskp9ou
5egO8/+9aLGZNRD51/Gzf3btR5dm1Ao4A+v+REzlqlOVf9ABLSoYA+4CObT3WHY8CwvXBXgXI1+V
4Uruj0GQeCwVxUWjooYWuvISPRCYaMmpYslGsnI3+0S70JSORjVX31dzLn4YDP81RUCuw4Nj0dTP
ZUQXPrse8PQ11OXzFZnTxaHTv8rF19x21KzULBAXMs5Q/T41GENOgcqG3nY7OrmcMkqJFRS16JxR
oYZtPykTQO1M1hlRhCfzUc5bVwOQ9Dx5tO3HyvM37D+qE1kLFx8fz+46KrQ6I6YUN91C9fL3cELc
5bnJGD03iDkYUYWaihTPkeFpr9K2NnIVxTY04vv4MOI//Cn5ZMUVhZgveEfpBEqNw9V2K3FuCOX1
e2UiCEMSIts7/t0bCuVhQ1huc70WO5ma8tppHZAxRlALQCS6vpN+oz5QZoaqcifje7PWqRgWTXlp
9jSQAmLfOqVSMy8t6pA/ydSYEhauvtSvf9HBHo3/c305vvCoEuBwik6yfplfQMqfWyw/fr0lZQqN
qc5DeSMnvPJq381utooKBuS/TWhUaonr+dfJfv47NgIf7QziNyRvvAPkngLfgTGNkUbEiJVqyBYO
sKCSZyIfxKjfobLk+uqgVU4bQ94E2urX7Q4afLROefHN6aB5nlgo62UI/G7obpsd25iQMtj3sNHz
Piv7qiTuCrKTRpicSpQ/JaGHVnzi1KXYuxkqec/DPS/zRm9qYXaLIhdWmo6OrEEjZ7vqkTJuBLRj
aITM+xcFln06NW72W9KknY3XzmhKjO7VimnZOxDVP6pTXtxUgtp1vFKysksaTpqhcYYhSzT52GOk
BEjTHRSCodcxe0lnhJ2OcffnTKMFow3npnVXZnJ3JRHx0lGRpMzB/v1kr1UC/KFQddCAS02ZJC0g
NP8Tio3nAgFPxY7rMvDPo+8ND4H0oe5hV7yzr9ZAFVKF4sG3cqI6gN7vSAU+oJx92SlfwvL492/y
xshB+q5KapWjVvx5YOeVvs0fu/1O4+uaFIKRLmyE+rDR30GOD9xeGJdkt/EgTbC+sA4bK8k6ZvzR
60WrEWNVH9ocWt58VgfGJ+gBZVP7krgKbbUmMGa5edhDrYWN+rObaWnuyx4MHOzxgizDw/WqRWKT
VPfOvkfo92UD4r4UsPZW0rz957HM7XHXLWc3YimRFh9mEGb/HGd0+t+JMoaEUNYPR0e7YbfC8v61
kyKUKqdjNMX6OhxTG6EAC1ifGPW0IxC/8S9yf12UEOGRGwgbpwCiB2UqwIwfOMpKgAT5dHTjc3MJ
YcqI4+1nDR3J7Gom82pZMuvP/qN97jPCMOXuiTl4bG11S0Jq9QxT1trqifFcgSZWRqQ5OaPSgbs9
iUuv/X7PfhBjNCrpxXvr7Rd70yTaURV0aed+lPbXr2EqvK5+UcHMlJBGbA62trYcSvl8Lu/2VpGd
msN8r92W8Sw2bRri5ASuUeMkhDObT0sPOAAoUv9ciE2AKUTiKWacb+hO5lm+PWJ3cCW8TaHG6yvE
8CVle1ZZo6auaX7AkI9a9oa7n8pA6H0Yy7zmCLhUuBWm0ESX7AsVC5CMLTaJFvehZtoR1DrhZgHS
M15hruhVG6VlUEV1PJTSX6w+DXoQyEwC/nfE3mQvh94KYO4AnxVxe3f+9hwDeNVjMM/dEUzhXLwK
tLxt6ijVCkR8+Wi0U1TO17Ocv8LaYpZqOMSsx+2/5SOmhSJAVak+SsYt/4bdiuZxpusftZA8aObj
HFFgin+ypbeTktwP/6g1B72KhUkUXuCKeUaHiFBO0C+gVMVPIMImQWw1GDfesdaByaNze77dHFJ0
KyE7i26wBtU+8nucGHiGRznMKv3d9Gj7U8q2canSDSgClrnY452Q5dzVOqcuU8X0OvLAzoH8mgz5
Sj0l/4SjKrX/OcRwVV0M43Ze48bV/JqhzIMsS7CTN7vIV9G05KARZJFxOP2yobX1b+5PIbtE3m6g
jbZl6rJ+j1IviOiVk4AAUHXrYA2dwAzpaNqHs2GzYn1oM2ShROwxM3ed9yXB4iUVgI3h2k2xOhzO
vhTXmaIUEiG9kTaWMWt47lQD0EF75F7/+8pW6mbdsIwuNOByet9D3hS1qvckoJsIkWrvhGZ2NcTN
Fv7l/s+KAtSE31AbEHmUtnS79lhNqZp29n31jAfmhMQsizShfLeJXiqQPZFYmblvkiVSnqnhcRbt
hJd4JTJH8wBbXJnePvD7gG6+KpeNdoWVWa2K7rnh4HQzPAogutK2HBKi+T7kmIcAnaWmtIiwwwi0
2nEAZeWZi45eflz+RFX+YO8krlAKpifu7UBzScPm6q2+lukUPEfw0vIcsNwcWsA+d4ZNpWwSPjAg
CRNn762BvXmwkwtHDjvaBca9+44hLKlNARPZpKmXjjqihLuYVnIGB69U6cu5RY6dScwIL6fxiV+E
Nzh7XCMaIaK0Mi0639P8CUAi/4+TTfNQ0mNmT50IG2VQAso8Nq0ZroK2RaX7oHp7AHqIihRwG5Nw
JwIgNCNDGMA/YiY3hW578kIKxjpqWWgan4ngX+4QQmaTGk8fRiNpDV2kj+wIwrhr8gg6xi79WZgl
Qz+ScysJz67iO4hCa0ruXzS9yO2hy0cKELGArs3Psz/3m5nP1eVbL01/E4JxnTZY4aMMW2PdEmF/
1bUX1CWv5NrydI2zTodzXbR5Z4WIXdYc3755ZYDBpC/DC7qubTLSPYe6dDtPEOnkN8vUJoZStu/o
/luyrXro6g8+nVHFzYv/JsG+1Oag79MBIAgWqdy6opu0KZLk0tBjOXTLN4XNFm/dY0rixvITz+23
JvOxAqD48ivEbvAGMmCuSabmfzy5caqKzeRMtrWYeIa/GWP+4hrgBHkM1rjQXSaUU2QEc5l7GEez
bJJLAKmPfEyL+bQXL7x/cAW+lw28c7BFsvBcT1hOyk2OEyCL/SmnVDzNn8DFA9ztet0Byjhg1pnC
TETN0pgqCpdVDSQwi0ztDkrx2wbcAhzrcQvwt4+4UctBkGlrxfjQfGIkewosxFdzjAT4SHOtF1Yf
aXTawXkjLJzW8Ha2GlvPpVFlqjlQ208dRv3ZzQQ9jwmEK7SMvuYf+CL+WenkS577SZ2ZIvateIvn
F2xkAko1+9DYuOv39N6s5eIjpQm0wLoM58fb1hjbvCV2VElj88qxO9sDq69RYkYD533asDX+pcXx
y5GX5wZDIh/xwVpRr8JAnaAmfAl10oLajK1+xaSXq/KlN8AXtbuK823yoNUA36xNPXfUelKGy5Nl
XI2FMGrTJtRiZveM7VYujSQ02w3XhJo39t97f4U2QRUCwKjDUE/buU0pp7yUhq0KqWQUeRH+s4Ls
IS5DbCbmqFk+aAbhqiFxCw9iPdjcUs1ebEtHt5iHDaCWTp+RBpQ3otvC8aK0VyEgmnPSS7G8+yIU
OQi4Ue8mU2n8kVFNj2XzVLY/u9YvCKIFB8bh4uvRJrkfhAgiILPVbUW6vcUVaWlitD0podC0dGqo
kD0h0YQAtH1ieKoQZi2AgvA8/NZm1tdX0j64S2Ac/UuT8foPYiW0WX3ySA/twe2qa+Ospk3bZUDC
pEAOvpDPICcqniEg1kL+aA/TtEfPjevDLll79ReZO0o6Uy2oJkpjCZEkQtsomL/DnE2DazeG9Hdt
PdDAVKib0mF3pzhafjzTGgOU8glBoL0PIORN0+wC5/BCfleixBvMJ/bNgQl5Asnq4jgdAgLGTrrP
wJsvXU5kka+u6yfWs/VkJeKs3PZ6VrGNsiv1i9Lol1/fWNSFVJjvtp36E41VH/eEP12eomO7xgd3
rlGR21gpA5Jfsh43MSmb4hm8nul/VRnXY4nABLK+nb2U05Eut3jfAS6TIIQ/FWTXCK9Uqr8qirgu
Nge96iFcushlUxYDsuFHvJwJ2s8h0QgavyLbzssUbNHiVvohGB1vSB2ihV3TaPzoXrQmwzGXtb4X
5BiNgPrLfXz7GkztvNXRXY/ZH+fMbQ/L4yfrTkHj35Ax2w9c4ZVN1r64ehOxSaRN24Hex1PM4l3L
yP4HpYO0WT8qBSNmti/cwcOLfsELokGAWZXEHyaJ7y5RR/+RmPD+TMuwX8HnmP6XXQfhEfh95c6N
UHry6FWmHsig/I27HO66Dw2cxqdl/IsqJ2YUo/XNDjiX53iIm0lWKID2dfptO6f+yU/bCVx5Qp6p
Hoja4ZPPPJO4T6kd1nMwVRg+N396K4yjC8Zgz7o2DCX0CAGHAk1YG2ls6UA1pxLs5VR1CfoxdCEj
pK1Wrs52XxUtk7DXLoAAGL9BzE4Euo4fQyju3Q2RI5OvXJ7/Lj1FCD3TVO0NDCVgSHrUUocRfJNG
TnmzplaYfdrzy5m0dlzqwJMNCkTT0PVph9F19uqn1CWngsHx4vmhLV4VPTCNGFVQbhF6Aai4JqmU
jGgLpGWRhLPKZHkg68rE3MQrFo0x00i74y61VH14NtUjCuvYJtRomeOH1ApJyQXASwV8t+G15eMJ
707VIfYDA1rB1N//c9dB5n545m2hAYg0n91q5ECRIZYGVBOW4sBoLTyUQXlgZRGJNnfEnJk5D1q3
15G0IhoA6ztwV+yAL7mA2kuCstRoYPanker1geSryfFTVZbo0ReRDojyYJsbkRNj+sMAYM9NWwnn
6hXCb/Ivf0zt8KAQmYDite2dj2zZKnC9L7B35/iVVUilD9am+ynjDm4F1SbodhWzYE3LKOVsSxxt
k0V1mqnGZ0S38RC+AEypeo6WdOSnYriJtRDqCis4ZLXuBpPxYJu85IzxqWRZG/2mMAcboJAfNCeK
+q4iEayOglw1Eglg5gOqj1RnL5R4a9sTVoLA0wC+LBTJv4gXevtAowRdggxQ0NXNsGg/9hkpsUi8
nNz11UPWDsNCJvSaVW7wEthzO0ITjZ2lJg0ZYceUncUebi9QlXirnqYQcvdd7/FMSE6i5T8kOSPC
VwPqGOUxEdg1niRpK4B8kC1vBcsSa+nbYrOsL4loqUzZxTstSg1R2V2viLkDJHRbZAt9QXkiwYIM
ViGa6tWE1tBI720BkXNelt/pm0TgFu+WD6cRVPFt9fz43ToqVh02Vdu3f5xqbCtXPFoNmeM8VaPC
u69d80c+WVWApidaVOj5k9Wxv/LaQQyQd6TA+Uu+ajsL2xtp8NdG9Xmko+t+lYL4Slblv20SOC02
l55pct8bTGhk76hQvQYwZcG9p/hfwavrL5xmLXXkJe4ZHxy+UwCdnXc84+72z6kH3QBOkdnHRTbL
WdNP6ng/g9z3yPp/LMVot+CKNh5N6HLSK7c8ig6CYZxas1Tp3OWgr3ZTrPQGKnrePxL9i+lATcch
hYgcGw/YuLdYMpihVcUzfkAQwF5Cu0OCXAHGI6bCFJBzsOARbAlk7kdhpmQuIMYywcR3yJqIJIS7
nmonWCR261kd6LDtCC7zsJ71J9PG7uV4UTl5y82G9mDhKvsOHXel2d07mA0SK3ntYzfEDvfIE3b2
WuQ21bi9tZpo8u8e+ZSdknT5s3qE6aICVS+LOvAwiDCzI9R7wFI0TC0UvPZ6W/2IcYyQ+6lOd5th
YB7POQeRNKlvbJqE9QFckF+05ZwhI1WLpBxKXXUlNv5tZzupx9S3qFcgrUTjgZ0xy+27X7kSeaa8
gLVdKWem0JB7iSKt1ZvB1tpkbh4hM4qA8Mupg7QOxD3wm1v5Pg6FQa+bRieoOe6ktS0LcK76Doke
ptU/BiLNElOv9+PI4sqzrL///kALq93KvOhhjhXu6QxqEhytYUDL251+nk1K4LkwDr+SWt3ZZ/9E
CHWNEz7LXd5jRfAAWswdXXMdW4REh9uWGnPW7l8l5F9p7UAbG4DvQJl39N/ydsMldVHbP5dCIYQu
2roXBJgaOXeg7MaAOH96xMhJ2Rhj+dCqwjET8GXPk2+zdkcvs2pO5RrfwFtME9hbbtoqBXnVAN16
iWWV0gCPOtfauG5wmUo3fJdBAduhMzu3QlEyGQsykvBZzdAFYhRhZWlSkB1PvekBHK04B7SphBy8
bg2sUwKDOsBrsMKgvJFV4HA3u316BdaVMEHaZzUZzTg9cQp0Dm/zKo5UIwxZX/qHiYhdi3slt5xJ
JcZYN1HXIuN21TAy+HC3c0Mt8h4Ppbmixlvdz2cv6cI/e1YdplzvCcO4yP54kFgBUUb7GXPwIux3
CAGVrutLSUbNy4CcC5HeAH34Mpmax1bwuSpP+QeUvrdBl+l0LiBZPUuGmo6J9x3aaLJWcbphYSaT
dQUrcW6vuMXItkyoH5NGTUeM3JeJQHUEuY8oOY6Y/6m67AsTZIlpFefMcM3oYAZBe/7hZbhkcq8Y
9g4SPDl4+ABhF9AWRcCeFYVKkm9+9vnzLQipGk0CgUd/dJ6D8RCNkHvFY6TyXIe78P4M/Rzyzsv6
seNur37Rhw0l+9g+PaM4Q7nm9fP73YN5L4BDr0bafQmfXGGLxiNCdcy/V225O7n/JcuhX6wR6sXp
1XfjmEKNwtKxyL5GtI/PECDKa536f3cCNPnFsVCXqvX6ywkrsGKgJuhvL77YiL2zHrLlgRCGLEpw
1tgldOsNMt2LqIiOXkjfFFxLRL9uYG8Nrvnd7869nNxtIxj9dDra76FMxUB6k9InoQ/6nTH/vA/c
S1q8tL4+i21iXRvdQRpknw72jv2fubKyNkNa6/BnsnUWmequjH+MqTx+Pdnb7MhsBWzFeR53itvm
UqZx53wWAGOrcd5wkN2lOf48wKL6cZYPJsVsW2SLw01M0J7UXmtm66Wjhg48V17iv5frACaMJwnf
0cREJzNiG8l/qfq4J2KvEjvyPubY6Bv/yDTQKLhD+xqN85a7FJYOta7lvU6wLRyPxc9h2JfDR+/c
8MmOa/nFf8j6U4BnhoSOPsokNOQJ3YjcqJqTWK2dy2FLGKAP9Qg+g172Jvm6JhpJvIyJBtnIhO4P
KapXvcqPJdni2BY4i63zwZWKVPi0O6Jn6O4d438fr2KGr1xfjngcoO7FgKzk3U9B1p+wUyiAx2Xc
8k1ciywAK1Kj2wswq+28lMyzv6TFE536kGKbeAagZPkT4vCtShDlX0uPRjvD6Sry8zF1Fmc18zTE
Z2k4DQzVE+1shukRblBeUjYIXCRQ2ke50Gl3bTPdJrqn7FVpkVvUoIaO7Sem7QUt+nnkKI0px+b2
h9FMEHFQzwmbxKrTHJ2THcmbWp4UvSZ4z9ow5LVmAvhJhlwiMRTTE4e/YYrZPm3wMsxptdkug3Ax
sMykdhyOt0h/A50zVIMU6XsoIYnbzBEyTegBnYWlRcVYSJ6wRn/ofRjdm0OVlLvzignp4P3pqgeP
FLhl8NTDweycROjexjsUsjHRBJlA5X3KQ38K8rWJJWJPjvb0MWoYALUe6hCprrBPnJRUSTF5ddkv
sChXaT8I3pqBTzmnP5E+FWeHy1glMVURA8kCNN7KJWbzKg/Mm2zUMO3ffAZvpMcZOpNOr9j6QHJX
9gFUFjON9L5dquRo8jwwNPO56J9aSFZXyamhGBzq929KcRUiwRX6iNR877gDK/aEuYtCS2s8Yow7
y+mHHnL9VQ2IhTDWgQSfvfKa3fWNj8Sky6B44YkhP0ZyAz7aEglCthw8/IN/+DQ09Z9k7CSjbyV7
ntr/6JpIE44VB/6T1rkXqBJq3eOZOTR2UmnRWsYoE9/gSHGRymiPhxaMvMWkmMtRhpuyF6ILEv35
EzPkX3RoyV2v+J6M+8LAZP0DWkCqvG4uUNTTMEP1kT191QMqZviLpwUf/oanOjGlBH0zPdtcQQ4o
QXrmHfrGmzqB5CRpBF3Xz0gdXu0aC7uT5RQvD8EX6aAPEaBRpjfaToWqtaC5HBavnvsfSPmf49Fb
FtM7D139j//0zdfejYqPlfFfhPW0f55/CWtV5BRhZtpqwG0rpjDMWt4v5PfH5THYDtl8pbCJDKwk
MGvkkfjdWMEdaUqLR570CyaDlmxuAvYIDim5+eP6mvpjETIAUwjE8q5ZgBnEL+/aaMSAycSDWFYw
JPu5p1zbxHbIn+uTtLN4g+uj0/aWJpszhhiI2XBb+jVJQEVooJ701jHcO2WZIRA5rGXf5JHQvDTw
U79AujCot3wpyVWo5msTH0npG3bLCwbvKQmHenwocBqi5deEvx9mMLXZ1BdJirw6iOzjGXreFrCW
cRgywYwu6kmM3HIWFTBAxak/HEvpLW8JbJPu22hXj8MbMc+0khcXBidTYCtxaWu/wEiHPmLY+SW5
apCNCHm+WKEANo5hLLr2G6Whcuf7LKi7jWnXOl4RidwhLxrnawxfL1ikL+hd8hyr0l8theFxmUPS
9/4DDt3jo/QWg1XP+crSGRU58QQu+VvkBqeT2byAENDkCWpu51ZYKbi/02gms+O/Zkwrfrn2YOVv
gcyMrawvrq5Dvy0u/vbwny5vuZqlUByyUwKxT7wxKwnrGlcZGNaS5CMfcj+Nsf7QzDIDv8cJUnY2
OZuFOME4OLY5gsp2j7ICn7l9EDgZ5DdfwNkJRR0wvz6VL8Dbd5jfKdgp4L83l4kJ97A3rDhc0zOv
Oknx33cB27ydLWZOoHwSt7bP8XR082RHmpTsvZ8F6IzFCmP7KuehU4TzOEjxJ73d5y+n46fHmkoH
zpMwXmfd2n2OVy/GR8RCwBu9W8gl1ZmYAvOnGKVYXqT08/Vr3P5VZBM//YkdauYRrMHQVo6sDfVX
JHRP1R3lHBrBYNOhZf9KtQJAeokVjU76U4vQ5gSFAo2qEWsWWDbO8A1ZGg6gogrwCMhTm9QFBffv
f4Zx7ItiOkc2RARnOExWxcPAe/aLLSWpZLSxiX+4JPw6NjBzpi6RCmt175MUUj8lQND4q1dB4AT6
iPMe3rViaCBelwDeK1Ny77s4d4ZjwUUnrS1NGCBwcRHNWbFpkWtzUZ3/G33vBLLP/slAMFt3kab/
dzvTY01AyFEU3u9+FNcumcd7LRlIeMmsO0p2VVKmVTSD3xzn0qswrvnPLQAwKzc1anZpGQHMlLI+
q8iQffPW08nkXrHpWSUQisONKbmQ525fm95N0As7lnn6Dz+MPavxQZ4FEs3xmMcJ4qYHeHE+wC9b
64kzMfeC617gDixid0j4FkG3VCKGLCBNKb638GENm3A41jmxGP74Lkhy2mhnK7neFMRyADZ8jga7
JUpzxuaKXt0pa8tjWO/LfpuKXQVYzF5ohUwry2+46GQJs/OGSey+GyHoqd3WGHLTNVGGRtQQSAx/
Zw60+ww/l+82jBoNr9DXwuOS1vbsXpXCxF3n3qDDkbi2fIHagpBqDSDYBL1WriZ4AStWp1JqwKUa
wWZzFsyOkxDP309I/R7S3Dir5Mtw9cHpej8WRIdpq9vdTO4ExbFVIs6PdLjgfKKfqqwwuTYZtWe+
WO4eyHiIzwn5GN16A8jIBgD1ledLjCTvGpGiSv4VHkzevKvziarscsFv0B3v2Mu9MwMz2tJf7v/M
Zm+1YzNt0B1aXViJo9wLzoEX9x+zzYRDbJoRrQIWT4o1X7XZqHdWoQZqb7/+0BUiaVvn94WkXuNg
DxY6wT5eheCGAtup3W/iI6jZejyCrf/1dWUzpRLGEIOgo+jeadJYbyGeJVEWNVAU3DvRjxhYEfPn
FK3jtf5I5274f3AxA2/JmunnN1JPHmPkIUAyT6xdP+kDnL3SAV7HEyq94LdX0DvVTF868yJtXQC8
eUry1JJ/DZ9h3CSCc1mWfKObB5kxrTAqbXLk5ZcGr0sw5Q+oRSoY/E5hEbEyazluNYNBN0C/70MG
v/u+g9MfwAlEU1bHgu7R1DCAeTgfuVcS5eWkeImDirHrKyiEXsx0Litay8NPCPWc5BanYmhGnBK4
50AjOte6rCOHr42WCKC3CaCc+6o03nKcePHkPATGESQ6Rw7+q9k3rkvnZVdzAYpsLd4fFx/Xow3W
smfQewJ1OFm32oxYQpYuqPiKr0Epb/6VH8OTXDgLb7TLPc1FLK6HWJpfBXwny6psedzE3awalXE+
o5l08LaaFdsEEHfQEBELn9hV+n0ngbuvwzYE95EZp1ElYdxC8mQbHDQTelWEOauFRMyxGC2ptBNi
DVZmyMTApK2b3fT1DXmrvB0N6BuGImhQVokGdAI4es4BzE7Bto9p2gFqKyaZHag3V33NqW+tQ7SL
t33A6AQovAJVDG+QEHTaPFCFZdSyMyKNekrDoT3YeFltnrFu0zjq44Q46yFJd9TKmLKiS1s6YISZ
n/KukHKn0g5Xsha6GPl4T+agdVqbm/kM9r+utNk2me/j8fyJFH1UjlY99xEKpZcArfpYlI1/bQN3
6bxC6ogR9zU5WEHwfeJVNuJ6jPDekETgduh0LCZ894bM9wcT9Rei5jiYnuNBD4zqlh16Yo3/v3Iq
rI0zJlsSjw1NWAT1xCAxu+sX2CSv822NcmO62zNZWc3sswEnRL7EvRF1Jn+sODmKNMN9Wxn6JWHE
2JwnIXDhs/09qU8emsHJVikQDUO7hfStR64etHKCWKe0JqkkDRnSjeEGwulmCUhfwzU8kB09oYWX
46kZjwWlseRnGgpiccO9sCSs9cAmzkXe9JFdG5keBjTE/puC8bJhndGMRL1cII4mwX1xzLNz8Oax
9auVYq1HEi6d6iF6lHq9twEHDGBweC7dIFTGk2f49mMjJfu9REAWBUZsO73cbe5IXDP+lHH3AQw4
Rs9m/sbAZwd/bpRoY4f9rBeRKhQ4XSCBy7lxXgaePWlAArROw6iGoNXgwzagWLHi+KVfLu9KR3HY
a8fXpW2uFzDEuRRQro+AsBGp9R6yUWBVV/yX5NI0TySgSRUm+WUQIoZqF9/4ekvscnRPgAzpClgE
fqZXcJCaOnQc4+sVXa+uLb4zQW5AO1T3OaKVCG66RybsQcTeXEMEZR9shCj3hehVQtTygjLCOVAf
I3HnzbdBWOHRcYiVct+ohfuW0KfW0DJ50g6S3T38f7+Jav0ybeHY3uqyRyoGONG395+6udgCrxiY
x47/8nvE4+iAujvHnGm/qAuVuQ85tMWL1Ho9f1PyGNw54afLBz++ycmVucSRJEkCRnQqmeadpSIo
qMCe/jf/6b1q/0n9DtMW/2YWTxo4zKMnipP671EQo2tmnfMuCzQq/WVmGBf+H21EuXhQQDnrr9Dt
kxW+TOQHkd8NTd1ntvH7a/ApK/+sg9yaq2otZTE6ZMJSPRUtThaSPzbEN40VoCsJA/tUrsLW0BTU
iNe5dxcUMrX2rJvQUiguMdqBEXIiDlBEPk7iMMxN+6SymCCSdYeq4kkxD0G72Jb/eX4YKcVsj6B9
NJRXvU2AUS9Qqp/EecMflvyY5+qKZfxbN40KU1LGoMkBm0+VDpcEQtBmHT1+nG+sEwOhCZhEBViB
BTwa2KFKphf9YChGi4dfW3BTUmfxOwqZFe8Pb5gOp73lKmiODk0eDgsf5ckDnKYSBlf+v7M7/stZ
Tbm1nZBQQWZVk3jsdIDXrrMHyJHIAmZ4b4R6BUVJewQ8R6RTr+fnORYeK5OmQXHN3OhE3i9R/rJw
wKgNNWS55jC0OmSR6TYbfN7Fr+mx2pvUjviHhYP0+Bzn9pYKDwuFFeEE/Tdy7A4cX75rtqZhTptK
Z8a6qYwuc9QTR7422ZgRXKObClSPP9Nb+RB8UxCayco33lu6k89gtuUAzRILkr0hvNHKopAuCQfW
qiaQwDWmfntenfjRuNU27cFJIYRbxpa/cpXrUggVmibl4zI0shTqSytlNG/f+Izc7PyeRmMrd3Cd
Jx/Yb2Vuo1eygo3dbzyfk8saITmN+Y7+rr89Hu96FhM0b0qmBB77K/EzXqNcI3970u8SQf9qvIIl
gZP41sKrxDPNUJozwnl8MyzUv4vuieakld6s9swWHRjmahNh+MJMhOtfBnsbpCf0PJ+QLE0yh1W3
seMYZka2fC1d9ZaP2TiJU68SRNNJiX/cnFfToZw2zBTIQKK3A5dGOWRq5Q1rFGLoIn7imMwNf+Pq
jNsMusAxAVMJiq5m47PbjqfTo0algZsnW01Z8Xb+Cj7bZEx8u3AaBVg+8sqHM6zczqc5moz4SpQc
5LGCOmzROJC/dHS1/TGu21XfstHjedimATtGSljqAMqSY/tdgqb5XbmWgZ2ajtMpx+QjR9AYc6Wp
NONgAR2o9GSu77GZwqAfMy7HOKOyot4yaZ8j1SfvefGN2qlC+TylWq0MpupyWfwOCjhdwBN+uJOs
Xxp5tlI+Nggd8SMWFU9zzZ6p+OMy4C9HsbsF+Vlib191vNany5FsbJtFYZHkQU2fTUlyoo05AikQ
FB2lxanA29NHOWnmnDPEFpF0V2kgL6Hsa/kayFoHcjsj5zzzPvjikWI+Zqy705pcE6mkOWqvqjx8
/LT4O+62bbREAF04XcJwdYMXeX3pZsO0W1V30/5ms+YI6/X68MkLeUkD/fYRk4TeNqMsuLdPwpbx
VSeWBusNkcsG5iHCO8kWq2CPvsEnj6EstND6pFr9S0UMjq5FJjvoAQh6rW1txPq1aH7iPscQWu0a
R9dvD/9Nb7V3+oCo1Nxz5LHODja+gB1TKGaY3rGNBQcWbEO2sKQe7wCv6L0EBEp8jvfdEvqjxprU
zhplAiFwpvy61uLJO3CYzNrA05mvK0gU/jF80J4I4mZtSPXL2lMxoyN7uMAZNWD2vdR5bqZ+zG9S
6HO3wxIlP1Js0fGbKZOsd+Oq1GZ6zbM8akglia++PCm/DrzUrX516tNK9GutFTSTqFT2JqrSkg4s
mlFeewxq77RAhyjTRB2NsYc3YfUsijALP/MlV10f4mwSP8cDfYHTKFjdmZ2mw7+eibIQWKOWhuxN
5x0SjKD9ORXwTXyFmmTxKh3IaGO7tuQ8mWRkF6x+FejAZj/cgEB071cbnOfSDAqlbjyXI0LRqlDG
e1kUAIh+guRaO9E6XHK0jpRxbWzBsD52RrTJh/DpqWycR1zWYERrS6zA4TqAyeVYDVHfL9FkUSHp
p6tCHaCfQ4X/qlrir+yrL4+l0rChMo5ywfECpY/YkrJdJzkwUet8a5tXYWTTjWjF1OXOiNzrAK4s
p+UuMhwO1zvgYKeoU6ilbTilTtCCUw7efLN7W6owB2xMo5UwxYsgLX87DEAlfXqI/K0IZSMkqD53
Ms/uFLoUsLZCb/MTWK3qut8Z9vViCTYIJRMeHqYCHskdauy6lPtuN1Anehe7s0sEtGbaSql4Jkpi
NHw3RMx6vsVD1nopk7RbHvZfAtAhe2aP5Y04SGcWjEjMk/rwG3Vi00Fop3yEy6ZNbiSCDZ3Qsas9
mjGmzQUw5lMTo9TKjHWjrYnBXOi4XC0htJVEdaWJF/S+9q/13j23i27HY/B03V1C1qPJSfdWFGEw
sn+GmKYwJQjt6dViEtXo+Ay3aCnPTn38dT8SLSIG+12PmGyG9YWL01itT2fbvEieipekKgMvItTB
QK879eBV/Pdfpoz/xVPD8ipl9BYBWM15q9IINz+1CGtTVfZGKMbgOERst8srxoG5eUtlFhOBcYpN
WCulBHYVEeXnOOOPlks60hkfhfMNFKFrHwUZLsn9FLq6Yo0rbtb16AKqQ2eCwNQ7mZmjZK1dVErO
7vMAE8XQlRkk5sdphSDXinREH8KIDA/ErIoISpP+bnU+4SQB/RcsWOTaNIj61SS5pFdOHmUk7Aaq
ScGWWmsidpJGgVXDljT1eTNYioqFAfAvUFkacYDoxqNOCbqA6UJvh/iqGBpNroSj4pf0GQl/cr1J
V/upA9mhxO3D68QxZ+mQwycnOeygAwpoV9n2cEBOQLyNa8By5nVbqXsvdFIVS9BKj/3WxbuaT2Rk
PgRr8M4fPJK0z+LX/9hRbV4Y2T9hdenrqpLEovDTzbQRPLs5KgXGx949ElUskKy1AXK9aAqCW5Bt
CpnZYxBiBTxe5K4oQFGduMya7bRCGfx9X4b/gu/+bmEUV23pGp8edvsPO1qGc9uDpUVsNpF+Baik
BjLrr5UGZBCGLAAAHNk+b3DDLvupP3CpvFgyyFbpLzDOhMaZ0gNSUgngZyFIy1Js3T1ABimZ1X9x
JzojhaDiI2XV2ZwekWBFsY3VwIKOdhhVJFPxKBWal7YEIWmaYbhQy/JsWaDlX4cG/cPF/OPWf3uO
/JRdeSxXld5G38YNpS3wpBTvIdDuAuIie8OGRUfJPe5QkJdtSe9aVmd2sVozQExSuojj3puR/mzN
OJbmZvlI16gtgjxVvnBGWAFZ0NnGrxPpPksklprRjsSO2mAkMku9YACkKz1ofhYdL+a2sh178wFx
MlYcYILVyPVvjFS1ikG7UTrfErYrAYbT6EhVCLK6tUxf6IxDCOsr6ppMONfySdYk39Zdm/iQXsy+
GVYcaYtKQyYTfVwQohvxYmzMIxFW0+QYHNlYF3NvMPvU7ihlLs2nF5ruiDRXC9uFmG1HCp0VnuAs
hxVBY6Ksets6W9wslOc5gg4dPFVPKau4X+yQeyoTG4QApqxwNQx5C00wzc5FvY9L7E9KeQyV+rEx
v3pWj1VT+yNcnMn+Ej1yvr+/U1qm2SMFTIzvxjnYnSwAQSbVGKvpCWiQLfkzeE8yM3KrUy2PRGb9
3wmIv1de5NTOzOCy4YMb8PDGXzZQcQ4NQQnNW16Hqa9fsjuj8wpKziedbDJmMx5aM7xI/WkoNKTL
O9NEilNSSQ3ZR9moBOLzDNiwaxlpJzgbc0U8G9s2cFVhyVvzB0A6xIaNtC2OPOWVxQ8LXQdAvWiu
vpwc/JxI2EUbCD2yQzrL/Exedpqww1bBwxs2wakffA5tlmy0U2LiJYlb0Dkc8szTUlmaqA5BZW0v
OHDepNRHibgIobmkt01ipIUfDethcajRDw47xLgW+MDFZZqLZSzB8JXu9DqK98d9GXfZbEoX5jsN
QEr3k+xHi9Tm6F5AcsQ+5TC1aAGehAtSQKuE3GWHU5FrRLFTxaHGnfFrjctNZaFtT/UY4PW676ei
mTHAGTOXUwarHPZmkGsQx+vm578nHTXfPS+Fd0Eu1qxX0K1ITuWnJ92+AWmwCQseR91Mn4Fh/zui
TqSo5eCYl6C1FzSkQtrnGOA6vx6P+jIEiYvkVy6qHunplxmsXjdHGKmc6YxJsb9BzwpiJ5RCEkGF
JGEtclv4V6xAeFDqUtStlSyMrfmBzPBYDqlrrViqBZxPPXxWNabWOLpRSSzRvLX+ZvcFgDi93olT
e5BQ/DaRSl8N5XZNTeMGjhVC6du3jIX4llwd3klt4H6MVl/fd+pJhvW6B/NSCMCwsO+nTYSbUqU5
gISF52kA+5BseuNv6uHSAXuSSVEF6mTkNw+J5fL0TMbyggVIuK0fjG1cFw/eTjQx0OcgiN69dWWS
YtavgxGhBHtlxoV8YHxEHyB0NvSlRyRreWmw3Os8adI71V8+eCMvSM9Gtu7LvMoA+gtUbgCyXsst
2hvyEZJk/d9NBeKFRNE54K+iTrSndKTlnY7I8eVHIEBtx7VLiGd4P7MuO7t4dtiAEU67JhNEYMda
HPAOVwSxGHLaAMFrbmiYkBkZPf/Wjo51QVBoQu4siVUXqouERfncgVZPW1Hgk+P0tauOI+ZQnwUq
tR7vS2ATJ4YvPVttTR+ZHAXmmMnNXl6OObEcUl163aS0g7rwP1Wm/oeYp6Ai7gtJ0sbw1fn2+qBH
PX5kLrgCzpQqOX7a7TifTedvNsCd+7PWjnB4HIVCAEp10qrXYFC/LF9PlKhnVvX6hNyTK/qYF08t
v7CFaQGaDzFjM+eBWhRzncxD4AZDEVNqisH+MvmyPSR/mg78QCb/g0K/IBQYr6Mxn2LoMqleluBz
Xd7tMZR0cc95mLd32HoJ6srpktjwwOiEro3HBnL84FtGxk+DUyZ1AHyK9mqwOHzMSgIAeGuN/SvH
bz5HH/PgQndau6RwIpQ4m4G5dNY/RzmO9lWYPEIcC1TRVYDGNq6FWCMKHljGbNS5cGlva3um+C6B
CQ6xWbOr+CMf/w/oH0NLMlgxH4G0LCXHQQ7fjxVn+z7x+0jlcTP+dQ8hNwLeTlTNozneM205Hc+0
3KLx+I6Ec22IlpMRK4l11ZEiP2XACONzLhwMGVyYx4s7m6efBqDWK8uTxgh+4T9ldswmJYIM6LcM
O2McH0vXpg0O68FmWwm2ZB6vgK1G48TJsX8E5gVaOQPH5QAVXC3Sc7cPwZ1JBWj+StylizLpt2NW
+2M2l1TP0YwPMXrF6fEPMdq+rTlAE/SIqDOqkW3XtMVfxELH3W4nu2GQHm6Jze5q0w1QlSvztKqq
v3ygLgi1UNQgcGd0mupsUcRAF8foH3pj0FmxW5TRO8YMrsC9sMCz6OTq34/R6e+g2zGtsCd1etI3
32VIt+J3mPs2FjkfWG1xw1T2YoyOfTwmavi6MGXnoAZ6VN7KfnuNKoQ4puY3/bDrpEdDZNzY7QTi
FQ5N8CKuc3ZUvpDudhNDCuR+U8oS4tT50pJVaauPqhXArvACsFN8sB0FubrtnnZYbvIuIThCmHNw
YFJnF7mO08e0aivHwLkWoa70B34lFhcAzAdz3kFRhPYSOeCt0UQfiUouPw4+HhzgWvY9tik6+rJ8
Iq/E+nlMAwVQxlOn7ys7avKuJsuGTurHz+zWO3hCkbe6z1Uvo1kQzRTVCV8EYIReqDWk5YTnu/sn
5/xO37kYzjuideBeheLo+HBsH525p3d+jEzm/RRGncMy6z5qPcfYt6qFZLxVAX0/kgQkUCFoMYFd
ApobIK2ZQBzpHFzYPV+TUPWTBYQL/31fIDXei8SUUfDl8kRBa3tQoMkzo8Ta8j9OGPckXxr6izg3
nTKau7bxefxR1SJHVKzLvsey6rdxS0KokJz+47kkvsW4Xcc7p11pjqp8G5NFYMXbbcVGGg63a34Y
D8dALL1Em6+aoFvaEKvR7Zv/9KWFU622WUq4uTNNZpM3SCIkUr91AwoTl5i56qe/osh5v93Vpvc5
M3vuAQTiau5J08ZuImzpqcDPqAyJuyz67k/C6zVeRgbayaG44CoUYYhuLrddqhAOFqUiKGb0MZ3a
l0QjiWu/U+sg/qGkSdLadj93geaGoe//qhfbK+TGPFwoS7Zcjcwu93TruJk+VftP3hl/iRf5EkUk
vb99HmirdyoDbGsOoz8fkLc4CrBop4HYdsmo60f3F5jyRJ/JmUhXQQakieLxF9AhQ1xdl2ukh/hK
DSkmW5Sjih57lORc4sW7dJtXx7UTbtc9tfu0O9ReMYq2s/wvuSCX9IDBYbr0oa7CQmvq0fvE1w5T
S0qMD70NF8f0dqCSrSgDsTf5r/52bLvkf3Q5sJKqwwnWFPzr5r5IctGnjMu1UWxArS7LvOfcuYkZ
O1kdk8oDMbAs3LYzm5FcsCyDAjeMP974G01HwkRUceu0YSC8/Xp910Qbyy6Uqvp5TOpJFzuNn+GF
FE7d0dcSQ/ka42tdr/2radJSDfPAUovrlggy9oSl8T0CFclNGlNogV4wLccWUZdpToUv3cTHFV5a
Cq4R4sRtTdCX0rpMlOgTn41xcYltsr5Aw+mPg38Mhuafj55DEygci/E9GOAIFekaz1Po9YothGHM
EQUOgy4F+0lnm+NhWL1FBd6FgOyiHeCHjbwqbhiyTJFPckKJ41T+3BdT1PCwiit4SxVOOGtRAr1l
DDaHERAY1jHXfwPbC8xFMbgAKQ/qFlmG4PRuk+Div0uTSvNnUo+lprLBFUR0wZsJBdgIFDcDrBzU
oaz9SFDc7xDAPMso7f31IvtgFX9vKhCuYMz6Tkm8aYn1RwFjUtESyBoQk1qheZuMF7mC+WV1Wh4w
QbBpYuedpEEuCYvV8icBDPJP6QcJqvtZx4apLWbjE572lBrpF4FYuxD68qc9OCccRo1TkxDxoqrF
I5FtZ4cr7hK9OQxSAlYlV8mWgIKA0zpxZzb06axRbLcfjakYDj2BWA15Co+244xQsEdSs9Liou9I
QMU0/iEjuTM2CxLOa3Jf0kMDajHngeyF9QpQ3+Fl8Ewk7HWzOqBApDTNeV5Pm0EWyAEENYIFNDPj
grxKfc5PNinsskjpL7HlqAVWJoOXzhgn7gylGuOjncM3F46xRJMVlj0oO7rXVv2E+sdr5XxATx5D
6m0hf688WxctZWRnb7bhu2WQH86/D6h3LXF42inV40oVElwjIINjxmOvPR+ZhvttIPHLFmCRn2sG
nahNUfvZZ8fs5uHUPAgWGdIasPNeISkB7y508g7L1t1zIA6uod29cg+/9iCxE1ntHCIP1Ir0Bq6Q
g6M3HdQ3jbLp77pPvGIX3vALdZIZyJocUkqPqgUkYAvUMp8GssJ7msGptvbjucRiWZ7DXT9O7ahU
9D8kxw23QPGq9Bo9KHHSY/91qPZOi27I57Yv8+avdYgnmheEDDcEciynbeyYvPGxmnW80O21l8FO
Dbd9G2ZCd0EtGnDJZMMYOG5wvxsruYbuX7NWl1iomJTvUHWySZaNCVPgcs+tghGWuz+JXE0032UW
jxEAoCBRpRzYUE1UiBh7BbL+qYtAV7oNQBLc1XCy1jXMGF+5FLXBZ1WZ35lSmKp/IAOHMcSFSlx9
6jYrEJiQntWucX1AvudeNm1I6pfZXH6LBlwg5rBKkLA4pTwt4Z9E4SMKGo9UL7wqVyfwtD+ChSLM
2apVaBqKt79rUdaKYe86MqZAwyQii9i5/Us581z/2aY10piblyMWCo1Q2Nox703Lm2DzlGkkSAp0
JR6k3tMiCF/wBnxwMkILMRNZY77TPvj/cPMZNJ102rfGHGoOAclq+vfpWFymuTIaTlqPG55J0yid
u8MmvrpdJdp1pu79QeodZ2M17ECeR7qzcYGuav49QrUmOKJM6vjAKvDcuum/OysRlXTk7Up7kBjj
mmY5dXg+ZiOsjHvUHKNeXI3kUIHAjbSAiXSOjuaiKnrmGHjcafgt9I4S0ZZ5ka+bhqXU3a2SKBFH
ss+4chYBoAUbS1YX1Yd8OP9zYe9hgjlGBprKYxX4BM0cDKWQ6j1e9k1LDcl3IKwo13flUny4VoGc
rh/ftKuFXC8YJ93kMnu0R3fZOKnCEEK6nzO/vHSRWScdtwGe39dALIVU0JakfX+IR8gXVPQ/uU5M
nCTpatqM4iornIrGfZDf/CCcFYb7WTkFjDev50ab4hhiJoEOkMyLyt1C7v7dkxD7JhXNV0cAZCJ2
xh+q+qeO7kw91oC1fpmtgzspI7qLEBheUn5Hm/p1w79LySimRceELIJtsHqZMVZ70l5vTpfSBhxN
1XtwuXaPPy9lRBCAWLKvbNyAPZe7vCXc6BIaYoBontmb0bzABEhqX5YytEhkZCTb7KP+6oYSUPd6
nHN9jA7NAecmPwaHysMQClQte2rA/ayDaEGERFl4YjZ1QV6rXK8eGoqIPgtTKAhOQK/GRG6ZpkwR
ZWe57dNinhfw5Se5rMiMyTUxPrj7WGMzeehCCsOQPY3vCOJygtbTLZtoDyKruB6BesklCItRwo3p
I2le4kzdtNLzakoiGIx8wLHVYTBUePrhGeuPsVCYa0IFG7ErC2rYb+A5PAy6PLzyrEeTJJrBuhKl
CIZ1TZEvZwuv5uTWLHUpC4TDGa461dfaBmMlKK31Et5rd/9CT17mL/qnbSu3gvlPrYKzUfceAquF
ceb/Tvnui7eu+eoBWeyJPV3haxeskK8TTaCWxEiN/ug05lqB32rl9Agpk0O+EjazmN2GKVh2gFKy
UZggnlfcKP2aj1KMaiFDClcahbHp/ZtSefZZhX2Lir2luCcQOzr7ZI95Onut1gCO2aivRQfp+cgJ
15iFTEH17yA0rDI88XX5tIEbUlRxfISIMeBG8MGgpOPHf7luF9froXBRLV1bvqmLt+PtkANzoffi
ZYUCqzwR75WJMKYFEQx8usQrggHLhB/xSwdkOHXKW2zenKgAlE5+gbuA3oONlnNy9JOHL7mov8zm
qjH1hFkOleV0OKSXYEzbzskX5mrYmP6ZapCw8SjGZZHBFsYvCkp+ZqOZTZtALnptiOaTaT+wkotN
KQeoh7DflrTgOS9OAAse3innZ6AYv9tIxi3ufFaBGCuNU9h0L5smp4BQ+QwWhFNTv5nJaWWz0qIr
H8X9S4/RBS0zuANbrcGRJaKoBhvQGXElXY9R5jKmGtYG9KBGi3kbfIam3LigZ6+SDCcRQv3pq7kR
jTMgbD3uw/bp5PW2t8glf7eoCjW63CwpgN9zuPVUrgMXGF2daiNcX9qPtstCo/3eXRcGTIOGYdBD
6Xp3KRdg4tC/FOBwdxOhHAHpo6LqXO756tl9clKBPguwZ/6GoGqr6YDHZ3MpYEznVMHI3i9F8HGF
lo83oOdQsVy6fVQj+voIAvVap5zAGXuDzs+Uu2oFcp5baxJ5vhp0Z4yiF9c17yRY62+lCcmjGwJ8
QoPrCNud7c75IAlVhATKF0JAF1e70YmeuTmKrbWsOBpT+UO6cSZtBuSi3n5fRiyz9SVXM4WgKr/r
uXJJmU96nBOB23zJohibKo89lmONcb/9VPwHunZfG2zxdHEruz7eTNU/FyY1iF5gLtWqRlymVpbx
wDATU2ySznjj9bsDw0nN8s6x7SAe/wSaAXojHldyVQSWb85VcuEVMxrufBsn8/TY+FZ6cNiEjTK6
+5tcgDwhiP+JszMZfAEBJwBhn9Ui7eOWOAN55Ve3Ezji5CvA5z7O5VLsgZ1ZS1KqQNSxBu7mJhHL
HPHeUyWn8QSKzG4IWEyLz0GW71EvOY/t/XT5jAV83RWJHNSRhPMsnDmRKakk2gG6/cB9+3mBJs6L
xKlVatVYwTZQvxYQy9N0nBoJyuivBJtrJfNYIaoZR3S6jOFx+Zt/44YAnGH0X4jLGk+KMT8UT8h4
9wt2/8GPaWzVUFU4+HZ8Yw8iy4EnU9O/vF4JX4l0t9uzEvViWBX9Pb1R3WgUBWveNsrLYQ19Exn/
PjvnkbCtyxgRvr0deeMQ7uJWtN5CQNj1PvinH+SkQlevbBfen8cEosABDaGx5vv6chZimLWFkM8c
xGYcgk7tjzJcw2tS7QfR9Z7oWorJ/ZoPJU1n8NSDbTO21ZJ6K00Pk6amHS//cSMWg+BYAqMXnWu5
DFqPTNLoAY1gYPH1RGuvJtreKDUIDve794WIM2OBy/MhaTbgscefmgn+eVkdncytiUPluzT3srYe
zAAtCz5oXANN10XBV4E01xS4ORID8Fc475Wtlo5Jxe79MK7r+C00jkN4vCzY8vovoBDWT9fERUSi
1ntK6MNJvE6rUYSafJpZrH6LYHVPTWaD9P2Y5s/lYJSiVvDv9YJLRNjhjHamoq4rGCVIzswkO/Ag
cv57Mv7DfjTu3YTjCrxsjTabcoz7RjT/pyM7EKYa7BJ2QcE706MiwFladq6UgiPFDjKIZlAEX9xF
gSijDnLY4lbXIP1B+owsqS/ey4OMt8qJI2GWoy3HE+fp5ksLG10VqB5T6xiT44S4egMs5JHORKav
DhXZSItfdmSwcfYwRpDhWU4mQ4zG+8s8VqXVk45jian/oBxyYllHtxcVmEdsvGJpSNUA72M/QoC1
q3x6nHEtT38PcVtm3yvr2WEzXKPxuvacXs6oZybgdIp0wvn/ZO8zUOBrhDsklFbKTdoJG4Do261i
kN34i0qGmoeLaaiS/1TmybhPd4o1DysUdWRECZYFatNYt2Rd/tiyv5Xeu5V+uytDj4tMWY/Hk7BI
6ZDDmU2XNymK9tfulE3J7HG3UgNvD1guQbXYg4pa2LCd6jeNuziFM8zt3cTiw0zGlsk7c1PNOTLc
1S6QxtXoc8SPNA3KneypaONP6AFXHoEgFun1BwRuf/wH3U4m4ZWKONPBvGVUFe7sBG8rqfb0O1O1
Xlq2NsXS/JTB2MQz3gsdDLLkdc2ymZUxXXMBfJqV7ObBE00nPLaucV3vPpzElfNCz5tosrKGXEZU
sqIQoCII3Ki79fXUzZ+of19v+5bZJZqmAf5pN7Ka4p0I7d1l0Zw616xjACRQxmUsD+GotBe/rrFi
jG9WVvulazl0NOGlEiFOnWaczInfxuV1p5irkz/LcwImjjR5EKtXAh6XrzcR0CkLv9q6HxLhV3SP
+ykcXuO0WPTC2uWRXjVG2q5AgXxiUzQEDF7ZUGftosrYp1/uq+u53sTIgWPmA0DO9MSb8fJfj3Sh
Gyu0wuuhXUryccw3LnIVMe93JmNUZFeGJprknpqE/ojkxFtDA+XfhtvXV2N3Cwr5EDlQsOZemFaA
E/8hpgVCEmkIrHjIltMeV3l/JbFPcwKuzUbz2OWuqFHT3Y35DtXd4B0rILhMdD6phDqmiLa0JmP5
3kTSgfPEKsU42d7S920b/ICeBfF5NHtd8DOqf6WItQezcB7y3B+ScnfE4myobg+IECwTLRXr1E/A
1wQ3Jjkl2hCBjl6bj/4nLgMFAGhh6iCbqvEz6D1rMeR3c2mNWwp622xOGl/nTb/3v36gFrFMkKKJ
Y+rCrNSdnnRly/x6Li0MX2tFJ5shuBrYF7am1JxMWQgwaeZN34N4jhsPwKdz5eOrztcngx2SM/OL
UT1NXd4O3m4RKH2KSvfQHF3oNQGXXYDOIzO+XTn0BTfqu3LuuIyYZbPtC2NadBIAekAFIiQj1BEQ
jdGCOx9ctHTD8jH+JIIZKgEYuHGZofRbdrVCf+m2TLMwTuWcRG+fQm+pKvyiG/Ifp1OTQ2sOXYqt
BnIJQyV0EX3r2vKgcK7IdSKTjLtp2Jvk64QIYIv/K5/a4hJsDS9szUCiPazBbvniy1eoKXkFRH/Y
GRy+vtP/KMFoOIASyPa1cS3fBfDaYzFgr3RtBXOtKl5Zm3uRyp2muIuLBRZ3PHsqdt1XKMTbrn0J
nII0Xmr5wTdxywog987lUGON/UIhLCI8Xnf7b0lY7CB2LE0lwXQVuV1nit+kmDxK5Bt8k+FG88pv
6gUbypbYSqpbtvUNm2ixY5lqu9nYncR/6eYGJNcyXHMzwhU+DuN17HxN5kVvrN6519CPTfz6P2tR
fO7/FccJKr3QS6ukMo/H5swHaezTiYBDrPjRFys0LCFua5R0CpV0ke2A6yYiFC+iwp5ztzYPmOeS
BkevGQknXLCKLU3Xv+xir1JkZKKXlM9VFV1YRnnFLSQsuRExPLXN8wPqThLhhLHlhKhIhB/3lvgl
bVS6M1ZT5mpMObSlzl1O/Xe0DF1djxJHJuww9LugCcZmZnxJ4wu3QDsu18V/YgEoaU6MK0sugXTL
bkb7NOqd8lpT2mpPPqgSW2bnk2jhibtWKYjYZnyi3dhkWUZkFvx64wpWYQplBTKvm5e9ubq+GdHq
emoKS2YPjp6jt5ZD/a+ePseYszQMhdUtJqhCA8gJcfNytT8zWHreaPD8PUyFerixNcDvfFgsT5fl
6JCS3ERKp+hoEwykzhhpP1sFrswi5prdmM+azZHD+/YWIj+9EC3WqvefWGZINOLhJNNkf4hf8hFz
/sqiJeYq6ukFPyuXIvqDSiLKwInPUOzc60mtAOcMm0qk1RURyR0QwqEybfsPlb/m5LDba+tV5bqN
4/IGMDJ0oQ03EF/JWg0grSVFzm7nscWB705117FsLQzupdaJyUcEJxlC98YpGtoWgzQ79Tmzgs8q
sOB+x3eD9oOozds7jw2esXMGzdwDDgDaV4c5sSUEgE6sfn5ypzAXkO445vQR4mJGaq7459GBz8fH
qdl56RlB2qcKqfbsodQYbMVraWKi6LbWzE28ZlP5vaDjU0v1AtQmUegWI1mkjpOASDwG9s/VTqb3
QlgnvcmdGCoo4buIGuLagp1mKyC1t2IxLBnlOsh7UaieztGh9nky1EQupKuRUckRDfuuwDOH76MD
SAe88br/Qt5PGF2G7pGn0TjLRmj5Jahqlp4GZXkvnFcNpWJ03l8YkXeQ1Ie6F1ZWzOQ22oLlmgRa
w9pM/GbwreITSPHmk482NK4+sSe2J5u4aAYYPgNIxLrR5RBTkOjEsMXrw3c3wtXGcFPuEUHH/jl+
8iEy2A5b/ja7o/PlChcXu+Vn8cn8tuTBRln9WpuLUqwodNCof/vN56UAr9WD5AUn6H97Ey1CmFaD
M6qelFdSVNNa8ZF/70TM67aktPLgQDpk504GTcUWXtukvmLidc0haUonsYvbdonTM0BdDqEMijct
t3LieowyCLMMgMRoF9KzLWi51fJMjxvv/HJesIhergV1oHO0v2wD5ioSpaXguV2LzvY6D4IioPTK
YjdAUK4q/AUVNYi5eo94VpRJ0bxY149obJ6mx/c2h54LHIbWoLOW/E06RULb3mOR7C61zxFZ7sxA
L3Jc/EDeRN+zj2PLEE5NXFqF2zbCuHqHoPF4Y8PSZDRLZRKPkrFY1u8pSK9LHx5LJyRohZU64rVT
ZYB8JXgd3U4XWK/f6Z+Jk+ZAolNO0Ch8RwOOC85lj6uHOu8Ux1/uldZAzsSY0tpYDm8SKU57PUpU
FqBlf1Yy5+Eym4rG8FV/A4tVPbdHVQaQS2oExicqj4JEZUI23IUo1qpxTuhxEJ0dLhww/bqxVATI
wunDAB/vklYF473XgC/kjl/DaiosCHtB21eukyaBwjT1urF5l9JY2H7ThTHL/dopkGcqNwWfec5i
ZKeBd3tMN0Wo/goR7sN+cr4OjHVujnXSC5c9Q3Y2bQ3BBIYFDosJA/eiZYPhnZ3VNZI5ZusBjO/O
vRG6fVz+OkRQF+8iRlTNsWnStyfUhUz+iSNiR/D1b2SbOzazYQsL5sdG4pXuqt96iZGLC/d2sBhj
TiCm7Iy2ehS88QbGA7mp4gXHdadxJyj9j0ZbPVG478c60PQ+t/q20NzOYeqsLaUYB7hrvmCwZp0j
eo8O+wcPfF3b0xi12NF4U0mIZ3y13aQO6H2dUwZESFo4UTMrxXWu9IggonRIbm8RH4EkQYon1NVs
sRlpiUNhhiPVVHJQIY/E/mUdg0ewG7EKYAljAylEg1QlWFYJ6RqBpqwF+hlG4Ww8WeBadJdk2Pr0
g+gyuuRcqGTrYqmSrVlOgOksgoaP9UYuJ0WaqwAq4ZV1J+6fLxoX+iqD/Fq+9EsqKcf/ms7jPqpW
vaOSKvfvFjUwbGfe/daXDVv16ACDM4QyWTJYBvdw1AcyIepIIaUKS5rjEx13z0ZW4Gi768/TyyhN
nEOws/0v1WH2f6vyIK6dkZb8rH57LVjE3veEuqGoj3f9IwrRP2D2OeMKaGTkPibgZO+xnvUrmWH3
dqFMG0EV12LpuxdNZmenKZwhPnhOVnowl0I5+XQ+gHxNsfm8xsx5aatHSZrjPEMwcYJaxinxW/yq
E3G2XolEoiQSZ7+cv3p9AOLFYOaarIp08lL2SCA56FkQVa6tMMPPhL9a8+T11BjfZnKXuayLSFR8
iw/5m7w7mN2he/epccGj2Gy5FBztKp+jVhGSFQ3nUKTgQyAidcoG0LUuW0WlNKs+agUVDYoC9v5x
T0UtkP/hmqbYWyFalp8zW94GK++2fJYASKAfxWv39L+UbbJfs6YkOvHkrLjWxHnSWUjTzD+b6OSc
9i72NHlQ/pa5XcI6D9kiJKmstywK0/JRobOoqBDL3Brr9jN9KCj3AZb1ZRHMHJeiVIwH+B4KZ/yd
t0VVQZvTJtrAnmUN5LfaXj1RFW2aFc5WCxEibz8wILH0Mt7L6ogC5AbuEj87NFrGgZRazojdqacL
512mbfVS0Jzf5Zg06N6xBOyxVofWD/um/awdqUZ2k0l0WJhF+q/8NitMMPI+Cbjio7wAFff/W77c
lisG0teGakngrg+xD1POCOo+havs9M5QEXssEKEpeIzTWbnWxVmQOf/gL9YwWC/vqLjJ9mLooXYv
OGccyqsX0Yz4ovsUItdeaTtrZF7Lcl+m41+5OoGkv64durIoVVvf2vpW16gGVvGrMDv8ybpOx65Z
QQ3LaC4wnow1lRKfhP4hmKuPIUPga03InQIuRtyDt0Cl/MSXSm7IETqefeXFbBICXWTH58+ginIf
HvpNj3o5zg957Hd6I6FMQK6uaEye/RQYMu20VTlqO4UfdmsS/1MevCHsjDh9gUwaDcxAS6jJzwM/
tqzKtFSlP/SyxeqLo/CSLFoIUP/8+sHWLUnitZKBLGX8QR1aCsxHhWx8bwJY7t9cTWqaD59gWs3o
5tZe9LsA0i0bSzZefI7CqcZQ/5q0AetJn0jqDZ/hWCUVri6W+ehrZ2whK17stJlm21e3TuuO3AUm
YMyA5NHmiVXC7TQI31peotnFdNiDI+YZ+YUSxz6GR31aFT5YRUjwjWwFtsY1FwNPsx1v4+b/+jJ+
rzVrNYDs2BKVWxCm4fEqbrbKuZpqi5tEyYx/novU750oB5kga1PaZ7cVZzw2KCFXj3JFDTlQZ/Ac
yc4ixkUzlKwLc+W2FLfNojetHQHxeOqgb3RPVc6xc3DIqYw2zp/koRv+tGY4TBDVYKCrUrXIgbM6
y91poIyHbEkCYozWY9ttDcNR08LqS5lbd3ntTo4Me/u3RkaMwno9wxw/US6QenJYdaXcMo080d2I
sV2OqAL5Fh/5kAxzwhqtEJlVxs85DWp9hT+xDP4L4+87KHna/+BNND4oHm2gbz2EqBPNZaadJ9Dt
N49rJqRYFZyxGmuATGC0sNHc14cTFxdZN4WGyF9kBBxO0qMIVg5sHfquaons1yKv0PJMNAkOhoXG
epcjEJC7RElmT3MPVIoebfdCxAkClANCTbNz5+1Pyzm1kCA6yIyHdXLvAvZnOfxDVTRd824464tI
DDH8EGYKelr7r9GoXszDwX6e07+HpWbHwlDcjzHyxF/YU33iVmKnlSIWPXCArRsyPkUFAM9I7PLc
VJk2G48wF+gWZ3tbaS8Uq+80iwapAjYteRTV+RphhIus/8yaovA6CFp8seWQJJ6bgku5Dw1BM3oO
VZH0CDJHvBCzluxdLe6vh4W2hVC1MPR1kwecM5BjkO/4QTOMhYPX1MK34fi2qu1tLDvT/ejduF9c
0jCh9BZHQfKtOQ/x8rQn2rJSTqmDkULozEqfkMrBEDUAz7JafTL/gNfaiVuogR1k2fruiW8i56Wc
cqcneABTVrEbN9ol6Bhfk06dQkJGVmFsqDSSF7/JWoeCfjNC7WjndmZWT+DgDcXrnKkNQ4SRdPUX
5crh1nLvDB8lTzXtSrGPrKGmNzJzq2eHVl6uOVnFkPg3Gi7F3QLESbkQ3PZjRbRVzWIEpi+ihbHs
uC4J9rKLQhFozhqUbwz0skRsIY5keZViVTZ8T59XnN2BmJNb3oeyZCgL7WfvhjQp7kYUE3+Kc8zl
jDuGwO1BthzncGEqxJZek04w1vdCC2lzmAWPxOsorMEciD7ldENqwakq1/DTxXoRc/HManLYn2CF
oC+M9yWJt3P8PQtUwRhoCPzror5OFgwWxtlzz+wkfh+a8crCtq+QNl1+E3IyWG/SSxwBlXMXVWc9
KSZqV+Lq7IBBx2DsXxtMcLS6Hi2oQSCqQywahepPNznn54faKKmHhXmfdfwHZw2sjlGv66XnjB5Q
D0MkHxSTo/EEdLtOuY1jY1o0fGfhkmDP9n8tsLmPIOhRniPesjNSlanb8trWbAbe2KQdAkykLfjH
Mmesnr0hxNpDZsfTW440ZNjVJWvi8lqFKIEtG/lv+979crfkXbQTmsNxtkL00UDZJ61mkneVA8zP
jR/kX2Kr8dNpRY1kE85twIh04BkWXLJ4avj7nvsQzSATGGjfo2wqSPcWvqcMBkvuyr/ebPL0B9Yu
phojEvK8ntenEY/NKDLbvwpqn39S0wGjO+7lmbF6wfqbXpb9L5BWybqV0CeCniYwWFkB00BcBa1W
dKPMzNAD8WgJ1OqPXFSm5sqgjBVx6RVtBN43mS6wgrWm1/IeBvqiWwu9c2FWMmnfdFRGqv9CZ32D
eF5U4CexMkt7vYcokRLfA+9maWkvEEGBD+6oM29H13TQvdZ7VOvMvp98aSpj6JTyDbK+BpI3AcAZ
cSOMpz+41ZGDKi1a7tfp/MHDxlO5Lvkf6q5DO//Dy8V+Dqf4P7fW61QMxeNnwNY+XnUAfKN+MONR
xX0YoG+m1QMitynNrPwloOf4aWlG17MRmFwbJXUofa5zEtHdobG+wmEM9/o1C0JNXks6pAMeiIgs
vsdcYW+toJyAe2ymiPAf8y8kBKayzBxr4+Zy2UBvNk3+dq2D3jNfxWSTjkh+yLAHY1mQoSnCdsVn
+YQ3PaZ0HTuyqqeljp7mWiz+j/cslwPBrQs87k3vLn9pcfgVDC2QlhHtA5kjy3GbwW+j+R94Ufyu
HUjABgLlIjhzt+96pArjDjTMNp65qhYtP8mxb8remfTJ8XAaNbLhBOFt675JxVLXVoXxIkGWVICl
YjOKFmhM1Y+wsUQOSk2T1/qkikqlqamgJD8YDhEOYos/ful5q4DxrJWae0Bgg+2G2XCjkHxdIjd+
orq3nc0PSkO+UtyRSMav1lyrK4RpkfVOBLLp4obSEZR8CGtuYeh1Aig10IPSQIrzXE0pVqu1xOMi
Rduf/ZMGeWc9lD2354AIO/0TI7PXM/RhTLzvUyOCCRd2NBfc3bO8ShiCKccbT6yWLUJiecvbOyuC
5VRKJfqTFhOvJ8zXpWTPg1cIcmwyafijkEfzBLsFuuxCqz5aHWZaowPkNUrbcDoa9KAst/kDX7En
KXFZA3BV//hxHa73BkfWi49n/5JvRM1CVn5uvn5pHbDqpx6rgNiZaOGHS59Eo2Lawus7/7JymDnF
3UbwxSnXUQw5nGjMCveeOOx7s0m+ayL+7DS4MW+bMLK0K8lyQZZ1Rx0X6OPtuLlmvnWsMZ92fil5
H23/LlqxX75iOn1cPZY7vx3OUvTcF8q9FPJaZ12RvM4yNFL2H3KaXYh6EHMtEXj9/V8gcQvRcIKc
odOw3KGKiv5uFjlh3oCfCqma5W2psOL2rRCdkxWRiLN2RBckP28J06n4OU63DD2dwET14PHHpNHq
GQK+aWRw56/kNb75e8z0WL9ZOMjq1EdFvSePtSKbTL/i8eYMEh3BPQWu2ihQh+QAl9CRn6B8fV4A
7bBHvUT1JvJYawln1X5KCc097Z55GbRyPBu0Q6KqSJJISlmvKHnpLRLFZOQnUWqorDufRKfR3nwJ
EUc8A8nQ+8TIZtk3nSz3ipZD3c3BxhMclDcokjswFX2cVZEmgOnElwN84bzeofNE2TgIw10eXxyn
oA6MM/6Cq+EUjOdzSCsD+oRxw4XfB4bOULluoP5NRjIs7pesGtP9j9q2KLepYKk9HRwYvDehYMx1
FOzBH2kVo3d25pOhr+B/ovn0aKLJnYAqh20mt3fH/SLqKxY/8kB3NyBr0vn6RhFtGbUmCSBcncTq
Fkhhz5WOXZyWLDX8d0JBzTsfx6vjtxUQP2Ck/yUBVc0UlZP19zbcmlWRggVos1Y66H+KU9ZaaCpy
TxtCUs5E4PqYr6PwePH2yn1PsR/wSt++ZjyceX17aBUy+/cNEx7UXXbMNc1NKOdEQU1cpTYeJNeD
AKdbC0dNMyKPxxC9Pg/CvGFUnzV4C3AzDgVt9lTSyjFkeJAr8tb42Wuqzm4BmBXRcWSBcnfYVRlM
fFnYXVjOapwFTpkLhBWgQPY/j8Eg7ZIt64UuSQ8pWtPQ8loVwoFkAnePWIxp9CFK5WkEm8dv8kRn
5ejF1oOxyl0/2vZ3KXADN5hePYeWDI7TXdHJaotdwSJpaRE7CUl5kOR7fpywdZe9JysTewdkbL7X
IKTbVanjQqBXhQrju+v9T3fFAezO2uoEbPYKjfpvssG07uEfj7jgFcFnBmP10zTPu6OloNZ1nvfn
2YiTc73kyoQvISSj+oX0Td8dHetBqLSjwjinVCrYK0PyoV69fskig980hmSkn8RIroYXWphg8S+V
pcAVGIZ3TbJqwxu6yg2hF9FTGN7XENKyg/jR0FJxYOCr3h7E61FbnRndE+ACnmmqne22lWmYl3Xx
//NKtBPTTtz+Z/pyBPvdqRULFX39w03qRiaH67GM8FFKf5x10RDGTINQNOXqUa8g294XidHMyZ6M
UvG36XjJtkEHbePW2XkEYyGTc/Gd+4wNRUHBHxjKMJ/rLk+GgyyJCbaNu+dPpuyKpSX+MAdH61dP
BgTWSk6J2FdJKbiuR+gErbfJAU+JVIGWy8FWc5jZlO1X3LsIlEdi9OxM0GiMhTrtA14mR2nD4ohS
BhIPh069Ua5LJgROTglk0NvcFraZbKHuI52d18y0h0XxAMpZV3HLrtezhJLgwQvSXbfuRdsvfGLV
TPfVguY9oQB3ZpcECGIOpDQKeylbSNs8EZeZPTPvnu/NQzzCW2dCrErLymPFs7R1PXJI6Ya6M5U/
UOMputZyjwHwRe20DRj4j4096gWDpz1j4pO4+f6Ry1/MP7wtE+9vNHB3fz3aaOsdnckf8VneHgpm
QaypfnSw0GvPTxL63Y1ZjFV2/clUYGzYSor7V1DeSTr5m0YiBmH+RK5ZvFAu/nI+sMwGHyTJfV2a
ONG3RtlPSOBGkYbQAZEnkxN1JcTSEzFgJF5s6X7M5ndOFjAor29LpGvVEPtKtcD5oH6v2jikaJCS
KGRG690/E8YqKYU2z5dIYRRZjJahNTPProbXF6SR9T6fFLFaE1k0WO4uO34lsjVwIukXhGpyjKL5
IIbgOgj9AP8gctM59P1zoN7ShgmYc+FTooWaWBQOKPzYV18xhWUOpN3g9YnXWcj+bEA/ClJtJPO2
NPG3OQW34RHhoe7XRWrFL6GiqM3zPHU+U+3IA7txIISkli3JEdBHSpfGSpZhfR+1EKfkjRT4vl0a
dbZ/rnUcbgNOvKL+mz0lMkUKZcT/6o1yg4mNGgpfz2WtZjdo17/fbVuBflqgjmtOWiZ5nvEBkEnd
bTCRQwEs+a/k1b74oY7noRscd+/on7BIem8wuxQulEMpq8DQSWIlzuseHrSXrzGVz9BvH06ExegF
CtkfptiQo/xroRT88vS/AHQW1u1DTACDV+bqA+I7V9Fs9t1Ya1ACZNinzvxmGPIK+xUtMpJFyKXk
FCzTnRUHgyHNZOUxfquHBys6ChBZdQVxWuYjLLRRD5PMgZUUk1QcWCSGXdbm4xrXQkbNOYvVAyoE
SRHRCfGKScUf3urxSl2SZ+gB3epd3CVvkdFOZpTrZznouBQspXLB/S6TIwDAbI4RRYuANOCS3aOt
oWNGKeQCpej9TagR9vMdNsEiH1U3Vam3DAXk9b64HrLGU5mc/ON867jobYw0Q2P5iCsV8Au8PaQW
vMDYPtLlyX32N448NQVUC6B68UwojYwmpqoxyrD+j8xSGweCHWo07Swpz3vWNg8Wqo4zLoMIjPhp
Vjzd7JXK5hOKSvN8I91B36bCbWrUHWhikaUIMJQM+E0paE0RLDrPHi5GniCutWpXgxRknRwEYK0+
lCwz8U4HoHRhFjtiV/1maCa2iJEwvM49GYEBqmMWz3b2OXY9G12VEauJvn/G/6OgW5BBJAx14oH3
mo/Kkv9FHWqcGwQqXqtADMzsjSq+wjtzge+xlk0fYRNa9N+op+Iye49D/qElQgp7qI+fiJ53n60A
ollvoFJ9RgoSoO6BbHz5tMNCL973V/L8sI7VkI85teLqU/EWuflQpS0UNh0To8tFTXD9vRar+3v9
xUcSj+27fN3DVduy88aXA6LjAseBbsrHAJeNPqN7/IpZZ4X+MK2IL3Yh/rdMw06qxDxz1o2wCNEo
h95cprI/o2cDAXGkuOI+SaX97FmemDuNOws/S7pmF/RUKWBXK1o4DBekN6K3JlTCzq1ouHpy1WjU
OZqbhr5soaFCfb9RJ6XlHPQe2BVFtJ6BlME2BgzFYsrk/aiij5FLYxUWzsoQdyceTXGrszmQWHN9
/MWM1a/r6D/udQrYXvOsYTvrYevOObmPj82p5pmI3insFtBFr4WjXEsYmcbhTMOfE/FXe8mzuDju
eLqP5ISx/KOCzrRCYC0Yw94ddmQBWX8btlxLhSryHg0Saf2YSdO7jDA+FWW79YwInPSNqfUMGjbt
tnk4JT8bmqULDD/rw3HuvfBSzTquG7c+5W7W4VwiCXmVFXEeHHLYGxUHQ0z8Prb7O7/WRsOXQj9f
3mSjJxQW7wdakOc0An+vu5yZ3yXBg+vionYk5gYymdUzMQjoBEDhhkSopik4rc5ak3A3gvvqD17N
rJ15tta7Su+XCrgHkNBzPAaLUAOQKGOQGV9XAwdgPC0H9hTjDkut3pu7iLZtJcATUonw937B5yS3
dg4dVYEjBo3gmGXPfSrILzSZuGfMUVjLeR05CqgGOf9OFrL0TL5ZCjAUantREn0j3yuRu++Kri+b
urwF/onE4s+LjMIHvhRYikhEtpObI2zTfavNSCeSYD4BEDFEWRJY369Z5ucm4EikP6ctnGrz/G5Q
UpZan+tsQKkZbjQKQZN0qQecyw0eqUBUOqwg6nF8ccZAZ5gv3cMEfaGEeFU8XvhFP8RvOxV5QjI0
/PYLmoXq/uLXOf1lsMqfECVa1w1g88n9md4MWYWgeeAqCfwK8bOlyPDzaecARx3LpWbwOwvT3UUZ
Aiy8Z5jHA2j3xuyecNlJFcBp75K1lJhdT9W3FxJMRLeWpJcKbl7P4qjOA7I2zRTcAAKqfYTqavf0
icAR+gVinV8dN3PVt+bevcxHS88C134lH4nQEDA4K89uTjsRRY7BYOQj7vesO3Fe0t/vRNWSfxiK
8imo+FgG06EO7pd3NmAMLfzUBK28bepqVnYGK2IjyJf4UViJYfYdCSMOf7dJQ9gt2R1W0/cx6Guu
DHzRs7+RTUxl5/GpPVmRfgoR08B9didsrAhwuqNeNekq0ceTHGKSmIzTOfZ3UXzze8q1g4YXfrdm
5Oot84rD5uUPNKLXsrn5OB8uc6jtG6TEqJgaHaBFBmM7J5E/KGxl6ZadVmlLoAjKVajJhzS0RwlP
SyA7kl/C+5eZGauOALO7lf1Hb3Cjgf6FNeoT+HkgdXrFkFYX1fxhTf1fn+E1T6/p3E1u4CliRPm4
XUc26amDbfiuEbjj4zUZiZqyXwzOyc7mOff7nEzjuzkZ9YTGaXBqfd7qj2xG3FabyAxRc5yi1ygX
l6/I3gXzMU0kLTHcyMnu3Mu/QHoaxjo96R4OXkaCx7iPRIBwqWviqFj19pWFZyLmm95wiw8RPo+c
6/2jQDGGgJMUahpCKjfiG1SG0PmxjfSKUn4RBD7o/L4kyKM88bpNq1zIYcHBx/wA4hk+P0/2YMlO
EL3261nAn4JANpxWraA8TwQTGtjlS30JZy6XS0kMV21WmRTXCcCPUhCMnGWReOSP3ELp1ZBsAWYd
fkJWMgefH9ZeRbi2D857m3fRccjeF+3ZKPstpJeVeaLwOWN+xYuNpMPBG0sKZEMAaen1y70cM6ny
GzJHBfmpZuBKIcFUfF9DPR87+HKPK+lusqcY52Vm+Dd/u6i+TofCv1toR5I3imA+uhuoz2cgvsm5
fpf+hR06acXd1ctQBFhmbuTLTk/E7aZJLS8vDk+jHH0E+GW1Cm5E1aOFoC6ftrt9sVwfTmRyHiOw
3s5fq7OFyLwE2cfrwCrCjWWi+WV7lD8jKS+XXWUIa+Huuu4biADNRrPpQUsO67k/238BqHHZLiGu
5tIIA/YtCaQPcwG/l9IM4coJUu/NlLs/ELW/QZdYvGCfU1b/UfZuON0IjSshFwvXL8OQizWRouYn
o48n+w9vvre7Ulfh0UWFlLMTSQrohZHYba6K/ZL2ZxkQv9+Nd+eRcsQz+Cxf+qnojZkSxyItD/ot
evCm9WIX37NNOAMhQEoLcDoava0ZzzIjIFomzq9Mj6+8bXZC6OZMRbeJ/02srJTLVGs0q2mNsfaz
mGRsg4VRRvlPatfO2FXrHoAw8gwml5IX8okDhE2iKYViJUlw6WvhC2Jwb2fVz+SVxHnna0ZktX8h
HrAR5zepaBsTezRxo3eHTQjX0E2OKQvfh5BycQWmfXl5KIamZrhR4kLZsjwnwn46hfGaA0kqladQ
dmHj/OI47joF0kidl5wLtWLEO8EWzhvbqy6wlNke/pr/jEHzANGOKxLSJm9Y2Rv1NWiNkcBRY9yi
a7b4UcDFsAIaehS7vuuOzPm7PJwKlMfJFEkPeMmxMW2CF+11KW+WA2DGMSxG+y9PMterqQ0r45hq
H2f0+1y0HjFxM8AXxuCypwbTTvUia/RXqf1TY/XhQ4ZjMlgLzZHP9S4SPHIWM9HvIeCbCycnQ784
AIqihsca6WCHQov8YkyNkDHPiVOqefkGPJVWa+ar27JT7WXPxCC7mWo89Oj6hVip4DE280YIfLAF
yQx1mcGFZ+ROzrahOJkCmKrMylqVtvgaXKU6ehIWFp6YTWEGr4KvnTFKLV1dUbEnCnqUAiTLJQhl
H2rp9c9+yjOMrA2CdHv8PHKzLCwVi4507etuM3Hfi4APjC0D9XMebuldAp31NdZz2vwSYYTNTc2b
XGZfaFnSJph7U2Vp374+Mg34PDjLtPLkz1NS7NlPOihjM5s1gTUUlqhvmTMWWLFTq0R+V8KHq7qA
Fc57a/RHzxa2IeSP4tBYFMK8NyTHiUlzyIeC+CIE8ciZ9Zyz3zPsMPkpkXPP+OeQERC34OZ94Ea8
m0FPdqI4LFn0TE7pYZXYyslgU/vWRrXPWweTh9NL2Id/LSavN0cK3p2gSLwjXRzjnAH8aT39yxxS
BRIYEzPsA38s83AsCz+IN3QB1fCPTcIEz2XXUNMOTk6B9NrAO3p19ufxhV9gGuSp2VTr5w1ofMBt
B6+QwX7VBp6OJRZLGPKKOB8HzxiRG6ehWNfq1pcvVknmpfm3p9xxwA07oyRrbrICbN2ggCbDBl5j
9Jv6T6kLOEIJFrOCjK22JPvZF6av2IYbCgphOKRjSZ4sqkXX9Bo03Vbk2nCXp+bL1tNLjWAupnsZ
stoBNXZfanH+T8YiBJXkbHy0DB8oldKgoGcByEHBhTNd66zaz9UhpUvA6k2uywei2uivV+8PWwPZ
9GjmYgk4yJ6j3ls29kpq8MQmDNICTmJSM8xOuHsEn8N6KtTlyG72L/9NpEEZsbKvPaFzTT1Vb2h9
5+doWwhToZ34Mwf91daJUyi2L2DqG3ajkGHM/9g4YMqBxaBbekRBmpVUOYpxs55QvR/PlsEPWcvV
G5bI9cgoBU28QO8nH2iyMnjUW17W1CTtAbDvsO9ICwcvCdFCijVw9F9TPb0rVOt2hO9AJofTl78N
P2UzkXxJnkDdU6Cu6ljm/SNnAl6KKQdFDyv3vsZouOcvcuuDnbeGg8p3Cpz70bctcDTaW2AA1VWo
xTEHLaeCFWlr7o0CLT5sNiWzdzxPqIZ1qv3DK+jiJeVkkqd9yu4Fai1FDw6YPYw9VGGbcQ0u+ZVY
2dkQCw58DojBY7ar9ulGgCEszLXXVYs9DhGwL7DP6c84v8iI6pthfS9b34ALq2/FhVLe3rdD4QHy
9jxQIU7obswcvcBK/Wvsr7uSZ80Mjb8C31Hhpn9wXJgglxSt0Fx2fNeR/eCGhougvnBTwBot5GhA
HebhP3tT+uH0SKqQrx8cfhFU6i3KJCWY4t9mjxywKvBwpEFYySLSidXSfYQCiss1sfieRytpNLDO
HK8WtioCujOBJlimz7nSAgzo02xS04aoK6yQc94CYXYEwk1nn828HO1HmWMLTY0u7rnrqYZ/DGNl
a+pFRn+qjWSw/P5FmrN34PIjXM44ihbilc/f/qdHP5sJldEGFX6sfxKAmtB8vwgLCeajlMpa5/uQ
0PCNDxSmM26nmQlvSvnYH3KL5MGC0wplc1NeWqJxlqjL0cTcSllpcLg3ziLqXgdJEDcK95Vf5iui
IbuklktOjxsXo3F8nMaIFG5BayuZA85DOiS6LRxWE/vnzgk//xrKuPBH5IodHiMtIssUzAePWUU8
fpvHQZJzGve6h7tsiU2yos/RTHx/gYdC7Fhh28WXHITeQtzerXyXy0OAJAU3bKqBKyjTzuPtOlY1
j4ePSpJLGpPhHSBcqT5mgEOjd48vs6cs1nhJI9nrtGAwg1cfSeqU7MWLQpebsyORNtoqRRQMJ9R0
9oLmjI9hwvk3Z1AFme+bYATwyy40cBe6EyiVnoFEcfhN6NySx6S4IL90ERIWEVkdCcPG6WjESV2M
xY4SHQv/y33LUto41/dVdODDNGSkYcZJQgiLE4zbmqtto2yAkCsuH+uXRTDmw0GH5HzNAaPRv+dz
6j9NhDfQK6weYX1My0l3nI0Hqeuv68MbSB3Jvv2kB2q5f8OsitgZ8n4HK3LZ3fZqhO+IxprY8Wxo
BCwtubvClStXbiiHcft6F1F3+3W6/vbs9VjZOXnLC2FfGi64zPKqoqxFKCz0MEqdJ8vu3mQBrL+p
lhR6pUY04/0si3apF2l9UmKKAipjNfS0Jt8mkps+m/BLr3C3Fh+eCc1KEfYlW1uFW3ICledw0o+2
FJW84/CT8k5zXSyiIzXziBEdAYqGNTH1Uw8nhUnUQLAfy1oAtSaoalPJb/CDlQfyuXM46aKRwv/k
aBxRnbi16XEsnZRCwATkFVkJ5r3WAuhyU5HEFe9pWu/66A6cU7u07P9gktf7Lkf5sW2c5wUdd3FY
RL+j2eBS1r14ut4JLqLSzL1GsU9OhESe0bPNBCxmZjS+8Ay6cuS5IdLq47luhPAD98BbsxzY8LQ7
RgLsXMlpDCYd5d/OfNiTXNpuqRZ8Fiz7uropMp1rXP+SfNCMApdE9ywBpEKiG0UHKs9KrAa0G2+X
GTMc7gw3hwTYeeKR2UOHvOZA50CudUYSmU8w+kTKvqwbHzN6vlkbURZ+PCKGwtt4eCVXCUf7iQBf
EUBbKVYEBbCKQamINbswPTwfLObKSSf4m4fV/arC0WwG5kyYlTGWejZ3Z40KDfy8PqCOWXzv2epm
sV1GsnCCDdBrRlL0YiNWOxjTtmBW1oZfP6dl0eFW2wCqAkwlQjbC+X9zlx5DxmuKVxIHL9Lpmgbq
R5O7A2FAsrJ+S0Ysv5t31F3dYp740XAyIZYggZY56c8sKPoGT2+9UXpGN3GISU054Bi7Nv5G3jTL
aE/DSDoyLgvEY5qoUw+Aiyg6Yb1pXf4qlgmCdJDS/benJKSpZAp9I4lvwIA+dAuGb5Hvxomwz7vI
bFoK721Fypuldx/QGlY+PviG4mFGUdOzCMnAg6fFQshtIfam8U8r4qW32bwFLg4W7KrQwRBMhSlK
lslUKVAw8IH1hFrWVenPLqxMCneoLtYifHoa675ZwLLn0kbUSolUmDbQGMQ94vdlpHvl5LsFtuN9
2PysYNRp7OYIYwiRXQE3C+57dnuHjCd3wQPO+ipb71XESDVPeq3Vu3hjf4gvc95jEdf47evRfC1g
YzK6fqSY2bQgvy00+Q5+zVtbjnK650AsGQDXXFQ/vAYtQggaVGYJk4R8iByePpWpVsBw6e1edz2Z
BCKDjTssHrKu0Gk5cCclPdH+fJl5hSnLjn5t+1s7Lyic33/LrS/ZgM6Su44LQspZbW8Sqe8RuoPW
1cJA15sKu613rPyBnkRtoQFsNRA4jLoi3Uf1Vmn54TbwzGqCv/mrLLUIcABP9Er+i0zYbkXdrf8l
k/kPnkYHOyqYyCtUL+TgC/mycafZSCN/PYgv6B2cMKvwb/m8ldkC+u4w4edyM0Oj7uuHbA+lrAAx
+MyVILQQedG0aWY5GcdFq4D8ywXMfTcsvUj/h13b6CejoRXg/6KdichbSO8z4jqVzJuntO4WS37D
qddALNfMCsyQaivCydSjw6HY0J6UMw2PlYkQtXDc1Xi8myWi+/HcNhXmZ2Ha4Rlsbg9OHMCTAjOB
Wo7f1GhqIbxNpwAHSWai9yUlOBaiFqENRdVbz+C/8t/IhTdvaGM2XVm9FDMblxN/gr1y2+Gk5fCj
e+aQb37yjDQ5PxslpB12GdrCcRGTKw6Phx6uEwdWSXmYcvNHlOuBRWrRhIgulmgDo0Fq25gxVKme
0rcahuZ7wpwWyqrxQGVa1Z+L79tNyZXO+WgFbiYWiPRQ2wcdW2NHiEo1lnHJZRrhUnTIp11m3WxC
VbAI8rz/e2OgK6J2Ta9KwuhAJEBvyUUuMny25hohKfqUAExiVyrvpzCAP80lwoLV4RTAVBhPIhix
qj8RwxSFXyNUNVG3U+YxCMSzZZHjwunK3mtd9dp2A0enYz1WxX+i1qz9udyXAIQob+cdMGyOt1No
jM3izJYt272a0BA3CI4UmwHltjRTAsZr7uC6ACXmsxk7tNEYHZdeYaIXpl5GNrYwRuq4Eo6IFgQd
ffCU1aGObC6zSXLRM0MQOzFJpTREJfx7XyZv2BmxXWR5PyYpOfobdy80hD/APFjfksoVrSJFeKWw
QP1/AlWwIzb7oPpkpBf85QpGN9FIc/m6PyLSqefIkodDDpRyshYq2nz96mVHauiEG5zmsOktucVY
pyeAUBtBAOVdj3ohM2Nkdx2h5ByWDzu7QfNdp7vEaVfVthJb2KkQhOkeJGsyjeyAAmQqf1jQ2J9s
17BNxpwcIkyk2pvDGc9ZuAGGnBXscSeMHEavt/MmTrZmMLvNEngoY2D2jqsC/915DmUqxr7KR3ST
DLjjKxyJg0091ZalY5TeCBP7E/ZbHu/TRlBXlPI147AV3uyWBKsUhkQthGyiEZSckZ3y2DoO+EQI
5KDvgNXLMHDBWfoQEo6Zj55yXwZRzxF3q3058ju9ctEHwmJE10qudzHKqa2b/QPZcKsK3hCp4dmD
ENsMc7Stt/agoRM2/M4Zd+fQG7X4J4A2cr4rLmo6eWg8lt2S0QvnCHJDq4gzo4Vm8x7URq5y3OKI
RlP5H9z0SBGGIXO2dCsBZBA4xgKbkUD1sY8DKW6AyGk2XEEgqSuNu55uujSOeP7+ndWNSVLlN1JE
2gC6W77wuK8RtP9UIHb9zAZrIKXkZYFn36F+iUWSm6KBlHztpyQmTIBCg8sNHNhtp6NUyl5yOmGI
nAMi4Lzy8aR/oIWt6J4p/ALwC/yvKKBWOMtcGaEmtjJpV0u7yOPwTrp9hs7V4wchybuGxr7kJbEA
cJChDOI68SDXavNa3bkbxnJTXHoGtemT8taFtztrt/7hTqJusLoiqsqgrU3yps/lmURGldaRtACj
MLHclD6Axv53mgyMjx+dv9nB8DCFPOCyALGY9iZ3P5aIlnQwIMbuY4xz83+DDW2zV3Gtrvs9bg8P
FnZP71sRirG8Xo+g+rm8beGGcz/87q2h9/usmusO2lg+Z1EissY4BsF7BgV7btVgTPB9EgyC2OPR
T5YCZK4wk881qh0j67uwQSyabTX4DUHe05JxbuskyrgdfUwp154EruMdi6H0APOiNRratDJG/v7M
OH1QMvuEe0iu8WpQhAZNazgwpFGciK7kn128h95c7gSWielNSpJ012Y2Ffv900N/HX/yB5wue3Li
ZZsS4o3By0HgocvM54h2pLqFCr2PALk4YK3RlRZes20zJfUpEbqQDISnrFoDs0WDYjz54KNDuFVi
vgXAf3gadxe95Q7sB+D2hJ8/g2YhnOjpo74HV7Hb/EGmqFwWsKI3N+Bb6S5qvfJvF1XjAZGtUyiS
rj5OWrBOItTYv0Fvpe84NA1CabAW95BvSWA/6uUsGq4okc83V5yv/HBPwiC2ez/m7Oqz2aBMYUzE
NVu7D14GZ/POEK3+B8s60kFOX8G7lY9EmtUJsG8iZzOVlv9vFYvtriGWGYH4d2atBzX3oUPjFo62
M/BgvBKGOS35QNHkoUDUP6R8xAK3Hw2TEznGRrP5qm13krwirqX2jA8sU5zlcg5JL2gqbRZGHf9A
gBtT5tUJc+zAwO4FTKF298jnAHjU+esu9/IzBTII0hd5ScQSNYoXdgWBu9VYGRq/kMfA3w5nGxEo
lKoLHbCmbXKj9AwQWwishhDj9gMPYd/5niArh4u3Prkdpj8XOU40+UmxY3LE9jcZSzlJbpk/vI0+
KePePAdCLK52NHgrBrDWoIQrPQvkSYUqkSPKGBl7bRJe7/wNSO2FAnDOBZeFzbGOdnAOv8pSjsT/
1mMa8EJfDpqkgaZ87SpHsbwY44VTLOCNQtGbzkyqo/fc6ycPIq8K/n+kMHgdXOKXGUcbFm4FYoWB
DXeo3SGNZTVEunVxxBWg2GE8TerYQiEHlwDT16V8hytQ+FPJzDBNoWKGOi4FKgak2fBtrCV+aGLC
re/7eyGgmqyY6SECA1Zhb9Ubwrbjl1KvMbeD8x68ENr6GiPQ6sqwUi+H8r+GENFgNZJ0HmWAPj6m
2gjBaq/QEnsW6nK6jMBV3kZhmaQBWwURPTpVjCzsbohBoH3pSPbacSiJQTvz3Ut0OB7pUen62z40
UkAWEiHBin2HG0KqXrsSPwdcB6ubPRkxJ6KvuJVQ/Bgazz9J9oli+L7Sw+w5GXPvl5IEoxx9Kc/Y
h8hFsyI9BE/IxHxOWI6iHYYDr4rZ1ejGhYnXC+p3x3eIszn9+xkitToCO59hsAJCUmoTSJVOsmHT
7EsAIScRMRs8Uueyf2AUFlwlHWZbVSHtwzceBX+qeFJ8oGt1n1kqEq5P2PrnEuGsuCfC9JPPskfe
pTFl1XmY7owXjiypKh89/906nRwF2ghiInH+o1OubtjkjxwDQab6mcCTuZ+qVRlcRp9eDOeumbd1
9uUwAlrV7SEH9Zept3+gg4eKjw+JFivhnMGIjYULS4fLDxm4DwNFgpnLwKyP/ET4YTL7RdKRSIE3
dcppFJh9ERDZioOUOBSYy6QgPp0rh3gmadfPWH6NpU+kZHrhPFaFEnETgK+q3OozQU0XcWaw3a6T
UyRtP5H3Bqu+hivCcoGq7BrKyfwbS3jrxjdBlCOGkZg1NXTmiO8LrYM1ddC3/cBSl8pO2qAeRkwS
sq2Xg2ZGpG7S8amLAIgpW+scyPHYOt3FUdFK3LxQfGgb+EuO/Dkx8oRK79Z6j6oMkQuWNOo7KLJh
VJMXDqqQHJWGNXibf/ni0QauscTJUpHEfbWFoNQm2P+OGvOT8VYa0WLCQYwVFgxeyMlp2QseO9a7
8HG6yB77WltksWba5jsPYxWBD4tfP9cdip4FV67cW+UtDp1i1g7e9z+WK9tH8RBsO7MiO7cVOJaT
0nNQd5u74BnnCTTzEdGcTtD2CnmkwDrVZIg5Xcq7VKxEeRJHtuhl4x8GMvfLTMXLr7fjE5mrTQ4J
4lk08NIfMEqDZHQvMDlLBk5G7zyjN+qT7mTc4E0DoC4Fu1qcexvbBaCGGEXr/gtRC9aM9sP/Pmxh
F62D9SlbDTRTq4bOgBWe7dcWyaYR6DAjHjU5P2vAK8zKqgxhEmLADReuM0Acov0UqAv4rlSl7muW
ZXdRZMjg0WKyqIKht9A4d4pAfJK2dLalsrWWUr7C3SqT/8l5ONnQy23F5svP0WpwqotRcn6sCZtB
H36RVSv7/5XOeyM3XJUKmJC2/1NkHLSsn/36fpnc55CtcEy0Qnbp/rmCAhylWha7niPV1TffNO8I
lkg7Ouy1/iCr/KqN3mPrG2b6BG3XtwBakOrxzY2dAQbBH8vk/shHJZq3cxAX04S+JeeVtjD+gw47
b8BF2E5G2zH0r63y/toENOYVskiEeqW4RYOTPpUxtdluceEEm+5dvRzxYi2vadU8kXqYMznAI8V3
gan/9xche0XmUF5lB4TBB6PRt/5noNBJvGAFQ3tPbkaeZotkdhQegNWGkEODGOTchoVZSYf746r2
VC1BhXKV4F7TgYs08vcgSpL9+I/Wf4cKZMPs88HoNCokZPTRdAVGBq/gSPW2Ayy18vrmZjzgKSEo
B0gICK8wrzQse4A3IsCX26w0iPmAwL6TmYT4UIZss2V5HRJnjxmFjO7835ebLsntAGZYD0XE+6Y0
gQxxyFOtUWAx2ydJfeOWl7IbXmW+mOZpdfxkY9xjpWleliN1swn13YvbKYnD2DRzZnikaNSlx6Js
lQUj65CN5+enk2Ai7F1a33kc/iPlUrAMCTbc2gMrUGBFYWwQjphTvRaCZz+kcgxxDYt8tUCyuPpk
VaUtF6dJ/FsiforNow4BkPCE35HKU2WDJ5+WdmJjtm++y07T75ikpzgoVgHyLu6G/ADkthFkgrKF
97h2ngGVO5zJXpVADOCCqOFxg2POgQVm0l9cUApXf8AR8cmttrMq5K3WfwGo4HFP4ZFNbBR592E0
T6/uYqAYhK6yav9EeHyE7wF2iOn/BCAWvwhNTTWd8PQIPTpLoRatBUMUdHSfV7ogRyaZiyGH888p
jiP+P2D93m/s0/jrxo/54yvoPrMKu0amlMUsHDU3fUJ+2RhXPlUOdTAyzv/nTMhE09w6SBG98D6q
TSjYpxH0LVH0ByUEEYNC1dZMEASwfMW/phDhSrXXCb/6UsQoF500dRrgAOiXTyPTqc1eW/UHPgS3
nX7ipdLU6U+nyaWL4dT9uaWU2yB0WLLWcF1ONQ+FJQL7S318L33kVVu1eHTBz+4zIZG+QvwpHmsY
3NE7ZA46Z1AAvBKgifTm+VUKr3Zd+6z/UB6YUaQQkp5DzEgU5Zy6yKR+CTVp4lDjT17hQWL7nu3Z
hbgIthW/9XRFthRCkYw3C+bO47l8k8D0P+uGOw0nG2Q++VBriRs5FfQkM4MyQfn1sUZQNXJDqWSm
F1Zo/d2lxV7VDr5K0KsEJ/fXGpGt0vD6u8FoJ1ZyqKgEouxMDMIQHnZhv6ViYr0zg2748np/hkv4
q9rh45jCWURqKxnIQsGrpumEZ7OhnXMV9rgveOZIxUh/0E0C3LJcSO9ThMsypcvLVJGLabXAbVhM
Tb8WZqYr1Buh6Flm68YUblHY37jKXF03UEZ+KS+nzAXKhsQ5/xjbSqqY6e6qBGu3dtL7A7m52ouu
v5kE1iKEkLYE1TvQf/4g4jyPMDqzrwLj27BmF4ZMYAtvLodWIU5XTqTlxf5s74GxpkjZHFvsLcNG
7RdNVZAztv2sxxNQx7AQtMAmzVy2hKHyXVpLYsmsddZPK/+/YyvTq0DKhirqnItN/A7rbhk7XSUm
gJ7Z4Y2ydGERrytLm+b+gQBVjXPMxDphzj/QS8kMXLx008gyZVRjsFFwe5xqkMDUc0DfalMVUMH9
B0HJQQ4EN+lS6cOevy9YVgx9y7zc4qnYAEpP1jJYX67QnTBnGcTnkIaNdS7XoNdLbzocqozciGLq
rclEMrxaLTAMTaRr0vyj5JOP1Ggbu1An6GfiUAQm2IWJxNsQdTU+41U7aPbHBVd1S0A7dNkwrax9
43m46NSAWeWlzNTnEgkKE7C5kgdPAPc1e4dFHfiG/OFGbAU7yfzF3301L5SRVYhPa3DFzTO/aTdk
axiMzf0Pk2MMs5ADbVl9hQ1d2VvOcr31TpZF7zhafHhFrWbmG4wi2tBIozj5SvL/Ah8IimGxClB9
P6oCxVF4M9wPGHYYYaWiRFTFF9UF1edEd9uHXLPPmmbBn+y8nzVDlQFlwUcDIfIA0IYjJsMH1j21
QMUfJmEEjvoPDPoeSKN5E4My4Fpjh05YHE9v/qqhVY3ZaSVy2WOJdJeP536YWesVHOkpxnkXjg7Z
1yQSx54+/jwYLPgQSVBozFj5pEerwaDOyoFrosioWV+4lX/nuThkxv2hUgz89VdYYTpQPuNzR+Di
BQm9G7aM+fPAc9SkcQxlxOpIJ2MLjLDDAW52yx/b753kdGWEGO1NIOoeaFTKZACWIlooFZnQI89Y
VRmbcUf/6oiHEYhSzEIYvTMRFfA33Jpq+hVFJcBrfilH4ZzJx2OdzguxBw37bX+ebVycmA==
`pragma protect end_protected

// 
