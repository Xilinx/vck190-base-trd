/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Fgcvq9yodAEyu7zsWWZ7LwHLqer2uRdIROgj+b6me/wmyj6mu+r4+a1EPBMoGlf2Rxb0wqrGm/yl
7FT0a+0gf6RIUa901Ug60cEq5l3MsNjnNX0EuQ9QHnbWnPHO5sk3W38XYr3s1DoIymcMyzWSb3j7
DAgt+R0iGXGbLJHe2UuAgwrybNhjpWacbybFOYZoLu5Z50wmOHt3p6J+gVbTwfuHK/f+KnS4VtSD
EJxx9+hQNEvkukNe5IcvkATvsJ495o97/SdF6+o/UvTHUZ0m3la3MPtrbbqjxbRc5d/SBaUYwJ/0
DSKgI3IBXs0nO4MGwCQX4Cy0xa1KtNy17Uqy4A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="YyF30NSJW4xBU1bz6CmJ7uDDg1utz4oEiyNQAWYk7H4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52624)
`pragma protect data_block
3JkMrY1IEAXvStruy6C+3vwvHqbalen/63me1McNKlT/ojlQBwJPVLe1rES12+1Zb920Ow5cEwf3
QcMXy4AAlUy+98HkSpR07lRSvmaVa9qWcWAzos7oapX+0NKUmikKUf8XnmvJTba6G5ezC5z4BOQY
qU7upcW9gr/vhUMsXfCAFteb7LidJm7XAapQe3wCFuw80VukcqacNSYFk6xZ9x5VmlM3MVuPvYoH
NuqOgcJlpP/YR8oRYJbQXPTvGBpqsqJ8d1vl/t8Hw9OgOiSf1jmV2+ZjRghCAYGhh7HqxM+3xDI6
GAYk+ga/zw9M8sWFrHMe4gwBTmaUlQkjaOxeR67VHBMDyqAJFmqF6MZNWKdj8Jclpbc4T5NzdCXo
Dha8Cq4YDLsqizqgqPX8vHfmxRjTFCH9TP5UXNxJOz8Luq8jGbblhepPzCLQeOcYNIuDrS4zSt4R
/Q+6qCgEEZQZ8T/a3U6XUyO7fGHl1fTfBZIHK7vd11gYbp5QglJPkpHdrsQ7SInnvWwVJsK+Nq1C
FqKIh5LEEH8lxgIIy4vVwZivpHaMNpPxaGc1A08NaPEt8Dcz/8R0YGaEehpZ4PlcHM6wE5l+5uoP
XH+r/+fKcMXlh4/7pSiFELN+cw9nz9F7Jc92HqMZ0P8I9yUgqCMF4mpstgIlxhECNKtHwKifbSOS
VvOz5+41/BksQjEcSVrMz0YtkWTuTtoEuCjaFxFikUruZlyV2bwn1icYmybvnL3bjpLK//qDoRzD
8AL0DSSMOKA5qqz4hJdHQoS+UmmUmMp+RAY4ayVuEH5ANUjx+FPhkktpp5KEfLinl/xwlFJc52Vm
OpcbEQ3tNuSx4Hzf955MSYqQR1jek+VACsYROHASrQePUIENrAQYQ/jIfzdNUeurwTFcSQc9hBIs
uV7doRwgYkXOzNf2U3s40wuk6JvYNaBzFeSw88OzV2//bfdXZ4N9L9yo0gav8nXRZyz/sTH4MSDG
m6UrUHki0V9Ox47HTk0owoHyULNS5EwbLY1I4/zUYtyVajH41peaOKXUThwZ/JyjMu4f0B29PBpA
uaJUF8m5pu5Gd3cQ8vG/d63YrgP0WMGtw17Q0dkIsh+4SBT38IgpMg9lCyiIAEPnDjB6HJbrgG5X
/OoujkjVmDcC4NxRpvLQeRNiXYM1vE4vNhjAVC9+AqBWXtFXXLTHkQA9h1Ku08lqUC0YVhrFG/pL
YByp3Xs3exoKVfZ5XJ03lHk9RgMd11B0YJA/AjoQVf0Wu1PNc9+JWSShAST0mS5vw+YZ7FfbtvTX
mwWIZG6E7ANsSTeZ3WH8WNIOGv3e3ftdadN9bLmCJwm8sDLrsArgWFZKIJOv0ggVRhHyXgVCyYXi
Hb1XiZMxqjv53uHliPnqLKbho0Jtwc5xXwDZE5PTuVTAGGva6mLdrqqlMWB/QG1I/tHJFKZ511gD
df6sNkytiO2nLUp+9cOJp9WpTCCxdtHBvpzhZX0JGSOP9kwkWuy20VFbcA2EOVlMdOaMkLF5RtSf
rVWLVNX3v0lezFjxYChtWVmNbqmtROLZX0q1z9OclgGE6DPdQtYkto6tmzMZ8YsOTxbNUBaN+NLJ
XgLTxfMsDrgxPIdUPTuiC9UgNWZDaS8V33cDrJlBEKiFwXkyhIlH/6su0UrQQLSmXSMhBAXauj8N
kg8pKiDDB80kWpU4Ep7BToa8hgb0Y36dy/43VKBlBjhab0WCTc7okgiGcUYBjdqJ1UlVK7hkefMU
5iSpKawPQJGPYALH2rhsa9Q/BrUX9lk0xVzYIczW/dHKPpIY5r870s1bJcPgtKJ2bqrJzOvVDY6z
XGA7HzhPZ1hX5Z3rRT99M9izLhw6EBBLDUbIxu+Nbo88xc10gLYHf4nGCNq3Njjo2BxQdO7LEwl9
bJ/ssrxAAi31Yq8QnFH6O43EMbf2hNkMd0LKvwgovYYt2YWGeg/kcIJ292VvuEy4gDwnSGl/7uH/
61XWzknJnw6ZAxbPrxoqopAkNWZwlF3W0FNKx8U7ezeX/CofDxubs4cM6edVSE/lzDBtlRqsfMJ9
J1iTDTG2twM0ARf82jHNQxTpPPP2Ws0UITLPehn6WSi/4ZhQSwTJ8vfMj4z4O1wNyq+vF4PgUJSL
a47gIeUhfEOEXYFpM792HCkhprfrz6mjFVmVQeQ+BHJEuXRle3+NFzCrDnH7BrPr4U6+BbcjpKst
jBSsqqoP8lNAQ3Hhcl0iwIlnnbGeQL8GIWQbqGi+qFaKcF3kdpHRQiEnV1S151FN3EqBX3OmwCeX
gyKxMsFWnPJWWxxEYFrlQRnKAKcLGqsXHM1VFlUIpYQhKmT0VzpdlLSA43deNpyua5hZmS+ehppW
Wb6kfzUIh1hA9E/XCoDUrpRV7q2j3oUYBh7IohFCKgifrz+rN15QukzkGs71vfrfGwZpsd39n3aq
QkGRIlEKMkokct4Ks7ULMEt0Nlk2Mz8JX5vTLYDMNkTxkBoNqGQ3fJG6E+oRfsLS5z7BxS77iblP
1Ln/Nx5Xzl+4fzf18iNkRt74ajWdbG7kkEvZyUn9PiXFEwHtOomJU6DsXfu1scTy2oqlfS8YjHTy
5hAkgiLAzQssKwIiJNszhj1C5J0sWUzHkKGaHKJE2lqNO7e6AKCqkpLckBpZEH6Qsb9X89NEMyWE
HxGdR/1RM8Lwq1azrVLDedVkqpSQg9M28fA9mH77RPPwNE+SoQxVzKDZLAust+oeslLaKD9yofmR
gLW5QeavxpXa2z0M4O+Ggm3FJ9KApThzXObFCZ+Fhturp+w7xloq2yVwaPF0+absHSyFgb/804a0
YeWvZ73Pzi1jXFjHAM7kV9MdfqO4aU4wzwMGL2eOV93lakLTHvMQIF5RV4p7/A8GYfGw43jz5cfo
Q9UXsH/omvET5cizVpKwEjA4q9zCOC1fl2fyeWlr3uyjtEJ368qmwQnhN0HAUW2lK9UJJzf9qyms
klA50SXBiWojzATJRNzhDwXQgS5FVjeCWuxqcQJT2y81ZC+Qngz5P6OoqDNZRZwy3rFTtlM0SgtH
a0uTk/r8AGQSvK8DtaNLZzCJeZW2yDSRHufwyT0ibQ6kHzk7EdQrMJJ4Hwz6US1WHpDzA2YlBP/2
gsMbwPMcD9EaKiYGiBlm3uwiYLDjfguB+9tXshkA8mgJnWRvxKgB0j4MWzv7RLb/Lky6EMOzgsAb
kH5v5vaxyMj6sOeWjUa7c4XFcKT/jzIJOg0zLz9NENqFVH/S2ZRu+xBHKSuGn4Mvg5tRZoSJK57v
jjotDxCNhyd9K+2Q0M7ffjlPGMw5GeAfwn9620GP0gl/GEebgepBbN5HjTYKF+z/7cShGUChSytp
4GtpYSgu+DFoAspdaw3y+aWMsspN3vqt5BdvB2+2G7plZcNuTZZ2vC3LHp0fT9MjJ1J9UkxOJ+Lp
ouO2SkbF+7SeWHYdIonUvchCNXC01d/dPbKldjAHlbIcYWuh0/r7XhKZDRU1FCodVLwe5RBnGoSG
1nV+qiOZjOwA59iuqS7gROhs22MZ7jAsRfaxNuGirQQPlS7ejUPMlydPoaN2jBzg6VSc4bowmCLD
WLfIl1xLqF7vH2/zoQrgxMgVNLfqMBjidP8rbyCqSESSVWxbjSGXImXwUCKCOlpIK5ynauOKAXBa
LGN2g4buVru9ru9vE2IAf+4iqOLNSUU5tadO0ZZA0/w98l/uCu392/0BGhZ1CEmoh2tT1/+jJz2a
IZSVV046DUD2TwBYKrkesAAFsOiSPLvv1klpUhu3zKYOEbRMTfjDlxgcz6dn2H0Cdp8loeQOCO8J
ISDF6qcPccNhLkHe31xpfBmQgWekz9WMyDAvwjFwy7mCJqjtMmCMCR9sXe6gmPs+3xGgzNK/iP0Z
f9CknO7QhNW/tB2btw/MpETC2n6d80P58VvRF4w998qa2t0aNHcalj7IAUccZY8N0gBMhgP0ODQz
r2C7NFHAxjgwE+lXORxvpslfZ2lbtV4CA8+JqV2cd1Em7sOj+Q7Dr8xpPHm69MFlvVkBLHth5Lah
PDGHytE5T9JFj4ud8T4mzIui6Eb1hBqY3x0I2i1VVbbSpAxEOM01dbK5vO4zp04y2qIuHrHZEWK2
TAEnEPZyWUKTk6te6XrmUWjczyTSMuVIQs5ljlWnVmCBF5OaI5WhmnUiniWcnj70KLx1Tfc+U5jT
C5SquTlIiC66oEtX23XVxyp2DSEknlJHnsMJBpYQoWoIn7SqekCxY0D36OS+bEqqo4EnV5V0tDA1
zM4mbxG0QJ5FGAzs6MNIyYwpS83i/sphYWjbSoJrlrRWpDfiK4i6HbGmdDxUZ76KFd4TG37J2DwL
FFlbVgMySA5RJUJLrg6EhvDDUXNSav+6f08pd0BXc9KOdwpx+af+O0AzkmKthV8lYNOX+p8l6Jpj
N7ZVOpsNKf6ksHNl73+ekVVeHPr2TfyM3tPyA8HgSC9tZP0Ey1jVbYAdL8K1FEGLjVQAX68ZVEP5
y02QhP44fpZdWxM02K6pU0kKCkomFbxmZLBpT5nFQtYiT8JuGE06DPCWBCXJYy2RkwIGn3mMwl4t
PQqovcrRQG7XrG+Ia9gJMNviilpRTKbqLqV+/HjCLtFn+YKJF7cEDWr3j5pe7sxC+FO20FVk6AXh
PkvdRmL4lC1z8fqXHtQssn74oR26G3CblaG2OC+I5UXJrHRoCXb4KgK65SgaYDkn9qDBUYsz9EJZ
1v7gWLLS81EGMeLAXpqNIJPEObNdPEjEl+G+KwxD1LqSZ7Xd9VppC01UcbRvO5JWGf7m6KdIjUK3
EgURMPdaiUza3TKG7L8atRbPc4H0xxLIWhWax+IBPS3cwNO9PDM0xsfoXLTG+w/vHoqiAZJzImQV
sZD+e/8lCo/zpah5KUcemXm5YNUm+AYLUXdvx8OaLHaS3Uj10LPwrY0Nk1wGFCyOsAElIYe9Mz5v
yKB4eEj8Y0hdJJB7VnuwyeDy9h5NFpX8TaZi8nERbByh531WECZkXZ8leZLEyaXu7eEkHk3cjgfK
1ANTvNZfZS5+DunyBuRNbbjiOQaHyZGGF1TwyA2Cf7FOtpXSbLXeMrgb7SITV6Fn5qptFwOPz9Km
JAGjEQIuJxR4OGmg+3HHFAg0OZSd2oJMFbgvGc5Um/HftpWjQuD1eu2UwaOCGoKYH8SE8ko9tz6Y
t56lAeZDArEkutQRczukYcMUpDvzI2GxhK9bHHNWULYN/yttSwXqpx9bAKHKDJUvPcaYanG9JpUl
zomnON3PsDK1+pc1DNn4wpDoht9mJYgBZ5hyRhVbIIlS++BMGtAQJYTtA48HHi4Yl+nmKnUUdQRo
Rad4aDfRb/rQC2Rcy3L66tZytMTckCUIBlbsU8CVi4ncbCElHCIe7AM/neG8zc1Q/rB71qB5h8hk
fS4bvvYjt4WeiQz3JU+iBiIpw02dh1QiQPWL6adTzP8L1lvY+8zFXU3VRMwxREkFeD6PWEYCG1+Q
6sy6ZfsK8H1Vy8wqryI/uSxekKHUWAJ1SJPRWmyytqkI1inh4eP8dPB8KyKJlPmJWMoFKCTNXlYi
5CmzvBskWzO6PfE3I41VVHpUne+6ZYWkvfd0QqcJXfNy7T7766ZWT/Cg2SLva6Rc/AwiAkll/exZ
lxNiYPdBEdQBhfJ8epmQ5paUTVpv9KJ+q4mKfZP1ccJuvxpHtPj5hfB6ABG1zcrMIxBGHwsnmktk
w14syAxto5D2vyau9toyS4+5KZMkmgEB+TI+sjElX6haOMXwgl9J127+b6er7KsajStAx49cOHsE
e6soHBkW31Ibgv7uiW7usPLmPLscCwz0NYhdFlQvDIsSBpZpaSRxYbdzv1lwLWF3B4+xxNtT82xR
vjLb89yeiUUY57iKvrJb8mHhcD9WP97szF+nW3yeLroLDsxbSv1bGOuXkzoYa6MK/SiDP6ypUuXs
R0l4oXFG1kr1LW2oVeXfNh0ZyJCu8OZIxp3tQ9MlF3YOFX87juJVaGL1ADWi/xd/cOfw1fxO0Dis
Ejl7b6n2PgBze/QwAbDxgeYBPi4W8fns7e55v0QwewnzlZ4voxZV9uIsCY1TcvjqOchHDiguwuog
cpCpadjpxYV2YIw629WSjgCUUTddROleQOqJZRggVNSfLJdYK3oWvqBiS03wtEeK1ELFt37wjy89
1tswkMPwwpX+lTtMoUNtzZu8M4nJddsMeizMWzAZAk3Mkxw9sTP6pOEy7kZJu3xgaUat7FzT5FWE
cVpMOOdOvPUNagJiezPkonnhIx5z+WLPYsAo8XGsDHeIymCbIvSDcsTlxkQpPy3kGyUDX64/kQjx
Xvxyj7my/kUTE5JcHOxfAODZUazNhh++KWUCcJo0Ughh+lyoCLQMCTkbIMPjHsX5DyX6jVI555Nk
qdtysvNizHCMqamrYiWBqKZ4f/pnlniWU222WmINRFQR8Zzh4Z9WUnh4bL0oR7Q/AoS+GAvE2jSq
PvyM+R9+r9fQpgxzxORY/u065z54zEeybp/3W2oEi5YrcVWynVVDxXB6S9qxtlCTuJoaXaf1QjVc
J1HKtcQH3XAzggOmBthBoOA+ml3okklT+86oARUy1aRq3c//NUU28d4jk64OxeXxNZRhzAZoiy7g
6t3ZjRdse3eJ5Zos9aYz2xqBCcqfJGF8c2rxl17Kkhc0ynC1m98olon4hbvCk5xAZHJ1ayNmLSGO
nj6R1F+ZkeTKnh4absQ3tDbUdZvcvPyBUxvO1xuYO5jRjq46rmV8oK6a84yWrdbmuHXLtVJtdvgb
s94CNt9T1kwkE5bSnY9xu120npuma+vWwh0lrPM+qIiLKmMr5ABo4bV9gg5InWNZlSwQdATfpMKm
pihnMWyWiIy+yEFqi4mSPyBA41Y0My/7DAtQBbdiwsnzRvbMY56kB8MjxY/BAOv3yXEIHb/p6c9f
8ASyuuZTAnnfatOD0QBqfAe1oTGEZahm/xRgRAeEhMLLSFpS5M+9rUG2H4trTd/rTjXORkajNxQl
1xZS6q5I2dFafB+xGrcx3VV6Bfon58wVqfqsduJRgMJrFfsH1j+yqX9xks2N8l+F4UZQdrgthJ9/
KP2EbzOAAWFhnUFf7pSEehBjDZYztQ9QVQu8F20mKELvVQBjAgfDUolPF+iGK/phqR9+8xxuy2j+
se7aqthHPnthvxkjiCKOTMtSyV7iGYxbLxgvl1lmHk+j/nCGuKqozfN4DErmq65g0xQ54qLtdEJ2
qJ6USLwBBvAjHpUQSEo1ie+1gZcnVFPVY4UghvMnu/PadZWFnKK84No8Td7Vp0SxxEJUU7wMDw+R
65XcT2kMTgNBa7fZB5bZFIB9z8avLF090ILiMtfGy7YXXUA2My5oNqWCTjFPOEcfzpNaNh/mq9T7
HgiJF/TZg/uChLPijWQ9iD6NQpteDzV/MIcTVDyvpMC8rwjaZ3aCzwlD1mZRE5+TZ4yrDjeCt4tf
wNqEWmZKzYmJB+di5kXfbZnYG5bF2XIkG2LjOt1tEcUAhyd1Ds5ldu0G05+LMeCK0VucuLovXiQf
fq6SqKtOV/SHvbMhVKVL/X0nxRuirjIe3hPQOuviQWELohkQ6T7PxMpuwzCh8FHKV3wEOmapzcsE
f7HxHED+gRdjokgSBsf5Rl6p33iN9qFVfkag+89/Hdz9CZid1i7SWmAax3R9sni0uU7wKd4lXzfv
IlXKxKUTZpLeukPM1vsuHMBs11/hhb9SdN1juoCxLm+fuyJJTnpNqgXGTbQAY07SAFINuxwM4OyY
kK1Tf4sML54ZZ4IBDtQFUu+YdHVrAYnF6OeIfqOIeumQHsGNa/Y8IbW4p5MAgT/1yqO379qRGEIR
zZGrFeW3iQpTvRC7vgYN9nj3hHaM9g5OQ0bdZJEz0iS0qxBdS3Xf0mw9mkbQpXoPxxHGr+6vz3ow
5TclBIBd2096Dhx0h2uPNSh3CaZDA4eqOHOltAW4B+TJGjPOkwMYwZfjwXEuf73ytjCfPwoFLzDC
2oMK5jugGpUik0aGY8kzTkwxBMwTnL3AuVpv19H6EY5X7/Ogs8rNetRyPMfTDLFbemqMZhQ0pWLM
G0I2YtC8GVNakjAmMqe6ThhxRBXZbDGOHtNz9AJ1JfHPLEdKlSbsqNfSFgdLEajr1CdaxmecGgHU
SJb2ffmb3QHo5PfXfnPbCweviaBtvXzLcoaS+prg3GiIkCkJUI6eyCbdpAeB28TFNzFyPF3Wjau1
t92Y0wH6yEjOg8ZPJb0VM+OSRPpHcIdCaNBRv5Hs25pPp6pMB0BmoAyqQ/RZgC08WhWCDCtbdgCu
NdF1BDxeVstIXBePRXagVdOcaA8ENoVBB5EOcKfmEX8fB/DhGqhjl+l36m4mOADrUSBBHRjdrLlz
WGWTy4FlOCz+XOTQDcQ+DmXPqLSHGey6V0jRZE6evzsvDdJU62M1lyTV54isFghBLskxXvFzdjR/
mrXayTowgcnTB8ewzNVwXaqfqYIaCFYv6hRDIko5QKBmnwt8QAzD8S2U8VL9FOwrZyGDhwOugT38
DQCMlPvmHXv2uSc6p6geD7xqOR0e/4g8EnDQR6GXvsAe7gKZBiDwk8m6aEdGTy0GZl9Nr1ufMObE
USYXsc23IOhauL6+WnUW6cqsemM0+I3L9a9aIOHHlGCzB2pC3ImlCdI3Xd0LSVRzoa+kPjxsxaz/
mkPXF5RhLtG037+YRRDLSL3ihhUzxBwieYdpsLVngQgyJJSmng5K315JuuQ3B8lmay1/pDnsGHEs
59DKnOR6MCChSc5J7b9rrEZLIBZouk5sAht2ItHBdvalQoJ94F+vW14Bl69LpMcMc9kKBlLvHYUi
hN7fhfSrmn1QK1MAbZOO0Rq4IQKC6Wvma/7zQlmg73Q97YirOH46di3KMKbmotgMTPvKcd2SE7Up
UoZ9rpDaxvW4pjy8FUN+v6IHEJsrxawbSKS0lf3FYCCHO+FP6dmrSb4pygDxqvlLrTYhbKLoxLb0
xIGlmBuJzNfB5+oJ4vZ401hraBiHpyBlrd7PbKT2D0T+RHkSPJgh05Ms6JVF9gl+ilmWCIdBY5VG
nfp/YwpKjW7cQ4OwBIgbyef8MYSYINnmz6iUg+AQZ8YOl7cENzQGVw30sEWudTUHd2xk2yLhNjyf
PaLN86Zus6zSAo52K5hojDCcHOSFgEhBJuyT2RPUjZ9Tu7+ybpI7pSBEXPK8oInmAKxyNsaCBXeY
44oqiTJNFLpPvE1yxR+RUFprPSJkbf7jBLl0ovbAQB35/6zagGZoi+12o9fR9drwtgMXsBjhYOoP
ZO3Lv6uYFuekpDygNEAFRy/J23CCGMyhgL3gTyJ+Klw1DQuxTqI1xw8Ic03VCZN2cWZ7Pq6XCXrZ
fpy0tkQasYkOgx6ye7dFs2+V6ANzrzEAfOpxZ8ZcJYv9Nbi1pJ/HJs8/PsZkwkxS18fOhYPMHOdo
m2GnQji86sywEteaHDbDv9+0xZsx6gIS6O2Q3pU0pr4FRaBBvTYkrwNn91EPNC9U8gQMvFw8SueQ
imvgNhrnacFaQhzbBjtWPt2wPDPhim8LuXXixCPVW0/PwQNbeibURv2DQtEeX17s+gDmiec+el+2
bWVydcjvraJw6UWgN+i6DPTBVu65+Jki5IkSRmdg1xrmZdar0mTa/EVA/Zb5JY39Jq592+db56MY
hvOk+o7wK7yD4BAV2rVf5jdEX65Y49/vE4e4sE4HEbVv7gvY6bbdJ2bxH4BuvGv94kRv5E6Bstpu
niLVK8GVg2N7u2b2Pe8XilPQfk8l7HaEBpAUp47AZ9aDLJwf1j3rGJqCSvOdO2i6uVVjeWmUIj7r
TZzeOTRjfOIFYEeAQcBuNHuuuaTNfmLgopZH09fGo/8IM9QhWmwW1ZV34GgPArhIxPwn0ru2XuHV
Q3qzCuAruiZ7W7vYU+Tr52S7W6zStOXhlh3cD2oEMbpR2W/JE+3NVQtliTvCh2DLVlGPqoCJqXBG
RvWHy82WrR++R0fuMOwgJ/ew9WuAbbTShKLIGeRYHv/m8SDN8MFFd5His/O5TTJ2kVMexN1io+Ks
8LU5oS1wvuD3JXgRGrZcX6qpkj7m+LAW0+Wfl9Ou46WrsasML0byzeYYSMXKRbfTq869GBmGQNyL
Imfk0e7jmMsxEK8SCR5rMPQHzjxRirNTh37Lruc4ffF90IHrXyZvmh8DY33pbeknqFqd7x0aey/o
pP64lUsEGNsbVa2Vg0K9N4gDl/P5ZmXsCiDusO2eBJ7OiE7wK3m+s8aechLrVU40+PYy8HNUg+Si
CSB/bSler6BhwY7e+FmOAhHHi1n3mSSOUUifEmWW6SIu9OK4HBRC/w1Cg0N2UXei08Yyf+Gtz40X
qbgKqNrzlL1MjwKxduIbWi2zX7zxo8tt7dckd2lDUtUcS4OcN7J45m+5BI1vbQBVFGHgjVS8LLjx
hiRVdA+v+FSZ7ReDSuBYxnw8Sn78aRA14wI+5UT25KxVJQPkBQ6FjzKbfiUN3yc5WwsOr67pa3fG
fTwnkfvg/TaX1NaKtt4LoQ9R4R8QFUgm0AqufIa3UfG7myPGCyiRlvM4wMlsHLusBw8Ku3MdND4R
Zhi5AKZq80L6grWqhhF42l7coJu0Oj1Q6aYmoT9MEDhulZdsfOFVK/Pgj+bVqzAqLW+rrGlLkwAw
AP11aMuPMGee4eS9d8MaxpkirO8EwmgOpOUojiwZChP6ie7SA7RReAqD4KYQlr8iKg4zKvbE0S7U
42tyDtFbVMxUuGBXBKQFJ8NV7EgcHE2Ai6LNzxDKPkhs7Lg7XZX4uJ8RBKBAkkhGf+5ei0Hch2hW
IoK8Q5uO3ptDlvBb5NYAM3CzjEZipRuexA+Mzni7i3GUAy8mMC697URbANCK//85FDlFgtE3V1vN
ll6psmf3iBvlaOOe3lQGdJLbJox9RGv6HVTy3WC11kMcwu0mh0jA2YcAbBAzvd7mPGDmu40O7si+
gYzXfATuOuxM0NmJda3mpqQu2ohGIhH/t7Y8yazvdxgLCFxaUCkLeCkXuX7BFeblyCW2yTxxMEYc
D7yjEUsF5CP/GXBbxVOO7GJRar49Vpjmp9fOMbeKseFr5DEp73T/mb/7AoDSABLnQOm6YlsJ20yh
b4xDgr6QZuHofYnFuEu7wpqzGpXpRg5jvcRr/uFT77/q8oQ3QXPeWmLpwpXCeRPR1Es94NYuGrNa
BXe4bBiitHccjRgWbzCvuobrdBLv6WRqpxCG0LvqsHsfVJxovgv2LjLJVLkPworh6BYiDpQtKNrH
2Yo/Y+bgjrquSRycKXIxojZjV9khWl9e8Bj1iTeODHGNbflCI/9PRObkFHNZH1DZrSHy4aurMqzb
cyQbu77ymbsi7+H97M7dWKQlVU7H6AeMMgBVxk6ZgLwOWkGUp4kn6OD63fWPZIoQMUXapdYD9nI/
gmxnV1jaQmrx4H2MlpNUmkZgOrO7ftZYq/eWTkKs7/FLUkb0gJOlqBbQNlNMfdl1PNvD5ni+8IXd
oGul5Hqpqp6CmkDOGgemdWcNqYO6Go8GuBuhgNaaJBPqW3eCNViB3BFujnAyQzaUfh8KBsdk8NVq
27pBLAmwveBWXqGuQf+TdytHoBTs3nPTw1dJ5JJ4mM7hW6MbFSxYkfFNaai4Sbsy6yEJ60s02vBF
MLUd+Yos8nsuj6HtrPBYDY1n6hsgTebpgL8peDIDKcLbrCujT0O4yaKTgKdx6HuUgBeIGvmK0ZI3
29e59AjbrtYY8/052Y4pY4epe7iC0NpPfevwaX1htV8T42Iewe2nxreGqA28bfUA2NmhulMqqmjU
cTwsltfDOabLF/PPsB0RkYvUlRNnnFCRV83KV4WipyiWmOk9fQu4ORoV0ypXwPxyRbV6XKVZ73Ap
IP9HVAR42wz7ioaLWnlKRkEBoxiOGXxZR7hcVFj0w7YSfnA2VcnJwjpYNgqXobEsi9oE//OQFJZR
A4SdZdX2zjmLlmBP80zfgaNsS7CIAwvxbyfV/q/fIzml52Th3QfjEC5ADpD6NLf3g7Wa6UMnt2du
h9/NqQx19lvkb/B1WvjUUffc+Bi8CegTA4J1SXVypIQkaZfaFMlxnY1pF05tHrc2bzCKidRTlRMD
DLkDCgLWElYrbI4cKe6q8ETjL7Z4zkuL/x4oPs8PyTPI/0uo5otsreNI7+fs14kh8OMiUDihOXUR
P86+RtDiGkEYPBJAEdZpbmSXzZiZbKssClnfw4r0gfY+NnekqXWFN7TXD6uQCvMEkKz50/3Av4Np
e86dIQxxufC/vv13QK+g736U/KnmJyp+JCz48axlO4CXCDkQpKu51fLUd1GD3xBPoOieRjMJInI1
RQS1MbBbfo3F1/DPmUj5TWZyLES/Tlnn7OP73JnqU3fGNt4ifowmlJw5375f7NuLwl/nCcPHvRHS
v2qfI+sQHC47/2ndOPKu2ozsT9RysjQma0piKTd0dhfooAyqh//VKURTQxJOVb+yG/tYmebmdCFN
/DRcve72bXdMnC0nhLOJf/ErMY+DLy6lq8szJEjrCClqZIkvuapVxYVJGfppQlzgldCXHCWbeGKS
TSUaGpaiwbsuCwgC5i2MQMr06D7YJqaO6Jd1/z0J0FzWg5tN7LhqKZuwY9IpTYecQH15zNsS4xfD
Xv5AeW4rIlotb/fFWRDitd6SMJWcZO1CUhdvIy7dwWk7P26oUus/CnEk6iYdXtzgPmTQVmx3RWGC
NasctlYeySdbWgXL4WP+gRaU9xsfZJ+8ReLnpUmYTEJ/EPrWGR/q12Fh6JZqzcWw13qHdXLggQZo
97g+PwrdJ+FD7HiQ5FVShdBIBtGlHkSZGRzvBLl8nIlxbMXr491/OwD4oQw8MyWyNJxRpjNguQKk
pS7oaL6DK1yc+t/aWTC+vAFwvWbLP17LRAwBIBs1LobxVvB8HBy/2NaoHEIF/32IWlej6JC2SDo+
z8W+h5Wte1Ku7YPCrpgLmC33WIBbxcWNqOXTNomtkDH7Xu90xGtmbj0OWZD7Pc5qmJFEIJhq5+rG
ytHRVtnfTYIVZk7zNM7Y4eD+7bU8jHrSE6qrX7es0lhVBNlOgGzgVFTMN9qcQ+/3tjP7HjBx7i80
XZfmdLUgKDWk6zooRAYBHVD3Ira24/pf2C8ZKYWh11i1M/bHxf9B4xyx2H6P40CmeWDNqMms0PoG
m0d9kjCfIQUuNQSd0YHyoqSjDsd1LRHa7Hvun2j7dF7YtEmOuz+pIxTuYkdK7fb0tqbHTCID75Xu
sqOc30SVf8pk3VGcIFLg+C5nhia4jF9tUULaYuOvBt8qtgjVJMnGUJpOtqNx+jOXqA2dfzvBNAOy
qTnOPfXNn02oxLhhZSVESbSdcb11bc//L3VW4YAEq6TaU2KbDY7/FkBzmLKO5bRSxZgun2KCgKFG
C6f5XZEV+BvUmlywc3SInV2jFDybqRW3y5bFFyFabIrCImjuchd5dHsBYIwxiBfnn7ZcD8qvTTDF
IhgM5w+rgFV2cHDRdlGaAALrg9lZjZB8P0VZylrzgciAJrcP9rfVC04unN9nvD5UIk6QBotnjsAg
GBA9i3LViS/tBiG4Gr0GYYjlIYwfISpSbIWg7adEsx1p4GzrGPf3PIDrjIZK0OT3+loyt3/Lz3Pk
zG1er1LMNq7TuDfBeplJKjEOrWSOtQxt1C9AMLj5KD0NcVRtB2QdWKvwYYx06v2YpL+4U/9vRxux
XrUp9dGhOFEbD6lj6uor3v3jqtfaN3AefQb/3AL2OBCeKF0LLgJyt/4XXPpEt7Xyen5Pj3aVSDGm
Fpvmlt98cF18Hd4/GmEUeYuHih522aP+N0ng7rSq5OJf4FgNAU2bsA7GJqtLt152e65lU/wqa8fz
PnxVu9+7e5V3qhIGXgquMX+MCz52d23LvYyH6WFAsUnZNwU2YGHEKGKfXLvuRKNml9VyWrSYHMxD
OIgNjvo3kY+8leyJDJ08FkX4Gg2A7vqYfB64vJMLwGzu78ueacNNNGOmPVsuuUsgES8dfsHWRP13
aJPWHKgB/QXYzk499ma0stKe9vCw36Nn7PsYxAPXN1Gu9N1H2ECTw1lacStOCksNsEaSuq6hkrL9
JeHgwxva/1NZ6AYmhj66in3dSqatEnuVLoUm+VccJQqJ7yaZzcmDpCNkePS/LfS69y4j7pNAmBx+
X/x1V1stK7o+gGmPbv2Z76WenLtLtnRAcz4JJuZ6LdAUVcFsHRZJmou/QVmbdMxb5J5T/lxwkq9i
GP6AsxBcgeLO7R0dtIfpE1IZVmHKkANB5OnH8gSjCUz2m1l84L5k0hyzi5fVeo8RSTki6Vic3ccc
nhQP4am1pyVQmVwLvtBhu/ftqJQ6kzX0gQH5h6bVY14jNNCB8+U6cJpza2HHEXIk1hbwu56pdAJu
TSaf2+uRphX3DwPkoOmZWD7mT+KmbSZcQ+ORGGg55MQljTesW1TmBK0y8TuO04KooVEOTy+i5xzC
uY9ApFKcGomcpRTA7VMn38Vxch0/lQ/+7ZonM5DkctndakMsEAWIljy6743Su+AQSEimh6RV6yH7
eZryOUT083JGvUtv8kIj/BSfgxX298eSEBsq4ROGT6Yp2MXSN6hWffTpLQ1tTP5m5AbHU+0pq3u5
2W6KsgFQnaWf1XQ8hEK3TKcIDaRj4p/Eif0WlIEvUGhEF7qeaSYDB+9aWUCWc9mgRN+gnxlYkM71
pcN1PlRWB5rYSTv76AaT/SQxOiaYBMcaRhfuH41rFgXo3znJJJYMp3S7aX/UOyDrb3zLB+TuZ1Gu
Z7JTBpNqF002Y/uZeSKh1VPL2xWoZlR/bra8bMHb7UHxGOzKQwyw+6ZERnT2R3MqU/oDvaqoa4mh
Ak8+KvCnwNceWTkVPuGIOrB6osps2i41p1BAHsMAVdpVrjXMLejGfkMP6qAMxkZXWDI9nNcflNRt
xtW/g4PESMmHFAJn7q+vvnEmx4tz9I7i6jC5hmgPfif5dKYLJ+nN3Um0xLXB5sLJ8N6riZP+WI6Y
gNY8HTavwzD9buLuTNPZeFKS1K/TDfYUAgrxKpRF76KjHCm3FwcpgKUUywU8fo/KAWM4EeCLayg2
3eRG1DjTicD8+4alX9tq9BnSCC6UuCPm85NnEOZ4BlVycIZPG77AEC45wkUoPVWuRTElbk/1sVsM
csI3mhFabohKVswAD40e3FPkw/f4aup9/2M4LOWDjQqWwNtyEGcwtcLtnPYMCcq3JM6vIqlIhu7a
4twVT0IZGy5vtr42ks2BjCvAxFGjEZ4TejgEs3vXcz/2jEmbDeD38t7EBHPklILf657nvzcystaw
4xSRq/IKZw559sjda9KhOhT5WzIe3B5eOwxxgh6LoXmyqRj5uFf/Px3dDHA5PL/G6Il0MJX864qD
f5b3CmqUVEylLhX3FuaE9aac4YwiLpSOXcA7nT94nm7VI0XOIJHOYAEy5/Jj01/73BNHH1LgN/NM
RF54qJ2fVZDgcj3cr239Li9uS1qSeN8zzbHujRFHdnxGnxb0d+iQM2ZrrMPe34qMO0evBQcP5D0G
QO7Em1LCHfWXNJv3Ub3EO3FYL9bCrVUGW875j3KvtiPdNFINgOIfXWuXT2olOQLRpJtBXkJY1OfV
vxkDGSM+TSoKT9QKV2Of26up2J/lSY1nnoHuiePaHl2A+c7IUbvqaMTO3JlFpo0hoeflK8LofYEo
Jm01fVf1Rai5jxsNkdqLgHfSnB7mChRiKCZh5Z46QOb8rHi4HJKheByvGH5esILYCo4+wFtlYym5
c0k5IwHnqrMg2XuNyIcBixL8jki+ki7a3BXf0Umc0DyoQpXiiSpDMLz763nPvNarz9wNycRrMel9
OxZtbX8YVZTwOPzqvW/A0t33M5Yef3n9TveupGA13fbskdvIQ1JDkQp30poY5GKOwSgph1ImoNrz
18ntObbCMtxJ5Bilao5HgvbJ1ylgyPEFhB8NRW7RoEDb6EDp8RK7nA8nsTEgB/hhtK08j8fYgLdb
xpWueWgZWCLEh9fvLVcMA6XJU4CIZbw92cJQMC5oDIJw3KaCH00V0ARtW4r5Pkg6uusJ5nv6K1Ne
eIW+71vTAJpy6B8IuXn29735ejqdAp1I5fKd5TktmjQUF9z9ZWj7uwthfsHFzrd1HCS45TXsxuYE
syaht4PMjSXt/rACpoVMLUtDcYEA28/CxTYxCq8Vv4HZOER0SfEfsx79Bp1sPkft7vwI0MOyHyUq
Fmp62gLFP9iEkZjXsWaJm9JXCDu4b7n6zC0jbMqoYYhUEPICvPZOVYmsmtSa7snmgI0Dj6fGCXyp
ThNXnieM3Sv6YCMgOwCCPe/PegMObmpjHAxx+DnIExkbqluceOQ/Z4M4aZaCx8HwHGjtoZKZ6fWv
ctRzv0tadH3W29H0TjiBajQrne00ST8iws0PgvOcEFOuZot7VjfxsiKNvjn+8uDZNE+BZ12GfXa5
8h5bpGVfepl+QYF7XQP5C/e5ZPt41qAoCUW0nnQX9pBaXnQ22XC2dYI7cBLEKPnxKrjAA8d+autD
J5IplKuqReYYdAgtbtuAqDXddchh0n1iWGrW0nHpjrxNfvGu93GDeWGqZMCCNzbFb+/7cLgnWYAV
lJIUeXm9ilnBPPZhy1cWV59Kcg3BmxZBzDc9K4fwMwkE2Ky7EO+ajAPk1Kdyqa4FpGAmmhiqBRPm
3hGxph5tXK3gJJvt/ENup6fl+ljK22tSITy97fbjaCAzNc9vGFtQsO+5iD2Q1ivtAzfIyWiE45Fy
HkKCGX849RU+SE+re2T9wxL9Pw8F7E26umxruG/BillePUm9+O3xrs9Yn7GRIaj7ax76IfDhq1js
N71gWE6mU9r1gSHywENI5xXoh6C+AKczXbg2OuWgAqwJKRvlx+vP+UPNySCJNsOeoohJMKDFahXy
NOELvNB7jX4r4MSJkJHPDH14onUuILUfcJzQueCefF+nUf/huCESjKYd8OK5XFY57cS5d4kvBbil
l1PDNF/A4ttalZSjoGU5GddE3+HaQNqXRI72eOX2QwNnoxGE1LxJC24vG0kTx0DsUKeSyO9HHTvb
pGlGLbcsRxHs9s9+xtSydqS4my9zn1pA0LkQQr2NfdV8dVKgCl1uK4BtbSRPJ9I6h1ydwYHtcNTU
2RfmFhVQTCJt/n6Vna/UNB5ZjZewjEdBKyr/JHiguifBVhvfFjAkoJVuPls2984DaR9v/0/DxkTK
ig/erv8zSUKMz8Ca13fY7iY1LP9vIJd9DrpyOuMDEF1aPauS60Y2Mk+HNrgNAxWIuE6EJwsFbCrf
aZLF8I6Wy9Xn3JRZ+3UnWZFGkHd5KNJN4+LWm6sYkbjAOh+2NvXebhGFwdlz5bvOUwjrdvc7yKxX
17+MqijQLQ6ZB06UtZVnxRD5Yh4Pvk3kaaJNPqdeWUJMugPSOVy66wH2y6cnZHzYw85DsTAr0LOD
bv5KH7FQVmKTpGlzX0JOVrA5xWUTdpJNHR++AZJPlY6r+HZuAkRLcTmHH0nCrXkuEkYDYGC5vCI1
tGKoLQyztpSKuDHda0iCKKGxUSkBQLKph6yrhpdT1+TIZpcYopkdLPwWwJF4wVxGubRhEi2mAjDi
e+HtCGOcUVSAokzOTyYRq95DXznZJimJLaMTsfSxsizl5OcG1YzuqJgQqWtI2a/uA7RCHiah4xc5
CFClp8rH5eJMrs+2vfsMVyv2BxfF2N5z1VXAdOpGPmcyqvkz8LtbmLMbFdFiYIGZOZhIkKlXuSu2
HjW/Om737csJZtWQl9oPWlo2yCppAXrEmVkxd1+jU94qNYAmA25R5mp8TolZvuOhmBe32S08+xzV
7CRa65EYZLeInkBurwqa54syif8w7tVZd+hx1QsL1PpR7MIRrLaOQk9Eb6Bnb9+ro1n8SJy1laLr
PYc1b/kuR19BxUmuuv/yOEPIjHchOItF1MBNSy5fcPDeRVszOrB8cPFkWEFQrXGE8+RaysMxKHL9
M/WFMmtAWA6uqHiZ5+hi/rcGGCj7Mk3aatcDHn8LRWxj5yGplenFTnPM7hk1NOsY1oRZGtbXvjQq
B4n/2UCPrGazQexKmo0YCKrp89oDNwlCtrAlU5gF/D07k1oD9vucVJ8tJdfUKRdV4EK+hbmF9vaJ
/FJcxyiLlnMBzb9LKKbVaSCMqJ8QfwUtb9rpUFjaAZOmFtHFpwvXZr8lZAD9nlQ6Jmwg0ArCYrMe
SC2BMFfBfkfHybzQ1YqChPpt/NnYAGVgN3InlVcJh1CFdgdGqL4/KJw4dFHPixaaaZ4HNKeZ6/TW
eZ4lmlJgAYur791hh5Vl26Zb1zxrJdGtcSXZIbn8v+Nx31USnQS4DvQPTdA6dk1VVLoXyvBpa/bS
adjeZrvDhi2j94H4pOUwfpprLh4AZYCIsy1F3H5z9UI3QQL7E6g117NvtB1wf1thPETpvD63hjtV
cGhZypIVijXpo8AJlfe158M1FNlUDXwzkSfUA6yNVn4qoiu/rizRyYPEX9z4FkcxJKj9mAhXHazF
lmPLhEhsVm9Lz7AP9CucbPEsluAGTB53UeM8E77J6bgJkjIzpQNSvnADWAT1rY6ht+8K+FSU8t+B
Eesvu+SaVisWHsEbBOHzfm1eWd048ruC6QC3RwhwzZISrxoBjDCkI4t65EHksJigDn1t9FOBBqM6
MJh8s/IHUxccRRWDHDhDt9DCqBbO1ocRC5U98MIQcqGF3ZylSs1CMcvemQoiRB1Zx8/VprEx638y
04wf3oHKHNWetBkoPjicQOJfqpfAwo3TZoKKY+7gKSxfctweykUTS7y39sgC8M3Bs9uTgK1NKDdX
RRMXlpsYgncLZ8aOeByBSda5iv0K2I0vYeN/yzbxGIBzl3Q+9ORNtuCjW5GZr13aqPvnBDoEANbe
6nI7XHdXof1goAVG6dZB7nL6AOR+tcWtmqSY/a45s85bfcXaUrIS2qVgObC3EuYEdGXBHK7br8RR
AYhRB+u0A32kp3LI3VyHi+CFq6uROZp0w/ao6pxXot1Sdvw9OFDPg2j0JDLYgGltvXEcO6XqcvL5
uwfNIJjR+NDirLLZsCKpMS3gqiyHWTGw/mDpIYvVUeGsEL6mfqCFvqvkhvnPTOnmjJT5UOlg5YnW
4fAaxaKYIBdxE6XXALh2F62FrXNnZmkZM56c4FUYMv1UhEbDu73UaR3CYQ3A046p9vs4l5YAFtok
HVVF+VnR39gE5gu9/H4SlV3rEZQ+fiMzvukVaOGRqXlZksv8Sfo6q+KdGfdlpj70Wo1keOD8QjnR
eP8UtYZjB73MzQnibuNB1FOgdp4RLZ+032KuMt9vJ8+Qpij3eqNP6ltgRWh26F3ymbJm76Vg6YUv
o9yH1MmASu3TBrxjGUYFFtxYKz8InnjKj4m/QUWz/XO7vSvlE4YQyNV/y6f77GAtf9X/jhXhCR6x
L0GfjjEFM2BVeOl4KxlHRQMfYyrvKV3hGnNg4HFSGP3cPG0/nBA/Pn8PAyIaE6i2rNvOtSCv7sih
B/zZ98O5eLZvuVXXs0X81gN8S3zqAePc2oj9k9qNaB7kEtNLkv8VNaq/FaTT84CYSmewG8C+ohPj
VDCueN1ZJ++YoUFZ69ad+NuEQXZ449DKm3MQOjd+MThjzRoaFWF8pLdhqKxBvgdvRx8nACeA9GRl
xEY5Fal9thuVSC3pJfWlmeA2T3Q72qA761RRx+YZFhU8fswMv7/+QdO4P+fwC2XfBePeBOMNE4TT
FnueztAndUj/g6kXDomlVLb19Re2ZgNSjUQBysUqBAtUgduvK2FWHTAXIUM5j4a+FWQcVxCg3oJb
trTH0+4MFtdT1ixMWqlLS/aLpgWL5TWRxlCN/wQhMudLxmEHDP0dwn6Gai8b6rCkk+3Bo9sBMcdp
IYjt2JVwIeytanOwcMgVxUDspVrA84xEOlBSYnvBDESPXme8IXLCejrWkrlswUXNV9f8xZ5sUUce
PQg/8HVqgTOQDfPKthSdjLEBlLjYm4k+KNwN6YMCK1UGM0jfMg78cqq8B4T7MK//9UXBI53zndRA
6k7KfLq13YBtVzdtwXshCtOGbFE9wQVWDcEjrs6lk+iTnKaFFxTkWyGgyoBgeIt1aHUwus8KXvsz
eoi9tLtg4BmYZOIwPnoxjGhHy/PC4QwSTp/6NxALy8ilmG4c8pOQDeyfslkbTy1urQg5573yjwmk
0C/9FWSgtosDO0DMyQg6UsPArRMf3rTCip79eTqjInpoSsyOcNGfc02duo7IqYJd8fwxDvsHbwp4
EfXWHA2SNlvg6M7JFd6sp1IsSxjL011z81Y/QpmifIQ4Xb+KbqbbWg0C8oSZL4+9siXzTXIcjKgM
k5y5wbEZht5n3PrifPRp7wWfMDNtHk7Cv3SEuZQjTROs71C1ulvv1MCSG8pQrrjuWVHVgrMD3vKc
HNOlBDxTYN3iIQmnCS5ZNW3MzyddfYi8CvomWgEo5CdfI0yxGj6NTHCotp6vV1zd3Pll4u+Ko/ei
KQ3/xhbHyoXIUEAzczBhQdmHwl7WEShitTDtUuMkwzo2b9RG8hfq1H8QIJlF0QoIzDV2jJ/RQ5cF
7mAOuoNitaYttliBL1SwCRS3U1YsEIUOZh4CHQFzHUs8DC0Pa61lM2UZHKAl8stKU8iv7ndtbwYR
5mdRHCfuuRsdMApqRXs0NsQFwhNAp4mWKk5JGWCwRtMfVnNQymDmUpFLygc9cNdBaR/uYDKogRGY
mz4FPJt3W+bfN4vGRiPPM3bLS9tLbsnh3l7DAVlbs3CCdBYnXiCNKpy7WaR52sR5KdsIZYuRRPQ/
TWQ1a55/UaS5P7XvzttkL18XfdQfpVK5Na/m7vOeji6BWQD4lR4L30Hw2IbUmt2dcpUzJ55Xkfgu
Tlulp2WzF+4g01YZVdtcVMHieHwqrIyCqLVSNRI747tUEIQtpT8JPHaDFpvyUyKv7RLJhwFu9NtY
pa9FeI9WKGPvtau0VJRuSxQgIGb4VGU4B3QFS86eP9cnv4OV2WLnIQL4YKhrHRuvCL8qkkQMmn+r
BCaJc7q+I4f4V55eNSw5JBqya0M35ZFAzc8wlm+3Jd0h66pnoNrmDtcRpboCSZcRVKhIGm6cLqsb
zYLefYssrAuGCiEegaIc7PSB2iIxU7wxYvPdG/7ESaIsNJQNmjWhRosc4/NXuvMpkOG5qB7rTDfy
vYrcwvzmd+OOTd90pLiDWxlKU5X/jUBnvQeby+oUzdLp582hqh3DmfrykoyyuH51bDvmtwZl8P9N
+t4Q9i8RzSj86tcX3OVnSVFI2u1+nFkRy4QpmJ+2tb7ujpAAHQgDSNs1/YJvxIv9uQegeHB4Pd2P
c4U1sm0Pgw9hffyISwDE84Vdx83gQYRqa9nS0h+c1f5ailTZxja5yjuqGpuQqV174O6fGDvynVza
oapmS9xkxEBtrNpsW5sb999GiUMUkDONO9bX2xUcBADOl0ks5a/cahsqnjSM4ry3sVfVlF3CwWuC
h+plx/JjFV/tcQYiTZY94tHCkNk+6r9bBxbTrFCcu6+Qzy1X1DZskcl6gOH46EvxxzjlleRZ4CUI
wvslJwalPhid3T/rlY/3Bj79AiH17OnfCNlrGNtPL2aOVEOX3W1IlpvMBFNCu5+u0IH/zA/TuHbY
uvPDDGGss6kd7G/1m6H44siWyNRp9RnUbmawZcTZYC1Wc899yd7pyYMCQzIVIKVbC5J/jF1ZThsJ
aSDIiKVHQoLmGLtvVtrlkzAt5WWtZNekL6CNNFJDZabJbY5hAolMPX/8dCPoAGDQ20lW4LNs9m9U
mDQIeMNUIpNNDK+FTBnVH7WZ+iUV3sQaXHmmF+mlMIJFCk2vYQPh4+AKqSV9nhx9u1jOOPkJsxzd
2UdOGEqCK28IhTnWz1SSlU8Ko1vhIg4mEPItyXp8N0OR6vxyphVRmJlJQow2gXeAwDKyszYUSqHd
XP98gskPu5FzRTKMaoIggkm0ysf45OZgIaEjNE+bq9vEtCof1nPOH5NrGV24EuZam7XFKA8hceCY
5g44k5VnFlivM4xzWqCtHvbZFJB1wjXaMU0Axu1Sk0r8FPfVlq65qBqwX4IA3wbFnxC06GWlyxzI
iTJ5Y++04UY4meH7hmPxyTWWaaXEfk9J0eH59NajM5LXFLPcQhzgyr1fVfagMhNDjIhkEpAkAp6X
5AZuwasB8uEUJtSWAKGZNeUbpZ9Y10A+3fdbRjnyBwTqLanF/+58twmZT35I0gnlc+MoOd0C7OMK
tadgdrPhtnK7VhoNjrNmcz05WuHHlRcNKKCCOp2S3NJldUCz9ieTf39URq46o8rn/jKMlO8QBlqc
MgjQWrrPEbOHW0W5IsYvcy56nz3d4NH5ffFJVHHYEqPniQ9QXU9IV/GJN9Py/X2NwCfZ8YEbWhzl
U9XslfDXVIMoUcgho0ja/Q7z2qdcGAbVqhdHGh0hNqnxpQIjsCQj7T4yFvrzePZPW3XMve0EzavL
1VBkXQADX8mPCgF9Yycurl0goWNZ9x6opn4RHfvFLQv56u/uqyIr/uUr9pvoOvUq83xHGqhrA/fv
2MQS2ktsCq3AqlckrXW7yA75RDEOSW9CzOQsENx3CGcklJo/uIfNGWh/o+kfcMzikNE3CGIHsTgF
EZeDDjzxxsEBBXaEfLVK/ZR28JYmyc5q04WJJRHXIjfQNlhcNK2201QfXOo4fVi2lhizsmCJ7o0b
IBEq347OOd23L5tKXPmr+YaKNQoyJD2uw/5BqRAO65uCkZgBfiOQmIDaBXpncUc/f1PWLCvzhjM9
4RpDBfsFg3KkwveW1wu0yefkWXcqRbRTC/24Phv2uTnNefsxc4v2/ybW0+Fev3eUA8m6n+8VfB3x
nQwo3F+ffHT/51vEdawu6qNgVgspcmadLN9DTZsNj4YGBJ16rlRux63j45/7xKlsP6OOTzi+cw3J
CFft6y4H/HWm6zTlRjeT4MmVvrmPzFeCUTP7uBoDV8HVd4DIwLjvyAGBZ2sXFWFQSxHrovsy9PQX
wJCrzXOLzpcv53PijXCZj/qYCx1T2LWnXgG/uFz947YogLYA/TuoEiGNjS3vtM1DrWKWPKEqaLjw
77lg0iSTo+z0BNN0Ckjl0H2/QVXUURBOCmpfOJpED9iYgBtjIHnvAI/h3JOOI/MM6Xztk1WYus+k
G+ceqXPlM1cqlUlrDQ1ISmBgI/c3Lcnf+mi3ZSIteAiMCtrmaUFj5g/IIBYe2cxoK6WwujwmN/+J
YyMkZ32mYuWqtNSQrXueUS57fUgt3qRY0tPXWcamSS1w59NU3PU85rIf5Gc6gu7TE8lPMe0cISAj
JF/Aa9ucDHeZoo5dN4S7fXq5MFusMyYjJyQM/yFU0XpcxTWaDeH6ije4JylKhJ60yZYeid+n/f16
DAg7Wj/W1dTDQL7hgzyJTg6STCXn1ILRRBxehoE7GRaazgAfYhk3p6Sxe+m6JBkYELh3WixEj6dg
9S+WzvAXt78dW+lCoeMRlRt0qjzzd9nNJoGvQ5oAHfNFDT3/M0AQq+G3S0B9+/IW6YStFqbWkQCr
nbiG+n3ydzq0n9qXuzB4q6Ym/b5nJgj56gjoIitgHm6a1MRyfuyUaRR8O7+v4fj6jJWL/et+SCD/
HWuYeYTKal8qHxIJ9UGd9Y7KHzi8JiBMTBo6R/8A9RL2u8juwRzPepcspOn9UCCbr2tvBY3q7yzz
gtHuEJ/OBomxGz1K1INNu2dZF98P0XIlmpFoAAQCKWxo4JyWcuuH9svRiu9JzetTz8RgPVfL8/h6
fcsTIyMTtcjsPtpVKQ9oZ7a85h7fBGCYDSZN84q8gd8/Y8u48O+Re/1t/6Jrv+eQ2VaOFmVxLyuT
Q0r1vAiCMjkEgQWeFaOBKA8XMNazWoUX8kvWXwwcAF2Bf1i8xECSQGjbnnbe4M7J/W3CwKQd5CeZ
dYsgniOK2+XzybcXn2zmFvVlnFestsURGjQjJq2G/oV2g1wK8rpDLxJXmDTbsajQSw0jo2fo6LDB
S/5z+VjGxe1D3hjH31n+XYokoeBp4PMxkzQQZWUFR16eyw0V5tbXmDArZWfZYPcn4tUf3lHVxaaV
CZh/hh7CTwFFVDdVnMO7eYO1tKB7vCLMEjjoeQ0KSezVYyJvXO+k1xwY3UlIbezBHXxPFNrCEu1r
k35OPDFy/ZAm3KQ43sVqEICmWXlfwX3sd+Co6pi6RUfoE3KOOYkusSGHApiExANOSjQ9y4n4T6TC
aQK3N8ehaphP3vzj45LqeWA+NcNdUjx7ors12DEcVXZpQhOAZQeB67wI/9HSE7gMR7w+5R57dnXf
WOMH2jYnRv8M8JvqyGRM6EjnGl5Q9b4I78heN3FuPXdYJUdvC8dkUczyR7o1EsrMoIG3CbfolQ6i
crKuTANLqlBSGAph/94vVJTyh6do5yidbfF9vsO9wg7grBbnYRAls/w034lbe553XOWG5myPhEmU
DOrOQwBvOqHV6Vf9QPuytBGX9uL2O5hJLIeALsDCE7A3rOXYfhshn1zEIz34yBL1tsN3hwAklxdM
mMqoVqyZLuNAs04ZxPEJrayYdLPqS8f3OsIuDZP0oj0G2iYxU533YzpDZ0jQ+4WsNf02Bx4/7xfq
FPXD4YD0jlWCEHopZ1sQa3/Q7Md1QcJhVSWwLeE5cWi9NlpFxGEA36+LFFOcLF0Rq06ScEROlhM2
wRXwGd0744lbhZ6f364KmyVvTNOmrEgdDgOr1Oxdc3PLUiQ8QgsSaoMqmIUuxoKzN/UgkMJI0cDT
Gmmcsob/xB0LhtCxdLzdd0wCltphX/caIfywRXrh8R74NTX7SmUPsfu3FPxljsbxBwSmY9lkJW8z
K9Kq4oeSFZO8/PIt+gX5sWSdQAdBkXELscFTTMN2WNBjG/QZZWnjz1MpV8cDEaU8ExLwg0u8B28Y
HcBPH1jGBAlObWf0gfGdjoqvMpZnBrdFvthiNXWMfOzhA6tfacPuKUR27rJoilspXH+xpTeU6Lim
i9fyrPMDCFWh57/+PxuzBHHaycCCdNEG8S5bwVBdhoJnbX7NPPDYN8WVOmHBF928sfriIlrRwPVC
woe4F7b//Gxrx7Y9Ml7lDv2G7MOY0S/Ft+VhORCFhMOVtoDxNOpn6mxHj1Ccy7QLEaoie0KiVV0g
BKGEM2b6q32g6y6rf6H+zPP+1h85TA1MVhK85u/d44AmW4nafbn/+Za+I0f+dDTmIOnm5RraxT7+
CHF+7vwtUPCy8jZaAA3GNOBeJ/AqwP+11z2Xd8jXSUfKVWWObCoj3pNYSPNt6FETgHQ0S7C+klY/
Ogool4yOeW8X1o5RkkPey6Y2HFQ6ldSUYIe3b5bu9h2Qiso29Qdkb4RRMM8cqUQveAeUtruRibLo
0ApQs/cMJGoZXw3/Rk0QhjmXouaS774gcAW4EcH9/jnNfBZKf6O1ezicGoRqpVyT9MTYnYhjU46T
IrrUexUAJ5DRecFvGYUeAmh68Nanq8R9bOtpu1ff0BHgHPtZGcj1ppTwx8QekL5kahsDq+lHqYf6
qM48UzZNfcCjs2g5/PByxy7FIgyjGYbDO9SmZIEn5AdqSkR+DhZPkcXMHRXZ0BnVO0b7Ij9fM72U
an6YjVK/oN5+IPs7Nk/LRMrPmOA4yo//poF/jCfNsW34+zs6zk34MY73R/wjTgLlaiWs4Pxjv5tL
krIS89n16fpLZAXCXqcMUOVbHLEbheI83OBXlX5U2QZN4RTNLRoy4SMY0+juL2q4lQIc5Pqu8D9+
glAl682wlnSoCP9C/6O7+BecyGcNo+JfauA/6STJccmeB5Xgwekt55+DudYZd8Acd7JaIpQE6zkO
k6c6jF63R0DxnH5s5Q60kT6WlvfQ/w+aO9P998Gk5rsJ7L0h1R/54/NTpjcLDIce+0Avbv1CgADd
gRLoSdpjY55nfbgllL+AzmFNXTzkvARW3MWJMHkAuRFtZGLPGZknYIUa714op4nLpn8pY0LGBgfy
UG8cgFR0BEBqBv5+0UPhXhgX3OyR8/cqDZ+Jp4OgGbBD//1deg9KElQeg2dJoDeh5JR5hNXiBlVb
NErZduu3M9IJuIfBK62Qmtkwsi6bsW2wtQqfPKOevm8G+a4/Xkrb2dtL89ByeuIiwlf3+fm/swyg
w0jt5aHTnAUAxvl/hHshvifQkeQ1DAkAgUMtQiBc5ndMpDbXJc6eZtSb3Z72miCd+oX4isfvbyJP
jPJvJFsaUcwFB40H5/VNC1iC+o+wh2IIUekLQsGvUe2sRB5NhdYMuC/5yF2RGHeBSEtGeXflzAmS
URcwMHGXfrX5zhH2Zskd0Ks1OGR+J07LUrxg+zNANj774Lphzl+p1rdJABV8iimHpMKiBzCLARuC
G+hGsVEs+9grb9hUBy+uYqtwnHY7Ry89uctLwkfNU8OQIUL2vpIZNwNDBKGtToh6zEBphbrvTGN/
83aQv1mW4AR4J7wWx96xbuHm4Uy3Qn4XMub/D/GChtye5uV+WMa7cEKgJv+StSEEpRPpsH0cwixf
WBPXdqinuXjNw5Dp9eRAhthCjIuQPF3kr24MWbcW9ECnk5PWeVjmXRbYd8dUoXuzlooGLCu3HfOp
Auid7FyKI/6ij4qZKR7AMhPFLk5HATDuFYYwVHnv/72iFeEfQQOIK3xUlCdsdqlKwjgIhGBg19jn
VhsP1UeLC2fwx657EpV6HSR8eNMfPU3aNXeGFlKYjzrhDwb55iubeU5egsTBzHNNqTA9h0XIi8tR
m3IoFu+W1qk/XSHgfy1jFSpeVttt160feZLQlPuUXgIrozEUMTc1lv/FgDrsTYR4ZzsORsny2O8x
vxFYHGHdL+ROQpbhoAI7PLbaeYunU5tD4mt4uwMseWHuT883Ndstv67++KWy5G6ryncjckzHZNWp
HHA7KGRRH+6ac6zWUMydP5KBJ894u912tjICro8/Ok/r+2Uy+CP1mHGp8XynsQEzOWb124uujasW
92/RSxMPofMBALEpAPuF0OFhCtPBTf1ACLxV/k1/zMdrRrX33afofoDKchBP1YeKmLSPO8LL+3OJ
WceTj3H4P7pT6H4CgPahtq+WIugNJ7mNh/r251Glp5TsM8Kunr4TtrKcFzRc0n2NyilLsjZTX3ke
NgMawh9aiDlYh886lNtn2i02qyXLNDOJLdWaeNQFItI7vbpNapho/aJcm57Xp0wukMRMJkd0AGii
RZistDqXAJY5Xe06IX6q2PvaGrl82J+NG0oV2tOtqeWDsEQtjaGvcuxl/DYSbph4WSvXp2e47UI6
Esnr8NG3BHpTV8v7OAxpzdKPI8TxfWxtvo3QrtDOp44Bx4YQEmgXi/iPO8ExIQFuDAGk5a4G8i9H
TivFOCvrGDRANNr25gJQr8+8CEXRhT7CnCfIxNiXcVN6S7xPtg1T3LZ7AFzDLljASkiRGWJ94hEf
eQCyDRFJbpGlJ3IISEDd7KX255qdXMqTS0b0mmJAOwxGkHvk+9IcBZnaVYlMpchCXIoFw3+iBv8T
tnaPlfDkCbkyc87DeW3FH51srq3s2fU7JR6/Bgg1OudEzQKjT0M6TGiM8WTeseLNeD9AgGgoQraK
ZeO3IqeRSpm6DtT81JgR+vTNl2aqInopJmlpUhsRZ7bhZO5wN5w0mDqu4+CeIMORBGsiScS63TuU
CaIV5AvXO5hdpCAHElqe+Iy5caKIvM1lWWANWMeiXXjG8UxcCWAVx71VEP7aVwAhEuOWdbJZ58/v
kSJwTw+xKL6XNzJ6wPSbd6N0wYHTuotUuxH7BPeDlGGnAVjJ2C6sFhejBMaiQ7ItfGxak4sCvibm
yuMavF/TbKocffS9Ws4Ijbkc2oM/0LHcGYuiryzIZ7J+cN2YsRJMzm7rIhLT2SqifSxp5+89o68x
n1OnhVW3HXQIy+8sCFpd8mGjK/dUhS1x4JchfcXZnRtK58zrHMoOQmdd2T6xNC4iHB7OgLWlb35o
SMO+JmuVl1/Z5HyzIHEhQQvg7uQDoCLFmiSnQiSn/HaiwK/2gvLJtS1m5+35+AlTamd5szQYFZI7
yxTTwSX8VnDTrmwHH7a0qxK/ati+qOle9VWUyZzubwYmEYwuQ4Ak6jzPcaBpThjo20NLDzOHA1OH
so6esB+XoHjNW9wKtrDV1AtbuPtc+Drhlon2H7epdG6cKRQTWvWpMLnGiYeuSmST/0s8HC67F9Sh
ZlYgfzMHXtU5LTGjBqoqXdfXC+gP7iea0e18YARNO8ERQ2Vz5Nu1WrAKFhodBizaH8ny371ZJSM/
3FDxwYbgh3L6kS8rbluD8e0WbbwrcphIt2LmSQ0Tb2ZYwlRWZopdd1iipTeMp4sfPTyiynTa9irK
szbRjgLTHD2ej0D+Y4rmP5tHedLMWgWspEHo5vOjvw1pEWp4sP4dysmZLDJarpIkJkPTDcBYr5qG
z76q1zZmAF7Bcbg0FsaxDNvx1t1JHvW+VEJeK76yK1R6xHAanwBdDpnlNCsIhvWbMAXCLCItp+cu
Nu3GvQ6DZ5mBG3SzTHh6MMyottM+9EDREa7X8vaEq6e5ad4TdPWwm33Ls5Sf+Q32x8ENFxI42AzC
k1+KC4ffIkXRTTp5YV2kWF0pP/ehJJLd8HswO59fU7JrKnUZTrP+bXFtEPGCk22H6mUT5A+nlfUI
NGqJ31ItiHHozYYcBSF7mkthzP86J4Nl7unCnwaT1znKmUSTWlpFc86cm42PxLiYanG8fV/+v87I
mkiHfwQMmlvvBw56b9KyB4sGU6NxbjDcXfwT0sdQisPSejIOGuRMMjMBZ+eoAK7bnzRcz+2EO+X0
dmpFfz18ghoYKOwEBzPItdQCuD2nWRO9gGCl2H9jejR/kWgZhJ5g8wK8tyMLO71orx9u8UExQErA
lRmlBfWmyEi6tRth/x16FnQPanECwuElfXBaWyUxdbURs6+KTEXS9wXULS5ZxIwLuml3XUtGrs2f
pUUldXSh7iLM6DluCFdm05u1PN1THcrpI6CtU+/FLfICmRmj7/BBRzoqjHEHRylPUMarbcdMrKzh
yPgSwprUZUpCvSRq6C3ew2qI/WeePwTvNlDnPWnIh4t2Jv5XfK4HoXf1c8AEIxBTbLIgQorCSB0U
Uv7kLshFZXl/9iYIpj0O8qlT0dNWIxcTVr8HLPmgJihBpff+D60KGvl+pH3V13hwVbK4cBpyrOKg
hZ7AMWmeXGvWqZWNuC5YZ3Vs/Z0+ZCVs24RVlYNEERMji+twcBXwBc08A2zzDKt5CEqwTfVQym0h
aYRuo9RB+vGI6Eta5BK6zT108jG3xeAaaMaheew0tYwdSK0Jypqi9yeXEqIpQyEEl05N8BXPsfTP
KI2xMCyGgIbdDRLVFhv1z8k6SgAIXhk7sFM80YgbuvazxGhP6SP6sRPYtg5n2fn68uKc7PsGiTFo
Kqyza4kcEL6cIOSOaed7iVrDq06FssCMvNsA77XI8fWFCzaS0Tp4FPtsoSfa4vTPYY7GJE6rZ6Nu
YqU6Tj19FFOkofPx5HBg3dTBA9CWl3PwUADbb/JddFUW5ZLlF2Cp3/cX09uCzRX5Xi+imbkbTIzj
TsLhk0cN0Ifi8PkyDmGj86KVf+ZoUrwvcwlM4fpmdfkffed5m2dsC+yIU3hPsKKBYx1B+Ba06W+F
fl+SjQ3iwAs/7UZ8Qs1yK5SwXJ15qV1go/B6P5u6DUtJDvb8HPTQsC5HJdKBjDNF7xm83WbP/ZyV
y0sKdTclUIyw3HFE4PZxppRA9Ud9m9691R+tjOCEYpN43seGGcJ18iuwgCYdhxZCABttbcbBFDRF
RUTFAEnOWGyaxh1dY4JPhE6EIYm5fjBznC3vEBgDiN099VkpYIdij1JFV52DTfe0z62ybxnu9W8P
HpxgTP8YPSXn0KaG0gMzMqqSn9Hjp1vAdUZXlX6JMbcQBTefc8Twy5aw246iy4pTFE+YPUN4s+mF
JbQaWjpGEoafAMS8U3kpZ6ZKHMIOPraaELAVY6/T62nZ9225DOGJkuuVCuxiGLm7os91fEgkRQGX
+xBHwbXoeF7ryVs/n4R2Hx6ahKC+kIQk/SiDOTRXnwu1DLVZWwwBd92vhJ4q8QH8z2N43nCbI9XJ
J09IbeiUtwuVyL5H6yx+DrXZbZr3b8rcdQ6w9IZKyEkcV26N3TwWAS0Y0oHnTAARPWk5V9hgcujY
02juXaoYAEbdL2P+wm+dPHlRSo4fvVBOy45uiILZ81GP8izf8EOTpZEk2wI7yTcyCAlKu49Z0ufd
eWspE5f9yflSUG32zOrnM5+vrhtN83AzhPDgPU9ztM4zf9T1uM9tly+TDIrcvXexSaakShAPozlX
dm2EhXMgMw2iZ7nkZ/yO8WJP1Uud4yU5Bg12cTkB4AkKTT4w2lGZYoYquVWeFHz1jIOJdpHJ8HAY
wI17Vqr4QOX0FdjVBqoYxl29AcUThi3fEazecOBv3aMKobQBfEhGV/bGNqj4HHl2ZJmGcBn3x0Ni
2RbzBsT4l2F3faiT/WwZFiK358a7P+8BGF7559OmOhtH+EyWlak5mSAQsi3TrsZMe4j78Zy2xWe2
0rxNervw6/JUXAUBRydHnRUR+VwMI7oktvo5brZMjHTH46JLcU7N60HXig/rSro+zGfw53yMLUeD
2R3UbHDA00YuIsK76fBRoerb/vDilU6jWKQcibHv7np7YO8O7nExpgr8nnT6bKVkrDh4nFmHK1Ug
t5z6hyhONokvrniLD9n3dGRfUyl+fP0EjEklKgSMSuv8FR1e2MTCWhm8rAcAOdmumq0aCEo8Q4dd
xkfbswHuhsdFffsIOt4yz+BUQTWeffK+kJS/O+L+/J4d8M/78Ts3fFNs9P6vrVF4GzyVqiJJ810L
B/JzV8SuYIDjF2AzeGHfKy3lbopSk6djEUXQE+Lg+/Drq/8NJN9WLSxZHcCBmLPMMHPMd4DXg+kW
IMP9gsoew9qbDDALr1r6+ROnm1pTjMniikxShUid+5lVAbs/WHM8iX+OZsBdSZLsP2rqOkeBnbI9
Wbb6yZASieKk5AHMNTKeothfP/KdduQzNcJmH88O7DHE6bVgAnEP0z9yuhl3DvXC1F7iaE9bFJou
pTdoaKuPTf6iuYqEHnwESBuiUvAQq/rVesOVmPr4VNgA8ufezZXShsKZN6TRcq6gdvBPpfTzL8Se
1CIKrFExh5aMpEyhU2hZAakp66MVI74lKlSWTkoihy5jsEbDBoOSa4v1Nr+BSHyFoH8YXQINhHPC
3YB99QrpliHXQ2SeUqgGKmyWJlHtxsLroFC9yD+TFzyqztoYsLJmH04/Wkyz45QRTgh7VqOwzAZ2
xBJ5yPiO3PJzEwf0eDCt65f2KcGCBnpTFLvNld+1nXQQNPtmU3vrSC6n16xrOTwG3bfFyTCRjWLO
chIupUPhOxArktYhS8P48RYzDr/8fNNQ01YRFD3SR5fuyf7kdKnZa8r5ODXtYpf16ZjO2MtdmY1j
3WzEZ4J+ybyAeTpOlhGXSJ6yUMvHyQhd3TQuMdhv6k7T3rbb20FsHCEHipGVXO/9B68AMoM2PbV4
bQK8YNGseImbNfAapesfsYH5elgRDY220AuYBvY1COVptvzplB7smlNnTHfnwvDueMwFh/TuJD6c
YjhpzvPdzkVI67xNuunXwiEGlqSIjqdfyPzzio/8tBy83ZV2LqBknrZjJDnUyoHZge5HrlxpPW6g
tTFqCIcsHXzCUnDDYmu7D36AYPLq+fxQenBh4mim/fnnUsuYN0BbjuP9DymS0A0xU6QelM8YIkQA
w8PcNqa3mdmUwVdjLrstaTHABZX/kKWf9t4fTwPcphkH9+yklyeRkJC3JMTR1SUUBNXuftm7LbnV
HssAxt9NOZ/7Q43oJEtHtp9hhH5O/y2kJFrCVsXGrumBNpZsESyMjSx+cBjN2gr7CkzHMvwhMX3h
1UyXwep9O1CvOilBv8j3Rkh8niQjH8ZPphYdsPTYFxlStYurPFepMKrO1AZt/CeW0OXaqM2b0xkx
excri4geGCV8v7EMGKJLR294ZQMxUQxO2oG2K8vXyVHgYrF7Gnm5QwEHWfsWSdUHgYLqFY8wqbSR
qzAT3AW+FJOALyX2pZLC+yR7cdbltY4WnN1GsHG9UMNBrZuvNAkzcnHkR3g7CSTc2StN0oNTvcFS
UN5ju0I6SyJVm8JU8gYOJqVSL2ztqgmoOChzzVRBMnv6Rzuxz4Xnef6sgVo3kU0jtGOoboSS0xvK
5blqpc/OJbQOdTrTar3WfuayM859gU9HE9W4t1TmdKTFqqHKEW0Usghd5eto0nwRSk2B4E73G2cp
Uonme/7mPy7eeUP8WBlLdfiKFVN6AmaeEFCu4NggPuRGpMIlpXgKHXMpXlRmLr6UgjUKr3WeKS9z
ZGcm/GpIaugEX/nM5y5eU9bJ9jeIARA0WQpvkWzx+2/LU6M1ztRarzKxyzSemYMS68fa84QS+F98
UXZVYXIo0Si5UHfh22Tb0/gTB/QsAOTWVcDEgoUDTVAVho74aLUakczCv+PrTibh3xClwbwqpCx2
oG2Kr3ptsWqYlA41FqJR1bYWnlp743UFxMNLO4gqvnNNV7ummnpRTNjcg2/1tmQAL+Wmhb/WyB7w
jjuMxslCE84myEtoINZCCN0nQDK2XprXZ52Rl1A/hwDWb2fDNFLf1mY6b6g6YeClDXH616NipEjQ
KuQ86teBQJLmlXfP56NtLPMIpYxi0YMhJHNkq9sEjvKSGUQlAwJl9MMbPtrSMHdsvCPbiM52sksW
9LPBLWvqn2vVAuzsImG/+xQDE37zoJgzt0W6LGsxtMxARl5F73JiKPJIoeAO59SslCnkfYEWY4yz
2iHI7eCt0KJpuxmZY/rib3immHsMPg/Y5HEiefFeOUQfRsUG6fFLmixA+JRQLm7h0nkaRdo9KunJ
riu1aQylzPlhLl6OJOfB8T+wv23Hl3ZOixotwGqOOi2yBs2P8YZfCdLH3tmzDM47Yt+gWzefX8zL
NXjL0LJwZcHVXON8bJyOAttSalDVy49glVW08d6hHE/VUgxwCNPBSxyBeKVIrBVm91/ndEo6sBlV
9tbsNxdT/fucRsiWm+1yVLhGPIIkbWI0oGKCu3/vLcP53rwFey7gUVxmon0w8dWAT2ekv8+fu1m0
AjgjUgaTqW8qKchisSD73VhLC95Clc+CS6SXp5e617bKkU+DE/1e/mXv1LkOG1tegWsw2/d1drhg
n1uOpzCGsWTNgNIaTu9hYKLpi1Vt6N9SSTrN/5MYCvsjeQysPP/XihcIl/BGUfmWrvR3vh/tPqO/
d7GUnwszDrOra+UqPh5JK6AP2Jxzyewbq1GlcgGQtVjM7G1W3rVOAfoOboIxUpS/cI1iqHJXXRL+
p4fRkwQs35sf1gf9j7jf4BEnq0q+ZpP1c+PFgvq6ojv12JKcMnxcqCcyNTiTyUDY5XDQN9V+m/J7
0xlc33ahBZBTKwG+hg0zX3RBMKJWAr1N9hz2eABH9qODSIaC14ZIjS85ruz85n7cYEBN9zO2SZLE
DOkRIVadbpxs5/Z+46Xaju+pufR2W4xM0TSr1LGlRg1pHPIr7E5cfwEl6GTQ0oxATxs91tTZ797X
GrF867TCBvTXn2wy/xAsaITk9TD4wxUIgscxhY1INWxAFpFm5mIrFL6DPourDXQ8E0wH6zd/wb7q
fPG7vHKPvfLDnsPBrJcyc/hfdPb+a8RH4vgtbAkw0vSCCcb9pmZNxbluEnLq2/l3ZdqpKKHh03RG
Dq1YfzEZwMXFC+XX/8sjtkqGfrRBDO1oRyQ+7GPBY3cI161OzvWv8U/+2FGmhpekaeEONJV4scCL
RYWGbB3UOwd/RvBrdLcFOyhfLogo8NC6G3zZaPn6KfPqK0hdaYHwzwo0qTrIMv+bkQYOx0rYe2A8
SYXicMAnS0Q15dcCOUXK/KJYqz0PLjRxaBPk5HIyfPK/NMCmdC6HgwW/Zxz+tsr6tbY3aulj61AN
wt1z2w/2N3VAlK2/4HmWakjD6uMVzlMwU/wH6gYkWihfNL8hyExRA5nujA4OXabDUGyY7GE9dl/N
C6Am5pQK1sc48UkY/fADzHGZb0WG1Su3HZ8VVsYi8tr8V+2539+Jz6PEiJxLF06wyEgAI8Oo3NH7
6qnUyIRsdmrfeQ0Vxg1evYkiexgo/TXiNzZb+aPyUqcMx0u4ASSmiz/4ve5sCBfTYKzWN3ljEfc3
eg5mUxKKFwbsE6Lto6zaqK6h5OYEFjar223+swETa5e69TlLOCBxnRxZTjNNi0JOMC9fqyA3GfqC
3/LK4W947MP9JDecWbOZKnD1fKfD6tKwQ6QdQWJJZibJaZOPS4R/UE/PoabblrZ03QWbqSi3RhXP
+DTUf7d6tTs/xcdhYk34S58L5Q0upSlFvZ2oK/uDzN7d2jec60/PFsUIFvEqD8DRbOKcIV8mGjyz
HNB5X+NLA26+tn9AsEQHI6vqmq7pQ0+oM50tcNvKHb+VnlR6Wik5JhpkiOcOhkPsSpG0+wMzg2W9
SJsPZ01FU2p8CZGarTJ4fi+QeE+kpGTILzHHTxX/3Uexe48lSdm2XXEgJOdNYBkLDuSCJLUdSgxS
sbK+aoBdoLQO2I8itAXDI4AORf7VvuHzQazrOvGIjVQMxW5zgsX7GUcx+Hsag0ajyOUFevJBBHtM
OeyjFagmV4WebGoNYOiDGhsJzvgHDZdafsT9npm8FvTb9gWzeodVxAJ3Elu2uC9WiTR1U+btBMmG
j4ybCJu/BR3Qw20hi57R1UVYeLszTiRdOy9Cr9cQre7nYF3cxrTn/Znbl4Zp8oS88EWUuqNePbJ+
qiVl4VV0In5vTfrRwCC1ajdCGBSgvEsuIiba2SykuS4qwK2C6mvl0OpoQBP0G2YuwsCTXZ9XWXHo
SpsS0hCrjx6+iywiP7tk5jnqWwf2y6fbYwsdTrk3m5RevtVx/rT8QFnSc2DKiSKEfRuVn10L4Eir
eaZpOnM+fg3LYbV4hbP32p5MaIQD1x3jrtOiHpBgGYg/Zm4JCGtOFIQKxP6iivfqE5P5+CHDBMbh
Zhf3f7YabWeULYNONIVNq0tOA1qjHn7toXHyfYJFmATgwNlEtZynH5+Zvh/C4PwXN1W8wnJM0RRr
5egMjOc9LvvhrGUaEdAeumDBTTZcEXCqQvz14ZVc0Fi9E8EOUupLYgxt6P7NK/68BXRhFIq+QdjG
B45I4MfNCeYLawV04ntePY1Z9qTMDeNIBBV/ehG9HBYeL3GVOIlefEJqH/LRnaYMwVYAAEo7gjp1
ZdSWbex2L3lZhL+9q8VWJZcG7r5u0nBRvvNiO2sV7a2Kqk1v3tI3qJUkmts5/1MYMctLJrWHWdbh
d9H3SEWNQo7STVNaAj97lZfy7RZHMj+Dn7SAaTC4tZIPiRxf5ac1ANeLVKjPitzP0A90kAWBI59L
s0bAnGLEgIp0yvClZQaseSCJTme1VHLM+ThHbQTaKnJhCISV/faEpAZWC5qEeGEzAsvgG0jL7lT8
Wn3Duz0NF9bKHc0Kz3Zos7MBUBekgK/BKtCR+dJeGZqSeUDJGOVGiOaoVIXRY3PaabYviGLgn/jR
Z6iEbP5yymSJXfk95mMk0d6pjTt1vsRtfHHQhc/hVx6m5jvK3gOYx5h+7lHQPgwxA/ldd3PayKGa
Bjzsky8NC4IakC/ILWbBeLKfPq8Jo5i1jzFK1RG3FQatQYrUxg/fiIVgs/JeMEMKKLnH9NJ86j4I
/TphALy5F5ic+5vjWO79r6T8xZLh1PdPpbhyqjznt5C7FdTZ1hTDibOKF82x4+BLIn2ZHKZAvQsm
KyjYgjwNKjmTkyaPL25goKto6REbsBEZPgy++3IIZSiAl8/kBEguRBTDcMdT+y33tGI+gzcpdwQt
ykgJMJItHCOGU8R5szmkasDE96OXGvgLudwMqyzK/T1T6qYWvPeUJki7BBMQCYlj851tI0iVRnUE
61JB3TWQ3ehCBx5xeJ+XMqk+s2WA2O7T5aVhkD6be0fCYPlWjx115avENm7vCUTz5gRvCN9eSbpN
hqmPfLHAF0d9+X2LUqnxcbZ2WecRhx9cLToK0hMCjLlvYv4LvJ5RXN06w0wWXfz1B7jdYby0mDPg
Y90itFe0uRCTu9o/UjdJFREhlRBiC5Yu4uXgC3BYy1sgeO6m4I/KuiPm45K9dIpvHQTK7g3Hj8A2
fGsVZTF4yQ1K03KER79cGAkA3ckIwmT4v9RdsZRK38+Vb66ZheWnCGtgjywYlfby3uabm8xan1Zc
JQliLc5r7EusFh+3Sfe+C5m2/Tqm0EBXf6KErRHIpfSRiaIxtPncG/82zsJtaUDWHLQMJJ1oxJak
PFtnjjv96XQiFQx0KeU9BaHkPIc0opCoItsTT2W3boT2qqweyFdutaMLgPc59YMk6jGdH+gdRKbl
XhtFDEBKKFJmTa26t++gM5LAqHhfMgMen7C9LhWEv2gQU7N/h+YlT6nGw+QI8gRZmpb/3BNJhJ+F
p3Ub138kd0+istGtZ3fxnRfYdxMtLilQypCGTVJb3DztHMuijyKRETTOD+SbVLQOrm9wrSpuOm6/
23Stc8IWRB3/XXKAFLbUFexiKQjiHePt4k4hmxpSgM6Wu+5aYsECDE4oCfgAN00e/NByHd11nM5W
yNV1e+g+dHTokoxJ0rhX/UWID+YI/MaG+OwvKyE/eN/5mE/R9ko14zvCsfKPZ4V2WJ+B6kDCCUj4
gPVx0+TWiAQHFKgnnJJPClriarufkgWT4vmH0t7TT+K4PqF8hvBdyczVa/D5fb2i95pPh0leYG16
LTR5uaspMTd12aP3+31Vsd4YvrhQwQu7SuLouL5HKWkIelk5Zdfp3R1DXZ4WPENbOmRi6Dj/Pzoj
1Qhu0y96G9aWgXLiNEkviMJqQBRNMfGAQuuzWvLA0xJAozwQ200rbpJtpJA86WjOPp0dh2kzOItr
5hnHzQdLZmxdNC5h1xtD+wwphQBydF1Os1SpmkoIufChMeDnDxMaY+rpH2Erpn14KkLWu9aQfa8B
4pzkOaWBu0/Lv1xpk0R+Ypr9qTY+ha3SoThPuR1hrexc+bsjo/oU8uCgTun2CfNlgm5+7pXEHm6x
erCe5GnCVJf6zXmbrLDIECFUg5exrEXHOQjaG0qCQCrlr82puKV+bg+ZefYUxBAXpdT+6FY218Ht
dbWY3ufbNdMbifYEW5avPiHdr95ZqIDZXFcMRIuqimYlPIWbAFwKo5l0mHlNQehX/joPg7Ki/dOD
ptkZBzgeGPw0YhC4ZB1PNiHcepJ9N886t4/YopSwkkrMlLeSwc8H68gFwCKDhJGQjK1WNYcJOPCb
Z6I9Ekp+FnUO0JuhB/4SZ0qxHAQRZ4DniTuaqAw7OjHeu2TgFGjFSFegA3uUTGHB+vGzczPvgTKc
+beatpA9uMZ60+JWwFbB2LKHN04SQimu+h+lNkHHXDoeRTdx3uK+slLbh8j2Skrsr1PZMIJhv6uM
OGl1XvMAZNuP2+yo3pKilqMjekX6AKws7Ctud1rxYzmp9bM2b54cvId3opE8WVxyg1O/HheuA7I+
DQ96FbcesDZ6GnHIfvPeW0vr+8XVIkUWu1aTSRiQGLxgEDLOwe8ckwHnR1csKm4RQ2q5uHbWfNSq
jvidozXHtmx7NaF5qhgg17emGfY8IRDOqEGMhpXqlD5WBnUZ3FRz4ym9OUbnYN+I0FhdvSajzwJk
hFIef5yNLHEokyC8AKPs30UtEM3noysg/KhwzUNatNHJufI04WZAL4btKlFDlVbgiJls6So+52tU
nwy8Zjvzy0JtVfdyM2yg8IKHZZ9UpP4aiEoM1bafjN45G+dedNuwUKCcSko4xd4TU1oYZ77P/OME
J03S3uz+vsI7kCWjL8AfLvAIpA5+kO6mwhZPAEqlNSKzS+XtHqDhFprp4ck3QsasqprxrkdRfHF3
CL6qWCVLjKaYBz9Nvb3G8/le13tOMf+uL6NvRr2ADtRNCh4bQ9J9P7aoSXELO+5A7eKcV4IO7Fag
/ezoSG2Shsxl1gmaXk0pKT+SkTr8nO4xwbWihvFMPtgdKcYAQ6m+5f1rn2RbxfkqIYTBa83yf434
fh5BFi4INFtjnNX9ZHVxDF+6DA/9YunKG+AlKhgv5rR/zengrTakxETGMd4gfHZvD30VQsiE7ykv
3Wfd93q+/Dvs70e/dTgV3FeqqPLn3yp8LIpiEh07pgQCB6Riwr9rbyvahZaiT28cfOHFVWPUDlk2
howDMUnG59VmpIviG7uTg+RtTCG57nKO53GdUHZr5M0IUo/rsrAOquS3VAn+vchW2qzt53QvBztP
/QpYGZqU/pcAwdzhkOgBOTKIdnnjo9rSzEiGD7cTiVB9Pje7c0flA2ecXDWiQCKWmlUJ/IhEnGsK
waFd74DPGK/ef96CJFSp7r9hq+kTmT/e9EG9DNTUAicEne2Z89zV+5U0w+CX2hmrYLnOFERrUSpY
dWV7CGYbHPNIuh2h7jD+pBKmSrepRXK/TZGjEOmEUvOvkdToVi5AUaACQalUDqbrgTg1xSYLrifN
Q6U9Qff7wLwfpP2K9fMftUWH3IZ4SdTgsmr3MC4XASAIEk4cZ0trfDy9SyMeyhjMU3iioBn1oca8
tzXMoUr5sQ781xuwPuY2o3fGsVVG3s5ABpCXu93zm/HofsWVB1DfVd7Yflb5sCkXdviRkeSTFh8P
qY8Bnw1cjtmfh2GjdDRTSHzw2mpOsZKEVUtsvk4S/wYX8R8W5Rl3ifDFj8Nl65M+QvJth5cYZ1vL
xLRtUmEG98PefifnyFSfX79uzfsvtPbAjkqkzwADxDg8g/kmgWi59xphD7rjqk5Lm1oHmRSi0FbO
hz7Xog9k2BR02N14RQ9Qzs0ZELfEhKW9wYRuN3m5k/PKGm5w2MzUn/9a+4wiA1pdHrke8cdj9PTz
zDJ0HUdqYhFZtoy0xKAiegKVO2/slEa1nf0S0hltMbbn5RvhMiccN/J5Y9FEVQyGa+rh6I3ClPS9
TonGMX3Y3htMW6TPDPlmc1NfAxLzKEBhSCH3/em7hdo2j15z85T7xge18QJThFbWJtz+83VaXhRK
la0QvuOHqvng3+x2oUMUC8ktAcbqcHAu8IcGUPdtsM955kdxNVkJm39clqTC+HQhlXYwyxl+2/xT
+2AsJp8DXInBW/Q2Zh8qH+VQg7jnirPP/tVfRyl/xMOVcYMYTLkDWUJAYJAan4/0xHUAy35rd9/j
1Xx1+G99Pw22RtIaho+f+xfvjVqHE0VC1zo2R5ztZuQV4T6/1wRQrTRh3DefGAz/66rea8a/s2mN
JpkoJd+XKX2xJUaKhG+XpdVUdJv2d8gLE8ol91JMwrQWw47T6y/EByXLg09v+6jVMKiKuAgResvE
CSicM7b1XEwtdxHXIAoY7lg4W3mfvNjPmCgaJXx/3OiGgm/6V1gXuMLZdZ2TX3L66F3efM94nE9s
yF7fQhhweKI4/VEouQh+dRe2+Vex2bPek3HvXA2ifl7ma1v88XB0144HrgegKA0bepkgTIqlAlve
/mVUp3oblQoQLcwsy9vwsPGIqgMOGop/QsEGDeVuyv60vn9VQZKDqMo67EZWBAb0VRzvXKwY5XOM
pPzkNsRhd52cT8U2Re3M2XTrDJcra2U8oFgnxlBRSvW223gZ0Yglf5AxXtXcgKDSNA1PHIcWWPMj
QkFScOIAx/qrx+OLgovyKKlBiQcSqzou+sa3samlLTgz2y/FToHVUFXfUgkbvvy+RGGcx+KQA3VF
/elQtb5H0c3ZUAlAW6zEYSwoToakz+dkoNDbWUHyNlrkS6ykmu79pnMw7ry1SqcgU8kY8xJMf2NA
kP4AFFo0eU11Em01Q3oDG85qUDUTQu4YdTYTCFhpvWEWaeIx4Sh57ohQ5Yp+eKP+fxxD3WxBQoeX
ExWFOzvKwMWuapZ1QjnehjFUi1dM/qYYgyRuFcXEzlQnq/oNAAMi/2/NmFZLWsmoCnx1q4JdQ8hG
3byP9RgsWy7e7cos8IXtSPJS87YSmKd9P8o2ecPptspPrRiIrGfkMavCkqb4gh++MRsfS8tqAZvA
hHPXJvyHh8jzNJOP1FghZTzRUmdYAKbD9h7ijbo/BzP6a45UEcq2pATd4LYBdhD8tc0okA/xCRbd
BAHJ+zZJZg19+uQXvUZ+p7gYCp3RbTLmVD6P0F6sVXLAX9xh6p/0iRzpmB9H8IlFGcPjPFbD2+S6
+/WtBw+Lj+cUfQaAbSD5221txAuYQbCi8kZILqF4jASpzQuPRNo/vO5Fa6IukqMrWdDVkKxqBK5S
5Q/2uYneIlCp/Tjez4NXFI391FornvgDnGZXjXb7lfimyrZ6PNay9pYq13xFIE2jYya/xZz7WhRY
CquXikHcxq5NYRSvb/vJZaQu5utD+uuxWm4xubY9d6/CF+ZAa6Tw1wxGMABfNKXAF2R5askHFD7j
ijbq6dL9cgsBb/5GlBRD6XdyrSq6KQOWAP5kG1azrhp1l7hzzfuSdFyS9ns9bzGwN/hmFGf64KZL
Lu4w14cbRlmd58gw6cJpk3XujslOepbvf9jtx7J+JpZDf30lxh0RagN87rh/yweVDHVTMZ7Sdo+k
X/va0gVtgAiXEl735nhjEtNarEBVmQtIXNmFTRZxwla+509YqOCE9YH9lmdk2rWCAk3L+askqxTV
pogzPVEi79DSVN1Wll9uGdUangukL3/x41dqNEsfR5WAdkDRAmJ8ZoWayTuLJAyx6bOWoFHxT45+
Hl4+qsMxNxv38E6X69ZGy5NFG0AudgCCvwxuchBnFF7J84nEvAu/SYOgQD7CDIW/BKlUMQkLCsd+
1tSG9o7v+dfWVdAwARUphDPjJDAVi6/slYClphffSTTF/Kp0aCssudjDIyT7nhNBOMGajcHcWzLq
ZIXyPjgcb2SrZYpnua6RUjFAlYMFlxUkKal8eSemkb4g1CO8VcyZeieb3Nr6hoyPCf9C/CRiZzwj
4lWJHHYT9zuRdjtY6491cE4UKUsmLKXTwzv00WE0TsxX1mNbantggR3MT3EzuoPM4TbRQh5oCGv1
FKwyJpKFlMhnFxdYSRdTaDNQIv43CsOglz25hdc0g9Q9ZTXtIYzYwcRNWe8g5+772p+lR66LMAMq
0X5fatZJdVpu/eIV4PsqkOAcAbsM+yLsx3ekIR5FebTOc1A09RuzPMw/pzHvX/NmocO/pht/bEDv
PcJCkhE7hoMNM+t7mB8TnfrZgQEKAEtBFiqUuWTCNb5XysRG3P/mkUonq1hiEYL3hfxev3ZiMb4F
2o30FwbybpLdH8RVeJ5tejwwlHzw/a8qKgXAEerVNDxDALahsKtCkFZ/eVrHviwuhWMcf94xyKN3
YKZ7LmV1UedaKn0nkbHm1KEQVRne8QuqwXZTahjoJOklcuWPffqhO+YdVYfM15iyfNKGICbXIuaH
rfvqOL68aCvhH2SvTWn1ZpNto/jprU4u9lWGrmqPrvMroxI9BMMs5XZm+s+xEd3wlhugP7Rcxj3N
5DpaLQFnvRTU1YT9EW5A7Pd0Cy/LZbif07ntkgrXHRtlOGhd7edokdXpx3vWHyisFm3umClcYz18
6iGO5z5yAnjF161O6angSpBJ1ZLiaXJBZHBCHvd77YZ9WhstuD5MFSVbRR2TXEKYv181ciFoyzm0
mu2fv80DzQI8dETvQ832N+/Ehv9H5C5DNJ9NOEHlyBvV2JHSxFgOlftK+9u87yWD2G5VtIfuy29+
e50Turt8cZ/2oAlkkoVMMbbPCLib3OIJl8I+6sgJm9j4Okyjkg+Lur1ccv5J+QKc8cVCJHmx9LxJ
J0N6Vl4C2ciTHJuC1pwAMCqEI0O4Hgh1p7pKb2mPGVzIUlxTdk6FvkFu4DukLErs2ApT6HMLL55n
jE0Z6NPQy3OwPy6+cMI+OAQ1+IfMQq62l9G8M/OuO4NkR7ZcaeZOCRso/ofd4lD0KutL84L731I6
mgqiQYCATYVYZPdvC5oZ3qsklI6bd6SEunkJZ+ncX9slu/Dp2k8TmASRTQUnvcsa8eeiGE7ea0xA
bPGhlNmJ1YbjeN4P/uvGfZAMgJNn6WQ1kchw6HPGZvWimZd9MHAZdCjrp5hIRCXhPwikrhy+KmL5
OW0NuBMC+KJ55Be44gDBPAGJlettCspggVJwUw/bbwAoTpgxsSsAsYiCsonqqtMzdnIxKWMJsBOe
jivSphhNtIV79SrKPlAmC4peJxx116KFXbxZGYx8XUfiN1YjZVFUmqwYkXxPkItFEQwpWez06mCf
PudVtxIh5p+KNWChU+t5Mk+RsjwxxjX26AJTk3VIDt48guY7WAlXfozxh3BDVe6l4dUL/HUofmXU
C2p6tflCmybJIGLkL/asM19BguOa8HLIG/iWMd6qXuVMAUY4nsfAsLaXjamt4hk7FH9BsOBlohuc
JdqtzmGqHdqkf5cD7kE7JfwN0dNGfG/l4W2bmiAS7uPpDL3vbPi/guAE3Id9bFJPSeb1lcM6n9BN
cleACW/uAFcoe85EKJHKlIvx1s3SAskp4bOLQ3xz1U04CxFerftQQnlIyv0fkZYkieFBb97iSjWt
ciqKNVv6mCNU4G2rC72oCJNpWbkOz32ihzZxn46v+IEoBK9uML9Ub/WYt6TV9f/jYowVPDSnE3VW
hpUWM7GYadhNufixxbvjUIIFn95JO5Di7IhkCGpXkfhE4JJiElRomGMXbrpOaeEv4RsYvlhtt4wc
UhmWvIdxW5U1aTOkSHG6wOPSbrF+T8E1crDM64U7723/DwdP6ud33epIdbLJ4djn3w7LwnUCHlD9
1X60NASfiQS2wlFSiGXgnAj6VVlaZhtq3V5VhzfyJz7aZrNwuOIRRFOul9KySjXalwRSOUMWMVht
j8RCceIWo3B/UawblNmk1JnLOnGFPeSaX7wbtggd+3pju2H/wLYZ1E9qHyPNeRXxcwddX8ib23V/
WY34mjTeKEA9pmGl5w7jgfLEbzDAvwOYU1cmpCMgbiqp6/2BNP2xEwQF29+8R28l8Z7opKV0nwWt
lY43cTE2flAVb3sQVLeEHNaZ21/ivWfhsmJ3Kmzai8Kmc1Rvp2A+hZGkHJIkA1npn3kJ/eJrLrQe
EBHWJHW0VbgHYrsVR358UttRug69NVKm8tpBSsipHBgTRraEL68iMbp6YVbRP32S2lx+/qrX+/hp
9eNsaHXMqbTNa2GCf/T7Gx8+G6kRueFrNGYyslDnVIDy5cvYHOTV8X64HHRStsvybK5BnrnQhJab
I0BKhPzB+tbOUYTutVGmyn4JhIS+zPe6Ro+0dziIdEH/ELJuwomHmfiOQ6xVuOToY3jeFbL3jmU7
5bNF32UP5Gvn4MWf47VBpoXEHxlMKzAS2Jsk+irEb6AN2SnITkUStsrFqZJmjZDMcRXYTaWEcKrG
uFanH/u98CbJdg0/P0GSHG0zddmNr43QsJMo9ZjElUm0oJ/I5yls30sObGzY4NuC+XVYHAe6mqxr
ZOgGpI8JMO4uT8zISfb3X4HKBrGpjKVr2Skic6YlK64ORCdbwNNWhzrsJ5b+LxFOUQiA6uOmgvII
XV2dpRb+G/eZPU5Vn6BTP+36hJU5B5bybwyWiOpPUYQ13l+2m2s3Hfw4M0qLkaXUh/HP2zUYcPBW
gjgMB+U/eADQLxPdboWhDWWrINAUfkGHQ7m0BzhGDFhW6dyvb87SIDuUptT31nslTuHPI2hLmsiX
KfeJVMGOCuso/d58DZBaNDMcHGc/Q5IZoFHSTr74bNyafp8r95vrB1oRtM03PHaukQtN4CDB2bgY
MLfYcIwo5OQ/j2n6Ll3dB/hQJiVCHA0nJUADCRfE90Z/32rzS2hCrejgZ7VqZHbrFDRiTA79eevj
75ZNrNUE7jSQWtIhdAVYR5UhMhAHhKqjfDdYu+LDHsJQqcZmhewjKwdeBsAV2tz/8Gke7iXIgplb
ftkQGXGNDfNiiX+qhepvzl0BWUIjBNq857em7FeO/v0db24sK5czxyOwyAlxbEons/jEDSuej9PK
Rc8DcAgZ4aUa9e9oK8C54SnvxSM5IHwJFPD30rUWvQaCWrAC+MWObCgJ0LYCQvG6qI2rHM2gM05U
dL5g8YJ/Cj9kDYzRv7ol8JtbvcavlECcBgFOelViWZC8/YtEcADftMCEE+BJzgrq1bRU6StVrfVe
nG/yfUF6lWMoUF4YorvAMnjZB86gOUFKxaiZA2ZFI00DEwpfB3EU6nI0e7D2EU6S07iJQLdZhrXq
5q2ZsMA7X52Iv7qwoGYXrp6wQ2AGlLYlBd3CpSDw6Sh5o2uhx3D4pvbSBYdL4Tv5YVFQ8x7XQDAh
tjIlBSdifsoFaVnMdK+aa9x7G5h505gucPhEXn63zVGwuR6FKogoJGlim35edVYy7KYjcQ608maJ
W8/mqkL3Imgijof8hp2t5GEoOi+AXDd4WzT6Cc/euk01ej5/m6INZv30SBTCMF1JbduP4KIpjS6T
YjwZ9yoJjqi2XN2EWxjFi/FcctXbS5eSrO/EaT0lSxLjvK/0aQtZ6wWngC3U4bNb42EEIwIgoC51
QbQszmNXA8ZIwkPNsHZ4XOUbr/gAnpoqq1ktjeA/tZc0hzbu9di0zfaxExKyZXfj0Nhvm4U7i0us
vKXi0qnSXCQ7CIphvC4Ka3Kbovtrc1rzgjBdw/qdNSNvWOZZI9+wUBPvRwKDIrKqZgk50zadZpud
qxVcIM+aJzCOjZAsy+LsPIR7L8B91ONv2Yf/08vdKwf9a5IvEwdCwI3RRrKBM25pxKpdfxl09VSq
N7+UsTQ6vSgFa3iMb3HWX/hwH6fmBZ/SkTt6qaOmGgJC4S8GL/e/KLF/bUg36l4GZctxlL815tR1
/vH/ZBJCNaCMewQNOEnL/tVcRv++UNiguK4YBod7N9FgHLiXwJCxNimGGshEn1JdxUylEBX7KHwX
PFXutcbdon7WTVCMem5jxz8h5qMJ8ecyi/B3hbqDYx6KESIPoFyh2LzPTiDGcFduPIdLvoTxQJnl
KCNTJ9AaJ5RqjuTiCzdIL7VcM00/l284ON0bjYTybuI65tI72T2k08Ik6SBQ6Sf74ilHP+ZTlQMh
SMDUqL2v15HpK5uoGscUBv5qPOFByHEisWLUlSgcjPRlztwriohUftL5ACqCKtMn9gdfNCXrcLIo
GICXTaeanTa0z5AEr0d9yZGyDDwMVsee03G3527A1ucfpOpJfiBwGQkXzTFPQcrLZyWl3bpPdwHF
r129nj+JxYcBy9Cqmgywebc3FXuRy5l9+2gI31zlR2WEX8LT+3ZyaV2aW+2014FxDqRshh1e+IHg
QFtZisePyBKVxoxxkm2YMp8mBBYzT2Iv8e5CjKhLfQKteT5rweP1gU+0qTKLB7w+OwnsjX1Zs/CG
yHw+0MKr0z2be58Ksea/FUkP7/Ras2bj4SV5DNHYPBvLpybyWG+7u5+Tdl2fy8aaKZV2tcD1M3GR
fSIXkDmPF9KlN+AkfqejeUcAUGh94fa9fKfkKpItWws6bIhV2/z/I08Igtz0FWKFdlGuF5oXGiXV
rnDOM6sBlo0JBWLl99nRGPlkPchoigSCnIGlwXMFry7n85EpsKMWI+eC21YXGTHj+AJ1fjAPSG9q
iqQSAyyHC6IxNMfV3soF6kk4GFTJbVvgJNnqdGsiaDu1/DRwCUbHNL6RTU1s6yYCuVT99dxL/xYv
BNoSJEUEfQsjgfQXsjkmGsa1cU/DGT4h26+EUr8l8mVCUjVhMzDLImwjPw46A20kOlBVz3eSNDqK
9CW0/Xvs1aFc2oFn2UhvpztxiLflrthFGjjC0AxzYPM55ZqIBz97mTGh0TBLkQtEofPfhABmh1nS
GK9IW9iqNDK4GoPe0HkASj4fePJcbdB2ACNOL/qeLsIumYlF1CtkagieZneD75BUoUuI5rlmco1+
1eWOLmHTORAFFmVA+yd87cwjDWjU8wRGhj5nyY1eKaiS/OQcttRA45uuHqj+bYJYKpKgN0Mh47HQ
ku+SQNjkLN6IsNu1T46U3EsaNBVKr09PwVPQTXQBypc2/kVgoTsEQBiaUncawsM2qlK7pj5CZCEZ
BjPAf7tCgEV3ndoVo9EYCjCSp6n87H8pBb7Kp/MU/QMH6w3/e92V5B7BvEk6/WKTc8+5/Y1My8v7
Wd0yGOkqJDkUMEjC+lXlh29E+itTNYQTAAUKfe+EcouTGS/95ZCWi60mzawYjEqf8uXyHY8Toqj+
qXcpSoWAhJPNxFkKjNKeutPwx1bkzW8osDJtaMHYUEpDo2V1OEzeLE1lzXEGg28xSTPZg05WV0nB
gVVlEiNdslNWbm2oVqxPgqywTCarj0bJjBebXv9+ssBDj7jQxo0q6z6IIybm2yZXsLHDV3DcxmLM
LOBEEL0WX0E5NYkqYJcFNyYR9d3SXZjCCONcPs1GdsDgFPhJs8XIFfnEjoJbipJRrxpx2WOIftTE
E1MuxQXcbMzK7usUkjtJ58r0z745ak4G2JiPxY0W9SYt7Ei29HqBwkwmmqe59BatTJJFSjfS7WAG
u0XZW3HVFTNiw6d0C3eiiEyJueU59Wv85Rd+9jU1rTumL9D/MlEbCUA9DQsT9NqaMOUloPlcoLi0
mqb2WCVD/52oQwVCO8Q2kd6S1jonAs0X4CIzqmeOtY7KZcaByAXAIZPLzR5u88w3aR+HMnre4qtz
OPCWSmi8iEsR+wmvft10ckn9sx3aztUB5J/QaBGyHrRlhppiywU5GzKYa0ITX0WYgKodUEqc1N0Y
9A/u16G5HmkXI9qG7a+wH4TaO2tYy9v2/W+tJWoja+K0iiWwL6FYXGt2v2Yk3qlBouAWc76QLpVN
vPtxsNahoOVHIwVC3CkvGQIoLPPl/Bir9+NW4dV2SrSr1lRW5T1OClI8/IcMIhB3pZGdeyaaNKog
Yg5rtGlQHYl4nMFuTbtf0TE1znJQMzAHZHcEFZr2qSX9sfKbYEauZwhuQNnBdd45sOcJGMim+Evr
6x7KFYdcjlOzblCIWwbcTnz/ywMeLEx944ckHlnAEGrRQGD/OX7dgfOHHT5xs4DabwO6fd1CGnI5
EkgPUeLT6jOc5gEzrajv3oZFqdZiTzazpT7FiNqO3c73Wu9r03h/LP6O9N6Z2I8lXBODp7vg9wR6
kUDYSPv7baChau8kcNahsKHoQeUtrt8EgpboHT4O+lyQ7PnX/z/SeeW8r7LglanDX06n+un9Vwyo
pOk3/UvdC9W8bn73ElNyIgg8WvyUZT6+DxUqBpBM6FhljHZD6fK1Oim2bDxIzWciAiaRyYuXz3t9
M8I67xCzOBgjOR/NRsHvqjeGAgtCeFB7BZyEROlo4WOGPwh3mTULaJfEfRdm+KOOUutdu+Xc2sfO
4lWzVqatsmoig93DgIGaalu2hduBNBBTSf4ZJfMzGWURKmjvKUN4QukIeb7iCX4jdmo7AQCvNPQM
crSP8F4QarH8mVhj2DPeBJYLcC+RFI/wBVZNaMdBTDt24mEirBrc+l1RxEBzExj8dwSFxj5OuI2d
+bhz1T2d5dHNhHvpx8OsfaWy2vcInna6+x6pYdhzYJAtwBi52l09ZsZBBK9V7xbW2cnDrAz6AoaJ
c2Qgt0c/94MGO7RTBAgxAPmZ4b2KwiWweRFRnceeGPafNTqO+rYvh5I8MGn1nfng2TgVa7RDxCZw
1rXf29AoKwzwfS294KViP8LvumPHjY8kHfa33MZzZzHT/O+nxZ46J5Op537wZXtEquBKRTE8h8Nq
KZ/ntvrFClIprDGqXwo+soLIIPENEmEoVD6SgFDaIAkP5XiTdqlhClIiwW7QjryJq0/yrDTKmNHG
N9I0WvTMK1bD6X0XNYEAiq+680C6gFnTfd/d2F/hDi53KRqyEy08cV7A/ssI7DuOCTv6KdT0CYSu
nJE8KaXGz3cfpP0a4ATe1+Kdzbiz13NqCt6Hkt01iaTcYomiNZ5lbmWjPSKfA/5++l5AEhkFAFRn
oTUEWDRZjcgkXLWQ3/6+W+dsEmJpqZYN+B1Rx4jjqL1Fpa8HG+1RZl2ccpHeV8m4nbZPrsQ7OU8K
uZ5LAeIk+nXGQc/JBYONVt3Y6Yub5PZimYQJH7gDIBvdA+auKe/6iggt/PBfC77KsVvGmLtByA7K
pIjm+VVBgyxEJL8XXVRZMLeK0kMKom+FLaWmCOHcAmmuNBCC6d0idoZn9x3GbEp03zo89nG5u/EN
fs5xhgQq3JxeR6Jrg4i2wF3/vRN5vMH4wXnwEe+7b9NDrTairNZVISG1ISi4xS4WemkPjiifaKLB
VSdOfC/sxvGdEsOQmuFgLbDFn9riQ4tHPyJhNsvE4uOUoM+e/6z0+zJSRtE6IXXY4Pi/nuXoIvy9
yK8puUK5A4Oh6CFRNoB+WDP+CB8BFtsJzQMr5PC/LGn+2fkVyNk2A++00m3pXO7DzlJ6CaBrtX1i
JI0QLs3gnCqaTQ99TPsP3eWC6y1yPuk8fyGmJtddyKlQyItUtqeSOWPAeGnPNENKCtGoAKmY0bWW
jtFCpnodpHxQ03p5kShiaOw/ZhVyTEqA4Tk4qe4iufPf53klJnbHfW9GKRx7tKYw5K1Rp6EK1TIt
d9W+4oCdTktxHYoxOh/LznthrSPw5E0C9Nnm5T04PhkAw/EvqD2m8iNyAgQ67kyMyJz8bZ3JCgyk
bPTLbaMvYB5rYfwj+beS1+GWm+eZTLEYPD+RFtoj/NZroQk6IAZL2bNRaNHKIdCro6A3coqHEf4o
j/M0o7jkbMBq2Xnsb6i8/XP138aefMm48EmLzfPTesfNCUEnNlq4GAddqjGMdC3SdILIWQ99by3V
0XQGCPkSOHLKF0MsRTlD+rj6LzkZ80X9AMTWyv44bxf7uEm4zsK+M9n0ZHNQzgUVFlPneQySPrgP
vWOnv5RHl4qYSPQu+Z4CcvbkABIoUHYAmUhfRzMwpx0chHu80TVN5vk6F5gmzC++D3Drn2kSScKG
Nx4sVRR5hqYSVlXYN90uFkdHjXBmH7GFe02zvvDzM2aFLdvYqlDRu9/9XjLe8GIT3LOdDvx4Nol9
0OvpqNXMFATlxoMQRwh4+DNT/zledYsY7BLlMX6zu/rcp0YShEgxFQCjWGCohYfv0DlWsG9H5mOM
7mKpfbCPSqkAhPU5tgrdX1o5zNREABU0afpEPKwX9teECsXxVKu2GNwzJS454841/zKAg75WljEN
ElkUcohTmprneTmVA/Ff692i/CAVbPEWk8aqRIxX2+jZSv04D2QobthCdR1dDGpDi4qEr4Gq+2Dh
k1LqILKkLbj9C6LIG25A1AYwRrvpZt6dG9Hj5FE5N+OqfPY6izj9+2CM+y8cGfBee7WJGKJV9iWM
e6+o0NxSIN68ZohEuvusnM22Kb9I3pZbYc+6Gf1jZz/hLBZO6nIk86/RYcv3AWMBeIyaQnHNJOQT
BymRXwZ4DfCftYsDa9ALeJCCIRkmZmuw8dcoPB+CgwCjGGZkI0uRfj8ov/RdE8/Hur/3sF6wlpFG
pmCrwCpl22XXKbno2ZQH3EjOUY5w1YBgFktqkQReEfefvql//5IZXCHLnKAtoet++uAOXLcIkb6X
8nPJsLnYxgPSvqxO2bUKOAqp0eK3z5GyhBE5vi855s+vEtNR63s1Yjs9H/noeHPkVjM9cn0ONxep
5t8f057YNHzdebWYu0VbsNrDeALoH704WKU0SsfwgvbruovC37ukOP9L38TcX0U7vV/5AydMGqDe
kFiQtBauUtuStkvVqeFu1AQb03Gc/o9XZYhRkWDhQJxDQpTOTj+UR04sAzKMvKP48qPHcbeo7a4f
OYLb7WWYx1D0Zv8BaDB8C0fG4pz/eo1IaxTxJ285f0k/Mp7ZTb4YFhE5ZOgas6+huTIaLB3u1EmD
sAWND3DqZ3KslbaEEgj31iQdHHBY1rTBvrxsV6TW6OzGvGpdkzNQllZ3H6XXFn21QbTHQERbVWQI
4LzCPj6alpOZ/Xd8Z3kiPSnhoX6MybVjQql5O2UCfue/fo24YhAExG08zfoOnBO9CeaLNFbzkcEJ
yJkKGbNwknixSPrymkWl0vHahQ4liv4eOaZSCcwFXOLc0mUlrPYGWR150TmN9AiMvwSVChSh1VyG
QmwWaSFokS26q+ABOs0UtVyeaY0yTbgXZBraO0+LmJ7z4iOlYAk8a8IrUBMtXbXBkGz2XQ2mPw69
XSPCk83jqR5AT3ipe3zhcHBnMPvX4nGrbcsnwFp+nuJ+QQte8hgZH8lb2U/YBgULo/8MHioAuGLd
MuPgEDanGp/i7PwrdoySI+N8/B6Z9FLuoILa0N19BOA9Yghpnpbyxs+I8cm2eRyQx5GFpJBbTpIP
HZktYtXFHvYm0JV6aLIYCF1CmkEQWgdtz9IbKCU0PMR+76Jdyc2+cU0sDg2fCTzWK7cf0WR/kzQa
C7RPvV0viSwdQAy95webH8RlECpGqEwwSnflyDtuC0B/lG+WMZIEnxe09eeRtN3wPa2LVo1c1tZq
7lfaP524igl60WuxOedwGQcktez3TT2Gh1rIF4UwzrUGE/YxM7nKyMt8QIsKpqHLKtFlOFGR5Rx0
Qe/epwBm5gmftrO7vad1pRas/lMHYni2+0h/ZNh5qQXusPp6/q8bKTMsAkgvdHbyhOnki6SbKIH6
+XiepEWhLaq9PykDW6lEtim68ZOBcgUPRcM0O/Xn3redk2gGKoZtG3MUlwSqDrxZmA8fftzMc3/I
QwWKJwkJdv8yJintwhu2a1PfVGb59+/dQUeViWKXzX/fFNKINuAj+Onh/DLl67S0dJzkwLOS3WQU
aMXshckHnBB7MXpYRjOam0UqTehfMeSd/nBIF6wRnGqLx8Tu4WZoPm7ypxsqaAi187Xl4IISkVpA
vlU6r04LcE5Of9Um0IGqBv8jqq5LFDW6sNVPVOm6u/Z47wFock6B2n/h65loB+q+Dk5108kYw/Ta
f9Y2KiqjJlB4aHtdmNIclxdTCI4vgj2GT4JjIpQN+q4RHTH9M5LFZ7VLjLYtFt8UK4aTGnyxfvQI
vk+hWwsY7yhrKW86rFcZ7pHnZZsh1VZc0EuVfGADHmAMOhRC85AW/7geXY8DtXdyer/GVuBmwQ49
p8NcRbyjJV9wqIex0dkBrzmrP8+UV+wZHWU9o8E3DTRhCiaFYUb3CLQNuU/ew+bM1FAZwEsd/URD
VeKR21GR1bgRJrzHA/LVhWwC7Or0Cqryo3l5sTyBxFkil/mhV7cLae9PomGogXNcu/5UINa35aTi
Kf3VXBgYEZZdOwNI1XJiHtBJVWkn1bi40mwyeGOrDq23IPXEoIgel+gGq7OJ4bD0cXJWYRcKtZ0M
U4qb0MTA9YX9k+oAFzpAo7VTW6x8r6c+gICjIDXeU3x4+25UPbjV9Ggy2I4BztrMfLykduIfj8Nh
DneQRJbIUTvpJCydtCkhyMIXDMPoJoJBdSvS00GX+YuseBEgQ7GcU/DfiqSwUsO2dgBoLfxlNF2E
ZgRmot9nonWfJAl9dh4CkL3jhaXn9XAQkOVJuo06jaRID5KoLPVJs+zhfs0ijZXVaSxhEfaq3+bZ
XV+4keoURp/rBap+Fx8wQpIktKn4+m4LXsS1ZvofvHcGUHKDBRrdjPs6VIn+gGqXYZPEKadAW8Zb
7gF2Gg5YE+f7rVS6rtVG/X3sYfSw8JG9skRbBKJi1JTcWZicWYopNgJGPVeJzvo8RCRYUIVp3jE2
Tt2yLwdaKM8KIuiiyIyJ317RWV3zc+7+2KhGZz/xfiVxlYoxwQBockqMW/bUN81zfZ/ENwRY7bUD
MmRt944zbb2zRpP0bdCvDYEIiCutY4IJZMKa/+TZeSL1cu59DpW0DXtSUWrecYpbxAt0dGW2pfD9
9AJLZI0p9VU0a4e5/SRFTEaS90ZbHjRUfZkdoa/E7OQIXJbthgr3PW/pcMW/9PKlU6K/LiyzA8S1
PncyWxZg9JbheWs6J0Z1g7COWZE5YAaN9cesM/lNVWndr4JziQ7ezrvJKKDCG/xfMOULLatESCBH
N553aI7PKAX17y5J0Pci6IGbLqimD38HnALMQ8lWxJrL+3IPnvd9MjhBF+1sjcuy8egkle6sf6YT
nmnw2Glz1WUQKtvEJAQJ4OAB5hntSDDZ9wXaPpvCKWJ5seoEjCuuNChM7AdZII83imwmhZPzaKBv
S5dU42Pzx4e6QjSWC3Q+QhHbJwxlDnC3xcGamiQS1i9HAC3F52AVWufhrzPL6ifTZ53KrrjiPSSX
jDpPh+H309s7J0M8kMathUuCWwP3KRHq+aIsRnsaO2PafYPHtD5mKQy4lNlVQXFDWKCkpEbL/irT
r3Qn1hYj7o+jLc75K78MTFEArgOL3dmJXhdMY193sFr19/BSd5Bw0eYFS5jsAHjGqrXAx/TBLX2n
qUB082s/jK7vzruqtmDckLAGB2LdOmcCfsWgINhAY5y+W9dJ40EEQ1L1RUTpHj3z0UTsT1OiKtfX
DOuyCcM0gtYkpkFzUNfQeEy2gEiuWISlji3QlX6WFc1cizzcUsuvnNTiPC540rrtQs3TOGTbSFef
4sT5bxeuBx6LTSc3/WHnBFomMj4e2HFXjUq1s+le2rZSEjF/OzV6ADQglrrUdM9z2gm361UFiw9v
Q2bLo2BxLcK7YaqbxiZ5wfJsvlRBpmWhY+zHRXuM/OJhF0gYCeU8K+Pc4z0C2jn5cbAzKPV15G7T
zX0y2yd2USG0KZxm44bpMZe7w8Brcm4xOu/xqBKgptRaquNydCGjnLBEL5usQik/fC/cRmutTkz2
tdwiOdxALDsYY2jY7DGnTHun2MBRO7fNSC7q/GVXzumPe1jC/bHUkvZVt80Pz8EKUyKx85sK/y5w
asuK9JINujLfV2GKuz38qnf3f/V3QP7H4yJB3EERSUhjRXuTleQfiHGoeN1Cc+pI7uj84qBVgJzH
1dnTirDKRzYtNbEKsniA5gwqoeyoFPuiI8eLxUe52wAjBRYyLkr5ZJpJpUybLlhtqbrXQIfwAs0x
8zQnQSwpNeZgXXdEYl46QUbtzwL4mct/odblORHugGSOeijL1z7mlzZ0m5WZfSlrpncBWs+RUDfF
+LbKB/MWxNyf6kVihJd2CINcaJYD5iqEk1lGpDkhWJVgDwxpecEJmEWhkqB1sW4KQ36I4eDIFHqU
YI9CBsqe1DaENrqJ+2yWaFLFAay858nnpoQ1axTUIB5hOqRWrDFjxBfGUZ+/87mMPhzVF7EAFObk
bLHPO5IBnhPTqbHswOnEWev3KhGLQ0DecLcaxtvjEl+3oYKTGgh9k6RCbhg5kq7uojXCZE9waaWV
3eX2hXvsB7661aBGT1e4CBBjIabh78D10F4HSyKvW+S34Cu/yJM2lATWuiDtOf29f6+0nc6mubV/
wQM+1u3A5mzzb47QUghbj46ZwaMIVE/xIcr7EcH9ycXhUI1crthOB4chHd6Mcw6Ibg3q/udIIkRW
HNyi8+YHs4hwXlisemYnjtCVDD8FuyeSq/uw3dYU8RzvJfVwPp6Toc60p1sTXNWBTXSdzWsj7H4b
bd2fsF7nZNNudIUSjriPEwBW6E3DMKT2DdvFOpSPNvN+pK+bPSDuHNMP+lnS65lVzigB/9h0nOl6
UqpwwzVd55qVS9y6k3AKnVvpQeysnxqBB5DfhVFjOGAzX77+m9ZRhzj+tzNsCMyOh3M/O2aYbbLM
LC5KXpkSDprwfs6AYTqwmvj0WAb1QFOOV/uprk4I7K+DeIwDWKuYv6WWb1K6n0S83u6U05JG+rf7
2rGI0Mf4TOqqHnFLUeLc2sLo3G18PafQAFjMG8ITEyRL4ffNuIFGcF9xUHVtQsvnmWOeloXmXrUW
Fmqzr+1sdpWMuLD4GJ8ETxRBFHslTA3XNzb+vvR8n6rs1Dw2aRdA6RoNPUNCCeaEMmFF+PxWRFOq
O55zDRyu+nh4uvTpIgDz98YCdkW6ZH79t1wvQozgnGkmoM/RGYjIq4jgA+wtk0y0EdUE9VGAaUNv
uzFDl9RPYfZNtkKNDL/jPFMrqh7dHiPAj/5Y08wcUvLy3CBPyX11t1BpWXOz4j0UX0twfAi2it99
uaBljom0SbwRTUmRKvQY8RTxuOrCwCVGZh5GT6CjUJxxlBe9zLgiMEc0F4sxUtVR42A9tCYbdWMd
bV3pqwC1wfaKnJ5rokVHP8beHDeBl6nUUWQjLylgtzj4+Ac0++6YDDcwq/oyqbzATTz1v+O8fpd3
sW+UMjCUnYNp/ckY1pdlHDSr8AqxzPymETm8EBjkG6pMx4tN3+GL/xOUT+572audz4VVcfkL0JgB
+ErZE0O4mObEiXkXXUN3tTs4nET9Hvqk3RlrwLODHJk5nOGsR9Tqdp75wJ+0lsk9RNpQW/4dWL3M
AHKU9hHBFlVDl5rHseeP6iioNva9a9xJEbfq8e2pFNh1GXmonbK+0oVOxSp9SLpXu00AoW7Npidi
ITpzvXZ+6c7Jz3HWIsxIF0xn1uJurY2w6ZcM9aRPspB3aTodOvJLZ28gJaBM7smwNye2tunfyujS
qA9rlr7m5qZq8LjvQSuTiL3w9oGheVc+7uC3aExOH4yp3hOTmO2Oi69dIOA9R+t5E13M+jvdq/id
DgHf7YWIvzpK5YeqcA1pwnidpxrFU6+KwskDNfbEZ+X+vjZIgBax8k2VPjpvQhydSfxfsEEHyx7Z
AhJw7yBbqAmjUvbW3dkTOrMOJIUCz8H+9vTL0K5gTjCKAd7KZfCEB1JYQ/MqspMEGcM1fHJ7r6W4
a3xmzCg4SSlit/G8+rvrWmhVh2Y/vIT8dRPfqafls9jMUckC+QPDbcBjqtcOkYBEpd4E5jTQ5+vW
3qFms8iiJZmF3vZGTbTbF59eTFZ2ZIF104bx+jYAZ5CidhF2JdybEq2uxIrbT1GHhiaCft8CyU4l
xNFmzrngpPavHVb2HWSUyQDl+Ajp8CQoH+DcWCVy8G+NEneRu+pnwtsrd6GuBP/AWVfv4bhKmoRH
fDrkP1jCp+8ej5nFDrbzaVKKYrqYK3DJh26a83F7BTEavM/VMhAzq/tIduFEYoibgqzlY6Gxef6G
iXXrcieixXXVRsGQq0YUXt802D7ww/Ibew+feLSruyH0TKf+siU6YEy/O3tOk3qCJjJoDzCaZH54
5uJ279FA6mdmTxT2eCQxB3ZLlq1uLbrnTE0LL09wScNiWIefQE0R+iqURCl8bm6JKYZCWXKn9+2a
BK3gtJnlxViph7Gd1qDxqicNmTriFRlMPeieaqe7S/oCoiufOeG7A84Qsv6G4Y40tTjAAqGcopig
dTniVLecHvq9Kc8TEcyKXgCehm9K6EnbtX2ffPwlII9ZcDfjoVazVnH7Nmc97H2uVsnvTvz9Dv4B
xhRvtNdqWh5b7KtzbITIJdN0iT9iD1o6bJEGwNG561AiRUiKXAmFnyTWQU396Xz8+6fA8rNZ+JOQ
qPQnVp7q+eU8l4lGWWvOxjP/9ZSHCAFfKCDZqVPTbps9z0uMxnUphbExwLJcEnYJQBQYkNzzmoyk
7FBN4VhrlLV4BCZJy/ZmzdDHEnXqCdADcF5Yt1YVaE92L6ycMUN72PPaW9YoKNfvJcQBW/+u3MXc
cPCRSQN0hO6pHMqy5yfH3dzKHh20XnsDIisOPMtY8eWpO3GMuRpfhlxksSomNULEuB07CqM9z7G4
Xjlv1wNWvNg2KGZk8cpu/XZg+JrBerY/CcBl10GGyTsljx/7LQcFlDksmyk1utMU0LZjdKu0QuG9
yX8asVFo0gAjpX/QfQ6cW1MzTbqEecttp1/bXgNSDtElJME8AlnvWjwPoHCnlqr4HcKa2q1yhDbW
cXx/A+8QQ5E9VewxZeuCTmvCmuePTqk33rb44SBc5HXvVo6ftTFTkt3MKW8ZkWsOCDm1V62oKhJ/
7NBHxmkdEz7n5Sjkz3OiD7gqIRIcGlGw7MdnGG5w4klX4CaYuVYUp3Hh/fu/hPrz2iR2HewG1yHq
LTGaXuFkHTyESL05GThwKMUg0uPjc8iI4BLVU8jKjsYthKQbiAIauGWjkWGE4uM074WvwuIhXviq
Pg3ryG5PhxjLptlgEc0HC4aogIlC0LcjIY7GcNF4BTMJlVGjKCW6lG7WutJLCY3j2jGFDd3oyXSe
4fthts4IzVWOCke1d/DIMly5hE2bkL369lBs0I/7bYf97ghaSQLdIUfqtsukY1PAy7k5X6mOQocs
+H/6FfJ3851A3vqAqbajfS3rDmik93jb6CD7vBTdOD3y67r5vJ8V0UBfkWcgP5fmuBSq82gnrdX2
fLkgwi9PxUbREt3Nnadeybke9H+6TGTwh+xUI/NpaD9zIo0OL+X503CLSzAzjxEWc/R5nzbk1oF8
sDcXfk6JpMB5YiEkMEH3IICoG+q+h32VJeKtzn6qd+jNHzL8QvMUytaEuMjIDbBlNllfSkKFJL3v
EbKZkbfqOTRXpApA9UuLtZDNZWcbZuU5CBo7ZeIaUlN8TTDpy1H68F5Tyyb5TrtL6lvIcaB0OQas
xeDANNpbGDqbYbOe5VfvNqwzpXvky3yFe/6ha5pqO4rT/8r8IlZMz0pIfaEcp3CHH1jklc/rq7Xi
xxoPkr6wlLaa3Vd59ikMX37XoAAu95MugRl5i86pXZo1y/TUfbF+MPouzvU7Qf7k6Ue8NwQgisW1
yTBCPfHD83ktW70KJDlMXKOAf9K6T0NPh9MG9hp1i3vjwg24WHDlezOOqMowMfU4M3pb1gTGdaDI
Q0vHSs0fX2LCQsXG+mAMpu20PD7eL/pk6wnDtf0j4/MAmd1ZapBJljT/hBlQLIC2OHkTmiY6Bw7w
d+pMXkggtABSiCPcXfECJytIf7P1+6pQKXDNct3Ojsd8aOXmON3U5yKJcelSs28cn0KuxPyY/9NH
fG3NYX3IDkNCOy9rkeecprYvMr5GFul76YpjIaxXdOxFNpSUkzz9ih9Xsw2V3HxXBPKeqQIcNfAn
vdsmEropL7g7S/jckFCfFXPLCMj2bTASqVpAYe7e775bkIsx9gvLA/V7jrAxDTer1DvLaB/aukMt
50O+rRgtAXdAv/SC6PFBSeYzDtizqT3c66BW/TWLbsax+IIe1/wl9y99qLoAxoQx2Rj4VQKQMDjD
8zfB7gHJW6MuAUoq+SKrdXx0iiFCgW03lFnPmmjjpAD1CBvqhE8PlTS/AJW8TzKwnx6YaoEh5kam
tRdEEuwCx9/DoxHeSWePUTqG6QEuexmA0cEQohPiOaCI1lKiMf2D3XuuS1aq/1HwQTvrcoCpcUxg
DJY96q43Sbv1bs3DQGe+eTPn9wNgEkNtIMvZ7Sb2UFR0Y3M8VvKdZgplqdxup7Ebx5fvmKTFVFyL
pxJGzk7KjIJ1hmZXKojl6t96HA6SoP9kEDGwEz7KFaekS9oVajUobyyOP7MFc5WwlxsyuKKAWjmd
Dkkhu5VlwlGh1UxAHBSTcAVLfliiOBykmM72K+sXwKqZlDL3d4dMC5Hw7EA1ealqVX3CmvcMKLKJ
V0Zj4sorCcL+CpBtSHubGnOC+KsFheUwVWh4COJZuQH+jQZ38CetctKQXLRDNtdvLWspphy568PD
0IsVSN53XBPKNlWAbfw/OqiGoaPAQrtW1Q1ZNnFaoozkUEXBblFqrvFQErXEAdgO15K4n59+MNFZ
MU4iEPyF2hhH2Cd94BL8ia0r1EJKphfZ2f4oFZoos/NY7tccCKEuXF3OMNnl+dTVGg7deal18rGq
3Jbcc3qQcf62y5xFYIZipoK+3BGOKhSFypvVWwVFCbgtuuRx8Wd5MnpmuX/l4s1ORGWd3FqFIMMi
ixSEJ0OMihcqi2bwzhy34ei1wQFNa0Ub65Gf2FrqxMPTgFFiiVq2OeMwuA3IoDUSymj5HpoMueTW
FJD7BqCLjeCwBiKFO5n+iFPFQm4ii0hgm6TXS4BTzCYFHZZv3GotFJRVZzLhv0oIvJKzeVs9o3nz
S8LbaUAX+GHB4WzfDuhWPKIJ6j9KMjc6tLJX8JPZJtT7ZMIqstkFl5WR3hX1O7ovNNGOm4I0M23s
NvbiBrXCD9LkAjtrZulCiyCTsewaAg4r6LqKmUV9laRQUkLdrZAUiCNvk4PhlxcsoRoTl2UooYUp
o/MYxBa6LHJvWlQeR+LkFtgfEbPLaO58fsY2ApgWyrEkOTC8skqdA29M1kpYUND3l9NofYqZlcpM
g2hekwvLdCl6OdOXKsEvCAPtLtLeIjFn9yT9bInM2sgOcvI8PFt4xm8qCT/GUJaBoGnGwci5kFfa
LEZVUPNXqeOqpSHs7bPUJFRtg59aPfloySN676G9hNoFPu0BohLA63+ATXR3ybgs8UNKiDtp2sxa
LOlC3vdrkKmSHcO7nH/pStGF0RZ/g7jZzKvRBsJAe/ZwtGaJv7WKQLRTi2izpvw8HTHfMjSbhgNe
xf9LW+kLl1qfWmf8P/8Qi/h2+52A9LvjgUJXrua6YdGw/utB6h+8u/a7a7B571NbJB7+vzH9Wcpk
U6DycbfTt2CvcFoQMi4451biZE0F5EzpCgomo6VD4j2n0lUMzyCDxaLUbw532M8URQKweyM9+vOV
oFEW5ortiPRPqZEKjlmJIRyXwxCdq94nAaezH1wbFxco7eRiysJsVBfaIufprVygoXriUCJ0pcUm
2mJNfu+MVKOPwV3nIBby5tdcg39jpP0PAK+t2k4rk1bfO/YO7fL2jg5NMBw/ZoDY+37TN2rzphPR
wIXBq7OI6oBnUEzycV0YUkGkto0LYSVJaJlZwigdoPR3bStBTOf7exT2X0Ok5iVMAgxCUziuybQe
UCqvo8M9m0W+H0oO7z9XF/PfqnXgwWYkFbmUP3tQoWFKf8tQxnc3t3f6HLn778loj6I2IJoA4f7V
o44wg1I4BSbpSSrNep7kjj1avqHieM68HcXwqM+Rjb6bPP3BmXkq7ffZAMEQTWzridmXtQm3TEoL
EZaOkbCH7OUe5iuMlHW0FXqFxYY+Nj/7q1hfs+sCY8Woyc+Gyq5KXGY0l501Omw6I4X18PKMP7Pt
lTiHWIx16PFUBQ4c/lqeQez6JrXlH7GcTAyWD0bMNch/7H3EODd3A1coZhs1IGSpVcsl+wa6YMId
QA1nEpo9CISEurFea9ehhkdonlA8nfwTBXXi5pCKLaRe0uKtqLdoGU6gJ+47iNSEsUPg568fU/B0
H0rgv1mYZs5JwA0UmB5o1C92G3n4Rf20g0RwB88Fa7mcVneGj0YUKjs69ZQe34axvSCi9U+j+OGC
t1fPK/KzTfZ7XP6D5s1Jsr9S8+EQrZ4hKULkZMJ9Bopz1cGBaDxhJSvgSpnaBA4p05IhSa7yasNK
vFee1+FHqXGdWwcpWwsqrZQHhmZpvNRuhdDOoVak3uLZB5IEXK77dzL43acp7dJzam9gAfPK8C4n
NeMDgwNCX0XPua2ljd8TJWAPxLM0Ue3Nz5j8nb5PAqMnsgJKu39D/Kw65kqv8svgd+vWLI5D+K7T
oBlXFZtu8TyGhXCCj2NnNcMSJvmlCBV5H9tt57AKEzDLq6Ne8mvTjadSGaSncVk3VVn12PJwsNhb
AS7gnf9JHc5N7smsim1pCAOG7gOH1yCvCo3U4N5yBx7HsCoMGSGwt5xzsBwe4FmsGmZrNaOvm6A2
T+BRtBBKzXQKmhsJpiULnilz67XedoXCgrv+24cKqJhFWv+hLwtLJLj2ZkXKwLnbNEifpRALtpck
N41oLuEFUOvtS3WGmD7x1c3/W7bwr64mWF2VhxlZqqIoBTjr/id/fLeoT39DtXyrQCFQkfsbciTw
+g5MU7HDeXSuDbDrzILaah/fW3eNFJ98sXsFDPG9V1E4hPEGmd6VLKv4CzZgmAmsKJfLTI6f8jZ3
28VmOWR6c1AZkr1bV47yJHimrn84UFB7OhtfgptkZuVmm30Gd309RMI4u4XmbLl7TdvB04OwD2h2
Uicu46l8nKhpZRxmUcsCuUBpo8X5m6ZWMuoQNfV4sKeuMEpxv8eUcg8+Nlblu71npKtmBHn88kJF
RZ7WTrWUyRD52WfOW4vs8qE/24RfNHeKjIEzQiFuB6WoqjILlys8ilfwisKg/DDwyC+BbzdikfHZ
GuMUr2CNerg2L3YXWByJoIXhjsTiDB8jIbUsRNSQbTdb5QX/64hZzPW2AnkYkxrqPXCcHGGqrR4u
HaJ9es6N5HqOqx4ur6UjbGWQj+QZhi28mJiEL3XtMbBv0PL4skbaswH/BLp6lwh6F4h1g/gk2Dt/
IfFbS1HkWQr74C4JvlC4UMTuVobjEHg63mwxTx6FVVyGuJ2rcdafoKT8lg3ueddMxg0m3dph35HD
pHfCnCovEFyTbmOhRdJGWE0uaGwO2sAOmTxoJbyQlqUjknrFfC3aqi7I7UqC2TYa9WL6eXPnSYla
KD5l10n9CLoaFIPKC5g9F3gC3Imd6Jf2/x2DDMTtZH5KfdQszFrVXEi7zZqHC/IgQjnkPBy30j9Q
IR2LSmwEErYqrrdUgHAwqo96MOGAymUxPWyWRjU2Uu4/E9GMG51TDOMYXLom88rrEL7cnOlogYKB
Zi9z190JbxSnNMDlV0lZVZyPznizT8ICh1hewJLf3IDDvkECkK1i3Omy5tVjmixcl5ghjyf+a3jC
C3VFp3JtwibDGl+o79EeXIoAS08/FufAB6gIN2dpJTeVcA0HYENgBv12wxct5wf5m0kyLNm18wtM
ksjZkXhsbLYpmpP1nNSueXMt8Z8j05Sx4+hgXIkEQM1EAldfcKQJOf/CuIFqsur2dh9/8tpwJRZM
MQOlKgt4Y2fNDaQ0wOU/aHg/n7TIAANDzho1+RmU07AOYk9pVSk2YgmCkwNLOOagzd0MXu3IRRbD
xyUP4LTWwAwBweW0kdCW5W1HbIzHrGPJNYpTRxp5TP8Uwz9OzM0JsQ3Eiu9rr5VZRZzkWwQw9y8Y
8iCLv5dUcqGk+sP+kVXDcRWvewzY56yq5/xgFGo4lLCHXcXSb3Z9TDJT9chxbkjrltVMAOZjOzzX
oVVlVouZmL6jP1OI03Dlv/v/8jSrJ67rj6rtM6ojWco6sCxiFC+7UBl/28gCImMRO0fBYW9OIama
Y7mEnByknbUBbFarb1HSleQ/yydkWq0culg+RUip2zUh+Zf57UzdqxLJ5J7EzT7MJqyoSSn8JqIe
psY8easlF0QEgUCMj7pPUBqHIk5yeXu5GNBKV+ytJ00GYKMSNvHkjQlzNGCvIHnbDTcAZU8Tg6Fs
1bsNY6bZiArJf6bmsOcgWtS+G/vBbK6GeLCWU4m2U53ypUvQOq+Ikv41wtr97Tr37eBOzlJU8a46
Zav/3ZfhKo9kkdjJhXcNGfnmyQGifYagye6hE5SLcG2rtbKMCCTDALt7mB70sLedRzBwBY4/FHkI
aJG9Eg357QsJefr9N4MfdsB/wmIi0RZ7wBK+lfTPIr+t55ios081c1cA4zKByRC5inaNpE6WzhvC
h6M4KnRG/4DP9ljePmjZWZNhocPF6lAWqJjALGyy8yBaZaLooN+CJA0FtCsTsrG/7i94XfoUR9fh
YMKoomFDxPCqXxzg9kCj3gcJJonx7RbmKMVZnVInztrJhhQECzA7OvabaR0nitaNgSnVsvwdN+PR
i/hmN89vSmRg5KQ8orXB5+CxVWbVCB70cVWqsJ+lQpOBTVgw+nGSoV9HrPnCPvHeG4AZjqPoqdrF
OtqHH1ybnf2O8zOg2S8b2Oa23kTbLKHVtsvYv3PsfufaZcCXKH3y9fbCEeS8+KAxHrBJJKZcy0bB
0mBlkIldmwDdJJs72f5g1d1UVEjsDWRIKBITMjJ2GfFni6jlDFw/d7fkEHoZ8B/FPhBBVjGkuo2N
tve4Xtydxplcb6L0lH3EBWu2r7tKxXvGzJi4V88TKl8Q+pKMQuqKuCp4YxXX80XDZkRwl1+7xA7u
6RzshJE7nAGnZjuS11kG6kBQJGMM2BASBsOFlpqV9TuAGnumCR5I4o1ucsXW7RnfQAMp8N6dwayf
auNao5YpmKQFfoFkhfgukJQPHP+ONca3YSe7Ie4jQN3VY49gLTlU0uhjuDSrAE24MiBN9bnTjKuE
Wuo3iszv+22vP1foSL9xXgaV609ogGoY8lFpXCNikEvVBBQH67S3I42kfo8Q6IdHgj+O5G5CyNOX
8dPvhKGyW8QteZ15DLM2B7b0LpqVitYHB/WQwaEeEaoe0JQQzGkqW6xb+irx8gc2s+GwqQH4EJi8
ly6S4xYFz/cVV2oWYmTd/aU+MFBPn5eSSGtZ5RQw+uxzEGLQz3C2TIi43j9smVw6vJAJkDKLA8l2
yXFIs3dzcaDwenpqNsOUca4BP5seoGNjGBveIgiUXPAe55BXh5D8olNr0lTF5q/YqUwPBGaU5dRX
mMUkXPdxxehpLyuukqcs5MnkRGlCHKPOdb1YZnN7U5Riziyft4vSNuKJQPhvFXObHM+Cq9kYiaHC
6ArZyQx2ZrtFCvtzGeUhylFtV3ntOp3lzKyvrJGZOV3t8GUdTNhso3yxj8Qn49O523ZbbqGPUUJs
Nak93SNp/PHIYNcaDhhbLWtWX3n2daYRA5zRHr4jwfy6C9dvYoFB7iwl6HDMWHywx1XYH+ehxMvi
j023yK7/IqhvI+zqpgfCNsJ17vcvqSNQX8CuECWbq9/SyQC0iIB4PGVlUf0FcwzXWQWOUxfwBaCQ
6LK8WpWN2AOvh8Ir8fUPEMgYmcnDlkmJ5LLx+EPr/+O/OctTcH6j4fMDL6uD1QwrBd2I4ViEQEYj
szINlnfscFJaHu3Uvz6v1qSy9mVXSs6cfaqWTIw1Q5u/E2SO7RBINnHPcuSykTzTqrMrN9oBcvPA
lUy1DkZcKS5cJ+Xq4OgvtUS8xQap4N/XSv8bB7dD00SbhVY8r+JST6p9OMjCvXKXP5Ren71W4a0c
9r3IPAUf9ym+erjUGWHtQOVRtm3ncC6RV+qd7V6hdcK6q2Rp7VcxTbEM0zBx2+hoaFNORAXhYCfv
meiwC9t5ZLUym9S9fkpWV0CS6C5w6pFiWf5ThXSaU71eb6OBCViMvc45UH5UCyHKyzq0ywkTDYfI
Q3ZUi+orCiW0HwyTQEwUEAV0p5yKsf/anNisGWK0K0QLQhoZhjy4ZyuhMA2rTDvsWYyQ0wucbggT
HF73uBJ1Dfh7dMZ6SYaa6FxxTk7R7IhFG5xAU1e2qJPXZXuN/uwduHrz5gJti0/hRsFlET8URA8F
mv8QW0g/qSk7eHoOR9Cte6PudWv4jdw3JvBGtk8MRfSJOv44btsoXIyt0Qf3Cpc5NrUgzfRc8zGD
hR3rJIrmy1fseMhrs7pX6f6cbxcZ8pra66P9wjL72mQjt/1i53wtXdjA0xihZ/4n05zKGwDpzmmP
cFErI3ZTAK6XV/JaWQxMTypiI3Ioj6HzWqc3V8dja4d+lbZzdz1EYJ7kBHOwvrcgix4PpJiiqA5d
UdOhSMjSfVl1CAM+xVKIoRUu511p8EiFX8F5NVWyDjvT73skkIK++k6/o3fo/okMQLtbP+S2tkLz
IxIOjsW1WfgXPX/G9C7AY78GLShmDSmNzfYjeMn23JoVFvFl4qpvlfUnI+Zi/YG3EEE9r5EJPYBz
lG8mROzmLNTNybdHQjeyNbUVClYhKoK2x/eq+PdSr849Dt14MeZbMApVzf/RDYqGNI2Hv8/h0V3L
kvnClSGoCPID56weqd414afEBa7/pFEMfnTWznDeLjOZxGHqXvMYYz+wnh1SWovEQkhs+7De+HNN
onlvPd3blyayLqmM9q8Qhq7kK4TQrOSrn0WfTaA1cdmvEmaIvejoXdGiJXVD6V7STBmjZzxNGcdM
tXhB3lTvNqIiCnseRKQ+RTl0Y1BRmZfHHyZSowDGgfEuLtryaAHNnLV0LbPu4eDZnBtRpEZ8fZ4v
zxrrIfm+AGuw21dwz1YAlNAVf9bmce6vuT7B2dMzYs4OfV2NE81JVFQuxEck/GD50M1K/P4bBqh9
cUywCWgwIXydsl52rzqW3m4PZIlFyG5N2VFdRipM3lNI4ebViNrf1qCgzfx35RQUQMbzEsz2m26/
Ent9IJ6eaWtIYt6A2YF/3funfinUdCYRzZGMTpFsPkmWQGXacym8ilgzxnEylknW1OaBam1U3EKn
0kUda1o5qhBKpJPLqmWrzMY7WpRn4RIe5uhSKjGYY/6zYz3vrTpCUptbn5R8TZGDLcT3w9ItzInE
0a7UpeJuS5hEbSe3aQEZsr37hWCTRWQXwjpF0/xmzqVL/TvBPNzgYCqJNwf95pWfR/2kYYjgLmq5
L8yZ1I42bNZBrd4bMvlteLxP7z9mKwOgpTacriHQRE3DiTkrKicOvoI+msABMUlHzOO0Ny6Oy5Gt
1tOQ/gGNA4EUA5k1Ess7FXVvf9q/e752+cvrcB17xTi8+BdteBL9CMDSi58s74rhmNxe97AiTaom
8jBfc8r87ICx1dnynJb1BNihEO2saUxqw8Bx2c7Q0/Xc/i7s8r6xF1R+7114MJgGSS8/TzFrZZ6A
T62xbpBgGVxvaRGVngZhcZ329tq3x1MKdCWLQOX3eVBZxtLQMWS51k6e5yxT7yXXDxtgzgsVy7Wn
eb6jqpqsx1bh9m5MYpkW6atfMcnpgzEymOfbOc20Z/i5kQUXItg3QxiOszQBdgyXRJxXu5R4q5Yr
muBcwogTIetcCOdvbQOaY7tdnjX4Dv1B3CJRHrOsRXtOJNkkYqbayje41s/xzHDnC14b1h16CvJR
77l/RRAC4HftpJj4LopYaMwxSWWtoFiKrry0X4d4AZ57aLTx3/29tgZCVizgKs7o0kYsyM4Ch53k
Xx+E1eTXJP5Ne+sRBDrKyKjszUJtFSKMG6+dkYY3oKi2pbjzTmoL4AKvXQrdXNascZ2+u/LYgA1f
d1sy8zfvKbIYxVgqek0eKFXq8/thFw9PQALBE/Tab4DR9REF0GYarLOOFFkmfJMuZaLWtqcawCob
FsDQqAm45F0NoMtJK5yrgClsZw48bL9EXL65F2l+zxvujzQeLRnTZHhAm0gzsQzKPYSPTslDuCMd
Vevz5cXXu+eRFbFolKOsVBmhgX9+iy0/o0J9DnNeL2Oo4OleBfPXYqQ8hkNiTLig976mPkqhoTbU
M05zYrwUxN70yXcOB/Bb9lgdCrHrdnG+FsckLq/5cMbaqWej1kz9QJ3neW748IpysnLn0ZEqIAGn
cEybYZelxv8h9GPcMRGZRqKX8ClozEVGx9ffIMS2MJXHlYz/VRzoZWbeFc8NgwH1AYyrya+04zjV
9Sto9IhS3WxsT4GW3dogtDKna/o4loR3VsSE4+5JPhDjvpDwlQyZg3SlDLMoi2ODLrOfHW46pYlD
jvsQbuo78b9ltHnpdZqmKQPKrPYuXoCFz2h/okjv2Hh8WtgUXIb3XdW4ofi3zeBNsdcrFmWFzaKs
bGda40yZEphWNZ3lpfIUdVtS55c+XJ1qecB5U2/i6yPqqBdhzhICbbE8WrJu8tu/tw14hkW+9PjN
aK0O+idZUC56beF/uFk66gzdVFWrEdS6WqXxl8+Xd9Re2fCp3TZ4Jy8dpLt7K+4QPpeX1lzqbzmr
wjXltF5cHEdSCrEXaUMUjmuyNoFeTXVbQgJFlnwRUQWLbkolrF24lEe11QLcAG7PeVliXHGq+UfF
M+hh8/LJehfR/gRfGf+TsoCp3BSb582wKESiK9dYvl1ypM0NuZptW1oWxUz+bFe/XL/I7Dg1WjKF
H4vvLNvlrVI+TOYo8L2IM3OE+lrkKJPuXg4gLVfaceKHOMZLbbt+UCDpPUDJZDJoJBFDRLW6cpB8
TVhSIyI3FPc66biYvdVtgTmjEQlL3HBLq1o0SZSaB9ULEOnjENwoEpBWQAG3dhno5X1c/Z7haNzr
hpeFL4+qISb/+b1u2d/uy/ilN92g6u3+BjnQToOnmsZ60mMi5USPqfwwMX1MnPtVUYerL4az1U9y
pTB/8dIn61/mZvDa3P8cS2sUotxMo3GewV0HWiWslBnsWy+kANhz8KgU+80Ftoyl0044V3Wfa87k
vsGj1hLRdhYqe5ussHF8yfP6prZCE1saG78SgwI+lVAJbKJxPK5xXw22GV9W0+CbTV6LOJHN0Eiv
0WRbB7ULXzSoTx1p6A6Ym/MtnXPy4bFqNYgDb+zQOz+SU9FNUnDYKua6n2upYSFQJ9z1MtDf6n/D
VSXOWI3gpSlQBWjdN80WurMGRBeZnZpBfPszOkus42PhlkWxGZ3NgENRqXQDqqQ8Bl7bfTaayWrB
q6Ozba2a9p846OotHYpTDKgiD8IH5psNT3WTl7zWW+nwloV6R03zvkI8lpGaBliBunUJjYqWPpcP
7zldUUyZUdWm88E/9BFhE/YcjxOw5r9E/AxxK29ZFyq+49NlICWKIMTQh9MacCVBFD3sfQhhV5Ka
hjckmFDlOf8jJ9QhM4DeDC6gVvew5+zoAvVIqFLQSQ4RpUdukAXS9n9h04FDLpsVAmOPXVeWfboz
AQXqy8eWT1M6xL7BhF7qfoNGUFGeivT+NOsG2wfkWe3BAJCyREdJZA270sF8wcmhwCBAow36QCJs
XMyrfWrbluict27hdfIIb/lxZmpDxzyWmhmUZ3JSzQd+v7PvhZM21NWEckJKAkOnq7anuvUMz8pd
Qe1hTs+23PkPJPDfCSdzUWmSPGYz01a+sMSCcth62mk3JilRgOE0X6Y2Mz4YXEyS8nbZrWq+VmbC
k6nTUmlS9/AzFrJvAD0b0L+DA20MsR5hULAuANaE9QW+HZksIBajuhlGdtrEyv48LDJrpoUS1W7w
HC11ZNWlPqmHur6bNrhJRaEgNBUhNThevqQ/v334prR2eObfbxX+XwcJYWXaZl9/dWz2RX6/d+eD
oxvZ1xNNZ65DaLzaa5uEBL6KZa+t/gZHBMomZGFc5c9r9aB66PKTT18P3MPXCNYsGRwI9NA9J98V
9bjzEJvhdFfrBVaPRXqupM5dm5XPTwCw5i1IW9b1EaGGE1qWNmU2uVM13wO69iHwF7rhHtmLIPbm
tXMhZk6k/1QS4EXhVUW2jrSayL/ElOeAdzZe/kbiWtZqgd5zI5Jr3FhWZdNoGvQGf5nbg3J3U/Pp
rD7Wx8bJ2R50ax2vp/50qAgt360VeJ2mXcRqQeQweBEhCfNJok/+FO6G+uVQ8uCtcGFtoqUTSS6p
gyZqyUn5SefL7zYGpz+S1xt7AzNZwL4hsq+x01Kqr9HV4NQ6Jd1OHkLYk945Sa+m78ds9CdbYO1v
XyUHhsBx84BnNECTr6y/13CohL77DT12WwhFt6TuEcCfklBDgOwz3OlcdZ9ZXXsPLamHrhSdVzvS
oe4CzU66i1/uAs9uXbf486H0zeHcd+uH1rUZ6qR0I3cFiB1Wjeofq7Ey80Jaq7uZ5hylHb3XU2WE
0B2Ijpkj6I+MJKyp/vnm0mqZVgcEd/hHLxZvwDfcv4SK095qJedSO1AudNtRMxdmtn5AGlUS4veu
rXZQ+3dEg275rK5vIa8KMF0iWUUp/nyvlCvj7jzYLFpaTr15Ib5gsKseZp8pjUlEKCfauZ4PoGmZ
Cho31CPQNJNxcWxaOR5grM6C7fgMHACNWL59/yltyKZvDtFr8HXYz4LwqpFdGPtUI9wq1mzcArc6
Rr0TwDJd01iRbEdxVgQxpPAx/eHtpjfd1lDxBC8meBOmaBcmHkg/D67iRBFjAW4JdkX89YNIcQkD
1zg4wKutpW4LLx2xCxG+kR7nm9S0Sc1VKqzhiquY3F0BuhDjXncpwb9+TIMjzPJoKFfU0q1Hf25m
kjOQL6eEYEwGIzgdpAV9KWNRam4/OOXth1TYIvtxOvQUQLrd2SDaVKMPnMbYI+e2qaFgImE/y75/
zJoUo0T7dfZHFsHF3tkRgjqOE1NTPXGccdXx7FIg9tWypX5fDgtWUQOWETD8awghjxOr/OabIQ7F
l00ArcFXt58BYDbVvflg9LgAGr6coDan/oQpZb/2oVnQ5wzucB+ValwWsiQ6AxIUexIoS/9l6baY
ApSsrnfDPxIJ5TMW2FsyaskVdTvh8DCTZu5zVeOA2Cf62dPj7qlx/RjuiFMs5/v4n/+LlwzFMJcG
33FSlmM8SQYuXsMwUng8z0hhITLhWyU92BS66cQjB8ezx/04BhKAt/aY9cRxK7lncnwj+4vEXlDI
jBLVh0t4usrgpa2Q6eoJOrbY6befoqyC7xAR+iZFvapkfJrGmoLgUA5ugOOFEQUR+eqAxsL9FsoX
28LCURpzkbUDVOSGe3F6y/k9lthqcTEwNPrHWVKmkVfQvroioVM6+eApcpxcFjhWCgnHbJoPIETy
IhYzDuJ3uC2Z9s8Ro3ZcRSZWJNmIifYgA+p92FYFgBv/3aTp5FK7EYanWmrLYlpDWM1wq5pgNp0U
rwUAi8M4GC0X1/4nx5IS/yRe7LEH/c8nfhGF0VZnPlKacyvrVmfIz7Yst+vOzH9T52CDjs3koQiG
uKLFbIRnxIMzQkqsZYpMFzVXW5h8aYIMCIkYG5AX2Q2X2FbDBMoaDIf6D6kwEJ/Ub2+GYFGFluSt
+KU6UUmh1iVWTWVzh6b8/HGc7W+jhW/iWbq1/VZ/b07K3XU/9wVXR8ZhFzseXAQUBeD3OqENRSjk
EMx59m33I3o87Tnd95aFN3tQa0YsfFRJ5x+9/fJyhr7xwSRpkZT8z17wp7Oqt98YRDsIF6oeLKNp
WBTpr/+p8LQ1rt/UzJqBXBzULwLgyWjUbxPNYhC/6JF8T6L8mu6BqlhcGoNEK/v4VLs+iBGiH/Mr
XINVwwOImdJ968TwRKsy5B3ZJ8q6CFK3uFTl7Xb/RY9JWm3grWc0P8BpPu13Av5Y0pG7y9bMaBdB
kn40D7Ofdvgo6/np3EnCC7ZZL0N4wv/YjxptK4h/Uk4xgecsNqCAkk/riR8MHn3kXChayHuuGcMI
E6K2/puZBsGFxpvMjkIFWT4TKSWqzHcpmWK3+L0o3Ay51YzUkUxs7pBvbDXQI84Af/ERCW7iIVcE
FhA6nKAA5jSW9OpMbN3zfhCBboSzGNezC0yP0N2vBLymyycbAWy6DSHku//11JjHLfsyO7al0kJN
mI2KvYiTve6s2AoqSAd4dTuKSI+xTf+vfCuPqNmkemHSG+ZitzePrb7DC9DBpeGGBICepOR627ke
Z/IiXCmlVJplJTnJ6tPPz45LE5I68RIWC+mqNUYqjExAegwRrycaCKd/HarQI2MPE7BLP5k7S8SY
xXB2qquAe2hXYt/i/SkSTa6jBMxgiNQoLC6TcNJd5aoZ5dK1sH4NtJFOk3RTN1dgFTw9JCkdxdpD
49Gn1tSmshazARO+Xm+WzYXy3FeW539DdNFDOzgTDLqwOAeRRXHxoahTSt2hY2IdjKlSEX0YyXnP
h9rGsR8vy3yXQQX+sFFqRq/HOzGcKTUrIP3y7RQ9RhIYiGc9el46goVABBiD5y7r6lTk6AfatMV9
0u6qm8AWsYf+XlwclTAFczVjcTInq5bln3xWqCToIHd+oj+Q7kf1LHx2FOLxYWF8sM7Gb1MayePU
9dQGX8295dp5adVQZ69GMkjZeTNCwcMDReII7ymila861wIQtmjTDDFY7xsCXUhtk3OWhzxh/Seu
AaYiCi76jZT/tqdzEI6Mfk/WDeucRvUjDdQB9JZkIr/2e8UA3EJXxtEmSY3ObgnpP02+d08tKaVm
v0pINL/0ur+J2PRGhKIb3Wpn1EgMsP+KsRAVkho2jX8HwuLDHEToB4+khEgUGNNbXqtyyK9nEEDF
8GBh7vqhhaQvZeWdvfnWKFWG1hqPjreRB+ytX/nzSBt9XfHPMdyk+69b1nTVXsC0hBsikKZFgxrR
1UzKzCceU6MzOQ7c2cc0C8ksppy4Q7lPQ+V1TFwzot239TeMK7pK/xmBGHLiWMS0lGBIrMZPAv4s
GQxvvXyklxn6CjwVMHuF8Fx1ZNhAdLKgPN4F7w5v+26lacUYaZrYDaGvOY5SoOxDT9HfcCzYH6Wo
lW0V+1ltmlqROGG2XXtN6TktBNgYM+/WtRWcYtBeoezuL18Hxs1OML3D26tYbyTFKR4G/biTM61a
ag28YuUj2nyEI1MqhoVWf3Px3ozUCkMoWKB9MtMCqtkdIzxPySqrPcNjBoTKaTpstgsaySCWkXVL
m4dAK88Ct3rPF1SuYaqKw6Y11DXu4BlXoyROu3ECH/oZpw37uZbx+lxa+TJTAkM+RRteSPNtCyzh
XQMwM6qjvoneWu05cIKPxfN0nxRIrhU8lARE1IzWozqCnwPOgcwIaqtUsEnARDeDr2TMpEHyG8gh
gwl/Pr3S6kYcvFDgdQ==
`pragma protect end_protected

// 
