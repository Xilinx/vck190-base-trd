//
// Copyright 2019 Xilinx Inc.
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//    http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
//Setting the arch of DPUCVD, For more details, Please read the PG


`define wrp_CPB_N               32
`define wrp_BATCH_N             1
`define wrp_BATCH_SHRWGT_N      4
`define wrp_ALU_MODE            2
`define wrp_UBANK_IMG_N         16
`define wrp_UBANK_WGT_N         16
`define wrp_UBANK_BIAS          1
`define wrp_LOAD_PARALLEL_IMG   2
`define wrp_SAVE_PARALLEL_IMG   1
