/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Fgcvq9yodAEyu7zsWWZ7LwHLqer2uRdIROgj+b6me/wmyj6mu+r4+a1EPBMoGlf2Rxb0wqrGm/yl
7FT0a+0gf6RIUa901Ug60cEq5l3MsNjnNX0EuQ9QHnbWnPHO5sk3W38XYr3s1DoIymcMyzWSb3j7
DAgt+R0iGXGbLJHe2UuAgwrybNhjpWacbybFOYZoLu5Z50wmOHt3p6J+gVbTwfuHK/f+KnS4VtSD
EJxx9+hQNEvkukNe5IcvkATvsJ495o97/SdF6+o/UvTHUZ0m3la3MPtrbbqjxbRc5d/SBaUYwJ/0
DSKgI3IBXs0nO4MGwCQX4Cy0xa1KtNy17Uqy4A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="YyF30NSJW4xBU1bz6CmJ7uDDg1utz4oEiyNQAWYk7H4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6032)
`pragma protect data_block
3JkMrY1IEAXvStruy6C+3vMii8x7xMb2kbKSKqbX9sBt7EEKNMzlKTbDh0HLsACCZDcjRcdDf/cJ
AZo44x3KgnG1ijjxjciLMUksUaThvOS70SDPtU1LsC0/jbULyAu6AoeA2Zoi5vbAEeABc+vhgtRa
6A9egV8ZQsJs+GoAFieYjbaG+yRSouBW8V097FAkWZ+JsNjy9cVKEi9IN9nDvYLsQ8/tR8TaUMLU
PSMbC3KQOY4GE7J/xEpgx0IQfDYKhFfa8Ea7iK9TSnxk+te7CO9EBwQ5x52ByOgyzHoJcXIBmRw9
kWOirgqG/LOD9vtZAxMvmOInl85alLvVlY+ByapoO3IlATuU+MOFyL6Tmxb+WvaA+Cz1upmMq4Lk
IiCn8B89Rc2aq/csZevzOgR+KLexDZQwUWfnw1tGVX4kueXHVl7BpG9YVizEzrwOtpp865d+SJ3S
PnK0IOX3EXf//KbzuoZ4UY0COMZL1XJqYzQImWRVq8YDCXTmQBwLPTCMWEfx7RJVSEy6WGmxRulN
BDtQOM0T5gSCb41wn+pa1TA8SFn7hc0MvcITk2FjQaOhASionboCogaX1nKjmwWN7QXhMECVgaF2
KL/G588sb5VFlYlnUpJRkP49c02SX8UgeK1S4EKmBQABkAamNhttLfKqEKJsP/HNHssf9awkEORH
mkaIh/9XUGoWxfs2Pse6LHX0vSXmlpjsglarVtHLruULYt/AQmqlkTw01dtWXrIAUlqJSc3p2/Ur
7RnFCQFOdRTH1yfay/3RXtmd7hnKNB3aJ8dK7cEtH767QGzJpEngg1vg/1Y1j6EGjLDW9k3a6FOU
wF35XdaBjEJspyTw/t4CQDLw0ogTW6e/Q9CVc9NV4wfuF0zogg7v/5aSGkac7AmVY6UGcppicxfX
instDAOEX8zyBfY4ENmGoccC4h5ef6CJBc+eQkw+fN1EPREt/YL6ILE8IonWpbkAsKdxXUuOhamG
L4WSNCHPFgiE1euxmEBNxwyBcJGeGa4dHxKKOPObj9FDW6Ux5STdHW7w0TcRgwZju/adTrurpGhg
iZcXfPC2ptIbvSVQRXvyY/FQYZc720TDs3IeOVOWQx6AOLA91EWGHR/jDOqrOts33tpQave9589P
KZ1tPxwiGV/KGMfufXAt80cXpH0lIiv1gtQn3TJd6pZ4tHTq81jDvONTRU9rW1wBcXkke8wpoNa9
5kmx5yTP7CLQVEqobEu95yrW2gU8EnA5DXrMuGAg3TpvkyTRVm85jnXaLptU/AGK3Q8lxYOI7WEZ
t3Zt9/jlvW8Q7uQoil3qtzpY7Dbf2GNCUgDzMBHkLPXTIseFASq3IiLoIj4oLAy8AVdPpydPq0GS
S0ukIJc3LkpkmIBuecfhSkGi0ZLkqyTf0IwWR7/8GdDLEO8iQe0E2nuFfCMfuQsj5TRkqjnDh5Xp
QXjtCdqSxs0WKIodEdugfA+zhRtfPMo/AB1ZzvTPvi3vybM02fuA241V/2DXZq+Gjex+hoKfuka1
Nwuj1AD/zHPj05mmiOAHxNU4L7YZTYf6kAIn8agEKY019V4F82dUflBuczTd2vGo9exQOHD1dSuF
YZUhJ+gis54+ySy0b4obAlNZ/KwL00yNiL+Y5G2WAef6KJ7NAtAqD01GTbfx4TVOp+qAYZExHO2s
0ZdcFQLsZ6kIhA5jfeE8StmaCr7vW5yvFrtY8zEE21K5UwPneopX1tqD58BJZlD1R2kK7r0TQRSO
qEYlKICqUix+8O8pCgmrnxfD3AQ2qG9sR56TKbUjOnd1WGRgqb1OuASrZYTkst+eohc+rnGfRCYI
pFmYtBiGVc8S9CYIbZr0t/4KkUIXODlCC9uXf4MCA5JGo+FxKPzDIcCD1okgjQIsdDkF4pRS/82p
KbcWiQ/m8XRAokgrzxnasnnlb3jfZhnkJpO7OgpUal8XFn1GVnaZrQCVlI24vPgx2YNlP344tK09
rL4Gs4iLooezjM7bBek52W6Z8b7p1m/6CPkePO95sg46C8zD/i1eUoT2mUgglVwCVk3nWp1y9+WL
7WVNkK+5/UsE3j+XFNk7YfPVwxrHyjZVGDl0y4RZFr7yXnGqtWHLYQ3wzYez8K06rOQEbYGS4WZm
ByNCxf5M/U382vFV4pNOB723Z6gNTtfYtGKzpNBJXby8X/JQMOnIyFkplGN+HxnRnrtzwmy1cKKe
wIJ3HsmiTvolAx48KCGPUYlnRALX8NK4BKH/WdEXKvArPK2okHJHYg0XiFzjIK2JGDQ75/jgt4UW
AiOT5BAWDTHzrGU3kscxQJqRnR6sBLFOFj89bJWfox15dZBE5Ipl7qn40HpIj0EjbClAO0qvfAUg
T9tcNo9aKc4IQkvotNMaGYq6K9KanKQ0dnSJFeUP68aNiWSog8MUJA8/2XuA9GZTG1a9NGMG663T
RVYGgQoug+gigwwjC8fALTjHrrBlNVOM5NCwgbRbc7wIwGmeGdAXqj7wku1lf13PLn39CYraPHkT
ER+/Tdh2b8/KLGkFPDfqM3ZWBTK839G8m7uPMIytnUAzpOpy1Ltz8+oj1XMvybrMB58YmfVG69ry
9sOgT3t51O0VZ6vy7adGq10U258ElX2fXf1rjrqXloGOxz1ZLmGAkgWr+qWb6gf8rHHjreF/iQXL
Suwfx8yjsF5YuaMkL0zJ9dKcV4F3ZL3c5EBs8LjTHCupYAIzKNOVeIUI4Yu4HfQZj8RyutKTH3an
nbs3V1o/KSZRR/3lFV7hoo81nJTWc+RwrT7sKk7rMGOSjLoK/r1vMIn0YAnw6lDrtKtIjDcPqJNW
vciOBKgzN+RRrigbYAgI3o/OFu6fqWQX/7kbEu/nUE1fwbENPP5Sy9GBWml0qejKXydSe3SPEqEJ
AP0pJq1QHEpJFQjDuVNbz7bSHOBDkzx5NYtZh/5JUheiUMnRLmqic5ybLRCstAYR6ZSAJ79eUqr4
qs+ggBw1puiF6a01sdfplOxD/1kGwcXSdcOWNuIyKWQac7Kynvt9KZX+OiZztaM1TmjG+F/cN8jz
U4vlolLTgu4WE3YHklsuQVN7tBAxMBBOdkGjc+uJQA/EzdKJuMBp/VcKpL7JuIalGC9tDkO1r3/j
5tWeFlYE60SsztBgMj+3jugc04EbA2dLj46IlK/8qSu97mE1AJ8UvgJQmicnCmn62ZtY9K2O2D9J
D7y3eUybNgegJFyHJu0x4tRx/TsKmjCzYoFUJVDMwmjn9tqyxqvfpBd+w86m68YCNpljaGt428Mm
xjs/3ztnTvpTJ9vX/sZ1/aNtncFZQyPwkdPAzkndFDok4fZu6OW1Uv1jVxJWAFpOuQGeh/aG3YY1
YabVCX+sbO0WhqeWm3XIrAOkfd2bKjiXbZLfB2vEAjncyP5VaTWP+ktwCLEXrs01KlnrKTFr5GbH
9fKfhc+Yu1T+4xVY7zotehYQ1aicXoMTeoZu9EstBWS/HMxWOORu69yX4Cqswy9lZgjhl4Ni5/K7
kgzwAH7uf9EQU5gLljgSPuIXleXoY4gk46xvoEOhjoWH7RBsrKbr9JtzgvSzSXAenZrhxwheMhV+
iUt5ELjtWGOE+69Z9Dm4SRI8cPfIebafpJsXgfhoSeuk04sImErmaMlahyDmgAp+A2crczZR2p7o
8/Qit/yVBfrLQ+QPjWA0bH3C0K67yQCKzUIP+EoKLBZhwvE2psu3fssqRR+QQnf7dQB2QRwmu24B
wg1crF/AhSvie2Ku+Qqjh9zdORF1l+EUUP/KDpTbW3q/bTVO99vKZKZjzeMmZ/v9rDRC2iEz9RAW
O6hVSmjNw2KfUsLK8VvFRI0MVYQrFK57EO8X5XXpgauGbx2dQoSmGzsX+qa8VvXiJUhVGwz57yzK
Omx57Ckki4ByzvTIv/6KEtnnXw0XaXCbfYRk8oTIViGeLtWVoLtFo9nMdS1q8yq6/7Fm0sBwKTCM
Va6owdxSP6VDHRiru4yDl/pTGbV2n7AM0G7WFiYEcgM9vGKMWs/qeZ4lX77W4iBgmaleVY1HYqJP
lPcyMas37F5YXZ/F9zPTrhtrerRji/WAYYiVsrxYt/OWHG11IDzEuSIvOwKpaRsvVtXievaSBfU5
1E4X9C1dsfdnqJYTIcjF8kbKXUTaQx+KJ0TslEMONlsiqkTh++M9taBDEniLjLs/rf2TAXOzfJBL
uazYoOr3RMAEHpcygA28PUH+Nkhe/anYXGDp72FbbjmJL2wK+pGtsIKAHcUQQsIi58ZU0MUgMZtp
odsZ/5tSM3WXID8vfj0bBEp4S77Qw5Q5YqWymwJ3RKeu7smpGBackH6C3BSQLz91cNwbZXpF4/C1
x5ZqvBDdTi96QtOCWFB4feJadRJt/3HzU6PwNznA1aVziqVyrMxbP1lSyQ7e4pAQShi7TeKvIy5H
lRRQ6l32CkSSQFEBKcu4XKNBoGbF74Lxbz94h1bloVz4gUnhqVhYUE9Mg+kyzzAcmRldmmqeeudG
DgNa+DtiqdNKDn4kLlolvw0yqNs6Fz/ybq2uZAiwIjGitZTE4OSWE004T2iBWHDhxPrZap7QvKjt
Ceo9BKRztd1YbDJgTxP+z7WVWaBZdhajff8Fqjuf9NlJwoc6glgUiGXFqS9ESdQr148vo5snjX4Y
RMMvVREO0dckmoVuIc2D40d+UKmwz6QbmkhHvK099XMrsNcZZM2q3/RHV3f4j6CKTS08o4LrZ15E
WDM7kaPUlHlerhmPBu82YMxGXLGufs2V8JCODTEVD/gggj+W7qOwHhpr6adERIZWZ1VUe8Svq0oU
u0RFQn2UeP3uY0shKx2wzXqlqmsFPOhNNLhe18Jp68uNSbsso6SH0N31exEmbqPWEMUKnAwDRRFt
t94zppodzX+bOJ36Yn5H8WkzZEgCVe52+9edJJWswuSQ44xp6UaC0pYBFznVAS+7IM5K57Ng7W5i
nE6l26+x08BCJDlaoYZYrzattVxH8naeANdhm5eqnTtdbxU+bp5bFv4Q57mpgWcmQXoD/ZYkDySn
B4+MKeoytemPptfRWnD+Sm8K4zdrGEs8hlkU3jL6hixcckoiYIA9YpO251tZsg/WyA8CILFz37J4
LD8ojelM2IXE4Ga792/ynTmLMaSFIhB2oRH0icMhulGRDjfrGWpTZywiHQRGOgORSP+YivH4nsOG
zefa0YCWZHiHJJpU78zY5UNNcnO1JyCngJ5cSGnAU/nggc+DfSBRs1S3w0S3KwuIGUsndNhHglvQ
xWFTLVEQCtMDWQXx8NBtHqjcZY9d739n6LVj8MqBbGSdwU8sYa+mkczYP6XWAMZL3y3KZdst0/XP
ep25+NNCUHUIQ8Zj+Tc0rbYq8lbICMUFSzPKwDqRx6IwKYfzSgmV1krXTGO2KBGTPDxVGarHwnaX
s7s0OeKc/A23pjTebm72PoVJlQB+JfvrEw8VNSKX/fA6aKub1qb5FVi8C/VyNmHphIyM9pzI8Rjo
08dd2yBvRjg66qvl33YoIYC7iukEOvzgow//9dOrHHJUN1CU8I7bAd20hduvz00m1toGVQxj9bH9
Ic3iNdxOpRHpNKf+FKUs2IYafk5U3AWAYxQ+EJrQR6rUYgRvA9rX7igeOVu592LosT3qTOw6BF43
oBL1rEcwJzgxT4xxHS1s/6l1ZFgmpiOZjW58UX8m3sPFkrQWSeNv3evE5g+Up0naEMYnv9EYat2H
CQEcF9tECM4pKyNDyvRon2tFeiek8Zgopidalp1mGgqwMlZTKP2GLu0VkfBN30D44+1DL4bTPflU
+rKb1pFnUpkvwVhZ2RVKEUi1/SVOWsjSvXKpbsoHbcKESA5sW3cA1FIN2a1HDcIpysChcPpUIGEZ
1Hgp0WFSN/v4uebc48fYR7+DEjrHE0F+OZofBGwZoQvtjn0vbtBNkqfsDd08okzzmBaBk6L0cXJK
mO/JxzSK2SvzpWJcHSzIBgy9SyRcBa46qjwIlAB+GbD0F7WMZotnAEQoi/wwsGKnfCdBlXqqPCyJ
nD66ob+7WvHp6F42esvr56TMOGMl4jey4KfyntSTHoIVK2ChGAkFj1daHFLl8497NSS6W0t9URQI
JyAnHjxxJyNl9x92sYhTzPCtu8h3aS75jM5b1h2/JaLd9tznnXpCLOPZ/XD0Z8pDOG0z5hSgVce3
Zx7QazQ2Uz5qmiFSfKMu7LDGIbgCHyE3/l6TezESEVNaYgzvZICsRnax0ub0XVR8USXco7JaK7Gh
EuQLRm0Y4Ma9vCFtb+D29uAQMLbSaD2pd7FKQgIp8UgLvwTW7oHr7BOIlqaCNNykW8LFabUnJ2f5
jWybi8L3md5rwiab2IAEzyBJG5ir6ED+HWVPgGxYx9MknBPwQiqMyiNSgvvlwxml39suIffZAtHq
Axfylufxh4VpNiuYnLR9XMXZOkHsUNQbz7jlyYgsf4JVh/hVnaUG++6+EMvqx+NHq1ykLPgOofRR
QsBSPuiXiCThTZFPlTn5yCYk5a/qbNd29nOXcMD6wl3X3n2CS1FyL/1KIS8wg1CoLyQV+AD3BNUJ
97KweUo0VkX1gMqNo5GQalf9EFIc1Get/bfLqpaM5d8MYvWvQZd850dDhq8zZA4zF66L9xnMHYe8
UM4+uJHjugjRW3xrrksNi8ExsKy+0au0S3olJPfCJZonC16WWxzzh4VdcJ71ZE7X5xdf8AJqrP1w
XYS6sKHlAizThmsqQ1W09n7xj2yKnH20Fe5XkRVk+P2wT1DzBck+w6fuYKcC1/O5eFnuMuCJJEUk
VbJttyC31bcoNEhoC6gRF6W/HFQR8FdfTFHtrjPxdLHFDNTqDyga/biPftyy98SKK91p1tPZ0Dyu
RIrnBcDYDj1hwPUT6PD2z/GrSd2lvyt07FZCIAGXZaFbArOoA44KjJjMOeAFDzaD1KeB6vy0oneU
FZHtDxXbYQzeSOjN47PNYQEviOH7e7oyRxJ5SdUeeWxUUJiXlfymdKIzflmnln8szZC/AU9lbiLK
gtdIUoSTAzNpczueNzytNrFCpfpKWncEIV3DrX37EwhXV5lT1xo/JeK/wYhglqPCZx1aHbJNmdWP
6o12Xr/WBOaW3NfVbf3H+dmKVvf8yM2gkfuS+548JNNQalV9HikwW14mU3xm12/zftOUxRrDSAZ1
m5V0CUz8Y1kxgmsQjWWRJHKnL2RxKR3/Gaux3+41sawJzcoI4YLgPRqtdYTs9oTMkRZF7+GvzbhE
PEZHC+48Kn1PN2FVJkExg82LoKRD6jFAH26LWkfiak4Ul1j2bXL11p3TtydDj/e+A+MqPAKZuDKE
2l4b0oDQr8L0BDN3iVcrFFWzmR1pFeUxZiCAKdjK2gsKPm1CzYUpK5yXtxBhlAoEkunYIzbViqTs
+/K2X9osaRln9fBFMWtRGWHyudF5FwWJBVMDnxkNsyppI8Qn/YIguoFVXkHW+AmXZnnBqe4kRLHb
9MTgsyApAX3mVaDUFqlJcZ8yGUKeibI1D5pd6cbyd9Hb0mclDRKcQ/4NTM8VSPB4i/FeVWM2+h1i
QjkxZEPvrTjbGQoBSP9NwYkGKw4Q4B13A4zNd8dWgC4BhoY8thqQwUFhumzOJAa7GBVbBd4QE1Xu
hn53ckktvP6REw2EVNexrpgDreJ8VCa0ieH+66KdzmzMYVjz3A3/vFrEq7TPwUAG37di1gNA3+iV
B/Hs5kkL1QKmqqZuOcc5vjL2A4qIAPkOKVnuAyyTSfKrMs7SkXd02PbMK93m6nJp4zbAVouNaPtH
KNnywmf5TP5Xo20I1LROLanNiR4FuRZinl45fDCxqIh/FXqT6kIxF/i1SuFM/BQQDxFB3UvEbMsT
crt7HPAJ4O8jUnf2DcsMCMaG7ZccDjRyQbMWBWLF+iCxItjy+5gLgzK0VDIBZxHVwajV5a0HRbIE
nagdXXZ0CXF0YDsIB+XE7wgljNVbG3EgdcFHg3Hx3uCbq9oB92sQfXHknTM+xb1troiQKfdX9vwu
1eZuL5eFpvF+LXPNs6e+9LhVrkXHUK2NdYo3O7pu3BlypOC9tEIyE7xTjYVg2Oo=
`pragma protect end_protected

// 
