/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2020_08", key_method = "rsa", key_block
Fgcvq9yodAEyu7zsWWZ7LwHLqer2uRdIROgj+b6me/wmyj6mu+r4+a1EPBMoGlf2Rxb0wqrGm/yl
7FT0a+0gf6RIUa901Ug60cEq5l3MsNjnNX0EuQ9QHnbWnPHO5sk3W38XYr3s1DoIymcMyzWSb3j7
DAgt+R0iGXGbLJHe2UuAgwrybNhjpWacbybFOYZoLu5Z50wmOHt3p6J+gVbTwfuHK/f+KnS4VtSD
EJxx9+hQNEvkukNe5IcvkATvsJ495o97/SdF6+o/UvTHUZ0m3la3MPtrbbqjxbRc5d/SBaUYwJ/0
DSKgI3IBXs0nO4MGwCQX4Cy0xa1KtNy17Uqy4A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="YyF30NSJW4xBU1bz6CmJ7uDDg1utz4oEiyNQAWYk7H4="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
3JkMrY1IEAXvStruy6C+3l0LKp53P26nc+uVJZ54z7Bbp4jWC/AZdd4ZbHsRt3FM29J/oDoZAF/s
cY8FBPMKSdv0dEVtgLy/N0sMzMy7Kz54fPC1/1Nr/wMBV86M9x94Ezbl2XdvAOhtjr/naHuqS7fu
bgfRDs1xKjwbVyFMidGggFiHdpIo9nO9FmnFmKO0tqB1vVrRJ57rzJUKBd/uxPlTMRx8yrS7XlNX
oHbBAoHfo8IVRnmRHb4jrtG/jxI5d5OBqRFngup631xQLQRhaCb4pGo+SLmiiMeQaNGvllBFBc7X
kzOQjk0FZc1UTKsvBec6CqSjxIZ7kEPywAEdFQW4222T2lyTSx3Gb6j1hhe7Us7xY4lxtph4KbNQ
bNm6+LtNrbKBOCBfqIX/Vr+NoS+jcaeV8HvQv+XeOQz9uxKgOpLtagWnII9t2Wmiv8xuvj4Wff65
AkccVvW8FcUtB7W66XWplphN0Qtq7pOSn+CgdGQqS53mTHr1QSycMVysP+i5FdbDR4jD4D04G0I0
PidkvYlAY7n3XhznEvqC/PrKsJwU/rxf9jfvLvVsSK4YjANW5CmrJKmoDHvydrTr233/eW+5hROc
5kXnFc7nYSyayfJf5oksqPOUAolRnR1dv/CGqwY8dMPQVo0tfhHmPfjpTDkzrVnjw7hU+SwlM6Bp
3i79tuKiN9i7AxVQzHBL8X3BjmmWHEyN/gR9ydotCD8JkhtkV/jbvSdywDVXSUjSLe9GYi1n/Rgl
7Ew2zdBoZeisAXliDNi4oDC4VXqlXaxGqs7Ctob54UpnCGxYXu5xrAHOWJxWMSeqmo6rQ9S7dwFp
AZBFBPSqknWNYLiFTBehx+xKBgASzp6lFgZ6K9zD/zR30mR8utYebtzDSgQA6pnzsQg2g35HmnUf
6bQ/MwangL+0gogcBbI45l78dUi2SBeQ1LZVUN2oNCfRCJ4zPs1saG1FboaVMK/KOS4B9Fvqv0Rw
UVUOmVcuRPUSL72boruTyjPG8QRwn6dPe+RoU/Wa9z58lYjsVP26Hr+1Z9+zCWWt5rcLjHyfMMwV
gyg27YFd7SZ4ZCg39R2EaKqxg11bP7wuSAD6F16ILewFpjim6I+CAt36CqN/sJa84cFoUtmKkz11
MxQXsqz030KkwM1yVyDV0F67uqL/UBVGG8e5Zo7NExDdBekgb6JgnJxm1KsiNrXxBmyswUF0mxOx
W50riM/SXYz2gXPFD5Nd8tph2wynCpqWgHXO4JZT7RQZ8rd9hhtTEtKwd6081Gvq13QzF72ZNofd
DezQPOH+Srw+g3BT5yt9doiDA4Y/FcLxiDrGgMDZ4SRMFXf4y5KC9EXgV4ZDLnORtlVJG/u67KVZ
0myJmPl0jGPxB1QKCZjYbUQGSdd02KXwcTmRMcMRqDJvJNRNKmhJFhwQ5HVAZGnTlRhg17YNUEn4
UigyIT0=
`pragma protect end_protected

// 
