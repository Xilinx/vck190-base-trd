/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_01", key_method = "rsa", key_block
WnUYD0g6/qDSYmWHmuZSsLHluSdi9+myTeKuKMxZY1YiclF8fPuiqftouQOib18cBMrk+rhxXYqY
YxxEMkXifSggXUrW22+E+kt/etsSl4zJseXz6n9xUwZYg3xlqNjifu0w0ji98CtnXurauen1JNyx
O3YJAh7IDwn6xZR3LTGYOPxMj1rA3ndIEld9FoiPlSfzRSRuhh7ozr80Ea1y9ZyRdn6UvlSGNFWa
K+qWQ9v0fQI5P76f/h7qmdvfXu9BKunBkypsT5BoGjV+yipSZpdDPJFuKi8ZALQ4AfQwwQQ4W9Ow
ic2MhxBJty6sWw08okzuCC7DdaVW8+sh3E0SQA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="GeeiI2S+0qmTuse/FWjb6tqEZItAqGIcIYeurwykgk8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1568)
`pragma protect data_block
1KvCHb5eogwPJFXkT9BIC3oPbz0yKVwognbENYETRekunzsRf6d5hLu/BcbHcMzgDf4l/Pi93Ods
teCT5zGHsNVNJZhXLCzSQ4mqQf4VYLK78+Hu4bFkwrCKLWr/MxD/IeVyFSRR4qPV15izfM2iYMGh
Fo5aIEjaY81T0/aZCWKc1FytSihsXLzATQXuPzI35bL0kZc/Xr6zmw7aRHoGDJm9h782UfnQBk6L
a79Y+6+IAycsY0ma0aVKe0tRgEy1TqPqVUy1e8lsOULHCsZAlv8m04+GafQA1lDwsiScsyd2xegY
OuC2r3t3Lhp/nRnB0D37ulzTDDIawn8nbIqD2nJfa+cNEV7FQ73/oIMugvzZrnCKk/51CGksU6g2
gR428spXsPx9EYnQhSEx1z5rpdnuL1tHBoZg6dOhv/sLAwZKiF1humLYj1VA6N1K1FxL23lNLfgU
apQ962xb3vwfyFZTTBsZTAIXgD5LrqMgDsYbG7JggIp50eoZLcZQCKeJGPQw4irSCCXz5XT3lvo3
lExJbFlZdRonwZFf1N64yXnXaM4fdTs9UNMw0gDkVda+Ozjr5AbDYFFNpnN6c5CrqlkIP7Jy4Mnj
boVZxcgJVoSr6WE3fLnKnQ9OMSHmMSD6TXkw+r0bej2EvSTbju5g61kJXgoqd+eENfd9I4JIJX1+
EqMuRn/vQLIkIHQlse9I3nmT0H1/zqY8/1xq3Q2AE504CT2FIyMk0PVRdsDoOgkhHoLMDYMIApFi
MSwFxjHnO5xqloyzzI1JbDF2vHJs4t3b/MUoxVTGkBBmLD58ih5cfG/WfCSehVsjKKgbmZWyK7pH
53evP9DmaF+1gc0Ix+9IvQK8iiJ173DXYTclVRae1/Rg6yfCtlIzMeRgkmd6WlJPd+dXmUt+nBpZ
HlaB3uxQoOUiLQTB/ppSD1+TJuDlpbJQ+eiD9LisLr+W4BT6UFU6vLUJLAxW0ePpYGoroiPZkhL2
wBW7AHy59A2UMGpJ+44ApCQS+UVggW/kAk7T/sQnVgl8Foqz8zlCU2nfgE/MqDoFTXm8aLJ++Lvg
IUzrK9Lq/J43iqeeNATXA5fDy1kRMHPH1M8o0Jxc9XEdMlxYveWHIesLikpAkcqLFQfXiBYGXY8s
Hy3Def88fhNSUX66SrkSCLwUpZdGp3Mlz/sxyMV8YSJUwqm209iLY+CyMVUQWdgVWVYULHgXg1Do
M7x/wHWOqfpsbbRx0nedd4yCSAyM4LiztkNaf9ialouH5qNbp5DD+VBB+lTEUx69R6DRcbOpgGeR
K3JWOpxISqZoU+sSB4coUEFelsVzwQfJm9nrEU7Q9ruCA2CjutZv4FqCOFsk8TfJcMIs6vODVV1+
5JyuJZiIIKrIEJrgpHSg12keNGEOVTkM+ZahmksvDexbJKcPLypfDrP4FYC5DTY7LWLTfVRgmJ+j
mFzsv2X8B71Jal40fHsPXMcLIr8WkdEm3v+0VwgRF9KsuG4ngCUgjzuOtIuEYM/FJxg4j+OsMutF
/ozOrCqir4J0iEM5j6PHmj0VSajRHpDEdkjt1ThQMJVCXWCQ0mRigLR2sdpUwbPItN6kSV3SodIa
YfgyHzRAB8zzFa23h0JquE6F980CY9dQlt3ow9IvghkXRYCXMl8CfoqDIS5EILHOl9+PdR8STjXk
nB1XVtNGSeHmuo003UpjOvMtv6hgJ8yCfStWt3XXpEkI+QhoAP/w7InsNlMMi+oygzewFezqfK+u
fdwMAksvO2qjbmpu0i4qf95PyXidQMxds0CIMD8rEWEISAAlIhVfkxJTcQpWccMERG6pxgQjXWWt
S13uCwoURuuahs9DhcD8FzUieG2NWxr9vusmDgOUbsOSyvO7biXXWgNGqaM7LrjIxsa50BJixTp2
LCZNeFBh6ZgPDnJqgtQbJ9rIaYrjXKTAHnhyJK+wwSCPbHskDk3bdfoh9djK8uK9M2wXYL36jRRl
j1vJxsipm+4ti9a8I00Gy+9QS8pu/PmRb6mbC3WX8GrdMp2hyae8hJlZVothkfNjHsna+bD8VEAw
80KCbSxo2yBBqkX0HMZYJRbUF1xc+Zi7zvzA1Nc=
`pragma protect end_protected

// 
