/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
l4gSYexUXlM7ifAaBP6t2MLRFhQaRe7Sma+zo2L28DiA8DDFN158h0/DaBr1OsRaQKqTpiBWurc1
Kc+8TD5uaOBbdGAOqQnBtAA+GhRIwIir9IbLuxBMnT/JmOaK4MUYPqvoRzrgYyXFE5yrJmMkU220
b8Arh6+dyt3Bh0bC5r9kA89v3D+ja9uQnY/8oodAq0Q20j5GmOBNL7A1mEvLof/A0UYhDRCv3pRO
FKF8KrYOR3RN8PBeGCM1EFnr+wW3J99nOfKe+v5+if1arByO/0BxWK1JYTBdcxntFYOrk/8juzWe
cyuQA25yLLNZSsEfw7pTdA4YqggvIwnYX+4CfA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="nooMg7GjkDsMTPG3DLODBuXednbZgjpzUjgowzton6E="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
OIw4y6hn7TeoR9JbrM9EZIsyONjVLlt8+ePl3cP6zXTjMftH6yGwKtlW4QGPAJbEefzTBS8T7hkk
sujASFY/ObXoIsBgBNQdTRXxuQWXxnAu3vjLPj1s6lib80BnxLb3+EO7el136o6xp087kK/sKiEW
BLC+pSYpYCUnt9V+PL6Jv2XfzhgJmPLkOVtpAL6r7XYCdiefvCGZKlG9NB6spzO0YH67LObIJzbk
kHKUl6JTqQI/il+RYr7yZJloq529zg1jveJx81FXdcFW+GiY3jlWTv4WTxjcsPc/4IF1SffMD83X
INff38vz0xV46egdqMjt7hP+zbfZplMjFTR2ywW/sT/QCt9AOguQUp6PjAefMVZC2jaJUB87VDN6
7+Zk9dHyDO4Tf/Ys7zErttmP+c7kOA1E0eUgdq8kAHWWe5RyDTnyC95LkjTqiOZv6bqzoIYwmEeU
sP3zfkf5s6OvovIIiwSk0a59LiHDYZSahqTqoFfBm/VnaCTqjlwEhB7ukFCl6BS0UwcYF9DPoVHg
WdQ01q5qIqUHSw7PGsTZHSkjIuabK42NsLE6BpZ1RPLs2hy57HE9/khcEMAQ4Z3Dp78XVipSvTKM
2zDWWFERzlf7FcIK7IolrdRMDU300xEJviG/wg+02AvSnzFLmsR6TOjpL2gG/QLvMg710JWg0y3S
n4LFXYNZPQYNM4XASjdorsWk6InMduK1vFR/7SEeZpb9rGt0PPwUX/m7iJZQdeYFCES10iH+XSxG
vm6fZfwrI9BHjO6LLOxbCH2Rx/5sWYU6xiCjYwfcIPTDHhw2aZDJoVQ27wPcnDs6wnXhzeeqebDY
trXSk93ESMh/poB3lfRrMl4Jh0SVjc8W7z0eLO4HumUzreGQY5Kmb/8KDc042Ee+F8M9uuxFSuqF
XgvKCxs941l9CloN3v91zxfPc/1n2hx1zWzgCRhn+UVLEmKKbg8ifoT+h2D3PZQvSJA+p68GYitc
Vn/9PVriN2MdL4Kj40QBvN/Yw1MXRjqGb8fd52jPzyIQwuq9v34z40R0Dxc+nym/T/EbKKnp6+gt
VPL5oUNDTkpwUuSEISZ0CI6ZFsFJyV0IyLSbyaaxkL4W9ymVuzdmNo+DXP5FsUUVACvC/3j1YiQP
rEmPhXL+SjHCjX+MUNrJ0LjDg94khQOqXZMJxrKHD7xaW8+DTXyK/qUI4O0Q7RRZLj+q94+/KfcA
IyObdIuWkD1dJB3bQ/LupooSScFimjSjPf48jwR3kDO29mpH1xEvuROArrZx30LZbhovms78FMGn
yamixCT010WSFdqKXxwW2crKyysLZyD2rSMpEmQAiLWEXETbYRqTwxgzStdmG8fvOn9oFburimz3
+GV5ek+4hjEmw7kzcQEGt3rhAoFcgHzroiDxCdXNecSOrxQFNJKzIK7ru9GX81AuplQfk/NFpRer
FVB3fA4=
`pragma protect end_protected

// 
